`ifdef encrypted_0in
`protected_0in
ze74c34e226135848fe16db9ffd31815111b6d7fb642c521a3f628cf6da949865580b22efd062a7
ze90adae0e65e66a2c36a587d0a790699161455169ed55a01f2084f11770a774ec4c588039b380f
z6de9c5084882a40b79a175f5c2114b2b6d78b070cb806e1c0aa9258297f4687ab308bc470f0040
zb0b1de382961eeeaf2e279e1462520fc31c119af8f2b214846f56c2b3cd2eadbe4099496abff18
z15cec83ec4a77b868344aa20ba7360908f5c0de2a79abf8b3534b883bb12180f68b5d4beb444cf
z3fba8f13afb0abfe8fcc4294810f75afe452434d2d0f1166236c82f76edf1e12979f04bc35693e
z32ae028996dd85737a8f5adc1ebb94f39c940246e887647b64782cd7ab429b0544c173176cede7
z01dfb26b1f73408344a52b7e1f117f12bb9c8077b34876c2e6fdc085981637012dc9754765e1a9
zc512ce062e0b8fb16a214591f5c81e1353b900a611fe1f4886b57940b41b7f2ce99a7b84b04b90
z916f717e73bd10589c81e207ed77ec660a8cbed5b487fa50acde1b055c8870bd8676023f21ddcf
z9c98cc47cfa2d654ff1365d1f45035a045a66c5dfa8279050262529d2cac9e64fd27d9c7de62a7
z731bc808811ded9016570962244887f98fe5440167bd0088f2f049df882af501358497c3b28776
zcdc5426c7f52a851c35106bb93e16fff984784050fc808fad15da330f6f0607eda2d0e0e4b1215
z2ac5b11453f6b6c5c6b428261a64553d70b4ab9f1bc235c2ceff4f6e3b1ebe72fceb7af9adc96a
z694b4bad7241bfbe775016041d7caaa74d9c0e7b507ce89e8b01980415bfa35a8e346f54c548f9
zda8767c02ea87d27eb7a843f4cada7dc3b575fb5cede69da7a4701b2d725c73f1f7375e85a74e2
zdeae70c30f1127407402c955b283d7b9512dbb3cc85aff97f613d57a4efe57b3c092e5ccc5b6dc
zd01018bef01fcb6b6afd138be37349905063433d6fc88423f78d0a5cd8c325dc906237be6d3673
zb87d9fada90e2c892651aecfcd04caae277f299df76d77ce870132e5e40888bd3b3b1b6bc6e799
z48a23782b89d176bd848937c64ea2b6938c5a6c2c52409c3721f00cb676ae49dbce756d647186a
z2d5ecb2321a08bb462a97b513b2f2f7e1913c836666420a662f742f4dd090636a3381f28becec1
z1708d87f1f0a00e76b7fab8e82c4b58a7479b0d3618edbc64d306b42be8b9498e21a252a9f7760
z4ddccf620c22105b64d3442eeae29848475b6321275c60da85fcc15cdfce58c0be67611b4ad217
z85faa32f1a391d7896ecd2d6a476653f33c744e342ca0bee6222cd817d247928bb48ab87008585
zf4c934887ffb02320d1f5e9901371c546d07491c6dc0560188ddf7660969a0521bcf06899960a2
z846b97706440dae0671d4d93134b115147c7d3bfbfec814d2c532f2bc7b5a866f7796e878f79fb
z6352953b57e9db9e47653b1e11547331dc0137729d159986fd727762f733f71a51abb4c40cde6b
z54c31b914f8117d35cf603a8739650e082d3fe6dc459f61998511bf1667257aa026b391e725e9c
zd247c1cfe5888aca95b9556c330b436327d8491de44b02f0abdb98b49782f878e8a0f3dac87de7
z0421764d2c9d42e6c56f714d56263208da0024b12aedf6170708d3b68853daf64392e3521f60e5
ze510ed798898bfe2e11f9f4663b70fd002046c63fc74725a266d2037fb955af755dbefd5b79015
zc7ab97320e34c78cc1d3f9b1e7049012d911756a26b82677698f55446ee4219b4ab15bbea7c661
zdc44753f614ebf8a58498348ebaf6d9fd1ec3f349d486ef45e3869510be7020889a33e22fa0470
zff44430a4f4429bb4f1fab0266a2a3b205388d778f21ad297c1bba18aadbbe8d51a41ee954da2f
z731fd28b2e99030912b9fbfb4d40b09de43581c736c2db28ed89710a930ff9475004671d6ea3aa
zc5cc4344451998766aa2386f7bde52166f76138dc162752bbf5ca18b8742e0f14c18505e3ab307
z8d90b7703ad45811f311b6d51114e8517013b2cf35416caa76bd31d86039c625fc6af0f6084896
z66a6612d10b17be683d2e0d392577c58d3a25d0afac0dc96ba317bdc8c6df1e56cbd4ad109766b
z0d5f1ae923b8133240653ae9df1449a6765282f89488d266bd2b0de8b4992a52a51219bc4f594e
z6127cc46ce23cc31909b73782b09f974e71302a5ae31381f06b1cf7c0e02cfaefaea36e15edf75
z2abbbc2ebcb8685cefabcb4426ae4081edfb6ba92a6d6b468b56ee53c096529d723b51c36cce0d
zc3bd26dd1f23f7cfd481d98052caf353313a5a4b20823fa3c600dd01542cdac3930adfb25a9341
zbe92efcfc5dafdd33e4d852a3dba760e50cf9b9af9462581d6318a7154993aafa3064a2419014c
z4f515b54f9612e3af0f1b1d9bd9bd45cac7358c8c289cd66a850275c06516339ad2381ee707777
zc08536ba9f742c5c02f1ebdd2b46c5f0c77334da2661635b360b820ac187f6018ba02265ce714c
z74db81d6e5ad74fbfe1096dda36b47608ec186dc3e6d22face6825d99cc2b27545f1f05161aeb1
zd7ce2d55f933a2ff3064bb0327822f9dfa4a6d7cfa6f3195560ea3064fff6419892c70ae68e50f
zff14a6d7d9ac69075b145b90177720cd3d3dc28245c8e2c5b33631b2b795ac2906a9c5b10bc883
zd206731cfbc4515cc7a7670ea6e776cde73e90513be9c6c260407fa41f0a87e5b266ef47eeb268
ze80b6b1b03eb6f7e4f80361776d3c860cd0cd6243b8c1217ef916f0396dfc2495a6a0d873e2160
z0628ebb99035f7fcfd02c4aa0979df7d751f0efea8885d14f2494f9f2b33e47cb3e1ad720fd939
z90d620b4a73759198043d43a9357e793f5c7ffd7258599ccaccc3ad5e13923228cba804b96234a
zcf8d4c63cce68193d5ba1fb71d6203d22123ed3ec68435cd5b48d6e1b9647447cb0d8d75ecb40d
z97e3e5be7946bcdda2867f3a82e1a0d6403da978c6513d683a38786845652af50ec68bda974a8c
z1648016abb5c0024d1740a4b45cd3eda57350976423cb156e03c7cc3fdc7054505f32127e396f0
z0e0f8cf7b7bc8baca317a27941679269df3569616c7c32819a17c43c629183c1b9aa8ef92173d3
z57c7d921abd5a37282a3d47930f2c5e3e489b16bb6bbeb5aa9a86e97edd9bf84a5141cc261b4fd
zb8cb031d9ba0dc79f35da478b3b5b61fc5fc7b60a7012c25c282116b1d1aa8b0ba82110040468b
z1b66b6e41d805dd1fd98363f7706896fcdc8b5ce7d97c90002456fe3c94eb7878bee6d5768e686
z561ac6b573d1ca89b3781bb95b4bbc74bd1bf8a1d9020ee6fbc4d7b7d1ec2956ea5ec3d13ff2cb
zfe40a927d573bc8b44151839334627d318729d94672a0fc8127d0cd5e1828cb1e7ab2fa1f2a16f
z48dff6c183e61c338b41f00b75e149c02786ee76a2f1614f45955c5e1370c495e182be578352cf
ze3022bc9cc3909ad5f07942e33ca1db13d6899c43cceb5f3a6da7c52367231c5af141b1a6bc238
zb7b3173b4cec9a65a9cd97884de37612a766ed0d886761fa9e07fe4159f95decf6b3bef46a7ae0
zf7c43c402f55831f442ee51febd99c3595d0dd92135586fae3274df55271e78e69716d81dc1206
z356b4834246a866faafa8f2054fef1d8f31478d7edc9d270126699fa6b29158434c34f9d1aaaa2
zbd2ce910740c7699a0578a5ed1e80cb36b7d64731a8868d39cc8e5b72407b7d1b2abd38acdd129
z5924eebc6f4363590c8a0cf20ed19f58aa57d8ed12965df00bbcf09a5e9aeba3219203c0fc7e92
z35af42a359b0af660e676260611fe6248f0af2c9c0232e84456c52436d16a74f0a4fdf96bfd2b6
z37e97dad6bd9f69f11f692daf542c2c4c69c5b84fb5e9289b807d03cd21953d2d67736cff638f7
ze8c79bec09a4717e698d1408ff4f05fa0880cbc74c9a65f0ee6bc659392d8445cf039f4c05a090
zdd336df5f24fd747ca20d2013d7f5db7625f66c3a65b4943858a0beba5880bd4e2f4144d500c63
za675f3eb9a50bc8ec07cde1d189d6e9f1ceb1e3cf8c455f520a74a86401467ba4a41cb0458fee7
zfa24fb19c43b5f1c4dba71213dce338b8b6388e7317c5954d3df32b5df8e5d492a446d05575b99
z1e98e6489c1899a04c78158b462974cdffa0fb1e43333c1fe8da3d62696a0675c23db9300c0c3e
z8d908e1d23d35d679d11602e93edf8d1966e3a60931d1961108014980ae6f0785bedce2ca313f6
z3029093d95d7c3fbc88c34864354f88322cce254427e96a7a98a68de14be340af63f6e02385708
zaee76d201cd55e5678d0f5535ae9836bacacdcc25229f2bd3d185478680fd4ad1e89b0426ab88c
z58c0b2f75b885dcf9766958cee9335653384a5c36610a49598f499903d6c40bf640349034fb5e8
zb9080a61a089606ae93e074817a044f2b395c63f66f836578bc55a929c60c5dbeebd393c0f3253
zca0ab55bdd3ad38bfb1ab4bd50ec2ec4bd9595ff5e208edc003e6ebde014e09e710e8d92fd406c
zf42e86e3959cbe6dc2ca21d7bcd005d4a742439d6105491108eeb336b478ca2652d7f138982b4b
za27dce5db55a346349a5db78d2129d140b72067e615afbb09f9d8830e68350bf464b5eaf64db3e
zbd9ab2ae373b00175ab82d749554320dbba6079b8333f540ae728bc4c11899952587b4206e1608
z1116b9b8d7ce26719e7f040673e3dd8c9ab3ecfc4912dcc704855d707196f2ccac17f2a490e782
z6626c3c1c51136c67411bc0d663839a2cda451ada7c5dab922032260acaa8cfb4b8d6406adafdc
zdbf4c5e4c43ecc7576564e484cc6d361b651cdc7fffdbccae8e081cba91c6662fa063f63cce858
z5375ad5eb76f5f4219aa93e7805f834c74d77b423f0c1a39c765844f26db4acc48d1c56064944f
z57aa979b17495063b1e8b37d754c794ffc6b0f74dd680ba783fb06af1f994bb4990875d09bfc10
zc1ba17f1f3239d870762c94f7fdc3dd2d06ba85aff3ee1d2cf0770d6c67f6b6d7d741f6fcab550
z8c62f4086290dbe2e6e3eaff4d951cde7948f9624cb4183e7bf2c6c15f8cf2f5ad9eddf418f8b3
z1b6a4aa75e48f3df26bed10578c144fdad70f765ac71d5771a86703efe238bfda780e8c95a6b75
z07ad61887ee35057ece65ce0d4be1cbd99cf45b141534b921fada088ae693dbea6949ed1f4e9aa
z32935ff43020279f95cb6d2acdc672a95ac0c0d31242cb978cfc7a6e40ea33d3018642147519d7
z493c08f90b886439a6206f610e99fd0d6aa06f7fb2855b87c2f6e4845f102e46d07d41c7e9460c
z315fc32b0b88e433ad6492c6e9cf4c1fa3d300d4a3fff95d750419fdebbd7d3fcd6b0b834bb2cb
z45354b64f258f1ed0f7e4ad66cec34c7d23ec78055f4288c8a834b6f0d1a3ae46259ed78b56f68
zf2a07685d9e3f8d7b0e9e76983e0c2b32638087e95030b85145fd6bda9ec428833ad32d4fe8876
z54bcc37a623aeaec9e8c0a8b3f3877a74e366326dd66c99e506148d8ad923c593464b558068cc5
z30ca10f5429b2b7128056f9b5aef587ad06a12c820fc4782d05e8842d09fe782be05c79d52dffc
zb12cd0fb7ea2753f11a63a3304aca7a26433cae5bc8bfcc71f76bc43cb5bcb5cf4f9bef3cb1013
z88d294e8ba726a6b71380fb9e72d424f19dfaeb0233f53e69fb248df512ed5bb9ff6e15ce7f417
z042ebc24ac6abdb93e90ea0f8007204f5133c8558761b687aa4f6dfed0ac81c2b6ae32e575c185
z29fa745a94e6a9aeb82ba2db9ff644faad99c68bee3bde317670e8e8dbc8c02a715f2b509c0981
z7367278dfc33a86346128b6c8ac2cc5109b509e30a7a62c6d411b372c02da0f88e0f4cb8eed73e
z81111401a595741644c7ddae035f3652eb8026d9df478187b8c944dff6e1f733f5febc55e8ce45
z54a11d09b29b4616757f3939587babdbd0c6d897469e04b3ecc3d4f30f42d4be776ee7441fe286
zae431381e4ec6ebf8b9c682e4511ef3ae9a65e2e1fac347b33546b94749abd98782eab4fa59973
z475a3203e55b94e3aa619ef566f226b2331aecdf57f804f7f85f897ae33abb9118b2f16cedd28b
z2419a06fcbc5a4a46e38f30e15c37c88bfd0ea59f6021ddeaa9bcf3bee82272903af0ec1b8db59
ze37f8fbc00e637eac7fc8f73140ede5fccfb8bd980df37cd30ccbbafd9416e99f259d25f76c53b
zec1044b386e34cb2ed4996092244ea97756dc0eac99fbbe54857d3135ee3344160ee8bf57a43ef
z1b72a7950aebce0a727a3fdda0c353fc2e9440e67c0cb8384ba42cff8f7a46859492106ea9595d
zbc5fc882e488d0eccb977a95b7ffe494f3a932d25182b406bef05ff979892a76b25c161d5b5a3c
z582b847c499ff754df264d774a3061d721c8189499cffdde84cc5fd14b5470b6c7208f76ea77e8
zc74a800be7ce5789d122e8c5ad9a0685bde53ba65f37548835bcaf85e2976d95db1230becc7af0
z8b5ddb1b2fb72d0dd779054d43ab324dc547ee5a51b5ccb3f5f57bcda36314ae62490a0cf36d9d
z071eead04285286bfe02cecaf53454c6a52317f7618f39d0dd259573624219b6d6cd50d1aa7906
z46e2828edbe56fa3901a62d69e66b7d00fed253c6a9cb0f1a08dc8cdbe7c84e70a1b2fa6c886b6
z7db1b8c9f8ad9f69b2b6c98e2140232d82687e1e888ddc2c28823851235161028ed0ab05d6dfa7
z39a9fdcc811b156101bd1f4764083682a7c1a0ffbd13e60cd40d6b3cece459b0b9dae6a3b7a94e
z6fbc02e5fa8707588a5a54e3716fbee6c8b400e1ef1d0beba22e7cc12ceab7c928f810163f07df
z7b0479d5977286afe1984471e19975ac3313e46b7e9524c4fb4a6049679755baf279e2aae01b82
zb822acb922245da793046b25af74dca7c94e29a83d9073e02cc31b17b568e2d1ffd8bee701439b
zd275190870c92b9323da4a66c596c6fee6e73c4b1a232e0808bbd93c6438ee1c836f9165500a67
z21497f5b7464f7df00fdfdf6894a09468cce93063b01731c2699e01cad3396a17ebdf882d73868
z1ba67e37ed95080bb01e8c50b8c27ca0faa3a6c28fd97af3e8727974017cf3635fb41859bfeb97
z00218a09e7551aaa73e421d984b11fd109f90fd60d8b8e2d4da89086ba72a743954eb586e0e24b
ze9f872630d51ddb7458c92d9a97a4280b06b9e5a10e7bc95947e20441e592f04f68e5863c89da5
z589be0e344bddcc5bd5bde5d654cf5ee8df964f85e72ea87f58df2c7daa79c7ffd80c798df2ab6
z6dd5be90c638de71495ab2d93631e08b272166a751b7b702e91501b1466fe7accab19af678a3fe
z50bdf2dec3f4ebbf9f8cbe74db89882ed092edfbec04b8df1c5efc277aaeb1d0192ed0a1c38232
zfd219ac79fbea7624da157ee39f321c00b3213dbc8e0bdbf6f3a2769a9d1059120a998ce678ea6
zab3fb0f415aa0a6385d4748214724f2007a550a5536dd4db13f9e44d338eba350bf7a09251dc5a
z2b3a3f8c5626f8384414bd03d91dc14487fda3a0149ea30561add38bbdbe95fa502b5079e38323
zbcfdc06897f5ae3aba3173bc91e53a7f99e466ab468d6b8e8256771b1ad706e6c2f499dd39b285
zd17ab04e1aec295c238f7f8bd540b06eabca0899583f66a322e77dfa4b66dcedbff98caced262f
z456bb2cd477bb3b0143c84ef9e8779879967cdee90be173569bc7cedc066dc200281430e0dca3e
z2477582351fa4b6864a68235663081d3a2adcdc274881ea79777595916572e0b20e2468400487b
zb3d3f7e9bd6bde1f67b027bd35a5d197390ead7ba048362a8754977403b023329443e2dcf9a079
z1578a08fa4052a55b773021f0fb88286b0c32143f0b0fb5827185b1aeb944e127862e7105b02c0
z64522b043f694d6bbf3310c41ccf46485c84fc726d372e6f49b1db7e917ab8890e42c2be4f047a
z24f9e05d1ac3cb1052d09f6484417afcde51a86bf87056f327f6e9025881e92868a0a31a2d861c
zf8f575e526400b342f88b1b38ea7636c6f72791f484be22b6471aba1c8922e5d7733b4603a35d9
z37618ab8030012dbbc83a2ba5cfc70ac57e7b5e75d1087ee7c601cf68103dfe59381f20c565406
z4f9435dcd5584928ea811dc7c4525458dda2ddd4fc5933e47fd64e0821fe2a75f2c1c303b65704
z146e8df08ab248265d7f3d378eced9b0be4ea0584702b072213c0614da4dde9f408b4ec4bd4266
zdc511bcca4240eebeccf25ba18cb8911d55b9857de01893b628188d3c3659957afa8ac25e847c8
z59ae71648b54af4c8c0f4d5a0c739ab5d363ffc49e7125e255b5b242dfad611242aa5b748f2cd0
z4fe3c277e9f85e627a2043dfaf6c2af8ebdf8bb3a25bdb10ca15bdb4caf0c666cf4c3aae8d1cbf
z58fdd2556b8465ca28c8bcb7896e5b204ba6025930603b83c9186e8456a6b2a97fc72ca5cd2890
z86f35549eca44a574e805db3f6c5130ccbf39679399ea9e1d4b9bd8e65b54832beee966aecc77c
z56b2d4cedcb4c79bf63f5d81e5d89ca0a508cd3c6edaa238b834eb6fdd9bc4b907c1de762f6149
z084af434711a462d9846d803e9daa2770fb8fb02f5c39461eb3071570c3a1f633d489931baa1e3
z07c960baae17c3cd166f728be05b72fa2817f00f049352b4c464913d80dc03a5bbda16c9a4ef59
ze8b5d5d54ba2c2873e5f8765984ed5a987164ca4da44bf5f13a1710a5824988a3bbcad237cb328
ze743e1785dd7424af8061f6dd0bdada0b39ea761719f98e8b53102a1d28283f615d8812ea65219
zf5a8204840288137f491575e6fe5c2bff5cb5bb0c47b3ac910e1c8b9fafea909254df723b50d59
zf760088cf2d41ae69dfa6c41f159ae16b9dadec5879fd04d944c0e1ece15e9046d1b054bad645c
z693ddeca63a59efe1d969d96d4b7c809375666f3e9ee775b97b329da1039565c8397ff8caf45fc
z20bcd9ef4e3baa96289cd7e344b18e6026f9b21b15992f3dd4f2420fa935eb7ac620e2b7d426d6
z4e82b2d2bf9e208dfe88812d2ca76bf014f046158035e779b2ff5a5ecbaea8f3931c6f26ff6aad
z3355a0bc0c3effa08cdad0e20859262b8383c2a439abec7e254ad22bfb08d108d15fb19fca37e5
z8b8e634783297f2a0cb9cd6cdfc5a7822e7430496e6c41f546877ff4c135553352acffe183fd24
zebc5e7bc98ffca2d0d56c319fb798ecfa22f9baf079745de7ba2b276499b470e98e7737095327c
z5e752376601dfe7db70e8fa867a1aea580ca9f3a7ec8c78ea0ed8047ebf67650c42577b35dc432
za191263b5e2e00ec5faefc3be472f3f13747a911626c7021a739bd82702e844be7932137c3477e
z041f8e7571e09f43c8734dbe4198c581f8b1f9d233e78209873a6bcae7379cadfa22483812c8e0
z46a0d1d89779de239e2646edf531a89a30379c7dafee3ed509a08ab6301dd5d5e5dc04083e82ff
z67a35529935515c94c5fdd80180d0064d3b0d642188ca337fa05e19abf9fa938a768bb949358e3
z7bd13767612bb4444d894a1455439b95f98efdd3881e886cb1f73c57d2a9cf8d86b46c14fe3a02
zd2c2942270a6dc56617b4f9f6c333b668b786528048e6695f7e7d1bc60035b0d6a54504c4e8e8b
zc6fc641841a00318a4eebed0f230b0697af76e31621b6825cffcaf8bfab7445355c3894b7d5e1a
z6da926bf1c3906ec3918323d08f06af7cdb530d5cc128c400c313064a5d9a40141d4fd5021aaf8
zc784ca5205a49055282a7f9c1ab00cc2484200b252390a36eb5c1e4e3f0923384af3ccbe80d7ed
z2f8ef43b6dcffb92873fdae6764cf38fb843826bd96ad6af391aaa387f889819116b5bed496653
ze73a86a9a908e9829a11421ed5b868441ab23594ff419eb3b21759d1b2db089f97504634acc9c2
z8e1abd9a0522b0456ee1e0ee31977d1b05ce64565e6aa9bab61883a71b77cd1aa947ec7754432c
z1e0bf4af9bef985421b93d1922aba1bd8dae5d41c5489c34bbbfa74b6c15579e0c416a514c8912
zd6a1373ad2d1a8152b584dd7d5fd53eba8d1751063e0137d461f6bd662642342d38aea4e6d0e4a
z93084e39400788995a46096f938b635aac6ebd012623c95a64de7dc29da3662d7694c77f24133d
z82219add46b2c0696b9ad297bfeece0592a73b3e7930a25ceacf49fe9762d4d96efcb2c9ebc854
zd1d850538ce41934fef380e681a526be5338c0e88ee591af451389e98b8ff5934d6e286b106fe0
z3ef3b03c3166d9686e4ab3939b1819468caf4b1310b1d3ecd5cbb5352227063cace4a33620b7af
z153b0ebe4929d0d9d4540ee826b807945c3ffc773b92aee53cf5d1c92fac8226467a15e6664a7e
zd8628b5a511ed8d99ea46c2b48893ba713b3e3711019624b93612d8b4cdd2d5095adb37d64b0a0
zb2f0018eae45db1eb46006ea28e3ab45ecd1937262d19cf8a7ed38675eae247d261876a3015d1d
z913932751caf2351d434e1756fb3987f4d54c1d4edb919dec0bb4f4cffa45abc64503a8470788f
z60584e62b9c430700c9cf6ae90671db36db1c2fea38c09922bec18b163ca80d2aebbd1f6aee076
zf816ef2ed5dbfd9e5b1a973cc5daedacf868d440f8362c2a22a952f6aec0215ce046011a20addf
zd539bab3b7dbe9a79dff5e2fbc61cbc596b2b1e862b442fb0e8154e6640877e2ba9eea57aff96f
z79affa7212d7b04b8fc87faaeaf3530cbc3d7a9e021fe755ba4badd545783d46ed0332c53edca9
z7b0ca77c96d832213a31c381535c13b733ad340f3fe96c67b83e4a9764a710d2563e5f547651dc
zdf4e53e754a2e4c1b65a21c810d729c1140fa21d22864ded03f4e23e01342a81f089b8002f124d
z9c3ef0437eb68979001982b9f10340d7a5545fae7942b53f074c85ffd4baec292c3ad0f254d540
z79e9ea724bbe7dcbb88379167b7a80734dcc62bf5e6d00f1c69691d42cf22b8cce0d57e19d491e
zc447e833b213d418ceb43abd7516edb4d6837bf29ff5ae1ba29ff60346b11870efb248ea680ccd
zf03309a2567b27e1e9f3ab85017675c83675259391092e70d28de784f0cac5ac9d0be4fa99d892
zc509fd902d011653132e14d53bae0a40ded0871944b1ce905403ac6b3674e096cc6eba15c85f07
z4a9bfd33e44b2f120164928b889ee5b23d18887fb4807b0679188a7c18932b5d0ebc7a19a85305
z926145b2d64270b13d9748b05bbfa5c795892827913a180086f5badd15ee4a2da3809936c0a6dc
z786886ac686d06a404732a1effcb7f18e6162af2cce0a8e657fe7a19106e14cc1c02b2e4ec9eec
z2d239ab894f9254ce28e8065b9ca8070daeca46dfe2d177ea57f854717fa2774373c1a1a741c6d
za17b21ba840783147978e186440cefa2828e928fbe482f43877850fcaf5c63f47a70d821527772
zad08b3c3ddcb5bd951af73026427e560678b1ef268bcbaf5645f9f85abe087dea77dc240e88c92
z7371425309e5b026ede9651764bb8ba538fd647fa73ed7ca83368dbb47c46846b26d329f101af3
zc6d042d183c2ef25133df273d5660d3416bfadef8664a2d1cb2141a3b19a50b37d5248d360fe82
z37ffa8763d3131c5de994cf3eddf5b600547345bd57e23da2598ed9b3d64eec45602d6c8278cc7
z72e3fd938baef9acf0e612ba02ad25069d014603e2cba6d6bd5d97e6351f81bf48c74b854560c0
ze9d6ca6c5a25e2b709c6c74727f8c7241bf0bb704111b2aa58aa5c06bae59adfe2e7afda572d0b
z78f41141ccf77f7aac2051197f5e9ae20f5a24a078d8fecaa0fe953eeaa9a2b9bc5b1f58d5cde8
za187e7095fe7a23424576b58d7ee1743e2c7f5f48595086aeaab9335d7d080d4bff921b40fba55
z5396e63f70ca040b97e9606784b80304e565e214b4a5b3744d219945d0e85a2edb77b1f19b4be4
z4eeeaa002f34033b35ab725ba48c6c34f4adeffa0051ed9bfe7c2a3c366f0784da2fd0fee2c037
z0fdf69e7e55eb7244efe9bbd6153b43e2452a9e10b12eda16456f90ae6223e5401d8966ca786be
zf9d5c30d07c78902601c9d4c90aca434544e3da42770f95e912fa712bb5e5044bbce5e0c7dc7b4
zc4144b5fee725e125bb21dddf7014a99af68921dd910d4bebbbf37cb8a0b36a6d312f1656bba21
z0359d60038e1c4f260785179dfc0a90337b82ac52970b4fac3630e315d07c9f7ce4d7d800565a4
z9165e133f1b9f7479bef86edd5edc0b33a6497fe0953c57430980fa48b1f47531c2251052cf943
z5a5aaf3be49e5a82bf7791523c51f2e974f3662d4411f18a2baf614a0907b3c7030f41f2940b7e
zf44dbca2bdfa2fee11431ff6ca5d7d4e9605e01de043e7dd29adadec2368185d14939b745faa92
z364969100b4b3fb9206524fc4e878bb43ab010a48036ed9dc5b84776fe7f23167a4a2827a27384
z528e4c9daf0754125191f1a7a56ce79d3467d34dde9bd004339962dae761adfa1d7c8cb35bd5dd
z5d4e7783ab8e177cd9116cf6cc2370eea7e29f54b8a2f57e40f5b13bfd4bc63dc34cf13d21a1fe
zb1da4bffafb0d1dcaa8a2878206aa85176f851b6c0df0e68ba381f31f28435756196c1646457b0
z83ef970a0176a69c13d6d856d02e851dd6d91393a68f5cb9ff50b15bdb65c510b0dadc0617acfe
zdb809fd381d6017db80475a7a444d7c2d265667503bacbeb1b713a55f370d81a26fafbe2830b0c
z51a08a476e256a2ea24178570a594c8b3c475c5400a6d351a13631cc96ef90c4758151159b0d67
z19827ead965658efa60404fcc07b549702f034d137d621eee33c881545c992e8c87903272b4d8f
z987a29f96f814008295650a4b3e674124d30e52c9c79037fca73ac93d9a3464c2ded82e0377acd
zb113e1bb8136f61f880f4193d1789316b7154e491465e49bebb321b2fd20de4d9555f3b3b50c30
ze7605e5f9df0db3aa4b9e78883b097371c2d6f6dea75a9e72ed503df87099e5e4fc00623c7dd25
zaee991f090bc33bb86ea374ea835417cce68135955312189cb99d5807cb1988d24b0ebf051c4ae
zf998a929396dbb880fec75a5879c220e568fefedec3e8b381d1531b9832bc59c2ab720145a807e
z683fc8660a63578ba502a060f16fb3ec214eeb84caf501f13210277b034bb492f1498d976462c0
z642db574ff18686738f6fc6c10d6c76e84676471b22d1910622d707ad7e8722febf0c63b3c5d76
z052d5a80fca257742c933fa99808c30e0e18b743b5a2f67e5f539e7ac1cee4bc4280606296ee82
z5264cbe53d37cf9f8131dbf0ab8f674c938921bc15c6882d3bb4d60f2671a468c28ab5be28645e
z0262c280c01f71218e570ca4a2953295b263cf367b16af0b161923900745f76844e2658a06c1fb
z381ab6def20505c6bdfc6e205bcbdeeb60cfdccde02f765011eee29eff8f28d65bcb3579c38f37
z455674858eb70b8c5f23372f20c15d7449ac26c41478bc76f5f4dd4eac911d41a0440a874aadc0
zf06b012fb0d863eeca652ba09b3f94f62da5a4462048be1c21acf49b0cb2a609ff60d7eabc9bea
z09daa257d578efcdd635d11c178594ee73cbabeea103aeefd6e59a01dc4e7e9f79f8e6d3d31386
z8cdb19d272be15ebd8a95be76976a02a245207cf13559124f66eca04b561ac784e74c324a6a2fd
zedc3ce963c04d34e8d38d521b35dec52a20b586802c806fdf2415d230d00b7e7e1022a4784cb85
z9fcb92b04e60c3ff509eb9790d27cf26d1cf77b131cace31e46c0c62164013f446a980c345192e
z6a460e87a0fee323d980ba02aa9159edb9adc59839e7610e0e47b5f0150e32545c3b23612fb534
za657d6234371ec489adb0f98b6e0f4616e799314cb71189f470d36d480bfd2b9811404ba3add1d
z02c5ba81d0ef8ae4722e8d9ce96411ddbacdeeb5da6f8ed7d4b9c619a84169b5edc50108b8c061
z8b01b580803d1a201146b2ba99895317393fa0b721dd8b413988bfacf57f6c7fa93b5b3b09063a
z9aaa244afa1662e538e459cf8e3378c108a615ad6085e56c1cef998a8db01c412d152c4a04dcd1
za182bcec66fd9166ced7263ac185b86a10759cf865996c7ca4236bef88e034353e13aaaf85440e
zef0a797c84c35dbb5f05573c5a8ca0a0173e3910f1b8c2c610e66a7e2325ce71a31b07376861d0
z578eb47ad2fd0cca5a824d4e2e50f1265e63d918b81101a05459f53f8ed64fc1fef48f719c9026
z352b01775d5556e3ac27385d4d2a1dc190c567f4e36e6c716512d9223c1802b38e276ae4461e41
z640db04aa4b1ec083979aabbc319c7512eabd20ddde00301163bc80a6e82bdad91d466f1486f99
z64c622be287c9ccdcfa170bb4dc38899996cae22b25128cd2a33bd44bf848d708a5914bd2dcaa1
z1d9d1f79dbcbc6ad08d8ec1bdd7a859f8ca0e9ca613f1627ac954fdbe7ceecd79463ba8b83b2ca
zec09d0415916348969d12ac17bb010eb6ab2a5704a73a9d4185004ca5061c2aff20169f6fd0356
zef54c1365425ba4d2426c4272d1d54ce4cb5adda3a95c87b30c380120b352dcd10224d25aabb1c
z99cd4d46923179b983405c04b71c8f49e6f010135848e7cb7f52a300ce17bf1d23d37fb317cb5e
za20940087aa48438943b4697028c729f99d00afd0a4541fba5baca397c635e0d52f5d009c8fb9a
z443470ccd083c27feece86e29435886c07d7305f77a0c915212fdebbe8340ed3de1bc03e2b5b9c
z2a7907eb2c43ee357aa504c6d97ba953a22340710120ac80850c719bc93859e6cfc71f90101bf6
z0bbcf3d937aa2bac0d0611c6691ac29fc7c4b6770a9457f2427a56f5e65c507770169e8ade2f23
zda89c2de9a97f070ace0aa72b80690a9904dd22fd6f2cabf0a1e9ee0c12771c81da8641fd89cf8
z3351daae2de3c4bbd3fc4407806025a6564d7e593fbd747ec012024f7ee6880ddc147d178bbef8
zd5a28313e89e6346d4063cd80d15e98447d4792ee39864fa938b8b34636fc559c24d1ead194c95
za4d34661ef57e5a8542daed5117973a4b9ff7416438b277f0e882d20b320ea7bacdd2404c10355
z0022201d669554be59fd80cbbe5795f7130627fca9f6e7739ab8d299a812ff117fdda4ad47e5d3
z8bfe4ccb77412dfd733cc2d0dcf56528207ceddf45daf05ffd2ec89cea3d15024a84413aa5c9d5
z32717d9fa29d3cc4579e54a5b65bbc3be397d4fed597647daa29b065c27f51be8ed4e42b8016a2
zfd3326dccd164d2a9cee999b7714daab01218268538902c671b18ce73d797f35940e937b283d90
z02fe36b9be8fe0575053330182c4c1b48a93a995850e4557c82c7dc036dd85c9679047a0ff8692
z6e1cee4b758de62fecdd486929229ad1060850bb832e75bc1e0876e53244ddf1d1d85473af4879
z62e8bf0412730b213ad89a621ad106894ce0d7cad7a0609f7e5dc0cdb102daa59aa388f9e05ab8
z450c6ddf3872cda25ff1e56d8612769f21ec96c1c3744fbad5860cba78a0fedcb664a8db59c77e
zfc4ed67462d3c1ea1f614bbf3acb7b66fa9b9c3d2c07d794e8907509f1d1e05bd02df5ddc3bdde
zdb261554f5737ef0282fdd31aee95f200a386e8f2772ff13b5ada74623ccde06724684b7c1512f
z2e99f6345cc530c26bf6edbe5b1e0df069c995396f36d4a4a13de44c4d83e7b3366484748a5767
zeec189f26ca08e1790553fa16f94e8771f4eb4cc322ff1dfea66c70b46bf03e6200eb8b5674527
zc38399ab13bc209ac527b5dd7fa7cb32a90e758c9cabfac6e0ae995a55a82260b46a3ac1eb0c88
z77e043f2b410984c16dc2c18c481c417a6a3cd6fe7891098a4fcffd641d71c1ff23e3adb53f122
zb0c86702bc9709f6c7dedd20ed8185d47a32ac1c6e5ca9e17eaa596f3beb99e302d7ee45e80df7
zac67d28c79f5e3b1b89d7070d3350215216e33344205a087a761e3d2786841151aa9dc987e11ff
z18e4c98777a23636d71503b3347e851df9b3cde852ded5e1ff237798b140724a7ff4f2a419a090
z4a5ebb33586751eca44bf76141e766cf2fb5107b3f99adedb6cda5aacdd9ccf35cbef676b6e1cb
z572dcdf7e3ed12b543752e2638fe92420b753ed6fd5a9bef0220f8f77d25461f5fd5b6afbbb674
zb9ae5bbd767fa4dfded70f0b483af6c4c284abaf1da41761d8d88c40caf789564d0f2be261a3fa
zb65dd9e4cdbde049d9e39868d9805f0773418ba681109aaf1119cbf4055994b3eb137fc24da663
zfbb9616bc902d6df05838c6897b963368c40b36f6353c244404fd735789af1cd32aabe846c1bcd
z4f31f5e6912180ad139a1038090069f142bdbc4c4f1a0280935b5387e4695bf588784b38934936
z3993f7149733cfad9248956ec0ab70d6ec103bd2e334d8eb5718af3730896a15af92856dbf8e6b
ze005d7b2f993876221e811cbc4f37bb72ce3cde4fa04ec0a6fd5b1dee300af48a47aefd4d7fdf7
z0fbfb79f554b409424be241557900a03ce2791fd391a11fb7933c3f77537baaeae951dd7c83fd4
z18d925fc56da7c2452f0e24d6e2d25676de186b758193028080def0b1316d08b018bd29b4f0ebe
za27f1c7f8c20d27286689f1c410b27a5a7dc419b123fa0d4f5cbf12e1e492b3636ee2eb41feab0
z0c934e9e8c7ca137612433d7c0d7dd23cbefa780a6fd37affe9236af879ebb58f36ea893e3dd5f
zc50b93753c1b8749bb9b5226db57809d91a3d4592bf4ff7469d34285c32e929bba998826f95ed7
z3807140010c8203a1849b9196e9fe5a9d6fea7cd4d9c3ced31021836131629e74c4b513dea521f
zde9cbc4e910539ad9a85a6255124024b8b737af068d9e3b6451d48526dec904f6a896d277fbb59
z5944c707859fb29530932805f7972cc7810648fb58bcb2c8eae5a8950ef78554d47fb22139a50b
z680441f2280adf287b4d46c7ff4da8aa8ef39be7575edf921161f6b325120229a0355cef09e92c
z1222541f71ec72b23e527dcdb44bad24c6c443231624fa2800b8061ec1cd6d61c8b84ddeb3c054
z480a99e2ec6858781f47b0ab19c4acb35d556d4d759a84b4a56f05b582dab168a6c289be7dd534
z8d41b51724c5a7c2209af14df16038b30a92fb87ca2fc477453bfb587435ed40f0f6a04837187f
z381c1d34e0e3ce3487d9b27d92298c5d5ec23f1b7590fa878751431f9a62d012870cb0b8ef70ba
z34782f40b360a28fdc05541653bd64158190bf781214285bc13b7555dba1898d93fc3caec49f00
z169eff633162579193f0682004b5b7fd5aca6e11ad877f1944411ecf7f89ad2a618d70da624d87
z1d012f36d34e6ffcfab6f64a3532f943574554495fc885c8e9449da01c929a644d9d5566669866
zeb276adb9f7951c068fcaeaa9e6181d5907751c99615439bc86aebbd0e38c45568aea3d3f5c5ee
z5ee51ebd1946524127bf01862731e83c527b47fe63f9c77fb4a8c930c53647ae5811b7728fbe3e
zcd85509cbd7e59ca5c81b6bea5bcfd5d3523dea5d48e9d3969abe37f4095c63b67e97fee57b0a9
z9c5745c67692cfba0f0c0edf8e0933787b10a2de2be1b5702cae12f9a2b8c9371fb67be41d708c
z1c1cbce0e555ddb0df9d0481ffa30fe958998f6a522693ca091cd3f1857864d78dcebfcf00bbd5
z59a6c5e36aff1cc3fb5bae20336ee01bcd38cf2a98700ed73b2e7ddae652ea1f30d4064afbcb47
zbfb17b082a38174d1b5350682b5bcfdbfaf27e7aa9f4a5df1076b9b9a642e24d688853c76a9c7c
z40cf7695af1ecd3993ecefac1480a38f33152f2c43e91ba34a1f4dd38731f0ff46e945c0176e5b
ze569266360975ac1de5101b4e7a040d88d38a234c090c5af450386ff227070d8a93f85c8fad175
z834edcfe2eda60a8d607a814a92c72f5601288fe093b009234501f9bf6e9c92daac24b471c5192
z660b64450fd09946608f73cabf2ae81c3368366fba60c91ac0c949a912eed81de57f40c205234b
z1bca9fc17285113c8c3ac07092f724fcdbf0239b3379f1ecb57ce18274d88c3d29a25a4b5a82f9
z86fda88015916b2793971780c98dc069cf1582c96072bd433432225133f0db359907bf80da0243
z6429a0739a99449de20ebd5f74f2f26145e4714191c81168e13fbdc4f622cac58dc596d6fd4035
z3593aba81ce1b9aeaddd9580322efd8af576641b33652a075c1d5528063bb34034f852eb2c610d
zcd1eca908b421828db432185a0b30ca33d292acc5a370a7d70bc208357fe5eedf856f8e5aa854b
zb9a9b7bb433185c6996bcfaddea6a9fd460c51c5f26d7376e566c7866da569fa347fa71e810115
zc1b9f3af3b89070e84eaf7172186491151b4a6cb0c5e0c0fc309e7af378f20f315f4e1cf6ad15c
zcf1cd32738c4001efe2fa43eca7baf8198220d6aac832a752703305981c3929c6c96fea99e5b2c
z5368c3eb14c3ac8b996c66fd85ae1c21041086550ba4e5cffdb7c506e29c60fb4a599b037d4547
zb6374a4cf8a480945cd8680a2072f9e229d4f80b4815cd69edd7c75628cf39c3338151cdaf68ff
z970c2e1441b02ffb48b2f0e70f6f45690b17528b88ab64c4f90140bb7022830fb1304e88b5957a
z128596e3a278d6bd7ffaba96ed2e417ea81174297a33487e3eb0d2a2f8184b727cf85092dc01cb
zc06c6286800b11073a634b83e5c4318004040df730cde6a841d1d5b8f29e69e0997a217af1efdc
z6af91e63a22d0a8086c7ac2bd1aa99ca7da2bdc3006798bdc75574698adcf5faa0bea6ad3fb903
z6303e2276be14e5e45cc9b5d15580c8ca3d928f7c4393c64adb3bd7816700d3cfba03f2ba1753a
ze05f679ea5b8284c2654720a0f9ef3519b2ad96c8e95cf86e58df6ad1bf2f1aa845a2c59be49ca
z62d72ee46b7b8cec3302bde952f9c35f08da6c0030f06a0d96b84478a1b20c532a9f8cfd14ba27
zdffc4b705f3189e609a19beb847690d74daa5b8ee0230f3d6fe6d8efaa1e035003ccab12380c0a
zdb51d68b30a3fefe0bf8e94b271ede40e1cf36013bef4f3c80748077c4fc5e85d4666ad69b640e
zf29d30983e0f18a678315c766423d77a7da6f36b70ff5c5a74bec353a4f3f7483555608f013cb3
zd25b572beaedf93501d60aed53adef4eed29d1c48eff903da0b637006a5bef9813704bd4beb21c
zdd93ee85c704b6e882200a2200409432087025627dd1a9885f9f4e8837d97fc6476bb4fc2cea2c
z3de4835c34898cac28c1af81723bcd0452c61889b1d9ae3ea86df7ac25a64dfcabd5f4a2119f93
zf3a2d7e6f5b0ffbef898738c89873d07abac228852c44ffd719351a216019606489fefb6ad6c17
zb9ab4fb4c1c492ca52a0ddf85e9b11216d22ffd373aa705a5cedbf72291ab214afbc0a5bb5f1f3
z630410cd7fa1936fd6826c682540647f1cfa29a9fbccf14d99672401eac3b5e7eef93a06691358
z949585adc9346a2e264d5d9525f6a319b78cca95e19bc51837936441060710c5ec7e31ff80a52a
zfa2865ec8ed9f46424566f59cf4dc417433a965da6c9a3e98b06526451f13b2fc9dc4750014ea3
zba4ceb07ad20f7a5653c4dab0fe0007d32633edb0d524c0adc84d113cf4afc77eaf9e97ad2a104
zbed8648476ce77c63fb8db29569e28f9d2fab26a7f5bf1664aece8ee6770116b2f6d6d75ccfd84
z3c8ff6cd3e0530f4511f53b856ae9529495a7db02a33e56d65a888676343e3ece6a833df739d97
z1d4b3ebd34aaf4cd895d0bb6a2044fe61c5ce7091c7decde3b89cc72b9a926854a349d48d6ab2c
zbd05b379a9a6ef773eed77ab5881423deb27dfdd34db07e348d18913b863689bfdb0eb1252db8a
z80f85fe0447fb421b50ca80af28e1e425c668921410b77fbed61a88a07fb9df1b2be721cd328e7
z411b8efaf02e111f7458859e6ff0cf85aa53dc556e58f3d25cd16d6324dbc6644a1fae0edd3ce3
z7892a7c6e441be697bbba8c9b9d632e346366f20b41cdb184033f872ce4754a48bcd836b3b18b7
zd0592abc99d57644c748d14c4a58ff599ccff914befebb48ed3cc0f8e2946179c6407232a8fe2a
z4195ecea0295a91ccb7f5b1ca330fb91d96b816cd44d2978c73332c7675d9cea864331d55ed47e
z07d06401a13914710fb2f2255f3feb2d137fa023a366dc78275f6d49498d075da4f480b12831f7
z1bd8af56e5537ebe4a0296b744aef142e957b03025749dbe9f3ee375c89ec944727157c4234ee5
z140ba03542c06216f0ad962ad0959ca4664c27cd4a81c95d8345257ffa77739520ef45d886d608
z87c87145c390b888d871ccbb8888efec7db90835279017a2559d1b3548e5c06c410158986833f5
z5c344fedf87d1ed5926edec6fbc8c363665963480061f302fdc25ad8d2072d44b8ded1e3ace3d9
z10d22e1e79599fff0f8f5580cc273cf509747a0496f6167cfc345f5d091c3992827c5d6ae80f1a
za930e1910d58d72bdcc21241650e4da60d85a0013f7fc01ed7db6f6ec536013066e4bbd62c5f9d
z7c17eb6da4be15c31453b62697c4e85742e91a1efda7ad73c93a4afedd945f2ec91164a2b690ec
z635f5c4cd7ef3e86a94e37088b6d4fb90d6e5302edc309a08086da544d3865f67ff3d899ccc983
zf0482a6f82bd63a3878c0afa2427cba5ce7ba0b6724ce4d23c438977f1b5f0056eaf3e93b434c4
z3aa31417ae5db3c6c0407d5f81e884c2274905e50f2124c95aa89909eadbeca6ae32c523a98262
z605cbf568956b08aafa89795d83eecd07153f913e6452552101e26c31b43828d8c3b5aa4118d3c
z9d16314ebe3029055ab7563ad9f6bbba8b09e4ae9f971fedf4849057c050f10598e1db6b8f8533
z2ed2ac09b49ebe8a1ae8fbc1a0891a57313aaeb14e7cf7e8242e71688195286dd5f53ef0560e51
zceac1691ca675a3a0acc583612715b0eb4c4e9ee47545de2ffa9c925c4ea37436a4186f3ad4307
z88fc85aa333d1442b44bfb405886711b6bb609303bfb8abce48436946587fe7efebeac0d6db310
zf368e6aa36d492e984ea0bc8755e77927744a8d889ef15311f3fe930de6606b1264fbbdbce9c9a
zf5cf0172da68d91b53587d0fae8a5efca607f401cbac5f898acf8e96f40acfef90b63fcedb2625
z000a93ead4054f3d96aabcefe7a50521a9f16fb283c0d28e53357292fe2fe8b6508a4e2a7d44db
z1b6a7c378b997f13e1cfae88ce4503a4472f698204f1483099f98b5eddb2befad1ae322c6c4917
za3b0c329ca084f8dd1c82c575bafca73aa0c2a669bfea2a8ee21fe72e8be0ca7ef52be85abb401
z58acf2e4d2c3b3b824f9fc7858e54f6a10bbcf7a5757cc7ebb544a0b7252db01ae3872833169d4
z80132d927b69e2e7501bad1ec7174f43234f1f8160a746eded42f45e29eff5b313a47cb8084eee
z910c1e5ce2698e42bdf56c38510269917b8f1767be63aaafc80e6f52f1cf874602410d3f45a795
z4da7379f51692e503cc4e1c2860a9b905e894d587a399aef56cf2e749eaeec351a90f209d0f736
z4a72f06ce57cbf0796175d1a2ee0ebe6244109fea17b9177b224985ba0e53ac06a90e27b39ee89
z5d7d319d6271595ee55e47ba4531426fc3860a456bfade0af8c9ee72e7a559e461ade1eb879583
z4561468d8aa228d4e5c2455fb7ebaae2cf73c948b3c44bb0a4bb611b127b251782e6b1c4e3a3a9
z9243ef8573d72b5baf78297c661dceb37e2fcb587dac4cd2fd8be1046667b9910b450ed9800784
zc2e342b0c5eafa8ad004475cb566edb1443a8df731acafca07c7ebd5fbd10298e2f3fdf2870f7e
zd29dbc18cbc675b6f62e52e927c3402776792bbf11eb86c256e9b4fd7171158a9ee30e2456be11
z919cb5a2ee095c332453511c7b52aa92dda1adcf943c028d0b2960ce363cf5b2ba95359f46700a
za4714540ced39a1fdff83b404e11f29d22f4f38186104b365be04868a0829a635f366719cf6dc7
z85cac42191a9d4fb3191d5a50dee4f883088f51634fc007a95979410e40abf1fd932adb363bb20
z80afc0fe964059de73f5ef06f49d13131e945a65c79cc3d31b34a21baafec401a7e17a10c1cce1
z3aa3eab82180208da64968316721b1871cb884d1a660849d1bc1f88a14c5695fb0ddfbf22f9068
z2f8a2c47b5d1ab3e71994a8341076468c48517a5793be001d8c44b90b9263d1782517216bef276
z01efca5f573a97f7ad5f8417237dd9f401d519c7ab49b7bb3551093cfbb642bce6f9b6ca98d881
z8a754c3326e31b85ee336c474cc280a000542b99e6c1f42ff93b2d70105191b919c25175ac2e78
z1c6e21055cf7088a6ad2a52128add061c1c8103f10eda5004810abe4c43d7f7fc4f79ccaac6d7c
z2b24ddb8cc89802fc5aabe3a739592fffdd4921b5cca54bec27fe2465e87d01f88a3c7407eb586
z2cffec9351f67e40b6b18dc2c1b8ee546ae38dc9bd673a6cd1804e9f3351cfe66b52605c8c02a9
ze9c78aa97b76f3d8d32328a2fea5cbd2547be45cff3ae400219b512488e34a39cc9fdb2f0322b3
z07a8206d86d05833d0adab1fa462b1e6edc3f104fef308686b1e4dd05e8753c1548f7d6ce88c7c
zf195fb98bccc7232f46223f2c219197c48cc3238c36e6f37022434a7e8cc00be7d389da13f47eb
z670a883923989bf2a772dd38cb26aeb25a25f6b89b88994c0b70d01682e68f2ccaf1a6888d816e
z715f5a28f97112fccdf9a399a0d35c491f6316c7b38b6c467638068c451b25967a51867615c6be
z7988ee9e3198edc86995988674b0e30b37d48f0ae13b80cc361c2b892fe7cc84b11706a621244f
z3b37f2bdcd0f1df230ab2f76e296bd60772d53d587e6674530c68986af81579fec7a97de81ed9f
z389ebab0ad3398fa82ef5f7336814c6a305d0a0e49b9f2c9358ef1765f7e901d50ad1adefd1d40
z55aa61d1efb1634663e3b9e48651c7455672979f05f000f24ca239959ca25943922e6eafcedf58
zb870cc152c0920a3ce6a62d112c2a2e4a9f0bc5df3c3bb83d9226cfbc920e79ca25fe3d24f9537
z54336efa3c380f4dafb89e7f2427d6a286fb11b1c2379a130b02b203ed929a80d03da56dc358fb
ze4cd118f0edefe1a737a8c0c5b0f2a6d5250465af7ce2e74ea9fac9ce07929b70abca5f7248ba4
z24a9e783c5b53da889be527d59b835f1235a6d6d652cd5f9c78843e5bbb62cd7db7dad0895acf6
zb365c5d313523ad044a32f4acdc4a6caba0b5d9ca14a7f705e2e05102e8390d60b82eee770e1c5
z1cf2941ccf49ef37224e920736de0edd76a2bdb856e8d7e6a170e428713c112747506ee0c06915
z80866a60406004993166063504f6e7c1d4931eaaf3a09ea46772011f10f94ed830d5c8d0ccbebd
z68b067ea1b2136124394ad3557d31254c4ab12e0d4524c04ed0ffec829cbee545df37d47605263
z943659e30f04cc91fda71f1afd4d9d268dd44976e819ab477266512de86a27b92d091b80186e5c
z934a6f26b122baf8c5178c31f6e016cd96d690f6e172098eee5344ead511c9d8a09f8f40e80275
z54861c375e4d05e0cf3ac47563442b7155cc20eb4b5bcfcb2d9ec9682c675fd02ad037cd18772c
z2f9a82a7c67b2be0a8f3e5c1d946b5508006782784b9017d5668749a9cd2bd848567489914de32
zeb679d2a56331abbb85608a4ec35db2cd739277d2202c806766ea22f5008dc8db7a9d71c6625b2
zd8f502eac42f963ee269f9410a11d97072392c0df030bbe248b6b2005139edd097bf0278c88b88
zfccf1d774ba9a076720a1463b40267adabaa6692f3e66a803a81d9e04c598ae75dec65382f9508
z57da335ec01dde80b07866476e67a8a369895dd692598d2f02496124bdcb9aa6d304e70373a87a
zb86d60e110110ff0f78e3d4471637f3689478a7843b8896082d0ddad3ef165272509bc549c3a22
z3dc177a640343cc301a797527bed3693ca721c8ff687e13390d46bbf15e8752e0e5d535480f133
z3d8c5ffc00a3d2ee0296b694b8f6837033d8c4aa72e7a18a360f110e4b82bf3b634ee14a9fd58a
z996cec080ca2077db0508737d16cff148f289e1abb0df634cc2fce15477bb3ec45f6d6d4db3028
z0d3acdff9e8e3bba9fc450352d4859a3361649e3181cef3db6121b65489b3c73dfbec7fe62c89d
z3ae882f971f61d8b861fa4d24503c490872674f30dbe086682a705408fe19394882f8486b28e9d
z22f08cbb7fb9f0df920f9b92827d443bd39f215416b4671fda31755bd133257b8c7b96da68a565
zd35a8e9f3059d2b83cd8bc19f037c9d783a485929fe60344be8be58606ea85b1765d6c1928b7c9
z2cfacb2945bd7d2659bfdfeec44aedff69a98bbca0752bb952a876c651a7e4701f61bfcf37587e
z0f42f640f75fe7172e8dce8f6134893148f72f2a2237cc200fd3cfd158eb10ab7ee28e3a8cc966
z6ffe35783e9a37e88664ed91ceee59266af47e1e88bb4140f9fefe8a41013813f65d2ae2f9d16a
z3c87a0815c6806c3f2874c707e8f745439495501f86c5632d9a1ff8330d6c33be18f148f7bd153
zdf682d016487cac21c0a94e0fa1c35aced5cb522b9d62af31b41a22cf4d55a402f73b2332ce9de
zef32613499938b7d991b1897b503b7c03b18be9bc0d698b95a961dbd9e772988f360a14e10854e
ze8c996d35d9a7256413170e1d1a6f44ad6dc70f62063845bdab27cc77bc0901da7fb50bb0a4b5b
ze8aa873e2e6dfa4637bcdb2231a9db57d1c6267c89f52b8202e86a732359f957eb18fcbacb110a
zdb2e79803ea657ae8ab5ff4abd2447feb32e164c085c839ed19bfead415744d56865a45df7c349
zfb89eeb3a4c72b6db4ab41a549f30f86abdf1e4c0f1c23396ce81d51c5d07031d791c10db102cc
z2b6d47170b85543721f95e28ef41b594c1aa6ca35f99a91380aaf2ec478ec1c3be00a6d97b9042
z960d2fa35a7702839973af04e9c7450098385c207541ccef1a19524c60690c1379b0d16d7be553
za9b507da4f54f7a9623a532f7cc415cdb6456fca754a1d694ef7308ee3076e780bd85cd84eb26f
za3fb86618582fd4016696b48292c088fb8715bbcfc6c0ed1c736a9e4c07a41451587e31040d8d7
z620e0985e86d77575f59c5fa6e1dc98c029cf02f2bad551d6b66aabbf44427029819af8b330277
z3a2d89090164e17d2b33cf72ef282c1e87565d65f7ce047a47d774d5c2f4ef395fa33043f87092
z955d1e742c26542885a2c3a97020132edf6a22663f2f08c7db92aaae5eea8bfaa4d778e5cb85db
z9c35806ef29793146f0671e537b9a919b8738c1b94c7aa6afabeb07cef2f6c891999cc33861054
z8bd6f4e8024b5fc103e22034ae1c9041a95e73386f1104ea290148699900a954e9ad5e88332e11
z6cfc6d17ec8c04a0389b5281b3858c47e4468bd1a08ab2ae2552a00a73d18832271c56633dd46b
z7ad1986a706dcdfb32467ab58ca8853ab2d908b370218caad8bc972a15c85b9235a5b95405257c
z2bdfbc48f5936490e749cc90bf26a02ca696558865c5d92754188565162c9e1d3451c53b026b02
z538c53bbe6a39dfc6cb47900bb5c8e0653c056feae1311497872417db11452b9fe3cd996650143
z260e72ed46e4a9f74b18637db45faa6795e9c7a3db0b06f1127dd677ae508ba4f1f1a68cf26898
zdb2d62230118071590546b7a4539a3cbdedbc2b3eab7042878c52e139b70347f993f01b80ebe39
zdf66f726045d2ab89e279de1145b92bc9a03f74677582d1ef18de7c82b37a4bc186bddf37ffe7c
z1ada3ff6976966452b301cd23296e5d422310a998cbb07a14345da8754de47e54e13bb5c8a86fa
z16e9bcfd0dc70dab1658b25e48650ed1d5a25255636b9fefe7ae88d9005b67e8021b07ee472df3
zee2bcd395587db4c430961beef95b41bf53e8dba77707d430213aa34f672dacccfe097649f9dca
z52ae957231120c1445a40b525e764988a097e934e9790a104729715cca26312459ee3ef8868b42
z2a38b9c284d748ca2042f33e5e594b5dbff9c183a8b21bbe3d50893f90344a6f7aec34935da68c
z3c9ce6f58f9d62ff1d36f4b4b91f3ea6c79fb4cf429920f2f028c08643ae72281799e919f343ea
z0fc3af47d7c05ee7f055afb603536b2f6a274dea747d77fbf2b64bf3ed6b889e8d43c5f94f0c77
zcc9ff4d28191d2a93d00fb7909584d4fea0caa145878ff83420a77bad7e227eff4f500bc3085f2
z537713dfb59e2179e82a330d63d57d485dc7b1e60e6a12a1894c87736ddbc958bd29d32b80c61b
zb6533e1605762463f035432a2f10744cd1feb43cc3a8cf2eaca6b5e8acf2083b7c317e85fc96ad
z6b4e0465715f6bd4d69a728db699c68e355ae6037920fe263121fd7fe60be5841695812f7d0809
z6d994e89f445b2138ce38ec05933b6d07e42382756c0af30a5eb2bfc45ba79a9153b33bd84055e
z9633d43fffd8610effc4f160a9d42beb855a8b8ea7da84bb3bf5340678b529de0482b4a9f016cb
z10f9d42b642ef2e5bf0ecdaf4a93bab3c9989f182643ac3b09f113be53c1c121360a5132d03a21
z16a3f95541eeffb9c79f6f9b32186522de78d76e1b02d8e2c0859c3ca66d51dc39e21922015667
za840f569ebf4474f67ece89a01125e44ff40965866766d3f90ae4e7169b93ae111ea99ba14ce74
z6d486a944616f5f7fd94614936acd804930b701c1d0eb5a4f97a5858798501c2d16d94cc35d1dd
zdb5f86f5b7d229de9bfde72f5cd17cb28bf73571ff7ee8fa038d323a28bcc3741d8161bbed03ec
z467b4b5d076673d5eb3f248fba493b41ba4a08f7b84f4b95275c753e33038944c66459296a4f67
z368818a85eba3bc9bd683d6d5790454b76282307f01780ad0eed928141e695f1e9218141732514
z46c7bd14b9e9e92abe43e180a72bb957a1775225ff6d0e74229cfe4d74f4de448b51e72fb1fb85
zbff6452205cf966553e09b6e4da0ad1d43411ade88714181ddcfc06a4c55207937e5a47c655af1
z8c796e1a3343e1063b2547e303d9810fd0ec3d48a0b4c045968ec60110170b7d27169d719a7ddf
z4228a01c2d500d83e98e6c931d2235644c788163dfa6838733da626caf8aed9643cb9cada64f8b
z796a03461e7fdcc04cbaa65336015c0113ca7d6485e52be425c2ff2e8da727138e005a329c06cd
z95000b041a2642fa9c93d5e359d1a24b71d3f16e2acc785fbd759f0b918de54e9c1db5af6db9f0
zd6d0c68c86f15a782127b24a705b2d78f6d30b0acf47d49048dab3afeb01938e05ac2cd914f12f
z74f8e487362ff94ffb999298dac6b42ffa353c09092ce402fa85280dd6a31713c75e74f695fc08
zb2a6f6a8aa8c86d231a9d45f065f33be40d0623e4ec6903c85771f2c9ac3a67ad6b985510b2835
za121f65937dcaeedd96612b29f0ef265d448dc12c94d1dc8dd975f18d63293a437540aa0cc84e4
zd8d1c4869a0ea11b4f8defd4a2f193c471a4e3df64850c50878739ae7d59d41aab49a35c9d671d
z31abcfaf95a24ae8c09b650fe9f4e56cb6a7cfe5164b158b584cc2654b6ac26fed15783b956d92
ze783cf81a149edd854382e6599f40289ecd5a3dac11a5a8ed82ee61a3e0b2e7e470f7c6b4a79a6
z08f4f61df873599aa6bd1ea27ef080ed966db9052ef386d723c1e6019652ad9447d25402bf5e75
z111c968925104ea2a153ab9dfca84adbaaf57dcaa667348eecad115044dcfa90ccf2af1ef9888a
zb47fafb11142daf730d1deb5f32ff763fe0bd217fd7365f2eba912209ddef2188405be426f2299
zd7761b8548c899e456f21bc183d78e36f89ee0ab3ecf4aacaa62fe60849c19a7022943e7fd7a63
z469c9fced458493a0935ee4f3df33e5c04305384718b4007c46cb40627ff9c6e8f08abfba5b291
z422b2c2014d142cb271272ac8800fb4020e0aa1d7600a70acbe222743294eeee628e7007e96bdc
zff4b5ffb01be216104fe65d4af2b7da5f87e1d9209c1446ddcf0d0bfc9ad2cdfb61c345a27a97d
zb47e84319c38750098b3e3935e88561ee3148f475f951e832f82870f5591b86ef1b92c0fb3513b
z7c1152ae848ed5e03c5fd1b8e3c866de019c33ae0526a94ec4d1f650a72a9aed61b45ef97c71bf
z7f003d090adf655edc3aea3d1ee57c171265f1e6745b88bd0a2562e3c833ba6e5ddcc2b51026a0
zf1c0956a37b79a099e8b9a961ea037743d45c4f3fedaba1e15d35c79c3c7344b20c74dec3dde2f
ze60c75ef293b53f782d1892cf31b258cea188024182a7768f4da6b6e8a97d6b29d5fa4d25d02f8
z0cd82a1270220e730be26a5737e9eb85d045029195a2e7095e403cecb2e6a2ad75d9179f63478d
z2d2a76c21ab6d4feb0afea6c550f7515052612c0bf920ba2912c09fba8ed1747a8d886fed70354
ze109937afaf4c7a532c95b2509cb82d6dd68e0771182134c4736b46f2b17350d40ff143692bc02
z3743a6252f7417ed2ee295b255f59660a0cd2ae57e370509ebf3dd4789542b8243f1d8ec0bdae4
zc5ed83ced6b6454838e219c7b30707c2494a77949a06787233983e360847e592b593c8b66c2e7b
zf2c1a4b696b38186f65e1d0d6d21c70a8564c44cc74286a9ebccb220f192f2e5d76bbca2a63376
z4d53c3ed5ecafeaf2b6f9f136a4492a4bc0534a123fa0c27e60c1b4151e0d9e38448d415a30185
zf66da3450a99d10327b579a5c438453bb37e6c92676c1240d6d7b6811f32585020bc28b7de949c
z91d27b2a4a4445166ca342aabcb2ed4e0da2c615c88dfe63e84494b6eabdf0b7c5c3c5c9aac469
za47eb7f5e51788bb112b8ef6e0d56c12e7f04652b819ee1b433f66249b5395c13cdd7bbbaafdf3
zbf2022da1e3959642fd02c935b96a6c83a472132c7019768a3183e90b8b688b28368cfc030c35d
z6da6bfc7f64a6422c56ebc69f84c802159e43dac435e2adbbd0592c9a71bbc8d31b256ba1ea71a
zd5bef3ac4f1302b5a0564cf6cd1c04c5fb8d7c29f9b3a6da33dc5515def08a550a18f3505f7ea1
z7a081bcc7388b2c6f0692b6e7d48253639e7ff6da67f12bec5b4ba0e83e4699636a1e3042121dc
z381a733c27572c05f046daac3cbbcb07e38b43dee6f1b70d87607ecf8253f5a41f3eaee3976aa9
z3eb365a73f9df7f0ed7f16140cd12f34af4eb5677e0e55e278b4d2a9a6d2a35496fadb0df6ce1f
z0437d9fe85262291ecd9fc3a2392bec5210bc8112351e9394452923a6444a59d6359d50869eecf
z9a3120fc0f6b4e60cfcd3c5ddfe1e17ece826bed5371e50e011c4c01bc3403788d6de9af75da73
z98beb5deb081ef48c0768ce299653d184f7f728fd1c436f0f008c977f604a2b9b37b11ed934bbe
zc209af6c92fca2272a8a3a60488b3a564194681793a70cb2c0b90ac658d9213e41cce69280a669
z76422a22b3305a2534a06c2ac1d6d6b9a73916bfa846c83969e6b9a6a90a9502693fa2841f38c5
zba18476f1ca2ff05900e9753015f292ecaf216f8bef6e81a8b091c0627ca0318cf872b99a0adda
z81c9e9465f6e733ba2dddcef26a7cb817e1ae7743aac4d3edc852af88250c1edff4f9437d37a0d
z1e2cd678e64b7d526a206d990d4e4c0be2342512cf8e406f709ccf92f02fde0cd97e868c6ed25c
z4c899bd9530275fdff3f4b73f95719c79e3bcd37b08c381c79fb4185d8d5e80397b5ed4eb62ca0
z4ac8fa4f28f4ed57353e3731a99077c3b324e259266563be273f83a9391d9af93cf21b614dbe39
zda2a1d23191d199f171fed4abcc7ac92df93677463c31bc22bd626ad3d56992d81b47309c03fc6
z7c1afb13f99725667c956231a6053dbf6c8cb832172e35109a2f228a50206705b75fc78dbb1667
z3d46a8acd6e2c110813df5de78bb35add5c02123154e859e2e9443cec64b5ff88c171b0e8eaf89
z77c96bec3a598a4025b2d56cbf99b3eb4bef11f0599584b1e1a24a0898a24bd2880077bcf18a52
zcb2b45aae41bed51dd3f376c96fd3b524a3f80a32c40a4028e79708a056f67e1b0035acddaf142
zb28a6b5d28b6e29ccd8cfa59c2ee10261f668ad67a2587033833af520b5035510f18f8e3f29f3c
zb2ffe579f5ea2148c01b18425331c96d8e55edff07ee4ff97df9b3c6766b302139ef52107512ae
z2689dfe57c3b2221694912aac7411009249f397267e41aee04f933550072ae1dc792992fb6c4f2
zb184ade49f9fcb4dc1ff5bfa259e942092db9f37dad70fabcc5e0e132015fa4829410257cb7d4e
zdb359be3d0402cf4952ca27e0acaab0ef76a27b92d38ff48e13e566bdeb86ceeb3b30621db205d
z7ad5db7ef338e230c269a43371d6d82255c53b2cb299c9136d663afd7f117079ec11ad83bb2a14
z4fabde83a72658a40d9f35099c680ad4b9347c6545ef61aa2ebd80aa74892fb5843d8ae94a55e0
z8b7dddc924c653647814c34d177ad248732c2550475dbfaf23cd7df40fefe58690e0e478675afb
z2c2c3e52100916d03589f4914fa6bc827ac1948f09dd27d24670a283fde0e70ce39f6058a8df4a
z1752e5655b63d0be93331b21d1a5abcc347443f11fc205e98c8611eb4ec17011365f3df58f349a
z9c945e20b7f85623ac8d6439e614c82535177601b61cc5f7b567eb31099da710b859e3c0d5ced9
zf27dca43682422734f365be9208184e876bd7471e04941c40bb85a829cc4c4395396bf381711e0
z624d2a9acecf6b371eeec1241c126b6a70bb53fec827b529053feaa2da3336652d4c0f0fbe49f4
z178d881ddcdd802a799615252aa60d7e3f80b18bbefb2f5c25bd9152806fe4a482fb763e37850c
z6510a6c86e209e5fe48abe2983b8d9e28210ff7a58978dc174c695eaac320c44497c20d4254284
z1611fd60af09b7e71b06157e890141b9fbe1e4d125021f76fea377a990bfeac1a3407099213d8b
z2e65bbbcc7906dff2981421fe602e507df3c96043a4637b890ad76d34a2397ea3b202ffd6b06da
z102140a61d42a5c09aba05a0f5cb14e6c805d6d9a20914f1da64bef0dcf8db69e4109e43d3e2c2
zccc96f1d7ce886c9dc9a1d03b12a2ae7689f3890a87555d7445506e7de7fbb19cf7c8a9e2c5420
z037866a6fbeffd4df50bb4e9a2180c0ae36cbb1a9e9d8ef50927ff94e20aee2a2bafe96e16315e
z55e776d49ba792530a01f28fe9640ab3a2659aee3816d1134af9fe700fb1e846a6df0442fc0b07
z39861a035e65b191a809af6f2924320dafb64882f0e0da593b42aa66b3e60a968302c25fa33e05
z7c850d582275eb2a7e390b7743c92e452696b1a74808fb823c6b69e7e607f15173acf54ed8f951
ze1f9d8e300c6a2caa78af82e18a81306d247fbc2fb3b4a9e6759d801c49526eb6164ce94ba6a4e
zf11ab7c91441c4ab6453bff848a0c6d2fcc10cf26fa6cf758ba5abcebb8febc3bf5053cda8cd97
z911c721beaa9eeaa6fe90dde3e2ea3f8781f630350c94a7bcfca6ea4381ead6700f11e535a28f1
zc8df4b0d986526da0b0ccb5a89a73f166a5be83275c811ca3b3e6ab1777cf9f1043f56f3b10e17
z008cd2ef127877b71c6ea30490abef50137a83ff7552ab0dbbce7ab0581bd6536c6e47c97da735
z0484c39564d9832247bad5f1f1f3819b5bc257790e7b9f1fa75bc7eb38ffaaee434523c9792352
z246e6df8289ce224c409fe545df8a591d56bebb7c3f56d16b695d3db55d2a15b85fa59613eccae
z7d7ead77c8f12410293bc92052126a015ff010dc45fe80318885542532ef5fc45a837e3479c0ae
zf601b6c7f02d81e1716facffc22e283a238a0c13de6d6c2542b57a8c8f3fc03362e8164c758188
z4e465badd628dd762aae8fa16da7ca2995ce4cbc690c9c8411a692032475e8bb23609bec6cb3bb
zb326ba52cf35735739a2e13cf97ebf36bcaf6da4ac1bf10f5049393ce6971f9cd1de62e5de11bd
zc05a8e41bfd98d2c4d8fdd55d04490428774724e07f314fcc9e2bb333f79138048a23a0af4e06f
z34fccbd07ec6814ae2bcf6ea3f491bdb1e72268e51219cd45be9234332d2f859ad2624024e9366
zfddbb314bfc373bc9f824c4db4e3010b37af6d9432ca269e6f7e27fdc30b16919ec45fb6446c47
z94f2982e986e4a200c9ee698a71e7bd3d99e3b6815f6713e5016219735e7d65baa22f75742ef21
zd823087fceb7d94117472787c9f003b1c02166113f9cb1bb555cd792a28e45fe6315f0e588fd3f
z0be914e3b8a80603d8d07d25b0b21c2d4459aca64f20066b993048a5b955727375276f762bc392
ze7248dd43ca9551a49b6b8da57f37dcdd74865400201bccdae8d626bc87c860c731957b7502279
z9870a2665ab7a442368e83b337912ab44a2286a5acb813a1e46f8c5f66ad9849db33673e9527a7
zf1e12012060921923c9133dead963902895b1db7fd1774ea37a974a7675acfe8f1f5e1d28928a2
z7bb98ffa96a43d57adf8404ff5b8f1088243092290ddcdab7c4f8de0bc28194848bf8fe5c73215
z800c2e9b16389fcf1faf5c8bcf2d0be77da966d7eff1f260820318e1172a9388509f47477f5b11
zc48a7ff559570a75eb17b1eacafdd376f94badd127d5a525a945739da91234224460d4935321ac
zfaf91f2163bbb73bb870b8adb9fc1b77a51439f00755d61b23396bb7ffe3e0e874036cc8570d85
z2b73ccb6dce36a14d89a86ad560f42ca9a9e60f6c4ab79cc96d28483af4047843e56dfb84fc9ff
z5196128333d72dd56595008d7057326178f05254131185bb0f52ce04edc40ac623993c1bdd90ad
z5ecffdeb0526d319d0e2a03dca326db4eaf1b405522a44ec6da9d98f3cb0fad623793441426cb4
z751333d2a04124a1afd96c1602440e7ee8b67d1e72fcdd156414b33d239895e23f1ef0876f2046
za64c5e9b67d47c24dbefa49ceb2ae6c8d7d2d80f5085030ebeab74f4f78f34eb08975062c53baf
z417c10be3232a4b2d04c336eba3f2672e28ad6e2c3d2519819647cf4497c88a7900338db874250
z718d783c935a810464777b1bbd5ebbbdcefa128616cc94ff28f461ed1c57aaf8a0aaba4c3e6af1
ze1b8a68181db8f92305815bd16af1becd7a742cddd1ea7d9be07c2aa505f72e4cbc50a7b5f9773
z967ef3f6f718acac1268e9cd71fe41838cad826212d7229d6e5d57db99c2d3279e654e67821efd
z75d0939a153d5854187c74bc5ce05813302a6dc8d027c6fa6cf14ca023b8af11230a8b4e3d340f
z88a1f36c60dd41f14206414228c7ac4fcce912fd2637aac32a91c71719f1214aef12d157f12353
z7e3c003b8efc4ce7416b0a8a4c2e08f541960c52fb0fb72371a366dac8ceedc791d5ab4e6c0825
z1b2cd60a885f31549e3308c020462b93d038687ca9090d00e97fb42ae752514537344f192823ee
z4fe0bf18395c9269a3a6bf4124b888a40259d84fd86acea76908fc35c47d7eac549b8abe5fe783
zc762439cc76c0e7ff7a2c3b3c5bd433e0d46e406dc7df1dcb81a47080e38e2105d11847de5eeea
zf8c9fed0456d693a3bd3fcf82f4695d162a1d0b475541868a29976a893067813dc719009c0791a
z3f0f544b12f64d1c5b21e8e3103c63e5b1662e10b8987791775889a58edfe6f1eaf19156dcfac9
zdc93f605a5a598b816fd3b4306da06ba7ce9ccf7a3ad93e8822a59da792f62ac337c3dab1f867e
z6d3ce7a4f16dc2d7adf3076b04baf0d273914407a77ca87e4ad55e03a6b6894374a175b869f34f
z53d4b913d18902c9c972bc0a5022f1c32de7c35b423f023d83f3525739a3de139f4b71f4f50bcd
z5da59d2c4d161af0a290d1184a1e0987b8c0c294a18f8eecd8c9bcd807cf97aaf6e47da72cf55a
ze12376aae8dfe9f819efc7cae9b5681e68ed5e693dd0cff02616ee727cb97746b88375059f11e1
zfe0af28249f3bf1d0ef2ffb574bba9872762d15fd9b97680a01110e7285998314395d411d385b3
z0cce24cd8cb3d6a8a82c775187f464b3dd26f3686376a4b72030d31bc5ab85ef0eccf988432391
z381ae83ff0ba9a7fd9eb56add20558cd1896792bd8fda8f0bf62ee763a1de8f09dd257dcc76a2f
z9b42a0f6026972f44a7c990ece8e4e48462055238986d26466aa8e00e8e4365d26d6554c71e49f
z00482019ba0761f4e766d6cdbd4678715ef364cebe1467bffd58993c6b000817d013e6b92ca30f
zdc0eabf97c918696e01a570d15a89cd169673df8395d4479d11b636939123660860e787c1886f3
zc017fe914d911a9540b08747671004a2075dd9854623da6fc3dcc1f74db5193be24f954e152d53
z1b25dea6cac052927eed0a6bf849160fff863dbd9e19e8681ee59746ae6f1c69f5f8cbb3bc4b85
zfb17221bb4c0f5d1e598dc01a3c7a9a7ea44c9ce1138a246e5f011548c51178ccbcb77314b2687
z124c70d5f43740db3107dd1ebe45bf3172d2acaaf4f74f80ea184ebc89c4e2493731dba0e70ff3
z564d20aee203ee5fcef0f89cf341891cf873a14dca6028c77c94f61269c6c106af274b97433c73
zda3d85e3159ede9356da39f0674c9b7cc45d4a66c465f29afc45585cbdcdf04c0a8ff0b9856bc0
z915f76fc05b4b77e04af7bd0c54ed7e9390124778bb994f6b00b9738f113acb4523b31282a890a
z19cfe1ceb46a6131209caff2da3c04c5f394e102244bca6e1ff1647de51cffb97e62474da8964c
z736c924ce5d14a5c705dca9f42b7286cdf3b74140738cb1d9cd5bce6c9bf975f40ac8221455b9c
zfcba8b3eb1d572163f828ad22c13aacca4b75af941650c01dabfbba8e66f7487f1719b725ae8b6
z7deed120b720416552d80dc1a8ffd9d728b3d3cfcb2b2d4f4d45895f6d4ccb0b9e9769b581a4bb
z1219c6462dccbb18ce1db581bd04d55c1f78841b22d4fbd0bcaa5f1c4e395ee4fc75e623d0bcc4
z50a4600388deaef958283832c7b1d23b7622c25856724485908d793594772c24421eb46f22be28
zb98a2b5859eecf2fe041cfa10b8db8fa5ba28bee9515aeee24da14e07453f886bdc1d6c8ffc51b
z5988fac699e6c84f2a5de826f1690392565bee1150849225bad59a43a0e38042ef61f12ecad321
zf0c65203d16fddb314c67295698f05247eb395df341ec7c2c5180a744dd4ab3e5d7207fe3b870e
zcd6148e48e119a8d05516b8bd91f469d46d751c90f24e29f4b107eb03444f348917eff2552d582
zdf89b79c4bbd4774dfee5692e1816e06756726ee7dedac66341f3ec33d93018cdd70fd282eed0e
ze024e03cf65015ddb383527f2713a20cf06dc9aae60806eb1f242e4938e2873f22950f907455f1
z24283eaaff74a249a4411507fb2866b8db8f3a54192590bd44fc5772302a7923e5838d596e130b
z9ba3d94e02dc6130066a77258dd24b56893b4779e4aa2aef2e58337a014034740d7a59b42aa734
z456e296ed3aaa272f6d8ecbcc3d70e31e84c2d0c2e9057ba3ac038026f9969c56536f86e58712a
z336c929e1ab2f3bacf9854805b5fd0e816c7bd1d21ab40f3a19408c321fb1dadaaa05a21188c25
za836c87b932b68d0bbc63651f692c962cae8c85345d6a2faacefa50f2068d412721729e6e989a0
z933315ef83187dd174235c4620585d7bb3b982c564ac726a925a4d7b2f42d0ec93bedcfcb11fca
zb80395b3c389c66e463150b16b1dfc0b31c92ea2e991f41698c3b386c590bf3b3e29765ef8b2cd
zbf9d6bec9dab05ad5334b221ddfff285cb6e58d0587aad5f6c3db6ad57f5360497e26b3dda7e5e
ze3f83e464f21bf2e99667a548a5e736bfa947b717e408c1de9fcc6b50924aa2a91fa137042d4b0
zf068e1ad4e8b627a7aa0ec759b999e71b69075509771013f4f3b8a49a3e10e926c15c0949eee67
z88e3b83a8d260df47cde6f4e88a0a494acd48966c071da4754a4328bcaf8718febfb502f0738f8
z67808fd03f0cc1f919a9cfb6dc44f98238d77e05eec274776594b60cb741607fe58ebfd3d6ce74
zc05faf9437750340752b9b5b5f541c1d0576c62926de9c66688bfc9154e1a4c35e07f1f9579b14
z23ab3700fae68eb4488835c7246b62b8dae75fcd9fa4552c1b0bd10c658b50692e1c420813a27f
zaa74b317b38074f2a3debcb501ef559d6361a641febeacfc0702f55cb7631964ce00964b7bc5c5
zec878ecf13914f125de1d8a2078fd227fbabfb0f5fc95dff16169f16402db0e94840f269aa252b
z35b7507db18f915ec8c99a0b1e35bd716d1402ee5a680a067647464696bd577d71bf007915876a
z37ff9c8725166ba793bc2c9dc675c85c172ed5f447d9c93abdf66d5949061b57e68a3889959306
z4f6b7cc500d2454d710178f58cf481f7980fa5b5c77730517c3ca37b3df97d2c9300617318db9c
z4eb5985129ef6043a0c894e341f090dc2f90becf9bd5ee03d9d04ddbed493b07af226c841763e7
z49973b68868f1ce79533fcad85a770f24c9ba55b4554d945a6640fad9c60abb253b79fff7ed682
z83836633d807fca3b64a2ba8abf5d5a5c72ab3ea951da7bfe6fc643957c5b97944251ac9fa9f3e
za72df65772ce6472fb1fae8dede4e4dcc0646029e643ee7d6bf6281b69fb4d40250612d5449fb7
z7ff532a1c2ec949cfa35ebc5d77ad6ad61bb964f768dbb2b527bba62d98f01dd9e711c55cf9d1f
z52cd4b6a7dd8a7c35ba68fa279056e738bb705b2632ac9a11f0f3c5954d56a00dbd6151ca9d468
z1f15cb698b8ff746c6cd8b149fd2933b15cef427ead2503f7886c6fd2428bc62b17722ee2a6cce
zff11d5050dd149c098c46eb028e9543d48938cc3b7a4cfa2b0c39b9ba0bac542b2a241967a30dd
z61ca210344dbc5c09db73c4f4ecdb743549c2921dd0886e2b0669a20f70ea3d4266d8c947f7305
z7d5cc6d2e625a18e1557ecea579b36fb713cf160a886fb024210f52d4b95714c02dfd284ef48aa
zf528400841859b9bfc9e071ecbc6371faf952e5b9d7c41c7d2a0560373eccd67a490723a3d404b
zadef9c8aef65f72d17d73b66dd2b1359272f8f370f5fd819b5e093a2aa058b0e09142e85646bfb
z9a4f7f26a9bda2baa5d83809bf66a0b989969de23482321c2229cd8306d42fa12d2e8f7bd2fc43
zccfa0f68e15ca6f2244ffa9cf00c5bd383a139609923141dc139ca9c1e004edb6de8ed5ee60ef1
zac8e3c5bd89d91bf3588da0619174568b3651138ef47df0856a625b66ba43e281950ca4399b157
za2137f82cc9a31af2761333bdc24a45a969e0f7755b73739349a1684335a5eb408bec96a35ad1b
z0779bfbb035ea39c841b14b692850eb2805f5eb1775bee42066efda0331f28513fe17938a34378
z255784f52b29c6ca9c3c52108992c8c08d829f7eae428433c90deb12f38dac74fd66f9f386c651
z7a20382248f0f87c80e8ccf1923154e04d4a95bbdb543254f415dc5df9b5bcbe60e70da46eb01e
zce9e197c61fe335715631798678c03a57034acf4c9547382e35874565ba9a8f0ea37c22ea2d6db
z79f8ccc33a502d844cc21e3885851bb864aff16f0c763441272c51fd7128733ab3690ac75abf44
z58bf1fe0700c03e6db04062d957086bc3de582ae09544710ef95c6ad832f26ebadcd66a45581f1
z72b9c3bba9ea13d55dc402fb90310ff737e4fa93872c65864b7cc7ddd8e6530f7ea8e1cd239d35
z848f62f13e299aa2be60a0f7bce24da90b10be5166db05e6aa0d1703d46d5f82602ae9c4bf227b
z73fe3caa244a5d72e488bdcc47f4dde7651f0f046f029fe8430e0c192f69c5bad29583f37cad2d
ze6c4484b8b1bef77cf2e4b6329e2722d6a4a873bcd5ba9ebd8b063ef95eeecc593c7e5ea5b2a83
zd0a99ced3b170984dcb1bf98c97e285ecada496393a362f9e5f561a02935d843958d7436d247d9
zdd0dfd23e23926ccbf06f6e51996962f446187b025cd2781ab096bac2e6fb503a3c9ce1345d384
zc76741ba3968f80d0bc7cb18e6c2e0e0c08bc00d524cc1674d2f298a6c10b5f8174cbe8a50f1ca
z59eca1281c6f457ea5649b88c937554c8c24919f50c8443c468c570611b91e1ca3eea4f6f5c7fe
ze5a4288fec39eb3432cbc404eed0fb72f050f82e3256c07e4bcc88bdf08ad4e2667b5212ad816e
zf556462d3a927060aa8a1c366efdb902e9415ae62da25f33cc72484eda7373a2372ac477db559c
z1960235090ef2079938371f15e22efa315e607032ef96d2cd6904d05226609b68dfc3b4e0c5462
zd182cee7ca4a6ee657106316275dc6ff90bf807b8efb81ee64195e3cbfd65f457f38d96dbba4b8
z3c651b8191362f2ba98f6cd2c08cc31add4bc7ed690fbda27ec6212d98be77d6101f597f4eb2eb
z4adfb8970808a7be8b373a74e34020634b8a286808c0c895197e7c32ba0e19853ccecd734ce516
z575724dbc94bcde0817afd8301fcd8a03f22696d45ccb5d9f21154794b88dedd4b3e820a13c0f2
zba32368176e63d466314fb8f7a74b29d05252ed16cd4c6b825b4a88ec5f439e47627771bc1709e
z4ec7e651f987a7b95e763d15e2a8a6c39ed4cde094626f1644203480b0706dfa46bda40615622f
z6c5e392381a90566be63c359489864df819270f5d36f8d9fa09190fc373f891462315a68da94d7
zf755af9bd9d388fc342833fc8540ecd299747c5113f28672c3bcb98e5bca28e57f9eafb17039a3
z3bb9c6585295b159e464130721e604c58a53418888241ebe2636bee6c94dfa6b462708537e8203
ze54455c957770ba66d1b179ad5d8af6cff786ad82a42ad2375bd6512608295b0a4efc15a18aad5
z92c0606638154a285d4bb1ca96a5843465ddbc52a05f77240c9f5c7183188bcc1950e1f70cb7c0
zb0ac654c2019ea74000355f667b4f4792a129419ef653bff4fe55bfe8cffda281483581a462438
z019c6ee716c9bd58d517816a0c77fc84264a6f84252eec0ffa7b5fd9d6384b963fe10e28c57299
z5c4d626ec86fc3c311b74c5f67ae16062898887dc99d64550940d42d63f7225804c0be2d7495ae
z3bec889704a1ecc11a1857da47ea5264d849a1c41fda116ad1b9c35755f256fba23c49279f676b
z0821a8e38abe121ff39364706d4137815664ae231a6469bbb334e61ed3975f8855490a85bd0576
z02f3b106986203bb48e428b0448956289f40d68f4ee47318457343490a1eceea8080424caf44a4
zb9c7bc2f0ebcde663934457da0df69a0f6805ab44f6e3fc5725ff0b1668c3dc8215ee6ba8c16fa
zc77d850ceff337a6b9ddd7a9adf5bbca49776509a9a8dcbc64728915fead3147e3d6ab4c5e7cdd
ze58a2ade158af91ab7446dfc79fe591927746290391dde072422d736648c4068572fb32baac6aa
zd3600032c6ce7e10408e9457a3ed5ce85ca99070355f9b3a3f1d04a1e48910a33d3e53d67b6397
z8a8ec8e0bcd256b6de4aac229414274a79aec172dd1836b87177bf75659811b1baae1e51e08b00
zf8a3fede9b7ab4305985e2e2d1ab67dd5582a0ff8c73ecf5162096a869f3e157c32fb00e55b14b
z6d57df5ce8557eb69298e8172efd3457fb10185b79a5b9f4f194af14fc7b4e5bb8f9ed4ebf878f
z9bc0fa030d8e170ece8991d05b115e0a82271e76101f3a32b722b90e70dd66d3f0ee1bfa63d61b
z463f933dadd47feabbf989717643c52f69478ac7aa182a526c76f77fe5473a40bad3a2151f6298
zf88f6adaf7e3ff4afefa923c794cb288cccc1897025afad064bb52cdaad39344bc864b6f0079eb
za14177bc069c97f39c7592a89ffaffd3100a4368bb9a284a4287c2e977668fdbad2cd285b7d856
zdb683676db25f03e96d4f8b0ce78c5a16676728829bcab64029478e91f49ed9b61da31d819e165
zd486c2910ab02da0fb11375be750c3248f2547e53217ffbb33cb9502414dbb00e783e569b3c671
ze173cf650bcb4f71f343afce4754ab77331c8b2683a219e3f719d6b2fe400c928e65812dc7e25d
z0f76b5de762ba36a57b2e4fe87b010986b3d2184f6d0677e221197339a0af6cdaecee70325d2d3
z71cbc4f7c17b556f78e847967537f9860d5c267ec0cb298bf4f76ae465adc69d431c65e546daa6
z1965c3d3511dfe434141b9095facbee50c49cb4cbdc6a0b63e011ecd1e40cb4f4ef36a891bea2f
z0115ab3a7dd268225e458b1ded6cd0aae45f073cf373ed157063757055c6b38d27502ad9ea9d80
zf15d02f4dd7594f9fd685abd035f22edd6392ac4761130f70f5a885bc2b89d21456d53693bb4da
zdcd4bded159c727df5573bb31c8e6bc6666ecc9ba170fec7b64e0d5d82bc9b46c4f2872a89a20c
zc1350b9a3e1a60d5928688d34bf3113555417a46e6e11c0175802aa508f15d0ffd07a76003ddb1
z9c78041e051b1a0d5d0c33c75477dfcf1b3a3bd55aabf1f6d1ad92a05b7feb59704c9930decd96
z5b5918eeeb72023ee259f7531d41bf66b874e59e595ae91a423743841b48cf41b8ef2d07e3334f
z031c326de19b3a863b9b7e9d16588de1ca8ecb9c31accaafeb2ef00ded797bfed760e367bc2085
zadd565bdd893c871afc839e23fdea9ddb72387dbe1d1fe88937de65ec95569a8a892c94011219d
z05a0f59df59bc5d57001c53a8c2944dc1c09896e6c62478a23d1a3b9237bbea97e7bcff742aa09
z3908917db52a507d559b090c1d8580fd399d96a86b6d30249571077bad8318af85b9a2528452f2
z7858d85fbfd8981a1936925d3101340c74b994818faee3f5596a76d22a028d45626c90da3bfb26
z0938b97554da2716b503554d9aa87ee7e589cbdfcdf102064cb933fbec862d9a050268ca2d5d17
z8da5fb9adb44d5e1fbf98da188e1a7fd26dc643d6319a3c8c4a2473eab09189491411577dac16f
z8adaba7cd99a14cf0e34aa7da75375e4ac65c263e54737d2864380f685a736461e4105a71b6ca8
za1dad46b1ddd2e908d21b6c2f61302b07441892589e7dca6b2621a46d0637ed7713cdffe228f2b
zd856917f4a419b2a399589e6349608e38965caf0ee8c2c07706f85b5504a181aa30b4dfdf06ba8
za3ffca706dd0437a50f561bafdfad26fce0d40950067d0d34bc93c13e4a2fc41889292041dd156
z935bace0bb0c0cc16034856f6d6cb004194f9177b063756b9e00d2fdd43e7b246c6bf34bb680a9
zb97017846597db0eff6852e0adf44f4bf001651c5a12e7840777b32b688787eefeb3d4d7f007cd
zb44a70bcf1d59a1e859fb3a5a4ee34aa1745eec5ff1879e467ab50cba5b451472338a4b60a2375
zf6e65651aa2b0c556a9dbe84fa9ab814475065bc68f8f122db9237ff51995e80a97b283dc64287
z4651699b133fe908d7c75dd44b08e65a1c5a04ddfdc28c2c10ff417891938816ef724235877937
z448dc17d984874ad070382a7d17c42a9c06c577448cdbdfd94c05b4e4d0256f5b6577bd129f929
z525aa7a1a6b35c52fb0418cc5bb44e79f3e23183dd3a0a4506fe2f9c16f8e887d23cea3d2cb482
zaf1b9d060155b29bed008f218e7d0ae3017d3aaa6dbbc7627ce96022421c8bd55be00eef880ce0
z331d6389eebeb24cff05134c8eebada4530a51719e1c3f18106400fd11cdeb8d4737cfe482e96f
z3c4570f6c6cfa61984c8eca8780bed2bfad86544832e867db88c1c15d2078233526470fb4f0edc
ze322be3df79bf9b98376c779bb5f8525b9dd48ca68875adcd1c3cf466b4f1a4ed1c00d5d925eac
ze4b3d53454b507fe6b80bbfd20d3ea444b1df821f2c2cb5f865a5b2e94dd6be160f9f6eb29d8e5
z84caa7945b3f0a742fb07915e55b2e375d6372454f4f220c8e23d8d1d4b04ffb801b50690bf8d1
z0ec27b1abd4a4cdef6043923512a797ee114af785a5c5aa04ddc1e88c0a7620ac34a3737c3f472
z8ac3da117605794892de0dc04cf82b0b33d7baed5afb6a47a44b3b358e090d7718ace6ed695fb8
z4d863ca77c8acd53998c3e660d54ea0991b8b8fd3a1042d7de75df7fcf106c4d6165c6a955b67e
zfb49efa9cbe674d2cd7d2d9c0ab565ae08022cb39b29cc2321ba8500eef791f4fc79f392f0ff03
z3e01b0c94c6c4a882f7d1bc58520f7076a015093fa7a970b0cc0e12be3738f0eda1a2d0f433154
z86c6bd1b04a93a5e39151d295c658d5ff0f1afb3611551098e0c1b2adedc1396e144d2daf0dccd
z2d9f688676997df88f73b87eed68563112f5e6ed15e807f6a2caf270d3ddbf5e5c22e2c25c0e60
z38faf2cd0f32c62c4b6cb9ef025680ee0e3c65b37d3da7d86b5dd043419d517e5277dd03ba5d45
zadf5ca16b825efbae15f63de181d1bc681d70536334d1f76c76d1331904b7bcabe02f84ae53789
z6c059c6b36957bbaf8cbbb641fefb860c073588784fa391495ee380667b163926fea63f0c0432e
zc875579c3391589a9e6bbc1aa098614bfc67a5e1ba1460ed0cc62dff1df8bcaaf05e522cc450bc
z64b583ba077770e1e1c850f5baaf47bdda9e0ecd2dcc4f69a316abec6a413b54a3c6a5cc84bf52
zbae083a28ee7d18f1092c0a948639c537fb2eafad72b488ff8f2845bc20fdcfd647397a368f6bd
z3c11f1b8cfa743891ee9e7d8268c90fc72ee721f88220ae54ffd83acf127286010bd6ebff0cea6
z3bf8c1203ef521ecdbad8ab509b3ef19c891d952b7bbdbedcfeb06720b67157219539b103d291f
z8bb489007a9169a5acc81ca7c1a74cc56ee4df034db34ea24c3822cb1879ba0f513a39e970034a
z1e5bf32b32589f2b9e98f542d0789fc3df5e66194fbf34925d2c08906c4063cfee18a1c1684a64
za81191d0c02aeb24519303a3f38b4557dac9aeb93c09bce0d8f752ab42787362fa6c0946e4b857
z9f7e7491a1e7f119ed10cc6fa36aed1d59031fd063e8955d912980e9465259ada8c5b4d5452d05
zc6aacefee7893e8c5f4cd8360f650b5c1a7c02aea822abb9397aa2617fab366c7c21c155bf1b6c
za0cd1951faf1e27da56bc1c79e1305cb6c78f0cc385c3e758a333ab64a2d8d05a6404ca8ccaca0
zf1a2ebe23fdb03c44e45486d9ed5060ee2bc5a5c6e4a76613022c8e4991a84a69b2dc5922e17f3
z35d6f11558b1739b4fd5c6b4672616936e2ed12ed67d4e8a178aa4db6520cfd97dce52e63500e6
zf5d25dfe018b37e818f2f3e3f5dc466fe5b254dd82bb3b15d3a03d0746bd68292e291ed2f52935
zbd32a86ac1ad4c69f925046d753e392c75e7c3ca421aa2455adc9560338967e6bef7f2fc1da5f6
z426c24a24d251f5253262d1dbaec861071832805347c08788f001549cc2c34964c1f8e5c6ca549
z41300604bed3e498f5ae7db0f80569ffd7684e65f6c690e530a49271328663078d92bb503eefaa
zd835fbfa0fdb8f2c2ccab872199b4bfe34a753ac8eabf46a629490fef1f865eb66acddf1bb8a31
zeef489e239b6b7027c737dd40bc03ae1a636ec59600f4b6af6e1414876ef737b0253e5c7d8f060
zdd16f510bb31290c94eb7dbf4b57e806324996e6967f2d0930da92a0108c094c7aa1f2b60fb8ea
z3ef6d530fb1e90cfded923cc04a7d2fb102a193086e2ed2a4f72923c31021876e263d70d647c12
z01d789b5410741938594732c5c438fac2aaa79323a4db4fb594f31dbae88ee4ded2bc398b44c06
z1e266ed99fb939693654ec8b74349792233ad6bedce155b3708f87d110c7548b0b855038c430c9
z1b661fd207542e628eec5f30fbdcf3eb205771889aee6909a1eba6a1a9c0b6eed087db678a7365
zf8e8043498605d30a8c10032c593d69f4287f80a647c67d7f572e898ae19559230d4f7320510c8
z06f426c5ab6c13da83874857dfca16ac72120395e3fb9d18ae7c7cf09b14877c296dd09141684f
z89166eabd0bb48c21b4b7d662dea2d27bd2245be963f6854a3b80f92e5ab72ca2df7b9cdbb4267
z8a2907a1a3218d9373e7fa36f60f7dd69842bbee811970295f3cd45960221476a8071b2c9bb8af
z2528b5fc32e6725560d47b659a499ca2a58e1dbb04ec98f583befb42d207bc35c957e74ac61c35
z1cad9d967c537274538cc86799dbb59bb8c39116a8c0afc2481554455c77ac0d163ef9d845adf3
z107d16ce13427566d772d9b0d961726f83979c4863bae6e8e143dd0bec31d1b7ce345c96598c64
z9bf4efeacd848a6b2b62571ece5b875b2f5a36cdee14ee4b432c5abe6ee0a9e4d2af66064a9bc7
z4a726180a3ef2353db0e23ecbfcc842392c22aacdb6fb437db753c76525dfbc185e3b4c9a2d208
z136e31ede015309006eea5d42a50388c77397011215d6a3eb6c82b016692fe4e3bd3abe53407a2
z12740c8cddfe6e270889088d4561ed12e953fd7a467a5a79e1ad7eb0b4d94515392e27186d8751
zbba4de32a3550eb66899b5e636edbcfe6ce3eb61351393df9f2b7df043d32c2aa568850320a148
zf267f4a6e93aa6abc003cd6a65cdafd46f183c94b7e8c689fe39a2b00436c1d3a26285f8ac4342
z810288c9708f75dd8d838d59ac6a938f8bac4ab9429efffe01b67f5cd252b03ff43c5e156fd99a
za24037c71de3256b6c426c69509d483ce6ca0a43f139ca20add6ea867a7750e32fec20a5f3c1e1
z885cdac32c900a483e45c4fc66eeeca7746a578d0ff69a35de6aeafc3fab1cb6838cbfb66637bf
zed8c5d475ca06f42dd3dd9f4c5e8050c2f1ecdc3ce6e6f81bdb690be487652ab58ef7771208f69
zb68973e9e2c61037d09a929f2a750ba892e9108cb5db50c6b902fbaa124edae9abfa95c9e06a6c
z5378898067201cd3a8896253993ff27d66a5f2e3ec50c3319625d478a797dac4ad226fc2119042
z7f01a111cd9a2bdc8db239810f368c081986b93db5fa2e967fc2592a1cbdfdd42eb8c72b89dc00
z985a2ba46fcaa2f63943cc32e4c8d85cf9747ba44cf7f813bca38afa9a3a803de3eb19945cc259
zb77cad786a123a41cdef649749cd983449473cb016e0ee799b6b218b00fa261e1db385f5e83931
z57967fc1f5ec8bc09d0c08bb557f1da85341e778abb18eedb838b0beedb00ce8aae54b40be547b
z2b6694471e87e90c0c1f08ef3e3a6a12f3c8a944d019ef9cf8fcf000f5a1db247abb23af226247
za8679f09ea818e2c736197457544aec26046a30880c05bcefcabe5bd979b1c3ea6285a2b12dba7
z0f4d2e74cc0ff4ccedaa033aeff02781e9e8e792543e6bde10b3e10e59aa136e35b43951ac17c5
z2b9adc84b76631be3a6d112f8a7e9b03593f3b14a6773367346c92c23191dc44272ed322bdf533
z7be642ad353e09b130f80bd72bd59dd067e841ee4c965d877bca73edb2201b5d0faee71ddeb78a
z6bc0e39bb9804ef6eb4f111b18f7a11304ee5fc31fbbf99d8d83ce3ef490b03da4e4d1d9fdeb79
zb8c180613f804c3c54d24ed063533faaa90824c6e1f043afe149deb7fab13e6e8419945e5269c9
zd20277b4b2994c17b5c9212fe0cd73b0d8835b49f27a7436aafa63e12fb4e59fc3a63c52fd1ab7
z71b7a765998cbdc91856472fec3c2f28c320ebe0b8cc13f46273e0e0c3f25d9ab8cf4ec2db0ff3
z94561a8bd9a22a081fdb74537baa465a806d3f466ee697c47d27149b8bfc92370b904ad79b4a9f
z658b12ad739c7411581e7040d59367ebbf8f6850a92e0167689f3c23cc6aebf07a8fefe1a6b143
z2e51b62c5eaba66357310dbf46f4baa2db113e01264a1818cd4047b08659eb9de6698acd5636b9
zf8c04d486c609c2cf9b25f00bc99feabeb9fed5a16aa32e0fc1c6b9f82d638ff6a2000d5cb96f8
z1e47fd08d0fb2ae4b16f494ed9ff1a291b2aa662f684db82f14e5371085ca81bf9ff5d9c21d9b1
zc9fba22c4c1b44510d8e583544771b2e954b893b0c74dca5c919624a8620cbe4fcbea3fea0e051
z048a0d6b809a7c1ac436254e9bc011df516d8b753334ec4fdc99e8427cff6b5ed4f77f5dddc819
za8bb0dbf1e2edd98cc641b25c7e205c472cb66f59ffe72e458b765b19f125b5f5a1afdc8068369
z599ed549d0521f2e747f36894321ec5c76cf6a8bf6445af9d3d3f1287806b3b9e13d096f6b8bd1
z9c3ea3b0ba760e18ace81e8214b0b75daa5a803e6b835d3cfd9131c173fc48c0d5771dbb0567d1
z86bd8fdd2e3657b3a3606188596f4fa3bde9fbb299b972ba790f51c613ccd4e2321ceb279deddf
zf1fab450e406682aa661acb748126ee7ed7a588d02318cf0df694a577e5b1c0434b80d540a27c7
z3c2a6373d6b4e34216752ca6209aebcefe18fc162cc550bd7d8c6abd5b589c629fafdc1c7aa843
zd6d60faa3d15287d7fd99aac3651c736efdda3fff2e9b24adfbed1ec74f3069181f85a7d13fbdb
ze7c6d5e034666b9616f4929d8d8ffb62c2fe59eb1a61b5f64a31bde031abbb126d9dda1c786bb3
z2ae7766637271b49090883a61c43c4e507ef7a46ae7c391f5e503fb950ce437d0373292ce98bbd
zd2c964aa82eaf4cefedb36d5ea5b155983dbb4b3d6d7be0f891b8b57e3f95a0dc021d6e3bcd441
z01200953b62737ceae5c5deb06d357f224540ad6f3ae20b5e02999756b64afb5d93285217859e3
z474a32c03835094b33c4b8a98232429c31fbd2afeac38cab636bdaf524969dd273f281dcd49119
z469eb2bfedb781ec458883d196fe4c80281b14704f699e46d371f794f65b8271c0b05193b9c6a3
z7c2e305114bdfed7169dc64f95e371a12f7dc608cedc7f7e816ec60fdd136cb30187e16de9609f
z5f8d14b2b6b7029f82e1b3750d302edd293e6e67e383b9bf1586d49c8f6518bf6f4229185d8358
zdf5d44a0d156aae43d3ca487b460c8e205a99ecd194b223a21551980459528dcf056cd172f8448
zb1fbe2f84fadaddcbfb476482149c644e176c36256b52b8724d5dd074c42a73b96cb1b746d2bf0
z10fe4393e1e8276a56b8b32b211877885ebdd3c782d9f369f0c87804f26c5d766991ff9f8768a8
zcd4c231e8279f30971e2e9df8d941422637f91aa9b60d265710ec5be3b88f861e260ad9971d7a5
zb71212a4f877c53ebb4dbca82b0535c9049a91e3d8b70efc558025dc713dab14bec7204f3c070e
zf7f830af4229487f3a769adc1106ed03cfb0f00357e5eb189d423ef65ed39efb17081e49df9c8e
z2f562f26a75383d3c934d6c0d80a09aad3102bf4bb5a6c2a147e1677207054ab3df390abc94526
z74d9ba56a790ed3ffb04f23732e9a4c90f0c189a715d192a0ccd23b1d7fccc02a55eb5b19a698e
zbfa36327a979c7fb1781b46afaa7c1c34d32fdabb1064f1fb95c877d0b1d5938f106c9b8177bb0
zbd1bb67b83d511ab7406ca8680865d48ea642b1d2704ffcf68b8ab45f7988a16b3fd62cbd79677
zf188e1de08709c4b466b2064d5abe2575c83ff74f0001bbd7677b8911736ddaf7b03bf136c5b30
za060b4fac91768705c6d9b16499be8e1feb3b8716493bdd2ba610d3ef36125b16f5ffb548b87c2
zde1515f558229aca98e67e17b1b0551656e9ff724b8a9c4ee851e332d8b0a8fa70fab892b2eeed
z76960d52bf9b244452150311111475f05cf7d2aa258740dc98b31f86101bf7b695c10af9e16b6a
ze0c03f4603dc65a76f95e3b60ef770be0c4b5976629899f5c154bcb3238ea3f39c66e27231ae52
zac348172a99b4b963e69b22321ee51f374adac7d59c4259c1731401e7142396f2155f477d7e49d
z8293e5fd19d8aa5a01e387d76b9f14f74b6eea6eedd2f7f938d5653814c4c1f1111c33e600f3c5
z2b71e91bec457c8b8ac6b18ee3d30b81bf99afc6d558dfe3a503441001a2a2035b139a8b7280e8
z54a99a5427ff17dccc17720b39009446dba1f4b1e7b5a7b1aa02d696dd6656de7c87ecfa17389d
z4290c1e5f66997d8f9bf2ceba01b84e88fd02c3b6aa4b32b7cfc75ea85a509b59116f24114b3b9
ze45015eba17bdb971541eeced6ea301152f9996d89f8e7b524549897a278861feb2d90f3d49905
zfbee43a88a20e900ddc7aaa581b39407ea3248edd357c90d16ca914d3b824e209e4ed952f6543a
z455eb3c5221ef22870d4a79acbb18b42e19b03505746fc004c9f0e61b590071d6942fc6934b567
z7dae756ab7829685a306f4a67fb9966fd9e91f4dc432ee529cef05cec4711f5965c1f801ed6e39
z1069c2203df8af3e0ccd8ce37eb9d69991155d74029ca3c261c93076c39d6c66416358ec2d7b86
zc292d387eba7f55b8b23a5907519d4b74e2cbbdf58901c4abf732b228646ca4415b1c6ed4ff7c6
zdebfa07a217266685231eb9887f67063820cea3bc8142f535e23f11b1dca20a9fa696f5cc0e688
z0015dd66b93933be3ba0b66ed488064783341dd3bd759300d55d76cb8af50f967800298f76ca97
z202393ece6a800f979eb5ee3846b6df137514620713ab4a9a57f86170fe2a4c97298bd34e64d3b
z61a20eec2550a97d522429c6074728d68b53a1d008ca74134ba3f14f77441f024a3e66f664c40a
zefe3a4fe10dfba812db45954b7be6025045223b1a13c578c9217050d0ad1ef82eefc8007a7c229
zd9d2db80ed24417065e054a64ecffd893242c9cb377d7ec81aef5b9dda08261705d96055536ef4
zd192804c530e03b98dea142e76f74cd8ba977a1c8f820be093de6ac0549583d177b712ffd43c17
z8c4177d885d0a397fd9f1e2de7244b5f2b2f169a7dcd25681647c1c840893187016c9837ad3647
zae3d32dbbdade9b7d686b11b5b85aed57db3c628856333429c5d0d42cc082eaee1ddd115615bc0
za809942be6a1bd7689a234ae6f8fee765665197fdd0790f4720691aade485a1fc5d39da03ed065
z6c3f22e8457c6c496ed00f0747f486fd3e7ff1a9177a3ec37d8c082ab825c769fb8f07602524bf
z58d363ff69608b623bb720c4c24ed582acb99662d14b6d9f810f5f4f5717b0e3cb90b964baf1ca
z20c2d08a239c96caf8f085236c0c379bb1089f3bd46c0f5eaebbffcbfb3df93b4db8adcd2c19eb
zdaf878ce4444d17153076599921016255e3740e9cb0f0b1a4a2341fad0ffe2885bba527012a48c
zcd6765494d4b240ceb8e4be47a72b9715da015516f373249ce29796a88cbeedf379435d9c4d932
zd170474eaf9a8a7474339b6b9f618dceeaadbd5d8857e803f276f06df70623ee6090198edc4c09
z245e0c3e5c4d73034d12539f2d5f4dd61af62c8b40f301a1430e7b38a98fa3e6961b0595608b40
z25ceb80adeec947eb61d5f4cf93aa1fc4659f67a07f16fcb1aaa74a351ece5b4dc2dea8ce81141
z8e8118212c52ae89279b4dc5c76821a212312c591e784092cd33206aeb3d3ea0bca661b6cc5af6
ze9125278ff5da259650868f370e061e68e0dbd9c993ca351ae29e230af1a240db2daaeeddbebb0
zb596e41f78854581057e20fa9d071fefa9cdf502089cdd9450b2e25e83d71ec3932c6a35c630b0
zb0b1a01caa7ac13d0d46aaff5a4da3c34ae33f255aab4263d763d1a9ab86eec5d306f368a5946b
z8d6eafcf6c932bef9e7d69f4914cb3bcd11ff8395ac2bdc82d37796a9b0958149e62b0417cee6f
z69354a356b6cc4d9416721bea7cf3c5bf7129609fb59232c9200358e8e4fd71183e933f1a0a4b8
z3cfd191500894dd2af4f1382e5b846e83d24563100befda025473ca21f0c7a07997a7d1e35023f
z7a07c7bd413bf9e0588445d3d86083296e9574df3fb6a8404ce299b8ed09033dc000c3524b3980
z366354f31172c65e64d5d78c11b8974017c62187c06d3bfbef1a868781450b43a5360cc34fee85
z41b1ca8aa48fb8ee767e2add617b0f357c0609830a9e8ebf42f12b7cdd77b3638135e14435b74f
za23a3d95646a17d98cf4817d94a7ea23a48dbaa64ad6f7378b58d30e64b4990c6a4db60a8529a2
z3af38a7fcb071c8e03ddbf8001153a5995e93560618b8b44c1c911041fd1c1a494ed719652c13b
z6bd7ee8f98191df1c387119be5dff9fc97e992d56f0ac3ba7d0f715df90d4060420ee009669a8e
z6ae547db87a1c1d8e3807a094a7681a491e143ec6e289c1db4560435db0db9ec6bcf1058b515ea
z3dd5f596faffa3c6a72e10a3e77d99415ecfdec519ba2463cb5484f9333f524bce40e8f7b2db76
z5671cd7d9dc8c08fc49192e2d504be62d422f2e92119ebd296315008c9852753d62b44bb479d9a
za17a522aa001002e9d2069c67994159ca8d2c08ca760ab3007eafbb81584d4c63f444290b172ba
zc0cd1bc1a316468728cf48cbf7acaae8c04a38f886de3e3be5d7d25f0f713ce9cbe3b83e9c8261
z05b6392c974db237d8466026a9ae89f9c2c2ccd9660a65590cab38920ed0736a8778a28641c0fe
z3a56c985b8aa18fedb03f515e31e9a5cfbcbf6314e9994d97f90e504096351cd81c922de5468ff
zac47d78131ab0bafeaaa2600d49d67f1d1e7e581b58d9f8f070b6d04f078563589e122b5ccbbc6
z5b1896ae076912abdfc83ceb73718824ed9cf6ecb5ca9ac4799a0ad5814339a9e901ac523a0ae7
za40202405caf2530ba1f0117655914b0ce3c9bb070f0d7793cf419e2ecabc5b9000777e92cf902
z9d7d841ecee6c77a39bd3a18a0674156ea398ff7d8e0ce01d41f63c6ec8f3d004f6e4da417c56a
z73151282607e9afb8d26417fa9d79c9fbd4a60b3db5e9dd1b43cb18642d37f181b427715d03ffb
z5b4bb7f3254838f63e7244ba550730ecc4fef40476e70268e71a3e41f20a8e65d58271f1cf3ac1
zdad8eb794b15a33cfd5437afeb6b08e6d59fa6dd48db42d5fa48e27e55aa5aab2409febf8032c0
z9a68d31304e75e99ba7691b48cd2346a0eeedcfe25d9952592b6f902bbce8f18b0a456596d25ae
z382188aeb80e7b71fb85cec4f67f7d0deecab3faa5a52427029db6e8a3b7c30dcc98fbda753b67
z2d90d84304807acec72767eb2f502f3aab2a609bc154865d34cd754f3071f539564d862c69cd78
z102ca0b4d6f30b0b84df2c73d3cdf1381a4e25a7698e15a64416299d84a81dac2a8b9a493b1b4c
zf71d0d39966ee9ec25edecea0613c805922377cb955c204e946df94bc7e2e95a24e77ba982b195
z90676a26a9e5beab49ced8f2aa034cc4e8075c21d347810e93ca4348cb47db5dd87910c08c692a
zbb9fdd03257c085d46d333eeedc5d27dcbf91b46937277cf05f51ec54737b9f4779164cf4ecacb
za7c4067d8b23e5f8c365acf7cd5db6e230b31de44cc312a55119695042b7604a2f05fd82c872ae
z294638392f7dcf398ff949898aec3306b50577200e96ebca6d3aa17355a2387070e3a166853542
z16c5add1fb862898e04bed5ddfe4b2cc33e9dec4c63e68bce6de5a75ceb9c55970c42261f1be3f
zcc75466ddc6f234c27e7ae8b783b2d3c1b5b7058abdc2f8cc82fe9dc2468d0d46378e2840a0f19
zb311da57ca36476c6f9c2825401e34994deb90dce0076cb4b387d728c0a480faacf280620d6219
zb2bafe0eb84c80cc43a12f4740878bd2d77a8facbe6193bf36c2781db177e0ecd2e188722e1a0c
z6dff56631785f002d32e8b3b497e2ad3f006c8a925ae9417c6d689717861a480080fc05f12ed40
z7981b49dd819ccfb871e939d919e64b0e305193850f88b4884c4e449d0694a13537fbb1454a089
z74e40070b0e57d89b460c2753a7ebeaa6d614372cb08b4f2806e0b7ded243a085efdc9f52da4ac
z42d195d01cc5293a07a80417934b29bd9facc68503653dbddfb3ee19b4439ce5455d28a817ca63
ze26096b5b1a68ef9b8ed056768d4610638d27339fc3de5a60c2973a0470c5aba284c6ecd2b28e5
z9d3a56cea12931561bc5cbc4b9b4953adfc9aee660654825d20e7efa630880cd98e9e79d6721df
z7f297d07d436d06ab1a1d64af589c39367fc7201d9d810c6b0106cb25bfa385d57356c2bfcdcba
z2ed3095a1399a19f0c90b69b31f2bed4c751b41d4883ea9bdb4b4eca93efbe33675388d4d8b1ca
ze61006b0753057711315b650bae9354619559a8653bf8f5f7a8c21e224dce1af518f5a856fd42b
zb1254aec465c79119d14c4bf976a95f59fef70aea35cfecd967857bf4ded1a9b2c3a027334010d
zd3ec4422dbc150c1a2ef3e78cf23e8d95d445797def3c6b8442bbe6c45820834d54df99a3d6f10
zee0dee5f54d9c1f8c0c3b76c332fb49121f94199b064131a1d7f5fbea02d0fb337e7aff4bcbc89
z8d45dc837c1b293224d1e5073fda8cacd4f5be593602952bbbee2ed5f57d2c48ec3909f15eb5f4
zb6d4c3ee8ce58a39b8a801e1c55ea36e62158c41e9671406f9a5ae98bc47a4449b55cce21ed0c1
z9312ea18c4ad175a8e7b7a0708f60e18205cf80fc79aee54bc5d1053d8a6dfe72a88e37e0a45bf
zbb897db2029cc9a365a6fe9a1a44e98a87ceb9f0e7e4e2fe6c9ec596576af94aed9eb4bd3fdc7f
zd9765259c553b44dadfc2968a9a6388263eb33fb510323f13851a9d86b77ed102dca5c4cb0dffb
z35302516468670986e3c338a3e4d9064025d7febe889280955c927d287ac3aa5f995da4e561526
zf321ad84420ba106bbd41b5c900a0d764af8e772d7af029b2935e2391edd2b771621a139cc6f93
z66f06e818fd1ac565f058968e91e599c272a754b5b8f1857a9e2ba97aebb507b6e4bb081aa51fa
zd797cfb5641f0d7c64d17d221ba1b802235294a478967cc60570fc2a6dfcf2bf77da6d1516272f
z63f063205641c8b1ae9c1988723b5991fe575ebecc61b7a951eb7ba73d1e874abb80b1a44e0fd4
z65f952275644e7c4615584f66cd8113619806bf8364616ca46f63a3237d84ff973aa5b4bf3fc14
ze09aaa96eaf59820113156d8f643adb0c6609b9aa5634601e162ba84059a2817e3a9efc1ba1815
zfbad0a8718a72ca82b161962c9aea00c57c0872fe6de30dfae32931ba85187ce7890b938834696
za32476fec8c6eff7b73126d5c37d35ec53118ebc866020031ae0937963869267695ff604661be1
z4a92db559d7645494f851e374e5279fda6cb06fd68924ad78542fad37273c665e3010d74bccebb
z7b75fe3bc50cf328735e579f9b235b89aac6a240ebe7eaabc4746c2f2632dbdc4f28855bdb3c20
z00a983a14ced0d13ff8c44210f75d0bc44fa1413314292ea8821f80c045892f0c36a5ca3743397
z535c6f4643ca8d02bbd6420c73324724f9fc5ddf75ac4ee39642908f56171c757bb874fad0856e
z5eee5d4e18361569b4bc7fd59e86bee2e564d9db9293c54fb3db0cc5174f0ce2963ae4b2f3833e
z677b24798a9cdd06b7c34beaf2c52a4b7af375615866660193815abce3244f4091d36203eaa397
z7581e319386125b67d59bbe91057483108f4726a3bb4c1a902a78c7800380a99c889b5013721e4
z072d0e06c582ab98a099270f8def1b02ff2b2456794522792d3581a90d420cde2dd25c87c18413
z2495f79358b01b6f12038103a08bff95587d63ee7a2e17e6c9acdba712ffca04d1418a571d28e6
z3331b43be63d31dcb6fc3863bd3ddcaaec21c17f5bfda57497d01958cbe6cc05a4b54824c1176e
z0c959e1f5da86c272574ac05597e5408f635b64a6e58e34db1587ee4110e7c9e83ee17e6d5963e
z5918828818922d8cc7f44beafd892aae6a17f0e834c4101352152f305f6a287338ea2dca057484
ze8d6ba5460bc77eec9d8bf9da6b4b3398e9e2654c2923d5d27dffda0035ea7fcfdd4a9b6eb7603
zfedf12a81637ae5bc02571f6314f2a45105828f679a9cfcd7663a5f21139b23020427b8ec36fbd
z7f475243691208cba12bc1f9c81b80c487466632696b0a3c03749001fe8ad342c2e6dcbbb4f90f
z73ebf2d53e681697e847e55ff242153a7618867a2c9bbfe06259cf363e36bf8eba3868f43ada58
zcf4288f25167304f142cc6c5764f128b0faa33413c8e3cd5c8c8064708705e495743cf37b857b4
zb4935b171805ab9b7786ceac622c17470cadbf271ed491d112013b81344874d83d7401c398da51
z55adbd19e3b146019e3e1bf04ced8ee594b38df32ed9b3a4ee697b873417e59c3a29c8d4a23bf5
z1ed9c42e187ba4454ce91f9be8e2b4789a8c34a20a8a81d237e685a6b1a65fc33ef62458b71518
zf6db5705cd8e3d0b164ce30abad5d8e3ea17d0202777f61bcfaddac1a6f9df405dc9f88c71534f
z3230d201c3f223f2364546ce620978c1a466521af6654425da6b53f843fdba17d0fbadcebdbc42
z481cf1befa4bfe97c0b1c62d14a330447659759b402230c4c22ed801076b1c5c01c6c4a9149ae3
za2eba71c088780e99b144365ebd0f837f03342160c0bf87ec9f7938abd28e02c9e09a06d21841a
z0c7724ae8611be791488b6841415dc4e8320d52e31498989d403bd7a036f2edc3c6b124ce697a1
zb86762fd2612ab20eaccfa767328e8d7238048f686673d8a03bce77f46cc4a4064c2e00b755e56
zfc9e1be05af41a13f685465f532e8c9f77d289fcf68fe4bbe289a303e7d8091b54f0923d36b159
z98d76a77d736ebf36b4b9bf6d7973838a312b3ea8f6d21e353153fee78ac2808b6d993d2e72d6d
z9354d14edaacb3c902b49ec57c8733bfb3d26eae734157e8314c48a26f0038dda7d2bfe9a0fc2d
z5b164ceb82279dd24dd8af436289d20043a9239e43d7784bfd6ff699eadec2e0d215170d7b05a4
z2e31077166284bd0aebcd99c51d5658cc2eae0b03c1f82de873954dec435ac7c515991710bda44
z3e9d0176f82c545ffaaf194e3863584e88f0e9280f08a6f26543af78abda7869cdd37a928cea1c
z8d6dc02793fbafa6a0ec12d995873ad0bdf1c92daa06197c882dc913cfb6c669bddca7f27d30c9
zabcc7ee09b29f1820a92d5b57857c982d83f7707aa6fedd4c7ab472ed718290ae0c8a7a130b7c8
z5d6cbc03f9ab719fd99e25d1afe6ba5b632495034b0388556cef46d67736628625ac279dc5523e
zd728351600b4a881965651bab43942d196f4918a4c8335359fec56b078b49eea0bda226d465e7e
z21b69b6f507e06e27a4cb1ee6bd72d330e3d49fc93acc821986a6c5b0faea0332cef44b8b8d2f5
z4d217e442625a18085bd245cb039ea629c19c891a87643cd59c8212712c5b384d5ed19161c2894
ze1d7bd6d486925f675b06e397263d983a2d9f980763141485a889012afb58bd84d5b1c906c6d09
z4fc5209a4025f7aee11581c54d39e9d3cf091c3d9dc99d4647cd96c80d87bf975c0ae2c2e0f385
zd5f62735077c0923083a212374da87f729f50d88200bba114ed6d78fee841769e7e64ec50fa239
z21280f11ac33a9e5d84bbaf7891feef29e25e00b52371b6124ca2144292d516d591df57abf84c1
z174b01d9c472b23acb3090350755f730fa6a8621fb2a966f83f34ca16c353b9b75b2a3cc2c0f71
zf2a92fa487183409e964d94055d99bf3a2eb7f21c67cde633626abcd48e6ffac29c9c3f3eaed06
z28b699f540a5b6bbbc3e881b09c414a6ecf4856d65e7a72c801474823a6a8482f7135252622596
z89a00d819559f7c9e59708279cd360ca0e003cb0dde9fbdbb8980e653dc83b02f841337e89ec93
zee68f94d1793ecce4fb02fb7bacb4dedfdefcd4742a7a0781821669cf8bc41dc94a792b99e32af
zc7e3deeb11f3e6426d1245f60a64e282cc43c69bf7e71bd2e1e22978df6ed21b1b6afa56c3ee5c
z57cbd35052e9d49a6082857f4793a503b421738e51eb680eb5830a9b450a98c7ffdd7f16a783aa
zb06033060479580adccf60138f1b6d388baf9221e42290e22a55a3a5a21e3b76f81d77dfb062e1
zf8bb98e7919c1acb328e47ba4b5a4ef0aa31c7d709ee24ddcd3a10fc32bb22e8d470aa40e91878
zb5b4245eaa909282e1a931d8dc5512f2d1f0bd46cfe9a1494e4b2935f553dfbdbd8fa30508db4f
z6c7d52c5c858328b02c93d8368db0ea20d8636dafcc996e41e9165b53fbf2751d5f68b9d5d284c
z9865227a8cbac6e0c4066b330a9b130f1b7cf1a9cdc4802d98b79137b94e76f29b062e8a0ed52b
z4339da5c2819a910b251b8506e154193005e4be3158afbef116aa6bfd9f92c2f835efc7941833e
z81a0f644b8d5a330923337834fb96627485a2a800f273ae3df0fddcf0c5baabfc7029102de3c03
zc33baa6c58b632e77ddb4f1177d8d4f9db57be48f6a05f9354000d97ed5c1656571aa46c6c0f16
z2e4a0c4ebd26971ea3932490febf00ea73abd0f4adefe0d23dda86d0ed86ea4e712cdb5f9fd2b6
z016e28950317d297ed8e1899d4b042dae48ef8224dc3b32602599bc03b849a1c9cd1c8ec7e5389
zcf40d82647e5470c246ca0ecc3b83e5eb0314d13c8157e3242ac642671766e113491a9db5e2179
z01755bf1e8f1a57b17f8db2a14526c8c937c8e660dadde63c6b8909104c655e8923a71fe147546
z7170cde9133ca50fe7315f4e9cfcac16c792535ab6ae70d7c04d408b08ec63b0be2d29e0e11b88
z27372afffc9060c466f6b322bee3ad5992663c60cccec2daeb97e701c2ab7d8d41ae14eb814ce3
z1e3d8d7ee864792a5e0d22aef8ce7d6fef2c2430fbcf37ca8954f9fd44a5044fd4750c238768dd
z5698378af48a97cb36f03f57e8b98b489dd471f197928347206656f31e41c87939fba53773bf3c
zf7df0eb7c8ab343c4ac88628c5b914d2482ee79270d3b33890b9a372f6e190d861ce6a3b59bd39
ze061d3c88e5c01179bd015999636f27c3bab6df35e7231f590bc27276524941c56132919c01273
z0f10b13956d5f76e1ae41ce9597cb9ae6be531a774d5da3c6070771fa47d735dfc4df771eeee33
zc2258de820a1878714804e83ff13b5f532711cd69ac4e273663978f65dd0c8102eaacc464c21e2
z5354d66cf924ef85149574d704ac9d556420e16e5a6b1612ea733fbe25742fecaab1d66506c970
z05a920bf8abebff5e0d848e3ee33f77acf7793c9725efb1ee56be33092faded1b1038822d84ba7
z2ef82bbae8f159e80119522a50b4ab6521072a00c5e8aef5cff2adfb5e2d8c8687819771767a68
zba5ec67f9531890903ffbd2dd65ba145eb9c997e4faed29c7088e7286851e1253bf41b5193527e
z458b757f25e37d1b469a4b3c9542f629771da5563ee3de584003458bbc27806d7e7f84e9c24a72
z8683bb743b8df343f7c7641e569145b1cf87fd17df9d091f523703399fc24c474c2e1a12a1bada
z10aa44fbc52cb3316908924e321b43974cf70b907882b1939706c70ab188974c2827375e735432
z5cf4738f84800da4416e51a58947cbf62b1d5ff14541d7f431ffa2311a614e240ac872743e80d6
zc45042d5a8dfb6f977b41c0f4ecb876939b1807cbaaeb0f6f0ade429b32ddfce35bfe1583b2b98
zc103d109166b4ec0bc6e752f2a67df48117d7515aebf26c51a289be2fe8979daad6893151f9da4
zeb8a64c46f41ca6f4ec62e369e9ff14195918e897c305b396f390d658c38786ce277b75a392618
za0be6ca7688805c3c52e7348d4c6304b96ca91d0bbc154c06760543c18a3a98f5f3adf9f999afe
zf4efea333e042dd999cfcb2132b6867160f78b3af0fcba8eff0fe6838ce56061a610148b630695
z4de4e3e33babf076675a5e37a764854cd6b62784f6d6ac642e3d378545458e777643fd6304bd52
z7e7586468c34afae87ed9e614fa72be081ac1b5db406b818fa29b5b03985a1c6f406e7a60d7667
z4a191fd3297bf00026018b30e7c94a9ff4546e475fb3fc5b3babdc4988df95a84dfb48a62dbf57
ze7a46d958cc996fa5ee6c6572cbf83c412bed46ec141849e82465b0cbad3e3e5273d6618f7272f
z2c3b49febead958a308ee96914d9b4e219a6daf9a39cb301b8fca062f5e4bddc2a8a964ec7cb4d
z3ee565fd57cff8dcedaa8755e26d4fb665e11170f16ca07450a7fa63c4c160112751c19180e885
zeeeab38e5e7c750e82a133c8a5208eae1967aee285fb577068d26f27a7099c933a7f27fbe00faa
z447dc420fd94275e36a5de1766f0a406672a9060f56a24d84a98b776d191706507b5a3d40b0942
z4b6e9bc85bd513cd41f3813c1a5f1e7e81600a910943c75d9ff470f01f6b57bb2760e30cab4c9f
z78b0f997206950fedbe4f2ef20d713a3d79df16e9b83e3fc7b4c09262427bf4dfc1569722d68ac
zf11127352ebb42c885c12b52529b012305a78593c4816ebd79e2731d123fa76c76c7def1856c87
zadbf76abb39831f5c2ed0456dec8db71fb03eae8c72e8898470d53194054f2d0eb03ab9a176f8a
zcdc2553223b2f579882f42158faea2e1ac5a713403777766f9b9250a65e5fa76211bc0e2a5f337
z5ed053a3b87d9ce5ac8366a8fb9476f57f558a2de599e4da9cc021b54731268b776d00bd3000a3
za4348d087c29269c2d465c8a61d105f97b0823dde5dba04cc0668af2f57f7ccb0432ee22a5840f
zf9938076846da44b163105c3f2a53411a76f59ef3320bd9b47bd3119813e14a8f2c96287f8d45d
zc003e808dd80a8d4c185725ab5849c9bd4bcc49a83bd4cb27f8dffdb4cd441b40a55b42ff9fda0
z9355fb27396ed066c651a6b3b6a0b45a0b741f1b0268e3ff7fec5469099ab6a0b11ea123fd5d86
z997b2711aef9c100ff8c7789e4b38ddbfbd0e666044f71b8484204e6608feeadccc3b5381920d4
z00990fbe94d44055aa33ce859cafa100ddb05fa47a52d665dd09980b8727085bfb39cba98b962a
z4e3a25487a4c92d621f033e5b7d8e411c872869c2fdbd2a59e8cd4e46cdfcf7fd216e42bdb653c
z439b007bcebbf4aebbb33c385b75cf75b743cfe7b1891bbf6e5e2935a7bb618f133de26fd5e1ec
zc51bcfc03969c307218dfe88380c1da9aa2b203d54989873a646ba7db2cdbac350e6e0b0f11b81
zc88479657b57f2bd8ac7db77460f564a7099e51f8d442496aa707a20402bd22032eb10e0aba6d9
z9b6f8444ac82b993aec5fea6e5aac54d651a46200572831ddfff19b02c2a2abe0722383d92a9b3
z60b54af0f0b4099dde5db9f4496d07ef087e3114e798bfe9716fec25ce3de7d5440be27f1c1498
z3b19513fe00212024e568bda3f20c045964641d8bc0aa517154c1ad06ae0c484870cf9c3184612
z09e60f5217b4f4049ee86c77978e5e1e09a0ed9efdf5ff9e24af4a114f877465d051c776d820f5
ze134189e902fb8c50b5f8f3f41b71153618bb4ad4a66507afa48d399b60ca94c33e6bb03ee828f
ze7e6f8083a2e2270a12b40da7f650e1d0cc4200d195e51571c66d63cbf9f7c4fd91d4862a45a1b
z743aec2c6b97232949a453ab523b716e40d8944803c9e2ec1169e2f4ef4ab7785b1372f0f669cf
zf65dfae9342321e7ac2ef5e38364c2f2563875ff313283e005fb817dbb2951961ec81d760b6d9e
z575d6463f379655444368ea6209f8cd43993988d572773141afbdf086a185530a0e50b6f037385
z75b8568c936df9ba4384e3a083c84bb7b6e5ba24ba6c9510eee5f852ae0079eca077a514b44ce2
z7259c4f95e0fbe48d68ef7e11ff537dd9c8435be253e584955f97cc0950a358ac622a084b1739d
z23a380723c1271de48005b8b2ba642d89b6c70a0e2ad3ef366d1c7d206b9efefb58759c9e09d0b
z566a1e4b5887fa9ce363fb508be2726c2b7c3b68027ac1916f85a40d89d15b670850f4c67d81cd
z248b782644d76c273edc564fdffeb2f0c2d9ef3281adabebfbacf9372ccd0e8aad8ce258205105
zb96ee0551e9aa5f8272d51f4574536a0f599922363ba6377d346906312c1ad9fbdb4625ccaf0fd
z9c943657036aec691561cd241500f05b3058c5f6b4b6fb768695201001c21702e4a9c9e9dc3d33
z42ea69694c6c890030d60a9288b91baaa36fe433c386d109db2db90b9fbdc5f05bfca9015cf54c
zdbe2f2d70aee9322c9c418576942cfcaa2d970df5121e3dc1ee8ecf39de2b7ad37b81b3755cd89
z534f3009faaa66c0fb6dc8e9d79e095c5329ec0edf9ad90a00e30e2a9f3339382ce95ebc834a4f
z6ffb2979b0beeb55429b3e254761d7d7fbbd22bfcbbcbcfd78d5d7109dd7f5e1cb0e0f28abaca5
z8d6251daa2b7b465b8a71f2800593010ab92a9bc41c240af4b429fce728d4653ca046fb348d5c9
z6477062ac650dc7798a97f38438a51b88bc5fa6a1fe0b2656d94c293ad794b15aa63d67421d532
zbfe43d2dc1374029d6813a189d59ab2afec7d7f7c22acde27813885ce101182e3d9d30e73f8c00
z2d74155eb0a6eb6f994989e9a6453f9a242ab9a907868da9fd7e8f5a610cc792d6b387cde713e6
za3da3c6443b38b1250ed6a7d9c700e2742d7fde2119c296507dd406949d77fa7a7b46b5de77d5f
z3549d37c9b3384b572a349a463b64c3e6332e51b1b8b50ae37cbba77c67874f1b7593037b5d815
zf7311d505505addf82519f2a7b3059d6e1bac393e0ecf12a27d3a71c26a8b670dfa24b01d029be
z4861ad7140c50f7bb515cc2f1315f4848b91fc28a6ba29c982f10cca034e2c76712db4e175141d
zc973c9c4d2952dd4dc92118680411aed60864e8ec72876a312bb515b883003527bac7b0ea881bf
zd8a9220dec79c18a31577ef401a7a0937dbc082ba33793e48964544be0354657efd7938c51913d
z05f5bcbf6ccd620ce2f5beacdd36c7a5a1e7cd44ae5423c10bd3accbadaa0f3ff7f835c3dc6143
z44145f55ccddc8616e8294a2c4542f062fff22286fa18528358842a89a53809d3832b89890af42
z95afa262b1885ce572ba2efdd680f33b814ca44f12e2a113567d157dd28a608f502e49872b313d
zf4f826d023bcd4ee72f64e9594e471dda496f2893ac983ed67d0321c1c7dd4178510a107d9cb2e
z5c13f141bb522518a9789ad0171f8ce2fa7517929cc408defe36bbe0e8c1cc63c7ad33863803fe
z2f8c5edf1e46fa76facbb6403b805716578f5d67af3336cdc6c8cbc5452770a001c1bda12354e7
za13ad9d23380c3bdb328a65307f8cacfe218cd1abdce56e992969449516a7d8e666e2e02195929
zf974b806a560bdcfff0f9ce2c42e293c35a2c7761f18fa5cc057a0625d0854dad9a6cbd59c072a
z45dcf6409f999e670459f565cbf5933e7806972518be6dfee02561b537a05ce44c6b66336df7a5
zc142a94554b7482507f376e537f46263d1974af507642ebb800f64ebd767bfcbec39dd0bb83bcb
z5b1d6c322c4412c800dac82eaedefea3bc3f6843750ff647e13fa21fc479dcd0e117be93c9b9a2
zdbcbe4652d9c6bf77c2571eb291e509f7213048fc48a6d44be44f1e7b73d914742ab524eef8c6c
zc99e7879159c07e53b91ba9278aee8f93e656191db954c0a1dd06babf12e1759d33a3335907feb
z34919858c83a897151c5e1863bc91b71dd7f5f30bbcb50a52fba2969ec05c8b11571d33b5bac9f
zee125933f4507888765277c3c89d7bec5b8696b4fa12fcd60ad568a6b91dab82f1ca6c4f2c2b32
za25ac800d128238c0f5921106028b878b0abb2e1dc559587d4025c6de3ba21730de9b1460b9a1a
z567113045412ebcdfa5199536403c17c0653fab756d8af3c7fc8535ca4446ec2c36ae94f39d5ce
z48d3922afcc5c38dba18118d2f0cb4b6dac87290b5fa668b35a10a642b51353bfa9339510c74c3
zc5ec3b612903fa9b6abad3d74c90eb498ffb6b4fabfc25c808ae4f9a68bbe66d67c7d61bb3fee4
z37d04e671a857ea8008ece3fadd8b901d0945c09b66c6a8d10895ac062cb5745af6f6df0b1e1ab
zfb765e8cabe7d70b05cd4f486021c22601743b47c03fff33bf5c5864afadc7ce3bf27d327a82a3
z8b2ce054069468b20ea862187f51383066267d6650e643cb1e5df4f58d10052b82fd85f8e68f28
zdb53f9a60e5d122f9be8284afb5c5abbb0a6bcdd613fd1b48d2b247ac14b88999caa0fa10edce1
z79a925f5524e523d9705b066237f91d6abd8969629e0ae5f51b0133a2d87fb32b7c4c8fc584037
z28320bcda985a52776e4b8ac1834a3f75d43a658a3f9a78a874fb1141e93fd469a13be00f2529e
za47f37c60f7d79f65817f9464dd3b9ae9b79e0948d43029110de01895796de30ce28f8ad688dd9
z21b798f1bfa994d7c9618a6a17a32967042c0e8dad21da62462bfd425a77a9169d2c95c528169c
z764084a0a79ca692a7f22cb38c27f0ee32d2cc3d7fbfcbee09500251f1d540af4c665420711cc4
z85323a7fa082148b3e69652c66f6084a83d4c7f5986d344ae4dd6d8b8a07db69b7375e21dfb3d2
zf0ec97687cd77f2614beb25fd062d9fc7f3ed8241f475097e20ccf8cda55d79016306184140ed2
zf42cf868458d7b4e4ec4fde3cde3e7fde48594c77ff517cdfd77a2e1c822ab39b966d5c73d709a
z8f945768ba575968ea49ccb1c698b8949333f4ccd8afef0a00f0843ea8e240837efda50b77070d
zc506664f0a7da4522fc682c400c4a187d771c0a7e5b6022adf33f2b0a486e8436b8ccf8588c369
z6140286b16c41b2683830170e53a083ea29f00e8bb15c773edc00f913194200ba984258a560920
z3d33206ec0e95c8b1cc57dcc1626807a36f2c322c8503e2b739a4b55eab098e65e473bd4345e3c
za3141c3ba74a0cb075f9ece929eada675f46230482760cd404aa4e929083b8f713a15e5bd9406e
z2a29be164374ea7d926ec4655190af981a7c4ef717867d793d603f8763803b7f2d785825d61168
z3fbb6a75fd1951213a470f0c57ee88b849cb4f47df7e12c0298d4d594ad7ea45d48b20e85f851a
z0cb80bc2075711f391d8d1f07642567ae13afd270c10000131434b9892a3b9807c788aa3834292
z4900e16d56efba28aedd8e1bc9f5687ec9d824524e9d638feac291679dce8600340051cce703be
z7cb951e15568fb52f537d0b09f33d1456db3d8eef8a316d72f0729b300f7aae21e2a53cd90b30e
za56b1d18e2356bc61edba54bff61c0402be0758b2345f339e2752aae2789baf87e41cb457fce0f
zd34e1eee4f127780af405289e9db811b9861c3a0ae1b750b5f51009ab27f7088c732cd936b3f5c
z587f78f21d4c950e78be1bd3fe888a54a2581113c1c5f4f4087b960e53f7d9f72f6206fd701b44
zdb45194893a3105d684c85ed7dff619bee596ca1f4b1c957d524e9f084aaa3c6c43b7ab50ce032
z255db938179a9569c4e2d8fd0b7ecdeb93644b0420bde75295409f425e3faa0324d5b5d1371714
z929d09e04ba8032bf2ff3942058835d74a1d203b61f6194f6c56074228434f6d2137c447ed2922
z78f84b034f2a96dfebdb820c7218336d348cc5b1e1fa39ec6e475d16eb9c9cab359bc85a14628a
z46992b1dbc96ab9ce75692f6a9f4fae8a1453917e85a8c78b22760f16c3a50b1ba91bdc6e86927
zbe3c296c41d60f9cc32b8f97bb4206f48ca5ae9f6f9e1ede870c91fb463ef528f57cd371185297
zb6bc67b65ae08025988fd04c18debddee9c50aeb6327d2563949c4dfaf3c62574f0279984d8e88
z2d6f1cf60df381ecf85fb22ce401655dc22f53c3713837158433fe8cee86137bad1236c9bad869
z00c5a647ec5fcf41073812d3c0621804b5441aeb7481092960a80a103cf159b3972a92862b88fe
z63abd7d7100dfda0f62882ea599139c1e2f3cbbe5a530a74bd6e2089f55db434124f223868df1f
z43da3eadb9bafbbce7304f4cf547029a6d7ffcf8f879f6d2e84ec3c02156d6d482a4a8e76ed096
z3967d00b87c06eb6a13728d31705988f32239e299f1da85bbbbd704366187e5b33a580041f3631
zdae684a94ebcb2c1f1cbdd311452d40b8be54b364e62ad36ea7ade34ed435ca9c6161f8e27fa34
z80cce32a3ff2f47006d494cadd80676eacabef425b4eda6cc471188d509000e6c0f187595aff76
z6f748a3b479cf1981f709f83a63c61ef3b517da631de09d1daa74e892574738f0b597b029fc966
zf923d8f5470f19a754cf5f7bbb2bca7f6564b84a444c056a1f193d044067f407df69a88ee5a82c
z4cbc9aa55dc5ab6e368b0030f0b5aa567110f8bdc80c852f932990efb39609f60fa1a268fae1b8
z7d6a2584c4b0911d26e5ef4532f8a5f1a055cb56133944c5a1fde34e6368c9a52f88a137f721b8
z5c66e004c84892659f3890c68ed0275d1b064ec9769f38e91c37124fcf3d1784fc1c3f54e7d04b
z805b12c583950670da3b508ff1a243354e744929835c6e89e52c63ea185f8c7444f5c9034e9b7b
zb8adfa0060f2798a590b863702bea21c1958b9ea3d752daa3f6c496c50fdd7c1c32fcba8965099
za0dd70b670d1a56c07cb8d8f1c9b0f54220eb80c42ed73da492d1ec545f7619fbcf6a9056997fd
z18bdc4bf313b82386c23f7cc9d4cca93f9433b76fc8c277af6f3003ac852359e1b2b4c1237f751
z0e3b63937d3d7113d2adef37c8de4fcc7b8735d989c87eeaf6e77107b66d69bc5f5f0a21370c9c
z439ff46947e39302a30068a16888a52efc264e978b2d25b4aa0591255b0e83036f1fed3d713514
zb1496cfa55947a5fa2a04fddd8e93dda5300501a24c7c73f62ad42b1b40ba7fec64ba41c5c57c3
z7f2d14fac0aefa45c21654235ebddc329d7acc53361b4d1b0eb104f3af817258ac30effe80d078
zfd96e9d5407c0ebaca1f96deaf11a69fc6438724bbff3051d750aac69c7050bc8dd633506a0c63
z9e44526003806c2b2c0c9139e8d13737b90c306f8dd36744ef0d94adad92af90c6df6286113386
za267d10f1b071c4897dde3b858cdd8d272560fb0260a55b4eacb165d89d21c9a59615ee0d2ff91
z1f040acdc1b02ca34c0df4616ee8d5aa3e54bd556b2aecc7472b025baf887aae09bc09c45991cf
z73328e847a94e41571986f5a31ce0f049214c0f961bf13e594be4e19e726c7c2013d4e50182e5a
za8ae9dac42b48e782ed0e3cc317797dbfbe88d726dd806ad10fe4d9fded7cce850d031e9a88a55
zed51a331b0d47f07087f70ec22fb0584998ca9ef62f209cf1813e31afb6750382e8f52d9e80a41
z7d52cb1249623aff40ffdf2ea3e454d593d4d4f1b81941b3229a0fc0284f6fb6475fb9f8e52d73
z01dc5f2d8621198c91b4362e1377e46a54cdb9cafbb684c09672da208f4e329e49d78969e4a437
z90ed73bfe201af979675bb80cf0122b4818f3c3cc2403d0969439969747cce4ddf95888c0a0e37
ze75f95bf7488943838de31a829d7885d5a75101da68bfe5e5f18aca5238d5fdbe421902b826633
z7e8ffd7653c24cab4080a08bf183e1ed1c5b5c88817ce565711cfa333d92eebc1f67d844dfb1d9
z6f6deaaba7495939625f3e09bd5a7a4e4ee55ac12d8e0a54c1ed36958ac2dea5d4c3ee5a90b04e
zdbba5a3fd2bb0e931bbf370c91c665899fc58e3acbd823cb54ba59472cda67f17c9b1dc12dff61
za99b8dcf994c000c0b11aebc92be48795e95bd0ad758f1db13d4b3b3435687889ed5ff87fad4b2
z1a11acf8cfe5ed86b341f2b7b9d71c0d1c9ab5ae55a5ab8e207b25db951e8a5c3e9350d8d6db49
z08ec255a675084dc4f477d6e2a0465a0021c5fe802735371086cfb0f86d98c83c140241f13c69e
za8ead5b715f4f166b2bec7a58e67d6c74cf05760466c8ab763e0ba343258d2c9e51f15e9df7dbb
zd16d1f673aff3c58f9725f6bba4bd5402266b8ec1abe218081d13d166a353c078268c6e8d20bfe
z225099b8f11852689e7c011f575b339c319de7f8984c318555280da51735e4a32d335881985671
z0b0ccc7bb26947932cf350d721764ec791dfb821db6da7871c1b7d064f0a20d747ecd574db123b
z8dad0f9f4698f30d3e0c2d561782bd56dde852d398bac5f3353bad24b6e99fd8e016b9f5d72a5b
z10c092358307694ae6c8f9cca7e6d52e15b2033b62f3e0ca14cd6c6fabb5c6135cfb611ec4d2f6
z5f1cd7ba8bd34a74e11286a0f948b8aa75eef4ee8c4741150dc2762229aa0e2ac40045a75144d3
za8821cac02a17a9c079f5f067af061fd91afa17ee6e7714cc873fc1cb2662b47fbcca3d3d3c2ba
z955d6fa5dfeda8a8ec1e7b5fe7f3cd5b57ca12a2321edbd67a53e1780526b7df8ea44c5c72af8a
z6c100deeb25d0424dd48314329f9fbf5fba3bd013118c4b67b2ec5b57891f6864c0544d18a6344
z84726ed7b76c5a75559f9b734e77f3ddbfabe1318ab0a67da3207ffa3ccb8ccb257f5dce803bd9
zb5dcdf1e666245a45c6fe5f355745e651be54754195425b66a57305e859545cf06fed59a327fb6
z0f41086967246dd6d7895edaf93828ed611f9b65ab53507bb05e67642d711971c068e49602873f
z5022d01d4ba8dfe57f1805d93151a6c4b2b3c7b3eaaceef1198487298bbcb0e986f2fce8a24dc7
z99f7fff19d2111c81dd967e97227c72605d6cab37e16f80a54d59c25249a0e932787eec6f3a89b
ze4da62100c7ab91169a292f063c7e5696c75f355bc459a9c5230b05eeef994be5610a1b99601f0
z65dab525ef37829173949b0618390b2ce373e264b90550356acd715820a5176667d1ace753dd47
z20e5e6ded38c9910511567539eab6c2e1c471836dcffed0678a724b9f8a72b39c55fb40cf349c0
z10b6d540269bab55420c4d537fb22658b981036644660376e49945407f221f628528ebbc8be9b5
z2e487fb9b8a244fb3e3b5a0ff536346e544bb689038dfbf1a8db1aceeb4f3400ab6e680c263d57
z542f6375f9e609ea59828a1aa65d902faac974f82e13b8fca6d3f15d1e32cce58fe095ddaa5c3f
z14fb84170a29460a1fb2e0896565e24119733e396939f2280b4363d075a4d274b3e7e74e6906c0
z43dcfac197fd012bf717269b75083c32a956848db895be14a7e4bbf77ce1760fb7cc6a58234448
za3a7f57c297a6aa17de63289a64e1fbbee48e84fd8e9491334234fa28561ea58af03d699d043c5
zb1c6d02ecd54dc664b0fe3216975cfeb8d1c97c41c305f4e8fe9d2462922bc351d435e90bb1e30
z636e9b16b7b78863ac39e40ad99c5821b8ef5dbf4a82689ad2ffe5bca023e282e4e98092981705
ze1952da49d421bacd7dba7222846e3b5e6e057b9ca0e5087b80b64c90bef68adf7b6aebb7a7202
zff4d1ea53cb4f748bc6515b99912a34d80728a445e9e22cebc0184a46bf8643962f32265070009
z56118b40e104966474b51881ed20afe89728fc5777c1cd3cda781bc0b67b42c72695c8c855d5e5
z598774d9eabc30b92006d774002e03d9dc48f5e786816b0b3cd4bb4287e2d421f5273955cfdae3
z19d864f2135dd13a07e776081f1863e7639d5a94f1e7e6cd529ae8f8908f4c363e9ebf020cbb1c
z1a0e5e73f800db64d4854bd7abf57d67147e62a5a3f9cac571a87d927c37fe82dbb7744dbb91f2
zb3ff06bab0335727d827fcd04ffa6e830533944e90687e1834444cbd625d2d4ab674cb7a736d9f
za44b411adecdff3dd236dfa8d3ff1ed3f02873c5458232b7890685f41070c38d12212b8f10326b
z7a75c061e3ac6b802d618b39b0e2bed9682a2e60e34210d2db9c268e4cc18000959a2bd5f1017d
z503c4aff29f2697b79f9064301622c0167f0c6bb1ae80f088ec05599ad3c25d0b499aba179b938
z059a9f91e0316a0050093e035ec3ad160b496b5ea8ede08c5a545cc957b643e36413cc9a851320
za75dbf63f9ae1e3089655b0fb5d458670938373121f38a0fa0b3f4e8e07f031162ce0da2acdcd7
z52a30d8af91b64c9b518b1a9988bd88e59d913b522b1130e91dc66f208f8c95c7619d4bf9a2e3b
z42d9772c3a98165615267e94471a8e4c983e7236fd461d30b3cf07a0dce4c14833f8d962e2df26
zce274b993162f2516cf7f5042addd191f97807be1943edd66a253db49454a5ccf7abe27b1f0dce
z4e5660982153c7b9cf29a605d334135417a9d6c68ee092d7087a398ef9c615df44d134705504b5
z42ef4832e5dc995653785d124c53ab5e64b838c613b5e31ed5e59cfce9ca0522305a24e42f18d9
za5935b9e259e97b95bd9f90ed75ff29ae61b7d7b5323f390cc21247b19011c6dbbfe0a90bdb1a3
za4941fe72ef1655e553f9c63a4c49ed06ce03e6bc1482e55422744c66bc9a8926556a99c457c08
z7272bec820687e13f462dff6ce7552cfcc45871138040856270dfbfb0acc986c4dec7a9ad3f477
z1df039fced3ef1a3e1d9f49b9dece29564aa2b3ad428f70a92c928bad392c794d18a428ffb0f76
z216a0ea24a08c8b58d941ae91d14317fceeeb2d41de1e363772a5205f9c0cef28fc6c237e3212c
z232a1b63994a4fe96937a5fa4501e64caa265a69556ae798abf3b630a251257f21d87efb6080d9
z166bae9c155ce27b246c98b58b642c01c88aed1ddf4644431c921bbeeebaa330e718666d796eab
zb8f8fbf94752774801dff60d0566e5d2c61f48f6952ea8ad67ff1265b40881fdd8d9a88e7eda24
z726533c1ca1edebd1d74d029f2efe2b76eccca841d890d8a5e9e9fb03e7d99261339f9ab4bd4b4
z03dcd972bae8722b603c1013f29d9b169f31ea73a81b1ad9ebbe01390cb1a54bd3fa1487620267
za1a8010de31a19f7a127c5f86d5a65e7a5880d0aa4144517a743006b6172f9c77e526f00bee0ed
za3b671016734481c5c2f9c11aff4b147d70ecfd9e0876af7be2d534f39c55888b99930e410f78c
z1ad3b818c92a9df36b1dd58f351c86b919ea3d5e54e1e8dcb2ebb27a7da36bcbfc579bbdd54d0f
zd1fe9f014e0ec8f4cb1ce8128759d0bd331dfa52112f5eafac4e609e757d0613a39a0d34cf7358
za985ceac4923b1e0755f6a14b4c58244d5aafadb9a9053ac1037961b5c3ce5a0fb65dfd03b9465
zb71545926379eb83d89e05437410e7fba0cba0e339d40c0e6b780542762d8cf91c66530f7ff8d0
z434dfc6c7b56c4852a41670cf1fb203a29e0d3e75b16018cc44356a433840a601b1b330ccf791b
z9ceb9005deec9c07402c2dd232380d29554303678dae060e16022c2a619ee9cff8146460a7aba1
z01ea396b9d1b00bbf7d0322d79ac419f3e1721762c376bc9229fc364ca4707620a239ade9f291c
ze2e2c1f0ecb51c648e8959fa002d791beda83f6c6d270977691366636464ef1d0efdd8efb27ba4
zf7ab330df6d443baf11fc72412f47361533488e0856e2e03cc8e9181a29fd61cb46c593b8ab336
zc9aa85c6060b610758d6ec9a14cb10c8d2320b6ac5a5e5eaf548526b090e363b94beee1b2d9d9c
z9a73dfd8af1208e57cd24a8086dc898544b7e06b98cda5ea4583aa7159ed51a0decfbcec90dcfd
z68e070d1eb1d634e182de8472a5d06b2fd4258a9bc372b2c1bcc3ba7ed0edaf0fe415fd26b4702
z6dc1e4aaf0739080145955c0ba7cf8fcb706e429b52fe1896373f9f63e9ebf9d2a768f312dd5f1
z3af1d683225729577daea47c021892300be5f045ff4f78945a1cb605c74a472070813dda992091
z5e3873dbe4219ea23abe62dfa64bd001e6eb01f5a16c1471a618fd5d34e85b2880f04fc1ecbedf
zddda5c6341a836e5822914f3da0be46dd24b346dff09b4605fe658acaae0212c011a00f1dfc54e
z28b3e84517c1c202527c6bf6b4e58b7f0422a1dbb82fae25e79fa446247279d9649bede6077a62
z12b9b1030f225e1c3aaec12559e1d831cf0084ff6f56fa01231b1ee04987514ae2b06a97817f90
zbe068258c542e5ea2ec1e4fb51cb26b9cfa2abb8d0cc9f03de6c3a836682e44da6cf9b8033dee5
zdaa978223ecb6924c493e844513118dba4a0f974eef58cd5648a0b1ba748f5557fc54da5ddd32b
z9ee1edddf9a01632cc1be9e98590232d21c9bfcd717675819ea18f7d7bfc98ce5c784af533f7d6
za9cf414cab2c24fef1b49b6f2509ae7756cd65014f95e4d24987c76b82a37c7972e10b70b8b124
zb5fde64d5db9e3262fa4119b94745d67909698b5e5f34c9b5d125bbeed71edbbc22606e08b3885
z3cbbd6dcc6c607405db1f2bde85b557b07e95b7423ed2db089ed55d9b048a4f6a71509a6a5c50c
za61a20cf5fdfd2a44d21d65b0842c1577fd7768070e5fca18b414fe88db73f7ddac6d7558b0058
z3396afb8c0a6693a44713bc56ed481547b0948c5e68fc03add0ed7a18be2a450486ac7eaa198d8
za5b248c997219ee107c9fdd236ceb92b5cbffb124c860cc7411516ddb9c77ba0f7e2a48d6c9cbf
z2b10516db9716846f5c62de8f05efa4b5f9d14e0512748fafae5d4619f8a998d9a3c06b4751435
z833151673de30ad252e2ccb46fe4d31b001de20377c0ac0c95209ecaba082a1da5771221318198
zf5c10c7063f11124918e4b0b8cfa784dfb89d585f1edc964473da8078d0773303166de13c4438e
z9d37a206e2d1c642201730888d5d442bbb0829d25eb7ee3a708a140cb0e16f6f59bea049327f6f
z75bdad1a62e271aafdf3c9b7d4afbb2cd8429cb9de5b38c326a44097478cdd481f4c7c690fc00d
zf58f2c380b8a823fc909bfd9f262f3b5d981145e9ea1eeee1b6c44844419a11b757182be8f096d
zf69af1fdc16b91f6fcca7577e2325d38ad427845d9635085da6bb3c8314ab37b0c3976b2bb79d1
z86789b166465b15735eb6ccb44cd59ef9c9c2e94cd1a5e0009efb32664573965c8cfba5bff9fcd
z2469da04939d4b78b504e6c3452cd710254b821dcb8b06f28763b3879dd8947c4d4804813018ba
zf1507110df4adfd10d1c71e5fb27c30e9f19d23fe6feab8eacb4336cb6e6370447dcdcd77520a8
z43c9d281d347efef6894659854b3b31120e0582fa8cbe2bc73e609519ad6e941f47e768ccdd907
zccf7410a3add71d98ab87c5ab09c41e7092d95604fb24b30e294ecaaad59745818319edf286057
zfdbadef0f639311e1909849c39cf0f85e559bf039d2fbbc655736aca729b6dfec052be3ea1c831
z85a8986cace4931317d9f4969fe18adcdac7d6dc4baa826d97a82e9c4d749d86280120f6b07f1c
zee088b5b4e258c31410c61d205700bc5e53e40efd67ebe14c26ae44cf0d901dbff58876ac0cd09
z0477d2272d2d63e9818920f04dc7cb10269999d863c16a51c4eb6e0a317c89b109dce3c011ec21
zff3cad26b3a25327ab24f625148ba386b992ad302d882ff89017e2903d82377d0b2fda55b33f84
z7f2944915d962fd64bfc01cc4659f57cf8fa941f3b0728c7880bf5e55f7327c22f2d9636175f5a
z9449f439befc59ecaaf754eb061bbe21217195faf742e8614c50e2684b36a0861c50cef23c715a
zf2e5ebd735b879a12f4148cc4ab740c52b51dc2df445e920bdaae2ebc700d24625ff9923fac280
zcc501c71129358e764d3b3c80d738c78fe3c4e3e0f46218be89b18939b6dcbda8dea08ae97dc09
z5ebd83ee6f4fd6540215d0129abb6ef5b21fff23a41d409ba3d6e03119aa8f2e43f0c0e7b0d1b1
z980f573c5fb50947d191e0531366ae98c8ab60396eb8568c096ec7d5ca2a9ec916a0ec794c3cf8
z3585f7b540fadd4ee1
`end_protected_0in
`else
`ifdef MODEL_TECH
`include "qvl_sata_power_on_sequence.mti.svp"
`endif // MODEL_TECH
`endif // encrypted_0in
