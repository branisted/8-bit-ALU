library verilog;
use verilog.vl_types.all;
entity tb_alu_8bit is
end tb_alu_8bit;
