library verilog;
use verilog.vl_types.all;
entity tb_subtractor is
end tb_subtractor;
