`ifdef encrypted_0in
`protected_0in
ze74c34e226135848fe16db9ffd31815111b6d7fb642c521a3f628cf6da949865580b22efd062a7
ze90adae0e65e66a2c36a587d0a790699161455169ed55a01f2084f11770a774ec4c588039b380f
z6de9c5084882a40b79a175f5c2114b2b6d78b070cb806e1c0aa9258297f4687ab308bc470f0040
zb0b1de382961eeeaf2e279e1462520fc31c119af8f2b214846f56c2b3cd2eadbe4099496abff18
z15cec83ec4a77b868344aa20ba7360908f5c0de2a79abf8b3534b883bb12180f68b5d4beb444cf
z3fba8f13afb0abfe8fcc4294810f75afe452434d2d0f1166236c82f76edf1e12979f04bc35693e
z32ae028996dd85737a8f5adc1ebb94f39c940246e887647b64782cd7ab429b0544c173176cede7
z01dfb26b1f73408344a52b7e1f117f12bb9c8077b34876c2e6fdc085981637012dc9754765e1a9
zc512ce062e0b8fb16a214591f5c81e1353b900a611fe1f4886b57940b41b7f2ce99a7b84b04b90
z916f717e73bd10589c81e207ed77ec660a8cbed5b487fa50acde1b055c8870bd8676023f21ddcf
z9c98cc47cfa2d654ff1365d1f45035a045a66c5dfa8279050262529d2cac9e64fd27d9c7de62a7
z731bc808811ded9016570962244887f98fe5440167bd0088f2f049df882af501358497c3b28776
zcdc5426c7f52a851c35106bb93e16fff98478405cb2c034d92a13b0536cf592c53efa2bc42b272
z5c52ed0dbb9ec35d0cee158298601da1f4ed68fddab40fec79905f12dc96a8110d8da442bed2ae
z163a3ad607d09d5a631332004ff962ee40ad88fb1ad2c6bf195702b896261672803134376ccec7
ze5247175339dacfe422e9e4fbd7d1adb9b57a18dbdcbb3bcf18f5d8846ecb4275215193ceb22e5
z98ca68fc05a3c074981f5e777b55bf3f9bbd22588d203a76377fc6313ddb151546e0eefa84f473
z85ff408a765533f621864e92b7ee7483408386cede999c577f802110b4e3e92dd9eec85b03bc6f
z4cc8a053d33cc32386da8ef494d24c33927f6a72552f22d1ac8d41f8c4afbedea8a94d26ec0e85
zde4b03e580bdc879b4ae42db2c5f2d039383571f964bb7466f382ad319d895262b4781780c1fdf
z14825bcf6f6fdef7df083b4f6d01246af7967a8e82c67aef1dd5c7d3beb76e2e0a251fd69dfdf0
zeb81e7a839b7c90e6fa72f331c89f21ea150f1e3c6949af27eac36f54b553fcf49e42e3ec12e04
zb6fe6b98218a3c450f754212f0290dc401bae67aa3ed9409c551af30c3b1cf5bfa8074158451f9
z0f4d50ce21bf5100df7d495a784ed4576b10d866174d6150dd4e0c798adf4d10d6940124d1a6ce
z8fa3129b2a8f4352d455148aaf4ac1fb85dc4981339fa7d67bb4604949bad28889b66a7ea746d6
zb403d00eecf7cff0f2667ba5b43aeda1f4d1b7b769bad6adfd0308b7108221993d1d65f4b320a4
zb7e28efaae50d3879ae8535c8ad9010201ba5fffb46490525a96a8910d3830e4ce041ecf381a36
z0652336b00c5d1c7d2babf02bac340d9713e960b6aa1e3fdf6ebe1a0d0c356f187d9ce4625a6ca
zf5f39f11847e5c85df10d88ce2e7e8830dc77383d9514b760a2bcc05e286671893232eeb916b45
z5338e99c04573394ff20fde7c316b52accda1558a0aed39f582779dd54bf1bb338c381aca93632
z0f08fb1cadef548d4ddc9875a3184e22629c7d969227434d1076b4d4c095a9345d8a654ceb1210
z1b4b2f5452dba083c03d4a6c5f4058a2f26f07e5054d7bafd1bb1702165e3792afa818beb1cebf
z6661021c70be7c8c74690d81048cf69da1dbe8f3a666bb3e7b02503bca83cf92ac4b7d3a05c6c2
z9139ae962308f568e20b0b67c6a1deca05a00f5aaaf83485b4d05ba6e4f176507f596adbc3d7f2
z11e48fa780bffa7989c0a378e1ea6a12fe3ec23648a4d323a64029e6f46dd875719f56ba1cdea1
z439127e05666301f6d2611cf7105d1a0c0bfae50ba84c63f3db2bc14a56e5ddb893ad096d6d977
z06ff57889dfc527037894c0512708a769e697e68f9d018574429bc3e8ae4a4e3e04aec11077101
z435596a0418ad8e256d98b57251649a488c61345b76e91cd0b6d6547750c28224c025a4b61cd12
z84a76d44995693e2fd616c79da43947879e7d50f03680198655169671643407e09acc649fc3ad2
zd066f546d833a6396485d518334e9778ae0ce1caa653035613e77743abdf5f044b582beaaee7bb
z0c1da327f092c17201bf4cfda168d925519964b2fae39b98b6fd3780e462a70b2c281206a14b91
za684bb1d63a8b3d71b6042a265b02cddfa4cb5e85595f370967e791e9c1ba9abd0f5d25d3ae0f2
zd5e98e92df5b57fecfc70340b6e1e41e4058fcfd72aa1257ff8c369950cd488ae82359c917aa29
z986143f7d6c34f63285ba0606f5bacf27609699f5b34b51726954d0f82e91633a2db23bab75dfb
z265fcf37cbd96a5c592985e4ad2cd9eb583afaa77244fec1199e769929c1bebe9b85e25dd40aa1
z69d7d43383fcfe7f013fb2a2036579b6c0246991a7bc76e146c349c47354508ba8783d647f44b0
ze8e5ee98c3895312dd5174fa885d58abd793c2a05df38170a13e8293e9babade7649ad7ee991ef
z97c0015b06d627a378ebe3f7f9f54ad62e90a16f9d5c8227c1e60b2c1f44748e2f132ef79a74cf
zce6a64db949a7f95f1ac60f9ff0990a2b004e164c35d4095e5a5665697ab87d527c6a64e5c29cb
zf81126672a72a42450c8632e30a342d94d67066466a8dba7af860c493d3ddc4ea6425f58b32aee
z978a26af82a1fda59137fb9f1fcdbbca438b0bbee805f8b24d353b0c4043d237a0ae9abde12dc1
zc9affc2cd0cfd7b069cd9d4abb232d5629371127c66b9ca6e2cd6f5e3c4becc36bfbd5c0916eb2
zb4a481b6003a74d9aaf905021a1989b6fb2032832336ded0bfd6e040131eca599b6d99f7c170ac
z4aa92012b22cad994943c801641c98c5a751576310bdf6cd1f2d11fcdb9add171b50932524c038
z2aeb9f566a9c9598da571145c0e98ea42dc09655d481cd5d818e1b4f5f66ea0315a17da25569bb
z8f2fe45942767c59802f0531861f6310efd097efe19226fa9dae19aadd2cab874d0bcda8814ae3
z7de359c417c590e4fa763b604ef67e6387cee636941e08aa24c7d3e13bba5061dd58fd0dc5620f
zdb7df643f1e5ffc053cd147624bf656fc04be1a442c16d5a9827eb9fe4ba58ddf98ac471a56fba
z8e9edf5b7ea3bfdce389cfd79fd3f5b3be78762a0f1ad636b3020b9a781d1ad9c2f495a22fa945
z469a909335e8111218f9d5be989294f33571438f01fbc302427b26380a271aa2e0469480cc6611
z42d8d1e8c09e307d5bb6598d17c8cee76492ed6962916a01dd378a2c6e130b83397c0fd519c3ab
zb8c2ef62947a866a5c435a1a035304000e115e90da47b3a366f8787d63be2e4610cc9f1b7f2d12
z8d44a4b43ebafc8e1c619c163591303af03e7438a5b654ac797618c982c4cdb4d39c011fa95ebd
z8678dc0624ef7772ba005ffde7bfa48cd16209b9a8901b9a5eaf87efc8a936b778b5a77389c820
za248db1b7e5a70cb3b164ce07a6d3cc25755d920878a9ff6f8c40a5a09aa69463a8ce6e5603526
zb64706351bab047a73728edc6e17116e014a489768351ac6f4f464eda834c037fcf2b5bc51552a
z05c4d64bdebb5f36d6b4b48c54b340e21367f7b911578392aa05ea19dc46fefb5d10bf08859067
z783c67e248cc1a772843dc4f9c724edcd61d9b5cdcf4f5fecfc77d4bbb0f1f34ad75e3e6fd41d0
zcec577fcb61b38fd4249ed6751c08da2d91851beb561e03fbb4a645929da62f6b2b103926f6402
zf5c2237871d7fd1100e188137340325d193a8d1c111636c10db82039aa61be4ca02e1367b0fcce
z3664d08373a35deca933ffce923fac314ff6e11028ecedea221096d73c1c35bbeb398c3bf8888e
z5c0033f1bde377fed7f3949c238149a93861bbad1a6a04d085664f6e9e31edae5ba6475976e0ef
zf2739bd9895f73b08e7362ae9644f8725e707182063fa210b6ce1b6e8b091e9ef8aab06b67a861
z191a51a1b665e0a3d10f947e0cded3a86ba561d76b828eea77a19bbb960308e12851769d9c1ba6
z7a5f68d4bdf69bc8c9488dfaaabbe79583cf436a3490890d95eb1b5614655a2893e2c055c6d087
z199b7af14a2cd821d2df5372eaa79ebe5219d12272a178c7581a3aa7bd8fb2a0d9a52b11c78935
z5c070d9c42275ca71194c8b936adea0b8337b32e49f93b7cea108d9482a9904919b8957f2c3560
zc2d96ecb3ebba55114eefa9b456d0ed7733626bba07422ed0fc4b6aab5d46a880ce7118edd346b
zd49a80dbb5b44956a29b8b1adfddf817508d229c6de462254a0d9faecffd38aaae315f81df7f07
zd95047d2905aece76415186facac86947bb8736dfd82a71ee40fbac8755a53577bd6ff57b70b83
zcde911138e5564e36a6fdff8591df7031ebdfbefb2bf9d8af6ac3918d65450939b04f818dcde95
z41ee53082e7ca85a68ca079bd26a52f2e0f56d38170cb9ab1a1ec990c9c662a7085be007371548
zd3785107fbb9041e7947aab3b3f20cf1e3575ee677b1dd2038eb3cd757149517478438271b52b1
z7cd41cc1c82c4e5bcb3035f13651482a615ea011ef12e2609b9047655fa9763c22410de6b51abb
z908d8055bb5aeee5c4ebaa304e7e1a9e98d9c3974b0c3447eb39c7930300d5456efa0f676aa646
z73166a31031d0c7e3c00750dffd3c9e3eed6094ae717292e342600528b6a9e4ee83b2a104f9dd1
z2c363adbd044ba191437d2b52be3488e1c833e5010e676835b016d6650af7ca3a4707359e37678
z3cc1e18b5f9f8525f170ce0e29445791f3fcef56b2c8211533b51d62f1bad0edb84459957001cb
zc9290519ca0bb7deaf4152c6f14818c78702346d5a87df0864bea2ecc089153b9ad832b2c13f75
z6f8f1a3103b9911294a6a314f937336ee7e0ed6250a9cd13742e0d88e63c38a998e21d0fe8e00d
z13a7a5f6b1f69e2d6511c7a5e52fb957d3b012a35350c5ed596e6fc5d21e53f4b16a22608ab186
zfa3762ad0a215e900b7c06f659b7135ecfbebe2e2f93540b66340a5cdb2e96650bceb83dbfcf81
zf6e6b79ebe22f829f96cb15aea0bab277cd401a435d2fcad5ff7786530d3c6667d1af985db16b6
z374bda1cf910a8a76d0c846c26db01773be74c5b4e1fd8529f2ac235504327b4e8f4f6deb1761a
z754cc47c5c9f9bc1514e25eede5bd2791a2d9286b1da3105e607160d478fc66f47a23fc5dd318c
z34159966ade1f78b8ab85e4c86d6326c9c250aae13f70f0f4e2589f0f91943975a99988a76cfc3
z1a91863dbdda0b917e2a85c635e7bb8dd358c81771d1cc8bf7d3206e2ef9f2b64feed15eb3f034
z3e2c09404a1067d512ce0afd7e61a8560dbcc114cd48519c04aa68d19e230f100105b211c6b68a
ze928fe6e90e1ef50c1ed00e5155648e2251373572b313600baf89cc67c13ba1005e04ab322a093
za90cb9eaffe2f4803176ce1d0b05ae97020d96ff27154d03ab330b429290125d32c0f760434db9
z39336ea11b7c7536d5e32e5bc20469b75d6d2fe946795588a4b5ef4d7fe76d3752adc4f2eecfc6
z0f2eb80cc6e91edd3f4d5355765b74dc59e7143617209f4a4cd5394c99b29d797cd8efec06d63d
zf5be366569c77af4a9ebbe5170cf175a09e0b15f1eca2e5134ebabd138883f10b628acc1076b98
zd96bd6dbf3410baa93994a29ca201fd820212bd04cc734c5b9a404eba84faf4bfe83a3f835eca1
z245e7fcd7f5fcae086c60a2dfc13fedbffc5b60143bf1adc86ea6253146de8293eff5d0d8d1795
ze7471e4b0d94b58fd34fcd34006b6bc18d67b2983a5262cd8aae65c116f1b1a1a294a9411451b8
zc290026e74e6e58306eaf9cdce42e66cc75143a60428c1acc18d2cb68efc034d40ff93ecd14e29
zde1e5e294a3204351c436d386639d427a4f3fccefaec134da254a8d91a89a7054b27845bfb0484
z2f86edbebe8b24f4a4f6cf9e085de0feda03c424a3bb527d24b707f950974942e0c79988ae6137
z6a23b5857d912eb2364452238a4c43cbf4bf20032be6de4ca6b013d09e1896c06d6983b8a4a4b2
z7d7e7045c99180df0406fc0a6edd3df56747175c1e207b38a519dbc75c12f62991d048418d95e7
z24d9dc33f5abac0d693c9752f9de752759188847d44add63a564867f219a1db574394d5cc1897d
zdd5fe973fc1742f7272cc37064ecb85ae008e3e8aee8eb041b300208554b2a0cf0a532c412c78d
z5c9b91b6d57167fcfe6e7f80086f7ba52df00bad8f68589935f34fedebb8b2a30ad09f5f1cbbe8
zcd169c6d3dde81702c66a5b555a5bd4cfb010a85cce5b5d0788e64d865badc784078de013a33f4
z948c6e05aa171d0984a076de19b9df448d9607ce8fa6b2268c5c3c7ce8929942cfb64afb83effa
zafd4ae2d3e1a299d8e766b94a760bcb1efa859dd259b28ebf4f6f4a8c6fa6ff3d2f7ab563d4909
zad0f53d5863450eb5c4e33c03fa3f017ac0f3c2452e10cabbb470f32bd9e458500e01fcf89bd7f
z195c2eccd43f4c788719a5117c1838561573355841ee2c1c86195336002b7f3c0c5d608a9fe9d8
zb553de5128415f0c6f8be8513d0cc536a74b4662500e8cf4e87fde2864ded4b26b2dc53be2c53c
ze6d9f4a361f74d444e3d823a053fa2f6f04c16c9cbce7f80a2a425526f694eee5616aa53ac6a2f
z577be64e25a10dde17e66faa5c6f51d64a3442b9e6510b87a7069deda40930a5a2dcc5f41e9d04
z0b2c9a6cc581a616b3862b5db9977d34b1e17bb3b025972c8311beb8287973cb7d3fe3c365c83e
zfad6d5febd2346724cf04fd8dd2f80192d1fe20ea242a5115b2236eb0e6b5bb2898d0434c467d3
z09f552bd5c5eb0b586149f78c989b86e359c4a817c12e95f7c2dea2164266623b8489722596c44
za191a05afbda76ea650f45467177fc9a3a82b675605813fd8a6ef359eae19ada684c0803bdc54d
z0dd9bec9295fdbc49b274f927758cae1fdb3840b06eca045e4f0bb87524a853ebda7e528d3809d
zc0c21fd1d8a447010b371c1b0496a68a85105ad86cdb80d3ab2867bf9f84ea26fd1514229ca784
zf6415f009ab6b0d90441cca74ad9d401e0c962b016a20377bbf20012cefc017a2b0e44436254b2
zcda84e4a29eb207cd8acde305e5115fa933004384abd71d8f3d116b10da4f15476f9f5298829a8
z3768788670a50dc9c02d781b34bc182f31f7000a6b9aa8dc5a2efc763d94e2b47c283073dbdfa2
z654e55f38c877107a0473a6c2448f11434082aa6cb00088f445eb44dcbed3c933e4434f52c01c0
zd62f48abeb4cd88428abd372863d2033f4d0e6c91b0a6588609aaf0cd327e7e22a5a149c21fe54
zbed9d2cdb2b9edfdcd64f276f2ed03d0bc64b753144cdfecdf0537f64338edc5fcf2692465adda
zbb11fa4a96f6a4bfc46608aa5cb8d049582e5646f833dc7e980e49b1236fee29e823bd1534c7e9
zae1c75999c902b7a6eeebaeaf72267e2fff32b32fca647ebb8d18e0991ced0a564db6edb0d272e
ze86d4495082f81cd100993853cbb52c47fdd1091c2b624c116d2ab0c0b58ff1d10ce9f30d0efcb
zdcf61fba33577c8355218f4a3a57d77c62d714db3409784787e65ecfe47c969337a4ea763131d4
z56fbf08a77640efd58fe22a908ff98df098081064f5576ddcbd151e6f2ae987c154da1091a6a0a
z8bc8745ce702acbce0c624538a65b18c675f63fd50138feb6aa2c70b1de1ee146e2811e88ebbe0
za371c7721b9edf50aeea7965f022663da418c0d18cd0a867928bbc2447e76c17cf8ada6c8c2c27
z662e0f1028f4fffbc40f17bdad0436b18f7a6e1f37bd5eb8482a74bb6d5c0bad9e95ba73d66ac5
z24acdcd95b0117c3d67f093d5febebafb07161c67d38b7111dc9c5e90778f7ae59ccacca6d2f17
z58bc91a8d01b4bdd9888eefefaa16cf19cb07b8bfffac684e7c2acc5a49da430707779398545c4
z910935e4b8c056ef70ee7e36f0a9a02f98d067ffc89dd773406786a0644469a133a033e056b925
zb14e87810de92b73692f58fb9613dddcd3260259cd76219894f10326868e76a7dd58a6c99f3f87
z403edc44e32b382c1d55137391e7542b80a86475729b1b98698943cb99d28a89c2cf81b8f7c70c
zc898b65ea703def8b3ba11341288e8cd17878e691882343e18e13bc1f94bc6d132c1c6a828255e
zc403db375287e32f5e0d354d7b1c3c7150f71336b389976111f10b8ebc7b618bc435d7dde9c963
z41307e91e4a326b6b620d7c0830e90efe718ff34d024b5ae02bc8be3ee934c1f71c7f1271e4d23
z7dcbe0a0b9e2e83393f8b78876b0f593ed142758d368f64b05b9963e9e743ea1a0c232dd3dca36
z3d6fc7b10cd1c45d800beed1d3358cdcb9b7a3683a46e4c7be51e64740afb78aa729081259499f
zef03eccb12ac70a8b2ee54a8c33a6465a3af7fc6afff39be6aad86d798f46cebc912cdb8c68ca2
z18dee539ab580c87de1d4a6bcdbd8ff07e180b05bf4a27b88790c988d4a4ca10ced5aec32a5659
zaf777b48ef9af960048efe53d400dbedd1b38379e7bd08db2f365fa96374ac91489b095126b83c
za652334d6830c140c7eed6469914d061af19db8e0a1c855b20acbdb25d2ac5ad78c48cfa9bb6eb
ze0c63c2a703f2beb87120b606f6383f94665c0951af3e116d7169de98b013f6de89cdc5513cd3c
zcebb0384f4ed70091c0e7f7c31acedf9e37ba03c333fb08f3d0b4761fab59c1a1fd2d97eac9e5d
z711958fd2335ebd0751f87cc5af207062dbbb18bb09c8d2a5c3f0fcd49cc8672f8fedd4b09d0a4
z627a2d34090a259665b1227f471d74c1b937203335f94cf6ec0b8be83b6811c427bf478a376926
z7b3ac37c5554afede8cc5cbcb7f2a52bcfd6445e7a713780dfaad8df1e08a8f69c9d47ee2b960c
z0581ae460467f0423f8da8499eaa2b6bbd0d795fcd0b3bcb1171eeb4241fac51a18841ebf8ae35
z70c236c962fbcf00668ddf78bdd956da470d4266eb0c09ad5342f0a88b6c35fa2ae7d947cb1864
z0f47ce183b4b0a75402ef49045d9bcd2abf95cfcc8143a3d15c525f1eca26c7fe56063f2c23dec
z8201940ef470f1f89058c8caa03e886ada16f24fa57dd5a30bd35d474ec27b0a046a3ff822e002
z7b9dfdc7265b9cf0cdcac0bebc74586d40b7d26c933b89c115b83568f1a77386a58827dce0cdf4
zbf30f9c323d5b8f9d02300b376b0560df25dc37ef7f15fae1222dc0bd54b5029203f1cfa932473
z589df07a8b0139a6b7746fcce8936695da84fee98744f83337aa7d1469d0381f861c33ea874ae4
zdc9f31f3fb70abc3dae62fc52a07b617eb787471ed4bdd1b3f08d3a15f386caabfd93d1e22ca1d
ze18b75074865787e4996deaeea2e5cb2f7479f60cc0a8bca25bfa370c20cedb6838a810c914384
z68b0284212e8814c2261e9f222fa153f026ded900e2ce8c4ed5028344b596cf07a5dd524502068
z26fcb52551f87a38e4b491d46f0fdebe41e3d10ec01a0d4846d0589c20c8941c7d49f88c382185
za3540cbcf333f8ae7cee1ddeddf80c460ac64a5afcd82e7789c08b9769cc05a1b65f2966e5a52e
z94821b040a01210e65762b6b8aa8d3d10f7c39bb13ad70b4e854306241531d0703aa92d77fd2ea
zea964668aa86293787618a8a5146e45747facf2aab672cdeaec21df7318afa5d9c28eeca6e3e1c
z965950242d273ae6225c321c28d8296dead1a58b990bacad5e7f74bd69e44ceda879bdd72760c6
z6ce23b40c12a7976fcefda852a99d4c1bb1b845199e6447e422f8907af9c4b333d5af1b1e73062
zdb6ba3d8c0b91d7c799a236208af94b99d00a6cfe40e534e7b26e845e6f0c5660a0eab98184788
zbe9461818aa212a6c06f2539927562040ea152e4b663f21fe619d12598e8cad2fcb5fad7eb4172
z65744762e3995cb99ebd947713a5bc3e4e733d6e0986a86d995425641c6619f56e88f40f8f4f9b
z0bdde8e38144f684b3d6ceab31f27fc4bf7e7b6d2b313fdb42a0030cc745294ccde4d1f1eddb97
z7c3c56b6ebc5450468b7bf3f6813d19dcecf6eda0865faf49baf1110d8aa16f82055e558f14966
zab04a03793221879b6d919a1cd9a51dabc26bdfbccc3b67d63fc2ff9ec2e7539305b0072113a2e
z67668835613c6018b075be5de0909074b173df74aa8a44897c321ff06f2b67edf2cd57dc47d02d
z500681fe4b5ceed932e5c2f2a0eb563e5699bd03d40bfa1382f8e3ea48c6905afaf94515b2c002
z03e9bc96786169574e8e4b1f6c87d3a600ad93456eee31d5afc77ae1ee3572418b738948c568ce
z3f1fec57110d3daf8591be970ba347b09c15639c37898c54263bc41b0d5a0d4a817fa79366aa72
z2614da5acc765b932cc4574e50c0858d95691d0f7ea6e28628e995cf4fd274a020d10384240811
zdd82f74a88f8d0830108cadd1eb933a9c2a5fc194f03ce09dba5fa92379ad973b10db312a8722f
zae7007c015fd97e7dbc600d3ebe6db66e5eda49e145bebf813dce78b70aced76a2a6a69e919734
z2dcf2367b10b58016bbc8cbc57dc3f25c64bd65885df4543b24e04c5ad7c0b20dcb35df1385ee5
z4bf827e284c805d2b82b874b6b28af3939fb4037caca44c4f8daf0e47607e7682662e5c7b5c953
z0a40eccad77b6e73c983d6d4027d3cc4d94af418d5b7624aa83c69a2aa84bb74d9bc334d535087
z6715c1283196cdd698659bc46e8850b292655dcbf1ca37affb36b6716f91c39e105c22242680a1
ze0356cec89b61cebdc5877937aa18c1322e3305e8e155d5285981f71820e18ef444a25235b3548
z9be906d6a6a01bc1611dc61110b77a80845447e347cd98e3ec39467c674bac12ebb9f9411001fc
z16af48a9019dc82ac654923e9fdcf57ad4dc0807b851ed06e0ebc0126bd10ca498001df874f7b5
z028529fbbe00b0e23861753ff3f71218d603aca07357c59d131dfc339f28766415479642e3394d
z7cba9703e4ad1be5f988ab7190e480e010ee1740f37c3061713fbacec0b1034874d19cf0a04f51
zb38ee59351e3f3a83dc72efe7b5f6a5b0242de6c5f617adbc7d197ed93487b717fbf1955179aff
z7e5b7aca05a210f03a605cd1f62b690afa7c83a41b7dc04ffab0e7d30418bf84dd8e71735f4380
zf22e3a9d203e2e1467afe2698f58d28664aba40e1847e1862857daa03829c0a199e53fae8c811c
z5b8b3d9094fc1ea73a875d0b48619319eb5979b07d4801114da81cf5f50f58b42989136c5a6818
zb855f44f65deeb85def6191028982ab1b49d36a493607cbeea92a4693898240f8a0316aaf0dd38
z6b3019ae5876248694c894d07233eab399a4f194102ac7791d7dfce9092adc81ecd08cf2ea7361
ze2b13bee2febe164c897e495223b8935c9c6e86406a9e83fc61e182ed9410f82107b85018ec5ae
zbd633a2a59191083cbb686187147d699b001c3625e14bcb21d8d2437b8e91984aa79febd6886a1
z7dbcf2f295bf8a16e408ba9a1ed604f22484de8a7b9602bad4585df2fcdbce325c8453b6c1b564
zb457ed37eb2ebed2941348c4c5acd0e7e76ba4b7669474bc389a9606bbfdd4625edc93ce0ff6ab
z021a9a88dc05ff1368f0725e62d4bcdf00beceb810b130d4431933f3060354aab299977aef11ba
zb9574c5efe3e7dcd950fa5068dd2c378a6692c0f495167efc8b9c63186b49a043c5b864b600b91
zf8b6e4e88b4bc9e794881811fbba993c7b58267ce18ca39a8f85934fcfc42b5b99a93a17ce4fff
zd8f0d843756bd5c8803b81f557dc6dc78a3cd7d9e7d3a83abb3c62ae7c2747b7caea56a879d71d
z873c18c80802a7fc2d660c7182fb40c85d4fa0f8d77f9db8d9996d6304c14844f21102f3cfd69d
z1d0dd50ade90b3f3db6531a4f4134b3b1b8f771db891dac3dd8c52c966d6e8e69bb22c91987647
zee5dc6165c444c94f51211d6b1a6de14bf92c6176ddaa38a2d0f97c6acf09f4be787b21e7c8c3f
zcd23bbf8a245c453da479212c8f56a000c1bdee13641c450898a4c489ce2fef27582d387a8bf67
z00a695a084f31cc5f5b37a0c1785b6928219b5e2a2e55a26cd52d5db1149b066a51a9fcfc0a039
z1d0c99b10f15f0af5e2b0a1b0ba372afed6e87086751ea43fb5d97003b0226510472dc46012da0
zd078b6337a7ba7139072b378da83b9b019239a1f89766ac42222120fe9e0b777c6e8e9bab2b21c
za9e066f5e992c4167a186d4e93a05315eee71292e35630f34958c1ca6539253e6fef998b8db389
z95414ac80838804ca565a8f505f5f9a204c97bdda72b806ea8c01b14c2d1ca14f4a245edb836a4
z02ef55062930b1b030772afcbddd8aa778387df96c34ae032c6d8090be8025e16cfb3e2d08993e
zea714c023f1fdced832229cdee6d3f4a9b2cb69d6cf920e3ec985adf3c791e7501c6663e8dc05e
z9d904aaded94461bde4f5b829fe193bfdcf5d98765d8b057a756f340034b50b41ea3838437b51a
z97369f848774baf780c499d529b290499d5b8e5550b600a3929e5e6fc0bb3455c4898d6563820d
z33017e7a07938abde54e8550cabeca460071747bc5b23aa38b7c6dd82ba7573b909b7fd9c43991
z966f2b967736a03dbaed56ffdc7ae808c0d732cfa655b80820c0ab1fac2eccbee9f3c1737d7551
z83368ba226ab4dee3dd92eebfa5de34b8db952814e2ef2d1a22fcfe3b2b56b1fcd53fece928b0a
ze504c8e4b56a5e3e9d34aa55839a972c30ac11765a43101ab20ad2e313119b920ceadd469d80f2
z0b80229dd9e050a063bd5efd669747f2dd071e621cc72c13191662c19087348b0d2d61ab1320df
z5feef4df90936fbfc1fb4af3b266570d07739865e393cf4bfe2a281737d5f22a5247d01dc1fef5
zf1a9df2b15851121f762b4749a73b2814c767db1454e022e9daa7c10ecefb129fe04789c8e5819
z9e1b480be2ea555c75c9b7c56c91ffc20600bd7ee9546a6285f5817abf2e2303e48bf4fb495a7b
ze1e111cbc8f07e89848747dd57f13fae3db5de87af3d4ea712d4e3423100234a087cc3aace7881
ze9bbc2b241ccefe0a884d0bc63e84cde93a8cb984feb0303d3cfd79010694e996377dd06b5e201
z8aed3f084f29b017046d92dcd8940b9e67cf0a614c1952b209e4fcd03569f913b2e5c0c8b4376c
z51487474f503532b1c4fb090ff8a2bc9138a97da3dc2bdcca5949f2b0e6d17fde7e861375faecc
z3e7eb48b2409abe39e17680456d7f1b994daedfd0075de59a895e7f7f6dc8afc63b7678d623286
z377ce6b9ad552c82d755cd796995e7d6b0481e285411eeb4499ff7e82e7f2c3301a2df7969be77
z39a175db5427b536b4f30507598e91f030d978ccc1cda79743c1426e69d3f1edb73e6134153db4
zfa2ccaedea03f833b86aa7b975cd95f8dafc56f09a2fa3877ff749c1fcd60da1036ad490ac5315
zb67b9ff80fa790162fa9dd58cc74823ccb9ed8659d95cbc1a9332f76b33891c65bd0d5035bfd7e
z7884b8123a25b03d08f29e24d9daf13f939924d4eeb31faaa4f0bb1b970f4af5e93656e6ea68ae
z9bcf33a39aae7311291852d124621c5ced7a8e0c0cc2df83ebad6dc9ade86bbf22387ab4b6d485
zc69b8032de5ac01e5cceb5cc29bc0bd84f57155a02f1ef0557a50637c2f56dc22e87b8425267dd
zd594ef02b0fd44d47d1059fe653be24fc626a52af1bc2d753ef4364b31ca3af64cde3280f39d5f
z9e27f79cd33a498d4edc87d28c3721978bb2c0bc7e17d6fe1f3138b09e8acfa954f0ea28621e71
zeffeb6aa79c950ba1c8d3993795b300d7aaa59795be0fa79ed71ddb80a4001b2d66a3bab47eb66
ze8acc583cef185412e157ef08d17fec7800967f5cc0e0222bf7a14014d1d17e540611a065abcf0
z9bb7936bec44b13f5a7b6211bfb87b8dd78ac0ff52af2796f120f0b810862290d48ea8f3eec420
z74db9f14e6fdd33f23a514742601c305b0ba0281d83bf89d7cdce39318c07c9cac556af0ac40f4
z836c24dd3487a53cc6ae8ba522127a1f81a3536197fd6a154b9f485a378dcfb480e7c2e1b63b3b
z4f748256524ac5e12418bc4bf153eb82cdd75664ff803f8b01c537d47bb8237acbbd433f1a92a7
zeb7e20da9db0133809055167a63b3d2415df90d6126d3b7b34991ccb5efd7865deb3b697f4063d
z78d71cc76d6dc150d4c4e7030923025899b429f8401d2c5ff351d991ae617d3523964442b2c46a
z940597a6e49a570b846597c6e799d70829934ddbeaa8a1e33881b494233cf86660ccfa94030aed
z8a40130b9b8574fe7576ea52005693f64a313ef8544313f0aa84c31a00efa060b6b386dfb61b9a
ze314c8888dac800d28078f6bde8489d457ef90468c3f053a16d1ff87957780a27ccaa2d5f455c9
ze13662f191b6eb6a58e5b4aebf9eb504e346ee7a1906e5eb26b50ca5ac6a1d4f62f9ad141f2d21
z984c66e493c3ce0ef493c746e96a05e35aa4eef6007e463f203043d00eebf619828ace95be959e
zb8b6b718a88e581dd626ddaf08bb01c3bdf6db9819aaf9a5a0688622c486b82ea3f7c1309f60dd
z8ac38c6724a4dd6ffd505f96bbbcda54582598f4c3359a0bdad3a6688353f8b0504b5c27fccf5d
z39bad8b26a8c37d6db67f577efe9027a8604c8dd9a7f3147077a6d61a3b342797a810f2df4c241
zdd4fc543409e23e949fa6a987e6f9dd929559c248588b81b10b4a733928678ad5c9e137eece71a
zc43d5883b024e76768b9add4d1fd391e9c357a20f8ae37d6bbc2458062a6f51b3232b7f7e9510c
z15954766d87b122242b849d8c930fad60616bdbc373c438848abe1831cf5261b30cd5737938733
z57e86e399d3d953dd2a500e7c40d0c5f0d86986ed3ee30a8c93fe663069ccfb9a4a458adc7ab98
z5e3461f01a2a0607c654cd075dee56e5be66d33b2499841dcb5c6375b699faddc0656c134e9a06
z4fba2515be7caa0f75a6aae84eae8a4fd4417b9b81760ef415ea74e0d7a1e8461019bc0183eca9
zd53d159822de377b371bfa6c735098bb16fb6f621192a24bbf103cfbaea573bcc4615cf94f8257
z79629e063a7be1701e4a3b027f00ecdfb5f8ab3c4775c25d556e78b3c407d4aa49767b7c224ae7
z6b6479a2cc12983b511bd26acb936b2ec6e268d1417a8272c62522ff739d679231adec9d00860a
z74590c742c54d81314b48309c499e200cad46872d5e3d0aace0c777b0707bbe02a7d91036061b3
ze6a3d631d3ee6957b5ac47ece286d42b3084c8ba0da4447cfa7ab0e736e93261e40599dfbaffcf
z6b53a21bdec93d9460099fc9ca2e57ac4ed470526cb65f42671155064120f03797a95b5b8d77c2
zc4b8682a6ed8f40457b323cb37a3c944391d0a17710fba7f3859e899f4e1dddeec1eb06fa95784
za071e2e13eff793cbb5d4e86450c75210b57b4100326d05e3d2dcb01d09fa2f4fa5d56d1a59a35
z51f9044d740619abdf943b4f90b6eec3f8754d95557bddb679a8887f468d07aeadac7425ff28dc
z07ce2698f0569e51564a50003f35e24ebdc4fbb04a3063cf28dab31c814bc51027f4e4d1770bd5
zff0a0d7c8c9d9d9ec731849ae21786e0d0bc06780b0f7e105d466d8a06613cd8b914c21bd56255
z4e534c59045c72172c389574eec1dfd44f9078a3300ec40f4ed0fe4c426753c7364fe570f41550
zafc9673c5abc1a743cb347de9cce04d1d512c43afdb17f7c5795a30ba2f07fed983ff5e8bd18f6
z95d3ad87da28429cf5514d9b7829b6f902f1060a885b24ae550d099aa54e394263898d4ba8fa96
z49b8cb671503967e2b71fd837a8ed67a7842b6af9ab8dce70c8b00a509ac1943edb9b0f9db4dad
zeb2928b7cbb0c5ac7b1a30ff402fbaf51f73122337c2f16d18cfa857f2cecd9040e424b7c3758e
z0fe4c105c6c87274be068903da19c6eb97c44e8db02e08de577a1fc2518069cf1a82d714f36cbf
zc9624a9525fca34d899963a40cf5d741cec3693ac7f922a8e74780e0f664498124bdb101e34273
z0e766ff7b3ccd22ac60278a8ce7d084e9e5647ee8b823d6b4f17c4a813c0e0793d45e4ed3ffb39
zcef95f3c3eafddec5c675644cc6e06ff03b0ba1af71f4f4245ae5e4473dfe080fb8b3027998d11
z410624e23294720129ccb1795ff201bb9490680d988a74c35ed3d60c105a564d93a7dc364e4588
zfae7272a8cfb5aaefb1a2bd0373766fc55177e267d71072e2b42a4e23afd255de13c07c534cbc1
za46bb8dd70b31e25bcfbeff2703b094d9db425f43852b8a8700bfcb259b19aafd467ae2d0bd404
zbb3acb1120a7b13aa837771048b259d2ecf086bbfa0500d84814c37dd00be4a5f724eeecaa448e
zc660833183ea05170f55855ac773be33d9a6509e37b0072a301ce79858adb6296a91a5b0bc9b99
z4de07092b41f327297f54d222704c680804c07b4dddf38efb452b643e35627b2def4e081726fbe
z51275440532a912ecb758cd6bb014834c50934c84d14c88f8e5e5954dfc5e8679cfc67a192a8f0
z0b6efd0b4140943649f4229d45c1867baf813a406b806b5d2fe5fdb95000f935841151638d538c
z2003977bec3ecf62fed4bf3ae1500b834605d97dcafb6ac435c7cc2b5a78b7da338df76d028a0d
z82b75ce59bc910dd57c246ddf35add78f8419c46ac4ad53a783c8479866dbda52fcf3c44ea610a
z0ce1ca1bf8a8baa89fe8214fa81e1620597aa93a571571de25c5108ad6c6ffda073ce7c124ef30
zf47eeebc6d6fc22420dd2421c9f00b9a2acfc738a1abf4cedc49d0b989186106c386551f2de6ba
zfd25a32d3d377b9903d7260e7740a338b25a90ad3b60874ec069b2198a1942aeee598d74188d93
z9dcf9f079ce7edb602822810e91022c26c5815c827a735b51a536959e9ee364e0e502619b19de4
z88de17c4657a8aa93d85dc6ab50bc7ffb6508af653d36c27d6910abb12e78b3c518527f2d955e6
zf96b1436465c658764ba8eef655363ca83a71c6350d41e10f22aceb82caec79b85d51825030e34
za8d3e246540854f45ea314bb9f5410549fa41af9a43ee2ae41da35ec9e129252a9089e4fbe2f8a
z5bb355da178eda17442e5375853f2bda4964b6b43c8c2e79a1e33dcbb8d83b75a1cea6fb63ccd4
zd32d47875a7e45776bdb7d9d811810b7d79c24cd340048222293561302ba71d92c64e85dd42d71
z2ee62ae73ee0867c8dcdfb0ff5dd15c01b2351cd5d815c447ee2ac826c921e0f1e719edc777fd4
z53b1b6647e1b826153f904402ab261cfc1b7c82044fd3b49e734d5f49c786563ae72be3e141ada
zbccaf3726b7cf997125afd9e4f1109a9a63c76cc75561396a7b626e3f594608131f75246a27246
zf1f66b783c59cc5880b61eb19c3f4c9807f956df8f8e422add836d5b8749916571a548409685a3
z90872e048a6129654babd8c054b13b9859d306439ff726a1a2e72025a37cb23851ce21859b80df
z58c3ed049d368d265b4caf8bf4ca290e1fdb93dac7cc8083203d1eb856cb6b3466669923f8373e
z5665b1ad41a08f567a1effdabb0d5a4cd99d5181d9b8401f3f6ecefb2ef8a50a67dbf27938a01b
z45997c9c490f637eeb073c910a1926c4e31d5f2bafbe4deb6aa1c0a4f081d268a7f740039231c3
z6fc5b54e9a4e6cb6b7bf9286094c8fbc10095d28e91454ac4a942947b2da877c054bec82770dcb
z8022edb6998d43ec987944c4fb585b56707d9636d98b625bebc600d1178b9cf4bffdf01904e7d6
z491bc3b883b479c3bf1c1b97b4ade2725f95d13b5b06373043b9ef89707332f280b0f5334ac007
zedffb52f3c67b57f0530ff943be9e3b846d8837c6e2976aa29284850ff8ab35e47ced8b03e504e
z964de9b83e220cb07fedb974dca083019cc8a747f0e21d5acd91802e6dee65da8b1c2592a4b55e
z3c65e33a67473541f3c7ded29e53a9f45460b862bd066bbf79e4dda7493e17251aaa2da51a1b76
z9046dbf6d1b2b1f47917b5f40afcb2474986c66b0613ed511ff02c6b8215dd58404414a047edba
z8ee7a09b293ccd09a7e2ec962d34ab8a557b02bd5dbff665b17f4d495c3ad3da40c7e9a6bb6459
z92368d0a0136582fca63cb3317abb93a27d4efb75cd2a0dd36d36572a15910342ae00d3e263db7
zee8cc8b434eae6fd7be6e157020a213d07be4620999b22e419b613fb1a32ec0b96bb0668585187
z1c820e9e05dcb440a3b68c9ba6453cdd5d9a3ca06c59d63e04db44fcd6f61b6b564035c67616da
zc083e842609f250b011e4252aeda65118309b5e7271e4f3d735c1cdc92822449f2d5f5154a14f2
ze6a78cd50c47ea578328fa69ac02bc7b9df2685c707241c2ed1ec6b22cee5c6b907fcbd6922ca0
z6985f16c55966e5d713931afb2d22f8e9fdb06f773601cd5edd9a902691cd98c1f65fb9a5cd170
z638794100d16beac0c7f60403c3a10e32fa833362705880830baa9d222941c2da23bb76cbf29d6
zaff59f7f48393a511487da1d7bf99910c76da757abd284b610be59c139b68e35e4e86f3b4f3082
zdebd5b8a00800c922369757fdc5dfd6aef73126c9986f2c1ed345bf299fb36a8b9c21630df60ce
z19c97133d15c08e8c89b35b70a53185084adf54bab3796897fd14b38807bb171b143fded704c24
zd5c8e3d3f605294b633465c1d56eeb045cf0d86e773e7b0382d33bfa90412263c2f2e43eff3497
z9343efc98878bbd18bf3bba1c32c6c9a3d406ecc43162bdd927eabcc51ebd2faaba93e459ca029
zeacb831bb8ebf6639fbc1a2de5aef06fb85ef8f59ef629b19a8df2743db3667b88d94a779dc3d8
z293214c03aa90604012f65dfd0933d7bae1cb783fa531b697d6f2577fbd4aec73bb5cd362b16d9
zb8a7a390c37571d1a131f66cded50fd76f8434ebfd4e4bd7cc85f586e2f5c7da5c54ee6eaa8a38
z8babb2af8fefa273dc6216232fb9f8c9bf536baa2a7fe5c8c82cfdd5507308c6fb202e1d1cba3d
zd447e7e76e2b8f4ed6b53b5a97ecea1abc7775c367d39e28051ec933ccdaf9d98d0c50055d4d6e
zd3a64b157235de20048d3c8c5ad1d86a57e09e92c8b032614f174403a5a6d5884c564f57da814d
z6a82382c8d70dd2dcb5eb478e795310fb26f341e8391f6a6b756ca669dd930c2af0d3cc1d6ef34
zbb33a1fe20b82212f12def7a4fff5d3eabc31a37e94bbf9247416ec2eb2962024c62f369612914
z755d51fa4197f505ae2d7b3e2811bf4c3aa28b564980e3b9cbca54c52aedc27f035c8b3f31c553
zd90dc8648637ce9e028727dc1f104a631f6d4d372f8339870970235713bd9408cfcc16b5b2cc17
z7a486952557cfc1707e8e926214cbce0ac32c7e46d2c42fe69d29d17c46e8525271a51155c5c00
z2582ce829efbb6de115f717d02b10a8fd69a20183e57fec234766a0600c3731a3d11592c750904
z250627fa2c91676c5e77eee3cd2388a2493d4e0d62fbb7aa9f1da0c666026ba50055ed44d89343
z05f65a1dda5da807f5d5c5affa989a3e5625c3e1bf060b78f2b055d505a430a31f76a34b038bdc
z14fb28a0af95726c920dc8a7df07f0e78a6dbd33a0ed879b7a8cae35d4d05be6524c7da3e520c7
z69235dfdb271edd06989e562370eb6c7ee2ef252b54827f59efb910be12be7e025ead210f44ba4
zca8d96c33a299b75f1929f2ee04d6572e862a7b9011ca10f9042bbc2e1b4dd10d1300ec7b47bee
ze7e8af49561b199154db1948c7d3c9e7576c11134685f5ee604558d6a8117cf1d614c511e107cb
zad321e3cf46610be032afef9d5140740846f0c932c589ed3133d6e8bd864ee9df6c0ca00a6bb53
zea069ce004704f85a92e94e9aaa391585dbfc05284ddfee6a087f3a6e6d60210f7b16e9768e424
z73ad3c2253a80abb6e998417fe1272591c1ced28bc3faf693d1c77e961b51e3fc125642343ca17
z83db6b36b49ca8e2e4cd34e2b30290d09829a7287126d4ad0ea0d316ec851b44131aef9a75f1dd
z66728a36b68a504f4f8ec0e3874857daac727905ec2e8c87255916f37154195dd5506bc842543e
z275dae39ae8fed73579c4e7e87ca8392aa9dd0064ea5261f65317ee81644a5bed61bed7ca8758d
zc24881a6ddad2e5425bf7d779a291fc722eba7b595f5208aadbf021eafefe8163f363cc2a2ccd7
zbf602d48b70aee1c12988c6ff4d3bccc70329a990de2a24e8e88d388c48eda39f3036d8cb53619
zc1a69635d2d51d42e758e9a23955d2afee8c35b94d748f65971ecd0ac44c677e73e577e1652e36
z247298bc25020d59677c65040a757779a91dd895f1e2bd0510335e683781ba69f27ca172b8934d
z4459720813e48caf2af0c9170617bc9b15595691c1db3704405e28871b4e546fbbff14178ad21f
za63b255d442b739968442eaeadca53be635e487d540561b647ad15fb7f247670bf01407b5a7bb2
zc26579ccf5689ede8b9e5e7ed129e40bac7ecf447572445ad04749633aebf5ff265ff7b1f006fa
zdd75647fbd559e25d15723d3ba549985cce4659b6abe46c69eed1b4138a964bd29f08e1ff5ce37
za542a7358573055947f7f9272856bdad61e2c1609600f26ef4499f80d1db481879c3407068f003
z632e5bc11bad71aef53648b466956d711c1381a072e9156bc395935c89467ac657b652af2e2878
zdeb2f7cd24e6e73f98bfc47ce0652909672d20e17661454e465ee7906ed7be0897381135d16a0e
zc29029213ec30c2a299fe98dbee39440967270e2dfec16ab1fb2292d0fef0047cf70092c68ae6f
zd8a2328fddd0baf4b072ffcc58a41a2153ba4c82cdebd073e66561749d246631daa5d72e60ebb5
zc82d10f2d540d796788045896dce3d4c92573ea493e0a6db4607672b6177fbeae55fe4e5eeb670
z5bcfe51de4e670f2bca1d869a7d7c2a2cb8988e9c7fe82d1ce95bae4f4027cd065a5a5375e8a79
zc9dcf641c0a5c65f5581699119f31c18b9e98c8909f59b4a042f23c846881f61e3ecd2dd2ea006
zb0868afaf1399632770c7fac62d1cf315d5e862ddafecca0e917c60a7fafa186d3a90808191c13
z5aea8d75fbabac25639b4f2c7be74b083c3814a48c511f335c416d11474e4a1afd8c6d4cb45b13
zfe3ee4a5a808ef2630443cf90142b0e4c12c6d34d0dc8d63ffa90d41b6155f79b43cb95ca2bef2
zdcd299a6840296abfb93649b888a6185ae77884e3f412930454ea71f532123a1729324c0c21343
z7a1b644becad8af5a4012be0eb68c726574b919f84ab7f14697bf2aaeb8a68ead9f8d4b402a85c
z98ffa118552a440cb07c7c1ba5b965b7b585075ce4daed4c3ff40e6390170a4706d76dc7325c42
zd186da3c82507485bdde0980568ec78357625bdcc77c4317979f292ec847460cb497685a7c2518
zf302dd25e2de94f0eb414deb275dcdb914d15128cc6f51105f582ecf8f81ca267b586930013eb6
z39d161f776f47230839b3f0aabe944469853ed6246be9251e69a23b16d53845f3ab72f12c15d1c
z26571f03e326679827689eb263a0843301fe7953185f9dea21da6f7ccb1805ebdd3107525282c8
z292a504cbf784bddb7317a05aa9be99aef93451f1bdbc995ea83a73caa9bbc46b7053216a9918d
z40c2f03eb906213a960e32a97e7eb0f72abd6389f349865b1227e243c977bf2f6c56f6261e71df
z1fe624b9408d36ac6dd3235370d48d230105489e37481c949e15750811536411f5b7f28396530e
z98060b727f25fa470908b6e56a63864f5bbb4de6843c9e2ade3d0d071920a5ff83326c54e12b8d
z12565935f5f75bdbd0249290ee1c59f276a25c9866f43d71c25d290e50a93c50120a9c6b496fce
z4d59ad333836d36baaead9887a03073e116e70861e2e8f9a04cf897ba913fe9b99581c84716f93
z3d42530bde4cdc5b7eeb831cb89481161a5e7f013b9c90a36bca9766536a1dbb451c3415fd2365
z5d72c513580dce3abf6ab36e253e1ef6661a31e09bd097c6c1e470f75a3402615bc62e42c4caee
z7bcaf002592a31ba92da222797aa67b93f9cdce3a2db665ab3c0c794636d732bc4bd709c2cc1a8
z53019d4be2742ba5845dd1db0ddca385c4caf749478a3a85cae5c51e435e25ad4943adaaa96cda
ze888b412c9d4be1ec82ae312efc623916727b7965612f4c929a7821f506628c77231866b07162f
zaa35d94040f7363ac05671b57b56488d937e16672d1f9e09fb63f11f77b36eaade1e4ed5da295b
z9278073257a80c88834549ed7ecce7ee0b0a144e20884b4c446269eee1c405673c303d1a87d92b
z48474a9e188ebb224d8d7bb7934f85be12a93edf060b8bab1dabf6cb5e113d8b676d9d4acb4450
zd7d381711f33a940008bb67a32a3c3a99ce14f015b6e35883df63e714d1ba3ebb0c7b870bcdab1
zc947ef12735495c75fb3b941444aad1bbbc96a19c554d1b47737a4dca2657fdd8ab2b40bae6b84
z2165b90deddc9e49237e2ee04ad3a8be3b97ed0cf4fb677e6cad0d7c476f05ff7422f420f3221a
z3074f118326cd5addaed1faffe3ed939fca60c5cb7feae1087d59b209f8ebd0ec75a3ffb7c6b80
zaa0e3b73c2522448d57ad6c3ce6b9d86c66f442a9d1c370d115aca3a9cef93cdbd9fc335eee512
zb7a873f5b55ecfa7f5bbe4d190bb73abe993469234aef661cb4447ee464dcff99b80dc61e95d77
z41d5273b8940b20313fdcd811f7bf9eafb968352d56624e5070f155155c06e788cd2e3060017cd
z1eac61b0a1c636518de88958be7699853b5f4bb9ca1ab2c3f998c64285703081227725cf007638
z70fe470df1964d42ffe079c1192059756e35be06ea44482ae752998bfc7917357047fa96b71f9b
z2284839249e409013f58b5c94a2165f630ee5bf0501aaf7a5457a718942a6169a75e8fa26be2bf
z264bef645acdbc73668512a2e1d13f1d7cbcf3b4a8ebc163b228a15cf1548add2c7fac952d2c8f
z15c96424b3b28c7e1cf481cde12db102013306dfc79f5b8f91d9b8771ff43974112c0b68861a3d
zcd9a7ffd734b99cd4e6a223a7c7a39ffecaac0cafeaf2d32d5c35cc887177a069a2c82f61d6c87
zb14cde189a2098ff5c3f340f2c288654507ae7f6a634bb2c0de65985621af32aab66a2997806da
zd3875939b0f82a6708d0d8b931c930b9b2c1b598c0e0e72f9b7c1720717ca5e844f5d172ec8769
zcf9c3cd551de80cc55489441bfad34125145e9755e94d62fb73926e02b01da55776148a190c3a8
z98e4fbe9ac31dbd007242e0b758a1796333a306286894a4efd0a0a5a2cce3c9ee982d3accc6415
z97ecb2fbf459a0ae414e7660d2025277bee10bdf51f679df491f2209cc69e40232cdc9e1f12c56
z25f2a5de2e7844c114308f71ce2a566354796deb9df161207b60319f1e075e3d2d8c4e813ed573
z4015a3d2e6e1dcd71564b615a088cde952a0ae865a239a4522a295ae534f1e3e18e634aef414d0
z88d712252e778770402e08221b11401239ba02f6cb911a62f809cabfc0a8ff2208bfd4d0427029
zfe5d7aab042adde23ffe6d743fdc138cb78895b5c80271dca2442752cbdec305785eb0db086d39
z97f63d27bdc657a205952447417a8bcd69c354fa160a93adb5c9882e3eaa24510183a62cf9ae26
z5c51656c9faf4e799e583b9b0d2d54d88854946ffac83becd80de28739c6a4a7cf7bced617771d
ze2ef7ee46dc421acc4483754e7f7a9804139dae562bd5df0e4ee55ab5d17d9897c77fb2385fe42
z9e8cd28c1f6d2b4a67bfea7b516e3fc083001b1d990c1ccce401de91bb8e5e552ebc2106535024
zc36344242c6f6927952e59a3de5e387ec5edf8a91b3eed338ac8a2d447f1a5c480ab841169203e
zfe594bbc183a68af711535fb3500f074f6b4b506d07b7a7d30767931508f4527c8b37658752530
z18a9dbacc67caa3204707b9dad34de7e63cb574dc65821fa66dc924958fcd4849709d04e5c5f57
zc4c8416e3be326df48e25527014d07c52f78993648e4094ddfc4d34108dba216399c0053dd16b5
zb2f617db8c9f9078391d2c5e8abc7c76fd1409109f4a6426bf444822e9d7b9e9b99b0a372b26bf
zfea109123469bf7f61756ee9035d5da52b8db285aa38d3203d64b82ac09c7f78bf97dd70785d6a
z1a1867d5790d9c33083b1ff5bd062252d59b9aa7ad3943a4005ab14e15d3c1c517430c8f7e144c
z575a7e591d2809134c3aeb72300420439c141f8cfe0e8cb89fbf1642650a122debf855e1ebe96d
z1acb800170769640b25259b47ed7ffefebcb60402025dcb26c077d26565348fd82b73c10e6fe3f
z6fa96d8c48d6044efd43bb9dd6d4b7c93728dd8cc5cdde43482702b5dce9809c14afb9b465bab4
za90c991462df85b2743385ab476a62d0e07a4c59b2ee3197626781bb6894ab6a476e72e079955c
z5c598b0b8500ae435a7bbf484fe790c169659cbe74c381eb96fdbf6e23d9ac24e24e320bd24f30
z4e7efc5639c140820dc37b7361b4d2c70485639576401df4d562464eb6f0e4e5184849a5d1e980
z45bb524b1a581d45092ddbc7dd58a36650f5afc93b614b3a6b12d60cb3fc452dbb3d6e2ff536ef
zaa67a7fadac987ac5154b137c9c30021f50d711cfa4abe1b60ca2c47bc931ec836f4d9214ac554
z4c1a512d16d0a5d885c599995537a393c23965cea22dd809377689afea8512076ddae1978320f6
z20ecbae0de76dcddcce488f28888b8d771d589107ae8b2540b1a5e910ea3d97efb78d57df13505
ze19183291544fa2ad5234aad48e8722e7796b68ba12feefd2f097f2b3386a54323696f5c15a6c4
z8053835e47e1e1c0f35326a63c272f8adf686c83f0d0316c89f96039d67cf6d4a8ccc35ca03c4d
z7d005c6fe871c17d27af3d1815c659dc6af5afbbf31d9c5ae9ae9f137170488d087b183d032abe
zacd923d2e3842c278fc1b68c45649a74f314a3679fea6cf7e370b40807c09fa912fef40d354f20
z7830763b0c83e2199a3ddda9cf01d30213c5977991ab2bf76fbf10f8bac68d5bcc809e94fe4e40
zad58eee0ec3324317b5e67c287ac7c9b102e565d581fcae3394009d88e4b0247d70055a2f70260
z48079aa343db9964bef91118d4482e461d04a7d4919de8b7bd1629d01746e3561139831950a09f
z28135e712a9ab31754fd4a280beacdace8f804dd91fc9fe3208a55b35ff0fc4b8303907e7778d7
z93341e3e14139a5374cf1fd1c12f80c8c6371f3c5915d10c52f02535d0cac9806ac14a020bf445
z8c38191c3a23bc3c0eeffcd20be8fe6a868bbb65620f6d6cc9880fe069037dcc7232f562fb70b3
z55c6fabc6a9b2bfc542cc2378f0305addb9b6036543acbc4b24a877476290214d481aaf6e2c3bf
z1a6770ca94319ed03f126083b3a6844e4f4925efaf225572c62b7f29d83798e8bfdb766fa58b36
z9def9c8166d38dd8b942c1b80957feedc60117b560314c2c81e9055eb455292143b12e7860b027
z9b2c4edbbe60e5ef175d166bc224470aebcc1dcf472ae74af6d83ffee1f205b7e7fce7871a99e1
zc9b38f116925ced33e0682ff94a41f3601f52e589247e8a31075d3f44b5f744d6f56abf6ce1e21
zc6921a7108819f9655af0c98338c1ca46d89407b2fcfceb201ff47e33c0ebee7450ef573592fcc
zbc5da21e64cdd3732f353df83a42e75b96491f6bdb703e8e41bb64e7ca5cc38de0e7e71f116a79
z4656ea512d98c740b988f7c383dc33b6f6226550de550ce884e9db74dadefd3ea90c8fc25fb86a
z1bf0999d93662e0b4a37d761619b080e0af93a69e5f179c5504b593d1496744b5b4177532bed42
z2c3208ea1814eb38c495e7f0ae76f33bfdf99c0a6b9189677c7eb9d667e91643d08c6aa5008979
z715b4bed05ca59e79affc07629ca652739a2dbd19c0462aa3c734aa29df3c9bd1c07a30cd64b50
z2d595f50fa8875e5b3d923dc6be3c2f31b89d04ab31926eef5e342a0a9fb5922dbd8d197496352
z29ef41172f0b01bf69f80b83dbe420c9ad19eedb879afa99382853f231e77d29e43082c6b65fd5
zdd74c58705bb80bfe6ee01871af72d3e9319c6fed5c153ba1b99a8e957c870f7b7c3b82f583766
z606e55d8ae3246ae8da08449d1d4198e10aede508fee8105c9146d52efcfa1a1c29a6232b77c7e
zebade165aa96bb2bce8b22c13fbac8b309c43af81379ab52f64ec463f35b69a234660f96afc293
zcb29f8f6b7f6e85344e1f7f427e715139628265da4061640f3489d41c8701def97de2723356c39
zd7fedddf53753d2cdd975ae751344297d7cdcb2d27cd2fb30a8aad27d1e175057942bc5c43976d
zd9dd587b5c1acc12a34438d9276369d86373e973457d098d199d93adde732221fb9594950f788c
z7b201ed140799171e18b78a7ef86db5c03e5fcb56b2885a93193059046941dbfa0c2facea5edf8
z3b50e515c99c9451892f4f23c028c48ad301517b8708077f4340baa1a27c09baff8ee23bfae945
z339d0dfa65ec6e8a477ef6ef3ac601eddff0e713fc4c564ff9183f267114a738dca0539aa243e1
z6e957f81923af54bd712eb9cfe18422b22528cae62dfd48c460399e090aa2ce6959e68a4ad5d17
z078dd4a12484dd7f5c0c99aaf6871a795528519231850866c7f2f4aed163e753cce0c924017c30
z423b62cd995627145344ad3feec90a94d8ca02e3dfe53087d87c11fd32dfc8ce559254298ac7b1
zd56a8c058ecbb7c16dc052f323ceb612dfec1ce08ec6b2a849d7b82d53cebde0bfe4264e9fd5b6
z7165d0840bb7e9b6544244d90828a1992af22b32a2b346ee0200f039ef0463f7139cb3888e9539
z25e4eaf3b13c3790ccb095d03e3a319f85b7f366db7cbee703d96507e7b6afae28b436ce9da45c
z8f3a13db39b98af348e5665cfc7fec33f279eb9ae2f7032df4384b18f2564e2dafa8795d1138d7
z204dd20d00c843a1d03d0d29dbb54411f82b538dd8c62ea5e348d7271d86b5763dd44132b9b4aa
z143ffd0b43d3a286b354ca530fb63cb8224a257b139b05f6835028e202476b0d7bf58dcdc4914a
zfabdf604773731e4b7a83e9349cdfa8377f53d09b0c09690511e8fcd39980c8055efa58e64cd9e
z34785daca2a34f973671fae017fdcb052615c9eb7201b8e32f5a44fd10c9cb050c3a2a3d38aaa7
z4bc9781e6ee817bb830e2a33f907b13f3b59de6f51a9a38e187be4ebcfc4e44bcd2bf7cecae425
z912534bce52464cba90f87f92e856cd4c72776b1105e936dd59abb1bb49b155ad118d008dcbc32
z501a386b0fef3ade1735dceb346da35a64939dc3c51a1a174db88f51a8d6535f8fb6728271a1ee
zbfeb874a6374787d08bf5ae68cb40df6cc829d64ff7f23f81647fdcc39636decd4bee1b10bea30
zada776152f8556fea3ae180a25ad0c0a8fc3be9215e7d4e422c67be8278c4e1d29f23c3ba7cbc9
z0e09991713d2c2c6b9daed173b6eb0e1fd51c200a8e567811f7fc12754686db8403aeae051c7ba
z251c0560f1a0314b8ae0f6b8c29569cdcccde77ef217e8f8653bee589081b8f872cb79fda6d163
zc5ec5160e5f69676e71d9ec0bc93b0e9ee858446ed78e20302c84092ba64cefcb2d91191152c09
z5a2f9bd1485315bd3545e71eda4c9c99b3caff8dcc89e55d7d86536b4985e106edefdd71a46f64
zeafb60be59113fbe4b5513b2bd9cc05af91db423120deb2a17237a4074dec338d7030b0bade175
z44c6a6e899962a8d30f126f8da137e93c3c6fa9d4e10998607d00a5766c179ad4f12b9b728156a
z451f2e5b77622578367500c1b48801dfc0a0b853108bb3a94292d8128723d7d3c39a453a367ded
zf6fd454e39cde6c08e25b759e76fe2e5a3c3b6bda06b2f71ecd813e6a8766a93bc7c0b92c610ac
z0e48f0211b92248c3849495887d6422f28db5425c88c8c971074c064802328db2f5aa7d70f1d38
zb2111b38b7b8d065293e55a881fa35734e57a777adca761bb359a6aef376e3d27effd71e44e0af
z37ef4c2e0d72b61b13ebee5ab9e43f43802277dcc88355de5a596fb9d0762c5c8fff445ac9a503
z806f342d3a2a92de25110e1f9d199d9e7ff1515ec24c2de865c3301bb46ccc7e3d45bf671a734e
zee4f23875ea67565663d1ec5b9de9889af6852b1b27da3c7df681253f4e356cfbc4613199b63e2
zfd5023a19824d238767439d2a9b7a37f64f2893414c6f49a49f9bfd3a1356ff78b7e023cdd73be
z3d6d1796778bfb1b6af23f6803de6cc6032ec585d405e2aa4628be3aa61ade9663b6c3681cac7d
z37504d49bf73ad0fc362ce5b26e3a0b40488a7057bdb1657c9ead064b17af920bece71b9c62f94
zd8d48f95c87eaba2a7272fbfb62c5c27fabd56ef5fd42725095722622bb364cb4f1fa87cf82391
zaab868fadf0007902a8b387664ede0fbc9d941603d717b396fcda251621f8930ebfad237de456e
zdb0a07700ff87060fa3af7c6cdbed9ad3e2ed5f7bf7729bd135ef33fca7114c62c3ce3027896dc
zb90d9961d2b56a0bf0fab6bc5e6725b299ae34ec9dfea0f1cfa74268e64880766fe803d570f5b5
zcec58d63d3409ab301642eda856332d8327f733eb3b83db26295393902377ae2f8fa9121aee1c2
z2c0373386e1cd6fe145dc19d4dda4c9183eb40e211780458b5724c0edf141535ee70ddf818dd8d
zb8e5e1a333296d31a77a5885610f1c02be2101714e0ffb578a3213cc9367c53b930b32e1b9da2f
z1cfae36fca0fbf71173b3d78f15fb3a684c4ebeb6a15fe78e48902deda78fe83b632cc2dae3107
z8c407ea4efac31bb50ebf4d14e606d7e238983ce387410b13f44dc54fb55980f840b069b592ca1
ze72b5db76ea1dca2da56e2259c5e2816668a5921fffd50f2ce0c54b41db8d29d849b7a454f7828
z0068e5424f9ba502f2e3cc1265ca056e0c72d5624a5969dc667a2b6bdf8f80bfb02b60e0a2b545
z7c12d3ae837eb51f2cc84790127ff86b642a39fab5885458fd3dc31fa54169cead3fa96b5d7845
zad270887dd1f94fbbaa5cd3e2767ec6a6c4f73d1462ca3fe488fef1fa863cdf1a20545df956e1a
z86ef23c8d79092d97f6b4acfb8aba08caebfde624e1e8ddad0edc1b3b85e8c30ee23f5e785359b
zd27cebc7f0052398db295c65e9f83684242555bcfee87413144f12479524aa5c98cc11a2962f7c
z0f4ddcd00a36b2f6cb276610615ed5dc52eef9e106e5c51590e29915a32a49dd356a02596373c7
z6cf05d842738b6a021d9b4aba3260b71a433de90c64c419f693f351446b23f28b94f0d43786130
zb5e28a202e12c69fc5ebe1bd4f914cb3ddde572f103ca881140d7f4002365ab76eaabb069e38c4
z189c70afffd6bc0ee0ee9360e9dd10535828840031554a58e00b343feb8a3ca01cd7cff14294d3
zd5937efff151feb242f4ce450371b06ce9aa57e26c275cec755e98b60bded2d8c732f7eb6b5b13
z034eb961441f645b85cc225e015f690c051740f74b4d94870f986fa1368b3e4824f1f132ab54a7
zf618a4083d54285b0c8ff3a210cfcf3e36640e8f8786126aae574833c66a45d7e23d7cb2a8f025
zd9224deab17fc139c83967449205582bc0ceef7a8af0389fff63b9e6b87904a0958415d3f6397d
z4a97f62eea98c0a8efc0a2c4042e5b292a923c84c36c18ba45fd0c1b28235d985a0d3f2d05088c
ze296848ec8b36e1b9ebedea4ec3b28950e5e3b60ca26e2b8719db64dc2698275dbeabde8e80cdf
ze204e668c2f950c31885abbd99bd1eb8e908cc0791aeb274cbb4772ed004ee39a50ce6ec1e43cc
z10603d1d60ea448dddfe6d76264fd8e3b432f924469fe94fac27784d6fe888c7db5fd125a013b6
z2edd05a95620954baba1b675403032a2003adc9cf264919f2feaa8ac0a57fe889edaa215d412e8
zdf4f460542232e40b393f7aa3ce41fea3d82b0abfe6ad659fa705d85e0d67cf482c8a760cf7539
zb0e088984faf30f9eebf32ace0e2f91c63c598be53485874d51bd5815737679c96b59102cb14a3
zb5eea9f1b1062d73c79d6031af9238fc50074904d775736dfaa6adc13ec9b150201b3763028339
z0f68ea87e122c07c02ea1c73f5469878a21aeaa76787852000839af85780d1bba462cba3de3f28
z7ce35a5cb4e1c6156cfa79ca7684278a754cc8ef90ef6c1188d28958785fb6a75be896560ff2fa
za37ba652731d3706e130b67d4796668cbe7d1b460ae51fb572191c2a7ddaacd9efbddec0cabe17
z13bbf8ee809924527c12680eb56c73c8f816ad3dcbd9a3589c0d6dec052183ef9066bc94258ece
zd9fcd18a06c1a3137a2d620076a21a786c28dca88b065336255d67046bb65d557a6bed6ba98965
zf09e4c1da11bf274f6986c94371ef65f7c3f79c9035f2f5f4467d80fd738ae73ee6fa8a658fa66
z5b3c8baf3692775cb5b572cac92afda35b776295594a86c81ce674d43dd573b2eb2f5e04bc5780
zdebc26cf642a3360c8b69abdab2da659848ce3deebfab6991d72abd842f0cfb99d8bc38b9c89e9
zcb133b07c6624f6e63335117a53111ba93a4369475c961dbb957578ca74a41e78c8ee6087f2e39
z6e35f54764f53112cd1732a66d361cb9e1bdcc3f8bd751edc5228cb23823a1d0d10904a33a2653
zc7725182817057969941bb16628b8bf18191d7f1626880c9a21bdf9a637c54e536270fe659eb83
ze58ebb0e212012fe666cad934ba6a24b5ad1069ff9cc44c5f6ef62734d29ff3a43ad775a538ba7
zbe33c4ef9b887654bd126830273711619d4a0deb06edd2637a744413274f2c97a9a89f1819c1b8
zd3758c969bc0a5a83d3a03b9069ff1a4af87f94961754c81bba37640620de410dfdc8cc2c62cf1
z86c835dc30f58c6e7d0494f5340a655e82d92b208b6eba8d6dcecd585909e68662b89595c8c4e2
z83dd9baf9d3eeaa5ec56e21a4e82197b304eaa1db68c3b05b2311662fcf5be1d8accb7fa660662
zb443a215eee56093fc6c45fe6b6b9599a084dac2d68fb28913d6180fecf76ca710e48c1b8dba37
zc5249764b6516987b237e31e5a4bacfaa8b15fbf5714535f3f7cb94d23e07a5097d3b00727118c
z0569f6dc86ae8ddfeffadc50089d381b23d2576f318adea5998e8637d8495761da458322549b1c
ze51851295c574ac5a56af373a7307a65c8a84a49facd77736dfcb06eccea88f82cec9321da7d77
z82766a93a0ada451baf91b5a492515104699fddf3af048bf11b39d2e69e338bab063eec599eb58
zd6df5001682153c591c3adeaa79814194d7bc07708f7ac111b7e741568f757827e0ee62c93824a
z058d567df166bf7debe5647613ff27d0a9a0c2a388a82774b6a3402980954f74fc945f19dcefe8
zede625b1e35ccffd37b2f86f61415786025e2bdffea860b41e09dcd1ea23aa54cca6a240e29a9a
zba19c60f08daf952645349adddfee6c7dece27026f65c191125fe77aa1040f889d3145b134f974
zc729885373a25eaa8a621d1b721932d101b1353f9d05802545a18b823314a49cdc27b431061567
z6d7e214db07b153f9b52d7b21121b7661030e4119b0c3658af625bf6560b6869ceaa39296173c6
z72abe7ac36e9e29655d4029a83b22bd272325f9866fdf9c63ff850fd0092b3dcc2cf12c03ea5e8
zc1017a14dd33f963f303dfb64f305b4738feaec8c0f7926f88418685535ec8bc631693d16bba36
zfb936ef0b4a968c22c3c35725a5d512581081c463113536aad0438b9d964a7244ffe157ded381e
z5cafe2311417dfe5b3abd64aaa741af35d19f418f77083a24b26b489316b80854a699149ba28a5
z4886a04b3cce932dd394c200f65d99b17ee91166b0c3a9a89c9a017dae637a817b2cca95289d41
z5a925c96e5d9f8bbb15dced512d725e8e32dd846671dd2c88cb06bc4d916608057fe44ecd82a25
zd405fde6f24d707187542f16a954998ced835efd2b49cb42541a219ac561e1704640fe17a7f492
zaf2e1c6df943f46fc2ff7a0608a6f1904074c02a9fbed1ca1706f44da76106636d41c26f236373
z84a370343fbb6c3c8550f5324c1ebb6cb6ce7562347f5b0a560d747c8c06046297a66f8b482de4
z96d314e66f3eeb7c26e424c01888e4802c66301bd84789ff947f4bdc3fb305fa76f87e6083d0d8
z83d4084ae0ee8dce84214dbb660b594bb7b20345f53bc6f73d0ea5a125cec1d7d757aeb092cbb1
zf21e41449daa5f3419cd46e33428a384efe5edb9c74e8b8efab794f8781f0f2cfdf41177e53dcd
zd3a5d79c413688babd5e658b2766867b7ecc7a165a9705e2934b549deba8c18cf293defe691b71
z380885be94ca653ae1e22ca22c1b1f024f4a18d924b438029a700bbd2452b1b0b41eb035d1f954
zbf9286af809205f810d5cb6e522fdb03060b859201189e5e8dee27b4ee79a1d50be61121013200
z1100dd6e5ed0440487599e2c36e270fb659f466bfbddba1413950724b25aa9ca8fac0b817fc11f
z867bbcbfd88b45603951c7590f582fd4da525a2ad1502f24ca7b18b38a4b08ed922f48f17c25a7
z734dac90211b49648ce20dd90ce23b862447f637c31f20c40b203e5727419a572d7966b669477b
z303c98d11c93ca750893f5aa336baa0c02d2ab9e5a03412d2a11db37744d2df6cc46623586f59f
zb14f0da6485e5cd4f44a11c54d3bf9ab35d3414c161ee7c7eb2c3d73551b2649ea3785b0b6a5bc
zd9dde0e17e7d6ef6503d6008121dae48adf74f8d51cc5dbf1b5ce0731a12d4b7125fa71c276e62
z6d702130bbb145a2af4011d0dc794bf75025e1a14fbe4bcad33921b5d3f3515a1a1fafe3ca23da
zc6f1e3ee1575f1331690b2ad54d01139147e3e37f4f7d2d974b35b186f412e66572b687f3cf430
z23a4b8cdbabfbba8b28db00072cc64d0b01203f05effe3507a503a040a0e54b6592e3e5a71f76a
zaa7b12cab498303f42635e83e474da3c57440330fe059f7aa6c9a77a466eb274c1645a3b2a9de7
zce57db001c532603ec3e62de14970df4c6232eaaa6e0121914dfe785f11fb56e3e93d03bacb9fd
z3c065f8335bf71c41876f452210a756a750829b773949155b3cb725c1cbe43daf0df7517898cfb
zcef800948325789f512cb3bfb3296a4d2e5736407828287408dfaa39af63315a8d7c2cf8aef4e4
z477d29881809c71498ae5cf2b917ec5e2510ddc6cd2d22d58636a6c1a7ade5fb916c2f684beb83
z1691b50117f9917f3160be825462cec79243c2e28cc5a79be27cd5d25f5b3fe93d506877d1d836
zcb6912a8e062fbc957f036759ba2853c932c3837d71ce6467496537df81e967e16f3e28be43597
z21beba1cac9fd12dd50f24b0e181698e80177ea28149f67cf663e4051f6ef1560c959b32f4b489
zb7fa4f3e677dfe2f188047edd67539fe74f4abb8a951a8ea5900b4e06c06fce7528ade1f848d60
zd5a9f09538f4ad1f995bd378acd80ca183b589dea15b54e748dca912e193c84b270c612ff5c751
zf7a29c5a9a3bc805fa7dfdf7d5541338bf01ef20a440654add23df35a28dd144805cabf6cab0b8
z953c5093bfefcb14bdb5580d1e4697d71209953732c2f212eb16420cace5ba15b5cd2189fd94a5
z9b69bfb259f0d6a0e3dfc59c2a769e4b74559653eb4722deb1486daeb450346755b03dba18a4bb
z23c954ee7187eef9d0b26723e729456be59a14c733a4489bbc2d284ac13d2a3477baa5894f6056
zcabba99d0fe49805163f5457faf8e6fb0c10a1a5bcba067cbc51dd824c668e312b2b4d750afaf3
z0b040d7691300f64c5c3464e94409a0d8c40181a24f40ebe4882a6d57eda47f841bec873cea92e
z1e2ec4377f088eb989cccf32207d1215aa33ce68503084452894d5de1cd0ada581f829da2ed8af
z29c3a89ba4d9775b579622b3d506583975fe710eb5f205bd49368f4c8de422690714aa26eb7ec2
zc7d3db33d445db395e8db54700ea0938ab87629a96efd1779c0a9cade138a171538d66a696c605
zb3abfbc07310cbbf35e577f8dff568f2ca817a5c948373711ee314ab54154ede0fe0cc78a6fce4
za6ab8f3bafa4099b5d484fa9975f5a150023bdf220625ae85ffe31c58ef1baca4bc2092f05e382
z3c9216e01a9c2d415c04110c10e49db6d516ae194e4428a70855c538191a910152a277d14f69c3
z77232b86bbc6b19fbea0a66f8a5b9b86a7a68b91c9cb3e52ec222395f365714c10a43ed9f88879
z909c2625a534faaaec81ca3e5ee977ed39ec3c218b66be89e63017c05a2aaf01564e3bb43c939e
z08606671e9e8f04c9e8fb3f5f319992c03133ecd1a7808060d81c5159739e5f98b34ca845fcc6d
z5a49efda2194f5a3d5d406d0c6aef3f8adfa19d3db10c977ab4ce96f10fa149c88bcbfc83be408
z2617d2862c7d445a06095b1bd7019b2bb4a12f3e7d2f0227d218a6e373e86747ae0ab8c1f274b9
zf918d8aa4f79a04d9426978b8594f91e5057e62cacbaa48648c7669903f7e6ffdb89caaed57692
z443346a818c43e703468fb89cd8e8e56d36ec40006844c00132bbe5d772cc9284bee06921c8426
zcaf4d623d67c8a5582d1aaa3df3ebdd5ef16c0a1d62bbf240b89419ae2c98e3803dae3fad8212e
z3bd17f801eaff3c98854b5f0318922a73bf86092e4a77e55479aef1f7f7380a7cb0c9101dad1d9
zacdec17e9ff15af7eec8cec4f4f984f50160242b62dd4f1941250f047d5b06a44fc9ebe9ec437a
zafe1574f52798457d46040304838795e1b434824c4fbc4fa1ab554057ffce0d18e45f3bf5b4eb9
z5d00687b7302b6bd3a8bfef9e6417df7a78b23d8ac555fb17732d31fc6fb66653d56c96a8fb9ad
z17e6e40db9eab45c6829cefc0aac86a9375d1d10c03468d6288bdc90b45b6309773c910ce2816a
z8690065a0c45cd6a47dca17ef9bf81157ad6508ca245931ff4d8e31b92554c24dbacc2a07c0f6a
z7834e63758567ef38e2a820273d105b8776583e5480426406b9e3ba5e58a4f6363c2b483195060
zd0ca44c29b3ffb87c2ffaf762fb90417555a6c23917caa137e29f00d41e30e45d61927c682ad60
zab0e8c25e27a3e90dd4005f9a689c52e03e9dcebbf9ea5f1c5e1115caa2aab2182890145338090
ze15f247f96511c603f97ea3ba109de7d1b0ad321f5ad5756929db056b4f3775a7aa5387c69612c
zc7c08bf6f974b5bfa7fe264005b50b0f826834f962b82d624a4ca4d72468baaef6f04d7070a968
z75af8789f45778a3c47c38966587c9e0327f60303995654a7dea0e6c32edd1b8106d41c3e811a7
zb0244a589de1c2bacf034b10a7ca99b705c4785cf236555eaf98d84ef132c7261a8786ef7ce62f
zf411f04e53fd177993e4829a3e7af5b41318a2d9df0eeed1b53d1e64297536d6f898bea038b061
zcab11baec7a70926271f80d7d3279eed88208a1e4be75446e34e5517216bc15849b20d4126e1c1
z18e0d250a34f2b765e5bf1e421831d12a9e88bede7fa957e145762488ec0b1cf4b97ba46d2e74b
z4920bb56fccacf2b571aedf74caeaa96b62f9298a66043cacb74f78e95417783709de1295b80b7
zc77530f5cad4c793311459317cb6341e6ff6e349b7d00864346866ef6b1264f43642d2edbb1238
z1b66ea2dfb9e816566598efc23d8df24964222fb97154d055d15025c1868b0711aaa11997e9628
z5e37046ccf089f4d8907df2adbfb11c448f5532296a67d9907c958bcf5f57f672647b6788bec15
z8d47c2a2f0fd798ff2a45792064bfe517e65d7e5e4e006921769bb01d4c9705e4eaa047e1c4dc0
z7de9da599f4db52def04f876012c95274b8d5739f6e8d6182073e43e139f51bf0d5a3ca7b917e7
z74ffdd55342ad796caf43914cabc46fa9203513bbda9d3bf2413b32278fa26135a34cd636a4c37
z4f0bb7f4ad1eb1818bbae36c1feb75ef5401b17003334dc6726e50d6406ba513a65504113d5780
z5d3fa222c258913b3606fe82becd323f329d1182b2d5596f84ceb6762b766f3179fefd8064fbdc
zff0bcb87517b7dc6920eab4490bbff3c74de0f6258eec84cc934d26df205de73e468013f8673bb
zc95ebaa06394ecc3e3c3ec4977ac16f33e5d14bfcd194bc04f576210a26085eeab0838c3ab3fb9
z220f087021048ce85612d8523f3e938eb6ef2608a5b244da7636073777ec972b31777e06550e37
zd2dd8adab822b1e967de57c35cf4b39426106a1337e2fdffec08b412a588159803ea4a4ea77d23
ze72838dc23aee3afa56dd4279b3e908e523a3b1fb182a2f6343db53e5b1902d0128fa3c0cfdfcc
zf4a4973731a9e73a62004d5708950f7a36ebea8bcd476c51058aca49a1ca63622f4174c4437186
zb8f0e0c2aea16d575681a0b95a66848c68e0cf36da7ba5bb56cb040f329d2b4b7d3cb5989ca4ea
zd9e040b1d2d39f98346fc9317f3eadc93a1c41eea928b76797d5e7d4c41a750b72b7dc8c4d99fe
z7779c4519aa256bf775b413d577237b00de41990e2f9bd7712f94b94f830d06c6fc3c1250d9d8e
z86f9fbfc5cf1479ecddaa11000a576a28f6845d6e4951264b6b5d0f6705ff425bdbee5618caac5
zec1bb0e56ac14ec663f768e35d6a8393c1a9db2ae60240d25889510dfbb120187a6e0864b912f5
z0089e56cc21d4ead63582b512c5e89ca26cc4e2a874ef9663973045ebcf6bdff5d694fa3a716d5
zcbfca9eda67f897c73f318959cab76cbf4b7624cdfc49ded15a20ef60830517c398e65bdf76989
z2721f0b4433b47bc278b1e9a3b1c53c4031673e23e52e6a1c67b0f20d4b9e8198425acae739d6c
z6148035ddd97341e40431b1883aadc0d6386abe4c1a276bc47de943a2a45be14c4e9254c62602b
z49a5c8af41f2c603c6c88f1a5bc3e20e9b39db44421839949ad49c91808b53ec428d54bcaa7f16
z164630e054a5483e3a54fa317c985b4bf2a97bf3f75cd33d3bfccef7c8593d4865a78dda757996
zc3d078ee9600e93ab739b84aca4bd31d9b2afb384458a7a07720ad54d527cff1dc858d0c4b2c10
z929a0cc2ea83d7a19f8688b7cb0334f6418054805fffbeabe3e283617907d144af5b5f6b4d92f2
z86b66638f81ad331b8448cc319d475252188a92b6f55c1950aafd0383b45bdd32a9a52755a331a
z99f8bbc1cff80f9835af07962b87edc1853f59e5b48050514daaba0b3346cc0f9dc4756a9b8bb9
z69b3e5565281d4170445d4e0497ce2c9bf0d089b36ddbdff452f489bd8ef5f1d66ad4206df7e5c
ze20b67ec63173016fb7f65097d87c5ace44e99ea32f773c4db8378730c4154bfb6441115cd567c
z95bb6033579718405709e2d8121508722539075ac0541c9fd146b539f9ef2ae3e55950b5b7b160
zf2df4b2f7a135dfff7f93f7ac66d4d468a05a434f958edaae01415da143ddbea585b0ad94e9c78
z1ff37e8471e5705f6d6b8fd67799ea11c00b63400bb41e7c96fc99b7386ad7a084f864ef584f2f
zf49a82ee62d9cbdb9970fecb52d806d0b10e8a88aa28d7f08b8c96d374bcbcad7388ca3f388de8
z78c6a95c1350cf66dce4b5d6371367221a15ff87bb99a95f89e0c1fd6f4d065b1b1575462e5ae2
z8726a9547a247e6a48c731263fff919472a41c22db77c00ea6be3c4350db6a43b0446abb6d6147
zb931404e6603a1d7843107f3924b9c35fbb81eab733106f46f51c83ba8983bfbd8caa2e415ee7c
z0c08e80f2e32eb99533b6aad08f72a5c7e983faf74dc171b7069f6d26841370f2d88a250a6ba8d
z2b9db0cfcc69d332ff160df6b947cb1dd873ec1b8e33f2f2b39f05f22c0f532e4eff1c582c1dfd
z05c13d9b9691ab6b59d51798a95047b1e743281e6221fca6a19b67c8906d0c71d8d50738f9d784
z3046ff06c8a558dcaf178b904cbb0f21e0904721a0c3afdae8a2f5497aa9c903d7cfdaf67eb272
z7fc7fd0af64dcd70bf204d3617524f208b8e92f6758fc2a3657f5174ff52ad033be61b8f8e2fdc
za810cb7efa8b2208534110943f52ed27446980ce8a417d4cfd1462b2be83f5e8d790035c6c79c2
z89693e8508649844cbe73e85928b19f60b15281bd75491613aa0859c231dabc9758d4bc86aa486
z2e502bba3f52e127b28eaa136ab98419a05a88ae86770f916aceb704e99d13b00e17ab3e40b85c
zee6d7b4d6cfae496a960e87a736be88e2c122238d69fb65dd3f9771ee6ab09f5b2b77b23de60ca
z25380f6be750d6211ddf8da1d856c6013a0fcfbbcb6c6cce3134df3ee6036c2303a13862ca1886
zde6df2588dcbd15d2fd5a0c8b900df373cda97fbe50478a996b2fbdaee4925cc9e049c950bc59b
zdf4e6e30e340670d3a1d260be0b7d180bcd0d701a3fc0ed057fa8984efc82d826876b2b6e68dfd
zc670af5d7723f3268c576ac32b67f0ef3f9fafce183b0b02f09da19a78eca8e39bc8b13efd7e77
z9d2e4548156ed5efe2a0545d663a82539511262aa368aa381d2e0e6a27d3c6f13eaa4a1301ce01
z2bb28e69f9e02aaea199d8082517d3eb8d46cb995a7ce0b5725b19d9676ebc0187a17088176fae
zc41a4c655926b2d44116ad9bae23d290c989da4b698028693b4b5b4b7a794df309dd4cf7dd3d51
zd9c99e69f32cce4c144ef791421c1ac7ab2aef384544dd693feb4aaa7dd75e93f02ad87dc42609
z85e9c0b60f1845ced96bc2cafc7c1206e3a1cbf3a2727be4e4122ad72743dc43467c88989e2b2c
za88ce67b53ba22bb83d88be5e5b9e46e5fde71d9ad4a0254df042e3af9b63be9e465f36e4953eb
ze32f7370e6dc313e1c75757022510f43b816e3a595afa4d0c2fbaf1f9d8ca4cb934291b8aefd30
z22f4cf77579e4e59f25d9a13c6d03b17f89a98d2d33ba23a860d28d7b8278d2dea1182701ca90c
z2b3db704018eb6f4f235fcb88335e996347a623d71bc7caef89cf47d670b117ea5a6816a0057cc
zeeee0e4ab61d803fb4e22621c7a9827ceaef318e6c8d109ba81bf1e08d7834e92ca8b301d89f97
zc0af79bbb78cee1243b9e0f580f58a7c780c600d3f87babf9d0e8e7e242b836204176b453db806
zc0d7ea5ef901053f05460b03d94601851e82af82a2f482e241b56822c4bf738fcf55de0d6a7eda
z59b118539abf3e72a7471c5ffcdfa7ce0d67ad17237c962797dfc980d3afbd7a5c8bfc56d0032d
zcd067f56a740903b254a3ac606728f53082c52a5571a9a9d9ae5ab8c1544d3e199c620a7918127
z71c7cedf122bf0ee111fd4ce4babf99f4e248de65ad94aee555cfdf6022b5fad94716dd816baa4
zeb5a3488e87f24113262ba342e2087265ebe5133c9619ebdbd012a1759e138de9cd56f2a2b670e
z2304e6e64c1b721c9a121476afa4ea7d012ddc516463daff677dc1cbea83b839ca74dc04144d62
z87bd7248901db9be18036850f4c88bff02f95ed95c517243b391b0ab62655ae4096f0b5728f34a
z98e41711cf6a632a8a9454694373ee3937646993c025447de69755f55eed6f2d34077a99def881
z77a6819375eef580c017d28ee90b85c4b7a1409cff27ada56fcfbf9a488357c4d7a1b65e7fd0cc
zfdf4ac7246c71044e231544b5a0538923770dbedb34dac8cbb644f67c7441ca0db9d726da1aa1d
z5c02efca4c2bf79f0e523003f168af2d8f14aa2e90ee34b6e42dfaa339fe3d5b0fc9333f8813e1
zd9c3fbbf1f1e21680976532ea7cf7d117cdfbc1cfda0a12e10d231561255255162c36dd85d1bdd
zefacd46de0e4d6e0ccdd585d338e70a72e47f61bf0d75919fce377205f2eeecf75e7908c8407ad
z964ae5ddf2d51789e981ef82ee6152fb3f16ef85b86d9a4897d04e5e05ba687b06903fe4fb42ee
zb1852d59ab1efc6d2afe6cd6f422251148ef45a4a5a727aa2e1dcfd4c566e687430c85529186b9
z4e4ae0608a302af5a9b7ec5f1d56306565fc6e0ee45f4510404c748f458196325a341427b608b7
z0e519d6c74b752e0f50c01d7d1f803df3a9b2a598e5fb72a0a50539d82aedadcf043ffb03159f2
z7e9a7823682e95bdba39876c0d506be3f6feacd13f89a244e4b4f6c1b1a56b3dc30af6c2e6996c
z09069cdee2faf515674bce741fda8c0741335845c9159463d6e5802d550b7cbbfb720b0e67783c
zf7824579df7381097b364ee333d796098911db7e25ac1df40f6fe339efc8095adb5b8ee2677c99
z95ad2823952ff9e3c416f513b33face8bdc229df397c40ca4f46519fc32cc79fd04351be9bc47f
z6d625e7433bfd330dec1421ceefaa8ae872517177634d363a0521acc24e85e610564a8d67227c9
z456d686da59be9e64f30169106c058dc4f66c8604eb1d0c2f532ab2ecc82bc8f190e6d01525943
z3a5840d3871551f4b5a971cd4a0936971d56a519673297e0a472b3a9b6ca7aa9dc0e105fff20a3
z026169c9524d2705b80d92bbcee5e013678146bc47e3cfaf1abab21ccb6947ab7701a5dd51f2aa
zebf56b97898fc28ba80f627558c97ee90f1214377bcb8a3ee8c31616ea0ed165cf2941584c1b9c
z96fb0277c9e0590bb5f2f650c6092bbd68ec8f465e7e4c71430dd73c6890439ee6529132f61b47
z6a2cc0f041f277b2a4e7310ca495b6c68ab9f2f90c143b23f0612b3600d6806e493c1c39139608
z078ccd9434b193f6cedb604c93ff1129b27f5a9b03c8566f2baed8cf0e944917468dfd24be4818
z14ad3b78ffdc0966b26fd1ede139cbeb967edb4cb0d5f868b0ad5fa6013076989752d956a3d292
z69f1de3b66fc520b84987d12fe5273d1e97a6ef6397460de990bad4d362f1215f4225a88126c5f
z8ce678cb189622df2c20e0c578ab5dca9a5faae0f7ef0f8d47a88b68e2e7ab3137f5f999234198
z4f0570757b0df4de40c56e9e80bb9ef4b775cdbacd099c7ec6739ad6b7e52ab52880a29ebc3686
z89724e3cd39ee0ad0dcb560b2246c0663cef9594e6d363bed704d8756572551fecd8b072c37a1c
zda38f3f7037ea3c882d2b5dca06d1acf1982b32bce7f80f2376cfa73f01215fda919b831c0c4ed
zeab29e5fbcc7f9c0fb2152b2a951858a3b3a944a2e0a2bfb94f2631b05e6604ff922dcffb259d3
zd0bddfcd29807de456b8f07a5b9382003b43641f301ab2ec641ef61510837745bf20afe0e097dc
zee4b82fd5033c9f08220113bce72f504c422490215d705c8b1633b50430ad0d44c8dfaf02d39fd
z22123f0c15c2823173d60c7a6a2c9329917275f4df95cddfb4fc0285d224ceaa560f13093526c4
z81a205ee92cf6b7b07b08704e26841317edd8ec030ef640dc8005e6bde15a0b41f1a8f1fb40795
z7982e78de1b1bcb18a5aa064152d7cf215f299d55c5bdbe6f69f8ed8c2fb9218c58aebf9aff27d
zc06eb3ee6f5e0143c201c87a06ff10a2437a87c9b6125a87010093018d407d4e27d18f83394f1d
z75f1b317e783a2fe891b2aea34bfe976bd1294094599529af32a535d3a63ef51e330f21f427beb
zef529e4babde5c153b4a8b3c3021eccc6a2609666e306c8dbdea0c8ceb876c6cba6793208bbbb2
zc74a889a287783ff2727bc198c13ea0c28536c2cbcc0e7e8ff3878ceb76034d2d87674f3b912b3
z9d4298f0e9cb09e5e0575b7fb9aed018a356f6e207c46f574fbdd582f2271417716143394573b6
zfbbe380fe9496ecf790471c0be768c9881be956050a3d94d2bbaab34b6befede8c3e3d500d9e0e
z1f8552415dcb9d970257ecd091c6c87559f42af5dd31b506bd69d8e53ac8af419d9b795647c849
zdd495886df66b89e6b0a6dc25ccddcabcada2f9043aeeac81caf89a2b7e0a56693bf483031af94
z0f446316340a669c943b74b6f0767a8330182c3f59d55e7ab55e03e1b4f1b04c28cdef529ee47a
z6f2cc4b12267710dbbe4aaa0fe46444a467484561788c9c71a06033f3328469a1d99eaa5030e7c
z9ca9c28a097f596a5babf1459bf981a9601585b9c596ec4e083dfdcb74837ab57c45ad805facea
zf2eba605936dc1326958942818026ca97dbc463814fedb052f1c8323e55e2d2249ca9df21bb2db
zcc6c2ab4211e03e5354366b442f8b620287f0fbe7b0e511e8155d0d80014e144d3922196fdfb0d
zed1689d5f0d71246c1b1dead73b4a6cc6cdae15a7d9ba690e7cca52e2e7f1cd0a62494b39d9e72
z64e7d74aca92caecc8c5edb6f5ce4e87ed0ca272980dde5f7aa7d8cdb21bf1e6e7a37e56034b4d
zf51009977c8608ee8b1729852f92a809d6fb2a12945ed143c129f1cca768d5c77b5cf96902b108
ze31b2c7ceb26353b4835f0001af69f022a075cb7706c11a21011ceb8f22bee2f7c5e570542630d
z281fe098829d8c9514764f7f8f82b90e91560d6ffeaf89a9aa888bb1f2dc58be2465c61ba1b108
z9d51c48b214954530462fadbb5f22c1d6666b3e693a6d77edd761b5abfd984181443c65a84ec18
zee682dccfcd513e1124489d48133ee73a43cdce6b5a460700666cdd75989a8aedc9af4a3cb2780
z9a73930df00b644bff2b3c81ea92b4d8f0fbe573e998e3a6684103abda0400b0f1eed8d229ebbd
z1d36a7ccafd7ad6cedc1392f3f191511ae154ecda4b1c4fc1ccdf405b47f953c2eefe39e1f5083
z91bdbfe655cfe38c07531dece5ada5365c2f212b2b7814b1241267aac55f17eadadfddeeb8d7d8
ze41ce9ab2cdb296be24e2433bff9959d8b069fe9a0ff2eb0f0c5452d62f1b2d373d0edd8300425
z4245bd2933e66299a746b59f1a930ce773322fb7c4430440943b0c416e5abc70d5ce762c106403
z698d8cde49be007b05650cff432164b93aa11dd2ec7168edab307beda92c3122821279af8aff1d
z33b1e7275d9245565b3c40ac46c08cedc2ff6cd263501a87bd6921ef19e2d97619ba978ec4f414
z80c2fbc560f961e86fa66deff790990b686d18ab2e580501c2f0a231855a189c229af0a1816948
za240ee96b40ae5461e842e45ceb91df9f0e9e3bcbef58dd10b3a544f05bdd856dca8635b981f5b
z3f0a0e468a517284be885e917916dff2d225b37063b6a2361e972df15efa1e7936381800d0a967
z16a0d5ac07b8fb29253009c840936bd2fba46d2d83d928d71a12ef0449e97a5a91c9a71e6a57f5
zbb3bf2e550d62ea56aaba0be6093a42bc1c92e1bf82c35f95e0f4a088156703c10592ccbc43999
zd980745e6782d09890427ca69e9e7edc4694b51a74a7e5e5c71bbd59fa8f372dfbd1fe4d2fef99
z6b824c052b79a32d9a0ea996698e1c8dabcba1522d98ff5d903fc29e8d85046b6caafdb9d60f46
zd33e15518db382a8117e8172f24812b9c858c2228716d3cc8a312e66ec459f655a4deaeb785d8b
zfca925ae59b79cf997e95af08f5dafc6e519ad0e9cd77a5a7ca1314a41aeafa88ca59de9faf13e
z8a5ac4b399d08ad30271c5d393449fcc5467fa81da1ca151f435dac61ba045f19e06a77ec77db4
z33db7f2cf3ea09fc0fb6cbd5387e53dc0051ebfc82bcc6b70f910491cca00b38b3e97f2c5e3d16
z550e8222178c707079097925f82b089d3e87273af4bfb18f47ed14941b539b70cf723e4fbdbf86
z515ec6892e00d74db0bee34ae3118c32d362ed522d0872d116831ab810e7f715cbaaa59dccc627
z6943457eaed79ab49b9cf1471fa959892a9ef9aae8be9aaa4bafab3dd5f0d868461f5a25084357
zdd3ccf4768f1738e6a6c53d43c98f1c5a2c66d43dd79d55dd25c1f4aabf4d8a1fe06ab0b77947d
z254f1fa02fc448eeea57532e2fd18fe1aabb2cb701db1fff0f40527d5183852987ccbdecbfda7d
z6e6399e16aec4f3cacd198aa7520304375e8ab858e056d7e11a253880a648c27d32d6f1cfc275a
z3b07352ddc66a41ae952c1a36819fb6ed5c13127b5de70b59b131f5e5fd0500c34ae2f5d99da7a
zc79ed85cf7d04a015eb6e11bafa4b5ff784880ab57d02279c88b486f6fad351830011eab506b3f
z89cd271d39b5650a0db5eb7dae22c1a9650aa81fd044699f8276ee1999e365d589200fa7a0bbb7
zf761ed5727ace6af0c45d5556d152e8aa201e5d1245c20c9f5872aa3b90efa50ee80eb2d14fc5a
z5c6c93faf0b93267a56aa97a5539bfdd6c150e285df1bf6b1a4b72d863861d7b17f89a2e9ea7b9
z5e79de129ed7eeb18cb912a9c01a7531c26f9a4a1b16aea0f686433cda5bb52a5c996eb2a7088e
z1f9dfebf1c0c384c5c5c67dc0b75a81af3299e7036aa88a56c48b52d27374f66774efb148378e1
zbe9605ef1292f668acc20c75137d6fb07b7fa1a4ab1542b4f20bb782444d8455387ccda8820341
z8e8c70232e1b09ec600908ba1683d7f5da7f0c46c50c8fbc49b3dcb594957814b676801d35553b
z5456c3863e255b1554a8af93f819b29df61172b13b0c4f3a215ae14246ab5883e233a93c58f98a
za1c4c817cb2417423576e6a398ff96e5e5b03d5b48cdb50d4c26be9ce40ef59c2f787e089533e5
z8649eebd6bc5202c3a0d4d50908c603e1253d47eebf7cc7a4a74f4e30514d246e461a96664d68e
z995d58f8c5c30fe743ae10e09d3225f17dcccd190e0bad46ce6e90a1904de416545e54ad6aa4b7
z254850586ceb0183df6c2c1ce80d11bf077e10193fce08f6b1fc165cb809a5266f4e5b59e9aa30
z632a1108e278e8c06d76dae914f8bb0fc856e9dd748065f643d3a750c5b84f43a2b89ecc34849d
z2de2e22590e1a417366c229bd90398406b48b3a7e5855371829bc2bd6785beaefbbad308f96a44
z4d7fe5c7326634606000762c178a40e5513ab160550579000efbe54e51ecc27126594b2f150638
zdbf26d69e458d8a48472f3d3482fc8c7c36738edc8928ea77e1c7128b46204ea366607131f413c
z1492e05e612966b9c8cd62a500d36bdb5f91bd49810586042eac6fabed08e27fe7b40fd932f3e8
zc3f03cc76dd1e7823a9f9c43869936c3954373d3b92f6a7294bfd2f063e561b5f9466a9fc096e6
zba88a545a670300dec7c5b094506f7cb64ac4f3e9183ebd5c2814d7688d6b99c5b7219b04c747a
z8db8630bbaf5764d312d6a3eccd5516efdd515eeb9e9537182351e21fce81808f4c69afc2680c9
z491bbdc793e05876e7765b7dbf39e2eeb238fcbe9770ab7b076ecd9f839e79d8c3a2d4dfe8c3be
z2946a297391688295cc074f0cd9a5bc8273c29a8f4e7bf9e67a2720d75db79f471cf91ff3f4b67
zc91b790aed1f99098f452a14e1d143fb80bd6dfe3efb2c762acda38022b6e0b62ac13aa02eec6b
za15ff1eecf8793344bceb791f47c132696b27d500c32eb16294a0efefc822086d85b33b369bb99
ze3482edd5d724d5df0fc5387d113dd27ac22e96a39a97f3e4b8eee69f57a9f4a1d946f74c70609
ze277058333ae3bcfebec26c23e30d16f6478ee6d673502b921356f689cf97b5d7236b878d7e343
z8c9be879d0724fb569283b6a68af14567726747b37d88f7d4d6a2010e7e62d490aa90481eb18c1
z62404696a3916bb580ca00e278c05e278d7ff65627a9505e9c6bebf5ff7ba6f070679351bab76b
z5ab453c03b575a84e47ef805b346c09229cac7aba7d88f1dc16c56c6c9e36c3bdd4b7ed3d8ce0d
zd9cafa8288045970173b6baf0a1770ced9ee2ffa7bded50400e5f831a90cb87ac548b27ceb92b2
zde4f656cf817f8eba6fa80a1dcab46ab86ab08a783d5807befa9ec69c44cfbe23adfc9a62fdfbb
z1f8a7606385bcd607ea88df9cdb91dd4b35b9b3f2a60529978107e22f1b64125a292e533538c60
zae5ebb21c49dcf34e4a56d47a32ff655ffb113c2897c87d0cbbdf56c454b5190b6b22464d297d5
z0f77357d0d7a8b5314708354932e8785d402f9ee7c1e4b8ee982457405a4ecfad62d3c73af4237
zfbda9624a51d1b79d0c82cc100b44f143fcb3ebd17182c291f11cda0d8b00c72fbfa434a213e5b
z4bc2dac0b5cf3867aac43d597723f7ee06816191d4dc02d62de883ecbd1b2b81963f889b096476
z1eacb6ffc797d25f90efa1d933094da675ce158a99d4c4c562625c3b54ab7baa724e7435ed38a2
z87d6504179b0e25c81925b2686fe2f577606bcb277a6fee8a947ccf5c2c0fb556ee4becf8457f6
z603c4f57d6358fee091ba6f82081d13330f882e9917c1d1d91db2f2d6cc581646d10ce28791b89
zb3b165eef0c8aacdd8cf87d8f97637b9114a26af0dd04ac2358fc7a453a8ac4bde25ff2eaccd17
zcba8fe6aeef0bdd94ec449fa658498cddf64e3e647ed821630e05f0eb05b88dc5de2d50e9d170b
zc736ad8540ea54a12860c3b61e243bdfa34e1be8ad79132f783d88690bd48f2299d06d4aae52a1
za26ebbc93b47a6f48e1a668e657c893efe60a2ecd1d4a40d9bab72e09a833c760a7a88480d131b
zc364a9fb475713d9e2236fa876bb6107e720f243f867446a493b50f434221b423256efa8058a68
zae6fe8cbcb6d78441f324f01764528f697879218c9533f849e3505c2aeab6e0aec6e2a9379add3
z132cb9ed7490a8ed01dfa315de537c04855bc7eef74528e9ea85ce02eca524dba59fca6f702112
z2a378e00cbc4dc51bed498401e2dd01d39d19a0e2696709edfcc12d6de947b0173b8b3077a1e87
z5f2899c887b9803ea998e67ed9250cee3873518cb35ff2da4c29db44754cf2cbbc842d240ae769
z5661c9f50acb8befee4177bef0452959b8c951037f82f10a499d19af67481bb9d4d241a73bdf32
z1b3721b033d98045db65117bfc3388a0a10fccd698eba015dd0d35fd3bf3a5dc3a414054828ba3
z92e9d5ad8da0d5e9e955c01f6a424469552333200a14eddd3d1b2e907baa04d836f49235307035
z2763def839871fca3733affe82a4f899131b96e456a730af77bc0383e9b01e409d0a5eae9cbcc4
z9a6c0510160bce47ee4598b6a09542562da276cf1820d669634e796c40aa57f93cfa2bf2899d4f
zf7cd900de6862ce237c813b1b79ab9d30ebde6af1c71089d6be4edd1234668fe9280565eec269b
z9cdac1bf30147c14ff5a88fd5e6aa6f4cd592c8efe9df8bb0c0df0d3c798ee958bc02c35ffedd4
z25d94e07f2c9db9f724ce2f2bab058b6a9683c70c9e10629513fe51c473757de6d08d3cbb06cbd
zd64157ae6b94be08254d4fda24ab3279199726b0c4642e750efa146f16a87d7c38bfe70bcc42b4
z91e2790e8fcf15fec19ba1d6747b680676644aa62c3e383c92479a1600054c51acf194f7b5d61b
z0eab27875ce600a69b297ff0761da09d8c3f0a6a2a7cb1ce8e4d42b011ee0d0dd5417e1f5cac6c
zd5095fd328a3e250effd7eee25416e28df592690ce1e7b74ae8f400bd3aed7392e60a2af6e809b
za98c57e2da6b314a4b39f7b3b5edd00dc79f4950a5421d43ec39e6d4d1caec92fa872123ef31d5
z1a0cebd7f25359b138c397b2c1c1de545c882a25fa25bcc4f10a26485d574327127c3f311792a5
z284bd8a564ecc923353c366dca34bab40275c91dff1fb9a1bd7c5e235480e60e240e663a37022a
ze4d49b8e6be8fb75df88bc8cfc81fca3f7c2233190cff542a5a0a04e0d2028df16639effd45037
z0ff2299b1573b86cc19c23b47be92d326494416bcdd6e196362412860429ffbf0330b98bc5e27c
zaae3a3349ebecba769bbafa1676e455be3c3b999f18aa7810d8b8189e08d0e0b35d8bbb32389d1
z7b3f33c5dc11310c78ac24bd59f10efe69338bd26ffc434cbc7ff9c4e0895b1aee723a6f4f0fea
zb0b0f8df59153bf96772371b6887dbb86447cbdce0f6f71d1f736b9f273d81bbb273e8a822483c
z469482191ba7aabcc6486a3b8c96d472f25614b4f94c9d2f065c0f5fcf06bfbcfa8456cd29746d
z3d1ecbbe3e584e9b5da4a997fc1b3de7f07b42deca5ea1429ad8a56ae9b1ae1e7cce4e4c00014c
zfbe46d52a1944d43de70870781f19b1b054c230b21b484b32b06a3612472894902c7f16324df81
zb8a274e73a9759914ae66e353a60213cfdeb73f8521a8465d5e8a83d414a14d979b7804819704a
z1b782aed8e2c49c71af80966a3e7e9cdf3adc3de31e61797af47043024fdc527305f75bec61e6f
zfd3769c76f71f694817132a84a8079d5fb6098f582a314de3a33639ab42557183915ccf1a61714
z78a5b33c00a83f8497ebe677fdc0dd61952ef56fd5dcfed1d8323af43d57d94a1fdbde8f446d81
z15892d4360adcd5ab44a2a88b1dd442f66b0bed316c6bfe1e21da7276e09f96ba67dc645a9d49a
zd2b987dcceccb9bac252bffabfd64d3aba86febcd61ef753ea445d3fed68b9436e73ed638cfa92
zbb0786ba376ff4451bcd2ec256211b492b94b57938ff55586eff6ac5a47aad8e035f9ac0e893ba
z4c19c0630d947e3f3070ebd035341bb500eef116dd743dbac6eb7a7de3e124b3c723e2feb3275e
z522c6cfe1566c7f65c00da71b0cec2cc402206fb5c3f9f6f3b9e09700a0beca310676fe1f933dd
z7e23ce0696d71775c4003eaf49da569f3d1a2f9846fcaba89641d4d2c1ca514617648bb93194e6
z13d3418970734396f2c4ca8514a2da351402344f00207083b103aacb1e6a9c687989b420fb8660
zceda69450118bd065c1e7602bbbdb8051dbd30c44be1584410bbdd1f5254998ca17e3f6356593e
z7cd55045769ba044085b2bb080410de1d0721409864636c3d195e39ec79e073ac9910e0ce2fd9d
ze1a3dc84f845a545cd874858c5dad34487ffe511cd3ddea84e1a3a04bb8fce2edfc84b853443df
zb36f1965d0fcfc1cac8ae184cf3beb6b71f9e613dcf9262909a15929c74ed454d35835a615d9e5
z180b1c51ff86d591d0c0df43cc216d1e3f3206e8631f8e578a45d72941beeaa8e72c1c2db825fd
z7c9139ed074fa28b679649402d2d4ec7c344dc8e3766d898ca1b22618219f45fa12d4d5df4ea49
z7a4c53b597d947752fee1850ddf62429c6944fe6613417d0e053abad903084826bca0a7985baf1
zbc7d26faf46825cf9ba8028911b0543a9c858b2f013b03d7f6662fcf00add537d7c3447db66015
z99689c860388a12f8faa2a624dc17fbb6bef3fdc6ec612cde946cb97813f07516a73e68a979beb
zdedf84ce0d49ca48df6bfe62258a2e59599822a06530adaa6e9b3d2c8ff62fd9bd628cc6e3f38f
zc0d4d56603780982026adfa87da57cefb72ea67d1250642c2534aaeeea8ac1ae0bcdbafcb0c9a5
z79aba80de96a805a40a580b891538f293b77a5c88229c9d4a2863682c551240903ce2dc15a2105
z6a3206b08031a1da54059bf20fff4c0eb86585fe6808e4cfd89eb51087a282f71efe5cfdcb556d
zbda2b93159335094bde1425df37f39d91006209a80bc92f487146fbd45dc5f41986aed555d66ee
z07b583e285fd54c440b581a487747ce354b3bd076a091479e843ea0732b11b447a7a34463a33cf
zc6d0955b196d58158d73b025e480d8a6ff1787df2a01b6617370e47d766bdc9db16e4f63a4caed
z9a3e77da6809134c58a7eaa8d0e3dbefa406b9919b7d403ee289e31260f2bf450f0ad7c4a8544d
z9fe14398001b8f44901019fcc9247bc3ea627e0920c967682ebd7025dba5586e8eb5da8298803d
z499dc6078033a37d418ea65e3eae3914300d654c9b510cf6328340569d4e50fdb8ba07c1b11c6e
z6ff27514ef775c597f9a89b4e8d3377f213ef2afd47bf271364220b044f55e28335544c231f462
z7cacdba7860ae45fb27052b22eb00fdfb795c146715da1fe703fadcf9bbfca5d5d02c86d2ec634
za2f2578d0d9f4b49147f0f885c7a97007be5c81635c0b04e5d0780a1b990eecfde6fe641026926
zd34008f866ac61ff3aae71ec92d29ca9e4fe0a01f999391a75e25a92ac983955266c5707315948
z8b04746bfa7a9bab721c834aebef875fde9bf470da1ec826f470b5ec1a1ed26c3e916fde889613
zb2aab2da39993296cd73a7e1d2c965e8ac1df1e890e252bd052efc015c829b3e9d3ddbbd9247fd
z7235617b5759d0bfcaa8739ba7118f4aed9216f283aaaba2d00b1d25fce5fca2d46ab6977895ec
z887ba6cb8415d008e2ffa3b6fe19ac57006a050582607a741fb83698f0870d6c1dbc325dafd781
z1d9f7d9f70eb11547c4649c7dc836d61daeed1375d8ec975391af2193921f13c33751636d7df9e
z64335de197c13cc89d661aafd5b113e2ed42887141f0e900007617382e47ac8436d9bb7dc29c6d
z24c38e5bc35cc69abb905a1cd62fa829cf89266d7e057720cf6735c6739de402de60a43bd23f8e
zb81038549e9f46398a6730519a4ca21b6672986959209f983f9e86195046cb8abb1bb3e0e33e7a
z1940e59af8043598a553f193ed48ccc8af92770b7f20c372664ce0945b25b229f168e55efe887f
z28f0a2e8bf30f8e7be10b86f0ef1b6aea91f91afa2a460f0346bed233e9b23935d1d955a1feda8
z57f86ea6f2ea8fa6fca5514e6ab389ca682da1f9e8c17e20a24f8aefcf8b81c032d76d86df1594
z587e10b19351985533673d57efb2f95eb73c068c1a50e46d77f07b13fa9e0fb228f6e16fbd61ed
zc13ad16439a90e308d0477df12e981116ff9731ad319e4ef67ff8e6aad84c771ba8dbffc1a2ca5
zd6b347d717dbfcce2185aaecf4c42abe237cd4f22ec98597b37119612668529c19169ceae7e542
zc73f8682fdc713a517005fdbc03e879bfdfdf48c4b4b6a2cc8b88a607201f3b61ee610ab2035ec
z927cd27a2f1b1f34610625da53e815cc6034dafeb2bb295fc75db39cd2358a3ffeaca87e75f30b
z62718a7043cc0f727f91c987c6571ad08f4b12bea33927f80322ca8760d1e6b860f02b61210f4a
z174e6501b670c35ead47a7431b0820cb60bfd618e3120c13c495ed77a7feba921565b3a50e056d
zab98237c657e5cdf17f1935eb2772c2406670c349998c98bba72b672c2fa0eef01f63f19593e4f
z8db8fc1bfc32b6fcce0ecacde4f74a6d17f90abfa1e7d38887e1ae00ee18efadb972493561c897
zb3d435748c3b4a051a1ba62948cd6b2df79283fe7858b80452a021773a6bfe57dd2337b92cd51c
z25c08f3ca5125712a25964bbdf1071012ae5311b37142a7ccdfa19a62548d1670672c57d12e090
z8ba1f94a8dde469311beaffa683a69c04abd1109262388278004e8ef35542e2ceb1953a8b0193b
z40f54cfd078e79417b7e0f402c19bbfef030126a09daaf0168ecbd814f8a5cc1e0c514882c5296
z39d47c684b239eaa311666168ec313f7c23b93b8e7e9e8354728d5e2ca5065d80012511908121a
z202ecfe81789589b0485740b73a0b59c377e8e21605f77a756f533735fbfe0f5eb1778ac207b9a
zb5c36cdfd6476aa47d0cbf41035584c02df8f781f880c1417d2c1e811a27ef745f6836640f11bd
z7bcf08bda02ec3e104aa8a4f1c29f55d679b632f61e2753f30f151e186406b2ed1945ca76d1164
ze133df0e2cecf4242943d5faf21b6122742f274936e3b6a38114560e29d37c16626e6e28376f3c
z2a4edc3311869ee66ff94ec217fb28eee18f41e270236fe4b2de23515cf4344ae7b1820a4e47db
z028004c311593849fe3a9998eb7dc1b74ee347b1e1e955f0dfe7596bdbe8b5d95c99a6d72aa8e8
zc8b8fe5752a845dc03cc0e8532d0b2aa52d72263d8ba23955ac53cc84a1f7f5e0681405969d71a
ze90450e5f84fe13ac96903809bb5db31bac46547ec86dfc4e53a898061edda7f0df4aba7921f76
z3e7618578f016838ac3243ace170813610df6bf85e1f7a561f234a8c272f133f86ca5b8778a295
z4f6562341639b8f0d9abb3cff158b2e33c899e5d437a34d09e9f639a71f67346b8f6ec3d098a93
z7bf40ca8d6d8408b8c60d2f7fc64f10eae15569c01016a8b227004ab67fd3c0e07036013886f4f
z98c95921b8db20951620a2262e93e37c135e32904d62c73d886d3ebce2312a4047c14a1f99271b
z6622cd6ea8d8b2082bdf9704a45ff0dedfccb1131be4b4b15589600f4b3ada7f252f03d8c51244
z213eccc3e88ed2528b5a4e94976c03058ba5a8939d0b6cc09f27c7e852dd1baaf0e6bc405af832
z244f860b2886a73dbf15f02f58fe26594f911ac459a110ff650e30438fcf4903789f091eecdde0
z3cd0594221a61800596f1b189efa776afd02a76e9cf0f0e572c6f557d669a57b4ccba49d3089c1
z68695ff6b6369e930203ffae16c517bb11f51a6f08f820bd05068822b647451e41b795c0dcc839
z06dff1c675c0fd2a2998f017174550e9c1ec7cac0328f27fa4d19ba0f6605780acb4de3ac32cdd
zd9c4f8f049ddd86c2e2062ac870c96c1b5b51c05d52ececb7c34ea85e388d6ece3872477377dd0
z36ebb540bc3455fd5596a15788e65ecd0261492517959e25b3c15e2a4ce280bb1ca06d24168f09
z607102c54984fc2ed02d924629dd3961eca453631dda82fc76fb009892946cad1f22d867515041
zff8ae84d7dbd569b09409e8d10b7cb87d1575a5ec48ba632176bc3b4a23e9de6a5a4e89fd1ffe2
zf33333a22feb8c2a3a8658b592943f7596c6e1494391f8167575ddd02318c99f6d4fd48bc7f710
z3b3e5b74d822f60bf2a57c991aa6d6e715e066a64998749fa76f5f1a18b75d949ae85780f2304d
z47c566df5c0f299a826f9ca1a57e70d38672ce2e95f004974c49f4a7f19c5263d4e3a5aed34db6
z7d4417147e157cd24d6ddb48493ecbf02666648a0149be5401af039811a3eba77a8c96d8651a07
zcd893e958def61fac5207ec6991af43f091b36b36ad6f44d0add7a63d81ecc18537c5105d9d9d4
z0db1c31cbd2a0c0dcb14a70a12bf9378cf4990231fef00e4b81d551f01e212991b88bab90a44cf
z99c10369befa13127c1b3b842f6990b556f14497896f3f58a9021ea8336469c448416155267f02
ze128b512f6eb85a3e254080a6bc82e7478e388022d6200c23881d758da1b9c085ed13c90de8c9f
z6b8ff1f60d30f1a3464377ddc05a992c57304cb29a94ebcc7cda5e0e2108793b5af86a7e3b21ce
z8eaad3df9a2c30b4ac51d2f4b4ebd0af5b8394f5c1687c706e7736a95e5b50a52e2051674a4318
zbfaf3593ef69acc1778780941240048176e557b711fc323f29fbee643d237c1ac661cfef28a7c9
z43e76c01ae7613fd015be81d6058bcc3d333e1fb9597d4a002da00eb58b6457b40b4d37b3f80bb
ze26179f086ab4e223d5d1fa038515210f2fe7d3a5a4f314dac5cd7cae9d8d8fc094a165f13a4d2
zf8ac583cc4dc9dd21f7fa0220b347d9caf742c03026a0e9a82a0413551d05185d84404cdd203c3
z4f33795a855b828882606ff9221ac78ff37b03cc8f989ab0351a23f08d7532e4de4fa0391f9128
zc6859562083b2ee61fd79b68e7c8db95e614729c9ccea1c26bc508325cafb6f3add2d356daf493
z79560d7b62ee401cfe08c7bdf7b057e8bd33af5113f043ce393d1b865a256edb25d930d90c2f4e
z6e2c167abfd8d219672eb030aafd3ad89c7f7e04b9430c77ad75cf2dc93034c47a27296b331b7f
ze54b89d874958c8086fbd920e51a26ceb32a775f30c2f4c3b9f5bd1e66a29020ce758242a787e5
z808a27673839552da6cb86bf3fddc77551306c24af49b9f195485648e12c8a9677e86279b2eefd
zb4b78d3a14e43b5061cf7eef9fe5460b9c29bf4ebfe3d3a950f24ffd545e6ac0174db8a7ceac8d
zc59f3b67d7c4ebdeeff08025011a0c3b0c480068dca83a36c82e81637c4a732885115dd9261063
zababcdb0355b078ca6d3b6f1f96fd158a336e736049e3d6ef657f992e4a71db375176c1e0cb9ab
z1d331fca2169841c719d5dc9b359397825f9f1cb078f30d988d0c7c5f3f99a1a9aaef9ada6c11a
z881b4f4e6b8c12e4d3fd141dc08d5c62e16bb0fc10bfb09715fbf350c65ad2505348844ca9da33
zfaf93950ed7b6d6da03cefce4a726169096b74d0cf97ea34d8f37671e8ee00592c0bde7bb98966
z67f51f2766fc65eb694e3d465ca927529d5084252c4fefed0d062c79f69e287d24858f05cdb6fb
za4e0508b0f153f577838533a8f140c596c42d9029808476dacc701be902a05507371247ca5d6e3
zc5f8367acc6fb292da97d9b9852314dbc4807cbed12c1e337e82bf12ba06ee919b4f4446acaabd
zbf1599b35810bcbfd819dd5e75d44f9486c0cc3eb2129a1e948cd14805a5464b9096de30e1b54a
zca85a7bfe0692fb04388d6902ccb8f17ba4d60e1f0732ea86f38aec7b019a8314c1b16a97e773d
zc134f91826e58720cedd39ff1be723453b9c140672633a3ded95e7ba8ac336e96cc6d193767a58
z8c97a642c4aec53720de381eabfec6938f00a46348d950b2696d3e7b75da4d816d496d70f7e851
zf0c0329aa875063f119a9a414a7f469764f42491cf787098f220b45c4c08dcbf2a226d35a88414
z867e3d63f66627f78acf3956ff112ab8fde35823c2d284384a3f51bfc788b3484c3e8449eef691
z5a9017ee9e4725aceacfe394ed10010925d0a153d95c5f08540ea4b232ca096d67333030cc88bf
z9196bed31a0bc0a7084a1a441963785c775eca9edfd607af033f3e1e20e4b1d459c91b8d893ae3
zcb93a1b4601580be05e850b50a59b576192d264b6ca499017d3a4fc1cfa3c0f2924009d1d408ff
zf821c3e817cadf23d95f64f4dbc493b7fe11aa3a0d5cf0d01c14f1fa005accc15fdcec4fd385cc
z808359ffac7f40626bd8dd5d036b746340854df05cb7cc45b245f11b1b67ce2d7990f2bf117e1a
z5270d6db26603418c56a73d1274751082670c82aa502d5eed0810f56f5913f863a333c3b57fc14
z39b113c3ce6b1e424af6b7ebc250aa958cd025eab6194271ff14bfe9ca7bd838a4ea91ad81351d
z325f86f4a80240b34f8b952087218c96c3f6e2d696ddb0157150b5ddf5c52dd35c75b2e6dd2b12
z39561cb5273337fa1d15fff8a525f6c9fd41860dcd0924f9053915329ae7fa0d8edf9c6dd6d4b1
z455bbd5190b683f12f0506bbee6902e211b05ebb727cf8df626d4b0f891f60c6b6100afe417f9b
z1f936ee30de29e30d9afde3048c23922b5faf739f9c5ef7d54d352b61b3b30306ff7cbd38a51b7
zec2c3abf4288bf0c150437dfe078acfb93017d28ad0955cc5aa32f706e82e49c3973a46c81d680
zd671d75acf3d1dda6aafe0f7d082e996e9a4b4ff585372079023d79f5d22b1983ea163249879ac
z9efa4812f36ccd06f6da9a5976abd59904c5a5c05b6c4aa364402b9a234254b46038eaf0f953c8
z67b6f99fe4c28375fe96152551e8855c30559da4b642074dd16dcd60dd71e66d88fa6eac12c613
za1f5fee3ee729055e2cde202013a7a89110a42b8e5dab88f81f9dc4ef2f8b612e649c42c5bf8d7
ze50f7f900dca08b8ec47c9df3c20928a8aaa2c3851dfcc2c5d3fc89e28ce1a3fc1c80b593c314d
ze77266a56f7355a3ac420a4061a88bd6358b3f3c6ee2e8895ce4bf19052517faa7ee6ae4add03f
z808d93c00aa8da9393a525a8e8cfb063484e1ab6bdedc355eea577fa58d2a55f9eb09c908888b9
zc37485b9ac66e76cd072fb97435baa6ffff54016498d282b631e370e009fcc6a31271ce0e0a3b8
z756d42b18760c33ccad9b91b211a7f01c6156a761592afb642a13b28528cc6135cd0f2cbf14c8d
zfb3836f8a3ccac222e8109ab06463ef7852fb5ce34f2f9397b62f4b5b2da38ff64dbd477847450
zc01a9024db05472382917d8a65f81d7c2d2e240fcadc831c6c8db0129b2872ecc7a2136121120f
z104df93148a37c655d923d3d5f9eb70e16cc266f725bfc1f895ce725d1bce6b6fdf4416294b726
z6fe083cec197c69fb7acd496773eb4f817f57d28ca71536712983fc700ad46c00b55e99562adfe
z063d2a07e26f09bba1f60c576e81dbc902b1ab84747080c4a44b19a961bccd2f27565136244136
z79382e08e69bebf5be0622048dd3c4aace3f7e99f579b8be7d38de908ded52849c95c7fb348e68
z8e9a6154c3c22bf440342b053164911918cad7ac795530f40f48498845162d0d0ce4a70d7b6182
ze2356ff36e17a57751154a074a9a3deaa2faf61314c280a61236d9ed35bd6bd21688d2cef54f05
z8399b48684c5f2fdbbac1111b79a30bd70585aafc2166dc1ee4a8438caad76b9ddfb85a890d29d
z314134d5e7a0a2c4500332fcb80f0ce6b2879293967b889d19a578ad5c70ed3c2d76c6671f0c6b
zd5d61ac4f665e4cb71e21eadadd25a93d55d360cd8607f0062db5ba8b495e4782608580f920e50
z254a87853f99e4e4481a50af49c5173720d8369042219dddedef793baa8a9b5c174e6e1c6c1f67
z64ed7f57efe4f825a744774630c2ab56f4f64433061027fa3e7f369c61ceba90186b49e7bedbb2
z1390a3b41d9219a947a14b7cd5bfca225d5f7f80579c2ea00fa9ec5377258de7de516d4c103fb6
z15e872979015b2daa70edf9cfabaa05f16e0901b425f23eb3f4405dde6fc0495d922736a69be3c
za9c7d1a266ce7163172b986a88ab7833d10903dca4eaa93d7ab96708f8320f3bea339b65b6cf0e
z618daaa665b8ae04f193b42a3d208ae8c5fdd4868a22f8883098336c13f25a829a852a8deb9ddc
za073327187a02549ed072dd5413a55b9bf121d340c34ed5969d4f91ceb98d297f46686f5af198b
z679adba671cae64e9bf58985f9ebe7a749f8e5c6925c543852e5e334c8ebfb6efc86d8e7369825
za8c5aed3463985c698121889081b7ab0440e53eb1ba3d1a574f092194ae0770aa9b2ba37f28d7c
z91331621bb4e883da0422e7d860a738c2274dee77a51c4dbb77ecd9c52928c22774a40938bda9d
zd879600c9e8e4a83cb3e3cec5e727bbcbfebe4f3adca3814034ee596ef4eaca5cca5fe849f6183
zc219e5d5a1391f3076ce9a5dd5c0dbe6bc8c4b90e430564304cd5237647e5c215d7b9e9092ec67
zfcf0ace1e11a1faac8e4498c68e10e2fc34708903f7b67e8508d50e7e1e20e46bbd9cb5b19b68a
z975f4f69132233a67bbef52b959c8da845370fac3563158643ff83f921f511ecd77c573492269a
z0a5542066a8d8102e619cd38d975be7ca24daa4b04a3ac51dbcd17643d45807b9a89211ee37e6b
z1e4f80c68b3a045eca34a07517351dfc14270180511e6a2a96abd86147392fa4f562fccdc2ba63
zc00ea67e908b85aa20c2420de35a33c2fde17a190c7ec0da1677f748dac1ebf455326f7eca15b5
z0de0628eefa4657ce77b5a98a8041969bd11dc306c2d9cec4f0bbf07f8a57317ba03509fc1839b
ze96cb7f09916bb0bb4a4a5c7224304e20992294cfff8808ce5925180e16541e1faffc491ea1f64
zbfa546296f00c15b0e0b0ba89745faf5caecdc6ae707f5afd1718739c975ac54829734f46601ed
z8fa69b3b417ba816bebd1ea47c2797cd6af60eda97dd2b21c2cad6ebc9646be906a6048af5bb9d
ze9ac4086e0bbfb2f50151204451f062afb662d1cbb2591f69737f134aa7269d34380532a985a3c
z91c8a522bd12c7a4c541ddf0d0be18c0154782546d55edeb3467af05586b25b68b7c3fd927285d
z40c62ac0801089fd37fa6a4ccc6d2e672c385bc4bdd34c7f6989cb98dfc5d0fa04aa7f67d1a9ca
zc1c7b1adfa84a281fd5ba4befd2d4691cdfe7b68ad83380e86d77bf70876d00a9f544d0ab1129b
za5d67d3378d95ef0f85fe8decc78ab0ecca05ab865aba2772361d5c310532efa603f22d8a7eab1
ze91159ba9d53676e2ca990d250cfeba8e0bb66097f8097ac93b9f55c39683f1aafcd0d04147b7f
z1778a0c00392a354df400c693c443f0dcf90395955616b1076b163f6e1dd0546481cf79e3e08da
z672875080854a037663ede034e33ced42424ee398f49041a95b00b3962a26ed240a2e6eec8afb1
z543d5dd965bea2fe0075fee8f793bc2d460974a825cec38a0415162d3de6486dc9c197cd306878
z0d544a33fbbcedbaef9666fa43bcc0e7d6230eb5b3e17ada14d4c7c0c1d95e22a83ea23fcb56d8
z6ce3372b19cf6e128e3ebf187eff63c1b9a4c19b249a395cf6244e117cd885c5889d8f8d31e669
z02230187ba60e88cb46b77b21a530a6d31cb1c0628147ef4fdff66f27090bfab42cb6b6dad7116
z21bde22f33d9bdf27ed73989e8a71c2028ed68e42ebe736f2bb43a947cc6495b80c15c9c4ea376
z195013267cc7ac11b325a2e72f61c5e757cdb7054773b92fe3ec5e959dce8454a38abb0fbc9826
z88b5947906b97613d06b7ff08fb04316c808c488b530880fb8abf55f0c846ced8b0ff8f1b6f3e0
zeb1f9bd8e7dd2f9308085544da5b3de4d18ba26daa006d2a89bd5943773123b0c28d3583d9fc31
z4d27d14d6b6807bcd4e78a82568703161cbfe582bda33f34961831f133bc0f8c8279968b0e4bf5
zce5bb4a375d5853f5cd97f0c0b4e06b1b763bd8afa6bcb8e7ceeb954a725fbbffd16ab454a1915
z180a8b2203f33e9e89be2e599e910ab94559d50742aecf28bbaf2ea60242d40f4a4576ceceec51
zca3b068f69130bdfc7d9b877a74b7a2badc69a4dc9873b4b4e0b763001f3c5b5c37cb944c1855b
zdde110e6d6241ec8105f5931fc209d46c328af7ec3d3d3bd198b856f8be70da79d46cf97880915
zd6bf7e6f478b75d44ac0e0bb398469f12ee7a23f69cde99d6c987204df47e287f3a452e0f8f3b8
z8e87a0fa9a53ba69594c0d6be3b658acfc9968cf02f0fc3e0c78734395f375327ac5c69a907084
ze25cc2a6c36a621744bdff98ef9e37626b2cf4729157430b7ba4db256ca244800fe9ded3989876
ze9d4b441905d12a5e1b2da63d083742f2d090cfc83c37d5003c6cab105611e82015ab2ad3b6673
ze2cf3bcedd01698e3f14a1f5167f80f23bdc370b6b0b164338280e6bb0ba7ea1e6bcb270500fd4
z6e0813b0c44c4ed8b8f25a183bbae3dcbfe6d4ebe1a75a5dff01aeb673bf3761268a27cf13801a
z2f49089dd84ad497f5150d83280f20ac72ded8e8174b6cb86772dc0f46a57c7f62b148c1a108cb
z429a5657b4db85425f80d02f0a039bfba76559cebacf94999a9c73b3c0dd9328164e46e2ab12da
z2a95e8e315586a89bace6abfaac2f8a42106da01bdd7eca115670e58862c0daef2754d7f87cb16
za835b22b2e0fc7f7eca628ae29219a48082ad8d5c26c445ed86584f6b46e5a768fbb4107328108
zc0254a410ff100b6d4e6834f7389c0aa6b01cdcba4894f9e46eb8352bde60563a0c14d85b1c96d
z182342d1e8dc9dea502abefb6d5ab8aa0ad7c7278bc6e6e2917ed579f4e5c6cf898ac4f1f3e111
z1068412cd848d78e4e0b33b3792c58f8bf6c33e6c11790b1491303408d32eb2f8fe3d90e051e28
z5e895b083b17023233eec33221d0c52281724c1e3b6e83aecdaeb53fbdd8c965e156f6b1400f45
ze79d8aab5b604464417db88ed34043d57d65f97dff08514e1e7388ce55dd371de629a866e22740
zb4960b2e594b2b3c8127f1de2ccada8b795aa2751fb689446abe69d63c11a9bdc0b34d4020d518
z2619e59d5930a080abde5b1162d2ed94dcd084a6333685480c0ceb0160abdd94a4ea7dfbead6d0
z91a9f51ffa88439dceb8a538908f8e3b572e355881129af625a75802db208be79ce36f822f7423
z238c07c20b17ba7330b1b65ba15e7744d862ce836e88572f3e74a5c2489e2fe1ac5a6db54dfc71
z3b07e4753d94e45519639f5709ea6e0c49706e8b63629d113163793e41d492dabedbd7b32ea93d
z7d5451848a7ac165e92fb419c644f65fc2a62e6c0ac880b3c1cdb82bf1f01df4be463587731a3a
z4679baa8c8fc7810db8302db94e507a528ea536a4fb6be47eeff87020e6c6bc0e2253144ee5a65
z709c1860f5e60b5ee9d7365bb1e2d50af6a29fca3151a7a08e7248c7cf7571363c9c5c942c218d
zd134d46e1582a276ea8a0c912951aebd4fc6e49d1d08332bb5417352545a8119d7d32e1de8d7b1
z685876b08afa84c7fba4acae0aff8c1d5c9cda1e55f9e8cfefd3555129dbaac90918c7e8764a12
z18daf329a675e5bc68bab8745cc6f8a57052f390d6fc2b42e1b806dbcc1fac55358f5698d9f20c
z9c0095ff31f2a157402ab82b6d1bde8e9a2d332c4796669ca13c3b811a183b63e548e80b986869
zac34241fcc006ae1be5c1d9128da135741532f442eb79d866d2e35b2efa17cfb4935b57ab2b3ff
z563e3c00cac188045a3ec94a636ca157f2edf4631710c3e8ac67c8c80579124574c7c6e14f39da
zfed60c56fc3d2bbf8e995c3a1fafdc889872cc862528b773a77de3836a932981857a6ae7e15fed
zcc1fac19dd8f9d10f26b2b750cfa82d9b8a2a74e8ddf5205d8fdcb17bce1d827b5d47228e27a5c
z6cd4818ea6365cb615508fd5467c23395bb40ca6e66fffb77cb8f7f2273d325636ad7f3a2cf13d
zf78313c674a3f452c9dd44ec1fba39397ff7355b9cb0d186a38c6fd0dc7af5f2d9be2f2d3552f1
z4d8c3e961468443534a4ed5b65b3efc0fa22b81ddb05004f5982be1a9e203a997eea56bbff2c5f
z524cd01338a001d0db5ff4f0c34583314f8b0a3a67ec0a8e6a4d78596b92f3e6ec44bd800a26bb
z92a3dfa68e20045f252d8de1353f757b5c57b7a09f61b2fb7597001ebdbbb5ae4bad5742ab2dec
zfcbd407fb83fd4aaf2d1a28d3f91b2c13405a08fa7bc97a18cac47bda4ae6e60fa751500776bb8
ze29d9765ca2a5a65d2c2dd9fd0c319e647e043df09eace0a6fd5a9ae90ae81b6b8f7f17aaf45ad
z12a548451cd95290c7c5d91aa952f95f8fd17edf10da44bef5853727a31a75e9ceed07e6c06a41
z718a7b6babf237fdc564d5df6a5940d199623b419d2b68db1b74e61353a2942c5785af9ae6d081
zce1bd4795430c1d08d1ec5987585b0ceda8edac2776f98dfcfcd395d258085f228b304d58612ad
z628a072874c73f16742544e5cc3f60aeb87604d3e5b280126bcc3c541496d8410361b6fa270bfb
z1479d4ff0f24187935271d54f0f0f70c013c22ca92a6181f9c55c31abadd64314cb04348e74290
ze8f561c3d1860cf25912aaebe5a2badade7177f5c2995e25b13045323a1176a9f175b564da75a6
z87ac109fa325b6f9e74ffe5ae7ca4984aa8ab2d2260a02cada93fb687d860e18a12ce97a528bb0
zdd9a0240991af2279e8d27ffd56861d25365cf7cdebe8c75adbcd6a681ce9445563119ccf60a30
zbd23b95d355288d51489af95ebf1eef5d07fa9b6560df0a0cb6083aee9e3cad44a557f3858d328
z8e4225be66e0d3095d5cbcc45c2185f8fa26ead2b3c30a9fd06f682743f7331bd03ce4785cae35
zae67d831f18ce3ed48e513f1c111be9845b04b51bcc481e9f35f9afa68d3dbe4e24019a7694da3
zf418045c898166176c85d040ae204b043506d2e7f3ecff10cac3f45f901a520bf709d587b422a2
zb652631f5226ee78b0ca8271fa63af333e4b3d3e61f69ae1d658d628ac251515742cf6f7dc3e07
z004afd63beab391d533e8dde15d157c75f74f8e5427460cf7855790786fd208bb697278afcdf4d
z11dc065bdd3b1b084cc81f1fbd232f56441cd2a6a01b933a8dd538384bbbb5118fe0eaa61fd59e
z20560dc8ff00cb93778cd24abf140a5138887b87e9068fa2f83c0671458107758e796b587fbda0
zf73430942fe9fe4da1bea269950113f9ce609bb77e27b96369e71a7c2f793c23865253c8a54cbb
z0b72c72e25172dd097492f4ef3c31f92105876498d66fb24365956ddcf6210073b75acbc4b4c2e
zec598a18e313ae7a2758588519608294f2d2d462474b913ef403c8acddec996eab368aeab29b55
zfb9c720b3a8194fb91dcc8c5ae966f9ff73896a568e8217e77eef4872329b74db905e2ce6c13bb
z7b543c738eb2420ed53ee3c90828db9ec79bf1c9b3073c628535882977d14daf175847633b7ccb
zc978284b44dc8cd085ea115ee10401909ef2cb3eea6111b9e943565f57e073c65b2de3f3ce07c6
z65935ac154c6452d408dad6b5e5b8e2744b86843ae4ce36da7462dc78bf7bf6399ab87e14eaf45
zd2b91679e957a229138b5ad7cfd9904568c737fbd3445549c3fa702ea491c093ee9f39391c0193
zae6cf7bb398d3e57936539b8c3563ce15fda94d34462569672ad8b9565d75f88c58182c06a314f
z11e679cf65b6deca0956098e03ad5ce2df5429ff7daa8bb6a2e495501b16628da60c6e296da10b
z4839b874b805aeacda7730cd1c6712233b0d286d1aabdb4d2affafe691b7e15873b4dc6eb7f03e
zfb51c9d0aeb8e321ee6d02fef41f2e861003be7acc3cdf63f38fbef4a4813a7a3186b4c592ea60
z97ad53b04688f3590bab832845576d1832453d36c4b85e5866a3a5ed64a182e8ff6ad001b039ac
zd4ace9d99862ee7a5fd69a1e8e4aed827666752b2cdf3aa2babc865431a5e60fe30eac07fb8089
z7f1707b08b243e3335d77c268da80360056ea7d9f6eab63564ec62c6d8e7b9dcde7f490c4bebce
z2324fbbcd4dc2dfc035c17eb704af9df086559c601d8a819b428e3f78d95ab59cc41a69e7f3d74
z03a3e1cc9e192b022cd63e6bde7d7a66cfd60a6f62af6dee662d8c6e2dc93b9d6bcf255e2948f8
z2fdf1d3945ebc2c3554cb186d1970d66cc7591a5a99b51831b9cdfe666ec7dc53ca5c5b6413efc
z1639d906f10ea8cd42ced3c1a5998dd31e0c78103746edea751ed0f9dab70f9e4c8b3f17f99e6a
z2ac76247a15594a29c41b371565e38125e4fde4b858f46ca8dc7d396246bf98219faea0263b11e
z4355dde04aaf23af48e75a54d4e4a8fadfd49ddbdfdadbd7887c8b70d31579aaa22636424ca815
zd9c90d53de7b13eef128a03356a4da5a32b8efa1aacc5c534e1408c6a65e1cb255d94462c2fde1
za2b47dd708180ea2b9e0373705e85361a16310add8869f1b0b7e5ce17e1f8db20143d45dacb5ce
z8eac2ac38f44f6d90f96093ade99efb48c8b5f53df92fa0ca5f9fd8938aaf6641e04724a9bbe77
z69979f2f82289fc2d58a00151e6a074341f0418f205300322b9424d2d7b48b947ab42b4f8ce031
zc26a5c27a42a3d7b650d89088c7f25e2a770ba88f88e33d676084fbaacea0adac1bc6e7d404cc0
z325fb733b347042bb0505cb1bdf3856a194bddbfd78424fa769f72e9a3079fba4a5c2b2c7f666e
z3cf26b02e77d15710459a7a92e9e2949444fc3585f7fa01cec398db47109e83dae4b9b1d599cdf
za0b996d99c480f5e803c4de0665329c8212c6082c86df62feeaaa3b7c7d6292872eb65371ea657
z165842034ad4d8493f23e8e9c9b39dac7325a547e9f009958b5610e8598b2443b719e6829b85da
ze1605c412598e9797e416e7181a2d63c8fc614272afd2a5de694243d94c1252db1d7dcf0e13a6d
zf09809268784212c0dac2977c9d4befe8e9d112b0421d1eec2fc8b554f3e78223febf3767ef57d
ze24bfcc746eba513cb95545e8be3c82f149281c7fb4dca148ab7374e31908ea812de414872c4da
ze7ad42cfac2d36a006184233ef65f9fa836e25b09ec2c41c832b083f9ba0915ac8b3c7c84e6f5e
z0cbb26b7ae9ca5793fdec938c53f03c5901908b867d80979153af7c53013c14861662adda04106
zed81a683d6cc209a22b860b8795c14e5e4d0834640d6ef7f98bb58595e767f2c0f6665a4984cd6
z81ce206b3ff1348ca7baf9a5f0a29bf601a4da83a5172631bc61aae5ccd8417e16c1d1a5c66f1f
z9d16e44693bf2f424361c2e411c7a64e66da7b24c35a42b83df3f325959bcad08dc3ee51db3287
zc99ec39c61ee180f1d3aba311e9314bb731c69b227028aa9c83f5651f3dda7245d5f034a09cfb0
zece0ae5a2b23be4256cafd9cb8ed4edc64457982ba84d824b224ae648b8e15312cb274f9d27fed
z1b46716cac9f1567c63b489a4ca66fc42db122a8f104b403412c712a9e56431503b8064d248181
zdd88a631609e525361cd8e93ef4ff99062a65edef9494bdaeb600f2c2a9052d5a8398651d4636f
zed6a283b2be8d69cc45d97efe2a982a979e3e4b0f7ed18a45286ae7d84adce03f78314f1e0f75d
z0229bf09b07dd356982c24f70c8943edd9b1881dd8cd85f9cdb2d91abe99d2fd74679adc76f881
zae3b34d1f07c93f100ceca3b4603ea1102b1a0a06bd4b473bddc2902bb0097394ef168c0923346
ze09aa654fbf87b538ae553548b97c8815a495556996de5b10cd4cf8d2a01a31dfe572a83d37b19
zb997dc5b5be79a30af65d73de1d731151f0391292924123afbdc09b7bb437d8871c5531a61a903
zebdc91d504f9a22f1c49abec39c80598bb62836b32180d0d47fa3a40069c9d2a38c107f9b460a6
z028c1604778c838e4704e445ab6e4fdc80f48b77a5615d4620ac796dfb14ed9b5d6f92d32ff466
zee766287ea8a499eb84036825fdda0cf0daeed8c27387d6d97f33b57d8ba19af17144fac411ee4
zf96b60928cc1ec518aeac640223c470ca98329a820c98f5de41c1277167f1ec10d10c36308176e
z225076e95a9c760088bb3286cde78f60a8fab41c0883178d9bd1a9e8da2737ffcba8ca7cd321c0
z1ca1bb754b8d346924031a9cde169e7816a039eca814f1f15483a42353882899b30e55e8550174
z3ea0ea3b70facea20ce4a4ba82ae8e608ee4a2a7add170303fe8aa483e4363ae09ef65b3b269fe
zdf5b90d2c49bc81c738e0f39f19407ab1ff576319c77a2207f04122440e92b650eaef557b6ade5
zc4a9f680a6b55ef3cd304a26e5fc4bd22125c0712990a84d20bb723d662135f3cfda9d971a7826
z03c2493b4e48a0e071e79ea60c96bcf533912bf7ef9c9901d8077e11d2e74ac5843bee380c825e
z096b11929a163a0cde05d7707b3d2e2528c32ca475d90304670f20159fdef7ada29f98c3d2c68a
z2d57dee4bddea8a49d31b98251455d4efbcebfb0ad0793584ada6fcb222b01d6f7e7c5c07adfd7
zec6aba4d831e6610e94a969faf33f32397b92d4fdd916ced68b87e7128fadb5f143b15c94a89ef
z4ba443cadf7210c472cdedea54320fe00654b604d6b7f1117f4ec79d326bfb3ed25b3478173fd4
z564c31a06cecea24d91e7eddc39023a32976f7da69960a29b64f49a3af654610be693a957de9f9
z1adaaa79ad02eeadb018bef6606356e867aa5bd0f6c9637b13e7fa0317187ce3fbc88c3c6f2039
zeddf411757e53260c0c3d0f711cb2a0146d00388d59d04acd15cbb233acf769315bf720a27dfd7
zedbba38eae537bb90278435bce6159dc316b3fbc0dc1eeafac996e3a04d244b3b60ed8a2a81aa7
z7f8923e8ec89a5d58aecea68960b90896205f7844266a02e4016dd8307624d61d5fa8c74f527ef
z0e39dc8d12bd6431232fa4598b04347638057ec4c6083e5b7a422e91f2ade813d6c5bf099cff15
z38e8c40f151ace53f3b8817b3aaf6fabc6e4abbdbbe754e87d3f83418b1aaa98bd0addcf1a017a
ze355e3fa951c8d2fd7e6f35684a57d00ed8672947f58a9d23dd978bb11cec1075f694b7c313664
z244eaf73fdf8ad5f2c411f12c813ca58fbab7cad0a357e828dc0a0f5bca6962aa4f97bc94ff83d
ze0dedd83262d5abea434680de75ebd2ff1cf45911964aebb4272a8b105a400d12ae3dcb4b09670
zf5b0a4fad9c9d2e810bd518bd1d8602dae430c10955de25d561fad1a38997c927103ce5640780d
zb4ed14804f2905ef5bc848940863a23e62756b5bd2d5881745f497bcf4b8bf6ee48753716ac51a
z8d0e6a9428c4cff81a7b830af169ada8babcd80189c157c0b49e8f11f88e0ee25e9521c502db6d
z76a8fbb9d56880811d33eba5fe5043368925a7c9dc7aeb58a768806acf23727e5bd51d3424d747
z1c2e66d6078204212babe8e6a956aa0ace3ea97720e9c4eb7731d60a39621aca0f69c229646030
zb37db8bef99ca2ae9a2633d1faa75cbb5896668d97b37135846cfe1fb329e7ab18daf1516c3737
za4af9a401809aeae9f2a0df249ec1a1ff9bbc7a92714ed63c9388f33c9f25fba3782fb8589a99b
z3b5b6f2e74fe234d777fe9de7be83051f74e747b0d77a0871132fb9959e064c9d004f798d2d316
zc748ca56023984b29ec19d1edd048e8e14255730119629f7aa4574f4c1bd387667989a19aa4577
zce6be31c6e5a9e61007b883097b5e5b72550c603aaafbd8ae3627133a301e70050b071b620be52
za59e6c0ded0e20f53fe3fae197c7c9703572509b4e7bb91e41b48343c20c711aff43f85f91ad74
z6e11a15a6a6e65147ce64221af84c670296c27d7322ed2dd424ee882526e74bbfa08aeeebb5795
zc4980d5f487a4e2fd96c20f0ee00c71d571af9b6aa8c2599af47a6faee346698538e0dd3c521e4
ze5d716093589ffac8d6b3b4b8fd8702fa0498061d67513c5e5e4e5691fe44274513dd06cede251
z1cf8afa98347b71381bf7d58c28b4244ca970e4d00bdc780701e4c19d8417145f36203cb6d05ee
ze82cbe9c30a9ed209671cf6826b8721f3e1cea1bd5625328f0313dbd3f30f38b3df1dadb7ee3a4
z5e1e3406f523bc8c2ba88c768b64d042a73c2b8f27fadd647544ef29556daeeceedfb3cfe37f78
z2afa698a55f51bd51942308c3013989030cec1ac416387768e950ae0adff05d8535ca68b4312e7
z5baab205e957caad29553576c1e0e4b0592478f97dc9b41fe2d8244736eb615b7d041e88374f52
z38ed7e41364d9529e640f23243851b25d88fcd4ef5889b873a3832165b47bbbca382dd750ba975
zd665939436115af7a89ecab74361403c397cd68d8fe40e36b4e2e82851a47b2a1f5c70c8bc4806
zc7e946278e0e88b21a94a9356633434c3a52e16429128cee98d188a6e14ea9c09a00804d1b1100
zf82b5c558846cab3f7195ac43e21f4690b3428b737d14d8da33a136a5f5e8e3d6668ab305d0f5e
z57b178d7961380e657b98372d34491b86baf38d52212d067983f0acfeb911a3e153193caf29813
zf73f7dd6ef542911af4de5a1e8788168c2766450cc9123d9809a5a8fc2eaaf1e160db0cf757f98
z31163a43f919d77ef4a2cb618a077b5fd826e19c7aba9f7251b4c89a71b07d92ed8444e6d2c1dd
z78db3a7eb3a3a669b0ccaebf5f4e0c47ea838a052ebdf6ee1db57d8329175119714f76a0602587
z1c3767bc1f09b27a34e1208135f5c584374cf3dfa3d257e38ee5a59d1f8b902fe669f8e2cd230a
z14e7f03adcff6cc38f6d301890566e37c8f9b2bb2ba8514aa310980f0d5041bde0796ee74c2fb8
zcee298101df76962444f63bdf19c36ba622962d6489f82b38aadf7cf97b76dc3fa7dc2ced58ed2
z0006a02b7123406265a08ed19d4f143964afe80bd42963f0b403d1c6093795b324d6a948ecc0ec
zd08f9d9101ad0c0fd9b0a72f17aee4f745de9e13525f0fe5198d7b64b60cb2d02afdefe2842e14
ze3ceb718401377b42cf886c7245d3a58d2bf5e52a98feadab717a3b67f37a8c35988d4e7f26d10
z94956d56ffe8bf7cb12cbfb518c330bf4c3ad330b832184693639cd11af70c7d71e3433cca11ec
zae7631e1dd6cc4652569421556c5f7a311c4e3e3674f76fc59ab9a9dae909a4b4c77c4dcb65882
ze6edfd15f339d5c9de101c7720133b01f8ab3081a736085f05e359cd3392e725f3af8c21398de6
z08579e64b088d3b41f3ed0c2412de38defdb752796b12f3cc3f075d95783613ff2a60141d3bc19
zcea6a685a1bd679052a097788e3125c1cf7e4f743c3877fb80c322da751f94caf3cbed5f354db2
z4912d7b5e343283c3a7e5577dcdb932d71d2cc12d6de0619b00138e0a9c863436d041a87d357e4
zf61a7f0ad7649a1c2aa110b76bc4eae9fb7933f266fe470eff25854420720cb1ab24fca975c51b
z4732ec48bb86b9e01a8c96510dc8d3ab3be204edc60d787ee89523350044a8328dc5cc84e74e6b
z107e0ec843babf1d1533d290645e3d48b0e2b21098d12de6c6dd0ea854719c04a5b9ad73bab9a4
z715f1ff543fa9b2b238536f363ce6b70bd66d0510544019024ca4804aa6777d16ee25e16876f43
z17ceaaf53dd0775f1667d0a1599795875cddd3760b9bf0651d22ebbc76f95df762ac86dfcf684d
zdd66d829a9587688ef90f17b93d02c42fd239241ffdd5b5b823774df1510b070e0c25c1ded9864
z99dbd52ec6cbddf6975664436540b7fc3d6304f539521f3462336f0dea609ef836d2a3c6106b00
z3471106e8c47741aae49882b2ade111eb371b7dc5e1ab7ebb8f3e5f0dde4f567c2aa133324d958
z909f511d1f74e21dca5755ac55cbf562cb3f11f6ba4bfbadbeafb245ee517ce13c6f7c2e546de4
zc59ce44d0bbe0d751ce831e9b9563fe48e626dd94e650a049d8470b56724f01410c5c242813259
z5e2e2938d1617fa0e1fb58e665461ca39e21f99403a33c831f0e45ec815d2dc827a7393b68397f
zd18d58b8b0046ee778de2a6e4542a5f5f5b93661bf50a75374750d28ef90dace5913611f4def49
z329a677550b4a8814ea2298600bfc5e05ca5ec2cc4121e19ec4a31fa2297a8387efcec2c380166
z8221c2e441243fad5c36ec64d8faf5fc358f29a32e1028526c34d8e3f7d9757c550af5429d0e13
z92119cacc2d23146650b7b77c8903c15c274d1b37bfe46f55fff1923c6974193874b249e2c926b
z996723e8aa7be07ec80deeff83497c3f4a7277cb62ef44444bd96a507f9852833e415f55f46c41
z8ab9f899912a703f8c5a9077f4034d08d5f674565097bdb58ff89de176acc08267a51497fc39d8
zf16358a170da19b309fc5be6b30b2645dd21c4d2419f4d6fc9b0128096cbd4cc03b7b3f29b431e
z3bd541b9cc35d7b120ea318907411994a5d33b4a13ea798760f432732c8e83d9ad83c782ceab10
z5c4b81d961941c0731d28a7ef573c5de10f8b4c7f0f52ea31ddf733a6cc701a0039adfc961db7f
z759825e1fa1aa2ea771f0bb9b1b3236937032a56a45b0ab93d05c5254319f7dd20085af15e43ef
z5a7fd4350e60eb463232d62a2811559dff3becd3b76e37fad87a9aede0c737fb2804bd56d0948c
z156c3a49741717428d837f41cf5a10897980372a1488d4d7dc1e51ddba6322226cd594827bbb1f
zc1f67be1bd2f8d335ce8c394d77e4a85d8f63207bc05c1a123fcb368985b1e81149816165753fe
zf4b1581042224df40c4ce9cabecebbe99c1724998766f16872a710660741d816640df7c5d9c1ab
zb289648f582c74a5a8b62f0d9b24a5bad97aff9b253ed6df873c953a8f1ba6e6f7a4d79dc58f5c
z051f08fa7c0a6b27147d918830260614608db67e413888d79dcace79b589f1141d59748a654ef2
z0579692458ee136017c5c5f465b16bb0b384e52d62e5e314d52f2eb9a76b45800c10a67367bf14
z5e5600bb397da8bf9722e7b4ce5c0b58a1124005b261f21f1e1fb53a0834e7e04d89d74fd3af01
zaa14409299904e005db595f69b36f3b8d68ebbe522d0f0a3f206b49a8b9a6985f160ddc803434b
z6baffced08daaaaf792d22b98276b32a0f3311fd1bb7a63fdbcbcb64ce3c1c1322ac041c4722fc
zf6f9dae14fb5176b6f9139dcc464f4a21d475314a0c7091a9d53bda5c756133590c4c25fe09b7b
zc4c04b4ead7daa37cc01a449e19fde8b1d680a80a0194b60236b389169dd04e395690ee03a9071
zd030d71915000d681cfd64cab71cd6a850cc9b8f8f8378baffb633a0cf421a387acd871e1ea2b2
z46417b87b6800664ffc956b8b09ce4518ae5c60b32dbd99c21b7b5dd31674c4b6b3469609b20db
z1a1a5c04b48663605853f703eacb6c0ae23c3b2ebe713fc68772967aacf5c0ca5f97a1d2010995
za49e2a081ffec173d6d45bb9ad883afc6a450b519d90998b31e6c00d70ed38040daf87e8bbb9ba
zd9ea61fe460db13ed2f2c302773c3c16b918de2cc710ae8a9b4a64b727a879fcf4c7764349992a
zcd5fe728fe103b771a5e0658b158a7737f24368e1f85c2c9d197dc692d7f2bde037bc05d909ccd
zf7e3513da41195935d24f51c9cdcd6ad432165fea891fd022eb3f70fa1491a24b387064f7e0695
zaa7c8ccfaea59350c406dbab771581b36e6367b9c6627cf3c46c54457c237dc714cbeb31a0b970
z6310de1fc4761898f1e708db8ccf874c2960c2d71cc6985ec63ba3f653939d18d3eb912055c424
ze16313c9817e979bc2f85f3998be8b396af84613ca5df2164b5d0e82c3086375617cf780ff6cb5
za58e45b96b7462172b3b0813d4265bf7df995df555397994dc554d9cfd0add1992d07652174eb2
z7935e482f510d7b146ff39c801c43010073163783657a5eebf515ce95f7679f59c1b292bba3290
ze30128d86c395ae73e4dfc49bb924861d5e87d7177fbe5632e7e22d5aa55bd3ebfc01c4dad66c7
z92cc6410a38e255d5f80c50528c6a26b0be9bf48ed5b53a8c34f9e5a71abd30dcd8d669a2c61b9
z18204419ce4ba5362408339440e343a42bd45c36726c884ae879f3bb39e793313b9a171b5800ee
z896d33a2d3f1f4961118ee7bc2118ef8fc0bfa543d950e3374d47500cd6bc5f7ec4f444865a12e
z5b021cc69407f5fe3b60a262516852da14213adee5c2ee0c8f5ad2542ea89c6a4c5626addd9f71
zba74f411aadb8f39d6a9e5153d2eaf47ff757b8b23ad882f29fcc2e5e14b9d60e4129c0ef40f4e
z5cc6358a32af92dd074846419d9a6f63e3e42ac1b7b4f503311b651bfb27a13fb4df5404b687ef
z79113c353d2cbcebf3319e2b22e6b5bf387f79d0930a61512fe3d7ce06e7bc7701841851d80762
zfe5708be7a73a3135ebaffd478ba4bb738cc9cadfb0e3384ee68a6b030e8fcdece51521bd187ec
z1cb2fcea853b3a42149b712534317482b5b0d32abb53c60fabf2ce3b0bf31ab78005bb547b3080
z8dcf5b1cd6ec67aebb279e853008bf61df9953f9df8a73e90ced10a4b19de8464da29aad75fd1e
zb242e1c1834b26839a4a09360cdda4a3ffea6ec86d9d9e0905936ebb146934e06ad08962459819
z7eccd235fbd696fa5dd2b76f75144a522f2c666f0b5f733ed31ed901347fed9ae3d2915d376394
zaf646194f8b4088c5d911e769d0d2041f2cc13f3c5371038b03f58a3afd039be3d7e3acdd4e9e3
z977b5bd024c60d183c268ae1e06ab2249ddb59b1fa5f4551ef54f129273ce951e4ba8512909f3f
zf721716119e10889dd50d91ae0c5737967212286f223c7436dba61bf519b074af8a6f89ce24048
z8a7acc5ec943e5cbdf35d8746153489e16ae49e50186b43b1fad81b88c1b65d62a9a11948a302a
zcc347b1794c38c380c7f816af6a7e906a143ddab3ca8caa4a5d61022c0d8e6ac8d31088ecb10b2
z750ba6b9ea4b5a88ea91e5e38dc26c3ac57b33321eaade1215ab7f87c0491b38d05ad5972a3773
ze8131c74e5c7eac0bab908935299a0730c22718872ccf3560f27fde5598f1546b48cb51ee1e1ab
z77861a808ac7a13155a8755f2250d5d53de2037fffbf169a2b42fff63ab4335a8a26176e5e99a8
z9f71b836d86c0171dc6cf6c58cfcd7e8ab1be056eeefbd342aac4b8d6cfd888976cc1ce2c2c1e0
z5332c8949bc997103fd56c1b7b77afd3b5909ddb1c211cb9861dca9bcda4a226a90e7a51465f2e
z198ef854bfc0a79b9dddac751630e8d41e782e0e7e5e9dd3c19f0930355d85432d42cb1e0559a1
zac6719015e57ed6e454032a927d8346fa63142da881564ac3d4cb88a595ab6bfb24143fc1b598a
z372c9b56c8033a116b93978eb7c8448b2aeabf3155defef94468da115278b0fcb86156c440e196
z33f4f8ce887222762953989b0615f110d438a26a27a1f9bb9aa409c97fd828cde55e9f103f77cc
zdf22f2753b0f6f1082aba43a051e8057ead88ab511ba7fb0aed17e6e8209cc8e9c463becd6f5cd
z084371bd90aa3e2d1655ef0cfcd3a5d72af25dfdac10607f77032b075fe285158d01e2cc8578d8
z9f1af7f92ab27d3329089e17db1b1f892848b2091866fc0f88bf371b525c59e76b5d5a06eaad8f
z9b0cb17ecf96fc7246f4b59883d5c6ac9d3fb6f23745bb803349c70c4558c215122b55a89987da
z7edc843e91bcd65968e35cf493c509bc9722f68d0a230ce028a6643b6306f06f3e62292bd92c55
zb7414555ca90a9980827ef81190e597361657ce465ef2232af3a1af5d74876ef8d378b7758ca95
zb39a3eac655e15fed5a59f906dfac7e2844dea0b1d849e35217f33f30eca221fcabc0539c9187e
z48a6fcdea637e8929b41da3cb84c2e3e8124d50de8504f5611ccda038256ec4e673c971726eba5
z8304bb818e15db19e6f1b937ee5fa07f1b13327dde0ceeb08ac54cc3ac213eb9fed56d6ad2e2c2
zfadfc7664c0949ec79d9a935534720682024628fc104a43208ae8605b79550f6efbc2a1da5acae
ze282e01719b0304d01ce6b7795275c7ffffcc0163f89bd4e1a1ba4de4d3334b9aa3a4cb0c900bc
z2e0c318fbf194051c80ab89a7b52a46fa456b7c07676fcfde7217d4912da1ad209762a3dae5113
z8af76ac4037b89889448745f6e24a6a3330ada3e359c635a270839bde86be6f59e53ff6f55bdc5
zfa47cf19a21d110baae902d8bca14300d633b1b2878b689d54b8917d97ac500cbbc6f82c547cbf
zb334283f768b839382c1d979e46e6fc70981eddf198af84e7729b4c8cab49445de0a8fd2922542
z8769dd08434ebfe6410f8690d76ec88febb1a226338e3708f80fb7118fe3b7ff444d9d83f2a54e
zd6f3ea27a2050e60da6bc48d73c6dc88d5cf75fc512ceba418547bb0a0c9c9a3635a02eb8cf1f9
zb81a9d5090421c996d02761e075d3c3d3ea0aa977e49349079c0d98bf28b8d7153b00603e3660e
z64c5c197cfd1d16a9959652b4f60241607af42dee38821188d8e92603ffaa5dcfe9fb653839a18
z6056ca15ba42150493cc6c0473a080428da29334e0d6e93a098255cb84868226be1e209b7849ff
z8f9296f6588cf919526e677a9dd15db9e620d7680f68d1236eec1ef976163d9b303a809ed027cd
za3789585071b437aa1a5507253a30995675c9703b33599940bb933ba847ad2e1a8c37d66667870
z16dcf434f75c50694aee0efea710a632d8c32b7efcde97bd86855212e5d47f45fbace4e0cd5ae5
zadfdc42c7d44f905d052ccd9ca0ab331577d94d990fedf5f9157924d156595419cce2930c2b4d4
z99c46aa52b783a0daac1207b2eb75059f74b9e033997967773c0aa8af562b1a1a4b10cf3d37dfc
z5d24ce71d40ae2d6f9b87e27e40e86854e500ef61b98b8aed42a619e3d764de35d65c1667c456c
zaa336afa776e203b7989cb6e1f489c9c03cf1f2551446ea71aeb02c2e301c0157990a33346ede7
z0d196e194e098907607f06446dc7acb42f762e82cd3786b556c4d3d90ac39842f1b68a42390169
z53ca25a831425ba9da3b558cbdaaab64dba0bf50b45f435703d680b2a66116e1d3537cf3803f10
z8402239abe094c141a32de7cafb4835335461abde88ad7d491b2d3d9dd98743f18bc6cee9ca633
z1e84295d81147e093e9147ed8c3ca13e7daca55dd6c49a114089997e167c4920f8f6f8e62ce8a2
ze3a67196589b87fb7d1597c0998fb11cde56d444d8f3ddd4383314d7bfe3816d43c60be289af88
z9ba23fb0364e811da338ead5cc52c856ee3e05efb12358a8204dda788738d11e072aa444e9dca1
zfe9ff98552ae51604e76c0c64d5fd785590e75f88d4a969e4499f73f04a71ed4dd12eb8a752d9b
z263b9e38983f5a968376e14d58b319e50d4a0c721524a88113833e48b18cb93c06e12f24a1b140
z27031ffcad4de7b7ab3a781062097c84bf3c3577f953bb510e49c23aedaa18aff7862981f53eaf
zd24a0eb614da3183f3e1778671af621b4e613fdf1fffa9d611ba0730ac9958ad40c6fd03b179d6
zdb9836520f19d9a739e2b53e0f01ea0a5a2086e3f9a870814c5f1393db11cba925ae6f31f84a5a
z56b9339b333e459cf9dbf789c94272123b4b6dcf9b452fd3d4ab796070a21191a4597d7dc321d4
z0922774067582e5cfe547152bc529bebed9f1c532c82e3ac50eaff7c7c99b8f53676854b7101c8
z678f3839e255cdcbc2c516cdc603aa7a178f17c071cc9718e8e0b490d9c88165da997cb79558bb
za05761cf31b8fdc87551c7439477d5891506c661e9b8e785f96c653117c771a0ab7c1fd59bd10a
z2722c7f576617a1df9f780b759d3d162cff22ba6238c3d732d632a278c0c421017e77363ef3927
z01a63440c5a5b2a477f6496c67cfef44ec1c70d54133c9fbfe08158da01058ec5cf092c13d9213
z6eec89821872fa64924e5f72d701edd3930753df14032849685f3516e5af092fce3bee085bb03b
zb00e329df41deb11ddf146a9dd44d16041336b6440d59f1be04f2462f9ff5a10b0dc0661cc9ed6
z096f05b2864e770d6512053d99286d4580e9b264048e430bf6fecb45c4f1349491c2631be8e1c8
z78fca507e1cdb7a4e011d756c654b755ac857e4811dac65e78b1850983c460a9550bd83f3d5f74
zfc108bb7a5096b6f39293633fe3e021545ba961cd7d1cf84f55282fd1c2225785cc0e1e5b100aa
z1a0cfbe3c6babf96d121a9162d332f44702c5e0446855a70cb9c3eb7a776374697742a612648ab
zd1d026327fe1287817caa3823bb896e059bfb66cd6f2d1d97e6bcb3f773351f802216aea319868
z2055f9f002ff130f00326d55a31040d8d81636badd21e8e35ced95bec4a607cb2c9941bc9ccf7e
zf655f31aff366ec130795856b83051f17c3f1584cae1792f38c40ac43bc199875072f3325dd36e
zf8deaedd5cb3172be0e967995d4ad15e75983b820475a6e1229b971bd0969a316c68c392cb3556
zff93fe139d405a5d08d0ff2a41b0230f77fd43bfc829cce9f95bffbba715c3cb9de4413a06b894
z3c626ed75fa4207020e3e7817c233feeae6d814592e853c42e3d04bf759bda5eae63647edbc745
z98b3b3cbc6882384d22f09efd1037957b8c38c2669a2e499fe9f4a062d21c48ffed5477863c935
z92142a4c7b7a2c2d305752d750726c743cc4cdc1f84068d83bdffb3b4c6a86bca22f218d8adec0
zd6a3b737d1a523ec54e8297dc516c4329d0ff0ddf6ffa937e2f9cd5bdadd9a1a18ba2f3867f418
z7afb51dace6d0bf86b1bd0eb6eb6f3a7d8848816578149ca356a7e9ac42c566c90944d82d79f19
za1b26444f21a424478ff440dc39564bf353fa59aa5284225641f1e765de079cae18818e5a21c7f
zc5ebb6e2c4f420ad802e20a2f57ea54df29db16df21ce15c3636bbc2421952e1796f3b307dd722
z899a685b9a673363b38029a36d2dcfa6197cdd2f7fcd8e537ae7e39318377bcdd6b390c374d945
z4bbf3644dbc5795c3649db1f9a1b428b8b435faf1f3c660e71e059d83d3f98a8d0049ae7e68f14
zb527bf5c160225636918ce500bee3715885f1bca24a540f9abf4465417bb2c3fcfdabad4085853
z6f8bf41bf434c6dcaa927cedf34fa4bf15b4b39376687c1f01b4d6e6fc2aa704dd2336be70a7e7
z8fc74e1e63fcb8619dd4de9e1302f48823b43d54348a7b1e5eb77bbaab4aef30a96435339282b4
z22bebd79bd5e3bbb49d7b201d9b98fb4b9e8edd47f499f1b00583c85ec4d0867843f4a0718b3b0
z0ea30a80a5ee954d17de38ece77c02f72a6ce58f1b489c7bde4211d05f30be3aff669d9ed6a1c1
z8746ceec191c4a29919a0b4448adf92906573afd9b32eb856be628e288c263b9903c7752d2a81a
zafee35c613a30f0faab09e15e90d2721581e49e373b2445d36892f9a8ae62106681c5ad6e4f183
z6acc18658370c93b6cfe9ad14ade0483c210117f8ad0102d3310cd487268c8d0dd1f8204e2e1e4
z98160ab181f9fbf868dcfc909f5874a0749f6eff0f8c88be0d133e0c5dfe72aa95c6c4267e6d58
z86438c13e70ca3b5c1caa8e5827f86fc627ab977b7b2248130647242d8524e1ccfd3932ff92b52
zd95128f99aad2fb3491941ca9451e0edbb3d510907f33761b0edeafae0009e9c979b3c5f1db216
ze9ad77f2a0520dca72a389518f158e59ff7628cdd012e91b1dacc22b2d4dac2b43de688c92b2dd
zf1853a9dd67cb89eb3638b94984370f0d060c937ddeb56ff5dc8819950661651722390c109a16d
z1088e728a5ceb013a5766a2a51d35bf73eefec87d0756ac9435a5c1878b02a703d0dba1f7e2c87
z178775d004f398da4bbf6aa180cdaa04f8705a492cb2492fc46d8d9f2bdcfe0d4022a8c99e1df7
z9ada823c4b7753343acd04cee5de6e561dfd878e1ad4e305aaa62ab44a0c021183becb817e546d
zb3683aae3b14f3bf8f94a1dc847ac3b39afeeac37a91701f22df19cf48ff48f3eb327140f8c2b0
z0a05190d064fc2a2c1f70caa51283d3a7a8ef366d1c17ce002362f4baf600c46c4fa3403463f6b
z2abefbd9bf09f68f38bcd0234fd738c6df265ce6a9b927b3a5aabafffe2eeab7529ebb250f5190
z900e3bf25acb4ccce0ac43d4d8e85279a48e451db8197139d5bbac99589ddbd27cf915a6401d6c
zd73223cbe8f61b655f21600522d5c4228aa289b3a61a276c99c26c8159e710a0e4287cd3ce17c4
z8b2a4ec1b5a2f8d6ddbd46a0693cdc1a160ea06127c152a1c2cb9870f729067e1d40681ee0fd77
z8ad608fd2beadbcd90497c5a6d8d8dfd07a403b0f7e8fcc6b0dad06a89c9ee4f43e56c2e47bc97
z2e546347a60fdca6c5a1ac24f3d28211bc6b6db89545123ad2a571e30b13c5aedbe29b2f186dea
zd40d76c49dc3600b3a94489472eade957dca03e086136372ef341fb8a7c1987c803e4485864ba8
zb3bb78e0992b78448c281b0bce396316a70893219c031bb9ff31b58806ee3d138d36505bda15d6
z022219e9a715fb025b631ee8354238ab74f5d9aa8013d5288d64e255442ae756c7d77a082bdf38
z010f3710693e8d95c298a9f6cdfe82d5f2d11d5511efb53ca53a89f70870754cf68b6a74000395
zca76161465a70eab1dbd43a8eb841945aa0aaa177716cfcac2ed32f5cf274549e53f858cfa762d
zeb43d6967c8f58d559d3ff6244ac8d605dc8da21b5ee09340ab1678a66593f3e686eda22fae989
z14bf33ced7fd34cbf75e68aab915e1cbd732dfd401deb657aad7379867d33e052e76ea8d1cfffe
z0e336ff6ddcc3f25cf613aa881c4bfc02adfe335a30c0d52e8b48861faf0e25712e8d15f23e8d4
z059182ff46435fafb1629000e6cde12eb67126f6b15856ae845f27e222b447650fd011af492594
ze7851060290235e421228b4777a7319020d786bdc90724134e41fc57856b472f911fbde81f210a
z54f0126ae5e9353fd1c56593272032913fed51a120a35003897676576585f44f4120c3eed02221
z4d25550a782c56daed1591269b8bbaf49b8dc567b8d033e28e31c4393eeb8c7e1dad0abad966b2
z995324ba3355322ea65c4218272bad9541b782223027f4085630d2a18b4b0338c0295d1868901f
zfab3064536dce19806977244e5c75ef4e16b1bf9021e8ce3adac99ea980d51848b24839840fc1e
ze2c8cab1161d495447d6f4e6a4f55c406928c0d89eb304900e5dee5833179dde6f916a67a2adb6
z95103a813d9550dd4e9a496df42ef28e60f1860343b2de624fd5484cf70b9530f5987731efeb6d
z9b0bbade86d86c634b4fd3be222a630b866469c0cf3bed6bd0f859aa1fe4e80269c1ca0dcc39b3
z79a9d8c2947ca01dadc63573669322fe98fb326771bb0fecb3aa7439afeb2f5506114e6009e904
z2daa3b3293f9fcc6568e2d6ad9fb2809b2f0cb15c2c927ea7ad924dc18dc53a54d374060afeccb
z154a47aee94dfc3c6ade1843945bd55f9347071a8a36e0b88c66c305fb16b64281e410141512a5
z334d7f212c9ea0d0169a331a71aa8c70f5e1715281803fd1c01ad9ae755a9077db0e8cb53cc1ba
za656e74a9d8dab548a03969c0d3a2c19370e50f3800666ad65eb46a4b6d6088867cde4b1f2211b
zd4ef85daafc80dcdc6258652f2e66d48676cb786f41ce2591c9c3678ab795166bca7f1f5e0aef0
z95978c742f2ddff5d7a425de253a0ec1f3bc1013b0097f50fc5849d6fc514549c419e43d1c6864
z3a0feb3b0122cf418f9fbf48041830dcd972200a22ec8f2d8aee194ef5ab1d5002cea157e41ff7
zcf9b8fde7826b3bbf2d09715b74a236b95917791ae2bde94ebf28169e880f3872be70fa980f685
z206ab4634226c0f872e598fdc79c171cd3eca1b3a69e1b582638aa79e26b236c27a6754a9fefe4
zb0642a5f217faf3ce7f3408353744ce39af4c0aa734266424f5a847831dc64b8f14c03a40fa240
z34e4d3ac87c159b4daaaf92d0a3d0b246c75170b31173bb74e614c5e47e525b04d10707dda0130
zb12b73099eac053293b58be8bf69df525becc0190a44dba66619b5d20507e02ed5591d0c2a1f8c
z969da2f1c430a1a32df4468c75aad747ae3a897d29df2e121d52c0c853541664f72a6fe5690f0d
ze39113d9161b39b0b88947a04d6b90e54aaf5b3082b86f153e202ea2e2003e7b983b4873275037
z96fe7eec3b7d6f5852423375a7d7d8e2b82a51d0534cf0d6718413a86b99bb89aa2e67349efb97
z60413835a725c00c571d33996cdfeb5ac9acff12ad948dc68282d1e63ae5c759d96a5abb440933
z8b8148e9d883161f9cb2bcc34ff966083b8cc9bc2033ff69c1161a62ac8eba4c1fecb9ef82bec6
zdfea24729e5049769d16815b1bce40a1488ae070bb1e97f8d132851f7db683b32a92ea601c6c6b
zd794d7e81b884e1cdf35698c4abd2e93417b04493a53cecfb8832bb3043c5ea759241647f02f4e
z1b22c0f36073a2efa4b5cb46577ec55a829fdfd9d6657de0bf2b9ef86b59022461430f1a3e3a08
z6885590d4283f34270d8fe3c82c9299c986aefc36aa51aad24b95db4a9746f15f705c349dd1370
za7664af7a54f78c2ea5d26474d54ede5224f947bf2687704405a8b31580f300c6265513dc0b206
zc3ac3739b772d7706470e6863163e20bdc94bf37e1e2da1fa09a73121e513c40472e7b89a6f27d
z6126190c61474b50b21c94161276e86d0a3c4f24aff42d43513105f69ad16906d71f6491a16488
z358f09a36168a6e8905301e367bd14c2776e7332880bf8a97009fe0bef2f1d659ccc20a9159736
zbb27ebb2148b4af5073bcfa3102f75ef8ecbdc8323fa86a13256cb500966876559f3834e3e87fa
z50eae68e62b16ebcd8c37217c168444dab950ea47b7e023c98745ead50062f1f6a7aee2fc22251
z2c36d27689c9b2c130bbe8acfc7c5660002638eda47b3376962ce1e227f9d1f0927938072c9fc4
z98629c5bdd3c2db0ea7327f06c98b71cea82e736c4581e8818635c2b45fe153bc387b69114eb52
z5bd36b7b3b416bd6dd769d9683399889b15cd3bb348fc8db7b79dfb1ebf9b1855d4d3efa928bf1
ze06d76e5e506d653b840220e79363911061ad49638af5d925a200d75f3e0cb4130b9b99316d00b
z2203a0bb596095593a0d7ddf66f77a3b8083e750a360c29edd59b5d3c75f97d7538bc37334149a
zf99566ac855f000549084194dd1855760f9b831eb71032f8b2273617f172b8abf3eff6929b24e7
z87ad253635f713a111364aee4bde7c79b8955b117e3cdb109ee886607c5cc2f5e49fef56c7f82e
z16158e025391d3a10144d48d63fdbbd89adb242ab11d2de7d7a4ae5d7b248358bea389253c3175
zff8d6a9ae54de7846c2f6e5e5e578a668558d8a184af822e7a6abb810d419f4fe18055b2e6ef4b
z8069354a993c80d9635eb498009154a0572a8f6cc56c15bbb3253902ac169df415b129776c6a5e
zf060d136fc4835dfff1e2f1084c16ba32c9e5f9ace682820538aa31a92b080dfae0a4e0f4d94e0
z86155f35e173f500756464bf385cfe3895cdc7cf162838de119f231e560c2cfd81dfb2d85408e3
z8963babb2e09135889a893ab7f69f4e61b768d44329967f21d91c1a50573dd9435d24c6a5d54b5
z9ebb5300ffe04bfedfcf212e4be60b5af76e897f2bdd288ca5cf8b29e8cdb6429e300bb4c0a481
z04565789586b582dbcabef5ed1c78a4aa74d9c08bbf1dfb28527320efaf91c4b712141f9448b20
zcb908d6ad47c728a947f59a1fcf4038e687df4f023576c0ce446889d175e8aebab3ea869ffa9c8
z13f02b5b78a3709fef3e60f0c5a379181bc5f1be917d8281c1121751f6e7193a680bb72df9e6af
z6e167642a3f572d04b7ef2c867da8102232edd4909b042c1b8f6bd139404337bc50071cedf2ffd
zd83b37472a6e61aa6e1d35d53ff942d4d9061f4c217f85b051c85415ceeef513aa76deb4b905ab
zde291152ce5815873f78c8d93998d4ec45496199a319b4dda86bfdfb55e940b92838b691cf919d
z6c5ef2f6dd8459d13ed3acd12f88ecbc4d8200297b0eb013d2398eab70613efa4ccf612cb740c6
zf21bab2a5f5d8b474817c401e54524cab13eea54917f499435e5c05fd1fee2e6e882243f1fbacb
z99b977ff11d80dca1b95ce6c3d6782a1bd7637f2b85c08bbca741d70b4e002619b8f988c767f0a
za87221182bf13c1d18c38084080851ead51de476cd6d6709a38f568b17ab4009765eac2b938ed8
zf4e734ca772d113c1842c214c634ea26e1695af351e1af495f5f888ab2511217f1cab005690109
zd0bb90c82b53b02eb4eed7bbae25d1f37f4c7962340ab5743d00e5f7475680fdddfbe8d70e037f
zc57f0a14ccf34e8d5a150c0b50bb40fba2f16eacbb6c0fca908047f20840d124abd577f661f5eb
zec3d22d64305d76c1e00cbfc676b09c2ae379d656d5659a83980e6776323ab0fadee5d01021fed
zc86eb7b281f5a61c725076e46f8b3088d6d9acacb823bc0a4d4efb43513fa525f9afe24a60c8be
z41ec4cc0479fa564cfcad11ac6c2dcf922b5bf94246eb16c814e743353e1d4a74b3d7df8d393c3
za6bbbfa4c54368e261212a5d43b36854980829fd5fe8d7b8d5ed44253269d782fb444f83cc0947
zf9184c40d544288e359d3174bf62a449c386fcfeef2d5ab5f499f021b2a02b5de4fcc77b1aee93
z3b0bde428202e1d592f96a4538152db0f14309db4b99998cf07c0e7e286557e0103afcae5eaf9b
z772e33bd4bb6383d58e4b39c128937cd629502c11a41e875f1d1488e820a46cbe9b40f2c4d8d33
z54ac367ec619ee96b5face812dde4179b56d65f4016395c088ff0a78a633d554c6d76f25b62962
z09a89fe6a3109627edcbb7d35500de541d3034a3a1da755fcaa793e861a12d683d0b62302b6baf
zd2adbc08cbcb62e9ff68cf27b7082ec8cd2fd657ec2294c811a822462781efccecbe5428a9828e
zb940703b9f4d9d7c176699c8c6972e73d33e50e6b5a4a7f5aa930e117127dc51e1d081bedff39c
z15e45765c92a5a91a9627f0a3f6a3d15749d2d0415715612e7a9b9f3a8b870a1864550fa6add18
z239016b7fda589556257df95f77717cea62edc8b8f91564d5736f4fc846deb2cebe4efa55466fd
z53d69cc84a1b59f705733a07d7ef13bca448c1e346a26e786437159ec6caf3188e0826fbe7bc09
zb93b9fc786f3834de6d1a755f026b64bc36137b47ba759518a24cada2a4e3d1431eae0a7b6dd8e
z266b4533c5a8872cc869308559e7f2def9530db7a36415487e2158d843a19dc3b5d1a43f34a6b2
z1abcb1e2940f697d58d1070d9eef3aac6122bbc3269ce22e1ccb6051424ef0a9b5bf90f48be80f
zbc6ef093886f7e00ed65389701ca7397c432690048efbcda6fc996486fb93223f83643c1e44d40
ze08c58472c3732055eac45cfec2217caec00ce418c4dec90bc9046e665fe3a89e165c590b8f1d0
ze394e59131b31b775e4ca4a411a3d25c658895b7d87f6c72f67925b74c7a26075f8f6dda237671
z039706bc84e8b6ae6b9febc9fbbd2946c3bc1adfec2891b5496aea20410837ccf93b60df06800a
z86a3c46ddf9cf19e343a4abf2ce48a8bda20c0c4669b913c218b3b649a4f3b1d133e79345923f6
zd433d2828023f006d387f118542bb134ca32295db5f91030156fe5f9c5e66d99e08f95707faeae
z6319f20b39a83b67549cc3a940691b4464aa7d083b5637384794a912185ba09372f34375f150d3
z3e37a0ac432a6605db112b5667d4830552a126689b69b371a94427e301d2a8ddfd7f2add48d08a
zf6f4e6482ff721bbf8fe0f18fa9955272bb3b8276617597b8dfdb3964a1b6895967fd0cb148259
z44aa23ddb68c36b3a676179753df42b58f37cf97e828cb622049c157beadbdf47f4f3be68d7708
z3eb1074c623dc838d6c13f9c249ce3360b0662c946345be6d761e34cc3af52b79b4a9a4624a4c6
z798a9c76379c2d476ab5a3555042b3b973454e038adf1c2b4603f01b9a14cc86c3b280286a7c43
z2c6d631f0f32fb3a9ec191d968bb5e9abb51c6be20116fe19600df465291e1b9e3516c1b7a72ac
za4648a07ae0e9cdea53e2ee118b0cd7b6cf6435a921b61f686ebe8419c3b6daff68449938c50c1
z253edb3489aeb9bd45510731eec19256146c8cad6226501a88daebf870fabbbfa4c295174f9927
z20f6d865754dc41cfb10baccde20b6a145ba3cba6d1fcc12b58a77f2f0cd0726a8ee2cd8f0de13
zd5d3c4e1ab42fb1f4e0d1b75178346ae6443b35ae32b2031650913c1463c48f751de31893639ab
zd6d17c790e921b6b4db51b17c4fa87dbb11bf93b4adf2fad76b91c9671b2ccf0c8b8fd582454ac
z9a6880cc8029b9f13bfbed627106c639c019ed788aaba534ab3b506120f6499ad8a9663cdb299b
ze5b91dd8546a4813543b7bf5a140927e15a7237ea8ac403e91ccbd4828cde2b1059b2c58e4420c
za3749e1363d46bda5b98cd9ae5f88980e11b1ee4aed822cadb215e3af9c0638ec82b939867765b
z267338fa9696900a5433b05cb55644258585086c52cffaa618b2b0a40854100cc33d187ce64526
z8082df256a747d83fb349cfc820381c07e58d3e524ee46ead963fbb7290b6d87e5b371c3c52c97
zcf0eb09fa50555198a30fca53aa5d896155ebfb2cff6aa49fa54c236449ae5537a6de2c9c52e42
zca47215a5a1ce013ee0c34dda5dd5fbd39623d4471e932ede9220534a7a6d52ab49081671a673d
z23ba57a8afe7b2c90cffdacb23b07b58dd9a49d80e74676bcd9158536155017a12b24783d9a46e
z8024c95b7fdf59a6d613ad1d4967f546c140fd24d91f9e9c124b1d4dead1579a84b3d31cb985df
z0bffa544af6d7fb7ff9058676ac9175fe89c983356946ee8fb62c3eb191175c7773375efedd51e
z91bc510808358a1ab508aadcbeddd8eb625d16bd77193c1f4ee39776a512a4d703eba1122ee770
z62ae67951128fd3a573e705c6887d0fbf32be99d069d45cf8edb8841a23775b65ed68c0caae76a
z23c0e582d6cad5c7aa2b7531cb142a24cbfc14080da9542a2750b9ebdf3dc8620c361bb191f1d1
z55e51898262dad7851b8087c64174ebdb274695fa80daae20a5b1efecd731ad27302d7f5b64f0f
z7b80cbc371a6dc03dec02a61ba4523a0dbda8f4c2fcd3c4cd44aa518a0f74055727c50e899189d
z4be8c41326b93f50dd011666e0cef94719ce3f8914479af2f61301d476fe926a06658d0c96d2e7
z1ffec1e66d1df842e618d0fcfd8c9727acfaf213c4c1a6d708c031a2d310df02e406a8123ab21c
z8894c67b78d04e66fa68669f6995d2839bc7105dc8ddc29a4880c3aca82b186bb7509db30bc3e9
z5df045eb96888ddd0b78b4845cd34e543d7376d84d1d7769e44f2045d82aa09ad7827963f9e844
z3cb6e5f965fe343316c62a55480a7cb6170dde59014b712394853c4bdc4788ecc68cf558606196
z861bcfdbe1a1541c5142d1a1bac492caadb76370f22e0504eccdf32c3a4678f6c1e93ca5d8c271
z83da7e09fb2699e1510692c46bcaddd8389914ba6729428d92e8a904669f6531ccffec10a562ab
zb0e56c006f1931e4151bf1a947aa6e355ce18460a806049eb21074dcd98e0d6c91e4ba32c966ca
z8fe39d5a9afde1a6c5669cc0f03dc2f1d3ceac148d4bdf86f03bc539fbc0f49c96c465fa1b8333
zd10636ef529e2396ccfecad67288139f583195d22bb313f96d253089811790074f4c3fe5ea830e
z54ffb6998e3269087c618a3a9c391ce982f919b158392de5427fdbbb37d012ba01e38a65612be7
zfa3344948c6118988c37ce9406c3afc80a4dcf66531d625136d5d3624ea0646c6ebe00605473cc
zabdf9a4447665028da19bc2e193390944d8c07072dc956f5457c773c0cb5f33b36358907405faf
zf2d951811f4c678685a8afc6865d189eceb1df9265be46f880d87ee3453904765b28471ace7f6a
z24b857672cae55eab00e1800ca580cdf0ddefeca2037f1c7ce4e1702b9fda73c79cad63502288f
z4b43d742b8fb1ff4b77dbba723e5031e9fc2d69aa34e74adf8b7679ff396f3e409acff4130a0c4
zc79242ddf3342c97a5fd3fe1f5a06dc872331a82320b5d5b1bdca025d565e68c53439e0bee3315
zd3e20628122d07e1f9c1665104da2f7b6164bc311e19b9721f55efc97ee0f59aea6172f29a85f1
z1a70725207ce25877981237795057e7cefc072b3dee4b3b8d17ddc8883b5df69c3af1a2bb48d04
z7cb1e21a314574878570f4eb6fa362cc66f0de3c240f243758c2f60d4ee675325c361f87abceb1
z93f941ec8266b1fe1e57684cded68445a206ca0c1fe29d8529225e337b92c8169cfdfcd445842c
z5ada1e10a653bd5baf335e2a2f5d52e2e6f70fb184b8f6efa6f4d01cf795b839e41f33cb762671
z9e25d1b3b7a62894de94b7516c93053f0900906e7e927299b14224e320ccb19b1202de6393f412
z7635da71539ff6712143723882b1e3733c05468860e6d5a203442431654bd2826241e68e20d936
z3fca06f49c79091bb97ee144c98ec3cb82379d39102d611734caa2d6521a58bce93ac87c5f0e41
z7c14d80aace492cca880bc5fb8ad2cd58b918985c64fd6fc2b5f641aaec9b651aa25fb3ec5004e
z9ccb08bf938de7b63bc16ee0f5f2967ea1447bd6a6401ddf4fef3e8949ad4732e85169b09dfad2
z8786571f1b40a56a7c3c07cf4a39c81c3cbfd283a080d712f461350f5fcead54ee6289e4e177a7
zea29ee7d8115bd900dc6ab68e6f80e4a0ce5e1eb373fdb3ceeafe24d5af87e0162cbac76cca8e9
ze464761a546ca79924b1cded1f7dff49dea10c482a140e4bb438e3a520e5c44d61406905fe3e1f
z8f765f0d52b5cba37d77121dd993c9cfe3d685a275a68cd3dba82556d28717ea3a12f0c338fb2f
z69bec839379a2ea18500305fc161dc64984cee4943bac06af7095d0b709096de5d2d0e8c8b8070
z296ffc3a7799d182b38c44c7659cb2d7102d6d6cfd21388818a6859fd41092143a944483a4ae94
z4c84ebf6dcafd7142c363c2baf9d8ff3cb0682c0abd09336e8e0287575ccf834d79ba69cf3725f
zc2124fab15c83b6bfb73f2dca32dd9ebff2600f68e9714f6fbb8e264158152bf8108f05a5294ff
zf983cb8890e1857673dec011b50643d650039dce77f5ba459e623a6d655f1e7100e6b3709b06ea
z9c1d6e937b2523e79a80acf51958bbc2ddbbddcc2adeae565d2c05dbb87eb3257faff97006671d
z0a47ee95e674be5d17d8651d53d99d3bf6a343e0f526da6f2f2a50a75455f7ea7c27574bcf0077
ze16372b5ae57940a30395089a86e69483c7fc1cff74486958901180a9f56e90e998eb9a94b3983
zcbdae9a83b0fb59225fa8ecdd9b0ce715ec5f9b8cd5496e7f18fa23ac5722c37bcdf9c6705b237
z68c4b8c0aaf4f53d3a01d39679b396b2acf2487307c4c5fd52ac77cd2b4668ffb1a322dca1a97f
zb8eeef23cc18e2e4b83818b392121063f54bd980bd5c6ea29960d91da11cfbec363ecfc0a8c10d
zbea925f36c87fcaa8bcb74de7d33e7c46a3b751e3c94fa1e9f079c32250576a3863841e33614d2
z7e996047f0151f64d1d9c5ddce543f52523c84c5de307e1320286c000dad0bfa34c62efa7c12de
z95e2da3a142997daaba6598f76ec863389d40deebec0de796e6e82f2b1633fa451ea3ddbe355bd
z3f4e259ffe335fa26dd422b6c8f2eca5904f7ed098e078fcb5fe9fec9e62ff25a4998cc5b152a6
z507ef669efc083907dec6805ea52521040708689e5de5d0e5c79f5319bbaee985a6a3d916bc1dd
za10fd3962152ead0d235c722526fd848f2a46e7edca726f026a3ee5bb5f9f8a9e04e2713c96cdf
zd9435ac555e7fb56347e762fa6c7dbe1e2e7cb9cffa8f94a339ec7214769661cf56ac8ad2600f4
z4eb5cace5d70520a0d62f0f4950cd5234dc01e87949c8f399656e7d18e4441a6e48be92edd3795
zdc6bd53770aa5054c2b9bce4dd0d18a43fa630cce334daf2fdbbb862f4873a3d24ff90e8de4977
z7b8635eb9830441cc32cee9f66e3f45d4968016d53887febc7eac6850c2d426f3106ff063288ee
za45aa095914b0505094c2da847fd65ebd00e9bb5288cb42f1e07afc2bdc45e97342963995e7bf6
z39002ef2a17d91b0c1360052a379657e0526fc26366a20661c378a1ff76d9d33a1e08abfb201e6
z42360391f877c6f70b43214a61132c0a556858c5a2df5c94b8f8e9a2df5ee0477d0797f6149e6a
z3ebe6aae154492565426e00a8441d0ed7645a4f7616c89a9953c5b79f88fb3ac27c3f5af573679
z2f5fec77a6a70f5a4e2417a31bf7874b299e88f9bb508cf97485fe9778152ccd18e592ea83840c
za5697b8d4cfed615939ca7267a1bca285fb88cb6e17adecce8d778dc92295ea553609609fc5855
z7cbd05a3ab94938c9237daecf6544830a3b8a684d83a89f2f0f5812709e7bca2822d8dc5f2f876
zd059aa70f79464d1b155b5a66bfd19a7e8cf08dc1b83148028c49e39ef24cdc4c30656dcdc3bf5
zfd99a97fa69aafd69468c66ed424f5adef626e41e32ae8b5beef2b8e3b141f7462f78dcc89fbda
zaad7e81d5525457f364c5311c466d98a81f0e9966f153dd3b97829ad6e1face3c4e654e9002653
z6039f877b4fb9192a7987414fb8f886613cd8ec4cc535ec8c8ac67ef2ba1ad8814f69e6402acdc
z12d58f98d98a5dab47ed079efd946c09ae388aaaf25503f9c82213c7a618031d0e2014b3d42ab7
za5716a4bd851d0e69285e660780a927b2b24b38b0a9f6d198330096b5e99b3d69c019ab55f2f8d
z6a3b1394b96be102e1003e429d4b895d82f0774dfd72d544022fa385829e63c011b4052262b079
z755c4c2683b847cc5bb5ed78244c451d8a6c9fb7d079c4978ea5b4e0632646a4fd575b23de5844
z42400942269da9a55b341e91f4521eb146261c47cbeb73a95c2eecfb9d29f5468834d84aaeb40f
z36a6dffe33d4d9d3e92ad03c8ffb2f112e7bfe9065fa78a3cb010eb39201ce7010b7451be7c28b
zf7acd46d9f5fad142ac37db0b56d791172e056eed5084378b26d5ff83c448f4a3162e750fd8d5d
zf8804ea004f5b6da2f3a5173e8b82717c90eb69f8df0b13d0e48e80aa6056f65c612a04e3d48fe
z39490a6093e2e3188d5dba500e8e415bfba0d56437e7c5f2386a3ad538d0c0725316b56099a4a7
z2f7e5c1619d052b4a425c25139e54aed7bdd66f1158920968acd8e838b41307f1d75cc5faaa0af
z1ffc96d3d6be408e94b0671f200380485ba43389074b1a4efa5e4505b3dbc1d6d018220ba0fedb
zdcb7280a4bf8f16cde5008bb1cf868c44cc062feba00b10638f7e61b82c5f2bd50400478ab256e
z85dd7fd30f69747b56be0a7105db2c30d2a31528b5f3ad3382e453730d07a19798c06f7f87d044
za8cd09c7b0a1c3e6365b5ecc9643d3eab986d7f3fd37c80bcc1417b24af0d60161567c1d604596
z7efe968f7495675dcfb90e2d1ef0bd267b5cd14007a865eecd9a58059fab3ebb9f34671cf9e941
z6d19e0342d337e5f5c060cef6b37c8be67d2f9e2877a769b7b936924c82a33dc635f92d726e741
zbe0b5912361dd515a530e091e56778853b145a826f66652dc496a91678e28a0502accc8f424e5c
ze3aa863682a04030dad097c6e046d621e4851dba15e0c9afb8793d825cdfa3edc666973093f4df
z2ea7abcf1bf57bf8a85b22d5bf2109880ca647a718d0e05b899561c5c5c10cbbae0f4dd7f56faf
z234023537e6f1f53a39164653cdf57d6ffdca99baf0ee38e9e0aadeb1dfbf765463ec70b1cc72d
z4d23f81add48d18faf06b4eb9dc2b66c38852afe4a1ef4552e88a2787d372635f97d9fdd3e2cc7
z77368d4159e1873dbc0b9df51d7c6fe8b2ca16a19e4721cdcb9beace107fef77be5784ed0cb23f
z5ccbcd69298c489ce6a2d8e0c932bc30ead98c008f233385da71d4a22a2a79b146627973484df8
zc3a42a1de5ae5c15b8122c41d1b69266c943b506db52a803f44d6beb87742a5e65bd99dfce7088
z186993232b16e4e6a2a0a00eae24e48613413e3cdabfee08889f5543652cecfa0c75d666601431
z1685b390772bdb4f51f7aab22cceb94e028478743b687ad9da089dfcc0156ef5483e252322805f
z4b601282cda5ebb0332acadcb9a2fe6ec9f77e144e93139c9526372a6c85151eeed27bf10587be
z8f3a3c7333713fd70e01bf55423cd792f6d86ad33db05a66718e2f6a17c47727792801b00f70bb
zd00fc4fa4701d64cb845552be75aac3c135b1a7ddc2566ae8f229bceacedb5dc0c5b50d090f4c6
z9ac1f84d550423d2b151c84b75cb5f04b19620ea5e910bdbe85e2aa37a9c261de1ef0cdc0a3fcf
z8ad61d3dda19be9dcbfed2bbdabe36d59982acf4f1fc1d101bb19331e3911e096fa6385f5c12a2
ze30dec09d6f09ab29d1370b05a27e84cc8fcbff03b2c853c49501f7c35bad1674a97a80a8b84cc
zf0c9e22c80772e2a12a318c3a7b6dcd1e7317c1a351a00831fe5ed49925396d55b47b2482a4a03
z9917ffa5a3728740622cdd07d74e82db116174700277fa0169994d4c57408552015ac00d59d3c8
zba838fd289f06095cce43804e2ba98ddebf7336eb6b027f308ae589470da79a9a6bb9258333a61
zb3097e9a40b663d8e9244ca7759bf2aab82b3897742d768ba1c58a90cc65d84c1cd8c5e897422d
z6ccfe0f9959337959752516e9bb311a7da72c7aa2f6228df5cef682c4320823b83b08cf8243a18
zb726614cdfad57d2ea2a3265e4e8fc02a430d98d55915ab92c3c9fa7b1526bbc8a886dc1b0c123
za1677291b81a4be9cb36ef25a6e6d4e56cc61dadc7d81fa18db6ce66e711439bec0f36521d4ce0
zc69d740fbcdf678974907a264f982292ab9149a8df89711a8087023092292ce53d84963a2655ec
zd2394210d43b400a4593ea0dddc717ed74b65054c448eb97b19e3c4b97f444fb9745a2a8c4788d
zcc968bc727ade91b0d87ba84cbfb3472bbb50989724fe63fd9606f5c0ff43dc9144f49eb210c08
z92852589af62875c4b032c5f8d0d8b49edf6aca8567063d98300ab8e979333436fe55467c84052
z3738ac37d1b76bd74b37bfef03cae455f6bb1c3bce40363b61631e8db61dc8dcc354abc95200f4
z6b8c78cb98be3b47fac332b818f483a00f76db56d4af0c49567ad9c12c36f90617cffa1d1975d9
zb586b77419546f3c31b14a53b6b7dbc1881f2ea2eed1125815d23a34decaedd93dd5c73981aa7a
z739a922e5916bc5485854b9d1937593ef76e65bce34301ed831441fa3aa0cd664b3e434e3f005b
z25565abe577c5d3a1f9558eec39d1c8f9145e0ed9948daacd359f898d5282f3ec27456f7898161
z36b372e78b7b370867c56446142edee1eb0665b3bb67e030bf726c7e0c729d8d305a09802847e4
zfbb78dd669ba028ae207213e38fae8fef612421c041a16d672b8f48fcc59781b0d55fb9743c1cf
z6f80e99aade2f0f3ed25828ca7f61cc2bdc60c759075400f16f369fbfbdfe4d98c7dfade9133d9
z3e0340e8aba1af766e2cc35271d5cad834887306b54f7bcd4006dcd5935eda7084ee1e9441ef7b
z85fbb089159a994015a0ad825e0e49a3e72a39677ed314ad5a53f269aa7da5c8065ca5bbe88fc2
z633a10040c1617783055b22e511493507e3febc46f31729b9344002e3501c368dd8c9055ac50ab
z09e156fb67cc8eedc3dcace28d6acb43950bf6d91318e2b43f904364ff3d25c34e8efff8bc1e79
z6492c6ad2ad7c612ac226b5d1862ce27b64e2684cf6310ffaccde1b6df0578a78c116137a24573
z6bf83c6d82739c3744c26f02edd1067d68f8800810f738cb4d0982756f8d0ca337a9ba8ebd2d17
z4ab2e15af0d9e0d4dce79aa46415c5cf01ed605bd251281a107c87d930e2c9fc58b08c0c70ee93
z6586fc41a5de0867427b6dc7a452ac68a47335c42577be08937db0c16df2f1f1e1cb55ee92b293
z71576cbd3234e84dc1062451157fcc37e1830c4dca0481e5a5165ae26ff33efd217969c9498247
z67f33d650af71e5408cce8007de46fb4a31dea875130a09191754389fff3c8ef6fe34e97490a4f
z03a1db2da58cdc270049239805e097b9ffac1d5225c4fbfc40ea4fbf7740685379688f059020d7
z49cf7e5d0c3680be228ae56b5d8a1ff914d106b2ddce450383d0b5dd11907832feb88b3b289565
zc635fcac5be46f644207c1e45f7dd83b18a7142cc76ba7c6021706649a88805e1bc390db292caa
zdef8de6b1e1e246f0614985f015505c0f932a99329b2ae3652bc6db1460edb9930f4562a5857af
z1cab811bba6da1cc4f7b224a15066d5733f95c655caddfe3ac7708be79f57c377fbcc1000691b6
zbb364bcddc20c5127d7d8b319a1a53e1743792524209bdc1e14e5191192f3cb8d28ba64b0ac90d
z6f9fe83f0c032950cbf6c6e5c752864dcfae25ef3797f21ee145cc175f2822c6125990b85f7a54
zc69d01faa9878440ded0b40574a8f424056e702853bcf90fd38fbeec162925edeef0c6e48e4b0c
z220d590784343b3844b4d4ca17d0c65e2dda32e9f8b8e379b5fc703f4abd067ecc95f9d5a3633b
zfe91cf1409bc53b2d92cba8a664c725063b921a3c1f2664613723cb9c2f6d9a7fc19accd1630b8
z2561c89384e7d351ab92299a341ced481d925208d0c04d46458b4a9fb19ff6c6c56c726f4039ce
z98864da9f2dbcbb4ffe5f0d3c4ab2ba2f0132afa6d5e1452283a93f475d5844f55e8db4a3bef77
z84786eb0fc43c53f4d72f1963feda4e04180518f4bc680b5bbfceb741519b2dc2d7cd7b7df36bc
zcc5189b197eab068c8cdeb9b47828960a890c8dc362dc4ffe48fd488429246c53d6b69ca3ecdd9
z7fa162db8256aa76f8afe386ff1d79ee6fbb4c1a5d098ad6dccf4adc05e8c6bdde8dd122872bdf
z0835497808c5bba54357c2aea736a012660d44fbaf55105b0e5decda639f25994e83ef9792ba9a
z013fe9dfe2d4c35361c16c4992b3ca7e47a3e68656d33e2baa34f36b0866e3e081a209396da1e9
ze7e889e695d3cecf4f553f2e704d75bb1e5bff3c3755c429b8ecdbc0a6c9e513547b1466cf4ca7
zf6d59f66559d0bd48aead7a1f50a8ccad70c5f1fad3c1a256d8814140779dbd9830c5d95699e23
zc659778de66a875903733b4ba5265b27658406aad89e07eec77cf6518921c8c899b24cf3de3d99
z631afc72afa0613efa94aa269440f735f4757122f2ad5febe98293c710a54950bb0604a55e05d3
z2f6d1cd1f8a960fed1f86aeb58bd73031ef85d36ff727d6b3de98e4eba73b4ba4f16b9364c6fd0
zeb839b57bcabf16838c6ab6df89bb000ea0d9b22331bc3ff7d2bced82b475c61128f9b85d750ee
z9a917430a87d035962f334b548ac173aae425a939441d842c89cb824558101fa81a35880f7cb77
zd997e65d41d842b0d46028a845f7d67b24daa5315c9011a3494afeeb780ea08ce34c6e09834d92
zba61132d55d4f88bba71aa91f4c39f058d71287815c93ff1b511d3ceb9027d19bc3db3e177f8be
z3973521f2e346b9ae7cbd4c87ffa343836ceb19747d1945ad04bd02f674fc1301ec6e1501b16cb
zc27bf88d98aeea8e68a6508dfaf4cac0f5b2d5ada49241cd68b4a5391bd324d103b26803cd1107
z3e7c42dc721c9481eef55ba628f620683a8714bf27232fc8067159bbc4dbfa934fc3ab6e5ddb21
z651f228f6e63c640a6452bcb60cf84334c6b02d8b3bd076ae36809b0479b8c36919f06386be0c3
z2d6de6d7021bc6c35a84db29d1a652410da05d7656c7942ba70deeb35939ac2909b041bdaf6e49
ze33204a67d6c0857bfcf40a88a17a6bf2f740a67dc6a8a42942b8757339489f133a1f93bfd73c9
z009650b0cab012f55daddd87783f8688a643727d791cfc1c44fdd730f5b55ac2930652de9125f7
zad760a1c17e3499e7024180a9b0cfe57e3ffd6d8d4a4baf7294a5b159d2294280989f7549281f9
zf48a5e4c44ef91bde9474675df67f41f772f296de6b7c247b6c00d79119d70286ace9c552bf94f
zb1f651cd85898b14a6b72ebb22bc479d6b27dce37f07ad30bed21101bcfc88b5981b4be0c6e0a4
z0546798f9fbbc1bb574a7ea28699a6f8953102c34a4e94fceaf3bc7ec7a056a2b894a9f62a12a3
zed4c39ff5d7cb44746aaeb7b22738b2ab8162bbe1eb9b697b65524b3387816749458847190b9d3
z1ef9b0b5b1154c7724e2593d35e8ba9761958f46347b5097a4c8f7dffc1e6c9086969fb256d8a3
z1f376043eb786a41650e0ea9d859cff6bd6ee2e9c7ac9d94d2ece761ef5badb771beebb25be34c
zf566edf71c9ddf10fe5545879ca65e5592eb915da0f1f364bacc323aee29d413de7f0a13d6f220
za69c0eccd2a63c8aef77cb4cf4d846d4e42ff480476db49971d0e13721407b099419130115ce7d
zfae93e8f6fef17bae1f1739eef43e94288c1097738b00e7859c6fd93a0816c56696c27c669f1bb
z2dac64de1e806ca9b6db835e2d4c8fc97ae61d5b9c33bcab4bb75ede2def5c491a38fde65c5b03
zc2cf26d66d262d87c3a932b1730335eda8427f88266725eac4b0f1ed03878a056f831e1d761581
zf163ae5a6062a07bd5e540ebd871d97c1f5850d7c7067f3f26b224c5f585477a1638cfc4e5d523
z0d3fd6b303cf54a9d71bb1cc071165c667be30ba8d606ed54a0b55b351cd6629cc9a117f6c87c2
za1f4429af0ce3e7d73a87a941ad81bf58286738025562f6de4f32efb0c57838ee94382c4966b13
zd55d976cbc86bf0319ded98989ebe5fd547a93f0d02cb7bf8ed506fbcbced3aaf32046218a6141
z9c6598266526983964ee1187afc4196503148e84e480e3104048fc692b9226809e28d7cdd5c0a2
z1d5cdbf677df300df8820248bc3f97c261722dfe44a210680b6a80ab81584cbe98a3eb25c86659
z8a253dd43f0dc62c9574ecb56d9f38a3539d7973de42cfd29405c2ede26c242bea669cc3f43a8f
ze05c38fe86bbc250a3fbb8fe5ba04aea5cdd95176720182c9efeae8dcf1e167ded5a4c44a5da87
z012de503ccc8784466d384bdcc2a059d9b16f67a0ffb834aab89ac31564f5999e2025676dd70b9
z22ca86eb99336c10a815ff2b76594279bab7f4d7ecda1fabe92dcaac303ac93428825b90aaf788
z79e16674f9949643938eb8fbf7e32619499427a1e572bced145b565ed375834b68a74df6c0a771
z4180dbd6ce3bf87c9452047d71dc61680ddcbe6b21b58ed17a83bbe14b3b66c305bb7488d41afe
zd7c706cf934ec735d5795b5b7865a52e377acc4b0f2f8d6cebea14dbc3255282d3bb8b7ccae3d3
z4f89b94bd4ed3e623c1e491ac3ceff1130c98661b7b1dc64a0f1a3d57a9a1b5dc68fa27e11806c
zd7a366f607bed72306a06fccdc3641c05c09e5cfcd6f0d627bebb5cb2069138df64181607136bb
ze1943f8638df86595d0723e9876f5531c4af57ff64727ba48b9c676a29cdbb762a7f266eb5aacb
za3d32bd0033959136eb03a07765fc60781ef7ffedb0ef420307e64cd80553e8dd5db3148a00f03
z512f922094e27cdcd8c70644936c3f39e6c12c7f2bb51d718d171f1d471d4ab8cf3a44d21077d3
z0c40b95af2c4d242f339502f7ed110f7b812a197641a505ae4d84fbd684c829e4dd9234d362645
z59be4d5cdbb52c6ff5508d1362fd9fdd672ac4cdf720c5bea4fa39210be7e60f7cc1ea2353e20e
z2f17eaff1562c57834bf99cd0fae7d3292e10ce881453868cae12516174b738c06513a4d4eea6c
z2a7e9ad522cee199c7386dc21c00985d0df09468ed312251bd6e601319d07d660ec947bc2320be
z2eadbe34cd269516e716b0e331a46a1a12781b779aae1f37650b9d55f9175a911499333a1895a0
ze56c903579c8856809cb00dc386e2b6536ade16fefb7280f6a61ea7f3d0adca223b2a22609544d
z178ba49d969301f0f0839c1d668794c7bd321eaa9d07415d27e65fc93a1e847b81c4cf4144bc64
zb55adde3c045f8cddf3cff0a20293b34fca5bcda296d5bceb2b59e5dd2d88b83155242cd23cc09
zffe897edaf9cd539faaa9507e1b1ac4f266ee6bba70e2156df0a24d0b6829e99b76f2b73d04855
z69ea3bda31aa9404f32b4736cf832c210b65aa1b735720ede3d46c71a086df3b6301e2aed7c5d0
zb54fa99ae9c8294d6f6b61b4564bad0355bc9ab89f8e437b6a86689b6e1ca941039d2c803b8a31
z063777a28e95b1526a6cfe431ac2bf2e43884866a5ed7d22ff6a6dd4224e1f9ea505727b590b78
zbec32d3a54e2b565ffe779f0dd0af127c9b5a95a4f163427959118c1930281b2839fc8e54a8596
z56c53469d5d47b7506e254fb820d91d3dd461206eb28bb5c4d17b515ec5e2e52f7569f1e376881
ze01e7c537f05d594cb02e77b5d63bfb5dd093c134052384abf2dec1673a0f832d14743c3940b46
z5c30be29ec872b43fa48ff2258eddcde0b1e183c20d2b1994cf27520e7c9712ff64de890edcdef
za9caab61efe8c5994671d4e72d0cd882406b08580283224725aab375346f8f64687a2a62969e6b
z8370733529f9a5d1d81401685ad3200c09bd71985aadc41a47a846d8a69dba0f648208d4c6093e
z87e86beaa3748e72b42733b154c4e31fcdb29c55f08b441f0531c04a4e8596f94be1d21b0981a2
z04982e3c69549198a8f22045564b224c4f09f1a36c7fa79a51e9b07b6a7c02878c4f8d0aa99105
zf37182ff2949ce4aa3be4b47eb5150634da83a9e9918a1635878a1133d4773ac052d6473fdfba0
zf24606743da80690967292e446bef0a4e6bd84e0ee81c8f6d22b4e4cd78f88273c96e24bc3e800
zeaaf496bc203b8671cdf43d4824faac5fbbd32a33cb918b56e866e33d8ecf1de5b4e1c979c2770
z6a9345936e01e04fbdf9c6c6668fd611164fc4a1b404a64e38b213ebea2adad48efe46b68987a3
z6c4179ac8f5bb2baf0bc9bd106371d104a0ecd388a91b33fa06b0e08ab6410184e8f3636e608db
zc73ff04154f1173fb2e5aeefba62da5f7549bbeee7d99dae241780b90e703d36935c6a27e47dd1
z70b0a4891fe411fa667cafe378f6b2a6f8d1a2cb69a3f7ed8f8e7467feeb7cbdb4909e06d58af6
zedc6556cb1dbe5b6524b62fc8e50bbe2043a0381ba9ff92af6a2b270d0e628df2c3ec830cfe908
zbff9cc032154ca8034cc520c0904610a6d59de6226e07a504a4db59f7c9c86b78184e71afe58a5
z4e8c0cf66f620776272939bc911886de24a3d8a80814fc83edd1434a406b016c3a705328378050
za768401f39c9f5535c4b35f514a0abeeddf39c261834b7263f6f08b902165426ebabfd3c445692
za59ce724ead8b2f5235dd1085b0af2b64e6faa8b05367f7a30d7dea8ea22958d41306fd5239f9b
z6baf4d5b2bd77cf8a2624a727525aed616858b976ea156d56201c782759c09f70bcd72451dba7d
zdb8a0b5e1a3adc7c92c58dd73f35bac145d3cdfd43c1d4cc118f599429287a09c031d434ed984c
z9d6b4d189742a19d627fdba83ef01544fd14041d767449699d3e6c0ea9c43611d4a5b2a6c123be
za9e3581baef7bc2a75ac0caf103902974ec8b9bac279f0b174a21ddcc5a53302c4020b12dd1e34
z5c9bf1516feab850c421803c5fd246bc74ac0b79b37e154f8e8cd92589be1b6cf04e7ae563a4f5
z450dc418b8e0010bebd578b6ae071537e4ef761ce088f1ac3693d1c56d3a40dc9662c74d1abdfa
z3fb35a8eef5227778acce31d4a5b8f740a7b060ca32c348d6cd3c9929f28a1d613d0d21e089673
ze6deab19b54ca7241dc459d784b9f80cedbc94d22a05677938e9e2cf26df9b0eb38c4358e47d91
z3696953bd357c587c2c51820fed0018e5037ce4709318c94289205acd27aa39d857a9e50ced883
zd6f79c94401785f5f1e3132d5cbefb91f20742878b016ed1792c27fd577bc0decd887efa43459a
zfc464b52e75751279f3d539b69b16839712ad483fbf95bd0ae6dfda767f066242d42679ae85094
zf38f79cb3d8d814cb9033ee0920640d531955e146b130d50a2e5f8cfd85520a1b388e0baa7098d
z319f2d303a24357a00275525e03ed2d79a2080d472aa30cbf70f161395519b3239e1f360ce185f
z3dd9bc207dfb4d8af13aa4096efbba65b3b20709eecb77a69868135fc4be238e64d8c000d9159f
z92e06e47a83d044df9e92f765659e80639db38efaab901ab35beee869c46b622274b02f1fbc59b
ze88ddc1a8cae9af1a5305969088ef34aba630879af76e3862cef8db9a36c9d9d08dd0dd3efff99
z162355605fe4b6080a2ffb2ef5fc938a8a62280f0674ab3d94a68a340fa452e4ce1b7d198b042b
ze88017efae61fdaa9ff118ec79a8b694c0445c35ca4ea85688d4fdf301b1176bf2bb0c88fc6020
zd9382926c800408ff01b656d35a57f4224c8b872b1c068c3b90e68b4e4c2aeeb3c7cf9e40606d2
zac1f2484d4447f1e3037a463c2422ecb717bb8a877ce1e55df0bece66440010a1e214a9f3ef323
zc94a49b9ca0e27a0e45c6f308c72baf230e50270e8af629e975b328fb8de29761912c4c6929770
zeecb81d70f789b1dbee3a6709705bda621cf06fdbb44e479e17d13776440ba7ffa57c336ca694e
z3a08b21f98b91fd28f4736b588709f9f64c6026b5e7531380781716ff5233fc1d5ad447597a350
zf21e2cf1f7c5b9c15c052c8451864e241d7f255129d77ba52bed5482396084bfe06afc6f93ffd3
zca4946c04726c25f27a2e4ba8012d42895b6261da8631ae9ca892967c13bfef09489e4c630e231
z4eeb815bb83da834044ed5abbd83df22af408df5ab27e79ee732f3e5ae37b9676d42786612042a
zba7f2742a79283f8b829f20e6013dfefa96fc41dda3bb7c036b64dc6f80e8bb273996b8991bb57
ze8d90db72a1952ffcd56c494738f07e1f7df47c16ca62b38744b5a147539435d0dcab5ec52b138
zcaa7337f089042e0b6f7079e4b7b598df54b1fbb08e940037235643e15ce9802e3538e5c7ffefc
zbfeb29690b344d6a9ad40d8b8e4d1982c45f44cf28ec72f52fe64517e62eff58cad536ecbe8f19
z659df389cf0c21cb0d2f553adb7d22e7b95a0410439b13993dcc841ac0ca86b5d853cae6d2684c
zb8956fbc114c8cc06b2c656ab85b701f75b95c680c2d83d2fbcad834779bdfa5a10ce6c6c8675f
zd34fd6d2117c63f8bb2af3ad097b3a9f0bec364c814b492ba37f21f553d95dfa218e8917149310
za3b9b6ccf2743888d255677e1ecca6187bb41696933efa7c0b572ca66038f4614dd31f7566583e
zc103e03e78d8b71600c0d7f83c08f7bc50d185a48b8472fceec2896c541fb6117c3681458ffa22
zb63f267af803997528959a6f9d0c2533521fe2ac194c2814e8668e501806dce4d0f09d355c7951
zd14fa0bd760ce0e237650909ab7595996947db166b7ec364917422330e95e9f69a835906cfb1f8
z65a8a759de0d330eacadd7bf87246bb51b1259f9da6ea5606981fbf8d3502bdc9691782ca59338
z099535dd7db6231fad5fbe28d0477e696b0c491a4978698135ab4ecb28b9d731a00df7a7afa73d
z535666c7190bbc73eb92ff8e148365368c36a720d3531cf08613b970fa1829c69491723a4da2bf
z0f8e6744cf6cca060e69779339d6670add8ca6ea9b31cbb47cfbbc28a5253534c708b472407725
z59771b17840582a7c07c4e5a7ef0cdd408fa08c278c6776669a25abb17d654d3a7c16e5bd590bf
zd35e6d2b46ce23b3a8d1c1adf57b24a0164838c3b0bb2d73d649fc30c0973db7c1ca1e47a4b2d2
z5739fb7ee33a902391031dde2941df6533ff9da1c7d1379fccb04a56d6681068e112f527321608
z729aefffc4ff3ee8247f6d6ae7105b189ab84d01548c5164ea0c21d7c742725f055b517b24240d
z488a9a5d5ed091bc11a8084c15cabd28acb390538ce7c014f24c8014a7cbaecde08dfb7ea7d309
z748a2fdd9aeab278188f9ae25f74459167dfa03b3d523d8647833e399977e34ee82bf42fb62f67
z7cf8c22a25aa09778ea8ba5d47f823480a8a2f8c729ed3a121fc36714d478439e6bcc64c4996d4
z4cd0e57c1e15e8d3a82c16af902b52e09338dc2ca96d9553aa83f31a4764ee0246b4f7863e69a0
zea30e2a04ad015987f89467d18a7c9c9d73fa4df65deb5353262b1f64cc0664cd476a01dd5e9ae
z7308180be33d4a26d4376ea0e389b4d61c34fd458342be22386360aacfb7d21b3aebc50ac1c9ff
zcfca056fb0fa236dda1efa7b6b7951b2f9b0eafda3818165af605f660f9ec69f8c788ec493aee3
z4f15070640c7adc1de771e2ef3b27a90f3faf526205bea09c8ad4c1871a68eb25dc9a33922e35b
z1ce091b479054ad4082ff801b488011abf345cbb30c280a726369ad2af4b6a864eb63dc4fee7d2
z9cd381f1999b8f066f5e3411ab079ef9e8703f6ce543ee1aa30a847463e6f4b8d1352fa0bd0d12
zd10d1715e004f38304c592aa4e0351c5c996ba5568e8d2ed0cb0ad27275d31a9c2a4c923aafe8c
zf95862aa7295617ae596410f15b6ef396768a455eacbda53ff4cbed0b38f07d9bcf460503f44b0
z4e922bb4bea360ae6f699f4e42178abf56f347f756382c99ecd4b6715e69a64933dbfb89f078eb
z0f22fdd9fc6da0cf35fc6716cc3c90e467c9257ecdeadbd146d63bfc4249979a91b9f46b4ff6b9
z4fb4d482fe17cddc6d5f663e103088b95ae64d7730a3e9759334ddabe39664d17d594d6d933d9d
z9ac2f2211226f2a2cb903a6ff784c6f1dc18f2eac0543a5933ab975fa47f207f89c930792a948b
zee94dd6dc5bbde856b16064f066933e9e4f51a97abb522c69a60dfb34f7d590df9e78d3ef66742
z16835d00f1d30fbbf378345c16b29a04cbb86bd711fc45792d609af06e9db2956d5d88d4428066
za492d981f0de63155717d7941637ef87cb01429e090573b8c53785723ea21dffff9b6c827d760c
z20a18b2fc227b60768affd30e2e6584cab1dbd9b99fa8138bd50a1a7eefe368c554bf433dabedc
z521f13d3a487c3717256663d08cf1fc1a2eaa86430314b129f830d0f274061a09e487640715b93
zed4ffa2d05eff308f2ca1ac2406a903bf79fac3e50a18a5d76ea419cb57f45e17ea84ed2a94c61
z9b8cb3f89231b38116500778a25522c7f547b4c08123bb0321db2d7b2f6582e95a809a60641532
z2b47400ff7bec4e5de1fcc1fb3b83f1487febedd291269d75db80360dce627692ff9218ddf2a6d
z706ab8c256d2edc3e1adf8a113719a1fc648eb7ac5ee817808f59071123dacae732c5615204ac3
z437d193c5d736192f8eec3535e6c0dd91a612a0209be6d720924935dfce5d6c2a87b67876801f1
z6b2fbff7c5e7e27a6329a0bb7aca69cb8c603f0a821f6cef5e39971ca16ccba6e9d54f5915a276
z7abb946555596f9212d6bb9e3f283543639e67f8be8ce4056f176910547096a884902e8fafd91a
z7f72092da185b985c8f2d95211c2d1310290a21c5c849c418e546ff5efdc21ec3a3e58f192c351
z96a0eb58faa5cf8c0a8e813a6a4b1570276419b1945fecbb82a0f65c4ade085a6ad5d66177df7c
z92e6ab0963ed430df8f650ab0fffcdea7c71e35d56e27ddfc5c9082f198df37f6100fd1963cc03
z6a27e1f34eaec8178135a9909d49fb9a995c5650037a6b918ec7946c95fc2838ed562d5c0809d2
z7f35eb89f91d666416dd54a0bad2cf924e256ff81b11e9c3d2410fa9e2a7dc576068c5d438219d
z70655eb9635c21aa2c502b6ef03b71fa05c205a7f3fb57230a5a27faa711fb90dbd6efb5f9aba6
zae6f06a137e7d72c083d59241db1da93f09c7790e34de2a82633beaa179cfd3627854f0cb66d6d
zeb3133627d797fdb35c87bd7a0f3af527050a592da422a99c7b569b5e237517826e7af622e54bb
ze229aa5762f43e3b665290a53b47e7640f7299803a5deee2519cbaf8fb7053e24e2f7453d84b28
z8a4337cd76dc928b0efe6855b285e0798b299b54d647408251b0c9359aa301d0cd52ed46a91fb7
zd1f231d3d0e824e07ca072ea3c90215683e17d6ef42bebcd3cabff38157d8c562d5b4fc5715cfa
z4d129c1bab6c7c1f2d777c88c45105817585c56b34d7b2298336d48f85a10a7da2b6b17d861ae4
ze9e01d002cd9e29166aa5bbc0cb95cc47a7600fb933c98a0ecf86c2a423a116eee5e118a186c56
z6f2d3cdb621b63776106e5555a60d21f4445da10b8f327a3eecd34bf74b0e5b810693648cf10ca
z70bd7d6cb38458f51e78de083e83096cf5faec0e015a514d282192e2d7e2c8ffb9c57ad8026042
z898152e328e44bfe87564637e710f949033cf6356086df01cf256d886807b78bceb6967e11d51f
z4990ec0e78e6353e254d94f3b1cb3cc7942abbadf975eb343ba63e83145806894e735bc81a2f29
z2674464d04921cb58f8cf0e37588671945492e051e4de4c8b16124ebda33de8eeffc9476acc79b
za2cc7f78509f42641d602bbb7b9cbbb619ad6e53e9ba8feba1537027ea431c91ff0889254a1e42
z689f165dd8a941a0e25c463b24b9effbb993ac9acad484c646928d7372b5744924185d9e5f84d1
z5c7d795bfbc7f8b6699cbaf3c343f4fdc0f023b1da0a8a33af76ff3fefeb7ae202113127fdc3e9
z55e5c684cac857311415fc5449b7ce95b3bdd7dbdd7339da21e196280af03c46d63447dd87097b
zd063a760dc2828c93f53b7fe861b3227e15a5be01a2cf87853564a3db28f7a597b8b9a3c319aaa
zb3af87018add7fdd11530cb09dbdbb84ffa22a5d95cb51f7a1ea6e7573da45c0b230692e148833
zd7f5de5611a295cb3c30885ba1a32c322622be0b15a679033fba8168d58ca41458ed551edc761b
z9d7ed7081766935ff8ed847e39e7d13e4db5005ab022054202a6cd33c0d26575857d16873b5faa
z2daf4c09b3c78f7b16bcb2e3a1bf2349e444edf70d5565cbfcabc77864df7e0d8309ea03a5fa10
zd68396f43766cd7fbf951377936c20866dbb5ae7999e436f812146bce0edcb66c5a88a31729459
zb18e6079a9a3b2aae5b735a11755011b6973e50512da1686b8f7adba9d78a11048596bac249005
z9413ec6bf56fdd61d6332ccf65a3006644b35db1220ad433c7265ec242486101215bf074a2b1ba
z3971c7b99f9e87dc20905760f7d5adf75e1b27da21b3fac13811625de06efdd593955b2c70f271
z8605cb12ff522457b4a6b9756d6e84decc5357f74cb596327d19e93fff13db411f1724201c6efc
zea9dd342be22f4f54765b32abe1b9acf92d5ea8d8a53770bafb81fb0c611f9c1dde426ca155feb
zd4839be4128d267393f5eb3d195b69b2c20676e91b8b53b5375936ff039951ab376e07be6d2164
zdeaa6d0f8f5bdee2a8688fbedfad5ab1ce9d78b0ec6c067e438eede52f9171eae4b33375faf93d
zd6d11b98b82f39dbd6048e0aaca7ea13955e90ce785732f8568daefd853a97eb927dae35ca0490
z4a08770c69d670547d18f859d3b810e288f5c77fdf928d01418bcf7cc06b93643f0e79ef0e8a8d
zc4eda86cc67e0bb8a39bd06e71058975f08fbec6e156a81cdee649b23e0fbbdffac0984d49bdb3
zbe8c6ea1a2a32706c4127b90cd0c1c6f217ac25a8e7327d4de56ec71e1054be6df39590aef081f
z7ebf8d091f5ffd3b9a361c21026460da52f058d7c2845f5d9a071853bca2883340589f151dc12d
z2da89bf346c019c4fb281d398e42dd7ff6c56e9c0177e2b20fcab7036647cc33936ccb2892a413
z8bea4e9faf3e1c230fe3cb1a64ba2feabd55d63499073c65b52c60c815c62daf0e3a66ac07fb9a
zb56d42bb1e8cd730253c2ce614d0ff2553d6b1bf4d57a313e220dd981c9bd38e426d2dcceb1051
zc28a84ae6b09b3568ea7997c38aaad8003349ab1d37d944971983bc60dbfab9b82a9f938b8fb68
z9439139d834037abd2d26b275b4c209d0efd022b1a69700537bfde9e915d9e9f5185f92c7cf16d
z316fd3f18626018134d3ff7e3e0e0480d3929135c4b15d965b1081b44aaccad86b3fb5eabcf73f
zbd63d937d47c19f71d5e4723f47c6713f2e465813f8f0da1acf1e330609e6e5769fcf62193d32d
z9f484065d7efe64cd9e313324b6015a207eabe57843870443654c0a3aaeaa1ac4025ce7a53a3a6
z8bec2f1df70eef45e7f805e9725b6aa89342ef1679ae93a8b43c8a9a60425e53cd0b2c5fb3931e
z9682005cc6600bb39a56f3aadddbc68fc1f740a2c2aaf35987bdba20f9283730b2f2654ede324a
zb5ee9ded7d67f7cee3d80885aae35af1721591462e1ea94d163efe03604251e19492c5b16c9f1f
zda976305521732916fe754543f4be68a85b3ed13b4935131f1a670d13d12e80ec786aa2c90f1b5
zb7397e75df8e5030c51761e4f6481fb5523f837a6812d218958646183057849106ef88260990e0
zc95c407c210364fd99649e52f963b6200bb9222b01b7844282720f863e853e13f637301604b4a3
z52403bc53667a13041670c5f66aec25b04646f8ba509e5ce170186d493b6eae7b28a8b19a75fee
z63e461595b57a99002f426065262837331b2b7abd1f24c2f7e6354361d6d8a6978e5858d189ed6
z4990f937cfe95dca0735e6496d3aad6f870ff62658279e1cf8b4905c7fef3fafc2eab2d2c4e9df
z207ca452fb62a6af201353dd95c3efb893ff7f67ea2604eaf7dedad44eddb37e6285253ec06882
zbe0f7c7d1108a939ae4e885cd1bfe3516b746f68b59466b013e2d75eb10ae65947bd236a07670a
zff075abd65b78db57208986ec6c75700c776d0e53204f9632ef14805813e4d41057fa9ede3ccd8
zc0b1e1c37e02a7d760019ab0c925ba813f79eb42d0d6951d7d3f6bd98d8987fc0d9092c59c1363
z8c8e919f5beb7f2f6ba8d484cdb32b78fe4160b0fafd0bd706cd55b8aae9fcbe62a861ede57599
z6ee23c5ce747e226e143e74fbd67f11182a5cff2e6343e2c2b3e447bab1fa70fb7837ad335b368
z387f45982ed35a963bd65ac85262fed436ff54b9ce8ddf52528d46b8b64c5986e7d19a99aa8c7b
z071cc75b95edc62c1d400658f83def8b358c32a51215bb72516ee12c6c25fc8ad879313ee9d054
zd80d385a3d538eabf0a5685a5d68061917798125998404598cfe5cd47862122ca2bb91781aa62d
z5b1be5d8b56f10d9f1ed1a9701b5b1131f0fd5c972f0a6cd9a2a477206d4c70c8a5a45135c4f3c
z3bfc794fd9d3751a833d1081b7d2a651a7f5988d5fc1a7136063317d884e571d17e772611ee1cb
zceeb1926a52af45f083df6b531efd6e201ad22816bb4f757db7dba3dc1cc5d605c2abe5148e1d0
z08ac7dbe9f676a8d328c762002e8a5e93791e7974173f8721b71d93de9eb8e4449ac30ec7632ab
zf545f2c63b0bb1c1687fe8ce6301376290708975229f23e0f91fbf07a4a3cf06f6deec58b192b4
zd520a3f4463865d42722fa8cfa4fcde8ef3dd5e906842a862ce894806be66a9310c94a41295e0d
z5a222283432045dbea7b11ba38a6c9fff42a01575bcde9ea5371d7fd928e4c7b1e51737a6a17c2
z702ce78ba14a6d5b22495d0fa87d2cf82de68ae35e896a9d60907d835901d2a0add00a64586e17
zeaec40b026a7d37a915d7809974b73b9b4b0de0f3a398d6e880bb83a35f293aa37ad420f1b710f
z4fd1ac5e22be3052510e249b3284820ca80c93e2f7445167b71fda9c74c3a35c3d27d688ffa555
ze4eb9c21f453b1b6074f597dfd254739d8f30806a93f9024ff08eb00c92b9fa53335ebd3c8ab9d
zfe41977ee8ac8a07ae0b991aab2e129d6fd20a6f1e7fedbb6013a8d2da2f2617e9965ce8e3e030
z1fa392f36898b85cc420e2c1daf2c0396e48c7649d43712e18cbc0077a5e603ca3bbff533cfda6
z4ac817b67a6c24be052d8cdd360a3d1618fef274f8de7e718cf5506453bd3c3415d773d35924b0
z1353258e4f441b9e9da70db2c4b1d138a16046102e5503714b3e5d1df5b3e734078b17764978b6
z4b661e2cfa8f24bc2a4ddf64ae561f267a7988c4ad83788f2daf40874a0173d6524c43cf43987d
za55a9a85090b3bdf133650c6d23d799f44b69fecf5a023544a92c56b79e7312f8ba8f634e8ab04
z50a59fb82ad63624238a99c072fb7901f9e5895d1477969dec606728077816a7e40a6f9ebffd80
z24d7426df2b2f9f7775c8ecd34f1d78e874f3cb2bee7d556f044931ca8d090d3d72205b7ac4ace
z473fea4ea13bf23d2966133cdca07185242d2813a4d8e279c67e504d384f3d91d23a7595bd753b
z20cd809b0d2d1498891a1e2a303448cffcc0ccbbff6e730fa17c2fbcc7e0275c1973529bbeb137
z516760d3912b7fe1a93b583e1b1889ab2b8a274ea3ed1b52ced67d1671735771e42743b3b021ff
z5a4cd31b0a501aea62c025a023e2ae10afe764d8df8b03391401cdb939406f56e66e4553ec2668
z4d24c03fbe5a8fa3c49cafe11e4b3d152d9ecf00b6a422e332ee0ecf2cb8c7a9624e72dcf4dffd
zce46628e81b4cc61c27d8ebaeca7293c4339c1729912620f1302c492c87821dc9dea95d833ea44
z4b9b5151c2a5adc7c16f4411ab82cb6749d677ca5654e8e63e4789b077e4f74f3bdde5470daa2a
z3de8e68afe5dde21cebbd79b3a707b3ced30755a45d3961a096713acc5e9be032aeccb5c8c417c
zb7137e4bb429a33863327e90890486cf8354a592a96081889f956bc6894441668623de441de019
z5e74d24f86b31d29eabc53441574dedb7232c63770fa39d6c76255636b43da5ea1d7847851570e
z9a1891a228d7fc71ceb94fba50b28079815af99a2f59a3d5908ceb6fd761a8a78f6c2440960870
z9c3a7f3f702ff274caee07b672c06599afd6ab00398a34a5b28563858a15dd5016c95c1f3b4dd1
z117c80d38f49dc96c2ffb339439fb9dca6620b3be3c1cf37733915bd854906a69306a053656302
z15c1424f3f696a847fbc1b51633242c4e77b2728fa2b2a931d53bd24ec895aedcd41f89eb042d7
z40c08278fb03d6b8c15da6c4b50a386c38a9f63c885e6f10db00595a70b1c97f75a5757f1ae04f
z74e4a5bbc104b384596998a929ad23d61d5dadb2a3d874bbb080420036f4714c7f5cc08c681eab
z6e5de54ff6cc40fa40ce86c37cc1dbd09abcb44535549d6e02cd43f98dbe317fee26fac1e1d719
z1aede251b375decaab1fb1ca890f8e9e553331b033ae36e54f51131eda13bcf61f3e078a105b58
zbe0806496cecfaab4a516b696bee507fbf5cac36d36db3eab43d539f3758bba08cd612ebdc312a
zdd03e456fd18b63d182479b436f961fcb3b9a058b933d3475deb2ad4dd06afd664e53e411e9fd5
za6d0330ea80879b52be93fb2b770ff6da8240007c98398f1a4757d7685505cda3a92a4f135f17a
zb194551e271cd15d0708964c7af120fc1a84323ecaf079c908f11babbc4176ed55aa780bf014ba
zea6dee51c09550f8941afd031b91892d8b79657f331a7251ce73f48a63d5478559ff888a21c6ef
ze579402d2f268b90c028313361e2b3ca846cd8558b269a70d78fc9c32dffdee125dcc53887ff5e
z3165b6506626ac1534e8a1044d1ff4e99c682dd518f2ed9ab9272f836cd95faef8c755408385ea
z731b0a4c886ad1fd06c8b5036b5c044fa6eed1ad948aa5e046dc8e53ce014adbbc185c186d4d37
z8f793d38b2490239aa1763b6f19d1df68dcfc023156ead08989d0d55c1e88dee8b58b256d28cc8
z33ed7a9509fc5ab79ac64034b4f2a1cdcaf3047451297e80f15dd05a7e431f1a42946041c093dc
zcaa1c84ffe1ef74b189e8fbe46594c2a63da97062f60aa59fc0b4dddad7e513715302f4a5a7671
z9b383b45004a74f75259023ccd56a23a1889625039967a255afe0ee272d946d47398bb9db4782a
z1e34db0d10c4dfcdff054e8312d1410a27c679a0656a4c7dad076352527e7c47f082644d9db075
zdfe38dba564d5b102bcd898669699492b4f459d3f0ecbd263e2d925979961081e9a48ee86f0d66
z22f3c2b920fb40319e6ed92084caeea93b530961a99b43d617c362e337913808c4dbf042bfed6a
zcf70a48e65877b51817f2ea94863b7e05fea1bb2427326c21e2c3095fda193daceacc4e621ed94
z23a14fd743eeb0413f1239067df456d427ffde7b3638d219194de34e763b2ec6a864d522c99f99
zcf14509ca898eb3f59e36b5eaba28731654a0dba1bb252e34035d8e45abe0bec5fb9efed39900f
z42ac69be26bab8c87211a696bee9bb6b140450b7435c3308f15e6379921093285bbec111798c83
za9842fce840a9fa0a02f2d15fd466c7ca8851ef88b4c990bed77533b16fe58d7d7be1905e645f2
ze7f7467408df84af6e36e4354a27ea2e3dc25a299df495e9e7895fde56d89bfd546d94cdbf0fdd
zf730d5661a876bada7f8a591fbc968c4c2ab29bca3cb3c75ae960860423fd8a6604f7704a8efe7
zb801bce11ff71d8b3e3a07a19f9ad80f79bce3d32f339443b48fba24bae4608c86ebb700124c9e
ze7d5be493750b707fe806de4124e303ff7ef458b1335888fbb744c05d4c4dcf54601674b17f658
z6ac4e41f68d445da1c568d0afa40479d5a499279eebfce0a876f443fc1ab77676ac979820bdc91
z088729becbd4607719b9fa56322b86eebb3875585b237f4b7d0265b13a78d2a0821d50abb36f1e
z041d22c4fd3b2fb3ad477357a863fe9946185d3ec938a49143540522d1eea9231b773b87191b1d
zf3237f014cd1445bc38a8289eb4acf2c431097d1978a1db108809519b9d5ff1a15b111b1274d6f
zc6a3ddb36dbec83a898efb976de84658bd1e668059eca4080a8944a4f1eb0af69a88ce8bf94307
zc14b9c2686507242aa81b7d377f7055656edae15880f3a34c28732a5b661bf04b1213f607a7006
z89965124baac300aa4ba8226ba91409aa07897570f20944881d89f00c5c70ffe4add54ed3421e2
zb424a416b330dbd916330159b28b77aa7361dff94d341c02b5b342a0a40330ae69c60ae2793a59
z914ced51fc71a49b699d277cbebc15e9e92dcd7f10d60e487cc703c147e44e716ef3c2f2892278
z997957408324a163864e4cb8557c40398c319c4fce010399e86215fa4f2b74c4345d8dd1584840
z42bf3729b094076a2a5c6d733f80c90dae2daa4f968aa8da8fdc172ce8b66d2e282b9d20acc262
zba7894625b4fc6d2759af7b797d00e3cd718e366255a493c6308eb1a72af673d17e798b61af63e
za5ebc2d274413ffa5c4dfbe7b01e5c68ab51e12c2c0aaa5a4ba4eda419b28fb334fd8a42b3c444
z8d97dbf28f870991cba12786de20770e9409abc70ba563ee6fb7166d2d95042f694f3e1cff667f
z99b0940159af1efcd706a57f36b2778aab37471a522a2125da9f840b6178851aadbf9ff35cdfd9
za65e56bc3d037cc69ca09d3f710d6dfea7292e220f6787254ccc213c68b869c050a432c6c53024
z598b74673071e76455739cbf31bcd8d35c21c35659130261acca8d601fc67a76dc3898e4f1924a
z1bdbf6c85ea8b4d333c6045fdf2aba3b77394478dedf12ba245371fd6abf11f120b3090d0d8487
z49943c4412e0ca373118b9767f419a74b7e8934dece7157bcadfc2a8e080cd96c5f81c00b22207
zcf610779c11871d9ed4793d2acf4a54c54157aebdf11dac9fc9426b8c3514ea8f4f1c37218cf12
z76162166d4418aa545e28cb24a46692f7282c449cc1ee9355606dc93e86c7e18922e3f91867f99
zfc3a2c1221ceecea2e6ae7bb1d4ee868b78283d11b7d1d411c648d5b1cf0e860d81e2476aa8a1e
zea28ce685bc1702351519e80f6d5d0cc308ed0606bfb740a4ebeb68e2789c13567a1553707fcb6
z300836a0cd6dc12cf5151bfdc680faace149f3c1530c3ee9f0e474d51c06197354c3fcf9f2c372
z23c5b1f4e13ecc8ca6fd0b013b33064f9eb9abf28ba7df243a9944b70bb79891012e4d09972f70
z5946b12a657b6e51136aa691224714b6155eae453f2d21d0d9a88aed1f0754c894c70af7103560
z6a8184af7316125092655782e8dfbcb3f1b1f83577be65b7dd7465970028fa677181460ad56066
z2dae27784753f18289d24a0759d4770f0a5ad86b58f4feb09df85a67e7fdd2626feaaf20454835
ze9fed27a3e07d52cebe08d5cfdffaf032fe612aa6eb0e7033b6d743db7d5d25a321ecc253f9ec4
zea389e4375444c552b4cd49c30aba513c8a319ebe5788f5dd7a68ba757c76d12d72c48b1986306
z3575de609bbe169d20e9669aba335092b39b3e518340b7f9480e8c53f32a7bd4749ffe0755b45f
z09f42571be9704b0a5b7921823c39314657cec6aec456c41975d21912b554589eb61aa935ab5b7
zdc584acfbd481ec348241c60cb101a47bc7bf0a2abe9cfc3271a67a88c9fef707dbb16a6825241
z8829f1d432d0825acaaa542fda38ea657fd435489feb9da7403535c8d0af6270504f9b06ca60ab
zc4a1816e76855f812c27f39263faa8dba051de506c4097cd5d8150292b8b9bd8bd69dc2ab4bde8
z0c22175f1ae6fdbe00376b9205e467c1703687eaf6ce0530751a05c7e56db27912ecd1db8d80e6
z2cd52a2aa8066361700d5cc1b26b89de49c0addb1d7b8c0cc4d8779d6740a75c18a4babf068418
z06106ceaa51088ac4a7ccd8d83977d831fa84ef42991f10b01b49297bfa010390a24912ab29477
za10647acdd6a38b425bdf5563a4dcc1031c4b90054b713e842a6fc7c3601dee58da36344abd1df
z47272991d4f0cc576b291e9ea8f6f1e1e000cf67266a2b31bf5b0666e392940ef63d7ab9d1539a
z20388ea87771ba2528facff85bb62ee18bd843ec553addc60b81a4f7ef351f65575a8a0acc8281
zf0c6462b2db4bf1c60cf94c563782c93641b83b8ec9e4539c8f81245b883a6108a90375873cc93
zd66771a694faf962865a557f7cff608dbafeed97044333b196410b8139cd35b13e4930437e8a6a
z8e8ca4198df3938649bc68ce53d8cc4908e5ae4975f81b0b1934d70d80a1f9c040c8b726a5a06d
z58ddddd5c0306ca0553717a2539999c123442530c75061c3f5ba6ad285f38ff31666c640cbaa2c
zace663d3de350438a3700e3d1244a9c921261e56beac403a8ef46d3d8a41990fbc1c18a0dfc55a
z124be0acc760c67e0ee574ab4c646f745b0a4f894fef28dbe6516bb4090a0ce17bdc057a04adc8
z7fd8a2f2349b091adc8010fc95af59fe87fe438098b0d307894fba73bcb644ce12e73cdc3bfa19
z5fa7b1ec337b71b90d65aff37b15de04551bd53650085dfac87c0bca51e39044d3556e40fd97a8
z1e01cc38e71fd2eb05b9dd5ab4859ec8a62ab30c886c2895e475b6b083820073dce369634ceb7d
z7b3489c530bc584024e1071d2d2bbf6eec444335d042efe2f3dff894668de66647558d8be94a36
zab3a95900f3d79746edb4584dc2f7aba482c03b1a8392aafa0a526b5d7689ff28c1b2f6adc3327
z2d1fa70f435171d2c77f351ab3f929f67291997f3f52291b81c2ce01b61156411d84fc862cb868
zd8ea7164e146ce827443fa33fbebabac063eea1d1be9868872a1c2085fd9ad11fd84980fd499c2
ze4042af5a319beb0a8a83b9706483824cb6e001844d3c4ac7b74653e47b349925c5c21f94b6ee3
zf137981a8c6b6500a17b70a9d62f3632f88e063d2dcf8b0b977781af931f6dfea1bfc252e21620
zf9dcdb9f249ffa521ee0b66488bcac46fbbcda3ab47041d220fb0e67b11eb706f28eca2aea5490
z6c59e0fbba7a9ba7394e237690dc950f5dc0dbf8a0b00f724265642ff987283f5a100d34f0c0f4
z4b9a913b533855a1d3f31cf07a024e0760c05692f23fe8a1e9b25c16db8429bccf4582744c2523
z02db4981c63e75d33613fa84b30d2d490fd8703caab138c31c43cb9a1f3dbf2d9f49b9bfaa10d9
z496e57a8df51112d864a308cf3ed76156b5b480d9563f4463bc2bd23e7408484596fedda801d24
z2aad453ff3cb18044895aea34b03854943282e9d946efbb4d750117b7c8cdd8157c93ad5f0fcb9
zaea3483fd8b5ab62f6c53f32e001c1dc1b79f5733e10d97427df03a79f1fed925ad607fec13a45
z7ec57a989bb8c559c69a2e064d0fca3862c52d51469161236b23150513c6e47fbdd9d4d052c9b7
z8a21c545663509166b43c7c4468243d33812c28951d15fe3fb4d0ec8f1f4e7a66da1776c52c495
z25671bb00e326ec1969307085de6e2e50e4f8fb994e8696beaafe583a9be1864b0a14fec62b4f7
z585a9058edaf32c00435196ae4cc4912b629e0dc2c1a685011042cba67dc76ac2badf989e81d2d
z5dbe8df471dd37d587a20710c0a9910908ef022e01fcf389cdb04ad1c039ad5cd0d6edccc0d854
zb21c4ab2b01533011c879cb8dd164ee6c54fab93827ff777eb76d8a2167f4dfc6ee7c40bec8d98
z96986a7eb74da5a91861ed47004f970515814995ba5956c095bf8a306c41d73a7e3f769b71b368
ze633865540883d462b6d43b5d7894eab7ba19871740a4a15a1fac9b84e0be62378b06e603faafc
z47e8c0dd99dfb1c41738bbb8edbd4a277b03572a5922e96b92404c269acefb964a840d50aeac7b
z69408256af26d1afe857dcfa6327aabc7d7cd08e3eba57ed7bebc3827f82344f1e5f1d566c5ede
zd0d3ae3181c451a956e50a382f2ec8e6d09fe58cd6e56121cc6fadcc5989648ab15754afda89ab
za54e79ee162b8558a5ab1a2a27bc59048732febb75d3c216ead9643bfd462c0b6f1e24eb77d955
z9800fbfb75c00a0fe7b8f233a0616c922ee404a089d21e725875e1c44ed33028e124f3d5351f34
z1784cae9f73b411f48f1a79024d7ba378f459aee03bdd873941d48f15072e41cb1730e3bcfd531
z6256d03efb6babe852105aeb2b00a0550b1f558149ded3905157bb081dbb2451aa020c825282e3
zdeb5440c57fbbd18d0b667a82ee0cdbbf28285892ab3511c46f66c93e9ab3dc173eee5623f6508
z0ead28dcea929492ff9e0bb434b8e504af7a356c130447a92551151cf6bbfd8c4a3ff644706f9e
z8c84667196b772b08449c40385b98e5a53a71dff4d8a75b7cc784b485aa948f03f52b2c8859b06
z583b71f2c841cf45b1513036750f78a3abb8f3e876de7edc83bd4552460b0f03854cc1e4a80862
z5db61ac5a5cf72024d859a0d0d5fcc8883e95abc014ded01bbe3fa2f1ae6ac59a7c450de63a687
z37ec0fb56821ef46c3737730d2c16acec6b18524f8609f28ea684417c3fa6322f4b95ca5759d2d
z82444bf2e5702577a685c31682c133769b40c4ffd03e96e0d05e33bc2f4ccbeb2fbfd5033317cc
z14778cf03b1b297f7ca2f7c8ea28b4979ebc52314e322aec866a32c0a3f0f738c83d11d0f7a8f8
z8b54625b83901cac252a782877551347a07766cff719f3f7fdb2977c5ed349d5353314745d6246
zbf1fed9a199f1dd57e80bc6bf3087341f27208935eea197ef7de9b63e730e58b8ccf1af3e10576
z58c9fc3c3361c7c2042bf937e81bf2a18119fd8fcac4febe36edb73c5ec404b3067d4b0ed9309f
zc58569956165a61a551c567035200fc160da50a57ee2baf249d100ea695a972751adb7fb5682b9
z08a789626c30220349966d9b7f0646eff8a0d6677162b18680e80828d7075ceedcc89d11df7ec1
z982b4f0b403eb864058215b3b4dc853d570404c857bc05f1b72bcae2added4b49014dd3e93b9a1
z4dbfdaf125200841c8664137e1a29efb78a6ceccf1e888e2b4a807a1a81a19d93af0a25a91196e
z46ec83d75b3de488c02dbf7db928b6299f049214f2d7eedfcc2480fabd924e69c564e2d6dcb961
za591b0508ade40981ded45494f9db98392f818e45871f8e35ce21d6c559545711467d6acf34fd3
zc6e72a699fc4e5b0f28bdf0ee9b92f95345f087fe1c6f7a814bbcba0e9586508b47daa0e84e393
zc92138da49e40e5da066dca92ac4880c485a265bb3b9c348cf89e25bff8fe0d101fa4b211ee2c6
z8c7280dc865063a0afc042edf91e91bea14075d6264ef11b4c3497044c3df49e674d2609d5acab
z73a309569153e0605b9e8f6572723c30e4fdc59c3c0c99f4bd545c9e2f171fe3f73bf7d8be3548
z0f58b11a0bfb7acf32576dced32d5cb9863e89e7757b3bd32be1c7b24e7f3d5040b9560f24e21d
zbe026c229f130b2d9f0de9a1d589f8a0871563232f19a6a03ebfdfe936fa288e5efeaa7771f51c
ze7f2bc164167ca9e306312424f14d190ac2b06eb57af027c7de045000e187f3d9bb75f47e191f1
zd5d24cba7795406256094d7767f3e58df2c6dfa15c0a8495ceaceb025280ae2c3a22d79ed9e92c
zc7dfe3ba5538754263adc0a6295b7cb095906be5cce007bb2e5da06cf9b0ffcc4116828044dca9
z4f7a10dcca1aeabf7ede01e9c4070795913ed141fc9c87fcbfa58728baf43329aa550cdf5808ca
zd285283956c377e8a1071707b44cd4688489762ce277bdd2cb731d2e5c4e0cd87c344137d35bbf
zeafdd506d95bec69d08e333bcd435f5b60c06b36820ae1833487a87665092e023f98588c4ddebb
z8d571be1acd30177e16171d914be92c9d3fd84f8e30f977d206fee1a0118d9de3fe32a40daf4a5
z64e7ecc004dfe59a92685073cc7bc0c17a2cf62a3c47b60e0fa2a3461ff32fe1f4c452ff0965a5
zc7f406f86f90e074f73c4cc71cb2b84fcc0904c791a35bfcec028da626053466ec8107d6faec35
zbd8ab705f3ab387e18b9e2aae1970a27c0b80876f3857bd859d22beae6b69a4b18356fbc8b34d3
zbd7b43da506dc3c46e68aaecd75999f30e428420c65ed76d11c66e734e5e1cffb2e56102fb78a2
zd6527532d88f527e5f31cd41e53348000786032761e7d9234efa1def486f7075852bd6ef582afa
z72740c627b37fcac99198a0be37f5b616f9fa486bffbc78326d0664fb69d2fc9d8bd394888601b
z0d18908fded56feb9b5bd47ad929a824818476ddce70dddd1aa5a869c17436e11a66aa099bd4be
zee231d133a3c2d5e8ca98db016f620a772406d87e5d20366ebf207197dbf715f2725217314e6b8
ze15a23ba83de59c9402f78dec031bb4ff9fbd5306d174cd3ae8c5abe0e5e2d77ace267a4d62d83
z1a35e2c7e32e63f40d4d22c06792f48e79215c41501225a46128fef9dfd07ec99de2095a86f697
zdfdbec34c3872d3346703d0a5845a9867be93adf974fc099c3c06bcb2891aacbb7f722a01eb39c
zd5b35c9b43402625c22085ce1a17d6ab7cc084b3a6a3d3db17d62a74e52c0b9e3f8bfe2a2439c0
z4b4018aedefc2b954358657b45ffe9229b3e11270e8dd0fd16b87b02ecebab774229df97854667
z1c66e7bb561665434f533a240e927d8dda23e718df9dab6e6bdedab4479e6b7adf1da6acdd3139
zdfb217086fad0c2f81ec62b1bacc0da5bb8f79cc4ae0ae950996f6b34983062c6b60eafc9d1b8d
z9e756958280769ce318872e9da0ea0dd654874d2337479efb62b30951c1678a8c5063a49ef92b8
zeccfee3e86d75dcd599abe4c4b059b84668f0c5ea7d0579950125056a5d000a5797e8f0857a9cf
z6816d48587aab15069039c14d76f291e79bef33db44b65ec4d25f0d3f669ca2984f5b39a16fad0
z8ff68db8e7ea6b5db638b8885d1b3d85f4b614019038759c5f42bc8e6b2414893efd1172216e40
zd3a845294f6f597092cdcff9565d6eab28f415f5494c3247188da6d4b4484a2adb8d9023098738
ze93fa520ba5284894958c3336c1d27adfe0cab1959f01403ebebc35a31d90e673f8804ebda8943
zfc5b27c393bf5e7ab24748020d695a634aa778b953a6a247ab589ecb850cf1091611242e88bd33
z766daf83ed345a3d74566ac76d481579b72516f9abf505f9b2bd473d305b68e2bb21b15e755b7b
z884cb54f3404a6838897cc92a228e67f96a9dccf761e18b9a9520ede9e1acb19851c5beb4453a3
zcc5c872221cb3df26fd0e013c6702923a73df1d3c3c42ade934d753afe368aed959c91c22f7409
zb7401ca7156c14729c11a40de36fcf279016c3473c50d1da6b8ecb7dca024b415e345f97a90a32
zd1faf4b25950e016ba7b920aa1ddb0e7aa8d8c4b3cf191e2100a9ae264ba937a2edeb663ba9b43
z66469ca46d3233d4ec4248d0a9d85550522381ba8f11f56fcc4f2abf8a025a8b7f2d1ebfecb148
z731ecb7f0f750bf6f9da5fb1ec7ea6bece43f8eb2c094efe8276f0be3fe24b9b1683bf53ed8fe6
z8707623a6ef9ee98435cbb4e09aee480043b74a62e6afd415ac2031522a70a97d852cb1e4c0c76
z1aafb4b3610291e21f0d8f920905ba2fa276be0d809d79849edf2ded81afdf48a5026958319de4
z2ab347b43a94cb413d4798cad425bf599947242b5f674c41a4e53a27d768e9b4937e8e2d176d36
z6d23e4460d997cf0ea3e2cd39457b2757801e8481cd0a5853446aadc5b732ea8df1eef10c3a606
z82a577ef1cc1a336c5e0d912a3158ff0ca9166158285fd59d32446caeadd46da75cace73f39ca0
z10de1a9276b2cae96cc0cc5879b1c4f08fadefe207053c1bae4a642abf398c1bd74f5f800d8e33
z761f925657f1a27ed6b0c93dfeeba98040a730ac8d02c1da1cf66cebab00fb74826e2b64b90c9e
z9f669f7d4ddde905715a8dbabc73e2a16e174bfd047f1fdb5b0e5728a2001523178bba8d2d2782
zfd5d956ea67007de23e559e23b2c7b0a1ad311a44ace9c9c0f9a509e7939448814203a1669cf4f
z37904c37de6f0deb933f9fb09740be4e045794ede6d3d82eb4990a43e86ebc7a863a4d02e19893
zccdf676095887345b02da5cda019a95052e48c6edcbeba83113d361b3f48a8bd553e75fe0d19c5
z784a44e363844fd215ab91e031ae7a8f7ffd53a956ec204e2fd9bceb2543dbf7743ca40111d3c7
z2911aba448ee70359f37a3b6c70b06f54875c5f1e1f74e17b59c7ed256f6bd759780d05fc014cd
z823c16baaf5b0640052a1aab898498b5ec4873b0eeda7fab125df32aeaf44a296de2ba375aa984
z56d8eeab18d526d62a588490fb83717d1e77bfa6d6372284235874e81da63428381f5a073389cb
z12d8a048f070991c20ae325cbac7760c73c40af5b380bf033c990fcafc6729ac681527b40d9a84
z72e85c2478fa5752386a49ae76faff2b4ea3d06fcbb468c01712d1035248e07590e58d46db1702
z10ec1cd876660a3df4dc0d113089cb997f9dd961d6e3b5fdf05c3174d92dbd50db05d5aca45361
zbfea1fa2ce97d1e8d50cc745664edfd526d08ec406d7b1f490692f2384a91bf07c42e7812d334f
zc232db0f33493ef2ea2e52d2ce861d2b72f7157f6857d46bb3f8af346fc4f109bc2c51d0c26af8
zdb7f79ab2030c667ba80016ae2efc0f1efa3b599e3754c5889f50e83ea5530b2945f01606e69fa
zcdd501a61d4912a383bf2470e45098c11ac4f8901ff54b74b5fc955c4eaee0142579d24f92a34b
zf047eb1b1e49341f8b2150573923f57d187128902f93d04a10cdd035b9626c090da06d5d96f93c
z5dd265c431c3936d9380473cdf8f77922c227d947ae06b30b40dd1e2a1da35e06b4357a05b0972
z3b4d338d8af66a78f562009cbce2661cdcf24dbde1bbe8fd8907fd7c690e0b2efcfd1657deb7e6
z0cab5584b7c88571dd42053db3232508dabd25968bce8f3ac6fccf5e9b90d3616185a82238cc8b
z3741e578f83bf314392ac0ec9446954bfeea3a03394fe6d6c7d6050eea7cf8d616db176d7d5168
z1bf5d1a08885d6f474f61d673726c5517dd4a2cb96dec965e208a831ab3c763b2d5d7014f4e70c
zc16a3b0fe67f62a72294fe64910b441f66836b36fc8d3028c96ea7bdf0a4ed9a83a7424ea4f02b
z9ae63537059f66fab3447b7248cd9c9f8efe1af472db0810a2ba61fcbe9e378941d465d7436128
zbffddc535a5d237d3c8b2e8534b4ed20ef83c823e6a11988d8cc3b7665aff78fb9641ba7a3e418
za18b32b97ca9567703046201d84dc73c5c1f65ea4562fdd26e4b097e61ab941ce3831658494ad7
z64c90e7059fe45fbe5c1e844d0be843d51834da12770c6bcb89ea805fab0b3fdb3b6130f11f27a
z3128b84919d0ba67e2ab77c9f34bfdf02196720c61030c889389751a8dd75220ba8e020b2cb2ea
z8adb3827ab4e5e6f66831d78fc0679b5d6262abd3b548079ed2b4e1ab9d01824e306c78a4248df
z18da8da82b7b5cc8d5d6be0c5b86e464556ed29f1a399ba05f3a2d7aaff63956a9362e8e91a6fa
z7fbd1a68d5760ff147075e30f7e34a1636f8bb10466dcf931bade1d63abfc03e66e1a1ff5474b3
zc8d9b4f65ca9f1e89670ae51e36c5910a96abc1f1ffbdcf510b1ddaae72021dfe3c07f3fb58c42
zb26eed464a911714dfd6785ea73ff8ec4a93513bb4f145e7442892746cc554fd70f785e484fdbf
z9f2fcc84b5dd1b3cb4cec914944a091933a36feb6f1133e251bbcb21815490523feae6be98e53c
zf170ba94049ccf9a3c33a257ce5498f482ba5613fea3d70a02da5f57a6a9514f77ee61864da8fd
zc268b49df5fb8362ddf500c274378f634f8d20780d579109668aaf6f6b5a9de44be7ab7d347bb3
z62caad178c1a5db8ddb2d64dd076f699f19f62953c54726039001d5d493854fa1c96ae75587ef5
zbed5acf6d9fe2d4940caabaae6c71effac97af637d695bece2f15b29cfc2384e2a8e868d176e9c
z05cb28af03a0c0c679a394c73a4b9da44e3bf1ac3e21a198afdcedf260339955881ee9c49a45eb
z75fa3dfd05dd3e89720530e2888725e3df0d5c2e790db34fd0059486097bdac36f266c1c881d8d
z723e2953f5daefdb13cc21d6dc3231d78d3637d1a99ce58108165a1fe8506802542c59e96d9fe9
z8e3445d492b60b33110d5ae103bb68796ba6ed948dad0fb691fcc7f3dabacf9924eef760d35e54
zbe8904ffb4121b13acdeee521f69aae06bc2943f398e86c0e8ca6d187e6983d297a64ddd08639c
zf097919c2e4e53467d57dc7a6a8473facad040576cbcc352ad7588da0c07e9340baac2b1f20904
z1d00ab72472c60bd2cfcefe935e048e206869d6bc28f2de64f1cd05a69b694ce387885a848641c
z71fec6b289b9fc7c45988b142ce126b3b1833b4485e0c04ee8001ba333cad4e1d12d565a362920
z39ae29782dec6ab61c18993aa267b95e8a910919ed67976c0592e27d093b6726cd23a2cd28d38d
ze0a5e999084c66296882e5e7a407dd6421b5ff7c68b233914b406040b4028ec47234c12a5d279c
zb15686d01f9327baa5d54e885b498228eff19521fc8871ae13df1bcd63466bfe3214256150bd61
zd87570e57aad6fc4ce2ca6ebc3a30e7c41a02cbcb64af175dabbb469e562c1584aaf9bab584249
z80e6996298b709ffbcc3c4777fbcc219b90bdcc02623891bd1f59ef34bef253c2103745f38c36d
zef8db55ed4d31b958c3cffc641703e8f0182309ba7cefba0475e434b3e89ea4bd166cbf65b2fd3
z4299ce6b2d361757015ebd57adaba5b69989162a0452f3dfaeedbcc8ec371cc00d37276ac8fa56
z2a59ea321276206a01b847e1ea865a6da95f23c3b25f24c0db34767dd4a7edd0747304ca9dfbfd
zc32659b25b366fbb39d63901dd359772640fa6a43ebacf84cdb40364ed183f14fa518afbd2706d
z07b9b0c27425055a542a48533ef2b79b0fe35e43c7b6e5f019d74c755b11032270a373e4678e4b
z319253fb9de0b8dc7ff27d7351421cca12aaa45ef5d7cf3ba6c95ccf9a089f276ed16da951d58e
z0b2826e938ddfbd4eafd52a67ae3faa2b3aa27e7544aefc2d0b1939a752183d6ac1905b5487756
zea9f32c4d3bc30cc9edfa54dcf9a0ac54df61c0f65025eb876176b93d47a263795caad4a1c28d4
zcf4047eef721ef72a82c873944c2b27266b667cd5e02ba746bb8d73bfc4937630a6c65f715c352
z8a2cdd361afd3808eb1b912c53aad94d81d31fd74595e8b4a4c2e5e3bff938f35c23123c120ff2
zc9ec35c997616c62e245ee31a1435434cc0af375881b0c43fd90a51955b1637d7493381f1d2e2b
z5d152c3af37959ae9414589ae6ad0ca306fd7cb669323f1ea8c2ac3207cd2533cbebcef67d8dfd
z4b4a036b07af4f7bc8cee856cd9002855af8cf07b965a43cdad624d9013dc9ab010823a484694c
z24c2900c1c979451229a43802baaa6c3d2949e19d305498205399cf83b8a9771a8cd2a3d950d4d
z52c243bd1d6895e2954ad0f7332fce28c531323e37f613f08e01da234b9f82d264a538dda68d24
zfaa666c811124594958770af68900eb38a1f93770d3923a52411b44c82cffbf14544a91df82eff
z90d9b68f3984441d7afa47cff9247a4b679cb560d7c72cf12d5d21bed7343a450abc7cd4618d65
zebf3cd8aef7e64403a8ba9d6ab0b75ac385b0921b6830ae1625b01f7c5bff5f7e882a821d27117
z115a9b02c0cb0f0944092cd0f0d28e2d4eb62500c38d78ffe097f128e99ac810e9a6ed5b69bac3
zdfc0b4bc742ae777f3ae04018f3e965d8ec1b07dcd14c61ba06439a49f86dea085bb92cf8ab5de
z3681b349b3579abaa89af4d7dc7354733b9f0f63f55a47a0373361361c4cbfaf61d218f2137c31
zdd255749d45b9612782ebae0240ec430ae81afd0a5c5bc0e5fa2382c81bba55ec0372decea6f2c
z8734330cdb8b7dfba16e29179cb7d1ba92fb1eef799b36cbde746f6bb202db5b57c72a925864ce
z69dea2ba41e38c633179e851c554bb9c5aeafb65b00742c495bcef36f7e8ceb82bc4f603a50afa
z1821219cb5d0cdd38249f4d89630558ae41006983a993d8907e77642ccac932e9a9cb0b1476bb4
zb1b2a56a0bb0b683bc798df22211fc65594558c6654381abefada60e3a0c6ec82a0d64ac28456c
ze3f228b98217b4ef4cb0e8e5c14c8a4fee37cbfcf9d7201b1605c40d447dc24a8a534f76b6726e
ze4ba851f1dbd55e9f356a8119db0f2fb4f5c585a3bc4fd18afd071c7441bc0956065f9ef513835
z9380fbe74c618ce94cdb646e3ea1a37efc6105f65d76754f5ec479b8ef74f2db103ae0205899d4
z1669568e1fa344cc3b3b7eebaa53613bc35b4d6da7bbe20d5a04a73e72752b2b69643b78e4079d
zdeccaa690d3850d7c2c5898ef07331bde2fdb18644b79f42d0a4b5dd1394f4ae6bebbffb9a7362
zd75bf34534ee3e26e178d64629cf5feec4477234064fc35ee60d4f073d70973f3df8e592cbe442
zf88f9503623fe397fcfa2ce042bb08844d8f14f698271e5bf845bd4300adf435d50e8f84b544c4
za3a8ca9632151e2630c9c3b14a2a305bcc2a0a1c6ed304a6b2bfa4cf97891c942efa76f04a7014
z0a13dbd43143fdd46d846f3e39bd9b81516fc12693b1ac57be0c8000e7ef1b27445056732ffb9f
z9b6de0a8980e9eb1807928818c35f2d23990a15be74b19db8ff7ef42e6970272831f489a712dbc
z441f29ee5ebc871b9121af8976040dc9328d373700b032101cd53c0a3594d1367154bc44565630
z916be9a5977d002378dabf48e931e56be806742fb8c95a50006f73e23be3eb07d5ae6b9cb748cb
z6cb40d4ad0a3de1f063e9d6b6a2ccec303c2331b90cf1b63a946fe6fafc6547b8f79b1099eda0a
z5d9f14bb1985ac1ad0638c757d8cafb02a3441dad5f9a4013e91dfdef5f89926e68a4f22a1554b
zc93296737e6f97486009c8c6891c54bf7f000247ba548a6e6e1de340129f1077d33b6c1ad05b22
z660e9ac299cc04feab2607926255ce4c828ff091f833aacb1aaf224fb7e46225b4de7248de36f5
zd8aa87680bc16a440ea905b7f06b8c7913eac750eab4fb3fe33cbb0b1f974639ee43919d6c5c69
zea0cb552a0e30be98a7939770bb5d1ac2df3ad7663d9156147f2771c2a82a7fa7e0d7b31afa37d
z7298b08d78cba06624f9e7046e21549429054c68397b038e17d0ae6877cefb7c70031a57ad448b
z8c79dd7456b2f3b55aa0fefe4fdaa06cab258f2ef844b5f75b5424ef80ac2a76bc36b72e98841f
zec0a981c681110620331cdfdb2cecafbff8fa03b8eb2b5b6345ffd517cb954d21f657561155291
zddd3991ac3cb18f83734bec905e808a014a5a521f19cba240a900751658f13ae1cd1bfb166e550
z32594c75f6432bceb29c8be8c31ffa51fd1ea9ab0a9117b0020b2f06d4adc3f431033b4e1714c4
z1fb2f2ead80590dbef321db3c0b2eb816a3474e02d193b02ca5c96c2a60a25e546fd7496fef8f3
z2d10996dbe68b1001bc3c86707dc2546638ca39213869e9822351e1a2fcd258bf501133709066f
ze1de553523f7f007586969940bf6d57fee891db311153b2fd260df1a1a006d7e695aa884dd6597
ze3e65e33864b604f986006df326054536c27d1d5ba9739f42b39b134c09dd5a56d6c5bd866b716
za7d6d1fa92abbacbeebb1be38dae0d9a25c6e1437c68e2e9309ce9f5d6a0d78951ba8561191bd8
zc3993aff2951554133090d1f76f138ce8ce81fefe23883653ed1ac0c93c4482fe481aa6615730b
z1d99ee72c49060d82f851f39d640d4f5f6445a12d820e9e0edfc902dcad5e03f5f8f86fa2f176e
z699ebe8173219abbbfffa78d8a1a7cfa553d9023b9ad7450c5d3fa61a96ab6a92ead79b750facc
zabe4fc466eabe227260c0c475410910193b14487f274bbf09b58f1259f039cf82901c5feef57e1
z2f9c7a60b7345a90daef5f1d16712e84b2b386802450eba07d18b91b1e199317f43d2e8131d169
za88a71cd2ed6f549ca7c1350769af65075828777bbf518a19a8bca3d02741e04ff18405e4c168a
zbda557edf9f9485785f2bbe3bffd6b98486e46e5f579607f00bafda24b9374e3b8870072f0770d
zd4644952da98edd965a51f414143da96e2f7de0614a7fef00065aa6034c773b6448b41d163f5cd
zb36aef4cd181abd47014d58e3007404bf68252b16ecc660c9b6981762341873fe45e6f4cd67cf6
za18247cd69e25f83bfa99704c0b3fa8bb0fd71c2733558eaf1e086d2515db0f6bfb16069c81f1b
z0b5cd0225671df68618448195133076c366fd90d9e6a54428db7655641f6db56b56828f28919e8
zd8a41e154a93393acdc86f46f705b2eaf8507ef01c8a93c0d096beb5ef77020379b374418863eb
z85988fc713fc7bdbd5146b3a52740c87dda8a0996acc7038f2f8434a27ab97261f333353b1524f
z08542e211e24c07cd47fa3522a12a503eacf04831eb292f4ac7ca1545cb92ccd2d39feb93e65ed
z122872304b6aec989fa316197dfe6f7b8b11bbeba16b473ec3642f4b3d047f2f2ce69bebf708c4
z9e03bcfd5d8257cde26b98b626a292fe053b9b5fb2e2f8247e650a103ed36192443c7491ed5622
z3e8292b19ef2230b573a8533d63d63d34909e848b8241876a9ba079fed39cceca7ed4915736482
z4c542285a0e47bb1096eaaaf1f8ee91de50770915ab29eb7cafefbd543b5bba19402b5f8bbd963
z6ac08ff2706bb491d2f3a5b76ca9bfb5df5901bb6e69545b890984a3236be60012c73b19ef028b
za678cc7efef8988f8a316562cbd2d92ece6b0ac76393f844913f30b7001e863e986cc1152ea3fd
z2b28498de254fbb653e7ac680c4a86396cbf156b7e3152c1972d8a08b5977ade8a1da2c4ae2ee1
z41a222ba2601299ab446ca46bdb69f1ca6f5fc5a11a7464172ec8bfac4bfd28ef0e35cdf718974
zf49c7f3270d319043418767b183720229beed566e14abcc1b655fd82260165041d29140ad34681
z262644f4356270e33323fc85066827fc4e8dbc076987d15c4306f86e0cdec2e04fd483d022d1b2
z78a665ca2ec6ab743c7a0ce11af879e765fdc31eac2e241ed3a2f930c4c5fb5f48abfef4c776b2
z1f2a48702903283fca5d068e3160e4e494b3cd62489e08cff7a4aa40380efb97dd7c035d7559e8
zb5e60274a0c7aeaf6ccc542857241255f3c3e7bdeba25c90a9e7cc058fbca83350b4b41d0d09ed
zf38ce7d544c49b36c9fab1a877ea0f5395b77e1d8ad5c3c6cbf5d25ede47271f89c359defef491
z043c8dc85af39c3a64df769794d04acd36e96eecfed7494baf39989b09a87f87c90ecd343404c0
z8dce6d0066c24a470f3703e6aecc034485141ea14fbed0ab26c43e206368d9e874d5377f47c12d
zacb6b70b964265d26e3d5b78190429766f348d5e468b710f0ad3222abfa8dd36389475a927d500
z53d7d6727406b3bc3884ca3262d84cbb709e0b7da7028f921c37761ea6ecdd62111782a4e173b2
zedc5e65c632cb6b3191e69869ebb8f8a4d36650451043b113b8d31563c18a8af205e91a4458ed4
ze5fa2e221ec8cf390bf28a8c0d985d733277322b34342b9ff48b4b20a457bf6916724c1e13b19f
za070684a1a572251869deb88b57590f5349fc24f29f75b0ad864cb0bbadcfd122d773524337ffb
ze62ef2d06dab5ed36b73acba0968f49993939421247e21268ee457aaadb8c25f496be6ed438c9d
z533d5295bee177e69e3b4df12a7013800d92de3aa1ca39f9889f5ad9ff3f01b03934b0de091fdf
z20b6fa8c98236079ee030818e7630891c8d8e30b76ac0ae5839b29201398359704fc970c881be0
zc2ab033ec4df90bb0415c7b0b1b19fc47df97f69e99a054bed9b7c89fce144dc74c6957a32435d
zd64db2bc2a8f4c67a3e2df9d8de674601c74837c025c3a4e51dedb46ab937899ad404b49efa58c
z0f53b2f6e41dee280ec60c3b97a275ea7afdcdcf01c669511ba01d64312b4872ed041e06f2df6a
zee9b0fb9aedb10e333618d7049d90d61b1efab3a004fcc9bb0f92a2dd1c2f9324ad0f1ed1fea19
z21503a53f39548005940b66440e59fe5b78108ff94a6a3ab7b91573be5a93ebb67be563244f583
z5bb15cb439df6f267e840ae14bde4fc77e61bd1656b13a2da1669051663785037a94a66c9a5e3f
z9a7c71a76d6392c7628352f187052a0d47476e5eed95fa3162091d4060031205d4c7a23af709f6
z91c5fc1f534c855864711cfcbd55d89cf88a34491e0adb46ad039215d8efed863e6c596db75866
z89a57957f2173ed34c5a34bd3e42b8d939e86d1bf1e43d4eac9b7a5c7486aa69a1281e79a21a96
z1cd74e868754df6f3a7ebc7f1e06b68fbe8161297cd003e6c35dda1188a8772cb2488564207b13
z59d316f74133afe742eb0a383fc8acfde99b382fcb40d6ac01523a9b7e940750011bd90d038881
ze51ff411738e8675dc25b44b6fbf7236af76780f50d7e7679b451d73d2f371f2565bf616b57061
zcdf37d4541b4fc4edfd4a4b29791b36d0da6e181f223660197da5b5760fba7a86947a5c39c71b6
za1789353727214eeb3f084d32a6644809a04041459b4ba4ea08fe1c59d40cd38c43fa1e997b50a
zeb2a0f2c1ad3b1f13d568df2eabd8b37b79a0a6215bed70d0702e59876df02ec975313ba09b6dd
z2c3c3f40351219700bb5d80a64261ad60276692c309ab0fea0c71713efd0213343df7db5a839e5
z21e9ab3807709600672ada8c6c5e6237fdc53110e175d700355e325cd6cdb6643bc43bf3b6bdf8
z00d72a21890b8728509bc163ea15feebf144fb11a70d66aa91dc72b6631a4e059d5219fe7fcfcf
zb26d99491ade9041113be043ecbe79976b80f1974d2550fed7fdd4cda7627206d1eca398d7c610
z5928168cadb93e0d37c4f862052c7ae304ac55d830770c69fe03de9c681560c06a5e4dba302c7c
zad7783c846a9b9fc9094a33bb1f1c1de4ce1fab25905a4e991de0035963b316089a0d595f74ed6
z2e5075777097de75cf0579b09a123e7585b6b686041192857444a6406b888642346ba295c713d0
z47f0e3f270612c1fa02cc90f393c0835af85ee97d278ebff7827be2e2501f659e4d6cfe16af75c
z8003726ca134470268342005b666a7c8af0358db3d24a85aaede3ae34c015522d19d1604f674bb
zea8fcdc13842a8ed7384f833e11db0a8e85aba6a5dde62df75074866d56291903872be5c85cf6d
z58d3a98b0e965869d0b3ad357d33096af891065e4ce073a7c733df60c95e31f069fd4a4ef6051d
z06c0daeb84a9d99bae7d33b345a55aa09e311309c8c83d1cf8e6d5962fb4ec584a4dedc9dd233f
z58e30eef0feb571b8331345a300068affa95576cb064585fffd5bd71e1744b0bb168a4f371a4f0
z78c2510e1064d16f66143d1b0e2efd69c9294d65e41690c8b7b5646bda342f4c3bed80d90d999c
za2e7cbde4f9769d04be6ac255b56067e342c11818311e2a05c5504b92d8e0aa54bc5ca934b7d4f
z094c2e6c99bf60c14c4854e88ebd9fb98e8efda5e084169688b1797438ac649524cfba694888d6
z1630f0c8dbdce12e73795ae84539ca47c9250be1026d6ac5dc12a3f012bf6deb27489aaf8a4e9f
z3cfadeb7177290501eeaa0806113aee35e76c0d1f8317e8af0cf1bad752a06a52780b38b34271f
z29b686223e8d6be69be5f5b24ef70b3a1095e30deff8a439148598db45e8197b9ff6f8f2fd9948
za129ce0a7898aeb7d3fe7735fd62ded1f36168042898fc6d4b04589c82014122d940e9a6855e0c
zad872657b159fb8973e0eca2efbf77b693138743c924547ab37754ddbb4b5ca64b751fe9cdd96c
z27276be214ae49080101a4bcabf597f99ec974e1e872632d1f7c25fd0f8bb001977a9f0a61c3e8
zd48789ad6aae8760aeeac826075a5f7d607bc3878254ed7af8b9aac7fdc07eeb107a34522a2dbe
z6a693838894ad2beebed46e0de6362a4f18fde240793da005a24330446c38c5e5738333ef2cb96
z46d6bc4ba8163da92867fbf40704d0648bb0330ff29d007e3330429c3d2f8901315b451e6af2d7
z372b260d3bea1d1f4d3994331faff7a678bad0bafa4334e9911302aafbc6962e016cd4b6504f77
zc62cf51ec1d495cee351eaf9783961c352cdf7d2acb5fd8f238aaa7c64fabbc8467e17d292cd9c
z4b7237d3b901059e4b6b59da99209346ac0448e559631f0209db66c9cd75d025a01821921ac7ca
z723230c73c90162d520340737c0df67daa424bdcfcab9868b0314f9ab520ee0bdee09bfa96b10a
za49f2b23e8b3935dd6032c4b15a8f3331bb5516e968fbf42e4586ec99cbba969e3661f5f8f2ab8
z679881883bb5aa720c7e824c5fc747a5f3f00ff0f45b3a52e896b6d49e4676e8d0ca9ac6c902f5
z52a67df3fced26554443ecb04de2932e247c5cc18633073154bc1d58c2d1957241fd22d64b4fdf
z45dc0911e7effa34f170bceb74bb857f236c99fd395270e1a0e33979ed4694373ac5901df10032
z89f5419d65df8a587e4f83c65780ebcb09ce679ffff14bf4310b676c7a7dae3481d0d4482e105a
z7a208cd569ab58ad409cb30729dfee7fb0fd124662230e1abd50f152696681131c63ec4536ab2a
z9bcd8a4014c1a326be801770334a089070ea79c219d8a572446bb476ec127a78e488faf7a97131
z6168c891474b3c87531e32162b6774b67b4c873cb4f3a2b22960ddca720ed096d2a5766f3a929f
zf8bb749e2fb1ebd692912ac7028e0fdcbe3600a3fef8a2ef0435309f84b5b4f0f7d658d7f0879c
zcd5d1e22f9c01c42f7076a264a04c03b8279a9e2c75e486cd5886c2c19ff1a6c964414a2ef8963
z99d71f57f8238854b90a5712adc61786736d0fe754d79665176be708ffbf16f78a876632463c3c
zcb11f53d918bea456f41df78c627f81e5a2472ef5fa343e537b04c263b8750b5f237ea7da24ef8
z5dd128b30fad963ae4ab62e4812072baf80ea074c0a9811a9ebe7acc1a752d3dc236a8c3375b28
z63464bf1be34a04892277c4c104af5de6770890c85856f857fabbf42ac2202ec50950bf0897905
zaca5f8cd307f4885c97f9460e91f4382e8328d9c0f96000d602d91218dd034dc2831bb4386f13f
z44ffc267cd1a0daaa69648a09e7fd9ebf0f4e5d39df9be5f2c4d2efe3a947a5ef4bed69b6c2e13
z09f1de6818db12655b6b6a2768a78c34090df81e627deedc6067f604ea1c2a40e0639e3a863ba2
z82aa12093cb15031776d952fff564a8e02b10a4ea07818659c7e502927a0ae8c9a23c578eccfb5
z4855e8c9ddc9875f4b25a170563456f367344047912952ec43215baf87ecd5446aa8876e3c2b4b
zf86e05df11ecdecbcabc9f792af3bd820af119a622dd66d968f5bad4e5dbe66045896f1cd69d6a
z910b5ce3aaea02ded58e1e8e31890a0504d361962c2c4fcd6a8566b4a6aad8fad9d6f0b2b47393
z347755b1987941ed58d06e9f6632968318350b9f854d5aa1c5a50230df5506bb68a93f0d60361a
zb1df3710de8dfbcc026e7f7da806ab183428e485d343e2fe2489bf71f067c3f96d3e97a40afa57
zea5088c85c451257246c3cc693a308bd12faa65c1f54afc362706cbf5785be609122246c2dc564
z3dfe1a42cd4df17d7ee5380613b02e9737f9f2d619ff7df329fe1bb601934a7aaa425f40b30406
z1f21d946ac782aecc8420ff7dd6c7af42a352c40669289ef28916f1718bd179333d17e8fe0c158
z36592867aea781547f0596287cdad8fbbdc08ddf09c3d44b3142e068d832938fbf6efa39d0898d
z4f88616701821299268fe0e44afd90d263a7a85d826619e17ffa86d40c580acfb26c5b9fb368f8
zc7a8af602e0396f59312a6e8df7fda5b5faadf7d1d678b9d7e744bdbf84faf6651a1a6621b4a24
z3e814835c4e6183d9e3c32f971af922cf4863fc2b4d440988210bc461b7154facff25ac96ab924
z4ddbda8df447e2482ca7396f6934b8c9702778d329e1cf6f676b195498b1fa57d23ec1c0bd1ace
z5b10fec34a77806335a7dc2255a3e76fdc345c6045d5b8a7a4e0a350ba2bcd67cb2cefd6806709
z8bb6ef2ca87789c94d544de632003572d953705cc0d96feb9d909c3c5cfffbd03523c49beeac76
ze8370e84a564de9c160e59d30dadd418e66f76eef627883ff43d59228f13d11dc2afaeb8f7b339
z78e663f67e6f42518be952066fd706ddbdf6a1f846e70d12b3d817330240e70cfdc39afe7fea89
z442f5be717ecf6fceba6dcd8ac769c559728bc6e0805924dcc0cfef3a16c92a25c95888fc16abe
z197783f337d02f0cf6ce9d8b169b7e7c3196ae0dc2dc094cb21e8b6e28609210f17809b798b734
z73b5dc5dadc91cff0cce438d752a9982b7eb61a776f4d4d25fab8e88fc5346c59ec9c2247bc8b6
zbda6d9f70c0ea295ef4330f12d2a88acf90b1013923e585f6f8e3f2a65f734c069766db799fe4f
z6e63d3aafd53edd28127d5eeacf7fe250c4fb988540bf8892cba88ab7ec3f68dbdf2c7341f3b2c
zbc819ba85ddf01217b91b38b64a5ff64563944efc44c3d7353134b303922e9d55bfee6fc455750
za29ea5f897586f30a6115c9c0448ed27e1e70bc829e2132107a65bb89a58ecdd4d48325d04d864
zf4a0a739ad68b1b08b387afdda142f2a9e46f0fdcb373a7311478402122d69c6cfb1ecef08f573
z3c76317182c43cb63d6745ae360c3cd137239caf8dfd64ff9855a9dfbdf523027585b1a1f87ca6
z96080ef0503a7da2bb62d1a2366e8071b5124bdf09b0e57cd5f8f03bd93b3deb50dbcf61a12358
zaa74ea0a3e5170c866ce03c09e262eccdd9444523bef63cc7e2b62dd97ea8486cec847d7424194
z1e3d8d620c78b27eda27ab10ca202f6a1af29d04df83c2a6a0382b89c8a11247d99435b8ca2025
zfad5af49c5e9cce2589ed189afc034c5fc79db06a9a83f92c5c997312ce4cf79ac9cb2128edb32
zac97e4288ab4b28303f114895b2e91c220b84c5e912f7a70672dd07977da14ef949d36fb5de278
z339c65e798299341092b8b171a2b35480c2a787537133b7c18a9ea2e958b5cb459c8f39dd76aa5
z5ff1bb9de7336662556a82445ba78e7b243bff002df12f1c7f46b8d50bfb3f927d97a2a929fdba
z2a4aca2d6dbd9ed2017e0fada0c19092a33f38c2183f7ae5c9f12c46764d62147cbafa65dbe3c1
z98a675a1e5a991e35d16ae4ead4668fd9ef150faf47e76341da7f1fb3ef9a37e6ef490abd4bc31
z7b1babab8e28eeb567d0680e0891e48fad006a77292dc5f5d0db49147d7d4a9124e5d0c9435e15
za77b8022538dc85e347ddc8839650194a2fb79d7b207df83cf92e9c39a146edd2cfbafb3198c3e
z60e3680f30d7593bc8bec17057512e602bf928814c080859cfacf3be648bf402bc8ca70ebd4041
z32886a08b404802d759ea5cfeabce328a81fb8b86bc96c2f3d34a79b8ed126222188842411cace
z3c553431a3de7f6096ccdcab055fe2ebca927bda78ed30c690cb72729e8c27ea89bb99c0abc2fc
z0f7c09b4b8f6cc0a6180e424c4c0773449be5f688c979c3265051b99903b921b75052ce108716b
z5cb7222b894797b8204084b1a2a99bc9b297ff0acb36fab058c342e51821b66c56ed1b0f59e4e9
z0718f278af9b35f4d1f81a9d922e37d780fe6930b51451c0c5f4dd4de1ce0964feb58bbec4edd4
z8a5c90377e0a300ec8dcce158e2f67d43ab70e5337b21081ef4ecea634f05fdb0f4c04a516df6c
z1de598dfa63f5eff15f54d53dcf1513d32ef8423f0fedb281063bb77f0d92d03275e23cad13c37
zd3c6d7f47a95cbc4a4343ba7b888f32359362e8738ae759c0807f04c7c1268167c08e36921f13f
z4e39f503cf202148881eb77f6eeeb027855ac33631e03094a3460416e76da4a52ed13e0020f04b
z66bbecf9ad622c9dc16cb63a28796262f6c7fb78ea4a18196e321d1b598413904396a060dc29eb
za367f2fa0abcd2c6bf197c9f1bb0f6587bf02f5e246fb009922f86ba98d2ba39ad3260606d820e
za48da932482c95b001b303d0d239a5a12d72a4dcbdeb6e5db83a125b6f62589a4fd7c62919cc90
z2c6437d4d5f70c572eea54301c46f623d6fef3b3c43c646c0609f5400d610bd06decc95aca4d0c
z65455f0700f43506f6e090c91a2a507acb84d7ddf761f5ae08b07ef59e1de864e6e5d3711614d2
z5dc4df65c04e5869b36772f3bb45193402fced4e8018ada19f59a5a580c6f079f0da108dda5be6
z1b76a0f5fc665d806bd80d3a6a3662949399bcf9518f9784d3eac9aec2b39c0428c6dcf494ef9f
zf0fb54693da4a9a47f6fe041ae3412f5400ee935c84a10e30dd06eb6c6870e2f2bc34933119cad
zb68c8cd3bdf6d1943ce708725ace6446439c7e95a7fa20fecc3507c6a7a06ba3f628d2940f5e6a
zc8255e5797ea2ca07513b43754ee938b9d2f8137324576e3eb8e46859b6f6ff4a0568d56401815
zb9e309feb9ba913b847387eb956e1f9c6584d76338e47eb624db84b710a494721d8956b0732613
z77d535cfca1939d7898610358f119e1470a0b28fc1c1b70debb34e86973eed5e066c76ec5842d0
z6203b18bfd1e6bf009891dad88e78d8827312fad2e623d261acb3f2184cfa7a72c757eb612c690
zfbdc8b50246b6a8c7cf0bd92ad6215d9f4b6940f3a82d30b64e1b5dd819a0478dbc582592cf3b3
zabbd146c6bb17be9b1b8d43d7ae6a89e9559300050ad420577c922c776e0fc6af4ccfa0db47e21
zf516d291d709febb1957c67b62afe73df6c98c8b89812be4b0afb4d2e20190ed1094ef709f9dc5
z46ed1fbbf1676d23dda6d07cc8a10f0c5042ebe51ed6129f74d0a0194c2567573525519e19a88f
z58e605602cdd976717e9206713368c920a29849ccef63befd2bb444fedd55068b7824aff077258
z23c050aa796226674dbcda703980244540d9c7b33dc95beecf3c3527efca1d14478da4fb53aa55
z8dc8cfe381d53da4e39add38149e1ef09c8fe943fc3a004c553f9187f5c01f1ea9f61e2d973171
z8bc86415c6c763ba104a44aa5e47c8e8fb6a4084e2a499e0cad67f6a6c4004c2266ef1613b4ec0
z07bfc03237a9681f46f7bd0b57f9b92b1d19f5ab2663e00e65eeb0f018607c6a1cfca8678db3e2
z31c1ab02358799255e28cd51a563ea59d2159dc3586bc68b61802ee61e3e56a457e30a945c859e
z46f5efbefb63bd28b570bd1f28e888d33b7c606e82c5daadbfe96003fb786a68c6ed8cfe0004bc
z2d4caf8c5a2218dba54c3658d1c45d1d492c10eb44d0c3565ec846260fe00fd32318bb3d152e9c
z1beb117ec3e4f451ff3724d05db0a0bca28951b61eb2fcdac6b09c4e3170506464546faa259bd4
zc881f0951bd7cf3229797d7d799a7f3cf73f21f9a546022b62560d8b0e7ab16ee4da0110813c3d
ze704b72173592d78b306f3cf75efdb0940a18b41411e00f0ef3f3447b1294b3bd0551356611da6
zff359f55feda27384cdabd37ab2b7294cce2c4bdda155e235cb5ded58bcb5d54dc7a152aadbaa3
z5f04d06485f4ea46c755b9dcc436851382c22df7ff8c2574ed6638e1f5655021b20ac97b9822ab
ze9ac480847bf42c89de7f49067a88c81d89f016fb3c5bfbe900539a51d3f6a1bc33b6e4ab7665f
z3c71323e4612002686a8b281e9129e4b97b397cdc81e6469a83169971377a2fe56b1a41674c2bf
ze695f0d94fa676919ad9cffc69773394bf797ec6c05d26fd8cdf34e5273b0e76d1fa2b1adc8946
z4ed3d5836d358f3a039f40d8b52e795547b8cfa01bb243799311f256319e920a6fa777b1ec8b11
z3a8129b84fcf59c5c033ab0a48f10ce2b36d4fe012410532ddc738c85af30f55d3745719efda71
ze2681492555a9847fa89eec96f2f6502b2facf8c213e2e2af42918034105149f8449891ada5541
z3ee50fb06cd89ca651b345ac8bfbe82e5067199791a10afa1a0f05ecd8b656a54ceea72933cb09
zed4682bc6e26c2d88ed7faee09d7398e750b3754e1e09a46e25d5bc5f06a8bc3d8a3f77b4a11c5
z4785b8b0c0a922483ec1a4b1ebb68e0d4a3b59845f37cda480346b0fa350804185c0d4cab59d35
z85222c9ecb460f0d23da3d6d4e5acf42fbb49c37f326da848425f9a80ac138fbdb0e5df69e09bd
zab2ba1a8e630d6a24967a5daaa8a2f503c6e71c0eb5ca5785ff7535db4b2262ec42f2fa82bb2fa
z193c7500744cd3a47443acb11c5e1a91c45d366828f0258c07079c6a1dd6b4d3895bd6ffd90b8c
z6496fa769c3898823732e7fac450a39b949b8473aba203596a5738ec1f5c1fc9c5571dcd4df0fa
ze732604719095509acb0f1c59f2af40af56bc5c1148b68093fd3e18a448bb9986f72a5bcf57032
z6ea49c704ab007bbb21645e283b660658e3db5393166c4f08a401425707453bd8b6ccc89994e20
z06f93ebba0ce6027ab2dbca087a35ff5503db6f00d6878ce8175170c6031044992f4e8144fc65b
za9cf6338fb6ea8cd070e9fb3611af5e864480dad714d13b465f3eda452f6cfcbd5d1d2e1a98cd4
z440462da1595cd45d0c3fd08a740ef63cd73ce7fd6d0895d7288860627faae74c9c7ecc1830332
z02407ed36b902fdf963b55878505c2fd90edbc2e3602116d5c7cd534abb74f5ef10dbc2104a836
zee6ca904eadd6d761cf50ea1bb1e5dc6f840ae593665144c7f005870e9b7041bcc8f29bfb204df
z16a04098bb062f16fbd26663ca22a6efac077a0465d368acb58d77f434ccf271e65b1c8d8f8209
zfe707c349940e09436af9390cc78da1daa8e6555f20d125e6c0ea323f5d56021d3721386e7e5c9
za39dcd257de19ac89d245390fb192595c31e300474869688cd813d6feac40a5ae1e6ed3e79a1df
z4e77e4596977167dc0586f58968e46e4522312a7c3ec58a12abc9e95fdcfeeb5837fd492c9c4a3
zddd7ca670248fcbd9ea83496cbaed7cd54e6998a3a0c054bacd546c32027e99af7b2c9b6fce629
zed199c6fa60724b847678d77ec38acf7ed3e2cdb2ca73cd52d57dcf583df360799eccfe654dc77
z504ce83002299c7026079cb28a855a93f437e04f834960751ba3a535fbdc18993cd5bd8acfc600
zdc8bb185f157d96d12b4f75b5296aa94c880fa59ef983295aaddbc99cadb2bb8aa1ce11ef9d467
z7cf80f2318e21d4589d35de3e6ec959342ebcc1636db7d3203f77d3dd6788928b7bf2d18af4529
z97b858ec1c205250736c157d523a0b74960ba836ddb04d1431e024e856a67ca4465167bc58a8eb
z0b254444697f14123745e60dc2937f137ceddc81638ab3933f87456583b0f198a95b543e9f4b73
za343052ea86ea6210d333b0fa938bfcec636e4a4292ee1cc76e9bf6edf68063760d461864c95ab
z6a73003f35a2eb74c9155c18609cc19be19fc42aac4615851d070d2bf22fa594826a7e28b77847
z00e04398f9aa0b5906e2a8c76abfacbeb334900c31522c1f43b635359fa544777e639e0532eacc
za947317767d90cb2611b46d4cb90691dae544e280716b5afdc953e2d51dce0fcf617660f0acb12
z6e5b1cf12a66e90e360f3cf55cbf9a0b1d67edf9b5ad894e8df832b73e547782a88340e1abe914
z55a42026b89802ca1ebd7d6a0668388e3d9c41f8083c843a6219e1937dc6f450c79e02ab9c3cce
zf41f3e8942c31564a8b29754beb44bd26a62df52af625710c09b89440ea0809f1eba0c6ebfad1e
z4b55d69f46b72028cbce47d78ec71d24a7e75b5fbe33e8eb9b761589afa2e8599353ec4b44d648
z9ff7cd2fc2f876ce360b522e75891da8d7f5d2e07a19622e47c9db546be9dd6da19c8fcb48c824
z4cb58ac8512bee2bc224ae12467f51eeb4462daa0b740f2e68df2d039ad98a0c35b1149ee6ace7
zb904a8692dd9b0003d800f011506cc4db9c502cae11d391d538f7e53ded567a73433b8ac3be60a
zb394c89187550d6dea0b83312641ab5ded1ecb8594989a7f20753243d39c8a31f4563f159486df
z5f892f605dd3490aca79e2d2e6af3f148c53d556e1be9c3076e958ea29939b1303dd509e860b32
z0a923e8758db376c54d9ad81f2161adb78d4b2bcc39c87b260c24780b075972429856fdb631bc0
zebb5bc5745399a1e390e4778ae8d9601314be7f5aa5c8442c52e3f5d049339109b7be613f6f830
zc3be645d09248b2cc6deadc42f6f16941cb6a51a0a18a0d3b85643f95212265d1bf61306507585
z86be64f80d42f7b054df06c4ff6f913c808fc0034829bd36555528707a4998946e95f55fd4228b
z14e0cb0463500eda7a85f3df3c8b86a2722369986080a7de2d9913136412fa2569f09b34ebd3de
zbd6517500d2f15f7a018ef5fa1451d978a685d118a89cf5e3652a999133b12ec7f75a1626b84a1
z83cc9e85d651c519592bc50ac7b67b898716e89dac0ca277da3e722124bfe93f53a7f123b89722
zb29bb059abf2f73cdd015b213aa80ab76bb58774cdff82f0aac2c348351171d89762f591e6bd3d
zb1f0f0808b344090def3efa39a3b767841d54ffad1d67a14aaafee7564fcaccc0820bf7ec2c374
ze510b7874dae3ec41a87363ea9bcedac744d538dab5fe37ca3e71fdf39a5379b1812aa49fbf437
ze3eca052ea29f965eb78b49829412f1e2627bda4d55460001a35bf48319beb5d48c66e64c84e59
z090e4b31cb1d7147ade88ccc4b56f74ab8212654a6689910c49dffd13e11e982927c9bbbc94d31
z99fa83c396550f6e60d2dc1df75bfba0e0f26a285ae17b27b8bc74b447faa90907d49c4aee539b
z7a64039bc79fda6c473c338a2a7e1834b0d8355d8996d916157774ec4e6c8e98c7d8062adac544
zbbfd18a6c93f9e757d5d48f01fe726a067cb0d199717a246d58c904fa534f0f0ca1c00a4541a6e
z8d76056fe950fe2cc505d3292094788a0efeef721bb76ad2acf923b89dcb050457865741cc30b0
zda65166f52e34cd9662b0b78d35660ab60886ecbe87d139c57c9a2ede11a515d93f1bcc2bc2cbe
z4ed1c10011539443c2e73b22b8f1f201f043d0e3f15cbd518242b6e8d226e136f611e2a07a9ac6
zc1a17b5da3f0d5761cf742b2e49621d8e8a066d4a7091ad278938c1fa645a804f60fd4973d14bd
ze59e648e8efca5e13e84f7c2199e08c33eac428fa78dbab834374e2911da085bc1f3481ebedcf8
z9df872f0b1975880a0539efc8d464894422b8cb799b4b33d3001fb4d957c617ec0c4871b8e2674
zd1501cfbc9d15b18efee8386adbc329db31dd5818af1d7105ce3007c433d1f0edd850cd285be3e
z0e11600b3f8b0b0799cde991a94897a5af71517ee2061e86de43f1ef8296adf001c6d19515d9d4
z8da1d86fec7527672c7e9cf834a6f18ade0616dd168e20c53fdac861fb59bca87df89f4be385ef
z19cb13740a7e356f31936451d8c5f3cb3dab8b79250948a50404697ac8caa9a07335fe7a2e3eb0
zf1282fd6a8f7a159cc68b7d66a30bb8d33d7c0abf0a61f0aeb6504ce03a5430d740fe6c44409e1
ze1645b4650b1f6aaa3f439170f042fe13296215490d2fca9b8366e392b3e7e8bf01bcd8275f88f
za26147f2f9c98326c0a8c70b14a11b474d1c15b8b0b326daf5f235bf8dc809af2fac768c963c0f
z22334ca1803ad601d8fc75dba84d76a42b096b057f4e13d647af89c585cf4c0c44bcb7ff5da96e
z9e31a913a0f1f1a2e5e7fde21c741a19d90fd99cbcfeaebcb51ee2171a1e547eefe5feae8bd4e8
z0183ffdb7b833339c237a9708f1d3d9842bd98dc9abcaf3e52cf040c077024823a20857fa31f32
ze18b4d89ba66c3762a51e62793814aab5d6cbeaa6e0756b336b30b0bfab98210a3c026fd13112f
z52fa54bdeefe78b3d633f2ad6847c4bb0206811d752bf7907c1b1a1044170ec6fac77c7fdb5d2c
z8ff301a018c9e9fb9a222153c48e81d70becaa93eeb5671a13c9c303623db52beaede4e78b66b8
z9380ba7c930bd36058df2193e928cc5d65f353171b2bdd50c05b0ff471971793c310b51718f05d
z8611a34260a1254305eed2e5bbfffa828a1f447bb18b94c76d9c857985041dbb7863c5cc8373d4
z876adc60be9e2d218f0e693f89fae7e631f3f34bd73e1ad9d5065ce4a120f1cf06861250ca74fc
z4ebe22186389609064a4712f3105182cdb4e4803f1492e196aea4112a94cf90157012d1c3845ab
zd64f77948130df447e109c8b9a9f54743f4d5389827feec4d10cf3cc9f84b74a142b7294d0eb5b
za5ea2fbbee003fe0bc9ade1e322eed157e79db249bc9e24ce5bd5fd0430e5ff7acc0f17256e1ed
zc04858dc0383c32422d0de6891e0af40064e7eb064260ddf4e21b3247633ac4153de1a3e8fe7c5
zbe62a8d191d4cab5f37ee9a8a157bf2783a76cfb2ee7dbda59d5d94178852dbdc4f5ad74275131
z3923d6c42e1d772441888f4e387ed975cbfb4f233b229f17f3a5b0922b5182064534de6a3d91b7
z171b39a66312c3dbe2998eff62bc52e7bcf9594dc8cca9cfe1b5863cedb460070d27ccb4026342
zdfc73f1575f1fc9efc4904ed505acecb8724c2b4d746d115d5b7d474ca4a89ebfe017d42bf3192
z3613fc2ac541abb7bf61422f47d1f8c68869c72fc21919e5c0dad36c41fbee2e4c2ff8f52d66e0
z2c478712ecacab6cb56568667e360c0f2cc5c512660267459c44d5f2ce3d97b4f1c3664ef26cbb
z30c8ec8425df250acb90a705cd6e523a0f5cf2dbe7e8fe4ee98526ae7ddd51a5e730919144e533
z25f392464da36a4eb11be33194917a7777ba892303b9029c8dd1c96dd97acba5d1f33333432fdf
zddce121b82147520f5b0930e27bf7d81868bc42bff8d9476ae89e70411f428193437aba6d2283f
z5442725d8bb70fe7d2a456b72a3da375035d2de718c1d3cac7d303a5795111ab8dc6d62cf8424c
z5fbbe896ad7d0c0fe3bb0d616f2d163cecf0b32d1aa3f3ca22ab90047f0f7d6928258128d92074
z1ed7fd44da13d2d6e41ccd76d0930c4ef998652773ff62236638ebee15b8b1c913d1da4b36ed82
z9a134fbf2e14b6784af32ca88e835e7b424b7e42c7a3167e92fb2cec6a1276fd5307de27ff76e7
z89a94310c0c03ca676fad5445d8367c4e18b1966430c92524b771927dbc698d0ff0dab31d014a2
zc73f289c6b7c1c3420c3eb0d8b8c8450bab37e1f5d32aa6d988e426e73cbd8c53b0a4871dc5ec7
z783abccb5e93831d52248ce0c66976071f0f9567b8ff5feaa072738f5bcbdf365ddaec71c42941
zfac8de081439dfe07c05e63cd0d12638540a17cc8bfb3d5711093653609aa5a851b9492ae5deac
z41c669eafca67a53e09c7b7d3e9b75f3cdc316943f403d57c62f6bc6ccd3b3c40ae336cc9d8e59
ze7237aa8d6529b9a0cc72178f6954ad7e7a17081d0c01d7cf2ccc1311b9c953bbf19bc4614192f
za8c252b69cd7e7e69ff2b433b3603f0b1a5764dff71485ab25a0d28a558edc150a0d26f92e7e6f
z2dd57771ebb92d26b2f3bcdf451c8a14b211a76171fca161cf3e6819d71178403d81fbda702e29
zfccb2354f9ec832c46779c2ca19f63ca848de08b720eb64e688abcfbebca30c832d21419b2005c
z0840ef478f5c53ff49653dd6fe6596bab4fadbc72f9691d925f2299fc348d4e3b0c5301af4357f
z97dae33f29c57e6873741f9d4325936a57b9ee4d33eca71628d1c537afbeb14f141a81ef0cefdb
z65cf3720b6e533b01131656785adb8822a994cfcf08172a61be60ddce86a6f3532108fb562d6fa
z67a300c41e818a62ce4dc795b6d57c914afb022e2a68bbfecea1b5f637f3ad065b0683f0af2617
z80dd2c9a435110a07af1868d627f62dcdee512fafa7cdac8d3b318f67b66b19575dd1d7656cb43
z0cb8d52cccb11d233b6c21f7fcd90ade7ff0669d3112add8aa10d6c20b618db779a5c6d648ff43
zb2db9519924fe0fe02522d7148d1c00a97b6c31af88def71b80b2a35f89a854a9fb237f9cfd168
z114c2cef76a6f155966aa3f832bf5894aa18926e4b1980ececd9431cbe42cd32b7c1fdd300158a
zbd0afa688793cd99878e2572075e2245a5af0d033b6c2582e82fcfbd5ec4cd3e5addd735760e02
zf9c0b39352d0cef7774f71ed33740221d17b15dd90cd93a9572aa87359274f294067e94c25336e
z5b52f00fa85d19a0ea18a49d8da229159eabc2c8278693a11bb086ffbaf3b14cebf407a5c84437
z1cd046858e49e1aa1e408af511d32d574407df786746530222c51d69a83fc04d074299a85d660b
z13e7d8da158118119b3513d965a1d294e321a30b2947fe1e34a1d2b3dbaa62c8e15352dcc910c1
zd37686f22aed6697dfedbd3eafdbb6fd478677a308055cb4a86c9195fe40d5107784aae8e99bd2
zd75148c881efb44d0b1aa1ee48a3f2e2211152647f27e85b10c809bb30cf89f4834e73ca5814bb
z72de0602a73f0bc8cc8935c5ee0adafdc1436ce166db2349bee211b5e2babb63817892241d86c6
z31dc3d7b88750c5b033286d9d16dd08940ec6468646aadf93dc1fbc10f964d4b3807cb861aca83
z70190594e59b0dc89948ae0663fa2641bef53fff5425acb2bf6d7b0e23b66f3d3e1f1e1856c4df
z6fd100abde5da7679375894493857e3cb6595fc09a88221df94b583f9916abe0911ef7dbb42fc5
z7cf5215c9a92f21678992faefe81d7a3ce309403a1d58b8f7403266722cae90bd9729f7764fd88
z1b153f12bec263c6de541006321d542942efa38e5f8ea773b01792ceef12524e8b7a6bd165ae92
z0cbcdc0cd472975c32ad4cbdb8e27a94d377e36796914aebadc0099021ffbf846aca71f8c47568
z5ad6a3303a98cf93d9139e26d31f990238a2a1b9262250f7b9409d59b583a35018f89a1d0df981
z467f717833d4f4fd5aa52e4e2154cb4ca95e2a173a1e9d11ee3b175faa56f2af06cc0a5b9aaf75
z52a9921e69b7f0005871ead1a93b63aae59a54d58925e3e94486a8fb432e6dc9c9371c571d70d1
zec976e5d25b3ffa14b045c55dafda218d6c39333ff739a31c1b6bb54c4f32c367e9a6ac0cd1808
z519d5687f101e0ffb8313da3652bfd9ead36c0a73f262242f1b457da6705fe6d02dbf8bfc3b75f
zb6a0c3ce1882bfade33d001e34f846d4826f150534a27bbfc5c113375084f555381a3997624c6a
z9a53343947ad70fad0329767dc3bc78579986fdd62fd575955674bd268f2bde48aafecb6267040
z41e58432f7bb8aa73a5cbe27c481b8bc1460c080b304e684a1aa08615e7521a9c43ab4e9e19359
z45a762938d1d534d7977db34937a1fae55050a113c109c1872dd6def580cf416f2a41a680dc3a8
z48cd61a2e1ce2e876f7e47b600029094868c4b8907e059013b6efd4319783791b54d4b45283985
z059a7b25c2ed68c5f18c3548f562e83e53e84568e89952de878514d37be38d154ab699b3c6897e
z06f41f59f4280c5d3305fbd66920190caf2fceed5f3bef8253a329c5f9c16876cba337a2d2a366
zb39ead954949bc2b60b76044c2a4436d41a9c1dc0b88a24c8ec0734ff3208ed6b627c0edbd8afa
z09ad82d96932e80b9c3dc26497d97d79fbde1a6bf6dab6d71b6a99674417c068fc4e1b945f917d
z7639a1328b48bce8bdbfd6c9c2d5c7d8aba6fb638c106f79d4fd609e1535b6829703445d1b7a04
z8a8af8a3d0b33501abfe5915c1ec190293251f3a1131c402357761dd3ac319e09e33e2237981ab
zed3c945e72dde4f0ac0affa293adb9ae03652b168072282e0b044d57e465c56c8a4c90265a354c
z23714465058afdf66f645c63b155194ed980e1b3159fe5ecf33e88e083ce5b0cad33980d302c86
zfdc8514c06258c203433f79c817221755df6568da643ced2d662af556d1292bc147d152810a3dd
zd94cfdde74a11fc39cae077c9cecdfd7cc38407920b845c7f115d9dc90a3dbeb249ebb65e4125c
z2c2a85d80e684cba6b8ff1fde9bc8c9c9fbbca65b41976edd81b6e5f74eb9cc444a467a078a349
z56db432212c88283bcfb1c5ad773e7fd28d132ec0477e605333754d56f869f75ae1ead8eb8f4a3
z18b14ef63444144b407f10940911c70298633e733ceb16d5e6b33990cbdcf1a8788724d98d5c00
z51d28db025f244c9684fe1f2f2937bb2cac94e1e8c1a578b99ce975ad7f1f68376dc87c473e8cc
z48c35d463a55ff2fc8f7aaa1f0d3ae5049ff25f29ec48e13282db9d9e58f43c6490e9d08086df3
za419bd5342a1fda85e7dbb33622ced6e2460d9c2b2e2cf884f0d504e415ee9753893189fa7add9
z08e475b54219d839e04faa705f741bd799d9643c0224233dd88c4c0d535b9c67d0749ff5dbd367
ze9dae75db559deb4f83daf086ba97fb731f36ac180b9b1642f902477b13d7f373941c815cf17d2
z8dc6f21b471af9f38522e412baea313839022731904dd0f11a2382f265290b2ca7c375e4aa4953
za73dee160c34bb9cee6a3631168621524f983ffd0b190a85c9ea283fa5f2eac1976a5b3728188b
zb681e7f8f93edfc091ea330c5caf0644a10582202f207b83b1c7e3f24c89216bd4836ad770993d
z980264402f1be2c080a1f708688702139956a80db1b30aeea7fa2f3fe4553e358559d46e60be2e
zafb10515552384915a9b7da7f04db43003febb2573a41a8f9a0f8ac66f13be85300a8b2ea6f84f
z4455da3f9765fcc85aa7ec330aa8eabbec04e7999bf17beca7eebf1a7265a3e89bc7898b61cf3e
zbcb0420d1aec31d6ca5efeba598d8b32258a5005e75abe10d582f9739be3cc551f5a7bbb090db5
z122199dbfdd63beb0d56374ee0f86124a8c537a49af222a1263431d4bf466652c5377a6ada458a
z8f0168c5270022ec4e176df3cf8b51d23fc43585cb5bb986b0625a08323efa15b39043fdddb3c9
z5b5a1d90bd5d2f92ee40290f62734edc597aaa1eaaca9d7e30860e08329a4c04438ebdb80a55cf
zf11aa60ee6de5c2adbfb768c892aea99e4606a640cfc3e451f22d211284e1cefc95f0c3edcc633
z5d50055f9c4f001a31d586859a5f18fa32ffd74abb763f977dc66d2d3142da6c39bbd651296cad
z82a4e834c889743b493e68f9d6327d19d63fe802ce541ed56344bf4dcc2843e5ba7bec0ef372eb
zdf9884aafb58b9e32d222b1a66a75df3db2a3c20725183b8b685111862abdd2fef5363acfa3d72
ze8a79c1d6b3815be1999c2f8d5f838b0b6a7f59cde6bf2614c4bb2077636b0c86a59b05a775f6f
ze6ce2ab359d2e03d81078d6a53b38c6eb737dca3d1121970076431c0bd96c2130453202c21c61a
z8499f41c6913270bf22856df8085d0a2a00f3dbc176cfbc98e4e1d6483e67763ada9a1a9c7f44f
z006ebc9f8570564550eb335ac18a85b8dd28e5f6527553d59bce945ed89c76bbdab9594dd1fc5c
z39540f73c88967ab3fb2c009a1871e479a64c90ff5442e6cf1cf977be67e6d3d69347db3288602
z55a814b22e9e31bb7be84eaf1f8a9b93d2d8abfd7b078db9659e2e104e09a5a0119a52045d205e
zcf2a4e551d8b2ec9dfcf3fa89dc80b5bb36d8a35dcb0a7cc160d76aa4672066d8593571adec015
z9f37a1d8f2a2ac2091ad1c060f134eb7913e924ee4807ee1d554064423774e9df3ad7d82ac5f03
z1c36e57587f2dcb780c7ea67e67901ce4972d732e5caf2939afbe1744a843aca88db641c31bcdb
z4182c47121693e279a5578ec072e104237ef8695bf0363953efc40e64170ee68dd6b80ccebaeac
za715a3dd3e1c5c59f869393d5826f7cd8cd80623d8502eb74528401d24d09ffef4ef4ee8dc4ea7
za5d2a842e2509803448e888083e107eab07b41c195ec2acbea6d1d8c7a7cf8d342fd2cd6192791
z131a87bdc7b6ccb2856677cbea83af41011b36d3998250b53e9ae85d7004a12881f3eba70bd71e
zed7f262ef4e9ac79ac2723c47a2df08d3628d85a05799b13c9524f658450123f28035e8150bcee
z37a62e0c9379587cd44ffd6a26b4133202f66c43a61246249d9fcf8477dbfa68f3d4a5d6ed9a6b
zd3eae9c16e6b6a3da388f246600b7882100e97fd6cfda80beefe154e18ad1ae64e3b9a4eedf1d6
z44f1c6db9b0218e14ea5ac308d433f54d6fefb8a5701798380c1173b38f2c1052576811e70a16b
z24a7856ab0acbd89005001184e9fcf3c338e9d7f7eb1523b20a55cec69664fa4fddc8db86e7821
z95a2b6e02ae6db931e0097d59679a3058601ae970b2901e27016bbbc7a05d9dde0c0e174fc67f6
z1017582d308d009bef03de0349bc342ce896b23af46ac10505649537216bbcf2ee77e60ca1b77f
zdcc3edc984714c06a56aedb16c533a746e9a489fed1f239493b2f5e7e1522d7ee9accb05cfdd03
z7de0d1dc236bbca40b3f88615a2b8f505b9bc08461d3d2fdf9781901d6a94fd75aa91712237112
z5e00bd9ec96ca773e0e23b614f7cfcebbe935935c648797a9bb0ebad0c0cc3c1b621c252c640c7
z819029275f23765a865d1d518b8db0f559087c314ff5504f5d4588dc746cab24803f7293419544
za1dc026465752749fc0daf6f1ec1613b2f015cef7bc4f5ea122d1ac9dce4088c4eaceb07af36d1
z30b0cbe9a665bf7cb519d2a7b5688a44e9e162fd56a8157a6aea8ed230106331eada464b8ab6b5
zd2e0561c89d151686078f8583de73c483b167016832b16ee11e31c60ee4ef289e241ea2e14892d
zcf127f51f1908ebcd1dbcd16e08b586de97982cf07dc9f30b3bb6e94cedab3b835f90c8a93a060
z5de5a9ac97cb5fb84ae54705aa81628124e6d50c4c20a78d75e1cec8403abfa7932d8235968877
z08bf542026fbb09de574cff572d14188b6595b25991a2e0150b7ed9dcd20ad6ad3e6e7251e86ef
z51075c0d98f94090e7ce7f28990c944fe070d4a9d80db0d8580082e6361c58b55ef886b67c8d28
z1841e5dc8afd6d9175ba194bfb07a5af721a82d6de12787ea66de370d30017f808698bff151d87
zaa27a8ca2611be7359fd35227faafbcd7bde75cc3b04ec317a1742af376602d55aef7ffebdd513
zea4ad04b2810557591dbe4888147d3a2efd750e51a56f6e87c7d111c703ad002ca525d59dc3395
zcdb0c238530faba89391dc7758a97bc10f42792127b63f40be8f1544d698fbf44eec44086c864f
za16abd32f00c4b7fc928e24fb3bb840d182c9008c5eaf87c917f575f961d14505c59c09f7aa86b
zc5c1cd43623d2fa9c6806e32c867083d7512194d5cdf4809946e462532b6e19c174ea4097ec640
z307d530b0a988de2e7066baa237360c535e6dc53d680808eaf42de1619f816016a0574b80d9de2
z6cf5491c372fb683d6079a9449948aafd1f098bb4782bf327a0e26379938514d9b97fd64000773
z73c8b2ed32cb4c6ae9ab8dea4a3fa7b89bea5275a1ac4a41658bbb8c2fe29df5990b00a610abf3
z32d581959a3316e992d9182a8f368a223934a693e1536998357d970d9e407ac5975a56214918ec
zcba239fd623f2a9e86166259e8446909a6e2d31e36ccbcddc611ad92cca2b068deabea52636f16
z1bd916db74f38dc776036079557f30a64728c6ab7c26c8f77730fe7fcd2a21d3dab52bd2219e46
za04092c7b37ce92e2e62be7e21f71f41ab663c7e058fb08975660f6bffb52d460f466dbdcb1402
z35407cde1ab5b859472c43b1a2cc89482d77c6bc3cc73c9bdf9ed8a24510b7b8301b457ba4e129
z26d6db2f37ccdfea7d7256f8f021110009af82efd4e07c40da47302b831792533bec56b8561631
z689bf0c58db39d49439055878fb8e1bac8e181441ed0a2fa22ac66c311cf7b476281c04a39455b
zb3a12595e0193a138be6df35e67edd3a45f33068b568d12b42165d51784cfdb859d6f18abbb6ec
zb1347fe58fb08ea7ddbf5caac0064131305c8b00fa2ff0a04c2bee0110dae1b5a39c99e982b2cf
z5d916d0b8e439ad9b31c803ab4d84ac353acfbc852f697b9d6c5259fa7d60dbfa68ba9d29e19ce
zdfa1d3fec8149480e0458f30ec7a2787998e166542d0dbf1a98a620f4641856d943b0c978b78ce
za54cefceca35f12435719f6e3b8172c019ad3b2058b338709e2f3b0fb980644deb6a38dfcb74a3
zf76cb4aead8f5b66e9e0ca3995f3cf792205e86cf0a4a11b4a912b151d8da05972ce6685b1becd
za89536aba824d7c7de66528d30194e89f6680b34ee12965139aad5c34a382f471404b5165fdafc
z14c5b29bfcef40b593fcc8f1d9fdcfef54589e9f2215e1eefa0199e6f54042d6a63d3f2ba8c10d
z8d93e4fb592cf4eb3d7df321ac3b6ab3e26d19c47f1a33049e75d04fd465093409341318960c5d
z0a3f1f2f520ff57d26377f5936dcbf9bb9af8be7691723bb16a7f2bf7ca71dda896fd60eee1169
z5ffe7d4ead06f64b08fd3ea94fd49560d9edd94e69e9b6b7eaf7c53777e7b4cfb7a5b97482e3cb
za69ccb77b6a7aef75d8023646a46447a796500a2142c253aad41e70dff5a65d0eff485da9098dc
z15073b3613b2b1594b5b99685526d7062635b99d2fe2690e757aea6660ee093360b57ba13ebc6d
zd76d7c3955d7158e0e1c34739c7705903fb286887e85491275b28335353486faf43d22c872ff3c
z8e76687c493772fdac5827807c3c1170287ef245ea8669ee173fa3c5911ec53f49dbe026b609d9
z25c7bdf403ce57557ebbc2c3af1b41e68f603540e0f31d16f85b40fc5e618455f771a279e75c0d
z731d90520025ba829d8a60251e797da640134099cd125d52c65ed12a421df4ec8e341db9ca77b1
z9377991e50920ed872dc5d909ad41895242ed2519e3504b261e5aebddc2383a560155da47c053c
z7514ee29929328ace2631f38f30b221a23f5382514050210da3bbb49b56f053070d2fde2529bc1
z4a5b7205ece849555462dcb9afbe632b358923fcbaa430169ca4f1ede941458a890f948bcb6311
z95c8a8da1e3a7948e9cb88ce34c73c81dffe9c23e95691a2a0dd3914107d32c0abe7d759defbdc
z5132aec7e5634a736b4b0e38f80931f7068c248564c2a3b9a3755937d4ffcdafaf2d387d76af22
z8766d38199e923ebd2920ef2337cd15d1fdc189506403d24e848a17a7137fb20d8ba108883dccc
ze4317b6eb04f29b57a7930b584d19400717c3dc580de7a2985bc49fa627b5d426d297eec7e8af5
zab8c09d4e0a6d9351441c2eb4efabdbb28d217506912597335a1b655841ee429da2cd4238b0ce0
z9ba9f68cfaf666612d5248bcfa9f2ae53be3598ed6dccabf6e7e31400200abc8ddee587aeefe92
zf405f896c18a1a88a1605a8ca59f20e6bf0bfe2c56b46412499098438ae4b251c9ea694d91e4e9
z3d3eebc330ae04ec8c06316f9987ab36552f9783d5aee2aec89732fe8928f34896826bc1589f9a
z1e440fc4c3346a4cec54cd812dfa12466fdab29cf872c09bec6323ff7915b9d44b7bf9d5da3444
z4da18870391191594e42f8f6a3a31b4f27faed2d9002ecc61320dbfc38bc3390452020a4d3b20a
z221ea9d5b563222fce5e80c86619d6c70dd22f1cd1bf7f2fb7bb04d0e6b7b640d46766aaa4bc35
z9cf2cd3187ffea6c9007123cde8f0c3900b5913f5d5ab3f099b7ef43a26cc0adb8ad7792d57780
zd369d9c370131f00c617ccba8324866a036044f0ca6dc4648c0b6f61d931a47859a5364861d035
zb71245a5a9c3c8c4655782a3202c7104fa3078d9375b631535cf35209baa0456b71d44626ae709
z2d949ec5a650d27fdf1896edbb38570c8abd3a01b7b117e70250da71216641b5cf27cf39e95d4f
zbaa67e7e5b09f35039e1d4dfd882d47b557cba40b32ee9db3087a0667096d554cc975f33b84e82
zd53f28903471e825874dbedfe6320f784a8a3811ba58724236e01ff5e6775252257031c88a3a8a
za5fd17c5019387dbce92d990d3b0e5bee166c5e1452fc6060cbfbfd0f9886ddfa643b045044d23
ze0cb9592f87093508f7cd383620769876df345253134da69b06cf2723ef522ae1004eaa3950c5c
z137e86feb6c74c7d58b66641ee03f84883e99d80e90f5ae8dd463de921b2896e851d0650a57543
z953a7e0509c31c63b992119079bb2243b2c308bb958fa8cb4fffc10ac7a28cff2a796bd284bc91
z8f76f04ced4af7730f5ee641cc43f21dc26e69d4f1db4f1054d8e2b78b9a92407c6ea28f11efae
z1bba0bb6818e0f74c6d853544bd8d19fea69b2e8a715c6b8eedd6719fc79d6b166245a15f3df37
z59dd74a8d7c9668550e57324d0da7b5e7b8b86ed8f9634a234b5d44d83b98e61a958f19ede7836
zf6649e3caf47c9e0789a3b24d9e20a94eb58d8cc91988723766ff2e75b6e2cd907a3a0238ac45c
z51c01bdff6b25dd328d9629fd9c0415aab14562cf322d51a7b552b29e39d0d751f349857fd8bc0
z5d8c267f37292e67ae67b65d58b9aab48309e4a45b56ea2464cf5e573da847bdf792e678b5e90f
zb268fffab8f2acba304b774b7bd636e39ebf644af4a1f9749c28f7d0ce7df256c460e12ad70580
z116db07ea34232845790e103fe6616713b96f95cd23e3477ea372897a5f901880ea0076e15c2c9
z443c41d8817efda3224dc7434e1252b5acceca8ef987677b4d46b6b93c9ce277535e9645a55a00
z9b890b0bf34d74636c20e0ea268a58526e47ec51800e5cca8f609a85b5170668d1589a7151e1eb
z7f14593a5d8d8c16d9db390be307c224211f8865df3cbd1a672d9143153801365d7edcdab6a120
z1657ffcba0bbcc21deda3d212eb1870e23c5104eb4d552dd061a5f47b6611158bbbb2737435b30
za48da8ab7ffb784eb85e0dfeae9dcd0539ab6c998425fdf24929cf602d9b7b939c4a46b31a2fdb
zb48eab9ccd8614515add47b9d6ecc274deb5f755a972630cf6d21b1b95052fda0ad69c8eedaca6
zb2ebafee60840b7a5b9647b4451b62cfb088e1bd079a107fdb36d4a22abacb21f13e18a026d907
zdcc62886a073c9debb9594ad228e3a655c4209b2529df5abb7f357e91a00568db3dfc1ced9676d
z2d872be1f44c7d2f1c3a1e83a5f0af06965fc97eb8e25eb5210aa495356d535095edf28d105b2c
zb86cc68f33f82ce4486e8df4a76eac601f2d8a7eb09d6f2ebd742a52c3a5e4f695ea05a565ad8e
z9fbf4ed2d8e55b514564f1aa7fbc51f697ae477aba5bb57024c0b9317cac3ff9e3cd1bf8a120c5
z9e53d035cf30792441a1c29bbd1fa1aef3f12710d07d4883703c014f8db83bf0e655f801a9038e
z9aca951cda8feb92557d6d5c8640c84c24757c10fdea9b98136343168404f8a5ff3894c43031c2
za4b3e6e6d9bd1e31664278e3487796041a9e95131218b71eb74368457b81c34aeb089561562471
z418b202540cec38dbf4078e589d9e1e65b2cbe9146061ee17d1cdee7eee12f758208384c1ad250
z53bb6cc6d07f2fd8c39f834949f00552f95d13a781e4ec4881e9adddf675aecdb84eb54ff1499d
zadf71ae9f0ddd7330da0fa7401dfc69f14bbdc72342529a22ab725f16fe2a8466f223b17a0eb6f
z06206ee87bd3a1a3b5c9fe15b66e40641f27bb051c5096d5d4125f827bfc0256df3bcb5160ac4c
zc38300e81986e38dd0e0641fda5b8aa79b075e0e61eee79d394be461caa8079fd1b4cfc16d6c2b
z86f3f253c48a9496e5d8d33c247906c4c7dff5e087e5565e05a9515f5ce253a3e031ecd5897dea
zc522d73aeb7aa83aa3af6086e98764aac87cd17642b14e84fa5fd2c32f583a96c882d39e61b365
zd0afcd49a5006bf970e80f1f8bf17f17c30e5ad4e751144e162fedd88f8766ae58d8473f0380b2
z25a40944642d5400545e90c2d8e33384c23f036a668a0865f501ab5c02cc8ef68173954db014e0
zc5c54bea264c1cc0bc78cfc889214c942e50469b895a99186e2b05ff9f1866d0f4bc538b65862b
z60f0d0dab91bcedd292d4ffbc9bf65077ea6d7525c997ffbb884037edaeb477f1ff5756e6f345c
zbe0a83507983f1b378cdc7beaaa5734933e8a0d26f69ae55ee7a5b949deac08c3244982d38747b
z03dc4b50f88a42e5dd38d88104540b9b794f0c4d383cab976f937aa0badab5637c63ac9c0608b9
z9101209a0a2998e18c26f1ae04db91e934f3357a524cb5d98683f01c85a4eb96bccea06acb8f08
zbc7f598c52cfa9ff9b2a90747ecf9f42e94bbd8b11f4ee8b2d8ac02fef253205e5466291326d76
zcd517008cc093e8fe8e668c1ac59f7341fc67e08bc1b87371ce4834fa54f5441f78037c22fa4c5
z9f020e6041fad28242ef5e58c8e9c7447585cf16281b3eba6190ed4de7801af7321d569073f958
z0e8ee63974a695fa0d683649e4b7bbd2c3448cd97cd12a5e2610dfc21de2bf08a901b629ae0eca
z1e0d723de190c70e82030cd042c583cd739a668144765cb78d2c4a9a71882c4844d1d172cfbe6f
zf3661b36a75a801a9a7c6fbd8bb86b91ac421887d8744f42b43d3b34a0661b85894d7061a25f5b
z324027c53a40d0e2e3fbc4a4326eadcfc4b945c04f6e63fa90fb3c0381b8228a9b8c067cce6df0
zf35f7cc713c2dc92c6169527b75645acefb25e0dbc24eb05f50f2d5bd70e4aa905ccbc3bbb9f3c
z12b11b6b1d64cc023790326f1aed3863261caaddeb97a9763cb11eacd42cb977f8bd0d11a3c571
zf0d54ae1574da2908dd5ed9334f48ea4dea35f5e3f43d02e728007efc69ed6a69e217b6d705637
z3dcc050a7a9d5a4b26a2f40c7cbf58641ebb677c71560381dab0d77c2ea541708e92a5593b4c9f
zdfe5d8ad4f5ecc6a5504f5276302b6dc57f09fe0289d4570852218bf6f9c16de1f4c14f1b0e954
z1e8fdbf7cf9ebb8ffd3a786c4fa2659d2f44b470f86823e39c657a4b67306e7fe357604f4f1763
zd8477ae021a249adec8ead152c1de66533e71c8a3b2bb5f9e86368bb0333c003e21de534e24fc3
zb5eaca24afcdca788e92cdcd1d8b9d53a33f0f01a2197f91fcabff366cfb42d6e790b485564adc
z9999641f03c812dadc6c3ea6e7f28bcc1c03e89c8e43ebd5b45e0525d5a161a7bb615a2da42e78
zed19bc63ee5ba68f82ab377b3f8812602408fad735f1bc9a73f9f0d60e94fa31fe1b28da05acdf
za89959a6c4812449a8c4c554f2c95fb2013660f9157481a4a8712e58669f461675a2b35fefc3d9
zd390f052b4dbb5d20bf7495ca51cf7bd7acd5ab403efbd8ba7094e9e5d2d8d25c3a7c3f55bb303
z0d31fb5cec7e9948ab31a91e9c377716c3a6e45e13ae9f60ec9bd66d211b00b84d08e7b214608e
z5050820bf688e19c8ccaa0f1d1ba531890473f332655b097cc67f9acbabc074d7335789a79225d
zbb45d78aefd7b41b20020b126e9e47575c8ee324f0cce7f5bbdf6e321ead3d497325237c567c4b
z754aba2cce424e7a823aaa745f63729adfd0b21de8415ffa7955336d810ddb704a550e81a5fcb7
z47955dcc093470d8c53f8aac0a67fbaa63d84808bfbee59b3f9e8b23a174a9f74e98110d0fd767
z26e0a97cff6c6c169793cd0bc21b7b40e28c4756a766ab277a2a41a15d08ececb713e64bde3e4a
z136a7cd9cc02f2359dd772a7faa1c35293788012376ed8a466f3976cf7c357c58b3256f3868e59
z2b8b682b1afe214f64b8717c882988df5e4a0ceb4f0100c7208b8067be0ca9db08fcc9762b0d88
zdb66667c78e620b9356b632e06d9bf46aa6969e7c47e38bdce9886c7b27e61a06e98bdee352754
zcf6ef9a117b83e6f1ef920474b9ba1a1e159b2a8cd45e5cf1c06e0d552bbd1ba1a02fa7a61fdcc
z3d756b3cd162c9a017843fc4737272eb77064311dfcfcae6924da3f95c087fa548e50ca19e60a2
zb36776630e9afc14f6418e920248d7ccc0a4ab0f9bb883d5e946e829b263d55e06de259201516a
z638cbe613da302bfac37c43fad8ccabbcd4751a01955c6312c25a7d02926cc0f4f018c563a5a4c
z13c40f00191cc1efb4305d1027655c4301e2fe5442ec29fcad6360e3c7c6271e7e772b775ff05a
z0928af505b5a45841d363b421ebe7a2161b604641712ff6fe171d7fa84fcac0a93e2edabfc5beb
z1385bdc28bb93155dc8f86253f6c0093a9444e29d63f66d043c6928753cadb4ae0ae5c72e58cff
za7f13dc8fa40c02e3a17349cb006ace3d9e19a8cf5eb20456028ad3b609e679a37cd753e44593c
z0df539151f6d9ec5a037c0f293d7b5fd91d5af893bf260d336e972670ad3e5c8e026e1938b3e59
zeeb25c5c957e976b4e0658a19c5b623c406c9d9c30fbe7808f90ea4495e04600c55953635b9767
z4c9014f5d3c0874a4da8af643ce4ad728ab8e33f27fd4dd5685d9ad9a176b3c090c72f8a3e3a37
z7131603fbddc720135bebee3f911bf04babd7229f49290d56eb3239036ee58886c8d5989a8f2fa
zfd7f260d047980829b2f9bb4e6d264c37e4c254c91950ec4237f9c49fc359039130b31efc289f9
z6c75804ddbe664f98477cadca7c3b60c24ec64db6a0a089eb4c88218d92dc24483fa649a51933f
zeb212b9b3bf85dc40b84f7e811d5d80204e2dad8b982c4440a020a692b1de1751ed6a90ada59bc
zdad58c00be85b26e5126ac9b8cba81623536bb33801ff30a0eee8505720694198e392b5b176df1
zee22dff19cee61f369187f626348d8454bd45a1c6d5f25656ab5a7021cf78d2ab0d5bf6a3072b5
z00dedc3ea7dc3a0c5ac1765b7612a4d5be6b89439d3ffb5004d82a5463d4b89af2a00e4841c9d3
z5146ee6456a2502454decbbebb83199c3694f20d7a72f0d1e0f17f392f9215e4f1e274a0d83c5b
z4eb696691ec0aa26fe67869f84bae7d022f9b42f30aa4a2404a28c9dde371ba62f333d4dcdbac9
z4939e64a996b560da289bf6da167eefc92de2c808ff44f6369556ace48b7cdb9819661301ecd13
ze7c76d038157c61947b7323c0643730ff9670cb1e009905d851f6610c235c5698d8d5b8420632d
z61bc5692978f548bc409d1127e6bbeed15faa8974a269301fa41
`end_protected_0in
`else
`ifdef MODEL_TECH
`include "qvl_pci_express_link_pkt_parser.mti.svp"
`endif // MODEL_TECH
`endif // encrypted_0in
