`ifdef encrypted_0in
`protected_0in
ze74c34e226135848fe16db9ffd31815111b6d7fb642c521a3f628cf6da949865580b22efd062a7
ze90adae0e65e66a2c36a587d0a790699161455169ed55a01f2084f11770a774ec4c588039b380f
z6de9c5084882a40b79a175f5c2114b2b6d78b070cb806e1c0aa9258297f4687ab308bc470f0040
zb0b1de382961eeeaf2e279e1462520fc31c119af8f2b214846f56c2b3cd2eadbe4099496abff18
z15cec83ec4a77b868344aa20ba7360908f5c0de2a79abf8b3534b883bb12180f68b5d4beb444cf
z3fba8f13afb0abfe8fcc4294810f75afe452434d2d0f1166236c82f76edf1e12979f04bc35693e
z32ae028996dd85737a8f5adc1ebb94f39c940246e887647b64782cd7ab429b0544c173176cede7
z01dfb26b1f73408344a52b7e1f117f12bb9c8077b34876c2e6fdc085981637012dc9754765e1a9
zc512ce062e0b8fb16a214591f5c81e1353b900a611fe1f4886b57940b41b7f2ce99a7b84b04b90
z916f717e73bd10589c81e207ed77ec660a8cbed5b487fa50acde1b055c8870bd8676023f21ddcf
z9c98cc47cfa2d654ff1365d1f45035a045a66c5dfa82790502623b57a3af03bf0f0c0d35b51558
zb8b5f2d29acf03737a9ca2a053b7a8f06800d50b465c41b30eb585f62f3d0c2c5a43bc21514abf
z7ac02451dcffc82eb9d993428d8e99929d06dfe4c7df23c439d3461190ac33bd7bda7144a72e4e
z44a02555bd042b3947862c7dfe7eb1dea15c73e0d04c1e1744cf67602aeba94a629a4058ee2044
zec841de49b48a7b4423c72fec39ac876c8ca70fbf0da6567d72386ace7ebb71c4995783a8a8ef5
zbb1c1378ba11f73605b21c3a7b9f78b6b5189c11ed3fd44e4b0cd5d7ea58afa2f46240fc1937fb
z3eab4061ffb535e64b6303bbb2b1ae9bde93b0354e550fa907ea6eff82dee5ebdb8e3d25f25aa8
z0a43d918c24118a99aeafe597e13ce16d1b17c556b5adac8808d66e4ab4b01fbb80beae2cfca24
zfbfcc5adb90aaac4fa5b8e7a33f842889c5e665813126313ddd2df318a3eadecbb8a4b4e2487ea
zd10d46e36773c7a71e55db87ba824e931ec24c239cc7b3e53ad93078265c8157e72269a40939bd
z39b680a2eaff0133c95370c240d8f85d675aa22e5f08f1c29c774c4fea5f4177ec7fad22bf5513
z8e41ccb623a3c04bc1f7a6c0851a75b328d95fea0203a26e6115f0d093bc5e3c1559dd4c8d80fd
z465a02c5aa1571be8724028ed9043b8e537b8a8cd08c083d202a7b3c209eed562f595bf89ffbe0
z906fa7b19944d93c8b53e92bceb34eedc1d88d0f05bffe42cff19d9abce86070df11c2a578e831
ze434e1f8af310eba8236159e1dd8534e6b2045b81b624ccb28bb8344fd330c10e9191ed193ca08
z67c1d14a56331f59988718bdda79bec2b3bd96b9fec6ddba91c052725871bf2a06c28b5d14beb5
zbe58d48ccc1331becb2dcf60c588983bf56c4dd5a7afabf3dc7ae49aaab6f09447d3fb7734243b
zae145cb012127ac9840d85f518a4ba27cc078f0d2e521c23530a2aa44181486a082542ae5c8dc9
zf2edd58e1edd45a60d75c10bc581aa3b47e43b94369d6adf22642a71c3160e30cc93cb88fc015f
z33e1791e50a7e4f8a9df91070e45809766c7b1e79fd432254bbf59920e723597f568e71edf493d
zf9a495dcbf7a7ec6a47fe89ea4f52440547373629e90cbf5621ae07494d938256b75967c9e64a3
za3e8f5befb7fca4455da6897b0fcc22b3d23da2c8681e0b735b3a5b4a7a919542197a3cec9120f
z8b18b564209690b99ef7e0ce0d76e0b68bf3c457bdbdb4e6cdad5b72857527b9c69acda8da1ddf
z0a99f131d3a9766b76fd6d3686d09580e13bb35327d7630319fbdb25a07742d0abf18eabbd0677
zfb39350d0b25e53a75678c51168e5893cfcffb4f92557fe27cda73143d45f005b3fced474276f5
zda9507017b782f26a50358344c49fc06f147d53c2985738b3894120d099e48cff1c74a03d5c41c
zc625ee918cd106ceeac0d65ff78586d7948ced108b009099f1535e70ee1fe8c3a0f21649f28d98
zeeb4b7bc7c2ba18e963bae7964a7696589e94a2c06ab94b892a0e002abeb67cffd80d4e8f7d2c3
z749ed6031be2e38ce4782c9bde46e6da18f5a17f0ae8e3bedbc60d569521fe751b2e0b48430d2e
zfbfeb920222b919c8324139c5080f6b056860718e906ab5f44e5e7c56974d3190c4e9972aa076e
ze1448896a4721cec79e0b1d9a0505eec38db5a732a5de0b4a0575b3d00d750413304931366f21b
z2391549100e28bd3f6559036464d247c2dfc26065ad128f7a2a1b47014f47d32bdc4bc1ac6a763
z7e2362491d1cbb45cc465873e53c345099928218e771ddc24860280887f217eece1a8aca69ef69
z499440104c014c57741be72abfda1cd3ef98e13391277c4786b82c1d3d82f8ebc685b0aedc90cd
ze2ed8084f7ba2c0f2118be23f1f98d085d1393a878ed3923c308ce5e4dea3787e410e49542b6a5
zca9c32f74fdb5f074ef5518b5056b0849de398d623d10edc19f8d22ae004bc20d5361b2fefa4de
zb5ea941a05c1da25c7465764b7ee4ee52e01be6f0858eb92ddb0e6e8599a63a1c213216756bc1d
z800d1a3e7a8e8edff750328b6599bda6e1d39608789f4672e1840f18616c582252c7b837d3b557
zac7f006d736cd226162235715b3f16746de7445d61e8209140ca5ec39dcb869f7d52c0c4f7f647
z8ad87850e6bbd6bea5a89e498653b3edb2d4bf38b3e7d865dcf5ca2814257133febd156768c60b
zbcf58b89f5f47b5723251c980dcca2572c8a6a08fcedc9d611a926883236846a650c245d18d531
zd4fb2fead1b334e3541cd5f55d1854833eac4ab92a0c0f6d6931996eb02feb5516932eb60ebe00
ze2be52b7289f5793e7ac0fd5a721f08ff6059ce9e2a430dbceb4c65e87fa11638b122c94fb362f
zbad51d8e1d72e6305aee671368e7fb6fbda6f6f75c409ddd4554f2822da8c51dfa712775bbd4b7
z0f2179dc0eef47eaea4a3bbfe4145e619be278c974e6eabf245d20328d6a6ee1f0ca434a3a5621
zd53b485bd7b2aebf84783d883577f6a1a2a5741b305a93adfa4249f19715af5bd4d57296f72cbc
z08ef9b74869e9e56ebfe57f0e5c20f5b7c89fdd54ab376a25fbb8a1b47ec6535d235ba527dd041
zb58330c590ae9a8e01036f2808bfd78cf00b285de609ab9eb17a6cef96acdc7d688273ffb21359
zce5490f997b7c8c717b1615328f20a417f21fcd81a012b357d8e130c432700a4b3b42daa05c0da
z575d11b294fb8086e74e85b45a8f065967bb1d45431b34c5dc3c845b43af3be3d85c6a024df8ef
z698494c7801d56d883173fd16c196c2f6124883bb4f60cfecede69b8122c60e0b95c8d442f37f3
z42ea2679e1d5449083244ad6f579bc3fddd32147dc62933af51785ab4b1bbd24f2e08b884197c9
z6cff369bb16c64f33f19bbaa531fce177847aaf4b7830df8f1debe783773da47e9db5cbe3d3d9e
z0668da6682028f8bad8b30d8be9368feabb560fd531eed4b4ad361f6dfb7a80019723e4d0fddd4
z74acad4a6eca868d7476098cd1dfab2ee2dc03987b0b1fd1f3466f5b702e8616814ec14cbcfe99
z03a69dbb1618c9433c1aa3add24a08791aa35b53ada386dd6bbd9d160d5ebc2fba0e358fed2224
z829987b9caef51beb39613155cc7f9ff14b86158cc6725131ee8ff4ef2ab31f2e8fffda1900a61
z1c2e38d222862b476636810b5a245c2a7bf6025e3280537121241a1a108bbafba0dbe05b06949d
zecce07fa465d74528fbb7ebf2401ed0709e38002f1bff8844ab4074ad78d5514abd70bca678a03
z16b0f574946522f147bdd6eabafbbb1738f80004560a515505c38288105d14c09b2e45d61cb501
z11701d2465cd60fc6d5a2d176d3135292636a428ab58dad43ac2e9fcbd3de858074139e4c091ea
z92aeb7d4bef4ca1a0dae8f6b1ff17400c1e97bf8a41a79b7afd2110b5b4ec6039231cc9ea48129
zed007376deb751197eccc576218cf8f044de6c22a55ca6ee60177b1e3fd1778d1791bc896a9d6d
zff7169335a08f5f774e62690de997ebec96b6156645e3a35a8982ee82721b951f31e6162d03240
zef70ceb28359df4c4a3cd73ecd0f52c50a4d24fa11327399f5993ceece9a5847c35a3122aa5a58
z3beb51c7cd3e67e751e9e483c81ac4c400ce0af101afac9e6d3459a8bf831dcbd29b7f70b3a2fd
zd6fca15f001a1fac224f40d9e3794d98327da581a851bcf9ba558ee6ec5aa4e12d0abd04e5cccd
z4185f4dc2bac6a250c7faa2987284f1fed127c1c9f11be8abc4c7b985c752d3e3d437f3afdf86d
zea0ce97e6c5ab27e5fe470a9bfa6ec8b59dd9045d1e611b7dfe759503f55e2c740b84460951ee3
z77739131fdb1cfe34994a2ace5d0372e8a73c7302ac1d936998a1cec2eb34d1b0210b6c49536c9
zb8f2c299be9c29f09ed8ffc7f8c4a2a48ae115159e27a0c355be9eec1ad95c0481ee81432bdcac
zb9e20a77e799d2b555ba51422f40f5b6f93a6ba380662fec22bbb434b64ee9c699a6dbe833562b
z3b20ef06104942644aca5b4062ad41bbba78b1fe25038ea2a591fe1988efd69250f11a407b5b7d
ze723e24bbdb8b3f8121996c4fb4fe585be1ecf1b9a7baacaecbc35387e7dac5b223efeb80a807b
z33951c4612162a9424d151605431a66e7a05dc98faa581e86cf20f88701a54ca168e7b2ef77f0d
zbe7526ac4417b0998f1c6f6cca1c75975be6b4458a9a1f653de3e8c828fb1491f4b9178678b1cc
z73b68aa38e56eaf2e9864d6cec0e8b05ff0377d4f7578b9a35c5fa4e3bb1616fe25ab60b15bb0f
zca6e944d75d8ec526cc21e41fb1c27c6e0a5f700eb88f6726491a4c3b940cf173aadd79d73f3bc
zf811056ab4f7cc433ec0a9da7d2242c65fdd1654e70198de9dc59e7e2d2913595cb9322e87b5b1
zf862d8066b440f1aaf1d6fc8ca3e972ed9e04f8beaf98307c6c66a9cda6945e6a0751efe4c8bf2
z5f6dfed3ad6d8c468674c133d44392d71ffba00dead30d27d15081edf1958a10d4675f84376c6c
z12d43e5caee86cc793528d4e09186d5efd154feb9d402d0b88a99d4fb864f9494778ef83c18785
zf6572ee274dd3fd1747717769c0bbaa6be7db381ed162415ef55fe817a279d75d8620404f2f358
z62e350946b2dbeb3612f976c0da8c3872e30aa71d416e5bfb287fa3ad3ca61ebdb0f2d32db9605
z3d4f64cb98a94c9b299cf2a38573abc56c8ceb0676513530474f677a6f3e9cff2804bcca4d4e23
z527b428dfa39361af50ef855f0170f00f02c6612db878c29f6d526eb3fa82fe268a5d70d3f5424
z8843d54e16884823a0ad541849a04845557414908c1d4f21e85b1235fba69bf0c9cb4bdc85438d
zdec9b51e0756ad3641c7dc8b5edc005f847e90987f3f298e9199dbdba7b8c7f0b0124a9acbfa03
zdda6c1bee88200f5e7895dcad11f4e2959c1d068ad29fc639dff192f340b6d3e73cb472cb65d61
z6a6f5df678c27109c1d787f44590afd6c760aeb5cfc0afc0538e39fe1e3943f2607dc9f95fba54
z4f3ceef35613a564f048b23f532f95d4872924c552b563c75b6c14a3f005ad8190d43c1e4b00d4
z880acbeb6f7a5db6b73eb458820b650239ebe59062e827e75cb5429ee97ec2fb7a61d988976f62
zd0a42b68edc8c02ba466cfe433357c40391823ec69894763e75f3e25f36737fb5f72b0e11e48cf
zf4aa93539d651fb4f94d8e0421f07184b52a39ff86596f1cfd36ce8c2ad9bc29dd5ee6f657f7e8
z624539111cc7983476012a3b75bba9a23735c8086d267499277cc441bc664b608499fe6ab16bfb
z174af20022a0f6bcee46a1afa96142f9fb3f42def678068f593e6b19b4c426f4930908163c7025
zd7f01c5556837908d0e25a97a58f32d311022b322b32e85f8dcd8063884cb3f923bd03c6d2692f
z4d9909ef3738e2d7d16ca789bfd3152db2018af7b6d6a54b8c6aaf0f78fe67078e42e6b79919e0
z71457162a73a16ca2dc00663ac2b80928a9d53c614288c72dc2eb193a037578a177f1686cd718c
z4e42b66ef5d32d2db0cdc15cf7a712a12e8e8ab3f41f9f89e22b3bad62018c9d5f594746ef90fe
zeabc56f9d6d25b45ad9060e006adcd5e5fbcfc38e7f41930d18f294ca0a2201bf3f9959d2028f0
zbcf497d0febedb7b34faa17902d5f2e245e4420f15c0202c933f7bbedad29bf1d5af619b3fbc4a
z8af4d4199351c50981c00d9a1ab565bde083f26fad6dcc98d3162407712c5b792923d323f66913
zea976c3cfd8b8ceb56853056d718f9275ca329ed2e2cc26ebf4e13bfc16a24c554d83b25db078e
zf693c431f97cf9b52e6b0e4126489c55cc293e44f87b93de06fd0be668e9d8c962e66433001226
ze9bd4cde3a47e28af6bb3affc265bd11211a598bf63bf3395f6c4b335e86d7eade755e2589cfac
zf74e2029aeb55b81cb576c3101cd3d70b08e227a8b832a76138eb71bc9b5eac127690ae7c7646e
z8705617858f1a7bc93c699155526f133d7c0107410f6bf1b399d67b0434166bb0fdb036deb21a0
z86c5264f7604ba720fae0163bad8d89381ae60c88f59b35a73109ed432084c9b466b56955a471a
z35f52957fcd9faa21d91292783b3378d29285618730577b2906d28e0b44bc3070f2d293a828fe7
z0e8ef15900679fb8098da4634893dd2d42f0543ba481aff0a9ae13ac545849c2cf97c4cb8b5c11
ze0b24132531518a2bb4efde6846341c64b06c5373d290e078dcbbf750e0098cefb74a1060f8b23
ze2a78f7c33ed1f86d846b51219421fbbdfc7657b7a2d7f9bd2fc0e68997fd905d43d5f2f3f6d32
z2c537625baad4b6dcfa1f87689629f6ca6a28a5d8830b2cbddbc07b1adbf5a2f734184a9326b5c
z6aef6e7ebc57427bb5daa4b7aa2a117ed01b493e4766dc3844321b7b8106e6ace0c923b8eb8612
zaee166870374426a5a31226a97b5c6d055396d8902f3b4a516c0ec61f27ee54a70e20f85bd1dd9
zebc5d3acf9c45097ca144069d59614d460079561b87bb1a2b3c4ba0ed2d76e6936b8e36569eee3
za54599060606e05d75d736b0f921f995212784350ae68fa23d168d6d20b0ee7d4c0f8a61e50b4d
zdf800d84c00bff1ff25f8d3e3d9e1ee89e67295ee1b66770db294bd89cd29362a7ed11c9767de4
z2588568347490e5f4b930b77d0cd98d3455fc9e973620f8cf65c4d0dbeff73d4550ed969002e14
za014d3e6b655b704fe8e98eb39abb31a134cb17dea045f8e32375740f546cfb9713d297b80014e
zff2d3f99ff3745ab1c945899b0b8fd5585abfac977d5850cb9c88e2614104734744d5c6e1cb3cd
z7b09de73ddf937df31817ec3c3fbad8a8534f239c5d6d9282034dbe9eab7896377a851e30105c8
zf5759777e8c38329b6a2327255d63adf0772d30886938f9ff3531cffe9b9e5abd957fedb28b5b3
za89d953d3e67f1b90d76b2c2cbd0b85d15be9fdffecfb2fc77930d87b68fc94df48c96a821afe5
z31823a6b7b3a1a5a2a5d6cd548dcaf7edc51679287e40bcd9df737e90f1ada8fae3d153f795b2f
z3b51a4790092c245768717c034cb9dc996b476fdc368645d6665d2096d9dcd1c2fa03de58acb0e
za2853757cf6a2ee9501658faae84545243a1a0c76baf96a66820aaf3d76832b0113641e0249bff
ze77166fde40c02a8a7c65df4ce992b0ffd89d83efcfd6833e2b28c960cda5fdf70e77089b9362e
za0a7776dbd9f032618c9e47937a0a17d9a5723cecd2125a82c42c2eaec8ad4d419e0dca6f1dce5
z775f498482736a7c8f9afa2de0ce1e15e304b63372be1ab96c2e99e5e4b109084a2a4eb6b337c9
z002f5b298235497fe6801dcf317c317a1b76cd96ef4bdaa72b824f40bc8922823a0783483fecb4
z6e1acfc5b305257b3a30c5c6a6a157c14a45c474743132d581a40bfeea475c760d5ea6eed74fbb
z4d335af2ef51d0721ba52ca8ebf5a7dfba439d12cd5937963de16f68c08d69b713c37e1b520f32
za6476dad767f7bc7d3439e7082a452c763512106e95002e70877d8911abc09a8f30bc08c95e549
z2472550a141982122f8c772577796165915599cad2bad5e5228f6196397ca70399ebffff6c1a93
zd188c291bfa40cf49b222f8f6bea52f264d2840010d03e0c90bccf3add5bba9c04e4c9897662f4
z0c5dad1ac5bed36569b639246a9b5974fce0840ac63783a99cc26a15e489d730f5c518ecfbf6bb
z1b4a7b3a6093d0585c4237b0f3d0b46899d29fe8d2e10a3e07a7aec8b29eae59bc84d73694fe43
zb20d90baae63ff4adc86d180c0d093b1fa9c622066f8d454eb94c8d3ac49a9b58c52e532ebeac3
zaacda42e88db2e64c5b98e86f39b3e4e40a5803a95a73b9623e262c7023524e331a7e10f40597c
zfc196013471a369dad92e89c0b12825ae7323736ab11e7ad084f2db4dc9de36a12140f98e2d55b
z0dd37d70d7dd3a4dea67e1fe5d6dda8767944f0708f2e345ac0c1fd2352459f32d262a37279773
z3eb32db60361436b0a3b3d3ad88e0ba5c55668100582680921265261ec0dc5e4159c4266121d2c
zb36db9389ccffa332f85a8766bab493e021fddd0f9848f37594038260bccc57d3209bfd823f1f4
zf1aba5b3c31bc3d7ff8dc83a487c5ae9dd63b0e79553dd08b95a76f1da949693fb0a9c04295a8f
zcd1c57f5af7fdc88499ef7305981a3c0ccd1d66b42844b53e5393572d3d3bf88bf0f4b518762d2
z1b65166c7f77ed02b86593fbb56f376e7c57041ae80dbceb4bb5651db0b60737c36b5dc292ee0d
zf086a65962ac6a1bcdaea7a7766f6df806a6de952a10245b21a42c7be4b3b0cc60c0e289a496d7
z710f3ae22088473bea855d03df69bdf6ba4f8723ad0b1d33a55fdd706dc77f1a5fea273435a2a8
z18d4ef813c1164d838ca054d80ac6fb6481336d7877f582859f450398db4fd27538321d7759614
z31fa725188590d22b90fc4034e3ccffbaf98d0853c22abe0a63993b2aaf5de4d83106f6fa64c08
z2a6b76810945e66494816038dbcd6a6acfb7ad981f0683d3ebd32e0aab586336903e123cd46099
z363f5d38e079eb8c8d2db17a158276648548e19cd8f238cd3d1b0683cb223b4b159c6858df9866
z1449aab6422d01a703e6811273897e945c0a0bfe853f3e1ac25ecabe151ac282d9fc28b05cc203
z028a436940da97c9c3fb64c6d93c09c03678ab3c790b721e9beed250ee87723465fd8a9400d761
z519e4fc18208fc6b56a8aaa03da2436557a67dbcc034fcdad5ec992046b648baae3cb293f5a206
z54ebbd360e1772c9a90f445be00b4d0bc8098cc5a4f3eb7ac27adda30976b0fc98a0930703a2cf
zeca9f5447cc4f09c6db097107784da424e783b0c92693426c1875f852b6993d673f42999cc0060
zc523e8ecd1d618a19487752267bdce1e91599f283509fef96cafa992df7f3245e81dd7edfc8101
z744566cce28ab0bd62b29868c3806131296dbe7a77dcc2cf7ef39cb1deec6b8d51961a79554716
z189604bf76f4700bdcd47bf99dbd78de6308e5065263429b419f66fe590717fc226b6fb56dc31f
z1166bd229681412231009b31e2279b37fa632178b79fec2f6039a048490bbaac925ab209fffb17
z45b823d09c5062d1069e0a4d503262b7ce51153eb45daa2de12b170050fb0d31ff8e00c6b14ac5
z594126c0430a005cc7bbc8d8c633913b5bf46b0c5fbf4b5bd0764fdf11b3a202d11eabc17d7066
ze53c0e41a833ce4499e52824131a2a44ec0e071aab35b86fd408c8d1530ea965083d86a7e31b33
z13a945fd9a55cf38bccda61c883a8bd2ece129412a0b2296bbb90c5d03dbd8aac444c5fc7fe582
z003ebd594aa29a715353ef43d1d730522a77c798ce4486a6320634712c7ea2211e4a9dec1d9cf9
z105e332cc65787ec867c7dbb50adb1b34ab0f126bbcf945dd1284ad59c54e60275d76374513a9a
zc35bfa4c13b6138b6453acdba78b9231fa0fa644d186ebcac1a24abb1dec865fd0f5394411c5c1
z98f591f9103d332c3bcacc35e5282066896eab852f14e48b2d6f63d51d93fbfdd286489ca502dd
zf0ba4a95a7f7f58404bd3c9b8b661343695971c1fc0b09ff96711c9ee6e738c690ac7eb92f97f0
z809bfd421439a22ab06f7ec5c641c5ac7908b863fc4fd3eabee1fbedd68531bb87256a9b70409e
z3b47a5ed620b1dd528e01d2234784549d91d59fa1231eb7324fc286ddbb60d3f5be43f64b38217
zd85c18e0bf79c68c6eb782a63b0601f5674df219c382e6b752c3bc996e49aa7f57f7801f0248cf
z52902c087ca50e6fded2a60d99de3ec21c68ecdb966b5ed892ad6e5705bfd9b039728dbf5cf070
zfde87fee411b925bfb84c8446354398e8de595048232243db09e97ffd2282bf7b07919d668104f
z57f119d9668aa42d4d6caa1a533c541ae172627fbc5024a1491c1dd40f2b07bec43aab9962f99d
z1fa45910097f67ebbe48dcb6df43b94d29a63ee7157a5e292c0c075d9be333d20d524ed8ab99a7
zbbda0c80f99d27e7dd6f1efbdf98f310256266492eb97af5a3c05b3407fb07d6f1c54733e48f4c
za26ebac6aefad3f6a9f7a619bc0eb9ef243f571c0f176177853ebaec41a09d965a36952cbfdb3d
z9387f11699e39255bd3fcf56126967433cfa599505c6bd59a082afbbaa20ee045d73b611649e2b
z8a91795af0dc2ea36936de530d3f50df4f545477d23369c6833823254c27fa8512b8db05939a80
z705e16955ae8ec907df8eff401e65c0e925c55dc8223aaae9355fb1a01fb3eb430393f7568703c
zff36597a7aed789ef67b2b685eece71f1f08af75e080af7f06e9cc6eef1cdf87ff790015fac51b
z1cce833471f164b10aa658185b935bb80c91183d16b85d0929cd70a7729d1aca04caf2835ebd58
ze8b362651989eca049eef31cb9002b5067b5644b6845949a78c88809289c1f8f5b857c12017fd2
zb143da7886100746942f98a2a7617b998cfe6f754933b288882226d47d3df5b8342161c395ab28
z7df22a4d1b572f389ddef4dc08dce3d82a2d72185346814beaa0f93a46faf91a7d6366d766a4b4
za6274ecbbb91d8e3973ebc32a2ead4d791e0d1d5e858e006c194565fee61c0c26d67112a8d59a3
z5431ffffd288d26b69525e578da4646c96f0dd6ed005158abaef5fd31ef3ee2f1665952eaacb82
z4b465254d0d254edcbea05d014df438e445066962ca03a64fb4cad1232eb45329a2adb8e07075f
z6e270deba470c806d38713ec19dcffba6cf792d0c94314d92ed2d13a7733ffd72e033fe023f094
zc20031a87fa140c9c793948a8b54062eee521f0baaf92023698e1de9560d40059c87978ddbffef
zeeb250c039450a3ab0abbc098ca37b4f24985cbb3b0f34a7bbcc9bdf09f86c6d8ea6df34fb03e2
z782877438b82b8b3a5c79514f0a04d0a9a530d55b48d4f3b6553e7e78af062f95288c2abf030cf
z29bd91a29067244b142e7c7c9f0f7b204bde81715ce56d174888845703e170884976b0603cdfd1
z8f0fbaeb0676b2a4d2e6f386d416363b20d0a944301c075fbcbe67d8ff74505a18af421f3bd6a7
z42c85a92a26191634f30e4638a2e0ee4034e98f8dc2dd0ea69b188147630a2b68cf8153899ca3a
z7ec98d0fccac5721461ba53b722b6d8df6c91ed4ba7ad47bdc043aaa297b1afc1e7781fbc5d550
za75ceecd74f39cadd9f6307bdece39218864e8e344dde3a8eca8f4b747277c66d291f1697b628b
zac25b65d2840fb59c3140017d7b20f5190d50bb769734415ff68302d844e0e6ae6678922dcd077
z6df4d9370cf0f0c43490a93cf865fab4817fd2901e179a6ad8d58368c3c7dc4fd010b9bf23f859
zf095643e6c00ae7edb55ebffd69fd1cd04ff1fdf829384864fc90988fab7e350c29b1abe49f089
z26f5b449c064686628510032f68a3d5e920082aec2696421ba89f7b0a5eedec5e51ef45cdd3822
z4c0b28e212c197f7a9c081ee4147c94fcfa4054b71d955a61f1c4be2ead8b4c7bae7b2983c0d11
zf65b931bba15cef91b48601f96c6fa1b089a9174a455a6170bda8676402ec9b8435f934dbe932a
za29ec2401d162ccfc5980b88bf1945123d50874e6ec5a5a1f59f632f9f0e34080422e2bcd13c5f
z80bb138e6d712bbfd41294c0a446686b65fd128fb09293558c95d9a109e573c49c6084499ef9ec
za68cd6986a5decd9e51475953511644cf40913a4b1e6c94b03c39015a77b2c31cfa5ed79ab3361
z9c53dc36018ea3600f5162d72f23a68da73d3491b498ae17c2bd1ae8fb4ba3123f193555524cb7
zf79ba528453d0a5a026e9b8c1500fe7016640b5bfaafe0042ade2f668ec3206676c158ad6c166e
z10fd6406c0916e228400df4a4d5b936a1cc29921944041909673fc651f5f4c833453280dbf3963
z59ceed8df4a0175cc7dfdbbcb725daa32444377a0c0c62574d1521fe083c23e60729a09529f429
z874de8103e4542b18866ecff57327efed8ef38fc627619d7bdeec8b35d7bf34c1a3956d86f951b
z60b0370d9a64334b6f482ea5535866bc473f8957c2f35c05f90606542325e1efaa3fdca5894bbf
z1366224b074c2c8a19b79bd65e1b147178b708772b93ec523b67f1d1fdfe0a10483db08b1c3e4e
z7308121c0e565ff6a60e33819662d6ff08861f0462e2b3ab8f7abe89da627f3b51aa72783d0a08
zd9fbd506e7d3aaad64c9085927a1a09468d670d5d700577acab9b5368c40ee85ffb3802a86c193
zaa7c1cc220feb3f2a526bb1f2207234c3f34ddfc611b2d9c42c44ffb8ca34174fc16b7a16930e2
z93f6a1a31de4014439bee176bf09f26fabbacf720d5801ba38a5e42402338a8a4e6bf84eb8f2fd
zd50c300010fd9ddf00fed199cc5b9928b8117e54e90a41c646e7d4087075d6b5b218656eae18ef
z92b20858c82510ed563aeacfb5346a646c82501763d5981bc9e7d60567c3aa362dedde13562671
z4540d0243e0cdbd98af2f7e4ff19e307698091c09ab9e84216e042e25998c027022da62def7e39
z3025b53da2d588a030b30f10a59687ec89a090064dbd08d8b94f21527179f6a54b816e0ddd01e8
ze022191a735ab387890936116967b218a225d0f1ce2bd0e7412b424ab471159ed2e3339b7e07d5
za58a2fb64f23ee516135b2c0cbbd39f0ea18c136e8dd1b47f2e8f5e6b485bf511b975b55169d4b
z01712d2c66e30b96cf4e5c8ec0fdf46c12d1d0aec9191f457c1162f4f2fa9ab41cab686035e343
zcedca015c3ab6544cd53ff51ac588fe2444f69a6614bfc61b009cf9eda8d0000f9704d33fc506f
z6fb221d74e237ceccff9a80a22d0f593d7985f53a322a5253dd691734cc79b0f577eab38deb771
z7054c1346caebf7736acd36cf5c2cdf3d95b84e18d8afc88041cac3f08ff7c893cdfa7d16bc97c
ze9ebc290f0b327beb3c3803de1e3b992922f7e42bc952655b8b40dfee871ba5b47c7e893c918a9
z1d9ea47597d140c8feac835e4d3350eb27d48610e00980d3a7fc62774c6aa0f500e8a7502fb30f
z0eda88df3eb4d0711c7a7277768a115751339a44c548b999f6627a03d30e3a63047f71fc613655
zce3cbbd3e15136e4a21b133a92c756a959bf296bfa264ec444223f0737e712dfe83316790673b6
z0cda861fe52a714b0981270c1605806e64234642a38c54eb6ec4faba0a60696d6b537c305cc657
z929f014acb687ab558f812298232f44e5ccf7b1b1adcccd96d973b88fb52f749c1648689be6656
zcc9fa08c81ae615d008b55f0e34e452e4b0770dc48f712595bfd123961e6c9c5b6a8336d04aa48
z785ae8a1eb1e892982e777b13a86871a19cb9147d91e4f10792b906dfd056337024b858275d256
z77dbf48b73874a369aa6c09178f9c511fecfa292433b9a4bd530f973584e33e15d9816b5cdbb1b
zaa388fc8e5dbe749b5e73fa4d3359cc5cb9a4949ff77fde13a7b8a764812d8ecba720cb88a42da
z29cc277f5e81d5669d7220683f377909424a1eb990d8cbe2ae4c98557413883eac8654fbd788ef
z27faf15364362c363667e04087b3b58e1ea4d0f1a19a325e25cc05487bf026bbdbf6fb0a08cd5c
z9aba428c37e8b8171ae010cd7d16f4378a8a3b4313cf5869347b20bd2afc9ce5687a949024f605
z3459e6d76e109570f39fdf48177da60cb6c00a2c9b31d3ed23ff49a41b298a2c9b84c79adc39fa
z0fea71ab052559f5559cb5de2e34eb975482faef30f01c8fd489e351a7ee3b22908dbd7fbb4f1c
zf579cc3e395fdf4b59c98d679682c78e6a47a04febdae45402add5a86011f85f077045f4727cda
z4d292094522adb962d3bf51d808e0df71fa632191b961e8e7688c369eaaf9adf4b2b66b0e54011
zf3652665e737caade45baef6a5a13117c28fd9fa86dbd1407d036433ad423b5c7582dbc38d32c3
zf85a6c6efd86a09d2c60dc6df26b92c511e80e2b318bfa18a50eea3c2f84cff98c766e891aa249
z0e802dd0852ba03d3bfaeed30f7dbe10fe1e78d4064cb589178c5706669197cb36a65135dc84c1
z65196aa802111ec37ab0e2d886f1151ef1748ceaf72b31cd84761f3a0842b97308562e5882e188
z85c96af0299a76e8b349bba6dfe1ebe29c8eec357a4107cd5139ca1c4d37e33fd463ec0be2fbb3
zf146018b57dcb4a4f1e5dc87b12906cb14960362ebba984c0c65fd432288f37524711e6e9108cb
z917f3ea42f21baf7441299a8fa10ac61ae166070a04ec5d916678c0c7ad21152a4cf1ce19bb019
z071e8ddf3eff9ef4459156d774983649b21798c9dc8f149898441f6d9c355a9097dfbe72b846c3
z4dbae14df1271983ad558ac745662fec888b169b673bd11f1b9bd6718a040d24d118ca5c4ac4ab
z4ffd0964c90918da9558502126fdebdbfc46f7efb4c36ceddfb07801c4663399b0d27573f51e60
z6b7493f8ed495f8120e13e87d5a1bad583fb3ea6dc6985e3ba1248471455eee38f82939a9b0bfb
zcf1760c6e9765e26bc5a8d01b6a5d5c421e52fd8f18e313df7db4f1b9babd385a0f0a898cefdd3
z284ee94d66f953cd8d34d5e442188d456c92906790aeeb6896c109fa8edbc686938538d1f6cc60
z321bda609220e52d8b41e3a610f495b3d189f50bf54e25aa49d5802774bff550c39b787f5d9f1e
z3508ffe7d7a324da1f58bde839418f539b21c064879e889e5eb477c1b3855cbebecb84865908b7
z96d248590d01d5dbbbf6547d46a5f163446d5d74dcc66ee6ead517c742f4f1c1912d56c1b8d508
zc0b698c3c0d8b25f66241c4ab8c7aff6e13f419b3663912162be699f7ead26e46ea4470b9ff11e
z95bc56351424252593db2676b74b6bcb28a2eeb403c88062aa890684766f4cd6e5e6adc629a86e
z5a519f135486cdd86e1486e8f5f42dd30ace63afab1b3d94a004afd82ea563ef8835fa9cbb06b2
zef60b9fb47cc93e3bf2578556a85c3cb0bb3e6ef78c133b665ca48a261b8d3c769a6177bf0ff33
zaba5d75248ecc6780178291098971de24c901401c9f7cdc563e0b763f0a9dbffd8f53257441f37
zcbe20d19a67fb6927b6e533d783926ddcd5700dc55fe134d25c2a043170e776c9224ae03d7cbfa
zd7edf4f124873452dfcf2ca5258b6ee4bddb070a6f9e8cda8268c17da18720cac4be6d275e724e
z32b1f2fa22e984ff1a00fce20972a1a9f4bfec3efa197b4051250cac62b723f8dad270c1303bdf
z61a9d67ef77be5cafc50cd0412c4a37e5ab3d461d62a92ffb653f5bbd41cbc670dfa7c1f0b0971
zc86b8af14e8aaa233f834d99339b40d49abd0631d6f1b5dfbdbf7592c4475bb6da2c9448fcddea
za7036af4f6174fcb0b0a0b442b2d650a9e1be111246c02cb01db689b5778f408a46d6fd15f4d29
z3bbb0e76fee4ab1cd1d8725ba3bc2b25b0c80df7455e543763eecd42e50f616ba9011ebc0cb625
z94ee157b8defa9b70581fca2dc23f91b659df8e5ba9932776618d0b1e3dafbf45db06d0df2778a
zed8ffc10d7ad927700b66da651aaeec9095f82f5f0534f8cb0a6f747a7c07eab7347a12806a483
zf2772437e86e4f61bb001b02380b8d9a2712c279caab0e15c29421ffaacd9ec333502dda521357
z81239114626b9ea41e7d0fce6dfb43af27d467b78cd346c936d14f8d9cddfb78504cae24914c3e
z0b69a25c3d42a907a39750b55ff0f53b298acc50bba14a3b01bbd9dd70ed1ec5b1f165c8f014ce
z033edc3ea6c283cb5f00f6ef7f0e2c97e2fbea4828ede3d65bafa6d54e0a5b728ddd0a4fd93350
zd381009ec68d81def87aa9710b05bf52ac4a1892ea969ee696beb9951956d4ab9e81f87a1a2f04
zb53b66390923037e1a7be8bb74132d94b82978f821a8d736f2d9c75d5d2f0ff4fa1b0c3b22b87e
zc9d1894125694c1b4af5d8da805bbbf42515c7f3454866f046ccd82cb08bdce0740bd5263e9817
z2947f5dbccc1cf76baaaf815058e596c4bbe0644ba8efa4999816fe23ad04461139367633f9746
z04e6c989dad4f8823583805af40f9eaf70e7a65209965dbf4a46d434e0255c963b103ddbc3e320
zd56e290ce3477a1138c911b1ba90a1e0390bc8a331b5a8e575b84a205d2f0adf36bb8c17a09d82
z8ebfe385ff91efa69049b8572fd1ade7d2cebc514fbd72514a20df8c368b1ef2806ac58f7823b3
z4c40872def771bc7695a5fd295e5e2007df9b0d9363bdade1c0d8c834eafd9b318a63bbe452cbf
z42a43968371714f24b87eb30fffb50e834fdedc85f5ad48ac66bdce34c40bed0134136f0aa26f2
z8543e4e6d175a50ece1722225e87e99b24af2db8f7e2186877c8283ba01c6ab546a8cc402d67b0
z4d1e14bc348545eac585f36f7db64931e7b1d656294b66f88be72f25d8026dc33c4e4f42ca907f
z92befceee7c82eee0217266fc2227223b294e583ce481c47841231fc28b8420cbf9e12bd69d0b9
z4c62fe9b6f669a64c2011e33a36c025c21fcc8ae883a8d1291dddc6e5110498d233f2ac904c9ba
z220b7352bc820ea9dbf416575dd9d9da732bd828229a676e9482843c6546fed1990b145e30daf6
zf8b2ecc67a8eca37c9c991e6ae6bdfaec808f858a61fe0e24853cabaaa8a70713b919cdefbcff1
zc9ca0b91d0a3f0d89d42c824d8666ed2fb528debe96a02ee3ade45f38a52b5b11571fcc607a6d1
z63498f13ae229faaa49827ea78ab4b258616472c780c0205961a1a91500fb6efc8c1b01ce401c2
z5837e9ef0f0a7aaadc911e2ab801d782f861cc68543be4d7fb343af04b4debf8bc66afad63f998
z81beb9cd1f357b36e8033a44b4c925584239b19c55dfbc15135332345850f955a1e17c86d31f4d
za8684e6927aeee9c129186828c860ca6095afe98bcc49d6eb7ddfd20ae6a62865c291956448ef1
zafbb09ffc1db8fbf9f58060d4819038804983f65f01587020b03964e6d3cd1915dacb4fde0c5df
z69d424a807969d11df0c55cb15b11fd0c4c9dde01d395b2c47b52d66733c800e60dedce541eea7
z0101093e7f013821b2d34e967892dcd1fcd797dd4eeac8585347f7861aa0abc0ae4c6f573f4e34
z923c54674a5a4bb2867e6993806b68f7eb7990dc163a6149ca993b3f56c6e6b55a46ab0e04be56
za5af1f53a69382d8b474ce7fdb37ea5d33404a88a1fab1164a67899ed8970f155233eb7b56682c
z27c22ea7ff2665e259922742d5d6ac6ef2935f9461922ee7730c3e19448b52bad988384d995774
zeeefeeece983dd840c3593572587d0198a6ec8a7a59db6c9392a4c93fd5e9d81d13872b9588558
z483964bae434b64547a7da1fa1c08b70e9e763551d82e9f562d790a0b3beb1d62bf05286460d81
z1319e27c0e4418dd2b89dc397b0428677c18d0719893531f96da5935d5644b4a8febbefbe3e0ef
z50fcef4afe7c97a758d32c7c594c13f4c2195392a3e7acbc2d6499129d16efe3bd598ec45405ea
z7488390ae5386f86ac7ab338b75ad0f29eaaee935b08cf804b071b1addf626bbacd3d0866029de
zb5c2ada9c673eec3ff647229dda2db0ba8fb95b6b9233c10e5b916c951555f34b16643382112a6
z11ac159479c295c8b2202ae4e4796d3e053354e546ea790629e54a0b4ec243f8f881777bf38e6b
z589a27ada5134162597c46ee9cb5264d9d9d626bf39a6e9127186a081fcf2e28f620a5a81753f8
z9dcaedd7e9b82841e918adfb78fbd45be76b5c97b7a048f6a779f523fc6698cf50663af52fc5f3
z7632b4a6c47cdfdad1ddab056b6fee1f73849a74fdfc1d66668998ef4868880a1c0676f90640e9
z07149212ac90a062d87843c4ac8916cce087f9811704a5246cdd8f04b7924f985ed0088c117466
z92b0c93039ccfb5d55b1a801242cb7017012cc7292bacef2c17296d0116641a4f474933acca58b
z949fe26f65cdebc680b39acd93781b8e2e00716a81eaabf1401b18c7ef40dd40f906db6129326c
zb7503da674073b9e003214e5a97d9fadcc2a06dcda452c7d58bdbf9dcc0f952afd6464b944952c
zaaab80f365c10e99e21df865f457a1ee071969d056e8c2a916a5255f25438264ad2f66448470e9
zbc8d8ccaf141fc917c6b37c13e917dad9054cf542b6ab018534b4ff3719a793d490c35cf975acb
z15bac4826938f97d7510d6795837d9eebc4877d0b0b744f9470e3d392c58b4ebd1a240d07a66f7
zfcb9a024668eb56ead9d3e6f59823c155a930ee4bc6caf61074a46dea8ac813aa1093bf7ce9b6b
z59f0b4998210d083419f0c6adee5838376959161fea26ee7afa5bf21f8c4c31c23bb70b820dfae
z9e6dd0dbe7c1f6977e9eacd12906a7d703d56ac70ce12fca9d86368662876a638efb91bdedd104
z10ec2031bc62e15bc01d36fbf163f438b45b9a7b4b54d520f582c186f04d26c854dbcf6e36ed0e
z1df2597bd2fc9b0606d37acf77fc6d946faf79faa41932cb1262976430d64fc7adeab676ab3e60
z6f432644397b524617e34db3389a2f279ce6b2c60f0591638591f5225fcbbde7f946df1a33043a
z862a8e4f1daba96e51bf3299d0179dd3e1d5753df72eff7c9ee0792caa1a2942fda2df351cc034
z209ef3b115a20d47129f522f65b1d1279ed75979d0aa51f206fe3d66cd0ec40a6c4537b1d7f49e
zb508f4687da985e66ec4b9062a6a43b15fcd4000feaee9095af5ee772a82d05e271d425cc78f7d
z1e709933a1c23bafcd6251de3e4d26e3de3eb74b1e7564a0d65ea6c4bea741a835c1a7d2ff5f8e
z3c4069f06389f259745dfec698cd9cef56c0caee6304d8a7c5f70c96cf9d72fe7ddb5335e245e1
z9bc0a05712322dc3f3e1710b331592ba75ffccc4db95eb168c8c2e35af222249d5c53bbb3a458c
ze895765cbe478e705dd9847a4f77cbf45108f3d87a3f67b5b4e43f1cd9dac4bc00ef62ef127462
ze61a7eb7b48895d56aeb0ccbbf9ed359c986015aa082815a2b08b67fd8da2abda09c4985ea57cf
z381e59d32554fb456a19fc1870d24064383650ba2006643ec3a22fa08e4864bf1d8d9c9d9ab54f
za9cb296b9b954d9f762edf79b9fce1bac24d54f777328d2ec254c9bec954361036125de2ad4255
zfdbcca755361a15ecfb00c58501f893ad915fd29627ac7d6620e8da359cba6402a3ec20773d140
za175a9fcff2ffd4b135c34bd4a057754abb8e6cd667544140379f0c8d47b5e391cede9e2842a00
zb6690eba386fe93417f2c03b29649f18b10dddfe03383eceafdc6c9706dd0f978bbc6bf5f38e45
zb38f76d67fca845f797ebf5e1be14d92bfcfe07ccc0c0cf50065bf3686d790c7393392a836c1f7
z3fdddaa34bf37e3e726f904749be8a0ab148db250e63a860cd97ce4000aa1d6a84fa53e332d1a1
zc0550fc4d0ecb886d2f3a3780a0999e511cb9ce36ea07fc3488ca7a7d4d51517aa8573f7c0c375
z5bada631cebdfe928b99b5d5165b45bbb2206fece19063890e5273a17949a5e46639d767395ddc
z91bf93d669c5f098ef5c029e07999eefa1a0893a9a29ea21a31812b87b84790d6047fbce58b768
z0db08b34b6b63285d55c25462a942dbc4d61dc4b7ecc1267636215487ff92fba75efe5ec9449e1
z86275cf7cb29510fb736b92ebec012fa8be7f637db8a1ed6994b53cb0fbc13b00b0f2ba49a8cc7
z65313904ed2aeb87f336d2e9d341108da83390126eac14558ab7c93a170a13b1aba019e3e6dffc
z5226e522543b84ea1faed46126356c275e0c2f583f666a0657e0b6f3e6008c39a8c58908296c12
zad99a8cdca612ad13efa9103f1822aa3f360e0276dc93e7b26e04734bea4d830a0843f68251f34
zdb453403de41c085b747cee035497119320b281c1046bb0cd0eb0ce626751bb1ac610c9f14c5a6
z1274a2eccdf13e38ff7ab07086d1dbca8b916f81e083b3fe1d369389972988ece04ef79e22efca
z4610e69db9ae5621d5984f094ca901397b59bd4a6eca87ad61376f04bb3a7884fbf315e3622b45
ze75fca84d9f92515eb4032c5b90dc319dba191f5b2c667827d34335b0b5f6777db63a7858d724e
zd6a2068f0d85ac5358e2b6b42bfa11d2a8f0ab0c0914d87a03fc250289f06a261a9f95a97f2e5a
zb941e135a2bda6622e2d7dfb19f7873e140d9dcfd539b66fc72a794595e400c2c47c2fe02d2133
z8093ac5590fa6bfa66c5e8435d755cceb508ebc65d3d542e7ba7b78e8e3c0ad7ba482cf3016fa4
z90ec524e57c2990236b867690d8483c9d927f1c96e2d06b9ebf050734287f2382ddb70291c82bf
zd7ac43c447740f4bee344fce7b8c49928afb66f7afeeda8aa66e926a6817163a12e91afb7cb26d
zf148d74aee84d44b1859ba16c524eee2d29235fffadba3e51ac4a34c9816cf973855c7332f2126
za2ab14bbf1494786b3ebb0b993757838387b6dd778855be9926c97ed36716beda91d0160cd3650
z88f8870386119d2b5b40eabd8b50ef88ee06363a64045710e7578cadc2c3305e6318699f043eb6
z790916365ae7de9bd1a20d45b10a4987802941da977971239d7f7a8686e51c7e4c00860df167d4
z36c5b8a5d5f14b05495f42c49fa2f5bbe9112e6c7ea62096c614c8f36f36326d995f626c7e29e5
zb73a5402db9aaa46f95e41288dd94e45f4bf9e8814f8602e4f746a76843e36185c1fcda90d2204
z9195d6e2dcc082baf079032ddb34cb5bbbb8441a4d134cf985f0602610102d36545bf9aa2c7a3a
z84edb79f856cfa0edb99042202d49444d3e7362e2484c83dbc05033b18c5c9f0f3075cd170e9c5
zee2fb37f2a4d8d680ec3004025a62548f6a7ae1fb0591a31e53148f27b7efd7f1ee6d1f872fbca
z20e9418e8df1470b8e8b9ba3ac580e12ae1696c9c393ff56550eafe4e68c2cb12bf5076205959f
zbad031e399388c26c7f7f9e79b14d63edbae88b6372f80e7b6b6083970545c00ec8d9779a84e98
z6ad9be2c563bead2bafeea3fa409ddf0a8890a381c268dfd2ceecbe7a2d0a99510965a4461a8fb
z29f62adc65f7ebb8de2309a8c0390b787dea5fb1ce6c11b9e1f203ca87a6eb9b37384576682eae
zf2b74c04e906c91e95845750be1678c1b28e370459a56e9990b5bc7396176e1804b4a2c97dfacf
z44f9745a3bd0b03b147f665563272461969d75f94a2b9287465f7d66ce210b5301023ea8c58db1
z5ba547cbdd29f4ae1a118296d54c2382844b310549be7da2451d42543ca9a4b3b53cee847eb7a6
z018ff7d96088a56f3878d3ed4d6941dad64eb660ea1969f4b78fb1da160983fb543e4478fc7e04
z4cded418e505b864e4c3a8e175957636d92c2a6b25174efa89152806be4ec3a224b9caf4cfe07c
zc4358684eac639bfe29eace2753aee6b18ecf962bf7a86dea197d1d53546bc9c00770a4b7d0929
z84918368b704d0d02cc9f0650bf07d7a6f070f842190f7798a2773c6f6f9a0249517ac97c8cfbf
z97cade3323222bff811cb0765416d2b0753dc0f9ffdc037a190332d28e5e6e77774279aede41c4
z4d9d1d8c7b10609222b858d9c561a14188e6217dbd12c3607b6484517d15a52d6499e731f2fe73
zaf68fa02b3bf355bac373501d371f08c88836af3c22869c91b74f37674f333102aaa23545ec76a
zeaa426d326c633e44c85418f8f4718cab8265344bd019ab9bf8746351dde5ee6f181a6f9c07b40
zc9370f5d3f6b027046b150231c9c4571b85e15c5f3c0cf26acb054dfb88766cfee3864ec750ecb
zefa4863c972c7c47f61410d15f8f63ba12eee75805d3654f4bebe028c3b8b551480e18269d95e7
z0e420109013b52b73a48fd7ee591fc09ee00f30692ed2ce3ad9787e5d208ae80709766d78f012e
zc5926bd0863dbdcd4b30e3cb4a1ac927d8faf436896ee6cb6c0f20c9daa9df7d004a3d2da03362
z4167922d2df25012aabbf5069775bf2e80baa82313e0bdd25e8920bae05fa3f18c03fc93418ab3
z01a0e58e976845c18db88aef60f0c66591b0f92f1bdbcca7a0a1f2fe9e2f0d9adf99190fa416b9
z43b1d1a522e2e70276a00ff2ca83466b757df4c9d4a4c11558c239d8ca00c7ae76d2f6776dc4af
zf83b977b34d2690995bbd8074cd588debc1773559ce2396d247bd2d991eb6807536f93f27db8b1
z52f95175467f54c4e41d26185ee359f97d69e9ca4f189d809d0a5cae9b6db7f40f145d49ba0dc4
z5a667ab2a2165d5b0ab5b3ed5fd9f1fdf28ec592ac7c3f6cc6e34850e2df45255b08edc158915e
zb3c2c5760d7858feb0571d932d39ef00ce03ff0d45bb3272b19219257aacfce5d748ebf56a25a7
z0e7a5b74f9fc774af6447e718ebe2a0f5acff45db2acbdfb3df0222240ac1037c4031eabf9ee37
ze643163102fcf49841bf5af12b9022a24237ea45b7687d6dabeb80a98e57f6c07b6d3b5a48807b
z10bf94e1ed6c108bbd9cdb6f8f350cb8b790453b831137a8343c52d025bea633700ad2f911d5f8
z78809cea3d8c9b1e6c897b07292e89dba3d687df54b6df18d46b6e36edb04e4bdd793faf03608c
zec187eb2348e649bbace45505cec48f8d54933c647817b01d2bfbc161054d1f3639ca2b474fc5b
zcf34f0c43fe6c7286c35b4becb47191df8fb237a01f8be4fbf02d4ab2eb9fe343abe62666c9301
ze0ebfd94475d12112282d8dd09ce4a62e14a618d56c9f98bb4c936b1b1380a7d637976112c7211
z9a84de0ed92dc271dcc48327bb911d79d72e14aa01cfda600a84e77404de49ca833718992be7a7
z6d8a2b276945eea8efb0ce2ca09c62b1c0c0e6c6455489135c7d57b0fe52ccd0240cdf9c6d12f9
z130c44bfd9b51b5932b938cb3a2af0db54f38c1483d5e27cbcadcd08b7a5ea4d311f9065ad0831
z4f6e75e5839f4fc21a1d5098f8747aa602467e0e9cae353ee42b443bb5d0307671536e3e717e21
ze2ccd99b64a0ba922795a16c6749fa96d8881c6a9d5e4aa478fc42671180a3c90087d3f7927cc5
z0dffab85dc9870c7148c21c29628adc082d0e39ac159af2756620880c2d63a43e37e2611b1de63
zf484f1db97ca313681eacbf322703a4a24737bb0245af61ae8aa4623842ed78f933566a1f8c1c8
z6728f44d35fd5f79ad3aec6176e0ab3786898a092deba154d38411ce795445328ef0d14a883e5a
ze376e64527fa429f5117ac3536a7190a736ae20c1aa6bbd7465aa6c22c811586e0e8c3349eb374
zf43ebadb75ee445afa6525a48d3568f9827358bf60649c024f713b4db1bcd802cfeaf2b4d2b23a
z84531c466f7c3fe5682c4b10a3c1631cf24a479c9c283e5792754f43a2a108f50e16ee4eb1796e
z4bf9e5cc1d13f9d1c5eb97b92d479613accf0f0f049ab857cb2ca1a9f039223e1e90a378a8f2af
z09d38aa017f582fed08b84ca6d2fc61e092d800bd69c32fec0fc495175664f97269905ac774c25
z17066aa1405b62d7b19f869d6636bb2010b2c4a734e2cf28f6690f8223ac7d6b5901ff8bb49376
z193694176171ebdacb31500ed0b67e7cea9cff4241b8840adb7cb057378876b3a8c24cdd3bb027
z9191f6fec7465f610ffcaaedd4050cb7a53729ba03a71008f936cbc3bd269731815ca2bf527c60
z82a60b5d266ece8b27962c9c6235069b7af09f67d54dd03284cfe1ce85398b545c34944e8304c5
z54c7ac59c5ae71b22f7e88814bc24ecc0b73818d03bc038d8a5302db334f34d95b87ebba584c0a
z7a744ca269e0d491d6247db9326a026376084a1721f24e703c311093872a92be0f7e9a4679f7f7
z0a34bd16cd3c680ba30744059740998e367a359f5843e62475a3731d9d6a7b9061cfc6b05284d2
z6755fcd846db367d9fba5855b14e2095a5eb74f62aa2938f288b0a331a89b19a1fffe1ef8ab761
z1457fbdf2498b2ce0361a82d6c1deb91f900d9de5c35404e665f98a27ec5b8c1679da415f8fdfd
z921cfda2f25066c57c3dbb307c7b3d459e79aa19f87205605f34acf3ba676b1979f9e88c764f07
z63e1b593840701f68812aea18f75b6a0c4400322373a2d341dac94c0903029d6651b26ca1e881b
z4e1570231aa269fcdb0939aad8ec521de6585d7020a95fede5cf15b34b1caca525ae2093c8b286
z66f4871896a4018d1ae0c52b66ea7f90f24d0049d047b8e2a369f7c25fff89da0b093aa273752a
z8f8df3393818dc168ea296b0122e70a9a66d1fd3734b7b55cfedee1904e309f8c0ccca3876970a
z096bccfbcce319043fa8831d972681c434fa00fd354f40209c8b092264f35ef3a17596ea9ca898
zcbd285c3f5b95e4a6c4213696721ea53f025fd4ca41c8f2be70d30976ab3b32cce21ce11b73713
z49d19f81d9bb517acc85a522cc8383127246ce8e9b5eec171892779abcb25938efd41061f80416
zf87942883cd382fe20a484393e6c97a04a078331adad8d21b1a10f77a56315bd2167b0485307e7
z8fcc955205f062825d0accef1f20e389bbcd5ad50026ac6fa9504b7dd93756b98db822129beb24
z8cca6e3f4ee80e772ac3ca40bc90f043024fc3de1f99df39a01a67045a74e2ca9d8c2e1c21d343
zf021d1a976568b590cd0298616432dbb8cbd5b3a871a8237404bfd693beb14550fcad45db18e4e
z3a40760d6fa177a1c59be992301cabde7971470227ef3399ce2b945a5da93f7eeb099db73b6b7f
z344ea40c6bb7bca1214705dbc73112d788a989c3a119f5d5aa932d33f421b652ee49bf8f41574b
z7edbde0acabe1a90ffbcfcc77f56278c52c7383b0f480807aec353890b817072015916ad913fa6
zcd427c57545430c75fbeacd8cfc6bfaf5f67022b226ed7e2c4455679eecb16db79e54fc6bc0b46
z9306761fb623d22a879ea186ec273acb93303e8bf6040aaa4b7b1742bbb36bd4819a7f13c9b3cd
z15799cac7381d4c21e04ba4bd5a3b6ccb3203178dfeb9c3c81620e36827ecd4b8c49991d4b519e
zc7322fa1cc299dae00410f09cae5e4ccba9e28c4d6813b2922a0f7403d2460d0ff25056b73ed1f
z5e570072e563542720ce266304539313a15980174de458a61e45e00ec5656ecdc69807e0ebb4bd
z30898a86e36d84a30a8fc242b62b3745a4e645b97501b1058c3904dfecb7313843f3689e2e400b
ze0f085196b960639f8382c86a79c61dafb8e18e5076ce6660a97665cf3af3eb810b6473c807cfa
zf54c6aaea8fb7fd720942b5e02c0d59ecb5e0066428329bba633ffe739368265c7d664f4f7a49d
z6f632c720f3443dc7d02dec9a5b8f89edc49ccc76e6734bc669589fafbb61cfb731bc0aca66c80
za608fdbb493557cbac5fd86658de6d6f8205caf2983b2756bb90e2df025f5d4c9de3c366c03f88
za128ec2851924135681d86c23e69442eb188685c0d63f32c90cfdda746dc9f56c5804293ceb13f
z3506ac0ac9ecabc1fa7a941629d1cccfa48ed19d58e9446d8d68cbe24f95d95b59e37e626dea78
z8ae95624ad562dbe2733ffb11e4214627a45edee3f546e193cc8279d2f0027ce786b889ea40137
z92437656f08b81bfe4280e56f2eea27b94ce12a57d775f45439aee81a25727f0514378d43a7a1e
ze0908ab6b3f59636219142018422b88b6a7bf96bf21599d1221750ec25c3946257e77c3fca0e21
zb99a87b1b8d3ee993011431a49e0a594c64b32c37b429cf1bdab11517f6cbc95dc032751d60c11
z13a2e71b1de9fc689b334e7ba855d14864c048528026dcd5b75b5883c6d3e1d7616b8971a0f45e
zd7e25dbdc5b9f5f58ff04695c66c97453ffe7075c91f16dc768987b0642476533e63d7d6bf0605
z782f274e693ef9b685b8fcf5e962451a15dee37a86b8db3eadcfe6918e2e237d975eef1bbf3656
zb16a01f8e8abe55a8a30ec78f937fa52bb162b1b023e99dba0c1800191a30ed58bc83396f902d1
z6ba4e70379020876f861b22ba9def5791b903f618b09b7820ec09903307d6ee5b9c329f1bef25e
z8e092dfe3fc7052b369ba8dfc672ed4ef14fc9589a68fd9a5f0a86e535c299189dd2996cd217b1
z544fda3d4ba4ae418a6b8ecf11222f098237cb436784c39a6db34320daf0f2f2211ae118f25574
z02bc920a1a7c17ca3c59037fa625dec0bcc5eee25996269b6e4b1ce497f0b709ad90dfa9790a3d
z107b2386b87084948232b19bad75bc3939bc6a79a1f4cdb697bd93b579a47cc78e6e39f9ac1808
z3ef4b69cb7da3917c5005b5c45f95f3653ec263de684a73d49aa9f04251c0e5174c5038bcd243d
z2d0f98d84a8195b55db1f9f814089d970106b26a790c818aeeb40cfe36314765784e72f96f35ef
z6cdeae90a799b8410637302fbcc048a9d2f82d3a8e696ac1b7c517859c3bbbec2ca49968bbeb44
z0276af86b97eda5d9e72edf0763b0d0569fa8cc0a59ae5c0081032b4cab4d21eb6c2606cc6d0a2
zb05f3fb3116b974b8caf1a1d692f2d5ae3e888719772490757e32b54095598c7bbadb7147f2c8a
z9a9eaab5773141622f1a773ce1d11e2e7d206f591b62a08f234626f159244c73f0bb0b1b32ae8a
z42c24db5f00fdb49628f14b1749e972ce2f9ece4208b72dda67cef31185d55fcae0e980b55b361
z2e53dd25dc8c6d73c14827db17227b52f0ccaeab5a7b3148e36c04291c010adbbf0315637b7de5
z54a16407741cc07637d016ce03d19d76aea733b39fe77d520a3d64ea1decd9c55113510393717a
zfa8780eda6e20b084b7a10b598420a6c4420cd972f9cbc74d679fd4909b8478a924df53b67edea
z4baa640d7203d1c03cbf5a368fa6b9068e178f3636531cbd62e78a6687e41b013a183d55d62456
z75969f5fcfe087a578c6563f973d418f27053032e4da07be02edcf3777a47f0ad621da0feb5f28
zc92a04bd67992fc3ca99d456419c4ee89f062c9ba4d47ce386baacf7ce74221d55ee972a50f354
zad193ef61c539772acde0c7ea6b04f4874632b231a308e361400751e80a43619b639028fa0c85f
z9368562daf09da2a3a7515c56542d7c9d1d57ebbfff9c7e2f347336fd0e2de2c9a5c7b47349794
z38b9c0c202054a32f5958aa3c4242b2b36c4c69870bd7451b6d9f6d2bd27afe5a078adc43416e6
za32a88786af5854a32c1372d7e17cbf0ce6be381545cd615412e13b1b94ce46608e18f569c574a
z9b2bb8cf5cf41ff3658c3137b92038e5ca5428a7f6d56ada9dd871e215988a51034824acf0b67f
z10cb0b277a1597a5b4095e5ca51d744a56dbb0ce8abf5153fd0fe83aab9040b127913c1c42bec7
z327eba2385457ca71ddb9c4d57d149433606b3249689b3a11946ae5e0003e985db6eac3088f5fb
zbc1574205db6b275fcac314c46a6c672c510978cf7bfa27c4d0c3e2bfba759fecbeec4c08e7dba
zb82650e1d4f76bb98649f311fab2d58e02c72a28449d3c079475c2aed68d587a9f28a6843ba1aa
zeed600090452df42a7578a0949c6482d3f2a0abb4b6a0f4950c14c1c78650a176ca91bfb3b3e31
z605a8d6b724a41e88fc112fbf68514a7ba87dd2739b025e50fd25e9cc9c8bad5ef89b54bbd20a2
z4c0d51c399cdc7545df107dcc952fb4d73707183243ebdb94ddc979a06ff1a57e59d98714482a6
zb80951abb7cf84f8d5b1a6705df3789b98694b4a17bf2fd9ad4b68c1eadc83858db9cfd853b8c3
zd5c38855f8978e137609232e398cdd97f1c35a9e2126149d9ddaac78b1b8aa14924b5a44480c27
zdab6de514eaaef1a497acb102cad47a97d38c062cee83aa91fe194763f12c45ffa1a85a3b64a7f
z2bb8a974fd8e5ee77a6cd563dd24012676e894808b867404bf3b44c01b92530884f6700364263a
zcc33a54ce8fe267aab3a2000bf9b97af860ac6d835faceb788b14c7ebba7aaafd3cebcc39c7bb4
za75c0e42b00fcf3145ea3879dfccc5eccf655167b209b9635b815e79cd3fad3f3dd8fd495d2675
za71932013efe21ca51becea9416c305562cb9f034af274d567f143b1668283b3360bfcf53fd4ef
zd66b373da7ea61bfbd6b2d70421df5644095c4f3ee2069e0bed38ae3a209f783cd4b92ae1cd976
za4e4baf0d38f9e7a16866fdddddcec181df7190adb3dbda46fe5304fff8979e6adc7a6506855d6
z069d1ded5a9a73651f9668d1434e4e286fea6d6530c16f480e3360f57bf67e1d4675ec9a284d14
z04fc9534dfb049dbd2a5007fcc5c8548de87e9ef4f71f55f37a5d64fb8aca1db408084c5717852
z4625ebc6f8d27261f05cb53a2a79b97019fb4620ce22a1e1361aa124b8575102b66757d4df46c5
z7ed97aa4ae7d958228b3ed9225bd51f5a68e133910a414bc5372493bcc67434582919785ad4cfd
z6fc018a02b16fc290fdf38bb691f366bc67dbc0ab6d9ad1f201355827e8d8e0ffe9b391fb21849
za04e3458ae09339aed6e4f40e831f173aa17972564e819d442050087e22d02d863a92df792c165
z59aa3dd5b741a331fbb32b05acca654a86a811b2934e9cc37583d208b898e98fb0fcbbe34f7c81
z0c73d5bf161d2ef6301977b7314c9114407e84a20268d6bd83d448b325261d06b00a1fa7a6af0d
z4d79b17c48563e7e3c2759607007f436bc526fd9e5866557d6fd9d2e8cde3bc0fa006ca47211ed
z4efdb64348a0cfe1624512549d450502d0cfd3e950260d59c8b836635e97568c771633560e9073
z46a9d40af68ca124027237234de217408e9d5726cf149f80cbd53d208e299fc0d2786f09e46e81
zd34e4670dff06ee7d7f414bee39a98dc0e00055fbdb4a7377adfb20556b3b78f96aa0b409a5be9
zec8ba5305989eb74dab111a05897f4896b06351158b3db78aecc6b6a9eba1c5258d586bc96c39b
z3831735c365df3ac06fffe6bb336ec69b61eaaf9aa2d11282584fd874fd7ca9dc2cb25c38d037f
zaead2d4a973785e45ae08e1afcb29596a2511ba58432ff987f47dccad350398c02babe56ba8edc
z6918fad5e2bdb36533b38e894e0d39aad9ce9375310451356f0b7a8e83900097175b346eefc326
z1ee23ebf33dbb6ca564d2b42dd19db7e9d615631ea7f3bb50fe7b04ad545b1c7f6d173371ff1ca
z9648fb0642d4145edea8504739b9c6e8f3bc4dc92c7bf18ec6efa0c0014693c36b2c93b44a826a
ze6e03e599dbba3ccbbb3a3cfd1642df0aa2fa32189a602a181ea71d20181cceac67b559f04ff03
z10ed9f1b2bfc0b8947d3c46813325292d8bf847891f1a283f915f6bf68cbca53d4b004092ea720
z1f743257ce6c9568c7d7b229be063fecba7fccc07d02ae659e14e311111c31248c67ce86c321e5
z99bea0e1254e26cd3771f0158595df1b30ad1c28ec88e21d8484043f9461f11e6a9c35e4195e9a
z3e197391741ded6e8b3ff05d10157eda8a9bf689a8090f7caab1313c0a4f8a64d9d2af2e5adc46
zd4eb7937ff11e51c6321e7872735e9be53f1c864bd203daace94073e29b272a0166b38fb76c9e4
zb8257b6787aa367da9e4c75c19be0d9d8859493a125b45432b72460fdbca4392aad2396fd9d162
ze18e32623be9afdd453ffa8f3fd361654b6e38c884f4a7e79ed9302e12a5089b7fbdbd7e2ad660
z91e17bfc9cb0bd4ac0be9bbe635079e85cc87bc0cd9be839cffe3bb437a927bc2ddf1b298ca247
z5f551d8f503eb7ad399a53ce237cd300cfc0981f1c2726d90b8eac7a97bc11f1db0a0eba0aa65a
z3f84d3817a45768bac0af9e0a0d0352539b82d86ea9df3ff3b72eda23057848f5ef19facfb3ba3
z84555ee74dc663d8899a67d514bed3742e24ecc67674d51b06f1bff5ce6cde8b4506c5d98253f5
z735166168757a98954cfbc90ba4b28964035eaf15e9aaf9d237837e181b070535e72f54014068e
z7c07481d5adc4b63db4caa04bb36d4df36d5a32afaed598e8d321071ea35388036643040e6b7c1
z37d2fd365d7d3c7160c6405d1ac623d85b3cd7516cb23198859bca76310fc51b817d29203fe465
z1c7ff286d990d54d6338e871e65f488c2545f9bce6049601adf5769515b4db2566758a9bc3e9ac
z014b4935a10b6fcf4d6d5c96e000c17d92085ca4b9b636a75eab02fde76b256ec357380e984050
zdfe789683ca0d4265101e8ba331189db9481ac1e2167512b411e0a63971bf923b651d84b454d2e
zbccf149e7ae076d141334b5f6e228e5f457e28aeb384925317589f5840843a503c3a61e83a9c44
z3d1a7ca3d03a60ef63d6b67631824e487c39cf999470b2c0c59deb9c366e13294247f54e7cbbb4
zb8bb62239dd747819a263e3d8a344f9ef586a29f470416d188982a99a8e354d19f658767fb09f9
z75637771c251c9b28910f071f91d23325a9c9ab23a0427decc6f9ce692d2ed9b9e7dfed7cfbf3b
zade2eab419362ad2d9fc4acfd397c198723807207e333d01f5dd07679b960ed3548b82574f742e
z66b9b9c004fe54ad28aedc386df7c5640db4fa6e1f0eacadd0cee7e650c3ac7178fb9310fe915a
z67efe473380f8a04913377fb6881bca056e0939f96968f524ec5ac0531c15214bcd0aee0d12d56
zce7fdb330e77bff66494d9de581e2158a3b07e5098cef6fee249d71501838c6832380c95ac361a
z91eed7c7ff87e16a8857cdc26045b8accc8280ee0d0f343e35a8a6f0390dd31b212ffa44c9b771
za1a5bdac193d18f905e28b9f829f234f4583267fe62360b2858f29bf14acd7b894ce809824e916
zfd482a2bd78a48087b26e2144d4b32bf08d40af89853bbfbf166e21ea0cde3c8b8974c85ea79e3
zd6c56cbcdce0ea0e91acbc93fabcad61a5776170559a2f88acafbe661372d4781f1337c020c9eb
zd8d8b957908557761874dbe22696a563f297573029a85069d7a24de92c845f3efe3c2407864901
z3992388fef91a1e8b88ec1e4fdcd5784b2b6d9705fdab318544193b8848727588e2a9f3a8510f1
z271dd809a13c2bbc68f68e709e884907cbb4916ad4628b9dbb8c99ca71778dc7141f2ab5f6cb44
z5aaefc2d2d50d11c92ee5d17e846a73c410126bd9092052ec499f53a3541877228f76850a2865d
z6c4390471b5cc7fb8fc717c48e60c96a5f79e33c80f29c479a2bd2af2d4200dfed7319bf81f156
zee4f23045f07c94c80552d31785ccb8973974b5785a25227361e7aecb13bbe7e4eb59007d47eed
zdb61fe858f0e00e8879b8f03a6a4a89aeeeec16383af5b227bf152b5957c01eef31dff29d8baa0
z3cc7239727645d372e89541e92d6dfb82e6854303312eebfc4b4273b3899d71d34f0126fa4a3cf
z92b8749f8466a16892e2bdb9cf056bd9d9d5bfc2e24de1952fc01d0352bbdc7eb0022ac3febde2
z6b008986f1e2353c9cfee0372782d8f1213ec33e284266073d839e5d9583288477521544f09295
z61c1c45dda809a1b52b33cd3a44a7d169776bf9c2f711c0257a56db1155c9b0bbe7cee6d9c18a5
z4988e86f2d61a698ba256b057fdc307d18d502fc8e3d9346eac7b462627457371159dd7c524464
z6f7f9defabb285a6ac42ba7f81e22c7dbb205de52a3834884edc352307a0daefc608b184a0eb6f
z0cd0d253fdc707e3be93c91cfc95e61e9cba8ff3136129c0703be7682d638d7bdb92cc04b056d6
z31f4bf98ab6839eb6683e18788f568a3a2f77aeb6f1ec2abff6ec4eb216a215f70086b93e66a94
z2addd34e01022937148f105f661a3abf79e178217fd35d38c647fbc6bebb1454c058cd41aa1306
z9d54bfb53bc8685a11958b2525fef0f7e19d0f68b79071131067034140ec81e861726bd1b56bf7
zb5097884b0c62eb2c2dc32c591d4780e906bd6193d8a90f3a63ce335dabe98e0929b537500c8a6
zf7c48d7f235859676cece95ee01ff32e08540be23a9cd155f43a2c457c723adc717b73fbf7a367
ze93bc81a00189ee3345868e48a5e1e8fa84f5bfd4e0cfe1a835e384c1141519d240463c9b069b6
zeb1048ff6d6cdb96f0ba73e4bdb6d7a6353f1d8a877e96ffb5746c9af6f07359c9c77fd38c749a
zdbef537219234871a43c538e3f392a50fa8e03e3eb78617c71434b7647e52d10585601bc2c6b4b
z4771a08af1c87c6c0aaff52142a6ccffaf1276bcbc2beb79c38f4a4b0ef26bd914708421df65c5
zc852561db8aa57b2e5caadcbc448ec682987b6392ebc4b1e7f085cca638cd2e031f26ee8e7d552
za2b4780c94df92d26023c4cfdeb374a12ab601b92367bc836167aebf3169d7b73cac00f2f81fc4
z9ddd18b8135d1caa0143151bdf2cb70cd7ea57a1c571a40f55659875dfc57f1c28a0363263dd5f
z6fd42afe4a9eedc084cef9af6e40c06e3216d31da147680dade2257e5182361bf36d92e2a04db2
z7e75cb77f7741e0d84e87805872eca9a8000f0e9f81dedbcae7ad2d7bf2293fc888535d3fd5edc
ze55a218b967a7b7107ae9652d24c2899329653b9410fd9eba67e333f7ffca357e9433cbf980ec3
z95b1ff65e6940517cc29ae92978c75d33945c30957e36449ead3423f0278dc3964ddc0f2715fa3
z8440dd7a14cc427798fccd2eb9b471102f200aeb287933ffd750b3573d14155ab7bafbc21cd3df
z43226faace4ae23afad09829248840fb89cfa63a2dca116cd23647923c804f609ebf1807254ee7
z187de3ae8275763cf523cb6bab3dd95c5ab33efa5475b4fc75cca1ea3b660f4368a6d57e96b7cd
z77e8cb8648a4222d23572fcaadbdda9fa9413d08709660ec321ffdb4d769cc97f12a96c427643c
z45da1cd4f70537a6cb850baa80a20ebc60421a6fa594e6b7a10aeb0180adcd7b45520bf2923947
z8dc6a5e1024fe12b9fd1e6e84c913565ce9e22d3c17341b2c2f7b970bb3adad472c9e45ed3ea5e
za291d1d9c86377288986968b4f8c7025161f7ea0738b40151561bd0a73b2216a6a18463c3ff372
zf4e5bb5ef4ce57c9196ad85f0d4e6afecb1256543e796e73b50b88eaf4dcd76113ab5b8588778d
zc27de5c06dc87ba6a21f7d646dc691437021bc49d515030248c93a37f637f4e2a91034bc193170
z421aec05b9cb1b1a7c55864f8c26824e18186297177c0a8a65b93ecef25def34458a6d0440ff87
z90f7119a4470742a69ffd4fd414dadc010940592615ad2a81aa8c062cecc468f8a8f7430d7f8fb
z1de87f622c1ef5345e5d86edf7d37bd0804a95c55ee969697a7b4d257aee581891334b1c944b0b
z38a3fdc4d634f4db2f6ba3f4aa47aa9e62791bab11c66e1c59c5ddee8eee8239e0ea9a2e5cd847
z6adb872621319122587e04e22a323e1f2376a7c1d3a3141552c0db2d0719800d12e66d4454533e
z49dd4bbab4f116227ce375368a1b0378d0c9ce6e8493e3ae88d1162bd5d6930a905bbc35197719
zf645a3af9e792081349eeb288606a4d29597e14e0f45321d3842c040767d4b40422c54b951f6f0
zb67a2aece4caf4aa095d665bd6373484fe0601de7d07632e6ac0c8821cd77e0cbc9c3af041694b
z8838968a58167d7db00946b09fb94932d4f7907f65c9646df019226caa0dc37d4bd4bfa23c7044
zca4f64165661d8bf3f7a71ade088cc13cc9306aa14e35984ae48831c91d477f69b0b6ee72674a1
zaf2b7fc76e78dd47d5ad568241e0e1943b90b93708735025917f5dfa428b8ffd39e1ea3abca589
z68f05198911870fb6f66e616623b071a4ce88b189d8270d4402a1dcdf380b9cdceae811e1c150d
z6ad5ddebe39790fca09d5ff075f1091dd1666dc63e42763f68a413e26e8d38db35af833083d454
z03a16cf7c1f5e3e07c473a5649f6de122faf7808ac78aae9fd7631cd3c976199d9629d2afa72da
z5d89ca2d63c7aaef901aaf13ffcd93899351ff9d28bc02160848fbf7d07ee266eb33fbc7975c17
zfa1681a0b6c884de070c2539978d3b4c76477a292b5dc7d90ae4fe8ae65cbce2569f1ceda42b32
z17360d31c54c8a160cf5e31782bc365db9bdb74fcce455403167e9a3e844da9cb769de363a9fbc
ze0f979e16a2fb64e94211af2d233c70a9a1206725e1cf81a55954543abef77ca624e5566eddd1d
z3c814a5ceb3cf12e8ae6f17f0cb16b200dc01b3a439a992e62d4cfcef57841885556b357c40417
zfac1816721677b3b8b4dd3b3b275a2028173981b5d1cf300bd640f6a76548b54521a005f642fdd
z97e30b21592a2d058c41156922837149d39655ec9af8ad2b7a763ede5a1baf13650cff2ee29ae4
z37dc7f9d8d58b12fd0a5c9490ea3b224e66ef0f135079262668223ca2bb69f9e4a084c0a25bee7
z927bd978acab99de4e4c3f39a214c3ba0f004f6414a09ae8320ec70e56ab4bbe454c10b1b0b59b
za2eb61b2191c1048e0e3be07d7e692ed9a8ac28802f46ee0eadf2a8a3a55be726c1d06fcfaf4f4
z1986231146bcac8527497cce3e04cde7b4cd29076f3c22fd683df32fe537038cfaa6cb6035d422
zd5334a6c14d48cf55fdd03a42dee08cfd6fe4082d5b2fada2fd437e8b365d8ad71b79d1abcfc23
z16bf670223a40ed70edde96a0248477a4055b4cc68f5d431c2454b3fecd0b1288af94165d4cf7b
z3245d24b0c5ea4bbfaee50e27d0fb882b90dd26b5917c8de7180a8ea9d532b679796d703b14240
ze281c62fd2535877f4c1f8ad781acb0bb79c1cd139a5324968d97e0a5bc17a2d380ee274cf24ed
zb7b12a658b1e4efb3992e408efca6de93f6ba0bb82d33a479b25e9744e4a644589fa60f5087b1f
zdc8e2b6c15c7638a06a6c82ce0e2596c9adc5304e08a51625d5fb5dc442e8d1fdddb53d2a612cb
zd178264e8b865ef90d6320973036c4299d3343fc004e3f3da9b027107093c6632400d10eef255f
z649528b68d4a20d4b32f720c60734a1732f49865e3be24938528d3f2b43f660a5daa93cfcba8f7
z4b45472b4bc0c211c45b53851cd8dd10c94ab9471cb448ad9ca4ac10d2a5a5f1ef0297c1721ba7
zd28e8df15d5c3687c334e453c602ceeca83b120e6f4b8be16a53ca29b4301c87db9be8bbbbd8be
zeb002f513d9039ee06e9a0725ac067fd05079c6ed5fe8a30bf6fdb11622dcd3f014053a0001ff8
z5abc463f37f352eba18d0a3ea05e93cb68aa9bb422e7c2eea3ff1a279e06cfa6d7aff1237a4ee5
za1e28b29191e667763321b3a1a1f9f2bfcf010352519f5347c4f7f3dd2966cb7523bf76e549281
zfcea8f899a7d00be10f52910e6af22924c4f4b06d9e364133230baa61cee6864921a6844aa71fb
z71f497158d57c264bdb77b8bb4ba13ad1f93d90218468b8ea75586e58ba423c464a461491eab11
z8df7d882de40576c06186d3649ebccae43227483eae925bd07238a14e4303a1c70147d5ccccb6f
z2e58b64a93bbca8addaf9d2f8e1c0c187497079ff9e36b3358f5f0aa530b1efc8a64a18c29be24
z2a5f44d466725be3db96becad5a174dbeff80ffdbac1e28d83d34477559d09920287454c4df2fd
z3cf906dea02ca98d6c6d61bce55102a000d9e7776b9b30259de8192a4a1ec9653cf02b197466d3
z84c2c4f331dc8c732ae561768d1ce3eecca72c51ade81ec2785209bd921368905e50597f7aa724
ze8d2f687f1b53bb32c0cf37f1ff7f83bd3fdee25af4023ac46505c92a45fae4827769baac70150
z3783bd95bcc014a2fb09d98a0076a8c7596d764bb2fab079b12e388e8724d631a6dafcdd8d7690
zc6c6fe6c90b6e95ad9858597ae0d1d10db40e7f3167fb303c2cc9cfc4e8a2cdc374e008a2a625e
zb7ff95269289decc54e5f9fac92a0da465be08ac9f0d4e21158c04da01a0173c91c8d8d6d7f5d4
z97835b6f658a3ab3e17c40ddb1f1c34addf7006ede905dd1eb28c3c6a1b78f94c923adb00bfbaf
z4ef49fbc2d5b931fd8e04b93da14520846516cda832cccfecf663f06683b48ca2767f0afb7a012
z5613af64654c15ae9b983ecf374706287e05ec57a204d0a3983f2c7237de96c4dc54b0734ce826
zdb08c4781a319521660e76b6ba8b074bffbd21ae9190e95b66807df55ae9160e10c7a6321df52c
z4419d4cf2fb46fadd193471dc415e244ff81e3da3ccbf4e60e0f1c77bb8063942528e22edf3b97
zedc1020d10a1eabe214d3080a37100aa1d9b2efe9cf01d1f6acea9c5835a8ab9e5b8f98f2892b4
zadfa4fe91c969ea0a21db6a3b35eb9d3df823935293da9f617fb744e2374c036e134661e27e6d6
z37545b76361fe9bb931fb3231650f1cff13443275d1c0918b0ae3fc052918382822e9dfae4467e
z35d1ba4b3ed002c4215d04ae0ce855d4fa7ff527dd3fc8e24466ff07c5a9625dc6cf297a165ca1
zf60c2d5d44ce16df7cb570c5d6d493ad570ec9265b61659785a0ea638def018095bbeac064695d
zb7abf228c5b8e5e235ec6277fcad510e97348aa231f7f387437db7815c157a09b3bb8bf17a510f
z15098c9a6c8e0646d0ccddb15ffd9d743ab36192c8544e4ae569c08a534ab80be0febbb199771b
z9dd31c5b6f689852824576ed37c597385daa670228899dd71b26b2b8bb457493269962ff4bf7c3
zf702c997c5df3a95c4054e4eb962b7f4b38037ff1733c8dedcf64a7d0b050fb6cd9e0c347c2a48
zcfdb16573f0faec2fa7dbd6affaa627ee69b47047cb2fdcc3d7a0625e318614f7c3c41bcf291fc
zbb91c811516d73f134258c00e1e2e2fedc8e376957c009e2f7b552492473d3a84b397e64f1b47c
z8dd9031291ef797881e9b8da2226a77958b41bc0f9eb478576ac10131b33edd548cd9f5d3e41cb
zbc1fdd59b7be56200acc431ac2ee6f99719c4c08ffb10ceebed22b7b5d1a2a7dbba699590fab1d
z7788b2b741f2c20ffd5fbe73d77c2ce1944975f3246eadc55bee8b6ef1204ada3ef41c929f6999
z1d744a9bdeb0986b010654535ffda43c670388c097c94b8cbcec5a81473642800b7fc24db7d87c
z4a120a948c17d48339be62a965c859a9cb59bb420e2ed42229eb8b049919045889f50145c5e5c9
zedcf1072b42c9dd06199b838396cabf5da2a87a9693fb2ed5e38ab1c7665b72d20610d8023b047
z1a139403dbdfaa0a99c02dcb22bd7c7d501f03303fe8fad741444bce7b046740272619762402ae
z044d3e4443fae1cd047340d30932a61696afaf859da1daf6f15366220ecb474c0fbb145acdf21d
z7e34440f6ba2ff41bf202dbc3f54bc8024f650a014ea8c9e5a637248805a9fa78d5c2ed0ed24d4
z9144165aa9f957488b554851e4134bb478e80eba8b73e634ab624459cf074987f7b91ebaacb8e4
ze46e44f459b0606d6bb1cd5bc1bb958c62b828bc79a29dec04144e4efa0f64989b33a04dac886c
z266fa2650afa0b7018496c164ade7b8541a9dc1785c307afbafa2c184ea6c151740322f57e15b9
z121fa32f025ae59f2678cf0828c94623af59e9fcdebe24af92e3dc4b07dc1aabeb5b8e22697991
z15fc1e08b2d4dbd970514264668af0679610f2a1f1c3d8489f1c0ff8412dba96ea3e1d8d6464a7
z48b22c0c1b297402bc0a2929b92bcc6e5215fc09472357ec5ae87a19032bf4f74b3778067f9505
zd2b725d7480c6af3d1d695b0ac1c2a865352c2d35f646b087d56576d5585c45009db54788c494a
z12736099bffea7c7307bb8b8801af0dbcd6b1e52df0027e22a6cc325a1ab48d292356a9810ff74
ze3e5351a6f52f06d6cdcc975baf9805a633412510e9706045cbb928f4e0089ce8dc75f3388ce55
zc16084f642c7317719efa4db0e17eeba788bc861a9669bae4234f37ee830460d9c3591b8492b2f
zb6624d6e10810728da12ced5ea09911f818eb22873ea26337c7dc80405fc279125f24c13933a33
z53567167dbf1c48805eeaf91f68969a5b8a3b159280e682b3fb5c08fd992347098a6d69753b762
ze66de7a13e6cc047468cbe0dbeaa32550d44f93bc1c34d2a60c66638e38f4634ca46563dfa9fe9
z2f091c5a1b1be2a00d95e9039dce9905c5dda05d390db4f2e892ccd0ce8878acbe4daf2a47823d
z19ab1671425001925bda286584431d9121627e63a5498dd1c634212bd92de78e2e921957f9e1e4
zceb6d228bb0cce8f34a2f386a9f433961999689051e6bed854eec148c3591313c1dd10e5125100
zaf9720fdeb69c1a1e32acd115afab716acbb67c974c9546694a1036622103e7c265eb3c1f706ea
zd015d8b77d7d7660adc6a9954e6b365512c5962ed6d81c999e5213abc8f4397fae6feb50625c40
z1338ea11aa427677daf5b34599d0c394f371355f26490e87a46c3fc7673ca8dad68927963a1186
z15b8e5ceacba033f73f791ec7538b06ef9f1b0b7372e97aad05640114d929a53c02af5355bf778
zebd95ad2cfc96ee36dab7a02e2b8c87ce1d3e0b5df11e772c0ecec85694c33906c015c3132b6d4
zc5492644a8a598675b723471856036a4c659119c47eb0a3289cee6d21894a6a40ccf0248ce64be
z5ad30b32440f8c4e43b458072b4c9855c8bf3965aa9ae0ac966341fe49c72eebea82c35ed6c72b
z776b533b30bceb54ea19fdd6042a03310a83a6b2d9c254551227d0d3b72bd3d6583d70ce0cd969
zb834e9f994c1d3f58c07571cf6d8bbbc5b20bd34f5388594b33501d0d9ae8a6cd811a9b8985f87
zf4de11cb91e2e4350564a07f1962586ba2bb804a3f4569df74cc81c2b09f4cefbdb4acd2d2930b
zf61b16cd604ab201b82e8b836429ba9ed49efee9ebc624a57081c033133db5110a2b02372d2c22
zd99888fd3c46aa622cabae81bf66d51484fd56fd76be1e67f29fdbb2e5774580bfe8789f0a8a9e
z2ff12cb88835c27295d7dafff33a469bbb8dfc6670b9c2fc9f17ce49065544aa7aedfc2bb37a66
zecfded42cf3f0bd6729f5fd1ccba29a8e688267a0b0ed7745c46f99945f17e2c99ea541b352e71
z878f0bc06c0deb0b89b943941e851416b33561138ea57abda13e81a53f8ee5fa8b8f1d45d0d6ee
z518ab7e9890bccbac138ef690c1ef2ec1a5fd5723fbd65eaeb5b4183d4618612c7c2dab105b783
z1e26237524047be103a2597ca37beb2ff4af821fbcf96b955d7bb0f9e2efbae820a7d2dad7bcad
z5371414ad4387e56077ade9ff269ed5cf506191dad243bdc58c00de5ef660d1f4587937875ac74
z145d3f449ba542340b4bdb37fc1867fec8e495a4bfb5b3e3a3f51ec8d7b870343f657af7988cf9
z30e88bebaccb43850c4dffa1370fed0310d94d9056289da55e7ffabac104eb66bc3f91bbf698c4
z2e9a8ee1e6938dc03e0d3956dd883bcfb1e74c3cf4338ef238b27d36d4adfba912f866043683ec
zf992d7995b456aa08d3d41340628f11b984ef242e19a6e77db3c352833edc8432e7f0e40997767
z201c45ab0f47323eb8b34c79b1bad4b86f8d1d6da0e59609c6a09fa867ef347308c033ce13dfae
ze01c8bb4c2baee15eae2786a0ea01db092dee08a8a4bd489ea268fbafcb25ff7f32535176ca896
z9f33a4a5408191f8565d2d9e1e0c96df2dbc139c6d400ff86db93f26b82b3e634d3f5e41d81a5b
ze7c305e1158f9d472e74270be09c49f12a0a81025d2d4abeaccabd991162be4123ce47e4fde38e
z43feb1a35abad7aa90748d8e8b32dfddc5c4c8c0dc6db582e8dd7311ad40261b25a0f0a56acc43
z22e2e7676c65723693487f222a98d900cf202b4db171792a21b45ba7cb24666b67758e83fff048
ze973193fac134b155d18da2126142cf10e78806d1d02c0fece8836164e35a9a56ff5f3f423d732
zfdecf1dcec250f4c5051aa1c1a733a665f01c16c0c819ac3e540cf3364e8b6f968124bfa8dc363
za0fef2f2be23c7dee03005df809493ddfd88c7c238a1bd26ee3faf557cd8600cba71e524fcd6e3
zead9bb50d6c97669f50e7f87c5ca455da55f4be1f0328fb356206160f1cc47ec40a6c509cf344f
zf2a8e3a8ca348f78c206c537f4ed478172ae1ee4c0a1eb3d242fd9ab37c76d3c8e69f34f1b3846
z2fc92d4fd71083f38610ee0c84555b9642602d6c5e4f75bcb94e8755565fdc3cbacea27756bdf7
z858267ec48601dfde24171d69fa84831fdefb26809984d31959f1943a5443aebdf9de65e356d3e
z7c662a84f8e1b0fb10c35a8af6535443289cd765db9902ece0b5f3bc7d5f967623d349e2fdeb8e
zc6312fef327a1012b347cab8167b534521fe8bc31740a8e008b4a5bd59adc77e32115e8cd19289
zfb4fdcf8fb3284b14f695e5494e4c97d6554b65baa2e618d92ada4fa494da25e44c13ac2db32f5
zda8ffbab22b222c578f91fb14918daefc5e1800810adc3796502c3fb7cee1c19140730e2b5c440
z29910055f092b3df5d4a167f0d0474b137df7580a7f21a3a1b7f24f34c8ae1c150db84daa05738
z0671aee95fded3e6ecf69d48e86a3f402e71d744e3ecb0e0029211ad0bc531ad22aedc09814f23
z71fa125894a2930eecab28185670b92af0237491841591c8c5d43f063e990bb8e7208dbe5691d9
z54e847ad392785366afda279b76f0d9f9d1daa95758fdc6878f3c995ed7436309c6c39d412674a
zc241f285ff0482546b46fb51ede8c445a8249d6ebd9ac33224024ffc6ac79427a63f3c4dff78e4
zeeba5fda1fbcb46228da55914fc46f5b948afda0d5d83d3dea7f97424614bc041f245df7807abf
z2b3f3ccddb52685c49f2521d75c9cbc379db48b23c3712d0ae9d9c3d8f7029b555c4e02cba6b0d
z01ba51cf579f45700002c480e69f812e02fdccc9817ccc6cda985c4432c529212605729f32a9b5
z94b379de28a85654f9370b2d2f8ca89fd63cff7bc2384e88ab7c435e0e11caa4e6a632e1663201
z91d84b27ce311d4e6748fa926de302cd5b0eb4149165654aa7de191068cdaeb3e8a28aae6face5
zae0656cb6448cb8ab89cf1d1ebe8278a5c86d7814ac04bcbef41d8c9f6b00982b84889092f3223
zdfa5ac23f549d73a54c159b85f785c8c01892a676703af4dd72d1078a23843ca9634c284b7b353
z44a73a00f584d67f746979832f5a73a786a16b2069813a0e29ee8dc8634ded5dc2f1bf39a66335
z2999d64c93ed1f81b4a3ce5d29ef2881619818deacc8fb70abba83b520dc1bfada7088bacf7abc
zd955cd834414692496cc6c32010d6c845d3472b768f474a182c72ef2dda1efc7f0f766c07bf578
ze70933059f88ff02647eae78758a0dcc2f2c23a026198d9c1138ec5421fd3efd6f289ad2019061
zb4fa82d9a4a8ea26a36a25485c57d1e42bb15aa7bde883cf196400ff156373c2dd05574166e16b
zbbac7d82a3146576389918ae1db87f0d20396d60da7b26deaf16647db434231b9a16b5285adad0
z6dd7dbab00cb5545db4369ae97f62b0a3bf06b42e762a5abfccefec9b65ad0fb0f5408d4f8f85b
z79bfc7ba446986e14af0bb91efa326038d6ce60b3508f13cdbdd974713dc89a4751267a9663a38
z1a4198a25a1038988460367bd63955eb5635486b769a58acac9a3ef3c44882a06e732a105799e3
z5c563e529967675dac315b6de097acf15fd7d4e955ecb2fb95e344e7f8e4121bbfcf02c16dd085
z746dc7d2055798339477edf1e2
`end_protected_0in
`else
`ifdef MODEL_TECH
`include "qvl_serial_to_parallel_assertions.mti.svp"
`endif // MODEL_TECH
`endif // encrypted_0in
