`ifdef encrypted_0in
`protected_0in
ze74c34e226135848fe16db9ffd31815111b6d7fb642c521a3f628cf6da949865580b22efd062a7
ze90adae0e65e66a2c36a587d0a790699161455169ed55a01f2084f11770a774ec4c588039b380f
z6de9c5084882a40b79a175f5c2114b2b6d78b070cb806e1c0aa9258297f4687ab308bc470f0040
zb0b1de382961eeeaf2e279e1462520fc31c119af8f2b214846f56c2b3cd2eadbe4099496abff18
z15cec83ec4a77b868344aa20ba7360908f5c0de2a79abf8b3534b883bb12180f68b5d4beb444cf
z3fba8f13afb0abfe8fcc4294810f75afe452434d2d0f1166236c82f76edf1e12979f04bc35693e
z32ae028996dd85737a8f5adc1ebb94f39c940246e887647b64782cd7ab429b0544c173176cede7
z01dfb26b1f73408344a52b7e1f117f12bb9c8077b34876c2e6fdc085981637012dc9754765e1a9
zc512ce062e0b8fb16a214591f5c81e1353b900a611fe1f4886b57940b41b7f2ce99a7b84b04b90
z916f717e73bd10589c81e207ed77ec660a8cbed5b487fa50acde1b055c8870bd8676023f21ddcf
z9c98cc47cfa2d654ff1365d1f45035a045a66c5dfa82790502623b57a3af03bf0f0c0d35b51558
zb8b5f2d29acf03737a9ca2a053b7a8f06800d50b465c41b30eb585f62f3d0c2c5a43bcd94e7ed5
z4fd176565031310b597fcf51c7a7fad9dba1ffa64d830aef3c6bb60aaa38c7dc51e09a4e7b86be
z1ec9d282ba091476713f296a6a964580b4e9f89419f7f9b327d59c83ae9255b8b5b5f72d2303d8
z28d4a5df8f93e74ad57cb5ecedec731e5d509030aa5810cda25b50eac3fcca05cb3a9e37bb95bc
z56d8f9342cc4d14389faade57e6bd75b961ea6a1c53a86ca282ca9588f79c3d40615552a904083
z87e533630742ac4c708eee0269ab4992fd3c19b91bbda7303ea36dd54a64c630e8f0ad3aaf3519
z7543a66e6c65ea33a357f341c26e7106da3ffedc7fa4f1e39333c3199da46a926423aa11fea88d
z9322892edec932cdbd2b954a8bb998a8ed73efec27da6ced0f27ab9dca89f41bfa94b76006d64c
z1a50c7934c29d5c6bd1e611518c3b2d82fd835c8fcf0c04e8060bab3427362d5ac3441c1fc274d
z261508641122c4498fd12d4f0ca9b3ff760d074a7b048fb07af8696145d7683d0793e2a60d263b
z0d9bc901bfa9eeb22ed281cfd581171fd992113a5f98e8d2a35632642ae6d288573ec093b31dc4
z32a434d5140170999fd97ab844ff065ad8171ecdf6414a9aee6fb0ba004860c5ccd2c3d87df070
za6e7b7a06fcf58b28fc6ccfcbfef6e3f62a166269a16717b5eaafe39367fa43c0a544032e9861b
z6858fa9ce7aaacd2393d7caa7092e913d2f4ef39517434e132c9a43206755f0795f68387b582f2
z6e05247229ed6435c710c1d92c51a0af303cfc462545fe74d8a829bc49b605629b5590acef5918
z0392988101b476e4626ea7b5de1f262512b52e771b7a1b3e55b903cc0a3ec381d72ce010bd1bc5
z983d60d1ff2d28148f2e9a789557d2d8a4e3925a6584342e7203bef5d21ea3210a38d51f65ea0e
zc4dc41a9f3c3efe69ef6a7196ef59e5aed0a513050a8ccc3a3f4fe780b8f2c380f972e2be5c5a3
z3fcd5d359945deff540a2d39288d2049c3a71d15a6df705ff50bf78760d1f92451a66693100f6b
z47b613aa2a337ce2d19d1c8979d3f85e7916124e59f821daced41ddacaf27b59139cf4a57fac48
z3ecd1da19839c094ca42542c28ab1242d5164977834a7d18479a19e06380692ace692eb971c02e
ze61bed23a8a137de91f5134dad5550911f1512b5ff0663c25f2891f7deced69911456c9aafea37
z0e61ae9a47c7f18c478f535e0b4fe7a084f5849f4e7c836fb46e878a875f9488f4b23e9f22fa40
z98836defdc94740be5dbbe37d1cf98a3dec89f4c4955331869814c971aff5d77b85fed5e6116b1
zc47af9ef1fe4ecf9375509ffde8f0fe3bf6fdaf799d6a8ea4ebd539525ceb98819866b81fae751
z3a0c7fd14bb164e85bfa0e6130f7de8273479d197e7edcbb3fe8d2f481cfbbdf195b33311be13b
z002c092df4a2c52bfb747061f11eaecd5f53fd6d02aed3c5b1caf4f458a4b8ff03c328b64cf208
z43aee10bf89394d01c257c982f544501822c836dc960a1e59cc7f290bdc247ec2b7cda89328b0e
za314ad06a65bf1411376c472f1513e061eb0d8c2cdbc4519887e1a2a1e556a672f40565883004b
z0af715a4f0f490e247bdd04676ee9d4a546bd3ebb1272c3b8624049174ca8b65e1f4f3da8489f4
z97c2982d3f8776c08530c4db61b59f73b930b7ee69d4d02e3d8a4a849a53af5126036c45162ff7
zc56baf326e2dc84cfcd56e13d9fc5e41c4d698aa3b81ad04d0e1060ffc4dde726f96c233bb6204
zc2d622f37dde4edae30ab8deb47a476a8e10842a59aec1bd3b411f0f851fe68c1ced6025b2ef84
z540382a3a7031a95e402e49a2af63b799e1f8795eb26acd489079d56b30b79f20a32d0e023025a
z054c67b640aa16ea0a38d88229cf5568b456c0d421ce493e23d53e94f36ccf9a6c8d105654ccf8
zeedf869e62e9fb11a405eef9db90280a6e9eae3174e5a9fbbea02df408ff791e64078ddbb99cf0
z7ecec37a4ac25599baa595f1a91becf74908ce894781142da3c732f84fe85e137ced5fdd054de4
ze46fcb189c33974f7be30db8b7a9af3ac6e6084f0fae404555b5f50bdc3227c40c980a1d1d74e4
ze763e2c9513c71199d550976b1fac625ea82d4ad6c7fddba6efb6c3e984eef13c02c4f5d75c606
ze27564e36d28271d750d3cd1268de0ce8ac8f41d74939e411cc7538d48fd28ebc2faf23dc609c4
zc99415b9a8ea254b79899f230d00614c4e7924d856618812bef145e151a11af96c5c3594f10c91
z9b0014516ad6cf0dfcc5ee402aaf0c4de0d1bd7f0710d42b9e0580084761eca430641f7c1a45d9
z67e8d15405382a4fbb6735b193e23a53379047fc2c6113e83f0903ec2106e1b153dcc885755532
z43060a540499dbe1a2e97e062f81c8fb83125755aebbd2b5815f8f2bc2b35e0581ca880d02484e
z38e24dfb151aaf7dc8b836dbde06566d62a2097b6aeaf8fc5c2920cb0031345ff61d90adbd5c91
z1d699b718047deba44d05cabc3452f36a9eb13ef805419fa2630bb1bcb20f8aa097041259b2a41
z793d90e22ad6e28a9fe4145bfbea9e2e5ed09107fe7b1cb0829632d0ac37d15db121f26206aa72
z00d02805847e5a382dd6f3eb7945bf7c652e65c85679155c42f2261b177cc1330954faed46b733
z5c18d352a65c5d6c874033d33de5cdc430e6c88cfa1a4ca5d83ee55e4cff7c20e2c792ecbd85f4
zf7329ff413fcc2d736b7b709e0a715e8cdc03df37f12590421491ffb62aa5cc45dcb2073cce112
zfef08e13ec8e13790bd05cdf590a3f5f88ecae0cc7de12304f47285a394557e4782c159f3a7cf2
zc82baba56da0e580d70ada65f054c2d34dd4c39f883b04a9ced3e597114c13b61f7c64c5940547
z11255886417056b5b6fd50a8fa2f08124cece60b5fa0697ac8b22587d341f18962273c693820ce
z205a08d7a3c90f66f18a81fad9ce3f58477c6fecbdf8f63ab1f487aee99fd431ec145418b47f00
z45a2e5d209bbe7f1ba6e30001dd223b78879499b852daf0ad3bba8f55116f6127bddca9450852a
z916bcd4c1216ec820d23a8f871f8ba0df4f4fb909bf327b1c31f4e41ada9d2be0443c3cf01171d
zaf80d943497a2481223622b0198ced0de26c17e2ee6fd0780fa45786e8e167dd19368856aeed69
z4a945dfa7084a76ec8c191d1c1b7a096a6e5e7e6ffe54ed840c7837030f2e1d2351ffa65b945d7
z7d87cda3c3ddd343a73ad0b1db84a3952cd5907ba92a734b2ab0ab79d7fec989fe96ec4c5670d6
z97c47cbb48195bea7f8032a77e127f0419b62eee532084d9edd43c03c0abb0d9e56c617dda7cb2
z0566cecf8f5a274b7e6c63eff32048bc1527ace113dee99202810b0c6e9983bfd3fafe7c7a7e2f
z0dc29a0c1f4d854da302c30afa5d821f8374a77372b06d173a68b23ea30c0b02a9f783fc21d5e8
zbbf0717f05f0910203c97d4bc6a72702dbdac185d6f16d70c82be56d873a17eb59d8467208bf2d
zb734ecca06a121b9d055ebc9589b11a1810ced7ec6b49ba71cd3adf747df6431dc3e945607cee5
z44671ddb7f58f5c4a34f77b0516addc2bd1db6e834a80db65bbe84c46186c131b245bacf384a11
zaa5c52a48ac092e4ec660bfcaab0b0ade080be47a8db0034b482316e9f540af810f809ce018c36
zc0e29f9b125f453645f66d48f9dea34b1605d1c7c64b90cd3bf990237758ca88baf945c9411f41
z8cb88416bc84f7dffdf83bf068d88eb127efd130d4d730a665a37b02e2def8bd7be9da1edf8af3
z86f52e5f5394aea468b1f593d40b4cbc8b90c8d10da5a299001f61126b98ba8a48fae37d66697a
z8c79dd4949b2bc6b2edc757c32c8ac204a71471b79c79a966ce34d8a106a70714c77fb200b50c7
zb9439cd960a15ddfbdc3d21bb41ae71fa83b47faa3450803d7de6b36263667c462d7dcb977bb85
za1eb3834a2d4a9233302b9ae1adbd56cd92e138370900652672fa42c047f4309356ebc850e45a6
z5f3f7f97f5212c707f699aa224996f4fb5ac9b5245f7b3a6949ad2efbdb7ca7949aa0b9b620634
zd77aa1cd930133f08b405ed3dad3a511b107629f77a336c605e5510e2d290292e0b1a0212ff910
zd55d70c925e7bd817846736dfe9a39467b8cfae27a4486432b5f8096b52f70a08903c1c972867c
zc73fa3b1b43888944a2adbbdabc4384aded8679b049e5901f1b3ddfd800452459a8325912ee2e9
z2572a46eb4f979a2200bb0786659b6ab8cb0c2bec29c3a6beef3c9151fc06c3d3e2147d6560d32
z906cdb5f6b1b21292399a52c9fc227664bba31e6e5bdde43e6911ea586cedd16a1976d96bd9977
z17f174b4012010f98705ecc90f319e9b83e1de2b530ec768f3d070c5fd876444d21f498d0fd6fb
z4683a8911ef0a3c863e9224f509348b02982fb024dc83e1242940a86974e35dfd826f609e2f805
z50a2506b9ccd464c724ea31ae7d22fc260e2b0aec41d3329eb8416c86da7b838f98dffa6971a6e
z9f95e0271608f5d5d08e75e25e168ff6607e853f8acee3b1f2d85d1f8923d0c4f62779e4e20421
z04e7051e1bf41c2ff218439de72ac8f316c009a4f68857f610efc40e31d368eb8c41940c21316f
zabd0f83d428c57cd6f5c854cd86e223fe46646f721e8b9f0858fa6d37cc0d3db8f50e5aa39d872
ze62785637db5bf8ab996b4177de83420c8ceccf0a06e6dcc7ba9edafe94ceea181f654c6f75ae9
zb4b67823531dd4b9b29b6c2443b9e32c305e271285785fdc0485e7882ea61994e912423b908bd9
zcc03dc3b11a5788e37116c1fa04a13f57caa92eb41ad27e62077cfe5da12b46cd9a15d8bee7cb2
z79857446a5a9e85fafef6a73e24ac017a0b1d2c85cd11c2ac6fc0f4262848aca0629fb825bd45c
zf1b01f22a9d206620bb5953a385e944ac4269e29fe7519ba4d74672c6087cd14b9fdf457305ca2
z4895e95a9ec558ad8f58c47790962123de273fc8d492668a46ca90752d7a9f1ddd029f4424d552
zcc18bd10a1faa6b2afd4a8d7265898e00bcbd9ea99868cb5c2d735027e35dcb75e718e2472d815
z6e306612dc1de05e10eec75444cad54d5a3ba5fca29b58ce539d9bbc00f8dac7dc30edf6e937cd
z400930b478b30178375d09f8ccd4ad128df6423ded4e5d638230e17bd770667e4519a41a7a56d3
zf1dcf4e68a51f0216ee53c583e12fd97178d40eaffcadc5dc2b2a2cbc64792dcaad5663de196da
ze60d77e9c7ed3b004fa29ac2fbf5a4e4bed87bbb378ed6750b12d197678bcf976bc1f5518db9c9
z12f9e7f2fa70e86aa0092593d6152ba8f5ce0ea7376e89163b0dd984c41c33c20da80eb252575e
z3e8e074cbccbebb16f7416f61807091218aeba172b7baae99d17d458112e97634022c601dfc615
z61766db4e05a09715b2554a89ada6a76212c1a203a85b9a7df333377a3ab8db865a2f1bdc90259
z8160295f1fa6aaabfd1ae81898ad8811bd0df03a7a9b9322795e9934358b1d2933f344b6886acf
zcf6aa556d2e1126d7a7742b4458df09bf1e6a198a3b107e91e6c929d261b263b5a204f1293edaa
zae73b7de1e6c47b1f308124f5128f7e3c418e4588ab253d68a551724f6585280eb1e33d335460e
z1f337f83af0376a621fc40f105b6646799a4c1cc21be10a833cef02947b10ab3b0d7468a74000c
z67d16279ae73c5ff0ea71a39f8700d9d74cc6e15f4005aa651a2d9141af479f05fba06e7bb30bd
zc91842ab0573759a362fd8b21ab9ac4dad87c74fee1b98683f0f8586ea6846336ea0e903842f3b
z540807fd7251c515b39d5f7c16897b0e07e3eaa00a24d885459980c16f8f297b0c9c592e3c7b81
ze1ff8b21e45b72c64364412e47772e13dc26afb4769da57e483522f32255f0fb49e87e368b1b9d
z8da10538cddfc172a83e0c01b28af17130be6565fd99dbbcdd73667199117246d94ea5dbcf5b9a
z10125ada53328f3fd7e834eb49385b36dee950a2202a4ac905408970f69c2f3e27544ffc429df8
z45996c095151719f1a6e4f19b123ec9db1cba72a734deb9c260d282f4bb93a3886b5c0804ae480
zb885f060b1c518acff287158f9e10b36623562e6897465c785b539b4d9457dac83179558a309d6
za69ca78023f64020c3715b7a88f75fa15608494d477c6269209eace2ba783335702508b1a67f03
z4d639f5d66cdb97ad7e61172e8252025d9265c5f607d4a695ff29a83e0365c00817043f74aae84
zb71406a2d0950f02892bd1250a3209f412642cb853dbe541b27b0535d0f5e88ea917df0d2775a7
zc6307cc3c87c51ef2d52ae38b560a9e4c05ee2660d26a7700cc4973bacdf01b4fb8db6809ff5ab
z00ec046b6260e603cc74527ee31c5f42980f1a17d18f8d12c30f6c2e6482752c6dd73b305a9a77
z30c1549618495aa15455bcd3628a45419d65c0e06a46bc6284dfc8ca2e251ef59da5ac99545bd2
zea3412386b909953b69489f24c3741222975ca6505a9f27e33dd2eab8af1e4931f487302af92f2
z20e4ed9b2b235840ca610b6852e76cde4d6f91573dd4cc281b0b3a20905ea6e4ec2623753a25db
z04e20534766832759610503c3a2931c5057323dcf268abf4b07bc109d9d6b3f92d335f77502335
z60b8a072ff4c8f0a30c18768534989ff9810bed03f56310d866256da07a79ea3fd89de5e446ecc
ze0a336dd559142e2202cee00bbd0ff8b4f348ee4ed5416abe103c1ee9cd71c124f4a1631042de7
z095f3fb824d061d0553b46d48879d1fd6d027af2d2aa185510d9610a925cf32fdbfc595a396e87
z3ef47655818bd6120d0fc3f06ac34feea6028d0515610e45088eeb6b19c62983f24915e150209a
z63fe9b8b99af80cc6bac77329213dd3b2e564165bd43b57eabd8476753772e2ec1caed7ee87f91
z581ec933bf7275fa3c5d0556f066c7ee8f0e16a0e86e0def357e03ad4c57e6ab23e74bbc83679e
z9e2b148df63a71e2c809e356f7dcebc0a2fcd1ca0d0b13cfe3660c9ec29e8f3b2f55a6353f80e5
z9975b38a25ecc2c1a3fd6aff19d8d5ca3138484749fcec7cb64ad770d172367da1bb93bf27e3a3
zdd046d0e4523a2e1d72816fa61bf43d15240c7de104d23acb12debf0ba67d4128ff994057014df
zbacdae4da8f382687bb61573ea930d38d0f7196847ac3c2e8ca0087603e5ea6b80c11eeb771999
zebd867d32dccc182585541ecbaeaaf4b00f75c5c679702f9080d46d4f63620e483e0e0052b99b0
z7b2407f08183aa0cc968c0e0e3c3aa2711352eace46c9e33cc34c2860be5e0ac93e2f5552812d3
z7f000e4f0ab5e44af5861409c857a95f2bc6cdc24e9bcb39af90f6d3e92a7ce7d67a5090e744ee
z3498e3154ff93ac2110a249f39760b59636e5acd83a1c387932b539cf4f78bdf97689a01670ef2
za2fafc283edffa56d1b8deb8aaaf11d207b01c0407fb3c1cf00f1b25bccbb076ed63a42c53353e
z0367bd011ffc002051efbdb71122dc87423d4d7bfc8da419d2c1686285178d4da659bb695afb83
z6a9de525c798adc579cb57b5d376eb093b61f8e4c0862079bad0662d42514431fdd38ae53c4468
z0bb67a50d5a20789c7a88424c1bca05f7b3b01e17329b7d2d6b958b2bc21aa7fa61b20dda60406
zd8d7c74c86044b4f710f21be3cd7f65be6a31a0c50c73675f79b743c8ca4be6029dbc5126b4570
z1c6d4e3e0cd24fdf978d40d7d86b84d1a13dc7ff8fa2dc9ddabf0fff8aeb16247481c206c6425c
zb8e92341f4854dd17432ad02316177a48c42e5eaa4996bd00c9f3f6512f1c8975c34a31c560dfb
z2194c56592fb043323aaa08669c22b92cf62795595b88c38776fc5d4a1b14ca3da66b1ea681817
zf6c9e19ebc1d347581380623cf313395d2db988af1f68949c8de8a3044f88a195eadc5b4c01e2c
zd6493bb2d7ebce7b42cba29f0e3174a79928225adda3379fc84305d4722941c4759d9219ed5f14
z08e552dccbac574e67aeb643c78399950033fed9dbc78d249704a6d13566c0861c41f364541f5a
z7a3250dabfc1c2da8d96ebb420e1d0ebcf3edcc4ff92346d9be601acd353bbea936e2a5791e474
zd6229f9ca7b71dd2fa5543131ee2e4573f68dbd56d8b618ab9b10cccb7940aea836bcfba16e86c
zbaab3f00d8a451b621e69f58c0fdcf255501bd1c34d32a7ac8e59cfa6724654fec1e1b0bb86dcc
z1d3e70cda01436a896c541d0e862b013bf0e3adc7daedff08858ccc54ba9f4a3ae82612f2f2682
z9a910cdbe2c1eb09bfab2c28c74ad3630e815e0c82fee19aee00dcc3516d796c588d2c682dc11f
zf1a4eba8edf7d48e61e3a74ad7d3db4d82d79d0e7c40fc898e126ff956ccb701a0bae5b04a5f18
zd5933341197769e4d8154a906fa941cc751d11ecad37f44ae5369b810ece76c6c81d3899a362e0
zbba43f594c69e589b16020ff30d79a54c25b2193ca5094ed74178b23e50afd5c04e6d1dfb45bd4
z9cdc5faefe0b2d5e9baab60bbd4778d675fefeb31072b2cd02ee3bf8349be8ebca079d560885c3
z480c58b2973b5fafccc5162e32a1648ff460bab04a30fd32c62fce5384774342df79acea6a108b
z356b9d65644c1f994d9565a7cf95a168679f8bba516d63fc33d02fc15182e0d6f2a558b10d6f8f
z903f0668c90fdbbebbb3cfd04f94f4ae020a4887aaa36136e3f82bdb09e666fe2c07ca95c79039
zaf99b597e706017276bc6a3eec765f0741ab6bc90594fc3e2c605f5537a1d7238aae4d5123db57
z85b2c36adfee859b3a260e3001e5f8805a8993f97b8d9144fdb6c21280f4812d6d8eecc33aedb1
z8c3ff8563e36a6cf5f066350225134da53266ade998bdba2c9e060915b2c2d39218833f0ed852d
z85236db81e4577c4760325c526b669481f1dfd45817bba6a5d202ddb11746fd00181ad047dd027
z15dad481e28e0391ae0de9ae33cc3755b2143cfd48012b16c54e9f1f8c4f5754dfa6596e8cee35
z584308c64d7dbecdce47400b381bbc5724843d75e1a37fb68b1e1ac1eb26096f21da34b8fc3ba2
z033139e73b2b384120ce42abd46fc225cc6dfd4c574ec46be1562bd2ee22deff9164b2d24075fd
zd7ce7ecd226ec468f8ba1def6046edba720fc617eea3c8e7eaf61dd45b75bc89008ea90127201c
zddd271bccb5cfe01a7ca5cf980fb319936efdc1eb1eae8f9be9ac2b96af9d85ce34b79e36c3e92
zb8eeac20987f1b6ffc3c053a8eb1a6dedd3d7cbd3669ebd239770f1e3549996497d8ada41c52cb
zba3b2be589f68a9fd9f4a583f642062fb938c79f8fe5158e33f2b480ce4894455c155b1ea2429b
zd6a79e8790556a464bf692374c66e2c48a861d59dcdbbaf7818662c53b5c6f14315480f207d881
z338af6773a39df550ef49e6033903e57e61ccb276aa70282ea6d5efca5aca23ff9434baa601dfb
z343fb1bc4edc1d9f6f6f8f630acd329b0ad0c5daf1d07d0b69dfd0d4090cd895d1528ecf8a5da3
z6e735d925bb7e7be1b9d2a05a6a2787442327d93ee0a9a3b2fcac7e8f25a01165456f1cbcb83ed
z9e9396ae52420c932344486dbe10857f09d5f23b11264225c0b177fefe10e2268ab9781d9e5105
zdbb4c37d669e3e8750f5aada36947a729b5d0b6a41ac0783b1f8d3b1d6f23d7e1f4d6b4fea8728
z9b85e4a1c2f344e5f7f9a8f55b88e9369069b714a75b8d640fe9d30ec73930185e1e089224f8ea
z8495849d5f9fe2525d69bd1c7a189c0bde8984911c0d766378fedb87bbe0586862d66a65f941ce
z438923ef3a0ecaaef739cac4ff7b03ffec6208da7369c15cc775072bda3e9dfec1005cd62dec37
z9e542a097f36fd072bc53ce46530875fdf166636a53beba35cdc2c4d3194d8f56df19058890c63
z4da857fab2213d2563d228ef7d6151166f58de0f39ab11f7c19223ea5ea5aafb38cb543a75b3ac
zcb5658a3e3a738df0b2d31397ff57c2e48865f4e690011db4ee30e5f6a64b78646394b5917b401
z904f97f29bd066e23e678573b8d815b3115f59a280662305a88cb1c52942f04ff600eedb5f6cf4
zda18444d673f2a90581953674310bb10fe1304053760ba65a79ffa865a6fcd70300d578e3d6ad9
z79ada840732ca6a6e461f3ba0a7838a0a129ef773b54d88eb0aaf47e33e54dc377184a207b0a56
z9c3a5f627d6f1729edb5a23be0d82b341d3a408a70b3d61a61f6472b7f7b9068beece7fb2f07f2
z29ab96f2524d0320a45882a0e4afd95e2a382213fb1d351f89e0f9855c1a361e4ccf6491ba9a8d
z3c9ec872b4e5af6c16519c8a3a2048f164b1d3f3869a43785ced983d32e1c9f68f3c81034a7191
z711b41cc3a9f77afea20a3bfc86b9aac3e6d300dbb9d58bc7d0424426fdd883278998313430aa2
z42a460a6819a1e954f133dfc7b66aa811d4ac26db1b90600c1aeb0e1c5bf193a3703f64392f93d
z9a8c74f260993fee9cf3c829c5244292dfa272f72573d05969ea33726201f2a0ae5a60b0669d19
zefe9d3df0b5add169cdd291724cbd1d685932c64a56cc17d26e48f17639f1e02e0eeeb8238205d
z9505beec07f69a4d8924ed0768b4dd56eaeec95eda0a9eb7088304eff43ed277ab7ff0a4429b37
z119b92086952a7a781422259e49d10523fc7d78347c3ce834ac13a2c6895e98f5f5727fd5c1821
z207cd2ccbea4afe537ae96ff33b4e5029c8eb78cc04952bab96db9b914daf2cff74338a09fa5d3
z07d3407dbabb2be88035d4cd7597d8ebbb22aa5dfd838e7c1309b6e047c38a73e0f983d3db9c25
z9493ead229eb9463019dffb0bd19230c74e01ee4db29cd7a478d2d2e6bd6c691d2fc80d62b46da
z536c7a869d7b9fae9d1e467995571945e2adc92c7efb5d0f0c0eb97906938f5d6dae3783815e84
z78ee15d5f9ab84c613ded7b13b932d31acf7e6e5a614fe81af14c25abc2ac3799b9aee63291913
z90062fc97e688c585d914e6aa35b10c16366b64bb53b35042b7ff770353bc93024b415e1a24d6f
z2beda59c7fb8829da6756ff5e2125646c5747734b70ea595e15c188c86e8a0b237b72b70b97b6f
z69e35d775cf6dd81cd95d8d040e02d59846bba5d71741cf605ae57ab8af6a0ce0e82b0807790cb
z05c8bb911c2bc1f2227fbab96598958673eb9cf8a02b00c150e3a659f046fd1d0194d7457d113d
zd636b64b0935c9e0abaf71ec9de6b6452fe48c5593fcdee6150c6f56123f5331e1667bd51de3ef
z9646a17e438a676f3e7732d50f7a162e2f1675370a52a6408a5dcd183513428e28e0b7fddfacc0
zbc7cacc5d91eb6d233b17c88621fa6b94fcc14e8b0955132f792921d9670dca0442ce87131aa73
z903408487b16b044ed71d125142172e589606cfc266cfcbcbbdef548655f9b61807496b34b53ca
zbba03342f3664227144ec805c6ad357ca7bce6d1925bdd010f4416cb289f07b8585fffe5f76078
z0040804bc5ea971d3ebc1042ad840c261d27d9dacaa04fb0281ae16fc1e35d99235c08a6d6f0b4
zd6d35c9faf3d1150678c376dde25ac76f50160a01b2241d7b665121e05ad27345e1c5c6221d91a
zb82e04bac49151b10fb53914fa2b344ecae5b42d974f2c90ad98bba57f0a36cc3bf76fe99f4c91
zbd9d535471608632847ab20c9b5cd5895ea7850c332d8f77d8489579fa7199a815d0c78854eb96
z2133375de3f0e5f6a0a7184b58bb23a67f14c8bf5bc7efc820a2c138a343ebbb315eaf229ded00
z6a7f338a71bb569df5c83f3bc671bc3025e1290705411b91e4dea240cbf2b45151dd8dfaacf37c
z99bf52f8a4c3a50023ade0b07090988bbb25b63297885446a833b455794ef1e9b91735c5fbe829
z907e184fc53932738e3b21e3ae9e9c1a02c9a21fd4dac626e8d7d69b393b3acbabf4444634aa92
zc5195141b17c05464cc44c64f6e0f27d80159f3348cdc2f79e57f50227fb8a6cfc97e172939d08
z384bdb7dd842339b8d319ccd3899026e689d311a204c2af48748f8aeb254d373c194382916eb85
z0438911818a3e6d0e829f2961bc77c422c769e262e107353448e706dbb90baa7ab07e28049f9f4
z8566b9815c3a24506e4427918e702b509960f5a3d8836e2728b7df83e7d0c5501f9f153058c189
z75a0a07ff41e8d1683530b12e5681e260de90a9a23355ff62bf0b6817a43025b47f50f0ba5562e
z1e28bce9854971f0f718653dd06df7f306daa7d49359acc6c88e7695a1510950a8389e21616d4e
z8e1a02b7356dcd2f9ea1fef6ed9d147bd34fd19108f7a5070a8648c58773303a9d2d0d30186268
z59681abfc17f53fd43bf31c14c2a8b41537f178789bd6483d852b595f534d89c006f849f878495
z07fc24c7b2d229e2a26893646b7efb8496165915679d57dde334f31e3ad9577931a3429292b5ec
za7bffacdf11cd8a3e9c2c63ad26e0996eda54c183a7b44f154e2d9b5b13caf93e3ebf719987138
z8f1442c9722f36af861e4750f381f8f0a6c8411daab410a5b19a89299d602f760ab9bcc9062497
zf251174d81ec792d879509457af0e99a19023d93ffcd71f90b8ce1e231f422b50bcbfd7cf3f055
z69667f6f4ebbf3af3b8695d0ae11542ed3e0b34fc251ae0f6165c8b3763b0f9738942e8992f64f
z8ca0432118cbe0874aecb6db2609a09036eadd8947cbb134fe764be08384d542db3d5417943af3
z61ae21ddab667fb18c2ee6b2fd1ee0d4dc3f0ab19e0c32fe9d331775f574e235cbbb8025ae5130
z2c1c6a2b577df3ccf083b53e77bf93fd2555f6a746d569dc2a97cb4dfbe848c888c548673aadf8
z00554af2fe99168523bc114008dff03dcbb038aecbfab8a128950b9768267541f4f78562245035
z6601ed9220afb4be2aaf08776b3974908d272149034fa64ae4c35bd5a65299b5e1c1155dc72262
z2f761a5d88acd0fa0dd68d5198f009773f75057db6ac87dc3f8b69dcc1a8e7c5e40d74620b26ea
z34fdc6dd2fd4fc7bbf67abccaa25019afe3e966e61c114f8b73ae41b7c7074c7430ddafdcfc539
zd91f5bbca11d4d4e40607ad8e570ffa4b1f0fe9b42408228caf8456d423091fdc4b831d296ca9b
zb08406c4d6fc218621e81eb01e9909bd15c6ae320f3d7ae7164325ea8b1e7ac2f2ea4df117b326
z46ecbbd0899263d7ba280055d11b940ef030691089ec1a51a6e5f162314935b69d7623817c624e
z7333fc159382723b5dcbcfc6476a3cba535b1d94bb71ec77ffc1fa0623ac4819a4911bf7c315ae
z71c8253e593a093c63d73b7cc8a7893a835dacb294f4e64acdc6abd395e79b7fb013ed8355139f
z316a17e28ce29f11067785bc85cc2929afe439dd1cbdd22a0aa00bf2e871651bf84202663b34d3
z192722bdc00119580c9d0a26bf087eaaeda14e2ae728ee30eee5423d11c6a9f8337b83ec5dcd7e
zb2ffeaababea6b0591522d2be03b12aa561b97e53fecb3c4e52b0ad85631adeb6a6cc2b9333e89
z799f82a9ba18c2f15e6456617354dbe7676ebf6485621d1730db15649c9ef4c621b022513d76d2
z8551cd1cbe190eaef065ed32b8d40443d3a7d48fea2150c866a4109ed8401bf15dd4003a747f90
z173c1cea8e0df631cea388f76a585e26a20f620de1c93eb4efb2a98cd84a674cadd7833b024ce3
z64d04fc60bb4859083ef02e586406580764edd6ba841e7306ef499bb56c075098beb1e0ae5fc17
z0ee70b0bf339ab02021677f99d4f386c659c3fa6c23e89936772a0d1e7d0884d6e88ca54b076bb
z207414a76c6bfeb9e4e5617ede2a72e6a121b53d72c05341a65e64a4e9f78516264c0def236337
z96dc5eab8c32feb636bb115e1a26edabe9b6cd4a24a125e2801cd2f4ee27e8f169ab07b5cadb3b
z32f9e8d70e118484d05cb4847fe504fb0ed8f2c937c024b62f2a7bb03243ba82139de621626e37
z7c0d73b388cca323b6c38548f48c5937004564b07de19493ea7d845be211f119c59a85370656fd
z8a8db4a4c26ea37566b9a0284bf71dc111520d3dabb6dc11947ec87b530f1fdaaa3923d7ed4fbf
zd2a85564ac6264380d51f8ef1978d890f5f15073d718e06b5d76c39938e740938f3609066ffcdb
z8897ef5df4fc8d0e1a69729136f4a4e12ceea9c1fa3b1bd4a5de8c4e2d0bc7590083b60586cb71
z2ed4345935e7cabb9f623c08cfdab3c41c974ff04b10ba2d7024b6cc3b6b223db52a975cc337d3
z9b7eb488840ea1dafd6e7d2348732b0a42d5bd6989df5fee51923cd982709ef7a009000ea0b656
z55c9fb046ce2ae423c56f72523d14fe0a46e543bd13e6d56d26f29724fa1fb5beafd3e4e9189eb
z22135e6ac38bb4168102363565eebb4bdf690e2a0dcd2b0a544728b68ef702df0355a7d439867a
z8779c9781ec78f71763d06e57a9f845106cb013a9c671cc53bead1856f78d5d8e87e56fe6cd425
z7cd3f40f273bd78031a612adf19aeaa793167601a4552d3783a1e519e57b4a67f47828cc085e90
z5955509c21dc7b18d6781a5d22593f9f10827566c416f8cda043caca9a88788dd8661bc0e0501f
za2ce3a8568b5731f37e294d06c00158ee8cce0c2728b4f6d3aa95dbe7cc7b04badcafc636d28fc
zc70bfbbf8d673eb4794293d1eec430b21e036a9fdff270754e4e3ee95ec8327eb477ee5882cc87
z9a2889ae6447e4a6343c2135c8564638f2ea5d35f529deec9265543588ea6da6f92b25fb38d4de
za2302fc453636ddeb1f68058a88a3b1d0638b11d3a966eba27614b8b853f336d07211d2a3b5ccb
z179266e52b9d84ec714477b3f0c7bcc80506b95a1b2c8366e1965bcec99c9606ea58de01473e24
z52906ddf1034916d6c484a42c311764c7d5a7fc102a3fec36a6a7bde4521238e5025f36582888c
zb5e656a8e9a85cedbad1ad27562c445b068e754e107ac987b408a41342ba40818106922122ff2a
z2379d05c1b0e214fb0a99ee89493ad5244c7dbaad9d4f12d86aeeadb4ea68f651f9587ff6487da
ze7f4c24ae1dafba6fba9ece0c47e63174073b4df0f1bf87af37204701b6575951b237630ed3847
z4650b3c7719bf0663b8f2daccfb2ddd9f70170d8e27ca6b455a56014af72b9ffa58a9c274401c8
z8691a6d5866d306aedd3de62bee2be7117bcfe5d7978305699c636d02185d6bc6cdaecc0c26aa3
z334cbf42cf5f461c9ad49dc9cfa50bdd634fba088ba147ed50c4b2ad583c8b0c94cca5f0d7942b
z994aa10ec0a1b1a59c51977234bbab5618f754a942ce3db260e838016eb96ab5cb3893960c29b9
z3264bc379b418b0476c8200530d219f38e0179e257ea495fa357e536d5f6f65bde0f09ba082b7a
z83eb2424986214fc632979464179d12b36bf16ee94a9055829b56625806ea6fb99b5b4c44cf6b5
z74caad454fc2ba2307289c0f9c078081b86a377df13c1d7550f15f81d8b922a0d5bbb4e727bcf2
z651cddb2e187f2e95277646d099c535756f1cf86cd79693bd4564350d3bde55833183ad8830340
z38f2be0f071e86f2dac541d5c38d6ee274b5bd57e83dee2aa03388475535c3f6f8b8a2914be2d4
z4d97e76518439862906ce0af7dc7ad54eeb4294fa6e2618afe5f234479f036cef1f8b093735cc0
z0e64ea3da7bd858e25381d4df28d728ff1942bac147edb806b637783fa1970e633737430176fa2
z0c8917d5cd9430eb7f85d026f78f464de3048658e09d12d4edb039967c27b73408d1ec986e9c60
z838106065eb9f04f4e50876c5eb1cfaf46b00c0d648701aa4994e5584f3ceaa97762529660bcc2
z7d8dd3c733399fbb9004fcb6dcb88a98ea6a9675f70a3552ce415edcbd0cb705b8c1cc72924855
zf0239b152c6e12f03385a262eb9d60e6d5eaeb524b95ad203ab9dea54840b939ce2ce8d6b19a15
z76a60fed973a4c6b50891441ff514002882549e661ce681d4d8628468985f98a6c3f3f41990817
z57af3e5af0caaf13628b6d78c9a71dc5caae2e4ba552ed7d0aaf6a1d99552175488ca043551a66
zb3e8bd171243061ab405392388bce11b7b1c06110536c17ffb40c8b41fcfb4eccd4db0479b6b86
zb74f9c02466f0734cfc64feda502bd6a955ff882312bd6eccad44fd3bcbae1e71f01b52ecd649c
z211ca382b3aafb996ad7fd056bf401a3b63b309d855804c67de4d17aebdc1d6ce79efc6ea7c0f0
z98816b5970687c433125af9e2ce91fb24f7144dce9ca2e1bfe0b940dfac784e83432019f028659
z6d649c8142e054af49f0df3c82f4d49cd3655ab84b4632b291eb45660d9930f641b5f7b38f3d44
z898ad3cd956540183bd55b6a9e44fca1a93a524f8b1e52cca1ee8038c9e502f410ba5c02bfe568
zcd2e22f07b97b532a7b0cb19b64a54b76b16aa70fb7a36274456db154763a345656c8b5e451091
zff7468e7339846daa9e58bc7f22aca343a4b59b31541186a583e9a715cf9f9bc262a4e172600eb
z5ed1f081097c8aad6140694acd6fadb89685502a445198c2c0f5d9f93bed38bd4e888d8eec195f
z6748bc016dab1b0a1585fc876d8349731060e56dabb42739be13219c4bd26a6f5fafb0085260ef
zfddc775d1c0781909264f75f916e21d57da41143a78ae2d3f7c572b7e942aa161d41da6d7cc3f1
zebbb46ebd6f1784667b49cc2b210668f2040fe9ce8e552e6e9a6da3d11d59aebf1d1af70029c0b
zea42eddae1e14293b11a24c4f7ba6441bdca84ee3044a1b536dcc53107c5a5d9d5050e459f9834
zcddb23d036c6eb534fb221b244630887bb9c32d01a656c3850d8b29fc4f5d1ccdafa6a4bb81fca
za0bc2d0435d3d4e69ba8fe11a866701cafc648021332479613a7c1c1bc159ae5bb366a7cdfd395
z1469ee59406173c205600c905d85bf364e301da5619ab0a00001b6b0a8a3b0ee25ae8b8cfdba7b
zbecfa68e21b43f0910d3c781063f5463edff7167d0ab690d7e36898a07aad8cab1747f6bd86af7
zb36f6bc9e618a5065104cc8cf005d362d407f4dd999831ea5325fb4dca2382b262fa39ad20a823
ze1e83ebc1fd2de91cd64599314921afb921e25e4a647361168b655e0c5d976893e2aa37531d95f
z7c23d3576ad266ed1d9ede948554e51e62319de6432684746198b6ffb8d8ba454b480671e2ef11
z049374e3a93638e1a9475536e0c6fcdd824c188100655a67d9820b0a6d1060d7feecf717ee229c
zbe9cf92a4b4d0c105a4c2d365c3066e3b90b3865001dff3574ad01fa23282cac83b62b236cd75d
z714f549f5a51c3e19013e9233f6169a29da3b15d4a48db2c4d95957f7a2cd05d8aed111b4c612a
z8bdd0a2c8f873e05ce8791eccd756f7e885821f1797a1593ce00877d7a07bab9129fa63ca672b8
z964b16403bd78b69c480e77de39ce8f5e0af6b37d4b0a97d868bc4bf9564a9055beecc5a3115d3
zc7272d94f29d424f8095f48fe01a898ef7f93baeb1fa4554fe7db0d9948073fe0bbb4ed7eb5fba
zbc0afe56fcd2904d8a5a9ebce87e20beb680417a70b3d8a6269851e768034d6b3ff5606987f7a8
zc6fb1ff299008291620750a50b93dc5fe96ecbb24c5ff2973122a3792782ad5ed76b41e848fe68
z3fd3281cdd93fdf4481e955a75975f4f803cf5e69fdceb6b993a499a7fcd9a1bc2a398e59de781
zc933f5c410479360025e73084a4bb314f4e44bca7f079b84b0a747ae447ce923c0d23bf62db283
z36f44ecb1677b71a76551a88a578ca9e69a96f90a54874f85ca06d84daef8ef33230694a6632da
z85516396a791656bf26d676ed71a57bc53172c38ecd0aeb819e2d826d9101adc5fd63241b17ed7
z9e683153598c6017a212f6bb268c76eb6d7563568c3d1dc4e4a420b7a7edacb4c27e8487228fa2
z5d0ccd8e97434b4983b5cf4a0130932f25f039d1fe90744a0bb077c058f02b8e591f4cc32a9c5a
zc91cd49d375a5cce3c4c68cf5bfc44db0bc7afd54c8f622497034e3931dba154889562d5c0d1cd
z6c785c4d127b5159d4ffe81611f9025493dc824a08acbba012c678b52f116e22af4e5f473416fa
z31977a2a0b07b2a4c124c3546c593d828fe1286a16475d1bc3dd9e9753949ed7516ecddad40b96
z92c1638e897c29ec32253566a3fd72e6f6d1c4d685ef2bc0a87dd56faf7d5893c2bf6d50789dac
z18d767d594b5b4b4d07fe53de632ef5f17c23d737e528de522e74c75f9a4f40861760a44fb71e7
z5a9445a12c0c61458172ff3a23aeaede36ad2f072512e7b7c1fafa2d6de05f04c756f9f59b3971
z10213e01cf6f67c464d502a7a0f84559f31d88d40e779d433a344eef22d467361675b5d8b16538
z13a6455b3b54a765692ffade43fbc98f0886fa1af80e06a4c602751879458356daae6b09928bb2
zdaade44a8a32d37e785c6c8621dc549a8f68929c02143ef12429133eb0c369fc0a98333eec15c3
z11b86899231f10b5c4d2b2a16f964ceaead8522cb916a0783f1d1061593070017da14674b07899
z077b58c2b024eb530c34caf5403a955479dfde206763fe12e35e8293c80dc60926a3db2ca3eb94
z68a21c6b585313e7781ba8e5cfecf83f18df10f68b427b68ce142113f73663b0c168581d0154e8
z4c22c40d057a55cd92661540c0cc806c6955b533ffef6fbb31c5a31f199846a786a698d0a41ac5
z22390cfda5f8976c82149fb9a7e026a2b0af9962948c9c8a22b17faccc9c9af68db215b1b9a7e2
za11818b5c7f56cc7ee3478f5cdba1f6ae02e7bbc29dcb45dc6a9b7efb4bff2812b907d2e4637bd
ze659e40eb41870976d810a0696e026fb60625c9e315cd84050bc56258da0e9f19c7475ed3a1e81
z0afa49ff65fc6d5352097d55988a5bc94bd10ee022051016c94bdd21017cfcd517a0d94302096a
z37d82dbbb774bf249cb7d2c3ee9096559070861ad34667c11a41a7ac30102dd531ba67246ba120
z5eed704ec34d1f571c0c62bafd75d4dce556f1b523c56c0eca4991a3af542ae4abc6b0425c17e4
zbbccef1711495fbd40d48f2ba2ceb6b2f5dff637d53258f9666351ea2c3ea9a26f15ce0d70b6f7
z14a5896aacb0072a504e916f7792cc7d1e32111feca5a383b84f1345940bac37ae69f1eaf5acac
z827a61a8015c091ddb8f0303ea1e5f9edb09274a6a4770d14cc5e5d24eba5ecec19f04b6df5102
z6fe4f1f69d3875ff610ba6acb1eb474f9fdeb12f8439c842ee59a795341f7e5dbfacf3a10a0203
z47596828d14a9f2770c44377e5dd9fd735d1b7a4941c6a13b45709304a1c9bd31da5108b3efa49
z6765e0bd7d524450fe0eb76d421ea695f11d9a5cf207658f5bf8ec2aac76196d41cc04d8e7b1e6
z60af031784d017c9465dfa2df03c124b76397ba4f1dee5dc9f878d9584e74b6bb932f2ed9e6d25
z3762c9e01da4ce1432f165c6a00ef30193d555588ac76866f13f4c6ea55799fca6afa8329e545f
z66cb8e4af8594fabaedc7e0c4e7bf92e986f6afd7a292d8f14879755b08175b521beccda260b22
z0cc1dcfe7bf84b0fd6be5850e4adfac4871de850b3a7048236f8a27a3429f7659530d2167b6e04
z9dcc7d690b49cf84f862b91254dd91d5473b0b28a94b79aaabb6d59fee8cac9c55424922e3f14c
z382f85e9fc5677a0e3e03be18b4d233539672299cef8f397527b9269e843cbb2b9ac22a9cd8bd2
zb8c848d948a513c9471ad7bf555f5a7af30cd27860ad6670f083002567541ef0482d372c6f0171
zf26999b4532392e580d0e7223e1ccc5480ab69359159db1863b0e6ee767f1a9bad52a99cb5aaa1
z859c799ffb193327689a28b2a3ffb414718612f9f9ceddf8838b8033778bec2380f5084e3626b1
zbdfabd892746dc74820bdaf44846a2067ffdda69a7054d7a0e7523056cd9a36c69c3ad60035dcd
zd97d83bc3622b9eda8132486b05f77558944dc4515e0838c79f01ea146ba0844dd22c4cebc067c
z283b0daa5b0eb789fe23e046169bb1023b198a8c2653e7972c5771b1fe18953ae4de1eea1257c1
zace43138393caa7baf5b9e9e6ac80b1932f6b940535ab20df566c9214b6cf2c1aea6b22cd5fa84
ze51bbe272fb0b045965c28bc11f8660b0ab363e703693c098d030d40a41e7179463a70a4da19df
z9e352e00841b9b68b87142a1a870deb006be8cb6979c65677af7d620ebf11afff0f819e09ebd83
zedce10422ee1792c58901cb126a354f34d42894f9c99aa03c80aa13e44c36796ad79f9528fee28
z9e73d7e7c83469a9e1808a901f198596b2fa86a7cff0cfdd409a61bf3161e467ba23b572998153
zd3847ba70cdd6905e50a4e6a81f877c2af7c217cbc0ccf90c0b26923280b09ff2a9ea57dcc4bae
z6b79bc590f267aba51ad2c6a015f595e7b82f53d555426bf85d4cac4379fefe9b1b346b25fb429
z880e80ee46bda2694ef4db8557421e6ae9be7440ad7f096479e9ca82ea8870982ebb6cb06a394a
z8b41067d7265270d09fd569b7f9d52c27a36ac1e9993d6046e56b531bd63623d711e255242b53e
z92174280f665aae9e6ad570a4b31790e33c1c3cd0568ed9ad9619687dac8e7a7a31b7ec6e99047
z9b028ed8a4b380307a881fd4b71fb9d26ea4fa534c16c6f1167f47b49e1429973dbe36eee60163
z10af67ecdf76014c1c30bb5cd074068fe70c0121a6bb721b2777b52b5b4c1cc43f93eae26d0692
z01130f179590c0eeea56315fa2927570b1f3eabd822b18af71de8a8d6b8d1ec69387d730cda8a3
z67e4a3c1f6e1fad6665d0443f21cb42c3925bc02744a201728183bf2ca4e53cb891f873335c568
z07c210916dc75ced7a1c8221d1889e39f992eb67809631a1420cff6c4a717b2619debc9b98711b
z6e2836294f948dbdd8f719b5d5014f19444863205f4c7efe0acb2bba5cb122543f647032e6e869
z4d854aec276995be8d73569a958038fafb00c027fd3d4b97820164f9662d74da8bb9417c897c5a
zce7dd8ce5a9376e3af145355b4d68483fbb8f850c5b11c6ec4384c2c67fbe9a11412ee0c4aadf3
z85ff8adcdd597b5108e4f474cb818f057038462f07a4a4375bfa0212075ab01bcea5be6f7ae2db
z6dd6ccc5fbd8608236bee49257016d39d43147f52f15a7e835db763548ae0bfa6e661610cbdb5a
zf9c4224bbdf210ffa9989deb39b78e71a5e11b02edfb3afceabe3e145923f6eb416adf9ad3aa05
zad6b2891d2d5f792cbd830991229912091cfe0dbe689380ca52e8daea8e4786a09c0c821bfa94c
zee4918724deffacf79a49f8ad2efc23ef6cc861815c53711576fb48e6835dd28c1b5fe6668d031
z36286503fe4bf2a4745f3abca1b7751ae4928de7da4ad4b599adbc04ac4f342342713edfe984de
z9908bdb27d634b404512bc7b92342c4bc95c9cb85e2d069a855a7a8ae5a09eccee9c52caee99d5
z1e56daf0b7c5e63b2bf8cd06b1f716b8685f18b404bfac8bafa408c9403946c875fcf443cf63d9
z96543fc8d4e3bf1ac3d10649d294664bb98cc04c0ba119a6a757393765eb0dfec4a294f6b9df5e
z490da7f745e08fed3b9818dcfa1d834146cff10201026b5d3881c1f356f1a71377804561d98072
zc2cb0cdf9265bdf19d4e2e4226c02f46e6fe5f58ca233103e5bb87972feaaa7b2675b70c2e5e42
z9c676b7740767568521adc4e547247603c4a0556f7f1049bb28025cdb221a2d7278d44fcf43678
z63bcb691fb4a7b59711ced90a9b014c24f7bfd5ea3fedb847e5b4deb9b130cfba8a71d8b9b21fe
z64769e4ca6acc75c72a92cf0dbd7f77d3c9f4ee5a0173042090d6c8b1bc6393a79828f09936184
za212e41e51228ddf187ca0afa95c999f7ff4b2bbd41b2a45c1345efb2665aa1af5e58fd978a94a
z41643a1bc99ebc16ad657cd4332a84d3b0404ad0ee88271bfc391a00225c388b67603e4eb8b8cc
zd327865c66376f981cf8163ea0147f50c8f4155c61f029010eb2adc84b8ad95b8ce232645c0240
z0304e558f0ba49bc96a56b2292949953b6564b49f4cfd7e1155ec6349e52d60302de8494e8e13d
z2edac19de5f73f3616bba86843f23c17e2ebf44eaa43c72dc4ea6c634792bbb31449dbc590035b
ze02d5b64e0f9d30595f995bf02e435522816c9cbf8bd25383911d548ce67cefae82b286e93db1f
zf78680e7ad117cfcbe8d682d2565e5b8d979b4abe2e5a2f9f58890d3d2529506c7e3a69734a2fa
z71e740514272aa76e5901cfdf5dcbaae719887ff05c0e146f98f3fa234dfcd65557a49a2b1fa47
zbb961e26f8152e8879f6293ddb7799cadd5078b054a0d7d55f362bb6c72eb237854418ad7d0774
z8f48453ca647a2b0726b3336d497d56f5ac57f39b7fd84c8cf942cd867c304bf850b770ef34cb2
z6269743a7d9d3ef9ddc638ec5a75c3a2503c653e0581693cf84e79cf4622492bf6ce1c41aca2dd
z312f5ed4df9b4a28f89e2fda7dfdd39b5c04706c834cafa537f3f3fc00a7d0ee2efd62de490466
z2c7439d11342150d28469142b7c472915b01a5ec24ee218b6b97e55934fb6224e82c5c26a4cd08
ze66182462ec537ba6689bc9beb818332fb9510d2a72de913f9364240177537227bfea4cab7bc17
zd4ca0845b4df7c68de0130222690931d8104d61525b5560b669a2d148f405ec6ec89a4c8f112f6
z9858f0ccf7506e953aded19b010d9b5e4c0de48bee0c89c55013eeba7995b89a69d5e0522a3703
z2a68f33935a576c74102b29b2abf927201f2c8766a9219c42dd73f9dcce7d36abd4025b58cef2b
za2c75449bdf2f6978462f72d37e3aa5fa2c184d754e55357dae174e535e092c46423f83f8d07aa
zc3895382c176869b97ca0282301b008144bc5b89d2c63cb4fba31ddd87e75fff4df1cd7ac6081c
z71f5b42bc7b28ae732e609d212f6df0ce10cb136efbed826f00e9c46ce495f6362116439fe3e5f
zf1c38f9db430a0d9a20a62b416232a5b61507683d98ea861f26a276d94426e9b1ec7d0f8cec089
z257339f6b680c035308895cc94192727e1a9ee36bcdd3dc7d533a5809b1feefe4465f8046ad33f
ze6159cdc3acc7f98de69b56d2dd4530efdd1c6073b41a7f014b3a842b850ad3e6aa108d5ce23d3
z98d13c9febcb8b404e185b19b93e4fa67f9540a27719c2010af117e0c8eb5c49486f56c937d14e
zced11d4c20a2a550d644a208df955b901ccc07772b5147772b3e8fc6b07bd3ae4f6a299573db12
z19d44c416ca7b17add8166679f91e87d9c0f7e29cc5f583dca86435d6bf90deac1c39064f8def0
zb9dc0b1a355d1c57f82961c9e3d0160ecdad94f3f0bccad963c53678d3fcf882ef93e16d0ffb8c
z40808c33920d076792971151f30ca7bb43fb60c81e344798b36bf8edc39ebc462baa3f869a0f67
z9b7884379d2c173c643bb80dab588b3b7f195d9025923a73f7789a0f6cd1a39618c75801213b4f
za97eb874189ff824653ff21c28fc48a0f973392b83bff9fa6aa52907e63592a92174738d3f99b1
z2c42dd2aa46881a563ac50e217c9d10160ade46032ee897bab5a4c4aaf6b2de1501132b5577355
z26f65a7f8a40fdc42e71512f2e1993b5d3e56edba7e0715a337e3f226c3ffd04e875fe2b473835
z4dc4e7e9670c00ab3f1003b7c12130a5466cc1f2a7c2f9b66b06393a2fde776b240f90d044875a
za8f9acf224965a5eab063bacae14eca43f995dd283cf961c78194d48ac1ca056e1b2fae987629f
z5e8453a223d5fc6d2d9c73bd61f5848848df91523b23cc80154d8a0b097926c16ba2fb8e7f843b
z0d6ac431e530bf51a0816ec1c10b4adae71f2760f1408f3fa5d2e264030ae977504d9ce21e7979
z020b91402669864dee50005abe5e92d87e584f0bc04e73d10f9b0e6b026c803c973f76862a513f
z4c0afdcc5785c854c820b07786ba5f6d011d844a6bcaa08813fbbb37947ce52745f981ce40087f
z75e8f301d1369b369e44fa29c21e22f7c03a3229c90c7d8a561394d07d4b93c0f16445a71025cc
z7f50621a7b1b832e7f5fdd76882a5a393ddbc1398f4611a222798f0e87de97c7a3a263271219b8
zf043509b13b1f2d4b36888f98c162596c6bd2227a27c2de8e12123ab6974c6eaa6f558ac3e41c3
z0128203a786a6f003ac076916fa6fc2bad8c61e331be08d38d8064116a493d4327eb4cb93e6340
zd5936d3365289f8a262a26c17811aa12fd1e58eaa80a816786bd76a269608a4cc4ff0073d875b2
z0113fba252fde852960a7c4445b0a8a276e4cb001e1b0f4db4051af28d1f848ec21a399d18a8d0
z44cf7bd31b7936c6179e2f6d66d3a899bc88733c23abeb55332b21a998df70c81bb12ffe038ee1
z0f33e784a45795dfed15ddcfcb1307d64c134e7bcf6cd61fc84ec3a985b0e81655e2baccab7627
zedc8a9fa7bbd644b5479452236538c256c35af03ce0de3420ca24e450abc8a193e41db114cd3df
zd22d096a0eab1af80795c8ccbe0f7de140260dff76d4a6486ac87de31ae3d65ed9317200c5d3dc
z3664fc53c5b3d7d55271b696e1c147b19e9f80e575fe0c2dee066674bfcbe565ac5277064348ee
zfc542401fd7c151212e310a01db2a1b96bb7bf944d0767d7862451b8799770e9a903ad326c670a
z21d6a0632662f59f1c884e50ab15df96038589302c88662b8af23089679589bbb1293ac83471e4
zc9855bb14e4850723eaf15f844d99055508cdb2a34cedf846a811c6137d339549e260462a60f87
z2f9cc5b535bfb8db55ab12dd5341b345b4bee6a2cd151586430976ee1c4732fc354d5e0ee7f3f8
z5a3ab77565e3a4b619509b0035f368879d2f2ff4444d2b63c688c938f7ce51c3172b10ee4cf2eb
z4c0a4ad676bb3f8b75666200d4fbcf67889fc0d9c6afb6ec52161349b5b11c83e6e393919f8bbe
z1fe826c366a86bb4cf2657e1f1e4454dddd9c940a93b648ef14bfc6091f08e7d6db54a0fc13feb
z6ae99a96cd802b16d6123b04e46c99d7c25e2dd3d407706d41117b8bbebc0212037f83d7a4c6a3
zdd480fb5d4433daa84e34446fa0bcd2ce11a36415cdf9a39fd51b61491e76f5528010f3a688101
zdbe672efe4d1ac6e3004dd510a436409946fe41e14832017a3f395330f0224683efa90417249d5
zc2dcd290af6e3701677b250b7a6f9d4b388acb6415e1346820588ee35a6e8a7dd480eff7db0cc4
z8250c08b54c98f5561b1480a61b03fc7ba2352b12e74621bab1462f4daa316ee0a763e256b9752
z8c4c29cc57201955236759940b7a5746855f813e884862154a5d4355fcd9a902e7439bc7ae0275
z7b4ac5f0d08e2a1cecd84fb5670c29cab829243bd3864175583c8d3df8ad9df59f6a684bbbb8e7
z053a0671e67c89b2bd6bb9cdc1b5ea0d18f7fbac42e1aaa751d2e7ed7f0b4d3043cb4558b5affc
za90bfed05f98eede499371db1c3a661e50b2cb946b4e3e30e79e1a837ca03dca1182a2140e4b6e
zd5a1d0fecbc3fd17c062a13bc0deae6d76f6f08974498ce1921790938b54c46287648eda53e810
z874c4c3b98dbca8dc9b59ff2f589bc3a8fe256dfb3f024112280b2bf6d9e5f8c02b2f8d4a13bf7
z96842f57810aa568fe0ffdb07068b8162bbdf8d91bf3415fde1cbd746e4cfb6fd181cba07ceba6
z0a896db23c8053ba96c8b403a51efaba1691ad998295b0a489fae061175d9b99ab553f0dcb6def
z923a035ce7621712e8cb93c8ed2f8cafb5e6391e85063d42cc8c4845972263e661c2c80113827d
z72078ef33ff76a790299d380b1751174f8f1323fa1477946713744d4210cfd8c62eb00d13e25bb
z943b77e8149ca9142e3630ac0813d78c382cb0fc1960b42fd5eb1df87b663fe7cac240bf80ad30
zee04b63ad3a75c1a656b6057e15df6d6e627f855f1bee7bc140fd3bb933691f57a94495ae54568
z150751a70f457ea8b512c4791bd54f797843a10830ec499b9d9add74b166ff3f26940dfa7288a4
z7fc1121c4a5d26e4f2d47c75b5726a15b4153124b4e3ec9cc19668a21b33c00584b3610578e5e2
z28611695e5872954638a43da4ffe097ee939b908148ee9e3891ec39f8e1c2d52e7ab250eddf7c5
ze979808bf6b69d1f837f864263f3e060d1f4b258aa64cd4a206179d439ad314cec757be683b042
z70d656e7e2e5470fd51720f8b179c8b0732264eb7894b9f75df38b15716fd13c53fe1f70e7defa
z691ec4725d4545c368d7da4a0573d74b30f8c89800a583b0b673612fc0c4873189a4429d186feb
z0f03494e1defdc9bf891ccef955c03d655f4aa5e8cdd38058e2499416239d6bb020497a244673a
zdf9c16c8c9c4b5b636cb376e6388e567280f4076186b783b459be82d9682aaf1c8d34ee356b2fa
zca037618d608a67dafda99f2ffc19285a95c07f0c954ea8fd5cc7a88995712a60b4c891bef8baa
zafa8e0c5b1a10d5d9d303655aed7f772322d9aa414d92aea2380b326c2048e8cc33639778bf4d5
zec1ba37958069a589bc37c6a36b846705190ec30a07dd705fc2e6607aff4c3ad0b908d81750135
z0467337436a8b1eaff47475810407579238f9c67805c8b022cc479b4520f9d8149cfed47d9eba7
zcc334d77a730c30a69300dda6390b16adbc128c9d65d37b1db30b1dd10d3a3651aa546cbdd28cd
z4a4b5d7b04de67e09d33df955d85c07a6cd508658d9a7a820c92ed28549c034487260d96f86f6b
zd4ea10ce9e4b80d4b08ac5f29846c8db06582f45648dbddf6d1e8fa20eaecfc0eabfd3d7cb9d69
z26130be9e1ed93d6b51c0681d2f34b45f3b3c6990d1c7374610af30e38c37a66bd315aa1e071ae
z805d3002515f56a05d5f815698fcaaf534ffdc5611310cee36d1e28e322e2cae12252a4cd61ec0
za711962ea81709351a184980ef62844a8e7968ed331cb7ca3ee4f1c5ba9799da44121be357cd9e
z09e09f56312e60f099181ef4800a33068482724c49aaab68c70f1874f77d39a46cdf122905cf28
z48585e70498f7b3c00f9328bbafbc5acc7e20821cdff505f58ff765669b3dd8d368892388adea8
z73097285c1397c851ae4ec61a2fd22f681f14590e6f11887c0a8a9d887a602d3b8d6f1c54b2a89
zcf5b4a6dfd27ed43969aa9908e5b82a00542c0b90b44b087818f4a04a3a7b33ec00e15c902f5ac
z830f95edff826101a99c250a4beaed1cbde09708d80969006f1b9f4ab555f79b9e22c95e631748
z156511190903c1f222f6c5de4b827bcee59cd20813898edaf52e12711d533c5f45ddb054aa66c0
z0fd0c5df2d0f27407631a6c84d96863c91138e468baf7ebc5684446e8f34a460f2a5c29c255be6
z94bf66a29ccf559a211f43cdcaded7de97b619f32b21c7f80fbb182ad022fdd82a590626f28899
zaecbd8bf3608655ead2e7d62eb17d03fb3d5bf0913b2e4bebf17ef9744bd826f68cae0baaf48b0
z5e2ea1054ece749c537e5fd62fc7f1a07e940d93f83f25336fbc277b309138971a3d5f722fa62a
zf203469a676a86c4bbf846fb2f3b9feefe3b06fdbf73a609ba33713e36033f751fcee625ed10ce
z3e64223c6bec158724e4c974eaa1eac8ce40003c8899ceac9e9b15223e3ad6fc909ea37786a1ce
z66ce1c8e42d63f968571c185f194274488ff6484263f0b6f2ad52defafb3c4f94df249ba982dbd
zc91623c69abfd97c36ca5c72cf3be199e312e2266e664cf470468b845acd483560acfc64f90224
zf56f7eeb442751d9b72e0e00715dbdbd58bbc765fcd38db19d31225f585ba56a98ec687ad80b04
zec5c867b94eb5a443ac8063e7b0e286315feaa1fc7205519c7d050467d5746516e8de608d4e697
z9703c303b5005e07c6467e564836b8b637bc1f512bd67ed421e4a7065dd54d81e5e09080cae27d
z5490931342c694c7aaeb5155e3b37a9abe7c1d96a001ca587d9718fea7d77e241bfc8f9523fed7
z87ae8414f8fde9cf2a73676782e225d7b161a74f9e790d8e9817d02b651f5413c0dd60987265d6
zd423e5f8c02f5e67eb13eb0052f62513d7cfe72f3e4aecfe3b21d2d56d486d5526a22a200e804b
z071e592cded70ffbe1dae6f2caedf49854bb55934e784aa7d7c78bf3e63e42fd66ec88daf77f07
zcda9fd89d06da8fe03b50cd39ab46e1b339510fcb77507dbcc12bbbe1ee4843843a9439dd9c98a
z7570d8fa87be740327739d34df109e0aa161b305da0cb563b4a656e083aa095dc8c640c2a25ce7
z30e9b12d447321a078185f532d1dd965923c646efd6997f44bd019db8528a8947216bcac35506c
zd1240d77cbc8b6e3059928fe1c39027b2b62745a24d3b5303c0f2ddc3a8198cb6f46b927fe9877
z96abadae727086136acf1cfbf236388ad84c8aeeac1cdb8a906a7ce1cc265bbab8dc3ebfcf6edd
z207dae437960628447ca97abe689b4636fffe46fbbbf522c538341aa91d39c4b688ef7ed2d8a28
zed894c086647e4ec87049dce8cd9107249c6a91b93b8076e0d116583770c1335afe0ab96dae284
z1ebe5b759b9eaa30f7fda2ceef7ce7172a4988f748b730aa06fabb83bf1e6655a69f17ba7736d1
z933a73c34b63a2aa4bfcbf1d88678cc5c8539c306ea74c1d51895cd259ba6328ad899fe4005711
zbd63d1d91dd6eb726ae3273099b70b2a9b83ae00c672663b436472d259f9e94c9ca35eee67d409
z0538368ac2237de0b19ee3933fd491786c8c775fc80f3bb217a56e51bfba5c77af9be1313287eb
z8d746cf5f8ee06b65188dde42ee883513e7af8bbf31b03556a7c69b50d60fd63bed106adc407c8
z43d86a3fbd9db2962a7bcbce2285987220b73f3bed1fab3e775ab442becebfc65d690969c574d5
zec625f2b5bc74e343ee52d130cb8f8db9733da1705bba74a450fd4dd50a1f4ba352c4728443c64
zde128db39bad3132ca30a176c7437857a888fb484e5bc5d00add82ac269c64594d04d8da9e5452
z2d39665c84ee0b985722dab33fda0a5630ba57358e09638f4c6805476bb786a4e313f1b159944a
z11138e4503aed009924df8499e60e9bcb1b2de834d5e2628e1488ec817776b5d964072e76e5988
zcf7d38151bceb84ca23216042f59d94674df64820ae6019772474ad7ae93026d5521b1d97dd7f5
z30091d592b8cfe7c0ec5af17c7444e9c08ea6b69a9f1a11c3548ddda749fe67d04b1467aa17347
za444c61d7e9eee37caabd796385b14ad43c96620396a4069b4fa2a55c0456e6d50caa7f365165b
z886e77ef26a3084556696490167ae849c52e16acec1a055342ae2913243b07535dc26e02f2efed
z046dfc44d2fb7880a5dfdf73fea458c083eefeaec39266413203284d57aff20feb95fc03a55adf
z437f094414d101a4615a2754d3b977221a167865a080fb8c5df4ad7a8663ec0fd2f3222a6e4f09
zd9bdb179133bb5302a7d887060e3904ad46502070873c1512a2dc8287174bc717e26802c7bca1f
z1a4914510440b927c39467fcc4892c09621012ea4a6528728bc284c2abad81a0a5c254747ed806
z8007c900b069b8fbd3ba576b645d6d111505fa417b5fff7d0b810e46d751a458d16e10dbe61375
z1f27d8d223b5b7e9c29e4e4a751a6f810f40afa7661acde5ada439d19928bd58e2a52d34b5bfb0
z323b552eb9140f9f0ddd4a80c0d5779d890db7788b45423b8cbc0bd722d2b8689616cd35278de0
z42702bea70199bc9454ff4662481a1012e40651e283353f7a7e48f761c0f0bdf5540e461127eba
zf8d907522cd92c34731980e03373cc900811d7e2cd9923ca5fc270b455bf6611af2a9d82236b82
z6ef7281e159b30e7a6ca38302aadc18197bc606ed89c3272420bb94d19d2f96d148e106e218a51
z5a79ead92a0d446da66502afeb333581fc970f161593ca6e4f6b932eb171d7ecbf6e3a56c74692
z0c9dc06dd8cdd875f55ab024c7561d0a00e5ca63435763ae0979b9596b716be021b463e4708309
z41b0dc24eeb0b1ab2f27827b07c5cbd38869f7956578e75d491dd2b17d62ade937101d1eef5b2c
z07b034d065582f0f0be9c2d3127f09548eed2df39d05807357d6356433d0f4256ac826aeaec2a0
z891c9aabbda63c666938a76e1bf8a652a6cdbab1bcff63606873db3a14f9423fcda7f9f8fee396
z734dc39bd38c22e0e57a8a285930da9e15ed830ec02c5816d8ef7ece98a56a8d867313df366acd
zb5e57b67182fa642e4bae9a397a3bf02ea166d5bc1db8936f63a05c81fbe4f6b9a5031f4983897
zb461af63419b81694a07f702b8346c74ae6702242d735c9ae23117a674d24dbb433f85f7626730
z0df7194d2d38dbe01dd74942cdf9546700a99d36af85bbaa12c53198ebbca4a2ff7e5493119733
zb9e1da3c9742a9a56b10423833248c6fc1a832e0fd7e91002979c3839585b8395bead32cb7b31a
zda80ca6da536bf5e175be3709bac4d9030b34dcca85a362e46742cfa1b007d4c58d26efb18259d
z7d1d1908307a7ad2e7bf8d4c5e105f18beceb97e5060e292bbfb39aedd00ee9a42f0852985fef9
zb8af07d4fafcab3d1876c114be81cc41f8b03a5efb00de15878a8520c1a21d6d99c035b13296c7
z61454178cd6552343b1d45d0a1a220570c9a9c9bf23a3deb4fd466fa6e13d3fbe4724fd7a73f17
zabcc564741e28e4a768c326d85cc1e41b2ca1115784c8bc11f652420501fb25f71dd0e6c0f4db4
z2a6418e1e3d6dc0a0ced8f50fbd4b14eb533eee134e29962166fb9405b4aa5da23864f15980be2
z2ac6d68ded0b36d83cab76ca6feb0380a7902fc1050ff5defeea17c164c055f6d0998ccc355a15
zcc63aebb19c4d884dafd4d816c92f8afdd3104c569669dc31e4765f219e5e3a9172608f896dee2
z87c1c5d9116d6f65f701f53de8867f8f2eaf307eed192c30375d763102a1e9a5aaeccb6074e513
zdf7ab856f5a2798851fbc069759dc85f0cbd9d1a020d52acc79e6b9b6a5eba1192fac07618e965
z916f667369095c835814fbddc70c5d2105dd0a65b937f783bdcdd028f03aaf8e80d4dd28b55cef
z52a98b69b8d5b433c8bada9260723a99860335eaf57bfa62c2b40306e3f3a80d0594e4c97268db
zccb3ea8a5cad75f97991db7d39edeefd3a5378837f83d4c07caae80451ab2b0a245d1e13b3a5d0
zb4d473a9a9e5b7cae1897e88e347357bc15b5725577c535f6f09d555b77bb20f8c045d85b2ae28
zbcd94c7930ea006ac6a3a6d7fd263b36106d756bb8194f441110b9a8ca0aef37ad16c71260f803
ze7be417f8079123be446549cb40dbe20a92d9c4b75bb878a841b86aceb4d52767ebbe1345b565b
zfee9d6a1844e2ee3e05d17f6b4950c41035ba7c710ce81f0683548727019242be0c4252236e887
zde67c338fb64ebda00d2c51a275fff9cd526fd6964b02b2c2cdcd0789579fc8fb2a7460faa8e7a
zacd2e615f246cedc71e82f697ce53488eded1b2cb74fd92072097ada180c41dce7e5abe7066afd
z53a64831eeb2e148f9f079d529d66e497921bc2998fc6cc082e53da43921d08238700df79edadb
z7ee1bad2fd1bb964c036dcbc4237cfa01e08985654391131fc4217b5f0ce8a5e15adc0ea5cca4b
z1191e4eee6ba5f88838a82beaa586fa035773e9d0adcf55155c93005627b1ea7472443fd34adff
zbf4d28688965cfcb75c2fd02f51499ec0c7e9ce88ef42b40ba9b8a26eb533dab21d214bf71b0f6
zd14eace360caffa7d632514b3ba010006ffd0ab3e51e132630017d999ea1fce1b4c5e66abe5f24
z05d5186444b78904ffe31b4112cbd0a72106277e902bceaa88ee46b1a0aa202b749f03ec02e265
z0ac371bce5561c4663da3df0c22090587294ce5041268e56e823e865ec73c928f8f409a84c91df
z776b99b511522ccd0ba39471d045b87cbaf898d68de938afe8dc46d8bfd6f4e18c1b898c75d9f7
z69b162f8c57e4c9558cf809d53aa238606688c503a7ecf9be868b1e41d19bdcbd61906543491c6
z72037b0bf5a355e5cf4de38731e81836063e4ebfac25655a0d854c76341019928325c8dabb4dcc
z563461485fb3f9ff8f8f5c072cb5ae2676342fd597345e27ca255b5086148cb8b780cb6545634f
z898830a75b497b5021231de65d0af6903774c2f84dff2e64f60316df3c2b782d71014459ce6cf7
zd43f8a3c626fa85bd250891a728084251e5180a4a1f84cec9ed6fae0020e266830ac811add07bc
za1bede723c35dffca212f47e3083e5f72628678771d4d6ac938c1f5d5af8269fc957f67744a841
z90b8f414d8c803096089681cb877fefc7fad7e17c703233d49fc29b045c65cc2fde313786c3b1f
z5d9feab64f7273106d9e19b4a2d49292ea0c00586e2bf7bd8193765107c8df893f7e741649eba1
zd3369a2b196fd12ea4a979cb331907ba2999e9669a7385c6f12e69187bc3e0aa83975be4ff2191
z8fc9ec9ba497bc8737a6de8096e7ecd2b007e421ae6d3facc4893ede1138435bd7b1fb7021499a
z2be5ab9ab42e3702f8bd59f11494cbe724808b791dbe48f737289ddd9332e57ea6519673f33290
z994d30dd73195328b0b0348971ff4c2e82f7da596936e429d87a2ab17c2181dcc5f08d97ce4279
zcfde6111ee3543bda14fd75087e86143ff42e71d697a8bc23272bbc3feec17c38defb985aa157b
zb5bffa0f2646350a95436551cb03719ce140c986cead9759bf6d70a0784502273819d11bed9db6
zcd42960bb4e45dccba4dc4266d056af77ada4795cdb846dd6c28280595ef8fcbe352035389bc15
z493782bfe0328fdcdd41489007e363f74dfe8f88582310c363a512f9757e798ba48ab0d2344291
z3ab687bbc2a686e0ab60b4f838923eef3a03aea01a8b39d293d536ed38cd9103f0e0e13f68005e
zc90a55d0231b36e83e93a38301a2e7df1da82d7398829b3d519b920149af31f85b591a54c119b8
z9bd32b64da2628563deac475929bf77fe424b52811165698c83fa8b3527840c1029e4e6c9deb1c
zcc1e97122a8968a1d31c089c020e0b11606bd5cd561d4d7ba6b30b29c87dfb11b4c5dc49ea4221
z4744bb069238a18e3c3a6c67f6e7648b0fd0640ddc07e57cbb2085d28dda64e2cb1b4f9ad621aa
z0e2945b5dde82716460f64822f25e50f22dc3bb0d675802390070dbcf3698b4636c2d59dfa6255
za8a5a2698140f3d12b1ae8bb0841b2f019042cc6312cff5c939bfcabb02b83bd4b5b197b1bc45c
z4ba450786bcf6458b1eb6101e5cc6c280e0b1e6705365d0466ddf0e220a29ea4d4720caa817d7d
zf23fe4d32e7cff6105ed98ff2740209577fede13ace0e46b6dde8b4a7219b86c7d55aa0a1c9fc5
z4ab6bc9f52d68cbea2b024e13b3e87d6cd906008c174c390ccbb42905750f7eaf3220c94772d11
z063a97d3a6d1ce59d28dff22ca4eaac465ce98ee6309ed9e5235b2869f74658f467630d25a666f
z2a973abef674d41e26b409c97f808f18c4d68e50be0e3340a5f2c343bbda229c9917b6ef991359
z71e63561996150423deaf48f3f3e6745667bcbb6088ed186af9d2e7743784add43bf2f2dd7be5e
z707b7655bf4f850829b609b593ef5215c86d993808824606cec7fced3c5cb564958c2094be4b7f
z8967205d506170bd94504002e4ec421181d9d850117cc4b0bda0f78521ac668af188c06b97744f
zbc3192cf3f34401e714a2c3b7a7a40be6e7ba5b990210c1f165cbfeb52cc4046f619d9506744f4
z51e8970ca612757ea278a204496d1701d3854c1868e7cae75947d7318b1783c880468e1c5f94c2
z339b06dc207f36f667ca80f6fde93b5bc12e0fe6b07f2c974627675d1a501677e950e952f6420c
za8d8749a4eb40eeef24c256e081083369f05fe92850b1849e1a67b3753f6c4807bb0e2bd534bdc
z5ea7532555671e92b978a118312f108071bd58a12c01ee5fa86755a5907387c5cfe99bc6067908
za3ba47c7cf978dac1840adf1281d0a64423212c8d71086d1fcde9e56a9371f9b79abcc7798c223
z065e384378997e9a70317e9eabe82e8e51106870948a3e51ac2373ff295c342f266b30c2431bcb
zbb931f6ecb7d2a281e30cc417868cc8b49cf9683ceaed75b11fa6c70883ec51bfa5d2446dddc6d
zc10a03bae8badc1e97b3b294ae074a4f530b92fdcb500d3a7fa31baa8d98c4cd15b55d7b0d1323
zb6da5bac8999279011ed22dc1ef67c5d60ec1be995c15ea0d9624dc8281badbecaea13b0e71273
zbb45bc6ea6f124e8ac2bfe9f4325d050867447659777cfc6a02bc0a6b37a607e53878b34c30065
z1826ddfb3ac383929a91c3d22533a4669abb1ad4885abc915dcda5147c06bb1fc73c0641c96014
z3cf971abd5d877a9cc89ba4028eca21f83d8a8163955608bc3d511d751fdfaa2537c6d507ce68b
zace3126d61602333515dfb22f5b5f62f7c02c3bfe70352191833adb0792726327af70860d67f56
za2f6ddbf42cd21b2ae8c8ad200e51f4c96579b4b759baf19ead8d5c537c2f5c8d04b8c79c867c4
z0d827b72beecdf227116b5ccf8918dbac3744973b3f2df25ed33d94c1bcc6cdd6ffd47be5c1607
z81b0a5c980bb1a0472b43b0bcc845add25ed15262edaa6f6308ea5ac5fe144458ba0c3a1cdfc62
zf4baf075c0e29c1be5f9071ecac9afc0d0df6da942162e9aa252c370540c338ba0cbb635f28bff
zeb18f16c0b3616938fc27e6ab4f895c622dca0502e52b197434be1c7cb609f93dd57a29811d402
z99d9aa122620a2200e3aefc1610c477adafdf71155f4776ca6d5e4a8175dcc0a4e8e2376a24011
zd8b371fc5ca6b61388949667a937e4d30af47e72ffede0cea74a8a12a3b155e23d742fd73393dc
zf8337158661d4013df687eafd1cb5447e699cc22a081a56e817e83ab1086b73265ae8d2cc829fe
z4a87f9f126b870877707a1e21f88e1d35ed1907a01f9954601e573ab0ec11096859bf554728546
z99a7263759c0b2e508ef11354a6e9e7b20e94cfaf276ecb85126c5ab50c10c20ee3f63c2a5930b
zcc6e6aa665b85ee95b097015b24f70cd8cb9fcbac27940709c6351314a15ad0e8275472f205aa4
zee769e6ce8947659bffbcd3ffcca3cb835a534b06cb74439b027cb744076d68368b0443c3ac7fd
z94f927df38669cc90ccd01f6c2593988c5197d71ef2948e87aedd9d06b86dc1388ace8b25cebac
z6ba269720abf42199da6bd4389112102735904034c4344a2a7e19bfeb04d41f419c3adcd9ca554
z411a8459e0b42b5f6d8a19f88d16902cf22d1bf69d46b1eae901c540afda5319e615399b376e85
zaad2d54b7f9d5c9e232bf69038dc31ae17295c4675dc611f74456639fc1f01a652e64c52caf78b
z6efd810457a30c36e5fb7b97b9949e695d09fba92af16ed89783edba61f111075ef365eecd11d0
zdf673daf8a08186b053057909dac586403d82d0cdb40c24d3c1cea7061660c4cbab2416f6d453f
z528de8ebb3b3622b141dc41c93a2bf59857f40b4968bc884253f2c7c7ba35cd5660b88541cc222
zd23c22af4fdf9c1e02d3bff51bb5bf2394a6044b09fbc14bb1d1c1153659a35d9454c67a2ea648
zaaf08cd983a26a8e9454025a1b056bda449a8b05b747a98a41b847c5e71b206e0fb6f3fc5f54e4
zac0b83e5e3bf00d4872c27f450428b48a2c46d5123cae192a1a3e8dd7d33b983c5d20093ffefa9
z69c42fd04e10cf1bd4688b59bdb5f114898132914e2bec89fee8b0552930dd4635227e5e57b8e5
za943b271674c3675ef703c6dbad73af685fcc13dd0eff4bf6b36bd6ab4d7ae29c008db6d8713b0
z1bcd8da8f5a0f2dfab41ca0c65edb1c663d9a7dee12c146dfe8bfa75008de4d06abae4103df12c
z86ce882ac1ef76d363984d88d953e0e937b531c34dfd437a30ac375ba69cd7dbda2a79e6ce3039
z59d58ccdceda925f110f2a297151127ebab34ca1f847e7082f58dde2916b5dce05f1320c795e8a
zf6d614a7198d0776346de9402d52ec6907ebc9bfa1d3fe286c6a6f1a224efc32b30af42d86005d
z60d4e742210ab30bdec033f37d9604487dc996bdc6b6f12ad516dbd7f3b8febba01467b90f43e2
zf9ecc688c93f3295942afaba4f519c8f9eb090651f23f86014d2f291470298edc711a2453aec21
za5093d214535e56f28d97a192e1db9231b1fbd44f1ffc3d48449412a93bc1b0e6f3ae49aa49789
zfefb1d468eacf24a70b5a4b8e4c1d5fd2f11aafeb5b6ed0cae8ac697d87b7ae00f62b79c616166
z34bdb5c250d504f6d73078b25b359bea911d84824f75ba4b4b57f5db1eb97e9f218d792a643c45
ze37d8427b9ab6479f6a7d4b0632857e7a84efe725b07d299f29149ac4267de31cabeda29256c51
z2bd2c16b6dc14bceb51c43d77cfa517722340f1c6f55dc2785ada2bf9eeca73ab0db2efedfe3fe
z34b4543bf20b06c90ec530235eeb7de57d8b0ab09a6e768db5236e26dfbcb599ad9eb2ec88c826
z6cae92f0c3cf92ca7bdd2ca1db10f386e386807608151aa62266740580828528f8c620239c41cb
z6f66d1eee9bb580b36398e3f4ccb7cfbf8c2a84deba1000d4c8344e3b46006474e5e4fc852a5ae
z82a67ada83206cdb4df29cf43c20b4543faef6c882f3a104e2469d93bba0082afe458624296026
z998caf87ff7104089065d22908738265ef7ef002676699acad8560e070a99fff50c0b22a0394bf
zcecdda7044a0378a029e1e078a6e49e435648cd1ae890d2a1fd4a3f2ef49603055178b480121af
z4e77e17b44dd6a0d503aafadcece16b2420d4db04a992037c305cab54b82cdca5d6b87bec6fe6d
ze4c6762b6a2cf2dff6a0769d56f3702f7356f59d0a269311652cc495ce69177fee9aca1f0f77f5
z95eacfb58f617c978090bf3c45f42284fb621ea62ff5e58f55476da2272014f61a51b4b5a55e2b
zce9d498fd7830bc833ea7fba5891e3d717d26b3ff5c2af88fe930d910aaab7fdd752e0426449a7
z63f4eea495dea1922fd3ef41ffa73cde3852e408f60816b8cf339d5c75a67a66c552899970a251
z8a67e6df28a0dd00e3ececa78e6ecfd485a89852395c74982bc96b3f52bbda5ce08fe3c0e950d9
z09c71f0abeb2d8791f7eb7f13f9e23e61e49b29aa1e6a66ce004a3f505ba3be3ba56b8518da1f9
z8827a69e8ccbd3d5afbfb167e6f2c8f81a46df718845bf63e8396b262a1715d795bc85db93a9a1
zb7fe16e8e9e57fa21f89adaf344832e037b757c2a56cc9bf91298bfb1294b01adcb625aec13a66
z42a5311497a235d9dc5eb806f3b594ca9a0ee8b288d489b54b97159bf26f2f2562a917dec7aa09
zc3fc40c4b3cebda832276058823d71683df251361c68eff19a77865a1dbeca7f6dd3989462a227
z61aacd36650fbb8f762e16955a69c10242b23030a600ccf3f73a0170f6706bf775d97b381cb116
z655fa54d35aaf5c8ed369b9d5b0eab87abe4b99db131e3937777b34da216dd0c2b0312b175c7df
z629e64f41b33349299147c514202d500d1b3879f6ee8ff8f91ed9ba01bfb3d0f2ab01fc2605073
z2ad0a5070ccad211de79bb6b009bddeb942fe3d7c949865df7654c307a5fea8b39cd0b11ba8290
z7fa0d7da81cc44cfae12d3283550b7f40080bdd9713c01c21b0d7d01c168d641922d04ccb4733b
z9e0786fab73b28bd0e6e318fe605306c779c86fcf2507f2e8c655b8ffd63b1137afe319b4a0b1d
z6b31e3cc5000629b467f5a4165d227042c71e19bb73b91d85a5295aabd08097db54e894b1a74ce
z1ab2bfaf31fc4252f8b562846214b11d9aea439d9cf1709ed4cd61733afb6356046c59bbf664a7
z7a3fb50489c294d760c2b9520f434a079c48ba6b45b61d44d841636c296270ae10473ab839d32f
zc7785cb685182c9f99186987f85ff5148051cd7cad5fefa054085530255c16d1d87149e030d347
z7be25361ba2d16dbd65747bd2ca757daf00801f2a122a50130a7204f53b47bb84b6123ee1949d7
zc6509926ea7be151bf4083c368f02ac6e6ca072799c7a2c6f2ee4215e1cbace5adf13747fd87c0
z7bee295bc1bb7244ba2e53ae410c560abfb658f4452fafa3b974bffafbcc341199bc106adec1f0
z7d591c322374583353528444ec0bbe24172ba7dd78c78399979d27f267f0baf8623c73995e47d3
za7cd3de5320309d2e3dcbb41fa758c68d20309f8cfd43411296d6f1cd85f2ee6bd78909ee59889
z5c0b82c91a7ddb33e34fd6649d2a8e0118c992803e5643d305b142f0a388103ad521a3244e99ec
z2f001549f86b61e617d231f21513fc460fa438295e548c51aa6dceb587dcdab2c53a6d2e4f9d6b
z4e0bdfd7ba0c232d84f2572c1cb09fb6e62642122d876618d4735054185210c8286f8eb3f22c93
za48b24db9326a5face4f6ff9c41847c9c9c2184ca0c2a6766370d61d30ab0e753b27e417f3d03b
zd56736a959ba86c39fc83cb0f9295192212871e3f3583868c010cb2012b4526d71ba65bbaef180
zd34fa6892b58c3371ce8c2fed2c6fe9002ff50645ba3f661038ca451de73b99316044015b5b06a
zf43ae8357236609653d63b0bfb1ae09cb73035158b89d5ea4ced6c9473557cc504a315ae285151
z4c6479859bfa1cc7fcd5e92c221630e8e6252105a853c8640c340d5ef1940eee5763df684960eb
zc5864fdf96aa1f616332695e44d26b9ac2f1a16a0283e5b89a7c5fe0f3750ec0e1ad581f4e6039
z131606857eb1dd766b38150269bd7cc8f751c429c3a5a50dd5b649c8022dac0f849cfe1f9d16dd
z932dc61c5d9960377ea37c388b8da15d6ecbfeb66fdbf7321ba8353f1e2a90d2f57a701afa761d
za5cd954f126ce038316f84a8f0aea30b61965bfbd6206978356c04517a49c5d2c2a6ad27d3206c
z211e4874d304ca55e44bbe6aa07037d495de8816c37f23eeae29e678a15fd3e8544a7bb283007b
z96e23527d06a32b077d42ace4295f17e0e64069ba6ba147f0cf4d5d1ea368c847b1f138bc965d3
zd2cc7154389acdccc16885156f71575929897740540fbe1bcfb0d00486b0da177b0bfe54524f15
z952255f65bde0f0bb9f502c54fb8cb910b7dc7a72605cc6e726afbf56470afa6915e213daae05c
z10cb933d780506911bd27bdf8184842a8b36d16791ad90cc8b783b46a80c18ffa4ad5152c308fa
z33bb2ad85f5a4b6e7b311645082ab71f4cc35f8f17348d051f6afb52d7fbfa3f0ac6d700b16f10
z88494f4d8f94b959fe5b5984578641fecdccafa2d7e78c362a8e5bd5888d5be954ccaaf3a564a8
z8d67f40bc7227228517b1060ca59ed77f41850a93b06809dba9da751e4a9c36ccff98c59a35199
ze89db811ddb6eb519f9ff05ce19990aaa9f44a36ce54b81c5481815e91560b1dff581202cd4927
z3e287046e8faa00e8e9efb23d6c498a25d335b9b5a434026a364a88ec9a028425181065e92a241
z8af1677c9422c85205f976d5a44884fe079d59e686fd0e3fc6305d8db58e22420d2d0648655320
za8e8b4bd4f083e54ddeb917d25c0eda4965f98045ff9c4de412777f7598dd4b6781a357073cfbd
z5b52ba91b8d0708570bff166c9d857d570fbbbe14dfab484de9debc508a0c9ef30e05d531af404
z55a0e489c1578116c70bc213039f8b7d771952bdfe91156140e1f4c889ab3e9b260b35fe90c80a
zd466dcc4a77320d4ca97e5449c44bb874cca6915440433e708d44e74c6ed7e956fd611cd8e80f7
zd64e31b8d3ac6af1bad852afa84f0ea9bda375ce4b6b99a1bf1eed9f0b5405c2cbdab7913a9730
ze36153ee240af4beeb60fe060c7020f03bd3b64b6f72e2453d76289909b441f8a2eea09af42009
za6a595430a97f07dde1956e319316174029d789415b3e5b12ca6c12b111c39465cb8efd8149c0b
ze8720e40012c384e46d717429ed392083c424b088f0a2c13e89d45f818ad6e922842ba0ab8d443
z32eeb4c271f435b1dc4e2a0441dbc3fb4fc379f038fc34503937c43e26b9ba5ab18a3126125345
zb58dd5339a5a9dfe93d0a0bcd52e9d6ffb6bc3f9997714444be8aac567131b073e55b337d5d592
za9f7b1860bb8287c4c8bebd5d290124aa2d6a01c6abe26a8d5d02555499b067001b69c530526fc
zb5c7cff1192ea6b3b75b1738b18e3ed07cad0266b24634104ccb30f5af1bc93db7669ccbe53ff5
z46fd52fef91e30e7f62de14a8cfaff23b8e99cde5b1687e846d755ee26d77378bcaaf420d6c8b4
z660bbf6e66e4c7b2ea2d21247182313f6dad2cc37f7858664b9217d5859d267c1998f7a95ca4ff
zca17610127c4a1e4606917821f5e43e9aa12311ad110110f798af9520331801775a5496ea3b3e1
z3694d4ce53fcce2610ae4823899e0962a03edc6638d52a20ffc3cbd1c1201721d8aa2358107ccc
z0783af6d9f1b0daffaeb98435e61cea61079d040a2e4b3fb65e2d9b8ec185c8c0597bde1635763
z11aa6d0d2f7bd1885593dca185d1ed7dbfa33ee24727af16d2114685310c418edb3738adcf663a
zaab6d03d1d72433c0e69a10b9cb153a9e3c67080d0add7c85f2de4321894b516c59188d16f782e
z8ecd0978528dd34ba32dcda32b80916fb5b849a070179968998e730d398217d6d48986b3253f88
z39ebc2af78e1cd9f4d29d046dfa7b188e184eae10fb3030859f7ac0504c526dd76fd12a53e48cf
z8dfd1e3383cd6d4e88369f63c327ef0b3d9e41b9678676c1f490c970297ff8530f40c7e7435bb8
z74ff6ab8423e988ca4b26f7ac67538cffe520511017eef83534f8cc7d60f474c3154e833a46d8f
z6d46644bda31cb89646261445e88505fa29075395d47892268872a9a030c3867e7ba40fea690a5
z44649bc27a0c78b2e5b6a6647b1c90580fa82a1d0a24341445b3208a6b53bddeec37d25471f0c1
zbcdd9c7656b62bb0ec110322fe88dc90ad6bb3a80817a0464417b5a7c91b3ea99bb0c69553c67d
z401a107fa51b76bec1251087e183d6e3e16ef9679548704e82053d6669ab9ff8a751e387beb532
z74680a1bc2a4c5fe34eaa8a166657a4c39be177bf751801f4b91bd3756939b093575754e7510cd
zbcd50a31c9037476e45cb27670d68aa9983f03e0a0cc4bf40db86a4ab90427f2b67b62f0670b99
zece41aeda5dc9544d71b8c98c53d5b13b52d3cc258c69843506155912b931ad37b6c6589560e52
ze2b0b7e02a9c3cfb9c2ef7faa3aed8ae97406108b3e9c92b83aa530697c16453ec9e60969e1025
zd2fae5f68e9c8f2473bc4daa5adcea12d410fd92b6d105043d3b963f0a96da1704c93b54a8ad3b
z3c3af3c0f0f09929997850bc5624c332640d43caec39ecc7ae94b489a0a484bf5444021352f074
z46f59464698cccb20cc40b1a25f31d69fc22e75b82cb29518c2cc4e59b1ae885b6761819f67e5f
z59c9d167e4bdf89e0f3047e811a5921db83e070eaab7ffd731138330feb65af812f3ce7f13b377
z6bb6036ab4b329feb1f537a19d965e44f5253fc312ca20ac5778129c9b25935192ed7b7bd33afa
zd01e0503d1a9a69af0d788dbe0dc706e310454f61e0606fe14cd12b4e44ef94495c8941602a8a1
z4a0f92e237a83fa30ceecb4030bac4fa75c65772bae633956557bed3c17a3c07925fe6e942721d
z8f71eecce83d3252adb3f65338ce8f8bcb866a14b14e6622db7004065183685abe75c62b73d6dd
z1eb83ddba8b7cee46fe71c4c6e3a8a914dcad74f452e0f634badb2b4e2e57aa82d55405434cbab
z00dab28c445ed1091c529ef14613e08099b90dd66f4cc654fbe50949a9ab6c5284107b5c183c1d
zf6cfaee4fcd821c5f0ae964b8346ae5591a5e59fef71071ade73987b1307efaa92bc04ebf7fccc
z572af4d948d7df4d2e73d0583fab61b82e033c317f7ea37d416a16f03c5c2e774aef24aa7ccce4
z1acfe945f1ecbda21025ee7b311458fb68d52cf0c2c1c6c8346258b90b69afc9c3447b8e70fd42
zc847d9d02a98dd05651e300bf7775000f98699784a7fc438287b2d62d935a94ae10fed8a070e97
za8b2c37980898079fd3f79c0151d2e453c04632246ecbdd8db665a4d2013c11dc22368e9a202a3
z0e76b661acd45be266848e84bd90561cc8295aba533ae78f3fcd413f9541afc9a928fbe21dbf41
z05bb84850d5510104ca19c32a77adf515898dd9b57ebd9e2dd2b2c27ffeb479354fa6773da675e
z2ab82f31eac7a74f2727bc53901153112eef7331c13debf4f41cbd005b105ca37a01ffb06086a9
zafede2ddfe4b7654bf752449402e95149376fe4c41fab889279abf6d32ade9d8790680fafec565
z909061a8f0decdbac05818f2fda8c57c6acbcf149d48b6ba004e02473686317628079c2d2af516
z3f187d55c26eb31946dcaa1249c77721194ec5ba1dcefe3286496f127b9cf67e67c53b4fe5d345
za5d355d49e486b122f369b09f9a10db78483a41ffa9dbe0117d43808b4b1b210ecac64b89c6ae0
z9a9fe4d6a20de22415119326a7782168f170f725003abdfb93a9fe3490e739879492fe9315cc42
z9b6aed01e34eace5eaa61f48466f4f6f9d4924ef16f7b76a6ef52260d7167351275566a925a08e
z0d1184c2ac7572b9eceffa9f2531cbf6d816ff368c6933012c111f8313b7be675dc9357c2da47c
z67a9e00d95750daac0603353c5bf6ec37703322b4183946daba954f8d2b09cf3dd916faf6d6ecb
zc0eda30dcb4bc71ffb4585bcfd65a3bc981d95d81446c92b48fd6423df7b444488efc2810f1fd7
zd883b7529c74f48fb8a510785178845a76d3a68e2f71788179e485e941aaa8f5dc7bdb021ef116
z57255fc699d7c01f51654f035d2fe07de9250f0009192315086d6e965cca4d444b2f0dd24d8f79
z8799ca75136091c1d217ccf72e9e5e6594050870286c787effeebd99cfd474ce6a1736572d4490
za84b10f763874a9b448ec86b490165918b879043db821ab7d81befd03ef4f12eff9cdcacafeb8f
zb34fc6ced3af9b3890fb2c3ac2e229c86a182ae00b23874c6b53a4fe00b6bb9532814fd319fbab
z96c43241434f4a07cd428c110660b28531ae273b3bf5e1ae1898700496aff69c2006b6aef5ec13
zbfedc5f60ceabd9de58e9e899c50445e986324e5476d0bb557d7a33c0c161f54aa090caea8c539
z94a8ff2b499035abaf5e5e4045937855fa5b7488efe26a101f7b4ff823b875c5b000bc695d1de5
zd55a6bea36300688bd7ce59fe331124ed058dbf24ae4ddc384a5b140d47968802a930cfd757e50
z86ff554a01b5bd8d5c670f1c384d5008662e45138d9176f53432a72891920062de643e808bda17
ze0a8a91798fd224948ef20019ba82499d5b0407ea2f0bf67b4aec59b827e7728c51347651eba79
z1cec0a8bdaa360a8ac6044606048f5738e3f16faf471a8eec01b838e13bad6d928e9b325d394da
z7836f2cee37ac3d2825aacc616f5e240780d39dad64e3784f5b0f717e368821d4a521ae414ad92
z633a93f81f2ff990faceecf6a49e442c8a53dbd8903f4a9db3f30ec18fbff6717aa514a51478da
zcc3e332478923cf8b00c6fd9f8b65948ec1dc75d27d39fe16178867de2b42786c90ad4c273ea0a
zfc24779ae756cc55e31c44a2048a43c8aaf77fede5dc2e0a1cb0cbb8cab9076365b75f32f23bef
zf60ab2c09f2924aa7c362658f5d4ab6a3c492b7e40f2498dbc1b9831a730f5decd3e968e0bc934
z874a891e2bbb4a549098723a1c752c6dd3c29d7297f118c1bab92f6dcb7634e260f63bcb910605
zdbbfa717b534ade2a8dbce2f4a00cfd08ccc9fbcfc60251f3483f60f1a94cd79925a9b84a220f4
z406f7a054ca5a8c58df71ffff6c8968f1a4152c1067acf69abaf37b8cfbfeff09718a7b4d63dee
z1b580b6ae08e64001b547271c1aa725dea34d58ad66c279668090e2d6baeedcca7eaa6d25a8471
zd48c24efe40676219188dbd064b91d4b9984650bda5d05121ea568f8ebc72c825eebf693302719
z7ec453c1f53421b310ae631e923f00431b0da0cd13abb7feed2c0f8ee781be87b0add182684f7a
z71e9aa8f79fae94101c1f0f50aaa13bf58a6800a0dba9562bcc08881e7988e8cc0e164f2a0609d
z8089f3ec1ea05650748aafed80aaefb115e44bea6338e16bfdbb201a55a03b6442d507f72177b4
za9b92f8127250f81491b4480a907bc99f0cc53ac2a721d7042cf0ad9c5e5f1e28f5f874923fc1f
z03e671c0abb5b854438e0e981a784ef68263dcc6a76d7fb4ce705266fdd6765b8ae67b77b3ff1e
zd19863c9ca199936e1fded6551a71bed40b47b5d9728ffd5c9761bf9b7ff2f044941278f22a64e
zd9a078a67b9bacc766363236741caaaaa1f3e30c25d4353f88a4c19d253c1bec06728a02e3a265
z1ce5098d349220dad3b5e43b9f9bf2f0721abee3c4df4cc08e80daaef73f47479a443913a32dca
z66d5263dac7010cc0cd6ec5753483cb597d2c252aca298d59fe374e78e4f2a790b7a275dac1952
ze40799770cceed09780c23eb3dfb15f70ffdc35f9b6344cc2c8d2bab76eff1a96590a13bc27c90
z2506bc0ce6dbdba1898c6f0cdf0c0e1ed02eaa26691320bb88e2527d6380cd34410d7039c69947
z4565845aadde72b1b390538021040caa8355b8edda35830e39201014ffa882fce86675079b1fa1
z38802d7cb119de58513d581fed4cce4e15d9115aa00e114eed77e1945c84aacf9760c28bbd52fc
zfde6d0004963aae6276483e9cb04e17cafa70b2fca54dc860761f3eed2838b441b16077f4c279c
z23de0af11bb731191182433796760beb1aa36f895e2c1c57bc022217c3632ee69a6ff0c83122cf
zaf9b3325c800f44d22ea9ec7806107f2186b6df25f42efa0ca5311d284aac6fa6de5db0b76b2e6
z951ce9f9d197c477a7ae49acf5fb0841a0529b0c9177a57e0ab1ac47af9b2855b64dd27982905e
zc53109c17b1123b2b373ac9b43d90105ddaf1b618879d04d9faf8c641da0b9a0ab6ec09b3e4b2d
zed8ca87582cec6cdee9d8eb8fe0e59c429114ae8ee042b1d210f89a223070112e43ab7c3bbd065
z7fe4e4c1c74e4dba76d8f427ba9c3cde1afc077b3e82ca03886ea08bdefeca7b602e17fe0c719f
z724f44d03688ddea6b26d27e4dc54ca9711051292ebcaf1049d9d36e25376e22c60c80052d95a6
z0c14b17bedf68585e7add67c13a8a6e73d048d8af79626adfa02d5bdf7b6a8702b4bd576826a0f
zaa40b7cf7ecc5287f0bae663368319cffca7e82fbcd9f4255df5723d8d006a96011420571f832c
zb32fb3b6713048be44d7dd953dda5a0b39ce2e48c3d3492e053fbb67fa668be6a6c2ef7151ba25
z63c87fa33e2835c9637a05ecb711ec71bf0628ae3d2dfdaf14d2f6431e1e24077d72203db33759
z4782049b365ddc1a466086bf584b7f6100081b73aac92ff265f271fabc3fe9b7f1a84b7031d10c
z88450567a93afb6241ab3bd562a37d81c4ef80321a7a4ea8b55d8c2360bc0e2297dd90a2f50772
za84475d59aa217c736425f1e0f0d6e74be3e05eb97e53d7d2264beb6b2edcad8f077e3a788d10d
z73a0fa00c86be2d1abfcce8c613c28a6cb5ed13562a4cf140959a65819401d37272b3e00ddb76c
z857b670e86139ce032a898965ad3314d2de945c0b2633292e19520b24d16ad565078a2371bb190
z134a7e0fb5ecc5715361c8dc1c8bd1187cb872a732b46d4ae6c0cc84b758563bdf9653ca03a600
zc5386e960ba76bf54c7663448fb08bb78933479a682cc15ab33e9cbc8f445935696673d986607d
z3c7cfcbd0d0d9bd5affb04f9520843ca3408abeba6d35f9a50e67afdbf7f17cb36ddc30005498b
ze61b645ed5980b78f0f92dd5391665acb7fc2a70db9059875da89fd9f255521f30a7733c542bcb
z3e1b13336bbb87734b825a7c48b44633c1d9744f79b913cc1626e2381528dbe2cf0916913973be
z6587eb31c89b2aef3258e5dd0e0e2959f3dffe4d81b825eb0326f2691d81fb026e886fbba137c7
zd66418bba7a4500d6a3ccac7882b6bad27f20f3c088e327923dcb8665f836d36f3516693f950d2
za467bb0b85c8428823fa98e8d44da6348d04cb100c74625a945f39ac8816f0e48133bac59be2d1
za3c5b0cf3d771cce854ab1f47304a12c76eff506c7a7a22671c88936dafc31cb4e530b1d808f80
zf2d8a174d1e9aa39d576aa6a0c126adaa97cd5dc45a115c65662b28faf67b4090302a62431dd8c
z8554a10ef07ebeb0d7fdc19cb6e10debf01f7cdade7f8ab1bdab2f7002234d96e4ba616f2cd91a
z8f3331a18907f2547459bd6567406bc6d20069459e4eb926100ace4162ed9e331d9a007317fbad
ze47bdb7a36cf18ad9451982a7b4b794ef37a00c3b5e7093da228549043632d660992c7071276eb
ze4859d81c7d282d3702a9a35ed621ef084461600a4947ee6a38b60e4b6785c44555b9bc5ed70ef
z151e9bafa56abb7ed00d29bea00ac5b61c991ea194905ac4980fa142b6b870cf2fcac2b9a6569b
zfa7feed46ad48ca6433727166318b5de40cbfd151cc4c6ec813310bc327aca4dba328177869a1e
zb53b1f9428ad3ca13a80cabbfe9ac34d63177e3bf8bd39bf7a25d7d75c713146cff8cba69bf68d
zf2351e1b753188b1786a6d8b1a7d23bb30c2d3a437cb4b8008b40f79857866874bf3fbce4eca93
z3d479d2608f328b0c7019831adc05fb9c20d13619c1350e150e5c92480546f61ea15768379afa4
zbdbc50936f833dd5e3a74908d94c92391b3feb43a0b354f69fcb10e06765012c71031846cebd98
zfeb0520b008efda4bad010244d9b2d2575861705b0a142417e6c1a56ab7cb22547b515ae37cacb
zbcdb131ceeffb70ab6cc21a0244227100bc154483273ac28516788451d201dd87951dc2747bf80
za00f550640b714156cb9a17ae3f768d4a9dc77dbab43a985a23f90f73c6157755053b57185a9f8
z38dd897f78c9c1e32af08d23bed6a4ced9af49534b1e6b98ec12809c370226c0fdd8069f34fe17
z38bb4efa4e503bc2f8c2d3b171da1f60553e0a94d34f01f6dd257aa104a27d65c5d69989b95649
z01c467a28263dc04fb22a7e7e5e1ca7c6c89a4603c68f5fb7c01ccc30979bb62a7de03dd9675e3
za76b91dd1aec4c1dc96fdd0c32f8939592939ecedbd0f4e19c826bf85d7a29102ab019a008c035
z6de2e79242da4ba5cbf0ad490d3bd802e3f01b674d84377dfdb2fc0af4964653992ae1b20553ff
z5cec627f2143447eb5eaeeed009ba6bfe6f55a606e88d338abe68d5c281c7b78cce8a855db5a61
zcc5e4c11adb2e0d967484915edae19b33d434726c8f242f87850a862adae544378232fdc5b0c8f
zcbc72bd33e4faa6b15ac970e8f54af0facf7a1a77e68b6b0c509394fd90a8808cf2d8a10f8ae16
zbf402495c8309f159e08f5aa07183f3483da0136bc452cfd0dc6597423ec30bfbc0be5186009a7
zd729b11b2d1da66ef7687ee0eaada73c83c2499755c76e4bf3ba54a25c244509c515d563869f02
zd87b219680bc8f5702795a1f150ec50e7eb9ac0856f0b211dfaee8c1e2073eb0fa7bec20883ba4
z78ec0640116716d47da9b862df66bb7d6b6e1d96b076ad01bc1f81a613336a46cbd843102cefe5
za1e8187d5a9cd15b2e8f45a0909036621101b5b89bbea13bc7b2160eeba2edd72206bb38ed70fd
z35e94135a0e1d8bd676e4327976237153c4349cc65579431ec0067b2d9e770d03c5f66f36e84d0
z1db04b8e2ebaac84a76001540c26fdba5302a6e74197047a18bb0b5f3ac6dfb76744ff33a6a82d
z8475070bc93fed7c341a0480d91ca755186632ac7bfc3143d22422f4df3ad374a1a47a024fea1a
z86b0bf940ed182ae8ef904e03d62d319c22744b77648d44188f4e070750b3926c5ccde26ab4778
z0e295e449e76ed013758f59a318a7312b4247d0400bc479bd12d775a3d2ac915f93a4ca17ef658
z6ff2d5ec91a2f0a83362213d29f3de814a5ff9d292e6f8cb6fa84243e8257e71e79990e06a1f4c
zd59327be224929d88d1495dd16dba448dde2f718443bc8c43140eba2c7cb9eee0d90283f6aaa8a
z8a50569bac1312419c0cc894cdc2a5d43347f48d4967b980b6cfa6f734038e73d9cdb50f926b79
z5ace0fd4ad4afa23cf084ed276615a864526e34f3094e312f396d3a50039def176ac72236407cd
za9923aca5bb26687fc19ed469444a0705a886faf964896d357c60443cbbb047f4228034023374d
za211044fb4f448ddac3192fa06559c9c263be518ca06f42e8ea911075319fc6fbd55a9ecf2b50d
zbd0e36b5f2b14190c0cf304f6e06e0e068a6f2c703470bd9952e95c080dc6a0a323e4ec2e8e00a
z8989e9deb18b375a5539e0f15b00c1332901c20f00e243c896ed6033279abe231470d67f86a2f9
zac082eaeb3d4b22dc30606f713df4a21ab942f59da1d1946ef921883819c86e0b15440346dcb0a
z4d28c5304b92cd18233918525411812d805d7c01287121a025f8cec83c36bfcec2338ad3bdd091
z0101402f0990a89370216a2969c60e6b705c6adbc4afde5623ee841350dd5fa8e252f2051a0028
z69be3e746bb066caff1c91ba4f3bc0e9a826718505557797d15ea2f5c4bc7fcce149f6ef906b76
z374029612a5fa3f3cfa3759c663d97b3cfd81c1612cad044d0b128eb8c5d19c66e475ae9ee1254
z83736352264ab3f509af3134c7bc2cc68a6b65c853bb76edaad509690518055e789b5c62c3efe5
z1ca95140f6556b31c169e41e7c520ddd977068dc57772777605be8ebfb0e77a2912ada1fb1a6e7
z4a3d7c0bd1e84e68541ea759cfeb270f9a0be7706ea101605e4c65b1cd82d03444ffac6e41b449
zfe0f7ddcf94ec06ea5e1a8fcbfb8d7562b2bf97cfe42200c72fd02b5959f67ae5a2d701cb3fc95
z2ea4fffa1246b1605a833ee05624ab75251830333d036b8cd9450b208caa2ed6236b56a3099fdd
z8f457f312412f52044905c7cbd5c2a234937bd38b765d06572debc3a60860054ada3689dc8bd55
zb3053d276b6d3d55308ce654c56579d1e6cba0b6c5ad0b5e23b0790bbfb5d8fcb873fe352b8955
ze941cd1df05fb02f532ac04226b35ef087d093734c038470ad60685719a8fb4e9d346b3f9ad271
zc7eaf2c4642d8467345aa182b8d0766dacc4e61c213230b76573decdd5acea33279880c3af8263
z0fed73743365e465bc3aca02ff6122798dd846f3449cfd864caa6758f5ac1584f69145ba02fa9f
z4c72cf8490cfce0625762fc8eb450cd91593a6e5638575d492e1decf3d6d362b973508a7e216f1
zb43c7545f9a3eefe2790b116276d86e9a77a0cc3c25197ba3cefba178abcc6f6abec9dec94caab
zd2983ef0e15e439ae711a632bfc6ce6f10d731b588635d74d32c4366e77a04c1239f4dba3f97f8
zf7bbca1650ee484e36de47efa4be031a33f6f04343acf7aaf7c7e63025f1aa7c58c6602a269dfb
z1b04b1a2e0089b8db830bb35e80050855c5149ff88b9cea3cf1c0ccaee1a5ef0049a44f55103c2
z73df2f76177436f468bdc0610709c50e963ebec2d4a8afb13dc0d354a3df5e4430100b5cd5a225
zc640a3423ce83c7dfdc6dff5d1dbdaa1bfbcc78ffd7271be89a72e4c40a186c447a40d7710e00d
z1240ae70edaef9efd92c6eda83e1d24336d04c396a93055c09fc438e7c443079193296aad185b7
zfafddb28807eeb1cc2968ca74a469e625c3c71c297f0e97b613530b9146b99e8057189716f8dc9
z11b52bc4e5a9fb334c805eb612bc837361a382720216f75fb4c240b0ec8afa4fe956805030565d
z5c6dd5a2fbe19b9940db1310ddc526a396bc0a2cc4dc07953a30ac729d8a5c0586bfa62c74ea96
z0f15de5b5f72f3a060b3acbc9e5b0dbf80dbccebbd8b2d83585309ea22c0f338f93b299005997a
z70f4d8242cccfbd8239f59a9fc29baa68f4d468375deece9de542e1ad4b3c7624296f9985b2728
zaebaa05dbdfe23fe81762d8eef91392d183504760bc91d82d32bd8125fa8bbdd1933fa7cd8033b
za5345be0c3573ff758f93b6c2dd063dde78d552f35de3544037edd8ea46a98cf30ea0578af8259
z898b9cad6df78f44cbc65b0c94776b15974f64d090f090b4d983931a44964297484655943ecbdc
z6b7958d71896034141fe1b1d2cb943242981d113068052f09fe95956bbb18398accaa2e783c504
za2cdb031602d4880e8c80a66e87b978fa871cab904e1438c4cdb0a4892e9368d17b438e73418d3
z9f83182d57ee5a1e98a679786425e9963f48a5f1dc3817169d7dd6c9e69fd744a965f61e3a578b
z686a72304d7fc23a34afef5e8026cb30eb9615fd5ccc7e7f9f7f06ec3f05da322c189aedd8f438
z405ee96f5f4993b88a2cd1f26f3c3b691ce3f43ca9a42ddb630d37a41f8441f81fd4e79b5791a2
zb99361923c07ddfabbb8670eb2e3cd446db7e9b609ce95742d9add98ca359b7d26f36aff8b9b86
z813e2fd41df17bee9e4a86a8078a1ab91006cea7d7962f5215c40693e8214caa26e7c18fdc1a1b
zcb0bf81078b2b324a63558ff6b9485280ed4074bf6da1341971dcdef90a15103e58aaa3944e2dd
z5ee2c8cf367dbbf6536817d4865ba4ae18b66648b912e8b26e6ab4c5517f5782c581b5cc470988
z3bb89e0df7aac374cd192d5d8502562cbe7dc0814f1eeb687044d4ef462a1198587e8ad42cc66c
z53afb35a6dd683ae4539bd7a0c47d5f21e9d697807f685951ad44150ce233b68cd12fef3129a06
z1e77d0d504f60d2e6f93344f722df49ffc2a60eeabea4d8d18df9da668b865ac573604bbf9eed2
zd82bd32800604b3b2fff03256bf7cd72a4b64e38b10bd492efff6905f7436686bc3a40a09692fe
z7977b1bd876a29d54b0f1c682a0afa8c3084197328e83a264d3a8e7bfa6edacdc36c8eb28c4e37
z03fec3f7e024583d5daaa71e0698d26f1b502fc86fb7887497095c436593c9bc48181d1a137ea0
z8295dc9c1677088df9206ea26c2076ab59587c9923af797b761583f0b612a7d83f9f33eecdc9d7
za28e6de459dfa076985e82f50b90342f514dd704d19610495b3db7d412a6a80ecbd112f02b4fce
z2ca6e06b188ee10c874b34351f84a79ec993776af5ab84c701ca6ad63becee619ab4e52b1f616f
za68758654a3b9165300a49cdc933cef9f0f0c21d9509010743848b4981d642168c16516bc0449d
z92588868fa86f7c77bd74d165ce50fbd03dd6ea1129a15e2afe831e1ab26fc270bcec9c11d227b
z98ba0ae46a2751fc35631dee7d7fcff4fc60ebfe4b622fda879922485ba200512667bf535d8bcb
za293a33d7f7268164ab1813e02c0b9a1b860310781935498e7844ff197aaa19f99a39d0ac7817a
z72281c2a4338dc811e451635efa66efbe80c02c4533e1e6904542d56dd5b80c6a2ad0e5c3891f5
z641f4785089f9e3de6b2e364864feda76afcc12c7b5f1d00f328af7f7861ef80b5504a63306670
z5859f7f4106dcbb0130e21b85ff2843cbf7a71b0591e6dac9705e44037c75a781e04a29f0b4002
z834b7d019d0c3001b9b81566cec746a648ddf85b20c1f7efb2aea70041616b33496df4df9a19c8
za83b91a6893caeea480da6a8322bc3aa6928da33c57f7ee81143127434a2498eaab59ae78fff43
z5de8107e4ae10f5e07d7940e110ba8e558b1525572bdf276f44f92ffb48c2055157fff6166495a
za6d79f559d2b9b583561d967147ca4c7f3ad9b060951e91d6524d1e94d2371bcc7f1021d6ce8d0
zf0c8b2651b36d03d46f49179d4cedd5196b427deeaede2f1cec980e1883e98bfc70c61f0eaffc8
z443d3e8f2b9e64202a2f83dcc3785a39204a8538e85279b339b6cfbbadd32f2e8a4f17127ac9c4
z53f8af7f342214e06d7e9d368880daaa308683bc95c4e9931e5db7b3a6b266159910cb95002097
zcd0f897fb01675832ea2d9d72f37ea0973cab0ccaf1eed9797fb8e9d3cca14f2fda32aefcd7701
zfa382a0a24302f72448418ac61d4195a49068963d045604db3dba166ed1825670870788e05dbca
zb8c9bd3fa9c7ac64b28eeb649bc4582a94dfff2626cf8cddb0b0bb80ff7a9da117110b45fec026
z045c5b749b93b2849be61de1a90a460065d936e709dedb5cc4303831b33bdf8618af19594da8e0
zfae23b38850a51cc244f2140129b6ef3831bcedd5a73b7d8cf7dcfa5caff956df94627543d443b
ze640a7cce1c7b1b8c9775faadce3d4496ecaf2cb9c41887454e1d876da314abeedcc0f56a5fe83
z90f8639b41b3556a3d3ff26d26f22b06301c3cbead5fd133b3a83e387eea2ebcfb81faed94ddea
zf13e8f4426b4099d31ef67bb1824da33d2362762b9139edb9c65a338f0281f1b7b441cef2d8867
z5c79c3e6c7f46cc280003c875be36c276f3e02fc6c7456ba5fd1d38e9ee11a4af37c51709aa73b
z025be448bd11d90c4e6f24d509ff2cb5735b2a9e98ffc0ff5e290c0430a218f04356eada056be1
zfd04d78eb64326ebaf6965b4629f720c423c0936c7eec72b08fc5c22b6e6ad9487fb1c3c6cd433
za47705fba236d2f0b3862d97615f9ac8befabc5a3fb985d605b4cdfc7a2bde10dd27e122166a04
z192033a0c15f07d3451fd925cb203fb9e1b3c8f59aa7991e5daf5c616d81e5479e02b510f651d9
z6111dfe4c5f316194c5ec0dfff8c2be3f0de5c7dbd18134d0d01c7923f0fdf6e796f0d7a54e6c4
z4348873abc74a706cea8522ed5b5b49f9980ee4a8e1273ef95993d556d1982bd3e522b60b658b1
z65d0ea5af98bdf58728a7977affeef300a02e334cc919068508ea453c3c3afca1b1d63474e5dae
za96431e86361dd37c74ae8c536700b1f002f68f59947fdd8544e372da63d548694bb2a265bf425
zbe14b43303db4927d582cb4cb621dda75b31f7bf63bd2d6ca892e00c381e7bb32876f14d738542
z38250c51edc94c00322e408e1447243dda51b46a970143cb3ec82c31405d5a2d8b0c36fbeadfca
zd34a38d5395a5b44c70c05a51c99bba95c128066027c32ca211386b259ac49653fd8ca0592861a
z20017c890258878fe0bbcd166698c1ffe9e9403f4a02ca008c5bcaedebce9808b57262479b5cd8
z7b7d271935c629fa21aa87b6d6580666774428e1d976e162e28530cbcd2b9d79bd7edfe6eb9fd2
zb30826e20cd884af17ad1fc7ff8ee03bbd02c2d8c04d9e197acb060d7f9a0eb46750d445478716
z556b0f1288273b39a8045b793496fe7dc63cbd1fd6e8b4520134191733442be8606ecf2172622b
z623922b7c66aab4fa3fdcb4c2c6bb2a597378965272b5a234b1b7babbd96ad71f200032a5a7f08
z511b9ac9d5f2a2f4f688df3d75015a39c894e304d1805e4d45ab377beb9a19ae984052e6fc257f
z760cc72f05341e0e283119d13430073181974f5ce56552dbba2dae9dd66c38de885550af5fb208
z4fba2a2db3709e8a5930dff0131a5c4c2799da7ebc3a18ab3b9ad2ae990d705981024992e855b6
z933c06e6f75898e93a63b863b020a4399501f09228782796a49606bbea656dae2ccf09f9f434b6
z5b02a910100db4dd3b49a3b153285b3a8b2b2f1ac447919cbc5efd372881124e9fe09125907011
zd64e1f2fcabab2194cb4f26f16deb60f30ab405e0ec1fbd8e608caecfec510cd833a28d06049e8
za93f3e652544ea340a4b0e5891ae5a7ec47051e08fbb5c868a3bf9a9cd0c1dd046d598616905e9
zb97c7703b2b300c5439245f7126183456267a1f9257fead6f0b4c1863ba7c41ce694ff5efe9138
z58dccbf1c1c3edb33d2c3bde5a476a8c15cfceda1cc4cbfd001bfef6c57283d22ccdaf2acf0093
z13e27de232ef53a6c1e77d8eabb5bd03f1f66b73da2cf2eabc68895d2732f0c337ea5a0c143ff2
z28ab5e9528f89c3ea5f4d0adb347d13f82755a731e97a0529845cc73207c92e5f7dc6574ae659e
z69ac8516c5da380f35adf25ce7d1d364ac719ab3cea4b6c6dc824147104f741d4e5ca071bf40a0
zb0d0733fa42777ae03fcef516e7ebb6fbcbf1f79b8ec09beadb3c25adc212f1a33af47f36daa29
zfc49f1981e47e6323f8bdfa7a411779d14d1b72668323322ba8f1ceeb560bf10d95eaf9069353f
z16c44489222dce7b34b25fdb26c1ac9c691dbb4ffdc00aae73aa5d534e553019c1cf9313a4f311
zdb7d54c0029c42f7e3ea26ab34d4ddf0ba8123a102f954ef410ff065c5161a4c8146e30eda49ce
z57ed2302e84c2716c28fc98e9e0e82bc6b8a8257fd6a4d266043e4b887667292c98a2f859d3d4e
z026d7329b0266d24d6511a47f02342526cbce20465beec83f2aa53f688346b08624348cee425c2
z6f71161f2b1749d82219769a5da250a4b7ce42e471e1e81fe3ca91fc6706427721d97592218e89
zf49cc5fe5d9f6872fbe176156471c49675ea5c435584c1894a2f2a2e37e5ccae703019578f7126
z33e77db22d351c6c830668b7d8ffea11d36884527118b284fd0d1642a746f5331f5e6e8dbda410
zb6f3933d7e4ce042120ad461609efef9f7ff833c89df314b61dd88ab8a9046035ca245dec5f4bd
z42fdf279f1f3eb222ebccf6c1b6f55d4b7f43148272d2e7fadea4a7166c1ebb2b08beda74e2dca
zb8f1a7561d01c2c0b0463c7404e20b1fb41dc42b42b21f935d59e5d60c5d20a7c24467d1fb24a9
z18425b9725b6a442456c00e7855ce250d1a691670ca2392efe4b333c4f514be0a94b9dd6951ccf
ze2802cac44791b7054cedfd088db3321c3716330164b46751b66f300cf85b41ca71a813e66ba0d
z9a0db4191ff43f94d1f156b2c7def1dcd0c0fcda5911bf8e82e1a6048916e1f9853b6d83b9b1e9
zdfcf0ca6e96b3899dd1b2a7a5fc73db6fcecdc5c356def9fd65dbe6f6b76e4176549c12d527276
z1db979348ec4213a9a8522ff9ff50e3af25b07af53f293b6ccd69b485cc3e21e7acfda4348376c
z699cab407672e4ada1d0d5f15b9374c7459955a914762795a720cb57a856670edabea93c623635
zd5ebd8d186340a4ebc46da29a82759c1f65920bccecf704fe481ff9ffe82c794f97b2083bf14ed
z20f5ebfc6e8b30ede56c716c308df770e63ead0ef25ef7eb6719593cd7cbf4e52d757a72e7247b
z0c7d48ba961d466a58e6f1fe42d6fc4a9508aba7bf18bc144fcb6b7570c9846fa064c617231019
z5eab323ed107ddcf71169e84477debbc7b5ed3c87d4c82fd333532a2c37bfc7fa71b95af1d1997
z043a7921204d7834563921be59ce409b139a5e784b7996ba3d670435f1faaa1462e28ca859f67a
z42437e40744d10b52abe52979ff8366854dedd01af9b45f648a9a0d3879eeb341c5af5970b847d
zcf62f4a195223b5f20e0033580720dd04c75aef1788b7febeb1a917d0b8d08f9b18207a914576f
zfc706e6161b6a7fc1e1896e14045813370d13ec2edf911fd59887c0acb1c7d6926c624ddb18ff4
z0c06557df42b52889f43325c9ec70152ab58e6510c0e8bd5b0967379db598be3950fc49cc2928a
zd4cc72b02b9eaa0134045f953c3e12be2da2e7403802652cf3a1136b2e62b376445cb90504a270
zbcd763d8e1a880a4c8b8e2390483c60ef96df52dd4018a5f4b21e8f0510c5a16d14af15199c385
z48b71f785370107e6f10f320fd5be400e71f14c5f44d0716ad6ef468d5ed59753d8ae245a4d581
zd094fd42c52deb7f640d408bddcd0d9df205e4486ca06d5b6414bc648dbfe5c8a618bb8ad4e3f5
z31bfedca5977257e79b305a5ce2f7d5eaa4ff2f5539cca5c65d563cb01c02b93b175cdd2adc0d0
z249cd46340fd89fbcab4688a644665db66017bdb77585cbc645ed552bb071f6b16800dbfeba0d3
z493e1f867263d4186c96300fbb8f65a8874ceffddf2fca0cd218abd7cd56e4f3eb462f5d178c7f
z15075501e4a57e0985e8beccd53a1ea2b125634e6767363b6d8bc625aeeea7831fa14dd6eb4249
zd4c2ccddb7bb34789e4a4ab263eb0e3b21242930af5a1859c152bfc62dd766132be2f732f20662
zc4b5479d4409813728c78eecc1914031180a31535b71179a7b30f36c28396398b6cc99d0e7abfe
zeadff144c118eae31cb34c18b3ced45e6f885226d2000abc45a071683d5a79b7bc7f428b0cbf17
z02ecd3075ac0b1bc7468280e2ce4b3d0df6ed3f938503469b30519f1b8b8dc0390fd8a0aa6b7c7
zbdcefbb07b83d99215afdbb2bd5b6993b58cd6496c92c0989abd67f88c9915af3673a440df984f
ze14d2b85a0997990b1e2f47a319c885dc4d9ba8316dcba7ca91671d0439a57a9f2df26c36c6635
z87e2d23d883bf00b9c2d77b592f5172b1dcb16956dd7e3d5eca8643f601e24c87eaa90b646d0f1
z53647d015e6f6f3cc7245b9d0241917f091431747715b06e79c89e895d239c74febc52c83f028b
zd468bfa386d529bf74518f4e0d0a923aa18141be5ae6aee6606ff34642753168c31152d5fb1b21
z3a533e2a2bc94354d025671d77a8da5bba10fcc195a4452e5230d53a36b17b5258dc40f85cc596
z163d9dfed55ff3a7e6906ff85a5e4fa6901526bbdd73de67fa281420abd29787523becb426706c
z3f4247e8f4448066444f2950d645d52d341e8ca79ff510cef55ea89957ddf60f666a7c7f4beb78
z86e8284273df3a87250f75ede26d572ea3fea0ad0ffc78e94c1d433999979f0e5589d7a478cafb
z9650ecdc95f58240acd552329e15694ff4afa50585887abfb3827e416a62895c51bdb35ff204ba
z915cd002d80a11ad0b464c605e7ae57d1db2ac8520e37f466df89c202abce60ae607cb28eb4c67
z0e213f2e8023a8f60a35e28930ec15fde1af3b21874e82fe3760c09952dd2eb56e207244b7fcc7
zc36d4122b65d92f527ba8329dd99264a02c5be698d231de7535e3fafdb4a5c9291878fa4559a2d
zce5d4a393302cce170d1256d998c613ef85d6529d025c5200f5adbd6cfb55648a30145926f1910
z77eede394b386af7d7dd01df26f7eacbf1afd7dcbcd29635f181e412b8b7c7009229f49a1f4281
zdc8bee81aa2a65218e90aaae7c0afd7a7a462c3b4e458b11c04499f67e509372d72287cd0f2c27
ze113154d1a042cfb5fde39157d965cb2e8f7859a3be147592f3ce01a0ffae30facd4890fd90374
z720138081ec02dacbf6af2ff7c922ea90a2cda935aea11c88a9f5d6132bc03ba9d3e5ea4741b44
z0563ff1aed37a4e79bd2ef0f8be1afa202767520959d07c143ec8673d958b51b063be636f814ed
z6c5ea0ab880c3be87fd3ed9a52f2447cc7053fd68d0fb1be668d6531a28ea9a9221bbb0bcdd286
z4884a375fd0b8688380da0118ddc9786f68523e78f151280eca3cef11b9fcb6ed58a51ac980ac6
z90c78498f93571bd1f2ae8863abfe4c8f1f82dbc1b0ded1cf7e16214d2bf25d4e7187cc33b0142
zbe429bddf188999999d1a5399228b283240552b15d392f893441dff1887d620118ef1e719753a0
zd8f005f7d5b44ad052d92cc62109d049cea2e07e683c84e59a40f5789feef0c07f0be8cefbc546
z8374b1d46f6b8d07a6224bf93b18729e8a2c08ec45805a34a6fdd28eb44f9bc024c1d141860529
z7ecc0f23d35dd7efdf68bb596a9fa37e4a90f62a52a35a57d8e17fd6d324322764ec3beb2c38f3
zf6ec0af3215b804e2278052a8ecb15bed69f422f268b580b6e70cdc6b71c07fd837e907b3d671b
z0ca65851304d319d43bc530b969233063d8c171a8839f67f1ad69b1c76c1a192fbe724f95ba901
zf4a2f17d86a424163c1ecd0446a58c347dcac60228a6e273e916554789dca696b0e25703938c29
zc134f2955690cf6100f1b06c23f2da79bafcceb6f050f1449ecafb8dc63f950649d113cd239546
z62d64fcec7da00f80961d41592297500edfe1cba596dd232672edfc738e0a8b43fb334c05842a0
z7a2bff5bc0fbb61423c8ff84a91bff32e2ac66abf3be674d14f07c90dbef3149090dbf0951ae69
zae83d89785b274206e4d3af4dac042683e0a3df39be875e4ca8bbd340999cc0bdace056cb950e6
zf670ed6e2126915e2a85c333f435607584d1a233fc1f4227be2b6a6fc0648ba3f2f744d74ddcc8
z3298cdf0ae97fb06e891dc566a37b43fb9935ad9daa73715347385a2f6b254bc90006ca797b789
z3889b57d74588f92aa3e75cdb9e3136902241a89b8c4bcfcb2d16288cd4ba113abc63811ad24f0
zaadb502cf8cea8b6cc60947b689bd53264f764b540650f7c5cb040cecb85faa9d7168c5a7e2039
z643d8aa7dfd553dbd50747b3a466cdda4dca16dfbf5ec1378199c85e646eebbfb85bb8139a6683
zdba34362bbf19cabe9bac5e19d8dbb4959f1584bd1c5f1e6ae6f5c82c430df0ba07ba22b31c6b2
z4e0713612312bdb3645db5783af4f3f9d860748a653a22ab35286886180fedbe59aaebd2cf8274
z340ebb0313650bba3ff79874ee6b0959882b72f94afbaa5303ae293e31eb240757f079c7d6d2f3
zb290c62d4e3569563fe414e4bf0f124e25caee7d8d4ae70370fea3d9515060935d856d0f6c4b9f
zba1c3987ef926cba9b5c39b1f78e5a76831f27e729c456048a977d06f2ccfff68be48196bb31d5
za3a3c19e8904e875d97b7f64e20a9b0b34841b8be112975045dfcfc6ec37ab41bddedf54eae6fb
z373b0101174322add96212ab91650b3d18326d59db8dda5c315cf27eac5867a452ac7b2b70159b
zcd229602b21190cb44889d8f0c8d1f6adabce265ad43e35f551f0c865542e0fc3149b6c21879c4
z85440341cfef3c4e3d5b01015e7f238d9ae8e2b1dc1bc0e059633355ac827647dc0c9a7017ba8b
z46ad41eed094833e63faf0cb3caa0256bb93b82f5026202846f6d4a3ff58af8390c21de896dc9e
ze10d4fa9990ceb6dc203e173434063b2bb03ed217a374cb7d5b039c5d077967ed2600164e34ca7
z007b0fbff75bf00d0f5a506f66fda151f24a56f2114225ef7416be77c9f0b82d62b05eb65d9500
zc6d632e6f8b26520ba1ea07bc766068ef6cd6c9dbf0926f45dc586df429413b11f3c665fca6257
zc0c2b850ee650788a8b93d4359460d23f5599d22c96e524b9eb9a3044187ab11131fcf25294418
z082a46f376a12a048728587ef8dcbeb7ecdac246e12d53bb1d983872c24fee6f91a6252b194a67
z183e8c8d14d81a26aafef232dcf73cb5c075ffb1edae1a2bff27ad246a8f24a1774d2f61c1397e
za57e015a199c99cf7318b00689d314a99e87676ef1fb35904fe17b9d82741e23690bc637074543
z6d3fc02d455e2e6954e2ee27a9ac5e49bc0953d07b22f6fecb4461cae77670a5a00647cfee48b8
z7e5e423b7f88a34e7737b0ebc61d51111539a4b9949758b03ffbcc974182eebbb5282295841f3a
zdf054157bfae54db489a23e765ea45948118dd823682de58df91cf876cdaed3692e17555b8fce6
z56c5cacc427e86693be100dbb9e479e08b203ea35ce1336f450dd704c053dc51cc6f392cb14928
zb50521d53ad0eb81fb93a1281421755b3979e0d560029a4f77430b149404360f51e2fe4b924f32
z9c69193efd03c4d699e504ad5ef0b685c17e9b590b7f51e4d1ecd0b9231326cd68f36484c20d89
z587dca56d9408bb13833212c41ba33d7883e498fb3c0a0789c88cb7475e33323328d1ad7499751
zd908f0c327cb92218a64c6cb1167db8e7c1acd5712be18995ad195809fcf491a51515f7bfef04b
z47e812cab5def266616f7133bc90807ce1fb72ca6da462510decc553b5da8bf63135c1014a2a6e
z2d529ebc340f6c18a4d903e26b1cafc5302b152743f7bbc8b5c22c2b4bbc342873b13512aba9c6
z0cd40dc3b2942a971d23c23d2482474f0cae726ed4319bd6b7c9ecf761f7f0051c10a762e5ca0e
z3ab523e4e9537d234c3b1b7e4bb1629bf9c334e74fee1bb1781a42a0a8650da56c8b8275a85687
z05f92a7f44a92d76cdcb06f24417a3d4ef0ad5573fd03bb32ca10d8ba901a483f476f3a618c135
zf03533cd53ab9686dd7918c051451d900e82148728a9048e648498eeb1ebcb514b3f0d609b62eb
z5010f40a547f1cadf92ffa0c9a655a091804d280cd1a65174a1b54af50987ffac114168e784049
zd2b5236f3dc301b30ad3a5655ece2aef23767f20fc5e794b8a4887b07b47753d342757cb778713
zf8817646ef9b963ad62b90b8e9badeba4c6a813e57326e5b716dbd8959963c4e21872cf6c0be3c
z09ceadb8b5448169818fa1b583ca0d84a91665df5a3f37b5814c15ac85bd2ba249a61b95b5db7b
z80cb20b1072606c6b17901496bc144433f914ec0d08f2c1bfbe8c23809112ee9331a08d4c331e0
zdf917d77dc498031bc7ee367dbefe03d1ddb5dac841e71187ff2b119f1ff3903500c4c91592921
z0fbf355c95192eb2fb2e7e16239ab2107a3f8928263e0cf4310cb437ffefe9422fbf3d410cf7cf
z0e762e4ab373f74e02beda62bba542f1f400d5fd4c0683de5f8ec569214af59b028db174bb7fac
z423aee9261037b7299597400bf8013f38e751f6487a2c90fc8448d4641f33f8b36c3b30effede0
z90bd22fc9cee410e6c14aadb8b581b02faf91313191a69415c3870f33c808430607ab7affb6096
z7c9572f03f470f2fc83dd1054802d4233147a8323fa9a3503136fb3e6c6e6df2b2f330eb78a773
z70d2153492cbdf874d8ec4d1ccaabdac7cb5c6430754c5be7702a456bd21bc1cdd1c87275ec70b
z406089431f7d4981d5bdcaeb61e53b949f9ee1764f25a17ae92c9f0c663a42766a62c3184025d8
z0b2a0f95414ba11c71f6b13ffbbefcffb75bdbd7ecaae1eab0a279526ae8da42f8cfd9091533c0
z90731bf2c0913831c75fcf7f0c6806d52897913e1f54c197b3445a02b4fac8892f8fa60bd1d015
z86df33c849b2b79a1f36ede341badeb6e85224facbba81226079a9895008eb038b6b8d3fa70369
zd36b30514c66aa45ff84fdcaa41ca5c53b2d09649748e13d1eeb304be412c7dc72700bfa2720b7
zd96c326a2a6ebc6c7af41d1bfabecc22bac486ec0ba5f913e2dacb762f4be8f9d4a44845268bfa
z6e851f7cc967f3cf58b58cb724d5816bd8e4edb21d663a24712804955869cb42f5357ea3ea387a
z669b5cc4f36acffc229fded97fee366d1c1610c9c8026a6d485442b55fc246edbea6877cfa77e6
z25460cb517779dd96f3b097f6cc2cc61754bb0ed4914688ceb46da239c2f4300e2fcc655ded996
z2d75eece1c00fba0e7cbe1881f81ba94da470f6399af64afacddae3ace4815554aac5b72c506e2
zd817da6e2450b8eed6d4aa88a55c80d155ed69605dd11c996ad3512edae7407ddf0c9b842ca90c
zc224c286b28c3a136f5c37b665ba1eb126f16c515e02af1aaa4576290107ff9aebda7e265d7eaf
z5b26ce74188e581d1a9518564afb7101287d1b9bbab013cc3472f473070a3a042ed40166296a50
z64bc392df851d84ef6a77bb5c3f7358406fff4536421a3de2ef523b62b11e6e50dea92b9465452
zb4ffe24bd3a10266b51876a35b4491413d45f56c5aa10d7013d512fa1b0acde0a669c586264837
zac258272915d1993843a8ce8405fa98355c8ce74c444003a539b231a86f2a46113382ecae1ff3d
z5fab57f71339be7bca26cb1fb347c6fffb4452d5867b42c07ba8b4f84f9d3f84f1c224f642e4c4
ze30531504fdd346c212a334e011e6d9454bfde3a0d1913344592859ef0639f630fc6ed742e9251
zb39061fffa65d6b020fa8ddc2cf141ad6ff0c26c8292e1e33182bafc318fd82599f16edbebfc11
za1ad2d1401d2fc7a9f83c0883ce63b582360bcada6b76183c4c30aaa69f3df9309434c8211e67f
z1cae4753d40315ab40c290cbc8c76e375cc78dcc81d019fa480c71a759f345f102b2db1eed860f
z740b6c958025c06c48cb2d75024f8e63fd0fb648a56821da084812953158720018416ce58ae655
zca65fe679249d7ce62f40262ddf15330810516d2a16be140341520d7938df18babb8c818a91a77
zbd0597aa01d3c0d92938bdcacbd468ce6c575d9d26a523fc6def89a5a5a5c7e8e0ad7297e15d2e
za80506d203cf8f2e4efd2137e20adc25b7bd8ff4ad4da52684f6b01bf1d75295944f84396c55ad
zfbc4b7bbd3667e988680a55eb6c33680efa18031cd5dd5d32af7a5dfb32ad6a6e224355704b728
z96eaaa17c13c7c2aef0883cccd5c81ee45e7a9ef662029682557aa01450cd85ee42fe9115d6c96
za5698c6237660e8bd42e037a27d9eec0626cce3c4a647c9fa901bfe001e4d9fc401efc72489b87
zf77c9635b049015b3896524906057125d6171c32820f77b349ea098cef7b9f0aae71e195ef13d0
z371392ef7b501dfd3f9379168bf641f644ce8649cd16c42f7b9ea9b0252f315eaa372235fd4de4
z0fcc37e4c8770685c1411e95d833a6b2b324850e31800d29a3ab64f0f57f174f130895da4085db
ze020d525a7049647b52fb994c1448bc0295ac2c5d7e3f703923e83e73194e886999381f1e266c0
z5528e832c72a9b338bd4d32d162716f1c65ac56db96f1faabe17ab11af4a459d095bb21a5cbf73
z59fe9af476cc38f0a494312bf6f27377ecd55ebc18b324562346fc7a83038ab90714902f2eb6a6
z3e2ac19d8f085906e40ce4ca5011b3e52ead7defc92cdbb8cdb94f41387cfd3ccc7d06f32d3b85
z5da8f500470623ada8a8029b851471053b3f5d61890db1318e7d997ac087a2aa114eb25bf00d2f
z9944c4bea8631c2ad238f97ea38f0c8821f00750c884d8e9e97ea9d753cd50a8be9e3205c00d91
z76ed12509af07f995a48e13b5cb0c53f46c4b278eaa74cc53dff619387c8f802e11ff83451cd39
zd676391686e69753e9b20ea811d071b078fb41c7fa48c5cd825311a4f6da2342307bf21f472a11
z65b7ac49332994d29e3c404ea3e8dc6375c2858a4eb377d511f5b2823458830b99773db38ca9c4
z9cf50cf2a5456f3787073e996a3fce47b3bea07d342827742073f93101d6429d38e6b0b10b4e12
z8389be42255d36c13a33c8124d6b0c983654f2afc7d908f36538e0dfd3e1746d6491ee8248095b
zc39f0948d3e0846db9366f6f13579452bba98d6b09193e864e975feec90cca849dab4f18c0b12a
z50bbb5a9b99309a11f054da2e6d688130cd019f8761b13adcf7e49e1ec6a95cbd25a9e3d576eef
z2c51f0729730b5e9cf856cdbb75774ae634fbceb11501e82d07148b025a7d271e74e03755794d3
z109d4a10ea1f73c7140d6893d33116f19ee38af08120b463994e2ee08fc396ae68ca4401ec200f
z52e54c2311f16dc8133c4eac95254bb2ee7c3d8285112c766b7eea308079c95d18634cae988ab7
zdad36d6377f21687b4a0cd528fdf5d41128c96902e52e2617a739f1edd8ccbc9407049f7106485
zc0d09ed18b5dff3a5ca3ec4dda239d5b42325d02e12a021fff010f097e9985ef6fd1effd98704b
z3562508326db64035f4a3fd2fa667d178da58de6e03884d61703efbc4d5dd07025a47d961ecf1b
zafe05c847aab32863a8d7b92962a0481b97acab60d437ae8eeb552b013303fdc121051d5c24948
z7149adeee7beb2120bacd829d9dce9fde41435e8325a13b3f50caac605f2fd629419a8208bc4f3
z12052be18ce848fa06bb64b1e979cd7255cbeec101cafdbb4ed2d7ee46c2e7a71b60e19e3d1821
z4470cc4ba8e95f96e02f0368419f3a7c0a18118add85a776ad6b6ec58006a1c29c3c618e3d445c
z1993ee7b19e904458617510008c25ebddfe9f6abe3d1bd0fe8c3561ea8b9282919b5346be361be
z94676e3dc05bd553ac2b6c750588dcae23b697cbc6a32bf719073957c9b6bec291bb57b610849b
ze5b893451f36d464c5ed6511b891cb9ab13d1cea7c40358042ff30ed2d4f6da6788d4505404442
z9a9669a4a72ee7357ec17b06bc8f61b171a0c5cfc5ff9653b81821c70775b94ac95de0695a23c3
zc5c12a84d6f5d0ff5949688e2527823d7905ee53807f5c2517da7a4c8253010e19634e7e58c53a
zc867995d5c598e090cd22070f63f75e0fc8e3afdc08962594001ca0a748715fdde5b8919568207
z4deb5992ae54e39a7764aafbcc98deb9b4f9700ce4b4f8574cafc0cacc1fae10079f0c297292b1
z83e308ac841e66bc6c9a53eeb2674bbb3855db90dd667473a8c01a106788cbd4b95e3112321e69
zabef2519f7cddd10aca8d60cb064792a5023763b526a9677c7caceb72fdac5efc70b2cc699970c
zda83dc1dab00ffb51cb964134201b2b75bcf90f1ac5c41c191d4d022159bf0c60eded3f9df4f86
z312da3e1fec012ee6182d79fb855a640caf7faa01dd9b2a42b27da006f8c98eb001c550566bed9
ze13a75ca056f1caacb58867bb6ef79dbe5438234e9f7ec49317a56079512593872c21f80b8114e
z82302183f3c261a5f53d38c5e69ea9e9a037f7f036ffbf0b44ece2161d2f4554046e602432ee93
z554355a74045bd0c4749494ffee63a256872b32d52576b0e615d35af41325a3b9f657dee0bca44
z439b47a2ec81b577d3a46db64d63be161c2296650143478c1f043f62d67d71a3a4806bc5baff28
z7228ffdc8786edd584ad3351127d99834b73393f09dbf0c53ab9c99f6a85472b26907ae446d1dd
z0e80dc1b6cb8d0f54bd515c8f39a8983168b406d6bc759759036a09a5169c93aa8ef57cfc891e5
zdb71f85456390afa2e2943f28aa1626166ea82c2b7d64a67e20723165f361f2eefe77c5d1c3d84
zfe462243b21e41e4bbfa8d5906bd0893dc1273982cf79f147466dd547ad5128b31e0a0812dadaf
zb5051053c83953ffe9cde6b70c16fe3d61271d04d2e410b37904ec54b46c177b93879414bfc574
z25f39e53abd769b49a4518875e6aac67d30357821df3ed2f84d4758267643c39be0bc56b97fba6
zf8dcb6cd8d6b149632326947cebdf5623c686b9adf3f09de5029ef2f73a1630e29c69784a72de0
zce9f73b892527cb3e5e0e04492bc3ccdf077e95cdd6f65fb0cb8ee0df85145abfeee592b18f0e3
ze230546714f64de649141680bf599687b1a7fef5282bda54802db1a1d15e69985d37c740f1e192
z7ae4efb43a19cba428d1378f37e6f99e58a6482d6bc011462833f168abb14545276fb9caa84585
zd25ae08ab6766ed6828bfc11ea8fe893bd749b456ceae867feb3403d6e7c04eda7856d0fd7ac18
z72b3643130ba28e8cefd5d8935fafa91370467c4f82bd6f583fa907272114b23d0c1486e6ef71f
z7a2d4494eafb9440948adf7c7ee0a3a32818a2ca1f2430d08095022946480c0cb6833545ceb16c
z65457fe5f3b266e70182d6e665266ca45b16a05527042b0afea3acd2608941bec976688564dbe0
z6890a82b5da79a14e99afc70d1484ef9b811d1bb0d4d2761883c01900a185111a560f211610dc1
z4bc3c66cd5296460958dafc5f79ace37290ddc22e5bdbe48fbd63a838355b2e3214ac7f456e572
zad97a9cf0eab156bdefba1646dfc979c7ac66b19ac2bfa2742eee90d20d01c06321d6671aa1c62
zf9c8d1b808c270c9c911380019fe153e494d6030b68ec8e333b1cd626ebf0fdc3911c47f379a5c
z744835b4f999f8ba4d6fd2289805f4fe3d5fdbc5f85f3246a0b328c1b33329c1b931be2e2d1b69
zc8c86c3558a3e61fdad0c27f1652ffb453e74472d6e9e0978a23f6b9d096e703e208127a388e59
z51979eae947c2bf7c49057896b30c5fe4003e9812fdcd3e55d3add15500832168b6dd4c138a84a
z66c80f080cd98e6eff3a497186ffd51fa5a93b49a7e749cf2f5b8b77715928ad9f890b95b770b8
z21c70300b149f86d448573ec84f9e0de0af031dc57b8597714bb6af72cbaa9c2bec61e0245699f
zc1c29c90705fbfa95e9140feebeab7676fcea31f18616dd129f4d39d19b2d362efe4bb89f12093
z21704bbb2b708369ba5bf9408201424ccec17655e22dfce9de06641388141a561ba27567cfbb25
zc932e5eb7c5e1aa07fb15bc5346a7fa384cb6cfbba89e2804837c341eb92c3773251e760b3d81e
z8dec86703032e0a2a62222f6ae887c35b6d56d8d26ed587fee974bf2aa9af0d092b7c9da971489
za6f11d57df787e14b29f675db2f7f73641563d2a1fda5842abf05a976f5078a2ef31a6c3b5bea7
zd6e9977fca83e7a0d1d0690995d81956b3d37dc7f0c964249a0f3528bd0bd16e8d215191ac0dc9
zad7329a96768799ec0b2b5fdfdbb64ba4dc8b5b1b9e504e915417c3f1b43fee7a84e4f43c461e8
z47ef995b1b627feb7615804dbc3e389d954006b97906e6f7ad4c524e5ffb5e9227369570c298ab
z2e1d9017dc192b11a73dcdbe18e17418e6f4ad71ede8238463868cdb739b17a4a20ac9f7e0f577
z51df76bd846a5a7474b9b7bebd67123d0a1f804d7356183a7a501278ed2a2ee648573a443d9ee8
z08ab0edddcd2e7a3dea13c9793f7d55ad92b38063a13f3c26ec3d1da58dfedd4f1ca9c298b7912
z911fdd4f2fcd0d75507a2e1ada017fc792c163d117c4179167003e560b052bc6754116f5dda3c3
z3296963b56ed9be3f17baf3565a73035996adfeb62aa8607990831642f989cc3dad16a770384d1
z92207024d94c4ba8fe2f73b33cd4248795ddad445abc82a570c0ace8ed481b6535e6053ef95367
z60b8b154b72cbaaa72d57e73263bb6169d233d1cd991fca93feaee1fff5f2890947c8e13f3c1e8
zb3db69ef2a30290988e0db522ab2a9edf125df2dc3b5c86a540cca8d3249af181cf43434748664
z63a572dc993e70ab0351d8fb877dff27135f578c8ae026f236cab9c8c0f445beb55c2171bbd47a
zc26fb5426d40c927214117ac282f275b61637c1f9a3bcc01e0e76e86c99b3cd24da79f939dd8b6
z0ac1b4b512baae17241306da81548fffc5dabdf86c1ab51bac8829b2671b0fc23c6cc80250727e
z5f8cb93f2b5997ab07809ea0ed873beeb28134b1966af53b09824af524770772fdefed9d72dedc
z4889766b29f57bccbb5ef30f29e40179e0b37110bb40bbd74d117be5bffa6776e52c030f260b71
zcb652b2ccfee1df087ce93f605f01f3a03753ca9d7197a41f560c73cdf564da0d1c772270ad918
zc5e0ca7fae43d85f8047edc60607532ea79528d2293bded9d88fd58105b37e7d05db318aeb6690
zf1f0f9ff401bbd266ae89fdb9a1b7df6e5464c0acb4808891f0e5aa71badb7869f70a199dbb048
ze30f8b26c667767018a25ac620230556d35190bb15ecfe697a5520c7de85b10f0c49dc346266fe
z8c9863cb1352fcf43fbe61ac2f50cd9c61c0383a96493f8602da0ea071cbf7b022ed913f22ce82
z626b36b1179e69d36070de8d5a6d8e5cb5aad4cc4820403a5deecd81f6d8bd3e0d0383015f13ae
zc22d59f0d0fe2c0c372b30459488121f20d5f3dda8e00a1db635e93da93f127989a1ba9f751f5f
z21dd67e97a6c909a35da292efeb99d34aaeda501252d919d7f114180b734473e04bb95309bebdd
zbd09f71a37e900739a50534f8bf68fe48458593a5db13d270a4f5743fd8e0f1c0615191414390a
z440e0369b48eb3d1a5ed4d2c39e0bd322c496a43e1b62b1cd3e70d755e962af8e39d093d9b9b57
z1b5844b3d777818d236bab1618a755ecb2944e2d59ce79a1cbe0bed333ae46a1b6ca92315bc2e0
zeb02ac88166b144760be13ea843ef69c8b3b4e4dd8ecc93bee9da6240fb5f3e1cd6d39d3a3282c
z92eb8de16127a16a11aab7b3d2a4b270b44a6b5d6828358e1efbf2b1f1875e459d6d49b81f8160
z67ebe05d94c4b5e63d8eb3ceedb63da0947b2c23fb199f110b8a26b6f9d0f36ee321ed5be81f87
zab9eb9ea36458ed16abc7bbf1c0adb4233753b71855495035af5c580f4971703d228029aa97d7e
z2ab23052c8218baddbbfe8d5ffdb9a8f91428450ae9e9f84ea9ffa84ca65120ca3df64c1826829
zdbd14da49961574b2627aa9d61b5944181ac94308d926fec6468515a5212e6b1201b189d9477f5
zfdea2426d3afb21b470e643e243d15339304e0f386f9402cd44c5210009e25ef0d0cf24b9daeb7
z50440441f52f43899e9b27ba65c5d8cbc8f3d5f75b0252a67b337a50c637066218102bf265e1cf
zbc807fa78cedd8d8d3c00b1ebea31dd3527dbe90fc7163d7e362870694ea1302726a8600eb6ea2
zf2717a6f798fdbd97318a446b31e5bbb531dda3e95ed54e848c7d14ac516b6924d9fd33dcf1d4f
zc965d636adc72de8c839cc1a097ed316445dff63aaa5289b5fd4a18a4edcc3d8a04d370907669d
z58b1eb173dc5ed244ac09ea9b7960c523a69dabefb56e3ff0d5e894e5aff3c6cfdb5979a08717f
zcb05cb38e4b87d2b16f632ca0209bb701e29993d6c8e55907fb0f0f4019611f6d9a28e201f55db
z2f0ce65367d00f6bb22cb20fbd59dce37e089f074694a3d08394c62749fa212127b2d4f7466bb3
z23a0d99ad0512c85f3aa860be7160fd561d8e7a7712e2e2071b38db950427c369ee9a9ea98b98d
zd3afbbe2195c2865202408c71f9b282bddc74ab5f159551aef5a4e445514d12e939c040587a81f
z839c5ed111863b72422c17ba6203052c3f33224cbb5f76483db73f971367fe3d58408cbe1e8691
z7b83c6beb549006959665fefb1ff0ebc64ad7684a91ceda2ead8993e3efff6a80734c7f82dfba1
z06231b2f759cac38c7d4fd27352dd9523b2c224d75bf18ee9cee072c48165f36bba5d1ea4ffc71
z9cd4edd97a12a143d9a361dd09209700c415d500d686931fc3f47a3b9a080e6058df4104524082
z5e28a62e3e84a132c4597c616f219eb9cf7265781904b80beadcf53e48eb715a9f42efc7aee944
zf44f95a32524e93963a2c0d65daee8c1dd57040fcf7e08e37bc2b858b1d0b89d8ef42c898a29b4
z46c17f53666ee3aec7dfdf685d0985add1f0bbb12f2c80c2c0ba1a0360db66470d44d60f3f5cb7
z9333eef8ba31328792c07cca82d93c40f2f14098c5355f9bd92016fdd0f4709ac0ee4f662452a6
zdf59c20e37a90a962698fca2223253c03f249b7590847282f798e9d1823d481bbb8b258e7f79fc
z3d67aca40018f053f2f45d651c0d4124b13a2aaba9418bff4fb5bf8c997d9c85a6a6cece6d956e
zbb3e0f311278304b03e08b8dc3c9af2ef88b22462bbb3b2c85dbe0ddb5672872f1ddcf0db03129
zca2530cf9dba5d71122e23c1ce8cc0c810d8bda69583862be0a34b27375571665ae93f469da4ed
zdf3c1519c4ba5c960fcb0c808c672be3d158f6003f2e97de659c998a75e5e0b17ebf4a49bb41f9
zf21c974b667bc0135dd8fa8363e215122a7679a2dbf2a9513a1aebc3d735476059e5347f70f2aa
z37161ee7096bb289436bf2421f5d54bd7d07495b7d171d124d9b868f58943c228b42d39f8034e5
za6dc9fec5f7e562ecaf081d8f8a489acbf31014084d84c841fc00c751372cb0d77e748047f4017
zb2454fd3d915bf33dfeeff3a660cc951084e6a163b80c62fb2fe9cedacc0d5925afb5be7c0e783
ze2701ff7a79ae593c6cd60564fa95829326907bcbc98a2a88eb5bdb2d6fbf66e8d77147d30b277
zc023bdf45ce6b0d27fea4e1ec5aa5e8d877bf7d1fc79cc696ec5cc941460f4c612615069d7cf1f
ze76800334b892405b36464876566340b85c05d1a62956628d602530272d559e45d56065e1a4c6f
zab95faa0f25fc80d4459c38d26f673f7d5a87a194d46b0d8d6fac36a5927767e161a17a3a3a814
zded94073965eed3ea9912fa008962c0afbb089a16d980a5ac94544c95a5eeb11e7d3ef49a2d466
z06dcfb06a0ecef5fe3a7192c87702bade54bfa39bee4480b39e57ba4773585b123268c77c1eac0
z6a7c72a605487ec52ef20628d9c16384db7311285188f418f72649e2655c609c15cf887770e2e4
zbfcac27bf3b86cd60e8a299cd7a31b8f657ccfe02a0c4b900f74ad3dd39384fa1396b82394c57f
z791acf4ccde239a63f119581dab74b42b683afd178edc47337ac31ff39094c07e7138acd0d2e14
zbe5803b72c4cef265d944c388e33f1164338d56aefbe21c0f0383c4a1d8bfbe71f8a05bcc4963a
zd2a6c10c29a29261d2504d19978cb1bd02b7972651f1f3de280239fe9fbd99ea720e30accf9334
z17d34c1a347302965048ad7a9efb07b0fd2ab65f27d3a969d5600cde8954518e550bb717918b44
z16f64c627494fa3cf8c413c499034c4fc8ef8d5cc4e717f541ca6db36b15d1c6253c9fb730bf0a
z3bc7898cc839e840425ace6d531d7f107add4203b8e2d007a8a24e6c0a2dcb42362afe75607484
zbf54db38c5a9295d58b41ff4e77d645e347db1efa795760d808fd7f68466d746f8b4bd2f7b138d
z557499dcfd1e914b812418f6e8308327051f455f5d8b3bbd123b53b177e14003ba812a3a766dec
z22f7244e06f106a174e2108e6fcb369bea43709bfa7e39b76e46dcfd236009f5dcf4ea2852e162
z7be79c11b5bc425df5cc74f595cf9292a34d8e67e00cd73741202c3eaf4e832b72f56088af3354
zf6657de4b34a958078f7c69df9fc12435279551a202d9994240c307bf835c449650fa7f927c677
ze804aa73978b1467688c9783bee4b6b428937b0aca47879714177309009864f99006ea5ad35258
zf950b1db00efc0220cb1c4f9697f4aa679dd6a2606dab337c7aa20579c2f95f88019f54bf1fff3
z006ce5e5ca7a51ef7973013a9d74fcef88f0819de608077a4fd09e5d665bbe6389fb7740a766dd
ze023669d52d6c5a1fdd912987ac6ff447d3de7a0e4628f548e597f1e694f0d70d6421884dae7ba
zeebc4d6f58b27848576c61747c55dd70f071780675700de95155b8919710824b3606e9aabcffed
z32f075f4fb31e15e269f0f113c4c317890799e0f7cf625f0296eccd70113d5bfed79deaf369f85
z39312ce2ba78773905e7ecc53156f1176f71dd2319017a8d6209a536fc71ff142fc52b8b451e2a
zdbdad6aec93c248f1094c5bb22b77949c39dc7d2549c0ffe4d3e54ad5f7f6e109bbb77180af167
z2f022a5237f2386425841c5f0ceb3a663d9aeb9e1ae576077903fce8e969b4f93f8f0b29f4718a
z6ced2b9b2f7b38608b4520ac0c5cff499e0bdec94e1883acdf2e8bfc7e9f7323bdc182c49d2fc4
za89b445647d59803cf6d93eb3eadbb0334f673fc8790131a29f39dfdbb450109450814699bf6ee
z9aacc9494de8362f83285c84303ba978815a6f4055bd448d576588a24d5ddf78bcc5740c2b8a4c
zf367cb7699f7782abc66d00f2c772ee873556850a215e8a41524a52b9745d97c7bf808ce627eb9
z8b758229e77f753437a5f7a004a232a375ac46bda7db7298fefeb368d86548f717f3e3266114bd
zc63deb37283823fdc3681453ab486f9880044e2f330a39495aecb2302e247cb7dcaac9cb9947d5
z6f9de1de3adc2486ca78d7d08f24a9c0f6282cb5cc00a5732071d89a2c34c6d34d0ca68a9be9a5
z3160e47bd8bd576a2f77401e462899c336a9589298a6b067526041520db0bc71c41269e355abf9
z82ee898c768f6b91ccacceb3905e65fa3bd6be1e669d0c9ccc9d75fc24d6ae9d74bc5844c52ef7
z99eabbd3373ecf41032e70c3db11d8a6e2703095660c743658bcea21a58424dd89b36bd3af5f42
z29fa2a0d6884792be2f448af024178a62ad31046c79e4897c6c64120b6e95c29620647765a1d30
zd7153f7bc4716c9e568fed75da000b5763e55d682249635dcf3575faa3c2e083d89e23f4e1653a
zfb1fc727079fc0526814403344e4870cb501fea263911b95fc25adf619d838790eb8418db137ae
z70a590eec5d19120da58afc6560d547b4be331b665bbc813c8cd41a76ddb0c9aca01b8191c720d
z5132ddfaf7f9f600c4e216c661a0ce8cf78e7fadd2bf71df104b37df16f076cedcf6627d140002
z33c96f9052ec0f14570e3b5f828633967b58c11c657bab0a449ee587c516da058f8f212e0f9c7e
z372bb285506d202465124ae2c7fa1e87587e95e9bdabfe92392a78143545bacf988df12ca0313a
z3fce1f5f144fc07f10b82af7aa15326f0272825a93e51f151ded2becb0b5b68f39cb0b6bd96bd3
za885036d049de776685cd5af839de6f5ba8d1f5342c44c4a13ce84c5924cd7e13220e0d7d724e7
z397cdfb9a9ee02643b96123f96b26d185169313315ffb70e506ba48b2f27889a570f794c9be4e0
ze6ce6b36503666dbeb88c185d579618421a83a26b9d4840098c3ba2ffe1cbdef9e8d09fd37cb71
z8f1ef6ba8b684c3e684f5676df62ced4348004384b039720cb3afa7924d21fb94a70b05d3c5fd9
z2127ffa51663c8d33438c6cea121d3eff28805e04371bb413ca7e8034282bf20975c591b6ff783
z17fdd84ac377980d86b17bedd36ac9cb5ae2d65cb4d179d5927e65e02565d0ff7a310126b599a7
zc4eda94a56915223ed9e3f64a58278179ee4fe4a2c4972316a216fdf69a7c501feee189db64c36
zabe663f2d4fbd23038616e783c4a6cb0f941820a61356891d2381e6d1c8b62d3acd26b4ec2b591
z9dcd098579ba11b6b6ecfded1d721bc8dba799194863c5fe932dceb991edb7226660a43f361e92
z7386cb9735837dde2554c529e85697477eb2ac9a0f12e90cc3fc73ca0efacdb4458fe33b5d3caa
z797846ce1dcd3a37269f5542371be36b1ddfae7c43c81902170ee6e945c9a27bfa41b79b7e43e3
za2061798ee62921ad4f33d74bbfc1e96c46fc47b798185ba1ba288ffea06f317aac216debc644c
zaa620815b4b6d6967a86cb9d8562abfdbaf2c580f470ad507835fabc9bc779bb8341ab45c1fd28
zb8d9a860b5797ea29b8412172feabfb5136a76e7840baf0ec60cd36d2ed4d5ba771cca17776620
z243e5977cf735d1a17de2f75c3dbae9ad2f9e773fd2fb64d84f205d30b06c33ec89613dab1ecb7
zf02e362948a36bc43def747705c0da6736514513226992180cec628a7d36aff2e24ebb44c4203a
zdbe782dfb2f6f0d49d68bef9e2c63422869bfe85ef20fc1fc8e0900dc0de9ca1fb7f4a07d28aa0
z3d38038d47039047d0cb1bba504346f1bd3752e52a07b05a0555e2c98da9425c2dba0fc513e629
zd55dc758c48f24db15db40d702343aa7222e929fda04328003e1842cae03e3b1228819c276c83f
zce1b11237c9d498ef3d678162becd74c411a5c209360cd1b65333b1ac8d8a4167b949813cf6124
z47ebb3610b7eae47c2c83f78a25c75ee015605f1915440a3273422edf1eb52195fbfb05cd82962
z2efab58ed21406a9ca6c112ca51f84532d7eaf0ff69fe6c21f33404f0e08ce405e51916a9bbe8b
z11e9ef902d09a1a3d5b67048017a2d2b739bce6d04bd73b712ed90e4179a5fbfa48cb6077b4767
z7f09cf7a7b54f6c2129fe637ddfc2eecb5514102ea45c9038e03286e6d9d4500b68d496d097cb8
zd083e4701a9ed5d16f5b7e02720fa58b06f648067671a977707ea51dd79297a3e0fe09a49a198e
z09455d626c697240cfdcc37da23bad9bb11485c2f35ba8df2d116398631f0b6a9a13e6960c8414
z8472142b746249ec508796abd086d76f29fb77ed63cfd99214ddd245905aa286364e927fbf2d14
z8d03014c587a66f8f6805e5c5ededcfb589b314f7e389b150c0a59d19162ae96a6d3df3db6c05a
z4902d6231f41cf26301f949bcb72b33ae506fc20aecc47bcf04a3ad1c7eb69d8bc28683449039e
zaf1c0f143bbd4055d6fb70a31fcc8a368af745611703cc0899a63f62b77a7068cd5ac064973265
z38f001e19e795ad0768c326e128f343707b8d6a58abcddb87e0f08b260e52e89a8239348b0d539
zfe4c623c59827423cf5c775279edd137e62c8fad6f3a2b92f07646089e75c4d794517643f2f1f9
z74f8daae19dd7c9116ed77c039a09816bcda3a987bb766dd246785f0bdfa0fb8ed157cbf0285e8
z7042b7cc1f91abff102f42dab9122b268bc70cb94cc0c28637f8e21b8e2889ff207019b8d6ad62
z0ee2686d5ae90d44e3278f24df6abce3fca5834a8f6ed157e4834aed7b29214af950843368df75
z6dd486a284a23a303e4d1ce83d4ff5d8dff259ca4d89c3659c744eeaf2880a310786ae63ecdd5b
z6b0358fc37a63ff1fff2255e4b504244b1c1d7f563085583731c333238e3bdeefa2300629c1f1e
z609a2ec2dc6128de19d7a7915ac9c037f325c704825d20cab4e127b136d4cd26bec4864ad920e6
zd4744cfd0ecdef145b3c0e0dff55f624ecdf48fef4ff030289d27ddbc976d7f2ba3a6ede1da089
z857f56ef13456005b60259fe4798166e532bca9872b17723b2f2ca7bbdc08da21d23bd737ccb2b
zd5adc066729f878e88f4d5515fe196cbbe048de166b748cb6fa259f31278f3f4878e60f566950a
z6090a732b6c62d195a9bc76b9efb6bf1cc2a3d3dcc5e1d52687735eee708c84e7d8dd0656ac910
z6415a7a4959b5d0121257d2129fa06a2084d76e69fd24d7a017d72384f16b278fb94574adfe8df
zd97c529b7a17db22b78f3eb440950f5d190dce99a92b76b041e8cc985575c8c59e21ec2a225746
zc316628811e666d4f556a9175d17678027a717a03872bf3fcdab9ae0827a00f136dc9b8ec7d48f
z149d47f3b9f0db01473824321ed6304bd1211d8d7a9a44d8225779712003aebb883256fd1b5c60
zccf7844403c077c6c3a1b23765899d9b6ee519e3427f12adf5e7eaade2f65a8cb8edcb078cd2dc
z0cc16e9ff56dd346c1dc17462eb71ced7424afbcc48d8547d04926179ecefe1ece66e6637f21b6
zb0817ac09027097f597ac6d2c537fe4ca000f0571b44ec957208cbcfc679c4edfbcf9c8434b541
z418d05011baec15d001afb66d428daa42cbcaaaa2b3c9d1d7c0e797e51946dc76f79d12789b669
z8a61894c274835b087787d70250823f5e5cc616639aea632f6f2b31015b3c6dabb8bc66967aa84
zf05a2ea7598935932fb0dc2be5556d25edc129d4c625a9ad74eaac3cb762fe019d078ba2ad061d
z8aca7e1c5b76f97ec9d8845f779f36762f7b0d0858c8cf0f3c9b675ab6488396c0d145f50eb997
z12d7077a856a3b75ebcda40caf6dea28e8c23315d5ec4393a421eaea4bf51160131c718f7bfb4b
z2cdc74ff4e37395de3c9fa94b6f45abb22a3d39b8328b93057db2435d3c563267e7a173023fef7
z455927cb4d5a9ff5373a2ccff0dcd272aa1d01cc32df274cdee12edce62f7116349b8dba446269
z1b5b9d2a5eaf9864a6cca0f31dee351a6615cf20c1549214452e1496f70615a44b0db06f41fb4a
zbd97118c61890501f902e986543233c6c9c67fec68a2e51c390d74947a9a1adb8f24b720daaa7e
zf90151cd8af9aa7a05704547d2f62268f3a1bcdcc3ed480386f8e7665dcc24ddbcdaf3ff0d8e1a
zaa10e8fd0f562b4a09d7120da7f22e4f108e7cedbdf3ea808ade2f3945e0778e02e565418c19ea
ze92709c40f709a2297717536dbd90fe5c18ee05204e7946ca04609e4427e8d7df8c146e9c51283
z3bfe2d9901c6c103bbf40aaf9f69bb7c3b38aec43a6db2ce17826f8bc9e2c822992c34a4596278
zb23634c735a0ac4e0e419f7de06b421aa40a7c0868e007fe60d3b64ac82f7357a8d6bb457b1d1b
z36304a3cb4200c09d59189bc20b1b8b30ea94d8721031cbae85aa0638c2205412b1cd85ef859e4
z510019075ee6fc528de464dfa10bd0e451761e7b113616861e352b7874ad5840e56825684b1044
z3324b1739b6da60ebcfc7128b2cf3a97c85230bfc8dbf380323b8d1447417ffe22ef9a1f2c21b3
zd7ea724e11972ac984abef3d4bb68870ce4f924b345a063a6e4ced8b3c0fe005a7b369fba13bd5
z3ee4a195db1d9a6693409ba7e82fb062507ef6bef542b9943a39f161bd8681b5c64544650c27e7
zbd4285a84b0032b150bd50a49c3f299b2915d5b256131250e3d6751df73c642841891c46263913
z8adecffffcd8ecf1e5861d062112fff97cdbf7fbe456da6a6c556fe0f57b4f22df04f812215906
z46bdacec80a1f7a57650cd91c1f50325c9310368542a9cd19d25a9c966da040981d0d6861c2ad0
z4dcecd7194917921caca93fd37c9bd9dde522896f5f584f26149ee1bd11ddc0c3015063f9c54ec
z6b615b81bfd75b92ee0ee982ef8e818fb7c0115ff13047ad05d428652e2234d11122ad1bfd042a
z1cec57d07e6b11e915fb89f07577dc1789031eac97fbe953858ad087ca56ad8d647f3585407743
zf3ca6d7951111212825a192187062d22db67a954ef9a970e47e0c763e1a8b795cf5a28cb01aec2
z6058918cacc2176958d0143741df6d1dd8004185a5e4aa169b2b8027665540aec817352534f819
ze2a9bc0c1f7b90ebc387695f8380675ee72a89ae1bebdd00bfc60637c5f9fc47198aaac388fde0
z4b3f44e598512ad279fe884dd1aaf25e277c3e088c35049de0e8fa4d20ef7edd939e7da9a02edf
z5696e6d8dd2c7aeaffcb85e43d806dd61b6ec6ccf6fd8885a8c5d5afaea26fc03bdd918ecfe8ef
ze600ac54faafd9f75a1fad588529ccaf6d8b50a9c30a3179fd142947045d7381878723a12907de
z3fa9f8403f9a8c62eedfb47480aab42eccabf755cdabbeb597f7886bf3c2d03a591b53593da38e
zaccb1428c776e370703d432361ea169f1b62f113a2bd47ef1b15d753475e8d86261c300914c48e
z4fec11fd2d50fcdf8888c06e1a112d7f5ad9858f1f8cc9d192937b030063df3d2e25d13c223553
zf4da4900b9ebd74f548954d8584c85d5a8665f300e6745d953a306a5f52ea4fa04403b0c8fed5b
z5fdfd27a802bebbb1e4ebc95b0e9a1c8945ae81cc8aefaf920ad968e9988c708d8b9a3860de0d1
z7db3301489e8782b284f1d58e0cde3b82c792233fbf10bdaf29554f3463634aa9857532e150e50
zfc86791b8736c2e27fe1c8f56dcb4d3a743b3c6f820a75c8c43df7b1b72173e706d44aa9433fd9
z2275192ed8303fd021c2e4992415a08652a0c6b78d54f89ff52c1517bd0720a2051a1f53ab1003
z24cfc84c551660174f84f502768e6078205c779eeecad5556d3f68bfab9292c894129f7f245e31
z292a7c940e21f93dd68a52ec7c847a36d3e6447b8a68f3cf8a5a832f666c16ad8f79d568c829c7
zc5dbb3a877100f0619b5e819c9e6bdaecde44263b2e1b1829719a45a6fa6606cc34d1b02b1ebad
z471359693c784af8c5a099767ae055741a8729ed356a07548fe67dfc51687345afd4c4b4087b52
z7a7003dd90abc9199ecb0dab68d2116e99597abd938167b8ebc857be1302233e5d16243489bb80
zcfafe4926e7649b5e08db12dc107b38aacfb16fd47533d21c70dd400e2ecfc94a6f47553291a1e
zd11a78e8b80e75d7033f4789b642f6688adfde2823217fab475aab9c00d9baadb782c9555dbd2c
zb77037ea741582025289c02fcc77ac8baf342c72932c48b6e98f3700647e359f66cc5889e933f6
z30486bafe062d526914476cf46c14e5f22d2dab57bea098f1dbc60bcf06d9258fc3c201e42d54a
z6008e37f0fa01e20a848f5795ee005e8867314053886d4884f7927ca4e7e3524af28398ca5cced
z599c660601aa4059de792c6b734fc91cec30dc383cf75dfc5a19977b507a7a1bf36ee22e13fe4b
z7c43b95d7d2e1f5cd68ca52b72f143d9d9002e85924b6754e376036371d2f31353e2a96289e338
z2b3f9236d4e91c98a6eb31a17e0d9cc6c9073a8bdd23fd78c1c0c0ec00a2c63e4ce67410863eb7
z347f3655cdb1e5c30cda702e5981d43e3f363ba30a939d085ac1e21005b0c02081e526e55c89a4
zb6672f2c8345ebc959ba2d587cf0cc7dd4a807d3062c366442dc169403c4c80b50bfb5ae763d23
zb6070b685a27ce734405d8b0050cd0fd43040d5013b626c1caaceb60e770eb60281f234104fb04
ze471b867c3d172186d555bbf1029fcc92cdf1abacabfd33a7e0c0a8df20c39c336ce7b1ff6672b
z20ce734bf2f6dadb5515c22bbf11c3fb0ac0ea3b42dd605f06b16e174b48956c4120e19d15da79
zb3f9a7bb4f9ee4ef9bdd56eb9f48a8f922a3825c94c4c93721762df79873dd6033e4212600676b
z0c1fd6b1744f543dd92c7583d7344491e0cc7eff24495bd9b26b50bca0e62460ff297b6eba4966
zef2b164b26320cbbd7d908fd4428db390319589be8a8433a88554b98136c1b9bb3b1c98965aa69
z5641056d94a15cbc8d94c52bcb7bd523ccf6bc0cd6b10e0239e245f1dbc20a771be2327e5a2a55
z8888a9bbde52dd0332b2c807386860a36e792ecfd43d9196a1d55061276905b4185d04d6df67bb
z480af4eb9fcb06ae8901554f3012c5fd30412597289151228e709d0bf522c4c4eb14ea4ebed596
zfdfbe84af715faf7322f63e9630f37a0322401900fc9135f2bc87c5ff3eb0df5c66e6387b3f8d3
zbcd4194602fdf122f8234ac574aae90118d8a5e4932b82f3bf1eb988884a51bd1c5498e0ae1230
z48c963dc1853272d6ce9efaf9f8e1fedd37d61e86e89698afdba71ea199257b4b66c4e04168d9e
zc8dd296d36d430c42f1892ccdeaa5bd56cf15b4486b2972837a1d520f504c3340f08d577a1b391
z09e2810c79d372c561eadc2326a5b09fa9975f03bf06d8af0a163dcefcd75085fd3467d4edb01a
z8bd119722b5e25e833fe3a4895a51773ea930a522e60f414ba879e274f27ce4434b808f3ce193d
z20c813d6da05dc51725ce82a05615402b7014cf49c88ee65ea97fc8cb7e87695d74088ba668331
z394eb09997876cfe8b3f5c01ad9308e231cbec57a4e1c36f833b9083850adb5a1951c538faf994
zeab73b25c0c6a05e92f8bd74693b1acc8b336e8083c2f27ba0cf6a9c63e304b52ed66b056c6de3
z3f103f3b57b33311bfac15ec56ad4092be25bdbfb0c3c60db27e23a1667d47d2816f451a87d838
zb485fa4be4a3e3bc4454633b2ed7867da8686edbdc3388396b03f54ed49d625221e18bff377fcd
z808ecdf9101438bd1e4b8f5470ad3e3708e42aad2f8badf148ff29c4dd90d5ca5407024a321735
zfe5e092f22e433dfc6a2ab4fdde004abf6a0432f054c91bdd457c039298a0f07b30943c67e0403
zd79cbdb6a26ef6c714d2d4fa000511e1f982e52813e7988baa88eb80c54d8527804245689adf9a
z23d0310ba11b14ca9e9ab6c58a4c8ec0231829467243543efdc005e3d78a87385359fcede045d0
zea66f6cf9cad57e215ab681d464f1b578f4019784691741991bec02bfa8978a710545c4d0a53c8
zee715693e86c4e32d65ddfea1ddfa3e7840bd020bbd579b43a6191380a675dc10b0c985106a3e1
z18a956c31870602884a8354281b092bb80453de669652a241987d3e19e2d2daceaf786361abca1
zc8f9bc65c64f73b348e0442f000117c88f237d47de8ebb0cad0e52dd888d5ccc70788b57d77fcb
z42841f4b2a23da1746fc9a082f7a83f3fdfe92b6154abf50b4543afb44b31db7bc863842b28525
z2a71de827af3958e51857191865e3435cfcd5929b86d0ed5e8d9b259be8d3d946e84b4458c3077
z4938eedc97789318684cb9b7c4bc8d3cc5084492168e42632a78e2a4a9a33369cc2224696a09ab
z361e54feda53b5f5f5ab8b695f6fc991ce1dfd425fcdcf3d04d972db33f059f8f4571df010a38b
zc5fc58e267bfce79c2ae9ef2cbc36fc8615d4a89deac5c810a8bda5290ee0dd6f9ea064bb1570f
z5fb390d08a4b2962dde9031a43112086b46ae4369c7f7d32a815ad84e37d0771521f834d4e9d39
z6dac5b0c0e6168fe4b7d31f1ed53d8077f5afe9c834eb359afdf7f55335227a0643a1a8f157717
zeb3e6c4b05075fe41d1058d9f0825915bd0590bfe2f76c8ecdbe4873cc8466042fb4cd743c4e24
za4cebea24c13ae43b7dcadddbe25a4c99e2ccedb7aa8b0d0989127e974e5f5d6d00642b5c02236
z931701b34e6b22372e459b01e6d8f2466da667a0fe8474840d67713904925adda551e2eda3efb4
z1ff8ef809902f8de9ebaa554087e751700603c629919bd93d174ad7a2335620bd5d568bd67732b
zb1400d9c98d4153758bdb745c8023e4b03823b9f767e5ed2675b4ac36a3ebbb3047b7e770124ef
z9e80cf1c4d7070ee5753c607292a198506fbf80bcfb0891ecfb299a5d5708192550f2df9b66491
ze340096c6a31c65c49df65c37468a51fb00efb60d94fe668fd325e036bc9a0b77087083b2c8358
zb25da6739e22c12ecbe6997d1c8065399f364cc4ebcac1e8ebe73fbaa1edb4c4ee53a4e69724f0
z1513a03e74b639b8ced1051a6f00c33f10468b22cfd2b817e4f0aef554d8d8d17c612d27c39ae2
zeebe5ee252824296ae68ea50439042c8ac87ed142d9ff4281a95d5dd948307190bf3391824b9bc
z8378857cc5fc428d00e410f500e7dbd26cd552df43c9683bc8a972fb4dc46a7f899b6c2335adb2
z817f4491c6e79949352fc12a6350fe748bd6b8cd86e97f7fce9253c80639252fdbf7e468cd6edd
z1701cf4cd201acc397f80c7dce5b5f768daf4ef100b2a6b82cf954f748f565c4400a18eb26ef72
zc779a516651f086e9f80c48abf77261c7282ede4a570bb1106fd84fa7ae7aa06c45b19126e45e8
ze60b803bf089fecf619b5e7805cf88c0ffbfa420093ee9fc15d645d85d0b2a3face341b1c4c0de
z75005d3c23bd076113d064756c3cf678b92c3fb8635599ac7b88469d96fe59c730abc92e8dfeff
zb8ca5bbf2d9d64c290f73816cd54c20c90a4d803332c733aa8f40c896685cc0e62334a4097a80b
z6b207a9edc9e61cf6d13f85de46c3ecf05028b672a79a54d4ac16932a87c76c438005192bd729e
z6326cf45c3a051ea171ff57753d115914805b58aaf507ef0f9a8bac9ba28abd016a756ca1d660b
z802d4ef1aa8c4d853739ebfc122de66b4a3898dddc8757eca896372591b2c6bdaaad60d3227a85
zf415fd500b23c99c00230300d16da915852ee20359c729cfd1afe6d4b1efbd6152c4215be56d4b
z0a0a17512e3b5a93361051970c315f9e4c77dd6ef8b01a7c7204bfbb89d8846e14766d7219c0e2
z427026230119faa88e262ae5e678fb40c03aa5cd4203ffd0b3520e1d5720612729f988463cedf0
zbb126745c4c0a57f56254ac49a87d3e2fcacf81568a96c9ea355b806d211f7604332030464cca8
z7394bcafa0aa8226729eb5482b9e5e2a3020d520b3ac0419c259af285452e755c1756d4b3b9302
z765b4915bd522dd3b71b43394b06ba1ce38f8ddeccd88363d09b0370c53bee253bd6710ae1ae29
z80935c39234237cc935038b4d505e2fb1ca3c5ace46c9a09869bdf6115594d4686b737f1816533
zd0155209aa929b32076f41bc30d25b22b0eb43f890b8e09fba5b0af8708c5f44fc686ec06c7f35
zfaad8f21b49bb9d3a54b7163c165c229cb2a39cf5484494ffd704ef4aeeada0c91f41472a04ec2
zd5e4bd21a7a6f45ed98584b45cc8bccb2a0c917ed0eaf73fbea1b29311db784370843943297b03
z23f45768140ff4082a51f26477ca74a72a35220d98b88f7b1a5c8db168166206ee643ebd32341e
zdecaf917ad9afd48424cd0329feacfc31fa7afabf6d3f7262ca9507686601cc94d6700d147d20d
zca440fdde8aa4d1dcb60ab67fd28704ca77b8227164fcbc2f9078e5c3bcf9a7e9e7763709392aa
zc53045d79a3b4f1dbd9eeb48d227da2b8e82e226892a9c26482e40596772dae335c15c291430f6
zadeff428cdea6cc4bbdc2a2e8de0881e547c9f2b98ab43c0f9d545bd9a0c17fc0a81f33da4dc03
z9916b5f9d1721a70625c6c7a2b3129500728e32c7ae4e46840c239f61859a716d2a927723450b5
z4d437be72d950e6ed48b667c15f198433bc823d63f5230faad6d823b4a21eeff811d7e00c32d81
zb3a9f2d8d3d30dacbbe38038e2084e0720681856bc36a1aac0a92964cab2db523a5afecc96f53c
zd6f916baba517f98994418f017806421dfc391efdbfec1eba94fbfe19d9bda97adf62ee2f8a223
zaf3a26f43ae8276578059f7494ca0fe78893539b1e6e44e92511c1dc5b21674bf30555c9bc6ae7
zf95dff27215ade83ffaf4e27a371fa22d0361b2759b29d825c6cdbade0d7730a84270337e26135
z3211edcda423011c4a75a8e673a57a3e41cefba5c7ff0600af52e2bd873180723a99436ba7ea69
z6782c312f4d1005b09859bdb199dc1093f4f493d0087e137e83a5082602425c86f998e8b715c9d
z0337bccd222cdc1044b80844973d3dcf0bf940018c5bd871a3a77e418a1cc6320d552c66f1cac0
zf14216bd02b28b6bd5fee841444714b8b443c64950897fca9f3341a706f7b17302464cf69987be
z759426d1510121943abf49a3f6b722842c6fd7e661881ac4f1280a891a6e954e4368e424e89ca9
ze7f1c3e3c7df3ef1dbac9493a53f2a42d29d1bd7f5e93b4dfb53bdc8cfcccbc26bb0709eca3029
zdc9abdc2d24b3e90b68247645acd9b3317588fda0154523d5072332a02c0422841dcc7b4aa2695
z17d77922e2cbcfc0953e822ec4d20cf7a16a5ce559ded6a4b705c44e508ccaccf255e1ede3c78f
za0cff1b9cd7b220e69b10485491f6a8771c303476a5544bca9d98d2694c7b5073e2c3e5bf9bb6b
z880726333b28f19a322151a84442b575a8807067530f2ae85cffc1dea3d2c8e5dc6d87bb51855e
zaa100f8f68bffdb3ec9f12bf6e624be823c1b9f02210967a000126c7de1166bfd3b1acdb4747aa
z46fec4b29c16ea70ea79ac7e7989383209d59d99d02ae584f8119b21df2bd0d958bd39c837fc69
z407813a7366bb221ef9789853a2102e6c221049566607bb2cde24480d30c3ad1110b1f5c1432f5
zae81ec865a19a8407985c13ac0ffa79239126725738f4f98915ae9f02d67612065d77ea9b59c8b
z137a8cf58af8b7e646ad36c2562b3bda75642785ea124e38b678c1b0fa881c45233c0956078e0e
z117308f81a4b59ab91d4105a8ff185f52de524dadecc9c4e55cb3c1218198cbdb19d6720ffcff8
z5844a29cfd64fb7a220219af7fc760311ea7752877b8092321312bc80143c0e71d5b47a801a1ee
zf23dd9dc529706a537d23b82d70dc58bb4f379e38a275b7af13575ab0af131d3e2be6d5729d20b
z3471a272e23d22d78d0c43a07c281118455e8491159004c910100f98970da1b2818815a8629120
z030cfd0ce6dab4fa79f83845a203d3efe74b5c787b650c1659df651121d0687849b2e3e8ebddb5
za2386555010d320fcd5693b6c64a72b8cf6e5f2ae99ec9ef58c1a3a96b81a1b727161080fbd518
z7df60c154d9f911e39b9a46df520580163dfbfb4b333530847f12b37f052741b548a3c8d57fc5c
z9b0c5ff345a5232678ebbaf0bf390a2b1a1a34886fec9c03cb3e48434e01767f169aa294d672c2
z73b20c70055105cafc8882e8c28cc0bdf86a89a5bb3b74d277c7fac277028de5d948adb9ac21d8
zae8c14b1650454e9943312f72749cc13aa719e5fc9db97796673323460eca918ff9e81c432403a
z5e68599fc03a2600499e9bdd95b1a1d50ad8159426c3c3d58bf3841ca987a31333a8dad77a7fb5
z59d749e8547a7fa18a8d312185f6538224021e96b598cf7bade733f3b323d054f4537dbe80723a
z8c30f2e816121ca26d4de7edf6653a9eb96ee6dba5016c4cca9b3717dc0fa9752dd4ab17cb94c0
z3ba9ed8aa4076d8525e07f396f4d702eba73e450c8555f96e5d83c09f488c177e59387fe0dc759
zf885f420b2969f41f2866bcafbe1edea7c9163468f79980afba2e94b0c261dca1e4cb73f3df435
z939a1d19427bd3eb14f1d0452275c28e41a380bc13a9b80d3317bc78cd4ced1f6d366afe7b7d12
z72e1997eb8ec023c9314b5002c4e8b2cdac2d8400ca87315b8c135c8736a171f936169fbb18f4f
zfc6650972d483d73b0671bdedd268c967dd289d16e1c0ed18eb45e0856883c7899ef25df79e2b1
z9b1915af35cb5a9f34459054cace6947f6e06d42de4fba6dad6557c93a5ea2802f301de22a7cbc
zc2e00d2e77193ef8758ee9dd75270c6eaa693f7eaa82edb8501e5e40c3fa5a794d0bac0b4d5dd8
zc4d1cc153e6b505532a79d5850cb8b93e9d00475fe1116e3fccd10e152aeb426c18bea31df5e81
z2fbeb29e643110596292592a38c3b4b96864bbcff121c46172a3a25511140ce80edc38bc4075c0
za88e1127d4a5342d56df5604df0202f4ccef78d3e656d340f18dd2e4c272306ab05c1b1a28af0a
z3167d4331734162ab034efaad7dd8858c5c0b36dec9589fc7f5fccd4e04a7208d42ae57e346fe0
zb2c85496de472bcc8f4ed11472815d7df3f0a822d08fb2f389ccc1b2a0502f23862f1f35983330
zdc3494fc8c5ea5ad659a3d16fbe6167cd1c6ff100fa197a85142a504479995b403e2e130b1efe1
z74738b71ed37e157cfc2b8d5895ebfd0faf896938d863f1acec16086254b8691dd22bc93386aff
z8ddc64a14e7f1c71a629519d1332db27a7dbb704910ceb1f24a50d61d2d84fc415ca9fc76046e0
z44cce5e0b6326bc3a7333b81487c320fb9cdcbdafba3944465c2886a85fc71729a6055d6a29e63
zf961ad3ed0e40052c628a83b65d5c4957e1f17c59300970dd6534d6f68aae53b01121eff318278
zf8aa8bda3dea0ba1bfdc2c1ff78279fa2cccf355f33dc423408729a73b4b17b2863bc709798ca0
z9c0a86b823209047e1c632ad2418cbc00cd8cce593da0172e7d304e0ebc306c187cc53ab1ce23c
z65959ffa13578af8b9019981439bb94e4523e11b50b0b44cfb462fc9c3709aac4af259fd9e07f1
z077fd51a86376c3fffce5cdba833d8e69123a1f55371c968941c417108e23c6f5ceb6009f3405f
z8d710643fe1303c1bbf27c211b9464dc0103d44df31ca7b6182eed17e78de240afe752cdcad406
zc54ad4243abc3d2b340d8fd07081ef6430986c73105d5b6e1ea548ffb057d3d8ed91ac4228af75
zd34c6e415ca05a65d4ea4d80edd81e0d2e7491b7ec633d82e9bd68d427ebcd17b0c05176fff327
z5fd6da4ec2743e17a8cbdad7cac5671dadaca1778248f96cc76991c8dde0f234904c565ce84e81
z4f4e6e0e5cd368a3918f1dbfed5092b2e3fe427eac882a1398646687fb077873e5980a191ce327
zf716348e18da65e937377f5236aa147ed32a01b3b6efee7ed7e58c4918626dd867a70a52ae8775
z4df681b87de694a12f3c6433fd692c711620f3f2d2f529a1d6da25ce00c45f3d97e10f41dc9c17
z314d8385e794e895ded9a790b5d738c38db1d7046be466610ec127e6821f43ae0e06af415f0943
z676904befcf6f13083af0e3ccc7c939938e870e62338bbe2ad95535938a0c53754c108e36b9a95
z3e2a1aaee76067d281eb3186455406be74c91cadeacf69b0777897c68d6f1edd5d5d5c93a7b61c
z5da59f5d00da9d511eb39012974362b008a3b601a3bec6296219325029990dcb856e5b2228cdf2
ze393a8608f17f0b850cc0a86f3db74960bd6a3b14b70c168cec6eae2ab81db85ad08dfdcb18194
z4a3c4acba5c706fe78b4e26a529d49a2bd1cfe34100bcf23fd93caf9c2cea6fed8275752456dd5
zc0a0ba96431ff8cacce97eaeb733e6bd8dcc20a0a82d69e19c2f0724da3888f826fabf4b2b4b68
zdc1d70d893942d54e3a46119ee330c1fd1bb6c6451f0e72b229ae93381e75fde221e11156cbf16
za47a90f51ae0b6b7d0c13419a2376d6d48c5c076b9babea3b98bef7c3967c5f5c15bc5103efb89
z93043c74baeb014dad9aaca840011d7e4fdfca6d6c86ebe0a9486c0740b5175f0bd3dedd34ae69
z4d4078e580fc625d0d68db72443fe661387b9c0953111f26c98e97caf843f2b27fddd70afefee4
z643af63cb18ca3f52d2805cda1f6ab261313bedce55289ed2b103b4aa365ac0ee8c3a659ecae1e
z5720e8aad8cb7ba85a4ee7bcf3633a99253dddbe65d8136bd16a15978d34f89ff44b0f5c863cb2
z9787f6e427b34d5bed9a0a4e1e62298acecaa2577a7b1e2b127f2ddc90fc0afb64efeb9c40575d
zfe93efac36111ae71f5f1ef2357d58141f54ecbfabe59406d5cc00215400710da0c3591d4d2418
z77e9a5ae3f25d411f003024dab7fbdde7c16856203e384ddc20da5170f0ccb2d0801533739d4d0
z35d158e45aa8d7a49e245ebfec905ee27c3f9cede3629fa358ef7267c997e78c7ef852e7696230
z3d49fb1c18a69e50f0a5dc5fe5c3244dfe2fa7bcfb838ac0b825c206b5c296b332172b1a0dfdf4
z83201711469a304f60d95221838c325d5b5e840fcc6d8e42270db1ecd5eb5ca102ab71a8a49782
z2d94369bb06e30e1bcfd2efbc637f82dad348ec3357046333198c49698eede1202ebba2017e68a
za245eee48fb661289eb4c561de861bfad540744b636d175a54cc065625c83f6fee37627b5ebeb0
zaffa0c16e1c941591945020af0baaaa9217a313cd8b32f651a2a9456d347885e688c3710b5ba07
z6c6fca0a96e000e048b4dabeb71b636d0c6a1abb26b8c7db2589b27c1f9e514b918dcaa546e295
zdce77eae8b7c5e1b64124d58dc2d7d569f6dd6b4825e7913b3a3abc39506897c2afa95b8cb263b
ze87543a1d53850d8e525fe836d1be38532a26c342626d67456549846d079aaf1c08ffe6216a8cb
z5f8202883aea82ae00b9a83053a96a170b36b9cdf1736fb2087978100a84bfeb092107486f42ec
za74c60a6fb6b46d0ee4bf617b9c3b415bc8dd2da49c0cbc68b51f1df33635d66b208566c731921
z365108792a465c5caf46b451931f31d1d1050087573c2702c739db242ff295028c2be41076dd39
ze48316f68978f3479bd41db93b79ee33902e76662de84aec345b30efa485583f71230c13e8481f
z35dd94ba6968633cf6132c8f788cdf242c4dc7e2c0f2a75c6dc6401f176e2e5d98083128cc961e
zbf051253abee8969ed6cb1d4f6ef91afab2732bca3d887f547e11b054adf5ef238742c4cb947fe
z1b90f5c461b40c7a2ae5f14093f0943cb52ba9c7aea01936bc550d5efb198fd67082de9e87547d
z79114e36a0e2bffe1c739e0122c46561c8e3fb0f498ebb68c75d7de6a81a72454a67c6b7050f5a
za57ed3732ac7c207d6124c1e72551344b746be4ec29ed0a0c4b0ee0940d0caa7be10b9bf8c4635
z2643e16690ac99d0d30d47251aab430432d09a9accc76297fc873ecb13bb0972cf014a87f8ff8d
z3bbc4fa9bd8f5521f10ab4dbcaea815203ba8b3aed63dbbed06496d722c2835f8773b68246545c
z12dae4415faeab953c7eeecf7cfe3e5345d6322917442225354bba117ff10e58bad179e7143225
z9cd967888cf59b7ac63eb27ceadb9eadb9f130a86ea07898d7006349fac0af4ba89b7344c2fd5d
z8112005bd81ee377df14f1a3da2f327be77cda693f7d9d762f516f34e605ad1515a9d0a1bac73b
z56c2861564f554084166fc5fc71cba8d781e1ff42e90cab4a750030522621f97b86efaea05369a
zb15c4e9b3565a8b45111e6a0de8334395bca73e88a90d97ec21075cd09ab491e4ce65945a3981a
zec6d7960ed43b7e6dbc00b10e6129be7c00f39abdc3034765e254e53a8d4ecfd46c8c95c79828b
zbfd7fed80d1f79fd8e7e72262d926d392eb08ae98834f07b5110c02c17893e5198d3e1bcc76dae
z2ba9c569b66da652526aa9693083eada2b9e2763124430b8bfeb74e46cd8c543429950887a13d9
z697dbe69b660de08aa552e22654feac84d52a4e5264db962dcc6b559117475a925a6f1be085588
z8779486d4826de7dece69c15f34ed08cbd8439d73f921f3efb83a16d12d7106122124388a39eca
z7e8b98640af2f67e675503b0038994de92651202326abb139cf0651014f535be4f17558079c222
za559e89bcacd71c3a5f7e7b8f2b5e14d8671b9cf36346f4d71226cd17a2ed28e7fc5eafd83a43e
z091e7ee0eaa07af6f7a10002b1257d20d1cb4ebfcba01265842579589af561e8b5faa0fd673353
z6663f33909d55233cc85316d1cbbd0456a5c806a2f4230ab13e0c0cdb5ea44801d730f89a3c301
z59305f25eb4461735feb6b109260c115a355377c75b12be620ed901c0a3605800da154ed7b5978
zb767d598b71c287a924d6ea0b4877b05144aa39e14b8fe84130782f10d42111b28bcfe958ec51c
zd5136a8f9a5591a6628c3d0aa633db91fb579d8716ed03cb73566fde153e34ef5726a95e75393e
z1282d16120901e1aa0d6342b26e24c929cc1f89c1ca495b57da7968feca33af940dcccc1edee73
z03849dc01101fefb98395ac00cbc0a78b62e59b837d2f07e0e4df107dfa058b929a0ef0a4e3914
z0d96f908e17b6a80944c1f828c5bacc86cc8c5afdfe70e552233bb316426181b2c5b5314ec0488
z3dc3d4ebb5b8310d2b230ad42a8d4b93457a8d5ddf646c77b2337552f8b8b19cfcfe55ce60cef5
z8dbd88c84b9a55693bdef1a7c1dfbdfafeb506b558133ffd29acfa501758fb39350712c6689979
z53504047af807871d094280440054171902de2ab922f3a89e482851c8b14d32bd3cdffd1b1c028
zb8556c72fae460606b962f433a98a05f62abb53cf67ade7222b229035de6595618d80f83385c93
z1b7faf73e301f5e834bb5b0461584b619262dd67569e8f41395607c3d429c349c8c1be0ff52625
z2dccf0f67f0160b235190578ed3399db4f843a5bfcf94bfcb83767c64cefc5fcf1135c03138ff8
zc731f1bb88ce75d2d2abaae22e33279fd2d2a6597f48e0684dc494674958946a12656fe75d8964
z6f85706799383318271a75a23acc52ce5580bf34631669267e2d149842cf4dc6e115afb2c328c7
z559d77f34c4f1502159f249a6432b73fdfcfe03fd89edb05f9b34399b2a2959223dba7a2a6d757
z3a722ae94f46302979b75775188995ea126469591795f8f5e5815d7ebea1bd56c6fe2bc2b2b9a5
zfb11c1ca39d0cc665b4694e69a35b6d9507f42495733a9a4976b247375d3e562beb88c2c3cc99f
za8c3781da7c51cbd9cdf920780444b6b43f8c2bba18301f7e805da8ec90fff760fd8b403c59827
z8cc2f983fdb2ff7d3a83472de44b79c0283bb64b55302c83b4e9e27f4968981e76692701a051e8
z782be45bca18eafded03709179b19ab314cf702a965f4f1ab5a775fc94be35822305a1d58b77a0
z55ecbb3b2b853a6e24fa1cb8357fd84b8b4c1ceda791deebeeb49370293c14a5470070c99896c7
z7ecf0ccc6df8251cc990144361bca390d6aed8b4c76c71df8ba7b7e6eb05a14b50940a46dec511
z433eb67c54bf19297bb90d4727a823293d3c5a65e110298e6fecadcfe144a8826c203771b47397
zf6bf79d396742da9787d2206e9c3ad4da94f3c93dc91e27229e7ef70f648946e50d49caf3ed161
zdc46daedc4ce56361c06dfe835bcae4f3a453300d9936b5597f9dfbf396de906eaeeddc4095d9d
z9f8d9dfeba118df7bf37461b98d5759a4acbe338dd48f4a88ccb432202279b655a127e2dd7e73c
zdd8bcef77522cc1efd0cba7ed8145761082c33f6073c20aabc1602991e04f4de2207936fa772cb
ze23c81234a2f07dfd5c7f9d219da8223ca478abad2cbe88f627289adfd8eed1321882f4b97b5f4
zd39b7e6693a846c735cf9cceef6091079602f7af84b85b6f4e1d87a06a8b95c36146d4f3ed43ec
z834b693c6c91aee1e566644a04e795177aa17d841439a5e5527fa9c280f3c8d032394bf2759a68
z20bbc1ce815656d6a33d811f87a75f4a0e9fb4302a0b2a018a9252187ddf2d533ecd3377e358dd
zef68537afef10754957710a1f2477d9bbaa8456fb3ed30b52b7efbc059bfafe39e2a2c37494d0d
z3874701cca1cda2f54b8d31412bb903ec854467b61c8dc79972274ab59bbcbd3f6fc106473b991
zd3fc603c59aeafbc80769b7b4f1c9e4726d101455ce30349b5de5b22fad81522e5cb25cae06d32
z68350621ae84bd73a845ffd1c0be2483c149e733ddd438ebd24ac46aa797affd3e3cbf8c57b07f
zaa1c8b6863d57ba62ac3f4e591f52b2713d9978f8f1dded8fb093d46aa74c332237b0c43e436b0
z42c1d349628252503a09561884d275821e0376d8f4ff9568713b429d8283611ccaf312e942d6f4
z23ffb76d965d152cc0b4c6babe033a3c07a38d152abc136d7851eedeacabe93dddca60923868cd
ze461f242ea072e82305ef732ae9841e5a04eacf1d8b710b84ef4c0dfaed1bd84b3dec4d5f6f38b
zc5fb586d540a03e190345e19a0e394503f2206d1ad4bfd43d5f2456ee4041b64e2c3649066a8fe
z160ea64fe3025d1b956c9ae17dc2026b22388348e26e22fb1d67e8eb3a2bb80bb74c4b4b356041
z3728ab6ddcfe6d5df61caea8203dd04003a4870c5f96c564a5349784388699fdc85e083b97a494
z3bf11756cfb9f3c6e4ee5fbb04441851e9fa09ed5d83a6cba710267fcc912724db88d7edf6414d
z5ab7e443ac98a70712558bd75ea3b1163c929cf81ab62a35d82bc463ce3d21c37be87cd6bb138a
z821bdec65238a15ac0c5732777b95b87ef139dc55ff65a7212a9132dfc5d1850ff7255d5d549ab
ze1df6b3aa2e42a3246146ba3695d659e99db8a8d229e907d4359d91662951f5f450a212747698e
zd4834e2c56a4def9ddf8f2a8f115693b7b913e7601a6959fe6c37568f151c493b51b19c94f73a1
z11717aa79ec9796fd6f19eb8cff5e25a5ae02867d1af730506c5f7d249ad28ab74626547febf65
z760fb10a155458462f67901eaa12ee5e23df4a77b37c0ac2dd5edcd1b73b7137ed687dd2ce5339
z3af532396d7051dbe377b442711c9e2c7024be659b132dab0ad1fbd16688abf4839e2474440a13
z9127e20deff480e405d4fe682facbe125d081da737dc873b982fd03221fae98ab947de55c391f2
z55bab074a135edfeeb0c4764fbe2c25813b7c3a4821827b09cf2261d72a0c74e86fb3c520b0e4a
z9fecddfc6deee819f11e2749bed98629dd79e43550391e998c678fda474f6aa7551eb6eaeb084f
z04b4eed98135ed74dc24377ec1f2ae80ff1c4ff952b100de79d12f0ce754b2673e56b0eb8867c0
zc5e46665897146f513290fc4658ab69d3c00502c5990e866aec08e7561138e6d5f844d56563eda
z6b607573bafe462b9dcd107d4cc4dfc2d51fff71c53ff7c6cfa422fc02b8f5b6ca471eedbd4137
z413178705bd6865b4f55c441d03d5db526f46953b9fb03aee6eb4da54c846da37bfe322c6ea9c8
zb506591eb1483bfc0ff078ef5c1492fed4c9b9b506f90d95589a7ea11297b8c5c48bec282cd9f0
z8d0a35618eb49afa88f89221c6cbec356010a23fd5d1864d9c7ecd1e5c970e369b50f852fffdf2
zb8d7ecfb830c21444117bfa32a7a1e46f34486cff764858b191a7ecfdaf0e2dcefc12326c572be
z6d2ac8e6a4d863c9188acc122a0190864edd9d1cffdc73355ca84bde33869c8169e8e53f7b0f22
za7220b6a7f5f10824856e4a8f10479c490634d93a2773ae6542206bb6c138543764a04cb166302
z9dd130bb780b4fc18395a736ce2f0856b4147271abd8206fa89de41a7d355e415b49925c829145
z599fb7db02f363c458f03f43a2bacd1968219239821262f8db928ecd707e66fdcf7f97489e79ba
zba1270b5d0a988ae979372aa5162246355ce2d4d07ca15fddd192f24c6a24f1447479f829b3d8d
z04ee75333e173e9541975ab1885af4c4ce672efae9800a82a9b274bcfd7f6221708b4fcd22e337
zf46505a4c70e20df95c2093fbb0d8f06ad48d7dd26afeaf1e90f6ec40f37b3874d2db5abcede79
zba7eb8f57d695185115913f2d032535b298cd913040d7be38d5e1946233a772e4ab7f2a194e749
z82200a1cbeb6f6a054e0bc2fd2057b03b0ddb7a903e0e794e38cc8c6ce92d96ac9b2e02b3babf6
zd59065cda53106932f2e8d63153c8ba068a4fc1d9b412e3478f5cfa3408f17e09bc712c2b10c30
z5071ca46d4c78c98711113a06b80c17eb7d30fbbd712682b9a724757de87793fd11ada63dc318d
z5362155ad9fe34ee7a38a906c2317cc293f5aff47a4a87b9d7d6ccd4f2198d227021f454bc16be
z07596e4922c69e44ce2f79878657a5f5714a300879c178e5ce9a417a642687fedcafad3bdb101c
z6d15be8a4ca9304eb5070036c13cd9a98f8998d6a1db1f1c5717ace96fde9973ee60c604050ea7
z07f95a37a010964f1eaf3a828fb458588656c9799cd22cf72ad9c50860bd71cb8482a6f31b612b
zae8cacf02474e83f9800b2f26806a3bf6020c7c5fd4ee3b44da7c4e5eefd44caf17902c052f479
z647bab593ce5e008cc60c0943228a59097c94d62ff6ad163f1875586c0cc3200e9fcd3efe36ee4
zb841509bdba868c83a653c271d58b9fcef9f4bfad103d525dbbfca2adc89e67f5e4b93d5fd51e2
ze8d6cde9a8981f314e827a1b70d58cce01b0e0bdc54d2eec4fa1a1fd031d8bb6e3f5830e5e7147
z1c84c22cb5d4ed6393f2bd20f566af507b950d19aacd97943f0ea6ca771a2cd30ad8f16b45e5bd
zcb497828971ad2382bb3dc599f18dc821949be730749a1cedf121073a09a04a5f7171e45dacd21
zd85813d1454ad971027941d68e77678e4f0ca5c50597276792f0c1d0ff076108c0ce29e11dc05f
zd48f8fec1b8202ec136d4ac22926f2dbe5206e0b7b27b063218e11ff5a3a55c06097e2a8e184a8
z3e036301bce2d2c4f2236c9118091f3c10d9c82e9fc7e58280130e502ee17f328f0746a53f73af
ze4917c3da761f4e52d2fb727713862b3568643624b0868d33183ac03ff94ed8be3d6f2960a8cc7
z1429ace46312d419a59069c2b123ded5aaab6f120eda0624091cf01a64cc68d81bbc18231e205c
z2dee80f4ebb5660438be56be6657943f4e220cc3665a99f29e165c485fab4ee97ce45789cbd0cd
z41b692a18da23e25557312f8e1041d5c97fd60884fa86273c47c0fffe70f6da19efb3f13e3e33a
zf7628958ecfbf2028c309d27119f9b842f0d7f0e993633044059629c96fb7b8e113048f008134a
zcaa3dbe7d9b674f1ec2d9b8070c2edd6e77c4a62cc986b5527abd927bce21f4543c3d0db5a82da
zf217eb6e9ab04ce5593959b8ddf0c2812f2cc026d99e7c06a4b679da15ea0644e5f5c632a199bb
zd941de3b9791527f121672a3d0b33809ad80721284b4af9fdee442f918201da5315e0395076baa
zde04ab3a4ca5f361c37044e3692bf59912b037bffc2de22181f67a3dfb541958b14fe9a8ffb0fe
z07fe2e1dbcdc5674fa3434373bcd07014bfa61d553edc011b9631253fc63a5522fbd0528010088
z574f6024ead79b56429800850faaac617123ce6613b92845494a5d5a009b6faca0546dac8abfb4
z09aec7c25937f2405f107adaa6609003637066b2b29826e9deb88e8ecae5393e018fb24f9c4a93
z185fff1dcaa722cf96edfa9eb83ee8aa217c3ef254180c27117d514e2da599f06af71f2c64d7b7
z10006d7b3819085fc170fa718a92dbe17fc38af2eb467d2ae72cb138aeda31a06eff0af89e901a
z3af8a2f0a973bffe3958cfcb1e4d58b448c5688fbcc6b61c2eaba32ea4dfffaa388345ac51b5d4
z290fb3613f1f7333dc17a2ba8a67cd81426e93a82f7bd4bf6e62b99aa2e4390446c9a9e6b37d8f
zebc592339dd0496b7d988aca7fb301f7a43fc1d86eaefaa71ed51bb87b109f5d54f9e5d3a4cb2f
z19cf650a9991dfa38c1cd3bee19966e29f377afc6f087a9ae5efeec94d125fb018da54eb71ce94
zf850164981966ee26cb8211759a5cb5c6aad2b6bc9153bc23cdd4af5012218282d606e5232e47d
zad2d83cb6a087c7759294d884334c56cc78bfbb78385f314cb5a182771e3866ec6b2ba450a69bb
z04343f31b5f023adf6f6ed5d80a69a7ed668523be9eefdc2f44f13842edc38d718e04bdb48eb20
z7c387374fcbdc9930bbe79bbbad50b442bae7a4d3f6180794162a48e4869e68ed6975489b79dff
z0b13afddf50af08eaf79f99eb381cd3f1689e5e35b6740aa276f06403c991a2bcc5dd469d82873
z929067269ce2bd6de68999f48ac1bc2c0acda66b5bb3904474de6c957cccd695a6992b8db2b98e
z7ecf8db80968b5cb9319239a7f318c09837b68fd5000686fb286961cea18779f7d5c4dbfcc6d00
z0e65add3e1672c26009b0fe533b8f25bfaeb2c33ac5d0c0c0cd13ef5902ce3f9cb6d3070c2465e
z2cf55b08cea425bd5a6e65e592133c6f06193223d51f7b2fc76b1abb07202e86b5c38dafe0918a
z7ec023df11a5f365b427d8c087956aa752b835425ee66d8296347e50f931718e6adf6e2e72915b
z55e42e4b8f82711869016af093db78a56fd5458b3805ac05f1dcbaf67ecfbefe9a18ea5999a545
zb21c1aa134295ff95a3a9c08ec7838e348051f4d883010fbbf57ccf0b69095266ef2e4657425c8
z658ef1b00a5015d2d503fc72db4fe44caa0d82ef222e6c93291a26d7ed5238eb23324a36d5ad9e
z4004f1460106577d182eaf2fc552201e6ba8f45a8e911b61faa0208b909eade30bea7a80ee91b3
zbeb2eda14d2bec09a9335ed7796e9223cf2083bf48321476179a26b00e32cc540d090043821083
zaed86a390a0fc542381aa55dfd46f5b4a55e351abf7e6065c871298bc416da705444e368807f4f
zfa651e3a750142f8fd8b7f478bd42478f961e52e30ba68bee5815a9c20d6376f725fc990a683cd
z30f10ae60f3f8c337dec55b066dff7bc450b29467db964b6030676fb4091b52960403cd17622a5
z411bca8b918ac26e9b64e0a80b2df353ba18abd420e7c17f0a60cc5ef91a171ea36994cd208b4a
zff8720a5bbba229b57863d049d0ceaf566b9ff23c80c36a3a1176486f9a39c20da9b977ae9af9e
z762c34c6cd005a325865c986f76a0a0d994fba3f83fba17858d4ac8dd9f5aede7ebf9b3b160243
zf4a88f6d68aaa1d32362417695c77012ca36588587e319d7966f4e1e3f58ae639c9b4a8df8a4e9
zadec7df598c55145714f7eeaafb7c35e45796809973eea76d5350d8d6c22e6d7e9b9326807231c
zf856f1d5e603c16f9a60a2a263857380357af71da70c707962b8f02c4c63c96f4b7fa1eadaca22
z213c07110dd983e9f399a528fdf3128e58a7ac916e4b80bd0ee97ffe79736d961c4250f94dd26e
z0ca21873b5fe36f52a829429fab7707541b4ca240bdf024fe2683a67bca439ed140777a83a5709
z8bf835b3009e5c8a459a2d6c264d5a85517d247262390fb26b0621a49043daf731e80817601576
z8bb43b07cbd2066ff2aab60193225116fe10c8fca9e2acc56b51683267dfd5e5191499ac9a3b55
z4089367030c228d8affe6c3efe73c7bbc5a975c0333065bbc1b0041972095881369c2b650efcaf
z6d241280aa7dd7a00a83f99c9b704ef082118e52c814fd3c318f528e4c1a850d1b25a10cb4e60f
z8fd710d1c0615d4a6422cfcae519217c5276b828f0422b5ceed6529dd41092d80bf2cd30024c8d
zb628f166b526a929e5594d790ded1dab60664d60a2af32e0041a05573b0ee1e387153d2c395871
z8755ccec8010d91b8f33b09a845c0be9b40e76835c566377ae980f727aae20b0401850edc9625e
zc80e829afafc44cec199a17cc31db48b9096e99ef47e87d3f6fa3dd18ef162a725232299ff3317
z5688520692c817d5d78d60d16dc1f1593f4e35bdcc39b3aba05c28bf4b0831f543e37e550ecff7
z84169e18565ef4c8c7b1a97eae799c67426b5aab84f3a7fb53aee5032ba2ed6e415bc2947a08b8
z8e4872e05f3b697a0c291ccd7165306c6eef003713b452da1221e5fee58f8798471508ec029f0d
z9c37f1684787183f3df4c0966e30723b9f8e0a6f7dbcf3673bd833b41e4c71bbb6caa0d16164ac
ze135f537929568b546c56f5f444d6938b1a31a92cc6d8cdbd8ddcdf26c5cfadca3d1e9a7c249a3
z510a21f85c58cadb6c41cea35306294e84d3147871677ac31271c2c39688b8953ebd0028ffdb73
zd05955c34eb5b33b2e825a2ffe83646e95884e6345a0974d10ad8383beb773350b19f22ac0d2b8
z68c21d6e0de196da6e5e33f4169e451019c2718c1f7374a6b637d5bcb993425af7617bc0909102
z644ef7c07e7560799a89bbb875c50da81213ed3b4952904c7fd9a85f2df37bdbf453df19a73fa1
z90c68e1e0c547acbe951f6234fb3b02d40248850e1bcaa598242a6415b14e0a1505d9bc0b7db04
z216bc0dc4f3f3ae560cd91a76ee2eb62e36146d388e3b8ebc1de3bcc6b9c77b56f7b33dd65f3d6
z25f7e8220438f6b1e66aa1d115fa88ebe0a1b0f6fee9b2201a9907947f258411290c3599910dfd
ze57e31d5a50b2d77aa5297a655ac376a7e74621a560c30fd6bd0fd3e79a130c0932d4277ea0d6e
z6de5ca5d0f25ef3023dee642ca8060740fb5a505b1f5a8ea78c590d9d2ac2a9d1b5fa8b19e461e
za3e89163973378789cff539d367e96484f8fc93ada74d3f3583883e40f901b7e50ca2d3651e581
z5954c18a0f957e48e2e0b35f8661767e8ace117144c2e08df4b6d92d337f4e271a4115249fa61a
z36b1ab66fa0c6785c5da20aad986129f8d85e9507016c6e700a61b4732c9984d2649f7bec503fe
z26174b4a9a0991695b1dda6929f0c62b023ccbe701f2cdeb2ebe5a472cdc1ff5c36610dd13145f
z5c3f4de87cd25a70a605a6157b1645db85956bef006bd36f7d9079207409d1a8e9bb02794f9d9a
z5e3cc3072276690df4c65e4eb23bf8e39735ca231cf35823635b8e9b42f054097be9e9ac6a565b
zd5e014acee8cd4122b3f5fecc2652c02083614e97bef380d833bd72167592ceb06f316b51c81bd
zff62dda2852422d6893c704a97ce1d2d87b5188aab13ce6486dfa5f7bc9e2eaf55b96593824893
z56a3ed2a697c83485ceb0f97bcd31a1afe99f4f047abb0f817b22875df08f5c413fa1452b8eebe
za496a384ed4bed04614e6cdb8ed49039a093903e40dfe0f208c98fcc2cbea7669dd9e515c6c397
z25ee8d8f871ff66f30827f2449929ef28f020ac38b22fcf347bf311c6a5adc4f9872a7838b6b65
z6cfdb7bba86d868e4bcd9c3d66f4dc015bee21ea7f584a783d22d3e9c0c5f9f8baf402b5f0f774
ze38c072f696b16b1f36ac07217389f825af2b88c9f7a25fb4c6f34a601d326b7386fa41820f0b1
zf5af63d50bcf320b71efbab2d6e652dec58166828c516dc54019d489177b1094c3b055e58ec079
z3fe009a27ce8d81c36ffb63b6f4cf932d226a8a8cc13bacb14ed3d78683fb1b2aa5dde577e3d3c
z7282291e7c328164016d1a9878163037e3f9618877ae0c2c0db738ea15f19796fb01c1bf17c111
z4d4ca07c11a7f8f0391bfdefb9f420cfc8ece1a536868f955355901e4bec2ddf86c8ebd0c72058
zc78c38b2ad3d0eba485bd679d12f965fad02e26def9985656e68181111a195079626ce7080e774
z2850e26d033d49b0da3ebc0a486b958687a4b3f7619726d003ecf774bfeee3bb4400aec0d2e2e7
z0a6ce4ba8a611249c70b9eddc91a9165c4b05d00b0ce85a5a3894dd416504ee0d5f09ddafeac98
z42a9493892704d3c2e872a1d4f39c9a4f2cebc6bc7ba9950ea3d41ebe0f9ae87034a08e177642f
z057365a4aba90c2a2579a535f78b86066c47a400aadb4dd914148f7fab4a864142c4cd3c2a6ee2
zb051ce0fe9e39d83846de6ea076e2be06c934a3964da76991602a26988608b71236a83ed8d857f
z40fbf8bf44cc210247bc9af981efd34cea08af26fe19bf194921dfae397c146d40b1c8b1eb9ec0
z3d8df78754b3f79f8f9e2400c1e7e603491fa3c7c1b7ab29f1884228c13388f8e34c18e6e00992
z951e4b8af6ce8c538b4973d967a23127835167ca8c4854c42131996c9281dc11fa6f6149cbcd9d
zeec5b9aa9d3177f3bc45b1482f24bb28a87126616a407dfde7ba76a4b9145ee8ced664385ae3ec
z6c432762f4528612dd91991b0b796127c00c2e58fa061e1b3c0d4b8c6a37a5e4c07210216f60be
z6e535e0dd4bee382c13f28b79607c076ddbc95a02496e0d68a8899fdd8ec7d193108ae6eee29a7
z52630c615f2b345381d304582ec295140cd2c07ecc9acf1e271599b9dcfac319ee951cbd15d311
zaadc5746eaa60471f08d8d08271bbdf2bee71f2ce10a5249182e1d1ccd70b99c8f7e8737aeb0c2
z4df4d72a077e06a9f50c5891eeffd79373a7b08642a82ccc6af237f8471560722f369a6c20d362
z0fb3b83ad7b5ecad2fa1d29e04cf80124e4df80da11df66f08d17b4b5969b0b6b031234fa41482
z88e9fabd64af1981f8607dcbba3f1d14a27cb7e882217ff19c81d4c619d4f1b5a8a37f61892cd7
zc340892a7a2af043550f3de2e4febb650e0a8a746abd8ba2aea1a3bb74ae0176d11dd329b8e73d
z216d83d515896978f38a6fec4503529da8295e1c5fbfe7633e6ae38b01b380f2c57b9e21923f61
z75f39a3c36733f7589cbf1078f8e7b6c76d828cd36245e547355eabebcbb68ab551f480ef842fe
z3d04e891df707f4b77c7ca729060475fb10005fb55c06425c0d1e860b93c73424e40cd3caabae3
zca18544802d0cd892775085af9927c8db452de0f1ca8dde01940ff4e350106d45f3c38fa31a6c9
zf7e3d84bdfa3e8eb8b33d6f36fd9cb2fabb78d8cbe48421da761065c5c5cd63c4f3f36cbd84477
zc98a77adda3779d94300f12fc51be8ded38117b4cde059a30b4b8ad40a271ab3d6a0bb7c1b581c
z1f295707646a54fe86f4604d4d4f6673b83e7113c88a70c54dadad513539c58e5fd7e046feeb95
z3b5d14e2a83c6015db31cd7579238ac99b22e97090c59d5b1aa787f5f858098d7e8a5744cee11a
zd06442a94e4906e74f7f31b7da2f1039811dc4ee3d207398f84895654f427a9303dd4acfacdfd4
z3d5c2807ee26b2f79fdfafdcff7334ca641253ca3986d204b953b017c88bb1f4bd2aae69985707
za138ebe36fb49dcebee5f3389d41e5a8e4e04fac787cdcd12547cb071de4f78dd714abf1c9c85d
z4a98165d2b538f19633009b99da7977b4c7d4b2956d7e02c05d86c27fc5d57d1c88da5c24f79b1
z125cdad9c442f1e10474ea50001b8275ca3c971fc00b93a26a65cd9ae93978be91ae72db443604
zacdb878f2bb56f3c16dc616bc1be0a2b047d723302c722e7533a6eb6c8c09f8a4af5b993a6b4cd
zab96c9c65d9b7e7d2be28647cafed862ce8cacf90b26224ffe985c7ebea81f26fd7f20a359cd28
zb687f5b3958450a7dd22d8d28ae34fc5123aefa0eb44e4989515bca862af5d81bc0cdbb53d41c1
z09d4f3e23c217d1535c999cac2e7201323bfebbc6e7fe81d1b49bd96581a5fa6b1bc577dd03c95
z3e9a730f3c07ed914f12273012790408
`end_protected_0in
`else
`ifdef MODEL_TECH
`include "qvl_req_ack_assertions.mti.svp"
`endif // MODEL_TECH
`endif // encrypted_0in
