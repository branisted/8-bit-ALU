`ifdef encrypted_0in
`protected_0in
ze74c34e226135848fe16db9ffd31815111b6d7fb642c521a3f628cf6da949865580b22efd062a7
ze90adae0e65e66a2c36a587d0a790699161455169ed55a01f2084f11770a774ec4c588039b380f
z6de9c5084882a40b79a175f5c2114b2b6d78b070cb806e1c0aa9258297f4687ab308bc470f0040
zb0b1de382961eeeaf2e279e1462520fc31c119af8f2b214846f56c2b3cd2eadbe4099496abff18
z15cec83ec4a77b868344aa20ba7360908f5c0de2a79abf8b3534b883bb12180f68b5d4beb444cf
z3fba8f13afb0abfe8fcc4294810f75afe452434d2d0f1166236c82f76edf1e12979f04bc35693e
z32ae028996dd85737a8f5adc1ebb94f39c940246e887647b64782cd7ab429b0544c173176cede7
z01dfb26b1f73408344a52b7e1f117f12bb9c8077b34876c2e6fdc085981637012dc9754765e1a9
zc512ce062e0b8fb16a214591f5c81e1353b900a611fe1f4886b57940b41b7f2ce99a7b84b04b90
z916f717e73bd10589c81e207ed77ec660a8cbed5b487fa50acde1b055c8870bd8676023f21ddcf
z9c98cc47cfa2d654ff1365d1f45035a045a66c5dfa8279050262ac56ccafe221d4824992a69d8a
z0056c786d54cd57e5ac49b6b8aa4fb7a6065bae21c146cc6f3a280ec9ff5fb2462d875d53133bf
zae8f4d22536259f63fbeae66512016868f4b63270445a643568f989ac09b3bc1139d0d92d9eb1a
z88c4a29c4e2d0f662661c665337037b0c0df7cd34064a8e765530589eddbb6721ce01b10a00050
z524d7a9f3dd3c68fb9ecd8e60e273896dcd7408b715b5feced8a835af3fe968b827ceab0ba9e7c
zae6522b7818761ee900f51dda9dee0552f02d56b9f29d80e35db30238a12101ae1d6271cd6dcae
z2751ab86bdba7e88a58177fe5fca2c4877e08191265b4595833b16cfb191f3b05ed40761baed6e
z309f1f341e8fd5c8d00520691ee5d3924ba313b1e0f7f07eff91d48ff90a9c5def2ef1db808a6d
zf4a33d4de3d33b376feaa5c24becc445df3ae0a2d7a34f7f66b66bfe11ef85ff2c9f989a97893d
z8565960be7f204a5bde683bd9395a8536ae0613fef32b582b0f337ed867d99d5eaeb374e9b0722
zeb2a823ccd1585aabb1dd45c25974b63245f2c8da474437f8c74f43776e65250a3724747814eb7
z6ab33b583c259b8a4718adbfef084d81b70977acc12d31cb664a36311506508196023dddad37a8
z5934b5fab7445af43f10b996fbb98de89c434d15e4d4f3dc62aa1499e2ad0a9496dc37188d342a
zc7aac8adc6145760019dcacb462eb887e47421c5df952fcd51e818fd28cbd80e834119570c8384
z63b69f81132fedaa102fdbc9657cf0da313709941e1331f986c7e9442f91ef082257a252558bcb
z22fb5ec3a7f4eb23c37b80710afa108bd887d457e0669e0e2075a8153f7c1580c0666f6373eb75
zaf7de8740dc5807ace95994d4eabbdd3a4d80b50380aee703381b7eafd3f3d666d529962ca4e53
z4c1755b522def4e32872c8e08034dca44a913accf9092b2e76bab508acc2271db65c92ea647410
zbc9ab431a65e6255c5615feb847b50beb058551a889153cfd61fe633a6174db8d806403c1158bc
z70739150cd0824f20a1ecbed4fa4df861948b5123fe542054dfb065650cc01735d503177145ff1
z75ba13645e855a31217f7c284d4d02904620172cf07a04a444625799e956fa0759ff1542ffc933
z9c5d81df0347b9c1b188f58fac67e8066dc03c6e10d6c0a1dfa5150f5a78f89fae813ab3234e5f
z0629850de329305753d3eff001c8b5da5a534e72d0608127ef279563878c2057542094a134a5cb
z06f5e7534e2efafdbe8b31e89ae2f4ad27f2c5ec891069fa9cb1676777444fbf7dd9db20971b11
zea8be9e22be0c75503af066ace45954c7691c41cd62089ea1705b69a43b5489074025ba2c6c5e3
zbaa2fe03ba1e2d27f026e33b6b5b4a82752fd96a21bac721ddfda1c27d65cacb0baf95a307e66c
zea65afaef88a0fdfd7b363d1930cdb75d487ae190731c0d6682d9915da23d9703deb006c984ca6
z607b57e367917f9bcc7a6e225b34b9939529accac43962beac6f68d121a3937a78d01151adc5a8
zbb29074fbb234bd4acb2f5bececcaf3ae93d75f101b64581f3798077afbb1d169b4aedc4ae3cdf
zdddc531efa39eeac1d23df6e4b0c52cae32ef5456125f28d63fa05b408afcd17b1e54c9583106e
z8ebec1aa3d12cf167a2a2f06a9e5e6e78ca2cc90d65ae11787bbbb12d22f9f78f5854110e12264
z133256a2ec497f4026d2137ac6c27d50ce0e56614d728e2f388accad8cd50f57d37d23ccf69432
z2f8b14815132701e8d956553b9d3375893fcc7c6b596888b3099428ab3fe2d30d8a64712ef4e40
zfaf3e5b130b9fdabc6948eaa3506f875a6cab837459a8a5ccf82b5d86205b3a536a09953e65fcd
zf17e2b384236874e27a3924e3515c9a4c8c3381bea0c25d0f41864b46496f2becaa270b8f4e4dc
zaf07f16ff4bce9aa977144829164bb02890aeb18b34c7f49c4883eafa76fb993f0352cc8a0a1b0
z8d218be7e07bdc503fe22087933a86c805a90cab9274879d1c379a667445878e4096960b58c34f
z103a3a663dc1254adc26dd75b752391f1b2d5f9b012fd85844de6074a14034b9cb2303576feb61
z77af0d3eef712156f054c6217a2960d476a15e9b38c61468109abf2694bdfef693ab084d4f85dc
zc4ac2373cfec8e0ed923087761febb6c1ca0b7062e392a0acee60051ee35e11eb00c60efb62702
z48e0b89082390295f82b5bdd3cad41f8a8b0feae4c314f2506c700663c9df80121241b16538835
zeb0ca452042fade28fe70d30faa6f2b7a0343167c8a0752bfa0aaefa145d79c0e1b19106e37ef8
z0dda6c4c3d25594fd1f2d060d88f584beb32d4358c832c32363d3997503ae6f77d9f04c048d501
zcf104dc31cf8f95baba9d5f8ec888ac2ebf6517d48f7a8cbb2ab0fce18633de2b42f042aa39bcd
zfa7ba042c955549b683112396cc242cbcf2549802ae706c53c7790a8361eaf90343489dd2c5316
zdff7ebb2c7e96442796c016d9a3cec52545fa8bef96a682d10ff5f692d794de7fa22d5966f4841
z6e6bfee4c8189ad6ebaef81480ff2c5412b02f4dfdb55829a2e9cbb7834d97845632a9604604c2
z39219b8c2f14ac31b5263f35a70b3d952987dda38c882d93bd98d95a10b0cb50e1d1750c770b02
z3ca53525d89ff89a930e20a37bad228c74fed2530a41ee2a612efb0cf3acbccb0066358f41dd28
z3e936d32181ba239ccf24a91902daff9ab48bca047af6823f581f9843d3030f84d1b0709651eea
z572fb1b061fed27e2c9061e36b144241b4112ef287e75efd5dd1e467059ba2e353fac6191ff26f
z14b018df03ee731bd54a302c26522ac68d313acce4093dba361a75c4b28d9a9f4429dfc0a07e7c
z2d6c7e6c3e709478f5c9db8461a788c0923d88661230559d560b4fe32c1d93cb4cec77dcdceff0
zc97bc3ce5201ca4e9815784dd41120f6e7edf6e3191a953ef06e680936716013cd7741de8a28d5
z9579b56eb4cddd83e0146c8d13707c42a600d0c2438ffd94a43fc4e847922f878ba5ae97de6901
z963ce8034d7b12602bc566684048b2c8d157bd4c1c01b4dfc69883323a2a6097e249bffdefee83
z532740d10eb540d00a4798d1b389d515c55244e7cbb27e31834a63f3b2887931b5b2d690238eaf
zab415b0221c3c18a0fe66ff3f79bd5aa1ff37136fc43d69b1b5f2892bbab29d9357429fcc12e07
z8895062cf00a34597f86b3c6b0eeec7a406a2565ba3f91eccad2f220f0a7b2171f86d565ae6062
zaefb9df59d2ce8b2b168a8fc5caa8069e4c7ee378139964dcd506407b063957d18ccbe9f244a79
z263ba824b440bb3c21eb3bcc3d0033cb2046e31fc578d40e459e223b0358c025544c3496c1eac8
z80bc87df0399c2c91a77360fe2cc97c73940bf94824a8f42066538ba38846fd32007a2cbf2a0bb
z15da83b75da511ad965fc4618f0bd191e034c81330fd46916cd9f401e9deb4ff500cd20673164f
z6c8b434c905a19da0d23caf89b45069fcb0a69636318ae164200b8b2a05c3760bc1af5a093ea04
z93883d306af3b34b8f0a5f927581ad39526b832f675704db08561ba98f3444f5cfd45ecdb6daff
z55030650f814f0aac452c61b8129dcd5472d4b9a4d0ca3bf5560cb6049b8c5d0374074e0dfe647
zffaa849ce25393eb8adc85eb83f591b36f3df4b9a6878e29f2af8460e7a89ed4f87053ef27bb28
zd3943e09cb66eb45d47aaab3ba7fd122203e59cf1bd15b291e0a902b46ae9638a71cdeb54c4c0d
zdd3aa58448b387704637451767a908bc146d8a82732f6e62368aa659afe66caba511cb82989cb8
z1bc689be9e00bb91168fecf79b4326a8a326d73574a08b0bb1d11ee79d61e25ae2a18159692134
za55cdb9bd4174793f0455610c70f68f257038146b4c2de33a892c0c094a0ddc050fe8797dba9ff
z94fb6f39d44e21d12a1ee9a7ebeafd68a2b2daf1e2a7bf303547255fae6e3eaa6159c2635f73e8
z3441a0b61a7fdd090c8d004120fc8a8f485067f575c634853ba200850eaa8f3e9a4b3b81db2329
zb598872a0909e5f4c0736d96abfceddd73c53ac1123315f3364fc0b15f36bb81b8e3ff9f6f433c
z101cd53faa6940c9fcaa5b54e29bdb3eedb867bf5ae68f9c9befd4d40f00a699421a6553501d29
za2157fa5d785ac78a4d5cccd110ca384fcb46ca3b731ddb31cca32554ccd23bffd436106866b80
z3f769e7ea72585adc268fb44b760bfd3e9c5a5e6a5f272c5755626504a3ff1316985347a33e3c3
z5a347871f9db984de1590c7f16192f0e18eb128cc5b13f2ff9b94723398f07f752f53fa76c1702
z3775e8065476b57d4393bfd7477dd0babc33cf29f1da627cc7df3ed33eaf4198657815a2f3a826
za68846484fcd9b85cb9f19298ec6bf2bb19e3cc143ba039892b84b99f5893121e8df0ed618f009
zaa35dad52f9b33dc123d617a980ed4d13c06f8d7c07d007b3a0a905b3a90a0387ce2138d4438a7
z3f3f00192ddba8f5f5e356c1399d840e3024e5c92d94126fed63796b0cdfb5d9702c7ab009c0f2
z8ba5d7d2033abc23db3a8416ffa1cf090b7a9e84b32cf2ef31ec4428030de4211aa8a98f27b91f
z767f2077442b7d5a35a06ad9bc8f307342abf4ba464f1b350db72b7278c6d374cfcc5b1e6dd14a
z521533a0cf1b52036eca9edd5ef63ba6f6a33414dad4a6bf61466d91bf1ed91cadc0cc25f5417b
ze468723f7c0765ca47374269621b13e2bcaad5aa300311f8f6ac46ab0f8a2537e887841e101087
za51c3378d4828ce834eea01e3fb2cc520a5d0dca963bab168c40f774cc39df735bd69eb33f4853
z53576c320bf6997918441efa4fa8d9b4e24db6c11886e6906a049eb750b354ce9c5e4845e9e363
z3a55a15dcd087cf530fc6ea745ce741ce76850ec0663ae5430cd91aafa401195a1f0779a5fe93e
z82abe883741651f0454e73dd5bcb0faa11464f12c4dd06d264dbbbdd53e2618c6af8c5f94e6cba
z7c0e08ea74feea4681c1ba78517ed45b3d2ebd32401ffd2c850c3769123322f65381fd354689e4
z530bf8c011ba7d3a55b62d09a8375ce45cf8b1cff14352ce116ceefb001e6c297321fe7834e59f
zf60ebb6afc063a61a50c409a97c1133b4b652fa560547008c6ef15c209bf2eb9a803d8e885fc42
za83eb4a57ddbd39473ba9580904cc01491470497e628fee1c3bd8616768849b3544afdcc2c5b6a
zde83b29619f323f18504f6230c0e1e8b1f4ded6b081856d8b2f51282afb1388d76b135d59aa17f
za9b666bfe4e4aafc840e9c8fd8b5a7a1a7b15c1904838da87d448576ae790a45ff62df9ffb4909
z867d626cf1010333d80b0e766b17af036b1580d663991900220b54cbfd3918bd09bc36d5adee25
z8460344a83f9b7c1d82d40f7aeefe14b7de15e612e150108ca796e92b47e0e3857bf9f00b48071
z502bdf12e09e68502849d3000845d5570a1421d062c9bbe9dbc588d129d78b4020da9fcc8a1add
zeb270a3b4ac08e11f36746888259f78bbf967eead751dfce4a46961053b713bccb3ca35e97323d
zb541d6a46b1803c62970ca296644d6e23151803ea2c48689ce7fd4ac091ff43061166720c356b3
z705c5b3f3595e21415de0e3bbfe0f577580fcc14f3596722450bca6820de07ca6ac81aaeabb8aa
z534d75e7884b27b925885cbafcc5fd5a4191de096abe9984dab6a22620319d50770f19768609c9
zaa69e797398e8543a8224512dbebccc7a9d45b688089a7648f590de6fe325e1349afed1a2b63d8
z36462504a9113adc7b42282c572accdf060d6f2b7c387e3aa261abdc3ac66a5a33af12052d221d
z2b9db6fec65b5f9f99150bcb144dc969fc32527efa46838f83f069c0c371a09f9cb3333e61f7af
zf37710efbdd9fcffd9369f574b796ac0f1142af13fcfe4eeeb441e7d99049b405c1158fdcf61de
z15b25fa098aa1e91041192ae265b414b39871d4fbddf416eb76e30496a050c9206864458acd6c5
z0850cecb7470eff6767d2946bcb2e979d2b2849abed969fd62af867641cd11d50e4c50f11d0509
z3bba7bc0ca5ecadb11a65c6bce7204c4811c7db2b337067fcecf2202874fd2403878056db7445d
z89c84dadacb2f65bcb3567b070398c613a80014b500faa2da676b4ef414de155e93bdd4250361b
z6ec2f204b6597ae8464e5fd437d0bdb84e1673c96fb3328652ad3a4ccf3db0a136d59131487cc8
z449e08efb7d68c108bdc6f84aedae0ccc348a57a8552d9e7424a76a3cfe9b0fae3c86f7bb0a8ac
z933e52cc52e750f52605152e03d54ea0d31c5c9a9e0922f0c1c3b0794670bf3ea942e1a9aec40a
z3305ce457c2d84496e1ac012f3b2a4829b56993a18fe87732c3ab4d661daeb1d993d0a35785569
z081a519200db71a88845c4f42e0883999b7257f39259fc441806d2ec92bf46ce49294135e068e6
z46b625adeac1320f6034f849827dc856ad58770bf831ab2dfe8c98f1796e67daa1713197be0e3a
zfa9580ecb78dbaebfea1069b018a95c9f04a0266ae6d8337817dc6d95d7405ab5a1e411d4c8476
z1a9a38e3b4fa0f81fa1aa6f725227d8fcdc75d338d59425cdc569275f692e4428f4915f80ed0f7
z96235bb362d801ecf450098f61af237a60631077877ea97f975fcad6f37f7a124540191e005706
z17ba88703a3e8c6136cff7ae0ccc19b9c68bc0cad7c419050455bb07e9fc329e87b540c5884dba
z749c663633de6b034c0ab7f0d6c74887aea7c7226d64908276574e664d0d2b4cab743af6b8259a
z61608fddb063aff7f28fbfe4c5ef1a21933d6a914eeaa62e330e8ad6118f37cbbd5b67d76fe241
zb7acbee943e5dac5554457d28b3a52b1d4ea0dfd22d85c6268c02f207b6b2c5327b746be4a8b48
za2007a58d37805f3233c218ef00de34ba4e623f630162a3e344cb7b4ac6325cf05b9afef12c8db
z0d1bc218b8f1257d9cf74410e5f31556c1156aefa805ecbe981fb4a7cd89f0081814d96bd31669
zb348f833708b87900848045f77e42eaed3c57aea1916626de373be1f73c925a4aa6b4d887f1286
z72543f019a58afb9ed9f6f7b79334c782e62c30c8e6e667f208f8aab6e72d5eb0fcb00f46d1561
z3c1081932f637187ccdd583aa316c99e16d3c1bf9f51ee6895dc765d9a33adf06c3b0ea6cd5734
z9d40e953084c82b0c98c86c98e41c578ce32f685fdebf00931c45a50b1cfa71eee3d390edf76e3
z6245d2bf45abb366715e84cc902d19123fa0d90fd24d0bc40069b12a3aff76a77715a1ae2c43c1
z69a8e16d4953f373f88c2e9970f07f495fd558744c8139aeedb33e5df63b0a33eafc949cbddb4c
z5a4ad1f7f1fbf0cd91cdf1e3d866a492b1075ff9377fbfd4df62a996c72850c3fc21d33c2f57a6
z581fbf2551f182895fdfafec41e661085456a79c9ce7d94f0f1593b69fa67902e34b77105cc280
zdcc9a5027013f9253ee8f103bfc94247af414bd85cde3c495fe18b6c0f7b6a4177a842e8d012d6
ze82bd7307898ca605a9920f85369bc0878009528c117c4ff07a3d1772707144e04f49a1423b69c
zf83faff9d97dab9106a579e2cdee626a36e118d843d1af04ee74ff9be82fdabf94348cd9bd515e
zb04be211743acb2c0fe2ec7cfdfb611e99f56e3394d70cb13411771e560184ae6472dd3934a981
zc2155a8f26ab45f7da9d439365c4bcf04766cc0d69a78a42ac0b1429e70eb9ed127745faf83290
zfdb5fdc038c444a8f6a5dd134ac45495a71718e3a10844a10bc68800c6c53c676eec4a47c97391
z75d0b82f9a2568336ba17d8dc72cdaea9c377d6839de4904439d8ef238e0cdbce5c36bba6529dc
z87323d95ede36e7374c859f556defb4e24d540f47c1273d0549c23672831af60481c069350a9d7
z007c2ad98f39212e174bd19bdf26f8e9049e37c2069c251c582f3fdefa1631069c35fd2759a9fc
z5d8b0f769a2cf7ffbf3f807bd460bfcf82de22c6f6916db69a112be2f1e1c8f958be499a5ec185
z43a2a240fd4e70ff695b4fb0ce4506ead984c6e3b559ae45d8c97a27ae8d324889825949ea094c
z9d477e31ec0f6f7e156ea655818ce1b4751ad8891bacc1511f4089616bf3eb64f686783a547fb2
zbbd5a69c5789ed51b5aec4ee822b1aea3908b8887e5c5ccdb233b95aab15534ff9b1100b6a5c10
zb1775f33fca9de54bd75162c179ef0b1761b4ef6c2caa1c3f2a83347f408a3929c19555da1aa4f
z15afbce01ca271533ad3c409b7b092cd4c4e91729ea8b066d21f7b8929292f3415310f18778238
z3d00e47b3526df23f6dc6a611d372ce77a5b4363c0078b3cb8a7d7e9e3bbe233d171aa13559613
zbacd6407eb8400cbab11826d2d679b5392a043715bf9787cf6284391f4941bd617a380b49b1a52
z3512753b1ffabb83cfe87cfa2ad49f13a8b2ecddc7f5fd0fb52be60097a5c6ec42d2b686448b51
z74660c52be91e511e73295a838bf387522e9420968fb2075388553e8f17ec9d0ed97802036d313
z8feb20863c0b4af3cc3b8ce2ba9fb0ed4edb6b15cdb2c2686dfdab31e858914fefa3af321a6905
z15ada83ce1411c597a0bccd834dc4e7439e1bffde34110c169cbbdc9f0de15c102c48d814c178d
z384943aaeb9334e499fc54e01fa8f63f10389a05aea5ba4eade3940a88730c4662b8374ef09bf7
zf3e2e628af8c0d95626d2702c0f5ce5b57da62392da9a1022f1351a92b1ba5eacdd8ddfbba6224
ze56b369544899fa6343916bc1aff532913adc52165b9693d3d25db903348e807ef38a015236840
z9c4996c61b6ef4393d482d73cb62a828c2084df1be397faf48d5abbed908763fbc98bddf29dfd4
ze685ae67aacf51a9713ec9732ff000579537880784cea44f0665e6cc632fc19bc7a60112e7a781
zc4f7ed906ad114386ce915cf7cd85e82b9b006ce01f6dcb4b6968fc3b51d7f716dd55e975fb346
zb38f508baa6e8708de35c4378d40c700d20b000c3f1d8bdfcbf1ce0ac26b3e07871afbab62857a
zf2175f8a1c3bf23b77dec75d84d5664aff01eca6c1f4ae0c10a8c50d618ec8f597d201dc4b969f
zc39a8fcb9f949bd0b01e391528e060899253805e16a5b401d968f8e9de2be18f99313862eb929f
zc07e8f95c9f61dade8dea710b3cedaca953e59c608bf04b903519c890e0d79618d9328ca7689b0
z93118cadc3f4b5af282a16678666131633cab69e066a14cffe7ee5a4918128978bcb31838b4747
z06aa40e451b32c612bbab167459838696b52849d8199a840cf9b8fa97ec2666d1e7532980f5a1e
z024e82ec57f3d98fbd464727a0c3398fb4996317ccc49439a0b30f0afcb7dda08a74c2cb0ecbbe
z243bb3f312c2069e0db6434eddfc7efa1b8fe89f7c29a40713dfb6aa125f1a8408d6717b1cbfb1
zdb0d253a410049876089992ce59cd405947ecaa3714b1a42d59f5cfac2f4d6cef789c12446570f
z07d77e72a45d8c19b106a155cbf8b3475fa7b2bb772c6abb25d92c708a2d8c54997add2e496bd7
z88452b958bcfc72c4db5c5a2f9385bc211a12083960ce8d7c2165b15d2311c68850c612677c079
zd9be5efb8f5e41191eb99aad3b07953b5f13e7ffabf40f980af68c5cd4e201c660eb873fb346f5
z320432b2f3cb351bc2ddb5c6d2b2332a03af52ad2f0818e3eb395078f9b3e6c12f2708ab0ac937
z035f56cb10a04c63ea042ea845f169f55c771f5bb12f37bf61e4d090e02c54e296bdf6f09570f4
zd141287ed6c451f2b920f25f2d3ed92dce883dee113e88be95b025fffe71919e093e6b305e2f37
zf312f8b3da4770ec9a907fe9917a4071cbdfe0922a2dafe3fa7afc0d6eb08229b10168fe3da898
z7d97807b9cf406cf2f1e72a282a22cf030a514c308f97315e68f9420a2390a53d84c04bdabdb02
z9cd785594eabd9e6c9a2fd50e5466cd5aab481ea2aa5b2d3b460a03ef1ed5ea848bf76124b51ac
z366b0b848740f9c8acb21674f84f6151506c69848db40f1304203e415dff097d9d481efe0b7d14
z22c65d81460784feb3cfd8b89ba770cb9ded96cd37a7f7179ff78b52d159df2ffbc3d478357c93
za30c300e94937c6ab4f75f4771f0a1da21a4423140aeadbd7b017121704806a3c6776f52acdb11
z97356f929f7d8012dcff8b10f030b3cf6776a14d487dc02b8b372c9a898d2ce8bf640731ef2197
z36b4697dfd320e669e23431ddfc1a7b352817d979802228439e9e4001870f6c448e148c7571706
z53175f6fb5da7dd717cf95107501a30a0bf040485e2c5ce2da31b6f15a0638da1256a80e1cf87f
z5a3f2cb153ec6a59f0fc52feedbd501a8be36c6e6007d4f2f0b89b9e4a267b66867205e8e2b39b
za384271c98ccc55f95492871209d5949147f1a99f21d89e587f468434f71f5aa6cc89b30251e31
z698bf850b7dfd6b13d5e99b59886ac07be1101aeaac73ab5d140362d1468fde19aff07c954807c
z865bfeadb37a1924b9db0883d2d5be4fc9619f0e1c7218f8d126399a9f23858972269c67c68484
z9665af890074108c99791e7d2ce8b6640587f5c0f4545562167a4a79719b5c658983198d03ff28
zf21fc5bf38f64515357db39ece0755f6c9bfffb9b7956c540418e4d1af8bf6358f5b88973661c3
z09c6ca7e5f33ec3ef7993f8e3ebc8ec488bc0b9ddda36e3ef555bb2d3b2804338f4d5c23a58e65
za718eb3c59473e38d222c875052fe62a0ed2181c200786bba3a66dab89e0f8eee23f1217a6e365
z735298d18960a27fe76013179bdce6d30abff8c949f88aa726192f04135ef3c22a772daacdab42
z6a708dab866addc46af6a406aeca645b1fdabb421bdb91503783e7d14339cba3b5289942fc22f4
zfdb0465f111fb7a06502ace5fa8628a8b1924743a7cd1e1caee9599bc92a086fff5a50e075fc61
zefd6ba1bafb9ace0ba4a8f3846c715d8682506757e21bd20564cbb0c2075e0503e2375473e4ad3
zf021f8f4fd121fbada4b76ecf65c96f08ea0f59f66751f5fbee12649d71ed87cc191e048a57363
zbfd3021deb59ba265ad70b85040c5262679773c1b59f5906328d8b97ed80f65d281fd18c4c5dac
za352f3c2dd88593837ba18f6d955e1fceb3558376bf03ee6383af5bad6333326c9b8416476f997
z1631b051ad0acb484da0d4928e77847b62ca7097857972a8bb131f050ff523efc1a831f0a9a6f0
zb29062b526371e715b0aefcc79ed3473372f37980127b2086cb545b279dedd4eeb5dee38b04c80
z9dfada112598d18398b184c4824848349f0433a10e7924e4527a16e9687ce737babefab908fa00
zb899cb293d2289b71394afec9e9baa834a238bd3cf1e561da972df821f9b14fdb8accaf6d49db3
zc287a796363143a7f0f8bd569a554b38b1edf64d1abfb9f79f32145dcd24474d80a95561751a4f
z28c59390c4023f8b0084fd63cba72ab5cb943e3ba705dab66c74f7d8c1b924327e5f82e9fce901
z5ae05d4d1f573703f551981619374fdef63ca64ccb7a44786ddaebc4465d5f062428c5b97c3772
zac231787d3d79bc3f48161a8281629dba510a6132ce50c625f8bcc90c921aa0e639608f14b835b
z31ece1bd43094881c70de92137c91f786d175228348e45fdba387c77ff779233099be12169ac1d
z7266ab196a038c4008e6fdcab30301cefc560d5f71946f7c924d436a22546f870c4ef046d22da6
zd0147133d85257761121247a8b660874435e1b30dfa2fec8dbcb1d574ba21c54bbc53f7ebc27d6
z385e68cdc4b7f8954ebb26ad97b42a1d2c9159bea2e6f77be9656c0e706ee9a21d6d92230d0d02
zc68d68e844f881d6ad7aca3dc4115f7b254930afc8482c3668ab77cdf6f095bdff1ba5d3bd9e8c
z981ea492c67fb73b79b8118447a150deafd716ac7ecd683a9c2f2846d62d3f93e27cf8aa9511bf
z8ff684d13bedd5052be0cd78240bd75ea5c713d6ca4a046f1b50d523ac2670ae63839e0cab5d36
z87ac7201c1411d0d343f0e44d5eca5919a1fea2ae45e8bbca4bfc86094f64ece3cb03d2ac7b925
z198a49a2521b45b9026d5395b533fda338703968d09f9d88a52d1a5ea3155c5a096f64c13676a1
z73fddffe564b9e686c65fd3ac44e192b958970dd2fbc124aebddc29624ae1e8865166c43443c84
z71d517df75dd7dffa327459f571807fb9f2ab603cf6b5445c1e45972f152781a63ebe209fc5726
z38bb98228ca57dc3ba8c35d4a3d48e409497a12168c6829a835759894b77985f9ec3e5b2462c71
zd9330dfa648fba4e5ca01af58bb0fa64fb2fdd56280e49c2bcfb1f1f856a48c4986935fa9941cb
z8263afa8a79bd37a2ac037b708d22696f4ade9064bb00bd4a7344cff40d2b1410df6bcd02657b2
zcfe40a126842636de547b3769c6516c0af45cf1d0743614eb157c5c4893017431666721d18a5aa
z0f0e040503074746fdb3eff04ad51b17d881bcd515c629873f665df428f028d14082db314a74bb
zc6ba132bd5a5d80a10fbf8dfe4ac3e43ed5a51ef74ea1bfc6f1dfcac310697ef96278f4f3e1e34
z2daab6b2e54e759cf09ae96ae06ac00679d166a63cc946f6bb659a7a7fcd9c91869b9cd128d223
zb042f5bba646a76924d12da5b9127d16b9bc31c42f4f477b98caf44186cd8a53db5e81ac60068c
z5236762a52882785cf1eb3e8743ba8a9101f486653482ec58d154a9c5897702a8c7b2dc7fada30
zfadb058b84a33191d003ed7af21e747508f13aa9c72617222a7d0031c67ebb30b3e9b6b65d80dc
z4c527b1fe68bebf75c4299514cc0b630d64472b4294eb6c7d252f4b6d38c96bd35c7d5306486e2
zb861cbeb0c882852ffcf573fed5b0742ffaf0c331dda29a0069482cc44b4edbe4c65244aaa9549
zd9fb6cc62443c977d80f67bc94e5dc780c642f74965bf6828791c201b59ac39cb807dc541684a7
zccd4e12e9c167c30854a7302b77df53a0ef42219d23b77d124011278ff0c61fb4e4aa7355510a1
ze38e326416395e90a7cae1cecbbead33b53a679960432e0c809e02c8d0ce7f6de1c5d10d288048
z3970ff47e9bb370a82127520c8f8ef49206653203d5c9f51dc85eabe5e06b5b6e56aa730c05cb9
z7a25a023fcb48fa4674ec8b70fe786ef34b9f41fa9e0afa4fd342fc669ae6e87df98939ecabd2d
zcd76260cb17038e33fa30f918b976611c129020f742aaf0da50662f3c2cfd4e82e87f75bee2bda
zd73f8aff69456774b219381a5575505ee933722ac7f455c4f90cfcb22942a59de705f7279b25f7
z641e54f69141e9c8e82f5cdce18a397df6c3608bb20823279492525fd100932dbafeb4b6fea47c
z86ec2e0a6c208fb9e9fc79401b1bcd69e72d54588b759f7c66a0600a4b0fae28a06109e16580f8
z43c63008ef252cafc25c0d403e5ac497db6cc67b07adaf9a454fcc6cdba4be0820abb5cf050c18
zed718fa6470dd31c27c91fcb934612f371325482381077e6c566dd9001214bae8820b6630aa53d
za35eac9249800204f4182130f4daec925f4b562ad50bf4b04e1d119b477488d2d66d2d2d7b05f3
z3ebc4533fdf82e58058b38afab3955cf38b18f43355865446d7b082f736997d2f4d123911b84b3
zc464eb0e2a18c247d85da3f8feb37cb03f8f61fd656fe16a439b0dedaadb4a0ddf293e258c9c02
zd764b2d499d031862248802979571a610456f9a72342ac594b78483d1a4635c0ac004026f875d4
z7b2c0e6b4f119c00f1bf6da4741f4b3b6653076b7d909a139685f39c88d038c13f63bb37797cc3
zc2e45090e8639e2933fbc3bb0caabfa7fe0c157449b26354e1dc19c8039f403f48882dfa37039f
z8ae0ff55a31ccd8af33e3235368f84dbf0ddc48f0a7faf2302b37981e2c61d746d14c630a81997
zac5e12388e5ed43ecc7ed3c97a8747e37cd7347533c4be20c14f97d23591de26e5748c3b9ff722
zb57797effe038ee849d82289943fb65ea0c8d51c772ca126161087106cb03536049e1610b21263
z9f2c739e08b57d14d659aabb5237aee850a22a8ce17b8da0a89e3a93a84752b3ccbc054ef7a501
z103478e584c592061b8ee1566d5fe2b8cf9f1197e11c8a3547c6267edb63e02338ea2044ada861
zdbf7d1cff2fdae606e5642a399f53c071049eefeb6f3eb771eb7d13a114e51ab53e410b193ba19
z27199e3abeaaabd6e3bd78d0f0da6bbdd10e74aaf579e431bfe36b5e8ae0f9b50cd0a2dd193580
z80ec28c1534201f0d50d05d70253d557a7578fc0ec2cd78a0c84d65542688292fcc9c866cfcb24
zc097059294ec03baa0201d3990835fa802915119235d6df8c8f652982f45a0de13df3fe04748a3
z6ae54978e926bc2b2a4fb4e78631f19420a9ed090164f1e90739e0f002525a9d582c2ed28877d2
z637fde29361f96519193efe58c87fc90fc999ca129400c719dcb3caf713fafc4ed381265ad78a6
zb28ba3ce1917d13dedef4e0ceb065086d21ad64efb79fe3d0415a52c421b76c79f7b08c4e4206b
zb30e9b82002a2e45566fed3673633cba776874597f145baa55bfbc936cd81e10a7da47e0e4544e
zeee7a16a6da0ecddb27863fa80e9c9636311ee25f836e5e7522b718eb2f055da93f006ca3bf81a
zf350fe1bf45095ad863b2eada91a1ee906ca799d083cd3024d75e87423625a6fd84a4c082d22dd
z74859f1778a863c2f87a2f66c2ba779bb5b32ffbe0a25cf74baf0c64f15f3bc43d0da557a685bb
z17a7ed59509b7f17d226c69ddf08b7b55a79ae835d2ab9d6d821525f37003b39567c6aa7d0b186
ze435eb148b67232ae0c7ee78b7c1bc258a2511b319e7d2708cfe35328ebcc6ba5a12f6b2126fdf
z56262c08859437e38257a6f54367721bf669eb30c187ba5035b66a3f199dea8ab754195b29141d
z93a47a799cfcb70a83f156c625
`end_protected_0in
`else
`ifdef MODEL_TECH
`include "qvl_maximum_assertions.mti.svp"
`endif // MODEL_TECH
`endif // encrypted_0in
