`ifdef encrypted_0in
`protected_0in
ze74c34e226135848fe16db9ffd31815111b6d7fb642c521a3f628cf6da949865580b22efd062a7
ze90adae0e65e66a2c36a587d0a790699161455169ed55a01f2084f11770a774ec4c588039b380f
z6de9c5084882a40b79a175f5c2114b2b6d78b070cb806e1c0aa9258297f4687ab308bc470f0040
zb0b1de382961eeeaf2e279e1462520fc31c119af8f2b214846f56c2b3cd2eadbe4099496abff18
z15cec83ec4a77b868344aa20ba7360908f5c0de2a79abf8b3534b883bb12180f68b5d4beb444cf
z3fba8f13afb0abfe8fcc4294810f75afe452434d2d0f1166236c82f76edf1e12979f04bc35693e
z32ae028996dd85737a8f5adc1ebb94f39c940246e887647b64782cd7ab429b0544c173176cede7
z01dfb26b1f73408344a52b7e1f117f12bb9c8077b34876c2e6fdc085981637012dc9754765e1a9
zc512ce062e0b8fb16a214591f5c81e1353b900a611fe1f4886b57940b41b7f2ce99a7b84b04b90
z916f717e73bd10589c81e207ed77ec660a8cbed5b487fa50acde1b055c8870bd8676023f21ddcf
z9c98cc47cfa2d654ff1365d1f45035a045a66c5dfa82790502623b57a3af03bf0f0c0d35b51558
zb8b5f2d29acf03737a9ca2a053b7a8f06800d50b465c41b30eb585f62f3d0c2c5a43bc02b04c6d
z3d2f83eb25581b21f29e4f4c1951d6ced3c36c01d835a6ae3bba5dd963cc9a33c3226dd92fa50f
z07d22d6e959f2201357aee021ebf53a8b04f72e9f38101154ecec297af896bca4aebdb013743a9
zc0c8a406e0cc8cb858b6767ad2b0b7a64588a2313895449186df7ebee41e5f2277d38d4fb8bc28
zbb309ba292c7fd75ad4e0da5b3ef58b8c985c2217702ae29bf5290efefd69a9dd7bccf2cf03ab3
zba6fecbc652156d6867a4846471f1e5c4bbd0f52b3712f04c5416288eccedeb1e03e56e10e9ebe
zf3f237dca256970a5a75198022cf667bf0140307189e17ee8c20d084f1690593b7350364c68c02
z4a2911ddb37559bdf72d29954fd02a3c167329a484ceca890e88aa12499acbe53841cac1747cea
z4a2f17b3e65de24f14d0bcca43a7f625137b98c7161ad62dfe9edf2743881c7f352ab0e414cbbc
za03fe50566281fba196ac6435f97bf7b161125bcb39672d15d11e9dd912844a73f03fbeb61e318
zc94e075f90808d9643bfa63733d29ad93a5e5cfdb29fb745fe67fdf0fe268e4bde6494be583979
ze24dc535d72408497fb44f430a70bae41df0836cc6377001efa59e966517b510eb909ebd240790
z6c0e6ec261895c00fc6e32aa344ba3ea1d8fd3d169b2727bdf02a7757196ba7f5de3624a2d12d5
z918c9e95c47f19281569fde70373e9a9823836c1a1c0f2ce928d35591fbfccd1623ff26f68a2c9
z1fad5e6d9d1d447abe9d33f01e86f31984a0448573db2e2ccbd784945e68039d2c97afd0eb98c7
zfe14696206d5d265674313c31f5de5fced3603c693a472a110812e1341df33b3fecc1c00a7b78f
z240574fd5dfda7a0096e0b672062f4130fa4ead4f50d9a3f69bcd1d8958aa4e85c88e60d578a06
zbfd745fc8fac5a8bb6db74d56ea056c66d89736988e65a1a2d9b8f46383870dd6de356955a4bb7
z9044d61df91db8853e7549f4facba39850c767e9cabaf83835b3e8b3bb96834a7c47386c48a659
z4a56761d56acc24d03622c8493f8c91229055176488eb3663d7884c4e121335102f41a2b274881
z159d110fe9d2186efca25249e29e4c83b0dcca7ed877485577749439065fff4d6327cf74f395ec
zb4561593ebd421a1de4de3d213ddebacede863fe0f59b02e01164c22046bbf5cc32a5218adef71
zb524366b390288c7b2af7dbf86bf2102037ec4543e1838f4939345375ec5c50905214a54f75a8d
za3dc26618be2421c52798f343c895cf61c1a60d5ea2994d2b895bb27638c1e3042890beb48a8aa
z03155436dc9620ff5337eafda9f07db89dbd74d26d0738a540454a5acf77a475733d4842c985be
z46f325afbbe018ec534267892fd301ea682e4fdb0e511a147f5e3bdd8e0343aaaf354f9a41eadc
zf5133e514c6374880ab02880071371d08cd8f4adb264518dfd18b42bcf539995c9d779ddecdd79
zb47a1b3535fd86aa078346f1c60f58d9ac73b754c6cdc72a01796e674c1eddb82b3292e7c0c305
zb33ae7b35ffaa3dbb74fefd89631f355ecabd7ad84f66a20ba2b6dd5063ba4da34e83efba2e2f3
z5190c28677f3260b130a6011654269f382f438942b57f7cf8c68039333041f228567396f668fc3
z23d92ac5e80c1d1695ac25736bc7d1afba1ad02213ff08441b56b051c906650410dd4f00064fc6
zecd1ebf5db5a413fe57cebbb6d05861026391e184bd47dd11fd8754425f6d0aa83284ca486e313
z59e86927cbeae52ea52ebd80c4f0129bef55849dde5524823577247c934643ddebda668fe8a55a
zfe009c30cab006b6c5fc7769f194bd9b240c73d7b765c76f66b37fe2a76d90653c408cf630f81f
zd9a04611a35d8c56957530a7c5575b9a861b240b4a0a1e5d71a17348ae90fa6a1cf7fc88840842
z21a0ff59a3a22e2cd60717d09efae615e8605395657072e5fa58e39a063c40635dfdfedd306bd2
z14b992e392c7bd4516b21adb14c66ac87059f6026b1f290efbe09a642ea1f65a194598bfd598ca
z4f9acd1495e4c46eddb3bd41fcd3b5dd40bf407541e6491923d5658df8d4133e534c1731167d6a
z16ff9eda809eaa1f746556fb01d661ad8a43b3b64bb4d8653942065598d1e9824c337de4ef70a2
zcb65646327032de9f6f28b934e0704311c516cbd1817625802df342bfc296525ad3238c01fb1bd
z8f9a6303ffef29707a09a6af4b8c86520a74d2f4551f5b130412114e65bbf02adcf6fb3415bafb
za535557332895483fabc2a2bc54c5ea7ac0654f2569745095679f79d4879b481ff49d83b478775
z2e8447e7f566c27670379b52e89778e29dc6c89f72cc0c843d5a9e39073c565a890053c5050890
zbf5534f5f7da8a18762d350f1193ca71fbf2f4c5e6ed1849206b4c514b0a9d76ab553adbccd308
zb59b2ad69f79b23609387b36f072f36d69728d3badbc31faba1573a316e9b437abd33f8991fda8
z4407939a08418d4ab1948d025a5f0fc06eb87fa941445d7ebbfab63299a9cf8bdef51587237ab4
z701c44e89462a0e2f3df721c8e6c79e7fed7f4dede40cf04927e742b64a890caf920f3afc6eca2
ze9d36a7ced472b024b0610a5f1064bfa88b276ccbe7f9ab96ed13fa5754616b99643cc58e66ee0
z3df66740200003ba76ab0e9babebb7bc236c4edf96c964a5235b3dcf7180e171e12a027954c4d2
zb6c82c62a21c710cdca76b7be585d135f7a57d36ddeb5a05b40b5a86d9964caeadeb3dd5b7ca9d
z77222d556260d77cac3d1e579bb29412d08bf70b1885a033b1b3265a0b364ec14d3fe8740a36ac
z803cf06d9fa22cf93f1e189b4192385456659099c024146cb5a102a237d56bea32a1879927514c
z16c2d8a0563d9d8610cb000250a4a82289b060f0920ef3fe4ad04ce96cacb3d5df23074457313a
z68f57d53efd312d61603fda50e00a1de18452bbe847416c6e3954ff3cb043d50c0856aa82a3986
z6c842d2663dab644d08b114091af56fdaaebc05700834fc665663b9adc975c2c4c3abc5b47d90f
z2450473e4025f5f884f945a6c521c3a362cb19d2e15431b206eb715765606bf627cafd2b134d17
zbb5eb396fab98a15f17ab06eb85fa1a835947546dcce23b3293ea9e4b133ea5b5a2c763392c4ba
zd1e802ac03e6af74752bc6e37c9801f76eac514da6ffa5da6348a7d8e1310b822a972a7a421c4f
z7d5a2d4c69fee2af46b5aec34882d8c8a34eece077e72b698397c9d0ef5a71273dc85ce4791564
z0d9d1209dd0dcc38f9aaa3262ee909f434d203f22c656ccf7f60596517b376717776a682d2bdf7
z1a3daee5099e47294e5460ce1edf6854360d53637b376bf4edd40423e8811cf54484b8c7ed6618
z3d0ae10e8c2df9329ce8030fb1048285d7a4ad89843c214450ec112dade6b90fd6deb14735c152
z0adb193515d4e27f1608900b9044bd77ac91f5b1f6c8e07e9e84a1acfcd6c188b966d93d3612c0
z4e9c966224a64655282f450e9033424049c72a9e4ce023113272a35d48546f1134c618933d5ae6
z676a9294d6187b2710f9614503fe6490f1c8e5914f1c635a121ad2203e5a20adab2881cfe9bbdd
z5bbe0c8f587bd4e98c682863f8b060ac58c170149cc366a6b145497987fc3c4477a93d30b438ac
z4d36916c4b5da29db47464e8566fb8542101996cda5e932c41897fb1c4d7c2d7e7de251125a5be
zdd20272ede0716cda5132ef747a016d05e8f71e0cffb2329997d56418cc4c7092ed468d5f142d9
z1fb487b65ed3608b1011bca270a5f6261c4842e806a4f56d4951fbad985aa58045de2df4524624
zd27179e965e4c670a90666376f014c2ad0f2398bc7aaebf668eecaa3785f5c159c2bff1f4a0df8
z6c90ee399e37a1b12630b32ffff83c26fe92681ea95cba2751571926c9a166ae658ddf631892f2
z28fc8ad757ea3ad37f29b0b80bc0e168ac9969ca02106d2be5e7a4d21d0e1f59d7ab7dc683d689
z41639fc5cb9e262007e9dc0d8587c9325ff36bdc18b282e2a08ea26edc21135fdcb9b6ba1abda7
z28e703481c97a797fa38736aa22aabf2b542d934e30f10d2c9624d49c6e29569150241e2f2fb12
z7bafe1852f29af54d7829a36503f683f7073d23c7628603ed2b0cdfa8337ce3ec4642078def130
z099735ef570c28d95f82329adaa396de4f9220b41d759c36ad11453029663d64a2a76f80b5ff0f
z0a837c23695c27ce61705da6b52cd6a4a14e589f88b165c45a4d5326a57b03f3fc35ad35c990be
z84027882464e4a9b636fe4a72b25b09423d080fcddf070bc5d21ffe70463388013a29f6453d533
z03fa8739ad45e4fdfdc55c7795f41f64863476315bb7481367e7c06516f5f6cb533decaf31d8d0
z1bf436b945e28576beb730c5df956a7faf78bb8be0426457b3654f07118ae89c1e1624f3e6110f
z618a6b419473ff65426a30537f53b5d687f6e3c7e9df2b8d708c4bdc79928dd5ded675d52d2bfb
zc4df12cd4b1c89f3b072a1a8955afb57102261b486a79501b03fcac358cf6bae942db3810e08eb
z4022eca85690dc10545fa900f6e030a95b686ff57f4d34fe1b5ba2fdb44019c9e49b143e7526e8
z8e86432a2656fc19eea23014a1966a64ab158b5340de702854da3b07c5d6ec5c980c4fe95f11dd
zfb30a6be606818f48c4158ac4d5fe5568879fb90ebdfacc6b1c1a01c34a3822746fc6b7c0f966f
z86938fa76334f6cf372cec5e3e721ca7833ae3772defaacd4389110bea21e076d63f3fe04814a8
z7c21126a330d24654912fa94d433d6a890f6378ae997c9e83749ade281ae5014687c28955afefb
za2b637dc25e23b13d36fd76b1e543663a7434e54f772f27feabdc0ec65f33af905f0f028576c22
z6dea7dbca2eb9717c647e1cd758b5a35098adc52b93384abc5cc13a32525552acf7c5a8445f1eb
z3e7b7428e985afd503a37fb11787ae32fd64275f2f20050a9f29d8b32405c4c44439658b595075
z45a40e8ff94da43b1bddb7c2ce0badbc79a3f5fdfa7fb7cba1ac2126fa435647f0f240ae975b43
z2462fca15ed4f904a27d9f1609efb0c5ccf672664d515b513ac71cdc67a35a0bf1617c552116c1
zcef049936eaa4064fd545ae413a769264fe9c011d09c6c024fc651bce47ba2d5a76dca9eef318c
z8310ffce923df5237c6aebd957bc14a9499f21ffbdc9f94c4aa020041aff62abdd9a3ba27220c7
z5be59f641064914acc5ab8d5cbea1cf53a70c746759cfebfc2e59b68b6ff2b5ac6cf78abd3da32
za8ab884dd23b448f60768349f3d83efb5409cc06dbafead10ed05c22a68c9b856f3d2722dab020
z9e7fdbc32404e793a4002fbb396d7953c8163b14414aa7386938022b9a53d43f35b8a365dbb8a6
zf656677b62ff88442a53828cf62414e5487b0a0e52bd40c10b67262c9054436d38e1c2016a4123
z5715a21ddd9818b61b33257298e8ed08193bb3e7e00c6dec394ad726b7a437c692f34d42a2dd98
zf0e6401ef5ae664d45ab0346c1191712ebd697381157deba9966ffa6117ec8b24c781cffecb814
z6213260a173c40012336756c1d7dbe683a5d30fa3c4be0e3f694c72219e41baa55a5ccf6ddaec1
za8a586fcd52c8a2d9422cbe84261fe7a8265fde1725a4dc832f78b684149005f510b36588c19ae
z2e8c262ea13b342d634ceb1780b33060e3bdb4056cb2d1e1872e7101dc400d6ce2c751600730ba
z3bcf8722f59040e2eaf9036a821651e6cf65bb8f346afd05bc7b816e2dbe929e0e1b252659e36d
ze6051664b63bc50bae07e34ae798f5d779ce870e65b93f4f69c5a498abf539b8d9497f0ee2af9e
z79244e4e154726ca22cdc651c293b02a617fac720032c0a8fada93b00e5cd907315cbd25cd3d64
zb8fef62ff276de0eed65be0614e0b0954a2e93cc9d6f6c722dce4203c9b5f7746410bba08327cd
z80aa7f75626f603d04b346173521b87284415992d7ebb08dac04d1d0ddb1b747a0c9abfffd367d
z02db4c59ad1be2244877accf806f87d582727f5bd5fcb1dd529c7e9455cfff7137194e59ffd4ac
zefc912c85e4bc73595f4eb180c67b939e1a31902aa6c89e5a7fc78ccfdcf1abf23674e05ef8378
z4bea110cd5aaa51648d1798d2a0977b40d2050dc3dbb0272f150bcf74347a1fd00102cf1858000
zf22da7558650c0bb8f29231e4b6b99fb158cb87ef9964435e7bec1436696cb5a3d7597d7523cb2
z18c46f6db29ef2a885ce3a2e6ed8547c9d1b86e27dc64eaa81cdf2f3e7556d16fa1525588ddd50
zea8692c7af2784aba786b4e0f45ea555b3cdfea7608f3f413006ff0327c1d59ec0c14910e60207
z1d4028afe1111787a028c59b775413eaf5977c5974f898b404861c7091bf6bbf293ed5c969ef42
zecd5e398a9d2a741d2c9b8acc38e2b24190128f97dfb7d09de866dac9fc1809daedae764ddfb16
z41614a4ad05cab218587bd2b23b509919bff9c4e0ce20aa91806d784a7059a417f51848a30758d
z2a1ea993fbfff1709e69f7ceb99a7fbcc6b7c18694eaf905470d48baf454b73589fecc91e518ec
z06443e197259e153eec976473284b5fa675adf2249f02ad38c18eba15d98a3a423a8b3c813261d
zc91107c6b895e8da74f472a84ba5b388a73b6e8cd4a69b5845aa319c4209eec5bbe0ab486af6a1
z7fa6bfe23a3a0a6db5d7a17d356844f40aadb4d44093a58857a796a29cee6780bf7d6a2aca9009
z10fe50e7fb6035dac706d2f7447079a2b358e319ee5c1b7d9a89761034e3ae4d1f3950e4a9321c
z70bc70a68e5ef1ce9936ea8400711a83db13ff1e9f2641b013545cd76a511011f68c6da714fb3c
zfe05f853fe831259d17334fa5969eea5c585580f24a9396af9bf618312a7899051bac4455438d4
zef87a7d07dc154520044d6a6f96acc7465ee432f525c507a2e0a84ce8c9523946f3b9ea885b9fb
z04cf0179701e1a050b389e814e96f71d54fa2f1895892fae254d276071e7525226899a14d5418f
z0e5bc98d7fa47142e6de24c31c6e1410f76214430f599801af55e269e5e12e88a234ab5a418d6c
zb5459f2fce263022beaa1a809e020065ead5e108e635f3efed9a189f57723bdc59537a481e0f35
z1522b5d4045ec5c03485de4037171c85d9fe1043c41f025cb5f1f6f9c44af0679934a93d295c95
z853d62152a35dc1075f5b07c0c6822856df7535d6cb9b82f073a12825cc3d04a83f26f68107cc8
z1da8563844711f1f15e862d6d0664bbf940d3a9488ad3f03ecc594e2f2254bd45ad4fa25d316b4
z689b39d5e820bbb0eeacb1bb0cd405637aa110566eed391e96c7514895d3d5c741499c8226d712
ze7397f4d84677ee45761789873903761c50d8ea22e440deb9a0cc2736a8b81a43308075cca6089
z48d022c98d24ee08e32747189db92f2747775e0a6f30a7a7b3902b28e2cee5036fb5c89e979427
zfe4ea2ebb6bf84f4683455bc4041c27264ff47981ac0832007fcce4ebd72adfad36e61fb15de75
z96d528c358cd9806aec92429f79c0b90f87da59bfbef477eb4f5a01e5bfb9c74c675ba6251e436
z484625d21e39145332e66736710da37bf67b1a0b79183125d60ef6d1dd7f95e544565a64609f00
zf7738eb69ae7a61816cc42d8b9d230c186f1da754c8a487b7ef4367f8157fb38d453891a72bb0b
zf6efc91bb19631c7def2365a7e14e5515d6993d61700ca9a84457efe390344877a227881562002
z36bc972583eba21f435471849c46ee1bf205073c36b0060d048daa125dc47e4c4c1016c4eca1ad
z0494ccb55b0a9a5530d74e715a2079c9b1e7fe560806ea3ba8160a3fdbeb8ddfdaceda06ffdb86
zc2a32b0849f3356af9fccc644697e428e544eb872a42fe6938f9a0c2ff2bedcce28a40ef8f01fd
zf8f060287644b7c1568f5188e0761d8dc85129e2c0fa82ddea3d3ccf31b54feb3a1125b4372d04
z67267a36b5d2c4828e1b44ce2bfb70b03eab2d3304e8262cae07bbd3957194a3082d2e493618b6
z46f683b4ad23cc6c50cc561eabbe8a2f83630a9b3672177fadedea9567aae860ac0913274e4340
z2bcf3e677f3b189a27d680f087a45aa30aea520f7981567fcb4ea912547d476797d6f962c1d8ae
z3d827928c4f11edd3e1d9465fa49341e21168e26ef095a784661b4ed9d3705e60778135775b080
z0f5d3d55f2fe7695d07c8709af33cc0c323919b02e539551e6ecf0d5a958b46fe3cbbf896e7bdb
z2d15cb62f7da40c167e97ac48e1d4903cf52a8db9109d3b2a38bb6370f01d5ded5c470e2522cfa
z2ab5f54df1f612fc9a5326080cecb911039a1254d28208aedbf701b65b32bddc72a1956d9568b8
z685b0d9a95481b395b9ff2647dfb966021c0e4c0045dcac2f5444e0895af523adc272566c3989f
z25816ddabe6591181f12f87ef90061ee5546f18ded13d593e908909238a99d446e47c00089b0cd
z621034836fd35b50748b03021d47421346375d672187c3b4d39ceae9fafdcda59065cf5e56c27d
z5dfe88d5b74369b50868f9c3f7a980bfb07ce434df5efe60161427ac6d76230ef3a1b91cf48081
z1f514519ae5d2b890b81295602742d0e8c71ee2537b577f381d6f47a3e9585464ee7abfe1461dd
z05042478d33999e7f5a707b4fd2806d04914c5a1bcbb5d4ba636bf3d582c6b0b60513736e8e25f
z5e328777da695da1e79dced934fc098bd9905a710135d501786a2faa985ce55ae2acf822f4d2ca
zcde98ab8948956b2a0c229c735ed385336e46ca8936bd6a654b22ff92a5b95daf59b92d11228f9
za4f2d346002f7afa4b7f9b24aa9e6f21299532ec7bb5a3757e4addc95965d7f0b698fe77a3a011
z6028071b9ffc47a9957fedf89dc73d52db59b006a63b97784ada72c4f3cf3c0a2cbb07f35f5749
z5536aeeb582061c2099f5c2009490c9e28cb59e63b69f3bd4a6a2795f3f10e51d3749de026815e
zd10e0642d23cac77602eef0dd2c25a17dd3ae9d6280fe4ff04cd2a4a5cdf99116e968e2a4f0bb2
z8c7292fcd277b281984b298ba713ca1e72e0ed70cec5d499ad3d157c924abebf27b40280546203
zd8864dc378f3d425835a8c624cf0a0eadfcfbda96f1bfc086b023ac54b4d044a514c624e0cf27b
z99bc0a78f18a5e43b7762d5e97ea1a620e28de09908f1f3b3e5a86f2cd1b86c2870d4c55fdc12e
zd3ea8c796798d02da35df8d0e13151ad36beebe9757f6891b8dae2662115dc1d39d85956486eeb
z35fee44bbc1e354526ceaef1cd81affae557e9a8187641048cd390e57180152faea87534112f2c
z44724a6c717299a5478721c19d888e9976faef7be6043fbae7ee4ce6220e54920102bd723fc2af
z695283a5441db428de552267a63756c18a6180273a16afdece4f09468b98649acc37e77d27a924
z907cf0e863678a49ddb111c80b03a3f891fbdc290d92d16425e79905d5e48570d4b1c2ce35cf0d
z79c22ee97d738d44ff89d725a22391777c12ca92c5f6c1b9edb282c17ae1a5ebf0dcd094aabbe6
zdb46dd857280b6105c42a8b1ddd24f28f33762fc9553e3b794bda9b7e407e4f2534865d2c37bcc
z15b22a75b6d37f5ed86fff346292862803a87e1f2188bc2620bbe1afccaae329cf96a28bb1ecd1
zb51e09bfe68599c6ebcc6caac1cc6dc56378f0fbb95fb5ae817276368cd172bb06899af744561d
z805d2d7173cc8b0dab6cbc6dcd793016c2b1165ead8c6fca032e9dd6c4aae255bb6595f62d42cb
z3c6d4bf965634e405de9bdb1fa656adbcf5cd3a8f1a99422b5be3317693ce8a915f2b77758c2fe
z05410e6673da467a1c56574484b6237e099158c39ac18f228d5f99281e31ac8cc6cbef54b664c8
zb0c16ec4915f8bead8fe512aa331055645be1010ae5e848fd636093cf45b9c75883459a3ebac6f
z109e328d7883925b28cfdb59da1a4a40163abfdfc484ceebc9b438dc9d197ed00f3f1f27c0aa2b
zc7b1af1ea2eabf29b01f91b66337274bff310a3390c93521f8d578009e1ad5350999e3fceb49d8
zd2150eaf1fe2f04f62168e19bb5283682abbcd23644a9ad128aa35b24e2fbbc86844e1e56136b2
z03965a4aae0c9704b546c917892abf1928dc0664e9ccd13c455b267ca0a7e9a300535a41667e98
z03b22631c7ff19631304e12f001073ad30ef9a9f84a0b1cb2503dc94ee936e4b5d4612bf24f47c
z4f94f3148a71d5105571bb4074a5bd8a82c8dbcdfb00e2966209fb958077b9683a17b82ddf3437
z54e102a52757ee661fca2533e208226cbb9a3548561b284d0ee27a5e3b65d9312e7025ae3da5ac
z1a3782dfe372810fc65d4233aa22d60f844b8a07b14c5558450b61543280b3da54cd147e820a6b
z3f4a2804ec7f78e474180eea894abbbb802f6880ce41bf36fb3490edc7ff6035cb62b61c6f34d7
zb1da2bd63008856495753ec2ce173e5a5cf7f20ff5d39b7a1e01b513266a9f4e43ec5031483e53
z6c043aaea1a223e8120b91d08f302f8af2e38b6bd181c1c9f210123f87cedb9207cc7c5ee00798
z853a60c6f9681b258f4549fcd3044763d04d21ddcfd76981dee79bbde33acbd283dfa51f2c34a3
z6a0e8491e73c806b710f3c1708b4b3373be4d9920fffe2bf720af8c89414502c225262056f127b
z706bdc4c99a51a2e26ce2e1f34c1acac2638bb2f55500acace759079567c46f8bbba98f2607d32
z5299bc928540c02f39d45ceac21633c842c7e76879bf8b92229e5079429359e203b2365d8ca3ff
za6d0d6675108599b865e60b43318ef3d5ee15c6633a8fd18a92fb4d7dae961e67429c533460111
z891f4f99fbeb6fbf5e24b00c3f64213e9e0e2fa459173b8e3a1a267ca8bfe1a15efb2e82183ade
z8643d528ad9fdcedb9d0f800cf0af8f6c1615e6a0c0bb98c16649d080f8da082d9bd086d2514c4
zb94c00e1b36a678cf9b0016b5750700937defa786737e1673db1d93fcaba9a09ac783ca6ddab8b
z6158a6c7167df0bcd8ee7849e9bcdf67a6f6323ddeaaba560dd97d293137fb8c033d7482d43f20
zf1bdb257830d7a537d70ff4177657e2c323a202b96535bac9cc6235332f9bce48c2fc1b2d551db
zd606ca4175a3796a513c7eede6fc1cc9e6bdf9ad57ca75f85fa7e0d4589bd5618c80715ac08d83
zc87687b58d1dc13e8e508d193fae81eedfa7742e1a1513454db165fdf51f5184fd86ee820bf013
z918f5589d2013cae009cd58c0c46ae9dafb479cce3bbbd0fcda0d632fe2e4ce3573659fe3c1959
za8c8c45f90319cd74f23248444ead6954938645ff987feeddc17e13d45916ddae14b7afe2e1de7
zdee47ea134a8f6842caf5e259b7afa17ab4c9ee2c636eae47e57ce4d5f625a23477895439d3f0d
zca5c1afb20e3653e3c100af1399f4d839690929e8614e1f0c804c94dc09bea353c8734648b12ed
zc8c329a0672500b6765f887a70cb56aee0d8f67f5009ff10426cd3190e65bba84a507c5633c9ea
zae5d1e843cbbf289cd54e61984538d4757596e7c272f53fece758d79ff7f2e0ec06e56200c1bde
z87a391775ce2eedbb258f64ba830dad7cd4283215b0a3dc77ac0663bed484cb0d7d3557bc25bd0
ze9f1783525f08e1f5af162d306a37aa14ad8ccb20efd4c5a8717224d644ea83bf351749eefe305
z9b9bb9e36502eca6fd66bc4188c67c0cbac1e92b26d3e620e6cd236eefa368577c8c8f132cbee7
zec940d011317a07dfca561c68ab978f5d6ae8583dbab6ee6e55d5b304f9705e22ea9ca78492c11
z197445a709081e5a179bbfba8f8ecc564bb154c9355956e0db4716e29324b7d3d62cbc679fdfb5
z3540552943fc72e8e6bfe4111d0507a71ff4075e90a274aa9b23d94ea72cc40ca160c3bd5c21ef
za2022bc3cb3fccc5cc2ac6813c7dfbad2786fd23a6e783f13e50aca4b669429752cacd95fe4331
zdb1104548ca679ece645dc3fc06f669f9366d09af377c47a42beafd5ef3b0ef9a1dfb05beacec3
z7e3c45249e27821f43292607eb74a778f2298e946326004315f7239b23aac92f30d7934afa5a0e
z98e3777ec096fb5831988578ce03325c9be4aeb7632e2ab8ca8ddf54fd8e0b6bbafd27e2542c4b
z3427a21e48eed5be69dc6d2ca74128f3f5ff7e9e60a911926ab3e6b3036208e80f7711f4e5f63b
z647fb5858b97dc4c7264b7a4bd136362277b56da264bb5091f4038cab4b0d663d9a28c86b81aff
zd8b88454bf498c13a64b44cbd8282330e9cffab52df993cc117925f2b6155ab201577882e2540c
z58512c17bcb19e93443bb39cefded0de120821f0b560036a936218fef105c4c0aed509380e3d4b
z3edd85a323b9ab1bf420e9fc87de37468d0d9d56088e04a0bf14e4e2e2d2acbff570f7cdacc7e8
z3c732551a49b37a39621eb154350ced42425cb7054c4f87b440e4c018a2b7e81362ad396e7dde9
z71df3822e3c4073fe86bee733951783df49dd6de7801bfef116e7a08e6bc64e553f79e259b27ea
z29519d6fa348cd88dcf1ebf2fd6f0502f2dd83ce80738f1620ec7ee60bf091ff5afd3a4df6ff81
zba15272b9d2722e79758ff0ced654f61b1d65e1162e0101a6e2f6f625acf5a0067e9b3a37decd4
z67d2668453200c077a8e8f9ae3c1449b09a464f0b7ddbf412261b2da3bff6065af1828b2e4a528
z575550cb37e81a39dea8cc76f3c0163eee6615d5d64b47065717895e2180f8a8e66cbcb28b0c8b
zc8c002d503b3e3eca18c8c6ac160d9c550cf02edb17736a9635e701ea92de021820083355a3d62
z0eae313437101ebd1d61d3b59fcc88bfcfac7c6d32156309d4e5c5745fb088e8a1efcc907f73a7
z86b6651a4ee8796bebaa1504dbef4818cd91f5639120be3115f26533aaf0a95457204f0e364070
z59f4592fcb35636ecee8f5a55a3cbc2d8e1d280a92bba0fcaa125bf9f14d91bf31ad59c2eb4628
ze60b39d0e0fafe2cd1ca22865bced204522b9fbc4011a09e848bbdb04bb69d9868988793dbce8b
zdf0c0d6284aa275af0dcf5e6dc1e2a26cd831d0a5e6a7227f0a7cf6477878a5c8ca32e560f7112
ze63d29dbd704448cc9bfbb2a529c5d54512db7112913a759a82e9a699dcfe4508c5ca0f593c241
z53e47e9606028304620a5cfa8fbd5f96897b6dbbea83872e007b5155822ee2efee1588bb7728f4
z80d364bd187c7c649d6495adcf2ecf07366fbad284aabe707947ac2cf8aa01233f65717dab8b67
z21bb2f6769d1f9fcb62fad94c0b452a87c2e6646d2fc84b0d6f1f5ed1ce4d902486c4f8f949a8e
ze009bcf02ea5218ce5ebd4275ac4314935e9fa63f15c8fa0ff0a5fea02d26c5608f2b2fde29dea
zc293f67c5399e5d12604e3fa6767d57271768413c90e0d22bf813a9f6bc83ab8a95e972fcb51e2
z5c219b0fef7ca0f470061d9a22a1f7889d41f11f27937d33e125c4f45d0ea2289b9a019e0b20c1
z7f2af5351092aed418772e56038384c7cf85c8206478409695052c087a0b43872d6ef845229cbf
zf862deca9be6fa995d538fe5c1ae0941a02fc0be8ff3bc62d27382ce9b9381a9fe04cdb7248ad4
z8e8630c33049834be126f80d4329a0d8cceebb8815c473eb908fd744b736b4439bbafb61d04354
z8f5f3f56e4a2f5106f383d92d457726d53014eb5974786ca587d860afb748169418aac8ebb73df
za82964c676f7915fe076425c401c13b457d67063c79034d355814576e917bb43c5a1c0b3dbe646
zc4ebd863c673b0f847a28bd97fd8838de3bc26b4fb2e5a86e236dd56ab945b61b3c819d02492c7
z6d605c6b86082837e042e17d9f4dc3752ba2256ac89dc9396fa708c28c75708161f4ac7bca594f
z7fdc7e736532dc8a9eed68e3874a9375f5ee64bf8c93bb79b70291de00cd5197d2397b7e38bca6
z83be769aec8926d207e961e78be938dcd3a24082034dd2731da90878fb9a1e455b1796738e2ef2
z89812e464a560d47810fd10755d1687495fbd5d8f7df336fc6919ed0d10d435889133444cc205b
z83dcfc00031b4b95405291b71980bfc780be9fa10cb86b18936b4f68604c3a6b065dbe55580c00
zb4422859b4800bfd9457dfb8fe43eb2bd3eee125284a2e67fc1b78e7fca04a601799ab6fb5dc1f
z4f81e0879327a49075b3f5c6d2e264c28090d9e162cdd8a45942e98e9fcb0e60ea6080506c8b0b
z79418d3662ab31e6c7863ed8f61fe6b3c030c738b6c6a75771e2013cd7acc113e7a1258153fb92
z485f030bd0f55f2541626585d44d13e1d095c49cc5a1b2348f4e5b37540f582a8c7216afe3aa73
zdd32e7056cb58514c3412b826ea90b90d1068f2d91a8389bdb5189678f308a78648a4d0476e3d7
z04e15da6fde544625942f6d925cdbf385d9137b571c38713f530f687a3966f131385bda01fe7df
za0b42bfcb0408228d42286bf668888e106adc1b6528d4fa1e025664e3ce3e057c34b936e12e18c
z41035f6b51a5801efae797a436ff12f624bf29795bb7b819f25b9553070cadcc86f932d91fc46a
z54de55e4ba83f77c41eae9ec695544ac76d4ef85308e56642b5b13283e570335f6f1be44fb3297
zff735c725dfbd982afb9b328e1a375f2567412b9a643103833d45ad21d9ea66b692e23492417ad
zdb9bb42799d123eab838a20ad12793d34857e6933f8df10c7a48bfecbc2b1266be290d73feb7ec
z5a76c9407204290c61f8d7eb466e49cb37e42b52b7b911adb16772ae31e07291a58f7b256ceb63
z49e3f1122ceeeae530bc3c9fdbd626b6558cc1080b9307ba9055f8996447674cc24e0d1a782184
zffd2ee3723f36694f7cada2c2d805a372a75ed8aa9335dcccf111baa396edc1ec6d6138ddd8804
z5ceaad1623f598ede5cbe66f39220b54d072fa8e7f720532012417fe5ace7803b9264f4b5f390b
zcd5dff13f0a6f8139b9d264199c71149febad6fef26660f4e7de05f0b8b2b0f6b647181bfccd64
z651761549d55a7641d37815eddf2c92827f57d1a855380a7149454a8ee3e75ff8a1c0fe378901c
ze3ac96f98ecdf9d87d4b9401f91d7f91150bb3bdc6d3a07f6346a3bf4ed2ce748f3211fe00f1f3
z79ae166ef81be19330c470f20f3d13a02d9296915613f87c597ee120b6f841080f9a5c49759d30
z53e8addf10fb4bf659d0632de7e2a0d7c7b5cabb701f204122a1126fed4a32ff3365486051a126
z1923f681e491cf0f1154204c0a983f4f0441b6ad6905933dd85f95373a0ea9b41eab29339d4711
z0fada5bd300e7bf2f32957aea65a4474b5f01512423b676488ae95f15a1a3dd397ea463bee4628
zca7f09c40e45f08e640b25efe3f25b4e9cf7952f471d8690707ea2d4b5c902cebf99a7f64bc2a8
z82a97c322c2a1202c59c768ed78329ab2bcc9dcdfb095a1b9bb4248ac1810150e9a96de34f7022
z2420b969b7ba7d3280a44f3cf62d2ed16f36245427af04aa0813be24ad0f1f4c58de75b952767c
zedc49d321026f116e296faf85079379f916233f7a4c88e31a21808026a04f35cb80c89776edfed
z4706189ccd91346eb2f7bdb4cab1c87e426dac3d6726aae4435617dc1f9a905b28d62746b18982
z212bfe79bf004382ff265a352d63913e3b3cf7998befd00204d44155c7d34fd5c6e65cb816ff18
zc51b55800108380d18b2aba26c5a6edf63fd3995991255d838077f17aa904f00cba62f26718e36
zfe84613d99ebd42b1593bbacb234aacbdcf3bfe540513516a22d1194669a68546c3b50685cdf39
z6e5a7628ccc753b21b06a5337c9b38122e091c69896ffb4da0ca234c348d2d64a2749f4169cff0
ze4a31cc886c957c94ad99011152ad3a4b885a3903bfa2cd9df17d379d6e245df3a45992fe1b688
z1956e41021e204d75e77a2cbd14deb8c755719093571970c1fadf9b39a87ba7c044167e011daa5
z1330b56d19f1b74950074b87f430d6cb8d1fe4174f0ea6fd20869f10d8b6c700a143176eeb9381
z8e30d2e37c7080b2b1f213f5a1a2c92beb1f9a3d84916778c96e8c06bd8c463ca4ef72bb985db5
z20f1c9cf7ad1c088555de3bebe4b7f0f182db2d5c16510ef932b039d400827e151734870c133df
z5f579170fb39363f6ab4129b8be568105fce095f817b4a5440865387cf37abb8d10ce20c82a549
z46c7e82a76598781c31b2dd3b18b176a11e77ea43a65250a33698b7582964a6d4a1b4f2a6575ce
z5fe6956c0426a05b77a6eae1ae70ce176ccb027718d40c457523e7a5c8511652c9b160099561c4
zc3fb458354371c0706eb0142d3e37844f2350d36cc3c2c5a0c139fd38d629ab5b11b511435b9ba
z22bcc20c6125232f14b7a9aeca3382131fdeaf3f19b45e0c1df280d9c454d39a1224af357d3375
zac7f2046c0538e238d6442cc67883d932053b2307e481cd8d1745aa6490254e4dedf56c0c6587b
z6ff8a39174c3dfd66bc4ba021c0a855b6894c759d3bef9942b70894f5c083f61280acbc43df2c0
zffc78f6569562422986478a4c45d32f1879c5b5a89b97581e4a7d5793a00ecee3dc0375a42441b
za3a258c9acef6f84ffb6e4c1064d1767045ce8809f5176b1014022e4a6b5b87ab3e5000d8c079e
zaca4f30a8850742f90080426d990fe63e10cf9a1fb59e84d537371c6c999f5bdd12af10b31ab1a
z0abb74887fb7f904a830080454231bf4f9d751a4a89425fb2b0c0cabff082c56617e25157531ce
zf017c8ee734b85d9d2140d01d5168603dfcb9819d036bfdfe6c8bffe8639f8c473c9bd632ff69c
z2f5ddfa4780a64f318d2eccf6cd853e32aeb0cf2afc58afef4aa1ede7005af32d20b4c003b3087
za237022965e897f59636ada6eb2d617df1ae3a99e9cdf9c4e50cdffa8577bdcab670c70b122f87
zd7e2d6359c50ac2008314c2256d5688b117b05ff78d397cad2f6cd717df6d0650c3cbd6e532444
z7b96bd4b4c14c67ab3c5cca9b2b818d89f266d7fd57b0898ef225b2acff3b5ea41a055d581e783
z79da7c70d8acf2fb8093aa9af61d8cbbaec0c8dcfddf31e3c36f3e9c5d97f2d6f71bfaaf134e06
z91b805eb5cad2e550332aa8f5bb6d8c89c5204f5986d73bd3a71314e13d787ff1c02065fd7b66b
z3b9a4e833194292bc14c768b03a531f6ae1f487b52505864a2f1c7ced4437a06eeeb469b085256
z50e4e76386ee9353780a58acee4d2e968497c48b5ad3ff78230e0040a30bd7cff45a636cdd6f85
z7df6885e99317f12396215446254cbd8990cdc0702b1523cab76ccebed7f997f7e4900c4d5fca7
z29fbbc2eb9d81777294913ff06409380bfaeeca8d62486161aface76173ea5955f8775b9c90c58
zfdd92b05ecbe478631f315ab55ea9c1c29e62eb1f2913312483cd10042dda7b25f68679f325066
za5110f8827c82625784fe5f1f306bc90af054c9969faa1c7a1a505d719336d96c2e20a467fceb9
z0d518d06dc833cdbd4bdea1af72bdf3a1a97e3b359bdddba3f021ef7023d32a5d00f30752b19b9
z9157bb95b23f755c3ccbdac808a4c78d3c65af2583745f3e05da0bec3582ced55240a386f49c18
z54481654bd0160fdceea6a9f06fd282f660522618c6910f5d2a9712fdd11201d063991a045e97b
za0aae95ae111a0611d1d2ebb9e899ac102824fdd8059258e048dab8a5f1b97a8405dbe022ed9cd
zc8f3292e8b4707aac70543a531c11659715095f38f4a80a4514ec2f261da274b0f952e9fe6c8aa
z74b0884e8e80697cd0e0a0f26d0e5261270caf29a2548ec36137e4d01632fa1bd296c6525f411e
z6a28fa7f5f9b37b3747adfa7b96f77b04339b7ba72a7f477c43d62122318c44a418c884653dd68
z32ac99c1e77eb05310f67ba8a3db1c5d37dee243ea5f11435a9133162a4c9a9c28ae58f465ac89
z864d7ff698e5394351d3080b6bb54177f35edc2c73acd179260957357c73b67035ba8e2788e885
z76e13d750107f4efd2f2440b04f3a7254ae519e52167db9161446c82fffdee6ded4b25aa1dacab
z516664e2bf7b18ff390d113b6cf647f121e7cf4c6d8a564a17d2387c0b9b65c0c5b225acb28271
z590d39ce0d77c036daa84ac3d21b191c2a8db1c476ef7156eae528238514998eaa856d1d798494
zc72e15ac126a8f56a46660efd574ea62d4dc94f48e85662c6efd5101a57a837a3de3401591c2f9
z3477796cb39787466829b2d159504097fd216dbe32f5119f4129114617e55a4ae55c75ad952734
z5480f8a2ef687f83835d910ca99201ce72ce72574fee2496394a5491972254c5177761fe482a67
zb6ab92323ba1ad53e03f4d08a6978a1c8792bd6e34f0d9bb77f60cebe3fc909557de928a6f6ad8
z6e2c3751f5940e38af50caf77b3b1dd1b7da2f1437943c44c8a3c340c11316577e33621409b1b0
za1c650c23aa1184dbb82078f90edd31c253503376ff4fe45eaa898c04ddad9f88454750947c38a
z7a4b48efe5434fc57524f86e5ca4463e365f4ed4661dffa45f0d7b1c81887a072de2206a3c7e0c
z5a334bf4883b5d5c5b09364d4e7c5d73fbc27a5ff5ccb01c9a4249c0b905713ee311020bad0cc5
z5d30036e7c3dd7d53afb8027cd945be3af8cabf0e7bae6c4c1cbb072e6e72cd3dfa7c4d994bb79
za676f733b822202ab7705b1011f9a7c9271f61fc38ff06329bba4afbe3c0c4daaf145ad4a61690
z41269dfbf2ee327b2b7965b61b68cbe53bdf736bee4703afb007e756d8f35baaea156cef9074cc
z0bba0f1bfd7cd4168d1a80eea59614f8800c7993389c85f7679d01338c52088cedc1411f5dbf1c
z579a0d1c96e4aa5140eacc58fdb0112da50afc73b017fe0c45ba6073c119d7035ffec05671bd04
z3355d8abf351a637a64a49045f1f1c9dde6620896bb4bad1affe7dbaaf451420cfaaddab655d77
z5f44f5c995749669df9585e891e22abe9088fdb1c7b1ea59480ac7d2f148f1aafd9fe2fdb32474
z73c0279d7baa7525e92b0e9f69f8cc2ad9f3b8100bf97ed2effc1d58a6336b2185a44069b5f543
z65e3f1bd741de5fb849c77386d9d03797adf46b2fbbcb3b86c3ffa08307274ad598f7517b8b785
z58b13e970c7ad24ec286303242cfbe5f0da98e2520c4a8ff7e617d45eb9716b9bfc5c54ffa6d82
zb7d55ba7a5b7f379339aac9424be29ffea680be7d1e97c856a72505cfee9fb4ec75329dfb32260
zda2631a665dbf0412578a6cdc022f4485f1ce3eb5d3d6024e43c25bfa3602dae58601e94f49596
z5ce5133992fbdd804aa2a3a0dbda799e8a10ac2fe2e1b925bca21a83d526658b4d72ee2eb8923e
z1fe2be8d25fc2951a51a453a58a678600f4a7b4137aeaa07609feac800bf65f3561dcf5f575dca
zc6a469f8ef7ca6cc02bd0df582803ea7879278f754fdefa2199c8f59ca10ea19d4406b7367f408
z8b44f6f59ac17f7ab6a485d20858600f3e573b92cb2f93fc2decb95bfa9f9f5efdae72edb28825
zd7363e03a9201fc4721706d43a345e0ddda7f87335c4bf4991777d29210823481849557bbe0dfc
z9f7430f794c12c6930a157f80585d63e69a180fab4957f1117a69be80e6ca5da27465ef7c60af4
z73cb0aac12833280515957ad6205f984cc29d4b3429bfc2534a287d37b68b7fecca203a033d76d
zf6102de2f661f23aa449db17f1f022a61706233de2f30b16107f1452203d4def1dc5a2f939beb3
z2fcddc21c3e8c59494bd8acdbdeac56178ed72a1676baa811e413b8f702ea80c7f8dca8fd3eca5
z952bb8a33c039cbfa2bdb4a7b3014dec56db1bbbbb7f122ddc838fd825bfb363807c0ae96869e8
z5d5b1aef34a2a034b5c51ea795713b69b4a16d6310c73ca6e4044d4110b87406bee597c959e3e8
z0bc1d67a592424ec6cc1472bdf33383c16a0ece04c990a5d49536d49c1672e198b138b5aca301f
zb9c13723ff670508ce1fcbab300fd8babd696df2666d627e4c87e3c9326ce3b13eba23974ac22d
z8628859a99a27584ff4550a564532ab623d9adb4bcdc26a55c041636c4a95355d3e1f16f747753
z32d65205311937273f51eda3692380d39a927a418f9e2f3fb08aba3ab06fefd24d3d072824f966
za670c195147e1f08812ba4d6267760e41a07206b364d556c5146133a1ab936925adb4a28b28d84
z2763060c992e56885615677b26cb5dec929d2923d9e061572480db5633b5efbe7200f993e3f1f9
z4383a8786c8f7293454837917a7f022f2bf8cd68e1b6739ce35561a30ed67261a08aef6829a561
z576e9ebdf04a8e116193916156196908bdfa37218dd215b7cdaab1fed21ab7e832c5b972937003
zfbc12a2f3a9010952f1a42c3f6c2d3a6171d182ed3e2c44b2a70cf91e0d5f1f54f7367ce1a7fc6
za74441547e5bc4d6f0ed551c021236b0ff552b62038f0ee8fed28fafbea2d921bad2b5395f76d2
z0ee711631d64702f3b60c18154fce8c910fedc00a10a3a1459548f3fcde6fb512429c908a2de5c
zb1fc6d802aa2918cd5b8f15d0a497e80f7fda0006ab5bbf31d414ca90679a090762d243cd7387d
zf69a8a3b48e56d21b509deafdb04fc83355a0512f001b454cb08046d323617a6c2a6e2426c42fa
z1d153fe4bdd7e95f448d989275c7c223a838bc20d7cda0bee8d26efe8e3676e127a212af49c674
z5ac5002a9ab36b04d3d50ec8122b108ca4c273d4bf9b9f02363d0ab4250e0b08383475adc06809
ze303de0803db301577f11c6ce8039c50d0f02b24db6f6351e62934dac3a7e815f2df93fe8e1804
z9da54343da42a74f63b7408ff32c323b70355d31c3caaeca13b478bcc28812737aba0c0382ae63
z24d1268a4f9cb475ddfd90640c2b061a747db5c6bacbacc7c3be66ee3fe1a1fceb58d22181b144
zf936f9895aec4582be171922e356d5592fc087bbe1bb9d179ff307deb32629bcc02859492fa0cf
z60911bf3d6bd940200453c4d16cb735d48f69f1f87a3387f9f8a08ad6b3b5775c7d708272af0df
z5bf32df58a488ad217994cb27d09d90fdfc65b070335273bd3de1109bdd5a68bd17a293a2a931d
zde489262b507d11faba14afba3423170ba324cbf6ef23a00782f6201e5d7304dbb42fcea29b5c4
zccc5ac32ecbc70bd8bcc08c4fae638a97bdc80676649a55d39d904e59e11a8bb39f48dc4193c06
zaa4372fe816764f4334cad62de97dba69725e560188f04262db95060598fd31d31112e5c65fc9c
z1cbf24186ff290dfd3032a4a9593f043cd7d48f76103da69455a3cd9b0ee4ecdc825af4dc8e0cc
zc254f28c784dbe9f36d1dca3fa9a83af67e2067ec52293836b630887decdeb7e604a96fd8c5094
zdde11be733e157e7970bb362c03bd1f313d0c5d5f7377f1db286f78908654d5c44c81afa1078c2
z20c578ad310594f20d4b39a997b7b14321f3e253a4f7f40007698d3c4f18712f7633e4301a7c14
z6e8a85165b7b06c3809b4b266a3725cc864f2565d5bb2a14de185e8d19ae696aedab1497ed7e65
z3b7ac5acd99635dbba5f34b509e0927149d796eac4964eec1d5db9b112158d663338e3fda09751
z4ead8bf087ab2eb52e5751b15ec131cc7c543e2e2761c4699b6cf3b0d44b8185659441f7d65811
z59a2da79985234c97c430881e6db8396a19af5d0855338c11e85fb4930ab2e4d23d4165223a348
zc603dc14065c16ee0d596e84fb84b4c2261389a4c9b64330dfb3e87066446c07ca0d9134210ab4
ze21d3546156ab8cb16a16f7d8f40c960103436b7c93a42e236f5235c2388010f9afd417f75788c
zc8f785a81d93e7afbdbe719e9b5925ad24ce433acf39aa1c18e8a850cc1ba9f3cee014494ef0cf
z55ec11e1e967eb15ac1df8ed17bb36d3565674ecca7dbd77f7b56728afb961f6098b4c7704fc2d
zae20bfc9c12692c3da04901069306565b1cb5abb9fdf4978cdd15560c54dbe5f9309524a9ad935
z34394b9dc984ad2c9bc361f6ad4a68baff17befb5ad617c5d355cc1c00259e5dfa5dd45705c6c1
z07b70d5b7fdc57507beb5379bf77a955ebfb9590ab568766baa9dd9a2504e45592bdb0c3281e88
ze759ab43e4cab04bd0353437dc605f04b1c9cccb5f58ba28a5278cd3cba357fca2881b57d40807
za1f4bca522b7f6d230ed641e8090cb7c66681b9b0867f2d203e34771983b09a11e9a13310be082
z1938e0f6d4bb7df2b862a3695af397ddf11f49906502f307c17412b825d252f1355a54f443d7e3
zdc4d93d70f58c21fc71ec4d4abd045c856863da214f76fa00cf6c998169887419acff526b804ac
za2513b045c4d689b1026496f885a0f9627e1f097cf77b9f504e048eb4e9dc422fedaece021f64d
z3f0ee0d14820a254faca53bd1e2a61a6e4bf0e66e4d266f3778222f6da686198be2543a4f0d591
zb49034578b714f6cce0dce33682b2b15bbd810a633cd262ca5d26f2bb4033ef4d3193ef00a1e71
z5f046dfa0c791672200495eabfa954ec575c1b3973726b88a35bf3ad724aa751bf878b5ae6f95f
zfba712646cd58e6cb5985e0a0e9980abe77bdaa3c48ff7207f37f09a81930c1eb4ea7672f1df15
z34577194fad7fca0ad8618f49668a69903f916cf341ec4637028146506df6a35e9d0090c61dfae
z22fea432c84650c61e94c9d84e5f2ccfc53bda2bcde10e55806686d2cda4c8add7f1d8f7dd3e4f
z303cbd18c6549cb48fb65c74764919e32312d2a6cdd84a5f1bb2813c4ea58839841797e047e525
zcbc9c58b03effba53092b24576c50682d4e5b5254136d0e661a045c93c275ff84e3d9e3a3db1c9
zc16e1c6407aa4c2dd0c00b3ea64bf78e2054289fb9d42aa1ed404268bc9deeddb83ee4a3b15edb
z0634d4e32a63cd01f31bbdb5dd2da320dcac4c535cad4a5fa93a4589fd06e68467cfb274f94ba1
z925530d303e844cf7417fcfe20b88de1436ea061c3028cffcd5b8f992b3a9291723610e0c138b6
zd6dd08dd2074e2cac6ea6d0f153e1d5bed0981bccf87681d62f47f66ebe29355e20753a9bb1fb8
z32232c20489d8873f62d2a8b04a656ad332eebf549d1c2c3a824b9a2fb7547236f8d01121f6050
zdcdfeaf40aecf5afffecbbf6fdb0b8563464015ecc9401a7575a7998e92bd650af8df5d31260f6
zff71b2c61021b80065d6f32f331ad83679a13f8c7ac72084e44ed0c4e506600be8db77145a8ee5
z808e48b9797b7b250e52b1e6470dd8bbe51cc80dd6a9995053426670038ab168d2d2486b6bfb9c
zb00d1decd1c3e8bad50a4ccfda5d6f65cebe33d141a7291bea0a0acf51e0f57f50dc2b7e5364fb
z86d60e6d8e39e717f294fa03b8d384ca03db334d4bb1ae439eb76be5e15c1fe19de4feaa92c90e
zf34c0ba27087846ef0d678e9b26b2730d2e4ef00cd80cf359ba704ef816c262703fb1c4d517075
z0ed44eaab3380daa7347cb34bb7857eb4d1bd6c05778cac660ea8766218937b44600998649111b
zcdbc2097d287afb8da9796aa8945143c3d1e41c091143ec752beb76b55f1efd6c4ad33a31f4b50
z81f29b720252d2990e26bbafb0ac9b1461b3e2792aebbd12cf87b05db9ae0d51c54eb54ef2b956
zbf85a4f0c637b49ecb5a0aacb4f59df6f3db6f8d6ac4a68c70b99eac0ae39c334aea05af80a9b0
zeb897cbed32b005df874caa69a0ea802e01f93d81e24351da3bfae959fab9a3f518cb53eae467e
z2bff9799b522e8af90735964862c9f4ca80574805e9df7e750b94c1edd5a056c2dc530270eb9d1
z0356feebd50b3dd91e364f5d520349d912e535b63899b6a9c07f204ec9079ba0173d0076e4e7a7
z6c4e982f92ffccb1586700c449fbee88b5566f62ed16c123b5025d15a85a1143ece16450dcd9bf
z361e985df46dc0914e8504fc72589164c88a64c913402bac9fb88bba81c45feb35585e6091563a
z34b52666ce01587039b820547b5fb2c3515ac98e3faec28772ca8e713aec6b5cefa05214e23700
z9b3c90119be30a88562b3d0db746c28653c5639dc9109d16d3aca25361fc436bf6640e4624cb4a
z314aba1c59a27c15d025989a61a4fecc6962f4f154c032a84eee83a844e0e917478a9d8baf6fc2
z8e716fb6a85d5b22493a9ae88a2a65681f5459fd426d8eecfadbf87db9f23ca7c9e1ceed825584
ze4edf816ca64d6c85d4b33892ac26168cedba980295c51e4d7d58c1e90d3d1daac57d5dc8d0e40
z4b2c4703117ffd473882c0d275aab7317b589d71ecf4b442e8bdbb42ff31fd091b7041f8ef4cf3
za882272f9ad6b009524c3c29dd5b7f174b27174b46f1e95409da36204e21be3c349fc0ff0c5b44
z27d7af8314246f6e9d9a9350dd3bc12744e579e4ea7e40c02f8f9cd8a61126da216529f2263095
z1df9302749f71449193c79367eb87bed9e435d9a353401d936e85b3d27d20bc8cbef73423fdb34
z676387d60479800c4476191f24d8876d782bbe660c0ca107e1cecc44d95ce56a7552c78e8cbdf1
za1b83ef64e899608ed0ec21c7c7415feb394b17a49f2a8190f42f832c3357d0d983118a82ed93a
z69cf29d4aee51262fde30d4e11da48fcdc36816b90cc0b55a80c15b49c4b6d577eeec262063b90
zda06ce2ffb0b8a8462cd7303437f78c0e9a669909d5b19c0cf948a264ba18e1eba7afca34f2136
z260bbeba2945254f7c0f17e860b0d89fa44659a5cb949449663afa292ce8f7a5ab955235fba218
z91cd59c3130a92e9d13b8dc64eb8445f7ae4503e8f59b0e41cb09430d1c0d1d9a216f5f2e21309
z22bf4829796d0b890ab3d728e0a61a1e1184b057d476bac1533d5b71d01069cc0d95320c47d422
z09ea9e9696c66019905c28cc88a1c4cd8810a72c70649f78a431f4ef4d953de48bb3dfd94c32f8
zed7815d8724b1ac15cf6d3ebe0bf0b933e753c56564fb9bcbd4df10199c106ba5a2ebae64c2870
z035df31a500f69114c85978f3e1fd276d5b8c98e53c477403dc8abbc6491dfb31231705f805519
ze970fb0dfa53d2b57b2f374b403515c2c2cbd001df8f6108bc685bc10b4165dab8bb43bba7c4ec
z060b2a3593d7de483f6ebea62eb14f31c197d07072f1a0d3fbd3800ac1dc801c5888fdf79714f3
zfe79fca4fc99d00561300402a245a45c154573b510573315996e4aa4f221821983e23ae85664aa
z74ab30aecd4dd9c9669b6a0b612ea18e5b926f8d1fec34a24c74bc2fed63f27f59e08917dc235d
z4d1270aab8740ef6d48aaa666423dd2bca4dd40e4770d04db2b93aafe02a1379808cc8bd12fde9
z74a854e93f7da30d7c5e6bf921519b6d7abdec3332a1909fbda8f819fb8f57c911d951c8163ccb
z1b06a7193927041bf4f3ec05dbea1b43fd8f10f36b425356e332391d15951b07250ca16463e48a
zf812730a99ad8349eca2c3e0869a2008df52d1b8a69d995a69fd7a27203bd81c78d0277d87d12c
ze0980db36f9074a2195b2ac2cba2cfc83d09e76e58c5da5639330b210bb9a089c7276ae19b0e1e
z699e6641ed54f654354a447b44e13d70c53a20d2f97908abf577aad0bf3e0694ac1a33635c5cf4
z4f0326ebb3f57a9c6f6ec6eab977e384269458026949f288c151260b3e3ea25c447aaf9a5e151a
z74fe450f91dd99bd410e59fea0c65d0f51dd0c0f7789489c23800539b13f71ab59ea6a3c0dc368
z58768b6836bab77e75cd70973566d22423bda3e07b7b4b8f0367fe33dadccb1d32b3ffeaee11f1
z76342e545cf42fee8c6cf03a66cb9a5c834a3d4c6323fc0da9241de2a958bc002ac44695cec1c4
z31d0a93f5bb99ebfbab600ea1ac2fcf622690219ff570cb2b9a3e9904a19476ced6b253b66c404
zae6b96392c7d46d1bbe6e561129939a5a44f4c19120f5ff1997e6c4cef25d9779d0b69d38c4c62
zbb726ddd25cb75692db0c21d6e10f40bbccabc464b72986f3a6e8417e2fcdd2a03188ebc365b20
zd8e238117b60a0420c6799468b0048213135569783b90732d43dc0490dfa7246e962ba834e6e3a
z09c23ab4d34b2a49ff0adc4c5f637f86abaa62f19c984d814363ecefbe27ffdb2894b785a44256
z5b3882e110c1342f51f8a48cf46556811f1d50b8d6878f1ed2213b1992a877a7246d9f978cdb9f
z0fba823a0fde97c0c33d2d3c8143a2f6c7c953afa6dd01001186a014ac65827140fb4ce5d8e017
zf5825f933937e0b3c9332f6a2127dacb0762dbf3b7196edccf6ef8bfa3d38f40f5c756449efc79
z301ddc341409b6a3fe25793a5f8479a6ea01a23c8718819bb17ffa40b1715935f00037b7b896ae
zfe33263565ba98f0c9ffff6238eb5689937884cefaf5643382224f432337535c83d58d48b0ae7c
zf39376e7e4d6cac4a464f8c73243bd1781f516cb240cf8f77aaa63f9bc01abe9ca86d959eed5ba
zd93eee0aaa94208e4aecf7025ce284b2b6028fdf36e6e2763483caf45b88fc7ae0e0ff91df6062
zcb0c45a958a0828494f65ef264c14f9ca8a98857fdcbc21a6f905692703af4f4c48454273f9806
z8d9c6280c73e00e8f39846b4124a16a610964d557342acf89cec8cb5254a86936020b71301dee9
z312324c26994a10396cc49799428313ce596418050913b9256f3a6aae5b2e163675b4929e47ed9
z73c32b7e0f6f5aa5bfbc678a4bf9bb583d2f8f7639a2669e92b2f301e329a877c03e544f8e4731
zd6803fd911fd78a9d6f545585754a58bce95e46ca779234d58d60defa736f204b1071dbf84cdae
z174b2e182b8c9ac40ff2a5bf1c591b9c2300b1077232dc1df088e80aa8a4eb62d37b2c995fad1b
z5a6f30de18ed0846d30a7a233242780831119a3f5237ddbe634852a3df97db875ec8fdacd9d35c
z6375d2ef318a5e34efce4cc2a30712eb2e7392f6414c451344b2c3e0e5762370b06951bc8c888f
z3da7260c6b1b127458cbb16656d7a579d061c305efb9ef58f04c900a4bc5fc1d39e2301ee67573
z2fda7ea569e592d03d1c51c2998373419343b4554a5c0ba1f302826c7d64e1ec90c5eaaaac2cd2
z0a62f24ff1bbd9a6f09a8a8cc7698934960f5a2489dc8a9d95b5d7ddc0384d59bf3226ee86a08d
zdb426cbd33d4326a0d411a373d4317d496aab4eb7901e0a1d941ac642d294cc8e0a2cd15c6ed62
z51ba55f484c272d571ba413dd3191a8ed906f1edff54dcd619c8a6707c60b926cd4ddc97d34310
z43fbf282aca710a84edb3e4d5140c7866a1d95e669b3d579f51f8f85215a85647082648bcb015c
z408e8c9260b992feaefc3f16a0144f430d3bffc60a8f69f76609d60fc67fcd88d9b305fbd28fa2
zc4e1a28bb8aac0a0937da81d29d5bed0ae1b67b196f6c92ef9dc8ff0a047708959d74ee2ee4948
z16ea47e0161fc33adfaf22a4bd2b17f59392db98a962db32e2895f79123503aa475b31fabeb666
z86df9cc6cb115f50d640de18493f7f48f5b3ac71c0c8e5c1d7f4fc83a63c64c445949a39eba984
z68bd799190dea8246a538ee6653eb27c0aefda48ce0e1084231f5f480a1bc1070ea3fc3285606e
z525299a00145d3ac1c7e19811fbc2c4fbb65eb0546590995917374a1c57fbf7a0cddb64cdc38ef
ze6a1efe5bb06f173dafadc384f9684d82f27e5e6d0bed9f64cfe929d82850f1bd287a23cc4cad0
z1bda089377caa21d32aa08be3e0ff7f5b8199675b7d26e2713c63078cce77b6aa652bd128b1423
z56099cd0b129634a5397a5fc1e802816e133d05815b717442b943685b5d400731c6994f2785738
z35784f55caeb8336832dfe8ab1bfa377ae7fad8eac3ad1304cd221c9fab66023abf7fd5e0be11a
z6404b06d3d5dade553876f95099df64a6f3700c7111757601c58912046ad8949a630487fa98658
z7e445f5f6edd149821d6d7206a5b04f89dedaae0661a7a46b8af3cebad45429c480ede2f387a81
zf4b26ac6aa00037ba114927fb216590a676ec3cdc0331230d24eb2309294b42c4cb6210a7c51af
z68995bdda6ea2ae862c9548ef8b377b6fb5a4f9f2b0854dfff5ed8dbc37a1f248308fb76a21247
zdf16edcf4e1d727e7439d049b19a2932fb67a1b3be458d942d13eb5b1a5a12f119052fef169a51
z6e6e095d361f5f480f2b687e0ce3e8e1ddc0b3bf2cdb7a2d993a29e54177acf5dcfe58138e7419
z728d0395110a2a9d47ab1875c41ab2daa7fb5b77b20f2d9b369eac824770542f248a4ddc0bd56a
z4fba18516d388592bbc620945b78dd9f9033212acba16503574a1b5c7699f15348325adb0e5ca7
z1104c3efba66be7fc055a6ef6cb693157ab643d8525e40e583cebca64837487db1cd72fff0820f
z8bf9aa087eed489ae1af90f203ec688d65b9e6bd7de25d2a8b8d729e51bfba0f572148c125585d
z5fc9190639fc650c9e80da006a03c7925385eb613c9656614a6df933d4fe128094b43b13bd8c23
zaaff231f3bb6255d6a2f9a57375dd0e7362ba1484967bd5c5a7dcb8c9bca574e490cee4a6b0bf1
za5fcd566d331dc619041989babc87b94fa8be091348fa06563b1a693da367f6272da1d5af5bd38
z44ea609c17ea6a10148ba926336a7786097fd91410bef1df6ef6916951d5c8070f41c161421d7f
z147b9601070c47c8c9dcb0ce9649fe5e4276ffb5aff287b2c5a516a85d80584d23438a523ba6c7
z62817a9630021e46cfa24739600ca70250e6a2c73df1eb5c35c5af7a2a900c28d96c39d97ad22c
z4cea3ba7b9eff16f26f54f320f18657a5ca35237cd90a6f7c2fd3c453b4aa52cf32afa4852c588
z71e3ab2158c58b8245c241fb27e6dbbfa0e37bb9af067f73b04b4ad23c22a7f8e092374457efdf
z287f39ac10f9e1c5c34b7dde9169873256ca97a310341e3d428a38b16acc9450ec611abbfb489d
zf0f07a7dabbafbaab5c9a479be854c585ef9e56c0fef52e615893481b7dcbf154df884fd67d3cd
z2a7c7b33a5ca9803b882ac5bc95c0d50ef04ecf1b328d99fb7ae22649a8af33de73253bcf581c9
z868388dfcbf0a8ec7c7ea10f98bbe15dc36d63ecebf04e826052474423cc27246bf6791db9e946
zed339b078c9c883bdc5e21c27a4a89669b93f5b6e0a507d8f7a65ee88c2d6a623064ea9c6d7690
z6d1b5e3c4b1678eeab708ebadbdb6151210450546b5bd6077fd449580ddba07cf8ba4d489c22ef
z26e9801c204b2fbe4c6e6bdd3f4afa6694e72e2f8ef98698d9d6cb3d8ebbf841e0d95975ab7bcb
zbd50a6f777b52efa33f2085d77542328454b5ce16c06d8e1331499477b77950de4bf92e48550fc
z18b86649f46cfe38257977fbddb17a99989fadf012d3a08a3fe016c549ed264918ae3ef0f28b01
z9ab744a9d4fbcb648413443f90ab005c2f6d43a16e9ceb64ad22ad03bfcee36e12c00118afdf07
z583be9c99143e94e2af6cc754219f08d9d7490915e97d83c37c9817bf433339b057e5d2e7038e2
zc2c17727a5b9766a3f61ad5a80a51604d5de4e78f71f46d3887ecf49c88bcfaced98f7f7be59a9
z900a98f1e5b4599cfe16a896a27d9b1d475010853c49fd9a10a58f98f6ad4b41f294608ee1a08a
z103953ffaa8b6462eeaca4d11d4cb527a47cb9124eb8dce1ad7a60325b2a2563dd6a65e4b2a189
zccd689a88b94df5e7963a64ba00e78263930fd62bb126e03ec8dbfd853624b83b31dfc36f5dcaa
za81b56d88995ca366e90652924857f1919798a587ce3a83d7c7572f9a72d20b155a453f53b1bd1
z4172fb88fb3b126209fa4b2af4e296099aa5216b69f0b7105edb6d55316c09774cba10d5da11ab
zf2fd6994cfcbeab490aaa30fa8d6031485544f397bdf5327e22cd85230d73c55f6a1ef123a95c9
z16ae718174971d32c9a7c05c342e2a9becf3942264cb9480af1c9722f8a4c4d318373064e50bad
zedf5f014391b4938e42f5daf9163d429454db76404da2b7ae91f6a0d936c62641a9f82e738572d
z9441513b811e72d702e35f7ec73c0d14d0a82bac0c78d5a92bb6b1164d938a9ece79bbb2b498e9
z31f90919fb4ca3c803e55c3ee2cbbc7b349a771bbea776d5018c10cd7aee4e1eb2fd7602d904ed
z9f3e49310b16ab02a8ed31999d42784c171e1832b14ef177244dad691ffe2a3044f150f93ca36a
z525822cf2b0ca0f065e31efff0ef322f1a61ff7971d6f7b2c715c8a816d12f76a746b1cfddd5d9
zfdafdda8ceeb8da3b2ec9fc83d2f83573010274a5f19b33cba4d597055b169c9027d2fbfbc8121
z120d4a695d7e650bd188bccd0f66a22541fbb864925663db29e8e9542c6301359a4d536c75411f
za3e06776ab1a2e329d5f5c803a71b55a5e295dcf5ab13f499386d818a31876850ce4ac7163ee96
z93a9d93c2cf0985b11aa2c12addbaa6ea2a236b8c7835fb1c9384af553245441b88fabad700448
zbe4e9ddae90b39d0648a7fb8029bfb5329971ef039bd8e38ecf2b5683b43ac0a9e967ac73def7f
z8c10bc80000b2c6425f9306e3c2026df14242a64bc1dc2f03f4c706de702da744ded325a8dab8e
z397b493a4e740e09acabce10fe0b2d2041777ab5fd7a619d7574aebac2d4495be8e0286a682821
z34545ac7ad040b4e33e7172a8efb967f0e6205cc0aa1d68715b574d99231b36a1f84b087218f22
zbdef07442f1230d238a5bb48ff84f9f04610a25d91900b8fe2a6c17ab8f15c01c1c0449404b5b7
z0703ee0e2050ccaf98c8e31fc3f5ec9f8e610c16b47f14ace63ca6e53fd21aa74775c729bb8f4c
zc614931da122c7b03441699fee153213cac7d071ab9c7bf982e99f22d196bb7fec950a66434a0b
zb7009b604f06ada40f9ac01f70572fe6937e465d1e544c26d760e78956574efa72a530d3d1d608
z39bdbdc51acf5ffd89ebc14d517e60c0442d5c0c09a4e9d260259f3513da43937740588ac99c8d
z9f15852012127378bf14c4a77a48b07f9fe8cd2f5ad4d29166866e583d3f96614da6fce9065dde
zc892c1e703df63fc705f00e9e49ba11170cf10cdd23a2cc6c2c4e39437593795335a5a76d2ec4d
z0cf499ddfc95b53f0884d37c13820b741e4cd7dd21283a9e4772476731f7af71466a509d9f2d97
z3326d776053d6623f61868dee2e0f0ce63add5e7f27917db5c93830917c8e6118c6e10edf8f1a3
zd74085b0a1445a87a55f375fe37794aab9a47e2b987cf5cd549b5f1d7b637079d5be3cec2e1898
z033698a0796fa237a9eeb7898c595f09fc55190c7080bcd82121823316a6c74673bd9404d0d665
z79e83a8972d96e1e12b024634d59413eebf219fed2d8f2f69567b122cd713d4ae3480fd7fdf6ca
zf7e01f82d89425d39174df2f573530c2d458676a385b608198bd0852bbac89abe3d369cb1daee4
z9f9839edee4d16ffd16344a8bca44e74f8bc2161bdd0623464e157a2c6d8a6b5e3f86b27032a44
z5f640f09c890ec9d67f471874eb7c6930c77ac6e2a8ea9d25310f444f7dfaf2d13ce8f91dc977c
z6930e88e3f3c49538c51dd8776656558a960f1b0dbef1546d7b68d90bcb16226c0939470b0c508
za8fd87e134933df5e571a406457ca7ff62d67a27b352baa1f428987cd4813d5dc9c7553d184df3
z74b0aa10c7c59258d1d686a158244aa6b2310fa395e07ffd8a6d389878d5c3956e51e226bcb1eb
zfa2274e502ed3655537e140a79eccd83181c15deb5500f91de978c73687e7f84cc153e3c871378
zd0584739e35e71132fc5cbe4b976053791d31e062bca38e7bb8755c0f6794b38fbdd23cd51cb7f
zac08d9320162d7cc665b71e10f87a055a4dbf9d40d87ef776ebfbaf21b6a195d7f576802706e29
zaf7439cf9ead62e2e72cd415d50cf05ef0072168ef96cd273db4ac0946cf54266c19f539a9665f
z4f0b9b6c9b9a17c61694269cb6cebd223e20f00e52097bdf973f7dda060ac0f2ce9d929736c0eb
z44736822580506681ad637727853fe5a6bf850e1fdaea13cbacd3f92abf078d8ac7c7545adf1a0
z7409f4415b3c92355566ee9f6e8e601e89a357ac8e42fac03b00089a830256682d516b890322ea
z1373f1e124959b06f9980f527b9a0f1c1f1bcc7bb8d291ecd88b710d8d50caa622334acd3448c7
z7ac4fe7c5d474090dedef55d91a49beb4e9ea5e59ec6ef40f2a52b5f9088702c82f03958a629dd
z31768af37ff791b023b5308e21940ed8b659c8ef765f330c4f44df1ad212d7bccfe61b16e6fe9f
zff5ac5c992b6239f744791f93d6c68c82c30a4877c444dcfe91a801828e2ad063e10fef1242e4d
z9e9bac98dae661d2b2badd51675139537ce408403b1ddd8eee04f1c913cde87cda4b27e9897b01
z8efbf17ca30cf0508d2a7fda2fccd0b647d7cb95215536d731d208bc1eb25178261353a2784fc5
za6c360ac39935c76ffd486f3f3042d2cfb489e612ead1fd7a5b4e10bb424a92151d207c85a9fec
zcf10010271592bcd58814c9864d97721fb3d08f826b3b1b320f33858f6d523205c757b9a30ad87
z970f8585e6e112ced677061db1f685871861347b166fb59e5f4cd169e56243a0719626e868ad6c
zabfc81b9ad83a4ab6da3c4db66428f7f0938fc8cf55f3e49b27069460ad3383475b5376761af35
z6f15bd99db53cdb9001350a9f6eb195d8ce2792689d1ba1d562faa1240976d1ae7e83a6c8da882
z1e03fb7ce954ec64ab780ef2dd47168d4667a33dd6fcb0eda8d5dfd2f42c243e916a6cdb480038
z2b178a77b915fa215343c6d27d38f55a20d6c163f3531fefc6422bce050e978aad831fad3eb61b
zf3c2b628648df5d315c7d7c3257799ba62f54ce3bce428580373c4987f3127030db348ad2fd49f
z40e4ee7757f3d2774ef833a40ddd8d0d2aa5c9ca98efb3eb0b0028be0c1465856fb666dfafbeac
ze766df974aa59bc63abf02a5c86ae0c111a8de6dba4cec680efa6034800567b38b80034d789cec
za65152b28a8eb33d5f36ba3a2a14d28bb885cb7e9d5e05a87e0f5fff60551b847c62161b0a73bc
zfdba8e8b1ec856fe17c41dd556f9275c3210b5a6e2b1576115de17d94c2d2f37ccbbc89ed93bf8
z3778fc986634a45e56ae94f3e315d997d98fbfaf533dbbe57057759ca6dbb5bc773eae7f7cca10
z85409fec17c70093bcb8b3393dde8d750d2732d69555c8396526bf02819023b5d9736ed21ae221
zc0e87ae6bf1ab04a740ea9c7f63cffd77f9885f757bd8b9d851e533f59c7ce55ff0726f4bdaf6f
z3ea8193b4aa23c6bbdb6028bff89fe213ef4fe6ccaeaa0c2d8672fb8a0402edaee2555e0176817
zc826aaf3964b7eb16d75d4b704649f3c04cd5ee5937a29b8e0c6f79a0efb9ce4ae54772b8d98dc
z6c65894ce002a416aae74e28dbeb60fa1edd6f3340de5b6403fd9c7dbe2210e582d2fbc9c56bea
z838098725b1df16cc1aa86c736cd5606da457d29458bdc072c353f5b6502ff2e8be24decbfee94
zbea380020db1da45607642b4e49c254dca831775a5f775f3c95507ffbcf7b3698a64dd80aa3d8c
z68e2564eeee3dd50c4bad1ad5c6d6ea41125dcb7fb62433b698a4adc9533cc3e3c442da8470842
z32e494ce9a606014a3cd66e99f3d05257228fdb135324af8b92fe49fd37a5f2b7ef066202a676d
zc4c3f7e669edbb85dbfd03f9d844d9ccd12e6e92d2a7db2389f46ed7af064c79f63bb60d8c8b9b
z0d566405aac20357756b1ed54d94987cf826dc4bf74029e0c0eb1794adbc524a609f62bf7b5d5a
z8cd72ec029264299cd380be162ea691dafb8f98095f65e78aa14a1db750750f565a780d5edecdb
ze24e8a3ecb539f63bb98399ac03954a5153b050234ec60b920d422f8b6181692e50652d8596302
z6a304f4e4c0d19f149a6443a8290da8465c50544d2299416da0ce7ccfb37081b88546a6a4a8f53
z6f6d6a319d3433720f79a8de4c7e185b2d6e6980b6487f3a6f2b3dc6a5e6621af8edc47633c657
z9057e7ead8ff595fc995a94ee6d5ae4e207a99adbcda161f69b83067126e7693602632ddfd012a
ze3b89384fbdba75bd3039da68ff96b56a81c7a6a4b28ab35c8146022a925848431655c423fcfd3
z6793c9aec99ce3e2e7f06af403d58ad5a36ae19757d764d9dc3702f6c76a20f5101c267f8524ba
z69ed0312c18e68de3a0b3e1627bc25a1c6ac67a1df5fe0c6861c290fbadba88e087962eab454b8
z0413eefb31a4b975221837b91fbd53136b766d1c2a29c831bc79913dedb8beb8002dc225b59981
z9bfb1c7666a4ca133ac81b6ec99086d3ca94d1ae1e0f0278c509c70ba8fc6f13bad9f3c928ce89
zb71e10b4b667acc8697f2330d24ed302150413a6f2c45098b57277634853ffdfc28cc5c7cc9c0b
z8d2d7bd52944521c9a9b4a45425954d9c40e82ed2f2f39ee683797da250e8dd47d56bbc6386b82
zffb8b1abbbbfa7e11dc0d7d4502f123ec81b25bc51c3f02d5683a6ed9eb97f35603c5d67b02194
zae08636c4ebc510dcdf18c72bb8f2643806a4aa20997349fdc17c2e7ba19636199481902a5145e
zf2a398586c7f7d6e5d5bbb827cfdd9612252c47dfdfacb1b906819223321d5a940fd9cc86e2396
z53117ab718bb25b7208a738882d6f61ad76466c80f4cbdec23a807406d3ca1db380529f4e3ea26
z6c6201571475db21513206608089d3081254b4ad42c73b5092d76ebfe5f108e267e04db2f35cfa
z9c7a768ab11fadfa78f0609c88769456bb4f2131743980d2d59a74639710f6ae4df64fc9ee0328
z7a2b3fc1fb3d0c5bc41bc43c9b922bfe4d8de2038b8d2db45cd4b658864d172884290d4960b9ed
zf2c009ab5d6c7484ae6f721784294a5bbabf31ac33f0c0cfc0886c1f20942c6f8b05febf804fb2
z8e9b8db156014b4baabc61ec3482768c00118854d0a5e62f41ce5227037d30c1c229f6bc12e6f7
zea22de2e27ea21a28b23ac00cb7141659d22039039b314ecb4a12cc583634940a4abd8d23bf9f5
z349e1f53022a1c6c4fb301d4364eb6ea5e437c73b503b2788b2a3669734fead1c6f8ac967ffc1b
zc43469a00b2399f3e29a20da495aa010d11b480c01e04ab9407d8e679ef66113c9215c699a8ab2
zc764f2a056b6d2b6c850b0b3a7d8d8c9e0ba2ed694fbafb6d369dbd90ef91979956f2d98c75479
z4eede2f881e51e054ca41f3a3b370589ccdb705b3575760a51578d81fce65373037258de8b2544
ze0a3f5ab20fd482f2b2e69106d24849ff5b0d3f618e5ae7723f849e8b3fdfa95dece4b69007be8
z22893332ff682b5aad7fdaac68350f8999f43c36663d290ef79a72046e8afc332ade0a5b4660ed
z61bd5b2dd491eac8f01f20173234043ad5d795b0e7925538be4d148542615218bb5214ec76ac28
z4d71278cac750183e810af3a16afdc5f0adf145e228d05a999c0fc0fa85ff206432aa0c997b8b0
z3945a6548098c5fe8fab4991077c8decf854c31b42057dcb4b905931d1bfe02937d2d5de2eaae2
zc4c81d93633588fa90072a8162241da94275cb0b0df332754999c0aae67d613f3c426c5374b1a3
z4c46eb6d18c3bb915a0e3d69f175a12b22b67ba6099809d308a013e2e34000b57abf1ffccb63ea
z9f81931af405e474bc968d4247ac7cdf9a55f76819b0cadde5d61a5a7707cc2b80c366baab5d4f
z044c87bc143b85eb33fc4be5ee60920c4dd381583b2b7da5dfd9cf11154813531af4518a9c8eb0
z9174c7164fc8e1d5d84de26e12106bd66e88f675861ff8e17a9e0406d5776ef72269083d9093bb
zbadc32af7816f643ede6efe31182cd3dd01709078d73abd4322537c2a265a4620f2bfa11c3779d
za799f70d86f2a249ca4ff478e2282da2cbb5c0ce1de567b77c51e69da7f547e7d2e57d625a6d98
zdaa976dcedada6191abc52353367184cc526536d5d8989dfa60f95784915340c7d5829a6beac22
z98e08b086471e4cb7224d87da70d171c61886392e3208bfd17b3cb8b67aef730d645c90b3d62bd
ze5631b7ea7ed92397b79df2a2d4681be58d7e884bb8e59113204dc53f71fb93ce9a14fcc59ac75
z5aa4326d27d2e4fb2f5d5549f2cebd70301d2187fb11b5afbf03f5184b667e77161c01765f7042
z18241b0408094f7789d5e6925dcbc67b28c05315a4113365d880b0e4556001b7e2cc7ae2153409
zef0cbe78da1bb936a952c7b348770d84f392831f3475e6023f2e13d9fcc6cfcb878fefaa69b463
z5f31714ab440f8741f4a09b74a406a32e490401211d4a41c1291c9d9adbec90a40ccd94fa086af
z8bf721aa6b72d4e325c1ad1041de642996c2328cbf3378f17f6b0c54561238417cddb981eed105
z2927073057a81113ff70ff361382bb113122a02ad46f9c0be1bfddae5e3ff66d83de2c1cb5c727
zeb7bb91c623abac37f3394b0f0e97d217c4e1155353a230097550ef00b9c47ad0a135bc2b5f16c
zd3819b3b54ee0b84c2eeb6531ff44b82e42520d7e6d59ae17ba544816372a5de184c2b9e923472
zea85ab9ec22876e9efaf8ac5fba0aea2e17e6d9bfac3caa2231d09ba1bc69a7be518f1b0620779
z82becec4ea671d0bfdecd90278df31e6142d133c21a329bb6d6c01eb2eb3b2d1dea8450634bda7
za5463246dfb5a1d3e8df0ea19fe36d6e7e71fbc9093322eb39b5e2013c3cdfdd6a27d00c612e44
zb8f2fe69dc63ac371d23199eceb292e6542317b02d94c6f95c7082ffa1556459b81c9721b9ac0e
z207a2b2673b55a19c801e55eac393a36c42e8aa118bfbe2e021772b943a7e920757ef548079a43
z9a69ff47422c6a6ddaa0111baedbf5bab8a54b06b956dced174bac06ff52ce19deebf02a5cf259
zd078bc668a08634a675e096ed1a1cb51f2571fdfa39eee2f999fb70b5b1426e1e7a47ebf6409c3
z648f7d19b16af46c81a746200031b0fc90bb72b03426b00318d82680f854569ccdc6058f312d20
zb19be6c96f87878e6f5a117ee37c04f71569190b138c4006817da7076826b3e63459c13f39f3fa
z4cb9e7f65593722fe61a432e51f2ac90d5103eb9b96d84b948bfbdd1d51e466e4fffb39afa2c89
z7b409f39a4b03a5c6b64568c7bf8432a44b83d1c73251bb5c8e235f0e62ddc183a79c5ae895bb6
zd02e2953a24ecefcf97341f257467975cb444466f49251c89452339a73487a728212e45eb0928f
zc3acebde7b85aa0ffc7104b117bb4f6eec06fe89789e3fd3a2d6b49635b4cea8c10ba95918ef36
z82257e2949bbb38becac18bca86ecff23f23f4d040ec1d71aa4bf1da65103e0d5f4682bcc59054
z7864041fc7ac757d775cdd9a7d278bed32f66edd5b029cd3f817999c90252354926b166f82a752
zff7594c678d18b26b51765cb0ef2f385d27755ba040d03ef1a22fc4cf3da9e1bdb4da6db163efd
zf8596e4e774d1662abc33b354a47532293be38a2f22720e2541a19261aa2f3ecdd073148a7871c
zaff10fff75911d5bf82efeb0a30db34a0ba44989d62e2a34da80d31c01b5736e16eed2a875bf9c
z1c5de67b8978287f16e6a4407c80ef4d7219a07b6940c854bc5bb5863897077fba6c409d952c29
z2ab80726a6713bb5f5d2fb6442d4bea27dd714044eff622ac4d01106fc0c2af654517fe90efc29
zd1573cb918d3a9c52ace1a9f6db19fff0c8b5e3555e239e49e1fc1e02adf6a987c68b3d19fec54
z9b1128c19142a01349f3c8ac107a5322cb5758afd7b00a6d9fcba655bf9c05d867956bbaaccb61
zcb4de364ab62055d167e21da4e56cbd98463562f9b113288d046188556917e579c2fa801672491
z75adb13821a53b2fdf463c80e97348a8f95317c0e3b9923ddeb2b74870a506e877bf95d73d18fa
zd2218b35f44ed90ea915caf7f50450eb70a66177b5fa347a38ba797b3631e7599b703a44043c4c
zd91af650fb2c494e04f790b5f040bbc9b10efccc7166621361044505ee2f0e64f0f2b45eca9021
z1dbd519a5e1dd09feb7f824a4236c9f78fba76a8174ae37e7aa6b28627ae651b27cf2e18df2bc0
z429ab2a9198a5b20ae4c3f95e17e59a94e2fb3578eb47a125d2b72f3f568780e23cf8cbffbb2e1
z02b3485f5b5ddf909cd71ba5431fbae70d6a6143cba9ababcd0e34894836cdcceaf9bf7c861af5
zafab20b45065a228d83d87971a28a03f65301302bf3986a168db0c6b89ea1ce36858758f3e8aff
z44777956bb3a25b0a47f91fca18919e379ffd49e742a256635407dbe6b73e317150c2ce7314e3e
z8adef68ecd3a6b7d627dbdd3de8c970855737f17b071d111a74dbfd7b37d6b54b7c6f0aa9ced19
z138a2c942cf1a4f9f9bbc2e4edd38ee3f914a6a08d19f305b2b7d0d6dff385749bf7b0f2abca56
zb1ea1abe7c8120c2088d97fe9bafbfa36109e78f41b16830228774f2d92896a557fd59d3c38bf9
z10a137cb672827f7d01d3ca34e28e69998163dd8d2fb88af45b434748a852c3c0d95cf98ef1292
zb13875176c27b289f1ffefb7e329edfc8e772b46b64073178693ebf1db50976ab92338fde0a2f7
z9b7f37e88895121d49e55b6d50fd0764d51c23f2061cb87329b7cbfae24af5fcf212d6fda21b0b
za8b65635dce85f47565c445a7b40f497d2ac5236f2c59462b97534a6c65399fd99d683f203fdf9
z7f29421ae6b1e085b589b26a4fadef11f686d43ed853e95cbaf17fc0d72f522d371071e1b103a6
zd2b101882144e43d9dc3252f6fe6e0447b3261cb7fa8a6a7b8d7c6d3b783feeee22133c66ba6d7
z4ea25c8ea48cb39906b57bb95f73568e23c9f47ac60bd1b654b949c05aeb279e14a03805cdcd8d
z4c446c2bddef51f10f78c4c0b680f77350de1f36e8ab70725c7b195263ef6f7252b1edcd597b51
z89229cb8903ff759ee63ea8d9c2ebaa4919da8ed2271497114938a908728feb1e65866bd9b110d
zd19464e9dbf9246e7a8f35243be54c3a6b6f740a6a6f4c516951427a64b4fbcddd8659bb28428e
z1ad88e096395a15e52e6ff0c441a67d17e1bda261cf78cfe33f0622c17884ad507003ae2732d72
z439f85b960f84e2bf22309b4176fcac2f502134efe501c938e4e9c10b5ff723950e280c09f2ef0
za170df0a93617e46685bd5265b850597bbc3696164c9032407986186f56814172583bd984e13c8
z9bd2134d1eb7319c9b6719dbb635638a6ebbdc062e5295731f17d1653caa895866d5fd0f787efb
z04e7590b306756dfe7c49b3197ef00c155e1a241230462295e6ddae117e96ee674deaedeff56d8
zbda47ea73f4eb9f95e9cf11c4e8c894dc48ca211ed961189db055f542122bd76885c8a48a1d1c8
z6b3230e9732ea784c06f8b481b1aea5920260dad16313d9e083060b23c1f5cde6bebc625021f28
z29bed87cda8eaef5ef0fb9a02a9432748afdcb6604bd736876cfee8c2f5ec60c32ee6d7afd8a93
z46fef1b3e2619280b0832a600980f6d2de22069ab6f6ae25cf14d4555bc375b32386481995a032
zf06d9a723f816e825f7d9f225400e74d1a0e82ae5babe87dfadbacbcc945f622c836c45768bdc4
zf4478496e921701fc50e062675166754fe413acf8a1b5c844d26fb8b8eaf33a95d24c3665aa1dd
z55dee269ffb87cae43dd68db0ed9625323d1ee89abda7b95144c957294354d44aea97c3d442b2e
z4ff98ebe0d6e28185bbd13e94371fb4721eae4aa2aa21e26f68ae7c7c304ae7f348740351106b7
zac80fe4707c702ad6ecadd970136ce368262ae15b60c99dd38dcb1fb629a646d2a073887edd62d
z873b5be54b101536b74120e855dce4f3bd29313a312527293d205cb200e12e66c8c8924b57f429
z8378a715b9fefc270cc91d80ea2bda3b53cb1d160ad11968e6a70a16b4e23c3986d90a686c2905
z2183bed78fd3964effa9169d8b3fd3efb9d2d0790fe5d98b1078b04cf2ed0fc61577b54f991c14
z31875110524b699fb7e3ccde1a677217e09818d3adc42aa757188d8d1a260506c9253bd404b3ea
z7af36cdb9fc809ebfa47a2753b82541e5994a6f0654924b4eab502249cc92181f1e1889c56d5ff
z86ad4336a560b6059b54585c9af319b667d92ae35441f04b6abb51693ef4b2e6023a5a503754d1
zf9a7dfb155adf8aec45631ef06a7f00966b741fb5175a0a29de99a6d6f622aefa77b28058f6de9
z5b490e735c635a9936ab23c5640cee1882bf51484842f6784f16f1442e9ec83b81663494293093
z3a77dd9f3405373136c87d51e6e7ec29383370a6f102ba319471fa9b0be3e82b3c67bce1eb835b
z0fff507fb39e46320e1c4c644041cf5cc74e53c149bcfb832fedd9b7d75781fa1526fe2c56a1c4
zf4305efb00998dfdb57cc9ff701019b62fa9b6ad3f3bc7deff7652db29ee3d9699aa5a89f43172
z844ac46b0f32c583f4fbda9b449711712ea588f6aaed70a4e0403a9cd64fa7c9c3d478adc14b1d
z4491a4b2339b4dc33d7b46d0b846b6df944b9770887a1655c79798f86322430e96eac5005eb1f3
z8f1ffdf911d69475647d3d4e67b6e2a24d450d8bfc33d43aa8de5f433a6e597ae9693eeb6a1c15
z934472c0e49e01241587e4ad093d303c9b00dd159ac744173e5c648de70311927c63e048f8d40d
z736c5a80e40473a25732ec3391eb96c2d12ed94e1ad136ae02836b29b0bca470e57b0847fad3f2
zee5074098f822fb1301096b36d40d0e4159a580e7b9dc3ae1f2538ef3d97a42739067156a40227
z7d62140186c867c53c60063d93155d90241ed1747caba1888977e79706992473066329c2d763da
zd236c37263f4d19f3c9db80747ed2ec33f177dac50b545abf6d2153bbea24cab491616578d6c06
z66c19e46003ab7762abb8c3b5fc005ce286b3b6f2be6a7bd25486fc20168b5d4518805560ca7dc
z3f9af4073ad79f3623c6d7971e2485992105f2cab22f282ed5a39e518b00365f385262ef18dad5
zf3622274a1b3b673494cd6caebaa24294c0917aaa1b492af53d5a7688e35b2b232dc1a7da2e03f
zc406dd8a4a3875fa4e7338e4685b6eaf93d5dcdfbdff5765245764cbbd016f2b4195201efe01cb
z76859582b6d71a0d37a0cf7b85a7fa0ae1728a4a342802bfb9c67eaa5967bffdc120c05cf1978d
z0d1e1fc34afc20fb3ddc3114d2a9b0dac2a89c9cde5f7ce7269e04535ee94c1ac500dc41b6c503
z15595c0fc78d462a07919a860f99a65b85f32cfffbbd201bd6f171154492c0b2aec01b62f0a1dc
z12150fe5d7cba30a1ec6223eae4dbbf2c5e97e089728648c01372c55fd37b8429f8e6b6dedbe43
za3aab084d7d2b37b6c585d8f1efcce1c06d8c54fa7514d457dbd99c1d421ffab03194128d42d08
z37286d4114937325d949dba8cef4cb6ed44c29c83187b94c71e45f5fa9bbbeb063d77c68e2a569
zf22b638c4d453bb5d557e5835202822b70e588a426c97f341ec4a49bd0f7463264f326f8e9a8cc
z686cfa60b8d9b26a6a011432244f6f121b0eea5a3794d142f30d001959847f38d833ce51753937
za8b91e465e6cdbbf6110fdc88ff635defadc34c7bad6daf6de9577ea6c1d6f9204eccc2a999d8c
zae233285f8fd4b57801bc92166d7271e359c5009960b966d2d117b6064a0e0be3489d58dd78f50
za8cc0011e8583e0984ac2e172558b5733705d3a7d5521f7b6954cf564e0bc28989bbe8a3a6c478
z9c26283bac5870c3cf1bcc4a070743e4ede93d0ef3d875059ec23980900ae3b0a3d06dcba37c23
zf8dc9d6f36f52ca76c2f7a36c1454831a2844aa5f02a544a57872b55b9425d6dd8e96f3e10e6b5
zf5234f190a8b9bdba8e3febe0480ba9cab2c47712e1ec0ab6831a19be827496eabef166faeeabc
z3a9f64c582d8c3fa27d5b5027b540ec40202456940f55856fb300b86ebc315421c797124e323ab
ze83ff35179f58bda9093965ebb3849855b6d1e49209be03e89cd22fd1bf3f185b6d26e62afdc4e
zdbbbf5a15f2250048226640b67a7ef64b62e560d1540e59d033fc8bdf51b55a007a2386cba4daa
z97b96132c6bbd3f972df379fce6beab9ba8b412ff7526daa6cee7e91702c74c757a64adc4fb85e
z3263b7060063bef10de8a56497cca51f74465fdc9c2f96895b022ce32c6d2fdd44811295ffd663
z45ca718136aa24c2baca49c8f3a1fe9f0977df8f8861358547e452ba06407524f673736e0de391
zb71e1b963ec22a48c2fcb83963b93b47dd79a51a3e4ae07677c5e1a3b6d4098369597416223ab0
z02bb7069489502c100ad3e58988c48212e247b65daeef3867c34e6ccb1e226698b6cfa9531bd96
z676473fda9d15382f4846afda7a48b82bb0a2ffa0fb4e9ccfcc0d1a02f3efc30e1bfb523ae589b
zb8192c2ce3bf9b52d857d1e01506527bae01c5d198e8fc28fb69c47a72444f7ce02eec0d77312b
z8d6af74456f61508421b4b1325c8d2cd912823f0f5e65777f0dec967cf2d526865d3ac3dfd3688
za8de15a102c293a71fab3c962acf0068174c73fd897f5dbdb821b37b68b0c3ff2c3e67be77ae74
z5cea856ee86787c2808880f7ec54987af797c542b8af9d0f3e62d7f242da3e9e03c8f32525fd55
za36c5f9f7034d802f3267e08b4d171e01daf4a020d3636924e78ebe711641409c1f3c8b581c77d
ze966b09677c84d518d72ae12c43e28f2d6f25c5aea4d0c405668a48be45eaa423225cb6050fafc
z8bfca0eff993ce0cce768dbe97dfeb3964eaff99de4ae7c12cd3673ff7883195008b766e383258
zad304c96dfd105a17659e1175dfbf1e979222c69644d518f60cec68727969e2d2fd87adaf331b6
z5c7632e4ba0fdcfce01946cab8900d58ae74e4576a567e36d7c5c1fee18f6726478a38d89ab33b
z1161bf14f1e3c039bb25e63dfc4457160d0831564fc47e1c383849eb083876a3fa0adff152cede
zad60e9e5837cf7a61cd1129f2f2bc78e9c5947891f9d3b732768f4d14684b33197939c010cb96e
z6fc55038deb29896877ab86dd0e95ac9f8217ceb9e0d1536af0bf8d70f2363e4c14e7e119f67b4
z82d73ad1fe0af96a206e4364abc63f8467ff5ce3788c6860a96c577b64671a862d34bb15a39c17
z91c6ee4daa77235aff5fd3f4f6c836fa2f2dc32a53d45050d9e44377a3c77f88c0fefa44844892
za81c8b06f6f957dc05dd158ae438622e527e76cfa00c5a21dc18f94bb1c7d0e2acdcca9cb8bea4
z7da23fdd11938c6913d24b5e6a4c5a6d4619c5e0fe202fa8f6f11a3550d504eb4e13c6b2e8de21
zbb7efd8b701b73ff3af1e9e00c2e31fd7de865c31cac448852586e0b63d59c526adc695a816563
z1ee946eb6a2c72c230ced3408e025f78b740ff6c6651ce857966b0ba9e1c81c3a952179a140cec
z38296e9d8028fc266e72e133fdfae7f909a292d83225fb621dfdb11792b4d2c80725097b941b43
ze0b5a5cef4c1eea41d97a277552f50b386e267eca1b415f6e7443b976bb3692b31cbb5da3c4298
z5a1b12cc5e2be2ed9a0e509d026446fcf1e1055214bd37492f786c62cb3a6b659d4b538b9f9225
z6b8af98fbeced3eb60f555edd9d6f049ac5483e8ac8555b21519fa9d46904719806f283873f3c3
z6c0152e1c46fb9d90beb79a49df3d62bd9d86f23426a14bfe71999a660715701cff464fe98b776
z912a0ec7cf2cfd006e6d17ecaf76a77e5cf75c8cf6f7f6e5b4eed5f862d00cc24b6d6a063ba3e3
z4a27c66dfe7756862caa72ea5324096a6acbc99a7db9a68c1e36dd888090cc91d1218ec423d6ad
z771630bfc3ee515b8d5a4cc5c1c7c017808817ec0a8c5f7ca6e2b13c9e7cd5e08a2ca22be18be8
z343185547f17b6d5cf9ad2f99896f41bd224a5f9001bdc80f7cd7b1515d20a89cfc8522108b2b2
z2bdd4ddd51b4f480aa9618e3844f273fd84cb0d763ab4f4bc77f7596a27063f545444221107c01
z219fae41995fa3a7698da81d7b7e271cd45d19cd8155e3bf964bfb2944433fd3acca4fbcc347e7
zc226336de45551514c3b87ef74a1b544529c8f36173bacc7284e3a7fccee015e112fb7c85c98fe
z79b70bf6304dd66f1f14d21ea2838fce62096e2cb1ec9b127cc029346637bce6acc887c666e921
zb39983f5ca4fb8fb149d6a1dea178e9b00a4bffab655a451061731dd8bfb49faa98951d65372f9
z3b713b53398d07cb109a198704f60564d5d8b01b361f72cc4f86362f808b4cc20a96745120ef41
zc3e80740c9197f6f1b4e50087f2da253cce8d251ca6e99fb581dd2cf319692e0f3dc7fe7842cac
zcbcab2b13a5cb3bcc0a1a904aa87171de5e459e67453bd535a43df57206a3d85c024a28b005617
z193a6cce23eb77347320a216a703133b8cd3fc456f082b5975d2d6cc3e6763684def8ba9cf13fc
zb9d47f8101fbb893b8872cd6cf2921d1d55c7f52acdff2c936b790c44ef8be6b592b9e06775b18
zefa614c6aca39ea30d404edc9ad369de2f282f2f1b3f8910c8437f1b9a1b84ca984ef92f1687b6
zc26951d8ed4c269ddd020fbb5bc278f8d7f88667b4e5397f9ed8792a4363e1dd8cfc93d68566f8
z829cdcf44a6d08fb3e15f878c892335cdf79753624e8994ab83b8cf8c9602012e9af3531f772ac
z7e21862227c27072c3ffe98b79b85922d895a81000f97c953ef1a37e1f8c7af966bdd64a605532
z81d27a42eb128c680e18423cfc2391008f581675261effc6af128ac2b6c30e10299ad69445a87d
z3f2d2bd70747f31074e6f4a1428ef88f47f412f06180e91d0c7e7fd4fe218ee8aee50e2ab628a9
z90af5d66494ddb62d46139d2993934dcb10b86dfcfcb7c69fe53b0f3478e390afbe240dc2e94f7
zf18ed9939ed6b37972cac7a21db7013986ac6c913d2adc4143d571cfb4731f2367a78995269ec4
zd823309f7a8faf116034c2471568e87cbc4f062cd6ace54ef2959e46db0f74e34c9970da2ffe08
zb8f10704920e98acdff24de10efcafe392a8063f6855e9635981bb6f6132f22c9644b1ab5b90a7
z01a58f53f5ddd44008dc42c44d3825d281606069f737410587b345300e35fa4f1a5b0ed2f5bc6a
z6b00eee6f81a11c12745bb8b5c4106f0c08e9d30d2f2164ed5cf40be2aeaaeddb379a03aef5071
zd47befa8b20675908151ecefc8a60af8acdb6d363b4b948102157034cb0f08cb1ab2b2ec8b4d48
z5dd4bab85fc514ea825398daec8e5d18412160c8760ff77b184f5ece8471296300dde3a5983ebf
za160472d7a4cb62918d9aac3c377ca951ce62039abaf4a3b8e42309d2982081fe39e191b78c225
zc3cc8abd0b3a348343418af62ff7c1ae2fdf5318deaad4df4c72400f5b41e20c39e8c1403d3a78
zbfb24fcdb794d60474fa699ee6a699eada5f0cbb306ee49f93348d3ec3c6994c04b57f36b202d3
zb6b84aaca0467d363591a9513882aea8cc32a80c5c03146521d656033206d8cca339fefbdcb788
z23a794c6cb61e3bc139243be23353c451c0d0b02a0cf71cc42f409374d0cbd27056aa88b13878c
z6329acbf7732af6c314db17be1c9fc4468133cf0d9289d531cdccac814185f1ebc9efde44dbb7f
z8fa564f064db8ffe9537e5e6f5e2c8dc5f555be7b7eeeb1dba909bb357c362701ac3cd8033133b
z78b72db1edb1b7e599a9d6480eda556e3987745c199e621932b6c3f8095128e8d574679960c317
z52f91d7c294aece0ac10dae435fa8cf5852eb63de5621c892d413b8978d577b3fdd393d83497ec
z8b4b483cd7d8c365183ad77c5a53fd55fa6f3bacbf7e9af576d1af5b73f63176072dc45ccfd59b
z9c636e481142739304b1b4a52a1b26f3e013bec4feab71d7d15053654362a1897c75c1820803f7
zcfc2279f8ef4f2c2073f3a161013bb41db5964379276191e75f3b3eb6bbd1b4d48162815d14483
z1bf5a13282b24dc342777997f6dd78f61b51d060807d7662f919564054ed4d18aea294eb6ea080
z4808893cf682ca4dbbfa3b20c64f971ac4b3357e1e0bc21e202ec48fb189cac3a1287a4933f974
z245881d076a9f9f3861a0282be02d17c06e66e29228607d938bb5997162be114ad549e67ee198c
z27ae80e72842d1bad2bab27c2e1c1bcfb58900b6434bb8d258cb6044df939ad1aee7c0f017fa3e
ze092428d43812dca921e0cc1c9a08d9e7dbf2bfb04e666c64aafa45f88d3f411a0cc090004db3a
z36336da6957b90d45bc8427580c0ddb5131adde015b268306350528887fd46f98e6349652c837f
z87c31f635583ef2c1a9c92ed767b26ed4d078c1378bc2c96612d36cfc8ae5d0f9fe52d33f42700
z8705b091161c1a8940ae63557d494a7dc000f3798d9c1ec3214237f3a9e8caae78eacfe5b8a9c5
z133456eaf1a98ff61b0f5a5ea7760d0a1f2cd14a49720faf2428b62c20a6e294aa82dc5956fbb8
z40223d29db06f657fcd6fdfd5fa8844c8b2c6875911f8875574e34344592374fd26822d5716d9d
z9ef161cc3546eb796e1abe7d44f8d68cba38ae9482c7628d2f50bfed3e8b6de101473c05606a2e
zcb24744370e6c065fc15664998ffb8f6b626ee30bfbf2203cccb8ffc0df5e6b92a42a5eb01d8f1
z6b549fdebf944d3a16b89474622016c7bd62df2d11215a7b981165ad4f30851516622dfc002e82
z5cce702edc01887bebcd7d4641a522c6d56da491a8df3e106c7393d405b000c323c47a8ba60e50
z647720322b443603bd27deadee577735e31a3e8d018e9e20433f0ec6c1d225dfb3e05831667749
z69e149bf8c405967b28b5a6fa324bf1aa240a33c66d98b3d6a4e3a57e0d3f3007e7628f9a1dbd2
z7c7127ef0007e1bc1b24d5b502ef7c9612d0fbd232ea60a60b73d1494a1e04a86dc8ad87c856d5
z558ed255e5c8fd80c83323b72d56d4361b073e283086b97f82071db055db4fcdf8f07afeede404
ze905eafadfc641eca437a50ac13c9b8f51c092cf70a3b202e58febf715d476625cac682031baa8
zda1966bb3708f562db103bf305efd5b0e5f9f214cacf5ec72fd885a46f90fcdcbdd4643f18d11a
zb9625a9fa1c195b668ef344a50fad03baee66fac46ed57b1e6aaebb4332aa13a44d8835662c3b4
z792782dd44add214c6d1aae4df61e90774fb8a6a9275e78bcbc75fd2447f03ce1ed4a73f75bbcf
zfd17a3bad6d5af6dc7546e83d9103ce68cfa84dbb68173ab00921c3e9f1e37549787e86551b900
z110f51270990b3a071a0332fc7230d9632248060830051e74d5fc1e708034983817c533f4aa1d9
zce6d536643fbc9916086abc1cdfeb24429555c4d83a5ddf8a6f52452812c25046e04ea2314dfe6
z0f55a3d7171a25d3da2f954b61cfc2e5b08e48a21e209fdb9c01612cc6ab70c25e8f1abc6f50b1
z8707132c25de92694b245e857689712befe97e1217a6ea98d3b0e67326c56482461dcfd649ccdb
zfe0d3b4f54df95ca44f44f09dc60f541d5d6ceb5ddbe9baf7e9b13748a3ffa52a9e1279134ba1d
za18080acacf077f9e384807c980ed17260f8fc28e2e232f80a26ca9c1ce6032005e5ce49c4a36b
za07f209db5fde4dc6b876bc3b6908a90e8373da476e01599e78502e2b1f209e2fa2c602ae2ffe2
z1364e003afaba0e4796d69c36dbfa8d9ac0d599415ce776f91fefb58118ee809a8b8068c2efc5c
z3d6e0a71a15ec12656795a8938c0ddbdd7c428e21979efcc02d68119035ab33deaaea1cee384b2
zc648f18ff7ac39955515b8796d2e76677dd010e2274a3004ea808dc3567bda544dfe2f8301b086
z481839126eb73103476224a417c86c8b7e7e202690c9cb877d01dcde6f3b59a3ba4dd4b0810218
z6757d166f89d1d5238005e605c09f904a3599342761a79174ae6f0f404ea17da6c6a37ed1a4fad
z48122fd8728239b1285a858827dfe751b5f3e5dc1aa2051517bb19046fc08c781337e91a3a704d
za07d7302aa3cb2ea54eaacc087f992f0de819d01ff86ed2c9a8f236c49512097d3c55f136a4bf6
z74199de5a10f7efa7b1a7d7c24edc7a180d6d8cd7c8bb51ca2e43f3738ea5f269a41f1bcda825d
zedbea64e06cdd829f0caa8382371ff5afd31e0c0dc9889ece4c3ce2cdd1fe881143556dc7c52f4
z45737368aae89ceef99c86cb8cfa69e4f2c955a2ec441303c4e1d758b401a23b0f9309ce7b4b80
zb01a27ea0ea3ba96cd8eaf41634d5a7e3160b17efb0381a353e6299789f0657abee6e97c610217
z784b079558b472d5693ada9b77c1ff1550338690f57443b4036c4a68d2f40c9636d965c5d5cd46
z18ab2572b110c63a1462cf3b44e53327bdccb1d9419096aca34a3a42c94372bc3366a40727b8db
z0cb46f3650df4a0db01cd634e549414e409a4dbc4f572de7474a232b000f3627f011a1508febeb
z428a85242278ae3f1afb5139afabb83cd40a708f5a9e627596cd1b0121bdc3da9861289be1d5a8
za99c78c158a4eff2c599c3f5c4ad1edbc64ad3564b9a8b5ec49344e1f1d71e41baaca248bbaa99
ze1e6c47671b7e09aae1b9c4666e1eb1de11edc4d2b057b4cd23b66d7cf608735d208fc75d62c1b
zef86b096b580af449ad663f0a1f82d7c05eb1537455014d504f9ec90b63aa3ec2df62331f36102
zb457393cec56ca9d30efdfca39945e4a34371402005006111941c6ee163fc28434594f5539eb73
z11985e9bf1e581cdaf5a3931e468abee7e1c8197bbcf714bdbc90e91c3f4b8a69ddbbd0456885c
z7a1fcc955afa797c114b97ba7d732df8d83fa6529931bda0948187e4d2518d73eaeab34efc6be5
zb463c3757da400c8907bd02fae43618c20945e13a67c00f3cc8a4a555dc8a8de530b6852b7f117
zd84f604c026070d57eb54917dbffe25ff0003e0a9e0fc1e389027c88ea94f95aa13d7d3085c772
zc69b2283b5fe885580919081960a44c97b89cb3db897a50a2f2e8c4554dd8519c8dde0daa396ec
zd7aacc80a19c2e1e41c231fd0581612a316de29a30f159f33c76a521d0e201eb1df30c37cbaf3d
z26c0ddf66a4565846651fffd1f39ee70ea3fd58b4ad065140f146e4d642617998adfb7448674d9
zaa3e4af02424aa5b78a83d9e36bbd9b48b96fe287dea8a8fa58011d7b0541c3c6ff52ebbaa1d82
z9b7714e389f7fcac180ceafe2b28fbde1c5c23b4dfe2c3a9224b98cab4bb6751fda3e9bf281dcc
zab703caf49463b2b53744b9918a2502db0dd49c31c34d0d9ce86fa96064bbb18fcad06bd5c4d0f
z68b8c7cac5d5440f1f084bd8c4a3c136f64846daccdafc87c3417b1c0213a8b41416c3c7c5af11
zaf77526def9c093464ed611bf6cb0a890b045ac5d5ee8bb778086addd3943a70cac2d93b384deb
z265c9f3f70b743eefd563e9a441ba29666a37ad283f5ab0d2eb64a2efaa1cdda1cf9b76ec06b16
z461e795cc7f6c7a719ce1b755611a422ee638ccf4ce1e2ef2e529c2dbfe17020d6cd92c2344a8d
z7324e7eebfb75047ea6a647e4913fafb9d421ab55e14c57ae4a5e150e51cd3d41e0f1469309deb
zd1a8a6272eb47e25e92b16f9adeab3deefb17cf269dd3b8281eff8bf94026d44414150e3819dbf
zbf5616d388d57d443913cc84a65b7b84052dd263276af3d096e9bf32d32cd377adc47dd2e2363e
z3b73fcdd188b8af44ec4da053fe317e4968398f986f0d0eab7a755be5388e89809dc736196997b
z1e9b2fb3d602d632a8bae8639d5e8b98b5f93fec81273f12fd873f9b2164c26fdb6b8b1f662934
z4ce0e5cb2e4df09326281ce3f37f5493aecf051e4750a3f8cac2bfd8f5d89fcb22a630aa9e2458
z0410121a4e77ef05668967146929e3d34cdaceab4b44f660ce3d1a8de8224f961018c5554b6e03
z780a9445800ebfdcf564a5a160f7e00f423074f15c71e208c495eb77536dc43d6ba606ce63aa83
z40e8b6dc850ea38cff9076cf4898568a2942256d4e002c5620dd87d00766a368511b76bbbf1086
zaf71d5d6450f2085d899592ab342c7cdbcf0e9fa2324e8c3d61b2ff329b5f8cc70b128883c03f6
z797e10abc42240b75b5e3719554c689564bffba2689e297990f6ceabbe5e05cb7181eeb2754d27
zd2f432b0b40c15089d220170ec2197e26263d5f765355bf729e5f08391497122e7994fa39f019a
zbf3a2d2e635ba1d8bce4636c0e72a2b71dae03f8170a1a688f005c673e39fc820e21deff485f1f
z9a60139742407dbda33227397e00f0ccba9fe43a1376045b915b10768d6400a9cb71ebaedd73a8
z587f07fd1aa09b8ac806112655af3b5410c807a78a83060afcddabd3161ad5beef3a4ff50064a1
zc4add2d27bc6e5f1df3133093a6b114ff8d179d3d11c2e9e354d142ca808c4d1f5e34ccf051a43
z1adc02daa2956191e5e330674ae63f6536cc3b2bed56d58ccf903a282759a58c708b9451aeebcd
zd89ec80a25d5d72938847e38cd1a117a9e692440c00cc1a342fe80f55bf5a48e2852eac397fdbb
z9e4921013c56ea9f8397c98f60f8281c66bf129d5e5a90f116f4f536d9c7e29ef5148c166ee3b1
z10e5cd0a8a76b9f62570d0c4a23a2aa7884fae7146515d2a86e2fceb2606d6fa3c5cd95f8f83f8
za4fcd9c75c845e8804da5a4b2a1ac942a5da0798c906066f981388b5529bee7b4920eb60f0012b
zb5b83ec289298d5e351a606f0e4d0717a9790f2c6d12e19969cc43013dce7117a80487e2acdc8e
za43a670ac2c909b5ff31a7a2bf93358d6424d92b7cc3c39b3dec8b94f35f659e978dc93302aa2c
zea9f7511ee65bc6159dde223db0906911fa5670d623055e61afa98893911f90ea6288be94bd9bd
z433c48a729de82612fc58d8e57a7f465353fd9839031d69f701b102d54d57b2bca2ea63cab97af
z3f997a30900c92293c417ec49bd774a5b7c86f68c29cf29198a64e36535fbfc3cc1ea490d98c1e
zb4d8541f9952229090639533c647ff087b2f5cc02052a3b1901d8957aaddb25536fb1778144ef7
z896efcdf5ea8dbca0c4644fe568ddb64a6d1467f85e1acd542d54afd0eff58a2fdbe9b3c6fb4a1
z9dd193cf7721a25df29060a08f4b1f243df049d9691ef53436381cbcbf377ef31d486d0395f02a
z70aea6e24a731d5f4dac3b3d4b78d550f1a463e6d4c2ab989df4329f8d91559fb92b22defc3af3
z44de70c2877cfeb28878979d5ea695e76a6cbf00c9dfa9cfad331b4939e1e31bcc1e89313eb359
za93c529b12fd734340077371cd545571bbdc77afcbc50ae579aafea0069d11c5fa42484b4b65f0
ze4a0dfce9710565167910d9932b94d8977c6371f876e5655c3978e08f995aa727091d5d87185fb
zeb9f8cc8f9412a9ec5596f8c74c70d17f78e4866853024597af6dfb55d646de2521c4b52c2fe17
zf1ed56d295770250d517ec30874dd84ab049959e3cd423bc2d686a4cc283bdc972efac31b2705c
zab975136c53aad31123d52b9140f3614b4e8c08a07b68e12bdcc635dfc062d716b919f82cbfb5d
z72055ae0cb84361bdb04408f67cade077720496e8663a0f114106dccc4cfd2593f0c4e9ec6b3a6
z5d211a42cb826e83de7836d24cf4ae14b3496e1098846e2b026ebc85c45a92d215eb44a8ee63d2
zecdbf11c44d39b48b789cd5e9eb4b8c04c31dac8b7e2324ccca9b49f115a598a7287f4b901affe
z506819a6ae13e385e10a2674abd0f9bf697e61b83b73cab7b00d2c427862341daff36b26483658
z835317dae6bf04f57495e6cf93013ebc99903835d133ddc33b0704e4718ef27658f3102db71b3e
z10a216ab16f9c7d1ee09e6ac886f3af48e17a9c8a99f133e73f3b1531742af18e83564eaa9fd2e
z7841293cf7f08ced4ac75e7d056ff1a522f125f3f714105c1aeff4d0d0ba361431ef512fb98ae7
z1402e0d4190a7fbab6af95471ebe6d4ea76cc019cf27f223c5ca79d9e839c7df063015b3f82fac
z0a32bc5d22216d36744035c46a474379756fcddcca4982f6e111446a50f07c6f4a311e158e5a7d
z54285e1921866ba39712851a9e5706835f3915464843f3fae81d929bcbe7233fd9edbedfc853a4
zf3913692d511f745e4a19acbf6dd9717286c75299051f49d3422b48ccc828c53f7ba09de03ff2c
z7e5d2e7f7fcc7a4057dc9d9ab806557578da116abf62e4505b2549c6a4b9a2f3cff13793f8e4b7
z3876250ed1976f2d231cd5adc5932873dfae2dff0757708ad717a3fbb70e7a733421c67f19b31a
z15d3b10b4042ee2ed4041ad98b78d6200a8e19d878ac7f5c1ab44997a3838722a17ca7e2ab894a
zabc7e177587314c0161a349017ebcbd06b0b89c571778436ed8ffb9e1683b3389e1c3e8befdd7f
z24cd18251c0c6cb745a051ae6674ea445833eabe6008d357c10aa88a72edebba04bb2e950e2cfa
z361dd4be57d0a43bbd734ab401a47a5847af35aa5bade8aa95c2fca270d3ce961404931f538b9c
z3f0e0f547543287e003fe5576aaf29742d9b3807a48131622a1ad48a012f714b6af216d8c69a91
zbe3e3a26798793e1f81c0d065b7fe0c98ab89f74a15eec8eb52eedd866be48f2f8ae1220b4f85b
z94737bfb94c7ba5afcfc59715d82c87e52d75e6be8c79978ca8aec38ce98826a64b9e56caae3e4
zc9390bf9a33922e5059d867d8f376ee2f6afee4ec252b5b35cc71174d34a9cd696805a99010429
zdf81e7d97541b449dba97f7f607fc7b403035f2d214c7ab6413cdfb7ce8bd797365a472e4b96d1
z7a45faec52ddd61aeac3e0210116446c1d1ef9413472ae0c09c5fb696a110949cb54fc22877027
z9cd1cc610db022ad440b0995f476513a4a8946bef856512298c7ef38ba7bb8216b8c19c0d6d664
z0b8d48d6c690e02154c326cecaf9461cb084e7f8c9a77a5f7fad69aa216f31c31f0fc665a2c630
z6ca7ff07cd5511dc5da87d4044a6ac4444809b845e3c5d5da054f957b5f3503e577fed61827ea6
zce72bfa402e76c479e6f5c4bda42541fc1f27f56ee2e885e7bd4dcd6620d3267b4005497425c25
z104d9530932cb3a44e824c39d5bd0f6589c2b3a0deb31ba3e77e83ebd866c03651407e83b31f8a
z0660344ef3dfc646972eb60013c3917dfcacc812b3cf42827aefc06e5ef5dff917437a187a4de9
z39893d11d7d9198fb246b8fe3b62eea2c13b03269493cfc91c8dc8de8ef02c87ff4b4ea0396fa6
z4ac1045bce4d50f53d973101e172b7a8e99ff3ee6061a808c08ace10bbcea1e1ff300c4a181d50
z8b26cb6b3acb1a0c4050140a30e24e56e681bee9319dbe8786cf3ca0edad9f99da5f6efd10971d
z7f7f1deb1876c6ca11cb4f0d91eb3f9f85f0175a0f5d8b61925c21b40128f3b290322b2211a29f
z5e57cb4a62f31deb526a56bdfeeb40e76eb83eb4b5c09d4055ae0122d044a9a806de64bf9f6aaa
zcd67055c797ddf095034c6945eb313113fda4fbe502c04c2d54d71db2e9bbe36b6c5fc944b5165
z33d180e0dff05a8d68a35bcce53c55f95c5e17b89783f7c84f95251c73c769be247a1c3c0322eb
z8703e0bee7c50e9fe7c0b2d5e92ab635c9530ecdb4dcbe8b605a63631d301d341221011a6a2881
z60058060a818d07b413b0d68e26226e9841688ccddd0bab68bea68764cdd11c6c38d705b54015b
zf1c683024f2f0e6e34ac52001b01e85f2f4f5bd1fd1c3658cb1663e2fec98026164388de61d1aa
z7e95c655242ea166977c6ac6aa8b88758248ebb7f5d6c6f8984820f5b5e0d5eabba5382488573c
z817ed9b1efdb244b6049eb74d60c64d6783f2b976ef89645b241181103eed0796ccc59d761e55b
z0afe9c009f3d3d839d1d938239336e0e3881a4e2b5fd857947069cf1f7f3574dadc27ca54e68c5
z36293733dd8a46eb9e6468f4695405ddbd0432c08419fec55e2d8fea44ee5176d9e350bbd29ae8
zd1202a9700f3174bd4802da05ea920eb04474bbe14536b8adae72c31b6f60d97366df20134f5d6
zf1295370cd5ca5c61df39d7529b46e813318c1787a2ad8cf45251bf60cc7c7abd5eef58a7f859f
z6c3b568faf9b0971ef01330d655c499a67831badbc14f7d07f46630e959095caae1f41d87d8a63
zea7705565294025367377479c57cb6b7b089292e1760b33ca455cb260629bbf39ed3d856d9d90c
z9051d94ddc53401f691a2b2a34e876931aa5075cb147723402a142c5c4b229225ebd24732cc310
z5dfbd4e31bbb1483d3292ff308ac4afa5201a492465278c3577d393dbfec87abe9877bcf0442c8
z8d5776f98feb3cfa242d3aa983797bed408b75fd7ec9b268635372c13c8b3ec26586ab8c99cfaa
z179dc846b628259cea4173013e0269963e5b9a7dd1e984584e7a34508e41ae5754dc440e3afc18
ze4f6b2f11585679dd4c3aeda282a44cf5c55637e67841376bcfe4df25eeb0a785d225105804d9f
z4003866c102dc64d6118d64faceabb34d6c00a8ed2b0ab8f80b0c49fd8e1c8cb0894f4d6bd12a3
z4f012ee5b8fb6abc702a13ec980dc385a6cf9df2e2cef8e71b46c9a021db90b1352b46540f4bc6
z1f4725e11b30388ad622247ff97f71529d6d9423950b0df0a63e8064348c725dc776188b9e7867
z3bfd6ea765459f549960deaff44710f2fba623ec4c2fbf30d5c76c2b78b9f7d891275a7c895e7c
z0b9a79cb2fefe99fe36566937a1a40c728a1a1d2b36e5edc52561bbc8af7146277fa8150a00dc9
z78daeaf6f7c8cb270007a56b0481af2271b3fc527d0710fc73d8d1264d8b1aa3d3fe03140d4ad8
z3d8e1c77484aba06b84c3c15ed24f901d6354f75549acc82a25d62e4e1b22529556d69b73e0b30
zf8380fb380ad442fed38a546b792ec692820e771e38f17fb883ab600b5ac8216d1d24bc433369e
zcaa3d4eb8bf6f78d98a52b09de6854b0809c9c84ffed0a8ef1aa5520966b0ffec29450b03454cc
z3bc33c4d3d31d593b2bfc8ca1209209c8de577540519269e95ef263079958eb8c5b137be4f92ef
zcef95e64860dd68882ea815e3db53c0be6d9acceb3f5b7c248bc0d85d46f915116a143e951c19c
z6ca2dc736b37782087ce87cc8b7f203766c1b69d2140ee606685a921bbfaf08e1a777a991d4171
zdc0f22b0c6bea207ca8d5a5dbb1e4c80c14f58e049dd8b955073a59399f8fb46cc664f41aa25bd
z0515a735ed6920408256e77cf2605857aa955829d6e76fa8ef5f113cdefbd735267dae0ac4390a
zd7a69eec7d7246fb61818e9598853ae08296d1fc5ae87d92100c5270abd00ad3fa1ed143fa7c51
zdfecfd6dbeb310efdc99f382bc071f2fc0326e8c6f1abfbf7c1e6c12506b9842167e91b7d166ca
z2f1ca4a8c0aa0f812338073979a20b9bc1cb5fb2e59c08258cd9c4acb168ffcf6dcd90e56230c7
z25e10868409531c7a115a1084707b9cb51460ff4c33e82a34db40d7cb786d65273c27322db5965
zafa948b6fa1555590d0ec1e64296cfb180782387699c40958d3b00ad27fe5de79bd13fa10d8e00
zbf028f678b99d6261cfb484c71422cc982252e36c280c1db74a925c03c934263d5e5502cdeea73
z191dd5ed2729cd1715892bc4e16ca0cc8619ea72d3ca6baecaec6521b23054f4c8a30ea3f5398c
z7eefabb642ea4f8f9447bceb9107841a74bb4604805f88a7086027ea32fb94ffcd020631c940cf
z06a39a61f52100e8613984b77770fb1d1238df2be12de402b8939cdd31a2baf40c6caa8cd014aa
z91a6162e1cc08789043f7e095ebc40842cdde454eec7b5f8606dd75a695124d7ff8c33609dc77f
z02b9526cbd789772e1963fff44df6cc8b6c6b28c33b7158686b57fd0cafb2eb78307bc7b15a3d4
z1227caea3f95646ea16598a261ede423ced387c337542952f0dd9f4031a0235325a6eea7d7f834
zcf4eab48909f09d726c4b30cc59f74682633fac10fe7d976e642f250ebf4618fdb2c4af9f124b2
zfdfc4d84edca9812a14a95b4047c4dfa68c774264d86e4ca46229075a68eea8ef554084f0221db
z4a5f3f99af824b434179f7ab11db45fe8789df09de5e6713f54af1b093c7be5a1d3dc7d63a9670
ze01f30d9d4232c80fdc97156cb3534105de0518b1e9667299d8890abcabd350585dd25b610b968
zd6f5eb63227599996b2523bc959afc1bd3e9f563de89dbabedc4dbffd8c2f2036a4fe22f9f59dd
z2da8c3b491d2b2f4a7f1b7f4b73f54df7f7227b5aee6b9ffea691a842dc4dbf3cc27aaa480791d
z7570643fe8f828f21081ef33aaea384102706e8476db812c220556ccdc877854c9c0b5498006f9
z27a956274c0117dad7796eb6ff7e9b6e9af02d5d9b46e679791915cdfc01048cd2271bc06a3194
zf96900b4398b97f06335b0ce0bf595c37bccaad5f9c66b7b417e43034446f793568f00b608ccf9
z9cc5a594a83d8f9a31d2272533fd58362972811f14900b0ca1ab4f823b8698c84ac0a2947a83b4
zcde18a269847d48d62143bab8950e2e2e4efc3b942394f549fc74111b304b1f62d67114486c0f7
zeffb57210fc3290738fbe7ca8ca34640d4da20f131b14c2c5c3f58cd8b094b1839ae3cd031b76f
zb5449f76d4bcf473ae08b563cd8d1ea18f1988f8794c454869f7d8a5ba21dcdc4250253dca544a
zb9c1a1d546dbcf73a72e14512cb5f17744994642a6aff6e35529cf1805ab8f7147431dfd69837e
z17360976759da46d6ac134327ff6a6124b8e44147c558e96c077c4c826666b6c156306c924f625
zfeecf27b829cf84a4c86501c4de93385f5ab0816673131bf9d3e1e166a272946ba8fd03d48ab9c
z3dd3d76d96c807c7bfe02c7cf9c8de1e73427e14eae9359c72f41ab4527a633207c63f55eb0b6b
z588e9a7728b5aa19ca0860031b929a808c1e4ee47b33c4bab952bdf3946dff9a9a2a2d58e880d4
z089aab46a84fba153adb282552cf49c5638f9656cb3c480639e7dff37fff6384c95250a9d4ec70
zc9a6cd74b525120b1e1cabfed188bb88081ed08a69e2a65fcfe1719b0a6f102d72ceaaedbeac5a
z0ed9916c73d4ffedd25f0680dba54663347610ba1e2657b6554117aacecbb9c4c42e30d54d978d
z9a0e76c7b05fa6edde4c3fea18fcca4815a073e3bbbea07ae6630a4440dac8c557efe5cb3946ce
zf91e31055a7d2089648b0e3790190a087fcc79969d5d7859d2015c2b4b4226aab910d334c68d7f
zf5ee42d9a2228b09e8648a02204d84aa2f7c0316e5e5fb66ef0a7f622dc3257b579b7d6b73f992
z7bbd15174046c0afccbfaf7ddc32d5278ca0b8e8e021453d99be008a33bd7bfc4416a3dd0fe2e8
z5e00b657abb885911f7cbf1061b529776af703a24fb0fa1b221d2d58579f52ca7babf9fde2c532
zf73aded8bf180ca2e46bc432083d4bb691155f2b277edc083e35250d52c370f5f4531af9dd5b89
z4b69fa7d7e499055554c1736a6a544c46c24de1422e33c537d26be1c1565fc29812f048616bf88
z5b386cbc173837d01d8fc6bf38c5b0bc3bcc21b5e3fddb95e1f975351aa4e50ef3df164c5bf5be
z412e4c8a4c29bd351bda21a2359b2c00f32f365795a03e5f17e67781bc7fcdde253f196f7c1b89
z7164b451bfda54e8d1c281c314352129b2f49a1acf31e7af813fa9909a91336da676a8886ecdef
z5bf06db8a0470b856d6464a035dac3248012b93373082ab06a7e319a1018920116e1638b277ff2
z1234d3f0a5bfcfa5180fc71b7efae3014ba99ae324931d12c485ee3685e4fc781b5469f3ddef4c
zfd0e927c35fbd67aa7033bc78fd84e46591eba3841f170a078a35145a510f0c933a1fbf3d8108f
z3c5bdb11784cb61b036fecfba7d5738929b983c24a5edebab466181ee893e78132251f57dc6c94
z60a3ad13c6f5633267fee2e403a94c9b3ca76fcdf4d1f20323f275966058a99c141fc4a1780ff9
z5d15af62a9ec9cce3aa55168b926d66d02269a81dae443ea448c7d11049d4903e8737a01c2e11a
z7a0df3b3a76c4ed5a2ffb2cf62b232f8be7fb2fec9d71cf63a73733d00560ca287153e6e6f9b9e
z9d1453f2e1c59ab49c05cbc5d67eeadedb6a5c7cbf7b2a865f8c704d1c690f368f341a1f6ae8a4
z5fddfbbf3195ced7b6452c6ed5729cb90a03c1003910d6dff9bc5a1b83d52da8242a56299496b6
z56f3369e7a1cb2a5a1eb363bad61dd03bd3fe97e171d8b170e961377d15bc80db6d3911d986845
zeb871f883a304cfeb5706689ff894fb56cab4d754bc3695c973dde35f0d314f8c9a61dbebce669
z8c00efed887eab4e5bc6786d6c45112a20d03f421f286009253e5bb11a4e139f875424b106d8fa
z3c64296d50969955362012ce17d24a56fc11ece9e933d43bf298c6c6213fe4992d04a632851fa7
ze3f8f701c561fc9ed7ea519a8475b8d5050f206637819f07f68cbf1aa867b6c2a71d1bcd32492e
z733d0d744fe48e5239d89a0f85b6084d7543bff97866b770b0b7aa40b744b95b39df992e26d5eb
z7d5153e361bd0a4285ec51a173f11ce20dfe12b2ff358d70e010355a30f6da01a3bdb59eb4feed
ze60d1ec1a6f96574ea1ff0bbd65aed93a331ce9b43ae67a8baafa157f88886ca494d5bef1a553e
z84a29f79be7ffcf1a800be9e44b14582a1d5d232f50458a86a71a6904a5f9925c675036f39d9e7
z8adb25e86eae5c4df6437e0cceac714545af3c2ae36adeaf85a021f98e59b62b396c8b1a43a28e
z646b4694578678d38b4f106e2dad489f75c1ef5dab83889b794b71454bd82f6d720112a387922f
zd41137d800e083020350fcc0ffdd139adfe34a97ba3ed105a40be3ed311364105fe85216fa88ac
z0581f9806d57ff7450d7e21996f86f54cc143971df368ab580a09dfba841ba5817f4630cf58193
zc4075112ed2fbd3efdce49e21bba72051fa116bd2bf301f3ea2d1b9131ef6014b424f2652ba816
z7d7bd091cc04a6fe1b0166468f654df3659055b1c3bc99bfd0dae9ad801287d5be6e16b286e2d1
zf0769ace1b173dfaf0bf8d533daf67c3af0f77fe9797fd718f8135fba7ac2063ed81ae848cf0ec
z531bc68afab2d070499e7a323682c525255cd30e9074cb81bbd210a16e8ec7604b9a8232b95d87
z5567140656d37c30ac36f6c8960fa7599d31530447b7d955e90cd78a5984b339a142fa0701628c
zaf4ddf96b3b1288e80316e3e68ba0bc0cb063c5851189a51b42db83fc173542b29aecab5064a4d
z4ef9450e00e6ea00bba205e54a2696bcd6c789ab83eeb43ef7a9723aa10ad3edf410a3e6075c8c
ze715572684c6653b4275ab728eefb1b2c5ffb086022f1eb12d07fe39c8a98838f977c5ce636a4a
z1b0741addfcef852393e6d74ae1f4f906be7fd81215e608458cdd4f9b633a8164bc063d2ee178e
z825d87d4d1b2572458fcbcf954176517776f85567e908463bf2f73fc62369c732783672d158779
z855bcff1c232b5e12052fa1e607f1eae4552889ac94f27e3440f65d522b43185518027afc9e6be
zcbb4f8a02827d6ee034bc57817322bb87dac81705ddcc5745e31dbdae237471ac0af7dfae81824
ze7a783ddfa6d7ec39cc99c1679c96842388b5f4b87577998272aca183f2237ea2693852caae406
zd754b291e5460e5a9112b5be71872b9f3d33e52588955bf23dcd4548a6a00a510243ec0627ac03
z32708411a5a79be388f4b983c45e0b326ac0055f0abe5347a92264d3e587f0cb377b244702e8c9
ze5a6a10ea2c7f6109ca2ba5dfe2d08d5da5f7556b117d49372496ac720311f3efcde9bbfccca0c
za3524041a697cbaa7fdf7fdc2d148462c5119a429badd2771aa843a19708a73ca75e124492eb5f
zef0c0b2aaa308acf516a537f880ed6ae0ae0c58e7f768b41fe47d37114bf762d254dc605175a06
zcfaea5e82aeba7a4bea810906d360041305238419757e64fdaa54491474b795654bcdd33dbbf66
zeef27883987f09de67dc80bccba1aff97099c88d4b953a15ea0c49c088afa33cdab8cc9a526b3d
zfab2a4412a3ed6f4cc71c2030e15a711dc07b2a8fc7d2425e6134b9bf274a4b52751d86beebc42
z7b958f4a8a5cf1f85c19c113c6f26d9fd389db61cadeef7dae63f25f3e91023f370f9ee9e7f1d8
z0f9b3cb4ba85009c3c51a91a20332f6479146a210d176fbdcf47b7a253e38a0524895c5c244934
z56b84ac43e46ae51c3f015a84d20c7f979f3a1f141214c1a41a27456c58a27433041665815dc94
z8f71f7323d9eebf1a9a613d8556cd4df42a3fde506d6a02faab69b4ef4ded6f25ec52021948d84
zf64bbcdb9436eb37fbc534b4df0b84e47bf9b2bf83404c3c82fcb9587fe6a81fcf06c2669265d9
zb6e464692555270f266c92fa7e351165474505e00bf7ff7f4f859faae6c56a781b9c08a908842d
z8a5d47fa19f258500f56b6ef88c4a4c6450c988912e08e9ac4e527f5fed63e10353e60f3de57ba
z4162e19628d277586b6a651cc0dbc6e1f5fae0e28b449e40c982930a2a6abcb31ffefcfe520881
z61065f10c6d61aca8abfeb5f27892c41087b0d2dbb67f2ff411990cffe600bb28d1d4bb09a14c4
zcfc94d247201c5b55aa6a681961cd71ce8ff7f215b6bfc636bca2b2dff1ad9c3abc5b38c548795
za6751b47cc6f6f37cfecb91cf860599a5134a741b958b7fe2819c33cce11cb1c1a0b45efeb1fa1
z741c8467d70a611b001426183e556f2ece37e9f32e236236952d31a2b6611235f5225d5cff5761
z8936616bad24a0ae52c0e863ad6e0f719a74bf1a771341427e88c265988f9fc460975518e0d38e
z699ff8c63b8101db5559cb4246b744b0ebe1119bb6263cc8a3ca417010bccc0266a617f3f3b8c2
zd6fdcaae92d40d5e2f5caf8bea8a529db2f40a153b38f7caebf186adf17719251539129a88808b
zae8de4becd0c5321162faed98c902f5c92bba7518157c7194539e6cc040253697ff66c2e3c5e95
z219fa9aa330601776b6a3fd2222ddab076d9f05beb057a6de8d2020b42c82bd478ca402bd1fee4
z214dd35fb5625a7ade7ac23aa5c82d0d4913a55538b6d6293ed6ca2e7f0100580e17d07144cb24
zdd15c855e5fa00c95e223c3ef06fd9621a5ab372bdef8d7b4ac7fa36599f704f5ec5b4776b32b3
z79935192736a349116a2cc299358dfc81801bd9bc785df42fa05cb9f987addf3c22f57bb8bbe93
zec2bd8d1cc819a8330d3be14303aa41c6097df42f4f1a56c52d65bc0f40c3d7936ac9424ce203e
z55d9921c563cb3120db7bfdd21ec1ed0379169553b9b7bbbd81709499d78a9d386eed1f991b296
zd8071954302abb002600ec5d04d114eb9e4ee477f986052094326fd03c1f25b145b4beb7c55e4b
zf5f1e83794774f1e8e9a83794d425b6331db450376869a550e8584eeed5a3e7506ba3171df23b1
ze4759c127a123d3def99fef4b41201c1f6146c20b22cc0a3110f6228bda46d745f4dc36df1c981
zf82018a381bc1443a3153efe9858e7efd3c07912a7131cec9c66d7091364c31edafabd2af3d890
z660b0883a121a68f14de6b177608c0292334b957da1ea9393a87f13aa3acc9f795e9dbdcb9f07f
z47a9a1ff991c9f0c34cda0cb434c5c86be1302c0d487b52335218c41fbb72c05e359442f66704b
ze6d4832ddece19222328d696453d8dd76ae761e4f769673ef700caf649f18da00c19393b44e461
zdf2e28430d0efb5bd7f14cad4590d65b2b31a005ff75e2a3419992d0f2c052f15fe1b0c848c86a
z372f8409a63336c264a6b7a56c7c759de39a6e91775f957a6de5c4d2dc3d2fee5ee71283c9bb0e
z43b22fb38adf9f73db18f575e5d6172a93ff68babcaa6263858b8a7c8b1cdf450e5fc3970de68e
z689501273b2378c68e4e2f089e99d961f78fb5d9803d322c67bf71b1a57532c33d6aeeff32479c
z4f7ce1773347b23cc5c7ce66ade7055372386194124b9c2ab9417c7dc0db9aa64344c1b89808bf
z901c0b351a663060b2dd6251cd7b19e6b263a4fcdb8a8571047a0adeb8dbb0ae24a4d6f718c302
z3f3f0e578960fef57aeecc64407fad8cffa9b45d40e4f25fbd71dcc6e4d1d9921365889b7dce81
zcdc8a8e555d2e87b8aab4cbd803580a39c149fc24f0ca7b8f1c1aa26ac2fa9ad5490326e2df388
z733b2522f2774fee8b4f473561f257f149f32ec50038b039147f757404f33053a3f228a6cf3af5
za0f354ffb43e99a81a9edf08b3972e4c80fa1fd9488a1927a9e488177940413877793c80fec138
z937ea70f8d75c4d50afde28333e76e211a6cad3ba78109b4671fa9970f919bd8760d65ff6763a9
ze81cd31d7d4ab8020b1ee792e512d5917c6407d2788a97c8673d876a5927d93c70f1841df4e415
z8a145fac97ba4825c49ba4f57d37ef6deda8a5b1705e1269f0d8ed9139964ceee5aba8c170c0b6
z0331551e694e3afe39afc01086f937892aeeb7d9cd9bad487909aac53ae05a809bfe80b390450d
z668caacf7eadf22d114ae10b5c33903bc998f9321a1592d11f2453610581b84bfc9e815c84e216
z69451ffd1da23c9d02394d454f26648dd4dad393237cab03ce7cd36331f46ee5f15f35fc8ee1f6
ze68da5f9c35eed55e319fd0f83f0dae26eba523adf60915570cf7fb03fa8d7fe58347eb91eb3a6
z0a84a58e80d9fd6eb26c1fd987f345b7cdfa6161fde754dccd996d2a58a9bd07a9803816719cb8
za77ee4b4028c33b8af75c3f2f4e5fae3580a3bef26cde756b9eb2472bd85c49dcd6a06c685611a
z85af01b6d3980a5bbbcc8fd54f1873777e138ef8032fec622562041a68da1f244f19074dec5458
z7eab1f43bf2f7c637359455d7675cd63c4bd725a3d14ec7893d05909cb470682b384d10914f222
z8e4086e377827fcb719c564078e6426d79557c7dd109c6dd9d769a828848b7b7db3305c029aaa7
z918353db3dc90e65149e71ebe62da98c7f61629c0cb87035c1d8309c2e11b748e7e753fb97cd4b
z1fe155aae7beb0d834ae885718608abf4dfa8e19afc8dcbbc8fa8d26be2693a74ff3815a9140f4
zc9b003f5a13bdec2efb8d285b4bb9f1fcfe11d73ed8ae49bdf29c768bea523bad548628d2117d8
z3001f90c3eae391270c5abacf2e6166324be15c54d6809e6a6507d37bf928b8957c22bfd832a41
zd19a1219ff9d8ffa3ac30738051e3aa81e00a95dfe430d2c571a3648d878a559d8718d703aaa7f
z30cdc0ffecf4c271c2effa32ac2a838d2e75b436d02bf3bf4f63a2e76f8a7e304612f10bc84017
zae82e1913c122e9eb17cd5e961545819587fafc73299c952de4432afc6650a652e12797e6d8d0f
zb06c31c0584a34ffaeda58e023f66805afa0c1693423d75b68bf73b8bd16d0451e9776a6f1d7c3
ze43dcee28acbadbc5d484372413389a3cbd0b5f2b52cb655d6fceef6df8918692df97981dda8af
z3570342025779cee4e55dabb83ffd1958d264d26ac696dfedcbf3cc4d5b1d941be3adca76c8701
zf4418da86341b720ae8514801edaa24434e1b50f5a0e3d1bbd24a975c49c71721224d7413e3832
z9cb76d01f9afef0211918584e4e04c969d328ace97047287f929f949fb192909ea44f0d656a35e
za36513e677b5dce78692cbe9dd8d1863e3e86713371d6055364b0d6a26e6175e669df70adf086a
z2a2de38329469f912d90eedf6ac314fb6cb923f0433acf0f565f1b6da07cb443ab3c5ea265120a
zdb3e8aad22b02a9c886f9de2ed9025cff540f0be4f6b2c4d8cb3bc723b4ab72e4abe91af6ad44e
z8041a33796e0d0df295c1b831f4d78557d0df9eb369a61f33ab46769f42503bb4d39bb9d16ae07
zbb94d7bfc886a41f68849a4c13953fa4f18ae9274feb129a06f22afdd08e312f6e48ed315eaf47
z082c9adeb994e275809706fce857c228deb720bdac1fdbabf0ebb79c6c305ac372085e390ec5ce
z5358832d5d7883599ae383477725f09aed1c8a4659dc24f8386a91c16402784fdca9884eccb2b3
zca80fd4d072c29cf2272f22cb4badebf87f8251a7929bf89bcd96b771f01ce6a2b96faf1b7f465
zc79bf6bdfea9c6d82633faf71c35287d96a22df4c20488e034f707760f9c5790e752e22b86b788
zf0e8260e3f38e8406cfc5924556d2118e42e65e222b79c7c8580ac34c5f48c6ba7e1bb8ef84119
z78b8060fa910ba56f2f2efb247eb3aa8cacdd00a14af0cf48265c215473b010c6c604e31004542
z273943f090bc15b49f8f6083eeda47e75af0540cd80fdf269569ad5d65edc45d82666d566d7574
z5b35edbeb39e6b828fa555749ea7ca2ae40b9a4fd8ff857763128f14c0fdbc49f211d972b1301c
z4f2ca69614a02ec5e16e6825bb0ec9c7693833493868844c3a0b7bd9ba58b67578b66e568ccfa2
zfb62394140b0f30feedf17ef461b23750a8490472b04c8440571c3d24e956c8c2d87c76f13534c
z749a6d80e89e9b18b660557ce3ea7abfc4c2a7c87373ad273f70cc2119025928c19a4a7f79894b
z2b6fa8c3623c7ebdb7b26a8b37cb99777c57a312287b238c75dac062a9c65ac3dd72c609ed2175
zed6ebfcb32dd1b7ceec69ea298b8ecc647985db30d237abcff801f6731d6a328cdce9082517130
z5f65852b237967864a4dd41c08128b8329ebef6978386afcd8619a4f4be98815e5b1a12477572f
z02f521ab6758bf8adf3f5cd2be28c371b39bd57f895cd26a752f7bbd2edf917370af9aea87d816
z95a091417cfa9174fce620a9365e653f621c186820551f2e4403ccfe1c60b01ea169b9795c0c11
z30c1e45dc04d20a2b18502e9149d7f62b998372f5620678c63c9efffdca737f93378b97768464c
z890f1c2350ccc46386e598bfaf711e1ff8ac5449edc1b6bd0886f91908224ccdfed34b84dcee9c
z766ef57936cd0108934852b28c6705af23158a00d79a5491991d644f3eaba7de3af8242b42378b
zcb9b14504bc56ce00dd654e2f17af97531cacc58af683a55a577bed6247f0d20cc074e0e6d266b
zd89e32e19f91bc01ed562b62092fc0b7f2b318b31b0655c9b803354edd83303af9534904beecc6
z668813e4bdd4862c91cc8bd6ad3f347c294b60e7708d1ff38ac1d48b3328ae854a2d22cc3daa3c
z160d8cf34116a76ff064291f6a6351abe7e37d968b03affc171378a7eb6b64504870763dae3456
zf5468c4b89f4190b182935ec725e3f24602b0024b8c731526aea3b6116540f07fa38832f96e7aa
z296c73030ac610f5e642e8fd6739ce020c6a9f78ddb608a61393ba436e12c73ad03f7799d3518d
z936d22a8adddf67dc328d087c7a1c9eeaf696eb0c5eaffda2bf2ff83ae85a15ca2fb2a2d08bfa0
z3119b259fcc24b422b4aa94ec9a39068de8e673e614a89e6dfb32fc0261066f701672c6b634ff0
z11403e3341fbd3af8d1dc54b01e649f51caabcfc12d46c42b5f4a2e9d5537ea687bbeb85d2dc41
z34b4fc4e1b4374081c4e1c2e036f12622f3c4cf5cc539de4a01f4389f07b13f0aecb6263c83148
zc256edd851e1d87f8507fe03e47340d93de963185745cb49ec122e19e8e9253f3ab63dfbed9de0
z075c8fe90b6cbdfef2fcb0ea20154577274b1c074c36a7a5adb36b4d5909bd48039e159cb773d0
zaea8e7a6b85d47fbfacc12368a9131beb1dafce7509421609f96b83de0e0c562d64c02eafd2dc8
z4902b2b4f4f5c8cec7690189dee987b72140e9cde3d849fcc5dfd7672cb13b89d6e25531220e51
z71931b6c0d42e5353ff4a903638f1cb820c88548ccbb1dd58a1dd86620b0384f07070f58cbe50a
zbdd1444ecd38f1cff881a063214d6d94faf729442bcedacea4b62b8d6b73dd2f6435b13c15af2f
z3fbeec46c0ed6ee18245cf765dde4996aff811fa2472a7697c29cfcabbea2d66303c15cdabccee
z66cb564eafb1899cfc19e5de4e4710cd4e1677654cb6f5b20b0b7f4a2437fb1a85b244ea1533af
z272347d85a78289001b8a5425d45f1825428563f239bb910924045592f5b70b8c3247f5d26a387
zdcae8dd844718fde49d2cb888101f4d095da080b9f0f4f94747d20ebca6d4a12c4d08c6dcd084a
zf18c28eef644857af139eadc7a9827e524d31452d793739cee9ea6e5308323d45e93d139ad9e97
z17006986c3813a2d218390dc8345d220347794d4a7415ea1c08bc3198936f1e6ae78077ee52756
z260b080d1a3196771db7bb323664643cc401ee76163dada8bddd2d94f0abe8feca8237aa7e1ee8
z96b342d3f1ca4a533dfb02f992ab7426879be8c23b771283e54441078b96fe014fdc58998286e0
z4351ea27a93201df6463e55014e25dffdd80854d718f434fbe852283fadae291a2cb10776548cd
z601f91ff43eba0fd6e447d3516252c93459e72f6d4b136eba1419aaef4a38a9ba889ec2d83cb57
z030505d9998dc8006851a744e224f8cd33a9f986e93f7f7f0fa9fa5f832abfbf83718283268afa
zc9e6d03878cadb1c1403f0e988ab56e0d902629fb3d9c7506b49b5877c7e48e2dafcc2d08edcb9
z4dea2017696cb4e2ce229a8fa9471a76351ae6fb2907253c5668c6029c5e62e5388daf167d9957
zd7b9165abd894fad4592ee01cf0f6ad3cee437082dfbcd1561951d032a71b526eec8806f9468c5
z85b493265e7d7d86fea7ea1a9e75b1c943209e0d93776dabe37ddbfcff7e287af977765f3a6cce
zfa73428d259eb0e31741bd46be973b116bc03d3be7481b42258ab0b341e5eec2188d11c4784199
zd940a81ee6d4c8b824bd81c5d2595f5de3c12828d0a2a940685b5aae12d7ced95546e229702ce8
zabb4acbb5ad7753e6bd8c3f17566fd0b145bd95cdc0701b25943595452ae5d08c2a043c2e811fa
za02221ec86d8daaf45fff40e175cab95bf16b6c078d7f6ac9d8d3c8b146573aa64256c3417ada8
zeaef736618698825e9a7786de90546eb9bb446f94c4df60582e7b87d896fc31548ef1f4f6a7265
ze21200185feb5b0d2cac4f76bfafa8731673670b18971eb381301a351f6ee6125e626f06347d29
z2421afff921f2763be99db9598cadac4153f21577f8a8d41fb91fc0592174e5d241524ca8d6bfa
z59723b383d44932dffb09e047a8f3c199f558c93f9cd81fc6013f030c56b9e633a26486a4117cc
z8733ce89af3012ffed554f2fe754bce7f68ac78b0f5854e13772da8bdf38877e47db34ed95a5d1
za02196b401cadbe450d3fa71b77d6a41d41a78592b9a556657e4859608931cc2b21acc76a2e710
z650c2bc1b7ee761d0d5ff9d3eb1bb91f578c4b7f99345265a5c9c7dfecad5960bb57cd19bad1a5
z55ec91b0d4ee4b8d4159df1fc4215c4fc9a456c425665d23c1df63694913254060e1e76bfd31a5
z9a9677a6d0e42c9d7b0fefa04e41f646cf045b4c6809e4791f949182e3f268dc308425342947b9
z886db16585a1f77389119ea2a04324b0c3019d3a5619eb7a6d93a6620f41096d6d6ac2d722f55f
z586998a05b806db41f28b0c3f650def469cba0fccbf1736c380bc8dfb72d150049848bc1aba600
z13f5044c50e8d08456a1998e1a849807e2f61d37ad0c88d0004c20bc737373b3113f97ed5c5cc5
zea0999b4acef7f7045d19b77d60f7bee15bcc5c46dc5610be46440dd425ac4aead3ff113d37505
ze00e0b4194e1e37dfe6126b2d005d64d315cdca87093688e78dec0f6a98e5a9e58deb4e2932a26
z83ed616394089d991c8bf871223fbf060af55cba85684f1cda22389e7a6c3c1d03569941eba4a8
z1e2f16d4d4f1bbee04417322fef3a18d53828dc479d196b1b18c6ed1254837217fa361a0b3f4dc
za3621a0cafbcd6465230054bd6a8d8e4da308646ab60633a5b26ad827691ceec2dd6fd3a26aa25
zf29d0cd9d5f27509d10ca9de03224bf1f2e12a63f90ccbcdb95fa5db6e63c8cb3ab1f82e91768a
zdc3f5f5494b379c372b71d3e46000d2434c4c3f5cf7829c09e0cc4e31bdb16aabdfa10b2ad13e1
z97d0fc08b57ea21ccbf34e53340effd48fa2366f366128917af66a0dcb5317d0c7c549178a6cdc
z00b92067b3e7080432b7180d5ad9343c362832f0a8a6606e8cb074dade189e9cad47fdbde83038
z8f0c0d4c657c76ef30420c7e4ab717f79fef9d30637209f024362eab9cd2bb2ff251cb87e10ec2
zd8b41b84a4af062157bb0931bfd4146a3806b2cf3c0002d22dbf7f4b30f89ad44b30a359aaf93f
z3cbac116dc3f744496ae4c598f4aff1df6685f0c1411cab9583bcc0c37212db87ec50e393da490
z20af915e637867bfe264cab4d4d7993a7c02d1a394ac54afdd20cbc132e2d5f28a6c5551954d4a
zd879422b05e8851ef095fd910998f5737d9e56a98d168332762794a40ea1815dd4431cba76081b
z2fbd31784766bbae7845115023303d9920a12486c905f914f68294da4414e4e731443e69ac8213
z32f71ff999c59277d2511fa3ace7a08f140742dc7ded53d97668d922db7d7e68751b6d6b8a5605
z71e8095f68ec815e7f2305378bd381be6b040aaa2e19ac20ff9f05cf8a40b6c6c1e8907c414178
z392d395c1aea556b4146ace33aa5c7ef9fce02aebfb98980ba846a1fdb1f428dae779dc38ec64b
z64364588f97e07c61158a2e11b67290ab7ec77c6d19058907ee526db1cdc28aa09712354b8d14d
zcd36ac7f3780abb8c2bd87746cc989f785e37b42a5229eae5cd82d72390e80a27ad482c19a6262
z4aaaf3295e7368611c4aa9c4ad43f8d35fe82072c521803921bbb21517146c3a70867a8085eb8f
zbd6d85c74e3b76f0a4cbcfa15ac036991d82b5e381dff0f4753a2345f4071ca7870086d1535236
za1ee238d6d96e51bae87e2ef514bd21390a9353959ae6428c1aaed7b2cccff15a6f23c9fab0f90
ze87ca045d8b40b3b0f601ebc25c46c605a39586cdfa783c5e694700af8664e9531a4a2c74dd6a1
za92f6eb87283d28a7c3719ca6d86867a2e7bf3894b108e4cb30b90f260050d804e7fe7d63ebd05
z86c7c5a913ac50d327df5825fb5649928b3fa3fcd282a52cc6de79fc93ababa6100eecacbf4bd1
z45bf879dd654845e49ba60d918919644efc4f5f7a137049f7d1118c6cba5f776ef721b554143d4
z25e82639731571458e01d98888b61721eec762c0cd6fb53d5e8c5345777ab6e0ac63adae032c28
z8f14f4cefc1b52da6a076a34cf5036f8eb23a5ab43c2988404f4dea2a662185313949e546b0d3b
zce1ebea3f6af95fcf179a2ee67c3ba4f1ce42bb293e10b5c070532de50dd30055a3e2ff820a185
z24fbe8595411372530d4e7825aa385784c1ceaef1851caf704e7f5006b5f132d9aa80f7a7df224
z07e779db3b6e314559058cf5cbf7ac87e8c29e47342ce9863d67e1ec418727178434533ce7c3ff
z578ac21bfec4e7685479c312d31328724934d395f1292ac5f244b7ba8793d800107a14d43373cc
z6d47e76e673762b161a3b8c162bca33785224b634a4b105ff880adddc8ba621046186151ab0391
zd68dbf74a7adef5d8569e656f01311d5bebc223285911bd4bcc01598bcbcf78bf22d8870462c9a
z862423e834be7f93428241071c972e8e03a3e8a74a56d26422be21867615854c8b344915e9c8ba
z6611a635749c3bc3628f66b9f2d246091166ee557ccc054ef2b18fab98c08ef51c2d059d069652
zcb03ca7125307d0606b234717a0ae7f13e7f00ef9db4b22da3845d86892e93036c5dc3acdb00a9
z4875c2c6ed9a0c31f41c603a13ceab2aa84beca0dedcd22e7d923087ea97e58e326e751428fcef
z9b7cc801f3858b5b493a64ff01f3e079afcf2650080dcc58f1bf1be1af5cbd7bd22ba04e24233e
zfeee32de6cb7bde28d601e3a51954a831452e66ce5f4adf5505354f7db4e2cfd67927c26a7c2e6
ze9799806b9c3156025612f1b45d9a10d9ef6f7b379769777bd19d078c8a0db5b7cfbbffa04398d
za1bf8540d8148ce9c4d955f3f206b1d8034cb2f3976a8ca188889d79408f0f4c0ce8e60cf539fd
zb1cbb45c1f6277aeec746d15224c816749e015090008ade807d4488b4775f905106009b56ac15b
zaa993541bdaeab3cbbcf833ace1c5e94b7ab892dc589d477d446c1c4e88fc4ded442a1cd711180
z0b438d2cbb6a3c55f8b6230dcc241aa02b8e701d88e334c5d79c62a3148c6707e8fa3caa4f3e88
ze237220adb61f0c7283f221b538b07e6b2a50fc0b7af1cc72f1744a501c5ba2a14681a0d100f38
z50201b3a41949270059ca128c6fceefa609e800682ecb52091d03d555d803c43e3ee76b0f25cce
zcb9a2ebf83c9b33e8f059f0413431a3c3621524b486c005ab9d3af9a349f3895668ef2b638651c
z5597a43bdc009e6e7e76d85f992c665ae759e34a946776be3b34cb74ff26593550b042659b64c5
z9700ee3fcb70d76672a4c8fb050f370b6bfa4df756dc01040b4e7959b684f91b39bd3c172d9925
zb8efb9af79c2744d9bb1337ec0799778b53337c9852ea1aa4724516f1c2c0e2f0bcc05f8fd31df
z53857e316ec45456a1808889266951cc0c1a6a76e076568ab7965e2459216dcc69571ea4d50d86
z0a7719a46140b3bf7b397901539700cfb5fa2dde246d1c44a31fe344cb179f152be30415a0f762
zf6fc4fc61bc69b0220ea410d48d56b99a7580d7c095cbf1a097bb184b03142190ac9c76be667cb
z3610923c1205b938c3e03f63e84cda697e5d961ca621db85f423f714c930d5551eff9009e673dd
zf5bf922dd2a5c6f05fe90a777cf95ad51830a0cbd9be1e8806d1d117d9cd157f6e094b53e861dc
z247b9c98195d9f6e1eed244cd142cdcdff583c98c3a01359cb6677ccdfa8c24e7d62597edc3b87
za8884abcec6ff2faa9f339b089fba433a1ad18357cd6d97fa04ed77a0223f7dee4f09d5489cc40
z8810b2b9596543e76cb5600a26206f7b63ed0d461acf6ec2bfe90c6c7c6e010e98a67a44b53fb4
zc7924a4be9bf5a098f499b2ea7d162c0fe8bf230a3d8c433553c1c10dec0626a285ca1b0ad8abc
z26986a1d06d214c8bbf91a4c17445c9d9ebefc6d08b6c8e813132c0f021f73937943fc2756a29e
z0911a736b29fd2d617cc65def4df096a327b85cb9e61e64a884484e29a712a0023225cb540fbca
zfb665b789f5abbff78469cee4439148306bb203906dda9ca8c9b6178ecd074d24cc2d5a7b858be
z2a1f803056ccee4b6c2dc8970188dee1257e3889291cba80479a26c1c6929288083c41bcb33f89
z38f377c04c5c67c9756f00629b5f03895a26a52d12fe69bb6a7f3d3220cbcf10750a02745c0e08
z734a38d32a6f3c35599bf433fde968d0f2a39638d4b0516ef83a00d01bb8bd36376d486b1d1ffe
zf70ca7bcac071afa87e10874b1456cd8862451f92333a1130ab66291de8f6110315aad04128927
za6e754dad55c19a82770661d090bbeb3dd0f2509c97c181015eadb0c3de1683e2f6bb30d5e2c2b
z548fd6e822f0ccff891237a9b7db61134d270794c4f2ca36c44e8f9454f2dc5fbd3fa89efee673
z38c7342f998f13b3a51b044cf7cf1d20d8f914281bf60b1dfb16f281faa47b55aa7bb686065056
z27d0b28c2096cd557554b6877866c49f993ff49ddbeefda597352c6f0d9840d1426ce9eb70eee1
z0558c9835a024d83704fb564cdbe79364298d1e3a86107dc8a95bd30f1ba0f38848a1237e8bd4f
z1c06817b768fed838d57ac20e863b5cb3c78d3c280275f0177e26fcea5f3490c60a6cad2f716ed
zc5be2543f4d8d5bb86732f904564d0879db749a5ba15034718537f3f8f9b2a380d450c652f69ac
zddfd3fd6d574cf2e0232fd3b3936eeadcdb5cf59e0463dee789cc127954d0b4163dd1093830e3e
zf7f144f85c54139119affef232c67167847b1c6ae2652da1cd3720acd391d39dae1ba42f09cff2
z862d5aaf1829beebefd4b5f35e6570fad21c052170c0168e741a80abb5c4e3800787747296c621
z7cfbaf8f62426de260f1377475b80f69aad0717672980450a8adab36ce60c48a3c6324827243a2
z635ec93649357cb26470205f9e33817b6cfe3036f06c45190e3384184982f5f15e24ec5a252286
za41bd27e0c7656d77e07eca25f492248dd5ee30140ffe39c3c2ac8c0923bec9961ce0c6baae5fb
z823490d10dca06ab25e044db2139fe9427c4b3211251b63a25ea76105e6d5f2133981267fd422d
za6783c99d8f233537c331453a1a128926a652e057b221ec583fb1048bdc46377acc76960e3204b
zb90daa51b69e083022281485cb7e3c6c46040b72a2244f6a654a5f66df5e858444ca6b2cd150cb
z4355717ea091da3da8546cb093399aece8a59c6988deb84308573bef023ee099c138a0d8677adf
z649337de8d2a7f655fcbff0c84c46c2a4670c87515e25a4f73b9eedc72fa8cd0db1c01d49b93b1
zdc032d02ece4ea3cb5418446ffc6b8d07227d62468f35ed4f5c4c0aadc84b24be1e9c7f4b751c6
z3fb7b52770b5a2454c2ea31743f008fbb6793f8452880b2f9c2bfcf8c336a1a75aac7baed80228
ze6a2dc35721a9f3f59ffcc91e351e6ce59e54a9456a3614a8784fe241094af47086bd0e7aebd2b
z9cda8bce0a0008d1757a3802d210bcb3ed4cfcb327e85a3d89f045a125143d12014f36fd14a6c7
zaec3d6123de4c2c31840a940b4afbd2d34d61043b877bf5c052ca9eb0c9a7db1af92786b273836
zc199690b18ea50b6f26d82d9e42645db2eef858ee8bb31b5f85e29a27b17963582038787c2833d
zf06e862a7b38e6800cdaca62e6e482586fee02b294f24b1b4af05f8d77b2eb6d7879b55f6fd0a8
z68ff9a31b6e466834b3bc34333c0c3b6ff8cd0539598e9c96e2ead95dc91b75e66046e552c8ce6
z844e35947aa308da0c0699f46f6d8075669726cc9af3491d1045c7ac9b3bbd232794cd77e57bc0
z79a46ede7f017b4f7e0950a9053a0e18ea7216ac80895d5f595820daac75964643d2955c52b2dd
z4d07fb1590d111ec9765ed19b93d817a619c213d24077bdaf505ce2754e1d601ecebdb5552ab70
za7e4a1391aa731454e670618a70da42caf531d81e7621030791dbc0f1e4aa5dfed6b21c4198b07
z551f7e859d1d0db00b11b9ede8e1f2cfca474be6bbe339243cd028acf2988288b1250e6c131e0a
z7fe720bd087ac6662399dcc670f98ecc5931a7b37b499234468e63306d36eebe08b8ef432ff364
z85b183dab886f28a85098289b35aaf426bc0db5239b0cfb5ae63267197e78aed10c4e434dd2960
z82366a58f9fc2822cfc17b9873c6186336a3eb895b22b822d6e53caa315a94c5aa242eb60f2fa1
zffb51c511e052dd3ae81e7447286df085a806b42d315bbec7d5d10f731fd49e3013c8632b46ea9
z1f50b7e02c61744c69a41edbd537276bd62f764cc84325afa2658dc79ccfe0f044a494d3317057
z823b6e7b0f63609c7443e3708085caf25b830a200306194598d7d79561705105fa51082c9c87d7
z19ef500eed4b4db42b61b8f41eb86bc595d4f93a87f01ae931ea97e8e9f71866d7639590a3a2c5
z4a3b2696e386fd9fbbf5b676cd45767e99232a7d0d74828ab9f301d6c79d27087a88009866a9b8
z652f1e61998370bb41ccf5deac0717afbf524913a4ebdb300995ca27328663cefb8eb4c46e6e0d
zddf54fd0024fb30185fc3e482ef23b26e3ab9194d88ce5db9b2f6ef3cd7af8789eacf320f208a2
z78172408cbc22d079ec38766c7172a0d231456fbe5ccbadebf55b1f31e3299c5dc269c6a82b0f4
z2a0c2a561f97c34f5ff3b43f45ea28e85ebc7aacc51b82ffe319043bc8a6d12d3e91dd6e7db310
zbf1202e9d5d2e3174cb318c3ab96e5995c956df769df61df447bc78685d0a5836685a9ae4f6b2d
zbfb08e892d3b6883e53081a5ac0a8330de504855959802c67560a06d6df823459c684aebec62c5
zb964f3d374d32109e519b3f5a5e2a8962491c7adbf3121c08c2ef2aae61fff0496bada62cb7710
z52ce7e5158d260107f2d7f41411d98f2f514815dc18005191cc6fcd7b872d3fab2e0897295733b
z0092f421c884092bc3edc774b3c38bdc4b2eee411d52fc0377bab56f5a81ccdcbf56361e9d39a9
za152b78269617e7db197155045b2a253223dac01545486390c80065e1782c2ebebdef7b5bdb026
z1d88402714e43362ceafb26c6ad3803e68f19bed64883c56ddace9feeb475fdbc095256065be45
ze409be06aa2117fd4da921c6bc9f2d9842976553548e1a72f1d5cbd5f0a4c1cc402f3d6c539dc1
z485029763cb3496db04047154204970ac3b88528c6a9069df0552c9b95cd7823339c5919503d20
zbe130d8f8fec5ef57dd84b6f3e5686c84779e3da27d81c431c0d6565bec960bbe44dd405f74dd2
z82cc10bb52ebd60f0ed8c02f7dc49fed59158a11a90079f983bd4484d34f12ca07e3b367f3f176
z0715c08011cb287b673f54b4f7d2ea121e7dae3ac3695dc0e55e413b8c51c8b35405218ed55e77
zf04ae7fe4543940694576bfa9a70b553e7fc9d17dd5e0d033ce0d4b58c4d0163870db25a6406c0
zcbaa10bc808a61385ebf70e8933446cb40a630c3a637a9f7a631cf73d01906bfe2643f0f4081eb
z26bd23b5385ff216750498e1dc662fc70322d9088890c73ff87b93a33e8d8a589d6f20dbcd0a42
zc60ee59c8a00402216fe8e5e2d914276bded4191ba42b35efdf6ae40baf16491f64bb181697088
z79c26ffb36a88cca82894d0b2eab3ca3851a0f769bc63c81593ab02471d48707552f2d2f047f8b
z27224ef8841337aa287c36203b5deff2c54466a2287caa7eaab85246b76b02a8e90c0d94e9cd65
zabd5ff147362c3f8ccf85534bb7b949cdcdb9cfe4892034436582a7933f2497216f89752114ca4
zb6c4a5fee766bd9bd30ff55770edd9aded910a0eb209c6294a53b4af1b2a2af69ea1b83e8fa94a
zd83d9d75f3b3cacdc845c89415953e0148ba2475f7c65b7127981e73160efe0ac22abeb153c7c0
z91ab82108b5b6a014d5c4d1e7954e9cd030bd6815bc2c49f3309277bc3030887ee176014304447
z1118c62a3e9fd4ea66ebe457bcf102f7366e975fde115ea882ed23b008c9a9a00a56e9c00c7e5e
zcec3296ae9c42387929ae4b398ab29ecdbf2cb88e6e41f8e46e4ff039c0efe01de0c2d3b507911
z5c26860ef55f0be3730a24151baa8cedccab15879f4b293872b1629be6bce52a31775a3ef47f87
z52837be235b22f787c76c48758a06f74e772f19ed6ee7e267111251231bd9e11df72702c63acd6
z9c5d9d26beaa0fe363f5f4ad5624042f86d75e0aac5c62da8e0b320262a6c70336d04569182a6d
zeed3674b9c171b0e59bc656363a0ba0cb6e3e59246e52782dd3a05e7285e1328e2cb398d561a3a
z6bf3d64ddaf0fe8c03e1001b816662ed3c28b015eea2b300efdd3f4924ea8877614331c353a772
z285dd8d2a428ec8143d908ca4e0054775649f03d7c5c7e22220a09260e22d07560f315f2304642
ze5c3a373af35e4db35e343265d3e704b4b24406a619faaa0bffa1cf0a6a5c55c862790a2776dd0
z61fe87969f40d4c4effb355f3e6d8186ae275dead05dee3cda57124167f1b07cebaf81ce1fd44f
z9226d890fe25ea8fbf7a8d388876f0f06eeeb2d6869c32a36511113946faf56e683aeee5a743a0
z9112fcb7634ff0ace75c99f3102cce1df09a40a3b43ffd0dc8a6ea0c6455a637e4c342637222af
zecf6ec3985a529de2a0c72a5c2f8d7f792bcb1a25d6dec933c03ac5c0169fe15a552559591c653
zc03f52026d6ee3e7b88de781acd249cda4c248d002076310383a88050cde83df9aa5059378d9a0
z911f18965775a0506be13ab0fd16cfeb661ea01875f39510450c38dd38c90cf970de5c1d5d8078
z7862d35b413876e2bc692bbb3301ee1996b2daf851c55d98edd4874f9ed06fe792392313c25e7a
z3bb1feeef6c5146f50d0082024847ce9c826d7edaf4501422b0f09ad5de26f3c1ad0276944b73c
z4c254381ad8a581980bdcd0aef81de91fa8c7c81db13b6ba419b75fe5f453dd5a3001f7fe5403c
ze89c2ce39e74eb529930a237cc2eaac09e64ecd14b472e3a2f298570cb8dca27e66ede900ac1a6
z9eef3c0bb5416830dd3e50ece1230a4fd84e3e067ec5dea607a6b7dba427b945119c6fd667e787
z61d3156dd922f54bd1c8ce7e2dd15d2360112c783c9a11075b8f5b94f4684fd3232a0849989f24
zd8821761465057ce74d9002ba0c06859f40969ded1f128f188ebf83072cfaac7ec1d69e233c7cb
z77eb62d0ac06cc380817a8e4f1d99ec14be375d20063471fe4a3fb27098a3fcd3c0391cf59b80d
z5fea933c3b60b9bab47e09a675394e985fa6515cccaeff5011dd8b621dcc9a9abe2d911832a319
z3ef82147e234268c13585d096ff480410c440181f27ad6a7d76b09e18c46e7ab89957251eda76a
z31790208cd9866ac958171d450eeba06dabc59ddf4bbf77d49706c821266a298fc0fa3bfd0fc0d
ze5910b23d98ef613fe0843be2c218ffbb719474e1efc2cf91ab960f2b6599b00ef3bdad6a02748
z6af3ac25a8e3d0b7e84b155a21809665ad860ea1a90f4348c81b674c0f96934d9ad119acf21ea2
zbe3cc405fdb54e7fda207207c7e3ce80d9011174a784904d03413c6f28af84b9c1951565ee138b
z496d0626e851d2fdd3cfa61e183b47b77e0b5d6610ed0d1a1930122f189a9caabbb228ceb8f090
z3b9b177472e4cc6e67518d39dc7d807f2a9da9f1972bed8d099bba7eca29e5e1fe8191930f74e4
z2af61cbb02fd2ccaf60ad7b24299a16cc73d2de771fd1aeabb5db7f06645dc5b67dd344a0a8e53
zb0ba8c826d2d676ed2066f88a37d9124601e278c3b3b0444cf4ca88b8346c8b98ef2afdbbf7e4f
z5daabfccd180517ff9ae8430623afec1276c8039e8d77a3f3d5746bb44ad577e4edeebd59bc4c0
z605ca40f23e0675b8075be7fff0cb79c93208a0d2bc6b422f87887139a6caa2e8f02533a649a20
z2c766c49595656a2e1f577ffbcf6b330ef7e16b9c0736a73543bed120ae3ad5bd30636fb190543
z2aacc2be424adbc8c5c419dc10d245f38c5e603970b0b8d36c96fae290960906d19371c49c783c
z66031ec8f40ed5857637709167a0718fa55c5c4d5be4639e1a53a58e29cc773cbb5b0fde5ba7c0
z8289b09105e6b2140730319e529ad3bc206e4482cd71752c7ea0caea4dd8ca5ffdd3b2b96932b4
z66e9178a18aa13d456768b86fbfcf918aeb5176c0b730df9424f1a97a3bd96350113f8c51a0fe7
z6e090f06390b882b7c98c0039c871b0d6a03c36ac6743ca42819c12635c7b054e9a482fd691a1f
z160ea68a121a2c9480438a669c3c9bb2cda26cf5523f50a3dc891622d1be542d0ad400a51766f3
z075fef9ba7a47a6467d2d015c8a01ca405dd8d30e04e6947561e323d418cbbdf8154a2611a35ea
zb2ec0c2d12d8f2dcc4f82a3fd7638c1ad33e9eff834cd89e7ff903e01526ed7640d8cc9500a7a6
z4bfee89712b490696e15ef2c02b2d054373e429d09037111dc8beb6711530f4dc2c941fa0c1408
z46a699bf45dc346a5105cff04cc4b566fdd32667eb49b0ec1502310adfa6d8d4afec4710f9be3e
z969b8ca535aad0e444188819f4640fb9da1f2cd7bb820ae9c8c0926a5d4126137f984e99ed70db
z316b49e7d129d650d8a35f73faf1bff732d0ab076966c68652e87af754a9022238869873425224
zac4d6f8a10fe5a6d5b136eae6d074dead9a8876258a2119c296b33f7374021a30f964ed504e36d
zd81b88b9a0e5f497f89682d6869a1c898dcce7bcde481974d4320b9cc3f3c653825d528ee013d2
z406084692a18cf484e85f6fdc16924490ef174671a52aa0392a9dc2b1f3716503f379789f8c1a6
z6d8b0cc48a3a3abfd33b898a6697519050be21f7d92e56df1da6b5d100a62e17ef047a37d6db99
zf71674221c333c36e4965ad1df34429d35de458bfa98590c47bf3336e91da4cdce8d906b19d5ac
zbc531f51e06dd838e681ee261216ceb71fbcc34954acd23f8dda10c3ef063f191fd3f896dbfe6e
z4af9c27fa5ce0c0de630afa3ac619065b97f7888294c3ef0106572d8b23e1c944d41d28bf7c26a
z2b6d2e64f5152527b1acb6a35884c2f907dcaf45e8e315b4021ad547a2bae33cbfc0c6b27cfb0c
za81784ae09366ca04daa74cf024d26feb2819c3de606b76efe17e74e963dd228856b0d8f40d41e
z544793de467d350d1d4a64cd1a0397a7500ae6be3326cb6eaf7688ea778cc0571b2fb2d09d3f71
z712421ec8716b1ec9926754049f0b1317faa627bee627e037439d0b8a66b43848821a19e0de5fb
z32420e1d4e4e2f72b0aac5f667fc3018343f0920541e2f34ada9326037a7331aa15058b83b52f5
z52258a305cde1aebd116385a020c31550d196056a6d308d8512b68b8fd286a6f22851b66ad4b27
z298020920614482f3bb92e0e7d172d99622651ff7b57a65f3acb8a99c35f6752e2bfc6f444e2b1
z3568dc9386c6abea3fb3c823fa3bf2b18a5e2bbe7618682dfa96dc27920d65528bda5e27e7a869
z0c7a3c242d9e314df87f40dca134b49eed270fe7b142580b6138380757c3abb6f674f0d8d94efb
za06e8634edc55f74f5500df38fa275ff8bf6f7595dc319296343d02497f753d36f91a293ef9370
zdea99b812af88d8177454a4b4a6d41ef059b5cc329299c02a30f8e5f08a9ce6e47764a3b013e6d
zdfb04ec9310a6ef1bc1d5a58525e756096f63fd95c9bbdc70169086fc1e0c927975a83b001476a
z23f8ef59d06ef38b1f949eb40dbe3f313d8b91a1d7daa80dcc74c0c385e593fbbf1697b488aa71
z82807c562e5364faf69a8a91add5ac20efee89103d453c2db580a5f9c0dabefe1775e34c72941d
z15a23d30aefbe0d8b44ab4c302af985b838577dd43c50f2122cbb7ac436cf3c966888a87741214
z9e4ada461dada278a2f0a8072eead26b768b2ff3fd4be5f364e31d6aaa05c40a0260b7387a6e3d
z1656717474956ef587a55d1d181a41cf8e159a5122d5ed9646fab26e25a7251f92dbe86a47e7d7
z9ad3232eecabab73cf9dec3938f527a41783f3d8d71ee1506a00c08a17fb262da3eea6718aeca0
z58b50155b4cf2bad85541ff657e8ce39f47ee96ba447edf7daabe220041965fbce76f492e008d0
zfd8803b6be9c2870f772233542082f9c378cb787583c927c4ca37e85902c63c255378767011f3e
z188af13484f90019b259a5a0bb8921126243e6df87f1f6535d3f3fb118770d63b02a157a61efb0
z5dd5c6e3682c28bbc0422fd8ca9de53a02d71243e999800fdc2c3a7409fb032c176e883e29eb3d
zfe37082e862ef583b7333800248a41e1cbb8fc25c1e3555c96e05654649c47d51cacb709711ba5
z9aa1ae524a5cb3edfa32fdb7e6a350cf321036cfb50a30b3bdd5e889dec0c81a5e8c930b1a2499
zef269dd2699fac4b641448aa8f6e1e98a634164e7a0548328714f427ce7837381a54387866572d
z29dcfa2ea7f3716fa57bb80202d9260746a4bab95488ec8e6c0d8b820d93d784102ea44817c9d0
z811d07aaf22769099fd24a6afbfc039e253e537b7740da8ec204f39cb80ba5aa83e3b8bb61563d
zb22db8df759bf7f883aaccac8bd64fdd9fb0f332774eedbc87e2d1833645cdbcaf154c61821eca
zde03ac59b8c5e9d28547f1d414adf55fd395694cc0417c9ebec381d9a2bc5b028a53d3b8dc8444
z2ddef92329fa9dbdcd9bee12dd4093869e89daafc2e109c9121673548eb4f4839599c15d205a74
z2aff81732820f0b612d314eca9151de0fff76b5a0759cbd29c913289edf9e7920e77e2f3387e1b
z1629a70ad12ccef732debc822f2235d5afdff7b5be9a11b646c0a932ed9ec882ab9b7c554e6a2d
z8668d7673bcc3331e67d1acc70a174647dfa470ced7d97ea3c51ab0a6d5fbd4a81045c329aada6
z9fd16bf15e4dd6799fac3ce85285ad2e036ae4e80c14c140a4d04a72a50896d56b472292fa882a
z95c2250466f9a94aba56a7ac3c5457b64e1fe95665892a0b2cda23b01cdda5e6b7427dd93b031e
z0e8d9a7d41dd8abc957f62def4ba27399aac1cd2c3ef01df43e664e14faf725ba17ecee0e87376
z6e45dc28373c7584d5b5500d3676bb84bdeee5cca365199bd8749e9f3d2d0fd5fb15e512e38f74
ze617b5991d1b18b0d8bd6e12bed3a6b5167dce3297532d33db72cc4004f2e5ae8f33a4f4f21d6d
z696418616aef894d3194455b63e5435bedd8340dc7478a450683ab63cfa9f0bcb105df12a08f0c
zf964dc425cd8aa0aadf372aac498f6d04955a1a1f3a94ad4093c53b8a0c0dd7b4b32b47e328cc5
zde661b5d83dbc7da6891ddff9e62b02d19a6d938476827e021e0547d70e0a8f5aefff0107d3610
zf9861cd9f3710d79e06fcb969494c6d0bb2eaf7e722ceea5f28e7879bf951f48a2045c64b5eb18
zd218d7a8447f445ed3b7383b04e4062a668809ba65c9f658224e15315199687493b0d20e1c2599
z0b9a57b47cf0e16d9a34189bcc13ba8d299aba3b8be6d01f3354f8c45184b68a385ae0956d9b54
z2e431592b2550b0cfdee7835da9b272b89dc4bf2e75c453422e421bd0ce93e1c7c578fc21b1127
z3a78b28ffd2ca35429e9e8dc05a8d3fc5a25bbd023abd7a434a72baa15ea2bdc1d0b0c822953bd
z45f27dc7bef7db26bd42597c30021e74ffd8de2b6be64a0379e370c0a0867ec386074e16b6b914
z152f630de06aa0ae810dc9ff371cc888702385196dba4fd90e217bf25821af2544253a7f507c42
z3efb08497b322cc93313693adb78fb41808712479239192112d01c80187a70052e390d6c39f94b
zcef9b3805d588ca42f182a3659e5425f8d9bb902d3b1d27b3dd4748792f63464b868e70a4aa35b
zf7d0f3fb11762cb2311a8902dd1e433cf7f2a365eaf87e29dc87cb15627a588c1bd9ad545847e9
za88ed7e594980deaa733a09e80f6085f8553f9489b7a4e67f6941bf2285294576f78118608da9c
z67dc2bfe1bb052964a4839d6b8e191e8576acd2bf5336e8a3653ef37453418afd4b9ceee13a993
z2c70e386475b2fad8a024a6aa7308ca7a2af5cddb15348492eddfd6afa57a7ad94c8ab1e7ba3df
zaa1366708ed0d48e823695bc4bf83121c0c028ef6560ff10f0ec07ea2d4ed616c43521f5049cf4
z801825069db90608887aaa8d15f8db8a7b75f90b85aae8fe661f5002334a0497eb0820e1c7d397
z88422cbe132c06813b90a02189633ae5563e595298980ca6eba48da5165b9cffa086a79990f493
zbb0c614ff379b023299255362f3d47e9560c4fe9d6bba376a6f753421e90e3c8e925ad6cbd5756
zc3834fa656f1e8335f8af3617b9467d02fe1ba66c7d38849659a52d0013e4452e15f4648a0a492
z661a8c02422b73a51968c07ff0d11f773b129468aa74e45e84c514baba78fc8c1a39ba515c0e23
z369714e121f08e70bced4c3252ccfd3784689c89e4267d5ea539292f107babe9abb7dc795d1772
z84d9ca6b75ba8ebd6ce8740896ca8ce6e6c8cbb4decf03bb1e211f8bf5db2f098d1b61eefbedc3
z9f71fee1981fcc74177944600b4a8f5da48325835ef843760bea09fc03634ab3ca9687d68315e7
zbc4dcfc848d7682e9e427cb8f6153634c2f9254f372115eea6361942a8c3999c68aa6047b6eaa3
z97f379063d00220c13548554b45eac3e5f7d82b2eec15ff44ab8e6e4bb69129f05795efedc843a
z3b5ed450c9018a3b8099aa49ae4640dc656cdb55aaaad595e0193da1d5c31d6be5eab0ff0aafe6
z54fb31dbe9669e619a8571464e78911044958a2d497eba00e5721986b4a848bd565d46d314b320
za9b479fcf3e3898db1ff6240f1cc810a000af440f746d74286581081c7dbb9c79201dcf98d8049
z3c846794fae3f6e98381273a5fd130bb49fd0d98f7a801b8e137fd606f51cbdae9bee19eb994e4
zaba9a94f23dcdde25c0bb79bb56e80321b20bb59b59306357dca149f0461402ca858ed7c568b39
z4ad9e0f5d2c74a1f6dc4ff021265caebcf301ac9448dceb04f12f8fcfcd1953f60b74651ccb9eb
z45ef15077c2640bb156a6c36e0e053843117afcc310e83453ccd5678dc18f21d5fed4da52cac97
zae24b0dadf0237c48b737e5cade764223be99ede318eee32cb9ed515664f20340e85ffb0613708
ze5a7a657bc2104b13b267db95b22c2aed055f8ee6e15cd9f1b35538d0f7d391736a5f620a594f6
z0f72d0afcb655401fb532693f8a9b258f2d5643e703b4a26e54cb24ac5a55aed706e6ffb3466f3
z7271520018ef9513004e155ada8e3ca1e0eca7f018348bfc51111ca848a8961456fde0fc6e9364
z436649beaee895344ebc0c46f821131c99d2ffb067606147457fc1e3ca81a6757215647e28be40
z31fe339a9dc261f31cf37205573221095babe43a6a6bd0f11888776c105b631a0f64938a6a9e84
z14ec8b76e038735b4b07810ee8eaeed6666a3b2881de27aaea53f917eb327e7ab8574b9b38cd5d
za7d04baf007c35e19b95bb8c59b4648955bbc597e12aa5e9eb443948d181273afccc1567ca0930
zfb23e25d173223262ed49bf3e38fba433ec4f6a610d92abb8ac635a91b32b2bcffa21d4ccebd04
z3a1c2d2c464e0bf364913bc4db04e54600688c73bb96aef31feadf4ed6d73d180d696698e3a3c3
z2e18e6949fa38b88b9296e46844cc2804c3efc9f7e2f9cddaef4c11cdf708c115f3e4189cbede2
z2691d67826c45b78ebfe245f6b4eb0bd370d4ba735bf7a281abe661312b9810ef59dec5003f687
za6b5a338de34d6ad1de2488f5e1e1c2c5228987e5038f7ae35618ac9b581d1c3f9a2c4bb876a26
zabad906c41b0fa569829c459b5f2280cba7aaff4781c99e53aac64f74f3b41e58ce75cecab81ab
z9af4bcd0dfb188c2625d0dad38163882711ad478fad2dc0825fd8d1c25f71c55b4433a4b2e0bb4
zf4fe38a45b26ac07c481bb05f52b0103fa4d0b553b0187d4cd95623050eac9f5d758c28476dc98
z65f4ba39db80ae441649a1001e268427ecc4144cd0407b46f64560c4d07f54ca5bebe64f78a12c
zc3ca0adb9a7bdf1a790fd29cd10b410ecf6b85f39de06e3f3458754049018436568271e10f7161
zacea8717038e4f61d4ae7ec832e9a4fe71429cea3099e32508fb0c83b518a82fb1d3246bd24182
z6903aee76628a6cb6765b6ced813776ab31948ba367c070ae7441e6e28936759a7f4f653b013f4
z557e9bfe1a7a696f55e8d422657aaea3ed13cf8caaf60855c42631c0ad40c2e8a2b7b941c55255
z72ceeb8111ab1a66d3311e601d45d31026676c2e383e35dac89f603b874fa5189d06d25291e30a
z98f1711e3068cca12e97334e7a1735f3fd384e0472e4af677cd130a393d1f7ad8ed6933365b84d
z19f1550ce293115f6312a436556f785e4412c6495443f4a4bf5b48d060b7cb2de11464a890a86b
za19d1a6e6b0495f58744f4097f641563188801f9a399160e6ea032dcc719180afa8645e849ac1e
zc4e5cb4844ba1e558f4f1ce6f0aad16cdf9f4903f04abdeddadee75e1437c91e6c97e47858c40f
z2b17e774e6ecb77e8fcb2b97b220c26694e60d0841b95c7d2ce8af9761a284187cfddc5d08dd9d
zd7f18f11c04c6e91f761ec5bda6a32ffa0128e50b905768474f6235cdc293745202dbebcf4d053
zb83c318b853e67dea7e87bc1e2c2e9bab8235f1337e0da121f28e724e45dfb58266bc4ab26a4bc
zf5c885e979b4e0a6ed9569f3f0079de223517b39fcb6e42f9f0890383580b06b96d54c7af95139
z418270097e58ec87acd6bec8fed3d300f152d4b43aa10954df589b3c2094cf201ce4888bbe7a47
z34f5ac6a136f5c46ea1edc44c549d8cc728b2a1fa34fbb8093829402d9d162a4c0a1be5c78898c
zc1b287fe06cf67fa0416f6653a6d90edb16b48e500eb27a59a4aa6307eda09606f9b3dbf755aa4
zd93c3ed3bbf8f5317683a75499356608e46ce029d1e45daec10001926ca4c5ddb29f1265737971
z734072191a54f90c5c87abbea065714faf56f7b989999f4fcedc896b28433aa79b82b8e805e902
z4f8de8567f3dd15f286c8189aa4d0d5ae5560f16920bd50898642789a565efc804df7b6e72ec7e
z23b32db3c470685ee532105f9cdfec1d3a7c341288ee3f7d5139b53195be758716570639bc33b1
z2865e0cbcd0bed28ab279fac442f83456963381c7d627e6ecf83c9a129c190fe32c4ad010b2ba9
zb6c08fa586c125470d9e5b2e7f076c1ec3a4fa5a31d3c4d3a56c3c5cadc7c0e9c9df94387be5b2
z29eff83e6cb1b3764ed494b28d6cf7187fc2e23ebdec7c20ce55d999a6d71996c9ef52bb461d91
z29b7af576284be90f3754cd33546a9f1de300cdf0fffc0162ca552625836be2ed2685c7c19488d
zd03df65e20847a30beb8e780e9f492a6dbbd6f4c8be510607c4fe9c05af0f8dd45b5e2701246d8
z75dfa0e60ba6082126da38da0cb55c21d95a9d5fcbb685776177c978b6ee062d9800a6089894e8
za3534862f13f88b187914101bed03736be7d7e3ee298448d0694e58a6c7c9f612c85660d76fb95
z1f6fcb00bd5dcfb51648fd331f383db5d71ddab05fee7f840df48a2c48f3bfc4b6e680e0a9ffee
z1e75fd05a77fe0b0dbc23080680a08a49de9c576659a77e9d7338e8c7a95f312ff69ea74088e23
zfcd159e5f5b6344dfee34d4716279a4ca8fbb23098fa2072e478dd81672d7924c33fe167895701
zce3f93d17f432ad7b9011c328ab15ea0af1ec6150de994860b9652741526b9fbe3dedb1ebe294a
z0a2563b28010b3d30a4967588b3f58da0aaa7a25a28fcc918f454d781f749bedd5d6859388a62f
z7fb1689ded440035d08bd72670543b534a14a99bb3100378f63f66a52ed27bf65076c358959dc2
z581f1c5910f6ea9835e5590d439557c037d74043fd6d2081b9d54108902248234c05e7b74ca562
z38a17b72398dde030c539a1ba8871441db174eefd597d6e2aba02a3624350ca912e7e60f723bb6
z89d9274a934d8e22f4f0e1011d003b84b38efbf66a2c94ae84aa081b846194a0691752e02c7635
za93f023afe12c5825158a49f6a2f27ae5a0f5b0c53fea2ab91e02090abd18b664645e6e026cab2
z081ef64e3bb9c1496adb47031a486609f917cc3f4277e07a32b5272386c6e2dae83e8d7914250a
z2e4688333e481c2b095c4b255c522f05714bbb215830b7ef4eed01f292dce187fcd4fcb87c6a53
z8f49a109840fadeeee51912f7965b04d99525ded5f7a7e8b33cabbfa5e3c253632e552c89cf474
z7aed9ba5f77a3d4a11d16ae22861c2d82bb042d284e07290d28e00985953b1fad202e78b959278
z3ca6d31aa20fb7d8c857b98d97bf3a6ba7d6f02cab8e7a7712f3db5e918a559478bafa83916290
z3cc7dbcacb8143a2af43b3102beb2373cd87865a7b330fde4bde5f649559b19746a676ac6d0609
zc0c73ffb014ccd224ee749954687bf6baad4c07dfdaab21ee8cfa6e40b9a074bed35fdb0b99edb
z2ccfca9f81c9df23224f2dae7eb1aee7b402ff6c8df5efbe337582eca1c878683f20b6c4cc1f75
z1baa96be32f44c3201e757b8980e65dbb919a4ef4ad4bfa39fd30be3e928ba1b6bf23ef25c2567
zdfaa1a6b42012a02a25fd08651aff775b69c1af35ed67daf1fccbf3f12decfdd8f25e12e508ff3
z13821686c96f6c34e8387015e5d797494052f346f9c6f4eddf912c29fd98bc9d682081f20779ec
ze4935952c9c580f148a35af91b8208097fc9d7b76e074895a21bff5dd34535d4e4dc832e24b92d
zdba1a06a84dc37d5c8f5d51b603649ee2347e9fa0aa470fa35d3277842ecd39764fc0989aa3640
zc901e9a7509924574ba5b8d7e8e1d8b246ee6acd0c699df98debe62587b4fd5192354725956141
z246e92e28f0bb601197a8579dc78a9995727e6e0c30f78af2efd487203488ad2faa5d97b675761
zc925dd305241ce361f44a535c00a74f5176e8af2858ebc6df361bc57f31beb1457ddd48d074c6e
z01a9549f6d1aa0098d2bc7eb4d2483c912d5b69b5da2723f2a07e61e2b53c6ff39148e29d9fbb9
z08aeb713f6b4ccf2d656c551c7778cf24975612e64431e7459438fd6698d2e3ab4f01ffe65cd8d
zff55f214a81e113d4d01b84da76f1823549f9c3a9cc7979feab96c7327bb592eba40a014c85c09
z14d948133fded3f65c44279322d77430805b0b335d479e22a15643266931e6faf328c454e2db82
zaf18fa1e5e1c3dfd814c6c9fba4b83b85796c629573b6ae2f380ec2e9ff2e5cb044b8b133d3729
z0f7cd027fed8f79928c88de819d7e7d72a24dcc9a8dba5919f95a35e829cd6f6389fada7723ac2
z60737e23cb18b6565346f13cfbdaca900046628accefed61ed2b155181d6fb33aed42453efb2c9
z22488342fc280570e4429ec54d1d41d7666b75bf9a9eb4ceb3a2b0d8b4751d1bc358953760f47c
z4fd6c7e660ba729c716cf31640d5ab476d80eee429abf027a53b1db1c5eff5136a8747b6ae9c11
z5ea4fbb0a912603a7302c1ac4dbf693569bcddb02303100497972cf24ec4cab52ac28d5b04ab44
z49c72df6966ce7f291bdb6ba2e2a96e4df0747c9ac68006655cd639d0a2d287953acf59739e7da
zc78254b749c0e5bb2a246d9743dfe610b69d7452a10cf4c1ed5858549ed99d4875eafda9c595b8
zfe56a097a0acc27dafad9ea27713b65bcb08a9b9e99657501c50456801bfd14f93731fe92568a3
z8cf52ce3b4e2bc8eb40ef26c022f111a030877940018b8165951574730b521c9f45faf7ae8e7c2
ze0da53e51948871cd78311e26141f106160f2980ba4099d23a2f26aa0112f61fbb5dd8f827042a
z21f6ad1f371c3810cb143e35452d769ac2bf9bf89aa5703089ba7d825a69a1f36b8e7ea6d8303d
zd54f38c1988c11f4546d7d6a51f152399748da237d1cb3a07009c22aac525782c75f64a7c3fd3d
z560c37717d01c8ec4c0ae67626d3d27c16da3362d64eef395040db01e2883aff580e1d1a45bb90
zc602ead0b4a9df749e949b0a630975dd6c58943c9bc67fd6176cff606a36d2f4d8598d6c24e092
zae94ae6625697db089696994a8f4024e39040bddfe01a88e948d772556dc02d31a8cb7187e2bbe
z13ec297478ce694374577daf6e47f5fd2c77d8af2e632133d0b5d8d8ad324e69e46551930cae49
za3d33da4f3448a6dccf32087feebb4b320503641cbc1d51ba522d6513da048f4bcd7c2b74fc867
z7d7732091a270070dce75b79f1d36460aed32783fb9ffce5c698f94676da02093ada41656c1147
zba6f78b88fad02a5463a244e68d3919a7d529ec21857db02a44a7fc99b012c35381ed8ab78ff2d
zb89a759832650f0771af11a72c655d90be651329ef7adbd4552e34f852592dcddba461718d588e
z430de1c8a4750b1666f2f1dd69c1eb8f8293b4eca11116a09100a44e409cd9875c880ddada32f1
z911cceb54dd88405cfd359698e4db942e39e7afc85f6f817f67720ba1769d71743b52ab876d7d0
z2a5d4448cd155da113fbbf2d4563af0724e3cc9f1e99a8491174a3105ac78dd72dab079ac202e2
zaa997a6cc2301e44581074291c9332799b5e022affef1335942ba6134e66a7805dc58bac563f11
z5ec98662eb9993881c573548d1e63f9cfe7d56371140d34b2781e1c82346da37295b89b040789b
z5b667c5db621c9989b8bc1f52e41d03120d4744f0fda5b74b332009adaeafc8e97b40aae3a263b
z6f22a31975b301cb6d668b5f29d6c71a4434109b7991a6d3f2cd412e9254ba1e59918dfdd17d28
z99fec5e93f5b11f751a09b60cd20dc69f9253edeef70fbc115885ccc0700be0abc736923a9bd66
z41d51284eebfd3cc2a357237a5330c3c3afa9d480771ff0d180fda18b957397225d41399150a49
z0a497f23cc9cc8f871e92bb95107090fa0636a4d4712a5b5c6e1876076d911bb661648d9df5f4d
z8a09c8500861620593577549f1bda6e13c80a1083652cafb41544dcf4582fb7d8461174551bfec
zd79288391a11692176757ff4b26c0b6876ff2eca73074612b64c76f8b43b6bca9079232b42a550
z96aff22fcf6075c4b6b2d5c8afdfead826a2706a573ab39a835c86c9ddfd5b9583707fa812d637
zd8a7a7e73e9401060f6885a32d515201b6d10eb2479cc79efb1643d6228c4bbcf8c28a2f9ecf74
zca1d163b9ee7c3a1485a9a92a394c075ae251d35894247937b8b3343d17d693ed99ac0efa58663
z4f3b2a9b474808f28c6d67f2a473928d50e1789cf3e163a231f75fef613ec996c01fc2040f868b
z736a44efa796b7e04cc3c88dddf8b425ef5d5a6222fca21100d728fe1c9a7e32226a7685b6570f
z02c4a5c0988cc9495bc93286e21b0076bedc4e2ea9a2d94fd58e84cdca3a862f46a556ab069e10
zb63e0fea0c1271fb84e8ade73da55ccc0ebe8f9d88206735ce69af55f76fd14ed8a1a3b38498e4
ze9a2c899039af34ddebf6254476e6c1f357cbee2b9b5d179dd17308e068fcf20d5c6200a22a0db
zfd85297167f9d11512c9d12ad37019fe093508674232eaaabd27af253a01b94e4ab188710bc1da
z1fef45ff82c74731396e31e78f01456811293503975c52f19788c00116e3adb5cf046cfada46ea
z8ad70e9ec00395dc17298f1d6e0be9e50d41a3b00e146f6fbbf9131981226ebb29ce3c7a130c5a
z469188c4a4aa951b28ee150577f0496cef78cc1898b80f0eae0ecbfc8ced9ea40a4af8b6b3677e
zb2e9213399b7140430d6e0ca3dfe4c13ae1d5efc009d698ce4d756e9d9abd5ea7fc4206efc8c29
z2acb8737ef9e6a67b01717a292913c5b392a5afd7bd5504f784b02c34dce2fb15f77bd9780632e
z4df37e805b2b733ca67702eaafe012887b3af9892259bd260070e51de382bcea7c1622d59608b5
z7fb6b8da0c789290b5cdd3942effd0ee0ccad421db9c2882198587af711dc341015a8976fd43c1
z750adc62ca6b049e2d7192d8551a11964d58c71aa64dffb7a0fe8f4b9d69e0175b485bffc1347d
z8eb2d4b7fd6de1faf63226c888cda50163e16c07e91ee72b9a533b9a5ce7ae733caab1c8992e50
z569e0d0d96e90d54b47156382a684cde1a515fe4ed176e03c93b0dda4b9610d2eed1e80f5c0e66
z3c67615ec99f0c1c71f41e713e4e754874bfca1abeef2e163a5e6900ca0254ce6eb3ba4d809bd9
z5827cc57023ebdc5d3ccf7fb7fcb58a971e1197750c49557fefb16ee34bd8342747a03c54e4f1f
zddbab0b63cc26bb8cb9a252c027cb33905ea57beca90fa2d8e371b9b6a4348c00f3569f7648148
za4bf3dc3ff02861388cd7bf7c57a9db248192373f4224ca1f1cbb9da7466a68e9a9fc54d041650
zeafce39701519a53a487bd0e6d969e7054a6dd56fd253e2e5a422dd4eaf5ed729e84ed59214375
z0fea5ad7cb0725c2bd2716b4c9769bd2bad2bca7bd753a124d6f70176643c6cb0c6f10257b36f1
z46305418f7cce85cbd2da8a321fd5b796ebe8931aa8742a604041ae18e9d8a9d76adcd86e703ae
zdda9f23867fd6565d064e0543b5616ac3e2719b33e33267bbdff45259f37e07f41dc539d7828f4
z48678b3807da0b2c3c835655fb0e696b280b852a2ab9652592e2ac94e01b6dc4c419362d832b4c
zf5b4c6ab1d9dc2dbe60db30b09e4a8fdac6c0d84c5f46203881cf788ffe31f42768b7993113721
z740a22ca99b3638774cb07ec36e7a885d100fdc7ad73ba86deb6321e04ab996686193d5a88207f
zedf964fa8a54ebc9f1ccca8ab66ec07867a27631bfb394b5de6fd265ab873dca0a9df8ea3ee4f4
z18b3576ffb82d2ce46af8258dd7b9e9ddd311082d82c2a54b26c5999c19427f3548595b011241b
z4e21cd8435d16e11be28bb73cf11fb8de1bf67a2efb39bbb6676d1ee4b81b7c399235f535e0b39
z1bb92594dc3cb131676a024106f3c8f04979bd488037a8d5f4de705b8a4db89ce90123dc08cf22
zdbb5306cd2c85ea534624cb68d294fa787e5d69e330c7be3f77d35ee496719111f0df5876f7961
z6c93180a47f7196584f08d8e486c0bbcee683f9f9b706010860efcae3b7c3d74b35bb945a4985e
z49b10d5f7aff4b3f0f316dc7503ec24952bf4c5b353c7223ddc743910d8ae51c06155a10844372
z2de67fd36c00d339f10972af6ea948b86ed6d91e35c86741649469668d52a2c7753016ea7e0b19
z6c454b7cdaf765eaf46672129c652421f9f2f548408f681e0fa93dcc885d375f6248ff57c218a9
z7adb3ff8fd80f820062032b17fcac0c6016e5ef610f270da60caaa8d63d9da5c375b877e184aa8
zda13b344f277509d45feddbc8696af41fc51a450a5307cb40affeea72c895ce5f3d6e62564cedd
z856920c5615571bcd943ad33201dc55347ce7db03beb44fb1f4fe73e1c2f014b409324682b6049
zcb1cead46a32531059087c488895986f555c51fcac33ce1bc2f004f38e2af1cfb4ed8f271104cc
za21c6f047c4245f2e3fd5117e4db7034bd7452d84935d352f1540eedc86b2e0ff7179af1ff80ba
zfb2a9592f3fb5c4dc1b21bdbf2195601fa8c375bcc2ec9622ebb5c0d5b8d945dfb913009b547a3
z26fed14b7d956e0aeb0f9c8d08b366a91c22801f4efb101b5c65438a02a092d913d59ba3eccdd3
z11566e88c3ee204276c5abf7c7edd8e77ee46f987044c574b9a2b2439777299d422924d2b5d41e
z637d5122ad490bfe13b47437466332e6801ad67f5b6aa589b8ef1d54918247d7b9a86b348a432c
z88dc243912f8463152a73d8162aa1d7a0b1affb3d6b7b96a9696b902e6782efb37ac53e3b8e130
zd4d46acd7b9f46cb5c95aab7ceff78163b8b7854e95acbc06637262bdd66dae80d1c46bf1e8cc6
zf1c2cbfc31ab23b9b2ccb12fa91d1898db96458181771577360e2a2d3f9c80fd8583ab3e6389ff
z850e85eceff6cfba8d9bdb8229b2aaaf018927a7f1823e2af38df902fb97bd88b98b043b133082
z13cd6adf3e23f6fc3adaf1e4916a70b0e6d2ad208762f671b0c7de4ba75bca284638312d828e13
z1891ae16da81c26e1b07e440f2f389699cdbdb5c376fb88272f89891380a215eca1ab6305f11df
ze7870e52f3bfb956db5fc8dd390ab120286dfd63913f4b0b6187b40530ee91be5ad0449d772862
zf479103dac97483d743f9016c99bd11649985ff42b9ae335aab7c628321320017a1382dff89c5c
z4da6197383d92332b57d5fb8699764bf1405457ae598480f8da22f525eb9b4e3b23ca1fe969b62
zf0c93e81d446459c7429cee05949a738a0141d505e7bbc026b17c49bcdcf88f64b4b852eb8884d
za7259e77443042458e74bb2f3d1c4229162dddc253000571c28ea97581f9811c9486dbe22ba471
z0eeb16526936095eeb74f1b29f0f06044d68be8832fd7d8f0d49ebb385fc2372c778b0842a1066
z1b11b4c86b50e1a5b1b54662cb977ef83dfa95490e366b38e43ea30ed1f071b962d8d488de51ae
z2688ce6eeb1786ac6f51c5ce60d8d4cd2f070e69280feb0a55042fb6f08695c0f448ff3fec9ea5
z884f1c9712c13dc1bedb7844223536bf211f39ebb828d954083ef0aedc5ea43dba2048044d53af
z26a8877e6e2d4f9a52bdafb8b07b29f854e0592024d286e21041c2dc8987c66aad63a1faab26a0
z32b92fa29f192c2ce4b7dfaf625e7191c6a72c14b201fb23e7da9a6618107adf6daf3284fcb032
zd3077a467e62e9f3739e1222d21902763a6cce49bc2d4e6d36e54ad24d8be5213db4e6153ff273
z5c051369c83442ef8d157e0db8823055b57e47add8685424fe3877aa2569d8c7b0c42ac7ccf767
zfeb0abdb1ea82fb7230356509cd3fbf0ff3e67d9b5aa6bc08fb810729b7ab09806768602082299
ze351c04c6cf08dcb9246cd47d51ecd03c9c90810a907c492e0e1041d3ff5cba0e49201120b2a74
zff8571dcd50e7fadf58dccdd47df5a4b670f0cda7dab9aaba2c6d45bc257cd0f2bdedf7c3b5413
zf623679839dc5dd21a0f6ab7b818c9650df665a7eba93dffe6f1405e1119fae49a88a434cc20fb
zbf41ab43964000e29dbb1f56a26dcbc8eb2a80d0ffc61f63f97c4aab2029ba94ad8e5359776e2c
z2cbb404146b80f98401ee09d8cff8e31dcd2424251808970811c81b7b322e66572cdd917ae4257
z2bb4c3fea246b73b3a5b6d842d0ffcb9710401b9b3569fc15777246dbcea04aff35d4ce3755ab4
z780cc2f2eb0969290f24dfd968b84a19d35d2149a2b7e230b063e99d090656ee8797f15b1a0628
zd7255d05a09b6a82072a53c14101baa57581dd61cc17a6560450b28f85a7af6547c3236fde27d4
z1bae6fd82e0fe7ff0ed2a271d30b376361cec482969bbb6419fe38f14c012838d934d3e464f2e7
zeb102a806b12880eb93cf83c1c07f366dcd51c6ad85fbafb6806437e30f8f9ca60e1fc82f930c2
z7be1bd6bc73867140815764e2e3eb962d2c11217eb29156c9bed06ae2a0f848c876d5551acc5fc
z44cf925855920d359f6e787c14d29c8904477d5be739f408a0cec0e261ec49f917c54c47c23d5f
z8289f65850d65e7232c45817365141b818ccb110523cb7f0c486451a0622dbb4b58e255f491994
z3d95febf5558e7368591a1e3d78428ce05b74c9979ffe91883024e0cad74c5e18b69735b50b6be
ze1d07036f47e28ce764272e24f067fe659e8da2b988ff769232363ceaa2a249e26f0f99eeda674
z956c86cfc2e59898cd833cfec27b2bd21fb0587c496cb04e6e16e69a71d2cf632bf9ce3d603269
z7fe39fee2d7d76acce01d6c8bd80ff9037b3dc906526002d6d182e36d035c6ebf1d4e3c0f487c6
z7c94ed0f9d202feb9f80eef623ee0d4603163ebb3a2017be31f1565ad40f3c2f599634df4cbaeb
za4b15fad8bdd1971caf316a686c25d11e2fda93d71df3c7dc289d96b871bb37885bf7a837a4c30
z5908668b8cffe1a387e3895b49bd5f498f49c1868d66593d9860795f46b7a3184fbe662b5746b4
z9c15144374f803c01dae8696bc4b5c96b4d3fc5def016332fb07163729003d5b883aad60eb0d88
za8d7e0648e84fb29861e79bdad6f1169c00be04a2f45bddb7ff87742f2aef950baf7454a5bc832
z17ccf9c5ef57bcc853b15f10cdd91ce66d55e126a97785f60e1f5b9aa738b207a66ebd776685ed
z4a309e7af95c8be0adab8f7b218da9154f994a1998fa2cec1176541ba816736793c3eb1ac544c0
z8554505f498d0676b9491df1cc15815eb3be010e2e42be4c4582981e8321e1c13f2370932e7288
z82ab2bf5390f4b5912995453e0b19e3e2e5c0c3a29a1814e28f391d0155e2338ddc149bbae455c
zf6c690e7b6466aefedfa2e5d99da144dc4e69c753e153984beae82104bb6adba0a19a036181670
z0aec19182d1bc7c7c4f0b96f4212353b9f4ba2a052071c611eecbebf4375c27f2ae80c2ce803f4
z331ea8332be7737b51888eb79ffb2e17e15690da811c403b5bdd509fd63a3c7a31899ed38bf961
za473c3c431a2e113bf19fce71372251a7ea50e9a673de8bd0a02b7f899fb90cbd27b4608b7d9f3
zac8edfac7dc16bb157be275393d05e7ec88ba1125505da38f14695e28da987e8f3fa8fedb4a37b
z4f3edac7502ca2eaa1667c11c9283b7c21136a313b22b5b886bc085d279fa25b31c7b7318d0063
zf5e927e4dd460956af5b7b80cbe419494602c134c30c7bcac8b68a874a0cdab740533d3b9e8b88
z591284368fc26c93af2dfab6b7f40eadd32dd0024a183257363b52b798e53f411ff6cfaa1b9381
z0e1d9094053ee3da1a4f05f0dea5772933dd8ac28205852f3e7cc50b511547a2a288624f5b5ff9
z3926846d45c9ef96a8424ee40afdb93aacaa3ba75581e0f158e12b9bee0bbbe726f04349010cd0
z15527cc7aac7ea90c5c89383d75d7cefc9ea20d735cdaa6341ef875e90fe75a35415bbf526fec4
zd801491dfec09c87171b5b32db273698c4eef2e1217cd8bacfa73a358912092dbd2a20bb6aad03
z2b96c9cc1ef3978a3abd46c8e6104bc0a2fe23c92501dcff4f5a8473810bbf31376e9e074ab178
zc38725b62e415c542549f6bdc30d6c2bf483cf1ea00d45477173012d98cd37acbe8511dc62a281
z67774f938e0a68164e6eefe7c005bdf77a4f7aa32d3b46c831a865c00ddec27ae1c3bffc468c60
z52df8a37c552ee9ef46f08054f6e08f4f19d40fc6a70b35a9f88769a1d787bf4ccdb676320a6bd
zb41fc142574a141894131a2d950c3d0f79ba78440e7d3cfe10a12506440da0e19edfe329e785fc
zb2230f2f8d1978420bc5129fb6801e10f479905ec995ea8718297995087fd63d63d8131aadb6ff
ze1ef415125d22ae6dd63b0a835e5830bed8220b6645882d89f119abf5f5990c2fd95f72a9563e0
zfef347b69db772093729f78a87107129a4c2143fb2cd2946a4c654308f873a39b727d66dddee11
z7fd2fb176aa10533d6dfcf144042b229d998008364ce3a602c8a2ec73dd3143d8c2421e608a0ef
z29593d459a9053195fbe5ed97d29a152affd9c6a24fdb011d11e3ad74767ce703068bfbcbb8a55
z14aaec5bda16fc181cbbde68a140b510c86bf1bcbcb34b4a4a882ae94acaa4ff5c670ef9710d61
z5f801d01543cf0f66b9981be82d28c8691b4acec911b73a6e651fd45569c4d309c175925f81df8
z9f11996d7ce03a943353d8575430a2512fc8ef0db8c11d85bab04676b1e437d8b6fbaa86e819f4
z69fef2bf736290235e6e3bc92d9ed58be0a1cf23c26774da4b3748493f3cbd12f8b2cc732d2971
z69b45bfee6f4ca67d16a280ae980c130590755979446b2b694af45e38b4b580928217f12d73d82
za1636bd5a89350305aa167b5b605938d9608608146e30373b4591708497e8154212ee27374036b
z18bee3be098292d01474d7c8501548fb8287aad551279cd866e035a0b68fe70e15393260656133
za9cc305035f123a5764afaa01b207d1ec8eb3363b561c0710e789a060296b099517562db36d45f
zce058090d51d3ea862100ad8a03da5af9ae19f4424febeb5011e9882c7a4d72c6355a6fa063b2e
zdb427043941ac694f2f7354ed293b63bb3a328f0a48e6495ddea6b69b78b2317458836dd8fc096
zd195650c3a2bb93d9e6e1e4a0dc07597e175099cd5c4f1954f30383c11753db7d0d6f1bb3afafb
zf3b84fbdd4cbd8d5e89136582811c04b9022d865404980522718e87f06f43516e46e0092bec332
zab9b0398aac04c5317b9289b4b9f81dac59dffd296292db0bb6e093685ec32b198ac736d672796
zad14138a1b38dfa00ee66026a585fbdf016c1a97f93d02a20aecea727e7e823a4a8d3794fd6cba
z1e1421eb2874bc206f401ed557b27e17acf5269ba94b25abc60049e59f65dea020ab8bcc23861c
z944e90b8d90e2dd37bb008fb5708ee07105dcd686f33b4aa1fcc8a5168069ef61bdb9fe7bd8bbc
z59ec67090a63fa8eaf126143b17e2095e785d796fc249a7c09ba8723e7f48fba4a8af6bbafa996
zc045e2dd5e1ebe787afb5081f8f8c3556b5e2b6c513705477261e8fc3e84a02ab08552a177b0c2
z4726af1907acc2a013b33f5f65ff9921086614ce2cb555985814b5bcff6fc63554abb0faecd5a4
z533eece4be024f5b31ef233aa6407402071ccc0bbf3790b9e7c24b0bba2333d58ae78a43aac5a0
z46c7d8af77f371c5f9d4133d9c07b982efbda6c87c5a967de23600702350cccc9848ba6493bd51
z30b0d00341fd5cc6a71fba59ba32337aa5f0a4a89bb0e54c17cad9eea51e3f58ede85c19c1614d
z3d6d6b32f67faddcbfb8a06bbcf0aa19882139204661501e4f4cabadc05270f8204bea08066e6f
zd5335495618357da925fe3d6d86dfd3dd6b7fed607dac022f097fa09247d2b042de7249c0724cb
zd07aeffdda86cd03f8e2fafc8d364ea23b07afd4748b371c2e19cddf250b92ccc24cd3700aeb99
z363634c28b64eea4c2c6cda559ec81884bd419b1a6c28323d1db5ec7e1159d06913cd377f659d4
zfbe7ddd79361c0346545a726187c0584b3b9ad0fd2f7fc64a13fdf8bf93a77fe69e25e11d37215
z814e035ee399f7324841788fe8a47a799be888ebae1d09421b3226118ed9df4fb269876b097a30
zf92042c53ffe923decebd82acd6406653c8a11fbd2732d0727925afeb45d6bd4ca19a9a69e03d2
z59d27db790ff70c539c0ceac424ffa951d12a80451312ff32c428d5b57154079ae8ee9f7c3c95b
z55910b70091998f50fd26406587658cfe574be0497b188b89738510a91d307507f4676bc5b6ecb
z252891973363f137c05da4740d9a5684e8476f968844063185e46a8c3240d53633aa14b70ed7af
z1cb18814215e31294139e0113cc9d88a13d721893baff5545bded13a75787393356e5f8c1344dc
z9c367d51d0656cc3d279fceca18f6b0332796f13da78af4b46e09344017e6f72fbce4c544224ae
zb4f2513035488641c10856f8380833cd17a46fe9af27e34aa1a8a4c39f71a2ecde2f0bffafb51a
z06f5f99be0be79dcd585d41d691975ac5d0ff52156d2643cfd001f4e5ca095a46de79e8bbc42c9
z7b1aa9602ffa8dbc1dd24ba6e77d4d76edd4cc22a1f193eccefc7b1e74af59b6012ab0a587d4e5
z353393e3fcbdd0f07e58982b99ab0bf7aa710a02d310859607c32e03fccb3f8b2304bee8546337
zc7b87fbe17c959cb266272089984266a5167b5ea824c7f2103ee3c856e56da23674e1234353636
z701c023df35e299a8bb6b9b1b743c595645ff1ffae675fcac1b12016a6a1b66a5ba8cf439d46cc
z43857ed4a52b760058495b37ca80c10a5086db14ec41fd7b73c6408ec46ae97950cac9e3bb1549
zc895a215dad70b8282be91a73b87ed0e79f28665f6ae95369350ac1c58267df852c4a21dc80ea0
z464d788ea51cd9c5a3be813a6452d5f2629120da57c290d5e799262aa22ff80c9d1622c24666a4
z518f89c761614faebc9e5f98079e4c2184c371a0102ad1e2c22cb4adea2e7b5f4e888003d8deae
z4b529dcb497c35da5798c8be80c38eaf72490563535c56d84f6e9c0c87e79b0a1da200cebd1fb8
z75c4b228633cad36ebdc61f34d900f578a9d0cab1d10e220c7f49eb38aba8ba5d2339be478fbfb
z023cd232ffd49c80258f19f89077309d5e929fdf8b0859800381cc92f09f1344320db19020b971
z413714f6a55ec8592417c45d6f187b0acd5f34220d44b07c4828153df13b860e9701b3aeb5354d
z6328eae126b5cf12beba26fbe823a7eaa9125f766e4fd577d372c4f21985ebaf5faf8f46e93bf9
zd8638ae4777a58a05e2f7a0a646f89118580166c72129d1ad8549a3884b44bdc3a0a1f16ecc6a0
zca46f121cc4e83abf45907cb14f03b9971121d9fb977786afe9f2fa22275ef66abd8050a75fa9f
zc505ba2afff31cfc8454d71221c8c73b736fa804fc3b5737a0fa044757ba077239c627bb71eed2
z9237cbb1814d3ee9286c1ebb14b33c101dc6f59977054105d3e79cc262fa819aef05432df631cf
z2f8388e3b0f2edcafddc960d9d57578899517d5b7890d73107dd81fea46c6f4ff841e7dedc1850
z23fd2d5d6651785b43e2df140a52e3268095b204b25953bb1318731cdae6ddc7eaad397f6d478c
zea9ab7c4aba6ccf8872e85df52567fd4ac8a2720d0d9c62578c19b34d7916ae2f74dea6a92cd18
z561e98e8a64cfd58df9be01ab1f1f207f243f4a61d2ad516000ecfa257c53856009f4573a5827a
z03492e21c671beccab8976b6f15890b828c39c5f105d3690440c5a547f24e2cf1ff9b0bfe928d9
zd7f29d0c756e3a41dd4f1f0c22e7204fe1e269d8314b976c4451fd25ff70e7220502853617f814
z9cfa7bd2e1ac0d6029cd8c52e2c6a994b8015a4574d8eae8bf0db7bf943b889ecbfb94eb04087b
z68d7d3fbeab16669e7d381c82a2c61397a57bf81c8fd300adc9258d30e85fb60dbf3df46d6a2d6
z6f9ad714994587906050a9887f859abd4ef1738b94e8f41c585ef07aa4298d06341e7ae5af409e
za1d2bedeb0cd04fa731f5f905f2695226465f4c8626bb42005e3b135122a03dce41bce4b6eef8a
z3e1c7db61b8bd03110c78a8d33a02de60ddbd6db8db4f0db6a0a43c772bf5decc3204d04d55914
z5bedad4c1efdc9062173d43d3147c6bad94d01e8bb5c86cff0bad6abd806a61d5cb71acf4059b9
z049286f37807a84a90858039df80277c8bfbee2ffaf1542e3dad76e8215e4e7fb8d619a51551b8
z8b74c1f29c831ed705b933ebd64ee0021fdf9b30d07515935c4a2aad067444c34e7858b210a781
z97184a8d13ac575098dbd5f3d4af5bc4f54383e163dafe86cdef36a66817499df22217058c73c0
z5ef765c5b60a98e860dc9f0a06251289c3366e8a30ea7208d840359d9d19c8665d788a7b44fdb0
ze0cf1db94c222b25407897a87529274cfcc2ca452b8c576805cc76725124015d1c2f5ad0f5b4e4
zc9894f02a03a7c09e42cd8c3549017f2b27fa5b22233b0b63eab1e5d9638bab4546c7a7c384fa6
ze2ad4719406bdc208f076095c693a473593373a2b2cd23dc00a8ee17f9b1da8d716490839c2d0d
z2ec9b13557db8963b5bfcd73686f72d7f2ef5bfb544c6c1087323518ae0253bf7d4b462df2260c
ze5cfda110bf7fb0123d7b1f59f11ca0a9bf309bdf214927edbcf4f843d4e21a0bec8ed39d80bd0
z67d6e83b95b511a975048d2353c69fbff528d931c7c66c32c6b27af4b7832ad8e74ed815f328d8
zf1e70d672cbd0fe5d338af1965104a5ce0c37fbacfc799b8ffd2a4da7ea27a0ad74d3820584c03
z183b747940bef278e5707b6895f00a07bef4f63f758cfb7ecc474db495f697ba35fa7cdecf159c
zb93b49ddfc662e810be2581e2591d234a1e7625defc8ccf97ab4532bf058de2fb3f1e8fae33703
zca5249db7b36b8f3ed7d5a503881403edc1006449429e053bc2e70034d361271a33de400a646e7
z8ce0b387188cb42e9a241907b0d2d9f432ca4a837816418759ae2f43854e00abaf1214d47ef7f9
ze6440917f41d924271b2b1152bd9693489bbd0a06cb5ddf388bc134229e48a76f7bfd370993a9f
z339c2878834d650ff830de11fd430967e13ea8d912e91f34b2031cbfcc4ffbe8e042b82249e61c
zbf5b562503207176d0bbb4f47dd3dc378cb142966fd769e90cd113d49a7da83e3f7dd63525e106
z7b2d25ee708537bf92110b40bfe5ebd8816d1252681b75755bad87c9164575357717c7951d99a3
z7ee0034a7027b2773d7ac1cf926df913fb15066c53c01ccd1d3347d712d530d5c8379b485f7cda
z091c1951f284bfd3c0fb2ae67118d44a5ac08c7376a6899c796a9c9765e36ae5a953fb5d1044c0
zb8afeeeb04800348054be4d27232dcde537625a77d685cce2fbacf3a1c71a0ab71ea3c0754a607
z7d35b1da82abf3e7d4764ae1cd68c071abdf7bd73a05d5753915d41bbb18e2eee0bb06cbcff709
z0fc25f19870c74fd5c043aea01c696ece5f8c9f55f175e8872b540525acca3857015da6ec3aa88
z7b3dd96e2f6bc39bca18ba5cad5d6950e21d005927485d9250561920a1a96b4ab8f21fee88d7be
z8cd7ff84db94bcc38790e871059980ec1947806e5fb940c5c21c3478fb40b6d72d144ca674ef6a
z0213ffaf64e2e0e75cf9d4236dd8f70cc92b1c37ca03b420d6fcb08c6658ada9e40b86e71eb017
zcc113b767c5c7146c57d061ba7646c4e0b8506c13657afafa9b7995242403ffeb615232b116d48
z0320d5b4bc005cd4f1150e0c8bbd6ad348473ee4c1a1b5f028b77c1701958b0f7c8b3908fcf8f2
z7b7b0450d15fe40b1f2ad4b3dd73709f0946ac66920fa7fc3adb5c316f49a6f05fcfbf366c7482
z25ae709870e17936321776adb0861be9b689159b3b2f0ba96319bf5639210d3ff695a2eb3e0549
z81cda33b9762cba7b27404cb3d781672fe5608b1c89a8d3c925956ab0b17f287610a9b678023fb
zfb5a468e1bc95761ebe609faa2218db5087f9cf1875a467946cdec706d658ac209dfd50d8576cb
z51247264ab4f97539aa7cbb7a54f3b4cf4b8b684171cd0080e6e0b72189ceaf685606c4d07703c
ze320eb0011ee82b63ff9cd26bf30870e996105ab315533a0ad3c3e30811bb6ee3854a977457720
zee6260158747eff641ec0c5ce5156ea2263e76f2a54dad137daaab26227a29f29725cb829f317b
z06547f7c9c607c3c3cca970ee8605424942096649bfa1d9146ddc688d2645de8c69e13fac8abcc
zbe929942b7c2be00f3475fe1c9d708aa092d316948f04a962a93380f2fcb4af69fcb739c307082
z993050c3234bd643e504c559f59a2b87d02dff10ebf223c5a1fbe29d3d1d9495096c73a20a0419
zac26166fc7c4c22dccbdcd9f9fe4d862fdea3d92502c9cad58eb04b3277ffae2a6b5ede703d5ca
z9099ceb208cc73e93572e79478eeb530f810a0a88de367468b006f0e68059c67a9c9412b536bf5
z9452cc094771cb3109eb0bc71b48c82632b25f3a5a9ea53106500ed4f751535524df0c44ecd397
zf72aa7b1d78f156b3c9ee92d0da70255f6d75d8b7b5ea69600a4cc084c482c661b389b834d8bd4
zf1b4ad8674d51f56ea64a64e724bd8648f316badee9453188f9479c4488222681137482e5164a3
z3484c6dd7260335359b2e1920864b098b2ef6c3ead22dedd873724eda3c629f9d8c115386f0945
ze71b5eb4a4605d34d75f5c03471ad469761961300a28ac0add1f416d739a020955852e11999681
z9dcc5de03c2f0bbef0edb3796f14c07bc1b627b63b8c57675b97dcb01aafaca8304773a6db7c7a
z44d1ec969b17f11f24adaef910428fdffc79a31973ca10a45bdf0df8e00685c3eaafe885346f92
z124880e95b4146c5e265454764653938c7ca91268c9387d0a4098608e19de74ac56f6f0515e57d
zfe97077ecc23b146311c501eb1b4e125aa7ee9ff4f98981866d2f2016b86b793b1ee07ebcbc474
z9caea1677a700b687f5ef7289849609514264df6dd260cad05342eb792ee0e761e25965ba10505
z20ac4b3c390e89323e02a9b1e46c32f183eccfac27b79e7c4c73ca85b7765ef5515f66192cd1d8
z25f0cd9336ffafdcfe8319082912d95bac6646d184a352728f3a31e31ebe8a6419b13def3db47e
za3d3c357d8cc76f0496b9c315dbd9a89b94354eac8e8fb2e89bf7d1e196f43eed2b8ebdcad4716
zaceb49d4fcd99328c9b5fba17765d8aab53dec3b24b75e6d8a9d6a4162b7993166807f7abc73dc
za8f2c7de43e5d8cc0517b07527c4fbdd0a67a30d25eaaaef9c44cad78223cf381cc8aa373469db
z869410dc49b0c2fb98cd742f7b9903d8af211fa63f192c5b37c1ea2746397352e72d0ba830c7a7
zd579d35e50c7570943bec9ef9ea752970ff1103d62d47987e82399737d4e5bb04a1a783ec4ccdb
zabad95206d6972e45657aebf41abbcad7dd6ec6d35e2155893b77ce610dd83d1322eef68858eff
z9d8477c3007c693b2a71abba6a7d3427e079b24a18447071d521ef612d58a7bfd4d05ca4b48462
zaca31b096357191099609927b52f6b8ff1c3e2ebe888460b2f668a31a1d5e6148e28bb2d8757f6
zc76480850b440f21da49b417021ecdc0ff26caad202c8dc01139589ade8e51cb286291beecaf1e
zcf811b044e829109df4e5046c759a2015b1a4969a50a3c00d8d9018a0d8c7ff29598dc961ca611
za712db7c168460aa498168125701467b93dc5ded27bdb1495f4fdbc81ca284819820b73a863a4c
zac1d619c40fa8542ea5121dd5cbbfb0159c9dfdef1e842a3cec3ee926e2facdf728a0ee6c38e84
z3568c64bf10227a3f10663f485edaa68bf745b881840d1205d4ccaf36159d3f1599145868b4dbb
zcc0b07a5db5be06ff7a6ad7cd5c096d5d3026f7d98999115669566e35d24483f0a65519819c374
za9e2a195c0b9f94e961bdb7f15a69fcd67f9b5d6da87fd1204995da1fb24df5e95585090b74ce9
z1f7edf7112a654afa74d9030466a0e095249c34145852f648bd56e7d35fa5a7f65579f91f88234
zc58168cd4bbfb046e919310bf7ccae899b6f21da8f3d8e835185f96c88fdb962ad6c9f614fcfd5
zf2ef72a5a3619ca3c4a343c62f2cc7e7f2c5b664698ac8f19c2532acf337fe634372e3306f2f02
zd6e404dec07f7ae32a672546c3817ce1baf97f70ffa08e98320854986a80fd92f5c84ee7e6c04c
z3edcec87a71e9738f25b6a36f942b6756dd044ca4c3f19cc4bdb3b45a15aab73ef2e280ccdab7f
z8072167ca08abe35d1b7a3d51167ede872898e59b130c1dfdc11430d00e74903727affc58ceb7b
z12565d7d2f0cd66d5a42cadb29d87921255947e03bb2c37b000054c78121cefc2db7daf43ae199
z426ae98eec05c2611b2fa71fd85a41b040292e71b1e568600927c8ebf91968025ddcc45e14fd72
z62c38683a0fe96e92393dd0972fb98957b5888bd6dfcacfed7f63b8eb66b91abf8937df7ec8b1d
z83d7a63e195f9fdde3e680339be68521913f9bcc5a7699d97a4fc2b3ad599564782fe463d0f0d1
z52eb11f073f2c65a6168cf0179b3abee38a2571ea633d72f38c929947a09b3f057c4da006cb6a4
z152f2d38cc854f981ef5fb2215c65450ef7523de1d30002771ec254a57a10925a570aa7f00b6bb
z19fcfda9ca3535f89a016a1676c49bcf1dfd8a39f14d142742d1a3e80b8f98f79ad235ec89d76d
z79acc455db242a4cde23e6fb98d585a4e843ac0500a6514d87696994c5cd4b5aa984bfa4f42b99
z4b44f447bb59f71c7e27eafba6f2f558e1693bb99cb0900330899c5021e04895b252b9f6e285f9
z4dea2b22dcac03bc7077c23c5aa10724f686e2f5cbe0273c43b2f67208472a1833c4d0a1f3a3d1
zf968e6dcdaf2d03dd88e1a29263329a3ec9959df4bf79b9db4d913d6df4ef4eb1d1ce72142eba0
zcd48e43ed32964cec63ea3f19c94d527f1f636b2230433dbde072177eef5b9e171a4a0d4075528
ze82423d70602441a9385da5811d89894695adc998b3eb2aae7ba5e94ba6c34b648508d1c2fff51
z48687fb33b730ec37aa235c97319d7894f3215af9813c3809b52be398d914ab7e9d781fa60e177
zf4366a5053eb158ab17e8b775083a39f297dcfd696b3bf55d81420d0546e29240c23ec613026c1
z682f1d1f430c12be38a3d3085df771c4c837a9e190aad9451a5723b6a0dec0a0e61f916d2096a1
ze89739dd596e622437956a96789bdb8e80ece432f1b689d8ccd8263168680d5494ccaf16c95ff8
zbbb4f6faa4abdc61fd12febd0fa56903e759594c0f81b4a6af1997c4bb4898b0e4691bcd7f7fbf
z20e4552659446aaeac87e743eae93d91c2637d12f97c736f67883bc6fbffea50cb9e7178e5288d
zd173d3dcc8b3030ad168aad8fea66eaec33b375997580901aaab42e7afccc20161531e36f15c50
z68ef4499cb24d5fd91b440329a3fe214b4bf80b06a6f9749c89e05359d01bc2b9500e78d9908b9
z1e711a98c86e6638528d51b959752657b5b739382b0764c8d4c57bd1c3d966e178419ad11e0f68
z2aaf10574456deba25f3695e54cca150e8c9a237f80fe672e695932e6c6ed59a3dec2664046bcc
za1486f00e686120fbef29219a1d51a01ce02e97ea31062418d4b75f6090356dbe673e06f1f78cf
zcded512bd4e39add31ab382a5ebbd28971b758f5c8466d393653fa6c533b511a3603b057aa7161
z9db27d7b6bcae34cb694442c246745c32f0f4242767ba7fca252962d205345fcda7c15e5d05531
z4d017538c1b6043795c0ea80094d2dc6db71bd2d8627930c4ac8e2a9f25420e01af3c241c543af
zb232baac034fb58a84cf858677b0d117b112b8dd17bb62014c39b680df2f02e55899fdcea3aac9
z37e6f27b64078039c2d8ea3c44fbc951ffeafeb9a1839307286353ba3f342c960c2a4aeb3e8213
z03e2a9649352b6d574c62bb8d7a4b9d688f0682eea2bb95d1035bbfe2392383c19aca61414fc05
z52ce0a804caabca6765ef43306ed1d5935c9060611298d0b61c8810ec91049a39299de5b9abfba
zf07dd16c1eb73a9d3e41021d57407aaf4c75c76145d9bd2ee2107551c27d834692220476565d2f
zc3a6ad6907da9456f03562faaf6ff5a969d5af67538763dfdb42eae5803488ad78e8b234eb27bf
z3ba9b955a81749ae96df8f7aa67c30044c7705eb6f1ef877679e8e1b04fe160c92d73e33b55a41
z883f558e6c77bc0f9652f7c0acb3a565d353302ef748b016083b074f2778b640704e1455144e7f
z0fcb56231206520514bedbbbad4f245c73fa374d62668274e186382985def18b9714ddcc43bb3a
z6bf6fa93375aa6b70c8d17c85c7480f87e1a1f75bc965e45358079bbd4d4a910a120390a5d0dba
z0f080c89215920d0d31b5af0c195ff19195a43404c0097145bb75058a1e4dc86c4851f8630b12f
z74c1997af357fe969269fd4e988c9af010502c0fa73b9fee74d80a14363a436d19281427301fe6
z1c57812566bc84593fb3aa6b31ad5e387ff7cbed2b2e00be73799950e7265c0cd37fb5851b62e1
z4ae1293a2605f6efaa070aef975d474b07bbc79a3cbb18a5ba9e0820af0a8d8d0c496271c3eddd
ze95281f1484e8f4c64510a4baa107dc3b3dd799bd1a2919af462834662338e54a3cdf05dc0e03d
z0c140ee70760c7620f101c056fd4bc1edd59283ed6250c2efb7db7d558ee7b37a9a032d17fe4d0
zc8680a0d3af85d7731f1f4b654c873d346fe2308a5b399b4489b72e96577dd6eaf343010f050ac
zdee6c9490ede94f453af9005f39bd3befc4d1184ebf3388b7d2e6c1abec0adca8c9d5053920b13
zd8e7f63c7c899a1c5c61eb52754650d73ee7fb980db0f09bf889ab2718dcfb70d1fb6e2815d55d
z3ea477e009afe3b6d4450da126e6dae2bd025fde891f14e5ba43ce1ca6bbd4e838e97e841040c9
z4353b9924517be8126af6ddd7ab06ba3bef99bab6246d1594b3eb117c3a558dabfe792b958f958
z43b3efb02c9156a46a1c9b1f20b4291d8d66b66fc4b3d531c613ebd9f2d3808bf7043e43879caa
z08eb99747c7c8f9b260ea0112cc97566ed647ac2bf38d5cd7249a54485bf0a8f74266641813547
zb2e9b22806f5d698749cdb43652af5456648e111fae564ddd264c602c65ff609774aff26f3d52e
ze6598f91089cde3537c1db207bbb49ac63842c10a6ba822953d78082eb36dd2c1a227d66230a3f
zb06b6002e5ed4c5b8e08317ff3808786f11fbdec2ea2a9395b54e941271a527a051b2ceec33c58
ze3a610c29e3c53d454a6826a7b3b9467623d1879bc4c2333c67bf9cde103cabafccf3c25eba327
z5b94e047bbbf7eb6b37ab0ac654af92461cef419dbb996c57730e36e73bf959d264ce7aa53a7b7
zb95153f8711fdb5726d1c311656a418f89b3bf69e331d7792eda2fce097f952d91056c7642b57a
za72f634a7257e927e7e1af475fee902738684722bff39197718263ea522d5b55b46a0a5e75ee4a
zcfa05031d26959eb87bff2e544b651ac9b30eee955b74bf0b8eb4c9c9962d78077296e32daceee
z3c2ba11a52cf0c2efc70fc3889852700c40d2eb258d6432dda96ca4b2c7f8e87eee6a6b2d207c1
z2ab236000a7edd9b7a2e36afd1b646385f97b2a07b3060027e20ebb4954fef8a5fa00882693c76
z40d831ad4be9f7977065e7f4720562577561361dcd83369c491f17831638a007e1d6c87709b961
z76dd7ba769fd00ee20f6a281eb5bb702f79136dc1a3e576ede135016dfbbe2d331c835e6a7f63c
zb9f038bdcaa2f5cb896fcba50723ef5bca06bfcf11bffd5513fe7cc3c303c135157be9a6d9ea0f
z14e03dd0b0b1d2c0f2cb41d473cb3f8f0c9f5a661ae56071e7052f6892440486471feb6ab85481
z3f1d97cb54410dcc9e04ad4b71df791ba2805b2cf8473b1810ecf4f5b8f24a0b984257be46b2d9
z15e0ca7d86b804c44b226a3042049d063d61a35c99d09372d36aa5547633d0c75787b719a5fb6a
zc82b7337dad294a4d9b1ce1f9aefa64a2ff560ed6ca78c55923f169f3bf38528bc29b078e063a9
ze655b7cf094d43d9996683979c824dc9629f35135a67724b963f292e2bda38bd9a79c2b08fd559
ze1dcf7acf59063d3c85311595a2137c58fe2b0fc05a46f8f2f27e05f8c093de0fbbee7ecd5abcb
zb32af9b49c1dffd64107411754bd69f90ba111cd2275ffeb1830c62ac6a3fcb70416c71328a25d
z2ec4969ff033dc11b64701182097bad53cc8008bda37e506f868dacdb530a0a06db8a6e7ecf72b
z574c818e226a3629c2075a99d138e46762c706692854aab4f41591ddb35cb5ee971ee8d2523623
z7ff3c2842ecf38ef9e91dbe8fe07bebf0edcd0614897eed39a1def3a1f9e5588c8614fc7df74f1
zbc4010e82a7d66563d90b7d800384e9f277c8cf1df87c5280309f784bc93b50aa0199e255c0376
z759f08b911ff427fb10d6551ee047889773de7c2d31a5af21db476fcd43d0b34169bfe191d89e5
z49bf238f73c11689525828a2c9d680c906cdaed368c014a1168cf887d9900b100ed40be53ca9dd
zd7e6ab78c00d67910fc1bade1569baecbeb427cbfa6a80b53f7d6eb62057e52aab9f58861bfc81
zec9849d339dbe9c23ac9c9ffe60b9390d122f926dcfe819cca1f13a31a57a0dfbdae4bb9183288
z149481a8e53c9d9b78acb750725057f458f80810f357b994e1aa1ab918c7f0bb4e3d9af022b4ee
z5f5e5d0a57136aeba5cdf8f40f2f1110308c6ab3b19cb4d03794b5b0b3d74d4a35e751e7fe66e8
z9bb041cf46e9dcc63171c39e64c44a6ef2e0808672a816236b702fe112618a4d34583617b4a194
z4e6ae18ab36489e463df804421ff5dfda46cacbc51a92edb01ff383463db143555450f48bb063e
zbc4dd58bbc510e08921e3518343a31bc7a45d1e82bd5a8ddf1ddc1020db206d63033cd4eb7407c
zdd5b677d5b8e0ef931edd0f1612c34a5365a58885added1f5e1085711ca1578683e03a9b17a2fb
z4147ec09fce3fc9438b6215af9867ea3e1fb8a138f70a3194297856c56781a828d4fd0017758f3
ze7ad383c67dfefb8291d517a9c27f86f3ddb0532dd18e38a1faa52409df42b54e1caee2ee976d2
zee726dd7fdd3c359bee6bd570363910e0feba83b1b4cc6380ea396254362a891efd785702fc5dd
zdc24e734688416eabe14f4b954c062b58b6e0afe6fbc914e738e4e837524a2f3800a3bf3f111b8
z8f7dfc8cbc9870d38d75fc1bbcbb881b36bdcc42334f3306dd66d506ab1afd11fc05ab4dab6d56
zd5397d7c19b207ada12f6d5aeed020c3a35b17aa94bea5c411fb5569e757f40e8e8e72ff2b478d
zd318a3326dd699ea9ade8fa452005ed210f1682c48950761085552b1e763827e14ba8e2b04233b
z10dadd62ea5be010803a96d90de564e5c5b574ec0d77a5fa584624ca1d83ae5f5c1d5be183e93c
zf3ebd0a8beff5e472c96253aa766ead6225873c3631cece990923267f9d98b9d90f9c16217953c
zd5f6c444ef5d8906fcc5540163a8dea284dfdeb08714fd607127fe37caee0ccfee55c3f8e43612
z92c417f3e2e903611004b8ddd0b8c399c783e847319b11149848d570b9129e81f49594ed2ac204
zda96789cfc8825b9ff9f855418563ec9a86bdc8bef2b3b7b4eb40667c17aecc80b52151f042139
z6fd0f3184b7015006a1b70d7d6a136cee64ab334b1afef78ec1759a58dd70ca1d2673b7b268ee6
zbae718f3e5c8255ab3bfc97637028b27db9c0f4c7a246ed977cc0d7e6838235e8f1e7f03e33968
zc1a92d2c62ea5ec00c89b50fafad7d376d30da89ecbc35fabdd53c6db80f954afa5c65aab2444b
z62a987e63302370650cbc1ab56100da152b7716ebf382dda7ac1e2a4d73734af62008a3ac85476
zda64ac888fcfc0a364cbe860f2faba3e1849a99d796b37cd64ebfa1c0f0878604a741a01ac1096
z5393e3e79634b56ecf8ea40aee10874461fb9813c8462885ac6b1dcd226b7c6174695df55978e9
ze1557a0e6d2a3eb66eaf6f16fe7b674edaed6acd547d3644107f6fa788c76e835b13f64fcffb4c
zba3dfa47164d81dbb8552ee601e3d78146f84d1c6cf066983f54f5de9015a64a2c93f2bb2182ce
z1e9e312f1bfb79071d5601d58c92340b885c698e2dd51f8cf57f88bf03f477bf845c9dff8180e5
zfd34a8e2379c49690863385a905020cb696fff807514516d3bcdfc727e254ef57a47c341b8be6c
z0ec5dee8d1b33eed96cfdb251490923ec5950e5d018e3ffe86406f9eac2a33b81c648926939620
zb280cf1775d273429872537bd06be2ca00a0f9597e3be32ab77360b117bbc0dfad3e285754fff9
zd05b510ce9d4ab0606a3a5684afc3f0b34d49d1f36489c3631b6c68b6877fa31c7acb7bbd63aa5
z7ff6dacd83c80516e838dfd9763485c7ca7dab44b4c376dbc0a7f0a9cdbcca6b0e376f9ce72ba9
z7ee16092933229d6ab8b20d8595acbe81e7ecf4d7e0e47538a23a1038faa0021f74cc760fe3552
z54bbabc7aa518018e65e38fe2b4c4a6cff685b518b0da43fd9501c20791d8069e4149deff6b718
z9a2a707f8069e9ca50e9c8e0b574062ddbb0a184ad5b025d356f61ab9f9cbce5de3ee4b0f4e8d9
zba71dcc42300d2aa76098b2402ee6695c6edbf1c1756f24266a43a68a233cd389e9fa8e5926695
zf0c30808454e8341784b1eb647c1cd0a7f13bc6e0ee1990bcba652eb006984f66baaaca027bf47
z576f353c44e19d62bbe74734044e12522bf17fcb1d849ef53af0ecb7a400e7b3a6ff6265126519
z995c43edbb9c5d435d04aa12391cbf6f733161abb84b5e7b90e4cb5e72efada5bfee13f0ef55c4
z285e06a42e80411e0dbe224ed4ade81039a36930abbe29999739aed20b7200dabcd2cb98bd782e
z0c32df6ab6528f7870d71783ea15f853adabad03b68e3360b6dcb203a661744be8b350608f3d3f
zce15ab511411655c5496ada59f94e63e747b6984613016ffb35f7cbaff1bf55a7b472464d5b2b3
zc6b429631418b0bd0d5f03913ffb39b5a15d3dca09a7540122f2704eb102587c40b0fdd9fc410c
z74e16a78f25dabac2c1b863757f2cc74eb56f6d997cf2478c2bc608d13792704d0bbebe4c12d7d
z008c6e0564bcb0715a6091706f3be260ddb8cb4fda836f40ee1ccfaf03d3a9897d62d3ab289b18
z73e3ba8be1da2dc28cc1564fb35d40459c31164f52fab598718806c1d0c4c5eaa03f95c92a1226
z9c04cc2f34561918815d4acea93bd6fb6ec5ab80c06569866a5ea0c8584d5d57393a0606318085
zf0f53952ee6156b71dd0e53a2a0b4f39e2f0741df2ac1516a05bf657f1c1b8c336df07900b6bfe
z252850280de73bba580707814271b7af50df2fd8b8ab9d6dd8b6f277298c4c1cb6e5f155187827
z7a807a35a125041b2d56e719a0fcadd1b69a9a9be22f1b961f6071dad9e223f714886b7ba7a97d
z747d51fda8bd3c3d43b12c312dac4165627d36e7bd69d2fdc4c7cfd796b59ff475facc973b426f
z42988d8cb6c7b117b51126244d8007d1d5c2aa1f393b77b5feed55ec682d90c0a238afb308c688
zf4f15af8f051f892db153a48f70563a3c50867e158653a7d7c28b866a939b2a97654635925861e
z1809029b91e0753d8a04dccaab10c48b0d59953a1220f80bc06ead319a5602a145fe910224cb7b
ze55266feab399c0a3aebb442be8c4c22900356fd715343a79ebde8d0141a811a241724c11405de
zc783d03bb644d65751b575578af8da822aed37388ad0b330cacbe6c21b71c9080e1a9eff9132f3
zd020dcb45c71d7c38daab56091adba5737b6a81631218544ec812c2c18d45751a1c69b159716a2
z96dc6aca9e4384db4c147fc940d7f14e27a19d818c435a6e254b1609010f20a0ede896c6240fbb
zca2d83203af0927bacf89feb52133edce000aeadc0c7f6e9d208863d68e0bc2079f6e12cac1d7f
ze12be687d7156b01f4760b319825b407133bb41d70399aaf7abc2173c3e522b21b2ddfe7cd0bb0
ze9aa2ddaa8c9e6b914903093ec183bd6690eb403d5f082e3173552476cc1478569e75664e58f89
zabb09fa4a731f262f965bed0cbc2ea00210ae01cea22b88f51b1b59fee5301767f3ada42d2fe92
zb5beeb3871e9a905d5acc8e827931f05c757698b97bcfc6436077e6fb79e54124da272c53960a9
z73e1065672a3842916d025500899f45376a81ee26fcb9e1d83eea72d1911327a4d42e730741862
zd5687c443646f122a042c282313297c62afe8f3546839d8e32cdd6e958bc6f913a15dd303c90e4
zedeb126b08037398cec737aced926f490a5b11b13f08ac6d2312d1d104fc14e1afcda42f6fe557
z055bf208d467c46c59e20563c9bd084f92739b2d1c32639a68355c9b100718d38b9c49aeb15c6e
z41378694df2bebd1b9f73521b5d03a631f120976068ad87e814af9cb85732d76571bdacdd1ec82
z58fe41952392b247ef1cb65c1d92ca22dba5878601bcbfe4bcb467e0213ade2d92b4e06b81e96a
z43893859aa4f83cf48150ec3983b04f11e0c08c1216f3c4b357535674bad6c6b8bc3d422067d21
z7185a37210754c3b808416ec8fb0ceb3d4017629e0946adcdefa30a6a94d502a8be8fab0ff6478
z64c63261c5a84e45542836ac5e665a213039242cdf7317bce22d045748d089f22e22ae0caa6b50
z4ac18f0017297013f4860f7c315a7c78e917df9b313f2f5316fa2f0aeb302d18506dcb2a328aae
z5331499272ab7d0cf1b207ffdcf0f3e08e6e61f2a4c695a5edaf38cb9b86beb4167a370ab3340b
z2f2e3b584e803f4bb1f3ac5caf6fe76e979dba1dc5bb9c4bb3ac540678eda6696b45b5dff29c1d
z4f1b7ee6c5ad034069746ed4004360ea9536df45bc8c5c95498e0498066423bc1cf702be8d0408
zace9c8e654293130e68885aa58c2e77b7ba1745cf4e736f928a6dfa9e6ad79568074298d5f8bc3
z0eea41ec9641c70f1be1539498986c0835221438d12c25f161c10fe338441ec3ccb45672a0da54
z6808a0f2f1a7688838863c4a348ebccfe6fac82f2ebea04e767f13b4fe30d1838515356c981117
z63ebb3682ba63613f7c17334b48606ba1575d5fb7f2f5990e100fcada5ed7fb7d913c3297ca4f1
za784bb8a29ed0bd48d0ca0b04cbb76fdec26eb23c93a791d6a46d89dbe0cd3e57761c5697f89ac
z15877e9b45d767a4f8d1d31ec4bad1be644239a7b4508328e377fde08dbb32d1dc3ec6ec9d7314
z4f4ad0ddeb661b7b880ce9e988bd61284f06596771cc6682ed173c1a0648875858c27799482f08
z6504664010151a0686d5a63d20dd06e553be8b69319339377d87c6cb3887b709c280334f3ddce3
z7ec783a1645fe9519dad660919e691b48d8fc291172c989b9da29dedc92284524fa920dabe99cf
zf2cf86ba42e15483f484e66f1528a05b40d80523956777c028abddcf5b37125f09b7c3fc32d3b3
z9348abb9a2ba7b9b44fbcdb2f0fd368bffa647306166a0bf02c8c2e62dbec7363030c926023f8f
z2bf83537e24c1096108c4d2b737afe09612f904c188434c18b56d206a2c9d79dc26378c16d4a13
z8a8ce158c2b2b4fac6ef283d148c58e8c40db870c2b97996bb46dd374b0cda9ed933ac7c797da8
z34a21878ac120899ff213f87978d0761ae308ecccf2ac394f5dceb9c97477e1fb2b330e04d4349
z189aaf29d75f5e8c5edca9ae82e740b4c74ca78be4f7b846bb20210d6fddcefe359505791b33d2
z7e6d01f94b93b54473c28ca55715e0fc1a7699bdc3d01e67750987681786e20ef18901748f704b
z2103b07a63d9076021cdc1bd3b62193637bd9f8a6d0d850218d4d501d39f380d1469f7fd85f062
zdc737ae1bd0ef4149bcc3e832cb99931e3926aef235b0c5956e614a126b283c12fef16f9d69848
z83606c04bc22eae0a6d8cc21e2e0465a08da2a8e3e50d4de97be9634b1140a28f02bb1b3590d67
ze3f3b9c334bdead97955638f62d447a0b53241318099ab133c832da548044afc2df303d307e748
z28a6827c817951edcffb2b05e30194800870b7efd7f27700f24fc47a7e2ee9a14b939015956557
z7d51035c786ed16c928423432f9c02ea91536174139ec121b8e33a76a081fd33d5f8325513f866
zd9a1e306a049548c3dcf11476ace5acb181ec8fc4bc23e74157b00b9743bb47bca9e638f3510ca
z26c3d1a54e88cbef92b4c6bbf61f3dcdce279ce3b5cedf9a524bb6af8447016cb4069a52f268db
z8057a4bfcd6c7673ce30ccf8f173c9608c0fe75acdd631ede17d81af2bad2ad10ab4e1483e9afc
z81065108db9660b2116c0afce9b9f705b187afb6097cb91b05716e360274d528bedbffde7e5212
z80196f880d57f10b5c854acf90dbb25b13b289115042e8ebe7130b75e0dcea6b8a60c000428beb
z318b5a0ec75eac9f29747589293eed087a0635a6163bafc20fb1d287c2b62b9a5d9317bd494b7f
z8fbfce820c8707d637d084cb7990d62d972a7afa38436146cbe44768c8ec3d8abb9d19bb46af3a
z218c514ee100babc3fc952f5a0f9f286b098f586ebabc12cf1b976e82ec73c8c5d5bc56ff050d6
z71c8a735119a9e41a3944160d296f6809e03ed76796fdab2341fe092066d66ffa98d32714b2371
z4207840d24e7b1233e597f1257af8acf23b161d16a521685116745468344a6928fb3384ce7f447
zff1ec60895b52c454d5b20a746c6a1eec2a628ffd40e9a0dc89ffee201d3611883f44e9317c15b
zcf2912ca59c4286e3405a2664b24b1d68d732f2759a179803df0c9ee98751e5710d6a097067713
zdc7164fe0cd20599e596eb0e10f3cc82577b459bbdfc1d5f7eabbb8c78a7ee4edee718b59debab
ze5745995d9b56d647076d6376e86efe5ed63ea372daa6872e5022ffcf69e921e9af4a1221e5ad2
zeae8deba2e4ba1d93cbd54109f4e1a0c1f027ef265901fa50abcd8c812e63b72e603413e64034e
z2e9cacbb0d4f3ee6d567e115c64d1b834ece303f4cb33537ae08cd037127004489a007e52d6c4f
z5756807cd7d7b57efb5d62736470eb571e6b1c3d7dc4f1d8f9010beb2d765e92e393e2bc3a3586
z8e760d1af72063533a1d8c3b1d78986c283121488e4e40aaf56b810449873f4771607e65f5d9c3
z6fed69c6f52a0ec9c29353f7d6eb55831d08a1f62175f010a415a520ca56f00bbdd22ff3ac2624
zb5747682a8650b5df483816d5617181a456c6f2530b2a27f77204f0eb331d7c02507164c17c1f4
zdadba66c997473752a6e15e9c523c6d12ed7fc2920897a2e058aceb7464a0d57907e078a61cfba
z03b94f6f1350052770cd411eb8a37ca420a64a13d9e2ef8dc84290717d79909c7b0e536bf0e9e1
z9bd4b296941f452ae163947374b7ea671ba9806ce385d92e6156b7bee283a375490119b76f63dc
z939cef4765152654219e5f15acf4a56eb54a41ce97eab23c33cf320442fdefe7aa3212a8cc104c
z0a42609073fe36173b4fab3e618fe05adfcce282a6f2b864fdfd3dc7210b8c15ca0270c94b43e5
z7f25983d9f65a7e451070ab2885a92a474b73fc66f994b35e8900b6d271f14007d45d43de17e41
z9dcf1e70f0c5d5927436077086d32309b22efbc2f6b77e6dd9d7192f15d2e2899f8a2e2a1aca34
zdb9dd7dd539446b135f8b1b203772abdf30657a3601b4d30f3d5ce901194088da56eebad1a8fe2
z32c5481995946592cc209b80a9eba8df5114beefa94a83c82a8fde912a4393b39c571a1b5df5ec
z9b85dbcffe765db656d7bdcda02c3bd86d1618fe1505e11aa82bbc160010666e9b29a110ca5111
z90e64eb29219a879e3343b1982aefd54ad8ffb6a1c527fbc582c3345468a78ac07b678440fba86
zf295a57c661e160a4577b456aa046c45620764051491dedb066c15e70af79f0abe346a81787a41
z2d37717230d66e0fefcb536bead7a50ec58a73878838c09481a2f8e1e69837ef0a6bddd2f385bd
zbc5c5cad494137ee91a1dbcfeeb30f1dd14536b2f3ba5564ba7763e94b834957bd6b9828a56cdb
z19f3d2dc1dd8e0b6bc12a8954871c1e7f3aa2fe043866a9d7c8b40fa04
`end_protected_0in
`else
`ifdef MODEL_TECH
`include "qvl_arbiter_assertions.mti.svp"
`endif // MODEL_TECH
`endif // encrypted_0in
