`ifdef encrypted_0in
`protected_0in
ze74c34e226135848fe16db9ffd31815111b6d7fb642c521a3f628cf6da949865580b22efd062a7
ze90adae0e65e66a2c36a587d0a790699161455169ed55a01f2084f11770a774ec4c588039b380f
z6de9c5084882a40b79a175f5c2114b2b6d78b070cb806e1c0aa9258297f4687ab308bc470f0040
zb0b1de382961eeeaf2e279e1462520fc31c119af8f2b214846f56c2b3cd2eadbe4099496abff18
z15cec83ec4a77b868344aa20ba7360908f5c0de2a79abf8b3534b883bb12180f68b5d4beb444cf
z3fba8f13afb0abfe8fcc4294810f75afe452434d2d0f1166236c82f76edf1e12979f04bc35693e
z32ae028996dd85737a8f5adc1ebb94f39c940246e887647b64782cd7ab429b0544c173176cede7
z01dfb26b1f73408344a52b7e1f117f12bb9c8077b34876c2e6fdc085981637012dc9754765e1a9
zc512ce062e0b8fb16a214591f5c81e1353b900a611fe1f4886b57940b41b7f2ce99a7b84b04b90
z916f717e73bd10589c81e207ed77ec660a8cbed5b487fa50acde1b055c8870bd8676023f21ddcf
z9c98cc47cfa2d654ff1365d1f45035a045a66c5dfa8279050262529d2cac9e64fd27d9c7de62a7
z731bc808811ded9016570962244887f98fe5440167bd0088f2f049df882af501358497c3b28776
zcdc5426c7f52a851c35106bb93e16fff984784050fc808fad15da330f6f0607eda2d0e0e4b1215
z2ac5b11453f6b6c5c6b428261a64553d70b4ab9f1b396e1048595951af798d8de75c23e123dcba
z74156e068eb331e95842c597f3ccd341bf87af84cccb14b945e8b236b74bac5b8a2e30b2fbcf85
z4440501bc40f64309e7a471ab1713c3d50c22d96e536de2d04cfd2bb0d83eb6aaf04a9877de238
zbb5caa1dd6b5dafe5c4877a0da5950b5aa1530cb9c4fe8331bc938271749f1da474b2d0fcebe6e
zeb86e30abbbcad3e690bb0afae1cc3f8daa978b294fa747ac1e61b40eb10e5c9106e9054787f1b
z551e763ce12a455e4f49eff66134be3beb6a2c4c7d7e37035bb6855eacc01199e2e8bf3e5f1f3e
za908e5ddfbc8a389e39dec028de75c97e43711fbd959290f8aef9804a45d590a6f324148150c20
z71ae80a9180fdfd6310b03d05118e69c73ee776b8a8cf7c11ee1a2235471441518a5980b786f52
zeb68c952f4679a6afab6d7a222d5359145498a02b9539143d54478e00cbc9958dd183e81a4c1a4
z5d46b5d3013d4e2bf526a832ea07408fab4b1d9dc6ac670b0c4aeac5b27e3ce626c6c01db16076
z62b221052cad8d97104463aca4c7ad53348293e9a7ae470c93e3f39b52c58c66efdf5a49107ea7
z53ea955381434ace56517e9a4e6464d7a18799a447e8ea2b0043129c33cce1a4f3175e5ad643fa
zcb3d50232358ffbfc9efc1c7d040afda0238365d22a25d54fc0984e228e137d259acaded2cd853
z79bdcfef66d4a608d2c4fbf0feb4f51fb273cdb95c6d8faba2a251e3c506aa306fb273e204275e
zfe3f6626a6ed96e7b88e9cdb2078589c42f9e3d2798c84a0a5ddbf227f1e30c5bd1fe99a04406a
z8d557b4e0ea37a3121066fbfeeee23c1229113856d883e86af74c34fe5681376c62d887011c2f0
zeefeaa7b707072050ff1910a63dbe44b3e199cd5ee22f5faa4aee9060d5d5326d54e9f34cbadb3
zaed70ee17fa5b869b537470c3a8d61de3ae582d900af3adb6575ece9a41bc0e6580b75e255adc2
zd5da14fcd88d4adef5ec4bc891f14d262da84920094dd5bf0044cd5e59a50c12db43179446ffaa
zcc382a658ca618dd2b59b1692c3f258e283766f13ecd75e8d60fd25420b2228c0a94117d52673f
z5ca74aef84a97ef9f7dfe86a9dddd1357f6e5ad76ac8efd329f5fa3ae379b65666771a66056793
ze3fb2b72f1883d7538148183a7ff6e44724f9b0fdcca75679d83c9aed92be74ef91983d63e02c0
zbeba46266e8160d810a7550adc46303afb2b621dfa14943ab51fc9617b3a3dffe2d7c6dee35b03
z66999b5244894809c34e2957a21d31baa6ea83620b80ca357a2e27dc96e9d68d4cbd3b7f26aab3
z8a9ecde402394e56a4706cb8810bb4b1c49618189ae9e885aecd90f7fc29515b4d34b87187689d
z39f612338b92554a57718a1b03c383224e1094fe6fd73cc633432db358689717e6009b3025d098
z6bea79a8b12b7f7cc98544def0cd4f39593f4993ab54247bcb44defa9224b09cad962900aacf25
z71e710f22acbdea76107528fa090045e6ad0d9a272e8f6707d3446ea4d7f58b5c05185da9d07b7
zaffea4faf5738030af96d466a3912fbf69cbd7c2dffb5118b130af18ed525f4dc1af66eb792e11
zca3c25ee37b529feab421c9cf585a48e16753327a73ea26880488dc82784c39ef29c41f9721a4a
z9b65df106fb87e9c938a811aed4c4178c35afdbfe2298a057b3484477145a320e0835bed433cf7
zdf079f02b0666223e7a86155b3d3483d046497419b0965989ce492a8e0b693729ba0dea0ff1e76
zdeed7373c35be0d34a1bb2025f791c0f8cdc1cdc6741c0f0a1e5c2ba4a79f2410a1cbeec701e90
z6619d73e73264bee304b9826e86c320ac746b52d219a8c01dd9f362019bc54dafcab69ea7ca9d7
zc9538a4320eacc8b4054aaeca4b71d9555a15e2b034e1f959f89417090c5e675a48c8f16be905d
ze07164173138a8165ae4fc0e63292a8b45cce6b18bc0b3256430929d5caf302dcf463e11e45434
z0990b8bdd4263e3f4cd24769d307c280ad342de44976e33b815270160cbecf8970985ef6ca0fd8
z58fa6086d1afb9574586eaba1fe91bb722128fc241b5d40213cb9098173a7a3179ba2405fa6c5b
z33e8006c5f6aacdb79280022a14f028eb681d4de90f7814722fa9ed207097f167d281bf49aab46
zc3534d2ce9ce6a27a62bf34b9b4e249c058e3342e217ccb4e08936bf86ca3edb8afaca245250e9
z66089ba3460ee8e168a474cb433e342b020b82c231236e54f06e6152c2abc3a98425c23924e34e
z38b83e6d1bbe4fdb501db41b5c3c8f0b9f3af23d4065c0ba38bcd0870dd810ff0accff0332975b
z23e7fe4d99541c3f1a8cac69bd81a50f7c198d2a24a5dc2872cf08154c9ab3813b63eb32cb7e67
z815c280bf45fdea3b9db8367de77b7592c348726ff3db90aee6b149b357930bb726e8573f834a1
zae25d5667f0273a434d1119c21d47545a4064a32205c6e32e67c8a99a2e80bd10fd3de88654df7
zbd99a112fbb462c675a38f21d4962c50e78ec0d49e6e7e920fa3954c3c65bac19dabe5fc4720f8
z3b525797593fdbdf3a7f38b725287213c16ad5f397fb539b16dfd7a8524c9fc45970a47a888432
zf5fe733dd902336e3ffccb8b1d86543e1ef90f8f41fa3b1e247124fa5d11d5ce82bad059d257d6
zb807ef267c09918f58724b39b332083a4ec714c892b21b054809a209911bd6a49838a0986f81eb
z9ff9247c4bfc109817d2e5f39f6b756eb69daad49ff6e2812bf1fe4663765043953b576b30ba73
z6645f27d903e4cc5f85b32f0eb31e47be43ec3560f307bfce7a4c1740920892c33b0915c5a36a2
z54b1f12e0fd006abfff57cb3ffbf6570db818d79fcbbebae93926daa006de030fc16438798e3ff
zabc151225e2b9b59586d3c5a40378e21a5b48b90c01d8322ead100f77851999979f84bfb0702b2
z546d97990e271b407fb054bf5fc310c6d92e6f9807ddad5271ecae07ceba1d4caf026883e645bb
za3bfa80c32ff56a5bd0e1198ca227d533d1c1f8946f73a97c7c3aba5629767b66c66903b341c31
zd5744c5f90fd7f7affff58de9a9d7641479715b14d73214923dc008e6cf2abc9adcb95fa64c072
z41ad9b640029a9c2d160d27216d6a4063228abb722a0f8996b19bc147f6ceee7927fa65012f82f
zdee34720df8251fc3b17867c51a48e86e78677fc2962abc778ae41cac0556840ca70053715f208
ze7866e284c1353484af85d0f35947b61217c275c6b8513309a056fef4882934d3386e401e21935
zc3986f47a49de06382a737c687e7e654517e9a6aa43df87fa5b29711cb17b7e7ee5f19946f29ee
z0d48271c1ade7a19f83db6debdaedddf15871223332d70b83ae7c85bf9fdace397ae681bdae1c3
z92442a22ff727e0f8f7fbd546585c5614c84bb951d02262747bf88e393893af1cfb6016802c58e
z9bb96b39133c42c2a5691d84354f355b7dad7e8f31b8ce7c7ab600f0a9f31728de8d9ef5928d27
zcadebad9e5194a6aa1ccd3911d3a10ff32c986fc34e3ac3ac543605bc696113d2c2e8725ccd4c1
z02f3758463132782bb8d32bcbea93e732232806e8191901f2c33a4b095f9882156daf574bde26b
z87229d8a86a54c8cba72a3d5ceec072db7f1ee996ada698b250235465465b001b84191521bca5a
z7fd2e0d2fc4dba6af3ccf9d3c387665f1d50d2c1c99e6c1117f9c7cade6cb331552f02e8a6efa7
z7ce268abbe74093b2007a8010765684dffc7f39cac8b082018584304eeeeef48fd1d1ddcbe14ab
z0d18f2d230f6b8ab03738b0ee90ea0e92f53f2b53b3a9668764846db914503c3d13966b9a71b99
z6391531ce88f04af68d50ed3373bc1e81d43afae2a4370f63b0eaff12dfaabd0aa0b2c2691ea6f
z8ec555bff81e9c588decf3b9ced0baccdcea5f6bf890818403704d8e9beab46ba519eca52517db
z7deb480a70e43fc063853503d1d371d0b4f4017731d513ffce1a5e0e24182f42ed852c51f26e6d
ze194ff63357a4b22767644f9e7102b0d43535123cdb2e1acfea1da026aae7085b83235f2828e24
z874cedb1bc54e4e5553f8a39804300d509abe4e58477e4e0030706e75535709a70ddf4b2e576d7
z2ecd8965780345712ef2f896ef32b9c7dcbccb36120851c02b1642e836946d27624ab423dcac03
z0dffa5927f6e841440c7f1de0c561183673f49a214ab1db9ad199f363166f25ffa079240186222
z6d7eed9b24d0fb0d1af4ab450db933a494e2de0307db95d2e889c03fa03708cb4dce097fb4627d
z261be2b92a0aea05b8d12ef2b0433224b862910fef4346678088b44cf48944fa1d0e1dfcc621ec
z524a3d542d260b69541c6d47ce6d6bb1bc2db20c034a197b84bbfdb7af7c4755b37e70f0ea9ebe
z4972a53220d6c6d42eedfca43f9ef0f6ec727453d7b7fcc67b0e731d669e4ac2297506a3b6b1c3
z3071603d132b7183ebdd9d24ac166e32f200db2c725cb03abaf4e8901365bb5e706642a107dabb
z30baec33d467e4f3f32413d6a1fed8ec934c46c8eb1f859be24b35e7092568fc6aabd5f16f7e05
z507cbe7badcdc536d209cf755648368575fd24d5f24c31deb0dc583bc9c422ae27d2a317830062
z53aae6c159e9df6496b0f8b897b37af2c6109a34852967ba854cd37ea1f655c338a6290bf7d213
ze157036755575b915c428ebe9647ce5c7fa621f671397a7a3f631ffa1c146c6379725a35a89823
z890ba9e6f33d7a3ab86dbafe91f6125f109c0fd0994ed56740a5cb991ce3b47bef9684f5d3bea8
z1ed58069e769665ddbdd4bbaf33153ca4c3b14be8bb8b1cad12c0fd28d07b7f83ae306f64dba45
z4335c161f1cffa0e51705a222e8479d38ce9af1d920a71750f52e025e743f913239a17306b595f
z644493c771e3dac6c2787a727e5c15a86a7f23171f11266905bd424bb5b98e20a1b925beda68e0
zba258ca99136a31864beb63261855eb33f1f7bdd1bd593abb189dc84a6c144e70c24136004577c
zde72fa4f258741d6b928fd3bccd0914aa0e30d6ccc0f8f7a860a2d9b06898f040b81ae4cfccac3
zb3863dfac2e85b7538e171e1e94863ebc98ddf5163b7ce2f95ebb7f88199636de45d00c1eca9b4
z0b87bf96e43f8d7a9d1d5fa72ae4931bd3a324d5640a305cbea97ae5ff075d880865ee51f9ec09
z02832b1274d8cb612d647db72baa1b7fc5ca8c4df6c220bc3f8cadfd91c69b7e976f1f3f2a292b
z43dcc7431d93bcd8038cdce2716a498ee6e6305afd43edac81571d05025ae66cf19b20f864f2c4
zcaef4568dcc70b6757ea97aed1f48c1f6db432fa6a78e0421079b33210b59f1e8bf6207ddb9212
z7cefe07d1b6c296767b6d6d2f03fd3cbc7b40aa4eeda51d0e1d2bf3bbc72287b8fccc6ca6678a4
zf39cf318a45d99bd7ffa5c2f23836e97d70576b5e1bda90f3e5e032ae326400b5bf66275107e72
ze8c3dc75ca8d11e121c61044ee13c0fd414abcc526588a44c64ebc7ca119506f69249cdccb4f16
zb674e10bec479d32741074aabb4d7537c1a2b4c55b18d9cddec7a5a484fcd0eaea286b20aafea0
z6303209bf715cac18656ba2e49557a3cfd415661f204a8ac30bd9c5c7a062bb42dd4bdefa93341
z85c3a273bdd9810a4edc3d380a3383d94078a9aa097f979abaf7866deca6bda4ed89b0a27ded7e
z18bda27288b207ab833d8b961690ba94a3e2e2992af364fe7d16cafa574263e05a989c87ba213f
z2b61b8abf2722ddca1ea74edc29706b49f3c979d15d656543493bdcdab0d1ddbea26503fbde5fc
z55ce9e1fe71dff7c7a304124fa49334e144ad227c8983776240006fe27593af3c69934a4ec0a3f
z9946b7aab7adc9315ec51a60800b11a89965b144c34b24a98df7ea4252ee963354537abb0b5d6f
ze5bebc7168bc17a7697fe078d6adc6c61de8b961c906ada58b2c7aa1de007a4a5d4e1acd8c178d
z5d936c43d58d0d68673582475b54d7e24fdb1cf88a828cfaf5fd26ccf9e83cbb945835dd02cff1
ze469401f5d0a736aa291a4d7dde97287cd5623cf33df99600563c0b43c444e316c3f8d6e50e450
z18c604ceff0ab56ee76ee9ef5a84ad2218b20758b2872d1279ed04dbfe1eb80c39d7bbd022ee48
z4457a6c6a30a86a4a52904baa144727442711d3a453670736c615f6676bf99196c279046f1679e
z75bfdae0aa221da7f27444d4290aa5069b520fa284f22dcf1ed4f343a45aabc1c6e4156eb47656
z7e41e116b2cba1ff8910f2594e33945d417b66a154e93698bae2f9520c86a409ba108d68db37e2
z9567d2c04cc382fd15043d2900a81b5f12281959bbe05a15a0d81e8537bbf01d7b7dad6ce49cc9
z7a20389afeef9df79216d0849e8b2f8ed19d6b7e6a04044d6d166545b1476af3095be0ee360339
z88dee922e46f7c044b997b965a25834a0e848b2bae0ef23382d098c82ef73e8b7b0ebbd2c4c87f
z64df2e3419fd1cf1e2de16f2318b2eebcfff569340a7bae6b8748557067769f848aa45bb344ecf
z385cb8cd7134eb533ab3269ab8032fedab034b42e5c1ee5260056c822bd0a2903ea8deca85531d
z648c71e681a3e283209122b512834bbf7b9ca6b21c77f480b589db18179952a0a936c16878dc34
z2ba40a4b4a5e43ce0e610dc5a491cf77f350f71344f1bd2bee821a7bace6709fb701ad58331f08
z5fc00555dbf62ed8c0ffc561573140befc75cb8ed5e49e1abc4ad3f960437c02bfa5493e304b1e
z09fbe3ea31bd7ccf678852ba7ee6d95c28c6305417bb68c4a0574c07995146708390c48bdee6d3
z3d4d32391b99a4f8a1bbb4f079472e2cf2aecf59cf10c0288776767f3d13851e52d9946ac3e8f6
z29f7fbd99567f2bd474471f2ff5dd4d61a9693a1f58b4189db8dba033fca3bdbf303d41d267468
z555e180194938d385dc952e894b924e928904c9dfb069f8f044ccbf8a2c9ef44750938e84edd43
zcbe8d09da685f7a3d468340115d15f2672ba5c44fdcbd0d6dcc96b4cbefae85a0b23e62a2cd099
za93d49cf5763b2380136fb7853499db5be5bb2e5548e044c065b46a15542f38e6fe52ed6a89735
zed42a6a0f9a6885210404b43f31595a30e1221c17d42e6b188274d80388e47aae832c47d830d4f
za2d5d2868b11bd833f95d1bcb89ceb1884619e9584958736b750ed3b5a21da253f39231accb844
ze5804142ec92ba0c9a32f0e5b34cae34cd53463e06e68c438269c50150c09befe37db7ead51c54
z6f9e762babe3682c21986d9da739e516348a2940cc1f7469b97b0996de2623b4be89de5c4b2a9c
zbc40eed0b73c3bde742715539f4141eba70007d2e47fcb699e73c307bbfcc7bb693501b054c88a
zff21dea8d540d84d7407dfbd68b1ff1090887180d1b27aaa0b1b78b9742fdce5aa8ee46333bc6b
z0e81972db2793399e5f164beeaee9fbb19c60a1d530b094326c7dba7fffe5962f6fddedbddec03
z16158a17fe5ff09069fb8c480f85a0516b23f7b9c8a35d2484a519bfcb4892c3c3a34368f15622
z3256fdf0578bd3e639b2074d15161f0380439200b16fa52c751696404a3a18cfc9cf7fb537840d
z788be9d20e418fdd7000d7fa59c35af429ba264cd0f08b12d35907838001172424b4a9a3548e91
ze9e95de9725b80c69b891e24c5df51a80479db245b138d024288feed8190aff11ad646b7fe7f4d
z988c6ba20d4da4d691f357c7d5b49f0eb070b01e5078e056358001acf492e225af847246a30e63
z3fec57ee7a01abad95b1e01f43b099b32bd03da578751dba906eaf9242a26554acb06c19e7cc7c
zc50515a547dbb1bc2a0a39dabf49cc689dfff838532d395b8a0c058bd7097f8c801758d8cc19cd
zbbd9907f08e0d7428f833aaaf4f3038ff36c7be29080b20a7f0ba727633462ac50477ea5b0f62d
z9d52b2a54ae01cb9c1f004e58945c3c8be105f30e14d99fe6ee4e88782622da3420936c4dbb330
z4c0e1bbe5d71d3e0a851c8ff696cb9a7ba5a5a759592cff9fdf0ac5fa3e3f014a93f05da3a4a2d
za4f1662322f2724c70b7fd92babe174b3c35c6b8cb50d1568804f4ab24fa24055cd7050848eefd
zfde78fd99aaaa4cb47e6bb5e766036f68d01efc872b25183865b4c47ad326080100c33fd255bcb
z608bdeb791d2ba34aa89933fed840a48fbe27376ff2b2d345940f9e0dc5840387cd3bc36baf2ac
zccda2f7ae6c184e4c67032c31259545e11287ac8f995cc92da8226d1b314d33c776174c0406be6
zd65ca5ac072653cdc7640528cfc5cabd57910afad0a4582388651e05e491e4bdf300b727942d54
z503030f2a334049e890ccf5d27baa595b626f62f602839e24f5418f582468825cb18bd03df0464
zb6502ba80ef10e3c13bb01baf6a02f2da26ecd401603a329fbc865726cbe97598d9b41581111e6
z7df3055b198cdf64e75540c14ca6f61bff1cc9a5f750ea735295ebb696b30ef87d0573850d9605
zcc09d4cb097bd6936c9c0819b092d9a4214676a766b5902009261374262c96e57c77630edb4eca
z0cd9e5e9f410ee7df52ffbdc439844daa80221320189db8d13630dda6b64845afd4ca4ed4d8498
zda1731595bd7191471945724b6d00a97964c41da63763e2275c49bb82ff7679207e98bdee772f7
zd3bb09a4d982cf210ee23596e6b0e3de2eabcbe24d0b894f78305bcf94e19671726faa5612c89a
z12fe46ac3bb1d70adc4d17e2e424c3ece1a890c32ef24ffe82b4169065761c33b68ba002767b5b
z5065300a579232570b02a6431737d50cb60cb1b5abe18b07ac82dd16c668a02592fa072eb446b5
ze4916aad009f602a28a1a97e38869b3e8eb526daa32a8d5a5db4927e52b5384863a5659bcd1749
zddd05675c37393198f94cfb11e8054e081fe01c4b0f44270ff874877ddfc41d6513f7ba6b3ccb8
z216431a12667f8231fa167f568e997d7387ce3493d4bb90aae4909e7b1d539a0057259297d4f15
zb9b3389703273e1e1d43acb549f5a22546536a147599e477b8098e704cbd2977e7b049dc3f3302
z1e086bd7d421c18ddc2cdfcdeb6e357fefa07718cd0b76877f3966e9ab9860101ee7923a93f5e9
z35196e8931a275dd41e6e24336c382f604b09d7c1f578f304160811799220f11f1bfdd53b8f3e3
z6b510c5a5bc00b62f636c3a4b87b33e93b2bcbb1f187b3ca4c8ca83e9f8a0513ee6eeeb301e864
z257420de184ed744d8b5162c76a804c5505480b7c8effb1f4edd1eb165252e39e7b9233237b742
z3ee7f57b04af4af21820ebf75ccb87b6ea12ffa63a1c44987a08bf4c8fd8bfcb54176f58bfad2a
z11238e612892697d8671806bb55d76de4b818cb94c61591413f332f4a0db5d518617ca35aaaeef
zec57c4e20f4ec617e6f7f503c0877d046373e6e59b9452768fc98f116e4f50c330fd5cbc0f9a5d
z90efd658026d84c34ad37ee3b9074cca22299c5658f6a6fe3ec4d4c5677db736ed142c94c0e429
zf8787eda1c28bfdee188e7cd04a5c74431331464770bf330f09477684d383cd1d5d43be3e81440
z0128af425327af1253b149ea1ad1e6493c4ae5dce8fb98c6b75dc0f3fbc1c83686cfb6533304cf
zbc679a35269d9b8a4ed608a17d8c1a812af807b8d775aa1356088bfdc490d6430f87f6bfac4bdc
zbca38ac8011e0837833f21972e364d52633a06ccafe26753ecd3d77e723995ee690374865300d7
z6573bd04064c6cb0e8a94e79042240ad86ee1e6d18413eb3ad066a9080b49ec450d5511a2c9e2b
za3a873671ac6b9fc85ef4292e74b802bef0bf36e44b1590b98a34bb8cf9a146fd316006a11cda6
z4d8ad71c6c873021adeaad548f39f8e7fea03cf466565b42e7d7efa1d877f2e06fae785c209b5d
z95980e958e0bbdfb086fbe810ce16b6396e9b79d07464b7d5723b90b479edbe2a4ffeac3c2460d
z506b0190a912393748086be3165fb8475d451edd5c18ea890780ba5b15dce1975723f1b4e588e0
z68b4734feac6b867f435bc9a89c7b3bea25d0621bab315d827cd59ad498f9bb3940d1ce559c7f9
z0524ee6a2e20c5c6af25882ae73b1715e6371706b939d44d777054a0f6bcac493d9e77ebeaffea
zf4bb998b856712ab8d6f5d72483c5c023fc0c1a553ffdd3948a222bd8a75924bdf0a44c9ed251e
z1e1a021b982efcbc22905584f791ff2005e72eefcc7ed4c126d91528261608c3901215d63c7b5f
z34a1a995fac7d0465cea35e73526c7b345bd7d3fbf2271b720c9fd12a09be4e0e1f61c7d8d2c6c
z2dd3aa0e4852d14e3c8c9ed84306a5690ddb0d9ff446866ea57ed112d52a3fb72851cfc14424ac
z8f9d13d2a4437441c57a9217dcd71ccdf9bee9a00bb7d8fad051e974452b159a50d2df2339789b
ze198fc0f7211b0db572d4f9852fe80c97a4de230978ad556d51673b27ebcff8b5b49618858edd6
z8d7311952ad0c227b855f12d2e6a1505fcc7171a90a11b8470d066c1bb2a2cb8a314a8c4a42248
z40feece844d6e8ace5b8374537a6ea377ee347208153c0a923b5d261e3a27e5e1fb026add7f207
z197589a39d37e3b7307a16a2af8d752a99721b3c8d310e9304d1c859f2ea954906e25da37ded23
zb00464cabefd13d85baf8f4a7ff590adfbcfb39be3b5827907eb90fbe85c779e1c4d36b8a4fc71
z70890092798b31fbdba7bb6c29a52a29a454d90b02e190c2536994d52404c47c0ae573d882df12
z9d31b2f84b3f69a9036deca5df6a7f7e407bc78016d8fe14af839a48e24b13deb08562b2332e5d
zb3611491b5f8e0e16b261e10479e7bf3640d5508e9b84044c19e4b2f0126b5e311fe484319f8a0
z686703466b5c6db5065ee4b5dc710530bfe36d478482fdb485fb803e54bbf948ddd03654436172
z5b130a19502cb1f7a9ee338e5e0fa3759953e4655e497f7ee07a9084ed7e67f337dd97dbe7c50c
z3d4be2cc65d3996abc50a0eabca6f1cfb11af3fd2d9353436c39f17ae6ab57318a5b1938eab5ca
za18764bdeb80d57344fb27339b81b69abaf58f92b369d4238dceb318130ce217e8f8a0e14f334a
z9259d30a6424bfe37189fe88b4d9c5fd0bf8d808ca8a8083f4dbcc0ce48d59a8937139a2db752f
z884668babb2ded65db4bf6d4515be22df60d83a3a5e46120ddc2503346c181a4228242c2d259a6
z3bcdaa5786aa29f4c754df426904bcc2d8ef0e69bd52f3a41355708a4cd3754c6e7d4a7fe2947d
za7217b6ee811f1e793802f74c953c90402bbf9f44bf205ea2f6ba1f427f7f39866a9d3e9cdc49e
zeb62d432c6db17a53a9f3f053733a547ef4c5510bb817b506faa01bedf64a0006f03b9cda3398c
z173c5f500187a10477e8718552911297861a4621c02b5f3da9bff4d4a1732403d8b09bf8371691
z4f42eda8f7c10da7e72eca7cb3b635473a8da5d31185cf4e3522560956ff81fc474fdf90a8e2a0
z68c14bd7a3dea9390cf09686ca4f9b8738cab78169e1923829172d13818cf0c954084d41ce9e2f
z17990f6e94307b37484fe142caec5bbd0012130a3dceb7b41faa1936decbde7aceed6b928d7eb8
za2e1c5590efcc69e7d44a35c21c13e13a3789783187a4b32c5672da6cf8b48462334b2088ce341
zaf00ed425b34eb14002a60a6cb3ea192b3a3ece0b28272fefc6bc17b8def1c47975ae7108074f9
z3bccd284c96ca73bf883f294cae5d804f3e9ac4eeaf47ec099e8c0a57fd30b79e4947363957c2c
z28ed49e4eb7097b79aada93f3e2e7c227f7d658dac481e6b235917598939fa0a42fc97e0d5e0f4
zd9564f2e96200632e4ad3c0e0a5fa0a1e3400e028ae7152fa4419e8f79529e63375ab168f61949
zb49c7d8a8b1d2234cbe303252d8f6aa55910328ab684508fb806ef83aa98f4cdb5ebabeb4979eb
z72457a2f2810e67daaa0cdefb6e9c7459bf29e74a2143326a66c2981307cc8b04ebe9c7483fd5c
zd34a42527c602150b182838b84c2e33b9d5ad3afc7603232ca0737c77505ab83513d3501a070c4
z3129594c4369b66d6c922fb841c21d44737f29ee7d57e3785e98a1fa72448aa2ad72830da82778
z2a0ef67d08c01ffdd3bbaa88f2d32c1962966a1389a4e4c365a7fb2d3778e69a9a27e5ad90ccd7
z2afa83e30c65ba4eb940d02ebe248fe43e1da0ab6818dd15c8be90964bd1e135827e55a12429eb
z9b48814dc0523b9a703389e6cb6797fcb20b872cec8fa6f32b421302635bd761f73781bc9d2881
zeec3ce25965229876d0a171bb0210f6219ace59b72cc1da746093aacabd1b6d58913fc03ed92f7
z96dc5b4e72457ac20241c9bfa42045613187b93b2eee204eef567931767ceb77461545af7ef3fe
z85a2e0d4b400fb8f0e83ae1fff778fd80de5feaab8d077f895c68325814989ca3cb8be1c806a50
zfe03b72e63570dcb4b551eb50e7ffb4683bce6051325348ed719c70e8778dce487c8fc7984bf53
z3734addcfc20dbc894f37d259eba852439b566033d1f6d79ca568def057b7031c0edb5ffa3a255
z61ba82cf12d5ba96ac9db38e7b87d8373aeea664684126262f0b0d05c5f405fb9f27bbecc3581c
z8ce90a850e03acc63ed7a5865b2cfad4ed2494b60280852b47f1e2ee37c8a7cf5bde22d747c997
zf33276a537aa66aa619457be79d1bdd7726620914d18b3e724ebb5ee52508465e5002d6e1cf16a
zff1849a33fe890749558574dd905c13af85b1f2c39949ef84ee706cf5d1aa3186728663cfe78bf
z6231ac5d1b7baabc0fbc17d35984d2253593f15894583807d10a680f538562a8ddf738764af440
z15949c662d44b4eadf9b84755e2b5071c58874ddac64bc6c4810bc138f2f4b3eab7d55d6148ee5
z66bf3097f4f6484b4de4ff0ae6f7835807374b83c062390a257d241d508b07bfbd465efc0d0e1d
z30adb1d5d8371f661110d02f6c011a7a1756132e6afd5a9d3e2a2c6588762c82e3f22381b5f77b
z2d826b1d9e2563348437440108a3a86667554b44b40d93fcd58826b59a43172f3c7cecfae881d7
zf3f56d95f4610a62bd7d4b83f9e4a10d49e312b050269607b145b1f03bdc5310d420cd21d41e85
za4f099e278faf05e428bd92191fead6aa161e2527e9db0685f657112a4eecdf16efc18e0083ce7
z2128711d53be7883b9bf024763cd6c9f4974fa12281a49f7e3ad32830e5cec90e1b0e3cef28af0
z182eba48fcc366e307e3ac4cda593adde7f7a08cb779a508e559b5097bc4c27e04005b3e4cfe2c
z31aedd0dab2ab716696da6780a472c8252abe15873681a58ceb2bfe87f6c9be4311b7f6824a66c
z6d22b85b8815081451e659136aa13a8532f90d8e9af98463850cdce5d3166619459f5ef5ae3866
z477c78fe815f6f643504a81a2cc943b054afb80e8c9345da8c1be1ce3869ef77e0fdc96c899145
zfc958e1d1c6dbb21b7c60d8824e8c5fe1b6d7575c53cd8777677eaa8c11d0a9b07a5776a2b6cea
zd5b205a59678032c7975128d0e9a0f9b5a5bd5bc9043664854eb91e1255f56ba522d257cce3743
zfe59a7a680f65b9b23140b87bbfd275277e9ed6b32ccbc4c176a3dd3cce9d8b9908c096fec016d
zedd582ae7cb657d9908dbeea9190fd9898b05eba78cf21f5d5ab36b095382fe459f65d091781fa
z86a01d02ea1f58218b76dfa3a4c7a789c5ef1a44fe227a97613881b076452f8009c64031593d9e
z2085d80dcc2800a79d1f3f8ce0e4d09f205b5ec86d8b30e21e55dafca25c5114af9fd97feb80d1
z64cb784abe39e0cbd5b81d0855c725f9e636b89a41a61061e5e8ecada1c4360bff4b747d47c208
zf0d2dc467e368fd4ec3c761c6bc9ee16234c5dc66b7aceb6fc686769f3e675c15c78c1b61f4f94
z0aa4eec8b04affdbee127d6983adc33f59115cc5d4991656c820b4190b75d5d80b048a69e12480
z7b9d9ba317eb0f5a55d84d18de2433c079024272629198d9615f1e965733b2c665a495ba64e8c1
z961bb25b1bc21aa45d0b1b67281737de96e73eac5a0d1ba9ea4bddf933872292e79bca77afd70f
zdbdba2f8f5310b236bb19712b6b6beaebf6c31a5e2be78a4e4cfe298fb7c5744e08ebd74b9cde9
z1098d20ce9a0f3153961b8a7fc25ee0f604cb71bd2263af24aeb92b917e9b35e8a751ce3e2cf67
zbed9f24a8425003321b001040149f6df4017ec6eaee25e5d6ac1f8fc0b947bfe49d9023662fa8f
z01da0c729e26cc55670909fd1d4daaeee92b08bf0d79ac711d96ab90a40caaf4543cb0faf1fd28
z80ad2633c3a3e938348478b6340f8f947558bd115979c53cf01551be5383a5f2ff2d52c07ea60e
ze94ebcdae77e036cfb12b543cd4f0a028934db19f450064ae733a0cbbc7051049d3550454e7d0a
zef59619f875fbfab7bb14f6154f48d6715b7adff4679b16c3ce5b16de75b245789841ca9351b33
z2fb2b25009977aff7944a1a9c45068627493b8e57bdb276780c2972876f8d72d8642ac2a5c01eb
z4f3031582cc0b7d8f1bc20a7fbefde2600ae31d0755c1fc887661b22ec13fdc24fdafb2ac07fb8
z0484e3fc022a73a6038716aa56cedab82634b8e1856621beb5d2e421214ca1c54cfdb1b4c16882
z499bab595890c4415f93e890d36c46d33a820c138ddebbed19e882104a811a150b714c2bdeb128
ze24ae0cdbffd1a4e4e3b892d4f6707ff4381d182887379d7dfa4b7252fb4dbdb1900839c3bba5f
zb955c176a82a46806e236d7a772cf881af5b7b2345c3c8c69357451d27807c0b4d349b606f69f6
z5acf1ff6f8012777a24a959851c583a5ceab8e08351047288c3c9ff9f2098df2fc8acc02797722
z43d1b13500963682557a2a410e6eb856aa4ffd94e53c1b243c527eb103bbd7e99db758d691d932
z0477a7dcbcd2bd3e1cb41bca9c50373b80f811475c3a341280a339b59d3a1fa3b57a7cf793d4a6
z471e1eb9a0977c45c0e3d8fff75c1eab749309cc1f7bde4fd3febea6fba050d888b573a1df3485
z1cb350eaff8bbe7cabe0a5c7c233501e936d20064a53787c5c81cc0c651ee5ac574ae1335e5e38
z863673f9d448fdfa9bccf91884720c9cc4a7077d9da84f44a7fd6b9f32897941f52135d117966f
zc8de021f2ef9808db6d2ee7f4830a0d1873197753373067ae552e012272aab4e9471029ac59dca
z48a6e88971b475552f2e46268c35f041615d0dc1cc4145959669ee6437a9840f1af114f3ea504f
z772626aeccc266435a8966bbdf333c8626f2cbddbd8201065112ca0f052fa27528c06b2e8446c9
z2183183f098860a38b3131ed09e827d06cb5f68b1220fb1131a10f1e61bf1479591ae4741c21db
zf354dc92c59803d14246d71a3b66af68e217a1097adf358ed9149ff07db8f8cac05a5d3b5e92f0
zcfea0c593ba22d4d8ec88eac08f19d48219522a73cebfd839724634b4b0b8d2ecd14264c547437
z3f55e08d950b4e0506f395f3a60caa81a22329b5a4578c8435e16b95821763d22031494e70365a
z096c0f57c787a8e6c3ab50a3deec4d961f657e49d2167954cc7387b1e1a93a76294b1b7206cf36
zcaef41a17c64672726f9123af0a80adc92ad581bf93423be459b4521191114c900312953d4d0c8
zbdeaed3f0d24b15759ea896cc0c37d5f2e9c6cfd48400a763debc13343ff5a6b1283816e420c6a
zc8cf0207ca1ae7cbe140c2f9a4ea674c1face5f0ff9af09f3e5a535b1b350922c3acd4e27f8384
z1c8c2fa92ec18f3ea331ef214b8243aaa01e049b73c68d2b7a6e09ef615251375a69240a509d56
zbd08c0610f94f1abed35495e136eaa052d6c8580d8fa7e0c8d0d0fade0716aa453a46558bf7855
zd159d0681a219168b2e74382fbee8836277fbd2c9cc15c49fc9ccdae288bc55b3db6007a38db03
z70910c3730b8e3a40497315c7876980bcdd6dc4647c930261ceae579b2dbf278ca34efe24515ed
z5a85bdc1ae94ad2701a83dda9f59845e12384f8a634632476ae6072ad187fac4c25f0349a90fca
z67474544876212e0396efd5423b9e8fa8328165440a5293dcbc1f0a8eaaeb049c95eb0bdab7773
zff11b0154bab0062c7d3e05a0dd8e1b4f050f88122e788a49e89ba77bfa728240b032c0db4c2f6
zeccddf5c423bb1cae576b34523e01b1699c39d8cfcba6e584edd82ef53443f39b4f58b3da65c18
z384d7e8e713dc4f5e3a7fe81b63b47fe348a02a7132d9f79bb7f7ec1ead120ccbe770a17bccdd8
zf34f46ad2fa76afb70cd3b5965ee4fa73602bd9566147d664068871c35b5853f0a2163c6dc3ce1
z7679105d07f0655733f65e00122b9800cfa734dac3d56740b904214405ed16d0102a39fda00031
zc21dc0f0619a022087ebe3b19141cb42d6e2ab6381db7a1327a2f971b99e0f5e6a90f259c0ae31
zd43699ffae1d017ff2313ee5b48ff9e4fd8944fa98a3a7ce82bdf94115e7078aefbf129d76e543
zc087a2615f495e2846ec33d912d1a8412aa90b0edcca3c93def3c4cb87519883168cadff3ef2d3
z3cb492d38ad01bcddb57538a3e2e79d6b3e8cfa1c8c8fc35591756ecbcee77f66ec4fdb0a0d072
z31fa60828d303eec08f22e9217e35b72c250f77b7b9817290b99771f4c1e6d08d50d3f3fa927f0
z397b1c90b1d196ed17a4dff9779d211990754525a0f2c23dfcdf2a33c136e177343701af784d83
zf84942558f63d9d1fb92c88f23f4eb963052ef2188568ea55049efddfe99cda8fbc551158a77ed
z911ded83685e428d5c95ca8a6441efb9dcec7ff82dee9c6a105a8f46152cc5a9dc745f4af86687
z0075de353bc4261580d76684c0fe20ba7ec4cdc4aeaf9ac09e17982824c6aabfc4c49bd7b7340e
z5e588f83c7b38c4f639ce7c2a2b2009a1f83cec68fdfac79cd5d9873a9f19c443a6650a7f8b680
za1a6133b2147a8fc7d394fec3d9fc14e8c14ec1714c7611122a88c7a0bc1ac790383258ba9298f
z0b5762e4222238691fc854896c3365ff87235a0f786687f3b6861296e55185bbf4ebd299400de9
za7168789edc55df0f651c7ec48da87f4e58858dcec992d84747725d2f657fc419e7a1e21e874ab
z1aed1c7dfd4834f8ebb9b4842e090a2c328d731cb07d8a2ac2b3099bc0434e223ba24568909156
z5545e405b7cf66616220a1b9205ffede90c97601d140ec5713f0645e9300c51f36cc2bf4623719
zbe170bfd455eb10754459a32052da35bfc032a351aba561565ac8a4aaf0c131a2573e35eeb720f
z71a4689047d23d405eab225dd9d279f693eb3ccafc3536e94c8fbad3020b966cea8b3546eb97a0
z7cd57ce592babe0ea09aff73b5b165bfd6b974411bfb9a0b857bf44aeac787c0fb453980249c81
zeace2b5a17dec076757796834dac9d8dcdac39b8d158f8b04129bd88a75422397eeea4be27e517
z2a645fd81d41cb7499a08e27a6cbe1151454f495c7b46ac55711e0ca952785ae8423f96efea481
z62fe334dca879fd826673a7fd4f642590088b73b99b3a47146983dc8e96ecd484f4289e8b59847
z83ee21adfcc46bd3c4a2e08200fbc3b7f443aa37d93a054c798490a788bc4bfa3e80233eb31c6f
z24146c3570daf7c4549506ce93f3e89a99fb094f2df7fcb825c33afa8f852698ac513d849d1598
z1419549f6cb9f1d04f3d4fcd4e860aaeb8b2a80dcb8b98fc2cd0cc94559808007a860afb3c945c
ze2e3a8826d502a6b1717713587df2dee5d956b097a268396772a09a9092d4916ae2bb35b7c6db4
ze69c9a74ef502dc000418df8516d79104e7d297d8a64b38063439fff8d46b818a745e49d197011
z5ef664b66f21fcb18698ac4416ec15d1e676598a596113d709a9a522679f9d4968858c67953c4d
z23a396a278bd164b6f77cecc5c72f97f2da501bbe3c057a60e227b75ca911aa7ecdc2aa9503d40
z5b9c7475333fea2201be09ac87ec0f49ad74a9ef9e5a2b5c3540a59a6ed7d6e24fc0b9f45091ee
zcca5960d49c6f6e9fcc9ad5e204bb8e65266512b0d4964353ba70ecff4647c34342e13f2cce3b2
z5e51bcf33125baf6baa1d60b4bc703f026565f03b423294848c242732d605057bef8daa4b60b71
zb5a9d3cdd20ee8facce996f9f45ff82f8135e311e821f8a0db9a5de30f008458051895134e7c50
z4ac56eef4ff1056c7d88673991519bd44f93177b772b1d84c0962d64a303282a1fde4d76bf93ec
za7b53f5a59bda0334eefcd954b8f3ea175e7ce6c36873bd167cb0a4c16ac5193b46006356fbcf0
zc3577e062cbc86496a81b99af697896d819337d151f9fabf8d5bb19d49c2b6bd5e961d82ac5915
z7d6a4fba1f468d5a34b0a6f623e6c62d2f5ef951dbf4fc23bfd00fcd91d099a5c21e879c780b5f
z70a6ca8df6dab9c083678763ac2577637c86bd3864f3574dd17228ed419d0eba5b84191a767b96
z38b2351085a148bc242568bd2d9e3efccc7ca826f20e1c919d9d562c98adfc2d93f53a89416f05
z293d356b0f3078370a8461d8ae9b6da855181573869522726668ae90adb91077ba24ab3877289f
z606557f0ad3cc1e435d40a20170c1aa30c54ce4e2354a4a57dbb7f45f3c5ff3851de3f9200dc44
z72a8baf32137017a8189a40c4110659bb1a83a6b79918f84fa0b3fd2c802b2f7c6e2a3e1c684f4
z5bc131cf4ebe42502ca6feae8034b49feddcd359973de624c0bc0fc4c8c84167a7eefee441f23d
z23d03422cf6e10458e51bff36d8ca34538ded21bbf40da941489cab32f75180e3cafd775929e8c
z76556382c0bd32504123db84a6f0c27e27c87e638bce434294359cf7e27cd7c2c4947082d261a0
zf9dd87281e65133a2e0b000cc2d5a1ca81e1331d1cf8e296dcd258a41a44db31ec3289ff104749
zd53c4d82ff9c06f75338654a810dcc42b963e68b4d78bcf370e56f45d94fc678d084948b8ed9ef
z7e2aec7582d655b6bde69db75bb471c6275cac0dc31f7e14b846c47ccc8824ac1196ff4c6f23b0
z507f74adf4b4bee4e64bc778a371df11168a630bfd6056cf986cea9905cc53f7c079d55fcde620
z3fc54879ded220832e002509216c02af563d76c772ed6f9752202e47844e4cf26e76b93463bd1b
zaca5ba9472ed324d3d75609d5eec82b547a6ff8c5467efbcefec5d4067dcb447425bc13b74243e
ze89258bbe18c53fef4a94bf269eb0239937f61a3e3bae1a6a5db3348ef4da70fe4b6b77e87e596
zc98eca9a771d8cffd61496e0f9dad65aee805a2fc121cce8c8b704e5d9316f0a55f6574c5ff591
zd1aaf68e540f51896e41bfa07775fa8cd5f1a158eca559ca6ce0f4d111feb4c9902c0c03bbf412
z0b0cf7ff4d0a86c39071a33371d6a18222dc2b14a1009682cfd3b127ba5af852f0fe28dc679f61
zb9554c829bc8e711119533d1ce498c34ab2334fd40f47ac11538109d8845ea90ab0b580ba48361
z837a57f6477c6fd0141d3210acaa9dc50f819b38ff20c77d50a96ac1779f5fac1d6bcd3a4766d3
z14a4b28c943bf58a3c94d80064256478ae3f4cc62f6e8c6d5dde5a1f7d3ae9b568491dbe39913f
zdefb6cc1f418f7f0ac24b51054a4143904c7a3c45109a1f60fb16936e6c855f3a716f380a48824
zdef85daa2d36c04e28302c7e842b8266dc23e9616eff835be5aebd81801bf931cea9e0c3183c18
zde018f0d50740d75bbc4b250249b997accd791b9044618c0b7161a48f5b53a47486fa5fe33d576
z54a981ec9265288170400715944472bba800619a76233df8fb3d7a134c98b97cdda02b38ca559b
z9ff646fca9a40603597493019e739e1f1aed62adb21734607243f15bc1fa0d42e60db123a0446a
z9a9d4db5d217e4f267dc87edea75ea77e394ba084b2d0265d5f8cd7a2369657550d009de2d406a
z2f0f34df338282f113eb44e14a9c635a7297c821fded7b5f0555d3c99a298bcdf9fa7571ed2ebe
z3e998c6930b3d2daf523c47c4e6f6f125c59fb9872a6ce7dafcdcd7daf43a0b4a8c1d42098d99c
zdd36cde197280fc106c57f318cac3c0518739c1c937d50f35733fd09d3bc0d9c528119f57b6d86
z8636629a0e4ddae13ff5638cedea700d188de8bb7629908e1005a51b7d3b39cdcce15640f2f737
zfefba7b216f17d46c58d1ab23c747430af65237cbb9675b974a376563242a4130644cc4165f6b2
zd6c0c3db5ebca7ce6a972b8d73892b4fd749a2faccb882f93932e76d4323022c781f5bae8df8df
z817ef635a3c680d47d6c305964760a4b489ede12289940e85c74524d37ff9f68828b746e64e684
zd89bd7fb6a919be702b54d8c443ead73875f8a3d3966101c0a5df0dae9b0fa8a1d005fb7121662
zf0ad3eed8e214561b7539efba084f289f74ee62d8b988432e1d7a8d9f41ee3451d2d7cb0dbd98a
zd6e0bbed4605f9e8062b1870b379f67ce790f786a798a331810d213f55cca2cfae02ba3f278b53
zfb56d746c9f0fd9420163f6f9680613be795b90508dd8ae3c3df1a6c694100134cb7d58b88f279
zc0b6c22eb26c78205f30b5faf89cd3a323ec4fb7cdacb8d3742dbbb9a81a5bc865b8e5ed6332b9
zbec8ad24c571feb61fb1c0ee4aaf61f93af133bd847ab6e52a38a00bfe201fba0dfe5291307949
z36b8429395867a56c38e402dacb3cb27aa34a5586bedd8bdf5d79bd81b71a909e055568568481c
z18736d85715e7a9070c7d53473977f84cf90be8b4e0a4f9c190fdc806b2fbb774652b40058b27c
z9e57f750a938461688243afa3e2b48c452764c4e39f42a29ea914ac407102dd6ae416e32fa9d0b
z975350545bdc6dda5f21294b20d5eee474393b384fa71c84ccb4c49e53bb5b50395b35aa62a8e4
zf9ef7e2824695c6d060b5a55d97db707c03e5cef41f9058e44fc4bf3c09c168cb2f0e21b00b149
zf7c7e7ed6d46d079494f9575726850ae461382d3771555f646e167b2776698849aac6c251f457f
z4406a6f71ef34760d27173dadefd88cb93b100da2258003cbfa56fdfd7359d312abc0a8fd0ca54
z779a6458e7b53a97804e67f29f30da31279562b9f11b41b33666053d8b0cbfd419f44f34e00431
z323d45d5e6789cac51813dfdb2d4bab1729aea7c1fe021b1dfd7e25a0ea5f6d9b73777c1cd407f
zddb4b070de8d3c9882e6c1c53ce5916d9fc1d8fdb9d3d9b75bbdf0b163da9c4de157a6bd1a88a6
zdee41bc6cbfd863b8555dacc1faa4f589440d82d8115342ae7d2e2cf8b7f1d076af0164cbdccc9
z97c61417111a8c14d081854d591696dd2d7c69767899235c6a4c597426f9d4d6126694ecd7048d
z198cdd38dfb85d34a48423727186e9e0876a2f4b32a7a5d1967110802454e0a3edadbb1275bece
zd41d6635d34f7ea1932ccc3590105a97c2c7b30e36ed048c5fe06472216b371cc332cc0e7b2eba
zcd95a3b1241aa4e819ac60b2e61e10a20e99cf417d947fa79389ab35276d7461b288252176862f
z4b9a4e4099f6225d708c70ccd40ccf6a6f0cf3203094e811552faeeb5dfe329b8765bb342f4894
z780e248c69639f9d8acec6f93392768a70b2ca0ef2f4bfed8a0335381652dce448c0badfa5c960
z02bdb642f3b1d9963d6fc85a27a48289e7e9c6f0bf2021bf05d7851c877ee97b207a63c834d2ec
zcfe498d2c7065528dbb64aafe49ea60c02420f38d98f548cbba8b8406f81f26f2c5da1380cc613
z8702e8cf9eae4d7cc84d0bcbf7d67ebde0bca7e67c62bc0dd4e42da599059143c1762c398bd4dd
z8267f69ff29bfba1443366e03f85d8d18e44ca0269df9f4f2ab9552f70dd8469de6364171d5769
z334fcb9e427a8444b369e0ab109bee3a6d86fb465fa32c723184fb2e270c378d0383dbf7964b3f
z607dcaf66b35204b76de9b0353cc06be3d165d0afd817797fb7d95f1b23253cc61f5fc88a5d684
zd199c28c9072336b96cddbbc5abae64fff3ebbfc57e1c2a0ad2bda1133af18a1b27f48c38b8222
z6ccc99d9c410f980b62039bbe4c88a70fc12b7d9a44287f27f56cb70401f72a656c468ce050812
z1a67162cb3fc024e70bdd53b4fbd20d92f972f9b1a6dde9bffc654fe5e56d0f7dd0fa382d5fedb
z43c21a26b4e4c72e1460af240689da3b3482fe6058c88e58a56317b89115be01f3f535c2c7ba0c
z6c786db01f79081edc8f69c45618859e19ef10067897c0bf8ebb53b350b960d3bf4d352c7ee516
z771542d9dd373ced34bc1800ae3bccc3b84b4e1e86999b3da9a73fe0bd052619df3adc3c12cf6c
z8aa33657fe05a7ed13be4215c0f19ad93be31d9082b712dc999e0e91dfb200881eec9a00a192c8
z07b888e63fcad43bc6a7020f5cd7747e7463c5b0a37c52c70caff7b7e71b9f8b2672d94e44dd7d
z8015574931383a3b64b3cb39e2b3d60c24ac0e311c9d5fbb93957185a1b9800252b1edf38a161c
z62fd5a2f248b372bd2f99761a6db3735989702885ad0071470a098e00583ff124d2aad7e6dda86
z22c3aa5b909a0dbbe04ecc7f2d1481c72fac734626491cb96b3630017ffcd0a94940f37de0f51c
z4f1960f9104dfcee4cb866b47e1bfb229382b6cc6ce70fdd8569f6eda7a7f3095144043fb4b548
z9f6bf308f2ae90901155db8b7c0eb9cd7ac660de7b64a27f0cf7e44d9c40e44958ff132fa9de6f
z46fb077ffd4e65122709d03f245c90af94fd1a65057561edd9916d8220aa8133aca74ae9ce3e93
z42f0e01afff77331cacea05838279cc726a7d7635840142a9c623eca91bffde9f4456184329fc0
z490875f3558c952df03d4eb1d707c71c36edac5d88b7e8fcbb990d326cec9c44fb59cb2054cbab
z05fdcce2e8805b2bd6715b506a38866ca0c53152e716fbf52d696806d80e1623ce992091a01f1b
zc19470842486c93cb1d1edde453d6a1cb30f2cbea4cbab53e0b4c114270a4927f83657e91ad3a2
za7c6a70ab8dbb72c0f0ed598a766f5d8687ad9b40b0516366a4a822a8391c2b82d01074bcd76cd
z278fe68b17fd7b692593568bb921d1105ed029af17161b72afdf9fa703ac5104befdcd26acad96
z86b9a67e4a50ff5b9ef5cbf4c219865ea99aa96f438837d95a98c4c0776885e57545bc005bd05c
z184ae62b34ba20f29c97adef3a69051f254fae0e174b30074dafceb531839549d3004ff51dfb5d
zf152d456f0456294c0fef5f09f69a1ecadea2451fd95bf3e07d5d08adb33cd9db93c59a74700ed
z35f3dbd8aa3a136b39237213554fc45f9e879e499dbcb22ec0c522e9437df8cea9242d58df50d8
zf4cc5c7f699b62fd521d76194eeee4562111800005102ce364674b2c9dbed6d4f7d47dbbae8509
zeed7f910122926f2cd0950eba4b1f3c35bbe1bc3e2498f8010c5aadaafae0ca16e9d8b7f820d49
z33a66570401599eb48497d1349110007d61d9687b85fd266c53268ec69b39545e629854c36eabc
z617362966d742ed369276594bdef6371c48e521bf1de99db49c7fa1c73a717f9a3d9793df6ad47
z42e35d7dd8d440a0cabd2408a20b35e050102869b50650bfc43fa6ba8af32bff605e9c42d1db3c
z7db6095875a788e709a1e452755a65fe29bcf47332adadb8e9d3e16b5576665c9fbdc0211dc6d2
zefc31f52fc14b02d889fde4c097c03df7da8d2ea567ee059d27c90e883be9ee559c4caeebecceb
z82585cbfcb461b36860469d7ae362cc67630100b3572e934e842d91a14ccf7f9efc0de9dfbb61f
z84ea45d3614e4e9d1dbb9a01b10a96b0b383044d20715bac57f1db270268369dc2869ae931979d
zfa8fd606688d4bdd9c8bd2106ac49ae9d0bd5d818d1b38e1e891aed081a60111a1d29cdd0a2045
z11e84cbbcf182d1e8bc8c399ba2ad43b7d4429a7f4040be6079c971bdb03074ac8e84eba6fd312
zdd05075e556f4424ecd501b03774f8e7ef860f7bafa83b490538a32ae42e0d37c265c42b3a0a59
z307f6e4f056afc318258102156e78bc9405a6044b28a513c0d19a1e6cb59085e7823b3be183dc9
z9a31175b945e05d7ef3cb09036afbdf7872920877f40383556aa8e4fd7a22a1f9b10332fd8b3f4
z305faa89d2ae7d919ca9f3113606fcd46accbe0dcd19c1dfa2ee88700cc41a2faa4c2897581e1e
zc05d106ba1165c260a27a7a7082e4041961c14f89b10bdee6fc6249e3f2ac9228341e7ef580a3a
z2b615701d94e56e5d16179ff7b78faaccf85aec1aac5e456853c8741fa90469501b9b783b5b114
zf5a80d2b2a33b69a188466fa265d569c703957a975a88e056e040f5007da1d3df5189be06962d4
z7d15c5ff742a934157a4b6775b2056ace7d98290b3ac26b15360d489a89518146fd48522132618
z2f1569c89556865b4739e66e91e01ebda5a624b680fef53c6d2e3650c6611df6330fd0db6c376e
z2253f1d5dc00a16027bd1dcd8cdf25e862226f6bde26e94bdf57874edf98bb6393a51e2dde4a32
zfe0254dcd0d702074d232aeab3182ad914063ee4a6fbcbd87946b0301e84d9c24d09c1800db70b
z0b1afb5bed45c9e261194172db21ddb3429da8362fc417fa2e31361bb15ca8e0597de2877ae0c1
zf2cc393e41a5f3b2138cf1e92b84d9e662b6e3c2a07ceb17c4f9be4870e6fec1ce5a32228917e5
z38f3950eacf63af5a0a25fef7bdc6210782bd49fcf33d593c1f40df42c4b450ce4b7cc740c087d
z8e2bb59caf772e4674a9235d634f1009f30dfe8903a1f923c027eea65b42f594a6009fab15d910
z4232e64d487f4bf46b2419630daf605e7910162598fe0adad54c1bea09143beff916903e54dc6a
z4205b32a3bf00804ca6000fc95234c03ca18b729442267d03e401df874faee8967a71369be5c16
z8f3af45625e319cf0613a10ea623542aed3241e6c69c78e5c583f294d5fe1c414ae8ca83106f9b
z1b0d720a0a0656952cd8e7a2d4e679078e578cfd38a76615f16278c3196b56de981a2e1f9ed8d9
zb61dc907365e5040a136acd00fc8ddbad83239f2fe1f141b36a204e1f13d5424b7ee5849ba86f0
z423c29dd27a686a4d3ff77e5a895860414bee48d612976f659e526e73d01d4733ebe2d4c9dbea7
zb1769c81ed7969188d24aac35dcead6a7116d51f6ff5eba312dc2a8db6296040802bb18816c309
zbc3eba4a9f1d9e9ac4c5b2b80390bb97db6e5831e9e105bde2205b6e85798418c89de107f9f004
zcbcbf47de789620ae6dfd49e750d36056bb6fea9759637750089f2bb5a065760f19968c1adcbaa
z30a057536cfb442ccb7e78d7e9c4120ef92a3f18af30fc7fb2c5d4d757c91ce395ec82d68b85d2
z464d8334815f64fbc93be976e0994de44ebbecd851962921b4b3e76168f70886abaa353ede13c3
z455fb5f1139c349191b106b34aedc8527da2d6d02eceaac8b28b8bc02d90f60cb31d585b154561
z65832fe8a422c8bc7ab6451993ae549eae7879616f3070df32f47ad915f6d57e290a17d3973c2f
z35f7c0d980c40cf5a700b1d9a9cd98aedc5e6eae8a11a233c4efbe6d770a57bf84c480f482b31a
z4390a4325afeb2c027e200e17a6878ceddd05202edfc49029fb54a54d62e93e07d174fe71af71d
z371d7495fbcfc0e90de7386c172e17d31fc3264aadbb92f3e3470a06877e26d84201431d97ef95
z97ac3880d9643bc4b10cdeb273a13a7a9f87530a3da8b73211655a4600a4fc1564701d7da4dcc8
z0e65fa5c824b704aab8e07a9bdb0f6c197059740570bdc2b93f4dffe830680b47c0d0363d0c88d
z0e51328bdaa8ec74f932bc866c1a90a3c75dcabb7955602f8348972cc243e676ecfda10e0e2b95
z7aeb31136fc852e1f81e9393058796cae14987555cc21b345f848dfeb43da30b3b9e35a3fd5f05
z0cbbdfad37b6d696560ef284649c15c93e574035a75a1c46af43f6be5c0d632336bf4a5621228e
z0586eaadfbebcd8f27e72fc717d23cb0d2cb7e9b01982578bed1846e5d0f2ce24308ad2438e724
zcc1490ea27fbcd3d602285392404a82e19d2b8f4ed70194c5b3070eea366d19670bb0e53e3b04f
z97d01ae14e21af70155ef5fc3b0b11efb9eb263c48e8dfaefe26fe6c247a9a583b6cc6928bb810
z868d6da176ed85a48414b870e4be1763cb28f0b836a4d9ceef0dd8910343b3d7cbf1c4a3cbdeb5
z23c788954a410f81294751f87f501d87eb3beafe3792c9ab0093c39ddf25a4fd6a839b41b1f528
z888aed524f8d62e63797b4c1f7a9236f5141571ff737037c91c7fcf7f6989a1646385cda1dc74b
z7a876c69c091d3658ef1586b0ff2d285127c38c8484ce507033d97d83cb3c0f15b0c50b6ed6dea
za1651c42291e5eccdb34650c76512ffc5dc4c67b4c1b4756dd7a0bc70aadc45339106cbe0197ed
z68e409cca00f699bc2109766014e8a7697339489d82e581c60d08ad0defcf4c6861089807e446c
z8da81f92a785a1d09b68931a1de1b1f8d620609842f82304b887de53603962743600489926ada9
z53df014a047bc360ca6e7bbd5f6b9668028b73f456570763a24457e95d75ea682d1dae9c3b3b85
ze97633e0b7187ce0389b2c803d770cccb4a944a537818c519979758abcdc0a9c7928afe5b3c55c
z5da56146f27a3ef868e0a1258cfbe94ba34d7a7b3782ede9ad74e937a0dc76f834d0ddb5dd79a4
ze9a5229293eea741e17e4f101eb800344a8efe0b1808d91dd606ce8e211d3686b37de7464d110b
zbfa7bfd7f8f3a410365b2b53b52aa1e90a5015f3b69bbb34d439548c30fcc7a3b1667942e39b02
z19147f63688a201e6d7f12782a42785b55db8df6663caa4622d0f260bdf156417b6adaa6c4d6a0
z0f3d5b85a2064f9173ea8a7d0ca3aed4177cf467a251db11904e29992656eeeabcb754a73f622f
z6b1255d34a2bae524ff201e5091f20ae8f6828595df241638cd7f67b1b6166433a6b1d49af152c
z514699874c5cf83f8f729909d0120f5547986c525d18abd38304ad384236fd14b44fa230844318
z52ea46c13e8151ffba8888238b6bb84fc70106942e835eb6582a8f30764c80b7369cb31da90acc
ze3bac2723481fb8855261e59823eaf957c5dae6e89a82eea6fee5a7dcf69a3f2369e55b95824f1
zb18351c1ef674d3702c874c76d6f9fbbbe496d2315636c2d5f00d79db45c2bd02619e58235a4dd
zb29d4b5ada8d963113e7a4315ec76720c3faedec2b348083670e8c013296485ecf396cdbbf68dc
z0aeded93202db794fe02ca08c3bc269d103daf82ddf967227b878168e0b5e36c1c62048e7ac2ee
ze64cd5d3fcc3b2a2d1288264c031f571307cc596e6dcf69957f325062c7f918f861796f076fd09
z72f25ed3a577fe67bf40e6dfc65d8c327c0b1790a081c38648fe9e9e6219f51ffed4e33bfe428d
z4326e1dd38eb02669ea6d110bd0e64b7f8017c66d644bc398a85763dd25940ec8e302dd82bbc4a
zc2d6d589ed42a3c2f36ef812ea8e1d987d6df0fabfc6fa2f61eb63afbc66498ca5e4210214933c
z696b7f37151f1a222afc4a1638f0d7b8073a2de853952a6f46a8a40502505c6156edbc898d4183
zaa4bb641ce53aad05b062799baeec9d6b29889ce7c46457c4f0e9e1d0a24885c9a676032c63415
zb56a61de680733750731a8577de4088eccc5483f732e48bdbf0a46a711f3e113260208de8b6b0b
z1e196196dd35484f3dbbf9e4dacce4a3bb45f84e460a69c19552f4bde7ec0360b53748d172f043
z53325e2423b4ea3856fed78ea654ea3b1278dbf0a862298b8b99f468490369275b5a3fa87831d2
z72d34c10fd4e643acdd071bc23abb37fe69b1cdf8ac6c1e508ee6761aa55b35a60cfbea8d30677
zbee6211c98bde92a047a8a616ea944828d11118895ca928c3c5fde73e74593811b6436c18e7e99
zcef47e42c8f33c92b6c00a0498110664a6106f2620d6e9d301d615d261f320c13c0d394f274910
zed31604a5e646ec82ed5070a6be89f5a7c2b9393d95932a84875ec396cc7b5453cda84b631362c
z54633480bdf7f1981f44a618b126451c6573455df85ef02b1e77dccad0653be1b1c2b0fe4fc980
z895b49f99b859802257e81e5af38b48830db133d3ead25ef1da48e2f5ec23600b396a75c8bb354
z61cfd9c5755e8d84e41800976189e33929ae0e75033a0b6349b5dda3ec5a28a75266da7deebda2
zda65175ef1a4c11f6c64e5e480842e49a00ea9f91d989cb73ddf2154a25d9d5da15de3d3cb32b0
zec9066e8d065fe79920074994515b321e8844b3a5f5226772e41230f89d27fdf23a06b28da5c2a
z20fffad3bf25eccf239d49f67b34288153cc24202284629c6df100a546a15f8f09f953e907c8f9
z2cf6d960c574f0056c72bfb48f1f67c1f79c6ad8920dc05cb1c697c47c9eb8aa21338dfa3e42c4
z7bd2b8d1449ae47d7ea6b834fd7cb9e43b83264d580b48c2b6b692333ad70ffe51bcfb97dc03e9
zc3490ce8fc77a1d9a267e44c497522dd8657dc1894cac79d729c82f6a155c00956b590380524e0
z2d3195d27608d84bf6f2313b399f886e0176e8ac9a57278f5c4d5ab5aacdfe732f23bcf1711583
zf89cc618d69a2a18c12d4743e84745acf5d3555f59c34318189dcf996c572cf0ec0e9e937f9764
za3926ba206afa005b464d457a05efbb28c672837ee5c051e5d98b5cbd288e83fdece97e3373ba5
z7125bf5e3a0f1cc3f66f7280e47124d48f5961765981857630b7fd7e83510bbb1684e5fc6ba233
za6ffe17f69e856ff5e0a6d9de558a96b9cdd48251b4246eb3814738351fc3bf6544fc9ff43c0cc
z67e905e347b624cb3de631efadd3e9a7786a93d8e0e9f6bee606f9573bca12b39bd5f0467f62a2
z4a244974891aa528a51b967b0cb233cfa8cc2ad472b6aad62753019c278e62852f9c0178571d4f
z9f0ccbadc9ec70404689bb961e6c4afabd370ddc97b75a431c212234e3d8006e2865da42f65865
zcc60e63a287a243642b851e8db713b26ecf8efee0747dfd69f6d009837188becb1dc9c493d510f
zf05cdd5cf4735c436035aac47b955a3154feca15009f4572266afe86da84749ffea8879dd93bc7
zef0aa48a985c3fe69fc408e34b5e9aac6b1ec044f5a283191db7424fbbc6675ddec9e64aefc5bb
zba15ca8108aeebef2a8a4c2d7929c49b2544718a65d49986077a80f13956c72a536a491fdac340
z06defcfeb50490483737cdb1ebd84746af2c0cdc20af8e0a91684ce35de84b8d5e8bca58a3a91c
z74a0cb3a704ae79400b93db29eac7447f6d0eff8d78e9561a46a18e6a3607a38c8dded37fd8e06
z27fc9f047f6c75a56ef2693a7ce63fc47811121e4a8cd70d04a1d9dcf7ec6619746ba83a32c5b4
z889944ebf66481c018b26eb6490524fe0024ebda1bb3a1e743bf532aabcb2d4522de1c98d098d6
zecd20618fdb9de4c56caae726efe6f4385506ffdd71772f9aa286af8f61df0aeaf3bfbcaa14486
ze79bfd6258ab44e91e97bd9a9def8a0e51320cb1dd0d693901fdede148f49760321fde0b579705
z9f74423b3399fd9cc4c26a7d97fae26a2a0b4c49886975d612022721c5b4914a7cf453328e8e30
zb988343bd27ab0d74c04ef1a8faca8059155b5815e4590f46562300d98aaef814590183e8f2589
z8a9d87d6ee2fcfc83897ce82bf98886de3ec88adc45000b727557fff35f590b85f85996ae32366
zabbe8ba653e2635d9358ba1a5bfea47471ab55a28052de124a240fe0be6652ba441b87b35e92ec
ze0ed0c4769f0b39c37fdead88bdf85f39c4a3e924d548a622de502aaba158ae7e5a60f94b1f804
zbb7295314e2ee6d898f900b2ffb37ad3536d18a1e0b771af87e629e8ee67ebfd2dac394b63c194
z36e33515fae0beb886da76682809d1192a2920bb4241cf03daa21fd9cd48ac1933a2147fa43da6
z6b70284430a683f0bffcc0dbc5ac191de945edfb55ef37efcf8c635cc4633816166d14b34e60bc
zb7261ae0d2df0ef452ebf4026979cde614fda69df72a5ad25031f04071f4ff72f704905bf1d634
z158cf2b82fc4c8bac32737186abdb199e8cd3f99b07d26a9123c4f6a04a37f38da7a941d377adc
z6928517b80b340880b8f1f4ad018d8e1551ccc77b0bca7fde2d74eeb0802247a535bb0fa69e563
ze4ef68c09949fb2b7a647c1a72b71ae60546f36ec7b7d9a9cef2ae4d9f3c283efb91e2896aec01
z7564feba3d041d40800e62569c45d21f43c722f9a10fae69c802a6447acb7779c8024c2b83eceb
z06f2c22d02eb5f308a0349ffce1eb66df1283cf37ddd23e31a2c969513ca81545ab0143eacf92b
z6ce0fade8c13c46e4a3f8ca2f1ddecd536e00014a0647f6a73487988b371d428d4149018fb07de
z16e0bae98406db83f44f3f341e9134513154284281bad37a36a84c9e939841c8311a345aaa6d91
ze99ddf053ec7cf78c75e0b93a2ca07b243062d5c1b3dfc0a742809ea85352a45cb4d04ef305eef
z6dab8929c84d61149b3575245e82c9bfe248b13f4cf59aa032e380315fe6778e91f90e4f0bba16
z8477dcdef16fd0305bfbd68abbcb3f1c651805dd724cacbd8b28bb9ac61cc3959a5c7500aab166
zabd5916cc89224c64508c11aa018968e56647c69554eaf0687d6357717cc01d09b0a429abb8e92
z49213a5790667befb175c9114529c3e366ec73681a79bf98258c074edfdab5aa6772698a3656c5
za999c995e078bfbaac7da2e2095249a48708c41d71156048164d221923423bd644479c40949957
zd58f8d36e53c1c993211e9bd561e702faed44bf157cc6558efae8f98da541aac5baab588d91d90
z96a124bcb5a2b03f85919be955f9a85612b89aa82cdac2d40837c3ba8018ca67d5b89d217e4c6f
zeefc73b88653317bda7a417cd1bd8608fb6480428f391e6c088238079b938836dcb0d7b0fb7f5f
ze01520caeb3c5da527289b40a9f90f266ff63cb3aa1dec39bd399a5c47910a1b0c3f4a40ec9727
z69cb07b9c5d04807d9717493819bae7bca4398bbef5ad5314bfd779af822a1ed86276ecd111188
z79f0e05c5aeb6ad4492992dcf577b0b087ca2d73d45485533bd6b3325650c1a3bcfdfb84b72543
zdf7a7045fc7c8b13f8f4b2f77df73bc80a6ca7b06d62dfd7c30abf94215faea17ea5a7d9284209
zf02e1ad40dfe14613c5b96d226758f34d3d51dafba51cf42593235137e82b861b2bd6fae7d7c8a
zafe7416d55cc9d94475d39b31363a7a5f0f7f879da2dc3277377781b08a6a0cf029a50f943b1c2
zd390a4d77967933039e16d0500623b1509e6b6dbcbae7815dc9c106504851e4e209e1a736fa62a
za09149bd0217798c7cea007074abf03401cac5c9fe7497b8f9ecd1bd165a5fb2867cf1d7f98958
zbfb4df7158d0717f259081e0249a9934c29d7bc5e502aabac323dd23d3541d7f3c9950a5586bb8
z07cc0ff43675db52d7fc73cdffa223036439277fc84a166b866da78d9bd0d5562aa5605c4bafd3
z8cd89cdfccb5530e8216fff041d7092cf5bf7b5a7c7bb90788bfb82e018783dd424188a31de60f
zeb5b3c92ae2d3494f91b7f92f1c8f232bfe0ce6c7032242eaa4195df0ae242fea932d2bd43585d
z8f136b77756270563908e364446feb9aed74c3b1d1579a0a2a0be6e8223cd034acc85dea25f8ac
z0f1a35700e1659d6d4671433bf70124c23c0d4f94730db0bb00d47ad5adff114b290a3da44dee8
z514d1718c70798bff5bcd6883d9d7e8cc807470404ba307cdf8a06fc603eab12f0f70f68e1f687
z0eed16ab679f69a5a38047a02c5f5cc8af1011b9666ea3480786f76d5a0faea4aef9c29980e20d
z931cf3c669ba8a54686f3ac4db09c29e60c7929791743ac5d1b73909aca7833ef96a6637d180b3
zdfd78398f9be3f27ecf02725a8b33445f80b596019ed1a2a91c3e02a8326e40adcc272a6596e54
za40cce30949f8cc0119f5b5efb27b4df6cb5ca3a9d2c4a831f39049856ad346a5bfe30701abd28
z1610bcb2e8c4f01ab61cea4a6b6eaf8576f54c44c24142791ded7bb9651ea2eedd7320bdb6259d
z79912f02a9ac3a89bc24520fabd641d3534a8cccfb83594af0e9f32c530d9386b17612da4c6ba7
z08f7eb2fbe439ca53ba8a99ee97c1662a6772a974f244e31de991af5fdfbc0085913655f0ff097
z5fe86b8ab990a739b54ac7c42dbe91d3b013bf8165ac143afaf15e49824469a8655f2ed89e5347
z55cd1cb0226510b796e82e74a21a50611ee4b65082b1d3b7ec03252842cc1efa413546fdd1d14d
z6d3a27570ed28a54dd94d98f9cc5d62eab52e6e0c5fab452106ab624f3b8163c3a423e93ff8050
zbecc70f096a7c8d47674bd8fc0b37aa1dbf9413a22ec5551329c5cfe708df137f89e1df9bf8a17
zb99d5e81c9e587a3cdf882b685c36769898420fc59cef0c48d56baa95d19b6a9c9c60b0a073079
zd2e3dc14a2b58333e46d387518fbaa848c9f73d0a335fcd72a621f061cfbbbe689d43cd3fd7b48
z531246f66f8183b502a045eb023af39c2c01693db5943ed5df8678bea6ed45861796b3cee20a5c
z57ba0f0ab5f885307f6c624e27913161fbfab1ef00a04793fae3bdfedb6df5039d91d14c164f12
z4a09043dd88a79fdfae84e196313ed68e36b1e9798aca11102e49b40679ef31840a3349dcad78d
z9bf0817deed899349329090a134cdf31e4590e29b5dd480a0d940a1a366d69238745baf066da8c
z4fc22dec9fd6801d52f8b3c4b1f3e44a6d09bd29b429903dfebc33428034ce7eb5c2d4132dce6f
z4dc30559cb91d687446351dfc50bdf29242dcea12fdb19b27acba7b5ae360b1d3cfe754348f15f
zfbe2f06825b6c3d96a612ad791aeceea59a5c157923827eca758dddc5a95c3f13aa16d0997774c
z6b887d43a57c67e45db09b294455a27bc582165c6952717108c4f9d8a819dca08559b6d2ae0a25
z2fc1bf93fb49ef7cc01b5e6d8179793beda01522ee31c1ce183a2e11514f369ee8905f85f34d95
zf5d151813295b86a5f1182467ccdcb36614c26a2f6919878553cdacf58607c79c0deaab32871ec
z5751885cbd331494aecdfb52f5af53f9ad8264bcb02d24f6bcce2262c5c5352a515d91642b5df3
z942463d079d717b547effb9e125692bc0ac0c39378bd53058a4ae330b12d2711c49c1706c3e9c4
zdece3dac2fee77e76520b9e4bd791a459069fe9f2bca58a72928194b36839c416de8ec0e131e2b
z738a3bdd591a22f9e6415e005f05c59a040fbf7e8dee188c0e6871975538462a77e7de490def04
z2af0e562a0ea414f84c7426041027b244212a75a758a084633d7f8ecef89dc7ac37918e04b50d0
z7de9cfc796ac4fd92ab4c0ac6062882872107d140e11ec3cf3fcd4ac13ce86c83d63ba3ceba425
zf7e387f854fa8560c58092b7f6e6d4c74253822cf5a965718aa669a868765517aaaee40db6eb32
ze75c7d4fa26e16275b2491275f4e94463290bab26302e2f36231eeb7164fc4b4bf19d2f9420f1a
zf646adf26a2359a3205b71892e843c38b4b37b6b85686aeada9e165e4167293a99eec9fa6788cf
z04dd11150ea149241fcbf7dbcd16eb6829a5aa12911abdb00d2e63f5c3d3294ffc6280bdba14bb
zbe43e58c857a2c39e84ae00e425b133fbd0ae999e70c11c5aae827dbfc0d92076af6743f5f997e
z548274ce0277c3f4338c42d7b044ccf9735562417f40e45f5b40a3bb5696279c36d1e795caf67d
z900feeb829d8f91d0f1445abbffdf9baa0a0e326d739e0709da95fa218ba9ca1cf8f504e175e3a
zad83d821f90170897d5468b5a624a1e15d1fe23c9956d0466e4e51eb1a717e2d8b86f5d46dbca6
z539b7d2070d6f1a121f0d9c9dcb60dc8f1239d2154d3d3e473a3c1df7a5be5c51d99af3139b78c
zeae98ef2fef07904d3ca9a313df779a279ad7e858270cf8ec3e2df63050ec3fc970162d008b295
z74907a5ee14101b8ba6a360e81e86baaf659524a4ba3c0d187f53684c062dbb7dbfec11783c2e3
z20b670c2b6cd89df428f1ecad54b1d8b079d0545c4fd5b2e741e2729db19efabdddc5275cd2eb9
zd65765c8321ecda253641d1f1b722c4821da75e23e8f4db95e5bd8d6f0ffdda3479f6d01c15589
zaa4ba647d995263c1fe2ee799b6122dbe9a73cad031fbb94d379da636e4b29fdeea908f421792c
ze49801c80881ceaf9b8502f076343f719c0f785fae9a6bef44cb1f0e745f542fba3470e78491f2
z750803717c220d21694534bd325335929ecbc9c0009f34d01f94921e4ee8726ac9e8fb9a25b4e9
zafa3182c7ea05feda200cd4d0cfc29eabfde56f19e89d6b6bbdd498b1024bcbc77b824c9498a57
z9442882529760ed249f3bd8819687bc059df72a18eb4e69d6467e8cc1faa832559a5b00db53e71
zf0bed69623950b9119f119944e9ed283708e6d0506932efb901d2b5846ef3df7a3c72dfced5f5c
zba74c05986ddd642b923412875214d595c471c2accaefc5614fc31993fb05447d2da4f9c33c54a
z4f86addce19ce4e349827b702acb0c6f3ac322495a0198a6ec88723eb798b4bd103430151303be
z75811ac8fb42504f5f50b9c7fb866c9a02fdc169363448bb33f555995000a8ad4923b0fbecc70c
z6d35b64bb43b92fea76c847e6d00cacf551d6e5ce4f65558acab0bafcfa5027f3cbfe077596f8e
z0bdf4d747c32c3d525b7d9b49a2e4f428f89caf13d04d87dd349028b64391edf12e8c717c2d5a2
z3a0fe8d90d28251156f78a4c756abc4f0544b89bbcc50f11e15bf550fa554fdadec3ee72218357
z938760708658285596f84196091332a9470df73398bd03558432a44d3ca43bc1bd058101564b08
zc1c6a69a6a8bd1b45e2b34e4ddfd5fc525d5fa6e464c95990809095c0b114d63f939d7c3207a12
z915883e1b2ffd5c88b61adff7ad6a97d2256431d718f988e938f21b1123d761a2f937ecd642fb9
zcfb575f6ab23300d52f21f9f59510045fd54d2e9ebed4e4fc263c690b72ab318c873979f35321d
z41ede91351887c7637e56fae621278bf29b73789cde6175f7c265c7137107574ce5e4d249e1622
z22efe446863d48725f7fb1ac1fd5aa36133a89228ccd354bb980bfb1bc3a56877cf48da63acd67
zbe2205eb86ca7bebf3e8da9162a573eccadd5dcd2a44e899fe80af015b7e4dfe96ad5edc885550
z3a922e1910d6e7f8a89d6a9b500e364d87f0de3876d0aa8f2e85d8e0c057b91910d9bcf33e77d4
zd1982bdd0ae9c1a2c3e0de8f0bbfd4f1b8198dc761e310a647a5a7d2650702ba1d39321d72e535
z7ea632d2aeaba20c1de58a09ef2ac0ce1c7bcbecb4ade16c8455759120ef914db351f451a4d423
z847c71b79fb7acf4b2cdad7d9c44edc0eb64675cb87784c25d07ada087f8d27d6900ca7de9333f
z890217e8072e8d53d3e6be81dc21f6e8347ac7fa535230058937bb3353e5da21aa960ca9cfb142
zd59be99635785c183a0741f5249c754f75828beb4676378a734bb44016f56c2c8625d55189921a
z5a3be6ef76c009838c9a315c01532811fd9af101dce18e12fd6c17a1acbab23054664b791fc172
za350ce77552b6da5e4233d750892e4d5b251e41480941d4c03883dd3feb6347a1dd918227669ce
z429c09372e1dfde8a0cd71a07b866d79ed8afd596f3ddc3a7b048961d02d46c5a025a66bfacfa2
z917e5ef1b71fd6d85a16cfc30b4932125fdb82b5f9a7365b6dcc6a249d0777da0884567ffc5c64
z9c77a8b29b2050bdef59e2ab63cdc783b3e00680baacaddd3d7c6e746d54511d9be938116ce9b4
z3fbfefc3b5dad4aec01a771cd5aadf9d0af0586446b59618eb2d3f5136c7c488f1a0f87583e89b
zc55cf04d5c2071f9f5f7980b4f1121265921447087ac762ffedb6541f25221bf1f7393dda2e9b8
zb6b879582250993afc741cf1718657786399d32640dd77ebab2f5ed8d83eb5652595a7b3c92dd2
zb52bbb9a9451e62d5cffbcb3bd47f5bbf2402bc5ddb577f5ca5d1d1c94c1265548adbf4ad3fecd
ze8bcd332d6d13dfc10fb0680f736476de9874d5209b8746fefdf3bb57ccde0964fe7577c69cb6f
z98d3008310af4d81e1afba4e445820db57d82699d0ba381ec88c879baef8981a73d87dd1f10de3
z98b26d85c485cd9c9d5523275b5d4f33229217943dd6c02710ead4b6e5059f8c7d73189362c603
z339702a9fa7512cc24643c95168e7dd584f6237dfb1c88262d189f6c8d5d2ba3a65c2e9cd1cace
ze032982589ef3dd50e4b3d2603ef06575181817d6d0b01ff0cd8af301931259d45976b7e62b326
z7e2c62188bd89ef6838c9fae5b1fa4fa3b39f6c8d875d07adf4cea4920f4d22fea8a049452fe27
z465712255f26df75e51a90ea58cab73b43f69e5444ae06976baa79739a34e460e4eeeec333c722
zf372ecee1c8644460cd62c01dffd6b6f4f52869da0fda3e6d0a0bbf602186a6db4a84a6c1ada85
z5b973ff7002c876fc8fa7bed289e9feb8f6899e45e22550a9029cf65306184c9fc8ba7fda59b1d
z32994be66e7d9da8de2eccba336765fd5af2ba13be19ec5f8f0e0c919677402074eba384c1baa6
z61da9a2e1f94fe55e92438eee2579db045fe114b51325485668741a7c04fe645936289c5cf02d3
z79720b8906d841bc56c033936eecd134513bd1803d8b5f660913a30dfed9edd4b6870e4bf86600
z29a8937ac974e40e2d8e8dc5d57db1c20662eeadc8067840a651bc5a09f60cb913dbc09951308b
z38141cc984ba049bd78d7eb5ecefaa5ccbc57a9e957357bf5169e87e76cf336090b4f06758a5f5
zb92362aa6c39667fda2a17b660ed425d19f8f7e58754e6a4dc9a5c387fd2489a3bdf3c974f7c8f
z5ee4fa6fc645e3762f67b2a283de27f9b0d11e55db380afaba41913343f33c2396b232c29012c9
z376b97a594e17f645d622bdb1f51bd2afe3131b07d9fd304a011f54df2df7ed9ea3345c9efc261
z2da98edcdab76a8daf235e28b4f41f96d17a81740e9f86d3193de3bae45591b746a66eabeeace2
z6cbb4cea697c054834fc00bc3ca6dae088d77973f0b7136529e888148674e7e0a59ce7bbc42a31
z6a6d677f05b6550e01bd29ab8cc090755b45d7cba4df091b7b4873565bec39574ffc412fcd71e8
z4f94e592cdfc6cf860a4523d0c1627703f26cfaebe877e30fc709a76ce888f7d3b43666d48a88f
z941d12acf679bda1988ae054c22ec60c96d26dd14d6e292e2b3687b1fd467110f04aaa238655d8
z32fbc88ef110dea40c5390a35fd2ccde65f7c0f64b60f96e5f0271d4afc32d58d46ed753d391a5
z9c3fc25fa3087224ce6be96fa692e0492f0f1ac7ed4d36b6e484c24acc7a8b8e4ede934db8a68a
za6fc1793ebd101b7a6a81731bbb203d258beac78b19f360a568ff3aa713ee8b571eefc638285d6
za5d13f99d791bcf2f6fa0fc3468eb91c98badc4172ca3bc3ac63770df42091abbf350e9a6df5eb
ze3f56f731b330826a505886263e709eea9e01f11bb944071d20831d8ddc46f22cf8f635947aec1
z2e5158fecde15c80e76983e4c2ddb5c799dce864c5c61e7b5969d5bdbcfdd9b1225aec48670873
z5d5b3a1a29df016c7af8d4be735ffbc2717d47fbb0d466f1d96500a50912d1ba9c8d4302786a85
z82c512d920fb3a603945532dec589e64c379a2341ae485b0170794935aac53719aa15c23e3e582
zc8ceae953c5737e6d088f57517ac8ea8639ee21f2218d789460f370c5dcadeaabfba1743b2da79
z239453db90bb3c8840c668a828130be0c0fa1f6b4d44442d7c3fe58da353304e6f1acdfbe9cd54
z01c2558f91fa5de06ded5675552a4f9b87931fce92ae54a5700b606c457f2ca82217b99f679a2f
z4f9ce201ca4a4cc000685e635c256fd812832342746828e1dfbbb6995b2316b476d33ca78a2441
zc68aaee91fbd3d4f9fb6dca21d60700283858ea240d6154dfa791ed27133357fe1c01ccfc8c5db
zdfa84fc2b70f7f3bdabf1968ff1e7405263437ec08be4334d7bd556e8ea45806ab459bd094bb4f
zc6e79496db1d67f250f059d5c6af9e24e8f7a09ffb1cef558469f89e266830ff4b1ef124263a15
za9bbde154be1b65fb19d7beb7e56b63042ed587221fefe2aa84aec6deddef4c106bfdd495f014f
zb6999181fd9b3f0f17b73623733ae4e69d6c8b377e4d42faa0e49c896207da087dee65cec2e58d
z05cc7e1b9b9d70d61a69d9d09d4133afe69a06b94f5cace22b5536c42eb575c088d3357dc0c6d7
z9f10207a8bb26485def53bd42532424b015a7aea926cbdf90c7d886259adf00d837a0991b7430f
zaaac3fc24dce6c9be6aa0b21ffb3ffe4c79149416322c19c5170dedb1b268d40a51105869bcde5
z225349f53f73fe868d6552a4c4cd0ac1692d501e4421499be157d2d621c7b44545c271a4439444
z04af475334faf88d0ecd73df8a0f0f3887036055c98acd308175d47f3d46a0a9ade91183e46b9c
z6c0e0826b76d24cd3ba65102965da9b65703f3e5f5362e37cf67104535d43e35bf7b88ca370b4a
z160aa2d725f197e390327b8b8ff88f05a4c6e4cc0095ad61067a8c06d2ad2f485700f85404a70c
z630003254e9172ef956983c75021b212385a72e88aa10efba003340e8ae3c2af502328d56551bf
z9ab34fc1988700e7f16b3806a177540e5185b9b2dfbc312d63263e74b863c3445463c10f989f52
z3d1e792b3d1be6c9a10f0c7c92e76ef099180f52fa47a8b484ca1047a4523d56c4220d9f0d3943
zee286adb729a5c073507415f09b36ef9f4a185dd38b68a2209e23976cdfdd761ef405da3f6bfbe
z2da1d34690bea58f7a4b85b9c31d4e05eb8c9f14df8b963d1f5cead49f6929548cbd006e67281f
z4293c7e29eaccb787712c36e2749b0693536c15f876dc98099eaafa10470f204c23c572ef37369
za6d1ea5bf2b395391f7026a99d4f8106dcf097523bd24ebff380bb9f5094fc0cc5604952061559
zeb86ae0201059f6ac7817c42ed3bce6c34fd428a8243655f603759f073bf4077fc6b8788216114
z907ae6d264710882ceb7d6bde97e12e6ffbe38b4a47b705a4486fe1374998a07c682fdb2cc26f8
z7edd1857dcc3318708e708964017b0e7ec0120c043b13a6bca997111d8dbeb796af4e29818338c
z47956ca1d9bb716cc8f12db8f076737bd8f3a917710ea0275a6ade4e004200cdd937998bc71e80
z765bdf85ede59865c6fd1cb17b26455f7f52354eebe67b1c8085a90f5af8ab0144f3523820795f
z7da77b8d6f352eeff461406107bb5375778c663a111e1f54f22777d5673dd279537846317a2ed8
zb223023592e9a1667fa6a2e1fa6912bd47c7e85e558cdb52a897b8467cdbfff8074be018ff0da5
z26c782e2c302909ddb9d08e9c067ef453e5f84d2886a6706054757fa21362e90da5f3cd39885a4
ze8a9b67b3873780f6c607ca7063c6053d4ba39748b2c676d47c61d803c22eb8a97546eac701315
zb0293bc6d8cf56d148e1de9f975d5557762006a89fc600c5a7cd84040f8c1bf4919369b1436133
z6bffcb52a85534665afa9a619c8246ac2b8e43c12d3a960cc37571067a2abe9e24cc68e385e903
z15355c96b392bd07bdc7cf2633b9719bad3c6c12af269d9664e3eb267ab63048efec4935f565b7
zfee9904ca5fef28d1d383400786fe46cd0856698b0b8eee0f46d519339165ef77292c0c25fe8ab
z8d245c4936de539a697f245f7b3ed63813bf418a1f3af8bd9e46cd8f3e08e12f8ddf0433fd2169
zb66dc07906556f2ef934345e0e547e747a48d7397aeed187283f46201da3ea450445c8a5a094ab
z7131b0f49abb466cb1b4027dda633d0d8c6e3abe8f62bffe83156599ae073c7f91b0edb35db118
z943451e205e8f0dff80007419ab173d7668339ccef5ce2c09bdeae5786f769dc7f2e1a32397b95
z840eeb23f36db6fdd7ec0a8e79dcc4ac47c69ce3d48a5ad38199460c42fea219095495cee26327
zab84c85682b3830e6b086915c30e98229743ec4f8386c2f8ff13023cb5b9c7d0478586dbd0a2d4
z5d08c703f1f595399ed4081f2294f144316d59eb22576c38dae3a5d57e4ce5b2affe99665a0274
z862cb901368ed81b2d6c43e48217c12067cae9b49befb7ef10355b48cd4c2c886cf3926e087915
z4bdebefa2699cc67e99efc2a00d13b6a1329dd809e982a019cdfc1801ccdfd74de8e5542f14754
zfda7a40965bd228973291fc9116e36df4f6b005476b8d080ba21eea5417fd452f293a05b717b52
z6781fd877ff3148d0d06937cd2272a9ac784eb3097a95d27834d2bbcc8cb7f1e7a1369ae1e7752
ze69170bf5c7573f8360bad825d95e03564dcf89290b86c909c9a351a49286b877c5c252d85a992
z9db05f379417d4bd193af2b95b460e49317e239f5a55b6d5f26b6a8a9e984c6c1418c93e93bf74
z80178dde93b54e201bbceb6ca59995e298babffc7e2c47d6e2f4699ac0d6cb7b90967a25535400
z789468d885d884d9bfe1cb60fbe6e1e4dd658ddb1ea2b50d2a969da4094eeda132acb148e069c4
zf06862df9bb1e5259905d024552d6e41fb2d6054b237ba428a8ea057545eff6489abc7c91f27d8
z3f118e79d383096f349133f94265106ab25007f43f511380611f1851d094f6c2518ad8ba0862d0
z504418e49a02ae3e3cffac9e8c14955e891209de715d915c1db88bcd810082e920dff553dc3615
z6f5e2b1727b1dc0b1d1a1b569e3cee2a0b4399351d7c165314e288f1b20e3e5107c9a43274ca46
z89728756ce476d704428f169ab3d46495297980b3a7f704426252df1a1eff25adf5221d86b9d05
zd99b4667d36e23ca369f8572b5614eb519c1013724e4f6107e5afb51a32f9f44ba671eebddf598
z9a1aeba38c9dc76e3cc0a34aec29f04ac7812752dcb3f74584e6a23c725577d4efd9d2a3d7d765
zbeebaea2facfd600845293df0c30cbe9e5e426551eb5fe324fcb4f788a9060631ef4e287f8838e
zdd035d52a509d51fd61eb786218b194be258a5abe51f0ba711ad27748f80b7b2de2283d8c5f532
z21bd78bc5acbd7b05524a61ec0f6f867075235eef3eb1a5053b18565ebbbc36111e60a9eb28b35
z87b0b353d4d79ae0d9f382bdb520301fafb5c1c20d90efe6282e797a98f11d54ad558357d753dc
z498a7de3734cb651113a12b110216c2dcca6154c17e92cad78c61dc75dc02fc8300a48f3b9f4eb
z0fcac033e2a1ef304b2b3a582b73a14847bd021f4a8dbd8be64c75bf9c84160a86a570a857061b
z0462afb557f2fc938c077f4877bb25380b31e9d62e0bbabc87722d5765518b7f6d47b55c48a91e
z0d45d83ededd04bd8f7824d7a833adee3a6c36c5741f5bf247074a6d5019d2b12fe058feb2d3b0
z84cccf7bdaeb39a9ae627105f0bf66097bb5905575e1f3d5a369d331114dfcdb5fefa89a188092
zc90858de88f7d0da3c2fbbb01933f7e21ad7c726776e992b44df926fb8494399e3dceaa0aa42f9
zf804f67d1c1e582bd7c1ed05e467449c6b8b1c3497f062b1d49dfec1fde76deeb35e5d99e8268a
z513d85f0e81e3237bee60e6ebc20de99eadb23c01ea918ba213e0230517aac20997e902ac2800e
z1c4fc6ddb04f72994910a2cf82048ccc554983fc49488ba4af4684376b726b7a77988dfdfc079c
z9a0cdd5073fefebf41b8c63df8dbe4010da65142cf1f59afda3b95cd943cbba2efe78e4a28ae5f
zd2822995171fca2658c0b7c5338f2eb1123fec9ce7c0cd338aa890bdd95a54348de820f72fa3c8
zf2644b74c8aaea199853dc70085fbb528de493f1bf48f61d71b562a00362ce979256074bfc9b17
z544640ec6e6f132fd0148f562b407c50861b6e867fea66bc1fd857208b0f057d8cbcdb20f8672f
zf93dd4f59b049895212f39d6e83540fbca66439615940215ad9628774bfb64d544ba11f02ac4c1
z49ca620f05793a4efd5b5687d078c4d2789d73c64c16def67068ebb183f139cdcc52d158d63446
z8b75dc9b0cea7ab4d3b7671011aa679f64fc33c3d5a514abdb200defd36f4821937a6ad38555a9
z311eb5134f911fe576020b6df197a83cbcaa453c2d4051f3ac648ddc2e123207ec222c70783860
zac424362b0ec7b77d75ccac44e37134f582f067e0940bd12e57232bdf42e278583ce3beae68af9
z8ddfb3b000df84c59259f55cef7ca11a693b06a48ce715977fa6f7edfefcb77fb9904c6c301ae3
z92992bbb882c72a61aa92194e292db2af51469e09f7428da440ac8b8a644ab0ed86753e82b0c3f
za76a0d1bc37cddbe4ca5cb829b1daca4b6ecd6554b72f2884108d1e566073dd2a38a1f9d1e408c
zc3d26ad4fa6699acaa8246e70815435c18c5612aa67f5d0258d569a00314e3be2a61e31b85a8ac
z7a9f20c8b3e2c384d1daea4e4ec4bbb79be6fa144cc832eb7f837e605b515742cdd98da4b3fb0c
z8f73bbebe7d093887b174e16c98e52567153ba8f78738e77b6f53d5e5aa2f0f66afe182465142d
z67c5604763426a841bcd40f7b7f17b87eb8eb68884555fc6347a8e34040b0a0fdd26842d4ea22e
z7604a3710a923d9d303fb73f886b4e967cec704f3684d100799b5dc370bb386dbb76b118ec58ab
z940008c592921c7855b806c81e6138048909614ecd3b6c3619f932b9f148f9a6166caf41f79d1e
z611b2af5bc424a99386ceccceac762a38d89a538006e0732f09f7f8b01ba330dcff37b96a237a4
zad9c46ecc5796d6a0a8f2c69cf56a6d23e8a8a3771787c4f3f507a270194fddec57b290bab2e3e
zf2d529154ab2d2bac912d2e50e7af0d4228bde1291854329434f51a05131bfb9ca7761dd81e4de
zd0f833153a3f0e3fb17590a63276e038ea1bdd25f8e1b69cbf1c6f704c539aa06e001933911995
z4f6e2d71d90c925e8b3a8a664c8ad3c4b8df5b33e5f6a38e2869f69fdd212a9db7ab5ba8f46a9c
z0c0cae68fe5a1f7254181e6eaadd6c903719782087bb54fff22fed10a9dc4f580b06bbcf901c24
z7b3eb8748ff19611832144e034e75deeaa4ed3ec99909542acfea7a175acaa3d9094529141bc22
z74c30e604f308d6dd53ce36be58556614d420f60f1b13b0570100eb30151e042e7a518985dee65
z320e4e7a1bc6934d436657286edf86caabc318d5efcc61dc05c7781f062542c6f30885e8dd660d
ze9b547ee0f514dab834ffe59e56bc8177f59f8fbed3c554308148a82bbba1b92b14f3f94a763d3
z18fd303ede1a6b6dc51443d687bc050ac88f5cbd9f1d6c787f0b3046a97d27fdca937f3594d3ea
z74d54ed9dfe14cbfe5f40eb15a82791455b13ee8a061831622b7b6e79680b08f3c90a179f108ab
z7f180b8efd46d2b1de187a65fc42c2f2a0159d20f80cf3e01f0d7d410e9337409e8e87c6ed7fd9
z3c1f6fc96bdff206a3f1cf136f85e328331e2b131183af04f8f03f65af5f0864c321bc61db73a8
zcd6c23bee4cb3a9751ef24c3a3e1a1168c3a5dde274f8dec489e16ddb7365237d29230b440f14a
z51eea6d4872b695f66b079fc09baa3f783eb8aba8d67aae095e475fd6b951c36c692cf0d0cedbe
z9a4360225894d9940dec67f739381b1a14233e54868edae93ea8daea87953a38838ad9288344e1
z370e4f54ce8c0715331425996571fc7ded06586a28d63313e8c96bbfb2c5aa5037c0a3a958ea49
z27a88531f1bdfc7765487e32e63bf5f1ed4bf1dfdf453d95e1cb91759a49ae9c5acd227e80aa4b
z601af47594570d84f516d20bca834cda171371c94b0f4721e228a3661b9776c0e3be30b8deff80
z7ff8f6672f7dafac90ab32a0dbf17cbbdd303a2995675b4b8cb709b9dd0b5d9e90560d01baca0c
zff64de97a17af033e9d87c181f3d1b74c507742737d8685a662a0cc8356e0f21b65a5827e2ef68
z1a6444b5cadf891d8d53da7577a60a401abdf8296f130b9b984ccf96909b5d38539f5181ade730
z9833eeef3489dcfe0391c9c483a961804cdcbb90e5041034e29db27b96f7273170625968d8b16e
z2d05e4c6e6ff6ee35ed11841dc59291761408b0e7b02e98bf00ba66b5fba98584c2b4f4eecea63
zeebb21f127db87225672d7202914337b9ac8e5be75d8628016b0bcf1604b5089b6113273b610d5
z2c83fa110bbba3a61dafe0fa042200308cb89849af90728ac812c069c8822344394bc41b209283
z0d6d7d390f9f8778d3d990bf107c800b119b51f17f868e757ca17aa8d86e0aa26c65e03acd27ba
z42e17783429f2aa290ad70e286b21723dab23dc9af254740c7833b347d4db461f4bd9764cfb5c8
zf5fca6af578b9996accccd682055daba0122ba35f23233c50ac020bc261fdb212ad7ed18f66216
z3533354bd1b0204e90b8b3c407c301bd7ca0a77e146593b357f1fbf4af0a98ccb99fa1ad5017aa
z0ea0ad59ba819bc45b75a4916a79e9fc4ddcd5c848456231032a9fa8c727e52767a6db49244fe9
z68d229c5b312e29530963d3e02e123f5f03a3402ca95f23f9e535f4ac992fa4514da5f61222c6e
zcba2080a709f4c7d77e566f7bb43b3b567a3138ecb87fc315115bbce03da933e197665cb8d585f
z866e22850de9efdf8c3974f131822510d5b96595033dd7d68fda00403d68aca20751a7f1b177ec
zbdf37ed969fb9370af6e4d7f806eff7d60b3ad47ab595f71791d5d3b2d4ab136e680d3341ad4c0
z09a7bd8a522e4a518727bdf546c727a984fd0172f39aecd6c5bcd73d512541066e715d79069e13
z69719bb5449be06bdf35a155565c6c9cc92221a031259c6804d49f2699519f47bae9244e1f007c
zb83db09f5e35695199c7ce4bd522d4ad37212c51a568f40b2e6ba4ba2339566f585092cfa6368f
z85c499ca7b1652a11b1cc093a90e7d4c511e9cd92547b6cf0bde7f983a929a0c746ebf8d2d18e6
z404a4455fe20b12a11e64c9d2f166560d21454117c744097eeb2d0f82fca48aee2bc872a7a329f
zd5aa19fc754a526212cc3bddc5680bc82fbcf2eb6c389fa5e8c107803757d626fa1df977763878
z2115fec3b695aabab8a6d0a6f99af3975001301560e2ba475d30a7715d621c5178c57b036dd2d9
ze0ec46be734f946d831e03d3479451ba260f7b31c36962139871b9039b23f44d57b21665c4cabd
z22fe0aeb53da4bb87d7b408c3ae1df3926f1c7ca72bfd25fed23426825899f0d62949ceda5017e
zd70f595a4fc57d625394a2c62ca29cc460db6e5833f966cf756788345b8433aae14777bfe83bb9
z554a789852167284ff97d3dbd20c35d440ae04e4577e8e9d7f7813f6625047bf1181bdbae6e1f4
zf029eebf47ebb30ddadedc0a65502f935e0d971c9829550bf8bfe1da088b490b3940d57eca13f4
z5c55562bc43fa460786630d9e03a06efb2353175e071d244d221ad0e5054a7fe6963ca31a57bc4
z9068b947b269a5ea1ef8475297fee603b619cf53d7622e5d89a530fdb95b422aad455ac208c1b4
z2464d56ee25bf5ffaf855d0631906daf58d5f58ba84ef5aa0d674e6d419091ee0b144382ed6e31
z3afd358354f0c5e73974224b86f0b906ec9c862aba4ab19fbd25ec03f569ba88a33c5ecf0eb64e
z832376a25397acfbc5c0085391701eb21053974e89256bb99c444f938695aac0ac92832496535d
zfcf52f6eaf36ddb9a0c39c921b09ae6abf2acc195ce63888094694551f245b3ab7af2e773c8145
z3428069599012c3c30b3699b2cbf7116f9112cec66195ecfbd178649760cd4635eeb6bde23a9ce
zfbb46085d7cc10112c388deed5c4824bc4b155dbd41222d388c9a097e83e8a41f53f59adf0ead6
z7e48684582e0ec7a9e4516926bb30ba7de771d34456438fb1cc7d6b41cbcb4eda67fc518001ae1
zc32d8963b5ed64a2fc7e17b83066282d188dc9c2105fd2608fc0dd1cf63ef1afb456b532b23956
z24f058a61564b40413e1ccfea699af3f8aa4ffdfde9c340a27990ea80f420e660c0f9e26f34a57
z78944bb3fa92edfc2640987df90a8fb053e10483d4ae6db2f0da13f451863f5ec5839c16c4de11
za5f1ebb277ed87b952119604d3548ffe6fc3d1bc0e56dcbfa594ccd52ebe2e61bfe6e7670dd48c
z8168c0e872ff978c4f366fb2f14f19f15bfdfe5081ae974f0d91cee7cfd4090f7cdc9705880de1
zb827b31c8661adfef75678707c0e9b6ee7b2f93d13e04d4d9d944cad3af42fdef589fdaecbc887
z821ab28611fa0041ce4ee61ed45cc223b6184888b9635f102d74e3ba0a7d3af5a8a8de135d65cb
z9f2d7128135f8d220027175de1c67b068e9f9c5f45f56af417e021f1466f66edccdcd94e90dcc0
z811687afb9a7c523337b7411bf8a9ade3db45312c81522d30a788feaf8489911af9201d449a25c
zeeaeb5a224c562386cbca29f9324a30d666341c566a7f102933aa4b85c0346c6d3edd76142e5c0
z9bc8cba69ddd92d0b3b32cf12db13bbec7d5df897fe0e2f77b1fa4438baea175109f0578358789
zad30d1a09a6354988fd53be6e56b357ca3188f2dc7ba5010f27095854220149964d6ad4f2b89b8
zb4fc1078b7e8fac2b1d4e32638006a219c8379866952387359f68b745f3db6e175f50fc788970d
z1d590345e1ef1b58e8d5479e018b181b1b49d8cf2e40ebe66c61ece2a5c3188aaa8ff03ba21fe8
zf3c2fc00ff5a7cec07087da521c5f81cd7b3930668f0705134848e78c9cd36c96397482db98d4a
z695e335d47d56db430a80bb9a272e993f7c9acee118a35d945b5f9f6631cd538cc6c3ae99b2f1b
z20105983538b4544c223ba8fb98c803ff8a2a162bf988ccd5900af3a55c5372aebf091fda65645
z15a185aa24a94471e3a209f991d98101487836d217f3863ebbdf48d9f0e0427bdf7548d4f985e7
z590d70238528054522de1c56511b64cefdc29680870ce2938a82cf2e4e1674a5ab61c88d1584a8
z2c0d8882bbae39d476775c5f02feb27e352c07aa13ed3bcdbf218075d93a787e9de5c0e55b38cb
z4b9f2fa8576ffad14f4041ed9b73299212a4cb07f2af393aba6a4de67a14d88f9155e6d9a88f12
zac1241f83429c5b506afcb98e1e30e62bfed65f980c9de59a76c36a62af1e57333a5eae4060f19
z154c501b582458321f942be2991b71c592217b74066d1f839d1df8b7a1993beb56293807b6ab9d
za89bc83eb49fd648105763395484d4506771eb95ed920a3908d1c162a1bcd02ea4c6778a484956
z92a97ae5f13233ce5550f3c8da08c65f3ec33def5293a84572532428a0132d6520308dbd2ed9dc
zb8d30c08491a0977fa928a6b703753d737e24f9b99593ab7a9400b5b42f3e847569de3736a5209
za43d5f86adfd812d1038187e2329ec84387975bb8cd0fc447fbc210c238d517226481cc898860b
z87825bb401197987efbb9a807b7b27935ef73d89714d10e938b33423f6dac36bdb33e6e6573fb5
z79d639363cc2eb080fddcf17b2936543b0ab42512b63a987d82dd8ed06511fb307fec9205b5ae2
z2560d6d65443cf457349194d1f1907ebd60c35335909952ef18cf06e5e336c9b757095e49474d5
zbf8105dac4170f4bdb78883dcc8c586699ce3698b1ba019bf90308c5e8a8d0a203b475647e72d2
za3c90b0f2f288f66078f2be7531419eea71a015c489fb19fc9f909987176dd1fec06273f325ee6
z63f900afe3c050386b1c85e636d0a87c3edf8e70571a472ae56aa8fe694657e3d75f1b84975e28
zaf3f23e7c8c6a798b3939a591ae7012c6067ba1298c18ee85e7ab2a8cf56d17018fa42ae85193f
zdc7bc39e91ccac869b6d9fef033db2087b6788271b1f7de8e036f9b7f154aac36358a183ad598b
zcab4e3694feff164b39e1688f50aa56b3eda20d54e29cccc04107a86b5a0ef457c900c27f62b40
z5bbddaff1971e4b82c17a51eae241556940963b1be57b715fa3dc1290cd78287e5674feee14c59
zb7fc867bdbc8062201ed0d0e40a46f868028eb9a01efcf55c17a350bb0a2ca0492ea2461bd8a4c
z6f3f182e0028531aae964751c0551c7b04c2b3f99f34f930cf794557e462f1a69965069958ce4c
z765080ecbe575bf003621a9304d01651f2143edff51c767bcb6f6a964d4dc84ec06b83191f8b55
zfc7180cfd209591349f3f86ed435433f860649ac728e4cf67e635b0012fd49232e14dc60ce343c
zd8251e51f045d0545c2339d19935a9ceb2b7e70bba99396759a56112c05ae731918dea975d5de0
z11f887ceb409d51367178c729f3dcb91c6f57ce490861aed443f4ff12670681c1d5458318b0716
z3da84aa600bf7cf6b707d855a4f03e67e9360657eee7bb9ccf182953649c0c1bfdcb183268e97a
z9cafc65a8b357af2064970ef1d075ee9b821a706b75df9d26307b613641beafdd233f15be551d4
zc8d80dcb85c9c658dc3eaed172a157de6bd8ce577edb9cf67028a6acbe2287ba6cadf4ef49d264
za18b6f302d535d8000e2ccc59575755a29fea769531979b0a0d56a1dd6647fe45d05564c7ad693
za61f190f958f51df27eebb2159cf375633ddb2491bb77956ce962c44d60502a0c653e2c08400d8
zc9543fc6c5e4f21b35d3a1248f57aa0acb274c0e89985230591835fa18cf9a13e365bf0ccf1327
zf3f331720dbfce3e93b4a2d44543eeb69895202d7bb10e7b5ae748d99279d137376175f9ffe52f
zee7be4328f270c2c48ef4627da324e9dc55bbdf999b193b5ebe4fedbcce7b933a2ae3cd6164042
z994fbb7231b3ba1783ac81c4ac280ce09347f833566507906a6af60290b107073848d219c1c2a4
z3c4a8013ebb2aac4e37753851e13903f37d1c87e751a24c05550e421828e2e3956492fc889720e
zb47d6ce96795c0de5f3648aec21e4a2ed78025d0caceaa4fa9f1425c7b6f0835a7281199c992a4
z307a4b61ae4df74663a8a3d7540d01e299d29f1991121c0c6b40d5c53597fe92e2873be1e351b8
z3daac31fd592a543f79b7891d71044595f72712706a9f47f3a81fe52626d8edcd887473039a3af
zfd7b080b17e719c41d9763632acbdf76bf3ae348da2a3da6a48a00b688cbe52afeecf48483fe17
z1983381f8baa9c45696fd8113de69d699b78b7febde2bbd2c46a156a9203dd3f732e49cbbec1d1
z1f6f90f77b4debf506558bfade443134879e9a35edcfdfdcfa71d35cc4a45c46eee869731aad5f
zd9217fd7eedd3912a02a0bcd48dee26c1152d37403158cb42bb5f2ed920e6be1ad20fa8ca37c4d
z4d1b82908c99dc81424391f1aaf8ef3f5c799ace82167f14b3f4be6f505fa17804d21ce9f27fc8
z4c5b14ac4889a69dfaebe92bb8e7df583dd567c4912ca3e89d30ed6d0e391390120c9486ec1ebd
z4c7706da6442f44fb80a6ab82851c089961850da65dd2b280704c4b55ce1839828c3badd307c4f
za3dd7b901c01b965fc788c02f3f232d655bda6895fec99d474d39ae5cc47c4c81964161c5bf9fa
zfe66b00b48de420abf1f5f4726b1f7bd10b164294eeaf9c523036835112e8e82294c0048ab3865
z7b1df9441c9c218cc9b2b1582aa66b119a3c815222438bdccb080ab78b55322f141de5ce0d78a3
z8040eaf69835a28aba53fcb6100902306b5751277b81272d824c24f89e65c3c7d5ff99266f6ac6
zff9f8e550b1f5ab1c88ae940c7f3423d4c3c4627347c20ce10dda7c744cc2b5c44cd728b490e72
z644fe75841aca69a844e38cd7f586d72079e30bc0c045efc30876eb3a9b8f43f25ba332baf3bb8
z9638ce19790b410275c56da52b63a55d16538e222ae7696a0e70a9095ecf8328a631bc164fdb78
z3789da1f1095119d165088aa2e64ad3e3bf2054f7921bb16da8e80e3727283977fa7c6a6912635
z387ca1f474b97d92d4db0203c74a795147ccbd288ec288a982293e5649bb4c39b31bdf7fcdb0c1
z1f2cc60801baeb06abe085a659f3662d17614674a2eb4ebce72c30c03d33e2c8e8b87f1e06563c
z1fd171d4611d7df6086d7b7f2366d917ff34b2b22236f744dd8cc2e40dd19486b9c52e895cd700
za4481ed512d02283cd3d348eb1adf17467a9e3ece2b499ffa3428bd6a5aca63e6d5022f9f11a6e
z242b1c0907009824ef4c32e7920531bd3df9d28e866244082b80ab786afb27f5b67fedf7654432
z6e84271e0b7996196383b2a4b8e75c74506ce126bbaa36d528b6c6bed8674f6552c85fce03985e
zdbc502b99006a519b534690e79ef66abc346d16f83d7aa81f0943afc80c86991da7316788b0e89
zfa4bd43c33b4285352b61cdd834c08d0e9f5a6574f5afb2254ad93cb31e1dbc3b047a1a8b66bfb
z99ea564262e2439677b44d36f0ed62f87a7f56facb75df7088ad62ba7cc88b76556ce6126847ef
z8f4d3f8ac298ba01c6f43342cebf99a5164d5c46b48615ffe2bb54c30901ce66db01b8cb97b7bb
z40c625a179d1c40d2c62f3f2d50f37d29f1f1b231974dbe58bc02e82c660952ee59e61ed1dc4e5
z6d4b582e2930291c1826f0a17756c1d3d599b95f5a12e8ff4df0d668f8fec16d8b391063dd79e7
z80c12ee1c899c5ceb96aeffa1758d7facc395aa5183a6cc0bc6113bddc2568982e8c59692a8efd
z0569a93a4aa37bc9762f24dd731e0f8ffbf518eef08edfb1d42a10325e92e1f73a7d9d906e1247
z2477efe3c177acdfb038da2287c536d215ad20eeb0b1cbe7625c68388c949650d1b38e34897f4f
zb39892cede6641e2d03c786593273312fa28df78bb2a539a7cf97b7409fe61f59559a1573ab963
z8a0cff7d5100b989366c08754b686b3ec377118a2ce210ae25132dd027ce67c85d39865b855dcd
za20ab05b9fdb10572feacb010ffe37564215e48eab4135fa6e550dffcd936e7084c3419b320b50
zc3744556b4cbb56671d4e461ec3debd19bb9228ceda4088a36bd89b1a7ba1bdd29f6fe4951d09b
zc98a3325f6e1b573cb19e145010619a6fef5b93e8e5960945f88b14d37e298801881c78e0a8f4c
z8ee804bf7b0de02602282ac6209ac52afd4ea03a8d06b16a1a49303503ab803dcee31878b6007d
zfefef1dc120ba76e3c63f2cc06abc9001ea0f13c3a2fa59e778df895e35f1ef09c797fdd8f23dd
z3dd1aeb33c6e1d6a95ecbda2726756991c6c75dec9a68189b823ffb8a092d39983ac5d430c7fb5
z201237e723a6e3895b022901bfbb499b77a913a5d1af04be6454dcca61167de16cf201f9cfad6c
z00fda3a1ea614fd656b69cb30ba27cce2414e554ebb22f4cf2cedeee7972cc26d47c3f5183f86d
z7e0e50e9940cb529da36d32ea5661855e9a0ab9979e3fcf5f37f73f5307ab3ad76265e9e2039e6
z96d60050f504994d38766e31b845ccd753de0fef882ce4cf6122c52720511aaef2921bf11fa84b
ze6bc716663a133505e4ae41228c5e381237ca64e383787f6d45534bef5a7b2140586117f8556b3
z5dfd7a31b24de2d28749918c24e22755dc75c56bb75a52c0c983a656036f4fc7a1e15826581306
z266e2b37f9103e9f0a6ec36c18be879a7b56ae84554f1d70fb46c13ee0278fda25c7131dc29fa7
zf5f1e96d95626c2fac46c64ed2400a37e22999f8b93268e01503e5eef0f47d4811cf19e48ec06e
z1958a94a136f968e81a73f7b0ad1dfeee06b63a0afd824cc9014549736a7d9fd09d59aed91a967
ze74ef1e622196322dc13701d67ed5ffa168b16cd1a9d0d6846a92c85c72d0bba961e149e0fb3f7
z27057dedbd2c135fb9215b85446a488aa98e7d3a36c2e33a78b95ea991809f8bffeed71275fd7c
zec1cdf0743299b770d0e52ac322058e13e766ffbb2904474bb7e4ba09b6e2ae5b5e1028bb7a100
zf3d912c2ab4ed77a138916be77a5402baf581b687c37ddd05df084c22a1d1d29b53ff35ed38ae4
zb23d01f8df19d6e2100d18396b5c5a2b5c0e6e6ce56f1b226edf03277e990b73d4b287469b579f
zea808ccdf9e3bfa878c9c30690b4ea4e16a51c3eceabc5992a6eb710d3ce820e606557db5507f2
z8e9eda8c4da8799f8867afa5a4e7c7303fd42c34423789638659b2659e793a03c30f6e75d4c624
z19e3b286c631fda42a9cebef04a9575b9d2cc80d065a310434c0486353c1e0bfe3d8cedf3609c7
zae1594a71c360867097a1eab178841f734df311cf6816a4a0b5b3ee889bfbc2ea2172463fcb167
zdc3baf70657a3cf90f5561f81b33ab21ee021be9de36df6b25e7e02c3f5fa0ed2a94d0472cbd71
z91099910a89e138cb7b190e3ff9a1e56e85954f2c341ffc90ea9200e3eb35bb7686de56c925d15
z333052720c16bf34a9b40c1ff32b3d1bd1d7ea7fb3bf3d30e80bea969802bb69acc6ef1edf6f62
z7d57a80b8f48e8f721e790d0feca341c7f1746c5a6a39d69bf3d7929e394f7a0de1ad6b356e566
zafa7aa9486c5534e1a4a9b6080f6a31c3eb5b522f45efcdbf659031ed7b5aa184a5cc3e5673edc
zee018b1097ac8d827ac3401dfb1058fdfbfbbe740c48c77587bbf5c7fd77d6330c498ae2889d75
zd55cf473902c67542a131119493924ef4e2a48fb47b2d06bb2f381b61d4ad552709bc6f5dd722f
za2770b658ef1271af26293d74c52fc13718a0fa70ab80524b5dd75ec8aa29fefed0b7ce25aa244
z089f267750c74de8718c3c47b6c32d30b955e0b052430811c390c0f6e39f0a43cef1e8db3a01b5
z998dae71c57803e51b4638c8bb589d8984c928d3618c3b4db1c12304ba3bbcec795c6df0a5a905
z3562e29da4a4b531b70d1bf8b49b21aa6fd026f605d530e8e9d45605b9b00c98fddeff252701c8
z1d842ba1c1f4e61d5a19c561d31b7b73909fae3d4c4577068ad150b51571c518e76f55413562d9
z0bde960b749d8902c776e27af825495cab78cad370ef30781c3dd02890f58771c99bbbc13e0784
zabce6f935866ac43658fc14e2947992623413a162e3747c55adb2a2fdeeac47d5ece8ba072eb3d
zda373b64ee3e762003bd923aaed3de804a67c8f103f7c4fa6c3defbc489783a342fb2ccccda5bb
z07e911a7f0e485fad09d7e1b0888101488b6581bb831eb5793458f597324356db34aee3c7cb9ba
z78c84d782205ac09b09329e7ed2ae3fd3d12cca1ef528d10ba8efeae9863f7d96ee8d2a4492c2e
zed3b83ec814b3d50d12f254c6d4d9cbef9f23a935eae2e06f9c1201e0180d08c31d7404f4f8242
zb02b5d21d78a4254d54098dee18fe0bbebd811704e33b6861ea2288561f26445be6551eeb629eb
z9bf04be6ef4d4ea4da3c0c4afc185bcfce204dbff3ce781b7c39896ab13bb3fff144474bcdf600
z7f8b0fbd65fb178eb78c7a99a3411f9d9d0cae291bd02bfe8cdab247117f071d4b211cfb2ce88a
zd880a8f1fc6e8046ac581827730265eaac431566439f58a720146506f43ac1c1b00fce2d6097f7
z837548c3f30f61f571e1dd88d1f80cb2c889af24b0ab811ead193b68fc5e6382fabaddff490f1d
z5299abb3f37362acb9d28235e04d6fa245b7f337d0b0b5fa121ff923e033bd8f842159d60da76e
zc178815d99eca98c5199dc4f6e4222f54fdb2383910ee261edeec151f2341337688284397a4a58
z4eeb921cd37f869c05085bf19b9e9e1234dc379f92d3ac6834b9ce3cd3cf29f52d6bfb6405ae0b
zf6812cd5bae871a93d4338b90214f9238f5b4cf223b7125cf0669f6ab010b992159aa0d7daae65
z97256955b54ad2e550d81d29018a1a1b68d76e23aa5c0e7990397c5641ef3c503414507b64bb59
ze66753b5f0961b16192132f06f95e57752586c9445eecca3161bd65c5b71341b9e0969391c03bc
zad5a695253c74b091ec82aa368b8ebf05eaf69a92818f5a757169775b54d7e3724990f362efc27
za2ba7aa2e39d44bcc04c7c0892f207460f82a9f5c941b301bb3897b46c34ae2ddacdaf14c7e12f
zdfa7ff77014eff98003fa8386c74b908e4580d655d58341bcddde6b3e99db855c265b46bd918f9
zfa234d74253941486c4b0acfc2ca18d143a1490a625266be355f48558fd3b4ac6d1774bb458399
za31b50fc446da886fe14df56064bfcf1117efa1f4043eeb072f74ada6a9fa97d2e8b1206ea4ff4
z065daa982d381b3988831975809395a21230ac0d79f0a27cb7c54f10cc9bbe9413cfdb24e0b9be
z8c14e79abba8be368fa5e6b65f77ee9ba668d90184ca47534e69ad7a6fc7b75941eea5b12fe244
zc4bd6c6247bc1b918da334e405f647247e4194185562355c7aa40c315dac6742bd76e27766e4ef
z17ce6174b9877a7c2961646bc3aa8b565ec8aa8ca9dc9a5d5b2e36289c7a0b865a64a7a4dbe7fc
z199c194cb35404a05c6dc4e1f2e874ef504f99590b864b79129ba6fad40ac1c0dedd60148838cd
zc3a635b07d3270a838bc728570cccdfbc923d441b23a03bc5fd352061db53484015f4a550f56c1
z0be009fe425fd539dc300963afee4c7a175d666245469c79ce659306fee7c23a5e1e8502b02323
z4e229a979788cd316cc0c3a15858f2064339b89a852d4232fb97c0c1e5e3a256487bf291a206d0
z63b80e78abbed741cb95f19505da922f38bd5aa609cfb358e2de692a5ced3b589af00b1599e009
zd32cf0e233aa73c2ee0fe0d0db1a8b623d7c14bec0c4fe03061c314b6f863693633ef6b91c8a47
zf0f84ba069b4075a0fc3df725a9223be60bf23833809183f440fb658368e0fc4dc859c5e47ff44
z6f4aef971bab942def48ee64d234688ea492ba9e2d0236bbcaaccdd5d7db540ac08b2292ee7104
z7e7a2b65586ef1c54cf1a6a601cb864787769f3f6a4814c672eb220c12e2e345112798ef2ff96d
ze38e58d62f24aa0e74accf4495a05c68216663fa5d28c39a2ce585d2a43402e29372ea05fbc87a
z978bfba87ac5a47fd3a21fee7a634d1d2add81844bb8a30ab2cfb4745008c67b1bc1569ba0533e
zbeba888ee8f8c7b94613692b787d8b9b86fffeac41cd01c0fd616e8b267f262ddd2348940a0a4a
za7f3e09070f482bdd3aeec8b7111da6019fefd17ac4fae52788a8f08e6468c642836049bdbd1a6
z0c2ec6b73ee5d8e488e4709cc5c3ad396de50ac2beb2f52c8d2a9c3db92e82c0bf6e6f669f19ff
z5c06af5c99e7a497d7879c24fb88d96b338317ef0f36fc507dac8618288c08de07f51d363fefeb
z2c0e9980882ee17a5af766d66f14cdfe2201f83d3cd98d3ec2ef19b289b824a7b92d23f810f5ca
zca4d579f0af5e452cda3da395a869daf21b561ffc7b0a18e4cfa7bfd544f94fd5fc85df7cbae62
z47e2b35e6cb576a7fff11bfbfa1eff5c46077b53d90f8bc1dfb1fd3f415deded7577199eccc765
za61f7af5ab840ce1d75b0d873a87cd2d26cbe0a33e4f4a60741e53d879ab0793b6fb7157e98950
z3ceaa245cca8b5a21cb14df76a28a8540ef53a10a3ceb64e14e3929659153dfa990ac26e9df875
z2455a69c72f3d21d2bf104a09791934220a7c5743947e27c1ea19c66516f35cab9dd2b5100021c
z6f93bc12ff5b39888e81e273bfb73a8f5f1c18ca80d591e0ec330f2ea7a62a447497e78df0f301
z8eee4e1a511945f3a96205fa3780056727f488e870b1756119ee23e7f499106e9a907354558637
zf62923c1c441ca02dabf7d792e2aed249b06b179e2f391f3b7b220018af5d360bc50cdafde502a
z22217b4cdd8d3081586ae8a717d8d49ea0cc68e82b705e4785c3546604c72e40a9e43840103c16
zc39f1a83d1ca106f626ad29928a10cdeeb51a236e0e42a6bb855623a0999f278646602a7006ad6
z656b9645bf083cc79a61697c50a61469d04aafc845263002b6d21596d4f2dcdb06c479473956a2
zcdf0ba8a0ce876bf0e7f4bd0d61338eeb1b6b11eea5475670ad5b2df33dca9ca5a371780e7f3b3
z9d39f0861ce7b0ee62dc202b1dc4e2d94aaf4fe5348692621942fb2057ef1159ddcd2fa3668521
z0221b1982b2b19a5948267114253041cab9758ec35e69823be55cce65bb934b537b09efe38f0f4
zbb5819422c7c034ccfbb6fac6e40729a9e6e9d0d2b46498252d8fdd0a109a89afd3cd845ad6f68
z6eb973f03812299b90eef0b914a8a0f8160ba6cacd3aa3140041a593ee58dc421e91a04f9f470c
z04ec25168aa11df3e9ab4eaf42190899bb26c6bb93ee9eb238261c6c88f51e75a5a618e2d413e5
z673fd2e5e0a6306c9e4f26adb3ba45e70f175ea5ab2fffe6e64e8ecbb617fb1dd0b61db4b6987f
z56a50340d2d9d0067a75d0e4f82794f5d61888e476909c50d7c2a55fe1b15fc79266719700e212
zb469eeb5e90d4124bfe0e513f83b9b2ae540e10e94109ecc5e91d2436fac6212113d6e6c15a6df
z661253ae15d5388e2f5c1781bff7db19f3e7cbcb61c3fb528550df4a6dd1eaa58c0cba592067b9
z6b3900227b7af87df13b92553391d9984aad11b10349314243caef1fd85881cbb4be30460ba28e
z7eb6532fe0ecc102794392514a1e397f6ba704f4f476a21c319473d9b65eff7126fab95b02ef62
z505623da8e0af32ba64d35a03fc146bfe7b7d5226fac9d6b5ca1626d4c6e525b75a8badd6dfad6
zd997f7e1ef5a3f67156805ee7efff0e8997ccc46bea214586b8513b75f5d1e0d9db296df571bab
za8f72b0c1e013749f459b03ac61f997c856b8eb68cfa744a78c7da7944399b09933d4bf408f1b7
z030b8813eb29a27c38ece9d222f419f2ba4286180b0b78fed5be8dff79fb6c1eb23789d92ba064
z57c5a7765bab79c4026eafc24e16572856e4da79ad1ccd8d8b29fffee43b10bf721d592bdf09f6
z87c2460667e2f0f5f69dd4b2b52eac27874b2eb8423f642d7e6308701ee5ed1e30986076196b9c
z7dbb9b651c6b8e44ef8fc241c0ffeb7c74d42447419bad151c134cde596b06037d8ae61dde4d0c
zf8925dd4a738e2cc9e9b68d37cadb352609c495c966539812dabd5a52b2fab588c3cb97e9b2914
z1e09c8e714cae47109181b1c3af2450cc897e3740b41b3b145faff2e54641022ed485d2d9d014c
z4b6794bf004097627879cda1670bdf6ade75cfc41d5d5839e76b45b516386d6ed54b7ed9c29d27
z21ddcc371856f6a7861440e7a35850f2be05b271a51a1fb8b445d47767e90f78c92b92b0b225f4
z194d93e7da0cfe02e23c0e5c6b8cf8d277906d032e24ec2bf9642fe43179c7fb1ffd3cdc64bf90
z5ace0728595d4da83859e286d7fe26ea17e7cf6f8b7570e9e333a592e717c146ebf950c8b34d55
zc5de3829d6cfeb4c7ba57f78fa23c7cdfd6fb5f7c74d5ae4230ba37dacd89f048528d38985722b
z68d921a663d1cbfafb55d04f3a3fef49fe454b0275d0896b2b2979fa9970bfcf1ccc923ff09bc5
zc32738d8d999d85bddb53e8f016d3d56d6e13c3a809b12f59f63d3860f38fa524aa81c5d1b0980
z34f5f42945376361dee7b7dc0d0c8bb0f52e5cfa2323fd97fb932634b6b7a5adfe3fa1596710a2
z513f56a970e1d45cde2c9d23ab50d95651117117a4d08db7735af878c4327a02ea840e7efc5b5c
za2fe561027a4181a47063682312f24a7cac51c55e4a56bc37899b3f02ad07f8ad7d56711095cee
z2e0dbd81ba4ebc0e1cf4b23f78d25eb873a00ca7de1f49cd359a5be88f31462990837330aa40cb
z7e243d04bad77ad24716f5e1b4546935a7add1763fe9f5327aaff28f56da7b407180bb5bacc418
z3f47f1b78046447bc7918f7155fc4965ed693f8ec4f0a0370cf82d67449155ae33da7f5b6f5a06
zbc4bc7d51af1c9fd7d87b6c94f6528af36b940691ad77494c468baabfd64dd0008d5737de0bc8a
z03cd9150b3c4f2252c3e52f7ca4f87400e1e597dda9025edebb2ddfde48d8687c93f0501e2d3ce
z4126282d8c7436ac1d40b827ef7690515fdc1ffdc4bad33c5fbe417ef522db2efeab1deb893c9b
za1ccea96d582aae6eb8d09a3abe836b6a9ba5fe6ef1fd3de3824d242560a0a48db2367faefc24a
zcaaaf7a11bd6e3cdeddd7534e27b0b543c3cd98203578671b8fc8eb5b31ad83d3ce82bf511e45f
za38544d19b3048b85dc42147e3122139eb1455a85dbfe41d6c45613d0f85997b69023e5cc27b14
z757df2e43b0aad94c2eda6d33144097be88f878e801e4cc674b1c8019ea8dfc08b59d2ab01f72b
z726102091a91b5b43fac5c89f8dbd55aa436d2ae7bd2bc20f185bb9bb338f4602f0888431a7a12
z69c6dc7b593a0d01647fb2af01324cb3a730880e26890a315e19286c2b3b6da9e0fa39ee4d60da
z36114beb5ac06ef1e252240b3799f752a31bc60a75c02e42cb06a99765b2beb07544472346d6a4
z700a2966f6ea45f6f6b43877ad2d78571a754b76d244c881fb6f68ac94bd5c7b6534e9eb6b5876
z011e52e06453a1bb6181e3edfc4f3a245dd8851b8720d90812a5c6dcdf9c5b3ff7194abe9bd745
z2bbb0027bd622846fe7d218bc7facba3882f1e6bc33a54353eaffd94a243dd3a5b0ac87b0ae7d1
z3bccb731f15517082fa64dd155c3e2bc59c5f11f6e9472b14b2233739e8951b2aa33ed08039b87
z539895cd2210954630524195d0c14647ae49c9771ccd03e48c0aba9ee7e93edad8de926325a76a
za1d8bb548688bbcf95bc7a7120397a74d18ac29c3cc08cc9c87c646203b2cbac03b8833e845f55
zbe06b70ba22b50ec9a433b2551427b53fc5b1a3f681ddd825f46f5b994ffe6131c78fdf240d6d5
zc95a49af4da37065b2bf61003ffe15d068377179d628abadb50682e77f9dc555dacf72311a6682
z2713f75008013d8da7124924f9c1921892fba3c87ade2aadd498d589f100b1a5d7c0b8802ee8b7
z33570c5b866205a504724cf72fb6410ea6810b33627b6d0b0b9d72e3c6d48d4e5779e37dc277b3
zcfb570cc2b13d536da7363f3eb7670a8af3c3ad46ce5ded635fe36b94d27dceb1b418bd6cb40b9
z77d554982df5b36f0ac06ca9d3dbd7c779cc7fd99dbf2b07ec8353a443d5bdbf305b98108f9823
z89ad9246b1703522ea4fd49460756f7bcc184309f1ac36dd4f91b7a30e22fb5e94284f401a5a92
z0e2e2f8a04676dcc2378b11186bea4c60956bd7d6ccc00158a6a641c8de430ae78e2915a9bdde8
z83d3bc65f27252aa76f97185e5e64e39ee02938888a05e116c8f23facd973c9749bb3e9350dc41
zaa1ce81de27fff5099155b4201c2fd6df3646df322ac16227be501889c71a3c0ffa1803203c3fc
z2a847d0a881bf9dc168ab1039f0e8a8fe018824ff4991ecdaa9bb80e0a1c0ae1a60195f7a8d870
z60dc69342cf4423a188da09f8e10374b0311fab9771aac8020af3fa7f36aa6c80dd768aa206d17
z86dca2ce06fb5607f8ff27342743b4116aec2b81385e082e6165e7cae3df50466c3f43877e5244
z7390366b0b3788c5e8d6237ee059577e422aa6cf772b40892f919f5985ffb8c4441248e3fa0223
z7cf0c8c63cbedbe262877155409539e4a06f546293bbee567558373d3a4d6d1210d1ac45315c3a
zdf1766f1cf3ec7db5d942694006f77c703435018928c81bcd8833d34ebb9939d342dd09db228b4
z312110c761f0d8b79aa1595d6c77d57ff286c82476df9e7edf897af9d83f85beb2b07360225935
z42495433f3260ce6252fb881da4413f03cae0dba22e87fa79c8924b15a5382daea8f441e5169b5
z41b9f18c897cbfdc52786a5ea89814051668133a2e757b897ecc81e55591a356e6b5e024a05467
z5a4b0540b5b784b64370c174f77eede8b19abb1e7137d26c9cf5c3010715d3f07b9530cd437f20
za3dd26c67794754fec4dd383027177946bc20e5a108ee916bbd15963718abf86001456f4615a20
zec48d69cd0b4521f6bcd171331f3d638ec3868e7ba80dde045c020eeeb39711dede5ec17fe0271
zb838f3f0136419bdb062175d5ea8a495ee85301dce26a7d36d006e242e401ec574e2392128cb02
zb0c6b4d1a3ef53bb50f4a70e3b27f646d515d9465be1eebb0ffbd95c50fc63a032661a378f03d3
z6cf7cc09736362319b7c62c8e3194c168251edc2324fc502c815374f7d265442fd7dab03e3fa57
z8bdf3787b2e14e20c586fe76d09dd0ecd6e920137139bf649aaec052e6958a43cf10b7f0f05864
zc252563fca6b06b059adce8b9ced179533e59094038f91e6ffe67712bf03f5c736f0e10f5b535f
zd534b325769a8ce36078b0de628c6fc0bff7168880cb90f94d51b3e026017d981fa98f152fb3da
z221d52a2fe5a308eb1b1c67ae336becc6ee6202e65b964928c0ee6df3202f7cdc91554cc73d84e
zf612bb7650ecd7a291480e430d00c79e680e6aebb4bb8b8f5d08d0f14b34a4a5b41dd26eae10d8
z21a9c085229d9a393ffdd07067e3390ce669188e15b04f8e94c37b2ffd36efb1497a6caeb59f6b
z7dce12743c3cd5e7784f757f4f1069961e5d073ce7c376a85f283e11eea6e1b78901d583aa1ab9
zeb83de5a6d1de68b07be148be2dfdb65b4cc11f440b5189330b37768f69cdb16ebba0e50c5de6f
z4420b4e1ad5574f948262a0997150fd961fafdcc0112593e114a828b8482271ef963bdbe4b30be
z6ed24c746c2c9cab37ad1271ac44b6cbf306c907f4bd6454132b3ca171d1e1687b8e294cecd0d9
zcbc92f5bcc4c54e715e1b11df9f11870c32fbd2bccfb31b86101dbcca22326900fa5d3c7e84131
z02e28c4ff9dcf8fe41a088002a60fe4c94e9d99c35eb1fac44d6c98897eb09492a9bd9c7532007
z152b6c63a707e5e7b7bddcd4364510cf169ac6c39c0f8b18e11f9491f86bc075d7b0df1235573c
z891c087c5868b1fbfb6c439329d5896f6671decd087cac26f9aa0cf8eec9872fc58dc7cbf8d5fe
z152b6680c37f7ce7dfa6859f473427adb00ed35b8160d4fcbdf232ad25a2e8bc0888ed1e271640
zb4e3df5b5683cbda6063a4fb553df16ea4c98cfe9b1ce8624b14ad9b1e2546494d5f605ff9f157
zfcc8e5bda4e4ab08b1ffed4f2e49ef6ac3b7814adf638544ffb2d04b74b1fd4b4880a028282ad2
zccfcb55322184f12f0497f83b7f16b31a3c6047ff60b17b75bf9bdf5a2048c95fb4cf8f9834343
zfd9e0dbf466e7845309a4629def844854ca0c2fa47ad9e849506093a5ef29108ae95ca838988c7
z68f65c45b431e28a468b07194db9a9dd14096e2261c118106273ce26cf520a663fb1e0357431cf
zb3005f8e43bad7b82f780e0f87c0a7e60b839a06aaaa098f6b97d68e45d252f9a46a104a8de98a
z9c4ed418ae93c8007722c4628b02ad2da3bc900c7317a5f08847a676d2f27a371deb1bc46c3aab
z23977f0aa74b26fc7c2d15b2039bac56e39330b3106aa462cbb7b6401a4a4deb28c8de689b804c
zc69661843fbf6af4852d1dd5a4c05a8c73d76b9896564bebb2ce6597db94661b87de3443f74181
z9f6d2099df7f56876669400341ad6b0d58f82d0929731464451f8d9047c47c5d154e59f1926e42
ze3560b72db0ed610e4047ec303d2075041f3951d6445c635aefa49c8626ec7e75e4060faeeaf6d
zc83a69c8a53880287fa7a4e91b7c04d046cc5b508fad752d17e5a769be0a6ce6d22a2ccd991eb3
zd8c2868e98f0b080d11d4d7ffa10fce583e3a64a69c8454e5eaffa5e02e73065163ac1f8aee88e
zfedb5dd22ab3aede3188abdc84f31e4540cfadef02afd7763bea3141be3ea8a23df04b1b22f15e
z9183069b6df5b2a32776944a666d408ba7218d05a3ef4fbbbe7fcdcc271a07e5af653db41dee5a
z18e751e3939e08d4a16dc6706c133831d1d3e1a57d5d0d32974b11dea2b052943d9401bd5f66ab
z964c6e9aae719c880ca1d2d293e1f8b45796463962c255e51cc87151409443e65b89ffdb6202b8
z6a49cfded80c5d8f19f9fe6cf41e40085467ada6a4609cd4128e1d60ddbaa7a24facd52265601b
zb8c5e440341bf6e415d01f5a3e6919dbc2d144ae84ee8b847414e1a05f0b26cb833278cc28603d
z36141bc5525a9768378aeee1dcfa74522582d5fdf3d3e5e5ed2b63502179ab199250961634af14
z245d03c5dd5290cb2f58d643624799fb9c57e17f8833ef797bc30492226e7d5fdc2e7c8b8d473f
z9f474da9f5aac196e60e409b64942c578caf79bf13a75f6247c3f2704798f4240e047bc57a06f5
z0bfdff8969c405f284bd6a6b2b7453abe60e6220e9b81683b4969e368b3f55851cba97f7920cf1
z2438d9a390269db17ba4c17b86cbf6fbf2b819d4aba47902124c5ebb8024125bb6c94ce7a1e998
za6c96a67afe10089294bb91f60c94cfc2869a80e823fefece3130afca07b15b83ebbf8eb154651
z13fc4a00c33657db3cc683802bc51317b9f4ddbbebc45d2b8b0a89906e8ae40d6c85b2d12a0348
ze99b19d81639c292e7ca8beb9a3b2927f26d3cd029ce6a145842143e2263cc3d43d3b7b5bbf608
z1f2e7bd62a519d08295232078fd862ede32247a224921ec1e6182e5e1b4635513228c2fbd406a2
z219c4b8a68e3abdfc28fe79840e2f1f1acd518e7962fb002c458a0497593d31f3f4d60253588b5
z57454287960c5dd8843674e15d03708dab21b91cd9540c69b486ef1e43816863c4e2375ccfaeb2
z724d1bde12a2ea32f7a72029e51bfe8308aaf5f2bf861c480f27075a1ebead3cc50cbf9cbc5d43
zdcb150713c3aec637766d9ebbc98f6f026fd21d82b3e3157460df3c46e847f98c328f614bda579
z9c5e4f2814bc0c41aebeafd78896f58d087d32cc01091e1dd9fcd26d47f6a885a0eb1ae68c2ce3
zb96d329bf60fc62d36ce2021adaa3bbd51ed0f666d86ade143abeef702a9672200baf03fc44deb
z20d974b28888e39e1da965fd01bdc1abc3ceb948c6c34dd50745af9b7fd0d71ef13e2222b076fc
z3872ed293ddc26f0fd6df052c23450cfcbb892c59f8ad22e1d06ebf43733c5b1e0d4ef7001363f
zb87f21c347da604572eae095cf82f3746e5089e366e127e6feaa9f44208466379213411729132f
z48a53d644bfa320cac0dcb20a09f06906a178f6a7a28e3cdece10d618e69223dec359d8b7f2442
zc716f93a71e61ab3404148dff82123fa17d7a500848299b7ce631da081ab95f984962f0443de94
ze34ba300df615addc7c1b21338e8f22652a19009dfd23a8c76437ba89390daea5f974659ec157c
z9694318c55e66f62cf56cb2359e80cb3b52c90c401b40e6dc62c0052071af6a8d772cc263fd474
za598205f1c3d8b40f86a643f1775290b7812fa9e137aeaa3894b105d7d1af4096aacca760c7d63
zd963d638a369a2d1fd149349017612590ad4e371e95ac6d24d5d55102b524b79fa244beff13868
z8fad3017ddef13e2875d21d1cf11869328f5b66ad87c970021e1a21400f67b29ea898d3f8a23a8
z804a118bd6710763026e1d024712094348afdc3a49eaa697cd254630210cd27958806e7bb082aa
zcbee796a318f5ae0558ad6d9d2c27d755fe0dea7f372778ec297ef5590c22bbc17306aba947b09
z11adf68d59f6166654cb905a48dd447e5e74304383d15bf4d46c102657a6c195534a37d79de3a2
zaa356a3d4c61d5b147fb755589533d5590d677b7090f3ae4b4f99f3a979b7f47f2ae28c7602249
z9705986b771c3fa51f4490316fab046c507cc66e84fa3fa9d8d707bfe3b512198892cfb5a4091e
zb539fd4a18bffcd01e4716d12ed3a00199348d7994ab23b00106499cbbcf31a4b8258fee408695
z88dea89a2204743836e747590a14a6e81f385767cfa5b1d1ce29a168d9485455293dcd63ab3834
z81bbeb48a56e4d03f95c077d2736d1aff53008c30a3a6e3e9be280a77322f07382cea1893d9b6d
z20ce7fedbf55b0fa513e11630ed4c3ae89cbdc26a410d4d14dc6317d6d2e6350456fe8a690dff9
zdef259e5812b0a7a6ab378b760da1879007974a242963a4d9978dad831f7a9f7090c4d46b54b72
z1c1f310a0289e08af1831611f3b611fa42c89662e87c3e79c612e0351086cde6fefc4d04337b53
za5a782e858d0164a5ed4194ca0a28bca4854b92b63e17167f8cb03823c49dcc0974d39d0d45e3c
z33a0fe25d7c7321066dec8d07a3691d2dfca718563275e4acf21e79c5d810e16399d5f70c9f392
z3e4e408cddddb863efb4f7755805c6bac51b60a5551cd6564592ab036207d41f74146b2f1f6ef1
za65556f4f35e1e12ff096be8a2fad29d7d0db5540d578019c861cfaa6466be454db87328eb3e0a
zcc24b9175cdf5924c517034826054d70de40606a754dacdc1f9ba883a13017220b0982180a730c
z47ac077829c083ee4cab1b144568e6b4c071554bc1881294fb6973030b28d37745d19312346542
z9857e1973198bf073c543904c53cbb3aa1da0c150ae3226f2658c3eb9acf82c8ddbc4fe221fe05
zaf60338506e7866c364f2a8a55cda8ca0fc05d2f1c10f7f86f9ad55dda0c75bc4568ac7f7942dc
zfa90cd7bfb5ba8c374610c4ede5735f368c3ae7207fd68337ef24dd19f98430282e259a5e77b21
z846cce0fe28de10bd7a0c1c482edcc868fd2aac313298ac2868f4ad80d10a1d3ae082e1bd3bd6b
ze61842c77afe57888ca3e9e3a6da7f45a46d48d2eae4841f67fc4b50976fa26052285fbb9f0424
z4d801743a64c0f9b37d7f7c3326c9e7847112dae5ce2cb6a303c33fae581439a484e44525c63f9
zaafc5c05ead4b9c4724e3fe7e7922553ae4a6f408b74a64a189a6bd615e5b35b8a1ce324a7ae0c
z7dbe0b7c1a31fd12ba6b419a00b020d3c28fe7f41c455090139b05e76a392af7c3f3e46f437bff
zb2507d87476085cc0c19dd6692b38feeac45c0ae5e581b286edcb9c4f0390cc12670b74b77894a
z85cdb9901841c1c4f494c9e6dbb62288ea81fc5353892200d765ad4fd9220c3479a45641aac68f
z35139411deb8b9c20f959f305c2dff968a4d15f82d0de0608424945d7ca0b05e8d8b633717f13c
z55c2ca5a2c81d84ff853bb119f2bda95ca035f4f847a2b6e11c5112508065c24e9258f784f0a9d
z362c0b9dce1b08b6129e2b79bb5f1cbfc35fbb439348f24ae72a6d0ed4d4c7b8a36bc55bc7ad35
z085ad3b05f5be32396fffba0bfcf822bd9dabd8bcf9d820bd6622f4bfc84acad9bcf408f1deead
z106d1875cd771e0d6c20d07c3b3db44340d635f28b5589bc3d39dabc1849e6a578250253bb5943
zc2a16b824c19c2378c8607e1ab97be00532e0cadaf13ac98ee6451e672181b6a18f5287622c0c2
zd20cf818bce0d86df2cac8801971e107e1e8eeab440ca299c67573c6daccc44dfd5b06b3d94e1f
z7d2b4e7a11498bc8a9c90cdc69d86cc81c85c6af197ca41d60ecb82ef5910ee7c86515519a2c65
za89ea6dff6bff678e8e4b195c4487462005282725e5328d4d69582b98b3a2426151f02822d81b2
zdedb8626321cda5002fbbfc4926e8f13475b67da847b3d190edb9cec23244661c2688d60317bad
z8e481853ae4821878a4900d0660d541379cbd4b6b22317a66da3f1b80c8da6be8a3aad9b5c4397
z346286c2f3dc63bdbc9694f0c4a4b020da2f1fa107c1a36e2aed824d3ae2e6d652568172980df0
z08f78b939f3031eee9610d6bd5fd74dac15b9d2bc382ded99a3f73785ba9932b8ce2ceb204037e
z3c13bb5bd98ae273efe27cc47bb016ee59cda0223b84b767de78c1b899fbfd9f9b0026cf92d9f0
zc9cb5ee816cb8d8e2b082d34159b6709028475f88209df608b33f30f918ce76878ae0084f483be
z1222648a8e2f38919d6a6f320d51b844df698c108e2ed97716abce9f6bdb4bbc56b8c29dcc47db
z9d715c71d28c6036bbcd85bcc955d1331b8c9a96187df57f8285bff9cbca629caefb9b13130adb
z5925ed1f24ea3b9a9a83dd2a732d825937d7775d52c1850051f766b9804f7d32aff6948e13d1dd
z36ca3e375d2f28e8ac4b1864cecb74fbe27062182b70b0a76ff9d492ae0e563efb790f21d1de05
z2ca9dcfe6ea88aa53e3fe0313784534d34bb1ce89606f9eb1c533bdbcea66197a9886a77354346
z4762c7e176b4a99831b338d98f2758eb4244f7eb94698bf206bccc46460577c71397c9e8541ffe
zcab49a4927de2e7f5bccd45c394e003be1d079738de1c50e46a38862020770a1109a372eac2f12
z41e6554f9daf9ea240bd63458a1e891c9d695565d5dadb807d746a81e5beb044c0101fbc0ed831
zefc0290d33e438c711ff49b6520ccead5867eee20755e43f021093f3a303a2ee68fa2ee20fefdb
zf641dbeb7c5f7b17374ad3c74068d82cb4be02664be4af06b26f42b9def4b7b44fb4a1d6a1ec80
z3dfa9c529a3da4471fcd9b704ea7602b479dfae1f24c2c8d9503e4f861cba46f25e14fbd472a94
z65abedd472d3af7aef325c3e3dc6fe554690888c4755e3aef2117db59aa78ecd7018832263d423
zf8ea37d822695107ff416bf84a074a441b1d1b5f6290e6af8c28414fd6ea10cdd5cffaf16245ad
zbca35536c8dd8c0a46e2697a740e327e6f6acdef294a6dbc335d7ec3d707fd85d6f976026d47b0
z64c12837d35a58dbbd95757b57bf27cc929d76f9593774987a0745b4bab89e84f8338b2a9d0ee9
z7941c0209aaf378f3c5e1bd3ce1b411ee51116b10b706f5f2895ce3a37181274b2cc54cacab79e
z9f2a3c843535ce787297d30b3275dac53cf22321b13b6c17fa36fa154a1a4bc29aa975ba12e0af
z7cea4ed64e0848e4d696fb5f7d98b25d8937cceb509d8bcd52d634f66f7b5e30e61c50f93fde36
zfd3dc95c1463023d066ede7dc520e3b4b610cdbace56fa89df2ecc0943168e40786dc804581f64
z5e43c7063e47ac0724b7f71bd2390c221f9381ff6cc9a3970f43afee63135d361cf4489bb0da8f
z6b167eb9b2772b19e37631587886ec5fbf0a9483f02da932bb6baff27cb6be11972aad99fb0f50
za2c4493b2d49e5a9f5ad34dea74d70e175f810a3647c6ac5f42ce7a594c52deaf5bd76fc3d2f51
zf0145326e9c8f70677f0ff4ff60953f3c15f14c5803b74b4611e590bbea2b641a2459fa6b0099f
zb79cdb3e8e73f9703db9a51eeac6418ea914488a81db641e585ee7bb620372c0dc4abd0a8f2c53
zd76771079df248303eb383f36ff9739258f124bd877ad2d3310a9a9cd1698979e023cf2d62ba1d
zbc1a89f4cf3d30d7dd8d20d54b83e9e9ec6819a12d7950a4dc258b77116b1970ed99ad604521ed
z8d7e5c85ede70b5427ea25096fd2de8562dba4b080b1004384b857ee554a1080efb9918c530a4c
z2714caff5bf9affe32d70f7129e3440b6e93d86dbe449a22b901d56d32875e97b1228e60ff44fa
z9e6a08154055b196d79ddae33f5aba708f94127bf3759ca505d3b46d10785f6dd8e9ee2444db12
z84925c4f9544ed4cb934a2a86171d04eae88f1bcf3e0d4febb0f7f52a9cebc7f7f2f2aedef32cd
z242b7ae4eba5f3bf7324fdcffe9a6f44a4b87a77b52a768345cbfc4e47e8962e069e1e337ad785
z9e2a5ba5f32cca405814537a3ac71aef2d8156db6ea01268ce2011a2936327d2ecbe7263a05b71
z79a2769c4ca38782417bc880a02afefc8f92883e300527c405dcbc8469ae468987bcb7c670c300
z5876f723c37524e11640ed347bf93ce44d1d5fc6cff9ad96171f62f048d7e96ef030ed8c699043
z778b6fd4fdf1a8457701cd8d41b67983e2dbe6d9327c231550427f1973b11138236fcaa8b66854
zbe027246ba9a8594cfba78797ef5dedcc6d44dcd167415e0ac3b7f7b722cfaa5e23ae0c944a8f6
zf17d436685699dfc72a10d47a1fe8c282e5524b0fe658e479513a84f7bf2533878f5eca272c155
z4cee6cc8ef99dbbdcd77866993a726e91b8e3ffe9a777e2bddad477d4361c76dcd479d7db538aa
zd936b2e96a1a3513d9d61c474d03638b502b57ee82636fe7dfb2846d2c095c7dc5e7d8ab3e4847
z88bfdb98def8cb3d2dbce4db2a46f585dfde52d3a052c6bacdf4fcd8c7907f71bf0530857f474b
zd69d868c4efb8386c7d2145282f923603617ddfef68e6ce64ba968dcc5c3bbb472fc325d67e554
zb1bb1207b7bb4771f10aa83ee05b4c1d9f416c20d32a792a71a5cc961650ead2cd77efd284bdd1
z9e7b48bbc5d4ba4750a06a9217f0136874f898f2eb3d8ef4ebba7c159a1fbdb96f7f21c188a8f7
z770ab8382641f087ed8d369e934495112477a41710b6f2177938c2b198ee72d9aee9bdc96e65af
z02e7c5cd23b78d17054b776ddc3ecbe2cf523ff8c2dce9190670b4078b341a6015f4762a086c86
z800a4ad627f81e4ef2dda11d5034f7666a5775e8f2c7e5575320653ae77a8b0b61fd1878978365
zae28b05981caed78f81261ab6b41dd29b620b6ae0f1f17121c0f38f843d4125e52a9804e078226
z07a660581a041d8c9012543890a53710e99b3fb3e400bde66d844d1312e438a57b6daa34711aa3
z36b683e26f2878fe7b5a2f86074a16aad153b0e331bb408b73a0122513322382c0fcc4ff5823f8
zb7973f2842c3e5a135f69d391200cbebef1234a09b52161c3e19500e37e3e1311a7331023dfacb
z045468c4ae3f237c1fe2aceca784ba7e013bb7ac1dfe8359a183d5bf71bb9a689657b3c23c6156
zbb8721da7a9deb28da7e3ee156c28b47217ca7a629d968ecaf8d0377f92bcfcaa43c4006006aa6
z230c9d4c5267e30f5c618b59afa7ecf2d5b6ab55116d841452cf231061e6f181e1b1dedd0824b1
z9b303ffdd5b8bd37ca2736bfac857135b307dd2fcb3006dbc3cc5fab2b55a8a070226cc6ce8a07
ze6c6828659d0f2469604c32f8717dcc1b73c3c27a80d6b01529821744873449e4eb94e75a33247
z3a005537e02860298249e590273048c296aa8d3c9ab6751701039f6416adc70b79be0b13727d01
z64cc5a79937afffab8e4c0a738c3000ab4edf6aba6125a3187fedeed4536a301e5ac3aa5c7728b
zcbf56f489820235c096988a84d76072c8d643e002d91b2472652a0b798eb58fbb9f38387517e04
z7a19c97bbf8aedfce6b7b8de8b0554120d9750cb93934b70da08b60586913794b6d4e48fbde9f5
zb7676367eb28b4b3d15841006d3b0245941edc6e8129ce71c5e8391250939c83b0882107681f88
z7b5e4a7a867e6c067f75412b5cf87272e44ba9d33dd5cf3fd13efa12756dc13f44e427fb3120b3
z29b36779e6031c350e537a0904b7bfadbb0e428f2757861154681ce807f84b5536a13847839012
z46fca8c45b8e31b34d943435e70aebf0f8df65c44139a9c03d3c03209fc52d4ccfba5243ec24fd
z9af812de8b21939df0efeecf75895ffcd4e8b5cc769970eb33fee59b9167eb7afd25d038c71eb2
zf1a0f33e27e5084bd9ea05dcb7aff4757c1c7a7a5a91a5b9f31b17e6418a290f164701c2b4b6a6
zc8d391a6c4ae78907f1d8a139d21bdf02c711fa0453f8bb612cbfb3734f5bea02b4d5148bf2faa
zc8275bdf3a664bf75283b9a3593374122b723b4d7106dbd63846348af5403740cd33b44558465f
z34346576b9a87bdc6853441fbea2384c4bc6171e271840c1379e6557c7c73d78e806a94b83773b
z7571e704a69cafd5cfb652f5840ce97b46b522e711b0638164fff0ad466adecf8508fd6c218ea7
z4400fa8767383d6919da2a303346aca66fdf552c7b4e30bb46f8db2dc9e5f14a5944a9010c0cbf
z99e44bc22744d71c6194acced19e8d076f222ffac16392e8761e072ca627920abf4774633a36dc
z390cb4743e3b5297a4f2e80d1af7b6f9ecdc69012aa53af946806c592fef31e2ecc3c8e9e8f9be
z6a0cc1a4437a837bde95698d3e5149f8728dbbed5fe15bb41853d8af18fbd6ba6a89114832b35c
z6d466f23b0abda852df1ee10fd6fdf05d8fed241d65d381235bac69285857244f044720b2c4b53
zbcaedb1bf1cc6506b66eb64a6cd8ae3a6ddc30007631d562650c4a7e5cea9ad94cbb5c7e19f18f
z78bd3314fe8cf1af15ae8b0bd9d38739c2c9f8d0741c663a740ef9044cdc588b930e1e4ccc4012
z4cf2b8b69fb81ae155ce025f6dc21a833aada90a953fc99e8197e6ddf0b57fdfcc3a32066a0f1f
z950243c2ecdb276a4b37fa48fb00271bccad43bd4913d435b17d72c656dcc5242d9fd581266470
zf08c94879ba3a3fe8a97261b690c526898ea0d082127088be9ad609e2b952cd054f6fe8767d49c
zb2194ec2984cb8b708bcab6334a0c4c0dc64aacdb2e0b101edada93c9cef00eaee87263cefdc64
z40aee7c449a9dfa882d518857396f600731de8721f6261a28ad8faaebaf5571c3b3c4aa076d6ec
z72f7a7cc1323a9c488dea8edfa788938eb48bc41f37c6b8bb911c8477b95845199a984572ba460
z9b6e993655f50203ab482648f99d7f0988647884f394c36f2465c9cc639f2133c17a4ce1abaa7b
z01b70dc33db649ccf3afd942263ae3f98ba51e7854db9126e99814a78ddbfeb5feb95007b9118a
za730c22d9f900d69458a4b676d1d24377c2f8c3e42a34747a704879a33692577ff564208669eb6
z2a843ce9d0bdeb09bb07229f08d9d431ad207a60d300b9de337ea828b08e951a2adafe4c628e6a
zbca9b663d802d3aec79e5d698887b6b137e4f98c8e65a87426ba8515034bc49dec98dd627938fc
z31c84dd3d131a68df3cbc69de006b25232a5749140930578a5b850dc05a3bada8f910740060bdc
z3797257ed3232d43ede0d6ac66b65d191c562be9147881bbcc857f486deb2649703df90f7b0586
z58f7e3413dfb02a514ad52df14a13345a94d2a831e3fe4f82f2a36387778912d8124993620c91e
zd613a09060c043c90049fe3d8ff81b0c4764d3b73b05dc90c972c22e3ed24a5b425dd035d83d4f
z15457e7b835479ee554924b5ffe059b363b353e8437f7d06ebda4ba870297376453a93ba8d37f5
zd49aea2e0940e308051258214aad2af2f38d0db7385436d0c1054dcc60e59a8f3171f8b7a27536
z0f40167d1c497bea65692173f87d80f8a2d514f0cb9f0228c1ada4d0c5aa164d30410e721c00bf
zace1988d26a8483e94dfc1e9bcb9f1c2157843afb568ee834a227e13fe4c65be9e0ea86bd60776
z4c92aebbc6a85a9f366e845e453f91877a56df7a589d43b0536ad668b08fbbdf0542d1e3a44032
zf895ec50d943f0ac1b5ea0538549fb0148e10c4f90042a0a051ad9e7eab928e0735816ffe80f87
z1b9e87249ba0018ba54e248967dee6ec33ce394141e8b7ae20c87faf09c2c2500023b9d6b2436b
z75592f9b0c7ddf5a22b8f2705b4289d0e67ce05c45ce4b796fd51cdaa3c238061d437ce9e6e387
z62beaa34944c222d7d99799e843beefde68bfb01a6693f30f398e91f705d46b535ff99a9237259
z3815bd3d240519281a67a5f74f863e27a124a9088934de12ff3976997af1698474851142732de0
zc26623d54bf5e02c3333597188dc82a039be6f836c617ab8c6a344fd05875447c459599b8bbd9c
z37702c10c1f863aaf10d973f49e4e1cf8d2e96ba51d21d3da949ad13a132853e4260f2c8cc7886
z2197c87183d408029ec5f0c78871cc29712cb785879c939e0df003e1cf7eeea8d0c6b05be406f4
z59b629481291bfe31b51c289c1728d3978bdef739a88d5eef71c96f6a5bb07f13517637cf3339b
z6fb487862d77b68b4ebcfeac89a24bcda2566bc8b87a9415005363c0f959a068bfbcf66ec6864c
z8d352c9bbd19aac2bbffb2b13334c17fbb74b01504b0b1b009fd7dd833c24aed1863fc92e87a50
z0af14bb793c1f90ce70516b1e44f39ae975cd72e0b900136181723dbb7db3af44e27bb1dbb8ab2
zac22a70ea0ae4a2ab86b05bf554f04a3d65437420aaa8c25602b5c41efb6da9fefefc123add3fb
z1bd7abe67f02f1d909088a98d85191e17cece5a072c68191d0d7f9e2634a6597c37136fe0e2862
zca67c05ad9952c1d9e2a47dc3591e8d133bd2e955787aa101e4ac5ef61969bd20dbd07b11de9c4
z4da37c6338330b234e0ed62c9b50bf8630d8b3fdb7dc80e7c49c9f313c544027c4ecc88446906c
z89905d43c1da611ff9acd67831535a66965b2538783e9bb85c1ab2e78beabf2b0e5dc6458b2f4c
zaa4a1685d3b75158da6ab700b49ea0fa195577f9b22c029d391c4a73a79e09b90c25dd8c367c27
zcc9964811e255249429befb06337bdfdab8bf6263ed98aa61df25b14a4078d029ca12c43afa785
zd76c5a75053a75cd033f813011213b6c9af9b846c61ced229748a304642673304abddb3362c22e
ze110d34f46f1f28ab34da334e75343022481b57102fc2cd297cfe6de4cab4c87afd63db7918abb
z9252481fd16f92de8a71a56511ac94af24a26e3cff826d66e4869664dca60cc83cf9e07d517ef8
ze5108ce34bc86bd0bc2c66bad0a1a5662dfa8a4d7f2018218dbc20710064a796ee771fe5c65a51
z5fa5b6cb4fd0081c823494a0f89c51738d6568556ab766e0c746926de5695a72e811bf27e912fa
z3ff6461e5d95e57440e361012ce9c71b60ff07b9b7944bbc0925038f1f3093c54d7b0bb31b876f
z0cc94a44e620ca26c4b6f18ffa2492103d2f660a614a3434a4aa087abf3d9eed043690e70f039a
ze09f0fd8f1c342460e803020d71189abe2a6349e2f21b081a57b83c6e603464aff0dee54a11989
z02b3275d6ec55475701417a21756dab702957266040aace0b993a1779b025ad9db4eb005b964f7
z081ccb66026badfb18f6e375237ba08cf8fc79220d2a015e4e53e972fe0cf46021e3180c1c8ea2
z4a61afe43f656afc83b253b4cdef41a974675d8e4037b61786382fa6ac35f66118b376d6a78c0b
za74a24895b4a9021df4e4f7351852f69b776e96ac4a34c67124d9801e345a974176b8ae2ab2102
zeee6cd948a30313de5fdae9978c4cd4a4dae3616260f021dba64029f7a461e55804d00ad733f2e
z6559572393eaf2223b71b7cbfd4ec034b6e889774227fd614e57e55eeec0d816dbeacf97040946
zfeabee3c2c4bcb98fc7814f9d6bf94fc9eca52190010131591d027db752543b6ed34313b5503bb
z8d7e0edbcff38952ae012296a3cff991ec904f679840d3c72fe421f8f338746afe0dd007881fb7
za4fca6fb3108e3debf0ca8b09ad69c54446bcb4f2bca69239f2ac98d364f46e10aaf546cc9ba3e
z48c0fd67c3a68c7c47bb0add96cb971231d7de208d0a05b0a0bc5150f377a3d747a42f6299d90e
z1d36e60773edb60b4ac383af0f941eee2489b21577c956b60219e590856d9ac088effdee202c64
z3e8fa5975ed0cfd131712dcf73a0e0ae9a36461e7825fc75008f76fe560dc563fb1613ca427178
z40a7414d665ad79ee417b27f5234baf672481e23ff78d957d2d93c5a164f9470513d5117084719
z57c73e116f3197f0d947c5032f3a486dc065f10ee691bd6b78876b0535410da4ab37e9210c5b60
zc4a45076f8dfd0f1b4688e5268423bf6282c2cf903be8f62da6287d2d9bd84f400b703b164b923
za51a6bd1da9d52390fa612adf46ae29926c00f8652e35831edd0ea4ddae9141f26da57402fd67d
z9a28c2d19c3c879ec149b8647381f665bd988861cdcef7cd91bd2716169e006adefe8d42a3ab00
z83af82169edac71850f8f47d4bcb7563e7a471b4802f1a52de5d6637c41fdb70dfb7c97b76a265
z7ef857cb2b411b749ac4b8eb7b78c370432d0622c1f9a07404419d379ed34fb94dab9252008a05
z46845f5de3ec2d598ca3688a74ed1111a624da7fecbf81649279fb64564148d9d70869e27de0ea
z3294d748edd3a64af49ccff48bd107ea77e9f4d45da89a3375240e4d1a9f2d5b7116f99ef2e1a2
z84bbdf1832f22333bf98d6c6db9873a287f87ce6b38c7e4b7e99afb86c8f195f90ca5e70980360
z0232d53835d56bbf5c8f1572f55c069b1c91d5102ba10a284b088655394f6cf8745168da6933d0
zc9682bf392f6108ef21465ca7c4fc1e17fd9be5a1e4bd98ee12c881c04583cc604f8736c3d42a9
zb65f26215346ac6c4721273384c7b378c36ca03517e3bcff4ae1a0b1a25a58038d0b53fcc2b350
z67d43b43e11781c0fd5971a21c543f128e2ca905f0b5b953ec1929e1b85c19fb86d0591877b19c
zb9a3751f03f12e21eabc05e2a59aaebbd9805a3397f01d5999a24620c9f08853ac73c65dc4c2d8
z94170f0deb0918edd91a22baf8762de7b519209a058b901392bcbac612674572664597fcd5f252
z7d5733a4a3ca54d65c836c0063617a6cd92e537ed7230f09faf02047c04f6a45327074f79575f5
ze3f2be3cc344672213604c93d852792e2d7840c71a710b8f81d050ab1d168f2af2c5c854b4fa85
zd1143e053a86206bb9e1d7c4cebb8d60de0eb308df3e01617a33868558bc0f0f07742d5490f59d
zf7dea367da1d3160116c84965f3d51d5b885bcb7e07a0dac2b61a74ad466514e9676d64e47431d
zbda8bcdfdd09c3c92a02b2e895801147833df2a24b9ccbab15ed123fd944a8a9edec7b9859ed8c
z05682d18bdd8e055474badf7b9abe77f79f604f799f8ac4c0d277fb90a27e681c52e65bd631414
z0437ea721c286a990012db0dde063af11676790939996f405b7c12c41e1b1124d6494f901e1502
z037bfe53a685133f586d72f892ec8bd37e6f4475f489692380dede2bd57a960a9a35e9a1f0b99b
z24b733a49ac57598ac60b7c944e514133026a0d912fac7d4bbf44c552758672b98cec98b3324e1
z1d9ecaedbeffd7e40de4d72d6a20dfff3fb8c52209ad02813ec65d65f3a505acab7ce7456a00ff
z2579b03a911e559067375bb9e82d073305f5dd667785a75d91b25ce2e883ce65d6d3dddc9a0a5c
z167da5a4f27bc1fe7e00a7928a805c50ac5cba00426737ee8b69b12a848dc02d53e29ba1ae312a
z32cf243e59127ecd2cd5878a230441b4ea3292addde38ca43e390a2c3ce2e618ae840b47e5cad9
z624f5d1eb720c1235d7e4ab83f234fea12e428efa83aab184637a0290ff75302de04c08c6905d2
z6517c0ea47f8e85865d7a7ed446485f24ccc955caa484c165afaf916ac2b5b1268bc1cc99a9299
z9ae878b657b58a4207f484110e1a6d3c69cf9385920d2faee421feca72f1b7b402880d864e627a
z1e4f4b9e235a8b271461fc98c8ae87d3cbf2ddf25cace6e8794321d89be6d1f4d6d7df48a1c90b
zf740cc8efc4472071d42a00b48f46bf31da82544bb5faa7e0731a6be29bbf36ee8e3d1911147e6
z302f574df64973468c2f06d36ea3e347a267d54d1b3f362fc03bb3e531794cdf47b2ca924a084b
z0388f06234ddf08ae984f1700b8b5d980dcab88ff3d9d15d957e066608ee942b4646ddfc1e1084
z1a4876dc5016644747761402d7e7f95e8fa1ab522917529050b16c7d974abe42bb234e38e2ccb1
z0e1ce5c0767845eff8fb55431625bc6fa16d05583724cc60e1fb8608c9b4fab8594ca73462ca6b
zad155fece1aac0b55b55444caad40ed0c96bba3d627bf36b4883bdd45c38cbd26579687736b838
z1bf6b852328ce5842a08409c1d0fd1c3b85d2ca2c44595452cb1f6a372aec13c56f6dfb9a4d7a9
z8528d4375800a797dc294ff393a6a7f25198742cc0fedaa88f259e9e3efcaad43a6c419f49cdcc
z4454cade47e4adcbcda71b249d890838e1082b3c90b88186732432a2f64b216749fb2b59e2d35c
z73715e6ee25ccf792ed906867d8dcd62eb4d79329321d5e951d9e15e1152a6ea8fd7cfb58a8bca
zf61af611b851123197038d2b00e24b9dd939f51040cb8bdffead395f31083a8bcb47cbadb5e652
z646876f87aa5d7384e613536e900958eb6bb990c7ccabbcc1c701aa475c44ca90a204f0afeedbd
zb0c6e827d80cf46f1e47383000ba8c46cd4411bfbb2c860653316ca89644ad511557d433a7656a
zc571cd9ea87a3e3e5d2e998c4603c8c13230fab1609918ab600144812adfefdd4f681c4ab4cf2f
zbae4bdfff9b830b97e21b89328928b6b0d8b96637869369c65db029c4ba305e51fe0c8d53d2be6
z0c499e1459f6d64e465e6d3c930306873206b03aa9cc01228dc7b3d510d08a9c2f2eb10ec68153
za952f8e0ed96e41af27460f1c06c09b8d3a2067613602c0358106f70c07ebae7e500e1c8734d1d
z052d80ada6a9254ab8cb43b764d09fc64c824d215763c657534d40c745225d5fd3516cb3bc7051
ze4fb88ebdd5631a5663778a76d2efa21c9cd98581d279c34358896cc63b4da43157cfb813a0d50
zb9ac1024f7776f69b22b44cf36ec09fdbd7382ba92137c37af165d4b234676a8648d942d9404b4
zcf5158145ee0affffff2ff6f36984957baaac55149cd331ee013c003753ab3abc2426e92e8d4da
zfbff850d2e460e1a6dfe1cd1acd8656edd7c050aec930cf69b0d56616d61f6499be847d1d6f307
z1d10e4a38ff6601b13d6ab10d772a5fdd06c5875ab2128d8a2d6c2a1f3ecac85bbd24ed6bce249
z11e108598e790fb85cc367e2baf2f5e45d2f53f5be726c82de00bc1463a4a82561e8914dd41de6
z6f9ee14ccdc899a3b07915f9e25eb136d817a75932d7581cb9925620ef5c3467bd8f0d0c93cee5
zeb5844fcc06007a355a3327839791d63f2f83f3832355af210d5235cbbfa398e6b77e3df15edc9
z5b447f96495e1636670aa4884dcb91ecbce8df496ff259393fc30bfe65a1d659c63c97b908a569
z4da7a1ce993507d9904f43d5663cc4e04184182abfebb3da673d67a191de84cf8520da3b4b7b0a
z8e65ec1ef68d68a2856b5765794687ddadc3fc9552db3bf00de443211163e2131b072b5425c761
zd5df97e3cb32e9a5a14ef87f6dcb675bc9bae6dcf485db0c769a00407b15dfdcb8817f33ede735
zf243f30f3572d96cf3d7de887342bf383211b30797c1971423c7c3535330947e850cd7d2c45c77
z376fb5886fd80abcee7b4813eb7b24986e26dc2ced2fd12915873c35091fd07742b9e9b668ecc6
z2af67d4b914616c847fe12637d2e3fcc8cd5c6ea3fcaca9a222de05c304a1677d44138a1a203c2
zfedb38747bd3e5aba9f61a7b8e7f131b6a8cb188b919fbac88c81eb2c3e0d4b532f3f5ef117078
ze1629c5ea300ec89bdca22ee6b6695fde210074d424862cfca58bb932dacd01b5bc6c2e3f4e58a
zf32b117c583144e63ce05ab43e797afb3f9871993221c8d212998ee841c2d96f099e6e40bdce18
z950c3a9ed6ccc22de043eb9eae131333af5adae10a45cb8124eb4f73932f1d63eff590f5f36a0f
z60cfe7ea474dafd460ed3c312e12a616ba5847d829d5f35164774663f4a60eee8838fdd38630e7
zabc7a6341a7fec91716a8b4f6473c53d5b6bf7d1bfd8dcfab5ead9915ec89c946a6bf20e8b1e73
zb693785fe49d43ae9fee62d5fa665f271e5ce88d2a4dcd0e7a2a7e4368ae1cff4b9982df8524d6
zf186a62abe2a48c197b49c06280745c8406fefd67f4ad4e280b59cb79eb5e8cd78e6644ada74e2
z662dcc8836077d60fd29416fe7515bb598796a672ebaba35b617cd03b5bbe0bd8d487240d16001
zd3ec53ec6c13949c867794809e97a0636d1da057f8c7b2ce0dfcaa0634a73496cb301cdc68fed7
zd308ffd2009a4675634718f5012b0f7db42298514a8ead1aaa356f361730e20622bfb8e3f706bd
z30b02de0b9a8444c1a424e4d4e65218396b89bd3b88c6595688a97618faa695cce188446f62d36
z168c21afa062fb7a781e0f27c0fb3a3178128446010b3a21245d04113c08cef8f1db686ff7ed8c
za34073525fb9cb0f5c6b0d11dc8bd0da9a0c22dbf62bead8dd514cbc2b46ec56599df3de193397
z728522b36567eea86b92eeaa5b1e47bd49faea26566c1e4d36d44921434fd5b53da1bd764d1d1f
zb0a14e05e4a773f59e430d54160f7caa64c5e3c957558e533e85d68e2a6811b13ef221ece43a8a
z9d9b9eb606234e9e804cd3979f70248c5f4f4600aa5cc847baa6f07ca98628c0d77c2f773dbe71
ze61247e0631a56664ef7568e7c0a83ff58fb8da5398fa80346e679cfee94532ef63b8b68934a26
z757b5d8bf7bf51dbacd59d3ef71c02de44fc28b12609cce8482e8f56cc760819241cb4f27c06d9
z0d1e0b62b0da67291a536f0b1c3b4bab8e7354f2455f50f9e73fffba6a612112cbbc83c59da9d4
z3515c63ca0b722afcc5dc66669eeffedc8914d5c5d336dc9aa5f594c5712d0800d2c06d4ddd07f
zdf177531a7abf4c554c43d30c922e8013e19de9a47150d4d866c63a0a9c03ae33155008f205bd9
zaafda8f088a37e869f95ed6c059eb31cb01aa090ae4900045a9e749a4397c2ca86b3b2d1fb7fb6
z4238eee07717d06cf2ad19d18acb6c25a573cbd5dbe850ce8f29910315aac836a3d78dadad72b8
z40806e9af6ce29785ceb6a07dee5317a5ced6819d9d95e95e23bc442d4284ba4786e4a20857ea4
z278598966a25a99f1e3309bfd787ac75d7ac7bd544514e5f8c371fb0349743d8cef5754861ed3c
za90bcd32e0e621e34cc8c2e8d683308e0b2a197f040e9305a35ab899e89a375a9a317fba7d6c17
z7bea1e21182d3712ee442bf38cd3e974068e78263a9bf76c0297732f7d4f48b51c8424d3720a6c
zcf844a025f1e8e7dc119b4e554e0153b8ba97e80f020c5a5d8bcfb4e73f9debecf529f5480850e
zb6b9be8413649fd8c44d6e47edd4a03dce7f60109a66d0acd7a365f3e5f58d3f502b3c3cb4337f
z29d362380227987eefcb2532a40ecba9f62139960c172ef984123d935f7f00ae1c7bd3d1d860c9
z296e7e4183c1cd3e6b900e1a7fa0450b31b72b4141e0098b8340c66e4cefda14aeb3b60669c97a
ze07a51f3e884b9c9459eb3c857d2a2bf7f0945f4e70efc7fa53181a120dbd1a49fa9f6de41da75
za451d154260d5dd9e60d3082281f8ddbf5bf4e6169411e5bb91f31471b3318bd01c307240c7ba0
ze32bf35e6c8a5a1d6c73db07503336d0bb02df1e1e2b4f59c2c175fdd33ae8799e3989158d9d79
zd915f9bcb45bdd24e412f7885c266a48a83d0c6459fb5b4f08da282def847ed26bec1cce4df5ca
z737268692418b9e2374ac6cd0226a236f531063208f625cfdbfe9884442e4afdc50c1233651d16
z3b4f4afbef0244a7a4f4acb208c9cc01f7cafac395ab1e40be6fd10bb63f3aaefc742038e10b1a
z4306003665f2c094a3d690e8fed2274c43140ef5b33474b332583f8c93440270235020fdb5cf5b
zf1a8adcd2f37b24e6b8af1d336ecfb6fc0d3ae75229bd526316f825fed76d4f0e61a848a8f1da2
zb53b3e5b5f858de52634358708bdd534606db197952881905edf7edd88a436c8979cfd96519bfe
zff13829f1e48ca3aa4fe3afb15e5e0f4f230f9bce57e3019618c3bfd619397a4417c30c08fafa0
z9358b6b4fac8a1be5afdea127b4a88697c8c192bfd94b96b93d2d27d3076712cdedd5a491e6531
z4e8383a20a90356c9d2e8cf74e0e468d8ae899cd3b0bdb2227d83a375edb745c04d67a6824dff2
z62fa650fe60e1ce04eedca5b56783c735110c1fb7dd50af1389f35f4dc9e11fbeda01f1240966d
z005eaacdc0c627656e93f01abea9c0c4f5e2f18f76be2a6905f6376a1a471b1f37ae378fca9445
z75fc81d86c2ba1f01df218545c01841df0b8a5a19a948f357c739f3e721b420ef4aa0d86a9b043
zb4a6ad4e6757a2593ce446faaefc2decdb7ef93df9ff4eef9fb30651fc6ff869842284aaf27c8d
z1c7dc65128378938854ceecf0f7e0bc9ed5a38e4bd2c0efa89098c81722d90eec35464b59c13ce
z9dd57c1c6e03ac4504cd5ade7fb4bef9dc7f262af7a99ac37fa58794242f22a14238e07113a458
z734133ed6b721e3972072012f0448f3c00fb8eb90716d1444d57676a92fe3d93f180f95a37aa59
z705a5bdf62047c1ba9d2b540efc2f28fb44025a138aa2ab182f90b0e33bfcd98534acc0719483e
z5b76b44030800552a5355b7069bbbf05bf3a87362d644349a8665d0da6a15fb8f0a29f28edea95
ze7f96f84bfb4aa3a4ff031e072ec47eab6f233a768a36e61ead71a8de00387a6ad01230ba0ad28
z24d58f93b8e86f5b763d1886b36052aa33ef7be243868a753d804126a3faa111cd4ed6c1d42eae
z096b659134fc56cc9822cea7cce477442ec41bc63e43baa216fc2538864bc6ed362e0a4d874bca
z0dae38d8157e597b23407c9626c2a85db070681be4e4a4c3e55df5411b036d0402eec1c0e94881
z356c0231cca02faee5c12990d077a23ef9323f3d20812b737a9fc0069ba91c17b2f7932f496ffe
z155fc5f571b772f3cff4d312aaf19140e5df025f68955f5e256f9c1c8b0fac5351953df5743dd6
z636ed9aa3832184d1f85433973c88e41f029b849f480c6820456c8de06261b93e6a15b229095fa
z3d33ecd4d3be26412d06cbf2e71223aece4d0011269ce0f2be1147c29f071db5641c0875fa1a8d
z8391c7aef0fa15cbf4d4853df0c185edd8e7f4b3a3e21e3241b1b2ac524cb03285a19a0ed499fc
z3d4e003eaa74199b661dc3f713e111554e9979ed2d0250281179568a7aebf11c44c5e15b939c12
z03795c7e30c056cae260279ea515b7ce2ac1c461cbeb00adb8aef9c7aababee5f3c446fea5c4c0
z484c308b9821f5f4ead1a847a8f8d9adf4bb5bcff25f6d6004f6c4fc95f761f295815af13c3365
z632554cf39f6eff78a3e6e6055b449bbfbbf719f07fef07f7d6dcc8a0efe50edf51b10103b82fd
z207365ad026a46cec650e4d9e46b457e48186d99a86cb67b6ae5e0eed2e97733110cf1342e623c
ze344457a01307058b699d13d26837a155f0906e353933efa87131247e495ef160b7099c9111ade
z5e2a178bd5e08882afc12488d28bcec2f1e4a5472c6ae8332594b1566edb6181deb62331433af2
zedf9db653ac78fe6dc91371033359c86fd76b13a3c0dec96a8c1362aebd4f67d81b42a6019283b
z921da12aa664c19c72a01578264b1523579f1a69744de4a29563dd4d831b7d668636d31a36722e
z93f2a7c9e937b3e4ef5c41e67fb88f4a28bb963d8f7c28ad6c36d6e260409117919db7e63f02ce
z1f5dd46041b62721812b3bf03f8fb66f2788ab608cf28b617275c9f89ed08bbcc53a1650deebba
zf94accccd32aaf61b8bd5fe4db5f29203ac66808f52ec5961908a50b13312a193d3b86560931c9
zd87a0f19f84047372c1555927f0e40097e0f86b145a288c10643c0f8b355f2bc328353f57cd88b
z340a66579fea9b4ea97c6d3d19ac1fb0af8b05cb38add963f8612256ce93d9bbc745668fa332b4
zc5e634d211553686ab9b2333da0920116740c10729ea7193742241934130e91f742df674c33ffe
zcba5eda231b47d7c2fd8919fefdd0b45fbbe3569f46acb6c9c028b0c21eb43ea212292e3cb4e43
zdc0daef8aba01b7a328732221bb24920ec96255283386eb7bfb2234ede4956c3d4d30c9a4d3792
zecfc195d0371463c9792f1ce4b3a538a16d279a77295eb6dfc58ec1cfea2062a210d2eec43fe72
z4c730c5c69352c46ed0588ea3594eb62b3afae04f69bf57e8bb84c4dc4a3f505c705ef19893f4e
zb8f16e57efc4576700bbedb2113bd13ed3f4336d790cd1fd20064d96e14c65310fb484eb52208b
zebfba90decef3e94d68c34dea2c3bccb32f22879372d2ff1302dc2d432ac37190153f6f8b4095a
zf2fecbdd85060d6a7b6aa8ed3c5d73f890dbc7fd1f553e28a7bf9ce7ced4aa8c8bc0f17d001103
z8ddf078138f5dae7a11c242c19a21f6e1bfeed41ff1ec03df6fab46614a1f77240a33b3257e7cf
zc15ce5b064a2cde77c9cba1179c540b5fbfcfc25f78a443dd3ab38663158f96224698e6b19e8fb
zf0733cc7acda37d3f0417be30d57a17c313aadeb0de15339ace1c419532af7dd96457c085947ac
z50bede2c1489f114e9c3533c4d753625aaacadb5662ef1f616eadd228116322c1346186dec8c83
ze75acab8dcab9c077382c3c4b1e513eca0a63880788ed9b55baaf3fdd5afd9e5586a5fddc47aac
z3d5b0565f98aa2810f9cbec32889847a36f32c14494fb8a5fa08280b9b9a6b5184c22fcc350401
z9274615511f1a01378dd40f4bb7d424565274521f906d777de8b21b2a247f8642b16a958169083
z080258bcea060afc2daf075fb20ea5340d39005da845863f480c4200ab96a6f079ad0560151b14
za26dd3d85dd0124fe7973aa92a4e087f91a47e60b8c3ababacc6e3f642adc98063bf1a694e3f7b
z0dff2c2a8f4de4393e7bd7300296dcf01b2236e5b70c101df0952cd568d03e5f155b11ac224560
ze73fa579d3b3389cc5dac25a3c99033dfa99d8dca24b4255b0f970004adeaa6000f90f5ca6d31b
z69cd95814f210924cf0b13de682fe5ad5801d4b6077442de9e8486fdff4f7ffb39ea1b392c2356
z54d30b2b068b49bf596e00a65f90f29871b5773df0198f513db6802cb5c78e0bda80c5947d37d3
zf47f5392a41bb927d3404e09f818cc208e3deba6e5990a0a4757238129c8e44581136affd66ff4
z3afefd4661bf2303fd4c0e4492eeb3c4d4e068219d90a883201e45ba9206ddde2501cded9e82f5
zfbac316e87d4835774e8b051b5de96fdb0b8acf09c010bad91b69ce2e81a350a63c7209d4c1aae
zdfce1295a28d0e7e1110cf5cb1c9dcf0a6a87807eee67fd2ae0c7a352d0c5605f8c111f3ff39b8
z63c7a237a75d2c098feadc235da5b00bc88e0091643527cfb3ce5f12057b0d51f498b64e4e3e98
z4a980d96ea47dbe051f7eaedb1962ac6ac7b8e2f36cc697580c1664a65d27ce63f842731933e7e
zd97212ad1b91e34271f5db3e21a0c2b33084f326d5ae0ea05404f2bfa62743936cf17d8ab22ce9
z7806af546970b79e412b4e5996a00e2966df9bc90673b6d4e0d4607068b3a2b37a5c26fcb2ef46
z4f19d3796cefba5317c6889d6864f231ec3d7caf9f3ca62297c8a794bec3914a8ee9911624dc84
z803a2ce585c722010e93f93668d7f6a0f14764b28d0ea709a3a02f9a8e75c8ca11261f930576fd
z026cad1f871a6985613e4be7d6705f0cb468e2b5d980f0b98179b368553e0c752438521e681345
zab30084da59afb6ad8da06c70fd19adfa488911fd041b0301a6617c80bc3a8163600d35a5dc089
z3075d3493881e9aa015e4d167ba8bbec6a61b18ea7b5ee99161aaa0086fd2ad239907966e753e4
zcd2fa90ced983fa766356660718049612a82825b474f6e8d5f78f5f88523a01a44646bc241819c
ze2d874223cf7fb72b60e6d8592b67482cbaffe90cc0db7c7ab699ac3ccb1f9d53611c9113895eb
zfd593d022c76d1e2a1d46dbbbb430eaa7e27ef62556b917328705bab1742a8d5b7d25547d22ff9
z86cf7a0e5c3dd8339c959f8f51a1d724e251ffd68c12264abf08fcc1c522fc0951d39e5cc6e2e9
zd066b8da97821566e69d52ee28ed1f18ccca3ebf0962b5ef4d41b15c76e4cfd77764f33bf2c499
za2b4d83cb08d127fd71ff8c21d71eb41ce05ba48f33f8143a8925cbb7dacdecc17ea594a7d166c
zc9e3acabb61083f0791bff43e999b8429309836e7ec1dd2938430fcd5a4cbc96cda1dc309c2f67
za1bf85d2ce60e08938bf25a150fe375d457f97c82cd89fc2c84e00cfca6436dcde30598f07dd35
z20efa3e14389fc959c11237b892d033af44bf5bc49f60391020b7446e89116f1951affd912fc8b
z32609a4487b41a71eea98e9888d83cda6656eb941c85511ad5a8de1dcb6e8fc07b82d1fd946156
z296e0460a180ad82eced4b9d0156da9ad86b08cb083377865e865d841efcde741b47f8a4530d32
z6e5995cac42a38169b3393e987f2e25d84e9a36e1f14a8ecef54f56fba1eff7a7b012c04747836
zc306c863637cd934dca3d87144d463b3d525eb2faadbff51c0206e4df56585bf0a73328e33308f
zef9c545036477441c957a48113c63182bde7f656865a144fd1489feca9cb123e2843858e0ee896
zfcb79e40f3aec0aae19f51d4b4d73d42ea3c4a386a388ce173bd52ca5963798bcca013724174ed
ze1e8bfcc4198b8d61a6268a56acb46927cba7deeed37ba08d656c833468d21888ec29229950e0b
z9b8d44e9edaec11d9cd5ca05bda17f75f114f54e624cf6f7c2dc92578342125613538136042bcc
z1259bafc39c80181ada1e78a41b2a5799c7ccd9b381c15a4560801fcccbceee83e9e6f3b706cbb
z7a6bb022991631db11081c8a7e42c2facb092fd983e2018496cf7058bd4285d0018464a8e9e531
za685cf1deb5e7bd7eac0cff6daf8b732f9782cf6cd8545959fd5eaac1a0df047c4ce129ef0e1f5
za5db3083ea1d3e8e25af5cb8225fc92922d3eeb7d1f3ef8f14ef46c62b41d20f7cdf628a794ac4
z5c507aad39979a253ec55715c60f377064f2f781a58898de6951340e392065034398a896d7f6ec
z7d265665a83f8d9ed3a5c4ce934b0d1bb772e45d8b0bfd1ec72b92bdf3b8853ba7ac3fc801b8f1
zb15fd6295cfe0df6a1d5ee4ed3805986d63a8c8261f013df503c14456099d8eab90ecd47304722
zcfef6e3c0a15773c5e3636a3704977cb43071ba3b4b7d3361b58cac60d556e40bec931e34b0b1d
z724dc9e9446df5dfff1b7627417d4233d84e6692fc310913db87cfb04346ed7846284bc5a96d9d
z0f9b7d1243556192e72c8eeedeb4ca98844a43014c53c660b996e3899f0062c2e8e95bd55bf360
ze28ec78f10c6757a5ac0994aeeb337f11770e740c0b6656c1b2b57b24c03cd7ddca981b6d7efa4
zfff25d612a2385f4c92b2e6fc8aad4df35698a7a5e83359523d1a289fc41d820c3bda11c1f0a5d
zc6ecaa06a2f6a4e766ebcaca6cd1d2732d2f41a197fb7096da2bad30977bf976a1fcd8be4e2963
zf566f57c243e5f1b438f066af377cd6af2063f873a3b02594bda8ad7f834650048b97cca471140
zf5b9b962194936223d56f7236b088f2c986e6ea23f919e670d5b606e2579c17056a831b888b322
z5cfb5a7609af2fd0afe81427a556f1dfd918b8bc6ce5d52716b881e05b3455e185b8a628bb6fe9
z56cd75a9981d2c172fb213984624c836d45aca6cc0d650d1e6062868f82d7798616cab771ed0aa
zc368d2036e22216f033a0b6964e2bad7dc8043846835fe88ea596cb67d4070b682ed5d871b0b6c
z6bba05fd92f717fc3efccd75b741243ffcf11ed339edf357c93c9b2151b9a1aecf47ccda909269
z39cd71cd1834d62baf420ae99d929229d5401ab0e9b9500ad7f833845b6b3a4ef5d7ac9fc360a6
zfcfadb31b1c41dc836b81f51e9dcde66b9718572c581b0438212a54e639a1532013eb364e5d912
zafd6012a54332a1a36a5950e403c870418fefce812d1542b8f98a3f8debe4470f783efd0b0694a
z1799b1100f858ba01fa9fd6187c0a757846b146974d5d3752238742671570db4f7c6af0b2fc70f
zb576c1746cc5ccb0e1644645d06d893f38adbea6974f9802b436821afb9f4f7e33aa328ea51b24
zb16a5c681e96e6192c6566a66c07439dc43865e2e2f7974da1f6abad9516a1d699ccd5ba0cb3a6
z7decd1b0290755dcc3500ebb056faf3be475ff5827c3dc2b20e333bb7bdd616a0bf9ef9bce4d83
z2f9256241bc578fd02fef5d093352980c16df515e821d7c027e45de0748f888d4a3320d58a8810
z7932f4bc120d689e031a2c73884443787e7aac37db045912a1d9f0fdd8d1cd3ba8f1b17f579459
zd6464569b7476043994449f26a027e8e7b3400de155ffcb32f28b12d42e61bec218bfef54e5aa7
z8f0eb60bdccecbbe03c08b2511ebd6cf04de579e996f106b6d8ce86e1ee160333e2249bf86e6f1
zca0ca2871a793e41c372564d667c37cce19d01590f4493c3ad3d2d86775a551feae40955ff57f4
z8293896ee6abac15019ef5b854a03816d67e9c084425905945d1e55a228a76b93d7c8ab92b94e6
zc7b26c3bbc683aa2bc45bd22c7737540bfe5eb879493e5cd6ccfd895d0a8e1c61bc0fc6907cd1a
za94e8071862eb38efef2cab9e7c66c2a7bef40e3e0b73096ca2b8c0471e12fa6cdd8b1d598faf7
z8c209c055dba49787c01a4525290325c6d122cfdc675498ba3cae662fee31817c629e04af16d70
zf5efef5024ae497e29848707d908725113fc9f8915d473dc78b3d50c94e4227dfc3f90842073aa
zaaef641c688a08525779058a96d866c485ff3f10a7c4658336a6e221306292a14b45dd06ffa49e
zc62a19084eec7c6ebb048c9d885feb9e345f4c5ecf71303e738ace916cca51d85377494271eef2
zb330a75fd09f01c44a837e35a27de98153ecba2a169dab6ba4a3cb973d6a087087a03811877cc2
z6da818b1bdb9c1e2d672701c59357dbc738db5fe14a2db323fd5e654b6b745d57bd921365ab100
zca2bbead9b71b949cfae716ce81899d4e4209827b8010b4645ce874c90219f580551517ea138c9
z87320073c4dc8fa3ad66f306bf91a3be4813e0f1cecf0221ac50334b71390623fe2d152166e72e
z5188b605d08f1d7ed8cb01cd1134e459a2d551a63d195b620e8cee16b2926d16c6cdf8eed4c7df
z9e359275a62be8c5036c89459b7c4963a04daf705d097050871e33dfa8a818a1e9568d53c9455f
z509d403f51513d5893ac662b582ad619a370bfb37765c1d3a3d276df58c65f0d3caa666c4a7c39
z5528fc2c8efbbe857b485b02bfe49e0919e1897fcca38248b5534c66ca7f760516ac4d3e09d18e
z4aca228c6b1ad0fad47429978f6d66fb771367588479da45282cd60755bb80b447872f8305b60f
z5e95c5f2285bafe7a0f2140743253d4bff96c555c68120f320235f2e5e986006893ccd9f08040a
z8b5c535f420436b849096a835532da50f86ed939f012d7fce146040372714abfae5b785dcfbe7a
z3b25c808ae1a7b8807cfb296d972505a8e9fd08d905d16b43c1b5cbf49e4980ae235cf808b92c5
z31babd58a69cb6cd501f9b37bfb48cf0ccacea1507083930bc7c360ad381004622f7fb5f7e0842
z4335b9686a6f93af7def9e609674ec51a3e5c3e5be2569e1f2e355b7c4916acdd5a41b67c7010b
zc8ab7317a6183d61c4ab338db64438e30210682761b344f42cebb488541e5d7fd6d698e61bf4e1
z136ac968384137ea5e92eed541e9936f57dc9aaba5431dd8a965b7178cb2c92d139c55c9a2793f
z8bf11b1716a61a9248ada02a26755f817b477e920ccacb83cabbdf5be3ef94341d40449da49897
z9a8c2873c891d6c212a0825fe6a3097d0cee8c21d4893b3776ebd9069b30e11109a34982b869e4
z635ed7b9934a8c9e07f225f1ded6ba0fd43c06ceeeadf6d14f0208cf13f72d48d277a7824efb2c
zfb4e5963308de8c05fb193345d9e481b3c2b4ab51f8a2442e3e96ca6033851c7a22f3bbebd9bbf
z137ccdf28c71a0bb2398ef61c94625e3e310dbd142748959cbdd9671537142fa4598b0034a9e11
z98e132665e3b6254260e8d8aef874c6fa3227bc9dd8d911d278a247778ecac757ac7487315b5cd
z52c71e10e26fe2db2361716ec30a7581bb0a1243c47174a17deb68218c785a1dba709410c22988
zf5fab024bef8a1d78d875374895929654638afbbf5ff2a5148c4ba0d69f4025e06352db037b0c8
z326528d57c405cde39e05c750a43cd5c4bc82ab1945b4ba49a72759591e04e291d2f7a7bcb5544
z6c4da7ab92af06ded22cc067b5466a04dce58326bb7a50a3318813a40fbcc9d2e9e6e7f895fd73
zf1e547a740237c09791f64daa7228484dc4e44abad111870d902cb3944b5662db995a92671d437
z92be31b50979d54c3bf845adb4c699aac971318ce6372ddfcba5a01af43f651ceb801767238b7c
z6cb1fdcab11591af48de1544d045b01038964ea2cc9b29a323055ba63356c076e5630e551fb07e
zee7cc62c31cf3f91d4c79de30dee0972019c1620c781cd33a9ec95203cf238c8d55a82464afabe
z7752ec9e846d8811217f428402485ff2891234d34e7056090e7616446d0e4929daf89f9d75e67c
zfbd1a4f25253ca2ed6c67ecadb1437688afbfd36f3a8c810bdd2e3856e9ae719a1321ac456fa45
z37642029f1a2ef24f3cd58f13893448838ed4b50a635f577f12ea641944d874eb424d4842371fd
za0fe0ae7291c6ac213456515d3647bdc833713f4352d272a001bd4c57c9899d54bb8e6b4190953
z34fad9d134cfb3e7f393506428af16db0e21cc30fab3abe7052c03e5103d8116d2bfcf42713e20
zab4bfaf1168ffe2d57783b0b137bf1f3e09287ab852584ddf29110002768ed349994d14749506b
zda703d7ad29a6ec56b8356900de77469c893e7050690b18b06d8e631ad667fdfa0715b8eedc84e
zb4b3d443db1164b44fe7e54438b206e77723f38797d34d1f78a4a27eb5ee4dc8f22d626d540300
z3b62c5b915c44ff63556ab9ba56d6b96f5f521073923c39ff3a6296a5fc662df4ffbe0f04d717d
z52640b0b306ea0266cc4794760a5461eea4e0639d186af540343828607660c01f234b5398e2cc6
zeb12b6f2343a287df6ab85514cf5e7a8931ebaaad3daac25dab90ae7bda35e6f8114127a1fa128
zd5a984dbf91c594c71383a849755709f2f731f69ffcb406cfd004a63313c2534dec74ee81e2bcd
zd47bb195fe35bbbc11c2c0a3341bf99c3f0b61f8dc9c9927de451617b55098edcfb30a0dab0c20
zf676240c8bfdeaba63a00482bcb248fd556c8b9af223960be5e0befdc6053ac6fd3fefce3882de
z145b8235773f1de3fca08e7d8f5b00f0f15593ccbaa7daa4474eb6544873a7bf9def2443319aa2
z6595855be5d1288d9c0acba476113924cc7b5c19ac4a37a0f28ea4fc15851d9825e34e67d90aa9
zf2cfe08d2be8ea0b4c55d5a4e69170063cd6216be67439cfcf53e42ebe40b984357802a1567183
zb2950a218318dbbeb135fd2702e2de11e797c50e2c41073d86e98cab86ee65128a3249c44abd59
z34b859fe3b92a8f2d92a55e0a1aacc086ec38ddbc8d3bb7e22c9b593674e71f7d27e78e765f4af
z815cd0ea9d3c21d784ea11ad98173f2eb14b02797eafc5150597cb4744d6503af016c3b5af8221
zd1397490af45fb8b2ae16dcddcf852a24665ebbe03f1b0d70a5f19e754f5c117caf6c7c4b14b7d
z73e2e47a105416f90e549fb057ee54c59d1c2f0c18b9b13cb77c2c3cad81c195b742c122eecac1
z11fe0d22f5cc1afa9e82d259af6e1f7234205e040ce0551ed87611d8f05f1523cf9871350b3487
zbe75a6752b714c1f8239f806172e76c9acddeb5e5ced85a3dff10debf4146f37d24f001f993e34
z1f0226b400da84bbe4d59a91d738dc8326fbe6490260bbe070a0e7fbc6b48cec023740d63c2a6c
z301bc1c3406e394dbd159246b3bfb1fa19e5c72f4c7f1f4f3df1296fd5d9f0bb03e391a6a56d8c
z48531565daf19363bd19814fdc4a20b1ef843daa9d78801cdc981d7cee53c3a86bcab18e25b15e
z388d240a416a3834aae7b9d9e8ba733d929d506f87865ff6c4013ce6fcea10487a6e36e9c28cbe
z55ba5063736e228733188ce839fb24e2a004f0cb89ba39923b555847d1e6c0082e52c583f8de81
z9979989d3db3b1a304b36949b9ae9a587a919d2d5fd5b963420355bbb09d2d2806f8daf2c4515f
z5b4c98239aec5666b4130e277a33f95f3c1ea1a88882593190324e993ed45a6e8583a2d3d620f4
z713831c2196033c29906578a4b0578f425e40b13f7d1c6ea57d8534c77c86d454c2e8dcf9e60c9
z2f1802e8d612fc6f2ded1377aac7af51cbc3a351d9cb93a95ee48453bd3bd4135169ff58315454
z1d3158e2094a7ce95a7093ae09f3ebdae43149d5ae02ddb04311fedb212bfe9618665175a3e2c6
z94f5083e8815ba5c0802f884b7a28c5dff3e2576ec1978d18e8aaa563f9186a029c3c6d73aed5d
zdc47acd17e66ddbd9ac5eda9c405fd19cd33a80d8c84b4fce2eaaae11c88a91d941a45b93555fc
z480ab6fd2619b2d058652ef42860be890a1247acecc4e31461dc9d0cb667afab1d2edb263fa12b
zd98b4fd20c4509590bcf4e5a9936cb6ba18165efc40ddd40a7a73f249621a54795fb68779dee46
zd80ae4f9b19a276f9d811e7769fb325be04b1902e0f8de09a8d2d15a272f53070675bc361e4223
z0c24ef16ae80e3c9af86fd034f0430a79167be6831306a7f123b2d240ca817af6f61c7a8f43618
z8dbaace52f1bcdea69a4247fc57b9a02b9c405e242dc3865f96a53c4b0866629727e5c0d00ea93
z43eacdd483399a2fc767df2e3a37bffe04d5343ce32e26605cca86320251196190817f1f077a5b
z46aa0293880d797e38e1ff51783c79df75ffbde2ad944678e30f2e52aa93c83a6524dc5bd57881
za72a382dbf7e264565ce27e7b811104a49bf16bf4dd62820d44bfc2886a6ce4ccb85d8df64bbb8
z985ae13bccbad50a62f829df44041176ff10ac5d593ae1460120bd6e597dc351df8782f2cdf600
z2b1407d493352554149bc9342f40df340e1bf07ac8536865b7dfc9accb859875d6841f7c019d06
z38d5b2e1c1fcba93003d0347770e16465f198a6dbdab48d5ffa53cd144f28c5941e5f50b68bfed
z06864de2545e7f07b93e30b58c21690a1498163dd7de51819551b32ea812646b7e18efef9a43df
z74bed1571f0229eda115c0464996f2fdaa582bb8ae74a705250bc0c50bbd5a5f585780321c188e
z3509967fb9829ae74143a81c170b43b179c3606b4c7535e242a67922998a7b845d8a8de521bf06
zf20f2b158738dbd92699622bb57075fb9435c60c2f7b7232c917846ee19877e2f38f30b945c457
z5290719ba082d46bb0885731c633efe70ca073d353761ca07f1958ae7e158b23034ab990516179
z0668c1cbb6a93fbff0e6e916062cfad92bc6f724a17539904a7cc16d4afd0f92a259be7f32d047
z9666bd11185acbb03d8d0652403dc3825ef1d5be04a074ea674e9b770b2525c64b8d2fbe572396
ze2094b0339f5fa7315c00f9e2c0e4033cf6aaea2464e5089afb9753c46b35b6200c24a4681301a
z5797a1cfad051022e656f14c7e4362e27be848f59393dbbf138ba4ddb8236c8814f39a43fd72ba
z140bdceb7c80210e221d68d148bb7268d883c1105cf0323d7db3ecdf7ff6f42290c232ea8640ac
zaca7f9c0ba91df7c34d5cc5b8ae6a1d0cc70db89fcf61c794a0c3b0138ac96b34d8e2669d2001e
z841e18609bb8bbfbd20564441ea16c9e7d503be44a29428a178ddbaa724b23e825e85919bc4aa1
zdfc956e016c7f2ce224335e602d11985e2bdd9027b8f6271decf35bb31b603cbbf7d4ad2aa9c4a
z299be90d5c50f2db99fdd461ca5bfdd03ac9a67b27241858dcd2088cd683bc8950df0c8a6511a6
z7aab86f1b13cd9cac02673a50fc7b84b3ce14cee8c7eaff1f9565cedf265bdfb8cff1f30c90f41
zbf075045ae9aeee003148d835d4c968e7d6c957e2c5da9a1b753fe574195448da7a140e67b32dd
z0b053ee3305914a1aa25dc2185385be38cc25ee0fcb5116129b801987d40fec28e0503d11f3b9e
zb4a31c853e0a09b1423fbae8b622a666b49d566ae2f00d9e4082ec0c7865a08985995060ca1073
zb2c2b3e18cf26593797fa7947e5332bdcb09007ba7bde6c31be2dcb41eceb78afc17e4c33ede54
z6213059c05ae5c2ce10d0af9ba36afc077266cf834638a11065805c8beedaec9577cc4b0bd7c47
ze40df9505f96b54d651d3f92d5714620824fced8e3c99dd539829d3ab7b708f37c84157ca50f5b
z6870f3a9451432e33df5c9264457b8bad4881a40b40c46b8cfa3d380cd9ccd4c6856b4bff9df81
zc3643c098ff07ec9e375634fd21148f5559d75641d64a2be7db5e9ed4f039ec608d9b1d4216988
z10e15bd0dc15268235c3029b689b541726f124c3b07a4664dce1267fd4e2acdb7ed7053d77d577
z01d61bb38b61e0778a2181cd0a0d9abfa899646857bb574ea0b9d295f9c5e487148b91063c277a
z8fba6289f5e5f27c2dc2cb90772c7a04ef32c0e89631d23e5766c209198dcd7ae981bff43cc914
z4f7a41366804edcece5e8ede1a09c39503696b7fa5cbbf34bc4cbb06b65a72336ea0e34df181d3
z328bb6697c53e61ffabf0c40d5419fbf25fdcdc1cdaab4f9092bc41f8728031efca9f6852601ed
z0550c972eadc4c7b515fd6c6c53b0b8ca32ac2ea22d2c23c3779031e148e5198ef20b1562bc4af
z7ffc66012a64d2b158073608b9d7f3d9c717ab99be14c442bc9009c168a7d181d2bbe95c409d36
zca87bc1f77a319d7a43318d95ef7365638cc305179bdadf05b5eb363da3d99168572188b111a10
z1d7578a89f949ef24d9e6fd0d55f1f7989ae88e327ad788f9b31340726adf1db8ad2c550873ee5
zcc79c3d9e724436cc17ae4741b18274ae0755849170173d0a5788fdf7a5dc96ae8ca5310848096
z2e0c047dd4814396ed98dc350329cdcefd3c13ed03d33e951c0ceb7c412c72a726496378f5a2fb
z9a41b98e999cb238f6d30f8999839cb3ea1e817a18e18a89e85d127b17cc6d189e4fc75493d36f
z1b639080d82cb98f8765e2d0e4ef01fd10eab337df5c7487745ec19281d57bc277944141ed0197
z480dd2173b78e0f23bc662908ac314677f39c80f0d60f6bf1f62ed458f73bcae0bc9cfeb73f80b
z43032b874aa8068a4a1f8ea734857081ecd54012d6be0808f2fdd0803b2bb21a1fd1fc93a6d12b
z239eb5c5ef35867ba50389dff35a8a5765450ced5b21aee8978300ff129e5e902375189bc68e0f
zbe0662666c3b12a4fcfc3b36563fd69b63e9a042369a3e4ad05f6c64bae833773a6b9152880c9e
z59f929cb580b6416f2e080dd6bdaaa56cdc659c088a2359694cd389875bfb67afc71523ec7c30c
z3611d7f79b8917d0c13a7d11999c320ba51507267f782bc7b079d7dda964d5779ce71c3bd555c4
z21b0a450f6300dac45825bb13609eeee83a631f069aa6571edd915c0b981c88cd07ee917555800
z6db62b1d0046782e512543feb96cf7a754040caf1e111d500b04e2cef9f91c2e06001967b57da1
zeb59998d45a7c58b00e0e265d5080f9b96cf8d5a6073680a55d4208e304cab57c9cd94ec3ad91a
ze4a3cfb13d54f35a370b93fb3670c5d6016dc931add565d800519490bb23bbe1bce7945d745744
zfa3ccdfdd7cb16d523df911f5b9cc2e970098fc8a22ca829f0a9757078c1d76e2c1304effe1f2f
z7dca48bc375398c96cf0be14bc648c5d145a22c8dcfb317e62fa1308dbbf36550ef730ce788f4b
z5525c968440828bd180f7e876a459ecd71919e36e2644c3120c7b63c90d70cdacb24767868b80a
zf49bfa1c8fc235f309ad5c22f01da7936f2d9f8ec62076e6a130d5e72db671da8784dd51b776c8
z8659f061f5d6ce0644c635947f5ff7b19e1f5bde8f56520d0a65619540032f743920746e939640
z845089659210c8a532b118be6b986a9afc6269531cfcf4727c485860e2229b3071097642ec1886
z041c3c1f94f30baef7a5e1cf0eec52620d2e0ec4a30407af938dc819bb1257c2b00979ee7efb04
zb5024fa3c3fa010aec5b97248e6be1c5e84ce3fe3ee7a34ce29b84098a4e3f79373005d7d896d4
zbf428894be6420c1f659e2979d0730179eb7c560dd9875f3c68bfd6d1f7987652555d1a4d6a4bf
z30f3f25de8ae6c71ddea1d2a90ec0459484a82eecb8ff2bfbb9ac657fb925fd68d6819d4d660ab
z4865dcb42da60e4304edd3583aeefff6e97bce306eb1dee8b44a79b8c6ba180d42a3c12ebeca1a
zd9af6e9cb4289dda0a117998d210837bfb02a92e7f6448708e7ff0e79b12e9a0464d95da708db4
zc20cd594918e76a8933e0ac035414ec39fc7f7151192d8813d5e007f45e86f283700104b2c7313
zd8e457192d301b32797618bdbcd51e44eeefba3965556f97f84c82be3699fc0fa6a39c0ec567d0
zf5c5954e5ce64420bc775b713b37f0ce47e9fd377468a831d37dc914c293a0f873e6b1b5d73934
zda8f0225572298510323b433bcf8093c57ed0b44f9541ef769915cdfd14e7dc0185bb30e57d87c
ze0a936ec00f0d48f1ae13b0173d163e204511e29387f1d18144b1c7e6fc04dbc2acd07dc85de44
z6f18d7c77311b6fc2c5dd41bb454039b74197fc8edd2dba997d3b223ff8402bef9322a3680d725
zb37f846584899e8efc6c1b59a7124a849762f7614db63c40f577e1625274c100057d12f9eca509
zfa0d875aa0ce48061dfffebf5ae799989c73d5a7bc639f50d924f9536dc68b57364948ae3a6893
z673acfd59b7092f49450c517359fa37555dc0f03a7236697a988abb9eed89fffd079b9273723e0
z2176eff028a7722b250b96628b015c225c34b92697e5ac57e9ef4cef595dcc1cee4d12633ea145
z36a543bf8f59a5bc89564b1faceef46d4ec71e19f4b5bdf033aee4d8c8e2c47f0ce183595ae8da
z02f4f3f6ebef4f693dd2dc5833dc96a4fff721d5f208bb6a705d7d44e6f3217657b97ad5acee71
z44e545311aee87fb922d61b37b1844948cb17616fc65db80ff159b8d941752abe0f8037c11bccb
z290e7eadac6a49fe62d24e22b21cec00cde2570a39b9f6ed92fe6b7e340fee7468a0e6dd541a17
zb7b5fb36a1f1c469222f26cdfa6bf7be60858c0a14797128a4798c5e5ae4a97f07d1b2d2b34552
zb43eea68f4ca308a814f6f23c31f3388cecc5601be7147ff58a64e56b3e7af35675152031b7e39
z975d6ed4ede5b7d6fa096f35b086e1f457869a60ec62ce3df4c12272fa2d359ed07256a176321c
z9a63234bf8c6236ec9d9ed1eeb4b922764d6e35fd2ea78f8c80b0bc76cb955bffc3b6b7b09a7dc
z8a63036a8e6dfe2f65da6d798f0776114f51884775a01776279974853cafa5e5dca0442d20c9d0
z9e352e984ca5e2c50c1f16f9a2c4d02e6b1ad134d36d61897e6a9e41e6abe7686556588dd033df
zd841227bd80713ffb17db91dfc5023ee4d6e1f7a7cefde7d530a2e393b954d21c8f145c1dfd595
z39fe6ae96338a22cfb09943dd2279937c9fa04ff3520d20f31eef647aea0bc26be3f165b7a5e8c
zd8e165919e2302456942c7a56981c5084d0d257e5da78f165656a1a7b67c891e9edcfe6b1bcccb
zeca0b26f09bea1f46c9cfac968a5fb7a138406272abb512b5d259890ac221919067f3e39279053
zc79bfab7eb9ccc69ad6400ae864f0550d0bdfe65b98647704ddd5b867a0a4b16cfef1bd652f915
za7e8a68c2a415505b0ffcff62a42eb74a7f400ceded69e89be966290890965b093d0fc05e7a746
zbc69f389e9eb91489802cfac3e92aec7a5fc1faeecb15dd1205795827c0fa3f7537985d398695e
ze6a721d73c269238574dd11e21f81dd321e5e7f94ce8cf436c92566b54c70ba6ca2e46a1ac4786
zde3ebc712e35fd3aa534c85d7708666045c7f8e0ba112a94a0ede54ea019275b605aab49203b85
zf8aa1e802c2145615d59cf4657f74567946a25a328942ce43bd3284219088ea13087ef00026639
z5dfcbe36c3a02bf8da14a8e8d1965d3dde7871e8e05b0aa5ad61e37cddd15769d5de71307d6b41
z7ff365f4fab1509f876f763b836e79537e7563419bd944f875512e56dc26cc5e03df43145790ab
zda780139833d091dbac7ccb2cd4983e427818d8f6801aeebd2917fc4f51a1e566b254b3d50d121
z987d2c5c119378e8c30430fb5a30fbc4d2ab04fc21456aff9e04a2cb12770e3be7b8b5d51e07a0
z49236490347c853fe75d7ae730e310794b4ecc74a0994fc47b398b484ab5bdd009fc4cf8d255da
zbae16cbb305f7f0e6c5942d1935144b21ecc270a77bd5218864f796b5dbf34d73168c4b7546df1
zd32b15c624897b80f8883744b88c4156a551b270fa00d93086e92cda722f37bbbccc9737219bc3
z54fc2f9579fe350a1d54425a4fe6a4dfd297645c2453c3b7ff51f954e315a37c7f81ae4785e775
za57c278d77c52a3c58de73efb81e062779bbc685250c69c613da192f812c26a48d69ceb98c9959
z2171bf262eef755e97e151208cc13f707bf03afb1231ea601757389ad42617543b70b0fedc7ef6
z6217642c90d338cd2c5eadfb355055c77c22fc8f7f099fdbe4a3a741ec79725116bd112595a95a
zec11c57910d9c92a35550a7f88f25a7ce6fd7a0b1c92aaf6734187be8959fcdb1ebd7c4f0365eb
z1f7b3ef6739b505a0176be7e5b050f338e477568a9cb38fd949d5cf9aabe61e2f5bf6032f43fbd
z66804bdb761302d06cd967a45ab2080c1e74bc687031ab146427af524bd78eee4f474462b67a4a
z0821e58da81a58c3df1e99d03e9e06ab7d4559bf67c33899e3db95b7843705ec3dbed4f701d35b
z470632eb611666f0f9cd9c9a1c3e9a30da23b796ad0ececa48851d2b24decff2af9fca5ae456b2
z4477e872e8ee2dbc86139ca4ebb10c38d4d55280a4b35f7aea271594e8dbbdc5ad4c01bc2db306
z41804b0c464990823bc58b2bc5fb7de82b1dbf68aeaf82997257bfda9b7bf94ee48268b624bfe7
zfbb56043f7f27ca861d1b75ec35b5fc784bc2baa018479534eeadbf68a0474c7d9b93174f1624c
zb93bc72ffe267bc4e9a26207da887588138cf02b8e35462937581c618f275a63965a941797b44e
z1c4bbd14acb496c23e25c233578df6b50c28f4e2bb4d2e42fb7d7e0de6cea25adb9d250e919e46
z044dd6062ac22bb6c6412739e6b59c7dba4cad55f7152f6df52d50ebb39967146181ffdf5f9ded
zefe859322ccb1540603cdb4da851f4880186ec32b0771f03e3774bb9ad4730af6135ea469b0149
z631f0c6d454c96eb4f805069a9841e21d8f7fafe9636b369ae72ac2d46cbc4e9b2e7604040ebb8
zd6124ac741dcb55a004f19c2d561b8c3a0f0f6535d71c6992b35088ae4d9f19eb0a306985516de
z35fbd7e8d4404d91578d03b03ebe2807b2986d81dd8aea6bb49216d2787deec58edc52a41b92bc
z5dcd019847be15ce786d085a0fc6278c7e4f69a071e4e24bc0e13417e242c92e6e8556e6d25d10
z9331cad27c7e8238907f5f26c3b6bdff0fab9710fe0ef76b21718206ee4c0347a3cb41415a3531
ze8da23efaa739b2fda4185d869d10334f7e12295a3496c5736824379dab7253ca6993d9723cf47
z29079786b0af0228b60d91d28c93dd8fc1b334110b22f22ccf7c9e4cf68d0124fcb80aa2de645d
z7b2a8b73b7efc2c3c67dd9dddced0682bf3070c5c65c731a68195879926db6f63912b291c78f95
z9f1094f578cbdcd664a58632208022168986e15962a552db7f4eecc981d8315a6579fa678672c7
ze14621f32361749fe8c3d6826e651e55eef05fd1557751abf35e19f09d08242b86c1d6941f9926
z3f38e7dbf5f3d23b5bd854847230a58fc48e6c453d1a3e7958fad054dedc31ea42c514612dc727
zcf72157d0554378306d009cbc00d5edcb3c411c9f766e4b7c8ec65ceee477812350e7de5f1a753
zea2c53afaf55dc10f41ac92cfc5c7cb69210eac488d95619bb0fce6f51a639e8f501ca866cc410
zf79d65fb7eba2bed37ef80701f836ffddd3baf5992d6201432aa67e4d67a22ea07bb2194f1f816
zbdc3d8af56bf13d6d624c77a72c9b467ba30613700ccf28740fdd40e270c05e19524a2f7ad227e
zcf1a1ba3c2da782c04c7aeef99650ecff1980133974738d2ab2a9037990d6ec9451f6fb59f8d5c
z031402569f5c4531f826f6fb0b82a94e04c2d82b5c37cfc4adbee3d4702f4636329f84acfbeb61
zb94033fce74b88ff0d0b02f1a512eda5ce1522fa2b1d765491e2237e46ab63556e612c601313a6
zec695eb3e3a671e7d0d0372ecf34482a46a41543244dd0e826dc4c17a795862a26961bbc647d25
zbb8bd9767c2973101314f5da5cb7ddae991323c0c6712ab7e20f8581a02e5c758d945022a9e518
z4c8bf134f3dd9bfb61bb22d670ad7af9052eb40ba5b3f65dce25e99a6a96f472e06c32459c3ad0
zdb78650c65995d532b0d3e59800ac04a8129862ff0a533e8a2a94fc332342c84b738ca131916a4
z37435c7668077f6ca2508db22db36460682cc3e7175a74e4b04aff4177f3beda1e56acf34e2531
zfc442993e43f3948db4709fe7fc40dd55f0dfdb9c9b14fd4d28f6c6ac005b4936988ce2432d695
zb2bc88286cdab5b15fe286263ef932de8f0874a4666051b1244aedcaf16abe1f3778bfa0b874c2
z93a251ae63f9ec5e09e44e38e50fe363951a3efd928325a2e01e02864eaa0111b92dae3470d9be
z4d4567bb9d539b1ce2d81ec9268598ff4f5dac53c935a6c55f22ed140ab69afb3fe264db1959ef
z4aafbfd186dffd3405070b32f9d5857416195d8c0ba403bf57ed2eb05f29c7459c65e812727ba6
z3fc6e1bc0d96c9068948c4cc773863ab91c0e5afd739d7ae49d5e502ecbb6e61cbb8f856a6396a
zf98d187afd7bbf66cc04a63507c6aee395f86aa99e51661b524447b34ccb2a4b5bb739d6ad5ae0
zec2eb8c922ac0c834120cdaf571299c83a3de89334ad8833947745f0e5a6cc74b0a445610836d7
z0b1d953baf14b6572ca2036a840d46ee6df5da47e78064bfc99ce7d5c4c8ff1e22a00496c33f26
zcf57137b9c7025b4fa42489b1caf2d7567985ba9abbc1ee5831ab3d87ad8d3a70eacb897abe7c9
zdf176b1ca306995c394f3b2cba9b77fd00081c1531f9d31cc1488e229ebcda0993d0ed517741e2
z14aa28e926a5ef53b350a1291f0fd3ba0e4d21638e676f9df463262182ea2b87bed99d822987c1
z068e6c4e9bf4e158bc5813a9c0629902f68a631b98beba3ba19e7935d5ebe9071c012ffd94504c
z3b228e76bc3e7c48da20154ca718c68598504cdbedca0e1a6ba540123f1e3194dd9776d7531024
z20c0196d31aaff3975ca63689724517fe67a4a4dee2c07d827773aff9eeab28b1491de4f3c0caf
z2d07340a00495b5c673c8f8264b6e576e55ba24a732bd85826df3ce64d39a183fd5d5d98b6161a
z26a48913a783534294e501c932cdc12f778c3aa8fc6ed1396f411a2e47baa642a7439429dba026
z6f8645948847c66bc454ca8eb816fa5f08c0d40914893ba027d71ea7f0b2f5aa4deb38d730297f
z744958fe0641a224129e1100003b030023ad5384a9435f90a3ab43b84882b64832ea76a0a47299
z161710f8c135cd83230f65b320bb979afaf41dd37cc7ccd100df8ad559e3dae9019f9661fe9116
zba2c3b11ac188e5229d24092b4024027bbe0bb922234e3c7ffc21c2724b9fe697e33028e947f54
z71d86e7836141f5b296e9adc90eb71c7b3d9841415c21754cdf43e0ddbe2731d29f946df2722c8
zab7fb2c47584794984640977c38321d3f88fd2d12f21f40040024a5f199a2057dbe1a8758970d5
z1c65de49707ede221a7239418c83fc93d49df806771b0631af43d30ead9f6d8c772e9207d7fc48
z0dce491de02679380de235d16bcff0b131c1d3411ef7108ebe0012bea661f1185a4f9641c8440e
z204ed0ee9142fcf05d7349a42fd47173a60340a040c09803bf2bfa6c9196d22b086d92c03960b8
z8baa33b782d252a9445ca953da764ba69197bb42c738e9b9e5fe536a875b7c48e8cabfa395bcc1
ze4886ea1796c1ba8d5c5514aeb9dc8ca710c94c1c765059adb6cd3f12894d653a6cc2f44e37631
z02716072cf0f99c5f6e4b4bc4743e52f5f19200dffde146b3bd6a2eb760cbdfc792fd2ef2ef87b
z498ea111e1c5a7e7916fcaf4934343473790d6c338a7678821bafc6fc65049793d55bc7e4bc40e
z00a46c4190165a35fc940c1620744ad42f1662cffad5356e01fb64da454adea0c76764e7659747
z97951b1db322ffe73191be0c302971014cd19d0e46abfa597258ee0fc4a59e5b315d31e1922651
zd1d63bc2d64e1ba85617562d7e45b9814404649fa062cab36ad5bb2675d0943caffcd6bf92036c
z0f41deed460cd7972ddfb9304e17d8b9f79293db288bc9710858ee6bd969387abfa23b1e3bcaca
zbaaf4a5d69cf19d48acfd3805c946efc735f616de17457b225d24b144c0d0a458adcd68aae5339
zf0e519f626b35acd69c49664d3440191047a7b0f264177186e5bad345a7ede5dae5d4132590565
z6699bb438dc4107277c82410548521918cc81bf9eb267755f4bfa8757400d73a5edeaab5a8ae3b
z7e4a8054649d1fefde84ba9e0c3be5378f5995f58b9b09083a61befe17dc9455f60544ed19ac7c
z02ce96490aa0cfcd71826914c8369674a79f1fd48287839817c343d66e39cdfde646ea04e35190
z69a90ce4f85aed7ad96d74b3787c541543c867f420482671a3f9144bbfd1cd7eb2a2fe6631d190
z379c6c14658f0d1ce034b586d3d745542b0ae06af972c08b1eea0506d967fe1db9ea1de6ab7381
z18bfe7eebf9528c07027d86e0fb872304c3ab00967383fe52ba842b3125c309b2c276a85a0cdb6
zbffe9a56736e70e102c3e56a1fd42e6f24b73946609b139257a63f54bb830198251cf6498c694a
z99dce1b11c030e4845082cf55778bdd7198ddef898d691e35a60427bb253105cfbd1e49219b921
z4ac31d7da7f1d31ecc36ac8fc0ee0559c04ad185a7bd38943cabbd21da3c6686592a56beb559c1
z1eee1222f5dcb061df6c0d67ed288f875d974f45f29cfe36dd8c956cae5e925553a7bd6b907aa1
zf7b3538da38eaf9e013a775bdff148d0e2eb19f151076c0d27bb15b8af2cde49e9f75cfeb8b38c
zc43b53b9df9a75686eea50e0a0e1f78a539c4cd41198bbce4065c52db49df3d0e12a365a4a20a4
z6100a80e7e46bdf53e8dd500fdf6e25b87f32cdba1977a5512bf7fba1f84540b39328fee9b3e3a
z51368e5d2cf68c0f6489d5804226270dbf5b8028ee7e3a5daec95248afd13aa746172a4e228f6d
z8e18b1519130818fc9cd2187eea3577a5d64f3a38eeb2943da58b898fbb30356aadf86a9a3a185
z46fd46aaf576dec9a35f2672bc172bef24cbcef0f4109ffe78037da80e0cf378d6ac95ac755e78
z15fc34c7a99450adefead36d65aac7bb72807a2b8191d0c7479df5dd2e178f2b0657e3ec174f15
z39074aec5cec263388986bf9fde4f031d1fd8949c20bf812cc10cd275f2f623a55e7ecfc416a4e
zcc15377eca0c06bd927e3f887992970ea1a7c4c770bb912fc353c18da6e0f3e8b0ab1b83ed0ab1
zbea57ddeeccc8477c622d3b0f3fd6e9968a87dbee3303db0ecf97e54641b4a41bd090e55b6d95f
zc463f4e6409c0970980629576264becd540b8b494e5c75460c25b4524bc7966f2f622ece94dce7
zcf461783994298e1492491ea110166406a197766193b5c07825786fec2ffa7ffbbe09f1987591b
z8ec8b23b7ac0b9d600d7d3f305929dfab17385f468deadc4b6a2cce38b7dfca302ce4cd887fa90
z7682951eaad58b80b6f3d4d2151122ae53382f6175d7aa65abf0f63313ee5534fdf482dacad0d8
z8f41db6bb6404ad66c499f41f0ecbb63c08b291f0bac710c8d90ccce619c7e2f8db88b920eedc0
zbaf61a21fb24593c57e0cef3e99aa5bfe50c71a32a3d54d63973eef8e7df452603aff15bcdfda7
z1068a07dfbc491babd011e3cc89edf7257e089882697e745a0c87d7c63175abb5008dd83e0f545
z92e709d0168ea734c5fd4ea4267cdb3975f2e069ccd8b48383d154519dbbb1dee71be37c36c919
z3a4f6c9354d46f2d99635a3c36c5d0ab3706c199d737f767c5c2970d4c4c0a0265cb8aa23e399e
z23469b5132dbebdad81c5db07007cca731c12ed9db5490f06765750d42dcb1b86a9ff72ac33751
z1873fb7edf626698335833d4fb6aaff8575dd5fa89fc6e0506f0ea0ca4eefc66d9eaf020cab652
z004c7c3893d1fa4564711db3f9bc2c3c0f27e029b0e0e0fed21fa4142c22da5103caaa20bc2e4d
z91b5feb13b0c4ec8ee6ac806acad3e1b285143fc5be53ae5c47175190d7f4fc2161c4e86465c17
z40935a3def6cb74a3bfad6c6d5f60a3d750eba7aa58c73a9f3fa73c4f819bbc3e7503dd1a62ee5
zbd039d810906053c6427728fb056649602fc2139c34c1fca09aa9525774ce5fbd086a64575aaeb
z047d21d7a7c167eebac3c547fb540fb6ff7187c2c811416d2b21d2477817474a6f3cb6b673fe03
zd7eadd7e465a69e8769618633b3d7d6c0b52cb981a5880c7af5258b1e7ad34bf20dc56ebf8bc9f
zeeb723c9968b6061e1f979dcd85ac31fbf258511923313b688ad6615cde7b6b16a7dea4b731ae9
z99cb6de2d527c6f6dfba142882a0daaa80b2fe9781730f954f4f2027459d95ce40c5548aca8dee
z47104a2d1274ad36c474b8d71ef352f182147a603276a853be463d2eae74aa62a663b201599f00
z4eead4243776f097e41e97ea049d17060ee108e1592d73e99e21dfef2fab16a9f84504322cb47a
zf5cf7e267338a830d3b6ad95d186e9bc6cca58ace04d318928f8e9606c664bb6f37d260db59b01
zd35d5842716ababe4d4e3451f40dd09051e3f82c8218de06e5bcd85d20e696f1c872f3a5858473
z24dba1758fce056499b8498a0115425a0c5bc3964ca36a7f3ad89dce0e8b50db26261fe31f5b01
z023bcf260f663183dd308ccdf205aad208a1917dfb4ac190064ca0c04b03869c63e2c93b19fefb
z08ac3d6d007e87884b632184c3ae96b11c3aa9aa26d702844f39238edbbc3781748cad6200ac8e
z1942fb314c0e11fcaabddde0d0cd6dcd22433c2dda0abcffbd72a9bb5ac3ba2342b0f9833491a5
zabf0134231a5d5c280c74c37a27991094a6c3544b2ff7c0b8fb23a9b89369ab560cbdaf55a3f79
z62b569ca809e591449b23c6ea4abf76cf6ff0b9381fcfffbdcbe0b7546505f804eefd615cf8f06
ze1a5dc4819788d720a6bcd5e75873103e599a30e3d6c3fdc454541cdd1513020272969a55df2fa
z0430fced67cf5b95f2a7f69cc9930b63ab172edc65ab3b94ef34cb07c4ec0085040c3234057dfe
zf0b25130ebd905971b0f77008a64c52ad8fd4268414cf50f8dd062b83ea1e93d7c894a29310b34
zce3302ebc2a3205540f14a03e680236f97beeb27fe3164ddddd8d9bf05b6ed4ab213bca32004d3
z04e3f577e5fd68893056d34e90104846be142b68d19a97e940ef0f4fa814fc0e07d82494a681b3
z746acc24488b9aa954de7feb45fef039cf52955a7d1179d82559b315b341cad35b19d5431de75b
z5bd4990ca0369d3ee4582ce6fca8bbf2be7e8be20984fbba3beb96ff5942da37f717b589c085e2
zabd34b874ba4859004458501aa1f1df69eb7815d03d7499b574baf01e45a536ddac6102c8f6253
z39aabe800b88b1ea64937bb26086091557a9cb1d97c9cbb09f4e443ab340cf983ac2840eaeef19
zf5ec10ee8b997d54c60afa778b7144cc60c8bda9b7ecf48d3bd4a5e3952df5b5a04eff84936486
za0adc429e7eea9f98ae6b683ffaa00bbacf3aecf32f1791fee27b19f2a5705e90160dce60e7277
z2de74b02960d33ab819af054770615e98075c2ee3efd2e1e2d0b16527c1287a56d13643337c9f3
za8e401282863c4a6845c56408258f690f579d174af709eafb155a9792f61aaceec4ca82c68250b
z151c6d8ab89231f48fa9abf80268a4882c15e516b5a35fb31b1566dbe3b9a09bc7293e1d411ac1
z9d1c6c73395a3657f02ee261572bbde765d4aa206aa143c52fa5daa7081b7bd6673eb87ec8e889
zf0c39b430da9b999abf35f31851d51b71d924ed345415a0daf289fffbaccfc4927f067c9141023
zff82b11b3ba2c750b16e5511a1341d0bd252f2a6bc89a195558a296c410187bf5c7f8461e38528
zb0ae1e16fd5c35c76464679fca5ab6e8e22ac0cf27e849c4afe629d310dbfa6e192b1415d9d330
z295a657f742249779e443d1a5fda0bc1024a0750c8fae03192a9751c2d0e0895a708f844377a5b
z9c76ad1c8e7b36688340bbfc74463fcad89444f2d43a8c88b12490e91b7811171e804ee2883396
zfe6f1ae0bd7bcdba6e49e7af9121de73c3c0b5f6ac68825bdd72a9d215a21add4b32c4eaf640ca
ze16d81f385d9d92409be843c105b468750df82a668309977219f76ea3d0544c05a31be8d62a985
z405854785f9feade2666408c7f76e4f1e13ecd675ef69471bce7591b4d61019eaead9f40d24321
z402a8f204f639da9858f9e83c0ca483d0418de07c2e88c6afa41027597f04e0f0379df4adcf1d6
z263abebe8f7cfb6a896fae959bfee40733f87cbed45a98967ce1aba52a2df549eb3671b05ed327
z704a7de2e8f10a88ddd7e3eabd15c0960846f0c5b4b3f88bc607a3777df1c4666bb6ddcc77f86d
z78971b9dc2f5cf78a9134f45ea75eaa9693c3caa8597a3dd6ba2b15b7153d4bf9016d32b7f9cbe
zfd93a55a6b3c72e5a8a0b48f962e7708c9a39cf3acb2f97220e9e086a756a18b6de9b85f123872
z1f2f2e097f8d36846629f90f3bfacdd07f1acb409271ebb2ece7a49786fe1547e0f7d2ebda6934
z083c1472567eb451dddccf105cd7e9156bbfeb7c600d731ef6cbad9b100379214d1f632c5a8023
z84f67539d0a4bacc89c4446a0bcdfa222dd1fbc25ed390913279eebd7bafe9eb8c035ab8d80a5c
z7fba8446319de784b662e208d7813b9dd5fd0cc7d4a48c4e991e388a0586608d021d2a4e84fb4c
z03d70ef2df3495ef851dfa21289e5850b22175e45913edca23b763352c9fd345f0c1d11c092580
z78acc7513b7f99b6c8b6e31b06ef31362b537ed7ed4de193cc4f8c53fcec56d91954756a30bbb5
z222e5f3a5c8f21acff070487e403b2fcbde5ddcc38dbced2c46557a59d154e1f83fdc261f1f5ca
z8568c6d7692b71cf7655f80c739ae707f2c0d65fc3e13a44a507e8c29c44322117e3b7d5437fe4
zf1dba7121e52ed096aab39c8589e02f707b1df56c9866dc9420212a9e6cd1df0c6f53a65a4efc8
z5b8a313c9c179bc638a73944d463141f5ec5b86a7062db2ef18ed2ce0c92c6f04d4ddb9355f89e
zaab0df08e9ffcdd7e1d76553a69a85f02fa9c467244f2d3e1b9d3241868e2fe1e779b0db75d184
z051f8d3ab60b5a78484518aa7f69832e5e43a63745f310324fd36b90fd73cde4a74835bb679303
zad333c2abbbeb5127b0db1b224d258ba2f1ee08a89ccb2795eeb1c3b215e0f467bfe74e38d43bc
z286a0e64af01c68e7d0bc207a5464dc1dfc42e83596ab246b718d7530e27bee3f5a0d605bcb409
z90b5419d6ccd49c6dc5843af783ab2edb5b5d9c2fbfb4cbe773e417f0c61073ef27b4c02e9c805
z065598737a36841bda2c9331df27b7a7e51c90e971c7203382fa74a7d9ae6fb4eec3a5831fe36c
z8a3638912c3b71dac93d46ecf62d5d4c4755e2c0bdb7ebc4aec0784e40328b4c33e30a8f447114
zd8fa035197c0214969cfc1c95bd38ecf8b35389e9d402704afa6448a29d2ca8b06a4a640d4c294
z9d8d68930b4ed3091042269304a3b52810d3d9ed4fad5c0f255dab3eae84b379c9db12ff0d9c31
zf863aa6eee967844832f8b85cd4f7263813160cceed58e25afc968dec3e72dab8b1fadcc4e0939
z74713bde572e3fdc107481293b97b5efefbef785c2d19ce4a05e9d635cd6549f648c4ed449cb79
zabc4c38c0730dab2379b0690a2b57754aa23d4bfec554686a47bf1f6a45295daad5fe0dd309441
z2646a64272c8e89b4eda3673c9a8876b750936e6e8373c4a84914a257ee70ec3333dd300df5cbb
z275d5fc4144c40d5000b598160b531081ab76626f0cc80eb6bba02c918478d6f8b50438cc13810
z3945b4b45f5c40493e123bcb080cf8f45bfe11b71f8506fc2f16cbe401f70c3c68a52e86c35742
z5c3d9354d15fe3e29c8d0b413e51be33e8d2a84951b5beb2f830ca08f669984ffb796027a30567
zfdb76319b87b4b2d31bbd7e2cb75dc57b417046388d36f7cf19dd57fdf5140dc966c805bf5bb35
zd7bbf5851531ac9ad504e8486c1616e54b9491ae14cd7fa06bef090f4a59cf0759f37151141219
zeb697d332a450cb6303631eb60d0fe0d90cbbb4a70e8093bb89caff2e11aeaa37e0c81a902b33b
zc512afb88f735b7e09fead86c92de32b825e3736ba058c13d515c04ec7248ef2215259e13cbeb3
z7446f324c4333b8ed56152dad6efbaf1c211d96d5fe429eff9aaa238d7995e3c6c62202aafc441
zb217bd66db000a773cb928a2b99ad045c7f359acaa2458e87425b49583b6a69fcb37256d717527
zbdeeea4420c8e782af7f83a72aa2d56269aca5a6aeffd27f4fdad57ed0f5a52447b5d77a88a7c7
zc0bf03deeab23e12c497f1b1154037ccb1d081c22b50aad35e189cf24d8944dc0f5505795202c8
z18ee0c5cbda3a20d8f0b225b0c7eb2e59be2e2bffac450f2dade775068e6429391819108744670
ze649544b282b99dbd39f22f927097c98b59d69ed255f12ed749fb8e31af45c7c920d6457531d30
z00182c52e933bc47ec724aac26a12bda4ffa32e320e024343ac9e3411186d0b649a54cf9c81fc8
z4978790d51e7e30fb71e346da6ccb2a6afee4296a2c57c0ccd488b3e9889cba499775adef1b81a
zb2919914ce3500748e9d70d6ff457b62415b8f730567d1831746f710611a3bdef8188c4642ba4d
z488410bcd152889db31369cd965b526fe6a6401505092cc52dc53d0210b8113dbadf06d0fa3626
z3554da03a9eec3f10bdb318569f4cf4196eac92146558f830b371be9528a1eb8257e2f84c3f3cf
z8fa319c2378c8dec4e95320729a406ac375e316461987d8bcfd26f5c9d633cccfe0615b04753bf
z9fde7d26b5126d122adc9359bd54754854530a582beeaee410365e48c863fe58d5f152e17ce8ab
z7c58034637946902b4f39382bc97dfa506e80038c9f4ef47e0f4f2399a1ebb1cefe0d748e2dbd9
z144d0ed96aeec3704e9bd218b4dc3c1df4a1a12c03ac96e98527c7f7edd41bb156b78f40731df6
z0c70d83699b2e9f47291ec7911f24ce8c4c3d20444497364d04ef45acd36cc48ff0e1685d335e5
z3a6a3cddb285f67e0690b53faf2958348751f7227c7e97d2294d20c3838f7397dd0d775d9e0b82
z7da5c6e1d114e3db7d109a8b997bc72177169a484cf0a833a170a2dd34ba374330186760ba6f09
z33e4f97b051cd13a2340246e5a458e76d99e3e8d8040bd015255bf2c5743d1ef1fe25556db9678
z9327145b61c796c81c8d9a63253aee954e1f69fa120684096e23b848e61a22265b8b2e2e17f644
za2ad8a9f47d18e1929ca9af761affc77d9dbba3a95862f62abc9ff897683ef0930674f46210646
zacf282743327818e3c0b33bf341a27bed98599b77489452bcc4dbda8775ee0cd01a3b0a92a0f56
zbc82e8e8c9bff21d3f421b658b014c9c060d858b2e813021b157fcbf3d79dd94e557503a1874f4
ze7cc9ccf4eadba2f23c055df8c5a2d2eeb0774302f78886af73fc8194b06d5039be83ef4e93c52
zdec4898afd3cae8be8644e20295568cac7a3a782e2a8f837d7e4697b2f41ace77b77ae73397e7b
zd90bb29b8fbc33d47b20403c638f7b4ce1c05efd7634b67efa99aa3ad415b6bfa66c28282e3afe
zf53826ee6dde37bfd0945f10f92bf5cfe436a5f07b4b2aca14c3f8fb0f8f482c5d5bb14c743185
zd99857c26cb6f003231a84f1f278428f93934df3d115d2697cb8b71479aaf471f7155cbf85d124
zb456de3db1949963a6a6d23ddfa42e2a50e2b96e81bcf1af07bec670324371fad0142b42caa4a3
z575aeecb443f4784c41decefa608ad356eb1449154eebfb9bf1a5cb37f8bf2cf7a09b4c0714678
z77e72ca9624e334c74ca960cce0889896ad249e51030b611bfb97e0842ac71e882c8fd2482caa2
z33e71a794c37ad8c36ed0467252c84c14d54a591daa1852ceee1ee39003c302004c6f9a4ca53b2
zd148760f494ef73547b21e8be9f4b25eab285d260b857f8cac5397ad1e3d8ca55ce3cd04a61daa
zc6f66670ecd436601cf3b24a788db406c5c8305353342a09f0535e87a6099f1a4b397ac93295ec
z4db6c921387e1b65e607644f3e4ae02eae12d2bea977e468dfb2a166827f29ea85e98db9e71a31
zdff90e1387c3f31cc9672b3dcf90385baeb165aa4a2c11e70827b65bd84b06dc159ca5a398c06a
z9eb52e53acb9a9851b56867838830f5fdda4d4449a4cc2eaa4971a5ecb2c029af5e5278c3a866a
zc86d0c6f00d022e079c738287e65d1b1e23a37cba554322665e04f779f42163b7bc5ae584bd13b
z5dc4673d7b3c56fe2feee1c9aa4003dd1dc09261d3df005ad0694dd36b73642b9380693432e638
z52b42b24dafee690448f03993cd454495817f207345db65a3436464d068c1c6ee27fe048b21e4b
z862683771593776a03456846cb1ae348ccee0c82037402340820ff8d0774914ee087ab287e7920
z1e3ffcf425fbed27b0190db0e58ce82647a523daf5c4204a77b2e5f128e4419f60a54ecea028df
z29b688fd621e24a65d639232eb46404530aaa1d9b023356d5ba67c80343aa8918ca0f6763a381c
z1b74ee070008fa08e633d21a49842856e7f817219545863daf14e44dff43bf5e52b7b39e1e5371
zafa267585e8a4a6a6cd5507671925cf129b54c01ce626c6d218b5df75cec8643e3a1bc697f40d1
z8955d8670edfc1dd7194581158bbca9a090cb98ed731b8c5aec815edb2e7f9c8c3a5816616f923
zbe097b4abaf7c78ef9ba85df1e35ba51d40c95229613209bf47b4513694cef7ac1532920d8d6a3
z897d6d469a3a46b0a81b3fd5a76afae09fbcef6d836f9e367fccc42acdb7f04e1161bcb6ab301a
z520ed4da1a5bab6495f861b94d43ecae2ef63b57d31054daa2e9c0dce1225b68d6f5ffb2068380
za586de5d0db7e7612e211885779988148912c1f873d848c0c3560ed1d78e30495bb4d9fd0a7177
zbf7db62dcdb1685c177f85e70b071002d35032a708a34a576b552ebe8ec8351c1620a32cfc02ec
z60b3e733002d9dc3ce407394891fd1346f1bf7604b2bf9d376f09f55296a015e227e08c6ad2970
z57b45cd2d47d4bb0f1e94c9e8a84d2f51d423f6ce564904026b2df37a8b612345b7470dbaca518
zb968bacee9ec315cfdea6d708e986b6c18115267ca008efdd0ba7ab60ca662275ddb920ba48879
z53b762780f4c9b63a4f393d60570039846f2d1174fc0dc555f611ba27fe568a3c83f6a204aeb4c
za65b00c4b8419e22838fbe3f4e25698cd992026d79cc37055442475897daf5f23110d26a0c734a
z010f23524cdf6a9b7ec7923cc92a746f500821ab5fe73251112216e20d6894355f7f6aa5a703a9
z8855fe1d74654448375ca7ee477a310bbdca379f9e48603557540c8f0a595f20bdef3353cf21f8
z940a9c560684b3bfe4962db5991d32d3654f195853a7791765a88a997214e39f8c70719e48b83d
z55a385dc720c80e3e7288caf9ed41278f40c93da5a22ce3ad9fbeb64957a015f9aff36e7c27601
zad12b651934bf512c4750625efa3e5c4da20a041db2c97ffc9d1376667bf195ca168bf5c58345c
z6488accc6f2b9d0522bc4fc2a355a6ceb1e8dd16b14c0a96ba18bb9f924b6ad68780e5bcaa8e7c
zd816f4f48f38eb3aec578e3d4bb10dce7cf9383e3a77098fa9173652b1e96d8a569815613c168f
zb820378209822b5242babed532e089c9c11cd0211634ca20a5a25eead166078378223cd385582d
zc7be781850cd2fe8fa6b28980cb66acfff28a28624bcefc222f35ee654a1ca887c352be475c9ad
z1ca8a71f8928222395b32e875b219caf82f403af710a89681666343f648e98b5f064aa5bf85594
zddb3e9ff47045c66f33195beda730f3958d9075d40764bc15583d738178e5960c96dab2dd577ef
zb36b8d03d8fb4e3bbfde787beb7a519232b2829ffe9f43b0800b6304640a3ccfa9aef23bb76d97
zd0a5a369a8ebd17f694455affa154afdd35d1463ff872ab25a971c1ea9bd0969b388879f9918a2
z305aab816fef10b503e3d9d38a41ca09faa015712a3675b79cab7e458a35148d79a4236b1b20c2
z876cc867bea5438a8d170de4b61c196027523968e11c54223499fd3aff4913326788810faeef0e
zf7aa21ef7d5f86ae54cdf616ed7b8ad5fdabf608a5c8644829cf4268f3006487ab67348837fb51
z0b63eca9ec4ccda18be15123f99441debaee09ce24c1a71339f51f2ab80454cf378ebb8348ead3
zca27fae3a27beaf961ea9dd06f35e8e070eeca9a4b1d09b079fb6b5fa8d4ee1dc3448f0c451729
z440a0b0b9489d6aff2aa8421e677aefc9285c2dc6801351d260b9d8423ab0883bec608c6bea009
z0757226655dbf95bfde030a97afe2a86842ba199d82b773faae0677b1b4647ead1c2a291713cd5
z1f348fecac104554852cd39a901c52ed12af09dbd21261812b8a4c094741041528ec7c7b2298a3
z26755216de8d2e766c18920638686fad87af2cdaa3696edede85191e0130404988ae2a9668dae0
ze2882f84947183158ec670fa4c27f2b2983fd3c487fe2a076dd49d0b1e703e016298d8e39795b9
ze73bfad7ddb3344446a42d5c5e39c13a16007c9d082f59042d3e4cef3fbbc4925bb92bb27849a3
z0f6d29e4074f8699d576c29ae1c58454f2847549254a1f8700f064b13495a0d91a5a27c6b9f335
zab420379493671640cdf5a6dca93cfabe8ab6b9ca66a0898bfc8358179f28049a045460b96ca7b
zd2166827c812ef3f4ed86efd4e68e0498b242101c8dd3945661c59a9e84d725ec8ef0d89a596dd
za0b8adb59d335212ca9638576fa89c5887eed35ad4078da053b51fd9fa805d6d68cf64f3174844
zf856e4cab0a3e93a0e7b33ef451bc697a4700022b92ae39101be87a501b53c4380e620b63c5a9a
zbbd2458b6d1da6aedcb29c957356dc0c23d98274e85dbb4e608de90cc2eb648cc270852c9d3941
zac09b145ba1a2a0e04db13dee4adb0934a1305f722faa3b96633411a5a88bad6021680692b2ae5
z1a76ebd7291766a0e695013e487d1d98b83b7afe0c48af14b964bd4bf21fa00744cec1ca9054a0
z2945b21e6bc4e2d2332d9e7060fd56c99bccf0adb96c9490fbaf12f6ba6fc8469b5fd9498dc31b
zefc7ea14461b795e65a74082906ecfe65959476231605f120a3f0f24bb7d24d43f8a4eb93df2c0
z75a166e9f6c1801ee16b136ead88a2c8e59e77238ff68a84653fa40d0f167a3418559a8252e28a
zd6a2eea98b967b32fe9d7091d3aeafa64c2b792d7f6ecb47070d4a9acc5cd2690f12bad1d92ea1
z3b628a7f771f2bfa801ee91f2da331d9c65276af7c70eae03c545f9d13769a560bed49154fa0ea
z1316bbdc7f7da7905ca9037b7443ed1556fd90b8e6dadaecf4cfc1516de4d1c2674bb98e8a672d
z04bd4f01b302917615e93eeb20459a49b811c1a326b74fbc3675c9eb3aebae9d6fde34d9d60c97
z46264c8a8367c0ad749fe1fe49a18407da1610fa67007258bb1be3d6d4922ace18e35bc3b6fde1
z195fe440cfbe3b5c3c50b7405b35c644793310c4c524acf956db81941d9a883329e18a08a8424c
zc608d75ebe1865cc03662cd51bd6f71e16727c45d287f807f1751ab6bf570d952da7548e0e9c68
zbd01990ab8cecac90e3e8cb6a4f4974c0d8c1d56b316f1693f2a8b171bfa9e9d6d7e5115a7a4d2
z8e280206c9d03815d35429f73a332dc46b70a90fd132f15b497c7ff3216a81a4f9c48d31f9bd83
zc5de7231c90b89618133024202cc51800fc3fa9e61c3895b2cd3f1de77f5584cbb4194b97e90d9
z49c7ba4a122e74e34015d61965b1cf770d9e9ea2409cf6c2c19cb222b78a0a762cfec88bd00c51
zbb648c0d1e455c8e48513cf8589f8d1dabc10ac7ac85151e34b5fe5199e188ce68eebb878eb060
z5612f660dc430227307e301a89524ca5465601fccf5d0d18b2c0edf5cb1b8e9eed27c9d2eadde8
zc826d4ff58d41c9b0081c4caea187b7793830adb88ea46a7aea906ba4d78e91250cc3d519f5426
ze9ef04d0ddacb6d4f6d169e5522dd3eb982a712bfc09e5fd1e4347ac998b3bf990a6b3d1092698
z586264261e011d88bae78b286c3dac1309dec72810bedb94ef7b7dad5b55f2d1d6a8a4cc468a87
z03dc2f21a464a7cff3dad3ecc8c6ac76e9cabd751193c8ddea87da8d5d9e0487f18fe0e96d2a85
za1843f756e69d93494bbcea7805fce8efe89f081b1ac82968e9ee56818344c806c7e5885d32c0c
zd9c66187a8d7393b03001d80d018570d7b494af55459ad6ebdaa71bec6c21830d334a002f3333f
z19bfba6f8f3b15deb2dd259d44b8df3a2ad962d06aaa5206c50a6a5f2ff2139e72c2c94acda700
z7cdf6e46b02fd15c624d5b32ff930d415419c01e6fdd0102fdc20635a1ad89c25d57f2aa58205b
z3e4eda005bc29cd5706060b6e6c9dced92674897a4942f66fd226a9e62e3626df1522c820348ac
z65fc3020dbd5c7761e428ac73f374e20c7e71fcf234ad481c17d45a1dbaf708e28fb4dcc7f7e3e
z09d2f2662541299009db3faae704e6b9db162f5daa2fbb8e4a6eb8d30aff8c0bc3edfba0290c72
zd5f913b5235b1b50d35c3083a80f29b9977c16005386b353db7868efcfa344413ac9658450d299
z9febaa0fae6e6fd23f86a3f82cc6eca076011ada205ffe83d3ff7cf4232a186dcfce0ef4f6eb50
zdd2267d5d3567c02cd4664fef1870bbe5fb714b0e3e898cfd5db5f41f3c408ff54cbaa77db8f45
z16f22672c650248f08777ae946f25dad838e6174a9130e3e264b4e525dcb808914ad5f49052163
z0ba9772288f0f4902f1357cd47ffd96b463978a18a92fb8ffa2c3c49bc795db73015b543c8b4be
zf4819475f445b1753c6108f65d09aa11fbc9ea69273a21f7b25a397238ae1de10095f9edeb3cac
zc735e004940454cfd9c179443a6b385720101a2a7bedb9fb4a52ef6e746f8d70160ab3f3b6b996
za7b3a437dbe65b8eb7e6591651bc2c96476caaec7524a32fd4118e67acfb595d85ab109e3b5bde
za2cfafd939a8c5eb8dd4add2f51e1787b6f3425713e44eb70a724d95ae21f2362633819de00366
zd0a8f1c9ada90123a0256011a505932b72d164d06eadaf03c26455daf79ec794a383a68b5001f7
z159ea3a0240d5d831962e4e94e2669ad602f5fbbd09d748a31c55457c86aebafe8d4b08c2c3409
ze2c07a8d09427692acf867e0dee24bccc59b0352f676e5fcadc89fd4b68a3247ba1ed3dd79c800
z39129ea79cee8dce5a464437f7416c510bed032d619d3470b30ad5a9baee5c0685f4e56c78a773
z1632ff9cc544cfe11c6360e89f3c31e8e08aa0aeb220e15062020a0ddcffcb21b3939ec3691a09
z46fa9d8d7d733ae9608763816c60a099797e2b00712331eb1a3f47498769690e980b704b5655b3
z6d5eb05ac69769c36dc267d732c928322f067ae2b9e4ca02954ecf9b860e1899dec34dd0ce81a5
zc370a5034ba2da6d812de73ace4fecfa688dcdc5b7a1ed247e0aaec66c080c096ebb84cec8e8e9
z818bc613313018fd4aa7497364eaf159be45231fa9ab9e2e07dfb814056252a78e773b6bb57e08
zbf0f512411d8b8d06812622235a4fe92c58e0b10690393b142c91c21255d77a44b32bcf6c67b3d
z4f55495cd0c84813f29160fa5fab7522d13059304a3906c55e8bc166d32e47750388892157e6e0
z8cc5c97acec5dcea94315e3d7d823cacb58785f4bff87f6418a3f91fdbb21cd5d151978a52fa27
zde07cf7b371f5c0bd90f967b2e2d455ecd398b87464717c0af4aaee60973caf218d279ee0a1807
z5542016d0d0a7a8db845d89654d23ef58c9f431b4d100e3647ed48de4c1b944c2c40da691c5838
zb49578e482b4d9977edf2ad2ad9b4b8fa703a20e809d09d981021c889f9fed9025721d43fba6a8
zfa56fdc8b19db7ed4da08d2a013ee823963e92742ce09a9cd0a2b3b4cc88318bbdadfcb416aaa3
z27e24b42fa074cee9697a53968a5b5e4416c5da90375252ba52f976a75e40ecb9407809995f722
zcaa04af2ebf02b91e56a0a99a33d1131e82602aedab5af7153ac5983d91d41124ac914e725fabd
z703da932a79e032365aaf2607496e0ee90310ea956f4fd490f38879de85e10eac985560b8ae5f6
z5f843199b7a66c3f0cf7b592b731997a1d3d623848a708ff6bc95e5f5079822ff543b91c0eff57
z0e3f6e6ddd6be28ce078b367ef153b3cf608007a565d86d38e008ec20c78c8e1cbb10125435af0
z3bf493326f4d2fc97d2db0e3ff074114fb0dcc838220f727f66eb5b6b042ddc105654b47c1e8b5
z7d7def09cb7055e2d3b879ab572f7f2e7a3935fd26482f9ccf6dcef1cbcd0606def1a7c18d75f5
zb113ba39fa9228a11788e9ce4072b7f80792f5cd2bfed4a650780396189cde80dbce72ee0bfa93
z89ff3b47d850d86367b1cab24d2f9a10efd3bc45ec34188d0bebbb728bc487fdf6d3514b567ad6
z91a985e582968c8dcc712ad0d5bb6289791ee2c725d42025d1b5e71cdfaa5530a080e31aa79e87
z9958bac37f9396ba2454a0ba522f327c3c12fabca4aab07474527fca988f08e6b34c31395b2a28
z5a32e5175cb92399ad348f3452cc8d8d3dd2ed05816701abf1a740c57d22e03ad10d403dcdb2ca
z83f4b58a0f7b6f715403266eb4a6b7867e82f05f8845e06ae9cfe54673eebad6c391f953f0a65d
zb5b005a01d54a87d9ccc35a698a20b948add0bc8c5e539509c9806775321a88c57769521b22e49
z68997c4574171e4e9d0f7e9af2e5c743ea50d0bd922112339ffc9b6d42c17ad3d06d16ad617cb5
z8e620e5658c5422e9ba166408fcbb722ad8ee9892c2639a9a14f4b9bc1f5307799a8e56e710cf9
z236b13185574e82bc3c3f2ca78d1a726a9dafce7f7967ad1bce7a4769f84876b19c56d00e2ba10
z6e9a9ca13301b7b3bdd4c356d2881f60de29762af08c87cd7f72a373a982cda5d1dfb2ca0c95a0
z99696d3e66920709cc362076fa37c67aefa4f9fb758d2aa54b0ba3a7fc683f3afffef9851bcb56
z6984d48835c2de9c5fc8ce9c77fb82658693323df497a3090efa4c67065dc80ed3b66c5e07d4c9
zaaa254c481927b19839a9505f78da9941ad6537211ff1df5677588b9591bdf1f65aaa3cd726c44
z27feeaed40df53de338a25479ecebe89cc86d800f7aebe22ea7d4bcdbc894ffcd8c3b6673f7ce5
zdbaffcea7887b820d4e74eb9a1f552cb48165e242f511821c3aada139373c223df5fbe3e79f6b3
z549ced6ab24c637210209be3e6532c305e4822a19f81e7d2df16422a29e4bac274e8486b8ce58f
zbb985a8c4ca542ade1b6ec99dbca90bf728ab2641f8872ba22a09f963a9021348013028479aac3
zc4c03bcde32068a011ec2257d9783978fe228b68be08568af210e5a75269157e4eee87014a8b45
zaf90214a9ba89867bc2fe63ad0e50816b85ea04dd04edbe0dadf98f8fa64c943344347a21b5562
z0989114f2085b7adf551dc9b879b4db281aadcc722d5fec394d9b61903f2c0e63d1d11b1f29d8c
zde119228614f3a87fe463411665bad88545592f062b320d045c876e70bb6c3abf26f9a72c8644f
z139d7c91717469966587070d49c27a7c442bba086529dc1da3d28d34e8073fe32e4b0af4e7559a
ze69d48ead70060d589e808b380e9615a4eaa79dce8fcc99d2b55d4fb528f411c7a7a30ac8f567b
z9aee3b50455eed0dea443f3047e857a3f00343a4cbf2e4f895d54c4e2c9fff770b4582d31aa1e0
z6e0d0d49ee6a5ab9493e72bb34fbe807e351d6182c0304835417dfb917dbf07470c04a7d5181b5
z2fa83de431ef4f61d005cefe6434789553463530cbb26ad98a3bf69bb0e2403bf4bb88cef19017
za55df00c5b513395058adf4d5fc78cbb06b9b97e24c24353d2926e23e2562615b3ed8efee310d0
zb1665334cb6826577e5542b34666d38ee71c9152542fcabfb0c1df3ebc06707700e9e0b848bac1
zf199f36080cc63453361249711912733b2d2e7f1502e08b356c2e4fcae2ad5351dd23a51ab437b
z7deb2881ab80abceba6067052cfaca1909e24357b780d1ea162ec7364aefb873d2ebc2139add4e
zc7164205281f27cefb4d100b5c033af93ef0f0946ffe2744018ed3d0ff81dba94d2d891209fa8b
za38415d05608233a2e24b1a48f9bbf6a4931ebbba661eb497dddebeb7e2119c24c6de46569b925
z9a609b323a4e50bf5a1173c03ddb9d57363093a8b5946328f9b51fa3fe4200df7cd694f47b64bd
zd66c9c1bd613dcde84a229929711923dec08ce9af05d312dd506a10e7b8ff916bd7a16c556a752
z54d61e189de2aceb9b2ad72f5879df83b06d48ce74aecdb1e154edba05fc792f552fc0f258ef03
zd88975a5b0e0b4b8bf17cd019d011858fb97d5738af785f4f2583b26744a88a309f8f4989d7c29
z2cda71681310f41314d3ec9f38cd6daabb92b5f435cadaea848e9806256d89731ec34a291f19ca
z6f04a6505414338bd5301b8da163bbc7542e4a60c683900f021246f3f66881a7e9c6f80d60773a
z78e4802ad5d591eadac734fbf18cd129d67f67f4c5d9280ba02e1b367715e27c0982e7cb10bb13
zaaa2304549658b16d5804a79572a3408da613a79522566b719e6a4851e759b9ddc472bde5c5007
z13bbc07bcd5450ca5b21fcc6d706d9005fd4cb244efb14d81c7cc34a69516355e2d5752f1692b7
z34af7ebbd2ac8d70ef1a2704f67654907fd95bfe8f266039ce8e6aef681e06b857b65be8ff7fd2
z15b9d36778c42b22a9ead92f1a0e1dac87af2911408265db36ab52deb7b47184f63b1099f1f770
z1d86342831eb420f30df486abd383e8b754c6f6cd26be00a7766f7b434d04dab7b7a26c9908fd8
zcb5196688e6213980afff67e3ce50445c6c2ae782b12a99e0077f84455bd4bb38923d5d514024f
zfa3d8eca0d184f9e8a0e08e3eb972df3e441310ccb4cf3242ff9d38c8451d6e89d963c840100fa
z3651f389cf59836370b59ee9dbeea2066cd87d9e95231da5e3ce4e8433415cc9343fbd95be3618
z24c339333d3e1d6815abfdbe8fc545a1c7f16921086ae76cb08aec3ac2f9941593d72a8040f7d9
z6065a067aa5ca27aa3743aeaf9571456aa1bd3560eeeaf26333458209ac34c76d4577752eb3c4a
zc20a50b843a32810e6e7345781f90b5c833c4ce005adcef012ccc571b389bfbab93511a61e1f98
z26410e85d746cc095d2dd3db280d69c5174835f20230f101ad6f262e6e8368d84eda679f07bd76
z9f28a4522cf9d12e4a96689711da2149003d0d3b0dfd64d239e7011a1633a99321f4e322df9cb7
z1029d43af92e6a570ca16110e2aea289e3416a38b8c1feb8a809a349d79c74a478ae95e4dc777d
zd5e848ab28bd20c44ff043d2daf6f5dc7e4ed2f29a4ff4a36f3804372ad4b77a21722f52793b38
z710a01c24c6083511aa22ee876f329daefe51bcc0b9c7834ae1ba749ef2791dd34fff130846c07
ze920a8953dfdc28f6756a5e637d284f372c3d2ffa8871f85699eee526db16da54a6b1156afb363
z29ddd423e2d561a5c31d69f2b8069eee5be77d4b6e54cdfe157da6cf7787943f989b7180600b8c
z2fe75f5394a5279e36f060e0c96177a4249c7e601a174778be710b429de5376e42054d7243ba66
z79578473b8febfe23eab53fcc3ddc0a54e9e6f069385b3a6a6aad509699759b5f95e16db659923
z17d9e0d3023d38070baef0dd9eb751de332ebaa6aa1a3040363c631957e7412df9bba8b559afc3
z5ddc3fd481e68d8b6d5795787240fbff2e6d3d4d27e8aad317179f5bc8b264f96b85b21be7f889
zeadf409ce678230f7b82159dafb8c675f4d95383f5e212c0aaed23b8e8e6806c9b270b508d00ae
zba2868fcf2b355339bcfaad02fea5e6ade52aca7f67a75e1b85bb1c60b9d007feac77a150bff13
z0171bf07c705401b7b3267909f7bdd558559a97491f83d4cae1b2caaaaaae6b22b48b271ed6bd6
z005b73c2807300332aef2bca77855e964d0c7e389c74d8ffb36b95bd525aeac14048d34d44a07a
z40e0ef9b676cbaf2e8cf39ff47c3dae150a2e424c470837c0cd500033ca7bb7768e528d3277a35
z70c9f9cebde3bc5a452f151a6baa22e107398add694c114f60a68f46f8fedabd5344319e7c708e
z3f45d4bc5e5dc31276f8ac9e5527ee4b9be208eaf754ee7702f6a7f8ab3ceb2899ea5af1bebe18
z4f617f2132ff322afe85db12b9b275bf9eccfd136b39eb91fce48d39612f80ee9128499afa1ff2
zd942ac58488b8c29424302278f3c26e8ee7ec92b97acf31ba7cca35e0d208cf66f53380264bc71
z305969f61fd0d6e5d3724bf34f1ebb1f19ff7fa9aa9537b7bb557991a6264c51def8ab7f0a1e8f
z70eb52a99cb3daaad186c048c170bbc05aeb5528464e9ec2d3527c57f83b6dc57f72b9e47c4e34
z0dcc5909dee2a16e71a6be949ae573e27e2d02a2c4cd3dcd947c3439932b2fd692ae5b70e41435
z34c79e0181dc0c308a6b4a5fcb77b5d0b3367d78254394329a0fae028e0ec465a16c8b478fef51
z7a3a357c9749b5050ff9402ea539853ece187f0f0192a23a26c456ee34a11d2e90b2f53621f957
z5cce78b616931c8161f87ed67117c1568fe6c4eadac53cbb2e5bb1b80c589975e81f7874894426
z920f89848c2ba1651b825235f7bf8a592597950af88eda32b0357edec7d2f5e19fd499ba8035f1
zd628e39a58d6135285cf0902ae2997b8aa9d71db9697372eb7cb814ca38045d17631822dcaae6b
z774e51a7cdb77175d7cdf0c21fbb8bfa0352d4ec3fb7ded58ece6ec7ca63492b26e600f82819d7
z365926c7b65c82aa7c77087945ba14cce91c021f6d5292d478507453adf71a4f3054d347e0f63e
z33afdfefb93afc58bf8259732117799980a907e0946581a6c0fdc4e589ee8908ff742af6522793
zb94bb0d849e92f5298f36e7d4c25d6c5a776da83155acf98ff58952b79189c7c39c4194cb51e5a
ze7889e091f1a963e32a67fec296a693c894d0a2b52b443731fe01a2d51a065238053f4a48cd23b
z967dd5eb332f6f07cca94bc90da407716c656094288104da5de3cd212b7260759d7be57a8c192c
zc0fdc5a536d58596fb1f0b5b3a34746857cda193076626b75569bfcf0bf4525ea9bc9caec9e9ad
z7888c412c0d74ac34da57be82ac5b2828522774c4daf6d71ee30357cba00e244daf3370b6aa951
z1759ff8bfeb8dde4757791802f3481f973f371c67467b835d2c6bbf10a4ec084f068d3a82402e9
z7f1bbaa1566d4c4bab4ed2f82dce51b9d2dce42664222044950e12db69e2a08b2772fd7b812249
z44bff4c27dd0a45347f02a3cf96fc32e133ad32d67d71b1d468baf6558ff7f661acef4d5b4451a
z63adf52a7e071a102299b02b919a872ae9f71a13042291bf197404047d0593ae28d2896e26691b
z86aa6514bbbf0f39218d6fc211f862d9307c2780fdc0ca2f4f7511f30ba478c80a6a7b5bdc0d76
z780f61bc3a13f45452d57675b414f68c940e8a3ad5cfe8fd3a5e7a498e42dd1021530e1c3ff666
z2360c25fedc6fa3057216d76105d8d1b3923a2795c6e6947ed07c9fa440c156ca573b1030eb68c
z7b2619b647936d1af3fb905c388695d110ed4d9ab39f82b018627977feec9a8ef10db90b6ea6a6
zcd937018c883ffd7215f834dc1b56ddb2e3ab3c710485d90472c9046b697a13fb7b38ef0884a34
z0941e720538326e1fd385554bb4f88b73efc28cde0f3b2c8b33e235721763c89b107f155a804a1
z249f94db29322bb17afd891c56652df3f3ab8b43f4e84a585530ff451b7b77984781edd457420d
zb433999701e7b1ca8f367c7d65a1e923043671662210a5668345824eeeda4aef42fcbb591c58c3
z63177f5b3f293dcdfcf473228f36b90c5a6276c707b90d669af7e1c5274d1a28826b325c9fd65e
z5848f61cef36814300427af4a83bc475b0721f6650b3716f99108119c55876b43c6f020553fd55
za2598c52cfe929241052ed3f221a70de190df6afd47d0653c29e40dac18e41e0b1291159273013
zc83b325a1ba161c12cb9faf007fb82566d39a4646fa878e1eaf5e4092997581a019edc3fe67b58
zda72f5282f7cab550f8272744f35235fd374a6ebd2e0bc9b5a3ede3b1c0ddb9a47d61f6a0e350d
zba29d8063ff39a203ebfbac60627c47998987e21cf4b27e4e5bf302d2da0a37614fed18d6634c6
z6ae1ecb9be0c78d4837ff8d255486affbb85939c05350929e647251bb8be4d70376bd2452b106f
zb5e2d8816ea1b9cb9d60bb7a771449ca88d6d98d3252ecb33c58d884c9a250c82d340b74c553ad
z43f1b7b6ce02740110782a85fb2187b5b514a9c928a8dad36f930d290ee5c301b241da03196f96
zc2eacfa471ef4cccbf27e56e8a1e0cce259feb0fbdbc781447ef0f9d8dea3293f708165c2942a2
z32e4add79f9af898a90651a8034a3a2f53af2b99b6653d1b8fae4758ca326ea0a08f54946fcb91
z8f9a467c8ca110882a0d931091691e10157aece3380b78e5970a78d6be1a03d367aed58a2ed8c6
z1fd6c6ad78ba9496b593a97aa86a5ebe1b9151618ef4c941b6b76946f0c9a88f2d11f7ac81568a
z0029dabcfe4b8c1ff43d2fe0212054b3ddc8247cceac76e1d998afdb2295e82d11c2539aa932f8
zb9a59a695963720c3f987f6c401017b2078eca61007efb1859e8a5834b924ce1dab17d07ad8f1f
zf25098504417a29aac7e391439cfe3ce12a9888c907f7b4f02ff912875a7221aa06ee2ae2a444b
z224bc935a1c4b813ace7df2e26bd02180f702dd873ac36aeb4fbe648f61d8cabe7c8f4da8a6f88
zee2bb60bf5b2157e18785ddf38a2e70bbc0f05d78009a2fa7800003e63d081967f11664d8dc97b
z090f7f2ce1fdc75a69247f72c25d41ebe341b7785e00b71e06152c8a5b429e4e0b8d4339fe2b26
z9edf0af44f4d5b54b8e7bbf0a2d3d0dcd0f1203e56ceaf54f8f0ea787ce1235aa06667682997d1
za5ea4b081e07082eb7f875378c95585e8cd28a56cb32950059c630af9a71fdf9957642a65a3098
zc7fa1a16697a701a13cd9f27b0862b99a09bd64537a7752f9a6ac263e7d61d3d4399c5a28d7518
z4246c345a7b3622e7518e4e45442c26026358562ca102bb7921e81a12c6d92135cd1632b77b8c7
zd30604dc44bfeeb996631ed7ed62ef9f592b6d1aea04d3b517db3d056af5c9c1168f619ee8661f
z4ebbcc68bceae308ba4b631fc347063c24d2a3aa2f49e471a260822a5929f5aefa2fbdb35b0287
z16c05c1e82f5b132bf9daebb7a7b64c368284d022a9439faa74eccd84757479b6bd36b016d9e50
zdfd9c10c9b18684592995e918815a304ddcdaa51219e1fc3d4aa047f1042f23e9f5ac2e6555f42
z2158cb44742bc0e4878fef8e041dafca9a4046151a7fff23c94d2dab209e82d0745ef0e4091688
z0c428a91da971f60a189ef9b4df66ded0b74f6e6ddce1ed4a137ba4d11b0b25d6f3c4795d63d2d
z07089a061272d01a2fb745e8c1ead38b22fe414f6a8fef8595fd0404ab24c4bd3a529d04bce457
z7c19552febff959947c1862591e850633a51d8f7878dd4811e8ffe6f739e6f22a88ea6a69d4518
zfc2e36c0b1609fbc0c17bfc5080c75d7492308867a09c20f499e0183a73050a76fb95f07561f61
z47fd14cdb5969224031b94ad28a69974565a2767a8df9864f15d3fc66db54f35c3a2cca8cbe82a
zdff8ffe6d4379faac6b7aa5def230be845400834eccfb9181d97375ca18b67c19c2c2b8474e558
z089a742cd21080babbe9f1cf54d7a3c8b7d5b8072533732ab81b7ca9d283c79c3829612bdb8ab8
zd048f5828057d850a55c1e2beff71461f154234a14ac4904b44139b01212d43438d8c9fb125b48
ze616c3eb27a57baf38aeb757cb38f7d31ae128d6d5e0660c5032c27d582b686cd710e9f6dbce9b
zfc0f14d06b51d946fb53a4d73fd922e82e43a1517154f7a2076d347501dd68e21c1ce41c8bfc7d
z7ad23c676302f509aff6545bf93d7975b9b3b56c4ceb28964762556e3baed45915e04ea702d572
zd6aacbdf821ccf66c84629b306d2abd5bd0473fe1a247b723bea03691215c1c3c20929df3f31e9
z3546dcab981994e808a795adaa6c21e4873f8dba53a3fc221d5753187c5159a817daf7e5904c64
z8ec912b891eed1742c094edd6cdfc99b873078f98a59fe43cb1f6b6f8112c25c1e22432b18038e
z0b2eddbc453c7c50f7e4a2567106908deab30087da430e3ea3b3a0d5a768a3e804281354a50ef9
z730a9332ea01b9130df1356ad02fd677a8fc96ea8fb06efd98a2d0dbd1eb235fa69b1b4f150f52
z223ca8070cf8e98ef581b9ae48c4d3c2bccdc30b22bca811170843d173786439965343da0e15b8
zec159c1425c6d1fd40fffd644975889c5f605093da66004eb0b5fc1507dff79ab661db9a7ef2b5
zbc442074f6b4b19379825c21684648562b14c5dfd3e3fd60ade5174656d8f83b74ceca10d03ed5
z335b6f0e8ae6941d48a279fe7004c57dedf0d97f8fc17803e90cc46d06c3c0050247d7fa4a7cb1
z42127e246098ed334f607d6e3dae9e3821cac6698a3c305e221dd8ac26b64d9566ae7f1c4e2fb2
z9b4258324448d3b2244d34f50ff967f073ff950f532841cf52b64289a3446fb77378c1096de07a
ze0a49583563722650cccf67310a5446056c6a88a085b64e547cacf0badc57d18ae0bfd28545041
zd130acc779b2055ab97e0aa5591999e5c96c3e75d4a08caefdc768bdd13155f423983c4fccf516
z6a64da8bfdb83f5d04d5d9e97a311fe1947e2bb95fd86ee759a5cbc21d9699e27b2ba3092199ca
z47507459ab280b192275327a446acea4c994d6519ced55a9f4314647c35c438031e87e24ff2d99
z8a02d6c208ba40eb70172dc7a60795613202aaa18501065f155188e1e54687ed9ed53ee878d525
zb08ed464b9f2d3dea29d18391b2fa824563ed538a1c213281918d7b5af072cc9b6f777274b5fa0
zb32ccbffe5aa0a5a834601e27a4cd0077c1ac0095889b52cc858121158b9d1b3305e4dfd270e66
ze4478bd5cc88f041d191ef12b5c27165d0ace464a51670bd0f61f4ec6ecec906d965b34d636eed
ze1f98d6d504ed1580ebd6bd26e3c78a939aed6228fd616285e7303e93a6f6377d48bd7c51a29e2
z0f7951852e69f95a720ab4c4515aef684b5f75fa7be92c2c79fa64089cec6fa080dd23b3d11532
z4de1e266ab00acfb438c7288bf13739b8259c32005226d226bb5cb2f71733580f56ae04c4ebf76
z5cb45a1511b92785a70d66bb5562025765f087762eb935f32d5199540ef30d207b1b406b2be198
zc26ae409857928d4d67c8ad1da08579b12c22da74ce4bf499c6bc05e3f6ad2b1bf9060b321a8bd
zc2a9db9a88e5a88a721bc01d06a7e916a1e77bca626311905ffbbb5f3e1efb626d35873b18e8d5
zb18e95a5e1db005172918ea9e90ad6c6abb4d7b1459c9d43b304acb6470ac3e5b4b378bee71a1c
z4abba4e1ace68c537342d4c39ff0b545e655b85fab84d98aada89ff8a84a7fca35888238cf038c
z42088234425dd4399bf4feb71f9d6b557468b362fb7df42036750e6474a0f19ada90da780b1f20
zcdfeb87a86f5872606b128c683c849daec6fe40c325c288afd939f972274a3c1dd001f5659e80f
z6b207a2be9791d210cc1ba1c07defcab522474f5e495843620cdd3b6a156d9d36617596e968ebb
zd56d313235e98988d51e4d66b3cff99c1b2052588cb65437eaad14e46413f0447ce17c2e66f123
ze06f4b98eeb8f5475362dafb16e35ddb53cefd7424ed3a9e05c15684ed6cbba88f9b163b975995
z0f1ecc591a2154369f8db6c15e2a9e64809bae418477f319efbb81f5cb20d4e3245564cd37849c
z43a8e4b7e149885d432a8d76930eddfce9a2e5735b20a4b98de6a33fb134972b9cef6d36d4a5d4
z4089f2f3af0e5f1963a95c13503df51783b9ac2b8af71db1cde07f8ac0aab1912326fe67bc6117
zd2296608978c0f3dc02b45f4e44bcf298d6482b264d7c3b2065ef60a240efb6c93c2bfa79a6396
zb26e15774e5a73ff0c7f8276d65c08621633f5a98a42a7531b4dadaeff6d75df5f6b4a02a36a17
z8fef1ed65dca92049d0687b852eb363b63e60cd1f3e1bd36b45ba3c13893a722c862b2a40c82ab
z3bf97e8770ff77c3e3e158de0936d810beb97e3c6b7f7b6db4e89cb49e6af7c162573adb487656
z4c641b02eb4ba97dab99fee2f516f37f61d5a64c272cd4bc815a1d81dff3bab3402e801c9c8813
z3e74f46b88d601c9d3c8b75af377aed9af2be5fa9c6278067cabc59e2ea015ab63e42da9bf7bc3
z082dee1246985f42bfc0733794eb8ade0584d576bbec3420db316b518ac7e02a9ce5a2497a2917
za023df42219bd33f992913764168e1853d805f45358d1ea2ea4d3ff95c23f4c5c2ec7dce0871b6
zc2ab02e58a9f0943d1f6895587e2011c51ab36ca6ce040ff1f75574ed18afd549d2e187299b646
z89469c103cdcd5fce40b3898a3f83b2b3422fd4b5a5484bd890c2b44834b4e47f51fdc15fad045
z9b044d923a2c49d74ccfd4e83cd41b6038705c6e0c40195b55a1cdd907e99ae5c459f1a54fe31e
z277e4b00266004f9031da3453fab863109a9bf77b9f4bcf38afcd24c1196fc7d9ab2168dd72d3a
zd38e776b4136a33d6abc45913754d748b31c1a4d2548aee81381627aa9361110de8d93ff6d8cdb
z6763fda0251f04d021000fd222a483e344ab7fa2db6654932821aebcb329a6adb6608f0623d01c
z091ce59416ddd5373e835e93dc7e38d3ab58cdbf912aacf98a8c24398121aa59adcb278c1df765
zbf89300149734472ccfcd99695dbe0bfbe6b1569454c300c2210efbebdc6b57906c3b9dc74a6ec
z8922eacbb0e1103348a9b3353daf91fc45337be0589c49499a4de22305bb59c702c32439f4577a
z0c431047817e508e701d678d6b542d7b6c8a1f92f0edd8752007f1b807d47dad3e4d43a64c1549
z2287603b5b91fc8bbfa11865245311ba3de2b95552e1aa7b88c9c79d322af2142352028c5a1b06
z5e0738e4485407a1c8a30456cc33056b41dbd574ead6dfe8dd6873ca6146962c56471dacdb3db5
zf4d55c61f8138632f1bd1f610a9eb73a329d3fa41fe8f4190886a0e66e544f4b99113f1f78dc8e
z1bad4bc016d2262acc811690f4f2efdf5a3b2c4232f208eb9286e5a54483f79a987d8c6ff274bb
z3d67009af11e5c98d6f85364c7938d0541ee1c122c72906cd518c9d95fa267a50dd1cddd448fb3
z2a317afb0cd7ca9f300a54d1be2d04ad270e4144b9d2220a2452cd27b453de4727d3054a883fec
zd063efa05e8f6ac9e563d6e9280a8d5813c7a4ef86511643416366a2ac4f51d2673ed6704fd699
z1bae17db1dadfce0bef0ab759fe9e4105736635b888d7ea2e407c66586b2ebeb1154546ebc9dbe
zbd3df2d7fe120cab518360f9052485f30b815d2f7c63be7e57822a31a6b98d82f52998f14f64b6
zde75097fb34a45df9b5b0dcd56563995b994b387239309f23280a07884691e539ff24e3368cbd4
z4ad811f459ead2998bf8d4c2753c313331c52f7c13b2f0c3f014b02190415c332867e200685268
z3e7ee5394c9795ff629cbf2d27795ffb3b28f107cfb2045af4138c1fe64b38c80e6a9569032d49
z533ca1418f4c4994ed44b8ec84dab3b0101ae4f75d164115e0df7e7169f103764810608481234a
z2bcfbd893ee54435a582e360922e1aa43e0ee073b0b8c2a85b2311dd504b23f9bc1706b63da83b
z0f991b93f41c9fc7ad58ed31b19838d44e812268ccb27bcbf6c9136059361b4958609f794770f7
zea5e6d371ca3198fa4e5807036a6030eefab9d52772bbedaaced1dd1c50ae5c8fc98c9401458c1
z333f7808792aff0fa5e62b605b732f2234a13439887feba1164690aabd81e4ba03cbc48d98e475
zb298bbd8d1a7082b0528da8d8e1455dffdc07378040eef66400697cf4fa88e47aa41240676e1b5
z0682cf495ed2757f25540444bbe42ee5bc5aae8b5c6f9bf33cc9b213afe19c050d46207080b16a
zaf7fb525d8ee61e8a8352c782056f8e2225361fcea008a5c0e45ada9994613a7f43a51c4bea3a0
z8421dadebfb44efa71d8d4d548a3f09c0454e018ce86f27f9e3dabc72861be35b8bcb88c5d06e2
z6718bea4d6a1309255d73f7f48392c486fe6c5d987316fd905571fba82877be4ef562ccccae576
z42d846f92d4f64e901811beccf0ff6c3d4cf48f08cfb4c011db3b7771aca8a9cf40b4e8776c904
z93d7ab3c51341270faaab47a7674b9508c17dd186f18d81c0f3469f43b4f17a30ed1687c70816e
z0ae29e9bf59b99d62d0b83fca185caaa972410bc8329c3b778822f145dc9bcabcc21cd28eaacfa
z50f0b808ab7bd8e8c97c299f59baf4ce3c1782d9606ad6b740fa5f258cbda313f762688fc9ff42
z3d8db0fc7867247f043c7e7a095a659933ffdd84e7180d12796768d988c462b3472b8acbfdedaa
z10ea74d54bced26fcbe1008a9debcafefb3d23a9e161f15e84ba956fd6b29399a45fdc5b97e48b
zdc476991ea9ccd00fe604628d63c09b7d4ab12e53be4cc0622e116c04ee63b66067262af789c7b
z35a597edc3c4c747bacc5244adbd0e32ffe13ec6fc39612cdda66e407d3ba5511cba2dd438e24b
z658079de356a5775929d6384ff07253db1d11790faede504ffa39b351d741b810535209b43f928
zadc7358938a85b0735527b54c9ab076a15f75c81705de8045eb567096eadbacef186a15e897a32
z2ef700032234db732deda7afb0d32507cb212ccb1e984f699e538dd118955358e61e814cfe64d4
z78d3e876fca3ffd5064394c303fa6a807628b972ba27c76dc8f4a7859447b94b3345835eb24dca
zca5669d519b9ad234dfc82ad318771379d27bc31b247be6ca44c68fd05103ca9e00604051c7f5f
zf056e276db7492c0fe04a7e0d64c3976d6adbff11f6b67516b43fa7fd7eb5fcc71d8d2a9b90dab
z81c9df3bc44e4ef127a7bcc759ace19c078ea8621d52c3d376f3fbf26907f59e1dfab517522097
z270f6103501458264cdf73019fc41b0b26be75b317c8b1eff48fd36b73431731eb3e73de38d017
ze7cfdd1474d6e6857f745fb6a4903eb6bbb192e6cad32ee07c0cf5f29577be1d6e04feae53c1bf
z514292a4da3c912521f74ae495a765705453d6473097cda56e05e427412fcaca15fa1a933e879d
z7e8288ea5ca7cfca9fa07f5f4d1c3e41dd3d7bcd8a0997361e9fad681cd3d9f25dba4dec4bec9d
zf642232ce2980b7a81c523791d94a28c2c2d16803287215d5f36b563916db607570301f966bd52
z128f57c7e6ba0fd58ac21b025447982c25f89fc77a1ebf2dbee1329da28448f93a624de1c0d260
z54fdc2da84683ee758f02bd9d7ff96b492bcb99c0e2b048b54a21a72e96f025711297b823edbd1
z458ad320541d0d8a82952f8b3097de0e88825575928975692523543d6916b569ac54f93afba270
zf97014fe60db76edc3adeddec4dea14b7e9e21c6d89a48c9b49abf570c9ed8e397d80289cf6a3b
zd9e14b2316042c9308a1fb25378b09401567b9f0debbeff09bb2e0bcb48594c8270993ee8ccb9d
z8973b1ef572bcb1d31ebe6c8671ac5e4694a58ea6b52fc8c734a2a8b6e4100306bb21b38d6e605
z09ee58053c755cca7993458aa8db8061cc3f47cc042e77ee4fbf610905d5bde8c034198baea8ed
z0ca69b37d65ea560209b660493a95984d0896d939d11e0cce8c001acbc7259ebd9effe9e74cf91
z5eae1d4f5dd6ce6a80b1c07a0cc18f948c0e084d3925b99194a9f9f0516cbcd905e3b6ed938ddb
z1c6d8e9cfc018987e5dbbed60925cfb4505edcec731d823e5c78349072cb327798be28d88e478d
zc7621d5150fe55fca64d3583db56d83215bfd29e3fe390a811a9a1546db3e27466161c0db9a5ec
z32cb66fae05d4bf8be7c4b8bf0a51bf0b3c0b74090f5d59145aef0088113b4b133113dcc51ac65
z9894cb641fbd1acfe67b487d20597b052c95375029f93d7e223602e47c7a4a5ef506778decfc5c
z2b8acef0e5a2ee12ae1116fc88503a6fbe0ae0561f5ab62ac65293cfc17f30653f1f071e286009
za4e0c2b43cdf81e8d392ed2716d47fda8d4edd5d6337639ed2988e8fc5ca414ee92f0365cf9bb2
zb6e25ef2120c2970539edd2870e675064893da9adc5fb47f34ab2305980df7952580521e790bba
z99789412a45953f83cdfbea44a29d6e7b039ba9c3ce9711e30ea315794e92542128c6305d9e7de
z5d5d6923a586e1c075ca342af8ce764956545254afd86adb60c6133deaa1d046524e9c6051239a
z341b827b620b32d86ffd3ed0cf3a282a8a11cdd693edd097d888a01a0b2604efa1e4119e761f51
z1e5013573faca9452e492eec306d1b7a7248ece53b2569bbe2e534a19eeb5606a8ddb80545fad9
z6b895922bff672e46e3fad7461899b8f67ee061cfdf8ac35871d6468af833579f9dbec320e2ab1
zcb196e9da014a3c07ead934ad1f16cc39f0bfd040d91a2f893da12b7d7e8402178672786a8261a
ze15d2a6d9377300e136d2627641aa8346f22f4548dbb4ee6f03ccdf94bcf80dca6a8f7d6df8cc4
z32fa22d8b09ae0c6db37ae8bdd1401a3c78df5dd512ccba1e0bd36d32295de7d7b70cba53553c0
zc0932dd4db1e88a2f56380183a26fb23483b38ea8beae4317bdd509b1afdd318064c8e2592eaa3
z7293bc6f2c05df91d91f22bd5f2830ca3ef8fcc3cb7b94c34885521350e19b8f284f4d94d6dc07
z92a08f70d6ed24ef4c1dd0c079b198f485e5f9864dbdf63584aafddfe2aa91e7696963945e7579
z097a0ddd7b0d5b76164572b68b42f06c9b52176daf3b720d28e487b834f563f74857fbe16ec183
z0bcc7f441879964a589cf477ac7fc9ab0bc457002cc747df12fc08e94de50b0fc126c774167907
z3721c8304006e3695c5efe6391d40b0d5fe747fd8fc1ce23e5939d4eba108db9cd6cadf51f80fc
zc300b2f0e6b4bf9a6388b5f8496b05fe6c1e7f7dcfd61e883de89e5a518a4760e31545d8a7dcb5
z860a53793b11397420282a7695e014cbcd8d35b82320f45f4ca221247e1a399012f8953f5d3db7
z124327de9e8af19accc5c72c3166d40af092c369024acb8bae45bf23d26bc13bea079f751773d4
ze8acbf6f30d5a2a0390d1dba5908c6e01eca8f0df67743ba80a2bd49853462750e5fad920ce19d
zaa2ec21c1f9673668dfc340f92372a504cb9a1346d60305b421fdf1c3644c17977619460bdd88c
zc331762e2319efd7d5f47036a4c61739110001c9cf99595437f552f2628e22203d216951291bf2
z87caa81ea6a778b22853751df0991a3a19aef475de7b8ec83c958fc9eda22275df43e2daa7c4b7
z2259a77b77ecc8dad1db4d33433b0a12e5fb26da6b0098049688c7abca9c9aecad45537212b728
zef8375c46d632ba668e1a4a45f4d1a60694a7faf99fa21cdf2e967dc8112ba566c7ef3feb04bd3
z325bf6a513ef0633a6bbeb1ea25a20a4ef44728d191ee4ecff4fd81109f14a3725db57c8f59a07
z4010295755aa24477a8049b093ae2b8ed68ffee3d73d4eae5884d17a1d86147e2ead9cb092084b
z92905fedeb77244f7eb649b3d78d76e9a02f38b0e1147594ed12ca91b548e1dfcaefae254684f7
zdf2012089bd30e395b5746d0ae57e740ccb2ca3d41bb8f177e0fc20e43d6bc9ed78468d94911aa
zab7e57f631be25c17e0f36cde853f59d1f4737680d5439b8ccda5bf006dff15bce50bdedaebd3a
z0458b9409113642fed57f91730d180b9f346d9a476b42e484482529e31d119808f7b0bed705260
z7f4d255cb50352e26689c88c04b9a14bc43ef838c7f6bb3b72a262f859daa7a4fa2a36fa7f1782
z477848a855e0f941f7067d1d377457ff2c02a6a4f55389261a3cf1cc08b4901b3a0dba69cc100c
z231a5562711b848df13ef06ca1e3b65e6b9a9d1cb647e2182e18a293367ade8f538e06323aa8c4
z7e3d73f9e876dab9f2c5e9a32b38dd4ef0e0f7f58c834c02eede5060379620b56ce6f1dce8c0a6
zacc1ab200b8a9617f0b0ceccd579b464b6c50abebd37e68807d1d63370484e4c841950331e3667
zad7287f193878aba43407b2fe2af928b3897ed2cc8ae5dbc76bab039d33134f635fe9fca7b0d70
z0485f480893feb02295458bea7f2854c96c0e0a43fce375275ede9db6b8deffce83f6acfdd94ab
z45d809c0147ae0fb1bb2b9730856d655ea8ab1c3e4d8bc89e16af3d1e6fb6d6a17feaa3c614c8d
zb1f7a9bbf8b2477fc8fe3eff445093e24968b14c7f5b5df7a290fcea90f34409e7d4d87174d40c
zd4cd6aa94ac9311c889c2bb3159e6838837c01ba57d9b8c76d257c37f864a6ca7c0c7eddea3afb
z339ee82fb26993852ce4590df4cb20ad6d3b1e11cbd8b51eee6dd6da441e1515e0c4ddc5468a17
zf502014b7b27330a6489e4c5336809e98f09f4b28669f136cb07bf026fcd9cdd87505679d2c168
zf46a2e1858307e7557f17d8a7e9edddc31c7ea2de4a9e055e19a700c7b24e7277a189bb693df32
zf422d84407c34d8de5476b4d4a375bc4df3938553afff91976aae88a5a684709038952fd2cb46e
zef4a0d5c3983f4e3402b4437360db916c588b6c58b4b64c5fc60be020cace8adb340de62725543
z08d7166d0d32869591680d6c1da886a9b9d0c9cfddf059637609ca12febf268e01c1fbbf6c1ec4
z8887cb731f0677f3e09e260f684c92c1cbd02130817e22ee6c8edd3d434b16fe6dcda26a598374
zead718fcb95ab7032bb4d03ad21832406348cea848e5ea2e87cd304e81abfa537659f88ef63c61
z03c032a14ecf23969d83b259dc8f2a33ddd3949adc0236c1816e0cd6a08da86757ebcb0707daa3
zf1e1d402fce92de52236c31ff81913b0f49929176549de56683aaa0033a2592fdc73f702f33278
zcdef6748d35e9a0c168e09d86f347c3c4610399b2f25503a0b9b4fc6f1e93ccd89451d1dde8a43
zb65ca494aafbea0733d130557d7acdba2137afb8d10050635aa0af8faa3c3b59de2d770df99b84
z25d7b28fd054e7e8642f28ef3b8656de7bc2705314bf9f2ede26d287b3296d232949e202b684ef
zee4c0d8e5a4b7d6a78fd975ca107d80876f61a95406dcb5120ed8164e0873c8a1c09f58ed044c6
za97f78cf497e6f2a3c529c6185aacdf99580c6990f75cc59daffe065c023fd19e67ba36db6c576
z87abaa049921b8b101e83a2fe4172b3b497b4a70645f8a5e80295498edbc3d34b7dcc0e3f2d240
ze09803a5e294585081effc6667bf1a86092e1b21575e53ca92d97a127324eb9e9d32a2848c0a20
z76e2a019ea6f4fe24a23ca3de6646b2cd65eadbeb8ddd5941f041ed57e4f5d8207379a30fa7bb7
z7f89619d5f1dc696e42fd5a5dc0c44e9eb17f77a955db1066f1652096c899e2ce73ed9ec8520f0
zf7186da1c5b2e4119002c6c934fbe386a11715d22db1e78849b5c1f48a90f3de3426f5f2804e61
zad98d8304e17490a1f71c549524c5a0c6112fea5aa50ffe22d3ffe29f8aa71d4602c33c889d7a1
z5b604e6875284fab69178f422244c89ce4c2ecae0515ba296399f6412a4f258fb2ab4b47c2c4a9
z8f03d76b09a78565a65e491d8d96146882b0ade378e4a9a4853f9b16585fdc334bde7189294e48
z1c320a029aea343d4f76fa2996f9001517e95f52749fa91051b66bb81176316803fad93bcb7234
z4445c41456e29edf0b85e17613b012bb813d6a5e61f78b04440ce713d32a916a71d08bd6021f98
z67cfc0a7c4ec5f67ca2a39c3c7ccadf814c3099737aa0a31b2c3f98ef1c489fb7f112aac94d13a
z93dad3e294621cde8cadeea32a9cfebbe45a6b8193921ac5d5fb8c4ed3d001c147282fba29497d
z815681ba051000ebfe9454504ffbe2a03473f7759a21d8b0d5a813b6f8a473c10d65badd1659de
ze4207a95ed36672bdada52986af5b43a903960c8950dd5aaec41999ff0f279d0b2d7d90b2ab5ab
z2efb80f2e0f05f99c9f147d855dea4ccb471f7ce2f09d4232e4ddeb5e6ed2c3e0868c5ec8dff1c
ze547136a92be382b9bd9aa7af577a7a9276e6fb016dafe81ea15a64197a9ed6cfee54521cd0d43
za0add9c8777f10e8ff22b530a4e2aafff6f16d6f27907800218aeacbdfad7b884184792802a6d3
zc142f816a95c12908421f72f1ee9fb7098115253c5dab17143173903d073eec5ed1999c929b57d
z941cc0b405fa2170c9d40fd551410d582493ccdc38860a04e254eb0374713a0edaf94b0ebf85da
z09a4ae84220b38af18d58afa0f4c1dcda662b770165c37427930e5f28c2db4031feeb67f5ee755
zf14a35cf2142c03f044549c5a8b9bb4be4db322f4e28e1b81e1fe8addbae9e12db3bb381e0291e
z6ba54331014ff5ddc45787e9f7077ad125cbc0d54e25c6008c935614c9067221f1c276a181b194
z6acb033b4709217d9a44b8d87e61424f423a8849d74dd8d0ed4a6a3dc8c751cf5d03486a0369ae
ze6c40e885e13bf574f8f0570c6b056acd0ee998d5ee9e1e17df3e1e2a24baceef7abc629a135ae
z7ffa49095a47fc8677721c9b78007767b8653ed40b3514cc67138e77bcbbbb10585670abcbcb5a
z18d1a274b9d7bd6ad07f1cf160ce26679e2e96e9a7a0411b273407099539fe2438495ca7e80aa8
ze0ac7b70949fda80a750e504a31c67242e66d0a30784eb5d5fb5f4e3dda56f5ffef4f6df52d89d
z385b4281cb5977ac99fc320fcab9c3e442623983a398f45fc900c2835beb836be2018a3c13b42d
z0faba69b2cfd6c4337c708628f91ab09344651e7663863cea3fe2f8d25f473770e366723638137
z8011e3ff523ec583093e737bfc39f599af097e87c6142b0a0041d860f648c9e9ad63599de3070e
zb504cb1e1ab921a1a85d8cf6fff214f9486f22a0e0204d592376cc822cdb6f6ef1d7c2cca50949
zbccb2bd4656672d5646affb7a89ab7a39421a013fb6efb6bc78dd0d6fcdc8413590c6423215804
z33fb2fc9bc731c81f4415194664accdbf6f88e9d6b7dd8e3e448c654a5abf336de45ec90bdffe1
z8765a58e334aeeda2ffae07e3de3aee0a612b80bc5210d6daaa682e1fe3d1290bc457464f99a84
z6f400dea2b9666a7fc288f42122d55670755cb89a7650a9fb541d444a28f5565a0d988fa52ae1d
z03a7be76d74b15df2065cc768f78237a9c7a3aac92a5b2d081a90391438936e7701392644f20e7
zda08fdfddb1f81c7d2397fff8a87ab4eb65b8ef174bcecfe34be3f2f708d41432296f30d9c63d5
z4351382560b2ab332faf6abaeba8d9eadc0f7411533f983a763d667571cb86ed16a75f80a0d17d
z4ea574bff146b3e9c974622f1d8bf05735f54bfd992c55071e24426d23693108d69b84a3c46177
zd47e8b48c782bf26cefcfb3b3cd275193d93281dffdc1f225e50315a82a60b6d02854559c57bec
z6a41c377a6779b4275be76b324289664672c2a0c3ae998f5ac2b6db7c058876ecd49be9c4cb7da
z5a50f701f860e4a3a82a9cd33e9a91cddf0786d8a66126b160dd91c1b0e7c981021b200d556bf7
zc005cdc0284b3f4518db42e7e5229bc7e165dd5f7e8e38108e6a3ea4042165f391d9a9efc54605
z6e1691512c15c937da5d5ec512efb12b91d3d4ba838e4ffff1b1a1857c2aef4b37f5a65bf34f06
zef11dbbd91627516fd301ddcce9bf86a78f3887b5fbf49c8bd045c12c8c49a42f739bd81e6c7e4
z2bf1a43a5e231499af87c0562a97857adc7ecab79408645f17d89f81de8e834b146d3c0258d3d5
z83d7b81c75d27b72ea76fab6fe19d0c193f3477f87b863855f2eff954b9a772c35d119fdcf6f77
za9dae712fd27ea4780dd5182935e323bce20208c27670bbb9f6b4c701c4b4a325d6ef781d783be
z99f58d293f4ab2b380e40e659c3a5baaee9286f64a87907feb6a00bec3b6ea823dd2e7bcd9069a
z409cde283dbbb7b2a33a4d69afd77d3f154668596e3047e79e4db5e3d37d22f5de9225f3c3a87b
ze719ddb7a76e5280446afbe08b21a889f27b99999552ce66b62c3055fb29a30fb64a794b9bcdc3
z2c5967d1e59044601098e1fa1658c5fbdbb71f57076074f2841e9f543944845bac80664c85b160
z57c11e0fbfeba7bb63966c94a74668212d02bb74bc41b6288ea92c409a9b4ba67aa5b694c5988f
zd32fa5b5c48beb7a791d580419d46312b77ccbaf159b53b7c5fd8732da578a99b795a40d50f18e
zc3530c410c8b5f3887208549fbb7c5537bfe43d468b3115539feefbf9c224a8f1d84d5947ddfb3
ze51f355ec746d013e4b7f00532ceaac9547ea56dd8b1881f420577154bba426430dc0eb848fa2a
z83d950d788ba83c611e214ee687132ccfb1bdd04382e1cbc19183917827f3235785b703ca1bb90
z0995a3c5359ccc1ca58d818123f6dc58f1fdd1c361cb45e4a6180dd105d820b5ad35271921427a
zf9ecb94b90aec74dd200bc74956c9226e89b087424a246b478aea9da613b27f5bd1b26f3f358e4
zebd7b3efa240e74e1e63b5013338c04f3841da253870c3b9fefb97f6984f8255d8dd5364dc95fc
zfabd7cd5c97fedcacb4e6cf59c7deb153ea4230c2f4000e84c63bfa61bac68374b1cfcaad5e8e3
zb05a07867972f569a1235539a36fec2ae7c0d4f61f37ae5bf807025bcaba33d785fa5f18789820
z0138c7a2a9aa870806425e23d66c099ebbf831da49f5b0c785595ce16caf9015d465d35d790830
zd7e7942e3e0838243d74a0b9412d9bac85201392c291398ff975ec594951df0c95b67979ddb875
zfbd6dace74d9def2873e705126c4941c01851c0fa7fea6d5c4b1e6d5786a4483800227cc3e90bc
z3dd3b864ece7bdbc0479108d2920e83cf34b6b98098cde7371ac868341a308dd742251e6e10a5a
z8422be38ad66bb8d3efff8078294927a89ebb8510b3df01d2e8df4221903b8d40e201e5d6ac962
z08f96869d39fa36464f5a85a97843b396fe3ff718cfafdf1ff708984857c7126ab3ebd85091bf2
zc6fe380d928616611dd6ca395211a1be0eebca4cc6b694d9afa3455d8fc400fb55b8ee6969ad76
z4eed242331c67e14420c03eacc8324c3741e80641f6a857cc015d8796672d9022b76b41bb35d0a
z2f3821742db433ba41418743ea84ab1773fa5d4f2fa5706e6d6e6d3e64c08ba25b556765f91cd2
zca8c8f718fb3fa7764d3ee64e4281c8bf07163f9a0e7b6ecc4eeb7792dfda8c566392226fde403
z74a3be8c2d031fd801f2ea786fb4e162ba4d453ba7d959b733e218f17eb12a086f0e800055a8ba
z180ea1320a208b3f8b8237c88583d637804560c670d1e46b26ea86f03e5f41d6fe7c97fbbe8565
zb2f797f51f6b6263fd429c81327e0f6a7574674c171bf3aefd4c3b0a038cd2614607d27df4201c
z86de5567949d2889dcdee9c409d83144caaba285d6782af4498ed21646f4ae2871d5a830843de6
z483842d0829ab8de44e72237c7b8a3a86c44764020d43a7e2a88ea7eba24e0ccab1085983e2a8e
ze344a78840e6cd08c5c016fed8d42990475610e6aaf69481d05453f2450a51d8061afe036f76bb
z4806fceb0394eb323593e8d5688a4f99ce10a2835cdf430b96e921fa07045ef858c64029eaec8a
z309a84a49faac564dbd1c9cda9e2c8caa589f8204e74360dff5826b986d0c9647282f7aaa470e7
zdacc4937986803c63a4db6b3fce178bf1f34e6b78f16da2af6f2d6a53bf34aa4a6f3582f8d77bb
zd1288dc0ad7ea831735d3ff4bb33e49bc25859c5cac6656ce6494d138ee02ea80735f64af76431
z16bf30895fbd2dffd382d2e08190f766f3a6dafcdebea3e24f4eb80ef37ce72852f09b14f87f8a
z4e002925ce0f3e3fa99045365298a61c6cb51b46d6a69862806a00978703a1961afabb01790d65
za426c53b0824bb09478cf5965c438b7077c747182fa50418d0bd73bfa4c5f34c91c5372e81f432
z1bf4d223c36957c6a764128eb94ebf0832d825f2adb2bc96ec4ecc6875c4e84572a92b351c3608
z076a5c4b9805ef78b46aa6680861fb26958bd2d97426d99f437a9c30d5a7f8d9768c908f42720a
z61dabb52023f078fd4233de92a9f781a070a07f0a0fd3cf99d436abecbf548ff790a37ea3c3a06
zb4a5eaef8bb0997b48cbc5ba403bc7d28aec1e4e0235f1747a3328e1f326c851b1c4e281122b80
z7ee7f604e3fb4063ded87d24811e38de16a0a8011f577cc66416899889104c414e4769f053fe1e
z622528055b6ecb64bc2e196682b279472cc072e3e7a5f271c177b0e0b99e84fd791a7cf8ad4482
z07f009bbd3215616e68ea8dec275c6220f8ef8d2330ac822a3ccd36b81c96838dc7e3f7f027fee
z5f82bcf7075ef9626abb399df9c60c3d5c5dd734ac388edd3bd78de1f442febe85f6d2b78bc734
z6b4981ef07263853e5c0a5ee534f5cd31279dfcf89ddf2ffbff3fecaf10594781af5ab43d43df7
z38bc1a52c8fd1ccc47f7aaba8d8f44cf559ef7969bae0b698e72d9f91353041e8804d5edbfb1a2
z694daf8645db89e5cda4dcaacec4eece8ff4077edfa69322572b4cee6b6218fa33473f6aa61003
z1aef3adca6799244cd7c816dd8562009ee43f38cd78192ea09d0125fe2d6261a692e06da2fa6d4
zf4a8017275511e6262cfb97c6ff50dd72d26dfa93103c163c4c5866ad2c92bbd703e9fadbaa1ce
z35fbd07167e19e94c26a0bea6dd72a502d396385612668835ef361a1327e544f939d594a090c2e
z23de300d1cae688a30d3783d5be746eb3db43ba587f99db70072dcf5fce0fb06749b94ca78184f
z0d6cad4d99f922b4c59cc42220b9968d8f9c8274ca7c348d84ae4f82ed374437148264031fe2e9
z64ed5754629e472665a5ae1d0e07a10d488732dfcf4ae501285187b314dee02b106a14d5ade68c
z60c0e8db1a43e2cb04cf66f831a88a0563aab03835dd2bd65ff56e346c0cc433f737aff3b47929
z2aee81c9fe2daf299379d584b3e5864129117b3bd99c151ff9c16190c267e2f5f4ba6a783b6be0
z22e36e7dbc9a705a2d08673282ff7161b02343d25a124b82ee67218c91ad21cfa6e9899400b72d
zef7fd01cbaefdedb117b41743d0c549e48cf2db3e46748214cc19b4a92a6becba97e9b79de4ad9
ze8e504d796b27f6a0a8148f4dc78090e2824cdf44262d26d9aad28cebbb87876e45e6e8c53e6eb
z208c96009350c42bdc21bfa22ac7ad075e576e6de43d02a779ae8f943dba48659773274731fb66
zd2838c8896cae1611765bd952fbea33e94fb1adaf7f6efb3844919ac1db98d8f3889bc66a7aca2
z8f5a95f067d9b8c7a3c4463d1bab450c45a0765ef4551f07036ce63111921cfcbb24256b027b0f
z86bd8daf133714cf8a36bbb388c1b58c80138088acd0c55e368a9bcf3dbe784e3bd13b9663e523
z234cf9f85da0cdba948a6961710e5eeaa8b490c5897d7c68d2b10764b575c6f75eb2757e8563f0
z32e569318299c164b7ff03f050d2a42ccdec5aff401c75b959908a3e631d171ffaaa06555952f6
z31e9f0093c92148264c8d5f7d360eb5daf43c8a40c879573ca530c5bd33a90dc74c0f310c5ee00
zd66b5648494029bd0954bb8b20d0cc7d1af1321b9002754890d331186e8035e46d4ecf611cb9b7
z4c4aa7b7532f59539d3e9300eea98fc73d1d73a778f60ac2527cb13c13c5fef5082ec315f7bd12
z04f77941f13da532d18a2d460cc25e9314eae7510ba2532839087052d1efa863f754e3bfa7b530
za9a127e5e9dee32264e28e44c419f6934781e8d9975c308a8bd7d4cd5a4ffa1071b4e6fe7039db
z27579ce9b2eb7d03b6642217e36e61b02bd88f024b94af6f914ba1ef973edf920e7a625df6009d
z395460bda5184bbefb826351bda01278a21dd7001e1a4807cbceefb0360f3f2cb6968b2c92f60b
z2bfff67bc1b8cbfbe8275fc159626ccab906d132ccdd424339da3f6666fa889b8549214a0c915c
z4c2a9f31177ceba1de96c074b797af2f15d301ed6f1b3028e8c7caa0e44cc7234562d64626197d
z5483feb4d077d5d0155db9785664d2a39d027e17f4cd1b5a953077cf5e54c5fd10c3e3995ab11e
z4299e999b19f78fa2e2a8edf4ae3d695d0dc80d415a9e5f3a236c58f451f9f1a22d0951fb9c749
zbbb648de9d045d32615fca86e30ac7d9709978a311adadbd80c7711482ff47818ddca20bf6278f
z3477863537e675f69f6683296860e4c18fd8ecbb3cce8eff0e949ebe1ad33ce2a3bb73ccfc0726
zc5d149ba093f18684504f4338bd0bf0e0044c9213080ea64e430cd828b41218aef4730873f47dd
ze28e5274c0a7f10ab27ed1d99c3d1e7b44bc18020eb21924c31273dc5df085747c64a6393a081a
z82d800f447b8373cb4cc8382a6eddeb903ed0a9ec3a3eb9ac3543694acae7f2d59dcc801c2d0f7
z86b5ffb96b53c6d985bd2195f734c9a69db8764b2dbb4e6dd23f0652a38c3cea089df610aaa00a
z26d034ab33909d2244a197f9204d26e5988a1d645ee6970445151d34944befab59380aeb09ce37
z21cadafb979f1cc9b860487d7e7658e5d846840acdf82940c0986a23ae952ff914c282c957e977
z38cfeb69ba9171b3cf810a125c41d478feefa42ed159b4121bb3ce706f5796852085870295a056
z0a79a9bfd26184ba8030ec2db6487fea9c1909c100c929acf14f22501d72a1893ace17755c9a59
z138f48da51178e0f28b096e7e22e5a6d5c8d7759fe10e1058f1abc56e07a159feb401300e0a4de
zb92474589ff9519ebe4b6961f42284353e03a769b29cc410e5e422786e2145e3fb91da38551c10
zd9fa7d3d7a46a0b86b2eafaa3a5566d1d83c12ee6e3a5d2b932ed65bda3748078cfe94732bf821
z64aef513f2dcbbf13e9bbaaba3a6c47581b480dfa59975a6293315f8d449c14d4529c0c4759221
z5e5234b80166fe29ad3aedda6c3fc06eb0ef29ed24efb2e69c4a04147f381c10c07eb4dcaf3ab0
z3d3f5d29bf6aa500b36696ba8d05afe99438f3bfa66a9851351c2125369f3c96339f6ade1f545c
z21f94926d39797f27beb1b465db38484d5c063027b41d39ca6d034f9493dec9ef47feffd4a69c5
zfb0e69326bbfe1b3d283a31fd617a0441014d4c450915ca88aab9e3ffec4428fe48f707097472f
zd6b2bd06f5796eabe48d43213a578340eac5d126f8f44fdab4cca6ed849b1bb74f7d44719015d7
z8d132b91b2e4e5fe837ac53dac43cc38a057ba453dfc8864c32e0e7685760e52be8a790b436894
z6ed5c6b2869c11f315b08c5f9539ae9f06864a671cabaa8504f37a602ce1fb835275883d1c7770
z0f62d4ff5bda427a3529ac628c23f01b679541e01708fbaacf3c83e52a4473d93d6bd92ebaf0f8
zb0f93764f3b8ad57e46ca053f64c5b2ea14930b695161f9eef41277d1062659b3cd803448236b6
z2307d8fb13fd4ede6a29e23447ce2fc7deb4e1a9bd3e6aa4e815a86af6beeb264a324a793836aa
z28a48bf767b5f0df20441a60f27e5063499ab7ec6f3c5b41a045c068b03105df30a5d9561d4d45
z119e0a742e8a203c0403128f189358a2610d8d3a4e82192ed9db07bc5dc9546408e12f11c0af86
z6b7d48ed4197535f3b55b60b62ff985368147ea1d027692b22391c6e15ef53a5a51c1c97a96cee
zf5f476c4310e09a5e3bcc40e8cecb5802ee25e68e65aa24a3577d43e3671de16065e8dea9b1821
z0e565af2c50eb923e2b5a3d13085a9f71e1eb0660735331b5f7e72c9c32d0700c85371fa814559
z0212e177677ced550ef972a1d554618fcc44c66ebbe71415a7f54b4701024626406797ef4e8882
z7b3a1a57ae222917d50f7b58b7fc1787da8faa23b1027b011781a19cf1bed281e5d864fd256605
z54772aa4b6ab428a9735a40701d4fb4b2ac9cbced8567a75b2ba214ccb2a57c4be33b400733133
zad5b59b4a68945afd33e6eee2aea67df4b907c32a6b094295714d51bbc32d7b0e98993a7a99a5b
z0159d3b74c8e93f3be9cd7567ca4e077766dcc831764619e3e3a9778cae82564561cb68e6df4d9
z956518d4815783b570476b01d6df84d9bc7133cad99faad6b0f791340c2a267d3c003e2b4b36ad
z998103136ac68f0a7ef15ded8e3186e3f51c3cb388e7d59369f9a3ea676d4905143aa51e5a477f
zd0ff1929c7244343a105455036ebf4f311f8e72427ac62c565c0282327e784bfb644bc24ae0334
z2cece35104b34c042b401a9d22adbad997d6175c2f729eaf5d1380d0ed8de0f8771d02672f0d2c
z62c1d882bc51fdd71ba511921e03d1a917a40f200a87fee4977aff63767240be104ded67aa78fd
zf0547d64d5ccb227624bbf5475f09159230c5a8c73aaf720a587d940501dc54eb1fd611b647374
z2962f3b7121a97b942a39dbcc0557497a77414cdb54a39a70b39a5d67f28776774935818a5b6a0
z8f799e95453a6fa537a477f6cd0d9310abd90ef446232eca4262718d6f530cd3466b70a930c946
z240ab4aeb8af0c6dbd1d9d4e17662c8deaa3823d5b270101ff438901f82abcb925125eec766715
z13496a5ba3df563c7ac0a83612c55b6e8dfd9925fe1e5fba85d81370cf220f6c1c48fc531b7520
z4ad1531a4113a9f362ac88ebb60a451d546c2390d98040ea3556c422b665270a1775323c5b99c0
zc9934bdf9e0320d6fd1145fd469e691486c9f2ac72f96cb978f8c44069b4f4bb20f4fde9aa1326
zaf378676b1f3019d034e659fa4f1ce28bff4e5417fa56e47b989a3c5f7db0f86c4cd7246488e7b
za6383254168faf542b1b800629c9415fe6d62af10c3094ba5e0c4b2a2a271ef6e0511adabd711c
z43aba4c58e2f26b7cc52d8ce278aaa5567350eb7c3b8b0cefe1631f53d8885cf4476ac2953d176
zb1000ed805e8f314aba86a600deb30cb6861226a1f92fa401e8f53d6588edb7de57dddcedf941b
z5947b811d578c446a160ad3bb66540622b5c5a7918fe3513081fe7e5142629dba52501040de21f
zfc0c0a9ff55f220f0f81cf3b830e1d618e7a2200fbc8a6bf456cf1e2752bc8b60ee2b80626f2c0
zd3d62bf270a5384e0ef47904bad68ba9ec88d5d0ab1b082d77dbe534de8d4ddc6ad88163e9d82c
z7b2c9c9de51ef8d08f913c1cc57b82a57523de3d6a68492d76f51e98574af599f4486be8cb442b
zc107d4e62d71f5b0ff5348a2ba433ee01d1cfb128fc09f11c49cb7d3476f947d4c8b96e5d009f4
z9b66fc4e6c96d7ff9f8cdb6a40d0aac7b2ae71573faa555910b3600265834ffb6b0220432dc241
zff11fd1c281c16b6043bc614e7c62625eb353a3a30c453c983bbecb9821881e15283dc03ca5407
z0d80533118e0a39b5968c06c41f185db03dc39d84549aed05d1509a07fd4fa093616437274b9bd
z6f0da829845886f9b2cae6374f60b63acd1f9ae902d00b7e26114a0369bda0f1a42f13dc66f196
za44259bcb646d4931667da07f56ad5f339ebe37cb15ddff11628f620177606ce6362ae34214ddb
z15cf68b13cefbb7a2cb57fc02ab8e002f5708d0961978a3db78ba5c7f3a914523442bfe9bddec2
z5247c644f9a90ede6f15af317968bb122a02bd4f1d927d35fad14d19192cf05a27ad41e54c82b1
z0ed86ed0b25a53dff0c8106ee776d7a0ceab32b1317af8b5e0707dc8acc74a0a6816f9b049e47e
z8e2be96fcb4e62dcec95425e068f0c1db922899e0fd968b41500e44d408bdc130a9e8259c47a2c
z4b840ce8292bd70e1c23fd5c08f7cc869ba96682c3fb463d151a746ee831d0fae8d5d4e8158d5f
zd5d58177403609711fcad5c410b1c7bf21fe79dffff1bc13e1431a444e5db953ad82ab99f458b1
z6ed65c477dde808104cdfc6c10d1be693dadde7d8dd078169f82f5e1814c9fb471ac0f55b98e66
z5ff08bc4630a37be8a93760a5bc0cee6594c9ef44dd48ea6a1737c25686d5cc056280e2e2ddd92
zfd74ed2b45bee8627b6f819acc0357485d1848ac7e83a5f1e70fba3e33e6f9d3c5a12376f0f07e
z9f7fcbaee077f21e6f79c06697dcce463cd2d643094e326ef3935f2c23010333b33ca62ece163f
z24a7cd8b0f1d485c5d5389bc2c574b87e8b76f2ef7d04e7149416fa3bea7c5f6777f0475216b91
z51acae1bc6b860e866db38c6716a0ef446045ca855fbc60a2c0069de7e2e76d150988ea9a83216
z699aaee2d730f165249741488d2912aae2f65a10673e87d7ff79965c87e71054e0c081fde5cc06
z3ec012367270133000e5ad97978feb56522caf618f648e865025e7a050cbdf3d3e7b62325159df
z60847daf00ed68fb3736af4b7c7d184bfaf42675b0a5662c7b4698bdcb071f65f2e065cd8ba3e9
zd24c2039fc67ff741e9acf4af85a6223a83429fc77497bc21979213b3658dc1f40479d8aeca535
z68ad70b62aee2015c15b15771054fb4342ea5a4915c8be8b54bce330ebe378180009ce5912213b
z08fe17b36ed8309c93888f1c16837a052603bf389294a5d41564e7ed86d23738b7a601b6f7ef42
ze1d0f2ae0cc4fa032ada4d267adaec5439cfda6e69b0dc056ed42482f1a70a12f98ae7f421f858
ze02f93f3b2752a954051bcec9fbfd9de58963494b6bd960a29700660923c5ea0e60f51f6ce3f3e
z675acce2a733ae69c553dc2c5bdd8a1f0887b05899bcda5c6d8191cfb66252112e9376ead88526
z182e0bf98a80a1beca5b4e9057c88a19ee21a9354d922453492d6a581f39d040f9287becaa47b9
z0c7424daabc81f2c67fa91f410a1c4282a999bacb22111c004a318ee3232c186cef3f6ee66faab
z14193403f8d927886a378ee1210532f5c3cc540ded9a423a2bdf6c41253f9e2ec741ca6376eb5b
zf6abc5fcaf2d307cb8c68913e0d8c10015fc2fa9e5809990cf83e8b8801aa029db774ced08a1d1
z5b04dacc7647c85541f6caac2309480deed2fb9629f7dc7634bb8b2a57099b485acfa344bbf1dd
z2b0c6e9e94c095ca925a7ed3a4e4a7830d6c10a3f171b067612707a5638ed332797644933fa343
z4e099c5304d3973f34fc5437ddf0832d9e3fb3641a6252e31e71479ac2f13e60c32c3c2623f8b4
z5d7043674761bdb394bdcdc1e677fc03ee4e02f06984b8e1ff0544d5a849dd26b2527a83d912a8
z9f3cb522782572243ec83e7d60ea3e83e3dc3e20996c74487884c7055794875dd959183fbff60f
z183d182dc923e6d2b56d46dd6fd8f6a0a8131935542266182863cf2b9dcb25089eb6e828702d0e
z60c34461b82a6614d8084b678e529b1842c38fc64f16794d94531407d3ea105641089bcc5f28b4
z3222854a06b05148580c77779921bc45e5e32c716456d445d2d3df0cbab7cd7f087a71376c404e
z5388d2cd706c201ca38661a7c6861c1591fa810bbc1a9818736e1dcede046aee90a8e8c3236a0e
z438a8d744cbe76d42fdf14f9987bce426fa2c61fbcb19d1301ca4eb9a904ac82542fba21871509
z5aecdb7c31bfd068f2a1933319dfe9129cdc5995458a198cb34f589cb8b94f51640304d99602f0
z4543f84308e3632e854a96973de48f7ca1770d4dde99841439ecbc8135ab58567855a1a44b3e6a
zc3dd5c73ebdfdf46a668b59f8c93b3adf79ac944987d8f672d05191d5bdc100af3a717144d0f35
z68b01b541d50b61b352ffd54923087231f8331d6f9db2643504fa4ee8c56f7b827fdeb9959f4c5
z8465893ab66a8726417ffb38b08c5549fed39d8d48f72f50fabc87e537825cb7923c8d4aaffe72
z6b3937ecb6c4236af081238627a5aa06d35e3087dfa5ef92d47c8dcaa58f5157aed169cb9e16f5
z4e3cba2797e67d37f5f5d4ed50b77cd2f9e9757d6e28e3456f151043909ba1d2b9c35b5995ce3c
z4b9cee47d0f8c1723475f62763db76e5ed54ae4eb654ff67294efd1bc6b59c4f3f28f85db73b37
z1ad253a3c8e783d9f4600d38aabc218f295992d1193e7f7477587f9572cc28dae51b981e98990d
z285225044f2ee2f2552ce0d8d7115eafff67334efae6f8cf90a3e8308be32d43003a9ffcb0d06f
z5f3fc375682b2fc64506d518afb7219cb6805e693ca2ee9ce9babe83988572c376c8e1ca7aebf6
zca0f61a995310aefd51ec5882c1cfc18173546080c4aec7200ed2d39e0d7061e1c3f6350af0791
z3e2d4a67d932972b8b4c3ccaae51b3e13cf17bc9f059b147cd2e3a050b841d69d5e5db6a58c01f
zf3ac602073c2ea47032d4b2fc7673156f5cfe9d62b8eea2198a037ac70b4896dd80cba25298a71
z139e76cb131ab80cd18705fb01043420d5e6e03d22d59dd10b14a653e37c00173efdf8b7cfc940
z58c9f863333d43caa8746b906925498b101c4ef4752784655a61bddb9b099ec9ecee5c1593d468
z134db69d8990c8390fb036e15be430e9017d929c460f3bc49ae4f0c5feb22b1cf1bf5ae7535641
zd2f24f95f64ba15ff63c0310b1843315cb2ab6b6bce604b6d9872e7da9ac998e6b0a19eebc0612
z9c21d18a2e0022d1566118c53c95fb29871b295f9437d8f5296d3036e769c17cbef2682ff09d2f
z0bda9533f4f7c711376947ee741ecdb0f07366fc6a5715b92720dada729d6989a1aa2cc9f76b43
z529529895a795220cf8e3db106d5428490f9694a42d624b45713b01c124beb2b7f69a5cc777b7d
za0e6c73948ba4300a570092da22aa22b68030c8e4bd9006faa0f5e490461392e6fe00f9f07eab4
z2f45fa8fe2ff61113d88afef7f04c10e56653195e4d6e5e080b42b47d2ef0307991f3eb1e6a6ba
z8203607a95fd8c3189fba3eb2366c032155503a87a12e04c18063546f0a814365dce36ed377e8f
zff803dd1a29088520c21837692a3d834bdb5c77b6af6e9e8dd17298dd8369ed487c394b45ebdf9
z2748fb1e42a063e47cefe7a6de4cb5ffedad28757dd09b22857606be846937e7624f6fccbaa40c
z9075e4b916213544ce7f27c1d5ce0fad434888d4f4e528fe33f1ad635f61a5c02ba419e753d2fb
z99e1299ade56d74aac86e8064fa869e5dcd1b50fd505e1989be4a30dd09e7ea14fa29381410a9e
zc76247eea6d9abd3f2e70aebe90002bf55318e1b5cdd89dc552ddeb7cf9cb41520f9bb11388ebb
z765cbec2e34ac12ac87c6ffb08847f79bcb254d27d7f175f10e0cab61ae2d0bdec2119ddacf977
zfae26bdf855c6b336192fb1e7b1ed4e0aa438b340cfefaf04b5e714aedc178527f1b6c684ebdab
zb7c6ebd7dac7721ff82f12e42b171da422be08a5201a0ab1c693ec6ac292717e29b73b16e375f4
z242374f90e32567cbff25a6a42c0f15d4aac7e2bebdd1607851e899f218fc8fee5ef37eb9ec540
zc543de466e34a39fdce833418462413c11ab7cc9a53e2a44bf0c3544262c8e453d8ab3871d922f
zc11f3b5741a5382ed28584e432309304ced338029b3a85ca913c6dde105bd83c0eb0035e961662
z2868890fd9e65202b6db8e30aefb68f2657e4759b07683df10a22742d677d8b9a5192ee4411a4e
zdf23b3aab4ab87474ff21fa85137b04a359674f609eb8b4f1094098642f29633bc7eb393cf7cd6
z8a0b11c8fbc7632f76d7f4495c854d32fb975980bd881b2a8d5173ca7308a19ca5b7e515243fcf
z3e926831af6f21b4470b05a99b9f09db49f8309966353b79dec332cff2366d58fa85e5b6da5ca7
z02e57513ca603ebb121e7f3e6ec65e496269ab2deaf7837393541723102218893e7a89dca31b6a
z47cb688173c5b14755f82bb9335aa2b6b0f6f9de7037b45e0b9f82d3ddd12df83e3ff54cd13105
zf5b47eedc683883bc52edd713b8436ed81048bd77fea750410a52249155431429afa376a76173f
ze039df7545dc8c85c394a2cd8b7717b6bd1b84ad3328f8d70ce4fe45bdc730c8cc3e6f3edc19fe
z0ca0e1cd87ca17e82e478849eb12145cd019bac0c87f8ccc0b9cc5c0b25e20ecece60fafd3a372
z81729db7f4444897423443cf7727e669061f795f0627857335f9dc04e481ea4b54694cf1155672
z7837fce37b6b6a8756b7077a18a9c5061ea3af0c7fa4f3becf6baa9fc129f0bfa3b312c5985de7
z1c919a1c2f90d8be517b52153d7cc535f0e6776b42d9ea4311df8e4662554adf9567d1b8f340de
z871f1834029a8e404bea5b609d4f4359a0de7085d710de07566df4880a6906a266f5e2163a0972
zdb90c5f9afbb61f487d0f213b3ef89ee7d2e4493868d6886323094d182c86c7eb4838629a73c59
z0d548508715689e84cb011e48af37aa9e9449b1872995c1d4cca56d42c2617d696ba36fdc04539
z671ffe7b56068e8b0df55ec3d768fb35bdac39f228956def5ae4d55d1c4427b049c8c5f7495f38
z02af19c8e627d6408c991878512329472c4c217a771d976c645057c408f4aacc5aa51cccac59c0
z8ce11cc34d7ab0f8ad1492dd57ad4e7912dc1189f275f049b3eca829b282d4cae6433cf790bf62
ze9d26dba2279a0e22690a9284f7014e686da93f38d007f1cd62af6510f210d22d97e8b726c4fd3
z9c5e63a318b4236737003ea93b37132ec2fec573ff0ccdc6dde9c0cee8679036e8e9820d013ecb
z164e2f2d8a1a687395d92b524ae949a44bfbc8665f3848be763be51a0744cc44dbbf90e5846fec
zcde1ab7551ac4dda71b906287a9ae965701399b7eb7e9b2e14c71f1e4849f713cae55f898ad22d
zb8243d349fcdc23e06ce10c5aa3896f3a05eecb98d1d3d820d13fa3d4ca2965ea5d9e565646055
ze5114f23831978ca4f86ab5f675a8f8bc9dd42229f8c6efa006c380e43154fa82f34ce32b0c783
zc7c774be31846f7568068f2e547c89fbc6f17f6af9c67c5a8517fca4571050ec18096267680df6
zceb80a2680d5d45ce98f227390a87259c03bde002d2b865aaf40b3ae2e46848ab7dd202098e56f
zc29cc73027ab4a56e71bad568dc5ad29f1d0724fdf998c07cbf5a8ffeaa735b14ab05dfd37f165
ze747bcc42b7010588c70d3978f1a38567a21aaf7488ed5b38f787fc4ec154f2adc1a135641d823
z099ecd32755116e562c1983c6f019f1fc7e41718bd07dd24bceb1112015399767df33e626d0ba0
zcb7ce550ed6b60935b1afc720c78f7564dfa11365387e4d67ec9608564491d2f95127db24c5664
z84dc07f6fa62c5c2badee109fa2c007a05e608a544c55dd32d374a242406a05a4f2d2bc2fa061c
zb445a0b7f1e36deb8810cd8ed861de1bc29e91dd429d9ebe2eb00b43488ed13fc8434b2c139d9e
z20ff6ed0a5970d851bf80df184edb4766a64936ee30177ee7e22f5f429d62a808419a620dd4bda
zf255412d8ce2e4564343cb801fde69673ce55405a6a172fb6677559c3f08edf2e8c6cd06165257
z8585b892299185bc2f6b45048a54e9c06ca6d8d7d4b2faf6aa8a55c694586c55d5bb31433e9ba4
ze935dc67d6568859439386710fe191442036efc9a4a6a44ef82c01c83e8e3222794e120a03215a
z74eb1c9a23e8322e98df6068c7ffbdbe806c7953af6d51815a9a2d8d4d94201831b2c2af61fde8
z4d2db413a9c0753732228c628d03a6f54a9d1e6e6b4ef75bfb6666def877b40e2cf56021421ee3
z7e8a3274d7d257170e46c3dc9311d3a984aa8814f025519fd587b2589173148c9c6c2c9f2bb733
z17b011bfc5e5d706c755f3e4c44b7636e01827e4b3138621b19a95c2b9a2e1edb44970b49d94f7
zc19b491dfeca6241daf45bf78c81b6c672b64316a6719151c91db5e04c35d5f56d359e5318c3df
z9ba335515f120df97715648d3744f83bef263c7666b553606736b5cce172e45e23b6cecfc5f0a6
z7160a092270b480b9efd2d265c241bcb1f73d81b0963a7a9545adb0c1800939e54b9904e35b0c7
z635f3902c8ed09e7922b7fe17fa7df7472c8ae6afd28102a3a2629e1e1e13272448dfaa7b7ef5c
z6c506b00fc32f1df239a92958a72714b75b8c1dad648f4115f4ab072e661469b116d769a7aa1e4
z80d2d6677a9d41bcc33d518777904472873d6388a3edb88a44215a01b0acb6f5305290635789a0
z6eb1768b0551af3bbde8fb72c146689d68025936c9cd0372c1db5175ce6817ee5d8fc29294f4c8
z842f4ec50cdd83567ff78f32a24fdd4ead7a1fc7e641496aedd56e3fefededf001855a600f0fd0
z174ce6b692383d0e7222c934812750538007b836d92b3fba270ad8e10e8a93cb81f0e550cb8874
z09ed9808816b86171650dc2b25112907584bf9d82a5bb2cbc31bc2c09be9574d22fdfbe3b5617d
zc19a63b2ea8671d772cc87de08755a8de2faf8e913e7fd10b60d00869b178ad0d96aab31423dc7
z7ef396fa0cdf2aa8d2483c96b667a88aa7aebd73f92928fe462ce22ee07d47e20a20224d69cbf6
z877c1a348411d16c0402446782a68135407fe4e11d8391dfa0fcaac324fc340de1a194726581f5
z4dea3c87c6fb76f5e396a955216019b6bd50dfa61ed6d57eb9d92ee259be3f9cae35a3b9b9549d
z464d83d86e3b4e40148267a885f58156a02c8bbff65bd4f9351c228581aa2888727e16a5fc1cd1
z421e619a91e06b58ce93ef5621efc8b2da5a0e9e30cf5bc65cdcb44fa0724dfcf2e2cddd30fb0e
zb685b500bcf29f893fb39d92700bf93b3df6ecbb899952bd0c5211ab2fd2fa5f4971d1c295f2de
z449b947521e972c4f01bcd49bdbdf67d1d90ce79fcb5476ef0f96f2f47184a6846b4bbd1fe7535
z1969f61b8100b9f8a1824c41e90d35336a529259b6b3f85e498fe8c42e3a55f5030d6816e489df
z65aa95eb710120eafd30a6b7e6c5666d080d840bcabf1cd0407efe16d25ca7d882e441872c8664
z3f402d6951dca43bb066ac6f119ae4cec4045717a8edd7e427b03e7425c98f3b36ba55c12b6409
ze9a2b740f379ad4b573aa1fd89642deb47391acf6a603243c815f5ed29bac8c35ab2092eb3572a
z03b9c3efb427a965c3d9c4cf08aa31f6d86d48e07274de345ba37c299d1d445cf6917521ea6e6e
z01ae4e65cb5773ff71533365392aa4b6052b7527df97024d55bc93ec0afedf1beb1c43d4884fef
z1a1eca09e30a6bfd3d7686123b9078165b1052abdf7697e6b8c85ae751183a602777f7b24caf12
z6ee0636dfc66227a8cc56fb14ef908b4ff83a44afc5fd88a910b1489fc48a3e7469e7d2d16fa15
z29dcdff3e1586bc19ab059cd000cc7e8f28141ea8a77139c6209fecf6ee782d4851b69ef45ca78
ze8ca57c82308d8e91098c6e8e0b397c06c36f77989899085750414c3b7a5c62ff581aeb09771a6
z584d88856998cd29f8bb90aa951d16bec4c8c1a3c252608485fb593d4ebbd16dd61bfa94e8badd
z010ed32581eb32cf10338e016b22019d7096e9fbbfe54d7635b69218eefadd7a8631f9ea06a388
z4dfb0f492eb13fb8b8ea4eaa7dc917b448dfde4e9dedfbaf766b9b8701b1efdc6d00f8d29e90cf
z46ad0ea0d5fd955ac331bdcd2d6535cda9c6e61d19553dae299664fb58aec5ea18574476c2682d
z8325739f6693d50af94054dd04bdaae66c818da883c1de35e90b5b5d8cd8081897ae02a7171af4
zfd3c8881156581a1daa5bb1bc2c81456d251689a7e4899c908873bf96072cd295263b6764749b3
zf6bfec28bad4f14d34bee9b8caada1cb71db7a45cce52f895ededf61bb25f4595d8f5d98fb12a3
zf8a433c7144978d52d4e2ea1185daaa34da3cb2d018fd24455516a7165aace942a43a8d520b8e6
zc0516eab01c9b12fc56077f41ec43aab74467616057246fc0b38eca580121eca5db15b1043750a
zb641ea82c6beff8aecfeb2f14521faf30c8099e5aad1a4c183e2cc19d605ec8295de83b2f4c882
zbcf45094f30024e3a09ae8fb77a6af70ecde8ad223af0b25f9b86054c899b59a53b0188cc0c983
zda314bc59bf0e8ec348f0b5f90f48fb1075eede7c2d2f30a6a3489ef7f2eca7474a03473e269c3
z8224c5f68520686ba69555c1ff5c04cb71c86fa12afb6048036e68a5efbd72627df2d7809097e6
z25002a759bb423c69c0feff1d18e892a74af194e1e09d7700c9d9fea04088262e985429023460d
zc81bd31cfb2265186ca2d696dfad36f56124d3a7aa2c54bfae6a1aae77071d427a80c5918e2185
zb2e509fd1b7c2161ed1ed6b6de2c26bd521cb10e510c574146a49b3097cef730de8a3308e577bc
z527777109e6c59c1906fa4fb57caeaccf674050e1779fa88efa4d154ff2ceb54e063dd01f09e2c
z2929815930851cd756089fe36736af3440c5f919d8f9aac30807933ef8385231e402289cfcfffb
zd123862bb781beb8caa6b83ae150616426e3b4763454d7418e2e0a656def91afbc39c8b252813d
z37c87fa2a2cab3a95fde9562f66514881d31e84c2b75572c9386a2179b8e917697e1a5050b4b2b
zc1533fbd13db543ad90532d62de2db978e70a0458a8cd893427c6704bec59d449e1fafdecc1496
z332e5b8332f978c5bfbc64f4029cca46c7f08f05843d78ad5824025b9fe51aafa3b464156bdc32
zb810f071d1b16a8b8ff0a85ef18ccc1a8826a8264662140d64a2823c7a417f5edfaba56260b929
z4c587f1e066083e14ab83f5a8d8dda6a8687dc0a12860727c001d16f88e280d8eac1d34c216cf2
z8e7992cae8ee454b0676bddd9f7437cfbb2a180a8367f223a8c18838a456aaab8022b2e36a5781
zb7af39136bfb6b88ef90eb3cf99e0f7ff381ad278522b0a9938a31ceb2de964587d1c287268149
z719cd05ae853838cdfdf7666a51d7b360084fc1d9cb8701bc98cadc7dd56d9cf3d38b6669c60b3
z457286d7daae9e0253419d8231e28f26374e773ae4347e67d196dd0ff56e08595ea34f2ef22647
z43eba8d7f2b4528c2abedafd93fe4fa10ea4b2668caab13c35e8a71bcec574807dfa99714272c6
z62ff2aee5dcf49f1f0019ad2c26859238f051e2a7705d2fcbfc0d64e9f390e4f328406b9ac6dd7
zc81e2d66db92ae573768575a8f615fc903e4e49594be346eaffb9dbc8c259877e9e3365ef4dcd9
z5eb3c2dba78d5147467dda6c0eb133d3e9ccd1b4c46cf4ca4f49876bef89b45f15e2261e570a42
z57982ecc1bda8099ca799df78888f408b63a3ce89ee2cab573819db1202da9250a3cdc6a23805d
z79a6db159efe781fa691a3ff3d4e6e1fa10ced580e1372ffbf72f6bfe1ca73ebd68f3d897b7e9c
z6d37876c459ac1d1c3a46f650f6898d03f5bd240ba70d40a032db1188b133aa74562130546be05
z97ba6188435d7718a222398ab263d0f844633fb38cf342b58ca8e68f2171939e81890b5c0e5f63
ze9b4d572b42bd3de3fbbcc9ca73dfaaaef322023c2b5a59d524d10dfc01726160b70ca0b7d7e23
zdb9bc1a45e49c1865d02af11a75a3a5cf76b0ebbba09dcf4d9191a6d7bc9560fbdfe6327dc5ba0
z689f6d0e12afff8efcb6f0c98589f5ea6c64b5bb6b8cee2d5f2c69a8239533b40a4d68b79f4121
zf14f5b90e56c4bc6afb00b18951e3ca5ae566a3fa7b2c971ae0c2e83ad4983f37ff9ee0935ae85
zc0f34887e7bd426eebb093ec14f3eb31c2f491ef7992b5fd0950320ba9569df8befb4cb4aa92b4
zfdf05b80a4a56fa8aa74a60d393bf7d9ccfd3360fba346667749f35fe6f1dd10b03c1ecd0a50f1
ze79a78ab036e9904df6ee765ce925e3caabb62e0c5e9c4a7990d8fe4c4db8b92b8ede430366f65
zd6a221f72465a65aee5440c3cb35557d9d6f6ed256d9e47ef07a4c85e297ab0f4d3b67c8a80bd5
z16a06ffe3cb4a48febcd3a230f05d7f38bbd3c457a803c0f6f73695c96bde4fc310066706b3565
z5198312566a15209b92ad29d2aa6a29744eae02a7ce2f953f10a2d1b116495fef8239a355f9d9b
zd32a9b474f507f9cf29deb48ec2e9833302a4a7b5f1407cac862c5d6faf15a362fc07ef6ba4294
z405eb27b609640d871b073d36823f8cf5bdc3652d06cb10fa57673f5990a3ff5f244bd04838112
z933e80ef2c19219747072d1a46b8fc870519c1bad9dca4e768ee102d591e8f17b0a1c5d258b22e
zfa8e697e29dced9ef5285f0b593e5413e7fc53e085397ee55bf303f4127f98f1800bc911009839
za833d7bba360c1572d5cafa8d272b815dffedd40acbc1c2caa161e83ce1813ebff6fe8a013ad9c
z419e63a533a1f55b25bc5b7d108e1317ec529283943f18127d08c15b695283cd4d4272a1324923
zb5f1342ca2e0e50ce8b57004446052f0908dbaa56d58e6cdf605e2a134c27b994572e45d9b40ba
z3243db19671dbf64cbe8641d932957c83289d0af045069d3a89d6c1c8b57ed5e3a89cc20f74798
z01c638b967e389376f0e113660bd6a19e002e00e31b27d9885a751fa5370709b4c66aea0969d8f
zff79ea9824fae0942353cc8bc37cf9b6a14f5af1dcfb79dd8debbc1505bdf9e93cfd7c81e896f4
z8e7566823b8826b4d2bd67713c2fc4fcb7fc0b855250596a00a7121aa7fb81101c0be229f33e8d
z699f4a545841d7d4920c7a70069cffca69f10de6cbd8b4bfafcaca3a46947aafd43b4c243e0b4c
zb5c9cf99ec866adf641ae639d44145972d128c7d1d77ad51c232e35921bd75bec0961d4a46f3fa
z4602de23434b1be9a327491f1bdaa4936ee556e352d29dfba5322dfa944cc074ba4b0271c8d3b9
z88f53a3f623153aecb86c40953e1ac30d4fca069137d541f402f65806a82d7e64b400370ef132d
z6ac214db06697b8b01905ac59c050dee31541d06777db5a91e884de37272e5c4072525dbfde5b7
zc9d228e3ec1ed6b5603fccc58f4fad0de4468659b67eb0ca9a129b7d113966269b8a007c74692e
z6d4f971b33e05ff50a8fa349e8658c73317e03d5816ce2517cc8b2dc8e34a295d7a199f5080a73
zb95fc8cdbfb75416b16b3359a9a77c0fa89e32bac05727c3bf3c65c9f766f0750dd753f0c90041
z9d65ff8b836d28cdcee54537c5a100eeb4148300fcad63b4b409c1b2e8d14ee8267153293b3835
zf9db06959fcda845ce199737d04abd667544416a13b925a7ef51dfce223eb581e5f9328f49bf02
zb046b2823bc6f68a3ee2c0aa40245be5ffcfd5353a6ee625e5bed0b360d7b3c616b01107c82655
z000dcbe53a9dbea9409e9615e872b3b2b12e821a1d27502baf19b620dba65e2b8d11c3f7d0eac8
z9520d70233c0c5946828c80356a052a01ef8496437735d71d95728ff4497184c7a168b6adb37c4
z7cf7b4ad79c91a0a522091494356a16b55190aae09c8124f5c9a8cde3fb38abb6c4be491f80a87
z69d34a4ac343e1e8aeb0266cfabb50349630b1257a0d7524df5371dbe4c29ed543ebabd8cf4b81
z553fc9076677f4d903258f0ea7c44ac97e08d37469fd9780a0b409d0d5ebbf315461abe23cf1c2
z426a400a22c0d4937f847b2aeaa5544dcde0d0ad1b1d6b1998c970afc10a58b8af3f56dc001e27
zb3e587461b53d70c25b5ed82759a6180194acdd856bc4d9229bf6a56b1145b82d1ee4798fd3bd1
zd613e9f39431aff1d0606324e03d2b5f90dff059ca02075561547e4b2ab3fc8f6d473b3665698b
za06678622dab126f40968e1c4b514d1af1c8bab59d330a3859b9b632574646927a8ca97e2b2c1c
z67e6accb4a3056741a7d5107c11a7d8e8e71a672dcb5a049d566281b4836343f3d14a2c806c16a
z6ddca9595cfc874d209b32dc1ed135da37fed1d858b85e296e2a287f24e33688a7ca5bf3890a82
z46cb91d3c7696357798a8ff4a43384ea0785fd08a4b17750592aac3563313a9a350324f3271c89
zbb3744eaed7386877cc5858787d01199fac6a5ab893bcc14f26dabc41dcbb00a5f331bb47e0be5
z42a24c15c8bc0b72ff274efbb8c1e148abb6827f5ab2ac3833074c46f6e83bca52e2de3e1f5080
zd964a2b55fe32106f584c47a894db7d9426e11165382b4ce4accb0b5eebb5f55065f9b92129afa
z48c446030dc24e61d7e6dfc191bce7130f6ff60239c2786f7a589f2ac5f343f7edae966c6af831
z9a712155785fc156e603da929871103fd952fc82129dee3a88eab0ce403ef1eb025634ab26bf99
zf940a75778b3c0f64c4e99d65d7d48106b3573d3267b396cc7f4d76cf35ba44ecdfa3637879209
zd5784d9c2a06b8b35e3160123298feed2d2d6f5ab0a5ee9c8955c384ee223f63b9e5e74b3ad43f
z555efbb79a022b43383edd53a93f5cfbb987d55f8242b8baac21bbb4cf843b5bc02657be6b185a
z8b3ccfa9b45e31790c3bcdeb46949c1e53361cb91068cc2efc5fd1c1645062b36e261ae626a1b2
zc11a623c9748768c70e35d69c0f30debf336487eae7e02eee4e2f60bc33a9a1faebc2b8c0efcbb
zdbfd4047dc9c3cde977205b7715c1fc6a09e20c45c4a0e059065481c231afe913f022cd980891e
ze251c736a27bcf61152e599f5c7bc0e1689a1e2ef30c85e90c72908e8b76671602e6fdbcdad4a8
z4fc35758ffea7cb544f361362a8a2c98a2aac490ffee9ff40afbf601e111a7c98c2fcf52c8cfc4
z43887961283c567443a65ae55f8e3b35c6e69c9117290456f6bf42f9a349a56da7b967d440dc3f
z96cfa1459c61b686048422d848a4753b98c85f4eafa66ad2ca9af58b00c4f6a26e15868282bb7e
zb0b9eec5e79c0987e7a2a4daccf5ad467f639eb987022676d099ef62b2ce1c0c214c2fd06841dc
zd341ffbf62326666cfd6e36c1b424c4d21cc8cb42fd619ff7a8e6bdb484581b03535acd931be90
z071fe48c54fc59a162c84c8782c01938fd120daa24aeee0e73d85e2506f0732203bcf83b0d4ffe
zb5f3671802ad22c6239a07d741ad2991896b3879053ec76c9df4e4e4df6e86196587f9b2456127
z7d2c2cddf80509a3a67fcd3532b10179bcbc8841339a80395c9874892bbb296b2b513da45babe7
zf6a654082972468a0d15a356666aca29a5c920c0e8879fb6a4fe344b578895d2a5ba87468cf6c7
zc092482dbe4222e03462f8637878bd162f490262c2f1b697b160e316da7127b9bf1c753cddcfea
z57d700c7e56f7d933c13a37217d13d4fca948996bfbeaae58cb5d36ad95e15bdf3355deda805d8
z1cc33a555444d6666282213b17c952db804fcb4fb41c218eb829389cbcff8e16873629d4d870a3
z015b65d2fd962a144b8c01a961c2ff7d4d9f24b7807cf3a94592b49ddf110c0874594073660083
zbef57333477ad48e41fca258fb1a996e8924aaf1b0defb05820ef888c6fe1d96b13b6adb1d2d8e
zfa3926b646be96fe199fc3977d2a248714574fb92d9b36b6733f8e23e5e3416fa091d59f0a6c98
z073a0246cfcd5e94ce33506fb640d06edd1bcbca29ad8d6a3bfa936eeee443b7f106283cdb8963
z9a71f42a60f010895729ac3d33faede85a73dbdd516f2968782824705733f9136f01c549e67b7b
z82b31de30a864c9b9e14b681d415922cc36d50ca6fb828ea7e1e39db5fb0a4a590dcf7273f010c
z5288808e13c2a697b89c7e307d8fddda619c9267d06b3d2cc064091c38fd15f0e0518580abb4e4
z0cd71aebf3545270b8321ae76148f6dff9211c79286f69869bb3b29a7a41aa6d6f59bb4d54b510
z81f4f562ec0336e3d8c7dbefff53c0d842b494a7b1d422d38bd5802d8fb40712fc7fbb1690dfb1
z60f52e290ce20cda9f67f63c7e7ea6e190e896f1a8cbb9af0d0fed1e5d6516f48ab505e744e99a
z17a53e86a02687dffa8fc4249e9d150a104ac1a1e7ed89ebcb23bfac524261c49b65c0f1aa8819
z1418aa7b21aaa4c1c5a4832d404656a2a402c6a90d01d5cc1149cf02137ea82a62052a5276fdf2
z27788e63222ecbe69b038cd9eef481febf520752ad60b6e36b85665142ecef0b8fc4ff037efcab
ze536e09b63e18eedd2eff7a606b28dd88e19f06567d69fb215717fc8a602fd60ec47452ef95aa9
zbfe9202a92ab86323a6389bc71f354468ea481d807ea1d68023f82f51c213cce4e528bb86ae63f
zb21806a6fbdc8fb88da1bed62ab0e7bc57bf6cfc15e0a297fc2a0861ea339cac390e341b984466
z1bc02299c9f0f799e54972762c9518b888e3e4cc09973cbbcc94aefdeb4b36954669cbd6aabdc4
z8abd82fd15549ad051b93a3de4a9e63034eef18c56d15d049cc859e54a8245e21418d20670621f
z4cb6be22a4bac9d6889b53e60a3a8616f54812df49aa6f9564f065420d57a582de76c1abbd4698
z8cc80e93a782d4d1318a71c574ce2936bb14dfbbee349017298e790df31e52cbc46e8464e38cb4
z24afc32500c551330db2a8246b7e1212a022184343889224a8b6c146f76d4c48266eaf655ba77d
z927b6854f719db94b2357f938c27979f25e8a7dc345e42aec7bd87606eaa5c424428f863a261b0
z72313bffd14934daf9cac7e84b45aeddb0aefcc2ffa15ee753b5a176727700acaa6fa1f292e6f8
zc9ff1dd7a1e61e02ae49541a1eb551ed6eae2e64b28e5c25603c60631231aea9fa1055a3f57c35
zca3f6b168a30482954fc8bd3d08d8a03a56f92cecb2d6d14afcee6adb57b145c8d67af78d867fe
zac4cc3b843f5aaa8c6ab5ae844a50807e3d331cb2ebd3e8ee5f14364313560a2932c7985ac4774
zef8371158f8b1f5204d629d177df27f90c4f6f0338807d2e710d2c4a467ae23b5fad7e936fc870
z8173cface1dfb0831bbaeb76f8f1784f1d271304be3c9adb9a0e585bb3c0af5a72cab962825c13
z86ef864bc724500c2e9fdb5d1e5ee348ef4d578a2bac0dac8cc057846f4572d48dfed141bef9d5
zac5e64eb662f10a77c52343651302a4f609b2d3b9081d770793f9b312dc97b15a00603c2e9b652
z1d0a4fd925b7d05e544f5d0a9f77da0a4d5c7e01a560b45124cea7ae4818f3ffcd3908e04e9241
z3cc5ceee4fa6cce83d88d56d4c5bf9131019298c00256ae69084a6647822500055a51fb93343ab
z9d3710ab1635b0a49af7399e760ac344a1992d5a8978e1c9a7fa6e90ac5022e659f907e8ff26cb
z28c327eebe5e118caa1d6fb14d9704e98042a81f31e3c1825d63063e22189f830c1cf605f920ab
zda9449b53d5b65f5d5df462e098ce9f061cbe30d6393cf7e4aab054cfc197b627d5e59f9c45e9e
z84748b9548b7d7bd401d21acc036a37ea993185500eb7d137817c2d53eb1f282ec490ce991c9b0
zd92eac77f9e81ab1c7db0684f58466db333497622a4cc6522fbce753fac3ac3ebe0f8ec2cfc1f9
z321de52f4f6b95a5bee691b4b5f927fd7e66fbbed7f1c375474072d5c82fa7ea8591bfc423e496
zbb1aad3d12eaba6e948bce4904c7ea0bfb299dfcfde72f8beece2c67e43e17935ba36b20b1b813
z3a134e75bc96af6cd2fbf0f9af0bb3ecd48997c1980dbb077583ac227e6c789deae0a332845533
z8196614d6e2da0822a8f6859643a26619b1e5bd6c42b11c592b3a5903e26d8d1652e7f7bf1f92d
zacf33c792f8eda87835d130df433991aab444f60792da3ef7039d129a322398a3cfdfbd8caf6a5
z9c762cf1b2a00e4678d7debd39dde4bd454f3bc87c6b151cb919df38d3943efec3b94feefd8104
z53794068771a0df7eae7a0ec08ab482ce11e8690eb0a38516b1328443cfe0ce7ca4d506a7eeebf
z0a2a2012125ef5c4f19900e0864b5a8d9ee0f0eabad97771aaaf3d809157d693ad6a59e4678d8f
ze16ddea7554c8c066e94f2a2ca9caa323942fb9b38f5009b520332fd5d5884e530a42c062e5347
z3656dfdec460d877455e1fb25e2e9dc47718c62efed0f6be313f279afb508bed8b0335bb6721ba
zf81ae39ade2ddc79066ef8dd660e31ed66c2b0b52195657ec34fbbe7b3ca985b0483f80cd3cce4
z6f0db3d211526c94f46007e86af5d335fe22fabeec998a1f3bb15c1e68c448f9a34cfa21f8984e
z3dab6c08d8eaa7954d11da3d0102d5ee653e59089ebf060c633ddee81f78024151342c90bf34f1
zb296d5506192f1884f4e70eed12452fcf395712b46439600db869bf854808bcaeff192332f6e78
zf51f08886119233755cfd0b4afa402fa5cfe215c5ee9336ee3ff1ff477bdeb8d28eaa9746287a9
za4583b05479f56934506d3a9241bcad812b33e63165661f18263acd3154e6dcffd2773613a5da7
z879333bffd874a4d75c5689d785c786f58f554cbaf0f6de9ccc7274edb1300885ee227745c589a
ze0eb7f17337ccf9f2879ca201f694ad0ac3fc1f2b0a2be489555637a9b4b8e4181e0ba657c7b4e
z1522ea686bf917ef2f8c235361c66a303bafc66f4d84426e5c021bcec3a4fe4cba0ee3499388c9
z0517382f3e3b1b10a269f62e54ea3c35e127cbffdfcce98915f0949cd5f70d291f14e3fa95d7b1
z58702b9ed5c6a867fcff3cc44823f74cc3b992cfa00dbc51c4561a8d4f12ed90bb00cbb13ac51b
z033630c844035dd9d4cfa3ffaddb72b01cb00df70cf333913707be380719e06b34b0bdfdc37995
z4a4823b57f1ba71caafe10259972eeb75c072b02a79db8718c65f94ef9e681497fe273507fcd5e
za1a2f366f0f621c33ca6696c77f6d0f85c663017e34044f58a7cc97aa8b70405ee5c67cba3c8b9
zd21e5773960cc7a61eba62cac660f923578ffe31343a10b4696b46e99851491e891bf011f534fe
z1be1c06653d100b1e46e9ed6f23489629d1b3b4ef5355f573f5f08ec0530ef49cd643026caa834
z2dbd135724e70366dcd14f3e58c264580d7da7add56d6ddce4a2b0f5e0a8ca1f57269d0ad70850
z4f25d180e0d6627b1453dd89e23eb7ae2978d472646b758ca24e949bd1a06ef8cfda26720e473b
za75a3ca48b9bdcea4c2ce818fe57a35ce8f0336f0e6a1fa163b2e16bb6df21c11f8a1086d80de6
z546cf85476bfdaaaf196bbdbdfe917ec7a59f8d0d29d4d5c8aecf96da2d01f12c57c8e52cddcb4
z2c50c45b369d57330f4fd8217d284debb0a807587e2681257f2ceaae24a393acd5213669d3955f
z84cdddf7631e78cacd74fe853a590c895d4442aba5e8b764df9b5947900886149577d7550893fc
z57a94ab8a8d0ef636360663d05e3137c69153aac1e52eb077bef047005a2ee9b253dfb22cd9cb2
z5883a4cd622e02b1ea8201752149b6b98025994822a379401378417952453dfbcd8286e12f1ebb
zc0e35ec6c37888e6b2493290a98156ebe3ea7f19853f8283a2191d1b505a06be64cd4bb1bb9bd3
zd0858fb736b4253d3b600d081591e5e885883cfa0196609c5a6c57d4d61b90eaad94447474ee98
ze19c5bae8718a715ff031f6b62e9d597d4ed265fc5a4ef26bf07106bd7c238dd87ec6cf04fa9d2
z196bf1e50a8d85ca1c607aa80b03223563ad14123c95e9ac0bfdc483d7f0480c89f75b0b8bc749
zd75a792063eddb9a2638306a812abec9aaaa81d47b14a0c223299669188d3ca6e1c4579fa26dab
z5b0a51bf426d598938036db52debbc6dc9f49af3e7b961b8c975b746685e03fe70497afccd0235
z3a57aa78d8fd8d54e2a8dbbf93ad07c1a9fc4f983249109d675c03a418f520bff62b65eac7caac
z43cc8717420ffc199a57a4ddf337cbd2e1dbc607e821203e4f8f2b67962badd092454b6115cf4f
z3b96d3454396d67c653c9167e2cce7a5f23e672c058c2990f016350cca3aba8f261f294b02be87
z83a7d6d9b86f855f45ae6040d6800ed77c3d7b8c1a1c93c4cf03b61173b1536a77ed6e196fe8f5
zbc36e5713ebd357d322155e3ab0137ee995bfbedf8bdf2d0a7f16226ef4cf8bc060e5a35df54f5
z68d0018b985cb3afda6099f74b99d5a23fe043f141359e9ef89c249ea0c5f08478a7181d154d60
z77d2041401a7413c0e6799ba5040a7d015aa9733c969bce7206743a291f14485d807a3c01251fe
zec1300ecff1e93f2b4f68209833afadd100f9b33317a692f4d8f75574c0a2446836b34416f84c1
z1dd0d0738b3204e686f9a51623cf477f3be6fbd8dd4498f4175f49e4995806dcab595098a88dcf
za9ee9ce6ee5e190c4d181412368ff1e4d72b9a70cee4032c6922cdda2b8f961121b968d0bbb266
zcdf8e320d9f35bd2775112fe2fec8741a4e0b4a7fd6f8fb69e4cf05f685b30107a4e3a7a5e25b3
zd8d9f4f32b0969d6fb72b32e51b6afca6a49bb3986a8fa628ccdf8bdadd759269a06537dcf8ee9
z07e17a0b49752c124916a44be365cbfbf2661ea80131d1c6914053773e5187c36700f0931beae1
z63644e0110631cef7d46dcec90544e2bc21f1b7f2328d20dd86183779e09a331f110fb5217d2fd
zc544b12aba3aa42cdd373b41a785ec9eda85e31e5cf31b759028039118c870bdd8980be323bf14
zbf7dd6809d3b9f09c1426a2f88d19364fb0907066b59917c8c402d945c0e5a54ce6ab9f1808f9c
zbf228f17a8c35140553c62d2253c9263f4c2019035e39243e268a755ee2f45ea3eb7b6caf75fb9
zea3fab56a42efdbc085cc556ee2997a2ba716255e6f823d4ce4bfac900f8d82fe4bc4711b9ab8f
z846d10682fad42c2a9b214db57e8a6fc085cfd585153fbd9c2e348f62fe8abf4d4a53c3760931c
z9cd2903783bb8a431cb713599877d99ed88e3c44f963f74f5086cd15639278948950e51abca679
zed1bf58f08c421079b610b58374b859a50587a4b08d4ee6c0798d7e3f894f021b3bd8ca31b6187
z519e2cddef395b006c388eea0c58e80411be11e4411084de886cfd8f3a31b4e7e6676047383f0e
z18484e1ddb1ab6a37c7aa20a74b2429b38279fa9117cbf72236515bbc858e07d51f8842e64318e
zee37c0369dee5e60df17c4a2d3fc81a60a59f3a977656d4bc098e160de37d4bc34caa444a8c029
zd40ffc2ce80e6b194d16ae1494f6cca80c869c99c80c28f38430981d1178e7bad5d77908f3a34e
za17f0fd682493d5d9e4eb8481eafbbb71591db1fbca80d76c039853f60936e4fa74fff66a118f1
zcae450f67cf39e186b97a7226efd1048c68aa76d32dd5cc4a79314e8c0d2087e253b13d116be75
zcc0c77ee9c631f2225db834443919cfa079b53e6f4e61a602e6c06404e17c3c2fea5af0e570cae
zc225b44fdc0066566e77ca853b2ed69c2c8e360b123043cb8e7a28f4689cd405a30e2e576aff3d
zfc714b6046f74f95357b7c904f09331d2cf3017074902b60e939bb175dd29839efabfb879f5c03
ze8a4d4d669c5777fc9b4781a13f0239b9510c076649675d4642222403c51ca2a63d5aace3c7b40
za1224999096f1ed1bc7e0109d574199c76d74123eaaac6e7b9bc47076a824e92c3431839002fe7
zf0828cd19d15b6b6ec965c897c52b29f072855e1e6318082489951ce9cddba85ee748f0924b74b
z9b80ab4089748c491e67b3a9d87720564257853fad965f4cc0526c6e49bd8465d2d4f73b260e8e
z68e654c7cf881528c2c37de4b8b0e2d875f4c3b2ea2a1b697dbbe87124ba55e96671898bbf618d
z786085baf66f7d7aea4735f4516f6d90d77c6c284ab3038edccd8f4e6a9246fa92472362871031
z641b2372b180c3fdaae83e438c7b0aaa0c077fca66ff1770861c8f460f9f450d4fbae556f3aeff
z1f7e023386714abb1ce2c75e80fd1508012eb1c9538e26f884f8cf063035a985a6cc71901f55f4
z463d4d18c218d8f9b0d79a38b9497c6711cb4f2b630a7a1bd29b77f45bb1c9891b28e10ca3b0d3
z551b47474cd0b6b1c36ce72a98169239ac81802ce8291cda503dd42d2ff02e6056e1cd8bd738c4
zad43604a5d12b95f00a19fd1cf3ef2d30a5306546a8834f76f8528c2cfa31464f48cba347cded1
zff9d059963813bf3a4a6e73d02641fb9e847b013519a0b4ed523f64fc32262dcbbdaa936458a41
z580665819cc582f9fb8e837f402ce7fd0751a53b17bbfe00adc9cb8df27d59bad3812a9f4dd6a7
zfbdc8de6d419e7b9a249a7837b6267f364bca5c643780d4918e0df82b0cdafe814a4a52106c73f
z73ab3b914cbb4c076e1a06e96cac617b611eaab432803865544b251e29660be486cd97db782c51
z70dd275ddae609a55371cb2b4840f7572475c382d6a1914a6b08ae0871319a5b383a5efe0197da
zd934522eaccd5e0d5e99c22e45dc540965564362c56d685c77f86e285284ccb2d4777538f2dff5
zf428e793d82e4d92208efb0c9ea93f62fbc9df80fc44a0a0b6d0507256d9b937622a0b98903f90
zdbe3486cc8d12ac716b34690d2a1d197e1126e534ad6640554954aa3d6f82ad809b982ac12487a
z1767244bd1dfb828d0ce90392c2deb2047dda57e3cfd7fa85f9ff191a4feb64afff1d4e3968122
zc1217ad32adf04f49a47db1c88540883c3334c459ef55871e9e1529b50902865b723e81e3c2d3a
za8499f9793006eaa1899d3150b1751fad58fda398b95c087f99380a7a281a2a2a7342292bec621
zabac470a1379d030dc3a1171253133cc0d6aa021647c75b2f8a5aa51ed7cb8f9838e73b0d453a7
z8bc4fa5ce7a2237eed2f751ce926f2b3b6e6b0c105c923fa5b15c017847ec3883570f54ac78a07
zfe203aceefb0e5327c3307ebecf97b809586d2006de181b590d65f8b5d2893be4cb83e326559eb
z4a6afa5aacc17491ef61a26d454eeddb58be6988e20ef8c1db9fc0047085db572b481e4c3c93d8
z600bd9568951afa32aada78e16c3c97b340b6b3dc91ca7b7f006e6c382c53f80157876dde074a1
z260049f342341020a87e2d53c6eb8c432149f1d701ae2594515004e9becd554eaa9799e7dc5b86
za492d8c9be7a5226e06d6d54b757bacab02205c5ff9eb9d9110a3f33c70742be6ab273d9d2567f
z1bf80cd4b10a213f81b6884b5520ca092f5579d6f6faca8c24ae67ffaebd4886a915166097dbe3
z040f8d284f449fcf8fd05b5417d5482d0943f2bee847e8c5613e0cbddd6645091fc1b24b8d4802
z4d0718e191c0d7a79e9d6caf6dd5d25894c49e79c6500ae6d82183da413f289403b6fef29cd8ea
ze1f14b98cd9a848a69536d9878c1d2e58d762b39b9f4c32fc61f193b3035e624c4149e26e455d5
zdb930160855ed6615aa5c030539b1a3d2d9608de35b653ab9ca74353494a8a0821f8e578961ca8
ze0ff5343c8178cbce5f5c2fc765ad05875a6bfe8be28304407b0d2f553f8fedecb8aa9104cc1c6
zb0d3358ee6f55886a2c236d74b9b2dc5a5d4b08632e6c9539ff4219030b08beba38c791e459ee9
z3b902daf4f5cd01dc0e13214cbfe6fc5063579f5666d0b3655060743c15f08feac6c69a4fb7a17
z448ee305f7c38ee77fba66367c455b1e6e4865e286c2e54868f8976c6e97c00128618eb18b4f9c
zd5cb76057b685001205840ed6e1aa390de02ddfdaa6b554c779e5bb5d7f4dee50be00e17bdd507
ze78e116f29c176b24c5a0863b755a16d1b3bd25c45d39b817a5af012d4796fe60bb8783f5d6169
z3fd6338cfd5f420db33183be885520f7cd1f27b2660d69203d08e01dcdc628b62f5bc4a59e145d
z9a01bdd50588fe8da6ea183be1694c7a7014dc0ac95a86c5d28127a091af1103bb553cebf9e695
z14a49f68cc1b028781abc9d790953da81f01740c36a91cec11eb9d4ae0a0f2a0eb5737d7ce3e0e
z3a6807e5496370473439208676580088f5ca3e2eb6fdb4b26dea31381248e4aea012f7d8082f07
z1ef824bee88d6720134fc685a1910ff627984c0854a331563a61ed8000303a96cee703be1bb463
z0f26ac924303464a8f86d6dd551be754b58019f2f0cb21a7fcbb255c25d6fd5144d868389389c8
z69547b693a16c4396af188e6805ac3331d911744604e61130675b8946e32f9a552bb6c167b79a8
z96e03ce9c930281aaaccc5d03df9ea09b3aa5d4c343143ccdc6c19062c4c4a3aa2007e3ac82651
ze338b4a7092195f8bc29a9e25c3ba8fdb1afa3281528849929ef60217a8181f37da238767ac099
z4f7fb5bb36579a750440ea18566bd53e76f5e3c750d68ace54c1cf3bea2b9a626b62660abde878
z9874dc9dc99cef7a545a8b77bfc16afeddb05e8a6bc0e8e16f34a9709e8f459054e50a9db5eed6
z2a0c3b0e07a8309379951ac9a7d884d659d096b30a80399d0d8a0ed396e9af20372f7aa4e56040
z2cce1c2106ff870ad70e766fcd3c6dbe491451bc9a8af7d304f589fe2a9ba34ef46acb330e8b4e
z006e456dee331e45e511066921935f3cf3f99414bc99727287fc56724ad9c3fa28ca7fbf2355a1
ze840f9d77368206a00c84a7a6816ae447f7c846634203510467e6fbabbfd2b21fa052f3a847521
za90c20d38eebdbe7bdcd9216626a2b2c2847f937901d41ae2dcf4a2d3237d6a73d46b483f6cafe
z64f657b8739e3a2cd664f019f6e73deb065402277ac6c6916cd3d5a56ca639a327f68b8260da6a
z6eca0a44ea8272375a80fcfb06438ff96e2a6f2180bd062702fd369595e4bc19ce29efa4dff212
z1a1fc0ed9c51ba1b009a4cb43c2fcff5203ec1473bee5f85e35083cdd6ff4cea31e463d34b1730
za0a8a802eb8fe021abb0efd246157e94fecfd0034a4921196dd52d1076eceb3e18f2140c2d7dc9
z27b8b036c8fc3e2a2d5b0c70d57d995166470acd75399904a30d7a052d2920c15b4544de0f9794
zd7066707c6ccb11cb700c9b910469728bef9a71dbbfca507458809604c12ac261c48beccfe2a30
zea9006d9e192e8a1e5fc134e67b6ae67a8f2baa8f8c68413c8edc6742e2bd2a102b2026285c249
z24fea9f3ae01883305314025b39e84494257129581ce0983387d433b9613fdf7f1c803f237c439
zabadcc0067dd45b4f44437cd072e19ff67c8bfc5a8877c2a42b1256fd29b7c8ef61db41e32f001
z33e3eb8a211b2b79292b9422993d713d97d2dbf20f9fd5ad61fead64e326a8ff96c998fb8998c2
zabdc36e57e12e9bf21117964a76e792e81c28c24ab20010e0f8dc5dc99828db17783bb8ee6779c
z07f5b9d8581a2f152735783bd1e2160aa20993956b5a57dea45788dee73def1ef5aafd4cff0d72
zb8bee312ae3ccd507c3b1a908283dce5c7906c58078cc35fa599fe51e8c219677ad171139ba99a
zff683a6d9290eb162858de6081409b79b45b3184afe7c7cc0ffbe3d4df82e092f4c43e2ebe2e52
z12fc401be27b09979a05a2db8680227c731822eec4c3d080ee05ff38e8b5d044c86ddaa26304f4
z6b604be69abfa8e9cd850eca39499a0446bbadf87d731572cead1094ba4f2cc751436a39f098ed
z30e56c6ad07f2761f11284bb1b510e2ae0e27f32ad48198c9dc00ba8a4b64b0768de9e7d6fca03
z7f1c692bd0b726a911f218d8f8b4eb525dbd01dde13c2d9f230598582eade6d8f588ff253cf57f
z0652c153a6d41e509afba98eb16facd9a5ddc552e1a180ff5321708a52124c551895e0474c4906
z8c98faacb83de44be1f5ee912203d3758c432c5e158dc88514226ea2dee5b4a24175a23bbc52f3
z7111648fe2eec497d3b29d258aee61ea5fff91e8c3c478e4052f8c07a0b9329690ae735d349c42
z721a7e94c3d65e6fce60ef6e4aeae22f74fd6646039dc85acadb85b1554d38a2ffeb32dbde9c8c
z8a4429940f9951da19abebdf73c37f7c74d88c41d79fef056f560a686f136ea457e9525f359f84
zaac0219270edc2f1ed5bf6511430a7f0353238cb99732c7391f8ea4c41bb4331bb68491b083998
zc28e52b2fd75e205d4059b129d7290702ab5aafe77ab612b3b48802266ed5462d18514193294fc
z9817824bf28f23c8dac650ef47ef95cf9e985b36b4b72e2ddff592f4c96c9888fda5f0f82ebb35
z32528100822802aa343bbe182364c28beff5007a67cb4a11140e50937e3e7dbdffef1186302696
za48e4b4eaa66163237eed06a8274a903fb788f117d9c23e2d1a627b920bd9b2ca1129e83b45fb0
zfb4e9c4152c94b5b8e59a14aad5b240b1ba31ab8553e45bcc68952b6562e45e0008789922a5202
za384a3c42ff30f0964c6fb7dc98f85cca4b1e37ed38f24e780e39e7fcc9e73c61ddfff92b99d5a
z4fe7c42ce2f6ec8ac20cc21e65e759f134f36d4b4a5da667657efca9e1a646842ee598ed2c33b2
z85b6a5a2911deb5f60d95787da274f3e6242819834a551fba73091d67442a25ae722683b4945a5
zabc0b5360bbc8a315c9a375bb3bd4735ff9584478e603eb81a9f409c01574910f36b27930e7cf0
z2c8f7ad60e2291fbdb7b682791e1deb37353bc8a4a950063bb99fef6af002791a3122b8847f072
z246b69a4ad49c99fd1f3f1d160962465e42353f497e90b6e05f8dbb6d873b0fe40b4c59a75926d
zc9a015a9ff4c47139cd168f84720f9d86fa079a3a3a24c8b43a4a54a82407f21f17d081edec665
zaa2bee37ae456e64e8f835f43d3e6395989fb5cf51419421f2e4e39e24baf41769ed3e2f62eab6
z1a04a9fc226b203c41d68c6d8fe4f4e85485fda9c651c342b73ac1e997e93717f650740fac52be
z312b13feaf073a1d6da58bc6a0140c302a1dd39492a554a281d13e3fe10c17dfb136c27b65fed2
zbb8e5a217f9a09c771a04ce61dd85c92a460055ff1acb17c3851712b30df1b3696df9999529029
ze57730d19194bc614299eca513ffc703e2000d2867803b94ecee7a5d362dcefa2750af453ba33e
z6a871b14ae265ac5920de685d62dd4c86a26fc1cdfec5ec18b727f60618f9c3224b0aaa62f566c
z22f484cc7b4f43147f9ed1d46dc879fb7a018ca6797a3dde04c16d2617bd979935dc9b1e56fd97
zc475e8d7af1a9cb2085a5c88a8bd396e087b7476055679f2645914ef2218da2c59a10e4f5e2c48
ze16259e89320dbdfd92848a902c06085f6ba06f5231d109e28fec27ba8f167434cf4b438b8f653
zb2b0d599e40d4accbb902ef049c933517aff43f16164db4992e0423e029111442c674edcef7042
z4cbe8596c02f486aa322fcf99f60e77dd397e403729b9c6d7a90a992f90cfce2b20e3af0ad9aea
z92a6346616e9d3066ae25e2e6813537706a4ac0a0dfa8d152db2a29209952786e65172383b3731
z35d9c728b1bf31bf4f331b155bd2bb2a40d7e6d5ac5da30d15a0cdf64cbc85e33c63f8bb8bff57
z1a83d9ece12c8878996126167911c9a4cf346f0c18601551ecdff226028ad18d6ce90b2a9e2e52
z8104b815476e133a4526a6ce78306644886e2403faaff8f45f34abbf7d398a745ae66b6a3a23b1
z6e1d7c82ff6f592ac7939ce9a4de29104a2fd77eef790023fefbafac6f302bdf7a5253fdf1b20e
zb156f603f03e2ff9caf4df7b4b429bb3700b84d930b8e623ada9b8cc2b0df55957ab9622245aaa
z20e21b9b37edf4a3efa32ec136eb5059cc746a4dd2867b609ca86d9022a7cb186135d585bc7439
zd30d19c7289cfaffb0d53df31ffaf7a6902df5fd5930557df6f71364fb763c1a8df53dec25bb12
z60507072447e6bf6801f63b06a9b0cf7da95aa160e4c8a04fea19c3ed0f90e124d3e20cfd0a32f
z8f4bcb4a4c20a64534f2f9f6f9a1ded19b58bf44586a13f8976762b0a87f80ea4e00a5e2428d2e
z3b7ff3c8f92473f9f41b75cb9e728ccc7b05cbe9011b23ac25a355b0c557c127894a05c6979ce3
zc976b6dc726f5f73a8d6b07369a9e7a257b3b8602f6c7f8cc88b267ab294c02b87fc89be30c55f
z41f536ad55a5ca1d6e49c775c21432a1f8120bd9b337ec7788ded1959519ae00fdeb51675b2b7a
z768656efee1f8e310e1d29cd4f6d84c082d62a9bd3eea92877ce35e816f3a8dd18a925d8fd6774
zc688c08968a0fad970c18862194377b192bab490c2a64f0aebd8b46f273856be912813d5c015a0
z7e18c8b6e07bfb5354a402cdf4790ca12ecae3c38cd88c3dd9b1ca7392f4c8637bc8aaa4616f1f
zab3750602df007e68813222f2ec753d90d105e91edbd395da945e7914e2b69549073c6cedc8297
z27dfe2daf3ef337903208a6f6ddd636dc5669a6cccbd15b867fafabc3e6363c9ba9bb446325875
z6e5fbdcb75aad5a4a3fc15d12545e54daf86d786e7e1524fa1b8483360a5720c096d7b9260b946
z4d7207212698a84c8d7c2c1c6f829963d0720cbdf45c541f2fd2032c8887c50fccf8bff274863d
z6053b4935769501c6dd21576471dd8b017c04b8f2ee7d078792793965e510f9971db84ef29ace4
z0637f5cb3772cf35bac5f9154fa8989286d8118d55234f69b4bd684993b5549efb30428fa50d83
ze9732ae0c333fb02a0933322785e9baad344f33136c63717496c35a1b034eab3a7ae9bac293000
z764f6a61ccc10dd392f7eaf15dd00954104210046929886193455ce3ebe68b404c82c14e242c28
zd4125f364e37b7e5bfda7fbdb09e4d4df62ac107ef5522a3c0fac0219849c144afd23940753e96
ze230fccaa83d2e899a422d541600b8bb86983337bc873caa8507a46fae21be1c583bdec5bbc490
z635d1f1ee0bb61dd903c68ed68ec14f9506a8e9ba4c762aeee69e7e29cbb664082b789bbf310b6
z38c3b2aaf8c54acf580fd3412d3f8f9176f1cb193872779829d52f96fdf9f624514b5e57d09a3f
z0eb131d844aba00ac74a15f2f519475bf2feed8c6804b7d633389313443e26f5e3c1f91295dfa7
z1636f068c1e458ce4f3606f656657fbd87677060402b5f3002aabbb6a1faedd3c030165651ab67
z7f2ef08187f55dac7209424d6f59ff02722b7c1f9f1615ff8377e134d92742e4a643d903d68fce
z6cbd0d6c4a54c83c3c0e1abc6cda4bdd8baecf82e7d3a989288bc73a8985f91e9d1d9d4f8c8a6e
z59a6ed770c70e55580af2faa408b9fc97888084bbba215f474a986cc267e8e459ff9a334a00368
z7e66412b704d21c4294ccb6bd19c688e44f36dd823085e8fbc8a10a422bea58f76cf93944a8850
zd923f31a05891a113dc482eec3dcf131cc3672b0a40007ace60c58b36f8df9c00f7d7d625dcad7
zd8131efde2818bda0c700a900207ba017a48df7ba590395b29d2af5895d035e0f6f30bd9d8bf57
z19e83ac47a228ee86142c162053750787741cbeb79555f00c278f650269e4c6c0083056cf5543a
zdfaef2d42e43ab92dfd69c5b51c4b0e58bc1d2486819870090ba715bab2c58b34c054425d2c634
z20b1c237b062b315a46105ff82747a61cf5208af6075fa0ea98cd02235cf0406db07758d09d849
z22a017a85d11ccb095a90dce9a7077d03f126d3ba02159dd169d3075c9de9bd5740c14481575a5
z7765e689909e6a592be3c08cfa68bd620716b0515560bd15795a57065a7d00072dd09b459bbed9
zb10d9524dd9f736c935d890d490ae099d1bb8a17ce07998676827772b63193e5de18e491bf477c
z20e49f52a7f11edecb662362e711c63c33a8de732637d95fb21f48a147b70f5c2a703725e39d51
za3055da2076e4f599ca1bea49503f9246964cc6ca03d231d52aeade0e9677c1ffd9ec44ea35c0d
zdc62baad09470bcb968cad60d4d2f75f43a869e6dcbec664c883f8c7caee2ab98f37e7aad6b0cc
z766366eb785b10d335d4f6708c9290d87431a94c0fe0aba7e6e060144629a48edfeee8a8ec61cc
z345f9518ad9bc104e69b855933ebd158f3a0ca3f853794e0bf812e91ec7bdda82cd115cc73a7e5
zdaa54d26108503239676b1560df13f2d2e23b0812009f6e4e41fb01996976858b3fb22d1bdc643
zb0c5dcfc02af5c4ed4f6e1fb73aa0756e903474f9c0f16144cd93300b6124c370ab9ae687476b5
zbba290ca67001b4227d317f8602b6d8f5f2dc9663a044fbeddb671d958fc163cbb06944dcc7154
z7a475138e8d8f088bcdc3f004e4bc54eef577bb619551a26e4798fa48434d0648ef02dacde9f25
zc8d47007d86bce336d9bba89ee0e7e824d0fe6d4839524fdcfac8b202e06b39ceb8846f85ed10e
z6f02ac764b6f679835f9d6f5703e605d9cab8478daf62dd399a63c2ddfdc81fb1190624d6e0d18
z7feb987bee3a74140342ccd427db2ea11a3c59e581773306f26428e4bbc14364f34694df6571e9
za031a2db17fa73c1bcfde342534692c96a6c6b0c2c0e966245662c471ec136ea71707c670ed3ec
zae0c654b75395fa25aefe7ffdb2e90981b51e50506e8524121c737ec02b171020eeb93a0772eab
z2c10e35525aafdcd14c72d282c2b95f69dcd6363efaf7d60805819b60bca930356cbfa39b7adae
zc14d24e7f0eec205580ef6586235dcf9d6a4053477728436e12ee27cf01e010f08d434a7eb8b9d
z0f9a017a1e711f1b5df82448580e0f05ff0589fd5d19403e837966464cd5ebc4d029c93b7829e5
z906495e2d04d87e7df64cb2f81622e959dc21f63df1b7c177e4acd24be6f2785bdc9c0237b182d
z7d91984b79a4f00621fcd48180daf064e8ece686799446c3289968c989458b968e2f14f485cc3f
z8afe603a9765973b58435c36e995ceb3f6a5f2dc6c680d7d6a859ac05c79e7320c00bc83fd5a16
ze70ea60bbaca28088f5503c7301a542cf43c0f95317c36fb4e78c017cfd9696784e47ea4a7bc66
z0f324ad6fb86f50389c3bd1c27c0da8b6221c09869b1c4084e509b8444d2a77f4aa1b1afb03c0b
z2ae4fc035224a4caf237799cbc8ca49d85d35511b7823a6bddc3773ca1ece1bdb83bb0d22a65bc
zfcb1e097d886e40240a8401a459c9b27d12a249f407db9c49df6a678d65c74f591ab56ea2fe03a
z37a356072eb5a25b42e640c9670f271a7233b1ea2f8e6a3e0067460c5a3b415078432a4d2df695
z529b7ae805bd029c4c85c0991e2dd04e1a6643cd388309fc109010cb9f7255791834bdd1a0610b
z2ae1783169c166464a4b91c97fe7cb944674cd2b40963e98aa4fd6b6a603bb919f82b88f5259f5
z95194d1bdc44147632bd0442d3b5eee08acbb23a4b6d1ab072832150f9bc56f09008bca1269b75
za2abb211e14a2dccc9b2e7736c921b6475fa14f2d513232aa8033d3eef0f033f4ea6c3b3718eba
z52f64c4039000bb29a7ae34a31f16d8d06599a55d8b6c8703d61ca42de8b4731a823829f2e125b
z39158e724f21878290f1aa3603006d043a5a306c911169751eead257493713bf7ac18b95dad887
z9e29b5c14e38158e8baaa23fda41eb01f6d1914e6554f9e33181c375a37147daccbe6c8d5f6369
z82363262230699d02d7a707c112eb67c43cd3fe3983230d5a39abd2dca43d324703085d688feab
z221fba9729685b5970d423f8bbec2c31c5fb47d1804ae25d93be7b067f4b2a8616ee14c135db3d
ze421b1609342488719abbaebb9e4b58c6c433a888d83a81bdb637a04fe6106b20975e9fd6edf3c
zfaf4c9af3afbbb83a12570dd298966ca2cdd534a2ec3c3125c38dc79187dc09e2b4ae49be90626
z249c27415c6404bf8ed127985af7071e9f9646c7425cc26568e79f17583de4c38462a2fa405266
zb5bc1b3de31bd311a365f2e9201108a2689b2428951f81b7f4c674a450437f4c247157917bf4a1
zb8b22ff6869045e321102216722639726fc119934383a5c845fcf7f7bdd7d5b24a99ed29ce76a9
z15c98473294d147a94960763df566efa5d8d259d20d8f63a5c1aa2c46abc20a4ae820c60cdb2ab
z5129706649b86e78109c959044d9d1b67799d97a0b3f03b6c30428765feb27de29cb760b83309c
z517bff9dbbc7f1b3244e8dfa087e1d0373c2790ed12dcf426c42c1560890ac08b88dc964c12c4c
ze30cc89d67e45d34bc2ffcf62320ff5c3b8a5f8004f3d5b8dbc4b78ddbddaf15103f7d348162ca
zf673b99cb754daec01524ad0b34acef214f74776d8bb91ba8608fead69779cf77b51a3cb50d7dd
z691baf20dce7403eb56d1a1f9edca076543164344465012cc376d568d34daa40914d90f1d816de
z623b51e62fa7897d45bb82cf14a98def6443ed9d1b6a712c2e6a32f71b8358440968469196a6e5
z5a9913bf8c914b4776a8c59d300046a91d6ea88cc5982bd8ce14c71aef96083ebd456597e52a09
z70efcc8c8bc2e741dd0f4353119a4588802ddcdce57e0a3b5436d8c166890d015e36dfc56f4d9d
zfd119f2b2aad5b16af52f0f4af5d4a3755a081222966a7762a0ba64b3d77dc52deabe3cfc15319
z22bd9478c35e639748f104dbaa2d86e44e4b2a93e8da62e163bf83daa54cf2747c7c5859e8d11f
z310255130b661c0d10ca62b4e010cabf272a1ce570fac68b3ef02b87be55fd931354bbd532ef9c
zd252f873e29de5cf21df779312a1f71c0ec1ece67131ec7f35389b990a8cb3eabad2273d90c4d7
z6139a4ad1284b03ecb6badd784a5d03e679add5706b00e98437255228f613a402a20b3e2fefd42
zd17abc0a8af902bc5a4cc3ae45bb0968a775147a34bb77224c1a7adacda6e4e6ae575130168b39
z9595ec607cfa620c07db6e552ae17bf186d1be56ead0d87afe48737755fcb6095573c052dc9f0c
z0a696db7d022ae87e2616ad6614627c437ed7e9f9ed8cff8c9384bb4e4bc1e8384b74d08490c1b
z9a0e2859b22885b06255a2b076837c2fcb4d81067a711b2c1120f09486bb98c7c593b3c8c97db0
z9c74006cb4554dc007bda8bba40efff31403957b7d6b0daf764e1cbfbd819465c7444c3f20edc5
zecaee93d2a635ff8b35d176fc3f2164967186d55d513116ceb23bfaf7cd5096be3558d91ac88a3
z23fdf706e531bd3fa3d11754e4f1fc08caed652200984d81b6df06f4f4961e9d0ed6df045bf1b3
zdd44c43e81053420ec0ff4b2bfcfbdeccf7314d5d8239531e00cdf5de4f68ca826c9c86da51e7b
z2d456f1203c440763302e745df4b81c51f6e6a49aa6eb1826f574a27e133d69cd0c974086fe0d5
z0f69627a195078d0e985931d9648df13a0f274008d14924d191bef5931a40a6e97639fb2a6fd2c
zd1ce21f6147ca9bd93777b18b98af303e1fb09fd5ef149662140d66057149d7040f9c4b52e3280
zf41ce98750e8d0b9e374b8815b4d0960c08536bc41fe2f081502c359b79df7068cae7511688414
z8712aad5b13b2720b87a4966d074eb65b5292418166ef86056af52989a659ef91aec5c66595182
zae01749c67daac7b344dac5229b987389c34745f6c9de955c8669a46f8ef7e1758a45f0bc8b051
z55949ef2caaae0f4860ea071a1362ac150df689fd37643990b68f063fddc22ef0b5c9faefa7721
z3f9f13bb657b7b96b2aaaff7869db797742cf9940c6f2fd131c5c32e2d41a503a216c33a38dd39
za72fd9f9d99006df0e1365c6c1d9eb233e032ba1cb433f48602d79d6ee8dd1d045768ef04f36fc
z0cb011d3f16aa820c55bb0c981ff27e582b9e6710c1ee1d8522640597ae87bda2dba3f84d31149
z1eb4a8f0dd9c65043e4d46e1fb4e319cb250cc07381cd3cecf4ee6513b0e580dea04231807aab1
z826e84d49c2f334903ece4ee3cb148c52e822f2636c2bdd44efcd446f69d665b652fe018e8fd2b
za34e29edbe7cb6ab66b864bb9b39066bfeac56887cca7a1f83355c403d14935d3943bfa0ae7beb
zc40cd385171f284e73f3a7bf31b758fc6d98471836fdde9624e7c87c2af86486223e615c3257b2
z9e8d303062e022dc2605cf773edc49b5074beb93e985a5a94c11f974f75a4caab5e16b45391893
zfd19842a68596319533087c47689dc7ece3e1870c35ad06de979b71b5d62a3c49cdff7604d47ae
z7b1ba093493fcdaaefae9bd7806d68de9a9a453cb85cffe30bf6e122b67b7b93f2e75fdae01e7a
z1072702334acc097a51928cdbdfe08a8224009c77ea1d618e1fa987553cf83cd68ec3936504e35
z2e9057e3079c5de06d7ba4c0b2db5d2daefcc2dc3db1fa66dac90a2ee5259092ed5f6cef512714
z16e80f0d74c3ee11a043c5c64f0252dd06b77fa9d73a161b006b6b76ae12759242087ca5a688a1
zb5acb5a802cd7d138aae40d8aafb3b740b2bd8f3de3cf8e2c5c3c4b96d0475db15077b64c4a1f5
zfacfc76555ea0f03b2e3654e9ba7815dbdec5d88f1a2bae390c5b34497df6bf2895b56222aa3ff
z6f7d36f5ad766de37539703561e25ed6b39d8cf91df00ded86500cec8813586ce4c33399e00cac
zd1a8a28177748f6900f3db7488e51a6b5cc2e7b20d2c773bad7ccffb2759c8715b461307fa3ae4
z370161507f8c63ed99de6f6cfa217bfb6c2e7267496201e455515a194f18cd06550af3bee3bb80
z7505024431edb31ed0df491f422c50a4179aeabed1c1316bdc742313a7966a9d49fd34c6519ce5
z46ddd5d2c8906e41e5b9d59fcae32839a2db247921e20cfd771e34b8783a127e37ed80cafe2fb1
zfc97fb93ff374987219c55bd9489eff444f70a46424ff6b36e96f92a813806b1cea730caee2977
z359c47cd3c5cd92c0b7641965cbb0d41eb925d533db7f5ccca2ef3cac0d8011a1706a9f98346d4
zb18079fdcbaca0d921b34ecfdb34030cfc659231883c68da617c0cff881fc7d2ac92a294062848
z9bce0fe03491708bd5e27b5d9034fb9e0b630202572616e5b48d5aae8a8d7fa4aef13797458d66
zdd5f83b7c79e616bce7ab040ec9ba99a2d0dd0248ab3add1f4b9329d250e6ddf2c93345ba89b93
z771e6cfec5aa4dcfc7cbd57f38db76eaf5ea14a62ba4085b3f52c57019fe5c494197b74f50ee13
z5eceb5dc0e31610ab97aba9918bd5874eaecc5d4ac342cc428ca78588fbd2066a4152aa5cc6b33
zc33b019a5f11c66c84fa412cda9473575728002d1ca33d4fbcdf7a78a44d998c18da25082af3af
z151203c9ef630c17e63cbd39cf55c4b01a07f8723e35a0e93bbf7a564a8748383ef53d1276d1f3
z7c03d38fcbcafd45cb88c54c806503658d898871bb9129506d69e78b2fc37eb700d9e427a86c52
z54b9d3ebd41845f32d73c906b3e8218054a447c4d60037bb0132e12c0d6ce6e9f372fb740f6e21
z3f0ba5ee4fd3c279897a8f4f79591c6d463b0a2d1bcc9d8ed1f69da550a7e2c890e4d452c372ad
z397ccb49975683c9b2b6d7c8ce2e08fba107fb2fb2de3da4fb14aac855c004b7077302971a358d
zd496e6c051e7fb88f1220809d5876eb352896fdf7718c4bce4e8cb7242c8238485987f489f43e4
z68c88d1083233e09ab1ad3837cb41b696f25799369b5f597da22e5c88292f6d813a3d4236fd592
zc4a4be12f0c0b667882b355b9e04a28dc75a21603836aada60718dd37a205b25e1c63d6891af9f
zdf6d8b7cc0e1ed2cef45c955243ab0e9cfc8c52a4e7b1f41ab36cc58635694d464bdfd9ad226df
z64fcb25814afc03521c55ae9b33ffd5cf2e81ec0b698b850d0763108c11de1a3005c54357ec2c0
ze19b11be7202606fe3dccbed6eb9263112c3f003f338b059c57a957f572f0fc5b3e37674b409e2
z6f5084cd5107dde8d480b740c4862d2311765e09000d9216503357fe32e33924722cd81aa309ca
zf94a2f7048d6e2e50892f9b74632eef03803bb97827be58b0811fded1a7829847601c8cbfa8725
z4863b17dc93cfe7d5ac71c0d1a07f07ea67be591ef29be82aef14af90752bf3a63747a3962b6b4
z490b96caf89f859bc105d51c7779d93db22de75210a3e3c42cd6b0c3879c1cae6c1e57015d0d23
z3826da018f09276f2c4d9c56402595432bc90b2b58a21b74bc9e91118c21ccf9d09d27222dccee
z6143a1ff87e418ae6e13b50cac9e36fb8b82415e24c4217868852ca4abcbeea035d23751ff9d51
za75e3096fc28ebc14c074d844350ccc4bc29965c6074fe0dfdde2d90b11ce9cdb3c025f45b05ab
zc8038f8e96c8097d000ceabe917d73e5b4490713ee9dcc72aea92ebb43f751f9b94293a57c2def
z0192ee44289154a2f3df0475984b01f6cd65bc579d3244fe06ec3e69c368747872f78ac7f79958
zf4c647ce18a731530427fe409c965fc7463aa4b8572ced96298f79b6c5de890bc360f4489712a9
ze3eb401979e07d63e2eb0f071e72933db480369a80ad8f03f540af76217176ccac41b2048ba122
z0283d4f6e0a59a66954d49ee356367a41cc7f34b7e3191fed10cadfcd046d7f04fc4657a063c28
z5a09069f06c902b91e4993d0fad02254b54cecdb006f643d193c4e4042e24f88a4cc3c94d4990d
z2594d9614c9b49a4f95c8a2d0b6da006b8e4034f1e96502d6f3eb3b654cbc99b1d1c3c74a916ab
z4b781b5c2803251a44213c421a4a16ce10f8c5902e31f440abd380c3fe7ac25934c5a0b66721e7
zbe173883ccba0f9583ef63c808bc2ae66379fcaacc7e602a3e11266204fb947af5228956e9ad6d
z4a2685b6b081f39ba8aa3f574bcd5dd80fc44d23dd7452302082823f3156140cb6d94e3452d8f5
z4c744cbaa30148a35d4550105f5750b457a41c17f8d645b74c7e75fccf303b6512cb1be9215de0
z5b983da1b528f5ff17552ff847d32363cd58e421d526218431bc510d289e81969932a44504213d
z3abec7a7b21e609c7762e01d98ec6a966fb4439414910a5d44c51f9d164d44a15cd7c4879fee1a
z5e645fc581c6a4c50f84ba2796bc1bfc653845b7d4a2f2eff107544bda326191355a7bac8a58dd
zf4d54715ac2d59ed5368e63f946d832133ffa6458ac021528d2bf8150ef74cc94c38bf826f8451
z057756afe84ecc1b9fbf88ad75eb6c2ebd56491047e2154afc3a3d3608eef818a79aad060edf7e
z4dae62283bb48e09a44c2673279dee9eeb7d9d48a80975cfcf21fa37d40c1ead19b22497ab8a44
z5c34451a4e77736ca0112ce9355cec3d66c830d9afdc34b23e1e91a2eecc5a161fbc707d73aca9
zc221804b49c02861a7adf394db5124cbc86b0afcae8033536c60852a658fdc893c22fddccb743d
zc33518b971100876a4735c5dadcd236dafb72abbbaad383873ffb7a27e106a4f309a9554e4a1a2
zd747f12712034e586f12b9a9dcb5ef02e6f4c160378370474d3a263f0b97de86cce12281e8ed4a
z24a43f5b4d7a4e389934fd687619509409e4116bd7e35ff891f633583efc592d1cdc7a41fd3aa0
z3ef68874c4d3391d7254fed1316e4e9f4e3c292001972f3004bbb5a5ee3947a243472c82f58b2e
z0be8d166d88af6b5a4794698d4c9c615763064f20d04a9a80d363e317e46cda7d22dffc4b75201
z914fa48de1085eab3251f660c009d413f77b9bc0cce7de51767241f0ffc7e3b77edbca94b46dbc
z08ed4d9c77eed4767c536bb6cb9a125b34b76ee533a7d437ac7fe0994bcd2926124b57d3cd652a
z0f9aa4e42c49fee4606ebb6f97ac94af9db2ad32c847caa8b2bb0f3e8fa7227cebf451ff88e022
ze171b5442a9bc28eddbe8265148acfbead6200a97e61567035cf92ee46ce080391e193a7d37adb
z2a9a820578e0d1b6419972d392a85387a242302dccf2d8228b958e57fd05a8077c73188c1653a4
z6b85a2e377d0339449bb50d7d7dbb365647c0f0b8ee72ff509db994517d8783625b51ddbb965d4
z27a2c06b7aa705401b4edc9558e63afa52efebb44e1796d44c1f856b0d8b543646d092844aca4a
z3fb1863f566ef05393e8bee5552c4a0af93116f5cca0b1160175cf4d8ee145622eaaa41bf655ae
z20c0e9b04fc1a11693d5fe0e4ed6655d2d67cc33ab21aeda99f3870c3aeaf9395d1519389493c3
zd523ff15fb5e7a6e3daa164a0c05f901624f27a5d9a693b5bae829fdb75b7be0ef3f75d6174411
z9a6a33c9c09877ceaa59f414332e45ce9fc448ebf5f6665500c0ddd6679727f6cf13cb1ddcbd12
z6354a4ade18b724f9d71827ff266db6ea9e652e969a84ee42526b9ea701aaa51ef981e5210a997
zf689f66680cf38a207f53b0725547abe4a6d1259a39c2c4095ab2e16169b16cd6b7e1237b531d2
z7888bf34b96447e36c18726d4e7c40f5915767806c8767b4730080e463da2e79d8eab79a287ac6
z1f4a918e4e2ce710dbf850f8221c7c31a44f564596da922ca2f14ad4c39ccbce4f0ec8fed685df
z346b412f7d4b9f15d0cd6ac88e519cbe93da7aaa4e2607642286c37803636ef80cd571689f79df
z4a0c4f65365ba8f0166525e671b765d275a6efc9adfbf176ec8c48a69e1c865dc6beb3f237662e
z1ecc3606c287d27ae8c76da243a3567788d09b6951d0e8a3dbea8d39f0a5277997c4464e8a7ee1
zfa81ea698537045881d0818a8a9d8a157918bd3fef6afb4622379420666a4d54322761767bcdff
zd2db83b32de0f2307792fc7abab8a157e4125159b155c0b6fa7169ca5f05aada6be485bc4ebe51
zd1ae040b5da0c34b65715e70a6c5e7797b0263c1b6a2019c0af315381f08e33ca1de9a4af770f5
zdadc231cfad5ec8b345ec270743941ec1a432f07bc86d4f95f6425fb51f632ddc214800291e4e8
zb75bd5087c0819eee5439982c2da9b2affbf5118ee25c0acf943ccdbb5face5a7896108e8bb282
zfbae2d2c671ba8ce82fc4dbf4c9220c9a9f16fa4c21f178ba0b6f752a73171d4312d331a4258f9
z4ada68b87f7bae498255a729935f1361adc17d3bd2cdd28344989cd2b952d946fbd1d828ff912e
zf81d4e7aa5b16532888ebce6263f66116c3023a1286ffbbc7b4e2ae2ba82c72232ba41ce6aea30
z89cb32f93ef3f40b1a1d31f54d873eee4eab284f50cd890ce386ebc25c8b2457b4efb0dfb7399c
z542b5b0b131c3c9f5daad5c32cf9b1f7eed4d3e12b0bba59318914cb658d1a3c9eb24624328955
zb6e025e497c51986918e50a0110dd6119705f38e3467baf5174060f0466e3c82a28b1a6b8b812f
z09730c4296f8fc391099a4221e5310b5e05795c75b66d6487f76ebec09a97bc45840a5b9312e7d
z413d989223c6adc6d553370520b2d630ce426de83c06bd495350ad2bef42e24e5ef03e6f3ba6a2
zbaca3d7b07f8877ccd7485557869135a70e35407c566712c8daa13bfee9d55988b1b48eb968152
z099dcbdcdfa6b9ab8555a72a03b714814fe5b48f5301428d34d8735343a9cbd66dfa905ecb5213
z745dd9a9a9e17062583eca4319df9c497a82fe02614e5d4f9f64ceae05e4d9da9841c3e4d1deb1
z3cf83c868ea68660933eecbaebcb89de5436c8b4af0320badfb8431d2d6d5323ab90791bc1aa0d
z6572a64c375c6c91ed3eab05e4d14fa77d24eb8bd4500b1313957416b9dc6eb935014c1d6b6f94
z00043113dc1e5bd3224ead2f8db419450112cad97d260261fb364c4acefac5d568685b94c1ff76
za813655f209e70649cfa6a0fbf5cb1ca7681494f4b2fa95ad7f2549e3e1f41fea69dcafe82a0b3
zc240436ea50f468d83284f8e3b045d5c23d14ef061c65bbd0ae7c704b1ae2e16c956279e4feeae
zd7d19786aa6b6ab1769214d9163477bc6fe5fd09574eb49be14af5a7c376cb58100d1f0360465b
zf8e8d6e566a883c8c1c2ba3bc3f25befca54dd4b5cb6e9c2db6b135238ca62e8a50bd68300db46
zbe42a8c86eaadaabaac53caf413358598437bb9a2e93d28464975800ab07c5fc826782d3996435
z22664a9d49e7afcdebe14ffc3470b4bfff3a02b7b4f9720797c39153c82fd0fb09dd99a142a57b
za91227fac52835b245ecb4942d1597d0094c4106d007b8964450f0f2a7775be3111646173a3fbc
z9d07d0717bebc3952bc38e16d7d7cec8a1b0a6bfad32c4c8aef299e4113617e16465e0667539c2
z316776b0c6085a99555ae5b2a273f36f0328bbacbfeed994d833bb65e67e28c702ab5528a0ad3a
z919f99fb2cac392c70fb073ddcdd376776b04bb3ed4e7a32412fb500e7f68ba1de84e0cee9a25b
ze74055c3983817c25c8e99329566db20a12b820a5b3de07978caa472b6c648336bd6240a1d4073
zf32b8123a1379702d7fa7397c1a890d70b71a5f37482b6f00d2b5b9af1175b99fe7d363b51d7bb
z878a0e31dc88bdace030c3c44ad0f53f07b176f5b584782832725f92bd5a252dac389fd882fdcb
z35b73aecf3400c92a8935ca9491f734f4c436056348ae309819a7b1add08537cda8177eea3428a
z70ade7e52fd6dea75bae1ce7af6290d9713265e8d75a674f0d1978b7f96614fb55cdac2f0234ab
zc291ed665c805b7fb165ab43ee395664f0a6bc78e11cf29b902714aebb66fdc56bf6aa70db7022
z4f79d1c961f85febf679fb87ba71cc226fc2a3291bc97be0c696045a6a77704c92d66f2264a207
z2e89d05c70e387cb4995fc889d015d44531d47085811da829c016c8c72c5750bb8f94d11d1c61c
z5be0edb356e601ca37b9b56eaa98de0077bd2c6f0ea351e67d350b929300a3fc98f9d0f099b0dc
z0f6e39ffc78d21056ce569b126d4c63c2da8d39e8a91d8a07aa3a5921062ed77187f8d9c85c68d
z148a9d9663e82445951fe7be137598b41f0c00c7424b2b3c6b930b5f07f2fad818ce8d2c00593f
z16f0ccf5b8094b9a56c0ff4315896fa6e721591f86ac21fa52b29f15a179e85c4ef23d64b54f7a
z500dd954a628946a327ff19d5212084c2226e4733452ada7ea0d6f63e32d23e18a7b4320e676ca
zb7d77655802908eec85d55973d87120cc1a771baf4e1c929b3a105e43c0111f02bd1a074f36b58
z97bf27df3cbba08237c1cdfc22b9ae9645859f3e338e2db53176569b7338c4a0ab62eb90efadf6
za32929c190d9eb772dd431a1ef3be8ddb8ccc1314bbd89e797273b17cb7f4cb49d76d7ef2858fd
zb6ccb267fd28fa1382df2a3974e7936155a629857fe3dae1da6eea6aae33e47d7c36e34effe8c7
z6ec0ae4fd9d99fbee2c1e4ecf03a80ad4f7f2e8bf452bfaeaa084624edcd602d4f7e1b3b170e1f
z8319c91e044ba33e366b5a468caeaa3a22b839124e82f702843704c47f0826c4fb9c715cd25297
z5abb98e6063e32d2ee14d974c66c95b1c84db6ad1fd907ffaa6464a3938118dbc9e29c5b8bb9ee
z227d4750284ebfd06419ad071318b1238c796dc4cae953b39d0760d2f5dde889d2802ffcd4eac2
z22c2099df6260192d564b6b5018321f5def9fce1682919f5de3a7b53c8058f532fe1e72a0a4184
z649ca82b1fde20ef73de310493d4a53550f84e0fda4b6edd0044c4c11142ea3a52f83d4d2f10fb
z58e2143755091b80ba4b0f576f8fc2a4a5ece500c3d2212ac91775c3eee8c53bfe7d80f1772130
z9e3075f532527307be9b279ec341f50d0ca38374a851671fd67b7bd54149a6555baca766cfa527
zcf7f56f5fc45b7900619f1c2afd338e4fe09af489bcc39b3a6d2acabc209e54d6ac653760c3873
z7c1164c17acf40115c898f72d3975b5d45afdd441f1017238b6da8927ab9cf2e020d5d63ec9648
z306229d31d3a71918632c6abd259d53d02b8b2eaf97031b67c3aba969a6fb16b6dc5e922bf8b6f
zb24173c6dc54660812fe2420c7374860d3d743c6ffac6f26311226bbb2a06d921b587a4d5af6fb
z6dfc45a127fe1e0795ab3fc781d0b6a1a3acf9047fc44045460021620cefbddb746b767960b07c
z764bc9ad259d3e1925159aef9787f801218ab4ea24eb6668678d947c33a30ff7807f855ab38109
z5a32988a16b5501c0bed36e8ad7879239cefe78c0912a2ff8a9aa59f0250b32e48591a8611dffa
z100dacea41bb3922813522a7afd27ef4ec9d51a10c07684bee9a815135bd3bc44dfbaa9cbf6ede
za680203eb0fc272e70e74e42ae01609996df7507ffdfe209ef189c55e788cfe2ee8fcb479c8cc8
z7c43be25047c3283156a2483091d3e745464f1b39038dc4989f1fd5eef8fdf3cd7e9ed4b5328f2
z45010cb4424b46e01e78b72286c2f6d1dc88db55fc2468d84ae2aee14e0770ea2414679b9a1d01
zfd727bba2cac0fb50c948259d1824cb5bbc1ead6ca52abf88c6dffd1a0e03259ca35b4fa6f8c6b
zba21b917571be14eb97a6ce21b580748fef008b08e33442e80b21d729230fa48ae5470c3ef53e3
ze71bd4b8ac78a3c088030a1bf8c06795eafcc35f34c3a6b49576fcccdeaab80e5cc84d9efa2598
z51328b30db357c0a4b4fe2b596280450fd4bccd9d36cc333d936ed78139a0451a7ce2dcce5a062
z1f59f555d51cc416ee6f676b3ef47de007e091573615d5da8a639630c62238ed68dfd12cab0097
z428903082dadc9d2e9e08627bdd1bef21d78219638916750a085f8160799005416fdd51d5c7d17
zd39ee3d5d20b5062b11f7fd835279d3ce834b8f2f0f3860dc01ef36431f241a216bf28f7b2e0b5
z6a022e64506cbb4055e6ab0c04830c18e28b86f7c24795488fbfd2ca523836ff58afd7a3b1c4a6
z850e3b1ae91ab528775259b8f469cec879366847a3988ac0c994d0eba22a652bd1830b2e1dcf36
z1bb1d182f314c2d5f4a702e47b7960e7fbb3868ea7d86bd856f8f50e014c8e8e4414f522fe32f7
z04e16c33dbdd6ebd32df1ed8106f8bb57a91f3176122760cd337ae4f032c7b1f375e44e5997324
z1c266f545dbf74923727dcf5d40709e939159cce808cf78b86c8e48f951ef38783b1dbb7b60334
z4f5b0d37ca6af5ec2b853be582359c9b47ac48c08e72c09006805b6e71fefee2c8503701019f8f
zb8364c59a043dd67c30207ca47b90148ab3efd9b09474d1b7a049977511f677e23d88d89c4f47d
z5e297e17891a030bd0b995a22533ce8e16880e4caf31647f4216f136dd772d13cbcd19a8d87123
zeeed0c07f9ab458e4c32a3b255c6b3c592ba3ea290a92f9a2dcf6231e9442e1b393cfe60cc7b8a
z2d10d53b45883c870a3f631c879dbd4d40ebec62a063d919e8932e262033eb8a47be90ec889feb
z69b622161e91f19370e924f91ae52a0a2b072bfe3dd57876c3379b1ce1db15f48656183351fa9b
zac59b4066314d3c7513cdbd462a2fa2da096bbf7d8a18dd10a71be350205a9c0a0c06ce38f536d
z1cb75eba146366addf47aebdca8fed976a577a614ffc6ef754eef5473556d704571e31f01d5954
zb0056c8f5c2cc786fdf5a3b04997649bdb83e030d1e607d9a297730d7657d0a45b0c71d621530f
za82d5e1f2e2aefe0fd3ecb833159c032e0383eb11dbf17e5c9501144929abefe1a6a813200cfe5
ze43413a77ad09bf259e112619363347395af5862489e43eed6a9bb1bd50e0e86cfeae002ed30d0
ze15afdb79ef843412abe7e50fefb8ceab13fcbbd6c4051a02d843c13baf812c7b8a438734847cb
z80b4d74fe6e68f27bf1b0f93075779cf0ad2ad658c2a6e0e458657435371e8d00b99c106ad2339
zf89982421784c516ab7df81e81409dcbaf536a7f7385e4fa1e7ed7154ece372bccc8e65fd5681c
zd7296b691c3982de188e05548e5225b5f1204f399f6b262d722a9b06dd1dcb4478e6c567089309
zc4f91a7475a1d8302030829ac94510b244d5737e4c96cc28744e551eb58424ebb3bfc23afee849
za50833bdc9fe88bb6265f280a5162e35540e1714ecc654c4b88f76c294622647743ed802e5e8f8
zea9165727f6733283e48168c195ac354273138691927624872f3d1fb852c9c57ac05ec01cc5fc5
z64bd78d4084b620a2e49d3e302d9e1758dd9b9e2b96b7b6082a6af2dbd36aa548e9f367b446883
zd8f15959fe5339cffc1731978e749e2b2e82af0c75e8bf310f79406d31996b2629751560b042c9
zf7cb62eec3fefa0b73b378b2b392d7345557d0372580e472b2077723c67c7b06d73bc15598ee64
z2727f13041a2e5f1de152c3000bb30ece3edb8ced0d1514750ded2fe8bd01e61d6c4d405f387f3
z544fb9d1d85ddc63d4cb583d2c1d6a5c0fd6d17ca116012ec13d6d336701936ea67cb67a45566c
z4ef37dc416288b1eafcb15ea5a122f829edfef8143f37113472a495d571447d37366a660e513a9
z2355cbdcf4ac8dab90f961800785f8779c3214a0c4a0074956d58fb9f8ccf34b818282e33ed700
zc5c4cc43394c8720c0d920692d3e80cde275dea383945f5bf7576efc59920b7e7c9e9e351ea371
zd04e94bd6da4a769af4d151d952600cf3acc523096ff29ffe06229b56a9b80b3ee527350602281
z26299a6e3d6063c6b68eb31876d20bce45edb646092fa42499310817dfd309f4f694663258861d
z324f4af37a2c8f0449fb2e0f6ec87fa2f7e58f511cf345af0e8964f2f660e5a3c0c5c665b59517
z44f149e74bc27890e0fa1039523e5e241a30a044c723ae6ee6cfe6a0ebd0a5e0a8c09e7f1f55e1
zfc3ddcca51673870cf99430fd122262a98c899443544d5ef30c0da2d2ba59508f62b9ca300def6
zd4444ac6f29df4ccaad15ec62c1f121243e01dc30c1fe92dfb35b5444de8e9d71115664e8e9bbf
z395b7c02c161ae7676c6323786214f9e96732ac7e72ceeebda9d633380e61138af80eb835c705e
ze9946b04a027a35119c7f0436a5ead22f8df630c545ca3d6b25af3e099e4cfca1c191035fe43d4
zc3c39a33492a4e93428d0bb0c201a9e436bc20cecca92a6ce8d6e53e48662b946fc4d2bbb8be16
z3a358aecdaad0f5f99bd01800a807348c41fc07cada5886fb7b209844418c74565c07976de3d68
zcadc09f7ffe4cdb5467c0c61405ad5885b18714901963b1f4e61d85062ced65bf5532716d32df7
z5aa531f581cc40fa019291701d424520086fb81deb3709fa1efe0a42447178854c75b6976aa753
za17f152ef60e4303c170d3fa50c336d308281614b7f2ebf2475e873d2b3e33b32f05fcd4dbe4e3
zf0607348465daa0c12e2f0913f22aee558c7baa1ea08e864abff78c7c8c93b9218ada97f1bc2e8
z795054ac00b857c6a7fe09de8cde59933d10ce15088a9f71a7d361ec21adc6440a92af22f33dbe
zae68a52daa7a1b96f7869fb1cc644023b6dc5e78646fd7a52f3c39fdaffe20275a4678166d116b
z235108f0199b6d844440be4fee03793e82163c7f8a477fc69516c112dc852d4c7c802b1ad5086c
zc6f6f77f9be92688967f3a2f4e553ffed69b9675b59ff9877ddfd00a718246cba41d621ecda3d7
zc93da324978cf30f494c222113ce4b449b9b2bb1a2648fc4ef8b921deb7dd308c71a0c76d6b3df
z504185778c70e843d64855873b0eea024a5dd5d460ceb424bf088bdf4cea7a5e472dde2307998e
z2a1d21f671c23a0ac209636ed4677b709ab43b2d1bca9f2fb50d31a3f4e5e2f617cde89a770b6c
z2af7455e9c5a75e0d5ac723fb7340178441134bf13811005712ef3536b150c055f296aee8ef601
za3fb22f8ff8d354858284035f40f6925136b3fa7cc80b842f6002bc1a20216d91db5349a0ecd26
z9efce7f793a4ed870949c00e09883ee7d9abf3e1469e3b2cf8434c7252a83d4f14a8608fc28ec1
z035732b2f33f23a08b45a8be205789d054986556db37b3b96c8f9de807364f0657b840975972bc
z7773063e1eb9ad9b87eff3cf925190734b2f43726078b28dd4d486443979d11e527271477c5766
z0d583726227acc437014fe9df3acc660b9ca13b385bfea49bbfb61b619476a426f9769341d5963
zc9fc9b01e9ba97ea071dd511cc1e5da4ab68a733439c47244aa0d4dd06bea64b3ef75b29633896
z4410fee0c0c7f9ca6c3ce5c4724161d4846ab4887c2e197e8e15d011203ad1873db912be430ae5
z897f81a59cac764b572d6ed5de1e04d6a0c84969d0740ea5fd0567dcd37f3237aa2a0ce326cffa
z153a5800200a3524da683ff6cf4abd6897a68212e7df90cc8914cfa6a7f6b376bc317d0f026677
za63ba2c0b187c6f4a2b89dc8d2c95f73d6d0a1e01a10e0d64dec5ad1be7b20f62570eb0264da40
zcdc7272559f344ca00dc2a217c576938c32826d43dee6146009450bdaba47019b46e1789c0ccdc
z99112b6444b6ffa772092b1f30e5fa81c5f92093d4e3ae77332a8f8b39b5840cece4efd11c9e6c
z9e5d8499fb4a8ae8fee0904725318d627dd52b31315f009e38eb8aea667e9b7ca628a402202e6e
z42a4ca70ad26253db7e62d5dc9563b10ac4e5ad0dd8efb2f4dcfc712255dc5e1cdcfef317d3151
z301a83d8015f8c4572970a8dd53d6eb48511c7f231628c5b4591a70a07f7bed675ba3814c7a930
zd0b4e54d08cf54b24b09efafc6391bdff7286827053dc5c406ed8d520a86ed4fccf087030d167e
zcce893941fe32b809a30c93be74827faeb550f6c230c4fd028a04baa00867dcabb6d615d5fb999
z77643987f36d54368a4419e500ecb116505ac854ccd70b5b7bdb7697c79783664f09b301cf94eb
z18a489de64c56009acf28ad7a36efc157283b5cbfc8535fd19b6766b4ba14fa31c331afb88fd4e
z169205b59ea7ee1f0dde3b519e8badb08d94948c0e747e38f3c5c72314ba4b6f6cf63d44a3bbd8
zb56aaa75ca2b2368d56cd1d535246705ce51cb567ce36c81c311b066331941720026dd30e715f6
z3bf66d0a63fbc99330fe2f6eac531088651aaf1559cc44b1261c700efe735d7ed5456552062ddb
zdf749816ce67452396b539d0d3a5c9337efdbb7de67a46691699c7d430c94f2785eba61fb19fce
z6b0a451baa4e5a63264b8db2c9be3568e1687fe483ca61df116cfd21b0ab3866dd1c246d913bec
z88e7f4680c6caca5d5118490d9e9cce87260bb9bb6312bcea3b8bae601546df5b49efaef094b72
ze811b488b6aa35f3cf6ca7e7b251c7cc24e1ba77ed595d4649e34095feb2b9f2ba486e8bada43e
ze568c5753ad33ee00dda3723049ff622d474628d31c84adca1ac4d4d97a0a7f4368264f9240603
z2730eb10e2cf01f2fb22cbf57f2608a182370884aa64b5a53ddd533c5f30d09615792e749594c5
ze7497842996e23d97277fad53891803edc538ee1e4d56607ae19280cc8a0e8fdb0dcb186f33a2c
zb6f1af97a4dae67aac465739c65502fb5da2208cba9db48beb9e59248609b31e6f7dc320dbab2e
z29e5eb8947ef962990e1964edb18e096bc886ddfec06983e0ec11460fdeac953d16676d2faa564
z9587d997deb7b485a71c0678b6173197adf66ba5b2eaddcde630567dc29ff85f7cb5b7eee61082
zf360bfeb3b053541543414b05e7aa5f5c7566f00686dc1057aeca9f9a2a776bdfe37e3755320ca
z6334a2892d7e30166f982af4ff3551d3e8d6d09fc6a1ab7a7be82b13358ea84d9305055a7a8a79
z82858b57a3e1db083b37afdcaf413730e94e2db7d4f2027bb0471843335235f5c1fc0930da46c7
zb2a70da8690040dcba9d69421bf1f64fdd3fb5dff43d96281cb75ac171f7306db6355444d60026
zec1d5cd43f29dde5cceef0b845a38c8909c3eb8f03867e9af7b42e90e9b6c6b2c2ee108816971c
zf54b9f7fb35830b64519ef603be657fd4d06fe0946cf81bb36745b93ae7f2c36b678520ae14510
z0f077cc9697021b0e7b8006760c69efe73f1321391e9bdc518804554dbb569989210a39a4c5063
z304322e35fc39ceed847a8b2255b1ec54643d5d746ce0bd95e7cc9fee67b3b8c7f823ced5156cb
z115192477e46008c4bd37bec71b97226b61f2035bd1345c7559f2884cef63e3db291fa6ad07a1c
zbf1f41f302212afc4ddd24205c1a73e4a954bf727992dade3c6c784702c92b77742e651cee7582
z8920e7c9acd7177180234784b242c99bc848ff4516dc1813c049c7a7b8e2a6fc452f25529de89a
z2e6c840976870f47672d0c11dc51272b75262a1af17c62071283d80167ea1078f7a2a16009bd28
zc58385598a0eabce352308c01bbd87070135512a86a3fed71e4896f242f3a6f2e45e98cb295fa0
z736f3ceb92cab1a0e8a3345cccf97e8f0fc397559615012ec7a0a7410375a08e5b9b6e8957692d
z5cc4f0fad830e53db164d0b12243ebc7c64794d21c9a8b725b34500e91e53910bb1db925e0dc69
z213f4381a4e06471e8b125185abb0a41b66bf14497c9145be3f6348675c5330c61a0a45abc18b7
zf37c02e728314dd0807f1e6b552ec1b10291dbf6dbf71499587a789a5b39f9410bdfebd94d8d1a
z55389ba74e2d045b7de40d11f04f77dcb05976393656588b3bb79e13e48d48f6f79fa243d023c1
zdf8d9b51a86a6789daa6402ce81413c8fa4789fe41f80a8018fd1c87d1e547272013686b62e4f3
z748916881437ec88fe0e9a7b5b4488ab84a32ee8a6b814c6e2067c5c05ba9257a37890482e6e40
z92b7e7894e0b42fa930e3f6a01729a64b26221e8bb82a50664b04ad1db06edcfb343e13fd8cc48
z62142f56c7b01d459342dad62eae92a2d10862ac8f615619bbe3f266f0ba2c493c1c5b461f707c
za454133bfaaede26a1743efd8620b623914f8e5160dfc455020a5145ca627121cf40530ee10990
z0dbee30d0de725ee61b124c6d94b86b985ee57f4dc02a529ab012a24fd47c53ec8869fa8ff0f81
zd200111de15460b765adb90632ce33b6cfeea73adbefc00ca9de4cb0c210f85f41d5153a146263
ze838486422645dd9c88fd892d1a2d86a201c348c49f8296abcd5a96acf3bd782bd7743fe12a694
zf66c39386f4cfb03af5a7ca46c73a510ed09d78a1047caa37205d08826a3cc2c03b17862a9c39d
z11bc85fe910bea551940bbe714e7c8a40d97cf5438baf4416c32a5a6a57274309ae49688693947
ze15071fb45e91f98d240562f5f23abc1fb28ef4c63d2b0a8ccf3867a8111a2535b950c48144494
z2f8bf33deb0ff5b9ed669b4ef25fcb72d41bee5a07e412a16c725f534eaa177be54e7255b8bb14
z923fb5c92eed872b6dc9d983141c4d29391648905c0a96639470632408624c77c9e40c1a0af616
zd7ef1026725c294a82d9c20445b70e8f61b3eb70f83bda1204a40620b9af09fe89f8501185c60e
ze2e46ff69a66a0f47f67f249deeaab11104272fbcbf9ba4d1f94dc072391d587126edd463cb6b8
z17bf9a46dc806680d5dd30bd9c7b530280c26d984a367d405b2aeb22fbbc92b758e90defd18280
z51ec1a2045c55e04d57b6432c92da419b189431513a90e8e48411c8c92ba967e092b9955a7483d
z6f860cfbd8caf9e2a8c017ae44ae2c97ad7406104fbd105550affcc415e850f91bb3f7b9acac53
z12240c80882a793d338151a8def0e9ac8815b59e04c99d90af302f943147041d230e1aa6740e2d
z4afed5c49aa2e045adff71f651b8add110c21af81e344ac5a9704f6cba9832f0fe467ca11bfc77
z553a6e31a01538244c4b0a717ff6e8587a3ec2b747f9bd5ebdbc24112b8c1c6323159cc769083b
z0f18b2c8bdb2d7f45a81916673eec4d33156ad1b2120726d226efca13f2e6994f06e1be45979ed
z570b3003ade7189ed287392380b337f1799359359805b0951cf2c3451fa477ea43dfe6619ebbec
z7a85bd82d2663768d420875e6701687c3bf2f59f73e8c52b1dc3f8a62df4f27f31d3ebb026a1a5
z11ccb3a12f607496fb38e13ba6159ce31702752b4146f72626ad7a808e0f00fd28e326bf32c420
z1589ce498c47c2451903433adfda85451e85079153d4796dd8358049ebee012b5d981ea552f607
zc37c11e102d1416e6798faed442b4aeece1ec2512b04943c44fcef96267af2030ce1088b2ca8a8
z8d24b9a20a4be7d9011241109197032cb50bcb751acebc1f4c58f50e2fc09aad5674510fb47c31
z5e851c8650e09f138991d341f7a4313eb88142062e49a23beb940ff1b8320c97bf8cbac4eaf66e
z037f3abd71fc9541a311558cf1c00907accaec5ed82654a2dd764d9f36e1857a3161a857f79ba1
z47e8f5dc226553896158e325e05365d65b4427c4cc362859d4a57339e52baf5bfbe13ebb556675
zd9b16bcf2e325ccdbae46d6d93efcd5e051f1c3f59bcf92cf90dcf4fe7492d1d6f80dafcfb1e6d
zf58e2b35ebbc7b1c39987c701e3d564df52440c8b8744f375b79a5d618e6a1bd50cb98c2a6c54a
z6e4d0c3f4de0605f650c0b193e3869662809635f49e494eb770f0149e49b55cd81579ce5f28004
zb6430c42fbc386ee5aef0537a523cd31cf68986ff174ed4f8064e1e3771ddf03f3297f4be0120f
zafb2982837e3832afceb82d697b42ea37d333e6a94336322fa8802649409f6fa6d3d8f6c33e6ba
z15e893d81da1e789802acd8e4a87d52c2ef71950bc3c1175d3df77ca81a7be7d11e1010220b0be
z47324d6500112def88b9ce0b1720de8ede9423aacc10d07d6980c763f07add36d9a30bc67911b6
zee534db6847c2ba877f4e5493c215d4cc07eedff15e291ee5520bc3e02885ce56d2b9c19a4a628
z6624323c6ea136df5c8469b1a89e11e9408ab5c642055102d6b0b7bd0161295762ae58e637e9a1
zb5e83782b7dd58eb42c8d91415eea1512ca895821b7fed9faecf08916953a4b4ff5dec91053957
z5de197849792af4c47ee145d8b5b06d55cc4d434af3920800a89d2149bfb928582a03e57b9a567
zb6c01dc2c4462e5484925f87ebfd5f5f092df45e8227ff8df16f9d43fc3ecea10846edce795054
z2b5a55d54a1ea2fde36448a82d9cdf5f68c49af84d4b60e20e3e8ed35f27ddc99ad024839c4715
z5ca261144c099d5cc0914c9159e3a9b2b35c7f39baca2995164d8e94d8b146d95e355fe7d954ad
zd676c0ea63556e1f07fe98502afd145618c3c90067fc1ad353452eb6eb077c00950350c3332db9
za21a41db2f514d6a04dae4fa3178e3e8b07062e3427adf286f8b13260a921025865d101659578e
zc5337853a8e34b4b8d54b68b37f01b98fcafd3341c5816592b31bc1f9eeb0543ca759c161327e6
ze6adc56ef8d6f53907ed2cb2f380f6c2cf5cf1e2ac8adf2ebdaaa580073e08f8ad64c720826306
z83858a7899078bb9830a7cc0281f6e5761fee46dc9b71a952cd084e0e8358c262838200d8fd3f2
z693a4b0be069fe5481af663ba2832afdf5363bf41a20b1ddb49096c527347074c92640d2a3f9f2
ze3c0f9959554e9db9f4cd9b5be5f70b5a9a364919944f8453312a817050e24e6d4204f4c853a56
z52f3d52ee7850582fed0ea380b4abe235850645e713de06aaa38c89a1aa4984741017ca9381c6d
za0caa8e37d065b08922020a41f61bb66192c497c6fc86be1aab57ba55cf76eb53b4d1ae69bea51
z4cae5bf38b50aee4a786a9ee447cbbbaa1280982b90ca4e0d27e0b5807268f84b51dc252025d9e
z5fef64db9798e160be3a0067760308e890f24906679ce0ba4acd56f5207ea08de3a6cb35ea6bd3
za4bb5e78dcc7dbfc8dcff542772ddd5aecaaf9aede76a4cf85026b35fad26ceed5cdf7cb4a61d8
z88487a6b28c7bdff3330f472517b3d52f53c61ba52b11d97bc994c741de24052a9d7f8a49d5920
zeaef33542b7fa0b8b0a75f1efbbbf8c38b3057d7ddfcb6a9cc67ee26328535c39a5213c378be8c
z731dde076beea884bd642185af7dfa355008635dc72751e84258924e343c98677137b00dd9d214
z2ea14450f63fe8b8212e8ba595f73ae90ae17721508c4c200fb04bd9319527849a79703e67bc13
z1db301baf8b9d5bc9ee1b7788d88b06619dd8c07a408f33dbf98ce8e2e14fff61500339c16ca08
z364473728c23906cfca02fc8012cfa33848ffde941dae50a5c118b33b9cf3d9cfb5c4d814bc78f
z1a27192810081b6cb250eaee614e70af3b68913a11045dc6ece9d73ff5ee731397f95291645fea
z9355e51bdfcacd0b40b2d8638fa5e60901924a4dde59217ee54f17beac29877bb8a575d43ad09e
za8f6969d0983b328c6d57e13019239caf5aff95248669ebeef1cb160ab72b9e280cb381645652b
zcd1ada539bf10434e77c712780f406ddc2791c5a9443bb3b740e5c650250762dff9a828a727790
z897f1c3ee1c05f3397924defb596d30603bad0b3caaaa800f5ff10b5a498eeb147e653bdc6e188
z13c7bed98404947954e620d1f1d8b3ee666f5f3c3347d04ea0a690b6817fd72846d076e6f71e0d
z8b6b33e492ee261fce5730c2410eaa462a8f3cf141ebb4ef32a841ca304413c4656185f93f3baf
zc370d811cf614e1f0a9979633deaf125da03a70860a689a32ef1f4aa520495d62479f3fdb3b4fd
z999da706ee32da540035b9c02d7bd386de0483e7860c26bc2ecba76f48395100117b8d987b1f87
z3c8fae8a672df44a32ffd7ae3a4a3b3242b89712525ed4c4cbf9d9b8e9bf7242ea9200bcb7cd68
z65b8f516ef9875800e4762b79ec9b65c8efa0e726e682ec1c1958f82761ffa702917683fff92af
zbeceb53756f291961c0f1488bf2935af2314889c77c2d0c23317a4205dfd7df40ffedc0c392fb0
z230d8324d391ccd210170c85af715be79b1f54f83e274dcf6df3d8e2705e82fe213d4a3028be4a
z5487673b21a78bd10fec28737c1a4f20bb89b70e1785678242d43c41346e847c7ba103c3e5b057
z889ff690580b708cd1f547344e9779c737c912e266bf914ca5160cff7eed32b0080067772692c8
z9bac9c10fdea330947df23d8204c693182c61426c3ca2ccd79faadfa8aae91413b5f633afe863f
z4dc756aa818f724616d8117562c33f3e6c2ef677b1d9e73bd49e11201c9da092681fc35a680e34
z49d38eb5ae87d988ad9375be36acc0f0cce1d18398fbe223fcd157cbde8917e5ae480213cf27d2
z2e0e53aa312c0271880ba13d789e6e849b90cce0cac5acaf714871265f0cfd39d4028388e821fe
zb640bc9e0c33794cdded057282bedd64167f8334617a09e57c2bea4c08c2086d487249dfd2b73d
z341ca616482f0555d5abb5777cb0526685b37b80eec81ca8deb6ed464fb8b7b8712bd5ea19eb48
z05577f8de889a6978e4abbfd235d03ea9cd04fd6827318532ec108fe1168f40e80e4f9c66c4aea
z0c8f7a45b86ae1dc76b9b19100dffc529e7c21544d5f311799fe2f33b4e411bdb2d3410e0dc8c8
z8ef3af9c93328c9338eb43ac91f4c29c561b0e6b74d694a305edbe760a9749fcaede14efbc9b9e
z279795b9c35d5633520b5f1fc4a2fb3ba8191e3e6397fe743ab44e1d0b71969069ff8ba7b49cf3
z91967ae4625f797b44b3269e82d23a5ec1b412a50c5eaebfabc80094a48af12c0ad567941f70ab
z53441ca66764c858ea659718ef1aabc2344b5c4494764bb8020919a2828582194804c1db10a63d
z4a02ae125f3858966a959a8685a8df2add669bc862a60053b5659ba7e8ab5beb323b5f9d66ee1c
z8361570e5d45a73b153d5b79424c42d7064fe65458263929697746938f91f9b73adb5c38ab8726
z0e44c56390b6f9519607bd7974adeab37e82198fdc4ec9da1f715e34db07bb04fcc339affeed2c
z83470b6aa01121287c68f491618e372f7f9b3cece2c81cb58ec42bca0719f949ecfa8a10e3ae34
zd52ebdd6501c18428892f42b79f74cd9d99434fe0597accd558ae83176154da03485a4f652cbb2
z88ec731c823c1e9251b44b100f52954f69212182d2117f43e553c1e15f77b4b8ffdfcfd4018ad1
zf2ae7444735a6a633e313874f507bb2778ab298b71dba33d361f9f33b8158174e41e7da7e0d0cd
z64d2ab8fcddbf6ebf7a8b7dcd93b1db4c62fdb57e20eaae47b82d6d5488c904ad7b23104f279d7
z2c47d25bb428a78d27a39cb7dfaaa189f9f6a5cb99c31741ad8e32c7992460a7fc51221eb09714
zab07b62d52a573571d84f84de752ad019c0d7cb892de34d8dfece76e273bb8d10ef9780b91fde2
zc1d6ddd8cafa088ef7465635b2a5510931e3cec112b44c3c9efca24b202f9825d01fcd9fe7fb68
zc15e83bbd2c7f6c4c2c9c4cad571fe06f30c4d62e7bcfd85f1914d04736ae84e61609bc5d6526f
z3d9ef257f0ce1075f59b142771e5a2cc61f23d7dd148b6cf7c11d9a6781555c3881356ad15b718
z51fe84e20a87485d032eb573e8f73c7cc77209b4ae79d5adfa07c3c558c88a328eb30da1dc25b4
z4b4caf8cb2810190dadbf8f51deac9f6c173d0c6c277b173ed44f799a0d7805f359bf9a9453400
za30c4e07ba7e6a5f3539c77131284e922f3a7a8ed9379736a1d0b140e25b1941c28be6d5637eb8
z6879719acdf12749f077f76afe26e495abfa535a85ee793989a3525e285c3e4c8fb94949a272c6
z8b365fdcf500f462bbeac2be8071c4db3f5aef07c6564e040b59878a20cb64ff198f09419db1fd
zd7cf14431de115e051d55ba7d4ac374dc7ac2683eea45ffe3e76f103299a7c540064480fcc8907
zb7a2f63e63c794bc872c467f9b661e16ce967696ffc54f435f5fa1f81f2d2475f631b4b0e234e9
z1dafce0e4d8ebd17a7e299c3d2e125e3ce58dc02af0f3452f594ace6b947a943af0ec22f1a4979
z7e5e1de8b5cb223a889c9a67876515082f062806ad7db7939962a79cb3e18707610b8ff278b232
z871bb5dd9a77c5a7fd8d75bad12e81eae659713d533545ba2498721deda9fbee29aedf3caf65f4
z9ed5c899f961d2256e9e1ec5c5ac0c582b7252698f35887c764d3dd8f93ae441755e24b5cf012f
z0bc17288cdfb0a56e8773ce6de92e287404b034bac7b2ca18b2079eb8d2719dc2bba30414f7c42
zc99d48b96cbb813d63bb1374cd62a432f972bf69471a66f509ab7f25d6fbc5d2da091d22fc8d29
z29b20a3eb98ffac4f59aa6ce58800432b90cd9be3c85dbbd13d1881749913b0954a28512e26b8c
z0a372b43cd8f18347f6f110f1b43eb599dfa2eb52e61d7a652f31a7bad42dd9e5a4c166cbec3c8
z117d34acb82c4e38cf1f925e36d7dc216a602a87da40ebb7fcaf9a797a91475a8d1ed444e13084
z519075f60b5b0b1adbaaff659b7337e893c08a446862a9d8b7b9550330e8dace5688eec1a69bd9
za07061db76f11a2ba78bd31fec0e2e81b472bddc6b819a722ff4742e7bcb85066394e4bc5a436a
z4142ec1a527ca9083d8158f017f6b5ce8e630dd63766fd3425e6eaeff733bcb8072a9b6c8cd6e7
z8a3d1621c64aac8d3ecbe1ae885d3dcbcd1873cf159a544fe9a121a6c12ab8e2cb86e333fde0c0
z0d6de3dea6f0dd4622c03b3cecdbc1b4772922f82331a66dea507c74f41d1321cfdd1a22f7a738
z81f6bc8327fe0515386fc044be27452a1f63ec1322734b12e44ffcf34e53dbf18d18d2a346edd5
zfbdbff80dff6aa4949cf73077b6066d2c6ab45df514b5d6008b4ab56bf5def1c10049e4be7c653
z2c5ee4aef01363e1a2c535e8d325e727750c7e4679d7fc009e5106abfe46e7c0457af0b93fd1d9
z57793cfe20753f49c3547940a259238a605d717412b27d1d1f3c8610c07e05ebb3acb0a0884df3
z2b5dd5e4980b376e0e59c4a21565ec97e1d9d2eacc03abb645b5cda10e831d652af3c02092ca07
z08ce06f8b929b936bf18515ee67488e38d5ef78bb6bde27d0d07f8f43ced6125478e05c6bc48bb
zfb4caef6613ca27b59430bb77bb765146c51c1bbfb3f3ca1c974ccebd9205d65582cb8fa2d26c2
z0c276e2ca4c1f8ca4da9b390501dff7a4516a597ec6a4ee43218c85e498934211cd89d4cf041d4
z3b88edf27253f836bc828872f3c294cdf8dcc4f7f8562bcea516cd2b0e147ebb3b433b49f1c909
z4fc5ad97a4ec6f5940e89e0815d03507a5243b13c7eefb3e2e657416d97db8e48b5255a44e1a33
zd10a870f289ab9aa551167cf8cfcac1ec801985201ae802ca3a2b41d9d5e630df565ffc585ce41
z46ed01bf14bdbde106ee99da953b5f2b4b634fa8168ad0dc2e862d3ac654f14b3bb93be4afd3fc
z71d624cb423d27eb24b55825420652534ac163678c8af1f28c1add78cf25189408fc1c02450361
z9991e6cef283224765645f143a5cc092d1adae76d6d61c3e32ddea33607f975c6b457dc828f098
z27791996f003d5e1c0b9b72af2a1de84bb633d309e287039a7ce2c5a755fb86fdcb013387e235b
z912a11b8f4107123d3179d77e112152c2484f4bf7041ab240e0f2ff488f8424b07efafe8864b30
zfed8ee5a8abb7b8c06967b8d103083f4450436b9906bf3e4add8e02255c595e766ae0b35b231a4
ze4e1ea7dd28b09cfbefd64633224bedd9c7bbfa95ea420e3e49a43294a621a6a55deac5fa54063
z648f92690ec1bde80dfec8658ab10d7f5e694872ead92e72faf968eae2d61594cb84e9c9d924e7
z6044cf0e4355ceb5a96b028070d84fb56d70ff6256409e2061938e7508f6e082100e1ede8047cf
z25e426f917367d79125609c0220caa6fe6bd19bdd6c94fff1a9904a13193c4c526f0973ff94278
z0b05e786d962635c98c57a9559b154a0f581287f419c7b4da9af72dcce77a58f5f0e72345774d0
zad4668109998b79212d368d546fcc30f87b21aa9d4236841b116c12cd0d9cfbb920a92e802b46f
zb11dd440f3f0187051f0c0bd910932f07cc84d23f7a5393b1d8882b744384dd7dd2bea35d89c29
z4dd26cbc1118753563b4ebe59ed7359d8674d0140390d15ed19c99d7629001a294f93a2a2697e6
zcc61e6f7a9f949acb762f051fd4ba86187e615aeda6737460525645324d3f9dfafbeb7fb8a79b3
zc0a84fdf3e2db64f4c1bfbaeec460b970466a1006782b204be5843195e0d14a47e0d3cc18122d0
z50fb48e3f533505daa918f4fc0c5da4d924e3740e1e2268fcdd1b1839749d7a67d2cbcd4625964
z662394c34d79c4d0c214f756404240996707cbcde5abc4ae578e48a8afcab7ed878d70140add51
zb93ca40b92f6f43ae47561461ccfdcc6634f9578d88a41b33defc3628985e283baf28655443d87
zc62396e1b470d79a1718bdb5a87000ce6bab72abb487fc498d3c44a4adc63fff727d44c52e04dd
z0d5be3451b45237f430b4b737740900eb0a0f3309c4017800a0011245bcd9bf597fec0dfcf3ca9
z16b415ac66cf50155ca6698e942faf34c847514f138b703f18cbb80374aba646b2ecb262107130
z5b2276c36ff345e24f4a6033de89feedbbbcf8ebcc8470b08eae960866b01f566a1aea22099fa7
z292b605ae2982bb67686ff0159938781d8dee0cdeb700190590734e4d489ffc4a37829565b4bf7
z12f92124f388b85f9bd67a64378d61f3df3da797501f68d294631fda54af39d41c422b81809c0e
z1b98b0d968b793844a8732d0a1f3dec7898a444ee99d827bae429bb7432f35a54c6c229e319cd7
z033f5ce028e16a68a67e4721029116d8e2ebdc22914df15d86d79636cbde5ebf0ace26b7f61202
z4bbf7496a642cca6193b0c461ffeb99ebe0c8215ba22e0527edec44989e4c392867d15ffc54529
z4abb5b33f06797dd20dba0047c44a2d5b0221eeef8dffa66fd6efe7d5122ec573e844e18190cc9
z28e500bed65ba65aacb606d9a41961f08dd8dcafbe1f5000baebb07d6caf9a86023444942fe71f
ze96a9bb3a3e3c3aec3759636eed41e749e35234901074a981ee9aba1e2aa08004469ef0584070e
z19ee8c080acef933519d43c66e0ed44f307a5bdc3b88747db9d4f3e9229e8b3a90f6fff5925901
ze984ec76e6a92e8789b71dffab3c7eea6fcfa44285c92d013d3ad75285bb12fb81617c088b20f0
z6f2acdd40b875e607703dc615ad1b0a7cfc3ddfc7bdc1efd46b9ddeca03fc95c8c1b7baf751639
z6744d1d25c5b2e44df85fded0b64874f9de0ccfd712fb9088199f360c02818e45d194644ea6259
z324257f9a7293ee1142a8ef119c5d56f07293540a81dca5b94a281a9e447c9392068ca2aad9021
zb30a4943d35c4ed0faff66e5a0bc49b38585c71d8e44ec103a47b314b0cd8e69deb9c1097ffbe8
z3c83ae49b60b719682605baff0f82317b97a13b379d7334137c213b75fad944dad74eec2706808
z9f695ea9a3241fb7b1b9e8feb4fdef590550c629a1ccead83d1be949783c88a9d3dc6fff93afe4
zc98214c0b30301774cbd411298d52b004bd5066572d478bab4f63594fd21b82abfbb2f07df2cc2
z186f2bba4e23109d878260c257dc2d47d652bf89a80678f22073ebc56b296faaf1768abaad3f8d
z07d08960d13cc3a6883f2f916a594155ebf4c4fd1812f92ccec18ae0c9f5be014b266ef065de48
ze02b5e6cd50a1c0dabf6b7866db2a6cfe2e5cc430610555c681216f7a772d711142dcdeae2b09c
za8066502771b191a8f2378c130f4194af256e89f2103acb4bf4bf551b0c92c6521040dfb82920a
z6d82a3cf009a190ec141f2bcbc6090decde908e4930a3cd28a22dc555469ea9d159c0e741429a9
z4e5fa7b20413ac6e7cb45866b02100f1e8876195f19c54fcf8cd0aa6f77b844f1ef890415b4b46
z67483f8335a07176a8b131db659dbbf7cdcddef7d60f6bab776d4281386d5fdf545853e4c9d74c
zd6ef21d3cf85a1768f829e53b910342cde0b80e9a53601b48c22cde54caa8a80358099d3f1d340
z0e892036e2a649401ff963cca21b37c956df92e5154629fa1fc7cbb722ed553e3a36053f0b28c0
z8e10ae7fa39f920126da29ad8d3f5a33ef85f33215fb4fd56452a11ac245dbd2ad850db281bc39
z1a7e606865a89704f47d965f3a5243fb904ed69d3feaa9e59aa15c4e8982a1b13047591b4b3e9a
z2dae70883f6b467b23848e60e067c4429742bf9544804300b7e3159767e8ea26c69e0fe079a194
z216f30d38d4d078b9e3c3dbff258ecd05f0478b3653d60d2efcd6deb26f91f3aa3ff00003ecc71
zb659efa8172e7f3fef1ff9e62dc4812314b22b1d5c4090d51bdb0558778cbc22d23e792b019221
za0cd2e8efa8beebcb94630d05cb7d4bccff0b39dbcfd226f9cd978fc2d63fd79ee229d5722dd81
z3d7db265d128ac1a4cb9033c1965cdfae8102f20c955737df3b68789df545a50206db8a39aa28f
z5c12e8214569ef4d0122235a16ec56e77047b25133e836ef71a7fb9a2eac04594feb89e2e45dd9
z53e9125acd7b2ad4486c4022ba4e5b68f5f9e64acd117e49ba321d179bbdda5d0664b6c6091b19
z5c0b218cecfaffe4a2c3a451a37c769cbafe2f887ae898096964dbc3d5c68985ebfa69c8d098df
z4f2c0dfa75ad328bfdb821ba9acd6459d358cab4cfb93e1798f0403d4c78905f4b3ac4b3aa8140
z3d00a71f992b23d59fe9d78f4b1420ec80295ac57610982b5a4825b8bd1c95ee62c47c23fb2bba
z55f7736b8499afecdec922be4423ab63fb81ef1032caea812a0fe5e73e22d966f1ebfa629906c7
z8ac0b8a1654f0488830cb63044165b64a1f4441489ca3ad6cee3bc7a57a9216098acd23092749a
z438b885d0db25281d79676d583a7d1c3a0e848cdf2e767b30748557c3e8d9057f9be866fcf1214
z75deeea29e41770344931b758c0c36a599e4c1834034a051417b691f12711e9519ebe945cbe2bc
z87d146fe4e898188f6352889db21b0edc73dbbe9ef0c5aec5f9f6ad4b250bb094e4ba21a2555f0
z419ffd7b94fc9992ec4a90be1909189fcc6789321dcdda4d75750ae420cb29b5aeea4a1b2863cc
zc3dc0ed821150d7351005f21ad7c568689236fc52cf0ed237ceeabac0da61a4941c6476de99820
zde226c3a0d590600ea91f9118a9e06f294e6222d4b725c48ac1e60a93ef4209f6ce3396ee168f3
za1efe2601be80b7e164574e65962926d15ab12e4929eb2328bd56f6f69b94d9de5a62429433cc2
zd05bf29f6d08c4bd2e2d506750701d65bc67324609b8edb783f29a5c184320dd7a533232d87066
za9f2571da2fa772e924bda9064d7e647aa9ef7134ec0f2e66ebf2b4f3229c8349bb6679893dc58
z2bd40bb5601885e9f7dd8d248f118a6119e834d9ce6956061d6917a186de9de1e5ba37dc409fb5
z0a14af2b8718476d9ed72898df53f03d4a06b0fb5fadc7b1ef6255514ba19d48a2378844f1e3b5
zac0341313cee0060ed7b8315d309420d0872042e861d8b478d2cf0812bfa8750867c1a40d4f01e
zc9b41de690751164369eabca5a1918db2e73ba71ab204ebb97dd99d57fe9cee51131941eaef3c9
ze68686cabb16991bce69a9296f453ba87bb87741030baac132780577f42a7f9aab1eade0fb4df6
z7ee7d514af6efdfad9f652a9113ca47044aa4fec6cfe492d2c07c99fe5d7175642d637cca51279
z72d1a515827549aaa1b109eb5db39f2d9a13b747e9d163381c56c8a9396873f4513bd3ff11851a
z15b5a05e53d1c99f170c32f429b857d24d5aba41c04061c9cf3bfee33190f6f72d4a413879bfce
za46bf732f0d2bf1cfb3b48a4f4dc52b7461d13b405f9a6a2019b2e13167e13e726af258b4ac60a
z573c25ec7972fc4943ce1b1f99ade08cbd8a54573b1ac8f4b1672ac304d9e0151b241cc7294880
zcaf51eb48a68f271cc2cb39e5c43e1839ce874b148803284f074e70814657aed7311ddf7d76329
zbb41e6d61f2565bebe5c43fda694683a150f4c7bfa744b47a2a5177cc72cf7930b95a2a736ae86
zec9a3f095906f969c97174707d92c84c9de489a0178dd86cbf6b6b49569324c4a7febdded1baf5
z070a7139111f7a694f04705094a60ca28770cf121a4a60caca3784bdca3237fc35cf92a07e5d4e
zad090a7790e04f1b393caccca9e0e773671e6ce3e85b223e5bedd253f6fb3df9ed618d46633a82
z4a8c3832899c3dcfc72c88c786b252d31c7d5e156c64e0fcd684c7f0663371250d59809b423c46
z52fde906a61d0d5adcd5318aa9865c5c33259f265a1a4403f2267712e1411472eeee3ffc1cb850
z0c114ebd91b1fdeba85accbcf3a4da6d8e4cdbed9d80051fe48f5294465e1fac757bb2d265dfb6
z972f7d318766de4d3ce83c150efd2bd53138b0a4280b7f3be9a6cadb1b639a40bd4838b2de3f6c
zcb7e1f3435b88fe0f704b7481816b45043798a9440f0568729545e628119d903b2715e3c088e44
z93c04ef05f9e15d3d70734c8521ce9314734e0bdad590a7c36121abee7a68d9b14fdd1fc82e141
zee559884298dcec0f103a9533c66e64c68334a664366c281a1c14a20162c791d6f60fe37fc19ba
z5d3009d0d855866cd27ffc28b23be51f37819d5416074ff203a411f39d5f95901082c7c64fcaa3
z80a55a33b214f8e4e1380a341b17dd4380b5c13a85ff387a3ca1e2c896bcac423f52e04ca2dcef
z4f225a56a8f59680d1f7fb785878f061fcee49e3b2719f77578cb1a44646b303fdbebfbf94434c
z7692aaa18e25545b01b62760b819669d26ac8786fa8e4677530a218e4aa63df3366df098600bcb
z877648a6d3dc843c8c41883e3dbfd0d9bbf859df73015b2e5cc41e9afbf50d84e41c2b13d6bc59
zfcb041b9e6b3771847ac490f2df7af50dd98f23e9906e246618e8791d1fcfa795584bf727caa33
z24135cf5875d28d689cd6a874bf5826d3b494a2e8a829e3a6cba4ff64b5cd1f11774e5f080b86d
z3b90e85e809782bc085113c5428d0173282a82bc59dc73cdcd793f458961c88ebcfd6e0293e2bd
zd2bc36e430fabb31388b3f4b89513b2c108266a0a3fd876b3c5b6356f6fb440647a163969bae0f
zc143190f34c9eddf429a6e2d5920c922d5aef91af49fb3ccf758ace74c04c5a758b160ed97f451
z101d0ff68dbded379e569e6a6a6a5c174cf611e364cfe0b25313f40e52be7170c147347406adbd
z87245e967246189fa727b8b0d73317b2d446900070ed348b6682b30ca33b2d72b89634930fe35a
za229850f07029177a6446122c8ff77ac734bf35f6db3de89a3700d5bf45a7e21f3771d2102fd32
z63bf90c20642b5cabcecfe7f5326843438f74aba49b7d8abae80c1c4d8979ee429937f8dbab5b8
z0dc0fd98d703a98b5265b88f4fcea6e323e42de58fa1a2f9fd809d4ba522722dc5b103ea6cecac
z705e7be4028896ec8c8c95c21b0f4658f9632c42550bd119a8503c68b3b3068e5a39af3f1a1221
z62a4593c886c210ca63f6d3f1299ad51b4ccf1c544dd2db7d6df33d6f3bf9f1c4c05c7286abd1d
zff76d11418b327da6931b5e7d54de6f761b447580a6e957570106b7f6bf4e8e47b92dd8418eb2b
zf9505d6fc7583eadd4bcd6a523d6fcd7d615a8812746ab206a05a96185412f80ec8c77e49978db
z843128c6b2694319352b507e093569eff883eb72cbf58ceead99456a7f8412c5ff43c76da50fe0
z2a00f0949885d5d0e5b6ec9f8acb7aeeb94ea780dba9df2b46ea4fa0f421c7622b713c96dcc845
zaca99f01bb9498f531919017d361a73b394c6b7f4ec0bb521b0015624771e16d627dce0fe4c723
z412db59ab0b8de8f50ac20bfc29b580319d0ba70910bebaa88040a129bfbdd7e38832f3021087a
zfd40091d5c282ee747b65368d3efca147d81a697dc2c54299da0b207cc3ecdc11741a714abdc44
zab905655773ddd0b60694febd893b085e761593835ca0945ba2f23d24bdc4e95d55c42ccb1bf4c
z5c1f40a984493be6ef4e547fd934c9ae0f6e753ec21cb312143bca2ad9e4f3622ff54baf36488d
zc2a443105113642b96e6eb8cba29051239959bbb28e5e4004c8ff578e6ca93765382ffe2b6afcc
z4c5e132ef905ef3bef85e50fb3532040045790a9408c7db243129d43ed54eaf0513c829a7eefd6
z836330669e92e769cbe6e9083008cc663e158c2a1294f6b9f97fc4e0cdb9d745d233072ca6967d
z6a07971ce40021d879565a0ce67b55fa321e166c798b25a792cdad18b8c3e514f68579cc1994f8
za3bf14c04dbe3bc5c76bde51b162390009c58c42cfe1eebfb14dd78a45f93b4ab66ad2ad50ac19
zc33288dbdc609f5e35572f44466312c9fb1505ee7a0293f2ce56b59ffdb1a2d1812b19e3ac7ebe
z82f39df64eecebc7b1024bbecf8e2b041f236ec24b28af61285a7ba8b69956caed5c4181bdc471
z0a8f2ac2d66d2a728074b3562f4c50f349ba00f4f9a511c0b255e6e6460db8a6f32f6d89b3e798
zd57ab085d981a09eec95643481a9c2da104bd8f1e41fd0a636218da6489bc12121f53227a71b04
z98adae5b4d0047f5d023e75ca88a4ca8d9e277d79ca9f242e4366f531ce00a37fb7857df325230
zfba17b7a5f228ea282654a500530cbbdb2ce4eb18b2c1f4f0cde4d74022a2261218f6849955e53
z42c209c341639258e0ce9aa6ad34aec2a0d13678148f9ea0ff60ee0fbaaaf15cb9f7ee14b2687a
z390e366f508ce15c2960dfe63d449c45fe3a7e464b012b145f708c15b6521f8e5be265a47d2b54
zda66dcbd3b128a814e00dff2824f1323e306e7b04b34658f759d8a605a2d399db7c81c0160e4fa
z744c08d680d5343ac46a43dbe3f29a5bbf1f7ebd18eeaf7be4326781fe04d737c8d29e10d8b60a
zb96dca91c11882aec10a77e03d115ffc38bd11bdb23fa115ba587df5e57b7fd05646183d1d30db
z78f399fc28e954974a7ad85a16fc7f36f6849dff826bddb013cbdaf71d0a952cd58c42cf02e09c
z65639d019f0962276873b779d3ac043a596715d7b2098f44a5ba0bea68585054d2927d22c24738
z2ae78cc084788b83fb9667f1668a0531c0cdc6c131f69f026e0fdf019a1b9a83a805f85e22eb22
za6f5a40a662176b484b7a44a3f0314fc715ee3f3b6f290f92318d1a6e2633d75a3ce3c94a3f193
z3312e2acf7074500019c7ee28c40015ba3b0884cc75c492330a9c2b90b1fa9fefd04bac21548c1
z13c3b6c0d849838c2efc8048d451f87ad1c1a328ec5e5eba83ef978cd87665e0ff27c5a2661bd1
zf1c3dd3d6a9e64d51238668d67577fc2620cfbc2b9c1f4fc9eadf7299be94265c11e2a7b6541a8
z159810284b89e9367e6ceb1898a76fdc9e36b6518afef582d44d1233b93719339953e4372780c4
z4b647463d22ad174e9916952e68a91120ae75a32c2cd4744f5a5648bcafeb1d515cb07a35e3051
z1faa508e56b0feafb1ab299d379b3c42a2be547f1f87528f471de2f49bc4cf40f9da57f0c01d06
zb2aeb0fb5f2c5fbc90be777786f25b9847f4d322757c2570b21e46071d88fb87b07f0f4264f93b
zadb218d4b5e010ff064869ac4d928f1a31d7aa6942715ae9a239c9c0ec2b2bbe0989699a877fbe
z7be008ae8bdf66356f6227e17a48b9c58ef205c85709ae8bcfe8f3a9c6c99491de3800e7a7e486
z41da956bab6a9b0005955d0dd62c6684fceaff3202893dc322a906bf9afec7eb02bc59e98d131c
z1e1be027bc5b165e4ed7d797d8ef85fe28327cffff2c56779e356bec6953d44ec1d245a5e4a471
zbc00983e1ce439c14fa8ad8dc6f3f795a6cec298d612a0f1434cb3d566571e1e58973c5680e02e
z8ea6000fb2ffc901002fd1140f43b22a13e011f8305f285d75b163c54977dfbe4ac9a5ea6eb3e1
z2967026b05a52bf006aeed0730590fd17508be836a847e079564f755d1a09ff67869e5592f5170
z464e7247885bf2e6a9d7c68bc103f59061cc9d7f1d0ea63c542bd530a5fc404daa63805cfd969b
z9582255c55445e83f637a3fd45f7ceb683661014fcaad50a6171e33e948f62876b903422baf04f
z37760bc0db05bb30da8b8b6c2f16aed61fca6f368a94eb195cc78e463297de97c37d2a6ea0326f
zfe63367c182007a4c8afcb21f79f1b45c9880a356157eee7ce4f2ac9ae58c14c60370bc28ef165
zc1cf6ab4080bc0307c10ae7ed621f20c42e8428655fa84f5ed9fb52f7aa51f1429006f746c698d
zb1f9d7681bd2f19db7a851058e24f592d2b5b183305c94e925c2515d86a3cb66941213e0607839
z838a5dad1c5295d739222defe091b9df74c196a59d0524b8cb4cf3a5d389d8450f14d0a6e51250
ze62534761da79cf5e37334a187e9771f74a90c4086609a0bc20bfba5c230127a1a71ca5dd55e8d
zd87807b64f506bd473a546bd6729f27285d4a107daa54999269c57dcd97bf1d5f5bb7ced982d68
z8800b61bf40d3cadf7c1d7f19fcc6cb487c76ca978848e3ab31fcca02bb36df1fdafb5f88ab9e1
zea1ac433b6635f78a766189c181e708216f488e4f297e249e98624c0f128017057c619073e8d44
z3b452e9c511db019fffc9c78c4eb92e1bb399e0d520f4acf0ee810bb775047d358df7ce0d82e86
zd1c7321a11e65bf3062f484be6902ec25a1fee270af7261f7008e430841d01344a2cfa0c652663
z38d3d31254ed4483c6282e2728c50036bf711f116ff0cec1ef7e1f95b4d8dfb7a5d072cfb5c783
za68d9e263798902c78cd12b6d5237ca95bb0ef046e4953423e3560e7042822672d49954f4ac934
z846176ca6436615d9d79d9c338d8b54d3844773e1db2e7b33274a5249bd4e20299773e0fb5d283
zae65e6a720b574f8b2e19be88b2dd5fede0f6076dde6485a07f4f8d2c25446575a380a80c2447d
zee2f09ae829afa5a1e143c6637709e1375c98ca3b479cb69e395388cb479d509e30430897b98af
z33b9bbedcc37f2c5ca24db4fe1f687f26f9ceb3ae79c0a7f751ec1be6150ed0dc4d1d855640454
z244b1950277646f4060de542541dcf613119a5df3764461ef1b302f580e31b8657b88b778546be
z5f6d163ecc1c3563544ef601a1dd0dc18a06de1738fc0db428b9cd358dadea8edc07a2d9dd139f
zb9c9037c65aca8832a4c428640bfd2ef1863c9c0a9327c40a302ff4b48a8cd308709f9f533ca30
ze9f925295993c387fedca14f2565cce1689ae7c9604363a33be2705300f0ed353c7debb6690c82
zb2ffdfdc23df4534f5d1e7ade9ef1aaaf0a2187c74d5836a81292493deb01c0745626ac789e7c8
zbc73eef8c0b8f1077c3251e718e899b4b02e99743ab922d4f65827bc5cc7de4bc0972fa4de8b13
zc1f80c35f21f17fb927b8e65d2dd45ee8d3c4070de42e122e310b2a158f0b09884c6273dcc36fc
zd11820dd77626fce8a2f6d3cec848825def2fe8dc2c37de53046b721690c0c39a935d0b275b768
zfc4bcb4742e913f7fa6e2ab37bcd0521b31e0512ecba94ee95eee2c1ecfa955408fcfb95182834
zeaa9f6a40c8ca5eccf0170450395f107946a8bdd5e69cb1173862834fde8bdea13ebfe6433e358
z29bfc7e5fae5dd48c8c2d2b0e14039fc6bc68a56a88039d32aa7a8f2c67131e942df2a50536d22
z591ab4ef6f429c97ff931d1c7a4f92d23ebb9f82f385662d7d2e033cc745cd74f6b24ad7367133
zde67b321107e77760f410a9b9a96d361348208646995e962400a25f75286f977b0d51058f9ff87
za49fde8781b22c83e70c60a6c775b4fee043cf3d55cdda9a2f0d4b3b79a0bc8f3de3cf01e9f0e4
zee8415871448ccee6546001b0c9e5f30097bd985359807bf22e424708b0c638afc53967d3461e3
z287fd313995aa31745edd857c9efbcd8f244a6ced883dc2e11f5d79fa73b261352f0c694ef133b
z79826f68f167b1d5205b9a1e96003ccd40df68ba92f4b0234541f56cd6deede77b04b56fe47aef
zd5d5f1b95cd6b490e82c5ab1d5ff4350d2e3241e3bd12d45a2a42487442265d440e07e9e69b9f7
z0ab7d351e7560f1f6e59e6c4cba61506b5f2f20238e877d0153afa4fd936fef5babc95b509aba3
z7a3983df969f8393777e5534b0129158bd9a1b78aa3efd7df5659717d47de2848429bd4b0e7c1d
z87e6061d014bf25e3e0e163314339f14eb46ef2134585f391cd58938c2d1c10ee0fc8a5d265233
zb979c08d9410beef9c6d07e0b430a7638f7c6a48b9249736db95003d9e4b91ee284d1129a11307
z43758c957f8bcb0e4668be8d134363fd3b90fdf05690b98a6c530fe736c7ddce90c026f0184426
zda1b1f761e653f152879466c4378fd42c300c2fd9bc543a0c9c3dee2fb66cafcd71b89b72d58e3
zd8a33584090213b49fe4766e6b40ea86217c506ae88ef80862fa7774e73458c1b8b5fc013d7c2f
zf430c66665d66cb5a668436435f193d8b0b40c2d1f25a616409c713720ab5b0d444b909e65023c
z9746f93cde30d471b045c9bfedde75fd3f4223cf4990eed0eb79ea6b40532efbbe0a456e1b24a8
z6a1eecb148f91227519480aefa7efc97a091d7eb3016713bcff2b2352a99953c2a6f258a492160
zb7798122bbaf483071778989492049131fd25382da8f1e002c7586aa79b11fa2eb52d401f8cd8e
z387fe2e5b0f3cafedbb5ef3f73f7dd57a8480a0166e62719a58611264c4d9e0fdfddef1a11eaaa
z4e02d77a8ad88bb1da7b553be920ec934f51ee3c3670f2aaefb8f0aa58d8e643cec6a75a665254
z6f89706b5de0cd3bf963658f47c3c03727b1639ffb28315e946f5dcb1e9afa7b524ad09e8423e4
z3629c1c631629700831085eaa87ca0c756b23e07c0c7aae4b7af8711fc5295c128523f7d962c76
zed5d6047641a12adfd3ca6a78f221fa547956bf70724da3932d058ec416ba5e5647ed51957de03
z48dfab395dde068dffea1ab627ab0bf02119e1dff9661c6c2df6c3e0ba30a6171cf43c53b4d1ea
z59c1369379a5ecfaa57b416cf4f5d63213e635cc5aabdcb2f6e6d2a3447465d4a44dda4bba8c9e
z8e7a2dc01a1f1cf026c878cc6959df85d9ee1e49622dc4ada2a904282c45ba454450f8e988ba9c
za8e4e9b088f5f0039a4dda9536d3bf32020c2c3d006ccd0e01945a557833053f7e6a2b87084b23
z707896ae38f2e0e88a7552ea710f0f9fcb5d57746131d3ef68b4738d71d2e301511003fa99d606
zed19dda1cd5640418049b50a91237ceddc65ce108800cbea064290e88e74b1951a3513bde2cc7d
zd30536c5295dc3e2b62f4888a0186cd6cefa2f63f408267b7ab568a70d6e19c15e103dda5af5c7
z4a91f29e6a5f7a7577f222e8d72b3780083dd725a98513b0d49bbc0fec798ae566f4e4e936859e
z7ce55bb57c03e0e42cd68a457fef9b4369a8f8e8e55e7f2b6c0b76b1e2910b7e440febc33edf3d
z210ac139f623fb5341b7a15f103bd25433615b2b3baafae80149b08c60881ed1cfe3e40f9253ef
z6dab74ac2b261969278d6e5519192f9b8f26d458aa73dc096861e5eaa1ffa68d0cb48f6ceccc50
za0bc7d12c95c36935854a900661501a5fefa4cd9e1c8a9d2904783dfdb78e963fd685b28832acf
z0366850b0c5cfa49300653c64a7f68bf7601b9865d28417ef5a24ec600d473ea3039d7a48ea2a3
z150c6704fc4934e4f946b60bebcc72a2fa274c2ae7319fe3c387136de6297e3647ae730bc23610
zf168b4e1766da2c776efa3ad3bcedd7b35df541ff099397672d597b9376376ca01fda7601b1e7a
zbb026f01e8932480d64e82e894016e58027dbd41d663de694dc200cd2f192781c4585c7fbd183c
za6e0c7f5588ec95a30f0a5b3ed246ee993c412660384ffd3c03022a262ee45494045a9716f218e
z44ad8ea6d65d5e3d4a313ad6fd21a77188a63c528f5721e38d5829e3cb17e7801b4394b01c48dc
zd963c9ddb51c3296ea0bec5ed830471a3997df5c90731cff315c8aca4f80be9452a88e06ff4cb2
z69efc110f27465c599a1f092c6a33ebac2dc4890eba43b5cf812f1c8626e6d96bc46daaa1260bb
zd493893fbe6f3a0e98abc124165b375b2a60e3f1a1c8ab1765b2882ffe7a069b4caeda5d5c5bbf
zcab6709fdfb2d12277cc2e69f5cbab65cd97981504457c8f9ed61010d62cfe608d593a7c157ea6
zac15934887e9aa521a7a39a6a7066c4c9088e243c82e7a7dfb27e54a9af68145962d25bb09213a
z89a7a4fab985cfea52f3a0d9a99f3c9a7c0d224909003132b21c83885e9e4816200628b0dc7134
z8f38d1697d65d9fce8fc5aead36e8571cebe278d6cfdb3d40bafa772da50320ed3670c32b2ccf3
z12dc2a7886894c51f929b97c4f200ae7ae08afb0f674ce906704598bae020dac98d3d1c2afa025
z04c977fbc1a6f8abd5f2c2fb693512752839f02f73dfcbd8572ce706d7ed8f93761d5748fd72c7
zd05023b83688c2dccf7efda2d1ca93f47e028a078f7d42f7cccdc7b9c7a805553090f1cdb5589e
ze5d262359f6875b6e7980dbbe232c37a6025a4ea5bb0406b044ad7222d29c8ed666f7794b3179e
zf154d1a610c707eacdc32f71a23fd5a77eeedb97e87a7625bf8c83f38d1af14a9910992d4d2ee6
zc95060973dadd9b3881dd5e0f2ff608c0930fc7b53cf1e4c51fb3e8e509ba0c3bba2c3c931582f
zdef67e7b3ad97cabac94b8fdae91f8a59bd848b4f5235e650cac2f463e7a837edc89d53e3a1cc7
z9185ab68d1075a330fbd2a424636e0b7f1215c521e06d8486ef3bf23e496ae35579c4ed4376dae
zda6f830c3571060a615fa00dc68ef3fc4270cb5ff3445b0a4f20b971c1e856ddc41f8af832ec82
z84d65cbaf317cf23dbb4d651b451cb200c8d8de092a7e8fecac096e42d65b10866f67e155a5d42
zb774d2a752f2821a33a1f2a3fe1abbf0737f46a449e42900822c3e6fca44662bce8c09d4eb18a1
z19666d194065d424547817758f567f7a53f1d189de6725a82efec384012641cb60c9c5970168ee
z31efd57e93522648fc3315af21e90b89d36048607fc3dc4e9c0ec0bf00a5ed1827d149893b8d14
z7cfc748316b0e603e35f2df8cd1606d26e8262c001d9934ca9a2dae1b18b88bf913959769785e8
z4e1de449b7d80002e3a32ebc8f5bf402f26b5f0848c5c761b8cced9e424ae2fbbb9fa10b69a4f0
z994030e45ad4f42a091ee1b51d61921d0441e32fb9776061d52c39503d9df2cd78421852a1afdd
z5b9f3b001b295d88a503fef9f415166d73fd099faad7206de88dc32e95c13a05b96831f74de5fa
zc396868831de56bb0b3f90491edb64fe65373e53714dcf1690ea26cc533534abb9eb8ca190f7dc
z77c9a0dd0f198c56a3c7ba070dde18a2f6a38b5575563dd2025c37fb15ca08a1d8a9c04f7c79d1
z4f17cf1babb8e862459067189320b2fdc65b91ddd62c2e6f727f85b3e4953a86d3b9df40133014
zf0aaaea90e79d14920d9d566429e7550d80fcc33c13eac67b5ee943a16b716c9f5fb2f9d9a3d78
zb1f7fe4ed0d809403ec805c8b0cd8f2f85d920c892e2c40ea3c58372013743991104f5f8c80c01
z8b8c358ce21817e79a11f456c6b9b65d189bc657b43cfb0d852e4dcb1aa9151497fc7b5e015d8b
z8ae0c8d1de02a8a8d0dd82371c995e1735c2529395ea884e37ac518cf767b571898f15e1ce8c57
zab8cbc8383ac76265ad37711ab7de10d011766e352c1897734f1abb9a8b3a551868a451ff3ce8f
z8e58f1f0bd482a552c306bb20e46756b4fc9a656d233bcd8f60c2bb1dd38e30dc867291f9c56e0
z0dc721eb753fece1f4d64925999810cf04f26c3fa0172a78d02edaf7799b7f3d517189876f38c5
z3854c44a1d6a9544a2cf4656c39cfc45cc50eefae2affb839fa5593daf28b0e972843a98b60d50
z9642b6bfa238a176be4f44063d5bf0d61a4e6f376b24ab14dd3e325307980f8dd789b297c77688
zfc13d429b3d7033da455f7b5016dbab835d316cc95dfefaab369189666b5d845ea47a11bdd4436
z162d93f6b7031a89778e3bd5297ead6960660c502f695531311964097ddc0fa58c00a21ec86165
z46188c47844036d96a891fb4545b6adaa8e893fff147d531eb000ea037ab7dcfd239ef5743d112
z89e8d6a6fae2afdff3fae0f4a2d04a0949ef37fc684517fb49dca28a87d9a8d1b8630484021575
z8cf00d91e95e041c4a558af85e6483b73e0cbebb0bee49cffc653ccdd1583b1255420fd4e1c394
z67744a78bd77070ec0aa49a9600aa056b54da4bd0caa006b9fde59b9a16066b05a9a9a3224a002
za139fd7d52c365a3ea461764858773d5ae72b3495fe77475077594e5ce7f644eb784af04f7e01e
zab8762a75099eb555a3fad81dd66d1d91f233a9ada8ef865313b06a7a94789ea121e2ed14cc872
zd630482d0c9d3a445eda25b3d38fbccb2da553fbcf68222efcdc4938539097a88e2af4ae3101fb
z459cd4ec1adf83584706409e1031403fa978b8b1ea77839b290830072911cc6a7cd2e14a625a8d
z44a6f7c3f8d851e2026fcf79d2e95aadecf6cb9a5a62fb2584cb3a9af4283dd6ff32d883dc46db
z20fd564a8327c4a862faeba90f9010936a30e05308de0e3401bd2a3f75bbcd0fe7a8a1b95dadf8
z9943f3f350f10e818b050640233b4802416c2ff06477a76995e67950a9f62e4a95607497a6a730
zb0bd4102f2b4f90974af24dbb5eaa2875a4e65eac72a41945521dca448889f346afd599bd25cbf
z4f58a72fa2ea6e91f195a32ce3fcdff42baa82041b2bde71d7b0079f8b6830ca59626ec2ed01e2
za07c887dcab03de3df14fbb24289195e033a0c939db89e318794242cdb205759f6f6e6a499b1b6
z5d2f998d8d3291023675be0aeb8379911ae48cd63698f533f3b14dc3e544202bd35638fb352263
zddce86d93248d19fd8cd93c08f2b80f94eee19f03710b1c8ddf790acc85e0b68536b659131c281
z7531fb69609a167c7141f6d9c8a0902019617ef487daa5f52a420683262945189c2bc04ba5b049
z074ec4db89115dd77b1f6731de2426a9deffe5d5d665a6e6a01408b30350cfdaba993120586eb3
zd0842cd2beee6d4c2f756e73fda55daf2f11ebf700b89419778679d2b442e992af2b919ec47aa3
za337d366bf39b982b01030dadeae4ed4d71a05fa41610edc7dc3a6dbb0daa5b56a5ea90d52f449
z7f930d947e2b6f1f7a53c5f6c5258dc063d3bfcad6cb7387c8da823c1f220e56ddb88195ace606
z1e12fbeb4c99a3304a24e733e76022bffb353001381ea53902e241c12807f9c769d3a65361e503
z10aa65c4fd61c46c5f3d67b13e424cd0476b5bfd59216a4599bf3782ddd89732f15ce49fa17731
z0f431a808b7d29fda6bf1d106c5adc505397da1bd0b1e1e68ef0f766ced2664ac333794b183795
z68012ff3937ae6dd28a7fce9af0f08c32b7221a8c1247bf7f8be5a51887ed29b4e46062bc5bb25
ze4dcf28d01ad7151945d305ed3e0ba1618ea5d6b38019c78ab2b647ff911c1164a92f9d365df82
zd88f43929c7424fde6ed55ed89ab682f2a8b61c85b4a2e9b6669af198e938eded09613caa9e17d
z4bc21a89356ae2e1f44ffe64b0c02ca017c48a28adc81a784eba72871eb28767e4bca99b669c58
zec7b68d464a49cee26a2a525e939f1ed2aafd05f40a76845e187ccf8f4531f4930eca6288c0a5a
zfe98ec61fce37d8e472da010be3c8fefb7d518d1c31738df031a4915b05fda4c06a8336b93491a
z6a0c85ac63a79701b0e2d7c302c80aac1680af771d5021a69d4684c9fb173ff35ca5325e71dd49
zd71c84b2bf8957f64cc3a23302cb6049be8fecbe107343da677ab4c1d20bbdc9d52cc9c29f5d85
z139a44ac16b18c3f3d98fd8b4bc6ef5cfd2d9b75ea9d38d9598eacd972e7e52605f3f073e500c2
z1614c086b0dc4e6d3917fd8afb40cb924d1b8dbb5f12416b59d8616bd68dc386d20ce6d1d29200
zc7756e7df4b836dd12644cdc74e3482260ad4f4d334ff8ee8c3efd728cbad25329bf76b275af92
zcadee0ca45bdaa9a26956d06316985549c04896c8e05b274b276fa0884a6e21a0ed83bd460e183
z74eaa3344df2324eb443cd643ed73a87cb98c4585faa6b387771436b2c3f1796106c9711ad4602
z7e10ef5ffc4d6c4d5dd6bbec7936ebc0098fbf690d53ae60cf5419cbef9136d03d99bf63bd67d5
z7b4c785e70f8c8033df7cb4d65697cc7fe893ba4f4d2a0af5c4e43447b1bc099019037a808041f
z2ce473992f354d715fc9d68c44e676e4138dcb42a81e60c978a976adc96f552929de9692f3358a
z7724e6ec3e96e25a17ed2529eac5551a5593c4bac37c3dd1bbf291fd413cd7afcaabbd16424d3b
z484578b5f501976b3e72bfd767427818291007eb231a10d525870954f212347ed009b4bac48b3e
z64130b9ae7307af672b1261111be3b67adf22465675b38469fbd01799eac5290ce2efbe1f939c3
zddf6ad005dac01efd5a435ee6fae3f82f3cdb189ff11b7a2f9dfa7bec4800d545f1f48e2f4b534
zb3f355d660cbf94a8d4211ce06d033fe827d66299569cf768158d199e1820e98d34f21c7fbd030
z4fbe9fcd5ac06391182bbbfd60f457a50c756a858e2a2dc45ff1fbaa7da849721b94a074cc6481
z734770d701016579ead19f6a851b15f114dcd29525813d314049a144045906d964eaca1dcb3cb1
z770e193717009b32cd15d7183923ae3002a47c5dbcd70d737e9d3f2112954fe49307b105ab6a28
za41ea66d6cf2b074544922f46b687b490e7fa4b4a2213eb9066c97c98b3c7c62f031f54eb1e244
z23d65725aca7335f1039d59172544ddb22eb4dc3a336b89d13c8b9931cc02332940c02ebe38234
z07678abc5f9fd782130be2ec82388eff07b6526082d73e13ab38d91c7bbb4f7f550bafa7f088cc
z62872ea2a93aba0b85af28ca8119867e0cb30fa62fc3b6fbaa54174addb1235e0ca77b04212e02
z2c301c86e4cee1005be1271797053025a8e8cfab486a550c03d5e574a232780fdd8f0a96558744
z279a6a9be4bddb64249b9839f2644352daffe857bc2b77580cfe9f7f945d04d8699391950dcb82
ze51c3caf12d72f2f5ebb28b9fced6720354823ae98c3b0ce513622c63a711e11ca8914dfa15a57
z07d6d71a2fd80c9701b268a5993efe24dd5fd096d3a8235ea7b4cedc986de5eb899f72613dc862
zb260018da0eca1a25ae02bd1da89b638fc01594922881fffcddaca807e976b1aecb9d86d7a17e3
zd5b05a68104b1702cd260f5cddd439851bf0a41cc97b99a2112e55773da7cae2bf4d6399de7139
z1213cbf6e7ba36fb0a79e9fbdd3ad0d9895a418c4d4e96e17cfe31733ebde946b225f682e4d953
z3a385ffb21341af8556ec95552dda4b5ab4998a87679b93df66f8db2b4d2eb5c081aaade427f57
z02c1e8e2e86b2487455fd2e13bd34fee8b10717ce855b0ef279383fc89f208833db7cb06487279
z92d7b0db54d81648524713766c6c6584e2e5d58c0382be1ceb5d02b8f2c0729a2660d53213e7b9
z44137ca5e998a861f26d1dd076103241fc53c57f6b0c04d292ed4e524680a58e49afbacc17b9ec
z6f6030cecf4821948ceeffb38c01f0ab344a7a2ab288b1718e30f0d9ff8352b77dba23e149013a
z321c79676456f97b121159675a6779cf8dcb734f87985d832aec017549d6687a026e4be120da42
z9f1e39c215aee6435f2d0bd1aa2988067b3c7830b977c1085c7516a885c616ae9552322dd97db4
z9382b7e3481a3bbc29cba5dfe3d5869352feb036f6ab32ac307cc0febb90ea985928e79630e4c5
z94ed61ace5d89594803d6ce17c2f8cb0d730787837c1934824e5c3182d15f274c9897b63075575
z3cb3bc800c4388b30ed86ee6e8fb69bcfe38423f40b334c70a76249a5f2cbc65d264a6d3e5152a
z17f75883e60da4fe91dc77ee28b71562d24582bc7a5deeafbb31e3ec1e46787dd1635db49d90cb
zd915489ac9b34f99647e801fbbda8a36ac452a52da60b72e372610fa614244901d7a783e86ccba
zb8bb7582b3135e08d668ba261262d1fea3983ff768de9c29ebee2dc3ccab1c12efdaea4621683a
z4b73b1032586b341839a08272d5536512555292757d9ce8dcd283a5ac0610012bdd523d8a4bbde
zb28d38daba7abdb6815cf830638fcd4dfb6a6079bee461f5b7968465964db28701aedda5838813
zc5963bccd1113d696088f4d467a8d241c5d1cb09a12039a79aaa63b9691534fd0357b7992cf029
zecffb3f864563110c1bff086ce797c98ecdcc83e8ac21a4b041dcbec5d665eca858706fb681cba
z9240fd642ae86a081900c4c2c74d20e99c862f80894af2840547e47e4b2666fc0a41625432bacd
z0d8d660bdc4d0b8f682bef5e9fcd0653569d1e2ed1d706b4ae932e615e97f95e4b388a6f23786e
z1064751da9f0545dd0163a3abe6df814e28277c3289cd39cb121d8c4c8fda0f7b06d9f9f3437e6
z66fc339927e9189ab86971c6c9ba4d1761f43a15d49341a211887b8affeaa7da8e08410caf7634
z020e77748a381009fc84afafe23ecd172188f383c4591bb7cc3466d6f636ab9bcf51414261ca0f
z33fbc8e8df8b597f28c9bc0dba6468908f3b84d2245d831ebb666e2e469ce123c96001665bb147
z457b7bcdd3575d1aeead370e2967a93b11e3d203bc4ac13907acc641f9a9066b71fbbb8a931208
zc03b83505d7a0ea85c7dcf883bf28b546a6817d3ee8e91696397532e3dfa05e4c52e80c129ebae
z80d7313b1fb662c82abd9d573b7ee02ecff69cbaf0fe1dcedc9961b0e3210cde599538f1e59504
z52d7068212b469fd9c75b1dc1064f092b9e41636847db21f18037e5d8b2f0b1cbf285e88313f39
zf22b0a1e534ee3ad234dd657d3e252198432b83c8bc9688d77f6626da6b4b300bcf317d8953bef
zcb9ce8e3cab56748ee5623d7ed2a52136a754574ebf956a71ba727cdb8dbc152b8be5edafe41eb
z127e0b67f18280c92adcab61e0d02930755b12b5c8ff3af6e19b85beb1f4f03bf5640450e26326
z0e1cb1c365b6c5f54969c7857545cadf3beb1ea24f37f97b1408f2955d1770344d7e3a73da9be7
za52979bb0fb7c156c9bbd327983db217dda10c47f200a46295c91f633e97c8a0dc715aeb02bc6e
z5cb17a505fff376b433dea67898906a99fa5f55e2f8b84ffbc7666515e3620d6ad149e9a17c78e
z739df194545d9507207fd5a3be07ffa64455678d8786712475ad07c93974ed51970d7acafaa004
z67eb5a2c92da88b33d03c1baa34bfb59caba62f834b8b9406a72c438aa0afc21b74d7466c13a4c
zf8b2c6e2a0a619f76bf1b0b63b0097e5dcefa6a2ca9f9825f11d23c2c23ede29ea5d6cfecb2cf2
z4558360caefb2a1f0d4b4e80d4e355fd2ef9cbadadb74bec39fe300168cefdb47eb4e8508f6fc4
z143b78847e805e45b12d270d35e4dbcbca4533736f37a1d6af1f5ffe5bd81a3f7505bf390a229a
z49c08eb1a328c7b90d8cc6ce8fa0b1f306145f0c11b7949faed730e3da003e7d05774687d8573b
z61cc6d21aae28a1ed2c0c11bf1cacdcc960f229b0942b028396bb430a81792fb84d036a866cbd2
ze17e11d99a6d72f2ee048c19b74b61109ed94a3b8b76f0c13f2ec4b4b049d65d3583781f5ccf12
za69d48f4479b76ad1f07fbe3c7303d162e94899187040feb035c58e4b9851547166d173ecc58a1
z5fb54fd34cf8cc577d00f6b03842b4ed63d973fb5d3a3ff8a2eb5cd9468f528d6f93cdca16198f
z635835f726b0123057c346edd68ed7765a16fff8e1452b95ebcb6dcf61bc28300573f703d8a6b4
z03be2da232bc1a7492a0dda17fea2c691090e37a69b18200c131322d846002d750aaa3848da267
z4b8034e1c886ba6ab28785347e96a97270bdd9835e472037c540d271a118e8ae520b70b317e8da
z3a790402bc283a63203125b7080633650a8439e1bb6c2c628f82c19a1f0763b30825c17374b8d8
z366e9c3f5865fee6d2271ac86f7ef2713080257193c44fac85bcfae5fbbef1b5277156fd379597
z41326facf56a73cbb272f664ec572fa3025aa579266dd77832d13a7299b6e540d620108e6ab61f
z402b745df6e1f8ed70fe294a832a30148ee3e7e2681d756fc1567487e6fa1665918c6fb5afeb4f
z06efdc95e5c57796ce4d683c8689d1ad8199e5b3cce69fb22a65c3e455431e3c7a0c0b44f8fc3c
z8b388c8fa1a572841cf1fc3fc5d69f43e0fcfcade1338e8e94e7018afd23bbb8cf50cad0f44cf3
zd9c51b80bac7be8855205e3dc9d391771766f72cc8ca0c4539c885ff61f4151cf8254e759a427e
zc78dd417ec51bab43bd044c27d8a33f2878f33b945dc5d139f8c68a422f8638085ff97026651ca
z3a1a2baa6de4c9ad9e15684469620d2c12c9e5c207bc1fb9f585a4527c989825bada08a7e67507
ze6078292881aa9e742f7e4c830b284fb0dcba97a520caa714c0fa7cf02a6506c1f9208471ba3a6
z74da0e375c5a2e4ee7d9035443221e23fd9bc25a2d12e55ac3711c8d5f513bfa8edccaa32f7e15
z0f2858711d21c93fac5155a3242748c16b7ccd82e981d8b5b82b98d64d33ff694942b61ea935d3
z9d32d19430ceeb55124a0c96bd5b0cd674e9c00fdd02526aee2d1a07573fee3f84c3e8b5216f4c
z8523c723550774849f4f90738510f9ecf08e138012531ab8fb6d25db108ade9afaeb96308bda53
z5446dc230c731c189f61b6edcc83df9c20742ae2faae69bb6534de659e3dddece268a0c34aa81b
z4cbf4581ba9ff3e3e3a5c84d4a8510e320632fd8fed26b8b214ef2cf320f96fbb1bf9fbccfb4e6
z1f53b43ef2ca11b2d12e16936efd0251824864ddc90ee021e345e4ecb8ba8f39f7ae723777ae24
zf92cdc1b0209b081f8932450270c977213a06092d1377ff28a98ebd91ab616a0340d9d3ed69a4b
z1e0e4e00202db14fa5678481b1f0665dd929bfbeddbbee5768b8bb2aff818018d533fa0017c878
z569890932777634e0f59bca39c3217c9b5624eef87b09cde4028aba3442d4bc8abd21e7a35486a
z5551997fabed27e3b04c8818d6ef903dae2a081c1180b2af5ec59906587ce119dc988ce0b442c6
z6194a28332800c59ee7ff561885a208f536f7f924a4f5ef9e5817358cd8caae8ae2eca37552726
z63d25b04c02250ce2602b1dfc9bed2ac0cde71b469903c45768f1f5b2339dda851541ed933ddef
z76213ca290e8cb1cb6c6c34dca2ff98ec12ecf2aee925aba5c65af5707777d19b4b341207b0833
z2a3cd50b00da058f11a00bcc2fe649e718defc0f6ff834e8d485441c58b89d64e85c5b56124c0e
zec70e69cab5ff3021698b7593c4575fd917ff8f34333a8d1d92b95fb4bd303eb7043b1680b08a3
z90278ea7e3f1acbde561b89cea77ed987819267192af4bb5b463bf03f957b65fe4764ddd9aa4b6
z99cbc3281a0377b10d67d7a3e0add28eda47382aa53088cba258ccd0e91ea1fefc648df88a6c3d
ze1ea1942377e2784012463ea6542aa82de7ed6eca29de9467f885af0ec69a05567fa2dbd1c585a
z7ee749437d1f7028595d095ccc57b3daf7510023c270f45b6720d6d4c73fa6a3dc9dfa964fff85
z51500bfe7def8ec135a530a9318174eeb9cc56116bcf0aea1d8029ba669756eec4002a1b1fe747
zdf69f28f2e9533aaf0e5e97247404d98c38c1404c81246b2b8c94f86129829f9d81c733b89e2b6
za919db3d1987b99aab65f581edbc44c70c4986b3690efee930b9982e0f48e45dd5e4c5f99d0375
za82bba7ec35205868b9913bdc52678468248348c0acdefc7bc2945ea1497818074f3347d5b00f4
zc04d18c34e606c1f5d99d9194b6d6314de8d764ad9f84f705fb3ce7ee070600e06732523d7169e
z5f4eba2495c1d0cb0ce971b7e70ad0b469c4a38a83f90299cbceca176547527ba45c1ac45f3317
za7e97618b863598dffaa3c0e077c81eb1f6b3fbb86d19cff7ec3bd57570a1169420dd8799ebdfe
zef7e4cd318b46082a4bbd8f777181da071448efe4631f0b3e282fcf2a140a2304e7a85172f54bb
z3b46e1bf638e220e162e659d2eb52a63f5d50629bda77b57cca01097f7df71318b7b2757fd128e
z247679430b3a16d03039ebac2e842a0d528577da57646fafe088df3ae232425b6329648137e611
z0eed575dfe0f1730ee76688de0921ac47b90a11ce815f33fd966178b8f7666f3451c1a07961e81
z77453aeed337bdf12a272e9082f90aae5f154852c4c86b9caece9034469f3a823c01acd876c7a8
z3023dbe9a341c36e1c8a29e5c371587a0b86987d2f2df267cc52f1d176e6463654d3d9d4fefd68
zaacb809535e4527a2cbe56d51ec7beea1715402106b1624e699fe693cc4982ec9fc11e63c4d78e
zefa5fb883fd12bf45de4e6016931a9413446441102264baea37c3136151b24be340fd5cb5ee006
z0ed09fedb64013bbbf5b968508129dff23921724fa95674433f5d8726f4c6db1bd5034b4406910
zd2bf8ce46ee390477dffeb406d81eb15665b8198a229ae10073333c154952752ef9d2506df7dd0
z0b1a2226b7596512cfe5e0a83f9315f91884cc15f81b29cfb0a049e7f3482595c58c4d51c21d5e
z0495a0249835f13b8795b2c40d4f5951a8c0b653985692dd1f820b78142b0d00c23ed25275ab7e
z745f6918a1e3290fa7731ff18466ca8068a3489a327b743385767e66d5134aeb8842f974a16af9
z1abaae949798f3230a906beec347e304ccf1213ba42dcdf519cc0a150a5d86cbd74b293fc5c0bc
zdd359e606eb14cbad49644a0907e3301880d682e4d5981df948c3c04740a1369719a5c4dcfdbd9
z5bfb18d1f6f8bd7100c0767f7e22a9b3d4eee8319455cdee34bda7e65e25c40cda410a9dcf0f42
z7f18d6e2720395a2400c3c88d78544d6c051095b4b999b27ba04ece67e0fdf403c056957ebaedb
z199c27f84b0e109e6e626ea7fa28f00185eba1b28e90d2b5bf0b43b7f2989b776c31784fe7d5f5
z4d7889ce25cda576d3e6499690592f3df3f0c85195f74b09333bba1bf4ae6d9b28c8b810ebba52
ze8b626383c40cace06c3ded50b17a565f9bf8cda7a49009ad0d54c008f6620d478c8eb5ce5a54a
z87747ae97e47e00d6e472b791fd661563ef72dd62c11190b2b62a17fb73ed71daa0a59e6a57f32
zd246d9371c7b1845a296171fc7c2f3e0ddfe4a47dc893e6cd835485858e5c645d4b043bb851b75
ze8edd7aed1fe5818b64ad01e756cdfbac3460101e960c2bf1a355692936225a209597e5302f631
zf4bc1f6bd4b459830bdf2eb6aaeda664a52959f9523b9dedea81e57dce330438c49676fe6ba1e8
z208738ab0fff228f57e6ef22676d6ce512aa4ebe3a6dd46d80d7af3482dff63bfcd948c8e9ac79
z487d81a2a22ba24fbb89b2f087d45cfaf4014b9a327ba679b01b6cb6567651f0bea39a7debba7a
z85f834ff283cc093cfccc703a99d3d60720a3ab7dd18773b402bf88b897bdf1d7d5c02d5cbb182
z0ff4dd4ee9fce2702ed311cb7446edf097171a7607f042a52e43b5a087bfe39d5d5df83170fee4
z2769228d35126233e6814a046b5f81dc1b70aec7b25e882c45981354c07faf58187938217a554e
z1734f7a26035282da91f08f027d4c5843b12d451c87baea7e4b3535fd3638c1500cd983d7e3f59
z8739890ac196866a89b4a70d92be8073febb2a227bf67090b31dfe8209eff54e625a3b264074c9
z12c30bda89cff4cee07caac5fc4774eba9674b208ebf4650ec4d9aa18675f3d10378f447884d44
zd3468e1c9fada2c884692fbcbb935b1ceeca36e377e5a39fab77413799e7a2995015aeac9225e9
z5b53c3b7b8ffd2588707d12fa8f9f02de8a33c405cbbf06f5766388e5f44ddd5d286f4bbec6b90
zb36929abcf6eedc273fd0198d322989007e82c236e60e18edca8c2adf91c0089d45f11d614182e
z3b4500ef52d6f5dbef2b4907ceea49c6f9fcabcded59e2d5147782adae7bdae44554d2c4c27eed
z4a2cc6e75039e06c7e09bf89bd66bad44ba4a88cb1c4a71160b52fbfe0d990ca4d7d8400059436
z2669ffeae9948b175c1ed991ea152c4f0767d04e8fe8f25b3cdff24c6a97589cc4b86df4f03ca2
zfdcf1018b21a48277a90bce94a748e2eb4e606b85d2105ac3a7971aeca77caecd13400fe39bded
z67b961251bb4267651354644a1eb6997afcbee39e1b6eed6aaa0d7149efaa74e20e9aad5b40e0a
z34819b94ec00bf4543d093a08ce399f222bb3271fbea81294eaecef6506b8bec59df57960fdb11
z087906bef338783fd58babfacf243ea04085bc77718b8a783d5111ff14999baef4ddd69e3b5f98
z489648f1d0fbbf36109055c1a29674bfc66bb36ac673f1cf7693e98c65a4d2be27ff07985d0ce0
z047ad9686af3044a02d234d1f8127046311e711c14fb4321e0a6b74132ea90733396b7cd4f431c
z00d13e053977619826aaba56f7536aa0ce7be34977b968b8c1151b77cb1aed0bcf210a62198721
zecb00a4d4500880b3f6afd728e053eb7588af7eb068398b59bdf693cea6f2bfed1c891058fe41c
z0118e5a6770abad721b94032dd306c1f98a8b67598a021bcf4ee571f6ba41871787034d24b84a8
z75fedbe7b441d99d2ed3b3f7f70230856bc0d0a64c3b06426af13cf5b9ff6c3257a0bd072befe4
z0d2e70ebf8777c58fa2eaa891c029c82e0dc238f6c3842a27b9617fe775785bd3e2e3cefb1ce29
z6ef150f39f95d9ae09f0b7888c8698ab24cadd6e975743b1659ce0aceeb9c434385adc2407255b
zd43fe0c5b9b6bdd742ad61704f4f4c28fe97e629d64938fbdb3458acd154974e52174ab3742796
z99af0784726bb486363cc075eb183f5360bd59da866d467786eb75f1e91709fb0ea0c23ff12326
zee4a13ac601f51ce95a91647748ae0851c5bab70b42b9223c0a11ff10eafff0564fa22a1b90bb8
zdab6bfe83e71c934ed8b44b2bf192814feaefbf1578952465db8672aa804c2cde3abdf0c32c50d
z055fdff4cd52d627a99b4215f97bcb9d73be0a48c9cadc95e398d68727dedb6c32814f762fcc68
z5f0b0e5e5e6a9ee858e1f01914f862529a7dc71ba079222bcd8400d2452fef06474652c1d94116
z66d6b41282894b8b07514196d7833bcd2627d0e2ea78f3d64e3d51f708cf23b971e737996e3c8a
zd3751a701aa5a7bd7fba1773aacaef6f7d5729e08c2c6bc02016bc4826148e43f8983a3ad6c63e
z01d33072c1b4f198902f9355f0a25b169c18dfe9bd59320c021b7a38e07f60b43a5c159f826e56
z61002b87ff1138afa9bc6df7ea1756e39bcb86ca826f30f8fcca098b7ebf0790e2fdf317e433ab
z1c2caac96de43bd581a6e9b2a265f9471248ef40baae681ad28b2c6eb4df9ca2cd9f975e421f5e
z76b455dcb42d487d29148851d02217044b272ad4a00fd7ee9d77313bcd3e237176567c06614d52
z881a198518dee0cf9aace0b298af8f9ca54badd50c775a2b4720407467adeb4b9809fa1a85021c
zc1fd602c522afddd5c896f8a099bd4065b4fa3e8865d986d84ce03293de4b5cf04cc075adcbae9
ze5e4ea0d9f3eae419625ae7c6dade7797e541e567e57cffbae14c0f666b19768858e218dc9df39
zf80f809a743f431fab9c87a6b8d00e162a4a094a52df55e1a40b52f07d19f9e189336fe5e01b70
z55b5e2e65d1021d1482c2fd7c91bac746c5d1735473113bd154da1266b33e0c4c2bd3e9ce0976a
z5cc5b30b482d7b2554b714acc5afc1f9bcadd537d6bdb1943c75656e4dd741a35acb86e9f886b4
z313c5b6d094521e90af333d9786f246b4fb6c22ea6f678a7c32aa6748b91f8a6290290262eb502
z38e17889e3779d3d5a77427a715fb5c0e3ef5c8d423cd9efb00d5021690041a3ae0609e8578229
zd7dc55d67d1b4d4aba42563ba45e7279057c17148d3e90378ba7b68a88a6383b0888bfdbe7b109
z405ac9e327faa113ccc3b1dc34d751672bdaf9dcbd0341602fd7f8b7e2911980bd02601ff3eff7
z9528c6a2e5320e3d4e33aba8de93622de14270977dd65f1513237a86540d8c526452f851e2d140
z36c13b58e4ad7c7b6145099d6e643fb0ba94de5d052819af3ab8216aaf85b9e9701449f909d806
zb647a41c9aa0fd9fdb3a1bea5f3aeba18a50cd65551f5d5be9dc4b03efe4534215ca47aa84aa07
zc1a50b0fce3875d6140c8c2c74b19cad88f84ae81e34f3ef96c9056740906e66aa6e6ad81a39a5
z31d8bf7784b813abe91f45d0a6322d8aa5c6364dde4e424e105d621877895d784a0c439429abe2
z6a27804fc4db30dd662beafb1db54830f372517aa4fd95eba799c20b3a8c620a893eb33a24ca6a
z67f7cb8c545a5ced479e3667e3fdf579bb458c893d42ca097a0165afce88079dafab5d8efd46e0
zf81ea54474c1909096bbb2b68a4b4dd9af75338f607e4fc28e733a4e8a39f77ff40dda1618ff5e
z6d5b833b0eb5096ef1f6bb4bf6336dd49a6cccef0ce547b2b4dc5f7d84f018f3457aedd32b9f9e
z1e01f1437588ca4f190cbb4086a1cfafe3cdfbcdf0459349eec551c3094cd4460dd48da8deb412
zc6df45b67b359196e937cff77e15d3449a207419e09a1facfda6293a80686eb76692d46c7bd826
z62437ecae8b8a3580cf27059fb2841183bb685433acd946e7c03f137abd18e08142eb767c3db19
zb5b68d50ef74c389a565c0c75b057f5c21060127eaa746e6a3bf702d507db130f3f637a976192f
z0d1d1436481b592e3a276cb7d78b8f944d85fcf14652a82a4ac9ca44855a0b9ed42030f661edaa
ze36f62593e796512dded7bb429c94003c89ae9d6e532e1b21a25565b0dcf589e27f1292da19f8a
z09cc21ba696a3c4843be8578ab6ccedca049aec6d0a41e1666fa78c0ee77cf583572322e67e4d9
zbd14b1a7d669251f09cbb03e7cea9c96da1171c0ca3f1144d881301be8f2a0b90c5fb87cee1b42
zbdb7bd9c010c12d2e0750b7501eeb5597c58dc32c7a16761cb4ed74412551b5f7eb05a7c69c130
zf5e4bc83a2c5d7e19de491e7b3c1aa09d80b67aa5006f286bdd1eba17c83d3ca4026f65c618020
zc4204b1c08f2e9f9dc44e450b2914dee3974e54855bb6e2202abe60321a8a3da417d953ab28fb0
z340232b840c1f369dd0145bab3522398b3ff9a44c795b1fb3cc57a5c223b1944379434edf9f37d
z23726c1308cdf0e86f9b603b11f2248cc78dd58de48c5abecd10876e3976136eb3c31c42edae11
z5e27ccce4e112511bd35ccf779b5fdc720de28299e05afb5755e962daf57bb0526ba7349ac5cdc
z6a8ba34fa0b5daaa50b1043033c426af093e3dc0d57aaea2fa47fd9a44b14de9d67e1ff50c6a8b
z0af772d0323534e4cee5c1a5c0b91b3f1be1a9d05a216952e0d66cb33f012f4757d4bfc59950a3
z2e90e02c54568fff901efa39e2ae08d170533b5762a94fdf6b5ba2604c11636bbb18baff2387b7
z12e567b2ad7391c0facadcb7d356651377b51f4a5e71257bdc5b417747cb374265d99863504b0b
z3206fe598f4c4a4e29091a1ba1a90d82222ee93c6fac49e0f3acf6c82e0f78d0e7c1dfe9662e5f
ze6c759f350c0f9ceee622bf55acd2dc068c493b95970a2cd1020d75b7f7e4b9b0438c2ae7ec759
z1c6344fdaf14a771f9542134efde0defdbc8689073f0d7e01e0472dc87de1ec2dea18284b009ee
z20f79b0225b8e9d139eca2184dcb1fd045074a91a0841f55cd57c4bb8b0d3f1ef008248ce64078
z4d393d63e45367124c3df2ca36ec5f5aaa944a6bd295abffb6f0bdfad58726f834cea38b206411
z2f5dc8847faa271ce84640eb82ef1bafc6f8408dd972d2c979613e5aa2fa1bf2f5f79bfa7494e9
z06cba42dec644273f1daa8da4a3a83f026ddbe727430bd962fbe6ddb8ccb0e63c92147f5b13e07
z7e754e7186de823bb13a41efa2ee6f2d2e747f31620a1b1ac2ddc600fa2eed6de0c77b5a98cbbe
za89f81475aa2c7bb850a5384ddab0eeecba52c33be60b628f33787efffe9589501bb5ff7033c3e
z21559d564d859bd5cbac7c673b9eef6e0d53925a8f08d786670adbe0cd51e37222189826f67dd9
zf228d512e4dc912834def34dfbba6a929798c978939733ef70c7b0d5fd7de6ce0527083f955f00
zd7e426eac743579a0cbfd1ca47f113d647973c8e745ab50abc9dd96acd27f9cae185d871817fb1
z7b78fe488e1593af90634975c26eabff7ce1c575abed02f1b2ae1574ff2ff63f1af69e9b23fb38
ze1178ffd9f5a0816b208356021f525786bc24ff32b4892a860d68728350e1aedba33e62c6fc0ed
z1c4b3cb5f0b536fe5fedb5cb3b9bd94873fdf01d2657793edf7da7dac537e74ff945e43459e627
z4bd47af03d1e2d7eedd2fb7a97e2731ff65c3cb704d5426e8d79938992f2c9f72fd934daffdd41
z45ba345a01736dfdcd5ecf9e06ac5056a415ba3c4eb7cd408b28540f334a6516e92e3e1b809e78
z20bd153d0284ad897b3aa411050236e6d140141a554464f7a97ed9fc45782b983df04e6ad44d49
z774bc2414bc0c6e1f8ecb512fff091be8421dfa835a4f55041a86122901b6412a61ea4acf835ae
zd7ba9debb0b3bdcdcc71331ba1711e5bca49955d2d6829e36bb4628f4d517243f7f35e123c4857
zbe1234268093a99181003d90333920eb919c4a3349a4ac5a80d6b890f973879e32e21418026482
z1f5ce5b01f1764bde66416e30820aac24c1d06dd99a44f42c6586585e6cd569c46f69822ea124d
z56c9e3c84116aa4f13257070b8f490e29ed00a6cfc426d4170fb2a32c50f60f51f856c6c939e24
z4a446c088771af42b57ccc55f1e25225e0ae2c8c08f350eb0f258fecc266150cb808a7b1afd63f
z2124bd0c9d33ab1d9693da8e357e7fe25e4072fbb1f0b0abac99a1302101071d2688d3538a8f72
z81f03dfbe0602470d08f3f8a244448ae09bc781a84d2064f13c5b17649afd66916bf1d97a8c63c
z9e46c6645379798cbf35460443b326b2871563226efdb537d7edc3adc0878473dc9d1d520ec4e1
z086142871343c60960b69505aa8646fb19434e78b4205bfdb7d75e931b14e1a598412a15a842e1
zba21eb40a1213da497dc62329dfdc7f0641a35d36b57a7da93455c3180e2e585cd7fccbf959447
z2107e9feaa04bd263912b4924b20b611544cea9c5a4529f38af5ab2794d16fc67e7e7bcfe121f6
z4b93e350bbded4892b8284035b1e2c28a89d712a39236a9e5fbe8091f20afea85ac11ad4584a87
z4207b1f3d97ea535cace52dc82b58c6f7af78f6b2f2521d6e19f298ed3a56603d036b0db9eb777
z636994e8d1e31d77aa421dd44f0a273e2c0609d6708028c607744e03047a3965dba918b6649057
z643f8844530cfc247d824d07c5351eb4a581fc75b1c97fefcbe260cf83f55ad61a910aac5f65ee
z8976de932033c07fce376b1bba00cfe04d0ca791dff33033050b428efcfbdec8ce9f3250bebfaa
z6c4b281bd01afd3d7b92c4de061434836810a2d27c2d41b8d749cee5c2438140bd840936732544
za14b27e0f01c3b6c39bba64a5f4fcdf84f20f9abc10dbee3b02bc252f6edc9f7dd38d995fb61bd
z613b475112224d9d4a75490109ff74a2c667ab701ed9e08f19027c96aeba8ff94ae74056dfaa01
zdd30af44c6fb9a88554fa00fdb44993cf066d8c2098904238e8daf8501be8c6cbcff45686ae6ef
z86cf838b6872c9d774762114b40c34a13c79f3e10825c6f5dfbb782d933f23fb4e783e5919236a
zff6660edb48403d90c877acb5396977b89b2db930597b4b794b4ba49f943aae7dd7f73c2ba5e15
z05473abf8ef690f4418e20b0589d151f83b4d7e7812de051a540032464055ef28341f4b6c55f57
z760c9b29942a170dccd36015cadd8b43a174f5d307ac79da1633fce00b7a821d665d4240ae7b81
zd80338e707636e911a3305cff6a3908efe232c5f0a065d6e7cf275d282fc7a988ec251a3561c90
z5a5fdda9f728cd5fac458787a2982b57e89d560b9ef0de367459655b6978a5f82b5bf6e87e28d2
zf9a263394a19c62add0af973099b5ca563b843dabd01798da3b6e8639e6e81bfccd2264b5d055e
zacdb80633ddfe47300022edbcf754e8d25d531fec3bad5143a3c13aba606c87197824d4819d4b7
zab02325ad275219ebedc1cd18a176544363a98eaaf1a456bb880b05d1cb515c2d280b1ddb0ea2b
z9bee6145834f05695e9414a65ae792c236ca672d3ea9fe692a615f77a7f27837c8a43cee363719
zd7ec9608fa7377b305c9a94512694adbe2e0ac763f0956dc592dbf31a802988d4624c9a312ad93
zc54bc905ed6387aff8deb65999c69174b9d88c44efe5bb97813048ceece7836f477cbf3a42355a
z6291b9bb60634144a6f4dd095c9b1d8e63949b74f68c9a9f4485367c3e2e68dd134572cd481b1b
ze467207aa697d7e2dd7d46f9a74d2990c58598d88240fddee4adc74216fea0737b3a19fbf37cb6
z915d803fdffd9ecbd9955587c1c1add49f26944ca9f03a59df72c4eed575a4c756016518c5e19a
z02355efd6a58f90b49796637878a068cc84b06eaa4396ef0e11171671af0a0d858b26f65bda3da
z812c00fb4f80f86611367be04ffd2ed0b69402492ca6d3de41abc4c50a8da6166e28f7c7a1b838
z9b491e8066daf5298750953a3dc5d5d63749c461d4a331db473a9caf3f10afb2f949e3f9b64cd8
z5b0971523e9ad87806cd2c4a709ae5be38fa0a97f0bf9bf1e484a4085574e831fe7a347b2344fd
zec2045b5058b8d04190ffb8eb1e02c4fd10722059da2a15b1c69904229cb5fdc77efa0939744cf
z70d6645751f29f9f445bd43fdaf437743fa7f64d8eedb9b82a95b40b69afce71052b3bb059e7eb
z86ec49bd7181e9d8971835c81ed93e44bcac89040beba2cb1d40c6a87e77b8896182dcf4e19d21
z3f72ee1ecccb3c2fb8d6eb1edc26ce93a62f850f6318b6c61cc7a2c8d2dd5452d850faab79a2d5
ze9e55d91e0ddc76056b4a2f02fdd1b89c577d54008429dbf62f729c220b6bf2efc5edbb5e312b8
zd588ce9681977c8221ff64f10007038409e341d949ea0f2334f5e536febe89a24531f225a3d9ec
z0a1f5f6fbda73243924d615b500249cf3365a70153bcd4c737fec1dc85e01fcb788ceffdc8ad9c
ze731bc770e024b69331d46c036f29f35fbe0ce1ca7feb5f9619c2f808d87be5cb9e6df1fba59b2
zae558cdfb66545eec2cca530ca99946a6c0e249bdc65d6b7cdfc5e79d1be9c5962cc6851f9f42e
zd72aa875593c1db8a79199a6d455705800cabdfb54caef7f1cc0021604d8be352162509be83834
zd8888722244f921d279359e776fd05f558e733faafb517906d3b354fad0dfe77067b83f2d430b0
z86b25a9ac57f869a9e6a73fee14940464e5f51308a7a29479c1724dbebbbe5eac23d87014452b7
z8ef1091238591e7fa1db7ab1e746843daf855307b87107cd05040c003a8fb1219dae95de009a79
zb7efd7b86cae2e53c9199a7c91a9bb71984ebe0c47b72ebe9cdab8ee6266e3601c827b8e3b17f6
za7b77760809a1c8b8495ed96af448cb2504203ca57497bb59cd7dbc171b61c267a4a9c4a445be1
za7a660126ad5d01bd767890253b313d51fc22ed107f88d25e4c2a9437c0ec99f16743a9e6e4724
z1cb29a155de98758c2e46331dc162f2916f5f10d1ea1bd0241171f9f9e92c7eb211e87fda25fae
z7027351e5af5b9294c2f527fbcc1054b46130329d21d1b49043f7945b47fb7db567f62700441cf
z1226d7eb148ec6bf80f8ee6cf4ee04f54827f5129ee80661041f0e7a40c3b017fb3770d8e70a7d
z6c27bb549953b31f2ca56f756a96666fd7a0d684bc8267a1d5f9f2712e1adfee96d7f32d4d6abb
zae4773ce4810997b5cbb80e3986da6edde7649cbcce8687da178000a2e6cec2c1b21cd9e7a2ea6
z01ad61133d29d71c092aad6c871ab257060959ce5577d866f0ceda649015505601a69cdec1b3ae
z723aaadf315ee2e78707f2e3ccdb920e08b67e3ce65f46b58225632c098139b3d4121bf51c58f8
zd27d02a0551344e6ccd3d8ff53dfdb19ccc2a249b28568ea7983094a4151bd3dc3c862921d358e
z53eaee3d21728ca41b2565ec89d73f69f50c3a6d9276e9dc4cb659c3635d2b388c7184e9304479
z14f84b8e965a13e147bc35fa65e4f9d36dc743bcf3f5cff393f9782b9f568a8016365457322122
ze1faf42c361b4715010d5c7c146ee02569811995fd06471f945c5666b9026f9d083fe303c863a3
zc999f43e5b81baee47145277415ed3a0e75f29425636571b0c17e51b4e990514b212c6df3f2047
z06b85fe80ad8e0c25e9507e10baf5f5aed3044b24945e2dc5931d0b7d628ba543c689c53ac4915
ze43f5706cc63484e6432eff228ce7f3384e107a5810331adcdce1e4834154fc18ceb46a54999bc
z912047363bc69b9bd93325115ed712d9d7eac1175ceeb8b0a53245a1fab7c3fe0de3fac61e4650
zc4f696d2a93992b36cf82a6f13a49d719632985d459e36233b6ed80c8f76eba26f7eb7c5309c6d
ze537c160fbe9257fe10086fe07d5762fb568afe4aa3d839ea78c5bbc9762224fb0c0a91465a21a
z8091427313fc673ca8b1b31d286a2ef78d7e12c7f850c82ea1af2814eae15e40e2c404c9157c49
zf5ed5e741de454869deb52af907cdae54057ddcf3fad129337b4d9acb058ccb22509c67228092b
zd56e9a79bd02e4055e49910d01cb0add89d42c0fb9a92084c07e2c080205fe90ea4c8e0eda70a5
zefde1ab01d0926b7ef948fb490d09a252f42fca98100a02ca61ade908c596a44ed124b9a35ad40
zf840d02ee24fbd3e4bb229268f6c95d725b540266be47d18b29703c840417de6692fa2f0aa5c5e
z56a590f95c36901aaabead06fd46988d154488f8e735f3b05b831087967bb25db8667beb598dac
z664066958cd28d6f5e091bd07fd080be91455b45e7cc254f1b5c356750851bd791c17876df6072
zae071c3e72a48abd264bdd3e6ed8853c552ab6079a08e768f3b535fb42b253922abda0a158d317
z8313d246540c3e953927e7de593cee6aa4c807644af43627832b895b1c64e3bd693ab95c24602e
z7b5b177fad6d6464207a45c4c5dc83a34d1449505eee24ad6ba3fa9139b067d6a03869cd2dd5fd
z9660dc66545ed4f1007be2cda93e501ee9d3fdeddcbb0d89aede930b0e4d8089622d6ef703074d
za97aebf092082a8ff388d729660ecccea4c58eb8006202188a11ba24cc7750e99c56536e689bd3
zad10b4eee6814b42a63342692dc7370fd23c073f52f611d113df5b535bf0d24a5a39e29ea170da
zaaa131db19607657562a4b7b48f60d84047dbdc9e80f42378a50802418152bd2ace645d6bf0926
ze58f1e6c3a4f2d834c6be10d6b7b3954577fe6291ac3c597114da8dc39f4099c9739ad5f1a1b4f
ze7f79b8c2611ccd64f9b713e8a85c2cc57b745d75ffb59dded09a5e9d4c270b8dac34050bf5cc2
za99479893eb628f8091c190834f1cc42935487317bacbc1e806551ca0129914b0354ff18318ae4
z80a4e7849908131435cdf3ecc6f81a114f7e30a8d4a814529ecb8db2e52d34cd7ecfafdf8d1edb
zb97ec5975451d1776ffcc9aaca6682ca3b505fe75e1b96c76dbd8e1d85c37c6a3152f1ea3b9038
z1902a5e3cb5607482b57ee44c09204522cac49e08b269534e7f1edfa8a3d1eec32b7a452a1d594
ze2124b167607319d79feafb7153677185812f9ae19805a925d9c7b39aab92a13fe3ad5082f8a03
zf4561f8e2f4e8def77a0dd850c694ba50fe1b3c961059f36a0c220ad8f0aefab05e30e55195aaa
z2ed67aac2103aec50023d0a06369879f1395eaafc16508eb08f0d10ef8f861169d33bb6f94fb1f
z612cf47063317a17b1c5ce0725d945e68be6c40dbc6100a97ba65dfb49f69703a1d1d163aaf3e5
zed5c0639268ca0be8c2d4b543041520ced715c579f7c5c0317f06dcc8fb8bf95f048802bf4e8aa
z15d797fb80cbb673d514b75ee19ea3d309cedc3644b95f9050ed6062f938ea750e4b51082630e9
z37c5b9ef4fb352d77cd55c1780489678395d723dd503dadd334a3586dacb8eb31a3bf52972c134
z044d0d13d7accb351bfb5c020e62a1073626d5de24ac07ded63a67cb0161e84dca324e64952440
z2e24bd2d8539a22eff214e14058fb61186d1aa12fd3697dd810f7f4da3d123cbcbdab7eccbff9a
z9f4a9dc1a24f1b60b1c2fa3d5279646f3448ef029ea047f41fb7de4f1af4a0f63ac690605f4def
z6c18d39277a44351a5ef1da2a73b737cc06369a45030d0dae1686ee67adf45310cb3047aa4a620
zc032954c7be59a27c653bd2e1b4879f5f91167aadae826ae02941e5f8685ab8e0eef7d3e8d7319
z7a50f487acf4a0d36c3866b45fb59b782b1479c104780196ddff93eef137c9765f21c60939ea1d
zeb199d49618ea2a3524ccbdc1ea990c213bea7d57b23173d5744c997a8f1c13d1e69168051ff3a
zda0a116813252e304d23317c6d2be2e00567d11c40f75c688d39f50999a39aafaffe56e8518df8
z778556c4ba41ad9c8d7db50d6806519b7144d9362a4e22abe6857ef8a060d67ee41c85b86ade66
z00dd1e12f3fe0d5ee0738a5fbfa2220ce07628054f1767557653856b3b6e34c522e7c102798693
zc361336283c818887df80d9982c4aeb66eb80c03453a06dd09a667b1b1e378ca699412777afafa
zef1ba718306d9b832f08dc2d52b21faa659fc793db14bf3a570dd5efb3a1be664b48fc2f105ba5
z032dfda36a7dacbb502b401f06bb1a2a89050e2b6a486b058381db2f19e0ab48dafff911aeb2c5
zfa8fec323ec3272b11f17c2282e7abbb55f851d3439129096fc049ecfc1ff55289dc133de6c6da
zd5b3289618afc9d0eec17606a5a764d59cbdb30d3903297a3ef610e388652050d17dfeb30d452f
zc80aca0d9c5835016a411caff6f45626e0535e81aca77a907d42288c1112451a6903b104915c5c
ze222a02164fe5309919fb5e8f6c379bd3b653161b7859b5f7ea3ca4501822178e7c28f634b5355
z5cb7256b239ebf664fff80ec385a727b86da868c59d689e772ab7b005151db662b3b9fbd7cb217
zf75538ac13b4346270220ffe261e2876e47d974abc412ddb0f6084efac976c171cdc5e0192f3bf
z36ddf5f993b3eb651d1fb8ab972e46147213197b0c77841cc3de2d930aa1c8571e9427a689ef96
z495d916ce50815e9449d4ad0fa946c4e5171da21bbc9c105be6e0b115cbc1252a8242c30f62342
z542445643fa3682099d0328aa566984944432407fa34a5984a0f7978ccc5f475db5482214f5163
zfa636a01f70039bcec960702c1b19402ec080b91ee3caebe11ec1514bce16409af136664005936
zc5bba4014cb9cecff867d29b50e28e39892837e49b3b050f57eba29d6940f34390501af3490fa6
zb0354cb25bb776f0a348e59f7038ab0b33098e582a774756cb42f2cb004233736a820105ba8797
z9b2510ad64e0f2df53c7c55173eadf419d4454598bb2c2bd14fd711df94d5af359f0631c75cdd1
za6689ffba358c9b07b690b2711790634d4f2a983922a3d94f2debdd5de2a8416895847443c303d
zc39c2cc1f7f713d34d6d495995aa243669fed4d8820d6daa815a259780408e245839b4e7d27555
z24e02b5aa1e4b483d70f77935e9f4587002672c54223f7534eeaff2a733044529b986fce31ebef
zb2313f60a822a8cd7538a35ca9df174c649d625dfb4314e46f8f065ee0976bd691a555b929dfcb
z1fc6063e5192b767fed86967e408d3e7a50112dcc6a65445624dd15c831111dc3fa4f3e18be0c0
zd70274b8392a5cb88ed1c02cf8c29bb75407b7e99905eae8b128c519234a0111362c9ff322793a
z02414f383fd579c843eb7885e8e5d385d61bcc92fb24f021a55f4dc2308b88bebe79aaed9f10c0
z067a132567d755334456ac89c6f07c79f45148a67c065499999cd81d2b4b0109596049e350abad
z68f58ad568fdf18d280bf6feaed6f5de2c7e1e97c2a2e18a190000703677c63adac13ab1409731
zfbc416d67d07e2d92c6eb7c5b50b370e40681f4770c4c461ead878f97cdd8ce11c23e964131de8
z165e8deac6b17dd0519b3d5869f3486ae85149e57ce709b7fb0328f26719b715b21871a1cc7745
zd8adc5aa88109ce29636077e52428a02bb3392767a0e5dead51f803195664a1ed863e0bf1991ff
z57c1045c8d7f48b7b07e52acd1ca6360cddaaa7c143f30eeb17c4c4a81673b8501fffa5abd8426
zd1d1671010eb86f5313ae7d5507ad7a06305a4bfd0386c8af0fc003dc47aaa254f73297d7ba6e1
z5e78894d631426149cde8a3075ee726e6188e4771bd6007e77ebd1fb40991d89f29949b433b5a3
z56f75d1fd66b5d60d72a18cad52948b8fed023c9666414581cc8d3458cdb861d8e7c9546a1d805
z378d0500a8079d6fc7868ba8f340707ee50ef819e0e5a94783d92bcd1da1fc351fc5aa5a89d712
z953587e749c9615df8b55cddb66e9bc77179aee3a49549f2a38ad255593711e2221df9ee086022
z916359ac06164fad4a45faa5327ebe8430a8c0d9e991c116f31fd545bbb163e557ff48122f7f4b
zb3e805309d563d6e7dfd236d7d2414a0a2a43dc7b7c88f456fbfa22711a13896f933b6407960ca
zcf77ecb8c7f4aa9b025ca5f9162dca44f9b31f860c836a941505ad975ad1f312a5edb573177bf5
zf41bca5e54348c52539cfcdcb218844c254148efc506866f2b8671f9ae385efe187648f484d81f
z4d96a85350ab8066ece3153f7f9b7a4d6d9e5155cb88d7e13f2bb64cade4cb33c5d67d7ef10a54
z2b568d24054dae95c12b9f8c11a991a01a2130b5c710387f5590edec17f52f074c75382cf3b289
z82cf96d4c80f2a9ef850b9d03af2eca6036b6eab5d8d7da30d90a8fb72a8a0f9e8ce48265c8ed9
z2d111f7b065c036a8cdec94fa0cdce7bc7af883de0660b68342d37f947ff0753331411f0e1ace3
z0286d216d5dd7fcfd0047b4f2235f164249a56647b43cac03643e59ae7df180665e5d5353eef8d
z2ed9ba3cfd5ed5b1d0ff5de1fa68f8f75695d829487ffd56c9646bc9bd7f6e1172983a637cc273
z3130f0221720d53ce9c364fc3cdf447fe8ebd9553ecf1bb9c4bd74a95520d626cfed4ba12fdd7a
zc2c7758afa2882668acf74b69c7706771967102450efbfb35d38187c239b703ae2cef7b26deda7
z1ba92889611e04f54a68c16eed208c6d9fe009e67cb0e3e2b3d62fb376710351d266de2b17ee00
z8bdae587194928320b67252764fad06ae27a08299c13dd351ca68b9c8a7cd1637f3b8148ea1c5f
zbcd3aeaf3f4504d76771e31f577b6d9471fb651c3ec4091ed3ee95237a956658e3e4921b773491
zb5a56e243259b9a2f321731fe59cd2607c58adf84d599976fd2ac499d0b697b091e42523140780
z7b533e5d0da8abc44d2cca2d14dc5fa5daf2c5e1c02b62b52509b295ef67c71e03daee0b697346
z2f9f9c757f4c759d0249726c51417bf2e8b8b117e39bfde54c0f370d4f67bae506cd99fede1fc1
z6c5aa9af034265432c9b48b7f2568a04e5fe00604ca22951f865d9915b23faae30a61d0df4b323
z5e9f5ea552dd88c19e3ea04491eb8de2eee02fce50f4381ec4897ba2d636c89754086880abdc4a
z191446af6d4adcf8914f6896e88d696f51aedeb13272483b1b5affeddc6f7a206c5707e0190b22
zd18eb776604b4ceaa43193e916efba83b64e7031881d8742c33e034cfc398d612a867e11230bb4
z77acf94d56e5a49ec869266f1cba06b6a42cbfe3809d73f434aa34df67b96471224280e606decd
zb5e53e372fe02ac715fc0191e33881655c990b097f3ece6806be1eb1309961e86afeaa12b76a73
z598c42e5cc260d62cc5efda246a21c25407092f4f6bebf98c88c8c5456a83d1976ed57f44bd00b
z316b61132afecc50760a588df550f998b4a67720093309362ded26aadb49a0efc9196de4007579
z6cc3d7eeb059a3dca89c0a652b2f8fa2ba60df82f8385454e5ba4b4d5d39e628500a9da89d71a4
zcaa1e3718ec49442e8ea076f36b8f7ae0245acf4b1abea88326a82bf8e4645ebcd40fabbca6d54
z2f595fbc25c81ca6279973aa5d9bdda13a2191730c525eac20cfa998bd2d9ab358177dccd1ef6e
zc253926d81f3373de19a0d8803c34d64d614a5cbb3a804345cb480d076fefc41746498ee6ca52c
ze5e8ebd97b87bc3beecec5deac4a006f34efe698eb39f6815f84b1da62811ac33e4f37c3b7d1bf
zc85500c73bfdb6050156d3b617eff7cf20cbc8f31ddd62d4b4992d77e1bb5c2ff246843ae4e813
zeb8130e0acfc80e42364e488253b6343183ab7501f2a7f05b06aefc665c3a3313ce6067b2c6e89
z406b151bfc70a66513b6e3e0842d50bcd9b42adb1be79392f6032b00707a84604ba03920049360
zcbad692b88133610b9e6a54d46b20e68d4df320f9182c15e606975c85a95c80d08f599ac1c0706
zbecd935d0546f0880a908bf163ff1a4fbf1ec53043aff406ff08a1b4aa3d9a54afb2cccd7c74ce
z71305e7d07c8c6def11db541c024baa67ef0b2e76a1f4dc632ef6ca7db3aa8cc91cde1d4748dc6
z4c9ae83d46dac0a41047f4b3004cf3b0baf3b826aebd8bb5e4d6e025c6a386cdc1232887911005
z09dd9f32d6345dd6434acbb30880f81fa2f34656a615065bb4dcd85b8d30f2dce80ac7d704f71c
zdd9459dfbb293c81505ed5b797565a2b8b9e9e069abcd830f4782bff7f490ee78d6485f6138090
z79bf5fc5ec9419383e740db019e1e93a166270e02769c96e475c12aae22def034996bba8c296ad
zafb484363cb76756c4b5069883b0331e9237d6f97ac25825dc2aa25f3d706a4e8fb78c43c80373
z4a66ad79d9607ddcea5008d06d447fc0fb7d7c5a7006d6f9d1b975d099e989d82fe5a0151b7aaf
zd6e4b9f37d7a413f3d78ec202949cbc4262075796ac7b83004e31728d51771289b667c65fffd7c
zd5bc8606989e31d4cb20c91dea9338f2d851a61e3f9121d91805d22d59d6bc69655684ac8d6837
zd6d91f0932e266398d4279d2c0a5c27a768b5a06e31ebc7215fb07ee1a15f003319060fa3f4a99
zd57976e88fb4241153a5734cc947f8e52cc1d557b9df3acaaccbb85c5fde22e902af53198d0def
zf6b25a18f541b0572cfdb9533c4309c72612dfe28736e442b6170ea1fc7f1b8dd5744fb32f0df9
z6e3417dc5b4a7c86a262b6f7156069f17d86d1433dcdfbad2de6c35ba3e097a6f2d6c0db2713e9
z1aaa53ca1b268cc1d8b014ffab5fa9f88fa0e48de44cb4a05b86f8f393fc7353deb36098f0ee62
z8513656fc5afdd6820d51f745c93d92343b4d7c28569b4f9e714edc76d5f2c21cf35fe8cd723b4
z801183532c4c5cc2460a8d6c8d2076a03e9c364f1e9aab6d4a39e19e847a9046646679ba6f9965
z10c4b8cde868d49df1c00c55bc253b8f36b4e7ee3795252a760274c77601d3d2efbd41a1fa5d8c
z4e2707a1474a47985bf02ea1fb627fb1ef260fabb2d887ea3aee394ad532442f81408fada0e1ef
zc5b0572612ecd57094dc5d30f70596b49fc5e1d7fb7f164649f4674b675396792a81993009845b
zfc05da11a2e7297241e90a8013634f8b1f8ee2be6794a09f4c31f52b1a34c8f29c3782553a3ddb
ze22f116b19c830a74a585945e19c16cb4a297b00999ae92027011993cca88ef3d6f641d12abd75
zb1bef49d12cd4a552991f4ec4fcb7df4a84fca3d2ef69ea7631964bd01d0db1c8637d4facd3a61
z0fb3097434a5732089a62e396702deac7ccb50dc52a2d31d74fce9c54278eb079bcca8ef8301f6
za522ffbd985ea5a616d16e84a1878e828d801d4856525495a4833fb08223b888246ce99b78064e
zbfc5953bf30fc53535927a0645a912b78d95adb3bdb997664679c739fad36680e4ef6278a1c04b
z0587e229c9e8be11713f66c7c16015780c51a3a10c19429581f1a8d28acd32e6686621b829de60
z69454e63c6eaab0e7288b14ecef8cd4f0a904738960705b85c1a3da73403826fc3304c8abb44c9
zd6b92d0757e402e8683b81882e7fa95acc348558892cd172f45a476eb8b6b9fedb9903cce1b897
z9a13b148ea0a90bb87c475f84bcb6969e39a96366030a2696d901e0a436063ba8980ee8eb5abe7
z76952fcfcd9465cf42aa5b2be688cdfb72e3a30a08dcb62a1b1c9a222eb2302bd3efa30771fa03
zaa237f12c10092dbdbdbee84fc0c9cf28627e1f90b4955954ef01f5e50f00040376c253e8d6d62
z829ff39774c71ae34068cd5ddd9b17b40319b6b042e2a3795a617c397dc42ba3feae25765ae1f1
ze1a937edcd888c8a193f77bd666778116ee68a9b1bbb1199968f5c4c459bc77edf47138d672ab1
z03fcd393a1c5799441027f457c2689f08bcb4a338304682ac16093f1bcefd92b4ff07ed77047c7
z068ebd044f2224771e947b1f70f73bdd6ccd6241dae2d5dde08b9d9bc7f4df9d2dacdc8e450a62
zce0d5c21d41eb6b5187c5ac15d061e0bf8a9de9539c2280b9c4a9e1c2811808e01f1eb4fd6ca54
zf3c2f1026ab2dcc995dae081bf4f63bd41d6560025c9d0b3f63ad55cc5cc4045cc0121f7108672
z849c26655a10e04b8f2f73c701dbdb217a6b82c9a1eee7cd71f348358b28e565bf813ee731c696
zaae76c0c213c15cab28cad731409c9b4ab6a24b429e7474664ba13d29e31a7975007539feb04ac
z30f676e6608b6ecd0fc030b3de600344da37baff3e77eca90ec5cc5067a2ad201a6f1bb568ce87
zd5d5b4a2a5b4616178168cf39a2d9a10b25ce240a00a171ebf516d6cca34283f035297c8b5dcca
z6a6cead804af3167c8ec6529ecd13658f415eceb8da62ccf4584409ef8dd7e6aa3b0909fb5b40d
z160281420e968fbe67c53849781526d82ff18712b93ef8d006d6a04db8b7683903429dc7adf788
z7c505d2ff3133a44a1576c6c928fd929ea1a69620902d44e247d823ebe14d95e84641580259b05
z3579d1665134cc92ecdf5e3f3089439f4121c7b03de2678f23b9557dab8007d962b61bcfe35b16
zece059b62c25784f9e13291aecfced4fe839bb1ed72de9bbd3d25277de54625d1bdcec81a048f6
z84a8193f0aa9b77840612eead9bae639e187ac2057b9bcd348ed0bf10e7cd94e06fc8e9820fd80
z0c541a273e20b8f3d977a9c82f460bb4b282fd3dc9b984f121e3d7266d19cc97337109b2fd7ae2
za91c6a0c84b41a68af6ec24389418621a2ada8c67e75e70fc2e518ddd348ebaeea840066ce783e
z2292c7c449ccbf8855c970c8fd91df43a9b7efb3ac5e4d0d59becfb3ea02290f958f8eb9144159
zcba79e8333bd0d81cac30147df593893fd73682d592d915f9889364c2f3ff2cfe68b84b538b0e7
zefd7e7d5d438def5d0db49ba675ec8b65e8c314f757bae6bec9d4a7bf138667e4cf27289c396ab
z72652ba1f6372e13186a1b5fb6a0ef021f99c1d85be7b5a86c914d76bf9dc79dc0b0511a49a817
z96df04a11dbdc85cb4732eb9b15527a1ba2710246d2e47dfa248fb2c15cc744335f3f25375d0f2
zf420afc596d8ef317dd8d9850a7713b7367b95cda111fc0e0388ba67b86f70d6152f99fbee76a4
z806012906d469e0eb426a4ea923ec833834f72c27814ceaf85deb7979bb1b70d94a5bbf7aab066
zcf967242b5e0311d3287a609f2fdc182608e54bb7183000684b0bccddad20406d921b087353022
zca729544ff865775073df4f1d822cb55fea363a6c1285fb4d87fb84ce8308786cb1648e265208d
z991ec8d35d80381606a7b509bbe908d962c313edbdbc811d475e6edd0ffbae2164d514869f720c
zb010aa4e0038cb06f565cea7ecb23a7e49c0bacee596ba5d74450d5ed304cd223ba2595d3961bf
z81810baa44aed78f6d509754385cc23edbdb86f2bac69fa66c799eb648f39d410c916ecc72d81e
z85f264541a687abde9bd62fbc73aa4b45659de393fc8a2cf6878eafc05b416e9a4fab015f56398
z8fec43483fbda2f7eba05e47bb838bb50c47ea5563904ab710e74fd1bc56bbb5a4ed2d3d1b43d3
z6ce73c6ef97dfb5c1dda59cddee64ea1a405ee77d7c23feebc7d6f38f565de8a7088557ad675e7
z899188f2e5684eefa13cc3686a0af4af1b92e028960b9bc86818421caa84b905bb8c039790f91b
z2ee96ea83743077b5ba1584ebc861b9dcb70555cb28a8fa90d7b5a0641b42fa3b17f2b928dd720
z462f7fdd2df2054c37a41f0f427b581372c33fb480ffb4e00cb6e06ea085f23dbc9ac31531c55c
z57aed55456cd2d4afed57b42df852bc2629600bf124de05d64763f50bb31c92eb64fb21820c908
zbc9a31c4a4df73da77a97b06601b9f9b94c7b8d7dd05a597efca1aec85750bd26926cd6ad02a55
za720f5ee93ffb482b5af4fce4731b9cfc6de3e1585fd7e66a334f61ac4f55616d1ccdd0fde44c0
z0244c4db18d3ddb4379830bb1a37c79942a8aed02f9a50b2e8d13f371fa1acfbb9ded4e7eef955
z8bc880b5b31eae313562db26c6b47f232ceb175962c4f11100c7788e45b1b70d9c39cbca1f9c5a
ze6cfc3a8b41724c312bcb61145a6aaea1a1efcb1333dfcce137f5f18d314797ce953e28bdfaf9e
z68ac72c7e8480c08892cfae305845f18db6a9ab4f3934a6acee6b54681ca8b01099505feeb219d
zad464fb5bfb6b863f23e41d611c0f7633f722d3aa68936f3f569f443ae8be8d5aa69b1ad26d054
zc151b9646707e46542e7af078270e78dfd0bc01a3c63c26625071cb929e284ea5db9543df60b8b
z6ad6841fe35d7bf736ecc82353351fcf5f455b276a1d88c3e14f24d0a2eb48ccb0689944da4fc4
z2c5d76420114df148154f0f879528a60ec800b3858b31687c970fd3243ea0eaea005335bc8244e
zcf38cbbbab691cbe16ff9ece704d72fbe3b07b9cc69b9a9616ca26da7a83a66fd30a46c00ee977
zd4b3af3bd18253a232429489ab9e396c9fa2fe9af11e19b64b80b0c7bf4f9abe2c8bd8e8fdabe5
zb88a1b26da2968a860f396f8804878b00cef9a9ec651906800aaebff5ae7a33ad5b026dd707477
zaa163096b6f88efdae4bceb5808177249816bae3d4cc7bda19fb8f1bbcb432b6f9f1ee4831e7b6
z676677ec392b5f7187132d5c7497a895a77ac184b776ab35ce066823ac675f0eba35da0aa586f8
zb10efb749ee6323099567e9c058193121a8cb3e21bc740d80961d46d660eed94c01a8db52127e7
z4777c48e48e46ae1d70877f01b94ed467cd263ff3eb6226f795e121619a8beb151ff2340ec9957
z105b504117aeb52cc275b2c5e5fb5e844d8bbfde911c0ca1dc7d600a18c8459946791a008ce0fa
zaf3cad5eb4d81cb6825fcbc7f69aa6807c204656093ac1470fece5f2118e72ec516a4c326e94bd
z52ca59eff338b1988b0f594d23ab67ebb63556bdfba18cf6fcf5f259fb13f644a83b14bb350412
z8bd910f9331d78f149374b2208a69c221c24832d327a0bc139b0bc2cb45c26392840499796e5db
ze40b48bb13e28bd2e14b975e3b2ea97e54248eb090174630fdd70ece14da2ff7e82eec7f28f913
zcbba932aeb1d9bd677e559a4a50c8862f86469f69a1e7c1020ea811dab2064593c338e6b01add1
zaa52f91d0f74e1a860c6e53b1efcae878c104beaa465cc2a0fbca98736cca2cfe5eeab96333ae4
z28b59342e4175bfcc420b457a16e539f1f26848a446eec61ebaad5f1007dbdcffca188d2b9589c
za691dc3d2a223b0916ed9f22f30632609a8e6a53bf3c61edea857231e7f72848a3d96380d52dbe
z2bd634bc123ed500013ab5d4bf23c00ddd360a12ba96351b3ad093d9e1e554977c14ef007c0aa5
z99ab299c79de2b1a590e94f315411e7033286794c2f3a828e42279b1d09466c88f44f30d669566
zeb1999dcd3488af7e2c4b624a2fea8a3e52a28ae9310563687ab38a0637074040b0b6e6a1172de
zffd07a40c824d03368d796f277f7cffe7d93145d5c465305d7602bfe02e0ad780e7ddc361f7d09
zc0397e9daf37728c36b10c747ee86b174a66d759e1d37ea7c1b90fcfff16e88f59baf44b03cfac
z82d236f49745541e157cef94ba69665932b81c9a43b9ea9f1824c0c0261d45f176151699c38675
z66e146874c153d200e02f1952adfa4daafed7ec46bedcf7c682fd816aa3d778a7e7e8deff26461
z2e434cafd803c14f7eeba82f2ac258eff9d0a2bcd49b2398e4f07ed83a389c8c6a1cad0496951c
z7705b510bbe875afb9ee185e3916c1187810383d74190b7d957d2ab2dcbf90b199055b1bcb8e06
z3ca5f5e55668082b654c39b5ba31bef3a0b0417d6240f8250725cbaceb17662a575cca40299669
`end_protected_0in
`else
`ifdef MODEL_TECH
`include "qvl_pci_express_flow_control.mti.svp"
`endif // MODEL_TECH
`endif // encrypted_0in
