//              Copyright 2006-2007 Mentor Graphics Corporation
//                           All Rights Reserved.
//
//              THIS WORK CONTAINS TRADE SECRET AND PROPRIETARY
//            INFORMATION WHICH IS THE PROPERTY OF MENTOR GRAPHICS
//           CORPORATION OR ITS LICENSORS AND IS SUBJECT TO LICENSE
//                                  TERMS.
//
//                   Questa Verification Library (QVL)
//

`ifdef QVL_COVER_ON

`ifdef QVL_SV_COVERGROUP

  reg prevent_x_to_valid_transition_count;

  initial
    begin
      #1;
      // This is required to prevent the coverpoints to increment
      // when 'x' to '0' transition that happens during start of
      // simulation
      prevent_x_to_valid_transition_count = 1'b0;
    end

  always @ (posedge clock)
    begin
      prevent_x_to_valid_transition_count <= 1'b1;
    end

  wire enable_coverpoint; // Wire to hold "when to increment the stats"

  assign #1 enable_coverpoint = (areset != 1'b1 && reset != 1'b1 &&
                                 prevent_x_to_valid_transition_count == 1'b1);

  covergroup xproduct_value_coverage_statistics @ (posedge clock);

    type_option.strobe = 1;
    type_option.comment = "Statistics for Xproduct Value Coverage Checker";

  S0 : coverpoint (!($stable(values_checked, @ (posedge clock))))
         iff (enable_coverpoint)
           {
           bins Values_Checked = {1};
           type_option.comment = "Values Checked";
           }

  S1 : coverpoint new_var1 iff (reset != 1'b1 && active == 1'b1 && enable_coverpoint);
  S2 : coverpoint new_var2 iff (reset != 1'b1 && active == 1'b1 && enable_coverpoint);

  S3 : cross S2, S1 iff (reset != 1'b1 && active == 1'b1 && enable_coverpoint)
           { 
             type_option.comment = "Coverage Matrix Bitmap ";
           }
   
  endgroup : xproduct_value_coverage_statistics

  covergroup xproduct_value_coverage_cornercases @ (posedge clock);

    type_option.strobe = 1;
    type_option.comment = "Cornercases for Xproduct Value Coverage Checker";

  C0 : coverpoint (!($stable(matrix_covered, @ (posedge clock))))
         iff (enable_coverpoint)
           {
           bins Matrix_Covered = {1};
           type_option.comment = "Matrix Covered";
           }
  endgroup : xproduct_value_coverage_cornercases 

  xproduct_value_coverage_cornercases XPRODUCT_VALUE_COVERAGE_CORNERCASES = new();
  xproduct_value_coverage_statistics XPRODUCT_VALUE_COVERAGE_STATISTICS = new();

  initial
    begin
      xproduct_value_coverage_cornercases::type_option.comment = "Cornercases for Xproduct Value Coverage Checker";
      xproduct_value_coverage_statistics::type_option.comment = "Statistics for Xproduct Value Coverage Checker";
    end

`endif // QVL_SV_COVERGROUP

`ifdef QVL_CW_FINAL_COVER
  final
    begin
      $display("------------------- Coverage for Xproduct Value Coverage Checker ------------------");
      $display("Assertion instance is        : %m");
      $display("------------------- Statistics for Xproduct Value Coverage Checker ----------------");
      $display("Values Checked                       : %0d", values_checked);
      $display("Coverage Matrix Bitmap               : %0b", coverage_matrix_bitmap);
      $display("------------------- Cornercases for Xproduct Value Coverage Checker ---------------");
      $display("Matrix Covered          : %0d", matrix_covered);
    end
`endif // QVL_CW_FINAL_COVER

`endif // QVL_COVER_ON

