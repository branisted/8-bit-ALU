`ifdef encrypted_0in
`protected_0in
ze74c34e226135848fe16db9ffd31815111b6d7fb642c521a3f628cf6da949865580b22efd062a7
ze90adae0e65e66a2c36a587d0a790699161455169ed55a01f2084f11770a774ec4c588039b380f
z6de9c5084882a40b79a175f5c2114b2b6d78b070cb806e1c0aa9258297f4687ab308bc470f0040
zb0b1de382961eeeaf2e279e1462520fc31c119af8f2b214846f56c2b3cd2eadbe4099496abff18
z15cec83ec4a77b868344aa20ba7360908f5c0de2a79abf8b3534b883bb12180f68b5d4beb444cf
z3fba8f13afb0abfe8fcc4294810f75afe452434d2d0f1166236c82f76edf1e12979f04bc35693e
z32ae028996dd85737a8f5adc1ebb94f39c940246e887647b64782cd7ab429b0544c173176cede7
z01dfb26b1f73408344a52b7e1f117f12bb9c8077b34876c2e6fdc085981637012dc9754765e1a9
zc512ce062e0b8fb16a214591f5c81e1353b900a611fe1f4886b57940b41b7f2ce99a7b84b04b90
z916f717e73bd10589c81e207ed77ec660a8cbed5b487fa50acde1b055c8870bd8676023f21ddcf
z9c98cc47cfa2d654ff1365d1f45035a045a66c5dfa82790502623b57a3af03bf0f0c0d35b51558
zb8b5f2d29acf03737a9ca2a053b7a8f06800d50b465c41b30eb585f62f3d0c2c5a43bccb0b7b82
z3a93cd6c1eaa0518201fadcd476c87f4109a0e3f6323004b1a64aeb50487c8991c0196054bd5e2
z46775c3db54805f307230c741b8da0c9fcaa49c35527b2db20219b9f224d3dce8fa90ab3e73f58
z98ff271bf07ee72fdd586a74277b6b004b9b15d85615f0bffde84e0c96aee53520e9185420dad4
zba952774946894f65800b677f485ed62936b3bc4af3b1d02c24251762dd419f73e88e740493883
z4c3175dc36268d95610b84c258fbb58fe5fac93131cde5db76ecb697868aa40b498b0dcdaf6064
z7601e6e917fe1116a6e443bbad04096b4e5d65b8c9ec849d7ab30ae640de42cd2d5f8c1de11cc1
z31d342e556a3f99f4553c34eea62ed0d3d62c6e221ab002d9189773172ffc7963500e62109eb76
zc0d0dc4826f3c4acc9c777e80c39d106101ffba63387de6c20b57289b959f2972f126047825856
zc9b2b7ef6ebe0f51cd9174dfa55842bff37d1713420239bf384b7d2d500c18d7867ff1630cfbb6
z9b4a6af3b476ea533aaa52031fe969b52d13482819f32fa1a4c644f052e9d156ded743e6bfd547
z8bc6e7ae600b0699558b54806e21322e10468188a0e02d414bbd7f4e20de597e6400fd310a6583
za702f31af931e29ca90b522bbd1630920671922bda3d09c9a76d91b75b407fbc4ceeab586bc86e
zbe2ce512c3061af2f7f46b6057f240eda8c3789d58681a6de8f30769f497be54ba39490acea930
zef4fc2e6509c5e938d87294889976c220c6f6b7e6276c2622c88df825d68cc797beff1f46f0043
ze0841fd6eca18851116eb987b1b78e705151ffad395e9e471626ef01a021d65bf581686bf2f27d
z1765227f6c917bada86ab374ca14574328c98d9f8a2b26b4c5c3d12d7600119d5f0727b0d2f183
z041c03d84ffa2f65beeba257c687a24f8b49c7e35214505a52c10d23584d725859de738a6bedfe
z43f9463be7f21f97d3b3d1744c1307cc07a15aab76702ffcda0358927fd5125ecc8a7799a02987
zcdb3b3fb2103a0a54b351c115db8f4671904dfccdd66b42a4cb54fffa595640717388ecb8ed33e
z3eda4157eb888561f216571061b5e7ed2d2237a95de31c10cebb2e503f039c4e5f9e53291594eb
z9ce98545dd1e1ad52f68154d0182ef2b44fbf238cdfa70c4ccf22ac6bf6c7b43246f624bb12b04
zb505fb7c54acdc2a3259e5deb21582ce605f0dd62db398473085f66b730d217826b43397738f74
zd44639cb1c94449f6122847733e3fea2fb17dd37c5991a54fed893259f1ae8eda7e445d968b2e3
zfbfd2faaeb3ee03424ccd10ebef9f787fe96c0701d86b0c806af5e56cc6a840198aaa7c7660ca6
z28b52067e7f22e9dfb48a550799ad0d06c949a3a05926ad49a8f57891263e29929bb13313c6371
zbab4bbc913c18223dbd42e222e4adc150b7fed8e64aa7dbb3026b353e7d609bdf03d3466483404
z0b29347d31bebb0997c8530c8bd8868679c3943ac53039243805359ba6c55c4aa54f1716a5243e
zc09ecdde0756c36d447a7e06870c6db88fe70fb5337be6de049984696c2ae2cc403001e77fe217
z33ff146531ba1f81d81ad35e14cf01175fc46a1e034a7a5091939eaecb7e3d5ccfe3c88d12b128
za6c3dcbcd6782dec3aa0617e5ee2b4f40930635a888e6be4466231e7c7f65d4ec52504a72887dd
za77463a882d07daa0f5ead56e90d0ed9d02a3a8f440fe0854d30e38c06ced5d59468c1ef7d9c9f
z4018b3b8d1bfc731ae01065e6aaf49f4951eae8b4193e13e449e516f3653dfd30ed1066e41492e
z140a06e50a1e68308baabb51f25bf810d1098f51e0f67ac11039e0ad7cf48f8c5301b2b6ffd014
z9b41c421326d3ddeac6fe723c8b604655a62ca00b84cf3ce2454f99f4dc9d4f74dbdc5e1f5efde
zbb0c6d14865f62d77b69b991940b37e7607d02fcf8d46f3edc8a93b9471100b57fdee5849aa5e9
zf62b7322624119a8da6571b677c2e2723732571d1091f06c27780f6a9c900b39193582fe441a75
z696222b16435568ab493a2c6351985e3bafceb44449cf41ea6a7b8be222e52bfc84ac717537c87
zccc4492924c2eacf5831076ad28ac3c17ef7ffce1cfc9beb90e72bc7c84416a8f5b6f4e7b56f66
z466c3536fb2b64e36e647297661d414fa402f4820597154e7203a8da71a459de384747c8e0c915
ze9a3fbdf8d9f3fd66c6c25f92c7e6e0db1d1b775f49afedff6b741773862b9bc6e89306a17f56b
zc812bb61a0c1ec8de96906ec0d4f7ad1a173b816957a57191a441b81768d2b25e9d0bb408f10d9
z45137d292494172871ffcd65e1f0e5f3d63226a3f7bd2ecfa3d2e43b39566db3dd58eaaffbb0fb
zce848c10e08452c5d35cc47a8adf67b1f3fa2e5e0298d1c9a222baa0b45357f5552b986af8178e
zb1d9987cd2ab2efe987131784ab222be65b1c9f96887cfde0bd49df5241d657c6f30d4fd82938d
zd8fcee934a105a992c8e39597114cb9fd63914a4022496eec8d984f538c401b92edd979af4fbd3
zb0a9f1c57fb63ab22d0a9b00a0479fe0cae23738678086e7b0c3ad7a3b895e0a51a8e4128c4364
z0f53e708310a55a64a798b1bbbc6c37bf2c67ef56c0c3749c52116d900b92b96c7304af6c4f195
z585f07f9435a7525ba3ac742e01e80028685913a31c4733a30d7f0d89d20488134fd7e8f95b47f
z0e6ea4888f7de7773b3f8abf785103658dcae19f632cf2348f2bb5e9e5ab70bce5fbbd9c31938f
z66c9f9dd0015592ff2509d49db0fd094777b38477b270233a3824cfdbcf31942737c473d5c48b5
ze74170bbf4edbe8bb50736bea559b31bc5b689cba202a701c8001e818c51e5cfe6e7faedab65f5
za952591ed173463c65ae18e75589831c2a1c72299cb2994a05ceed5cfcd7b464876108ae6e2b0b
zcceaac8ffb578c60f987303b46f164c40a498359d07e347f682377d58df99e3019e57fea8b36bc
z8d92d71b4a0b15f4a19fc242b8d05eb16393560c540140ab5970f289c2c28d90a7f6718b697f0c
z794d987a10f9bbcdac0caecd1102f68d043229e68bdb278a0401a17ac22260df147cd25dd35993
za4ecae08ce5e299d23d345d18ecac24404b11370717f6807eeb79cfdbf5d3abc6b6eb387a0cbfa
z751bc3bd134a3787bbb90a8b1b8fc3c9849bd5acff64aa163b799d9ab45d0ac4d35273a119dc93
za7bd6cc9834217ddade95c9ddbd33ac363ef370801112d059f932b64462add577df69ded8295b2
z77b434fa268cc1eb13b0b233613e1552a712d1c478b89ddfb4a71cb4081bea3f4fd3edf0a255e1
zc688e22e6f674809bea15dbd1b6b5eeb5240c1e734e2ebbf28604d0a93c1f5ae25f9e3439e674f
z577826ad60ac7c59a18dd6b25ff43bea5530d9184194e5656f6fa70b0259c8eb9ad78144716388
zc0891f0cea930ead6009b52b9d4549c62711dc10ab12e4e41adcfcc907ea07eefc7aef7c6f67c5
zfa8923826648c02e43c62b46964c5856acdc9dc455aaa65532b33ed62f2fa22bbf9ce3ce6c94b7
z8befc8871f723ddcd9287d507aea25085fd6238c95138453569eb566a980ffa7275bf1506f77d4
z7752e2cd232db07ecabb46a85605532fd5299f1c5e0d031072700d96f1db4b5fb0de3bc6330cbb
z6b60c1368de35e4ad592e8798437be23853da7c430fc2f43120b0f2c4ecb1ed3353ba86f61b269
z8c92ee15568adbc1a7be688448eafa2226ed68a42dc4f66a0d087ab93459ff2a83bddfc84a6f75
zf4e78a1a382f57db33bf31f3bc96fac57e590c27f9ddaa8442df2b16a7a43e9aa41d74ca2fa54a
z4f344d15e810d99b95c41fdcc3a3fc3a5d5194e1ca9889f80676b289073b4ac9a4bfca1a4436bd
z3cddf119de9b2831a88e414eb18898db3aa585736c2fa33c7328cb2325b36d3531e859073ff5e1
zbc510e84fcf302a22baea03a0c9d76e3a0fe2f4a0a13556089af06e75806eccf4059219363f1af
zbc28db2a92e77151f7384f8aa8fffa26e6bc7b5943875c9939bb2f2295d5b939e57cc071c1f456
zbc5aea947c9bbc2ae54f9e4b27595e9042289bc188269e58da5c4c4b3e67adb8b0cc7934a127b9
zc045017ea0f74d67d5db41aee2a7dacdfa8f2926d98bc8206b8780b93db35ca8a8c1643158a378
z1250dafc517f04d57363984fe48b05e2a9acc433016f8589747e1ae749d0408b89de2489d8f78c
z8330de79daeef2d18063d30ecc42ed2c0e6bda90398da7ed4993d2f2bd78af57705407abd4e1c0
z73f6fce6a4f189032fd39a63781e52ad2e9760e5f5e17bb500c6baf42cbe5929bfdfa9649c4bf7
zdeab40fb14cc896cf9903f9e82d9e569e5de24681aa6ae5c014a08ea91247c9d529c816fb3bac2
zd8fa216eca8af60fb46ca31c9c21fe1be11942ce7a179b97388185439c55e8f16d948c4b310adf
z94898c412d1bb6f845d05f70079fde603b6a648ce55aa80fb8ba02311fae1e8d28b1220c9bb9d6
z384ae70f0a7ae73a2838e7b4bc8977d80dfafe9cd81ff2973d272e11b2349b40618b22661cd5d9
zc759a56809da3f5a219e7f4d674053a076c34d8e66b76b820cf017ef14a0829b5ec8025c9e0292
z574a3bfcf9b7932207fe7bbb70751d55e7dd4231a2e90c4e940b679d2cfb4ad285b865be29a06d
zbf3279b4d7d5cccd668ec633e90ee35d2e11e8cb30805dcee0f5bf6a07c3e4e4b2e2480ec798e5
z5c2bbbaba1f86302368c225d127d78cf4c86a0a24eba35d587bd9eb28ea3e71e6278bb4ebec4bd
z4e8916e353e78786dfe80c06986c2b5db804a5f0df7e92b73b9da728e3f38fd463fabbcf03ffee
z88a6e98450cf3ee1b0841ebe5387e27e06e9c1fe0c26b76157147459fd8fa43c9dcc6b25428524
z72122405490d93cf0b27e6d4b488a6f3f6ff655fe9f111946c5f5938286f26899bb252b3791df7
zf4eb0d5a9fc91dfebd67fc727d5f17f9563fcf99921317a0e492ba3925ba3540d0f418f3181733
z92310455af6fd65e3f98a8d49f76784622baaa268cfe9597f00ad6b9ecbff991925b749e077c76
zd962eee833db15c87d4678ed8f7db75c064be29f73bbd9c135123925b16638dbc43b3f0ddf289a
z42fac985dd543544eadfd07d10250fba6808d3aa1f4475655b3ae85a97c13000e73c44c248d5e8
ze70f52adb7505ce0099c05de4edb7a5122a8f5c41902415fbfc7c9c0edaa1d61d599d1f3702a8b
z58b137ac7223b8403bb70f61a7e65695d290c2713177bd9e423b802ac24844ae87071156ea80b8
z7d560803dd055ee0c847454d31cef81d35844934215dd467411b302bab6a2565ba65829a4090e1
z4afa1429286805e2137783bb81a94fe689f26675482aeabc2ca8b82218e65762dcc6ce96e5c759
zac371ff94f9b3eed5c873682ee7853fd427d8a778088286d4f97d34ca13cba198716e03103022c
zb1b2e9c13bb7ed87e2f5ca474726ecd7bf9778c2cb697cbcae5793f4d175e402dca92ccb1ac9c4
zf1635e791b574b9c07c030371fd693db6e17980d6f5afb12085da5ca97596248b2cd9544cb2770
z92790fb09993180e8adbc589a030ba952c2db5c7c11dceb048105c9091ecbacd3c54e04c7fccda
z3dd5a5df765feb2c339b626b7d6a77398767636542d778b6e88019f02122893af451f3de4efaff
zc459e750a776d275118f0203ad30dfda50bcd1e103337e1b17a7a83636dc6cf04903c90241b5d9
z4986d309c200547a90160227fe1dfbea1fd723aa59d37ea494c21c87ed8b137c8129a285ccef35
zac80a8279f0854b71efe38435d4985be5a249719d4d14f49b591652ea3cce9047628ef959a9125
z176b14e5624691d4042f8d3af5cc18d69d956c26501846194cdb1d195bba1ab3105b4e372dbbea
z534d2cc172b26fd38f5d728fec169eb31d5eeeb6294c5aa3f4e548eb2142efd281a9f0260f37bc
z23e8482ce2210880a49ce24c32a6298bc8bd2e01701d8727086496502a71ab682a480c2d3401ea
z68377753ff9a3a6812e051772bbd6e0edf6d4fa178d3e3bf5608fa3487f8abf2fe2c304df21841
zb9bcda643cb864494956c742a8cd529f15f9b40c9ed14c770771c6c307fcf8dc2a1712c159263c
z6690f1c361280b545431b02e8faf44d93e387e8750431a689cdf36f4efedc9e161d5e10ea75ca8
zc0b4742345d80907613b63d3b5f1b404191f9222ac1ddca593d755e2c57c031c916296bdcb25ea
z34897b17883c4713ae2dd19d7a05f8577e4747c088f530409737c1f838f9f3a92afdbfb3508316
z51702ae87e8951579e097f7888a04457dfaab0310360aa0f2fbd403fbce210229bdd249edd8797
z87824b99c13b87756ed8519911bc7cffa46cbaa20b2848b32bfd9df8fa5cf3043be5638325821c
zb6923672c7273532ecc50a755a07fa04a08e02db12e091e8305fcad348896fa131a655fcfdad17
z8c85dd43f552aa6fc71f640d07c85ef9df05628440986b6737dc9b3775ddc905852bdde49770e9
zb780d248b20209fcab56cb38de9da6c102c4b3adaf7e454a09cb6b52af8f2476a8b77437df53b8
za49e7b2df3a2079cac29eecbf14f2b73b7ebab54db6d1af33d6b7151d07f063ba4307450e78efa
zcab952473d3b4fb177a5e42703cbf1d96f4f4bccd5a6bd91bb27e9905335ec731d2bf2f8c11285
z06b66d9104f4bc6de087aa5bb82da67e90a9be6503c6c47b10697e96c3131e3a164482edb45249
z8c1fdfd97c94133597654b5a5a27bdf4907631da03a97feb012cb8addec438ad76865c1dfa155a
zfd6bf22873b6ccd20249abcfbcccf85310e25c8e3888e9ab2d7b44971005dc9df04d4f0677296f
z661244a774e6fde9637eccbf01e608055385d014857eb2b0a8fe2b4786efbe22224b875d93df8f
z26a61db0ec7e8928e94fef8f96ce1387bbb13d51952636fdac0a360a5b539757aa41fb20fd304a
z6e4e55609a10ca65d18ba2edb26b3b9ecd6e2ff195e0613db38f57041569028361c93c1fd02791
zfc39e0aba6ddf6efe2d81a85fe2009bf50d6d69d51d1be1298e0c0cbf938d9bccb6f6a726be74d
zd18a3b2d76615467d9f065642ad145deec5787f86bebac21dc06cb5f56102d69f09fdd1ba7b352
zdbbb296bec01da36549bf500dd30355bf9563ef25ddcaccb418845cbaef065a055b73e1a0b35a7
za047369bff6f01b04547a82179ec080820b1857c471671deef3961d411d743c025a2e479801b5d
z96c163c899e24186f95f16ccd4f3ebed4bff6ea601e9968ef6ffc5a12e50ecc5e01b39d9d48c29
z2f2718ae2f6dc8b67edcafaa9a9ea3c90c0126ad40d1cbef9186e8ecc862e54bb6e22cbd59de1a
zef740274597e2b860b0a54542a59e74fe47c5d344a1914125ea9ddba46ee9e1313b10c2c75776e
z7831d9ee86eddcc0e0e68ca98b9c3d189935cb20f4012f29a4577474d32ef58cd9a90e340496d5
zfd2992bdc809e6167d3078cd21d37b30e80197034f62dd99dea272924e3a4fa2f33ce1a0b37517
z4bb9e31b8c6c777bcfe07e74fe844106d217cb2cbf023856b1e097dccc505b6061e9337bfd09e0
za77bfd68e8916bf998e6d8bb9557ef115e93cb163f4e2eb6d5b95f764a85bf84073b0cd58b39d9
z9a8195094c932cf897551efce28d9fc43b96ca2dbb372ae10c0a405f5ce8271ec7d64f62eb9388
z4122af990e0bdf2eb9960c283a7c95808fdfb4ba804513aeaa624f6fa536bbb9af44573bc9de97
ze72de73356fcd8092160bbe2db3855db054a5e62af9dc47ddb04b86957c244cc07e377011dc6da
z8613c2213384bf93ffce180d1fc82437184a989807a36cc14836f79b95531a95bd20e6cfe600cf
z839bd9f6ed645d73d96f9346aece227a24b8d4ea46c31be92592c23a9f2d6e3d9cf035b8f4905c
z90f564dc2c95069d511aed733411c72c9b9adb06088ecbeb7f8735cc12e778b97778014cc7f061
z369fd2c51ef2f055091d11a366c2879ab692c4b2c640f95d553081e95e0b9e3d95275dc67e6fd9
z380459e680702f172f698879c2ffd32786ee5badafbd95a03f4850cd99b41002d1dcfbf1fe1a7b
z2fabc4a002a55192dce44afcdb3e4cca727c48b0a2eaf394c4e93d03c03b0d09bd7c60d0e6e77c
z6cd22b8e43d4ca693851d527b911f90439edbcad44725460699ad3d235521c53b7f8693c366945
z1186ccf02b27cb1e035feed5705fb41ddd1cdcbe496874ab00029ba598d673bdc8af8fe2882401
z871c64f81ad818386bd2bb375e70a8ba45d96b83139d59c6565916ad2004dc0a5ad692fcd5fec2
zbfb5280f7311671dc3eb5f9eb8b387b6e1424f829ebac1b075a7932857f9d2a3761b5c786209b6
z7219f3ade48795bd81c7a26ffd16a4fab6ed66eef13aaf82e31122a620813b68b2c8630b251d15
zcd2c2a0ab002a2f97cf2562beb1b00b478f4d33c40d34c0016e48813a27af9ee30453c1567e6f3
z1a43805556f972d48d06cc180e3c1d826f0e4ed00cf6591392270307741ae8affb5216b55faf94
zfc6f345ea588e0f7788cafb69426da73d912106b2d942c29db402e94f2481fa0cfaeb64ad490fc
zcd55b0ec26c544c208cb8201a5f35ec1848ee030a938ce8b11a946473ca7313d6270157234673f
z69d17a237d1ed6dc57ceb39b03eac26269b8ba1f453adb33fabcc5cb8ca1e1f29ca4960af8014f
z980fe431b80a5e8456c09ab223d5db789743126aaaabd35cbdb9c878b09e00f2853223b1ad6ca9
z707a41e6ed8f0eac6d06ef229cab2b07c5d263c4e3297f16d06d513a9930ef8f041e8e5c069dc8
z9372da23045c6f2098e87a65766fe76429c25e9b49ee401ef26ab65905afc17f532018fbb1ffcd
z16c6ffa9e66c706c3fe1add7071a1e315108aed82e5757d4bd2ab997f95cbbbbf80b2b57279c06
zd1aab44b6bfca674a513763882b616e3dab8cef800afd93e4c49777461b23865cec32685bda507
zd394c67444793e4580fab9d851f27ec1e58c31209a5d754ae98105a5d492aa83438c03895dc8a5
zfccabc4debf29b56b318ff95e99b81f17678d99b070f8e0b035fd3133fbfa6f475ec56b814b165
zbcc74078d0da3610dad60e5be6cefe345622e2e37365cc686146293bb90f10424f0158b613da50
zb06cc44b933f11015da1f49573bf13ae120d182908c1a4037fdbfc8fc169053138c238f5dbc93e
z0f10881d4da8943d2bda20295327a9286c3f73bb6396591b142d78a485c2cce0e5183748a301e5
za5dba2a5a504c2605a0a33148d86ebc1206fdc490f4598316e633b9da426a307f04f1619eef23f
z96821c5c6fa25a898b2e0b9a87795b97719ac7a1db0cd1a8ce099deca1d97bdae8b8182a8ec6c6
zeb9a903510be4d50fcbe25157b664f8e37088a536f7ab16891c2f2241c1b01eaa2c1433572411b
zf9a5b247921d5d3e1b7cdd6c548e77a355043bac3eb4cb90363b477cdbc97fd2812c57758d5536
z185ce82f9e3039c7837d089a7fabdf1a74650fb0af4ad8687cf5aeaa3e8377abd05d0777a61d85
zb5414105ba756ac5bf6e3cef2d0b52353af41609d186cccf9cafda2fcac0d8bf5d50d748c9bfc0
z17d660ee1fc865019013f67c06bdbdd1e0e442a60a986a82b977cfaabe8c5b3b54798055be3614
z4a7905fa00f025b843efe75c4a75735a278e3592c317772efe4010cd201f3785b680842d25737c
zed76949b5059e255687bd2d2dc73442d3270ce2c3b9a9a0d0f3a5e7601e7cd06c03ba71911a1dc
z5d6985fba897f574010e3bf689986df93bcc6c0c0cb9af62dd23bfe783c640d48de21736a4ec0a
zdc5b993fcff0648b8f48d4d2b725754ab2871e2835e97aa5fbf736299fee6e61c230058c83a40e
z0b6d8acfe09d189a3aafdb023158e745caa5a2fe86c132f23d80150c12c95c4362c57448f3c124
z95a2eab0eab7766cab03143c4986c0a21393d3da65ef6124deca58480bd82d429a8a2e86b18a85
z0c829cf84d8d3829c771313a7833d5a30fc8167f1c73ee931eeb1b44a6a1c2db23a95fcb1f54a4
z9b13453e7768bc400402bfe823eacac99d179eb9e927789c8877ce552daf87fcba14fed8744216
zd067d7d0c9861d811fe65efc7c19ff0bd2dc33378204240a388508933f50c6fbe0bc20ad230cb7
z2eab417a2ccff1457a6cd7aa53b5d6e0bfd6a7d3119ef3e02e8becad003b87b26b3cfac669cad1
z791c4cc53fae6b4f0c77082afb84c8f3aa528963b3784ac0d48bc9cfe53894346ffb1ec596f5a4
z509ac124a4b8b357da403384f0d0b260f7b4581d64b526a319106de7dd1091e6cf24a135ecc35c
z5c24e36f17e136fd1d6e135de334577031593f2a56ee6501560cd6459fbb773365f6c48c52760f
z2a771d6634ed216a2ca645f73fdd05800c9ab6d78586052832fd94b8a6ee17c0bc680abccdf22c
z97a90cc45f79e7eb439e7dab376d97fdb3a1ac8299652f6c6c2033393c79f94fd29aaa9fe45775
zb10f8039acf80c1b02055bd5a2cc6c39dc7aaa8a1f97d1b24f928c8ce298c562310b97abaaca8d
z0873afd0548c010c663bf3676eaa95d530788d8f751d7b98b65bcd98b76bbf9d9159bfc96dd237
z9f0463afe1d3ee2d43d78135247e01a797afa7ba1507351fe390c463d4e1c497d969c92d1c49a3
z00b95163345bd4c443be5d86c2d82d55b1939ba7801f0a0393a1019d048e9f68dcb76afb7e1de4
zf456812c4103d1c3766a211bc53b941448d269aa2bc5a427e544f10d5982787fd5e40cf48cea5a
zb0ac183291f7a7e543b763dfbe8d624c5f3705c1935f50fdb966cdf366e6258e640b57a796ea08
z8121135cc554d7602206f0d69c5dc4d6c840ffe243a23168af4d899818b63c5a9ceda8e8f2f296
zd947556001b9049da831bfabb1e9f318bddfc77cfc3e11711902bda1d1d8273887246e6dfad6d2
z5a69e3fd0aaa01b1f7d64c98c0785d367db49e41c8176fd40927cdddbeaaa78953f9f9975e3221
zbd20681f534b6c2152f27993be3185ac8beb9027e652e91092277830895271b4dce09d1c1e366f
z865f96af5397a6e15a121dbeb818684589019da0c13fb0ff73d49c5a1a65fffad253469cf2a2ea
zd4e76f500774fba3c6ec68296b5589dd7e43110da1b8c3146d1030d40d20ca0e57efaa0da62e88
z8a8e2b3d4b11876e7fa4ad6c8b1457e294da14dc2f4b9b43a2d8b0d75dfa18149e741e48d8f52c
ze7a9f36145ffa003dd07a5caaa73014ba2194d4d5e0f7954a2e43ed50721746562b52d52bc8637
zf9b8bfc3a07119949a5112ce590ace43762a5d1f27ea273d3ac655baa4adcd6148521b2fc4d56d
z896dd6fa8938be537e85c80ee5ee47a5c20838ebc60c5cd67dad101330633883273befeb99ea19
z2abe85abc5e1cff4477fde403b5e2cacb02dd326b105ce1c6a16974048595590b5fe0f26614fb7
zd3d79c4bd8fc00a10471668a735da431f2acff84773ceed7d5fd9639aebecb648514a15abc2acd
zfed03a6ee4365db98bf0864d903411c83e5295e398f4d9a788c4edea89ebcacbdf20c58cf1d250
zf4b5d399bf09a145e085d3462983ae7ebd999011cb9d4bb2f774ea9fdf18b07e8fc78ed45ff2a6
zb3b2ddf38d69b84bdb8a9790ec10494300120834450242573459b98ce5af4a0d482f42e75d977e
z2824ee303cbbdcd881cc8754b49c0dc5fe3e4bf91489599123ff1434651e4572c8caeb419119a2
zfc97e380ff8922f5bd5f489c3adf45884b2c67e517fb431e4950c52e7cc324a955ad5591b14149
zb3b09fc5eb2a4ca3c97272a8b2cdcf6c1f7463496a3416895e80e799d8fde1230e50196990cf47
zcfde84adcb1db768477eacd3aab10d9ae625d7f998e2e8d6fa84306320ebd2c1a7b672d510278b
z814e34ea1fa47f74645457703647b3cb304d1f58753c0e17f53dc7c1ff1f9844b1e8268280b1bb
zafad1b38ae84b3c85e6abe4890a745e6f650031812c3580c5f738262377b2eca498411c6484423
z1fa8d328ea5f206875ac0da6fc42303205b7a1950942cd2e156e9db6b5fbf057b7877f21b343bb
z091cc133bd7d48bf04f6dbd57d1b7f16601ec7a596dc51480bcabe5b8382dec09d7f19a3bae8ab
z3d73c14206d3d26353ca512eb97a03c0f2c8a9a1ffc4b07ed137fe8dc4dcd6d3220094aa49eb2f
ze7491ddb732be1b67f153badce9d9d5b61bdb062c33a873cb96436179f2f041c2e6d7c56ee39c7
zb5b7edafbd28cff513a67e9af845ad070fbeca0c384e4ba5e2e87f3900d97068f726186bbb3900
z06b531b2fe529952d25902c82a5caf6e6b207e539385bc815a92a2a485243071bb7935c841a31e
z3e0269fa58feca9034db88149b71e7b8873f2884cd5802c91a33f2d93aa01e60870b528a26855d
z40940004a11adec7f4e4114832ec014ff2a6ab19df252845d975005c154a3dedca9ff255949640
z59ab38fc8678a6c4e08d03429502cb824368f93df3a73980c06ca0d98d534b9b2d3716c54e0877
za6615387d9b0a61eb3b57b79166cc2b3a9a99e754075676127afdd60f2628db33b081e230b4b73
zda31233d131b86739c70d9e3bed2b9036576df2227424b2eddcbf7140f9fdd9f2c8f0805ef138e
z38a9a782fdba370b74614ec7c27009214ba07cb2e03cc9b47ea0ca373fd486424308626bb5db40
z353f2937520e97c4ce00f4a07f1d665b12d71634ac7fc91e6d4290fadba63b8b2f00d3756a49bd
zb4e8a282c4a6dcb66207966e51426da5a55203ffc30fde29a4e1ce4c90111ccc974e5cbab2d3d3
z6a01a7ec5f1daa4c8d76f1f80388c1a03010151d3a53f4b219e01118ee76112626051e1c4840a9
z2d4f2f89df4876feb7fb77e9b9bafb45beaa8748445a209cbf3ff5f7f6704a1e9c73eb60e4563f
z74e04eeb9c7aaca8793e4cc4911ddcdd432ecc3c98289feb6b7997cc398a2155ea373939e68ef1
z81b4417ca6d175351c7c92a74f79b10e3878901fb3b8685cb3d67b491f8221970400519817b6bc
z2c0b4e144072b0b4b0c47092fe8fb32519a54207f0de903d49be092a08679df0443ee1de9d389b
ze2e83c9b8c4ccf8de636097e576e5f080bac4d54c0419e595878129481e1c9e60ef226b8112898
z8f979f92b33b5df879969c487d695da45d0a514db6a0bd79d45770826820315eaf8fc82bbfab7f
z6624afb93c22256e96dadba609e9a80937b668af972424583d81c118ee7b40cd39e59beea7f2ba
z5d770627c38d9329c7b5560ddd48d3a51931e29d56b049d80b4efcf88e0dd2750617fa1b9566a8
zb8f62a24c9b629947789aaf3298d41c4e31bc56510fd7cb778d50f989d78d7a078d92331c08b61
zb2ad9454a4c345d84e9d76c235808537436a8affbeeefbc9bf49252c3fa79eba28afe8443e9270
z398f073c792435b4ca26be37fe6512ef231ed29b6cb6d306111a42f4534786388646c6230b6033
z21b1fd7d5839ac78c1360ebf75fcb187ada31c62a0c6b0c7f44a4c1b49dcf0c40287a3c5178933
z185b9a21b772985d8b5ee00feaad18c73e80a18ad3df8005a680829483f4315585dab3f4394385
zb83b13fa3d3adc91703d15d267406e8e5290e244c6bc0ea35d95a2d86e165d97ca7c3b5a5a5055
zee7a872fb816beacf34bbf9f57c42791e1e32bfdf2826ab5f0ec7c2d225c16aeaf4582d7b87a76
ze3bd976aef2d2ce8cf1cfa43c73806d4ef37c8e42c80316b06ab82f2d3d2c30c506e269731ad57
za8a4cf495a53fe4c3b895bc8b268f3ac92f4846fbada4a1bde79c2f75b986da224ecdb6de68d93
z9213e1181762ec8de214e655d85d1e0a23f6b9cd1b5ec214cd204de1fa663e97762e8e732596bb
zb8ca8f019832f3f53a6e609b669bd5dd7de928db0b0903bb993dbd62fd25b6326c2c31061a04f2
z5ff329455e163bd3440f3641b0db94c3ae6eb70b63a7f52f2454ca3d45cc84aa8d4c3cb5b6da49
z194f218e3389c0a0e68443ce5a5946a4ac7eda3df44f55ff03d24dcb2466f38f49826b38b4c196
z31821e82e8cd3bdf58373b92dc901006fcc10f627fb7d2f539672f675cb580d5333062d023895d
z8fa5b6e2daac100674e72b866a4f14beab50bcd798160c08bcd53a6259e3cd6a35cad5c4c037c9
z304373c921c5956d4ecca9faa7cdfcb45d3143dc782576e827d027bc59e2a5d10c664b82e41336
zdb325b702ea9ca1616c52cb3a04b5c4074218174597ce6472c9318b3dab6d6c71db72440861e02
z8ea68bf54ab6493544f25890f6169651bdb75dc274a65f9b8e5ab5399ed760df906390ec2a8bb2
z5021c6cd108aaa8ef0bc1d8497660b9c9ff86a3499c269c42a7cb8a31db323fed738b8d692bebb
z9e3c44bbe3e903fc95e79ea2822f7c4d8d4ce9f2967c6baada9c91499f215e7cf1ad5b5bd91edb
z3376a02a30fed1b395d7a87b95f884e462c62fcdc6c40ada98f1f196b4bdb7db461cfe0943878b
z4c0b095c09095625157d469a05d7800d5cd65f54b1507eb172f906d1fedda35c7577f43f5f20ab
z66881519caeb84f9a6ac192e6923a6ce6058a2592d0364fcf5fc3428eb548145d2aa81a08e8754
z32494cbcfa301ee370a9edc6251dde045324ad490e1dc48cdc31a974be1deeb22f9cb5f06eebcf
z196ac266a7a15ec7a2a1dd105080b638af6405dcd6ccbb25dd6ffaf3757e77726d8ed0c320dadf
zd31b2df404ca7eebb4334a52baa81610d2bfb739cf8eb2202cce41cb6a969ad114440d3092f6b9
ze6372e5ba410bde2781aed188c7c1ad2c483fbcf8487616e03adaa230bd4cc79409ef2a1984237
z37742e78d66d1dc29f8bc7c61fb8204f927a607dbd250da4eada2e7e01feacccdf54b37c30a26b
zbc5f8d9142da1ecf5bd630ca28bfa66f83fbb9745703484835e433e158d4272c3ef3a9718c0ded
z62e11086001333b05f6293b1392225826544975128db8094d1f9b220829868357c1f23d6c94d58
zd28d4d8db1f7615e49fe371c3029dc7de033147bfc5ec2415d21e1611762890726fda85d94a3fd
z6cd5fd11761a2d2821ea1f4ae8f5c82a331412995df275839c9a562855c07c01a251387e20c18a
z842bfb6d76c6a73cbd7089c8f066afa6b1e1bcf444114ef461365bb9232861c5258be0290aabe1
zfefd456f5b71de5052c15ac9b4edf6c28ecdb4a55b1e9867b13a7c8cf65743d5372da701931228
zb0c00391e3a95d79f84b77a6841ce3b05b1d9ad36479842791eba1cc22db80b9846e3d8e1c4c25
z852dad8e744e924e81a53616d48eb24559caea99420434ade7727feba103d3d70fb42ecf5f570c
zeb011ce7ea09312ecdda56dbeb8cbf028589b7065c3c9e294d3fc578492ac8c4d612b37dce81dd
z11a928881088081ba7424d31d03ae299ff00f87b63366dc7d7e5c40906013c79476ab995d9f94a
z1e2830eca60ed5afda75bcfc8df5a7c4e2b9119270950c3cc8f0dfd197ece1ca32d27e2e0cab49
z39e40d19e9e0c78f789be9f8fd11db6445257a3652d7e10631c548cc78e26ff43a21e55d356a65
z967849af5edcc33bae816d2396e770e333f1edeb4f67d7d58bc542926032e58cb3a85ef1c3ba8b
zb99475d576ea8ff79c4af0747fc5a03c4d242c130a04bd1a57b12502506bb2c9f572aa541c3a5e
z0e442a0e8b8a88acce58b97d48565daceec2de7a669d5bb8659076cfc4e4aebc2ea8c2fb95eded
zbd7883b03f7c9f7fe2ef479aff701dfd967bbbdc5057ba49b233aed9a3f00eb4903320d254dc1b
zc0359e9b2de9b88803fd4dcaa049fa687df7d78026dcb950366795265c1885054a768e2d56b15f
z725524160ed9ffbb1115fb5d29e0390ebd2372344c88f56ea74484c03a63e4b1b01fa211742228
z9aff3de388d343735b69c6ce09ae79143a32d3f6047336733e5cda5dfbc25592869805ed0bf086
z111dcc69616113ce9d9226a60bd961021ed8ba4cd4c8f8a62a8eddf49a2a5431700665c2a3aa4c
z016eaa4c2d918c2a118817853318103aae023c34d9ec1ba90f6f12293b02374a82711abdd1ffad
z30b82782e7eb51074bc260211cfe55efd52f83ccd516774b026cc0c7c79233d65b538d022c6fbc
z7177d7e41f08f2b152aa5669de3d013faeafcb30064673f46fd8e461e992c53793c9bff6dafb08
ze43300d9c1f6680168ce5b18dcf9b1ee4b06fe648eb2c6cbb38b111a0b5d2757b563b1348c6cb1
zb2a05ceb0d85186667618c3e0c5433cf2cebe3488bb81bb00a78cb0fb533a180e08f7ea077c4db
za2799087bd10f1ce9d2c288a2e5a1f9d3c8628128fb80a838f46ebebb6ef4f5f069c10725f4e21
z191bf9b173cd3a5489f1b61d929cde334ac39aa0e1d3bc7d9d78b973f01c9a863de8f9399f26bb
zb5314bcbcc82e17c27d12acb762cae253a8bed7ff0adacc680a21dab1de0799b07757be3087279
zb51f45a9223adbfa073b9709f8d277987c4b8e7099fa2bc3847bd17093a44583644d04a07ce325
z5ebf8754a70b294f87ea413498accab4c37bad4a15f617baf462f963394b8f237f540314d378d7
z65261301dc9ac14cce83766a21c6fa4a27197fd8af9c6f57b5147a5d0d72b51fc72be42ac6961e
zdfffe43cb4ad9b79300fe2611e14843297451b21f01be4dc6ef9d891b1fdab4586de7a1f895839
z18790bc7698896ac5c1e1830a311b43dc1664af882817410828a74678480b60e3461d66c7c4c45
z87ee985a055c23b550966de82faf592fdd0623678a08347fa0631844c7f22f787a6b2e3b9ee08d
z7640ea3cf51d9daf9a1461b0efb676f473c9988001606e9928ab136af5d2dbfdb49b06172059ee
zedfaa142912b3f9a27350d22c49e25c6a3947dc71f20904d5e0bd2dbfe2bc83f9de6c62ec7f30a
z4b84ed8d3aff50c02d1b91dcd9c20a06171966995305169d29cc3cbe0146db1f326d84bad583f2
z68f1dde2e44fe142b2f086bf08a4b450a2d1c7b265dfff1ccb538b08d9204facaabaa0de2521d9
za9eaff857e5f20d2e3f8713cab153515fb3983affc0c3169415e3bbb9efd089e45ac6435752bef
z6e1c1c911629f96ae326cb8ba0fd8bf0e0a98fc936886240b75f1f7d1efae028bc4289b222677b
zf9fa1e69d7e56dadf3ab0e6d84b6f0061bd4b2574903204daf64b985e3e0bf994708f5c3024466
zb26dbadaf7a7082b9c023ff2be237fffbd2e66997681e05ef252a127bd447ec31ae27046433b34
zf0d29618326d826bd01999590bba4b5e5f9bf46c3da79cb77db368662282e5570dc43edb111167
z4b8fb56333367172adf32834bac043f1024892cadca9f74f52df728bce010d704caee05dff1351
z549ed840c1606e0a26352cde8f534908eabd463ef3ec1a9516d928bff8a5c801f813fbd78b37ab
z6bc3f96d8dfbed0c09e7f18d516ff7aaa3d231f82b9bb7e661a9c9124f43e4718b87b0e399694b
z1455e6fb3d5ed389854ad62515e5ad16bb9ccb3a6b70b3ad17664fa5364afd065804dc570d9f9f
za9c5d71b69c0b3a89cda1f79a7cc7627d979d022ee9d7c9fb4d96b20b51b75b87b455fb9919b1d
zb3a77930d45386867bba5eae64bc20bf362a5ac7b8f45a05902d6369aac9b386dc30093cb2cec8
zb60c2ac98d6076e6583f70c0c6ef834f9b4ae2cb11348f2509320dd5bcf0a73659c7a3208b566f
z597af137bbd8fdad9502c7be61d80a609d19af665b17f452c333188546c5d03cf10c8a5a07b6a1
z5ff2d49d0324765144be9f3a74355cce4bd50235b37db7616b5f367aef280b73fe4b6f97d475e2
z596fd6bbd24712c3ab9d8e4b1f7fbd1814116a0a85f24742e0251da84124f92d693e1eb61338d5
z2f335edd83f3d7c614ec20d188ee76612e2dac3087be0355c33f61129a8ddc7b82570a7f4bbba0
z3ed3ae7b7a50ca328b653c92a46b21610a7f51ab67e27d5a5cc0c4efcb53d783b54b6858abc0f2
z8feb0f24c3043718e6e6431c49cf434019ca6ea827f2d4e9d57e005227e24adb0f5ad9411ee7ad
z57d04de952bc0c62cc8f1cc4cc23e14f7e811a27116ee108a5fa52fcdd67cc3c2dd0aab8258951
zd97712f0d5395f24d8f7cdb0b9dafd4745967f46b1f88a2ef7a9d3ea4b25566e911fafc0d30cea
z366ded18e272e57988c9e523804e646d0f850f9723a94dc48ad32095fd45453aedcad03800bab5
zf37f75e730e71c62d15b1013a344ee31b2cdc4b7dc2ecb98bf65d34b42b4f9878492d57a79dda9
z6414bd9f464b40f196afd163a7656c23908f2d196cbb84b84a185908c2cc0cb4b7c542dca72153
z0b829549854c81f594cfe598e071a9d6f5a71049bc6eb166016a70b959648fd34784d8d8dad7eb
zebd1a1541f6a06990389c868554d949ef80d9d42441c7301d2f8c74e2320a812f326a33f8b456e
ze00c93bc9cab521f31cfb8eb8dbe1061f29f22fd806dc7d230c68d44100db4db102d9c30a0c9df
zc09f8c97f873d64c44c45e5b12ea9bcd3d1b0d6bd06b0b47a89e7054b379bff639bbbb5cf5e176
zfd2e765dc73754069f6f4a717f3683fb5fb1c99b1778dd9502e03a8063247cbba588169fa513bf
zc176ab6360073be3d29631fe2330580c2abf7134ebb1fa16b43f15124d5e5188ffca010e9d8934
zb65a25d49d1ae11801890dfd491c4f248ac289efda9384714c9e5c7b90ef756c0de0c0601d81ca
z1212af739ef6d42cd5736f3355ec061905768d9489a16057494d998e84204d2b02aedf1afac8cf
z1730c84fc5e4d1b406d1df51ebd86d4757de272ab8c62a879ef08bd07747d46932f691218efae4
z0e276c141877b1928e592801942cb2a74fe8fd6c19ea6a63621a1461165a0ba70e6e2fc1c29f09
zc8b3decdd38a8abd7d3c32add585062aa9e9c61f7c0d273571838539b143e071fad4df3aca31ed
z4533497d21f851732c0efc45a98d49a0cb3f9bc21f8165db48e2c32927ade7653d4d450ec5f3de
z807ada1953a744292595ca5427df6b0ebef47c24b2c3190673e4cee4ab9db5e397b4b5c7bce00f
z975b9323af5d9366b0eb3de2cfc519de978a2fae1ede91954260d49a3b9cdbee4fcab108ab8bdf
z9f4c93c25f44c6cc8b0a2ee515535ce58c7c4f3c83aba8a2cc6557a963ed226989b3573d44bcd9
z05817169d19e0889d0ef52f5603cc6ecac79fe19b618a3fd92565efac7c5f6125255bc17919dfa
z56983d12ef35efd190ce7fc23f01c72d4812b31c0de422be6d05e69806bded58971b7fdac36c16
zd3b93daf2e36ce3ca450900d55f1eeb575621055e261a2784ad12ecccdd696401489c0ca45de10
z3403258c26e268acf15c56b02541e9d16a77a809cd6cd7d194f1e917c97d8e648252cbe084aa52
z764daeee703d9e8092a7c4d7286d3e6fbfcaea6259b2f222a756b254e9b41464384921ddda4af5
z876e3e082cde5313cfc7b664a4100d636a9d750b34234e99e642a570b933234e885a7029c3b1b7
zfd379fc89b7ed3530b05fc46718bcd79a00c6633fa4e24aceffe1dee2d3f48d048723600c6d208
zb3f61b91c57cb48eae726eed67273acaafff1c50b907d4ba16c65dc59bae23208c09c026f1e327
z258805318d99f2ffb98a357a2bb1e0e33d179994f20e5d5e537c3f04002d50b891962cee907493
z075d7e75da31bc5c9a55bdce08109ac47bbddcb40d93ee34ab90bfd58d7fb4c6d10f7f1cf115f3
ze4688dc650202d1d2a01c8278eed2051cca145936e71161653abf37016fbfb88dff103636c7afb
ze195035c62a54d7af1ba36658831fe75aa6b1eb4be159da6a0260817f9fa61f0f7bc451150fe8a
ze503a8b85374e038063f28731fd34e22a9062c244eff106cb4f130485d5f5383f0424fea036f2d
ze41e705e5ec154b70590eb0bd0a8f4b621e5ed0df17d2cc3f49c9de2c0195f8151f40045218d12
z1c320e24ca8393ef58aef45a3678030ca4277d0a0c610e00366bcc875328032525eafa379788e9
zf4833e0307a29fc44e1553842051c655ef2c9a9a48745eeae428b34ccc9c1a5d07908d22748060
zfd4f9333a69da0a8b9eb56163d3fb331e90b241efa40a4880384242e975ea3d3f174e0024a0528
z941afd0c4ef4209469d5dcc3aa82bca94401da7c04833566bb0dcd59e60882b85ad003bf34b5cf
za9367173eb57dc6204c8caad7c8f82c47eaca133d7bacbba97f5b3748c1586f087d1c825ed3fe1
zbc852f21cf48e5b50b07fa666f44df7fa6483e26d58476917dff8f0a44cafd913b7f09dc1a3615
z466aa13eac135f8f8c4e612d462aec4e94e9bd0cf219f3ea4a011700a4e742a87ca98625eb2c26
zb12ee337b24fd60aedb78aee1bd3c67accd60517e55895f95fa41046bb64134567037cc3104298
z62d2214dee4b4e499a9c48dfd4742955385286bc3430540527ff9035370bc3aa189172aaa9513c
z23aba52402bed796fc58c3ee723fbc1982ab9e77f8c93854fc7eeb61e38c07724f07a34cbf284e
z1f763e6b6c3f606f9dd4fae7f350dc9aa3859283f0965060ddcdbcee5be73c86a7f670f5a6eca3
z3953a2079d4610793f8c95f876566c73be00d1440a85c13646f8326f126cec3588c500731be5f8
z718db4b3a68c7e8f35ca9ba53b8f3e013957e5338c83db7d1ad35d536633340066d373cb798d1e
z9c9c3f4a1d4a41a91cc5c78f03a80f090c86bf8b60ad62b139c2a72840c9e6d0e84026833bd988
z8d17655c1640c67d9a6454b3edba9ca7e85c216967bea00fb3b013a07ef31ec1273315aac2cfa3
zb6c4f0fe4e19ef577fdf8960f571333375886488e30cbade875f294fc862b7b4ded618032f23f7
za35251c769d3557333efd8a19befb858d17972a9adbf6acfe841cfc116f2ae6e1f5f0c6507970e
z68cbee9f6da38914cae640232f971fc541e3fe88b402400df29068fd32b7982b0e51c775a44cc5
z6fdab682328ce35d4ccfa82bf4e1035c29291f87b34ce26188272c112288796bf17cef66513232
z5586393394b54c933172925dcf68c4353c31043a9ada7c98600a67148ebffc98627b60a5f71152
zca83cda6401295d88cf2110267ba471f49de190eeee947a4a8db568d983248fe3d250dfa23e1a3
ze6e273cf01df5451cc1e7e0ec8aa8d64f4428c211bf79795501d7f32dcdf79e91773de0da9526c
zba99ca8fde3bbd5cc5778cd954be4bc9b1ae0ff7394f69b5778f4261ac4b3086c8e5d289578793
ze80d32bc22a79577ed23e744e441fea821d828426d1ef7eec57e11d115e2e29b6143a9745eb662
zd5150b19eaf945e3e736a5ddc03c0698232ca274fa4a1c605beb691bf633c977de4364c081bc7e
zc7af3bba1c54a702a07a9ccc6908a7598b60c450702640ed0db3a6afc8824ae04b4ce4c5bd3e0f
z0a768a02d5836786f7a7ee00ab810237ca90d351eed574292abeb65e4582c33d1e26e9089cba3f
z52246adbd27fbb97aec0b77eb8348119b0640bbfea20b80dea599df0c3518ebcd8943f847c901e
z563e6df9c678d5fc73ae04694d3c230eba04acfc9219a533977189105d1a00b62211d7514fb1f5
zeac4e877c18df6f1ba355cbaaddaa5f974105a7954a7aafb8b02cf8181ed1f4e6438c64efed0b4
z863ce9bc2026f5453c05ba7a351340cb8406f50ca98325ebb642b6db3a0e0e489054e52b6a52aa
z84cdc16c4510929a168eb08839827d7cf7281987bbdf5cbaaa504697c56d513f7b169f86a3857b
zbef6fc66c0815df9ce3220eb6532acc37f3c3a6b2755e8e21d1ff5bc90b2595b90f931c9dfbce4
z435f83676bf57ad938013719066f81626789f7c673e2930695f340e0da69cad7bd541cc025fe0e
z6dadf3b27bc6868b68488c887200e4d41144ebc140fd7d1d6ed34fa090a9cec8e4dd0dae2a0a08
z5ddc5fd868fe01ba835ef3525ad6674068e4aef0153603a983df429e9a8d7bf0ba38fc6f0a8e37
z18bd682dd59d90a3c782596083f8f906a725740e4b08877a144f999e74fc305db885a833ba9fc4
z26e95a24f2bfcbcd10d1baa69b7212ba30c78b44453850c775fc1ee7c2540620f0c5aa98df6bf9
z3ea26b8ccaa4eb453b6416ddf292a0b40744b1b5dcd6bdb6730b3920113244bd04dbf2bb358437
z15563fc648a9367dbea8a18dc4a2b178109624601bc57d8018f6ade1a315251a53ab464d8bd780
za0c786c01180281a5058643e5c37450d369a4798e64919327b11ed369abd662157a0dc90095bea
z5aad0ac92b61f485838ef0a51cb7f0c8817e47e4f0aac398e318bd089cac396477f578cf9fc800
zafdf42bca2a3a187c9408051e3e0a731ec6a74aee55a02ce0516f3994d2a77198ca32af62fd1fd
z64b055605c319f78f5aa9c90d9a48b0b8f0858a6600c3dbe660b6523620c199cab29c4a4c3b316
z2a9dd7ffc760046e554e75bb1e758a64e7ea8ab2305d14bdade90504775d6de5f87f2b9361e564
z7116d903d7031fc556663c3e5db8924cdd89878dab4ae0a1426b9b615c681280f5d22ef9b0ece5
z365377c9b6ae0d896855cc98b6ebf35147ff802b949ed602c1f896a9a7117d9d5f201de567865e
z4aa9f4821cc238218889a55a28f72d7b85634368bb042d130519aec8c3cf6587bbea04e807d57c
z11f9a214481f20bc5a027b3013f722abf226300e1a9dac419a620c328af918095a77dccef834a0
z09860378e3c3ee2ce8a7a93dad2fb6b221fcfe2bb37924b69d56da81c7ccc6fbb53ed27b0a7ffd
z21124ee4060c3c6a0690472f32910da27d385a4fed1d6523d6f1f110401107170f6e0f79894234
zeeb947a2e8a897b36d356ac3cd0eb0d2fce3a69ae274f6cd5719f5d4ddc87a0daf2fcda7eae0b5
z14fe08205e1ebee602437561637cb70953575ac22395d14cb668cf06bf4608477912d8987b45e7
zbeb90e553c8ece5a38b66398b0428f0cc4532b9ee48e4f8882e844bfc155a0f3a4f5da726c4ce4
z9a45c84fb68403da8a4723b8f7c879123065aeb3ace30a3963742d2af306dde61e60fdba2c1cad
ze293e3eb91e65112c3fa46024a8696205186e220c4b5b1a01deeabef99c0c66aaf9c1e27e4d3ba
zfaa6bd78108a36fcd7a37362f1e0a62e73f4388d80e0f5641fff4c60031aada82bc663fc44947c
zb90ccc9589291628643dce39455e42b8d6070e2331c2034491fd8cc4daa46e904d47546494b34e
ze816ee7c1376d757ca1ee11b125ce63f7fececbb394229677e68e76b544a8486bef0925f82a15c
zc8468767bc6bd4c0e7310a06067ae90de5716b2c5e4a80aae4bb2e34922f6df5f5712f006cd3b0
ze8d4e98d73486acce3e6370c96533d2ea0e536961485264358298bd5078ae3b7a12d4ea2ff10b1
z2754069b0e75288791e55d80868741c6d91242a74a2fc0bb8432fff803f4643ab47a65918d6a7b
z2db920959168e32ef79b66e81ff48418ea51fe784ff30bbd45c4f6dd13c1fc8fce79e7598b6a82
z3a54f1ebb443effc66b1844735150ab711030b63b55db4e60c802026701a45b1a3f05036c01bbc
z4e703dde6bbdff01e0856e396500d96f08a634c2dd0e75d926b9eef57041d4830a782a02b9597d
z21f1b3529c320ae577a684ad6230e06ccc5a3b86befe707cb3fcc61e726abfacf31c8c15566139
zfd578eb81a1013f8bfba4ae7a5a38ee1158297feee954e8daf98144664abe8115da847ad80270c
z460f74a07c9320c11d062603d199292c440bed2629f6f365e9dfd88991e6b6a11dbb7736decf20
z6abbe81fb40c20c247feb8c1ec318c164b2085b4d51fb0dfbeaf5c981a8bb716b8a34123d92da4
z21264671ce3c5d4b1efe2ea9f57195b2781864b3fa907440f501a0afc70410829d38c91e1ea25b
z9561ec36b793771b3f52bc58eb46ef2de9a2eb856c38db20b494d66dc04618699e4d03b9e02c00
z0ed5fcc81a8b550899e444378a27fa395373a56d3feee9d6a0a740c80c8b798758d63f27bc1254
z895f562a7850a7738478862d98b34d9a1c052e49102f72659c283e6b60b3eb79403f3353c3b61a
zc3896cfab2006741f25132017ca3be648e932e0610f022e22d1cc6294cc420cc7eb3e676e9a800
z91bf4ad068b7cd6d0490ccbf47666ad5f90537fe083985ab8cbc2d98837840a266a0a66cdf0c14
z37bd972cacf101273b1de0d3714e090a1e8f074dda3ac50370e9a26465378f817977af5c971790
z8691999b06f11a443ca603c01991ea83f7b801477c72aac97e6bb1cc4434e359dd36dfffa11d5a
ze020595724dfa7e7a9ff1255e772ea36aa5f3841224496bd7ca1065a6952cadc6985c998b3521b
z20a1e463cf875f61321235ac6965fff12281f28e0d4a749aba8aaf98eeb1d18560ac5f5c36b5c0
z3715105df48f276ce0b0e14ad43997f437dda285f9a923173ad86f819b2721e72f8c6df8ab840b
z3b6e6e35ed71a2e8928d16806783067177c05c497a2ccffc71b539fa93e6a7b59004493e439247
zec59639153ba0382803f12a0bcf091dc621cf1fb3643f86b8b153d4fedbd27dbd7eca9adacfb52
zd04caa3eb076641edf3bb8e957d6ea44afad0d2edd03a6872c6ed57a67cd82dc789e541d3355c5
z048ebeccfa88956f6ec37c91e33e11270ca60bc87118f02b9c02e10af086008eba37f92160f8b7
z062815e566a4a17d316e526e12e2ea69afbeedb075430cc928558ec55ff946dfa77162f652d6bc
zb0161ec935552c28fa6543a43c4d925a56e396891ef5dfd460f5a84f2010a8d076b9b7439a2cfb
zaaa0e50f2d45c261981ade468fd824d25d8fbe4b9e598dc8650fca7ba0c112f99ed6eb87a3271f
zfcb88dda4c59679dca2dba78346cab7016178ea889d36a74e86a5fc4c8b9097b7b132586ef4e44
z5bcd33db153baf0b10d7aa600b6e96e5986205ef6af4bb701e39dc88a3365e87fc861e7c3145b8
zb3bcba2567808a65c81cfc73ea821212620c026cae5c0ab804b9e25908c49d68cbde2e71647052
z1dc064c13064c781d16f987fe1edd05254d32550b01d012fb1ba13497369fbd0a8ee678595da1e
z62acef17f717a985590b86c145dec130c30f8ba10c879efdbc7b6823b7ae9a00ea50021dfb7754
z883e44286d6d6854235e8147803a42cfc76bb9f09987905cd82c23e2856d56e75792b52428816e
zfc8fd6aed786567a9219be64a18c448a91c3af594d66cb691ddae7b9544a89b70b1136e42dfc63
z7c43bb410635f84af6f7e63ed6a9050b612e12439e2168577f31c4883e91ebea16a298bf4bfcb7
zb7d5ae0e8128a3698c5fc7fce70037f2944af475f48c79f73c2132a0e20ca6da7043c5f47896e9
z9fef1a00b66d6c36bcd2a082bad733dc3efb13f389f2fc293e7e82f2ffaec4214686911a747261
z527d395276f2f3733c330e2576612b3f5eed6b0270348843271e8fdbd42a2f9bc1e727e4338e02
zb96f1e84968d0e566284fb0517f85370fe37f75f32aecdd88cfa25ca92d9e409f773d2ae036a0e
z7ecb4e1a73debb50888f5693b864e039ae1c30c7b66fc7e22105c637fd72d697f2461d8ee21806
zee8e7978fbb3520d200c3cdc3689ae083ac1d65009d922f4f06b1294e122a1cb30e4f55fb2d842
z015998e987c017022440d659e93ce47dab8d465b452ddadce55f232e5094554022cec9dee46ae2
z5ed29756ddca8344f55490c84c1367f9311b5c320a5c8772b641228ef884f3199825b264ff9d2d
ze43ef2674b05ec78c07f8bcc03b3a73db8702b50e42105b1c921e8c77e9da09e29a2be5b6f8ac0
z69f45875e064a3c15bc6782df6e6c07b0bce5117a0105675fbfda84a550defa04e05d8f8ff542e
z8f3250a042db1e5d42917696079b86f1e6c2c34ad48c5843f9b75eb73d399494e53541592b644e
z2044871ad5619dcfddc6ab7093f7cd88a43206a69ce31a9034c87cd5c510129132d61c315b347d
z1395fa4453a43ae2d78dad8bef09a28018e132f4abad5ad831323514540c2cefb5e12d347b995a
z752941661374d39979cd67a2d220cec8a1362ed41c434447c930cdbc05501cbb8b9b06099f99ac
z08de6d019ecedcbc94221868acca4b440efe3074b90c42741b84d2ffcc0eb0478f2306fe4b10de
zabc061c526ff8a3816da5d3f31d45f38b890f746896e525087220e97c17086d0b2692856b8f370
z32c8a63d4272099de3539eba62e445fc9fae6cdcc3bbe5a3457d74934522e6ce93cb2d5e666937
z9087245f88ce54e466fc38fc95d0e2b4a75265ca036fd83143cc9f6114951330164d7d26e477f9
zada668b4fad95e2eddb55e85ab8d6e6dbf5b38b311956bf9b523b0b474ca1d84a5931165abbd19
zf012036b6dd89065126bb8663f608c42be14b147b6d1ac2025be174923bc4d9ffc77a73096ffec
za34e3eadf4bfff946ea3c888cdea4d78b8e287342993b03e1175043f9f30011ad814c1f1ee4365
zab55bf162d5b0705305a55d9b5c58a89614ec32575025ab71ea0592883ec97eaf9e73400b14991
zdaae1c709ae00f4f751390c1adb1944bddc48ec40a0d3132e0acc95a71777e83744ce7ad776397
z0bb6a527fccdb89de15b9607a8ff5c51223986084c645848d718a5294383e35c6aae3fdfa47b1c
z98f6d2181065de9d24aaf32571b84b7cabccfa57b68a7d3f5817bff061939ef02e5b524e4c212b
z5a426d556cfd5a9481b8795b1b39e09ae62c63d562421009831ca3ee585eeb4189fcde995eb7d2
z15b0efdd9821dce356256deec144b3d19857367b26132c3374073c8799aed24e8151f98efa660b
za6db9f4cae4da62d5b95afdafbe524eaea6bb6b185e3825717f3b0083071782ee63580bce3428a
zb26434b0cf6619f8e14da09c453324a4eed0bb91b63eed360631c11599af027af900749b75dd39
z4bb92f02cfe055e1fcbc1a6571e2e1020925450bddbc9b77259205432437fe628514e0c11d887d
zcc92cb9059619fac7ce60d6843bbd66c76d5d4c54488ea70f6dfa5fde1bf1f7f7b637773a6ea78
z4fb8488eaeabd7cd928b7de720b0625d2f637f4da15f2fd7cf9be6e18fe2721d4bdfe464c2964e
zbef9ecfef7db72afd4a4765084f83e103ab42991037e97b1ffc8d4027e4e3f49a446e9cad92160
zdca899dc64d084d7c1dfba8d55230fd02d8c51ec0597040afb83212ee8b5a25b2195b19264431e
zc85a19bf3bb602f15d46805b5dfc4793966d894b47884672b0fe0286e428475057db1a45cf690e
zf77aa80c3dd3ae60cafeb85b4921f4663be25ab1287fab3da358f59e062a7ad135f70f180538e5
zc644fc87ab2f3806b6abe0165e2207c33fee1d2685b256c02719ab84560c543bd01d661cde35fc
z695c615a3d78a0c1eade238cae82f8c03bf5d1704d62c49b08ff6416b619febf287786bf4753f2
z897a1c372ed625529c7c5eca6a4d4922f41c2dcb330b56ef94623d693eeed54553005bd8260ce5
zf4630c5b8e5abc3227952e4ca69e34a175a65f19bd1e5857efae3429502981e6a2e392205d04d3
z89f95c174318dcfae7aa8c67f6cab3feaaf43bee1d8b1cd7cadfba89fcb7774a892ada4a076348
za22ba60dfc100bf7184dbd8cd8c0bccf919f9249b76f8a1df5924507763a3dfa2eff17eabae0a7
z038a93d153bf54c2a5a48755d3e2837fece43336546c792efcccdab6552d2de584c057ed3f5e92
z0645a8e6d969d7b771e6e0861b9ac5677798cdc9005d11755614e986a64f53b90d0fc01b2018da
z089006e14f574bdffc026e9bd272e80cfe993e5630d6955dc235f2cfbd799b446109ec26a8b6d1
zdb567f49a6ed8319d7b9b8cb1dfa9376cc04e7d7ec845fad757f92d2b3b467af3d25737125f77b
z09cd98777c511771e054bbfef0f405bcb2495679e24b15835b1529d7923b3e986f7d58460f770f
zc1829dcf26c29ae3633de893d33228a32ea277604e7cc49a19643c16b0c68951d2d023a0c7358d
zd838c09bf0cc16dbbcfbbb03bb123989459eb2b446db17b9027d72ffaf70b9dca78ac34735a2f3
z8c7954af34d6c34f455854b02eea4dca11594e50c6e13fda3ac82982f1409dac0f504869637d3f
z869d29f9f45a662fd7b4a042eef9f0a99c0f46dea01d9544d99257dafa9e3ab140070adbb3327b
z0821ff41f83b8c073dd7413c306bf60dbcd1caf8937e9647d01b24ed16dc4a347d49bcbea72247
z563ab8eb6b2efe186ae5b703079d2578f1fa27e6c3fc01c7c3f45c94de9d135f414c1a165f83b6
ze22d35cd72572c0c3b39d5824112b64557087e1dc1bd931c56a475fe28d7b4de6f0dca7fb1e8f7
z1c64d32d5895120aa8229e1a4bde010df0bc5052f96415fc5f7c1867cfec7ac0663b289a93ca07
z72bcf042e25a1d25b74d85095e13e79607fe56cae2cf70c2eebd6f52d533b074383034998f48a4
za99e776f099998d6121edce6ca956704ce1442f1592c5aa5aec9c44d839d0231190abecd642e79
z6727478cb42e50c3af419a7c62b54fb5dbe24fa7f1e06fe1bb29dadc0a931c27447adb20b001ae
z0582684da28f538e01dbdbd433049abc0f9c040f41b1a80689773a2925429758afe3769c780f73
z1a39ffe3b023de6cb6adf6558ca576b0eb3911030e9f123ec0d996c1936a33579e071bf3b2dc8e
z3f0d5492c1a7f7621e05e375f82bed17e350ee3ee3f89d0524cdbcce0f6ab9d52a46e13fe682ba
zff36490f5c223e8ff6f8dae21061c085c221399ddbe8041215a4469891254fbfe3918ea8c4a574
z770ae80148842439a6e99ff1e66af4a9aea45c7db72d54d9adad95eb9ff6c795d618b474b6f9c7
za655497afe0022050ed2a1c4a655462c61b138ba1f1a57edcd7c87a38b8b005b43921b04a8b921
z873d10a990266d52366cb75dc1b0a21dc30253fc1cd5315495e0edaf1b9edb16487cd06af2bf54
z720df8eb6ffbcc31fe5d7ae9e97e24101ff1f9a22c16c3ff919ea938dd4784459d71419240bf55
z089942e1f2b39863c4eb447b58a26761b2e6df9abe4e70eb0427fa3a55d550c4f6bf68c85afccf
z559f0680f50cd687fef21b3669258b215e6fbbc6400ef912bcabda5f4a87dbbaea213f862e2f8d
z85f120c3cd917449417ee09de6798e628877e46c041b22c2393bc836cbc70d6bc191f888b66401
zd7f5588567d1b9fabe2ababe64082e1e065846004d7917b8225312853fb6b64d8e81af8b49b0e9
zefeba061ebb154f2adcb9f50a044939db5e8b2aa7ae0be68be3593847447f88079f98a2afc149d
z86897c741ec9932e419fa13e5eeb2912043c60a079fc07c108b307019fafc91fd509a37378273e
z1ffbf497fde72b4f399c027edcb21de9b7b582d204a01bc5eea4e703cef700e43aee9fa5fe95bf
zdcdde46a1d6a2bc0352ba17610a3b778953c4ef5bbeecf3d036b77cbffbdce7104fb20cbefa3e9
zd2275c949e65a77632482a89699971ebacc42f92d123c8941c0888d76a1f93159f986531a97fb3
zb94d86ab2be5608132aeedf75ec4d499cc5942795702e7cb9076e27d8534d53e52aea867dfe6fa
z810b11d9ac7174582b069bf8723a2ab1a7616396becabc81ba46ca8fc5d5244526ff2b6d3bfabf
ze9c6428428d1f7e09fb68c9ffd94907e3a4ed517c6e282d6417039e37bd2b9b506dc656d2b1b1c
z1bf312d4683defb2a19f8768121119585f351f0886d766b769ed69b1156eeb8b0a9107bb621ac5
z66be338f0cae5300666a280638a6e42397838e04542a8154976611197687959a309697fdb11099
z96141fe7d4624bb48808982c98f930590f6fe5d81479834ff2662dd4e71ad6bdd0f364cc2d45
`end_protected_0in
`else
`ifdef MODEL_TECH
`include "qvl_data_loaded_assertions.mti.svp"
`endif // MODEL_TECH
`endif // encrypted_0in
