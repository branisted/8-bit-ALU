`ifdef encrypted_0in
`protected_0in
ze74c34e226135848fe16db9ffd31815111b6d7fb642c521a3f628cf6da949865580b22efd062a7
ze90adae0e65e66a2c36a587d0a790699161455169ed55a01f2084f11770a774ec4c588039b380f
z6de9c5084882a40b79a175f5c2114b2b6d78b070cb806e1c0aa9258297f4687ab308bc470f0040
zb0b1de382961eeeaf2e279e1462520fc31c119af8f2b214846f56c2b3cd2eadbe4099496abff18
z15cec83ec4a77b868344aa20ba7360908f5c0de2a79abf8b3534b883bb12180f68b5d4beb444cf
z3fba8f13afb0abfe8fcc4294810f75afe452434d2d0f1166236c82f76edf1e12979f04bc35693e
z32ae028996dd85737a8f5adc1ebb94f39c940246e887647b64782cd7ab429b0544c173176cede7
z01dfb26b1f73408344a52b7e1f117f12bb9c8077b34876c2e6fdc085981637012dc9754765e1a9
zc512ce062e0b8fb16a214591f5c81e1353b900a611fe1f4886b57940b41b7f2ce99a7b84b04b90
z916f717e73bd10589c81e207ed77ec660a8cbed5b487fa50acde1b055c8870bd8676023f21ddcf
z9c98cc47cfa2d654ff1365d1f45035a045a66c5dfa827905026201628cee5aae21fb892db766c4
zb5b1406e11aebfd6dfacc9da5ec03b70c276807a3eb15e28ec7ab1dddec42388b9424ea285623a
z248195c9f894b36317ca6e59c86f11031163f5f5bfdba36b10b435d36514783bc1c6e60eaff7f9
za2b8eba90f8fd9a9cd7c932ce34efca1757e6b2718aa68644ba032b1bdd74efc688b935cf38d81
zb1f311df3e5b8e4d46dbf459c824f309500192485674c175e61de609f1c94488da73614dd500c3
z680b7fbf510ef6c68927870992ed3376661d943d2a929d90faac51228c485c2005ea015bbf306b
za52b2ed3688d7ece69bc3ddb93a45ccc73f6e00673486a8bcc92acb7d4412090924945c1f1562a
zc5e0949f06ac734085ed2107e4aa9e39ce4ccd2716381ae81c00f915da3dee1704ecc26765111b
z37c91301861edd467e17bb93d5e374e1e91c3d7ba3c326b7180905901191f995e97041dfe92a43
zac13264e5f9c269b6e7a2b22e5cc8b0ec5aa75177e1c8a2d5c5456d5269c1ef0d82494bce3da12
z4598593f8470c230d8cb82868e2e8926b86041df29c6f868fafd01b20d15e9158055c9eca0eb1f
zbb75e94bdfb4e336e8888b859ddc98e14841807274add30af47330407dc3fe4317c3617f953577
zd4f5e2050846fa11e22136fe1d04da49bfccac468a90087d714c5853724d5847e1f7891ad9c470
z73306d6006d0e807052eed0126c794c03087ec8ceaf31379819d317f9fd5324fc9ab389e92c9f5
zf87f11ffd3a7c0bad30910b0a9ea77952d05e3fba0d239dde3f9125ef3aaead1e1207717047c73
zb189fa783b565c0b5b80a8e5c3281139cbce0dfdfe225634179911f45e0cde88f30c27de391149
z382b51a0eae4d2c9b552620c88057ab506bf655c16dbabccdb73d222fb33195ad5d88137daeded
ze8768562c518640df73740465574dc1be86f73f1a2e6f160ac27789bd73ab387a4a5b882e9f759
zbc93c683fc934b63308dc97e65d7f7ee1bab65c25a19e9fa02b58d7835ae7aeb9892e4b26c83fa
z73e703e4bcd2932b6335711c60c644067a80c1373acdfd557f5c4d7aeac35376b50d7cc7760000
z277d4c95254538a49d0a0193114173cac900f719d72ac0e54202fc99572ea3eab96659b511538a
za3e89d7b9a64495b4e97359ab47eb6fcb5319403c8fc9f5cd6801e2e3a13913d1c481987e81cf5
z073ea5b7384a286591342a5d2f35786d6d66476e7b7102e8384907b2bbccc217a307c4207563cc
z0afd6c20134d4f0351a85c8537378aae9b6bacc3822d1f0f990d811de2dff0d0864b1f7809501f
ze82cbdd99aeb4d0be407bb283494ba9c047dc7ebe3b7b1a4946fbaccb15cac06e4d314472edd99
zc658a3651b4ea88f3facf27093d9cb560e28c04aa59d4b6dcec2d5d0ecb8fa95b6aa37e114952a
z747959d7cfb9bfdd51b60eaa90ece423fcc28e71c96924832338264cb86ed46dbac8a8fec1504f
z3579f2e8340af11f48f042b656e761ab191a52dd3861bd6f9a5193d82b396ea8e3d7dfc7b31870
zecc86593d01316df27402231070d8cfb01213b2bb6ccdd5f07b6d0c3f823ad0b65fce7d1ddd9ce
zb54cc3f24876246973151348d7446eb6944e36bd15d52c06827e96bd6f0a12cf4469fee6d4ebe2
z6b290ee4f55be5798ad8b8d51354b0f9746000676a7bea2b4b48b645e175c44b896f14b0e98b1b
z3bafc1b82470f9c90c3151b940495b70df23b76f7a95501f45e28f26029db6a444dcab02f0648e
z125270ca3ba49cdd50eddf505c9c29b78c7f05538af3e91282ce8b77d44978fe2d84be8d231434
z3ba5f81ddf669f5228ad01c1422ac6a527191375e2c00cd7511b10fdfc23496a32bd5abcae338c
zd8b85faf8f37fa228589b13cc7aaae04137c5887206787d517c41893d9ce5ef7058d32be1d8dfa
zeb537940e411ef354afd4f2a3e0ec534ac720e1499c8dfbfe9180edf954cb66ba1d1a3eb9be8b8
z00ac90ea28cc37d619642188378a0211675a8e307d3a9583f23b430e7afd53c5afa6e32aeb3bcc
z6317b460f1fd0f41aefd258011e62e2e5adce40350d7ab4521f0a2a105155a051465c8ab2febab
z74417939597132e29d61ec3c3902717c00f3217f1e1ee14633d0c6749db5c4451e251fe423f32c
ze8b2f0c752af76bd25acb99d4bd5ac7a5262e0ed3082000c910a3e59b2ec163cc98b2f906b87a1
zf5ca2c2d5dff30e41ae88ddb0cd75dd9479a6329177c1ed32a34b88d1c44d7788972f963c05f14
z1b69f44ef838f8ff217640806bcbe34f20285235200fc8748704db4abf0294a6aad4a3e9ca492c
zc1fac03e39b0610dde9ac3d8919656b7829b2ac83dff081056679aa54ec9851e255b69c3b5d19a
z7e798979528f9f63bd996af4af67abd07a4a27fa2a9e0f5737593f139d8435aad0f7ecd8ffa3ce
z333961b8053c994c893594d7eb143b21ec2bfb1fe562127349ed87bd243bfd24e11a90a4cbde57
z3be54a5ccc5e7b5ea45c80f37906088e346cd13322f3cbd1eaeb3aeb9b049e75be805808101512
zdefc39a57534adb76d29a6456748a7e409479133cd69c92b0ce4882c5762991fa6f260fe602b59
zd2d2a7bf4d4f08707536cd9e6698edf0ce08ab9a81362057139258dc7617ff5a9bb6eaf1aa24bd
za116c907ca1fb3abc9dc25113bdd1393cd7e66e4653e642be2b774bd8b9bf6ed744bfc970c8979
z38452675edde38dade9a4f528c80a691390f32abbbb3e07bdd2ab75a668d9a0bdc61ae6bb65ab3
z300fa9eebe5a20da234d5ad6a724b6ed0d5abe7de4f3340004a0fc564cf194996d457c329d1b58
z74d7671f9351dc714ae2c0f130c111c0ea6de40adff0750a11f11755a50a42b214ec2f9e04ead0
zf699cbd8618b2deb7932b5b8dc4d981a0a7d91da554b99201554f5cb80e638bffcdd30dd426caf
z231d79f7f68eaf0ec2e22c53aafe607a27c8c57b0b7612b2f44cc723dc85e3711b7e8725956464
z1c0beefc23f11fc7afc78d6067f54405548f3e0ec1e43ed012c372cbc9d3b4c3d226bcff38a7f9
z62c9933cbc9b5d06be7f54b8fc28e8ef6480f4915fe50824db9edb806042315e6dd4583c308afe
z6ba83ad9799183e8a8d29ce47e7c861e8b99f21a9164e9cd5c3c382f10e878fd53fc50cba51197
zc3b2457b524f62ecd73fc3741a57651bd7d9782103b57acd16b8eb2a921bec861f29183420974c
z183e4ea12c60a2cb6d163770898a168017e52ddcad0f16a8a237d1f4fa273b17c4483ca73fecee
z785ae70df2080362e6886e6ba2e6239b19a6f1a01dd8b4641da962f9656dbc40659373e6aae62d
zc30a40662c02d934c6afd4a7751ce557e21c0507266fc02b605e7f5a64460c59d297ad357069d5
zc2ee133eff3aa48f54b72259552f9dcdc26ac03bdaec9bc1f2f9bedc130965fb975a6bc8d33bca
z69f861753a6faea4bff73dee7cc62304feffccce2ce4b0b9ef2385705c24d2a799131cdac8bf96
z447d2130d34dec1005ba1f4e1bde2974c173b262731607f8170cdcde1481ad27272962a8eccd87
z5cc493423533162e9933c67f5b9e3e5b862ff3af05f28fdea39cb89e35db6add63577b9750126c
zb5c7e7b1d81f71d3e77e9be4f8e0e526d546767e0fe7a3b42e58e3aaecd198b90009a0a295e7c7
z9e894a1857ac79914261b0317a792be7d02d9433e72cf8b597d2edf057c2e1eed6c9f00b6ad608
z66e667ec0e18a4276535ec6121e9e7d49acfd3f3e8e28aa704597e10949f9bf3f416060fc4154e
za3759852ffbae74ca38684e7176f749794d131917af7a73515bf51979678d38f2cefe5768ebd0d
z1b24bce4a13ce23ce8b516785041c0c64b21dd9f87eedb408bbbde0c167d5a911cacb896c12a64
za9e28b20b440fe3b95a140b3d736532ab7ef9b1dd031e1d84eb3c64cdaa773933e5a2215cff8eb
z6ada012409e705c880f2ba7d4685403b5ec1a93aaf99cf80827a7671e10a83c0aa5f8e22058bce
zedf4dd21e75c23b0e93c2f6bb941fd2f09b7a6f40b73368b878d1190d5b4d3276cfea14f294023
z6d9c0d4b1e021b3dbc276b83d5f4eebbef9eac679abf9e0c67d6ed9321bf481c58de0d5951bd14
zb52b37f1001d92da0cbcdf753af9db5f6ffa071786c2946f3422d1cc889d333d009e13a1681a0b
z9ad800bb98f39388f673b078daf21f02851633aaa88e4411990837301a001786e1b48dc6f4375f
z7f1015df6d5fb69ab5b29e394f9bb0e8ee28dafa42b3088bc674a6bd0dc8a697edcc18ed1f48de
z9ae4fc125ff9fded82604c66d81f278e46608d4c4fdfbab27dc8ab0fcab97d57dee52f18ff1ab5
z7115180ac3a191b66929f6c29d0ddcba69782ad49c9bb5219af88a4f8cc0ef847b15da8907edc3
z2996716f358de8d17b48e6e60a10ac06880a5e2a376902827a2176f6593cf98820d9d5a1517295
zbee3b14c74ddaf8e2dd9d25c8440a2d06eb2314f7d664b787fb65f235ac3c075529f60be788e77
z6317fabc9ec682fc6bf165fcd1d6730ffa3719fe844706ebd83c859455a87028b1af01918e3b33
z158f6df059f0411309b439ccd08fe7151440701ee0fb320a3d4a241f670c6e76f5236d53b867b2
z8326b6c30a6b19679a9ad3c840462174a20655d0c3c1c68458afc2f2949e3ea0181bfe4d2235e5
zdef59f5448cfda5f24a0805b68e6906ec0faf7d63d16e4f9e3e9f74431c2b8bdc0f9d27f654959
z0d16350245ad19c7a3902d34f16a62aca972c37dc574a4627859e37fb9a58d4ef34c9839f0a3d5
z80e6a68bb6d0b7678f743071ae718845e6f522d758b6827cbcdff54edadeb2749172c0f20366f0
z311e019fa1e64ac9ddf36898b3da96ae3c5079fe2814de2f68d8fafd1f6883f9256be5485075cd
zcab87d82df6d37a0db2999af332331e18e3d82be863759229052e861691572a0133e43aac9d128
z16c755dd1f06a960dc0328c8a631c583c2953a47d1332db21306745f967cfb8d369623ddd3ca07
z54f60761bbaf1932dbd9aa83bdadfc4f6ebf831537ec56f4de5d5e536e3ee94e8304abdebd5339
z9d8ca88059c2176f2d6493c1bfaa0a8c97e4b0993550adccd641879029e8def7cd26f13f7ed791
z2271643214a2822ba01c2647e72fe20bec3af1cf0650af2cf6d9dc1535b2f92b7f7bd777801daf
zbdc6a65e9062ddf9fbdd89fa9a17e854fe782e06575356e9c076d012555b3a0fbf34557a14fdbe
z1d1721356751ee092ecd254c119c9a0c46b5bba67c446f67288d9a2dfc394f527ed82ebf62d6d6
z87f9d6808ae34275fc81168d68a1ea207aa592feb723aadb6648c0b1aad608fa9c392d0f0079b1
za1ec9bba7397de043c369a7a21d163029e06816a5628a6e8bb9cec97f99a8decc4cac5ab6c6de1
z409a7c3795a139d692869bb9d721c468388204825accc7aaa6ad0e765eef6b9a3b43557968b05f
z300eab7e9b1cc0bebe55725717bab5ed5944e83f6e6ab0e6550dcdce25a5bd4dfeed19ecb7a182
z1df84e5e58e8d7ed15927c87931bca0ad05f44ab9f79f4517a5c80f36b18553751e1ffe0d57a5d
z1b5e7d53616b92e7a88c11990a8d94087dd5a11eb25c7fc1a597bfe7aa308459146894daa29347
z67e6800db3c6d7653bedbf1ec7bffcca265621089d99fc44fd19ea56e632853e3d69e13e4d260b
zac7bfc73d81aa350fdf7323c43e00b4bd91de044641e991bb939b965413695a45aa6819a659787
zbbcc9f98dc1bcb1ace3e7d16c94c2db1e5576ab9e4a0ba873430278d26d1e8b410bbf4899d0ab0
z5d052886b43071df744a34e4bb99f73aa8502d3f774779d8bb84f2ad6e4311ee360e1edfd2178d
z7076d02c1c23f73358446bedf8f13bd6eb0fb826104271dfed31873515801972fb3c571e4e382f
z143725fc822dad72bffad75c1930ad2ebf8bfe0f32d44103168dde6a3096e3915bdb90d35ea1ec
z1cbaa2c73a4bcf041bcb7cf1db2ac9e73ef9076396457944b99036f41c53e0272a1f50f816ba13
z261710180afb30eb92a3fdb24d2e190969a744c117c36c5df80e4bffb7e5535d8fded71b96a5ce
ze77225cf3829111bd48b1e90e1c68b50ac2a014a5881b0e2c50dfff08e765e2e4795e8c4a6a4b0
z8121977d3ddcd583a081222e11787dd8a8791bfe2189f83650043e60ecc0037b0762159d20b5bd
z7dae3df8678129a702f31da337b2643b4a5a227fdac81c5a9277ec9b3471658f2f10869571193a
z0c0ddfd41f78e4c08f64e4cf67b04ce33dc4c53b6e3f68081046ad144e6447fd9db1b19a62a2b1
zc302f004fc5c4b72f5ebd1a2754fae0d64df115d14e935d8fce4d16809754ee2d5ff623da3ae96
z0df65179bfbe35ac71ab319fb5fdaf4b440128b475592bee5b13d31d3489a0ed7b1621addf9caa
z6316eeb5ca519b8284ad7809c7007c569dc0f75d88ea5638ab2ee6401cebbb5ef5e4549ce2c991
z53801f898f6bdf3631c4301ed65198fcc877767c7997aaf48cc06d9180ed8bdcb6c05131acd124
zaf8d5a67166fecd381715c1cd944713da6e7834981e1fa30b843266f009cbfe900f3d581303f74
z00186848e20d394afffc85525b1ac0fe822cb22ea16b88b9c8a808ca3ed1b2f6b40b624c6b12ce
z31c6b5bf23c14a7fab58db1c7ca9b993430839e9ad29eb79c18dcad53b7d27bce1a6b6addda5e7
z84a71c5d1769786b7b62bbdd5006db7ce13290c16d9fe0c634e6cc5e7c844cd7270d9fd550a2a5
z5bf00ed8b9bce513e708f2b20b87941b649514e6e6c3adfc90f5018b4b9990d02921b84420855e
z5085e58aacf8c0e82d21fcb0a51ff02d891ca15972d29628732bfe07dcddb3b8ce00b5d06fb018
z9ebc593a75a7efe942a232b65087730fb3fcc9f2ba777fd969bbd25e66b3e2a1296ad850bfc564
zf00574d7fcf6fa2317c9dde451f4ba6e5b7321c9cf87ce7c1524817a2254270102b9b79ea15849
zf520dca91e3bdaae98aad427f410037008b9ab3acbda62f7edfdeeb0adb85e862afa6636a4151b
zd9d421392a3a7419684daff01870dfe89481b4b236e669885675560001a55b37016f1349bf6165
z49c13f8a218c31a624662ba5ca68f038dfbb984befcbf311fa70e36f0db28d0a1d13a1e825050c
zf600195c11c21b4a835505549acbffa646a72e49ea882e9f6985d15928bdea0e43a8441b5f482c
z6addcf7c6395d3b07cbfdf7f6e882c17603aa6ba1f99f43be18c02b1088f84c167591893c34ae8
zad42188b0a22f84886a6fedfdbe19c70b24a0cf3d33714db575564475657f7952ecec361bb7022
z8e71f3c3bf9d5ed4681944e8e63ef781085beaee8583947082f63d5c2f45aac768d3a74374fb17
z41b841ff7b759261659920e502e5a22d5fc3b60e29e369971fef5a2c16e226cd0ead4ba32efc7a
z27fd8863b21962fbd682bc843f57a788f8c10fcef9aa91c03154cace9360dc6df5fec44a953c46
zaaf7e05f9ba2caa73ead7eaf3fc95a5a803a90fce8cb518b0b3572b724c94a6aa145eaee3c3e47
z8321aae07b0fb26569858aee07bb1a1d8635262e9739e77e93e24ed1c0d946e5b4cb3c9f56ef77
z1d3e3d87f57647df390227f8fa283edf64128d009caf10328c3ced4d1c842d4a0f6c935506d175
z201e4acc67de6d3741daecdf025af081d3e71ca7b2288704f29e895ca24a5a74485de1ac746a16
zbdfa4ae267d4f1d767c3b5902d5f2ae4f9f7aaa4c63144de71901b09acf83c77e90ff792f2bf5a
z0d7a5e7a442255ef9d1b9dd91d799830ac9b5b455de58027bf3e425a2456ce1d14fc0f7a9fb844
z4420ce1835b15b4c4aa2590b35f42b4be45908d9c0396cc6d9225e5cf5afe681c314678f222031
ze619cbd1286fea2861d8117273694cc825145e08f9247d0e95879bb96090d167804a137e91e58e
ze2cd57dba88df146ad24e8c5f9f2e36bea2e36551796ea9e0b01757288bd4ffd61acfdd6525da3
z51926f87eaffabab13b00818434276027ef95e702befc09b4b3df73768bf9a13367851fdc91a0b
zd04813b3437f023793b022dc482a47c7ac42cebebd86840bbe58a71ec69dab8bf9f266001680bd
z491fbbc7942720ab29b19c299e7c58a21a5b0b3841a025b3a51eab0ccf960344b06771e2efd30c
z0a51cec1267922e36f7dcaa7dd88d5736fadf3ae701f35b00128c6275174718f5d150990fa61b2
z6d3606fff595b50c0dd0201e68c472b84006a313b7c52ab37f5ac3b15f52e77fe2f770f444185d
z14f681a3d29f873015390100ef979a6f80393e0f331ca750bd3e9d1f157a0a387f1a190f3789e7
z3230e12fae06dfe0edbbc8441b4e5383a3ddc9573a19e93595732b51f271505dcf9d8ea0a9ac7b
z91168d547291854508f39593d1e7d05828c297c50826850346375d3f903d9b2ddaad316426c4fa
zd531b846e09bce3bc250b514a66951e0bcf5ae971f1bf70a0b614d71e28f76914ebdf0ded32b9f
z740262b654fd8159698a0dcc7c7f4b837e5825c36ef84df0eacb4533eef544565678e169f9a4c9
zcd977a1c0a24363cfc35b53c900d37b48e8ad5b5391bfa4bc1c3a36dd870e849e851c3144e62bc
z6fbafa731fec183f8198d76269f95e3b84f76f389f6dde0855f11724d180993cded54c45efc539
z2f95d31043d6e0f636910f1be43a2f5db9609c4259c19be08977a9fe6e67edfa5a6ecb6eef724e
z6a7ba12e4b60f53c3f4f6ce30ace96ed35e3e68d8faa3a4493ee57d57ee273192e7eeeaa0fcc86
z6feaca23e4d82619aab253cd9495582dc82eb877dc11e956a14373f4beaa579ee7ef451802c3f4
zcce06d0aa8c6bede827d5ca4d4b836fbf26f25b964b301d48e61aac7e251a5c0c12a09f7b6c67a
zd8f02033a205885282a9f0cdb0b4751d70ba875d5e43a349a13c0b8796b0fb8b1916a0e50ef25f
z3a2d526fcda353a2401d42449d482974ecd2e69b943f13e81844bf6584c760e77d6061f17d3a2e
z1f686baea08b6a4ba20ccee915f8ba2f62c2ab28b85c003f14f9be2072e4619e6ff6570d9aa718
zb7ff9d6f92f6386e9ed3dd12f67cd583f83847f831d16db8395eb13b4e228f4b11179c4dd1356e
z09a8ce92230584d775b52312066071399f922f12197e70afc05f8c8f0feb579c0ca0a4f6ddd713
za9242833b5e01871fddbfef7fd5efc130095e567d8d79050ab194fb282fbcda659ea0db2d4cba9
z228a05a4e833e6de7ce9bcd8de4f56e4a5d2c19edf601e17909e81684b2fd46dae13e0a0c5332f
z698b9c6085acc491804967ae630a76de3375cb99572f7b2a25400334aa58a5073e74fa3e0b0199
z346a353fbd0b53632a1b41be1b260dd48aedee44d77e7418d729e126abd9538e57fa1d54bc7d18
z0b322a8cdefaef941cdb967bde958e568d609aa1fc0d5d69eee6cf1ae365112f2fd028b2d719d5
z08fff510557319a7135104222d0c6d49db6eec4d4a4482cd6d71c4f19aecc98120f5ceb805255c
z225310c0470c67d367fd3330561568cd26363e0cdd19fa38e9260be6f0350d95d9642e20c7879c
z55f0247fb5b5621571b6b8aec072955045e4da764ab8cd6b24e963f4659222cdd094607245b9c4
z8c058fddc66db3a9d72848c5ef4eeecb7cc0820498e2174d0b7c66623f1cd5be63713f1c850a06
z004bdaf58ee71dc916670e657e4107d1258654b51ceeb50789ef8473b0cac4a2944891d80f696c
z3fa79b7e54927d2ad7857166268367a974c0889bf354b86c077353e7bd80c79d99cc74e2dc28f2
zbc7ce35d5a3bf4656e5472241ba16b7c358eb3eaf6cffd10c5c731f977c0a60cac49b79e8c8fc8
z80ac1dc8183ef01387b90732d2741f090ffb0b73365cfc6d0be89e0e3c2a5d7e046391a774d083
zab13471082359410463a10610cf2a0dc78974c043d1f44800f9ce7fc61dbb8b52a5546feaa5811
z045d20da00bd9b8b2d3f3c0b07b67d76f389495f59978ce45ff64f1fb3e5e9f49f357989fab159
zcb8d27c3c05a230037e0e02db40d16025bba96c485edfd72cbe87cee4cb5d05e6e0644e0a80db1
z79a3e9b2464e7e1320268f500dc17a0e9bfdba169d4915d4246ec8cb4c1dd6b2f5ddb457440577
z65c4ec1655c51bd46ca646a4d271d654619abd5894833b7e0d955e35b8d5ace28455df3b4e5dbc
z2bac04986368d455861725fe4f9b6e6eb9df3c88e2af5bbd7c5aa39d8d458f8abac438e880320c
z386ae495901a51e90fa96be12d225b7dd49b98716348c289280567369b0991b0dbf1d819d7ee48
z4be41641e5c78659959f2660ee7fa0167b985add0344f453d8d4e3125f68cb2c6ef03502902177
z913b43eb7eb03e7ab2f127002fde2171e1c33c94b4fd39aa1db0094432f8f3cc6fbaf30b7b3b89
z82c68d7908eaef56db6b832aacfd40594fda9ac9f8c58c454dfb66afc91a705e237bf3d12eae19
z864f6148256587231524ea667bd8ea6591df5d636c7fd49f951f60e6ba3b5e8301ca54bb61301a
z536ad8260cd7404582824b6832921fa06aff9597132bde86e6f595213b201d2451fa5e3a6c0642
z13ce17308b43a2edb7469f38b91fd69710e34e4d90f8679ad674991e619bb6a609ed34c9b3547b
z8d8ea5e2f1ae3df614ce7a8085b391288746b3cd0954bd1aa2f5b8f73aa30c186d14c149a326d0
zc4b78dc737a6d60e28657eb87eae3cb701e97ed31b14822cb479636e38466baa01c12c89e5ec2a
z04591399c3e9fa86685e82810991485b98a7b010accc99cc8e358685ee45dc8635e97ed8f410cf
ze51d94e7c22589dbd332d23bfc9aeb202ae2a349bd88684b25dd4a0388730ee46b8b9ab881594e
z11671fb9a009871b5d09680dfc08bd75908f24ad5df673e4c5fb09ce844737b4a00c2dd58b1560
z958e352e2147dbe0cf6cb1cb3f0227f3965b1976b39a2bcf79db21c27f17c4766bb5236f7cd2c8
ze2979b390e6367e583c2bd3946fd4c67bb730808832ac44a40f68a6f2a2f29655e8f3204f46a4f
z05b8341a9f898f710599fa0eb3023ca5eabbfae9c4fe1212b1d3ab516289bfcd34d41d64dd4401
z3801a04e66709efbea7c6eb6ba899bc5c989d61a8176774c8e85f14662573c38c27a5df375caf1
z3c51a37b56afabea9d360bafe29bbc257ad884150a31b1cf13dd6cf7e7bed3eed0266815ebc831
z6f4c80e9ddb4ef828742b4ff165c784de5147aa545275699326810e50e096ff739b82210197e7d
zeedc82debf56fe7528927a8a8cc62fff99abc8459a9864a725c7a4f11f8984b6386d65de1c5cc0
z7b368cf20c0fb5f0382811da1b715aba3b346b7d918b9d6b4c35413c950a716acdb5f7b77d8a24
z14f9189f5c36e1b6fca668994b76de20d7fcf9fbf556ad39535d6c27dd3d944c00e559d34e23b3
z0f6f093088c2be32049d74f1e9529196d0fbb59bf9e3283c0508c90dad70f50fab77950cc9cfdd
z57d499123ca4199bf1d88fc618672d2e76d7c75f85e23cd9a535c190fe492cf76e3fba41217974
z3cadef94f1269888d4210b6561db14eca0b0cad9cde602965223ec607b760f2bddf5c7eb691a33
zb265619d4c7daeff77bd5eda8b134d1f9cfd542c02de9d2c9f013b81dcff7fb31fba2a4bb1105e
z384d613313cb640f0724a5bd903faa89426371a8b41584e6bc8af25538112cf2ff4fe68daa00f1
z17b430ee28d643f03f7981aca72bf312ff9bccd3b9e774e3c9bfc9504eecee452804481b056e2d
z466d842f5e89e9e4172a2aaacda3324a7392065276df8fc7c0b05b9dd045db9693017ea26c636f
z2d3cafc247c8ead50a67538346ef261b91a6452104c4707949ae979e084aedcaa233c4cce06bd7
z62c50c7d559c3ffd83fcfbfbf71ce4fc594dba0b82df3ade8515372762ea89723f5e5f691dba1a
z058faffd8e0936241f8a25c2970cd5ed5156785419faddae5c8e6607db4833d6c7ab9907664958
z9b0e1b3c085cda5df328a8adfb674d8fef9f14f6fa24f7c663d3bf35070e08af6284626724c8df
z7351c436b37ec05966882735c96f56a5ac3913e051a805b078da950a50478ce5529de51b6af1c8
z00fd19621396777b9ca4e509954e5b174fe8d663d4b8cea2b96d896a8f378530479d58112eb063
z646419aea00033fc6b332e29554bbb67a14d095f85ea9822cfff2964128cf0a1c3c1fbee58af60
zf5f524b653d38ea66193e35a06e809a044cf0ddfa165773a66fcc7e70b8a5e2ab392ef1a2f1a78
z010b8a3b468b0c78fb1151cf4b318064e107220e5b739eb9a44866eed2df9cc706e9448d7ac724
zf28e01d2bc77132e790ea17401545ac1d1e923ad4ff89064d1c9757d8f6cfd1a5860bbded1d666
zb67c6bb08e7ec2efb9ed9c6c40d96866ba8e4590be5f643aec16b4d948e693e45e115599a56af4
zc64332a7dbc52f9b479a6f1a8c4b119629a82ff8395354fe1f9fd8a239d1a92df7e8a0f721a122
zfa24829d1a25bae76c7182c86732192914fec9b49fa5fc85ebee4b74af09e60404bb553da95174
zd579388d594bf9314ad25bdb493dd7c17fc661441c44cac3a86bdac8840c058c6653f21fb283d8
z883d9ef7a574758e3bf141f6293cf0afbb5bb0d1937bd9677e4d266f83d71f672a795a873264d3
zb194b5bae8b6b78225d1b531a80a740de568b100434e1a9362733478f37b3d962c296e132ff56e
z330dbcad5ba8e6c93873e1d1845010368277337fd16e1e0be3d86831a908f9588e9559242271e7
zbf4ee9177660534d9cac9262f623751e27e4e4ec73bfb0f1b985d6e623d0822ab30e1f17375e24
z68d4e9ad48430b35f9904c1cda0ee2fc0cbe44cedea6f92144c0c9037b1b7f89db42c8120bc997
zfc5387ed425fbf46bacdba6c5f4991215322e72133254c56529393393fea9d706640133e1504ff
z1e6c534f8eeb558c259787ef7f8861b21b67c345a8488d2ea41c894d1d4aefcbd17b960b4ea072
zc86fac2477f3a8f2f82eb70f5734200253195f10ab1074925acb642db5d3fe1c99c57b96e916d2
zd55309620aee239bfa037afa1f7ce53e49eb464145bc308a8261d8c0c0c04ce3c8eb15ca3e7570
z9bf8723bc6c751910e3d33f469794f35dc8db0fd249bce19d7d107e6841e903514ffc06dbffcc4
z1d7433742fe550ec4438a824c54744ce861809ae7700a624d130573ce4a0b66b2593cd1817c44a
z9af52308266179e5f3738a1e717f006d2636b697b026c87a06038cc30b97a692a953f75d0bd287
zbea32721d33c44f8788a1d3be4c0ec2a4ccadf92c9046bf6f79b98cb83f355e694a77d4c5b97fa
zd30fcb13df7dc6fbb6d2e1a8ca8a03f8bf808b280f54f1f89649bc1ab559e7bc94c015f21513c9
zb626202af477ecd8569677b5fc4c228ff1be502a5c87a727f9cb7177109f286ed1c623f5cfb0e0
z77549984b4e8c3dea75cfda5c1332daa11e65695794c19c071caae7c58c78c9e3c120647e8997d
z022dda291a4fdb763d160fabef1d02731a0732f6a4002735d5cb378f2dfc3d614534b760759db3
z6491d92fef6a5a17fa3d8ec03d1b6b143bde04e9c9af7a7572ef19df0b090fa260949e141160ce
z2fe423150461aa912d443f9cb69965c7496e18fa24173d693b472bb863f8887b010efbd9020817
z5ba3e67b0883cbc41d68f7ab393f7db2449d2c7d09fc7a35b67f6322b165f13f918d0c1cac5bbe
z0c16b0d4c3cff45b1665db6f92cd67866fbe27f1a1b13033569aa18303ab2126dadab17cd0bc12
z65d837bf64bbba7c87931fae5123ff78ef413ecf95409e29a445cdb256d10ebd9f2d089ff0a533
z2e47a98283a9c43e4d9e10797fad0d5ad2c00245d6a521dd60d8a5aae657fefc31dae242f2a132
z473636eac23c11ac27ab1b300e47b4763f1b094c4171a64bdbd76d56f2dd6da7733b486df33b8a
z9dec3f8eaee0282b47fe95efcc109acd2b1538223c9374d45141b65b6f317e490f912afc2debeb
zd67fc6410f1b242c37d645486fe1bda9284ab84cee13c17e77655975c382640261f9b4102223a8
z38a1a1db35df40db13f8d7adc67f3f835348b5d0a5e594bcee7a66043abdd99e92dff16d014fda
z95e0df64c1271bc1f71fcd6ffd0a47fae5e0185972713e53e469234623473f58a6e63257cf947c
z0c8d3eaee23e8b54328bf56fa97a9d5d166775f883cde42dd14b9d46bf18ad93c94a9acc5cce55
zb06367a070fdcdee56a14b0aaa97cd0df4c73e0630f8039d98093a705a1f18b1823a6da094a66c
z7b0d1aa0baf361c9474311973bd8a246309271d4505e7d323db1200ebf79dd3329ac28867b224c
zfe85502c860fbe6e0bbd259f7695137672899f48a4212f46de4a5312e2c9fdeadff16282e4eb31
z9221663225214515e725ca28f29dfd7b69f0e3ee15551316e26f49f1ec8c359f13d8f0ac86ae86
z726b8566e3ff2c5581ba50c79059545caa1d9aeb6b41061835519e0d1dbc59a837596a31c7047c
zf7561b899b96946e3334e1de53fbeec18036ef5a1a8a568221abf8755dad0af2b94601c5c7a17e
zc2b5abd4a49933a2270bac89930638910ef408805bd433ec47ef2ac9437636aa914162c4dc3da4
z878770fd882459ed6cd620f9e62123ff9fbf4b5a88054d55d9c3645172853baa6ad341dab61482
ze33f67c466194303c3b80a0528208174ab74324b1529abc87c94e22d43d0c57e8c2542b5758ad4
z4346d3a443f8eaf83fd7676de0cab66d07af9fa1ed111676272f84daf51170510ddef30a4c32e7
zc355966d07fe374673157c67cdf8ac27e970cb144462754c44c7cd97e79a8788354d0cc06ad4d6
zcaed27b70e03f048154ce538d2e88e0f559115b7d50b6712271964abf6c593625091c9f043f584
z5d5bc6b16dce8d9b6e3278b8ec5c7624e5aeb801fe1a277b1013c274aa2ed417c5d139019b39eb
z650a6c2759b4478840cd4832e24a7b34e2bfface1a160b47716b7449bf1517d7e97fa34b1f89a7
zfe1a5f2ee6137b5ee5f13288f5c781999c26080490d44c34bb6f50cd0341070836c056af5f6cf6
zb987e1adbb200dc6ad30106de9584c2257025baeaf0854b6b9f1a4354832fe28ea9aedb287140b
zb9735483e2cdb8ecaedd0e04566decb875decfd7e9ff9893e0bc60a60033476921784f803903f1
z1197d3d1340fdccc7d77b255e0ed193290e18b3b64b9e581b7f65ca18e061756ccf8196a109bf9
z699a2f4e677a6d08d9f37888a258be0720978f1f45d5e6a7898c241344fdf0f674622f8213fbdf
za710bdbdaffcb538ae1262f1e7c0600f75d486d89183bb34fa383978c018b037f6f304174a192f
ze1036f07d178d013df0ae360acb09f7a626e18909cf642f092d181e9346d8107776ba35e98c385
z8f84063cbed4e23c48508ef33cc2ec54950ac09ce825134f017eee2a4a049cdf8b910071b6c2dd
zf2a2e2fb88f5d16ed966bb122a6bd6c14d76be6755ea79336eca0fd22bd633995e6a567f28f52d
z6593835aaceed1024c8de443ff88540db91ba818a1ab980e6c4d0d62379509ef37b1f7ff23ebde
z4af6c956c385b45d8966cb23696fe26052d80224154c600908e6f8db975f318a624cc09a06d2d2
zcc1c5b93598a568395d3fa526fb00266ce8c358122db317d5ad8f77f7ab85b31dedc9d7cd83fd1
z909a445bdc96c55a4351665824e5b161fef708c9df188ff7845ee322790743d7970a1241878144
z2c3c6a7d5f21e51ff9990b33b1d1a0748c9691a615709097ad351bee51c5e7c6b80d221da54bcf
z9f91fa3904acc36209537ac5e6d4847affbf4707d625a78be38a884cfda689225b15ec5ac4dd66
z1bf07d6534e4a59690c444cd932a0a55d419b2059bb22a8be02288d01b9f142f747f354800769c
ze04ae0c53deaa158783b2c4997f04983dce0200763071ff4dcd32788e75c029ba2a1b777553db7
zef0fefcbc606c360a2067e975c4bd9f3882e3997edad21e3d8b37dd8fc783a90f613d481e6e1fc
z9b917e738cc7b7c3afc3759ed6c63551993886bc00a482b1f79babac434d156b42510987add0d5
z17dbebbac841dc58ca5a1267267e8e721ba2e58ff9bdba48781bbfd027b54c039045faa4010377
z982b128905625970d14bf6f7cd7267029773aea6f6a03d6462bf791d3c9a7a2a560350104e850e
ze4e696485d80faefd52ac1a1810e8bf8ab99ec30410187ffc4653996f2e61a5b3a85fd2905964e
zf6a5c9bd749d48a62fec03ae96b649211bac0aaa646dc7d376a768bb9b06dfda37ef62852ef89b
z500f5706f6cb08a82a2d04a24e70df4b552107c2fce58d647b355367d4f0d893c5a4b890652b70
z6a2d1c9fd02f39eefb2bd660fef0055df4a93cde54b3ca3bdaebde432bedf69514f2264d8fef59
z7b73a3daa1730c80e89bdf1b765b215781b9fb7fc311b4b1196ba93e6e7172907b024baf67c775
z4e7c50a3d3b6e843a82d99c9212de1bfc8c1104f80e80ad75bece275119ac6dafb8f89de622ca3
zfb23d15d52f1b2ef08f06417728bff3c8a74981c083240befb62110db88896df928bff6e1160b7
z72d199c9bbb95016c7220fdb2696207159cd0b6a1f3bbba20a0e5f324edf18bc12402ca0731ed2
zc140fbefb6c15106268e7a06e84aec7eafae60070460b5f1513cdff22fc2fcebca16f965fc0613
zc02e4f4693fb0a3957146e8e1a07ab0c6edc00099abc56ead884ea0333dc549a7076ebb6a5fd9a
zf67501a56be046b8f9ce794e04389278837a309f80ea20655d4bb2df4d63f05f62fe242b7da140
z3b5d322dc90b46072ee5d3345d65b765f5186f06074ea76def7b955be6044fea30d7ff444656c6
z2c739505f33fb3ac828e199eb7ff1c5188aa9254dd808d26aefcfde035ed07a58e702127711f76
z6acf47923d787d66ec89af205b13947c9463e39e50810246c21c210eb68886ed745a991bf3e135
ze15c3fc8d5a0b8169f7fc3bb029325019d9a53a5273267c6b377b04dd85bdccf2f69830b3154e5
z817c5a3223ac4e020365467a07bd17ebd16e827f5c427774422d99998ce6df96d5222a0ad7b802
z4986caf0d636fde3d3740ec5be992b029ed806069d92ca4089730c016193f523dcab0f18a31390
z4cc2549e6ee174bca0fc34ae04a1af5289781396b00d1ba0ac8ecb3ef336069b3d69ed99ad995a
z74d471c6d9f09d971b4f5cc96258f0e4b3831972e5a6bd16baa4887dfbed84a0254eb676359658
z7fb2654a34513013eca535f5b9f828c6a15798c87a8b9b5be6c4647099beb953ed6096972de5a6
z9b9a499564f01bc17a5470729fdbcf258ccb796e18bba9678ae7bad4f151a2e6db64a99830c2c5
z1db0653e5b49f32846e015c620985e3ca2d74c8d0e0452848953805ad517524ace7ec4c86ec117
zc38a7b39606a430c8905c0f5e27cc210c9f436bfb3073556e17c5689d303b22d63b312a990bd86
z8a9c51a7796819edc8f2aa891faca1edc8b82f9bfba8ec7070ac67bd2ff3349d05b81f311d83de
zba7a1c9427f01083806540c4f3625477d36405b239b373349cc28032884220af5c78a5f0f796d0
z96e2e7bcf7c252632320b3502d97c651cff9ee3fcefcc24365e3cb68a0734faba926fc47e9e695
z41bcc922406c640240e35d7ee4085b9512c5ce479e36ebe594286fb74307d5e1324cef4f9df324
z969c00221039c94125a34ad49212de1b3005201cdd58baf5d20a767250b0155ae08b210a9d6959
zf86daee05d31ec857823d128f5ea5fe6b38c8dcac5047b96e9b00c953a305863d139f6577c4299
z4ff9595194d2e617a4f2a679251743cfc8e2bff419969bb17a01fa3118a7972b9b4897243c07ad
ze95af50869134f5fa7ae43f7e07c5d5ade10f53bf704ca40eaa919a7464f88c9c1ab4b0968ee50
ze610185a8248a9cb4a1f69507b75b8041cc67c8e292b2b795f1d7e375bf673832da8ef7ec6e6bc
ze4f56396c365d27ce9677c63b552ea945811be118e7da202403b693e95a394826c7b49a6ef1853
z21cd9fba4addb49059dc2ca0542ab06cb89f3a9d784ef69eff087836c5539b76821a5e6c9b5f8a
z7ed27436ce67200d19aa4ec9702389f3bf9d2c0685e32a21744e014072b04bd01970555063b283
z3a12b572c29e25ee1fc33f78758c658ac5ca74a206bb9b5bfe6ffeaa0694e1b3665e441cd1f596
z0849a2806dde981f737244a94b5c098863b8f13377d1526ea90fc236e843223d9cd84cfa648332
zac8d8fedc03b46f5a30905b6ffe818a2c1c51e4a49e26f1b03860b608e6dfb6007f99b17ab85c3
z53f301fa32d706960ae67639187062b2528e7496c66ca05002a0bf0415de737e0de2b169e4ecbf
z7afe2c4cd46f229e6c751d020f12da27c101254a66e2fc37ae77cbba1d487625803417757eb376
z9d6735fa36751ea126e29ec2bf7ac1ea4f5a19a3458fe8164831f4281079775cf1076639470dc8
z2f996e5bb0f296a074b1cb0761b360cd0b15c98eaa661d056538f1445cf1058ea0a7bf1dbda85a
z49af75fb6eec486eba9e7a6b93e1fe15aab36602116f9bc4fcb39177ada8a17e8c8689b77fc210
z03ae4e1654f8f22a1c373998bcf382cbc425ed052ef71dc761efcf1eb5431af85cbf0a88180c5d
zae37cc730e5eb3cbfc702cbc5e5b8f444244872709b659e795aabb22ba2511d410f9d3ddf016e5
z693e4ab55b64f54cd4a2e7ede1756994c023353e1d6f780e0fbefaa97518fa4a20418e92d3dc4c
zf08bb2f9cf750f5bc93a000ec1b39b14cac74bccb2d9f1cb3cb866a12e1fcef34018c2f762f702
z1f28284d7060d271b611f3993354d6351dc90c4ad3491e49c2ca797fb262ffb351c5402b9649cc
za45ee203c78b86de28296ad77dc90dbec678e7cf5a8176f9cbd3c50688acc25f57d97380b5568c
z4d2e796cbb4ba236160ecb4d5e5f958bdc11ef5716a598fd66b541b89b51e0ad6e10980cba4ce7
z2dacd7ed45c8bc91127cff5294d696ec740e514a98831ab0a813637630581ac2be76d795f47904
zcfd344d349528fcc2bf9621b47f79343fe96ce76a8a2fa80c033f68566024ed81406a61cf6526d
zfcf6b85523926daf5402f13ea108b770e8f827fd3d15f9ed590a58b6c9e7e4af6abe0ea2e8fb29
z91c901a07863a94abcd1f9ea3a9708fd903e5ac191b9d4d10580fa984577c257faf6ffba16cbc1
z6f4bf53dd27a785a44a0b5e71c1df920faab40c5e427ba6788be81a0d3f73cd9f6cf92af7de473
zd3763d8e06d5febf8ac3b5a81e7c1d2410941cda7a27a969a5f12f0954db2905a74c2f2d5e9c24
z93bcc0c6e20fbbbef783c921f3d68633ba8886e48d9906a139c55bfe6e9a658c6107132a440de8
zc22fcb9aea0f3cbebb4ec13ada8d6acd4d4f6788bbd7fb2351300d4829e14555e44e356314ff1e
zddf218aea8fe00b2a54a1e3d59566a350761eb8fe53682cca3eba5b223ba75e67692cc1fa699d7
zc1d5ee0b08bc8fd57f5f0b5e27ea85c7f19ceb1edbbd328b5634c3a7853c84a2ee353d64ea9309
zdf7447843cf544e38e5919a593b993814325cf8ab3a2de3fdba6b9ca6041581e94adaa9b6e81f8
z0597f1510fa3b785d3116b5b1eeb5b9ae052fba57e14954aa568c35dc46e9c1338b3b6a4497f1f
z094e4046dc9771f22013c7cf65d557f09f4613ad1fb4973689d2c9aba815bd59c07b2c68201a9a
z9fd4988408f62e07ce3fb1ccbc4fa11472cf967f0aa9264c58d0485eae5b9db54077b54b5ef34b
zaa756e8161c93b5a7b295160031bed6a0d5ac3e2d12d7ce782ee64566b3aa9ee418cbf9b57f6e0
zd004ee254cd6e4d3b7710ecb2bca4eaf6411f8c489a1a5383b45db862dd67b98be80613e478140
z6851116b9fc044e724de1954b7ba5a84e44d695eaaad538f4e0e726c6a0b177d1f858cfb139114
zf5caa7d4c41714bed9bce4aa78273d88e2ad7b4b040d3106fa6df54d9288be32dbe82f95001338
z15117e06a291f4af874a22e1e75cb87d32ab9a107b767201ceb581a7fc258d6f6ae186f7f01b0a
z38ca222daca189f36de5babbe4139650e8443b9702835990cdb2a9bda4cb2eed724d41f026890b
z3ba5408866db098f6abd501c0e2791c2b80e7a74eb1819e44e777980ab546fcb82ab754cd4166f
z3cd6c760afaff5db9e170ee51e8e1497767beac465f70e1455ed0aeb047aa9bd59dfe924cb87cb
z62b794a3ec437304be66869546dc704b4c599cb36a3434c59c1db73f8217b899c2eb676f4bcbde
z8fc6aeb5119f0867475ac2248f23c4d897135e16428a76322edca909dfcc51b419aea6c490755f
zfa3dd1661791c94343ae95a91aee746846a3727fb44c7406428df673422dd1047bf09f9a0a4fb3
z496cb05f6aa6c944f7152881530c62a2f333f7a49c3bce2c14d7d6d8b02d9e3532e54ca9a12f8d
z4bc21d78d7d434b64cfb732f855dc0d7552ddde3e28759521da4969cc2e453c20b64b29c340793
zb5778fb61a54ea62c1ead0d8715945b5e074ac2227215d1091c7bb33e8f2c2c1b96e8cc6b2c514
z2b1b5c3ef1c9d0b9e4505b219dff9f8645499e192ed4a5241b4dd6ff5628336621d06352b86424
zbf4fe5dbc37d73069135045611ced0611502f250d72ec73582964a78bd206085b088b514d80b02
z191ea0a82acb3acf6c309b0ca07ee27ed078456587b1bb8340447bf82d832a4bf285877e916ae4
zf1a9d57c75d47b1a06815b5342df09cb04af835d4f996211de43c9155f978baafb68abc0a38f34
z91a85187a30b0554b624464d6af2dcf06d892cf5ec8663eeb5a2b28c405bf6d19ea5deb4d1f7de
z0b5f696fffcc7874103716d318afbdc7239356edf9562e8e144b275f9ba915f5a4ae2909b6967f
zfcde045428e411b6de4e45ced322c90b97cb6b3beb05e9bdb6ebb66d4e2d3857d09a548024564b
zf6f8ee5348f0aa8e4c36bd1bfc083c96d18466cf146f563399c909854307aa0f9d27da83a3895f
z7d8a2197daae1f49b89cab2acb16a106ec73af7549227c5ec0e78dc87ae91c27a99dfab765f4c3
z8654a8327f8602e0ca017409424e990257928b2264ea6e23af40de2e7637ba0e102c2f0f8bdb17
z1dfb2580a9bf07c293832942a71d973d57736f0200e42b9f13dcf3bc2b0ab02d93f698dea0fe93
z799a28d9f6f0a3a1284694ce8afdea26cfcfa60631bc296aa40a1c9ed7c7d683d3e8fa9aedb136
ze4feffb06a55a03536f42283566891d9d1f4993fa14da5c9f76278cddc2e95270a44a6856f3958
zbfe5619a71ae2e796055e02e6b44cbab8f3ad439a0c89c466d038a06ebafe0ac10c5e513ed77ce
zd1acaa6d87df320fdf53ffdd4bfe4897094140fdb979446682dd328a0b512355c3dab320fbf005
z883bd98d81b7e75fd493db0f7ca6d10adcb8d0b2069d3285a98f92f8e699284ba46d021bb6d278
z2995bf0fca81969ca1c32686c473895e92aa5fc2c14f7e7b30b49d3adc44ca772009465a31ae06
z8316ea82bb27ca9cd872589e6a44b1f0fe763864b3c40c427bd703d301220b9587f05fbedd5d65
z63c4bf3377ad5ea861a6132655d013da38ec648b3602cf0ce1dd50288c3c3684f3b26fa279e390
z3adc633b50133e0935f89b7f6272c3e3354ec73e99ae8132ac8e703fd9686ec409f65b76551afb
zdd063a0be32110b4a798c42a1147ff42b9b5fd18e7443d2c5b8a6f8353d373f0c7a9cf8c05c762
z32da57e518148fd7031f4cdd4a981a2f1eb9f46f2d90a238909e770c34897c8ed856325310ec9f
z30bd23a03f73a5821188cfce76f4f7d21dea81aeda39d9877fe453eafca24ed0a25a7892b47325
z08aa455ee81fe0673ca145b3bc1977557c4f39ac166fc103c8366704fb388c25a153f7549195bc
z67e71bd7fedbb6c291921327d71cc82a29ca61debb62a2214b46f084ec5321c94fa5880a389a97
z458767b41a86d28d05b31ce1b2c1f3de77edc6c6f5c1f69142230cfbec2ef7f265a77fd95ca6ef
ze0cd1c1c55ab906d665153a1a601d29f8aa3951c625c9cb1284d76077fe375f833fb1d3f1ef7a9
z1202316f1253130b10a085f8270824a118634e54f53301828b6fb03de5a6a7cc412be63a2f589c
zb2b0d735941397369407dc18034c92420ce37f8c6f72c0ed0e6f731c2ffeb83e29ba3da877cd0c
zbdf10f84173bb6dc5fe6a8e2fe24af2ca355d5069367ede50c1caaed6cd60926511a592681d44c
z945d7b7bae172d09a5a5dc32f771b935662ffcc8b4ba764122c3b451cc5815b8e3c1c2c08aa149
z528d7b7de8313345475b3f999fbab33eb245f692530752831a1db0c650b53b1d65b296e2a5c6b7
zd8248808abece5119c97d6aaee7cfd71ab27f707e236254a5e9f54d9e4c7ada65c2a7d936081c9
ze095e2d870b0a977c36d992cdccef0e03bb2d672ad45f70037bbab50556e5cf24c816378b3dbca
z347180521d05f08c5a606679d2a03e42455312c775e489ee8fe2f7e5caffb17ba94d7ff88e24a6
z8d44139310ecfed8ff4abac31eed0484c9edb8cefab7ca3aeba18edc188745fb5668c99f1d9d4b
zc0881895a885e4e97c1f7233b688c83de52220d2b036f743653d35f15bd075b15c9e743a0701c1
zfff2d34d8573ff18f11da64d7d26b0d61ecef2bc8dc8e7ea24dfc44ce5c0757ad5b1473b8451b7
z6ce9cfb380a9420fad57d3d85f499e70f80135b866b021e5f2b443919c627c3f8f462bdf8d2693
z145a8d2046ba0fe4248db529147693ec2a6f38327909cbd3f137eff37871eea3c2a2ea63292b9f
zf89fbcb53364995176971077fa85d2d4ccdbdc5a014d06183346aa50cdb75537329f5918a69012
zbeb53a750e99ad0792ef7ff9444916a2799e6e4b18f69007d849563d09d5ee489ad70b062c62d9
z5a363b6f342a021eb746fa70cce063f6a12510d58e904e83967673335501bf5cb3c98f2e8f2e52
z73846efa752759a821eaf1e04a4265e59ced0d60dc0203bb4aa44a07c4df329f9bbb22830cd35a
z04ccac07a8461b2a84d5ae7e1ebfe96459034a82fc7abf038724c7bfaea113c3e517b5f87efae8
z4302a53df30bba21e5fc8ca4a94e6b59a4456d71028c07efcc63f641dddfeabbfffe343ac5f3bf
zcc332041041125587b60153779c3be760a1a7886b43f47837d7f2585eec0d64be358cafcbf4f06
z22e919d421e45348e094f6ccb6fb3a1421d29f083079d548560e94f0e3298a30d751cadd2c2c53
z66588298eaa96dcb237dc9f6e6e03c9371200555de5f52bc88c0f920f5a7b781c5074dd402db9d
z871185d50fdc454ec667530790f175a9d132dec94814762c0c3254abb4961f98731afea138b2c2
z7bdcc368e118871f1a325c8bd225e3e12dc8512ad775a64880590da51e3afe5b34a665ee0f509f
zaa1d1b54c2fc4d8a0c9887be797b777595b6cd0b3908f03dd58332717d092f958288695bcaec85
z029a83bf22f48416ff63d8cd7b9f533a03dca0d643a77797bef9586aea1cf79b61da88b76cd37c
z4d2279000dfea4ef62ba179a0eec3b5b9557177f877f1ecce028e0addb2dd2db11ee3b5b23f086
z471e437fd49c488f7f8e59f5332ec3b9e12ffbf8579f7d58e641246450a844140fbdc754bf776b
z2f6f3fce5e6dd4bdea7afd3b5af99af0d88582f4cd28aa1b53048dbd1b507f5de1b97c4b733632
z17e2b19a5d9a22fc1b3d0bb9fb4f21feaf3a63e5b3b0b5b99a63c7b712f34c0cc658c812cc688d
z8a6df58a7133a85e99dffef740dfd41a6f19d7480b67b1a3da1962e4a5f314e998fa60b5512963
z4bb0288b3822645ba90c7e2d6d7e395b8571fb73387c01cb98b68e76161303c62d799146405d66
z8be0bf414acff303c1f2b5b3c7d4ea33de20aa687d0ab460033b8d486161fb7bc8bdf375da528a
z51f037e6df2c7b85ed7f2610af650efbc461c35c94a379c7f8e9fa507166a8f9db877ddf736706
zfb69efc3be0f8a246a95fabb5c1c50e1ecec3922c9ad35a6d03e341af47fc2d4a929526acdeb12
z02f0b3b0439b9d204ec74f7314ba1fa100068ccae4945e4b083db7d52dc6e551fb8ff187f647fb
za1ba6608d8ef64cca3ab31412209490e7990b83e3cdc02d57d40d56a294e6f83a1fdf7a75b4097
zdf9889ddab6a82c2f49b79aa5a7c33ac52b693a6541b68baf261414903081c9693bc63f0fc1c6b
z4f2e125fdd78b5fc79a5085d1e440cc718535395b520954d81969b910ef37c5511a88344561b9c
z264b9a3acdada4053e05ae5e628cd53a5721d52a9e1b398029f481969d7c7661e4d02f71103d94
zda21640ca10630255a576f5cbafb5928981a82df3531216bc9939e2d0e10f0e751a2bb1fe1fdc9
z4387f6df9417e8cdb4fdd142befc66178f00b90a50a0d35162b087610f1e6fa6499577e04b6859
zd367c66cc5b9a37e240849651aa52a3955756d18093ccbc5e5bc06b073165ae7a644f5397ff39c
z49a29ed1c29c0a9f03e788acb06de5e2118764eb4fdafa5a4d8b6928174c0a5fdfc7ec4fa3a940
zd7573af20718e5a24e714d95bfdf96bf2aae6190dbcc589fa8243761c5faee4efedbd7fd8a5ace
z6dabb19af651a3857b247e62f5b0ea4dd69311866cd902de01ae63a5cccb0ea7aeb564827c1648
zceb4d5473e2486445694e027cfb31fbf3e8007a45632e91d3d96c40aa02fad9336dae32126cfca
zbe44dd36b89a21d025e18365ada278e532d0fdaae174d75df97de51fe73918f94e5e9513ebc53f
z5461a7de87d46e929d244dae70ab6c1b8087e95164425f47ba5472c927f6252a351569830ece00
z4ebc29cdf85bd97858fd7e4ffb47fa0e95614e6d66bab0001773b8464da62e375024ebf14f91cf
zcf149379c4d9fb5f9817e3893fd43330c9ab30b9e89d70b086c115687526073fb9b622d7129b56
z8dbde5e500455ba9672d96a9a286d27cd5502745fb59a9113b4f5d79834ca4e48c2e65cc01e641
zb5e767813b3f8886f548b220e2796dd05a64877eaeb49a4d823b2721cb57e7e25fa8ac39c34f70
za33e871fc8deee358439751eca2deec4b1519db890f9e7d6bfe5350a1a5f9bf1b0405c0f7222cb
zaba45cfbbadee38d3f4fcbd8e8f5b95847b20333ab8a00d4ec0628900c155f7854f04d7f22b540
z3ef43645c5389a5bf62fb20ec307267bf8aff045c09e977a9159287aa6a2bf727661983dc542ca
z6f32f9e5d5478f5096c2e238e103b23e65a2a3544fb6c4e93b568ee52c013e8434b1d7b2c8f9e8
za4b66f8767b46655dbc33fa59029074b5b2d0280b3cec4ad517ff77a55b2c31157305c118f8200
z684be3522eba81e5179f90410ab2a8c1213eab745117d417ac4cd92c6f50a84ce8b7886cb86675
ze2d910f901a2d24dd5d6e695b79f73033d3e06900430c7e36fe9834a628c25e87935dd0842ffd8
z4f3b9260b438fd27aa8b297f89e0c2b082ba94ad6cef1779dea8e1a70b8608f4152e7ceb21a6cb
zdf6970281cf1aa4cc3e0d9517da2820b73914feb8c828a109a7c2b1ae73a3ab220abcb52e381ac
z139a92e524bd70a1aef78f9d23369021e4b42f10c24adab7d227f5500eeca9f8dd7c671da3f235
zb921bce3f5df1ff13f979cee79fd598f63653b13a6cfca818078293cddbc48241807fd7a1ea5f8
z6f0b991106d88707091047330c924c3c472d756e18e0fb70783f30c8b84b30ebd90754463c19b6
z9196dceacaeb8cd972796b6229bd39f518c5d754b2ca288d7d872d389caabaaf7eff6b2c45001d
z5f96c50b80a76a64fed5f1012bc1860710bb4ccce6749ccaa2eee318369b6c7616d95c36fad678
z54a53eb515c7595e3ebad00f3fcfe6ee35eeab8b0534fb3480501d859e5f199ffb0433319e6387
z760b02d2364a37656e4dc0fd3cc73f0359c805f300759eadf6dccac652401f0133b77cab1e6999
zefedb4714e6f31c9eecc2e05366fe3490f5b842d4aad05d58906fcfaaf5238308a7e21b1193cc3
zb6b2d1d697e4f26f8bb6e14c6d94f91a0d415d562879af57404631b06bfdfe6e7b7fa58d150f11
z702e025c1dd83b5c74f7e95cffc72a8a39a8fd886c44b37eea3c737017fa1b2a1ddf85a874975a
z102994df561743426bbe559a1f3d8bd6a99c7f9979c3ee914445bee42bb4244bcd87f5f37881d8
z89dc9b929fb4016ec80a2fd5d8ecaa88034d89fb67715803427b4c7f39e1e918e34aeafcc2f71e
z323bdd092dc59e10c2f6e0356d118bfcf1d2eac4cf6073ed0f4e4799d00ba4f4cc286fd021d9cb
z1d2660715b67cd70c7f8757e0f0cae944f0c245b274364a469b6b30641c645fde3d5375e657682
zf6c1af9bac029f445ef20fcc6e16d2de451ff99c29c555fee2605e039f75d7cf44789bb33c7f7a
zc9b0b7fa815852a4eaaf2bbe912e00b6cd651517a428ef1c983785006e30c26c776af25069c47e
z54e067aaa8519be04d1e07604979295654488eb181e56db4d6b04fcdcbae5986d5a38be87c725b
za2b121d74d4a45df68a6096ab5cbf913e9ebe994042115dcfbca8afc84f762ec1f0135dc93ae38
z87e9964a31f4ad83aa07a0ff2618b06b7a60f7e00da25cb972f55edb2f6ec1d15a53b689fc6cfc
zad78fa1859cbff9df373774a2f5ee371a1eb7609934e287b88027a5341d86ee16e3fb9b707262b
zb9216b975bd8a164e04908c6482511872877843a1b7a1af2f53d4c30b30044bffae88becaa279a
zd94a00b2e8825a98abe20b0dd82c5a8301e3145ec5a4235f350699a7e8fa4d4e8c78ecc2297008
z47f16be4be73168b6b1746c9d34607caad86b7be6264a3bb0dc7b1c7d8e0eaf98822e6ce67d9d7
z4fbfe22e51cdc4de04b128472c086f436004028b7b99842de362fb1e9157af08082acab4ddbff5
zc0c147fb14d2f0f9190dc6f53323820acd92b68c3360b6709e594836f575cac7efbff08d8623cc
zf1fcf99212b9b1186d4ec322118201c2376b3450d0c7f1c33bc26c260f11d68be5b0969e371c75
ze31e681c9f981368001f5a5336a9cc4d03214ce6744dd8ef252e9b71b4bceedad56050105976b2
zce959cfbbc8e181463ed67ea56e02bbee6ee373ee3daff7abf7296d6bbd63e3477cc2ce483b821
z19ca2a61b7525e67e1281ea10eca73f88df9ce0f1d3b305e0cefb4d5b56fae2122598101216700
z484d23b188952669ec8f45c5aa893e53e38594bd7906d89fd8622956479c8b055c33e2d87c53f8
z83e7f1a3e529aa202986998097d4b2d4540cad2035e1e69d19c4b50a17624c0f9f715923b859b8
z491b66f8a624686cbbfacd48aac8e1a772eea9ec7aed17ef16eed93c00cb62b9cb71d2a5e8a03f
z79e7ee8f266595b8f863060afb3cb60ccb6f710bb538f8d204701d79fbb21bc15c85dcccf536c1
z5aad90c53453338baaaaaaceb8922042bbd4171aa058c1611eea1baa16009c783140d0842128ec
z5bf06d12798bfa5541cac71d179f2a34d889618242e3e24a822d03737be00ddf12eb1cca51e04c
z181ec7001c6da54c6adef76f4723632bc12ba98e10ce5ac5812a13fd7b0747c8b64855c8ab6cda
zb2450cf85748c3b13a1ea777e93a638cb55a909c68e19326d3238e4a4f629cbfadb06d5ac3e452
ze9bd98e736c3361be9da352037da4a4152c0d46d66c001ba8386d7c6af04a9f77b4bbd018fc77a
zeb88cff451c29728d29f88a195d2c42985033e421008b4b8dbd12f29b423ca8afa46a931dbb904
z17b123fba9af073fbcf1c18a2ba835ebc4ee4806fcedbe39f5b592e49af689d008a6ef309544f7
z43bfc0e9d20cabd11e3bad9c96d3103eade165dc3a85414e9892429296a42d2129d72f148dcf88
zff0a16273534efd3375d85daa4631de425274a6fdf6a6bbb37eecf53cf17a86bf5723f3fcb2eab
z8aa02a2b6bd418ab5e246c747c4af7a9f3a26161addbf1276df499ed430d0a2c46b27131487333
z518828e487aba873bfcba369222d3034a84f744044df1a64016688bd22ef3755b63091f38cdb7c
z13209c0a4dba9b70dd91b574d78c7e3d5a764cc0f3c899e00a6caef536d86009c5026b8150881e
zba0b774f6775e571f38fdb444926bb5ef96b418dc88c490d3ecbbfed0fde7297840b9782271fe1
zfc30e5a6ba640251a779e12140f925091408c07bb715ecb556df4c0816b048eed3bee565c44d5f
zb3fb535e20617074ae08163f2b4b6ef9da391e5274f61acfc442459156d91a20aa701f264378b2
z85705b66ea3ce2791c5a3d40896c1624168f5f3c858dec571287ec43c823d4b3fbc5457d68a2fe
z7766b2e5140d02c67a75275672d999be54b24bde19bb386582083a424c2e8d37463a378c4257c6
zfcfca1b466a6ba390bded3e5ef8044923a18aa206fdef97462cf1d6f810e48d7a908538c343577
z9d51054a5ae97915517c1828d222360ddcc808eb29c13ebdd8c8636b66896834e1aad986e6d44f
zc738ced522d3a13551040825a8cca08b38743b41f07f4304fe4df74bd5191c3698baa7d2b19401
za4794a1f3c6de040b59ba5abc3547e8b54b8ee925595a311b68067c743d92168f1d1696980839b
zd92d284706b1bc1b54e3900064e6ca38c7e3515709710aac1b83275fdfe7bad8fc8026b87ca776
z0e0d502876920622dcfba8b2aabc3bca7306fe5e74ecb2e9bea5eccdbe9ea862ac75fb9f15ba48
z07ae5ede2ae0c09b3ab90b6bf9e6a830b54d2a163bd824a9101dc1f35952adc2b427cd7f3ade02
z33fff0d7c7766c5e4d71621d9d08642e2b63eb4576d68d9ddb7ab079bca657527ff081c673aafa
zf136c466fe3d43af5cb11e3b5857dc7465baed302a3d0d9ed5a91add2e65f8e3326e08994b851c
zbba75d334a6d2c3d249a8f92c56c52e3bb9fc2e572ebfedb9a9b7667cf9c78e9cddb44315a515c
z318916d45851dbfdbc1dacc67f599b80c02473338620ca696b885e87b24786816fc1a3283f9279
zf007b42491737ed607df56e8f12e807a86d10d65aecedb07f83537f5d7df513d8dafe1d6f3fd56
z58f4725de74daf151dbb8411e248b14b3efad389c0c4852d0d2a1cb63fa96ec401b1910323b6fb
z92191cef2f394238fdab4daaf93826ea594c7e193a9ad36df1595daa5bd1d1b2f77d9a3e58c41b
zbe7cf2078c85b570d272ff9e18437bc2fb174ea69dadf32bcb3cda65b6e89a1d6c7629a75a8bb0
z5e1dd1372e9db8eedac9c9360fc29ae8150af94298773ea785e9785e72345f8553eabfbae1287c
z1f5e0ba63343cf511d256e4e4d12578253d4154af2a319bc863d704ae876711f6349aba8f4c8c0
z2fccc9bf1f169e038918a6a1795775271e3002f5bd1cce9d53c49f79b65f2643f53a2e2e4f0400
z50f4e5996487b8f9e4333591e50a5cfe279f8c29cb37692a19d5994806ef493c855f78310e5f73
za56a5f8de1e0dd3786a50f5e05efa9c37794de9a9e9a542459d4c2c3f6ce75da391cbfa72d8539
z371e733109afefed63ef410235ed97444ccd449982b95f05c40b271fdc06a90e0c539e7249ff64
z77d417e3895234185ae1421724d8ca8b301f7cff1a8043edec71692dc9cafc4d3e81ff485011d9
zf1fa9dd4d7d12ad824153961fbe445909d238a1168fe8e04bda85ad8f1ffe8a20e5c0f7857c8a2
z517ef92109f1b1aa9ef472b667d29cdcc84a23131abfa11eb231241e963ac4658f9db22fb61e0b
z8ea19c4eac429c26a10f86b71dbe99e795962f0c59c4cc6b549759fa9f3762dbfae257ba1672aa
zd73b3fa5e87a461cbd9187da3c9350ca8951a46cb611dd10e958f8d188a58ebfdb251ba01f0263
z0556798ec2d127f3b0a78d7f2138225b3af8e9436d1f0675b56832e68446d8400d3913859ec3e5
z9f7d81b81da933c8b1d89a7618ced0a4320339e8f51fcaff58e3c0d6cf40aaa23f402722a7f691
zd80a7e85952b0e37ae2f05f9f3dbacd39a427d704b73fd2099533b64df995790a5b6c34c3659c7
z284461315be98e4094ca980c0326b4c9ec604127e2fdf567d3ef488994f8a29f9e545ff1c700d9
z4e61e5514d5b3814f2ea4a70e1db3b613fcff50ba9e7d27b44e1d8ebcb0896fff47bda08335788
zdc3aea1fdb239c354393549b6670f14c5e814f56ec90e1384b27e94950b379f3e8f12278ece35c
za97ff12e39785162de07b8da5bf97ab8a656668378ded9b72a0720714d7356866951f39c8330fc
z3b8919eddc1448e07bc93468e82d7fe70ed0f3b4bda606589ba99bf97ba21a08379251d2a554be
z4062d766a9f67a8d45ecdfe36170f668460b559e5a706eb7848f47794801f8c57bbc1dd115a313
zb22575af55bdeace1e4b1cc22c3406e6d2ad1c10d50bbce996013da7066c9c0459405e375b3cdb
zf41847380a1332387b9b842aa63d4ac53581622de744ad4fb40158710e9ba25883a4785bd38e81
zfcce20bcb64091a79525c27de2c92ec4f422e95865ff049363d4adf67b285e7f93855cb7f57d29
za827b8e5fa9ed0941d10dbcc15895fbd9cdd654d87cce8abc262c6d0ce4f324fbdae1b8f58442e
zd883c63222f6b15edcfcf520bc771cc4ad9174777dbfe0db14c4d5f81bc83058463ad8223c5732
z00f79135cda2efec5fad10db1ebbe60630b1906c0e9354926539bacab13c7fc3c51379c8fca334
z3e5ac85361534fae5041a9465d80f6194787e08ca1ca02e5e8b8bc47be47eb9439a7ffafabaae9
zaa6eca6b419af711ff46230f9bed17c4fb54a4fe14415b839c43be65185380febb92c81f264ff0
z2459b76531b1b4a4ea2ce4c2a1d1b0e31a9adccf02abb29b65fb0e53a4922de5cbf4fc7efe831e
za17ecd31b69396a877afec2c41a94124dc59291f6a48959aefe4042ac26db40d8263b12e8e19f7
zbfb0a84359e7afb37c5be6e17f2b47edcb56c73ad368813f59d3cc71bce60daef67b7699e8f158
zfe741e420bd989b646b4ae1f666533e00577d353a54321efdfd53e863af030fa417f4f8534e7ca
zec181b2317ab4f0151124c0e3748fc80585bea11ea2d3391cba4c5baa0fe5578bb9de44d29594f
z9e109139d397135b6408c2758a144c31b653a5e334ff02a12a326c0f4530d708630f0f1862d967
z737bda2e2499aa356f5ea9b02c4f2369e1b4a5d01ca4c4914b5fac5f1eed417fbc664f538818d1
zfd7578a139393af97986cf4660d711ca2448ffcdd3dfdc7a617dbac723c7e12a8c26d73fcf3483
z7e30facf9ae6a5b8c7cc261b272ed0489fa6faeb8b057ed899be02ebc884b061c0bae2fd265a7c
zfa8177b0ee496cfd2c25ab26f387dc820852a4e0472a559ea80ee5634da5991e6382c956cc9c72
z6561851066eadf8a03db694d0feb0a9df5e5946f32dc4d1d7dc12f88b4d3c5545a77ef3c64f260
z5836edaacc195af30ced17b4d4608831770706ed2946b36dfef1e65e81d2d2e8fa588455695eac
z5768338b7ee5d1e46662494ebef08f3dab71499482194469443c804c904c2c939eda18c255c210
z44f03b4c8b31c4f56a255bfe07a089f91882d53437cb4bd8e72b914e7fc215311a310cc4e5a5f6
z9885b30d6e08c8cda7a89de284c61c496bc104f7444f90d60a928da75743a0c7a87bf2d2aaf1d9
z334ba5d5cb7aedd8bf83e90f3c7548b1c90aed14f0fc3074cb86be3886d67059ace5a9a53b1925
z3a80b7ece8201412bedac47b7ad99266218ac0b523f46b78f925ebdf5d0b4e304435ef31d79b40
zdf37bcc42702d188f9f40cd5eb97f1e2efd2a89cdee11afc326a30657e52e88f9311b92073da30
z043992a24cae11ce9f0bb5ec76cb0d3400f1a26cfff0ad4809eccba7942c6b37be93131d7be6f4
z88064d956e760d8dabd0a6bc03287155282415fba2ba120b5e996b4e9d60584d0a5618da804951
z0da55648bb941b0aa5995f524d40d961ac5a94ba386450f3eb72463f4e6834ba8986f3e7852ca5
z8e04a7668e4e33bb301858cfbaa48e1ae0b69bfa7e739318e7bb51b7e1a7fa04c90176af34e3ba
z5f469746c79884ba707cebae9d8590fb07e18dd58c79e70796ad0a4650d398a362754f3a14d6af
z4c994019590ed1ba0eea6f381216ca99fc9323e92e9e866d35b7bc152d70bd675ca36bbdc66727
z63cedf23a0c2b50cdb390b9a7ef52f1c02a604395596dfa69ec4a223074e00db57b4d549fe3269
zec583ab01291251c3ab3d1dcb6bd7977ef1dff0d99e8ed73febfe89b373371db4c6c986410b263
z21b17bac3355c1b1478191c320ea0730658237c609fbd30611cf92504557aa66b4d04778745159
za8359e31891053b88a91e0aed844fa8a31b3ffcb7ef874563b17b583aae55d625aed7c0563fe94
z3a087e2b397d14cb47ee4401be44817cf354c3b1375325e00af8ef6f8c77cd41982f49857c0c2a
z6b96370a32407eb2c6213aaa0b7ad56860e5b84cf27b06e4eb63626cca1a4d55c9bde1c6034ae6
zbb2802bf896f8d5f1b722bd56853a3392d70bf9fda6d86915dc406e134c4701090560b4f4610e6
z8ea73eaed283ba2e58ef23bab2784fded922762b252b54aa51ffd866bba2e2f12eda6c542ccf40
zec5da16cae4c779456c94ed2f16e62858055fec47dcc5c5b98e6808c7a289c180587df6f942572
z6eee4f4a19096632c3944ce6717bd1df70066f04c612fcfb2f5a94bffbf789edcf5a7d75562a8f
z7a41dbf74b8ab478d4779711fbf05a394ba0c2e39397e626bc64db373558adad7f762af4452d10
z3475b09673f9c5b33a24def9cb70f5ab11ec90aa58d21ec6542c0cd5e484799eaa6b9b35fc674e
zfe47067a6ad360414da17a4a3160de76e9cfb92b4fec4b906a36b0c977033bc0cac38e644d2176
z3b3b536593b525489861735832b815cf3c110646a4d7e8e622608a817db3ea21b6ffed290fa270
za8568f1ab6ceb544e286db77411f9bfbee057af49e7e2583ee7b87cb92423ee9a562cb3b5a0000
zb7548a546eefd4cfa6fc9bc92801480bf72fbdbaa5333b2e60cf7fde7c0d31bd077656e1b4df49
z5b938b803a6d03395f4e036b6768c25dbae1619030e8abb30995e5d91b8c015243ef66b626615e
z47f15e6d3c136eb5374d2c55794d928aed519d4cc08f13a9d46e3471ddeeee7b824dd6bf5252ff
zce4ba93941bfed611cd386b1be1f4e9a94e272cd1a6c6c5b1e97a7ac01fdd7ad3fd48edd5dfae2
z322a2c7a229ca40e6f69d9b743a8b462204cc7026f220b59d3f79cd0de9197fd6253fcb9529d96
zc448b2838358944371bd63da5d8a2de7286d3625189d5d05eb6522f009ac64d1ed0573245890de
zfa6805fd5a78250cca643400ddf727285da42152472d96c351c75f08f9993a743cae549ce94d4d
z757527c410d58bd0b0c4873c6c33e137a3cdee2cf91c08ad980c3c8273ae13bdc49c237996cb2f
z50d3cefb283ffee88d3edd2f179008fe58bb6c648fc71745814be05c996ff126cd26a77fd83e34
z6a551d70872ebe037e880fb1274b57d12a2a8f57bd5ab64d07e6711e5810f7b356615ff39736ad
zd35a487ac6005905f6df19fada5784e986694d823ac99a307ad8773f2e2c3152f670493d053f28
z29bdbf1f7b9f83c5cc0cea4f4faf690f7b642cd5e94e94b74816c70f74f1e4b30a4ea1f0ea700b
z7bf2ec14ea6ce11cb2b4a42c2a493bb578364dd5ec824ab56995743afa681afe10ef4dbcfdcc0b
zebcde24c8a7dd88dcfd88a850a54877a4887942e18f542852f2c822e0013ac62cafda689ae586e
zf925d4600db3775d6e592ba599b6ef1457a1d9a8336c19ed71e888b1e80adfab1c257c425d63cf
z79787022fee69bef21d9e0f8aedefc51b1b42e5b09065aa599a08e457c1c7080d53ec499a7b805
zc84eb300bb8a579f434fb2d56e84bd74481ed8c5d808d5bfbb6c1f8b3cb087023f5722bdffb990
z78531a0add2c3a768201d89466b1697ec434ce077ee58e89b1b08fa621eb7c9dafeb3f68162b90
z9515bba76fbee6d6becc2d6c7cdebb783e8bcc3400451726f42f7b66c75a5b933fc7c83ca000a2
zfa3b32581bb9ce6ffcf10737eebedc40a8726db96fe086b484324a7d2bb91472927d8eef53bf2d
z987e14551adccf9c3d3d32731caba6f903badddadb10aa8eefe9066c6e296bc8d15ce067a3498a
zfed28c0a8411bbcaf0923466262243a0c6fc6ad370cd47191eaf01177fd07ac81bdf8c17a49460
zc1d137fbc212eb0259ed8f92182555592c70f1023c3d743197b8f2ef9461d785e9958f5583b211
z8ddfe16843b0a3c8679ac1283ef2d7e24b6f291783fff5f06b5ae34db13a101e32b6c94a763b4a
z290782f8512503c04c1b44eeaeaebdb6bb1ad36ae42dbfb7160518f00d12ca5d6c790561f3e0db
z0ed8bee9eb086871d19092470a6f041ff4893743cad373e6c450a3f289dddfaf3bdb1bfb32cfe6
zb3ac8843d41f8d045384bd09c82e0a3b217b363b1acf3ef685ac619b57092b7d23c11a54b34854
z59d043b6024fffc1569e04e8184e385ed762a8d8601eb4c7d2ae8e07507276f348c4d304cd24c4
zd92a91758d2f14ef8ecf1a0a25a8f21e0bda0598d7d8fe096030a99c49c25eec50138f5037b022
z957f82198b5e1faaa8f4395143fba0bbd217802e0f364eb59da3af910d95f9bf1debd033a882cd
z8189358576341ec4c661ce841aaf2d96210e46256ae45121f5fe9974420f9f8dd313c472045915
zb303587fdcb00740b88b1fec60861c263844b5f3acc581d3ffc3eaa0f38fdb46daaf702bdec742
z63157f66ffd9a8bade6d8c680e05e90ebcb6661caf89e4f9e5673e19206400da72f53e8190809f
z702c86f177f8ae4d44f864ffcbdc06f25ce70878889ac25e1e620d3300fb4c14f9d13f1bff5ad0
z70944a77288ae326c4a04ce7e7e5669e07f8f9124661e4bd147a4dcba82eaee8e756808e0f0265
zbcaabeb6ff62ca1ca6427c37952be34016ac6eb549eb801976df603aca286757d96423715871b1
zfb760cfb45268f70bd7aa0e78f71926c26c2dbf5a092775ea993fda26be545802820ac4c0b5089
zd43c7b0dd1efc77f40782c6843a3896b14f9f6362f42ed1e1bca83e406395ba6045986d0cb1489
z7bcc67c82c6fa431531fa9f68a080c4a1da377414f8bfdd8f015fdd2b9b88388d2a613e2835ab7
z47e3387f317a5694d6423ea94f773cdeece67f893f333d90a1aa5d854ceaa46fa5d34d6cd0e982
z50b8765f561f4634e8535c880f3f0d51e29cb5e03b5717c0c7f1c3dcc9513430f3c38650586426
z36546bba7cd82db80dfbdc6fa14d9a775aa95b32673ae90f1f4bc5e637134bacdd6f9467e01f53
z9fa3efa64d0f3134a9bf52b4df111b5d0083b076b5719b06185a384796267380caed2ffebc484d
ze52a25a53b79c60c1daad280a03782ef8c42e1f10c6e64ada6c37c6be0340fc13ab7de906d9d13
zef7dcdfec17ea00c0e0e38ccb1c5ee8151010755b727996a81485209e7661ca0955ea88c9fe1a3
z8c53536795a87bf9720898d81cd5f0cd90480d27f2c9f221cfa63e265fff482621fd38cd9a3e56
z820191cc13a69fc23a3e35a5fef58c1ea7f38995c914d3bd81c9cb4945ff94e4981a46f7b59652
z6d06076210651ededfff24cf51d32581f398f339da1f1062e7e50dd4f21b98a2cee964a7d4e52f
z0e106f43b1ae072a67be44f8e628a5c7cda759bf878a841309fd2a46b28648aa75f38bc1b9e3fe
za4294e9fd41fc13be46532bb36b449ab079ebef86234ebabb63b801ca1cadf11028187f7b99e61
z0c4b2b0ab63546576cbf85975271c0c6f7c0f7e5c6f69ed79d130fe8fa328358c0b00036f86554
z81ed2547959906e4a3f18af782f266c22539660d62667b0f7a0ef53512251a9867a8160790528c
z8f847447c9fe2d39ae7f40cd12c43f76e95a1b26990fafca3a37de76abbfcd021e9d381f1240ec
zeb3f30f176e8edabbe94cd02626635f2aa7841f2c7fc9870220de2a0c2921f3288e6b4e73d5815
zc5c90ee64f8c05af950941b2f3f928d7135f8f11f5a81d782d1d7ac27b177251c4005a2c472597
z9d2435bdad2866bb392991f053a58e2c17f84e72b3384c53f5b4cd7e7af774cf163b7f8f78de33
zaa08adb14caa8bc848f76524f206f62c26114cd21c78128ccda2dbdd1002022f82eb5df8b7bdd4
z6b294d837fde059db3c8aed8f1ff6306e7e552c275dce83a7092e9ff6ea70e8813e91c089a3816
za9b27b953035eebc3a58a6977b8afd722e0689d60f104d453e2d4c55671025bbf023cc565d3b2e
zaa31cd4f653c6a21028a6bda27ffde74869681f957630e732055d41592437dad7ef5610ba517e2
z64060cfb657fa5cf5b34bbcfa0c0619ce45b2616a04705e5a551549a41412b3cad6d51fe1cf83b
z734b3feb2249f1a2d54bd0d0cf67336e9374a27281be979fd8ac2595a6977e72655ee790c403ce
z2383166f7275b747bde68cb695172a5e11e20c4266648a914864842ae8c497698b1b2e842ed853
zaab39db64fb5c606918996dd09aa22285c4c57c629cf475ef201b37c74d04082a433253304d7cf
z382342457b2a7a22acd5b522c0933f271b7689904d5ad7b3fe4424c74574527bf8350353aff8e4
z6a125ea2dc2ac88c135b59e36dc3d02fdf836d3ac6685ccc652f20748a04f63fd41b35580ae2ad
z19e29f00a0857f2a872abe81eb873f59e4356227a49ee1e422139648eb5ad50051ee0671eb7a52
z538d3905bfe761f48ef89f3bcc5c733883e7895877c3611bdefe3ca68a97c752763f396a32af61
z31f28f58cd90921723c25ea3a99aded16846e9a71712721469aa959fbe9e1183dc779ade811d03
zaf5f3dbc544c09360a8ab022d39158e403280e7946f446ece38ccd7b3fb9df908ff8811b6502d3
z7442f30f691431a0faf4a9514482fb1347758c9f7e1be469342f43876a2290e44da1d65f4d44ad
z31aebc550a6c73ffb2fa7dbdf81e80c9627e098a911775a7784ebe1ffcaa75d7b0a865ce1d7c1d
z13431031e6fdde600fd965cd8bcca3b18955f14126eba0ef0b18b41c5eb0449b90864299c45596
z5efd413dca321fd19ccd81ed6820679d0e4fcb3b587259a3e32ab210307cee49b0e74f201c4572
z4d5b97b8498fe0f15ee7c4732cb96bc7e5b3c40a75c4f58a57ead30f680bf6c4c8af4ba6e79cd8
z205a9ebc0918260e4899c6b9340cad2c55835c0473133c7a3652775e260c136dfaefb6db27d8be
zaad456f436716144f35a12b88f9019cf6005f0b89f774cfe65a0cf67b4adff489694e23212cc06
z401df0bddbcb71e54c97d5266079615ca9d04cdb39d2ef549be7f50c7afe2288d19a5b7076c9d5
zd32e65fdb9b2de4d4ed9f74e2546114ce1966803b0d5a24aa8bfbe661b149673bc9e26c8d4a7f0
zca27aab3db3a37422aa9712ff975d67b4dcc7774194deb61efa7d83c57228268061fda00fded22
zb9aa349ccb786f027335c8e1f36373c4a91eb37f316421015d26a99a8dc8daf3f24376c954b81f
zb3bfab5b26322fb2f5ab0db7417ef2aeeb14cffa5ccaee7926762087365b35eec135d9e03c6db7
z33929edc15d86d3bcbd2d3c62e996a7c084870baf37345da66a91c5ce56c0def590e64e5c7d44f
z4bf65281d7beb65f0c711436eca80e5f42038bb01cca25050f44837f80bc958d38dc1270a6084e
z24d6d1a5856ecc6cd8abb958bcfead940999e93ef8920ff0baa496b7ccdb06bbbdb99dc5682343
z3a3a7f5b5982596e9771db64c70ca7dcce07beff84ea4be0a432883bd67e70b814657dc9c4e947
za40538bf40ae5167101c6b37005de7ef6ff1f742b42dc1f49cd5b6a1caea1e080220415b1d17b2
zdb4d3c56cb27935ea219f98a92435d8866c607a7ec25e6c3f763b912ef844a11b0a1f412693cb8
z3209a09c950e16d15106c11d3a7b8c697666559d67eec2f229ec90ffcc49b6d4f35e74cfdf2db4
zf89dcaf19a441d680e008c6f07fa1d47ff45b1fdad416f97e4ccab3dac86b39bb3908bde49c7a9
z5b1d51764f48f263c2324fdc48e584b91518f644a5bcfc39cca70d77e868e14b56bd211d8ce465
zd0d771b65eed6c48e75376b9bdd9d1ae95320fb0bee352d2e4fc70d6ca72ce045240eb270df5af
ze59059adab92d4a699f1078e604171389030ed52aaaffc35841f135a52c3bc71305283f1e68c07
z753b161c9e069d753250f0d41fd726bd72f00e31aaa519bf889341fa343acfb5a6f18e6b4f7c17
zd1b4b68ebc8deb20cf216239bde29204d6ec5dab35f831c6f59fd8dd670eeb2654fdb3a9deed6e
za1a841cb6495fe687ab17df58f8877be699a3fc3a0eb166a79aa993a2c0fb73db548985bacd43e
ze537edf375f952c7c37df813afbbce9a8393539a6adaf90628636ae3869a2155df79469f06aad4
z72083db2b367a9f08810fec479ae5dab76eebf947116dc4b84aa8792f14d1631da757262dfd163
zc38ebc380250eb12f15b1d1ecaa7397bdcddcfdf9e7eb2d30c039fb4f69d2576a6ddb3bd43ba6e
z9d46e1a5203bbb48eb9d7399b56daf1182188370cc567eec912732ec9212034e5c2e7f86408387
z0db08edc146ee4b828814d97dbdba53e165657a4ac4bb871874861b3a0cfed9eca4f95ffdee1e5
zd1acd3c7bade840aa0f546fc426999a1d92734889716dbbbb3b9c901694a27f2e78b8e90c167a6
zea6855fb52b81c02a3d180a02001731e47660ee6ae4cefdf63c6dd804adfd5a6a6804d0859dd62
z8b5ea3f9352ce4ec4c574cae6c996685e80a4f03bde820a4ff45c82c8573675b45c189459d3b2c
z434eeb7e15a0bdef849ccba4c211b3fb0400d34e69bba848113e221971c53d1b92c82d48a284aa
zfb46871c66170365555a22f73010fd0cb30a891614fc3990b308e0e2e7cd3e639f3faaf077bd07
z7d4402ccff4d286dba86907f7a86eb0d3dceba6ec781a814a668bf4599ed124204974f01ba9c45
z74b7fdb3aeb1a64b96ce2f40e34c59ecb5ec7e32ce75d48718e133971b93b02fc7d26cb9262d0d
zefb245e3171dee1919cdfe672e44b68a617c13bab030a56dda4c0f2e8cbbe313bb0cd25428d159
z9f22520597ba89fa465307448cb5678f46eead50e94122e5659cf226e7c21abeefb0f44dde23d4
z60316a7c514677017f677e32e6108489de868b2692c60f2a1d5ceef6730cd83035c6fef2b4b4a1
z8499c4e9b8edd9a5590048bc3ab3b9b45c0d82f418cff8f051197707375a6b19fa9e229856df13
z1a3efe09e5e47acd82485fc34063f8732c3d9c71a2994cd935b43eb89ea0c2239350752eb5dfe7
z3421c05162161c0f215782ff8a16e4c6e47aea100d65aec480ef43cb4ee58a29f3e221d7a32494
z406a4499b4a07423f72f78afaa8ffd15e6ebe479a06776941ccb60d39fb6f2ed20ce0dd6e897e5
zc1585c25bbf710f0299f37cee00af1078338ba2706d17a9dee6bd3330d5601843f792747f5d312
zf50b322aaeaabf0ad1f439522019c7f0ee515229be125772601c0aaad054cd41e04a0d20f4dc80
zd3dc5d10e2ab86c1283f62a522879f466faab09d464fe0ba899d689facbb50316f46a868dddb9c
z235c718ed19eea63e1d3a175a79ac7741c6cdd489c8c646355ebf4cf802b4f0d03147eedf4b371
z223ed2ad2b80896722a123c06e4d200621c18e66d565753469fac1124418bb02cda867bf780139
ze2cfde8389f662dbee97e18e28de6e0d982fbea9f3912b25274c23abfd09b6282420ad5169f5ff
z8d41fbd4de3e000974dd70da496c7fdb18757582ddeba3161d30535bed143b59d2acb10b5e603d
zaaa36fb8715fc3971f1caa068a6ae264c179be07546ee088f86f221fecc8acdb1f4404f8d10ebf
z7f1b326a561173d5120da454ece5856b6a99f767d755320b9237b104db5ee5e98252419d743d5c
z3b4bbcd349bd4b2166779a483fb74f06fe72d6b61671dee78f8cbdb98e2d5961cf014def39db1c
zf0358d44591c62fcba0990a693efe127ad98cf45ba68737ccd717a8e02e3e3f71a8747ebe33840
zfa5fedd292ac8a7aa74b67e1ce0e43da1b9f569628d3ae01b5dd7c0c379b3c194f73cb095cc2ea
z0c0540a3a95c4fcf9b629ae6744b63593d42debb543eacd9420d1f0982df0ef5c2270e7b142549
z133ebafa05dde2481c0f2539677f91ca3cfb7dcb3067c138540d4a62ec6dd10976f170028b7c8b
zfacbf77d2b745bae84ea7dc7cb1dd30d9a817b477a0086e7b2e1f56782ed88cb857f34129e0cc9
z5d6fe1c34e29dcc4fe6818449bdc27f6a6fa012a51a2920a43ef9dde70ddd5198ef1809e3f106a
z60bfc618d7cdca888cec9a8feb1d18d60c7de10cb8423810027daafcb0e9da52b08551178f79b7
z0b5ab07d15211551a68b6054501b1b9d487e59db231846e37d69e1df2e07b2f30b5aa63b9b39f5
z2c36ba55df0aea49bfb356d05354ddd6b2de61b1d0faa6abb973c410f5c8f97a627fc4d0d37b32
z74ba9e048c6ef01f31569475e6c2ad782b9db3bbe237a3834da0e7ad6dc3f8638cc5b22d798854
zfc4a226fe9ce4dadfe93f11caa0c31923c1f991c13a4a057fc3e9b0937edddaaee2665cdf9bd1f
z8d7bc1ae3fc2b4d984952660b7cb1467bfbb5a57939fb6e05166da3f138bd211ff9051cc6e1094
za94d833bf192f9c783393eed990ead977c17459342757ddbedf323e2f71187509923e7ca04e87d
z5594d38914f685ec206a4890e7c171d7fb7e38ae6fd3a369f2db46d39cc9d31692b0cccbc826e7
z54687290d85eddc503de3048e26427764c1571a87615aa45d031d8392e7a13c924e883cae6da54
z2d0268911f6de7bd297957bf961101fd460854ca677ec85dca40f6550f7928641fc5bd98ca334b
zc6b70b17d05c0c636e48a8ab94c3914f6e01151da9afa060b50c3ae5e04903f6a6149c553ddeec
zb7555ce5f0cde307ac89160828cd095613bbe696f892334ab0bc022b9f84b4ba1772e73a21700c
z7a0b860bf462bd1d87d6329bc9fabf266db6e284619438ee10e51bdec4b1da0e3ee9d6000f4f03
ze37450407e5f9daa5d6913580fc7f0daf1081a7374323e071d6b9f93ab8bc46e2e416a3fae1552
z42a423b827c1156ccc46dd11e1e38101039d85797e81bf24eeac41f51e502f0ecdcfa65d0beff6
z51f9a124ccc3687c79a1ee11b16913e3decf916a4240cb286ed3714d74b783aa31f11dcb633d1e
zeca1fc49624be434dc7d8a8aa16ee672bf3def8d128ed09633b21197fb47389f1cd89993f0bf47
zca556d921aba6c80c495ffd96af5ec1d366297cef50f47239637641634a10e8ab756375be6afc9
z4e8a4ecbb8e392bb08e527e200e298a6855e85389a2c5b276604906217c350161955911acfb44e
z65a842be1c386b2810b8c54e5e877f89326c2e8e26797f199e54be525673e9412bbd490978535a
zfebe279928fcc77ff4edcbc475a19d0ae4833938b200db65d3850111c09708ced293076fec67b9
zdc70859cc761be8249a7ddbdfdfdb36bd06a50ae5ac13321b501538ed274ac3af9a50837803f94
z34b5d98d0dc5e8a2d8c001f4f88588a51ba0bbc5656baf1efe3c1e837376ed1998520ccc33e1e0
z22ed4998457f74909b71a67ffd7f05da60f4302e79752a387f02bd4b721da58745456f24a777b0
zf6faa5afaa3059e22225a81fbcd515246eb967620294d98cf3be05c2b68785777d7d6ff027ffdd
z115ed4b29d469eb41e72ae5b17b9809ca2f6223560b481764fb06677dd0a0b33533be5e0381018
zd6694b0dfccb112f3afeef82a0ced88661444310069ebc4173aaedbdb2dd2037929997980b4780
z170bd47846c137269c9113dcf2faa37d4ceffe994d60ce3784a46cbdbf5a1c3b933a62c4b81dff
za4b4dfc6cce7a06f8f27dadd44c6cb382ea90a11efce79153511145500781911591be7f208f0b8
za1d4a873dc0385e2ae6b936643e0793e35060d0ad9c913979b05dd862435ea166d6f8cf2e910a4
z6471cd9a3fef30dff7f4a6141d20e3dfc6b84932a2b0157e122ca62d7ebd07537381c4de545951
z96eaabef7cfb5e8b0178c1394c7253e28e3a2f3d77778d02158fbe2aeca4b04d8795dac01a1050
z8f9c3570d314cbd7186049d6e2bf93175ae6b713e84babc887180a2126b7e4a42297582d0f6c8f
zd3dcca130cbcf318953904046d31e1b21cc5da41b7b430092616fc07c811f7deab7761c0d34cf8
z5e938141ebe02935a909e0a41d57c1ae43223b5189f601693d3a2cfa6dc5e9f753e05c9af627c9
ze9c2af93498470860c33241a81407a481813359db59090bddf750364af1e77271ae74796ce32fe
z2da298d3dd7c734548a6ff541b8ffe0f0a3f0f4804af7941bf7f950e469e2164e2f77a5d5f04b5
zc1a855c1c20ffc3281750dd48a5c45b8f1c3e2c1cb251236a66ceaeeeca0b713146e4c5a560abf
z481bc9d91562df97587ca038b59534146f73533ea2c451c5d3ccbb8ff8162706134db61629d3ad
z7fb10c1c2ab104840f7da2f463a808d92cc1ae81dbce5fa7b4abe436b91fb177532c94aefb17ef
z7c9af9526e31973ab0fc643b22438bc5ebeed0b7d85b63e444b4214df6425b24b26b60af1f9d0b
z4b81b553ca008df7b28ce16aaea6da4dfc5a46a516c377110fa4b2e97aab7f1702e58a2b67ffd3
zb43e4e81691dd7abf7fc6ad2ecb0ee69104c32ef817c94fed82c0de5c3089edce5b2a37a293644
z490eb6daeb05c481d8c718f56158c1f3df106d25c96589cc45897d663330626b20d7dcfafee4f8
zf8fa343529a3d2811973f166cce4682f9a59018f08da4e4129adbd75281c03e7b5fbe2dc5021a0
z789fa810f5e7855af4875d75404c9f5b19f8173129a2b2debaa1babe367bd4501282ca7c9edc41
zf9dd80177f216a4553333bf48fa703b41dba26a8fffaa20ffd3b3c49592af544bd4abb9e1fcc8c
zd08b57a0041d8ce9862667b34e761aece703789d4ab4c00918e55c949344820aa55878f24281f0
z4caf3bd78f129610b00e046adcaed7265b19ac1213e7b106ef087f1ca5c74277e5dac2c9e254b8
za213bd978e5717d5d012e02e74a83d2c2f7c9d0010d7002eddf059503a8d15b9684d8fe177cb3f
zbcfb554b093f443b5422683f30e7c31fd6e400fe4b225dcb8eef5c5f4874193d8bdbad92ac08ac
zabe0c9d3290c7c36997febbcf416b80a609290b75c76d6b1d22271c90b87543227604e0b6c8451
z53ea19e311974bef49b71ca017b2cf4cb27bc63d8456f819d651b82b2980b14f511c657d7969de
z6c22af148fbae3ac68e9c3cbe09e6d33e7309f239f8a624877452ffc46389bfccd3f3b78442c7a
z85a0966cd2fb7d340ed829f78d192551a49fff69e9ea16001efb1defaa0c2dd2aca7731936bcfa
z9839aea055fb3408bbd2905bcaa1aa632c989e216c774e632b973aa883db7095fe29d3eafb3690
zca18582505e466b3182dec1212ffda8ed94d41878a7f4a229d7742e483e0d840fa2aa2de30c8ff
zf94d5bece964c26cd57faff74954cbee766ac5daded446f7235562a71262fe05fbd7cf1f349e42
z781f966e82cb835d336e86fedd63370f862227684600d8f007291f73e81ea81a2200d229f15bb7
z45e1c4a1507e345626bc0f6c88864a89386eda092acd35414e53700d76ca129cfd55bf3dae37b2
z574fdf634fbea578cc3fff6ba5ad2e473aae1c8ad8400a472b44d415937da3cf2dcb15fb9febd7
zeb76ccfd3cb8575635d37886554ba95996196f6021f51007058f2deaf7d505384d8312e6948048
z1f6b12c9eb087aa80f085dafbae5e3ad8764877b5ef97b11cbcff75583777506da1f3edeb7f2e6
z59a3f76cadb8057c1544bb40e03e6bd9a7c684692cff1b527828e87eb92897c74b720822a3d67e
z4cb799063d4bdf89f8bc6dc19d68b892474b48b3bf6c28accb82026de64213c5c0551790bd5960
z535950fdd18a270fbc7b374afb661c82ce8c54514a806fd494edb6edfcb320fb7f0babc31111b5
z298c1838c1e9475bfc9c4eee7e138490e289d2fc343172c2414aa914694a371e13027d64828a0d
zb7091493dee54cdf224d327b4fc07f8456d9fd60f2f45f944fb01fbd4922a347d700c2550bebbd
zf17a968ec132d095131f4a84a013a6c824444707495528e2b8d348bd377e9ae92efb19d17aedc7
z435bfa7656870d64ee52c6ce883e6c798c1f06e490333c7d137c720885ebdb3f5fd6cfe2c2b071
z91685c724f353b5fd81a5873936c2b777bf91939beac7d04b295da5e82006501a53cad0ebb362d
z8ec2be4b6fe37d5de2e8bdbf72d54171e128a688d1479d9074baaf812101f031f574fb04c2be3c
z7aa4543105efd8cef339883db96e782c74cf33c0c5e7c17d670844e63cf475b79a7d719051747e
z84856ad2e6ed7425e7e6747de7b5c0c9e6773c875d0fd66d93c1d9f3d3016882e44282ccecdc4d
z260fe041a46b83f28c8351c630c0429e4ef901e937caf7a9199c68561e3d344625882a7846a37d
zcba90082d1dd01bafa268aa19b956a1515b91670fc21ff995769e8c619250577609ba97dce334d
ze07c45e70e5c860cab9803e347d45be3b6d1ca11b59fcb219e98eb52714d179ec8bbb329562901
z40222226ee7199e12a07f4b206b612d7506bcb9ee259e7ef1848b7e21d49eb8ea8248ac6be9ba1
zc4a55e3253489fcd67643ff62a79d18b7ad42161c37d89f0373d8d33291063a0e87e99b2df1b12
z87fe08fd2b1b97e54e379f1e38e9c55826f426b63b697358f2bddf30a2e4e37529839c6758aeb5
zd1113dab38f8a7466f7a23cd88136a9ac29b947aaf81a35ef0b9f5a3b31a282110bca8608728cd
z168a41188d5e606118186f00febfb6151355f6eae9d5dd9fd1b3a34651b51b8ef2dc86e580eff8
zd9e44fab1815627fc548ba4e404f3d5e9d0eb970a8101c650b5b41fee2511b1cf9e7fd0d8e7c49
z66bc25228680d901000fb78fb9771e857a3a8416dcbf2baba692168d0d38148198daff251a56cd
z39c6d01f399415819b42f2fc2379d865ccc1a4e8371042d9a0dcdf24ba736dfc6e9a35322ba521
z22177fd75fdddf5ee55e49427d6be3d07ee5b95b62d3fbeab71c02be086091f1c1206b638e8c82
z808769aedb2cbef205f48a914ee73ffc4e5bccead952d5ab233bfb209c9edf532729f87829edc0
z9eabc5f594600a93d18df095185b26678dc65bf53ef1319d89f02dffe7de3856b5e004f95ddcc0
z109201dca26d40cef1e6e2cbf61cf9b1700728a583656d01bc52b74d4ee3cc98c2e4f7a6017a28
z61979d1567c167bbee127f041265fe3687d138b11623a7590f2a8f038ab921c58be4b3ee3925bf
zc5a75e30d29ed5eda0448c5dafb8c10b10edde414bf1c6373fd9bb0e74d8abf0bb6a9b0ad59d78
z89e42a963b3692f8bbf48a99fd8fa4049e64844b4cba86e461a5684d9d548e5bb0fb4c99f498e1
ze9409c37e48f301af7f3c5fa32ab57fa54570d71b3bd65e5d0fe0e3a5c46ccaedc97e4a055737d
zdf48f0402cf48adf3f9e0cc8a246c1f712bde9efb7cbfb580a9452375675800ab84924b1e9ecd2
zd5e671d60e25d36585ed435f4840f4a244713a27edaef09423bb94ceffd8769178e89b820e485e
z8c134aaa62e574b05da2b473513af270424448bb64e45dac82d6e33afea4c0045029b123d39e2f
zdd2c3264a989f94744d47b5d56682d01e57cbb6e9d20e2aba916f8c42f99b8a9b83551b47b6352
zc8332e85eb257041a5cddd5419fdb1b7a00375e86e467abcce76579df8095d3898dd6c1501d208
zdf92304a899201af400bd20a3c9ab1907524dd59a66544b2ea67d51b7a2cee0d462b868553e4b3
zff4c7ac6c3c5e9e34eba9f92a62ceb320bd9bf351e8ec97d1c4cb8507f2fa57ebae26b9fb40988
z069fa4cafdc3e54594d44ebeef120d1974098b988309ed5285ab64185daefef1ec33ba022669f5
zf04c16df21543dfbc9178b5e439aa4753dcf6040aa138ad7f03f8c64ab46ee3c8bdc205d6f426c
zd6965f55df2204768f0e5b32f3ccd8380247f5ecd709ef52a1ee2c9b5f1292611b9dc1d3082f70
z177f13d1641afe8e88cc7cb6fff9faf5d03c9a1f137a5c2dc39fa68719ad5120657f005aa43874
z2963baa2eb8826bc97423b328c884e734fb2c358e77053af16475efd7c5d8506e6698aa8574ed1
za98fd7277c06498b586c7048ca4e21fae24e1a0a37414a7e80be502127dc53368feb03eb0c6807
zcc5806a70c502e31cbae7f74422119ff6f1dc5bac5bca905b45656d4c8f33796bc98e24dc3445a
z069cd995fe1160dfaf0faa2aa878ad411ed1b1ce82df71d60a171496708ae4935cc9040476a249
zc31e17d5846f7bdf1b1eaf8b3b304cdaff3154ce9340c9261a5dfad39e85c0f0a2cc8e097b6bd0
zdd7a66d2b2775c1261fa103446f8df909272325c26179b6106edc721df5b002456441069925360
z3243e366c3982434bff4c476e47edc759300f58be5b1a0a41c35d700df656d5d8247a6219e0fc6
zc68474cfcbbc4fe763bed3208917994629cfdb4e849e74b981da110d03a0677dab176e4aa8b6a6
z80df0e9a29c076a0054ad4133fa567e01e406dad8b7f759b7e769dd7bc28068b1155ea0572fd94
zbf7a9d69358308b247e827a7d4c817d7cc7ecb3dbbf736fb9b24ec1c31c3d3c1edc83233ad46e4
z0be258236a72c4a92d4df46b59533e84982dfe794429ca07fe3cab4e68e11f82c880051b3add74
za8548dbf7850c23617cbcebda0bb531a16a0e3a8b8abc74e1a03c572436b7ed2b3931ad847fdb0
z3793b2d5b7c8f27ccb80c7090e154e2edddc6db532ae8038b51f0e9218b11569d28f6da077cfc5
zc3e7aa16d31cf82873faf9f1f4380c4830e7c68c206fb383557942858b6b0fd5d0d852d76fd358
z29b6bcbd6f8f56f971ee5d5ddbff3aec2a64b7c3ad06e87c3a71ccfe74aef34d0399dbdb8da332
z31461ceae337d8d59a2a6af7ace0d4deaf584dfdec442f47557fe74c13d2a8388717cd2e6ac3d7
z62418d8cc355b7efcad4f6921a50564fa3dc48b905852338fb21ed81cef1c027d2866e2f1feaf0
z36e5a5735fe2915c7904b1c9f30da6900d44ec2c92483881d7d543227fc0b3509cc8e0fde5f424
z2f2d9a8ba3df8d6f308d814f4ba2fd59d1f9233706e2731163e0b8225abc66fc9eb8e5a48d8c6c
z85138f96b35176a11f87252c6437d8c4df8a4b96995d15f2c2dd77239c6d262ea55e6ea6ef55ac
z7bb02e4acc2b174788be2d867bd71b7aadd052aff43ef2b0379c168ea4163697749c65eca692c9
za84a7ce062290a5d2c8caecbff69498666bb2e11acaa4bbab391e59a3de5d7a58fd3ffa9db69f1
z869ef47a19e30fe48df427ad47d876ed433c7a5057d045a1a15124bfde09a68b7afdbb62e9b58f
zc5085bb90478b787fc36d8fea6790f5a9881bede492f649644518fefc5c4c678739c028d1d60ef
z38d5c8659dcd542f0e3a21d8f0229c8dd223f45308a3256de1e50908101c8f08d1f9ca10aec203
z2a77f6e43f2b10a881a665cbd7e4df57abe83aea0dfd9bfac159bb504b15ed14d46a4ec0dd08cb
z15aa21e8f942fa7a94b4076637dfc0f06a67b28ca398245904b299d0230be6e8a0c64bcebcf874
z51523bf42d24a957fa98a23d4474e05fde4c46b3c26ef9c13a24f5037d31dab102f644e8204f3a
zd661e6c3a1393c84acd5db916a1c9da328990f9f432bcbb31022c9ea62d159bf5755cde966e42b
z0050e4455670246df333e128504b86976e17ca2b617dd93cdf47db441c79d363bb0335a12e1b43
z9ba92cd6e4975c7ddaeed17ed30cc22b8f4cbb8453b0a7192687b0e8fabc4f50aa7d7b1384e257
zb293332bded3573ab678973f77daf48dcf4460d20cc192fafb3145612ac5179b43323d9c3e326e
z32d335478b64d4296afd2700a80aada493218c377637fb7b8816cc99f16597ea953385b86572dd
z2d513d5efa79a7d501df88f91557a0af65cf6d209599094374461fefc947786a429ecfcd80ae5c
z7d87442644f4d3ea5a420fa9bc3a7d4d8e13275bce53337585c084fcf61dd000cb875d6d72b6d5
zbdf247db873abff80b89f908c4f20860c7e486129e2cf2ffc6775c5569129b876e94a5ce8915b7
zdb5f4289ee396a9cf9ba094594d9dd1729be71de5d2e29fcbc11bec90eb3b3c4eab236710a87b4
z2d06fa32aa03f3e6d0ffe4dbc240707ed0c567020eb91841ae675ca602416d008e2759328de9c1
z079958785ddc549d2c238d2e78dd74eebb763c484bec381e9092e7f37e8381960c5dbea0260d48
z81fefcda11bc0157b9d89f2fd61b568ac666ef59a0a7f5a28cfd82491f4d1f8964c6ab5775e406
z33c3f9b178946dc1f4a36af21a4a8ecf4ec29653cfb3a4e0304bc6d17a70ee8e32992981f2072d
z64f0c86c32c6cd3d6fb43dc58099b66c930a56c3bdbbbd97fd98cda2e0da5b8687067918146911
zdf71af6f7a06334c05d92d809cdeb164f9fec6d69d5e7b69eee44c0ccb9cd3ae2a8ce8e2d6e943
z79818d8cccebc33092bdff9e95c12419dd72786073601e94e13d1d9dc443fc37eace5883ec31ea
za6233a5dfd522c8e14fdbd180fc831eba05353d643bbe623f10c4eb58715a997be1d7b72ef85ca
z6ff0100673aa79f869376e4a211d1e60fcf861f8a35e61262362126841cfed484487b3e6c22ca2
z9000ae21ec1908f164a97eda96b8ff1a54b53779385e535688a716e61f4716c3b06868097d787d
zef32fe2ca8430a1c7bb03e4fc7986e2d3ec456368877f52d5b915ab1210c613e16d114c175a8de
zc72ba8d9650226ab887e5211b96aea8fea2ed63b08584d8bb4e9b92ca613776488062eb3c31976
zd96097967e05a3f7fdd01bdfdb9dbe1a0ee7170bdfbcac4770969edce5f01a739f0ff9cf2d3e35
zcea5e6415195a1668ccb9d35768db4bd6da1cda03f548524e2d7ae7ff5816abaf83b62ec40d015
zef12b41701a04d51b5c8a6c97b6bbbaf63cd475824219e1c9cdc7ffce2602cd39b90de95cf0148
z4d4c0630f5a94f696c1d4aabd6d835913818471d90abcf39583ce2932ce2deb438b5bd28c755d6
z713fb6624ecac80b0043a01e8b531381ba602983329771c033e7d37d931380d09878e77f451d13
zc6cb92359960919baa29fa7f2909c8f0f15201b0fb1b5b768707982b03fbaf7fafb0f8cffe5399
zf95e7b21b5d40cc244f028298fade399b4f4ea53195723b37a822e955db812ad147a81f3540727
ze3e0bd687b5652c3b9db86273e2a3995d5a1df92596da2305b32ffcb414765ce8537bdcef9800f
z69fafc0f39fd4acd63c7571c23feaea5e5528399746d5e9bd7a849d16d9185acd496dadf6db4b5
zf9a744015ca08d92c5089f01518dc1a63d1d1a81b28bf7f182fbc6fd00357110cffb6c3d9dd47d
zd739a41ab838406ec4853b79e23a3ba9ddb080fb63c4cbd4e963cccdeb5b20ee05701a613ef6ea
z8ee7dcbdae40dc73b83eb471936f9aead3323e67a1ffd83e50de9510c7231e7e70883e89167919
z40258fb8d6d084cc1329008e5ada049e02e9d279ef56b9bfd422588f713220a82ec75b26f136ef
zb2952f351b52ec2e831755ae572719dbc7bad85a5bc64937b2873a79e6f953b66aabde43dd1451
ze761361f8620fe84fbe1f48bff31ae0eff1cc0c2ea36521ba9b5cddb13594ec151ceb577264c20
z5ec9a8350ad8e7dd77163abe451b7ec9944f68092b4c5abe308b2e616dfa692ce592af29f99011
z4a43211b57cdc2c940bd6493e940754a3bb5331478d8f5d54dc84c31d4eb936134f5e3553b9965
z6fe1f27f7c997572c01bee308ea12ece244c74ffdc96933b11e5acd9a1dd4e38de32d87c321efa
z5ec146b233da082a0f2e110348bc9a21e57c84ca5afaba4d1e2cef295398c65f2b502fbfb475ad
zb89b6bd2deaa35fe8940b6b6855150806a65d36b7fc98e5a16ce3904349a196e230cf1175e4bde
za0f38d1d7d1f1c85a1c98eb7a2b4155a91abf360fd6c2cb0898e6e3438c254bc57230006f7f747
z9e2c3bf2edc30cf99e418ae9545a1e9d9659aafc012e7e76dd2a5291782d38ebbf189f123267f2
ze1692f1ad33a422415e48d42b4bb9fe543034374b3c0a0192586ff7758bddf81bfbe9d94ee79be
zeff397533c1b669c66c2c76133e50225ed7583cc21b4df0de8f2b25e870848a91d10ef738a7051
z5bad38a64ddbfcc6b90f59ed05178a0b12280a89cd38e10199677055781899e91ef935804ccca3
z8f60a131682c13d9f1e5e8d621c882da9bda17298be43e0998b4f4e800d7c7ae8aee9a573658ac
z75c22eee48e7a1ca880099e4fa6023b9dc4a78ff11d41c5ec1183f7b08f546db0d60900010f9ec
zc27b304d17ef670e56ee748748d5483b8efc607fb9f22dcb5aebce061965e6fe93faf04b89e3a0
ze879b89a17861ded399170035690ed057eb422c5ce3392ba7069c61a72c55b4c2284981a683caa
zae5e189bc55d9cca60f8d4f7e1c3f8723267afd3e9e4d38feb24b26ab56f0441132d4d4c61dd5c
z5662c63261ad628336f510a2dd7b2936f54c6023734129cec173a3aeac63ab80647bb519de05e4
z1cb74c0308d5066df77216fd18d63d65eaf0b2a5b7b0a803f08c0eccdc879aeea4f94d2e3f643a
z69667a6acce5f0a849cdf0fe99791f06d80ed253e70422910c1bea2f1de10802892a7302920cce
z4b5c14e06661161c00f91a063fdb69ce8314c6cec59c34f7df54896a6c2fefb0b4b48e5accb65b
zd3fe2e19e86c2100f3d07f63d72dfecb1afa169790f5d1dfbce959b3d23b8570ac4444a9951ec2
z275afc18a63d2cd2af6f6019c0750bdc01f63f94b46963425c7f9c9e1b9411f8f28c32e5e15c57
z20abafd9dcc000c91df2ffb9612f8022aeeb0f14027a685f49d9d4872c16136970b3823421ff2c
z661bf4c422a5a30dfab5e55a4c1f14ee1e6ce0ee73ae48ec7bd86fa116acd3a84994f650141405
z7fc2caf85faf1fdfc37f85088134ba2ae1389ea86fd7dcdd50cda9c0e2e1565b1daa0ea6501ce3
z3b531c30a596240f0f05adfc604a7edeb099df0115f9d6dbc270658d8b9bcf72aa321b802203e2
z82469fba012bc32c33fbbeb48470e7dbd6524800fb9ca7682596c8bf33c4d2d90db8e31b1e81e2
zc2d972eda23af8da528322565e284530e79bce50051a09cf6e3682b590bf92e37f44f4fa4b245c
ze46efe805a40b6d97769befb06a4777aa1f27cdb93287165366747742266abdd304bbf26a5948c
z64bcecf4b332659d005e4bd944c66505203842e7fe28118b9f60fbf63c9ed7dd43e81d1ad0d904
z6df95a0cade773d0b5641b4ae26cfd5d710d7ecfef4870e78f84f5bf24c9fd7e890e37c16582d8
za08a9bb3194d453731901557169491e5e86d09e88f774ef72b57401f4fb559ab67c66ada50827e
za2113bd9e0320d2a810087bccdecfd3a37b48c87f1aab56a7dc30b869b2d0c2bfa8aac4bb8ecbf
z9b835a032d320e27f07219e4f5b807fb28eb8d726dfd0544c40ddbfba3bd9f038a7656ab477252
zfb23561d678b8b8da46b22c6c26e823274976c7102eed86d13f26c9d24cea6ecb27bb223c21279
zd5d44988db19f31eedb35cce4871bb8a707c7aa8ff90c71601ef98ecd697f094c5c7534a4b389b
z85899284be3401a0061144478309dfad99bf03c1b7fe322c29b12f83118c6ab255dd20a5d6e81a
z99b41c84a1a6ef30d1fd1ab816b2afc79ac0b203aca19a50838d643f31b21b07418414409b9973
z42d86e5784cd8285f2eafb7ab50e34f78575da4d2e92574575cb0b9f613e3057c99310818dcd72
zcc3b551974b274e5563a5575d5e32f289330af2b0d66912761bfa009addd3991d65b1d1fb82386
za571b77033d6fd1aece0073ee07f2a0bb9aaa8965d9e6fb899306d8a31221e9ba04a2e75e473b9
z4cdedc364fbac3be90163fe15a74a02356999d12f1bec56d3cacc91f9cc69ebf3a2478b45fe9c7
z25acaf37e291ed67353943267af16876be12820197519c95b034818a662d30e3c747502ff5a5cc
z09bc16f3da1a91ee1e1988467e5ec4d07f4f95f9af5ba7ab855feec4fa4bcbe3b930e3f2989ce5
ze661a6300bbdc01ee97d749705907121ac1a3022472cce2a673e9af8f14ba376d9f0ca0b9c3870
zc5abca48a1f93c8b0770714e0054e6e7becb181cc782086a7dede8037d041ba6463748902fe37c
za48b0f7bdebf25bdec3c982ecb8381896dfebaa95331dd19950fc044061fdf2d93e339ef4b0667
zbd444b07aa926761cec96155f7f6abd0c9ec1ca407d7b98d459dfb0495c656bf64f349d8be4884
z81ff8c1214ca6ff1757cd3a7ae29bfaa49a068d31e361effb4c98a5bfb91df0ebefda4fdf2e39d
ze78019d43e37277f6bc200edabbfc97e72c9d9f7ed20d7d15bad0563f666e7c938217ea63e8e94
z20811f544664c55038284ca0f0013f197bb59c80b58f4c68b06e7c2b7dd21318761a8096ad52b1
za1000dcbd64506e17a7774949077367f24a649fbe24dee5bb49714ea15f0f07a81343ff66d954f
zd9e9a65e836e32fd269066f7c8205eaf62b818acbd1a1e8b23a48dbceed503a3cf7b20b274b06e
zdeb52c116ca0bd7aa91f9475ed23416c317d63a8e87cc80f44d7e645c4a7569df8e47d9e0ccff7
z44d6d5d1ae74c6c6428dea71fd730e2c58cb4cb94d9801ec5848edadfa72b2989af0cf7249d7f9
z5173ccd23d81ec3c6a6d290e148c90fba65138132c822ce72e20b759fb1e45733a12cc55ab2635
z81cbc49db9277b3c3ec899ecf27f0c4fb7428258a7a9ecb8779decbc6d1bc662cdbcca3edbeab6
z9b194bc670ee7adc31b4ff91592d1a97129f00e979be22387e2bad77af8b2fcf3322f71184c260
zab6ef15f7ba42f25daf55619124cda483210dc3181e75ae666dfe0a5805ccebb1586e6d16a39fa
zcdd83c7461b146888e85b4a2ac770b08065210b8a71cc6fb9a7160f4abbcd08e1f18dc10f279d4
z62bf784549add006594e475ae4c7955736de29e335bb2457fe8ec9252a166ef662e6a7db59f979
z2346868277be0e7a38f64d79fc0178c99a8bca5a1d27d1075fa59e7a26104e45e955a86727355d
zd2eb5946e6ba47bed7dce9d2bf020635e310896b254065cbd600a40177a747923c3aab9cde17e8
ze62f26bcf07211972af384fbe5dfa472eb1ff1f44bd46583a543d8e1eeef2cdc649e8a10799593
zbca26d77c1ddc9bcae3f4765e907327c089850ac33724df08803953bf517dd2ee1fa7e2f3a5913
zcaa3b5e06e10f15783d0925762925c03fe6fe693d22ade1323d12d214a70f20d67ae9e48740acd
z9a5e926add137d0d2cca9aed3871318531b815d66a27c19b8eb8904e3362f3082215984fa1dc81
z8f9e6400e2cbe794c87bb645f96273b902c9fc18adb80fd72522efea2053015fe3c6b452a3a9b7
z10d64101be047b1f472f185aa8741c1450eca4ef1540838ee180ff942eb0a727b822ef4e71314e
z64db4777d4f9ffca2742297de4656b043fe41af9634780d52c781d0af083bd2d0e31bdadc51932
z361d3999b3b9972b90359fc76bdce722cfdf5a7a475c97749ed9296b2548f499874d2916bf85cb
z3d13012f66c05dc82594c7f29661bc61b9c553a6473ad83734c6c3899b7e5fbc33ab1e8785c1f6
z2161974840a8853794475a78e0869542ad5a5d7fb62a256e196e4d12c038e6181f409d69934ee6
z30a9a9083d8aa7473f36b5eb51a6bac32d56211721c653056e015d22ea72d1dd169050ad6ca0da
z0d5d12818a757c71f5a2280e685bbf35ab567a11eab310d0771dc5f57c96e2e743c48f3e86ee93
z07c07c10efd51bdbbb97f9db26b9755e5490b9db0f2212be502faa77b83c870a00e81b4b25bd37
z12473ca4b715060307c23f3aad6cd7d0b742905fe7ec61afe85302a8c80f263d8796e6503b816d
za8685b3e049194d3fdf5c2082e483407d06f1dda57163163867585bad9f6b674e8896796817f75
z57b67b688209fd6f24e5c3b9323e258c75a7153677c71410f4f07a51e1b2bdbf4913cb6efdbce5
z13df7c523e778910dbbfbdd47e07f1ef6eb1b051dcafe4701e10613d75466e2b22624dae0f51aa
z50a97e149dd70dc071a08ab4321ab43d243559345d06077d7b2e2c1ec9035345f5c7570ab363c0
z32b0face3692217e05df7b21c933eb1a33e3742d8cd0a4ce5669c9031dec11a3efae94d1e016fa
ze733e4233d0f059a86c8f7b7dd9a87fc7a9759ad7e3f99c266ce9ff93af9392ed8a23664a1d4b1
z3e2d0fb23452bcdea6611897f66b7e310f8bd3a0ecb10c08967f834f372e7ae634b5f1590bc145
zba8b22fdce927979668f3ed7844fe432a994ef76ff188f76c80fcf602534e65c716da4f419914b
z1b7f94e0b4bcf76191352bfb450b023e1dd2e5dc38ad94f7e2420d1314d529c59549d0750597ff
z2aaeece1fda9f68eebbf5ba803fe741d370d57e7c13c6909faf9e33fd0fc9f2453cf50ec7810c8
z7f541ac09f9f63fe86d3f74d22c9d2be031d2fbf482d602d30960a69640e8055f0d452e3106abf
z5997b90016f162f345fa0b2f7457876e76c888c24862d2adf47fdafe38cb54ebdd808259b73faf
zf642fa9e77c9aa8fd12d1aba7509307f978fd465dd56452cf9e116e4f2c42924f57a0ff14bac8d
z2156ef49681ae62e63a6896d3c27f6e0dec11b78a9f6387409b7378884063f3fae4a30395596d4
zde225260e1cd3a4b9559d2207eb0e5cef3c54a01a88a69d36de70d4aef358b4042fd52de3b994b
z07bc480c06076fe29e8a9d14c13f8736dcf14e8bf9fb47b5ad67e916fd4f3b5824ea22a2ea4303
z872292c4b3bd265ac5aaadfd783ef1114441d4908ebfcab2b228b16be7c378ef6af2d81bdd4fd0
zcdd53c7a11c28dbe6107c0a29871e710d2493cbb091af356545a70d769bf1459ed21fcd257f9f7
zeeee4887d31e409fd5358ca2f9f3168affffc1f8e9892dd492a3d05f25878930e5c2760b7062e2
ze7867b79efc92e6000d580495375dc71ce8541f5f1379b3a35a3c73c51895c867337e26f2d4ac0
z6f3e43e1c6dbce378b2f29498fb8341bd2d403986790081daeb9562797a9cb70b3b23945c8dcd7
z6752177ed0353234d72ab03d5672c58d7313f0c81d07d9ad14a3a0fd62495d5333419e7ec8cebf
z842f2ea34abddd65c4e0fdfd8228d53a398a6c6917698be5ca06f7e9e212b4c608c4eaf47ab407
z5e50a0f1666a2e7b569cc0fbf2e4a8bb0f636fa8e4899af11f3b0a53166b01d91b388563402f78
z8656bea9ef9edac37c0a3357c82131dbb4dcd92dc4457f60613fd263f729b621305ee6c428f386
z9371856b379bd3b8a9db6fed0b642af99c522f0bae94d03b548793fd6fdd8e983aa2ef269fd7d6
zf15e319d8add0744aebb29af4ebcb38546de214a1cedf1e4f9087fb8627dd3c11af9d0c8d14e7a
z1ae8cca5630d5d097f83288d2a2d0d4eaf3d88a6c55f4e0d3220885ce024bbe52acb1a0c575a2f
z4f46edd650d6302b1b0584f3ae78d69f0e10c5fd842d7313099133d506eab30c7fe8438b89ce05
z1abab17ae7916d00b1dab151fe55a0a16ed9f3801bef0e6c99ef8c77fcdfaab22a86af26733d3e
zd234bebf083533efe60b1fe8925357f3cb4fd324341900a087c6ca4e4a88b9dd094d07a09f6499
z585230663c8cbb42027620c0082b13569cd619e1f71f0abc8ea3b685498d68cddba60ae414f329
zd436fc5616c8284ab5ac23cc5613d442e493787090851f66e2571f0bee51f7b2eb40495aca074b
z1b04f13f498797f2b709d9569864f64f5f44aba364f04d22f4417391c96f8e7b189cc65ecbe616
zf05c1669177ac2cc7a9da5c8ab98436ac025c84baced013defd6b77565ba9855504b85fa91cf88
z2ae880f6684957c6e33f2d11a5b45449b6a848f9212f2e56c86cf0e9db7b5065a3db403b86ffc3
z74c75dd22b548ab693cbf86f709ab4a49aa25587b291c90ad946a30d218d30d9b4b99009eca6d6
z318b76c617d6a4f6e2297acdeed90f3751539d77b479603bbbec4728245f3cdd1b6b16278128a0
z191fc074a3a45c1e1ad54f1ab3def60f8b4011fb28120005ca4e958f7d36236540a054fef026e3
zdf3e32f0cd5ebea6d71dc5f4d418f6893a479129205e8282616d2fdaef4caea0faf094d980d29e
z6e681881da0e30caa2e5786a850833d6b16f79aabd91da4d36e2fa4196c3151ab5f82359bbfab8
z6d9691408b90fd8a88c20ee3cfe2e27dff874c21ab030167e895fcd0660c3700fc36b60e5ca3a5
z772e9f983f831c7f22aa9ac3370f4abc8236de0c6c76787e4a288941b19ab3f8f61913815d7346
z5955934efb06693b1a937ede4ea875548337cf5c346cbe8059eaa061f2e6a60dc980664d243032
z2bd4de14c5a38a8d3bcf5c5bb80f691862c422512ad6f912d7afe5f123499e66aab7bb87d58d56
z079fa17241d23b81534ea8f7a9357f7578d78b9cfc34a0e187c5110a2776f8c1fff9c292207550
z3cbfb4684363cd69bbf833be7c6c62bfb8926c809284abe42db02dce7fc7ef747acefff8bab25e
z5bb2358e20d4592240bf78bfb5af8010db96beebe637a95078e1d994ce7c4ee66fec1c17eec4e6
zecdac59b1296b9a3f79b555cf4f31435855bee09733222e270d378a3397d272a96e6c67f487179
zdd0e0b694f655e1b151dbc5c989cab3211363051d40498b24a014ae84dfde86372369f5b5ab770
z444825526145bf7d94cb61dafae14e2ef63bc1d2a0b272f976ebbfe645e325dcc811b9680b241f
z9f887c1536f46351c40f95017d3bbea948118148274bf8870c0620a6e0379875e8c3614ce0772d
ze7f6be9cf5ab9b64ce03c72c465a64432338a31a183a7e22000b2698f5a6a0cd2ecacfdb6dc5af
z1e726a9adab68c5291d94ad87bd7abd7c2ac45f56ece33f36ce83a88a44c4a0a228ae890208473
zf518279b4fd51fa0ed3950429358cc88ed5256d2db08c96fbd3b15c78d22ad44b41d455c5efb3c
z4348e1f3a0217b0a8453ca89b3f44874ef905352818e442a1fff1200a6c5a11d78080687f00c97
z10f15e8261742562fb3e2660841e905474549aae8c9da7a6b8698815c986585da8df3d83ac728c
z18e22e5cc54afadb9785e6b8422665f9cf1bcaaa53a6340c908bd67a1bc2a2f3ca3ec6edb6a91e
z6de1e8511391aa60d568d7e58c3d43e2957281ec76beac41d7c9a747da54ab39fc3fd96fe0afde
z3857a0e9039f8dd1fee09f5e3ab39cf6291b104dbf26e23b3ba6ba94a5655c4f5155311c0d3129
z29cf37a17ec416d407c61860f78361041b7c0839675e5bdc442cc233713e681cfe8995ef5d1ca4
z7a019bd4cb26ce3e9dd2ea4b5094c3a6f483aec87c817d8bb539d0ef225bb7af4092068a60b6f7
z83ec95cfd2c4c315cd79e335cfef6dbb004fa005dd9a69d11d0be75849b1c3c21efa7e629f694d
za2bd942f834fea579b3b343f82b5d93a1861e648ee10700e08591002a9abf73012169e36973ec5
z47d1c4af13ab46665af3b3461f405f4b51fdafc9f6b76f369a060fbaa5f3acc830e7bb7b660f27
z48e40a170b1c6836fa7b9c4b5bf463bd7e10b993f29d07e22d0f9bd6a595e1c31bd970e85e7f31
za9cb6637a744215d513b943cc383955881094a2c46faf332f97f5d1d32bb3f94b8cc79f8255b86
z3ce0c1dd56802ede941f2dd556e4b3d499f41664a3fc10c4098da05a1f3a0abac348f152320e34
zacb36a372130383e76253bfe6c6bb86a460a426dcc65159ade7f62daa2d769bef067610411c116
z65d3b04335957b964b5a8dcab24470635fa2459bd2e13860fb1f08ed8ee5dfc081532abb0297b4
z280c07f37ae1d9b7176ab8f0a6b24f6f394bd85e2eccfba3a70ba6150fb824b82f8ce7cfc5f3de
zf215c63b2c99190b7c59ab3f960dbf761154efec245ff95ee53517835c695222359201b110aa8e
zdc8c730b9996faf81417d4fc39640a9ca7a85acf0c9d52a478eb0ef442e8ce2d25862c64ca5b88
z9e3d8471aa9faddeb5c70efb9960bcb52f1d5b7ed1030550b47e5d599955031d54ed604548eac2
ze4302e09a66a8e7998411cf8c02c0e61ad61b33f79cdf4c7dbacfec93a0889599be8359d570d3b
zfec235a3d53c754cf3603b9e88c6f8cdfbbcb760f3ea87380bc81dc644655936f3604a62a1f0d0
z8d7c7e831baf804865e48644d99639eeb413bb06dfa06b3cbe9af3d8565b2a66d728ae2c4ee8aa
zf51a3164c31ed7f278963ec42afe78e0dda3240b0b606e44e72bc0b901a1ebaabc496c6fdf47cc
z5b716b0dda3155cf905a637a747407d500729774c1e41643f459b8577349fad8a5a76b9ab69356
ze112119f1236872f57b64c7abe60bfe441a50395b012b0e109460a82d5755c30eb671401943386
zf8922b618562bdca8a4dbd52a33d87ee59c3da5d98a293646b8b34bc9e3235cfde4f09ff661619
zca331d54b7cb7a573a7a34ac8bb9eb66c1d4adc026ad805663035ab323d22c0609f94537b89f5b
zb0a24572ae47f58b37ba23ec2f462406fcff35d9f0639df9fa320365eb9487ed83986b5074b6dc
z506edb1df9235d0c488ef3d142ebbf1260766d9595868f0c4ce7264d3007a9b5b946825803e371
z0cf34f6a53a6d516024debcdabf0463fe092799a6a12f6af2767a8d461039f5053fd868071fab0
z1103066ab744bfa6de9d1e63baff3419a05319a4e601aa8663402374257687e56bb8abbcf1dc3d
zf77fc84c237a467193ec191997ca4644c03bf5cfc12a7c7794bc18eb68fd8aecd25b66386ebfff
z9ff9a23312276cbe1b39573afe6929a274f5196a2a0f492d2fc9cdff510cf94c199d170c185237
z787cc37d655e4ac8bde41653e467f821f74c0cb4419c8cc909122ec422bb41c3d209b692047b1d
z666cd2d34226b66648b3b2187bdcde27a5cc31be1da95f93d99bd927faae902b5a6002b72dcc4b
z50cc82deb60bedd7783eb8b8e2246bca912c50f8aaa791031e8370e2191f8b7b5e3362a494a76a
z7899c0a2074f28556fa5d74b0955ea930a9c7821ea9549b98d1e71ca1b8826180b431086f3f1ee
z1def9f664dc1369608b2a9d9eed6942eca7a5d5a72cd3c61eb996e50245f4bc6e8147a576189f5
z45ce5c83e121eb6a9a5b16069d427bb0c6720d008e8ce8d963edc4c41aa46c76210d09866fee39
zde420eb47a4cfa598830e5f91c322dc769a022c09b0faeabed8f193d92a578f824931bdde02f90
zce19d10fd5875f90152b984a9a25375a7ca65f1c1306e2046a94c6deb1870df2c3e5d33a168168
za00c36340cfbd9ff14a96c6abc6bd44fbad2fa56b8d0c2c95bacbb862c7a67bd2a650a9f65e592
zcc5b63c338ccdd52190953886276cb702ed411bfce7f4819e419adbd2119488236317d35f8f8b3
zfa3e248719e1893fec6173f969465a2be42ae4aa99dfeffb177e577466a76371844ac0d45bbf12
z70786d568a458dbae136448f1219cf113e85cc80676c59d296f1068a1c508f389ce9b8ab52943c
z81a24e19577d08ff7ee381a89fedb8d4f34b914d8b74f67783c5bae05ab44e7f96dd7ae7bc0776
z63377b83fd514ab236a347e2e863cb1bb345a1d02e0e90b9d994df8ad36a14eb8a410ef85d562d
zb8f8c1de91526237b3d1dbb56d8e0b9a2d96baf6b19d74fea723e663bd78aa0f9c0dc1e1a6ddbd
za4475a6cdde4466339e882b7c1ed68daf1c2718ab6108176dd454f84c8ab4499be603276cf9a30
zc9cf6236f36cba9f7dbc9f6958f99eda9fa3da0f0f9d43d923f6459b81707b7713aa2df4794a19
z2a6c7d68ec7652cc148a9705cca9df5d478e4a13e62e4d1e9ed85e8a5b1091ccfc727bd8b9f551
zfe00c92279c3cba3c0453f428dfc965cd2f153fd1612e94814da3813ab0a9d715120c57bbc4790
z6047d48efdc7090ef72a182a159a1c8695acbd88d9c19f723bd6caed229b4511523b0f729246c0
zcb67f827da8e78071db551640df90b0ef2d85c7bd9a0fb90abea01cec263a4f108b905a479fac2
zaec2bcc5954808306f4541edcfcb5f0711b7d6e82a9fdf8572f02591fcc7e9ee10ce3bc307bf22
z70a735c0e3d2575f652e4012740e3950a48ef4734e18ca06fcd71bd519c5e14c5e5f6e08943f5f
z158c94da5b8033b96fae8572794f50572cc663bcac0af95ca7f9046fe21f05a25df1ca8f371edf
z1acca05e45555be86ef8786d4a250363671962d823c67963cfc45534273ac7fed9c3d9bd5a1c64
z6bcb1a8ff7d62904c2649abab41edc6d18779e3a9f3f37a3db6a10d490c817647299e473306e7c
z68af5aa91e295b99aaa7ec1da15a70b76960d086b7f0e320e745ee0960aa97abcea723f7b1aef6
zef1be896fb80bce8fbedebdec831dacd61b46a192a6e9145b2f36e7f24e70772cb41597264cec1
z7c624715b9c807ce545390bf751d8865516e879a823140c407ef77bab0325a00e60d0693b7fcaa
z6876e5ab0898b8f16bea776906dd69dc33674b4053f396484b23f08c0b5177d6a4ff5a042ddd69
z68d2a8b1485f902032a5c832cd8d2930ee63565edaae3932f66f6e9096e8e8621615f41798b4fa
zc17d04294e3b58a378cd1f74ad2576f57bf92e637fb21752cd7ec0b2b410d1d2054af2303a2368
za103e7781bc90172a11a65d75a1fd9e96104e2c1e33baafd83972b61d09702d59a248bea58a658
z6d66a19c43bbdcd80f7f1324a1136f2402bad20cf8ec0e3db2bbf3dcd4b33c93eb066f3e602989
zf2c8db42a047bf10c4e4a384e8d325116595191bcc5feefba06b268f45292ecf0bc9c2b1ce7e9d
za5f3ec6cc30df19b8e9b5c2e02193ba322a56a84e3318cbb629e412c9ea57c5ac3bfb841e8768f
zf510ce8b1c1f3a6fdae6b5987604c3296c2c47eb0332a9bf2518ca7610c4b7fdccdd8838a0d669
zeb8e11c63551ab9045cce39d69eac241706db42809d34dbfa6b02fe25f0b34aab2d8c0e4c53adc
z1a8d04bbbd1f05a209c129fc5e4cf78ee2cf2f9ce2f39eacbfc588dec709a8e406c4ce89fb7e22
zeb27652e113f1d2d95e457bb69ad323447b5ac127a5aa16c4ea3f04732fe595c8bf4abbdc817db
z544f5d23e3abf24fefbec0404f48a49845c5a211975bc3c84b7b1ada5f6bc7b77f4e985c3a3738
zb7f17056084946d669139afb5374313ef8054141bff97e451ebd367cc379a5fee864aa1c3fe983
za35b0a787e9aaaa90967e4d2152bcd6c1c9cbce97d90cf54d28b7c8afc3f524528d2c43f7fdeef
z26a36655d420d625a3f116e096f564038c5b9bb1976e6346e6fa59b26b922713b51d413e47efc7
zffa53a53ce0f08686dd4d16f5e922ba55a641e9e007b199152378d8adaf53ee939491bb1e8a0e0
z56830d0ce5a250f41bd3da6af3e7ab8843f653c9e57f6f933e638c6e44b2b21fc8c89951bf9d10
zea3ff7003432a04a437e59523c91a77256ecbef9b7b3837fb71f7e49e3de312494dcaffd064287
z9ee136d2b50918253f460ffc8ad0a1f476beb93ef52ff4d22f65e4eda5dc328e662fcff11b7aed
z0e17dff4d8345d05bd5cccb7a51d0b1a766fe80cc1dc2d3d6a3719ff950cfd5e4a452bb606aed0
zb9ff8e9894007ce3d261580fd25682e057710b083c4343240a6a571ca828dfd396d8246e73f2be
z1df7db4863e0f0c0642fd7d90730be42cd649e3e4097b99f00a419ec97a0eb0a3e2674fcd2d767
z4e74c91bec2aef75daf9782fbe89ffc6b067673dc8078960b1d490d86fb9e6c750b80ec5d81bee
ze551aad9584782818f03ba568277c3b651b83c02c9b755deb272915cf9874ef9787fecf6a49e30
z47ba1ed6d9778d6078726fec17a70631f89f9327c5c87bd234efa12ef0a3d79577f25a8119e44e
z5b67487ac7607cd693179fcff7b8de3b6575db4945f0039314ba28c522a014fc83f1874ef55b80
zfcc49d6c32a5be99120bcdbec47502415c071311e28647e4386d3a66c93a7a959681569fdb6847
z466d721030a3ef044eae1fd2e338c232df014d26801ccff2c3800e94d51b230b55632c496e971d
z3b1b84298245643e79deb2a7d041a0fc54c15dcc23e33af0231608bd7adaa877e90580d91e87f0
z32c12945201383b53e397a8c059c951b61343817c1b4b7f8d80b9ec9659a8f102842a5c6f8104b
z029d5442f0b1a03f633aeb39680e0c33a54be11014a3c4bc58b31d4aea35fb508cc190a22817cd
z0da92542a56d002479ea0f4ff43d0927bcc13876b29700c9b6ee3f1ef1dd467bfd5c35d4bec419
z54ff2e0ba85c298dfe6f178bbd378784d31cc4b72926f2d2e67f08ce171de008efb8a6a5d54ead
zb73a279553b13f5126048cb1bd2b7936df0df3d5d9fcd88e41c9ab6e887d68bc00ae84242c90aa
z31673a79c6ff7b708e6206190c1a48cacfc3b1353af5c38d8a7e065e8c6d0846df6fd7a713345b
zb18805d75e6a43393a97344b5734214b3d50cd4246667c5d03c46ee5ebc0aa1688cb105ccec2fb
zab7f5798b6c1c4fb3f5cad9d395a161b3ea96ba09229f55c12255a73c60398557343f8115cdb75
z79414ea64a13f85da011560dbb19e7d5ea045aae11754976c22884446f383590c4e4c19afbe4b7
zbfdb352dc09397bb3dfef53bdc063505a93a2b1f8109a94bd4c1b7a193ebbcf53873300607d05e
za5469f26ebe48b9fb3992f62bc6d8b6bbffeca47ea6580d996cdf0e3e24506c8ac708dd612536b
z38b493013516a3f2b8ca89fe2d7cb77e2a720070e3c0ed72bb5435cbaeac8dedc7bd39bf8c44f6
zc76581bd44a0b424ae9d82cefa84301c2b872242c4ea558668ce56fa514890f17e95bb4c3ab6d3
z32bb7314c980bf8e2988440da8d4148247b7f4bf9cb647092de3d9dd7a60d4bbc33a2462227db0
z928f8e8a1e545c355bf1db39e9430b0a7e51584fc0d5b7549f9fc081dff837a1c76fe2cf232374
zfd6f795d7630de30f16330dd4f9bf60f732b81d50bd0ce1de86891f56f59e469a7b4cca2538327
z9fe51cd44123a311f3623584d6e396559d3b91b512d799c190027e4798a32e5b44ed3db7f463dc
zb239650513917e21dd4d9dae063089ecadbe61e127916ee52b1a3a2ffe3663fb828891b56ffb58
z4e17d2598940815ea50ca24e4852cb0ca6963e900252338255fd23b17b86061ec2ed0b7c0942e1
z6e49311a7c625ccdd61e0955253f57c1b7bd8a1a08ce448e073ff51efdd690feed26704ed20395
z880a62a1bd9bd56d03cf924b11b46617654eab3dc552dedc7b0c0852d67eada74447c40895d383
zca3c67e330cf4b70330c89dcccdf844fde1053a6ee4a80a93c67eb50a3dc9d49d74dba51f969ba
z87a998f380820da533fcefcdbcda5960639b140b7c5efe90f9838cf865d521ef19f81141ca773c
z10fd000415289fdd973d3f951898fe21e290009ee7bd5ff3688cafad935553629de460dfdf0902
z853153e03bf245f479d8f9daae9509c75d74b4821d73c29d8eaaa5693e5342e02dc46d7369f9ea
z27733ed495393c00cf7cff183a43d509c2bc58b3da415309a3c5a7ebf5b2d6bb46713d2849dc63
zf63304380916b2d2e2e2e737caec1e00aa2b9161dc5fae342d807ab54e6ea619719ed4610ab74c
z7772af50038e57cbe9a9f74b735a6978a58a363de0cedeb460f33ea927449af17017fc359bc6e0
z6a814c2bfbfa1dab91cb1f01e1ece4c2cf9fccdb457aeeebc93ff7b9cf46ddb26584c728d408fa
z216a90b09d163a9ad3435fdfcbdee604305005d3f857823725a2823095333021f989a4e0b44dc7
z5ac375f4c5669bb0499e042c2ecbf6213bd09254222f4e78ba56fa993f5faf3a33983100f10684
z6861c4bb644baf9dfc9bf6b96dade6fe5de04a5c34a116db30f6c945f9ac6d876a3a6e4d02151c
za4038ab0e6dffbdfd23586700ab010c5c2de20de554443a44f3eb8e5aec2aab31162f236803229
z385467b1f0acf4b4c3e96cc148f3a5876e436dfbe17a6548b154d6bbad5a1a31c88a887119fc13
zcc7a2175759bceb62f772c2d1960fe3787f5d798dc856ba79eb8694a9337a5e72e22f82d0ab220
z075eac107569480b9aff2c773cccb13300cdfc71580725b734470fbba92c732c40ed263719ac06
zc464e8ab89a144cc46979aaca73b5afce39ce58cc6be6bf5d248fd94af9f1835182db996fd5a7a
za103a53d410dcec702c943ce7316e2c4615c0dfa06051a0b8eec493569ffa348090bc83fa39a17
zec4505766c05faef1358627382f730e8695431b7cbd38475edb3bad45f48591b08805e143c68c3
z8856b7a55501a0fbb610f1824d6f828504e1a13c1f2526558179dd6c302585b4542db135d3c916
z48322456137d1f225080eb4541e3f80cbd95d5d09be5a23f4e0290b5d744b65ec74882dbfe3b42
z7de4b86e3bf0bbfc4cfa3de3cd15a9592b0527fa2bec7dab639d4c72aaf6ba007a65361671055d
zb8d931fb6d4cc4534838590948c0f8a624f24fa7e47794ceb61fd76fc442469aaf4285d11111f4
z438989f1e33cca492d603d450f3a5e6670223a443a8578446fe30d3bf9ca5de5ee0c562ee35e9c
z605d53bbd3b25ac7d5c7c69b50280d7502e44da150e5f4cb6ce51e417708a21f554936719d81cd
z71b8d8eaa407460bd2a731119091c7641e0260f2c9784c6d9146210f1fba8b0fced249b0d8c4bf
zf34f4495029b26263b1e6499e3c3f8bfd00516a68f8cd85482638171670463aa4b3a8e66685479
z8f33723955788f32608255b21391cba82b940dc36a32cb2694a178fd1657a4023142e32db0dba2
z0d2647ef7ec0d73e191b7cdfccaca720b03a1dfbad13877742f8e018057528a61a1210399b518c
z7ada33b6a8307d058309400a4bab9a3b51c749ba55236a81c3421c9c0ddf21ba88b9bbb199d8f8
z68808d709afd97954511d60b888eba0359d63ef0306710041ccc06d92a31c487b4dddc3dd1c049
z25b88c3e11d06dad34456b76e7ec5282d120472f8d52de82751ed439d5ab5a37099b665cad14b4
z4c22f6c2b2e19e946c0511cfc99b226472e5c5dc28670b4a7c4f66e93c5a8680a858ee2b844e2e
z8377749a5e0150a6f41247e5c914ffdaec466682a0a579cb184b2b7b3d17bfe95713c47da5ede9
z6d9f4817476a54476facb5c5e87bd8e2e10ba5262abe87a0444f5ad753e4505f4166ff235a1e34
zb08fffa179f8813a838f1652d092975add5e346c62c3f3d47435d266bf4c0fca24b475bca5416e
z83877927d29f09083f9c6d78235ea6be0dbb9dcfe07d23865b77760d34fca45588d3455fd76d4f
z70fabbc51c124385cec946b32faee96228b72c65cb08b5df77bf997e24f9c49f52dd0dee2be5e7
zd3925b42e42321fc5537c05edff5b4103f6d6fdb2c7e4f670f2346c2b7aa33b48d4439740e3056
z7f0018a12d98b2d3c7e92e48b85d757019ca76ed577de486f43763f50fa6f7610419a0429a2c41
zda1723ed14402ec1fbc8c03e6a325c9fc9b4c16c62858a0d1b8785b1184fd5e36cc7064e210fa0
zbd3be3705ea6b6b412cf3e38b81396fe9a565044768ef7b2aa4b353ea3fa95d19f48cac4fc1f26
z5407e282eafc8323d41283f2f66d423d8a503a5f4265e63909285bd6b0f8aa306a7ffbde03b257
z34c869713e6fb18e5686d18c42c7fb58cabb352da64104edbaa826188858ebb20d67a96d7db3e1
zf378699cc078dbe984a2cd8012873cb9a8e10422391b50bba1f37e712e96b5761eb626eba62ba2
z8168bc9dfc6489b3da27e48449373b1694bb4dea7c0d42cfddcef781bd66976c49e20665fa7ad3
z1371bf40a396b8886ebb908bfa64351b5d651eabc5f814fc44ed3d30deeca167c51ca7064fac48
z885ca385f77ad0e1fa8e6a5c61a77c92f13a4ca1a07413333b0f226f71c2fe7a1ba10ae8907410
z3426fe82e7225adcd6f82479efdbff0f74a35c71bb751195947f3837fa33262816557ef6c8997b
z49a0ef161163de36d947abe1e61e995faf82f290d626ced425fdbc24c963b7b8d48100b5224ef1
za7c8d341814d9597f5c5499e78bee9b2f5b37908861f42761e193fa55157ca14c00a11991feac8
zf956f783f26f545710d4070f818d4efc0d7d34afced1c9caadbc869e7fb3e250d2edf392519454
zf52fe16b92524714957b3234ce0e1f6e871138c2e53c92cb579ca46c21ac567b63790e8c755564
z0b1a4e4bd334f50e860e2c8856fcab676c8533fb998c1e1968c1f016984d46b7ab41f1bd30e38e
z5d13b1c4e1e886c11cdf3204840de89c0d460c7d68e5ab45e3ed6aaff6975a786a031d475c4cf5
zcd6c5eca086266afb827de7281dcb315ac1db60a91d985bd45f6b7da7d8f12ab641c3503632801
ze90216f1433217b3b92c324a826a2410df52fcb4e73a310675d340770650aa287f62ab78751abd
ze25dca259b9d42a2a382c731b9b27ba44f7f3595c4ece0920526be68159c4ef82c4b8cfe48fa4c
ze49e5672c55ea7e901404f74e30761c6a53513fd2d76c406ac47b8cb08c3df9345067d60a88c71
zfd3a1da160d86af398402e7c1b14d3e9634bf8c9f315ec5829b6fab07d18cf206ffcf43b1113c0
z2124198ac418a0943c7565d70923f2ca5166eeb4ef823dab4e46e39599546ba77ee84a958e5101
ze88e066c6fab08e670e7fe49b75f58786896aa8d529ab0f1ee9a2f899812d3ec81bdf1324805dc
z4a6240c3837d3496d0e4a5be824859280f480940512ffcc9e0795fcaa65b6c0943499800f07e9c
z32d38f5a80a9eea5c9076355955bc62cf917df427f3569db478e76e0342805b0ab88bae86a7f54
zc7219720f49f5ff8d7d8a63f46b19657cfcc8e9ce4619767d901e205c0c49f9cdce8d5922ef3e4
z8a492037d8cdff75bd403f3fd5fda8fd1a501c8a1d00090af5a8f714fd37f8fe027e19d01488bd
za399b1569f8fdd6577421bf7ffc6ba284e964862ae4d50f58a4a52f24e20e779cb4f24eb54f02a
zd6639538bb07f45f7c17c5a29de823c0c700b73e1e5c4978191f9c73d4acdeff24341812ef2c7c
zbb562848ed211a88926b86e6972e8a47f805960c34486caca5373980c843a3993accc82b6e3bfa
z5199507477d26875e1b5759be289aab954a5319a31d23bac9485475e2037ae2a57174fd8204450
zf5015c2a72ea3aaa39efadf6d48d78dba9a414824cef42890b14345189da98a730e5ece424f84a
z0c8ef277545d70114c558fd27d6140bd99e30bbe43143c070223cf3a428ac9f2864524fa349087
z85a03f06567c109cf16954267fe86cf159fb5504e14348f8ffe2915d401161db5ff2e95e5e684b
z58183ea2dfdcd51c8748037988cfd120be4498a8ddc057393ede82251a8abb86227a8da516bd0c
zd857f144af8eab3262222686529fae22c968b30019820a3151271b002a4ede8f23007ebde64791
ze7f5673422fb16523e7a4f2a08d978feeb1a2de859be333fdee8a78569e1cd2bb943b16d65a331
z6fb04e386b6347ed06f1a9a5dfa7704b0b45183e76bd988cc5b2ca6a2fb6e2f2447f9d60c38911
zaaa67f366c784acf40e898d5a42a5235105857fe08da99f99c1f81e5cafb4be4669a38e10d8470
z7b5b9f1eba7859a39272a90a938bf581af322b79c2bc077fac1227fd38033e920697bb48abfd0a
z9de835f8c6784635357900ee736d2f61632f3c93ec73d75e271a149421a70c773a8e6e81fdd547
z71384cc9ce85e7b58b91fa8cca7643baa30f237443142802b752fea45bc8788abbe3467865cec4
z9006136e39f7ca65d95b30fa04cb5b9e1a6b6e52844b97ed5af975887392b60382f2b22297a503
z4f3b9bea460603b6c655bf95c80d1a5cf81cc88308a7c73bce9548bfc8422d2634ef5202bce1b6
zf9ac0f92af340ba4205204553afdb02e1f95ae7384a4656abc9742e51892442a14f3656a226ba4
zdc8e40a43853a16f705a876b0b3de413d4d1a4cd542145ad499a49094dc2e3cd754bef64d3f000
zf900b729baefda864560077b3f1486635c44297802c4e01803e24d540bd46dfe0983a12f448e78
z525be2d59a5dbc49dc7b3d97dc95bcb723f9b4c80bff11209ceb0214c8d481afc3af93b1be5889
zc2108ed34c4a8694f6163da61798c46ad36294e1f7240d3ed2d9eddcffc1521833f41894c4a125
zf637c6ce31c933887cd810adc0f40dc0acc0e1967f8fce7daa8958e4ea22e30095e2096a7717d2
zce8b882f021a42af28aa593093dc6364503d4f97d61676d61879df3da3c64ca5093252417496b0
z5699a98a782a1c10d702f667c1c0ce014d53db9d1699f399441c4518705eec67e53c80321ca1fe
zaa3c40d363c88fe7cefd84129ae6f620b896bcc88a776df1153fad8798ab36575aa49f25f7c2e9
zd52cf277d68d07a54ff49b87ab839c36f0a7afe57e37f0585d4b143cbe2d5300d0990a5eb648ce
zf85db91382fa9356fd3f046afb27b9cbf6250c10be8886bdaeee4b6f0eb042041a9e976ffad40a
z595eb75cf51461a50dde164fce6b8f9d351a8446698f9cc0dc41b1d78b517124fe9b7f78e77808
ze3c4a273306c43383943094f320911286bd1515503bbabf5286302342798a7f30c98f61dbc177d
z3b4e91b6eef247342fc89147fbe5f5978085c48f7f5e0bbf4c2854f86a23036b7a85f4250e7f88
z6a8fed8f9bce515bc71827635751a36f80878cd9b18aa35ca95e537c3978b88efd755eb87343b7
z7f96507aebc7583498b9afaef7400d8698cd13ed038156f18d5a3b0a283b741d652e5531e5e75c
zf9396fcf53ced824880330a8b4d00d1e302cee99c5ee301255c5b8db465b23f999819f841e1f2e
z30b10568845ee388724f10d847547d6402d800a12105af53c3f3e11916d2bb4002a3ecb767aee5
zbe72f40da9a832e0d2bfba043da7f33cc37f223b978a50c0f845395d10ab8bf7c85a823052ee17
ze4e91e3de6aa8c8c7dbe8535af684ff97e9fa998f7739e3496d0007848a617e33ab63b5896631b
z03f8519dac4306d1b9b80376e68e92cfaef26401fe0d963325be1930649b4ae6d1f2113b10c35c
z7bdb8ca86de5f835d7bc0f9f61b989988312ebeff4c103da60c1963aa0206086cd18d61328d46f
zf9664d2fe5d51b768fbe86b43a2df7987cf10141e7a02496217f5ba06e4ae87bf5432adbaf9deb
z4b9de0e73cddd29a35b53bfa5b7fb6444b2962d2cda7f90d6fbdd8ef927dd84067f51a920db1bd
z457811866bb551f5f098624b454914669ad41fcbb231ce2ef0be3f8c29955eb9c904f2a56aec26
za087a54c60b8e0f496978dee8f3a4661d9f62b5df00e3229130a515a055ab5a21faf2a478cacd4
ze6f37d161b098a9d633df9bedfb660d3d0d348561ae578e8e5ee64f334b3f885c9f03f150eef1f
zfb758e1645b17cec348288bb93ade5414f7531e254262ac19d3be2fd37279a7b500c22597dc03d
zf89b0f9b76426e0436285b1eb7e7ef59bb053197f09d0fb9e53afb1e384750b101c6bfdd8febf0
zf05bc4cad07560c85a6b2065c63b4071f7fee94ef77ec6e6490f032c7d4a1a3278ce9e411e1ac0
z11548be203df9571dea4dbfe82d01a6d75d682adcfd100372f880b6b53bbc9be8c65fc33be3eee
z73f250fdfd04da26ffea00a3cb22275301d06f0b7a431ed3900068e147a2007a3e3945da9deb69
z376efd2766d96d23fb7a5e7bae8d5762cb063e8567c3005aca6caaa5a24e0e39701d1f84485918
z38fbb0c0be4cf0eb6d3221a637a31b19be5c43eec381f128eba4576ce03091e096fda1a8df97f7
z542884f8e322906c5222435f233633fafbe968f6c7e56f108266af5f6e1bc86d1b760e52b3060c
z8b25a42132092e34d121d15106af8ab45e272afcde8ef34f47f25bd54f912d8ab4c2d8d85f49e2
z6ef65964f106439b2017417d0a622588adcc396c5196ccd9c2ecf2129ab895ced92324a1ad6a8d
z3815e25e0292f5e8008a230c323c007336c4c2abfa51c383db4b0305c2bc17d85706e8c80eeb13
z2c0bc888baa4c22781afabbc511f453dab57f01c17d09fdd809e20e9cf403698d390bb14b4a6f0
z3c0a9844a9503b60b64ed36323c6743d5fc5d96bd454a18e1c155c9e1800ab68730fa20f818fdf
za24d594771efd9ea8791a4874471b32666d822b22f02e2c57a0bdc5943aef6daceb6d703a67840
z2e3f8918d16e8bb25f5a9f5d3ee4d82ecbddbbd93f9ffa58508029ec9233a49d728606eddde7ec
z7fe30ae09f985a0252fe1dd4ba453d4b082082ad6e06a32be8822b4ccdd10e6913339019982e5c
zc8d07b3ad2920447aa3816cfc27320df3a81cd6e1518903f06036c93f60d988b72495361d7b1ee
zabfc349bde1089bc402fcbd1d68ef13fda32c58c86663a0a8e49bf715a97712849482c0785c314
z4420d5da613fa9b0c10ef47d7d95a96f682f53a0041d1391ab23ee6655b382713d4afa8ad0e7a8
z500d38b13145bb42bb1ca1391865d8bdb7c6bfdbec20239347d38ed484c64060693f4888e199f3
z9397b83bbe7c996180dec03911d14b2fa468775a55db91b41cc9f25cd91cc2b09ab7eaffc7f697
z8d93cb1f38a8b71e13c52063e13113bf6724d347b3bfb908ef45aca2b802ac96bbe21da3bb2d0b
z95c148ebfb7542bfdefac4405938b8edb3f11580571c1832e67cb781fd82fc6a7f96dd2849f327
z474683b6cbb58804a1ebbed21ace7f6c2865b78a55616f3b3263f436f154c0531f452ec4d108df
z9d5c90dcd4bfc1f92afa0d2a71d513327e19a5758fe758b9ee7c4c4a7a8b2bf68fd36a68eaddd2
ze5258a371ee99ffffc7b07b154bbd0d1b976adf2780011fa008451ceb748ac848cda9cd5f1b8fd
z73fede75d5d9d6cdb31855d61d52aaf35607294d9febcf68b08100a189d76d45e2b3a8c79a1d99
z54eff91112b2bc77b40c7ea6a3602a2afaa2bd86534901e94f548e0020b3543d99f6d3a05f2d5b
z7fe108cf82cca623465319b4cc470ab82f5454ece910c74b68947ab34b7c0055afd1247f2a5b6a
zcadab5546cc5d6d49b188d485eafebc8e1dc10b2112b933238e83582c0597372ac649d4055f52b
z580f8162fe29245444ccf914433afbc16187e6c6757005d7ad8a5f61bff69bfefb95ff60e3a35b
z75442b2d5f8f4c0b89ba801e91f8eb144622f5de430aeff74420adf72581ce8f674296d1e821b1
zb811890475c26723d0bda6351078b245d4f7ab9bbb25e4d3050f46a4372174ce798111b19c6ecc
z4b96bde713cd25de18fbc10f669c9f3a366ebec98a0d6c7569d5ed9679b677e388b42f444da3ac
zccde55bef5776cf7e794be193d29d467aefa0aebef52c3bfe341ad7d8eba8f257cf0b27bcc52c3
z9c7b8a7f785622084cbb1a85a7bd3eb47c98167fbfedc9f9f611fb14345607ee5ae30b3f56cfaf
z7cd3cdef98e34bc964fbaec85f27b589946dee746f28ed2d3386dedd20d1bb0a316c43c5129856
zfd9105698ca0ad43f319b4d1d6902849d49469bba1c2fd19c5fc1f32e85fd00a24503ea20e789f
z2de052224060a6b3c8bd2e6f2b82b86e2fcf249f1818650e5de9869af8074cc744e24612e2f691
z7da7ebebcf042ed107f9c5d99834abfad874f950d16662bb0c12a47484699dae7ff71cfc0405ff
z32aff4b5e8b001b79cc974222e4bcab1cac028cc1e6b96eac1205aed09c8dd2b831402d8abbeab
z96787c112f88c78f94ebdf6eb4d88f99e7873f5e6c4bbb799d7ae66865a7fd466267a7ff3ee96f
zaa20b10fe7f1f00bc96889a6d462aa6afcbcd00de27a547f303d69b4f693e6b560fe535d71cc14
ze23d810ce80f26b9ed98dfaefa99a1d8fb9de0b183f50238d78813389ea0add32fa774a6b7503f
z82ba3991ea194dd371442f3bbb0e566d2a87cd75c8833290106034b2b86467d851da11ee1fb9b5
z193f57a69ec774dc2f2e305376f9e050cefeb273d460143c38ced83d7c00137061fe2bf484e158
za88bc6e7e1523cdbcacfc1d55cc0ce26ac8cfcbbd2843710881dea6f7dea37e5271044d300ad42
z93c37961a66fea8f1d6a3a06078c76356491a04ef058b85e224d42b89163b0ae66e6a2bd4fb23b
zea7ac31e5ca833c05e1fb928040cf9126da5b517e86f03ab16c7d80a80ab0afd3d28d854b84b1d
za2021008d563ad5c1d2de4273bedb4340075e6acddf54b78fd7c9c0d1b073076b35abb2ee10e0c
z408a754b96c090af4a3094a11786a25038a59d5a0037ee476647c7c09560ead1a3d3d46ca198c5
zaccc14b22eb2a542bb0daa211670c01428e036414f7f1dd6e66b2428ef3753ffc4f59d8842e2e8
z3ddba7a75111ead61fa77eb021ab5a0d584dc03263c3aa283214a915e492fac589ed75769f7f9e
z66b8c463e34d06a58e1950ebe91f9436da4a7639f2a8b77ff5f4d581fb79213b75874ac58aa0a7
z4494c6b0de09bc9de5119dbc060e8304b2494c3a862ee5137b20e2ef9f3d2803883fe98a9e3bc1
z6a2242ed841eb8927a17380dfd1c600027982745f6973b0b819d66999dba23fda9a018cddb0526
ze923ee6280ec51bdce86f77e46dc007755ebdf1bbd6529b0d2d95a5a101020baef0effc6c38a5d
zcdc285b4c7ad1fd0412f63b77766ad7545d0e0b86a6230167d6099bd80ea3865e5f870752a4873
zbcefb7efd96cca8772f75a2f92544a22dce51697f0b8b03a5b3c113e92de5679d1712062754fe0
z234edaa812afea872eb20b3f4145d7aed641df57764431ff75e602c0215182390de189ac4fe70a
z7ae3e8d453d27bfca5cb0c68feb124f6168ba97c8022d42a0bca83add21ea6239a13092338edf5
z2712db5d86ff902c99b2e4c3788e0a3c2c52147af101c844efbf8a0e2898ba89be9595eda3e333
za18854b9c8679ab5121641d8d7183c3d04624b4213db5567bca8d203a2014a4f492806ea5f30ac
z6ed33174e69e2ec2650b14911b42cb621abcd95149d658db42d6b53022d14a9c6ffcd2c1f266d5
z37927a1c9b24d36e29917028c2b32a7cd1047c45e272a12652c843f47553d2f3756b87ef334a02
z8f2611c4d8cbbd47eb26700033fadac9d6b175c71131e646b532abaf94ee4ed3ce32ebfc561fc2
z5bc525a056aa8b383d529c27e0beb539a208bbccc30893e3514fa231bcbd955798ad1a3cea0507
zb77731ce1b7e4fb6f4b00b3214e98fbcdd23126d762ad9194356facb207fe20077e30c9fc28e82
z868e057fcd733c3179617f805d22aa9a5575760a716cbc1cd8d6057f488f59af380c474b9da6f1
zea65f715edb5542ebd110da7e75e5f337f6dff610832ff51621a1610b97b6f7fb9496bfc2ccf8e
z33a87c3e0e3884b1b135d28c698a40418e962c72e7212c0f6995c056440fdd99c0131f43cc82ff
z76f64848b8cc99bd703d94553fe9611cc80d447ba3c0c123a5ac948db45f27a8b536fb294fb05e
z2ed106dc5cb390e9171f6a7a234bd9030470fc5b1eb2eacb0fb99b08319e5086c9ddb4051d8192
z9bf366142496b1c6012b46a70b9907f2175245520f34426d0179d6d354d3ee56924bb14693a9d7
z1b287a4b62cac96f9d136078419043a7f677b7ff952c9b2081463cd9c7d2f480a4b63037518c54
z36b1b9e683e75134076bc4075c6b1151e4be83c10b14bc38b64bade76adc966de8b74af7f3b62a
z74f45801fd52ae8b56ac44e609ca36f49fee184f80c00f5fc1d3ff1b86e1d21745ba35d6a03f82
z954d46303f51e7153fd7325ac8b46000a3a5669db51b31dac112bba27c1ffb038881c4cd162c68
zc4991b04d8832df2528504e7ce8da61dab21aad39b0ed1f650df0f1f76fe1641ae663f05d6f94b
zf6301edcb85a1613b421c94b8acefc5a183fe074ca7a460dc08e4fae95f984deaa243cbb43612d
z7364330c832c9e00ce39066f28296c40896c609e4d58813e14bfe335eb20ce7eb0b4058161f529
zfa88bb5ae553052061884ee0dc9819c007353e024bf0c82c57a3a1221c802a4a2e6f53c1c47d07
zca1593759e5329c6da9071eb74fe7366a5b0e1e6114a184923ed504fc3bdef4859fb3921e1d20c
z1f68076b692c2abbe81ca2211d37e5d5dab880adfd3221f498b5405a62e3bb28199ea9bfe10826
z1bb5d22255767f08a9bab77010d406665e1f6f3f04c6b71f3d7f974f3fe11dcc52d921971f46c1
z3ff2ce8b091988305e2e7194de8bee1744595f575030c30122e84729c62ccd0ce3bd4306210920
z87d4a9ee1639c4296f3bb9d890c89cc98cf760647da1cd06e181cd859e94d4be21df35348f7f19
zf2bdd25a3b403906150edd108884e76d4827fdc39a44664d193002391015920922d5e2fdc1d161
z29a79faf8fbbf19db97645895d3b25dad751a548a47f3195bb894db8723384f08d4865c30c732b
zc4efd40e56c5fa8fabbc8f783676dbb085511c40e13b6e0eaee231feea37a240be9f071542cf1f
z0d38072b5211c6b6a8a66ea5398981980533eb5a8f6c12b2430f61676a05c2824748b226cb5184
z04dfee286ff620e95c282dc62d62c7067541fec8b472b18b97b7d276276ce4dda4ff6b11ceb712
zd36f79eb3f7be639ecda393668dcba0920730a3e4f870f5a31d60db76d657863113c62fa3904f1
ze3b900afa96eaaeb29042d22e6aba3266ce7944bc774de4efd6b29bb11abc784c3726300809b0d
z4899cd758b9f18083932308d2d10c44d331b085a041a8ea01286067e5bcd6664bf960e1b0a3ad0
zfa25efde15a3808ad876d75a594f88fa4982bec6fe190d33e2f9b30257f104b4b87423c1a6b9ab
z3198ce8c8ea5de558db6ea86556c753c84c61108cfb554c9ab532a72d5f80bb2d419f8cec3accd
za8bd294db941499eae70a022565159480f5d3974df61669036d48b4b45adaf27448116684c736f
zaede1cd8e47d9d9b2de6002355f1bd2f747ffd5959702944faf5cef7f88c9a4ce20ae7b3f2ea94
z15f0923fe118c5be81b6b5661f7c03d1aa6118da7b766730a6713f65011feccbd88500523fd06b
zc07c8f315a46620e104a8ad8630022bc6ebe065dbbd5a19b580a00c5e70680fbc23c4eb0e37fba
zf81c41222897f7223676bd3ef3f2df1b18266e31e65aadf13a5f0c8700fbe86c2679dda1083140
ze51d1da5ea8591b836a714713a23f126f4817ccf91659d1a59750207dca6885c19b1ccf2992de4
zb219a1fdd0b1c04320ef720380dafe233bdb828ad033453a940a5142d64569440bb2b5cb98d40d
zfcb10312f181c8da239d0f09a44e55e74cef163014186893b843c08f1b700020e90dd3a17287ed
z9caef5e347241a2b0e530ae12aaf001d088e6d9baf24db7bd6b891c3fd073a96e5c5588c1d677c
z34011ca394975b7d0875fa8b8f76f1e5fa1fb1f42b3c21b69ae837f6a50aea0c4636cf3d354618
z7011c730de93e7e8fb663a93bfd10ace3165b4097c1eceff20a7eea273471ef6d0b2894bf8734b
zb7cb6a9e1f9f9cca6c7c599ea0ec0a9afbdb815d5bd3270e1feed4f3e5b98e8492f475f5614eea
zd6e2d8b8785ae77f8296b80f75a5f56f4f32c614d31b207f13e4e9f8ec806e6aa0001f81472439
za1f51b4ab3ab86ea74d9e54a07000cdfc8d38a284610ecd5968d06a2ef2d24b1cbd9d7819ea8c2
z020d0e898fce49cf52a7488fd60adb9397ebf2c47715bc8c5ae54fe1194c699d7b1734a3df0af2
z64b234b11f46c0667766878fc544d31ba5fa6296e7f8142a0c9f0c9585ffcadd6a13bb5617e409
z1ffc6d1c2c1021270ea56e11839338b9c61aee81edc4a08deea84088bd469514080355bd0409a2
z4f2fb76edcfb729e5c63d897fa0d0f8fda9d15576705ebdaa9a9458c48a2346cb6bdab68745dab
z7e84658036568048391d7b16ceadfbbfb8f7d20b00c00947ca684b6a4b055aee2f4e79df8caff1
z7015f63b3fc45dd40ec27bcec665719718495b20123f0e4e1cc4641c27cc25de86366ede0aa8f0
zb100d0d50a22ed23681ecf96d2dccfc4122e647a011b2aad75c641efdae8b90d884be47420f652
z6b040f2a437816ddee461527fdd8d05789dbfa389be806624899e31b369b41cb7f19ed5b5e6d7d
z8e66fd92a5f3362b997c5669f7f9b84d1a924265b429a9d1046a633690808e1c34d58788396305
zc6944d46856e5c309da464cfb82a8726465b007f34ebe15aa32bce61df502e35b34457184ad23c
z294284269c0098c36e27ea602d50171fc42826d381cf70de8a5668ac5bd559ddd3ca9497a1e995
z4217e606f38a8830c48bf369603fc4d99b347953a52589f083fc80ec2cd8bb355777ca1628c287
z2e495e400da041afe5f450e45dc456462d6c0179c764aecbcd0e4525235a28e8f9c7b5fdada01a
z2ab02893859f12b73121a5c27c9aeeb642503feaa7eeeb484098ab470517cca906e938df498a27
z3164de82b881db58c38e975cde6719a56b64b731b9896d5c4419eae1441fd7d1c8bc5caa5e7590
zf75df90021fd28eb53ff2564973865140044e4c859564b3fe0482e130552a1567504066f0216ca
z7ff64071199a6e4e7ac39890533db85d7c00ef6f9093df53200e83c75cb9f894434ec37dcba779
z077f379b266c6bf99fde2089613087d44c5963094f45bfee1fdf557e280f4d3359baae3277cd73
z9cc42c5bfa83a14db0a0e543634761fac4b32de318e2f281fdcae200de4926f281d1a719fb0877
zf2dd9fb19bf237aeb84cf2955bcf68f12e83eb5f7d144b12d443bf2203dc3eac7eda74995f07a4
zd5f08e45efb4d007d0bdfcf75e4a13cfc261e55018c56b9fcf827016d353179e79e0cea33338fa
zd583a16082aea80191ed8165e00f1b4515fa563883d96637237eb2424bdd5c8e9ce66674bf1db8
zf037c26fb76be7454cb13fd438c370de6a666d71f12e7f71ff409623d232ae8e705ced574c04f8
zc04542d67537d71114ef4fa70203c335947688cbac7065f26d92b3d439312d9d3b149e88ad2d64
z520fa4e4be8909b4f6b4cc13dea800301d6ce6845471259fc028d7bbbed2380980dd3f111374d0
z9a2c9a582b9998562bb92e2cf474b9483e4397a2e2419638db58b229b2ec22bbce07979e627394
z9c7dfeb79471e6ca97a8d994b23069004668e895b1a7460c0b24497c4ec10be8a9aa4d4657f8f1
z54c3fa58cd19b617e2c453d8868b8a4ec7ee89a2c7b4993b92f7c918c946c077ea6aa0f4f5c864
z444b45392375b8396e15ab4773c01fec7e64412913ce2b923b67350e9d21fda4f7f0f3cccdc335
z496a9475d4f03c55438d2a0e6f614db7e0dc3fe9658a60d6f26ad6eefd4144df9f9f0bc30056fa
z5cc71fea840cad3442b1765782fcbd8c4aa86267cae20d2fa551ffa1951e072ed0091d17c66dc8
zf529e1fa9b27c36489dc59f19503a2231e60db6cee1aca20841ff843cd6e6beaca048e1de45553
z56e38ec0874fbb954216396bd6d134c60b891c54c7f795c1bda7b818fb6ac50ae91185ee282a4c
z9d9960475782235982f7a6d339f8ca1191583a4f1839d716044c611cd8ea482c85b9cf880f8f74
zc1275c0aa98aa8b3d373ea352d4d0f771e25312854939f73da85ad68ee5b7d54ffe40ab57047a9
z048ea2acf9b1acd562b31abd69462358ef0d89ef0be8db2c32bd9139885d7398b132959dc4d543
zc37d916ac793744a20693df5e101c1943271f14bcef6a5ef2f030c573a6822fcf63409475c5f48
zcf950742119a7c2a5725d7233eef1c7900b915c7ad1dcd9a75a37edfab2d94fe26b391ed4a571f
z0047d8aa74bb0e80fade20f80441280a33b91ea60eb9bd360afacefb206291720b7c0e2c575ccb
z958e8485adc814da3aec5adce301aeba4d6da6fddbaff8ad480f80f06e8c4b5675dc012aca4ecc
z0b86f3ee77acbc9131a7fe742648a975e6740c30b30b793fbf28a1654a27fad41df5eb44bdd7d9
z75ac6c4956c6f1add6cec59e8842e68558aee5361b77434aa6f2edaaab110ea68129ea79eefe4c
z6925103467f31633525fa20a51e6e488930615e2cd6e362ab97544245f6a1c1a258ef9b54dd99a
zca80bc7c6e72a677f7403d3c9ce4e6942a7512b7bd9c16ba1c766e0f28732604689e23b961035f
zc81bb62c4386c31a26207b023bee49800c7a0adf7b14f60630db5335cab36bf8a7a5b1955bddcf
zad6a4e36382c036d0bf6eeb63f25ed0e6f11e13ab0bbfe9bc7e1de2d509544986de7dde5dcb2ed
z5ed6b7833d389b3a7fc051f5db5b25f79fe4c7fea4edb0d17a64552659152437dc4b4b0c1dcd66
za1507447ac64711b718a0a1ea76547dfb799b7a0ddea872f03b2d3a98acab6674db3dae53f63d2
z4282ddfea7dc55ce2d72f3d8a72f63179ed0a75714cf766305b7a5cbcca436f0df32d5c2af5893
zaa455566cd5cf0e18b9b252bc92c5a20d8ba058a4a9d93cd79b7b61064a5bea0b5b9b37237272c
z1f44bc5eb379ea0cb7363df3f0e3cefafb91583b4afd5f3eddcc7d2a2fd16c1612bbb9d4b3a060
z7539533222057843919f060989485207ceac0b2b16b8ec8b84d731a1a3050b1a5257afba4c2290
z578efd8a49d1c7ae82fc6f5084bb82fbbde50dec42dd81e7029cd1b075e71c97de68bf0cbddc83
z50f12b00adb99530b27aefb838734def1c3fe7a7b39e58aa7030445870a3320c3d5ff7eeedd5a0
zd5e03eeceecb1a1928dfcd3d808daa8277435398b51433909675066dc5f56cf3034449d0975986
zb3bc0b33c05dd70520fa248be5f5e090f5e0b2b15744c183705b8b0ce93526fde1836476d5c58c
zba403c3bca5b198fc26d31c83014bd2a3cb6e08a0118da4c7cbe678b68e6a7ee0182edff857db5
z0aacd31afe7c44616ca95b41ce2d2eeb3527993cffc1be813092976f4036ac5115d579e544cbd5
z3abb2956be064153c78b14cb5787c1a9c4061f97517a7925be2fb804abc02db58c20265a59920f
z18236133e10a5ac4cf307f3cfb1a83edfa1c76404a5d8586899167129d48da0e5e6fc7583b58e5
z207c134a62c9eacf31bbe759be29e2aa7bb7f22f5569cd0e43160962709081eb464b613ad90290
zea35b2bcabb2078297c906f511f3bfeb152886c8d7639bb96cf39239b880c3fda6a6133bd1acc7
ze09070db9e232312099cd06e8e42829ede65fc3e58fbbfab318d94d51b562ef7da654fb776f437
z358b9c0169abfc9312bf76de21c561b9ccf4524ab6621cdd9e071ac22f7d685dcbd420b498df38
z843e6188ed0031a395ed689f3f6bed4d231245d0298d6602f2d252c3fa37ce009cf662939bde55
z7c796d2812b76499e40d2d06f8ca591d8ecb151b3da69de03b8fd1c0fc9eab896d2978b52cec5c
zebe2694ca20dd7860e2074f99f461243064c760241d727b1770ed58189493d6425f5bb786c8719
z3dea1385082c9149f4dcde5af39bfb4391d2998c1e6a7029ecd57ca8a647aa9d5a83e312e26c5b
zc7e9a4e774f37b6d2d81de25ef9d991a86538f6cfb3a26d95f0fba43897cb350a7f359d0138e4e
zcfb579dcbb0033c658985dc620349a623cf80da3625f1495a4fbddce481bddaf823cb3880425f9
zeee8412483c36b4c93f41c5891a327755ade72968fc27732d7aeb62c8e96af6deb7a1c92fdbd78
z9245669571a3c323bb7b1a4c21ddde78a3e533ff8ff5855ec51d1f65b082ac64666acbe45709fc
zf3079d99949c6b38092e9649ee5ffcda9a90e7c9a446b63ad84a2ab23d9dd828262db0c14cf97e
z8835b6605554b74a5abfc217472012ab3c34cab87a108615808d02b254c5b06c3c01258ca002a1
zec9fe79683fb89c189d1887c0b22d23ff74b3e07724f11f2392effc40bd9ed660b006bc25faade
z6dcd07fc1158b171169a7ea35d026352c05b9f47a5de392bcd6d9a121dcc38f078c76e43224aba
zca0fac4f425dbd44b1f4fc3ab744305948cfa410404a42b906fbdb92dfc13f4d29c97525a4ffb5
z5c977736c6be853c2ce60481d257c6836a23d079d6361b2121b22c102e0512a61ff35c5d96ec24
zcd11a2fcc8833a8c545341ff1146e1eec6edf34ec7d5dd4b3b8cac3b55e4659058d8811fc48d27
za73d4d5d76799221c679e7cab01ac1c2cfa821de428e0642d6fd38f90fc71b572467042b4071d3
z844ca9d7716e86e24a511496f6b109f1cd5db64ac7e005b544a1941fd6d54a6a3f450fea085964
z247af0a5ee44551aaff1fae058af410e647834480bc5e603728e38bc9f093fa253b72b9ace8ffb
z4122b4f6810a4f377ae3a442c6164c9e4c9d9fe32472fd03fd4b682a74d0cf426f3e6ed5fa0953
zc72a347b1fd6c89d5f00ce25b1fe95e083ed9236535e1e55026296badafc56ebc0f38dd49462b0
z47c1274ff1334cce41c4d194e8e5df277a82c77c4c73e4edfd65698ea38a151839444cd520d637
zb3550f855f0ba2006173fca03d14a5ee9d4e3b1734c9150852dc900d6189cd5ee97f071f50dc50
z7173e21a53e33e772cdec0566f3a390d0e87bc6b587521ca4fd0002f48aaa9705e68baeeb06fe8
z4d2531c48a9722f4e9d1823b714733b3dd2042d0b767ea057ea0b4cf426f070e70a16763fc5c92
z0a40db108e63e06b0133989d1dc4540db3432b5f31e0914831cf91dc13ebf050f8e16e495e7497
zbdb56a52a74457465c1f9d0963df18e9820532fb53a7199ef6e570aa4adb3db663905e3f191937
z2a381f0cc7886f4b67142c407774e86103d1e3e23804040664d36e0ee4bfa3ff479fd8fd9c214b
z739829d31bedb4c459ca9c03aafce899f3727a63a5d53f50e4e078f59fb40cb15169e6f1fb0595
zb00c04c947391433e5338dd07ae9f7d7486aa84955fd34c99d1d0dbe1e4598368165a83ab96bfd
zee183529eb43417f676f1cd02f8e9bcf8510db8c9032b9e1ba988bbddf4ea5dd7f516c034802ca
z620c1baf60f91809128a436988323d8c2644e81a504aae02e9dd83545880488efa91efad60dc1d
z1f2e4fe587d81c8aaac5adb43ab84a32b9c7865e5d2f7747337e2821bf093072aee2be91beff0e
zf13d0fb877f52cddc8c80e1fe94e4369408dec5e715dd021b6471bb90dc90551ee167382d0a260
zbf14a7628b2253f8bbdd38e19bd56c83ef7ca1f421ae7a4e5671ab52f8aac070f84d0b2f9c1539
zf9d20786cd3069387bcd763ecb352f6ca70bdafec44741d3c42b0a572c09322f364d0f98031828
z2daa77ed855c7a2374c8653629ca251ca9134b3b10d3ebf14a47feecd87c6eecb343382ada5616
zf782c0129776a675f3885ebb39279c54f885d7c05a8716d582231a1cc5de36f8a6686bd7a005f2
z5ff5cf7da92f97d0a32f59ca61685eb95f589af819cbb4075547adff8d50dc9b9c10d42ce5d4ce
za8b882fab9d6b2819627dfdd7ff00300fccbd91ec81766cf7819722c179cc1ba71dce0026294ec
zb1be522892a1724a72165619dd5fde990830adb16df80fa55111073fca5fd908726f3fcc31195c
z554eb549ee65194ba59b84bfd105b32ac8722aba11b23dd4b90bde3ec8c8dc66b953ebdba33aff
z708b2b4d92c8d0891c7f17c0b785b911522a2a0eb05129083a66cb0e531f2073a56bbfd928bb86
z8b7c00f69e8852a7483f73257dfae90ad4ea2f661a15e6a9509c2d6827f42dee62119f9042ff72
z2c366662f59599e65ab7b69af1bde06611949481af082c78e05463abc6fabff2f676b3ffe2f3f9
z236c4835afd4fa7217c38dab72de3df0e3bcff2fefd0a556513711170b54288261054781cb8b90
z2d729814b0fcbfb5f6687bac1e8ad4b920542f548d77a2fd32dde2cc0b24c0403bf9a8803a16f2
z50d783b0e2273aa1ad4580af5431c5e10570b7c62c9a388f11fb5b6de14ac471438b970b3b3173
z22b3173b61fc95e2e5ac72ed9ff5170b0806f113008b511c3e34f2fad20e6a7afb460556d72444
zc0400d2b77393a127dc46d77370a4b9a39e6798a40921f0211d41d246c4264a368fc04b5728596
z9df1f0812fd6389b2cecc44c92f6a26d348e4e530403c57ebd6f0e9d496ebc2aaff71b5b6df1b0
z4b215b40613035f2d0d466cf9017b1a2fc741e2ed465fa5bcb7ff34dcaffdfdcf1d0d230e32552
z573831d183b031ec2ce7dd0c3541565ce53765cd4f97edb59349438c5fdcf81cd47bb4f76f8c64
ze5de27f6c69184c5e7a2cd8e5d357220590573e8788a46458da6cd075e29b0ff930c164e02e4df
z0fb7699cb6fc45ab1e65e79898337fb955f8d0b2b133a8a3d30a4f813c344d90c35d981dec4da3
z55ff0a5434f0cfd6fa219f890b122e2e4dd2a2cf6fa163db4cfc35c9017d6b09b484bff0bfe89b
zb845fb410dc6031d9a8142897a7a85c48c39b68c622ff823f424609dcb31c3a88bf74c4be7b36f
z50ec76897558c56030604d8c4144d5f2783cd17f8d094d3dc825742a514f89b24a98a92ec4154a
z8399e5f5d199435340f12b53b7b27cd6a5170cc13989e3097a77224ed140df363ba6dacc507680
z284a91aaa0de273e82e6a84cc63de84c1aab46be89c283bcbc67b39df5ee4d047bec2f19218efc
z89c0fbe4470bed1dc88204fd008439fb37b27f0fa2fc00922988d9caa44fc81f368764bbb5341c
z2c5bfa1ebb196a48b16b20de08a839e249a342a3e77d83e0d69bf9abe4add44df97349d1f617e8
z80f74fe19654353ec44a24ce09dab31ef48a58022f3c8373b35d58987cd11c64cf1400b50e4251
z9476c3e511f3d8bd50e087b7f89cb9b1ac5195b30062785bfec153609040de0b0481d70cfae541
z00780be260107d60642f8d3ad50186b68f4c7725b50c16088ec7fb7033f1e8faa5312ea8a1d5b5
z1933886590bd407a8098d2aabd34923e16ae6c3e662a8ff2a3610b027f077e320d8a2b42233d26
z01ea55d83b4af2b948a3f38c59cf7daed2f9d9d24ac886436b07f810db8e72cf44655338bdc433
z4de03b971ac0f9521cffa0d2effd7ec6ff0bbfb2b4d7f28644e704537158a573bfbd5189c26e92
ze423708bfcfe0115245b782596a9b9a4cab6c803a2fb38ddeb3028374e105c995bd58d18fbf946
zdbdb0afa7e26abdc8a5a5ffbaa8124d157470e4ad7900de677d24eaa2acbb7dee88c442511dbd7
z795400aea4a3219dd836efddc9c38fef74f4a1ca4cbafe3f83c0f2b51c3db1dfb6980554049cbf
zb90819cd6f4884e702d306781d03be8eda15c78ebd02eddd3ac917f223bdea4767c945331086d7
z34ec90055a9b92a6e2897ba35e5fb3320e27d2147ac714a2d784da989ffc0d3f234e578d1977f8
z1ba818a08677700b7a8d8ee3ad0dad97d8b237638d8de4e70d0f14ab17bd7d7365383837f4871f
z3612c716d809f6f963d386fadc8794bf72a566e3da77651489447312688a12969aebab8984f0c5
z83104089a49637d35a3581a9eeb5503db0deb9b7090cabc52178c76595f0fe35ee6a37e18c8ddc
z25e8ada6df3f5e826474abd685f58ada22929aaac4bccb49a9d750c6c66005e3390d20e380af20
z7ca7a0dcaffe22586d2e2de07bf1e130007f81dddc27cc61745826d015839abb302aeeb68f58a1
z1ed7f7cfa7228e0fc137a4cbe06666a3a1a6c0b23dfa0027f23121b67820bf215b4b40893a44da
z5275842dc12e29ae47735bd4cee7ec0b194b00f8510826017889a57368876b01f77f4192eb5b82
z02a2e5e820f16b431af5b05a4ee360d340435adc7b683e1226ee7543cf1a623d115c2bb928e374
zbfd95956092f33142a4f19a9b2ba695487ce3d9ffc485c9a16fdec93b780302d860b97a276500e
z9dcf5ea3d114c109ad740fa06b33475be116aa2206276a0de87df6301cc431b30fa73b31be21cb
z2ff4c2f3e82c5842e67c500620cc3d3b5ff59e4f417d2175e81a031a7ecf47ed48a86badb3a5ca
z173045586ab3f60628a44be30aacd2ae78b355aa74b1a84103160cd51481d50b04c2e69b063e75
zc285d8ec9bb1a928c1a95047c9a532dba325920b5fb07c201f2d9b16c4a7f83cf468ec851da737
z7c6eaf1b744cdc40ee2417229ad96b685fc639bfe3f3becc9429c18c5237e80210b957a5e72dc4
z8dc6812e4dc36b60bd32fef2e1a0dc4846dd35997903adca53e55cc014ba7711f6021b82018312
z618b981c00fd8e9943f598838348d2cef08c62f343d74764f5e8424e83101e1a0724b63a822660
z1ec0f2a920a5c991a2443257ddcb1c7625b68e6092e8e02aee7fb216cb941d93ee2688199ad16d
zce15a1d5d06dbd0af87b92a29b852356bfe3b09d665ea4e690412be483926c51db45c39f2018dc
zb64bafc4e648ba84638cd48c59c300a21fa77c7bf4053d37e2de1355bf9bcb89e3ce45c4f90f42
zba1b96a1cc712845c4965c40c0175d56364d2e02b000451bd506ec0f7e25fda3d56c8394fdfbb2
zd5e8a676208ad4a1f1ce924f20d0f5cedf9aabf7836d0011a1a2b9f2e21c17285fcd51b019a3a7
z34049291f645d84d1df09ca8abaf119f7cb9112dd744c6e9f212c2f0858350bd7395c9e88e16ee
z4222db5a03b7693c773073b23a41baa6d9ce00b827c88a1a1397b24737e82738809a351ac94e1a
ze2e24cb46e42684304a16d2c9a2f064a93124bce02ef5cba25a25ecde304d4be9e2eaf672bc5aa
z27730217170eb95e305cd8184d0baf6e84a3ded0e4650bb9ac0c7a80571e472c4c4aee0ac7cdc3
zabc960652ff47b1bc198f8ed534e40e9ceecb6d782923a0114960b8767616b85b07896fc7e8d33
zfdb586d5a0b104f0e5ff1cd46ba28a7adf5e3329e03ce0bdb8ecce636f150340059e546a4673ec
z9e4762ba9233a085a8c05fd349bdf4e19442a5b58ad494f8d8a1d7ef4e88b01873f535b79cd0a5
z3ba3032e148dfb6e3017d4f3a61bfbf645c5989507737e0301ab9f9bd029fce7ccabef3ecb66d5
z14f0b906250e230b0636327e278418838baee7198b8fdf591171521735fa7870ac7c4e594ec297
z29b760d48241d60f621e41fe08b4784c67eda88a7b130aa01411066348cfee1de0df05d0b36318
zd6251b579fb2ddfb9bedfa97dc96cb7a489e3ba57129afecc051239f86dbc0cc2fa62279c2a8cb
zb1e0de06189b96e3165801305655afb747651f58040bac40acdeb58d5bc1e29ae123175b4b3e2b
z1ed551ff8829009c1eda1035c86c4fa3151759243358e4f65cdaa4db6c1d2b6740305ca8725825
z1a228c763d85bf1bd680c04fb57845ef08f42a2f7f4534c0a4f5255623e42642190c782bc4bb5f
zf9e1697840e40899d21081d2d09700573e54dcd1c080443183a33adc9eb26a036972b9189dc997
z8a0e9d1a492f2f7971a9596e2c6a021b291adea9f54f14b9d16a41cf0e5f2378dfd48e03192992
zda05590039214ab828d28c89d953f3c17f003ca4a5f90688cb5efc560508974dba574787a5723f
zc67569affe663f99258f9c9663e78ff4a9935ec7f3eb5f78d3c475bdb03a5a7f8c998308ed59da
z83afa61adf41378614ee6e747125fe8a0eb0e2d876a5ddb379afd6a4aafaeeee562c6665072bca
zbc58b2764a8dff2bd52181f9411ca8639b1baaa98ea5a42680aa52dbd78c08ddad710af0c14213
z89330d2dfb1f1cb05ddfa2b108afe0d67036e55fccd8e8d58794c6bdc011d1cf9b68de22bda737
zf6677e0df3cb7cee75b05ced775cbb722a3122d2e8d0ce9523735c827c0df740d576435b9735b9
zdb5e6b1602dce0db43829cc9c972fa5f714a087dcd8553ae77338b3bc81771c53ae1eb137f2424
zb8f7808abb4bfaa5ce8db458145c8a18168ba59b62e90fb9b8252195732d14bd18ea6581406d6d
z33249d9e6f5795af247ae73571b9613b69bd3567811871406e5937aecd1f037365fd049a60f8df
z0680101e93b3a76494f7bef16a379c89ed254b445bef60b8e506ccd00db04a493ddaa57c327a8b
z4c90506cfcced29d8f060e9c072028d9b318f159f1d1ab5962bc8193eaef11b849734842d0977c
z225080ccc6ee5bdb3666357004841f73bc9c1a1b2fd61a822d698fe27aab1070fda49dfe189610
z1783495ecb38d9f018b40b9bf024d7f8247f00ce6462898de0068bb85034f0a59e7ba356bcf22d
zf2ede3464ec2ffea8079d717f7e8e47189a92439b845d4273df7203f26ce75e03e5391b5098f06
z7824de99c634b4081f0910564440e988267bdfa16c059b1b83555d5f4bd6459e521204c240a64b
zedfcc3a15f359af78f79b2d99233662c73fc7a8f47e12c836f9d281b6194012ce8221e6162a84a
zd9aa45e6e18a4e2d3a72999b69b100a5656eecbb325a28699536bedfea1db5d422ac5976173e6c
zc4437dee5864ed79fcfa846956a2d838d528c4d3186fea43c3600bf8f1905804431453de1136bd
zc7e6bdc27a8fc7e103ece530580e1b45535495c38d9b3e7a701fc17997b866b0386ecc5aa4f25a
zbc9e4d07344fdb5472d8afc1df752ee074699529c8b607a3ea56cddeec51fee1f00fee12888012
zb40d7c5b9654518dd6690d1ec425e36ec511194b3fba37b675dec47d02a3e85965591315c1d570
z203a150bd878e17e7310aecc282f991af26dbeccb307454505fc104941beedcaa155fff57cfa8b
z314328593ebc2f39f668ee4478d52fdc7e1cc2d1338fcacdda0b16a46e0256ae1f5b863f4b0bbb
zd0072e380b2b2b2c1ca3d94c1fa065e73acc686d527551ed405d28de4e895edd5acffa32c75bf5
z80b4dbf7b81fcaaccd77439933557016e7733c4dbae3fbda65839eb33b08136626b6329ce556ad
z6575503b605ccbb7b506e4a9f774919a28ca610aacfec0657d4aaab5346f49f22ee63dd42af3f2
z242aefab8f7f57f68d5f71723d83534b1b63aa53a95ad236174611dc08b9110bc0140dc607b2e0
z125aa4e2e6957ae2657ee58e7f4cddc243a3d49525dad6917c566473c19440e148bf3fa3285263
z1b36449b64566242d7a5418937fa6a7d0f01bebd9fafd4ddab0c2dae02fddfbf761b1e0c61582f
zb550e9df5d6edbd35ea3a0320ecea8f09dd3d7fb63249aa1bc19541b540b1f04cf3c267201104b
zf1fe3b3d98aef7c0e1a31ced78f48db4c801c989f9702b7609a47a6fe974957ae9d51882ed50c2
z0553f0ab8ff2851ed9440aa74699ed22a0599418fcb37561b15d6fa033a6e5fc8b0a988030bd60
z2c2b3122f58e0476d478fe8965988729d6b85ca29200da73e3229ed07601e67750c982aea9ded5
z55c4e164176516d508e4b607889cfd0532854ae500de22907bda4f5115c52bdae3072c2a9a5b3a
zd23a898ebbf76f8098d539beeddb7021dc4b119d537e34a90c1301da1fe4c96524916f6631ecfa
z292e38b47edb48dd8d68b60dcf77cb8fbeb37160ba50be4ddbc1a4cea79cb8a010d98cafea94b8
z6761dd5ae5baf018e42204d23d3cac44c5a816067dc0c678c97874a70e620a31e4a7e2b06ac031
z1bfde519743e18b05f15a7212a8e849828183e353db165e3030752747984480a60457186dea9d5
z5767ea6664875c85db27c140e10bb61c17c0df5c83c9ab838521887f6609b355ea1e3411690378
z3b2826976e8450574647747ad2929ec6c29480810d1c4c3d38789b47ff2d917bd4e8c5f236791c
z395ff1bf89c25330952d56472faa0b811562b142aad536cee3f5716992e443b6b22b4a36aa2751
z71795c35dff02e7b4dc07f6a2e76220edfe572002ecdc9db126d1d6a1edd59e218fc41f1b0fd40
z17af0ba6adec4621ebe31da04eb6530d638da459f536c4251be032fd1dc10128d9c5f2bcf1e1f0
z768958b82ab058e724a3849a6f1656c3e833a5c8807fb83c8e81d56fdf51d0e948f33f47f5fe32
z77181188e83d64d1b7ca539da6eb3bdc87aeee8a7ff190f0113440f78e30fdc8a56f4a6c1c39af
zbfb9c9732712425ae38fdd5a4da8576b8034bc3a3b05d5ee0f390d65bbaf0b62ed15a64986e678
z6a50d3b9bf46d0c013025c43fbadf50bb7c0ba885dd44e61628051b8e00e8917b0d17d61857d16
z473809637244b738d8d54468a94af1e37c89c3f4d4dd471340fb68fc05a6d723681ea950d0bae5
zf3c6592229339f0889ad20552a42dced14347ba0666415f6411c76ab014ad8604de851f9d9cb75
z65f94778ccd1246425f4aa150663d7c36131bb934acba8c14358eb6df76454208971093b1ec079
z399bdc0306820669402c36660587973e644f1c2e5a7f50a95333f796f3ec53b28bae57f961d3bc
z20a6e17a9b1d56cc0751c1398675ed6c62008aa698799ad4cae4ab981bd31bb0f1af35feaafa41
zf26ea11f69f1b181415667405aebea3009467ca90d151f39d89b59f6aec48719ce085655ad66a4
z54c13278f7cb69519195c45d5004a419e8b70e88011b4c29a3419381ae42b8e229febee7b6ef10
zce1e7f267da621dc5d40dc5065d9e49e117ded83c33fb52de8b540286a272666de62dc2f8b9b59
zb201745dc5a29b238c58ea5a4d1d5ad3d03e11def0f7e1b12776bded07676bbd7ff53234d0aa7d
z017430873f2cc78b7e07aefd8829f4d3e24ab18f849e8c577580a00ba30513dbc70259de06ba35
z9dc7b4203fdf45eabb5b7cecee54f2e0edf970444fa2ba2b54e483c9232610a9a375c03bc343c1
z72aff3a9e6760618c24f6feb81cd31753c1bf06c6883701a11a46a874cde7e3e8afc8d7a0ed544
zaff92956b9cf6878fd275842f5c2e558837aa13b31266c1f44245fb49dc7574f29f6a4d82449ef
za833676225fe1521e6baa8218c6f62e96d14c1c2cac05eb82c7119679e8d067346eaf086bfb4e3
z01e15b7f92b47b6297a56a20be1f316509c1962dbdc014ff00fd0d8316e5f324e66e13618dc690
z439a332d29e287060a4880b8faed0971cf134eff3c443e95d1e3ee72d8c8de668b282b24f943ed
z1a08bedc3851e140d675e96e75c3e6dcab51a0c0ec0fa01f10873cdb1899205441369a55a3a2c4
z44d6bb5e5871e9f9d77840b111c956ae702d2572d8d4bbebf8760012778942c6439c7cad7fef94
z451830198dee260701f99e99c9a4550f8f822143550e855ccb0e26e97063fba6f03e16995eb730
z5ad54e2aeb874a2ab08cfed2aa704408aac928d11a9f7dc2ee587af74af6949a41cec8dffa17f0
z0f802a3bd88001b658906542d02d14a4fc7f7dbc6455706972b84850602a4be7f03728507a2363
z7e331d4f82d5ada1ec1c5faf3900f20e33ae84eb05150a9d60f986f793e5e73e1958a7ca28b856
z96e4d4db6d3d822941d1059dbea60a2ba41c0afdf630a83c0d4a67c0235bfe292e8432fc9a297e
zbde77ebf5ffe932b69c6fa697e637ab3666c2df5310da0b9bff0ead6e75553a8e8e3a3735f998f
z7fb352740daa98f3abca85ead039b31fa0a74d6c34b637a4ccb7b89ab725097477992936fa6ea5
zd48a5c78313da76dc7783915d3b1b178c78ffbf7e0329c4d256c95f6b6d1176b7d87232f9e912c
zd44223d0443c738e6c7fdb74d1dbe339f5b7787914929575811acab8ecbff5f35741694fad64e5
z3074091c52256d62e59de65719630ffb1441dea6a516d14ae4b52e76232ce97b0f09881d1da15d
z5ba0999b1794468f80ede28248b8c945480fd6f347407d075d2bc1900a3910b10da7a7fcd7f108
ze379d6df4ddc9900afb17ac9e4eb2d216fa0538490d7051c5d0e582d8cd59218a84c01f09f3799
z7b337ed4436d8567bf7b9e692e4a2f564389aa5a1376fac55dd6e8a49003559cea94d8f2319c95
z0c60ac09c397ff43e5dfec51d318d384bf055d39f283f7abeea13073138ce0d188b12619796b40
z38e1fb06966499119a03cdc1aa26f169c7ee7a647e42d192c49058d221df856b90570329ca7d30
z38a97a760fab98d077d6b9d767cbe5e43abc9f0569305ded57b36dcb56515b1f665f714ff470de
z816cfd9261ca1c250423ea41d1a0e20c5f71dd65c25181af725d4b68eaffa7a6a8cfa092a28ee2
zf17043cc56c7d95856a9787e838a0aa2d73b85df39d75377514a804922064ad93db968a4419a9a
z620cb82c1431a42eadde3af87d69121b0bb87903fbedf7935424b82281c4f0366d492be5448c11
zd2e8fe24e7564f9bb48b949dccc0b90ef81c3c15026a9920118611cc0b3eb25b0069e5f34651b2
zb5356a02fe49e8aa90c0d254d937b8d1d35990007710ba4fa2181fa45eea51783e35a5eb043168
z30e58bc90f226d8bda55110ff1d182fe412bcf174471b18f08f4d8fa925597cce028b6d1ab8b7d
zff5e5e9556b664a73e2f3d4073f285285535de576d955580415c796d316ec5e2a126ea641064d9
z4a5495a05c76b97dcfceba4cca704c4965f035c678d6872615f0d22199fd80f1f3c09ee080f163
z371ad7e53f2925763a5dd4e930c50c1f1fa697cbf2c283dc1936cc2975750ceaa22f63667c2d38
ze12812eb587ab264f157a9fb85ffd60bd14d42b8134aa71733067e1516cc6a398a59052fda211f
z68f99b39cec2ba74b303f1ba257ac59d8b94fd1797dfc83edf8b52bb39ea2c1186329e86f6adae
z866606eed85ac2bff0d231483acc43daa186f279f4695be7ecd04841938e744edef25ba2448253
zb414910b5a2b499601b3b3e8f31e1b72cd791d68865df0741e814ee7988197b00ec9166ab67b33
z413c11a5b65659f10a4c9c31495857acaa1f57d1cba8e7daffe8e06b77842f23aa50edf957de9f
z52ff7397d5c861dd15e12bdfe16deaebe95880a5bbdf429b36b56a85568ce8b8883dfccd5585fb
zb0d090c4f2545b9c82878d3a561d219c77c70c102f324ce3c893762faa4a1656875231535f0543
ze7d4644707701cc7fed043a341fa762f1cc584b993a5cfc32bc098f31009a600baa472c8b12d33
zde4e50fef5255ca6da83d8d63160ae40b70b711c470dcd26509493209e666c1bd7ee165bf418ed
z4696fa45fa403760040e36e9f29cf2ab6e1911dd44784724d190248fc569be65f185ad8f1fe95d
z67fb6fcf1b1c9c0088de4929b634b02e3395852d32d5ea12f0f7ab20dc45c2a3dfdf3a9a6922da
z462f50cd41f3a9ad7613bbdd2bd4f2fba3801229d059a224349eb57841157f1931cfa49963210e
z8ea0c00788404ed8608c28d30bdd50032d1a5b2ef3beff77c9087c39883e71d4913b7e609c2c5b
z8638b83a8c234edcf9155488c1a798b335240734760aedbd288b94f89442297cd7415f8ae77753
z8c326005c0f38fa9fe2c6c1ae74b80bb75f679485faca4b4379d0bfc8f7f0b710b769e25567bda
z50cb65b4615c3a1378cd897f03f8b42c90a13fd5e4a3ae8653d48b9ee682bf22f784c6908c16a4
z12d37ac3ff9c226b9be6d201dde132ac2f3143789bcae26a240a2c0e7aa096a82ff5a746c6a1a5
z7988a721d5acb7f75a923c44356354b522b76cb4db3846e5046ce61fcdbef0226f897d2672a4b2
z107cc5eb8332ef27b2970dc88313873cbf8aaa7281c6158d4487bd8841b5509e577f887ffa7054
za7fea55bf69e0a0036169e1dda379c40616c0d54d21fa9fdfc5431e58a653d2afe19bf31486c01
ze06d16681939ce4077c1798184e72a1662c28d2927dae2f9ee2cca6beb6a87744536e5059cdcfb
zeaa4a2359d6fba496f646377170f9b52e8a147375f6cf07563e62e4801360877fbc33ab8baee8e
zc9eb3b512b0d3d3bc18e116ecdaeabba657168e029574e15c579a29fc99e344d89a2c89df01dea
z695d541e315731afc09cea4f49d71bb5b5118865603cd8bc0403575fd602fe1fc314d49619d3f6
z18deaac364819c165eab272fb097adfc7060efca68ddf11a53df0978b6ef9dfccd82ebc8f611bf
zdfabfac5a980b64a099657e6772a3fc48e3d0e342c0a11ac49502d19b3b58288df8fcf5473ebf4
z6488fd8125e3b5a568457857cbcddc96d25e74c2cab406a04803b96260a3a389e2f670d88ad7c1
z0d9c1930d3e8e7c79d87e5095eb76dd5b576193830699581b09f7fccedd9c298e2bf2dc6250d91
z569f560a0ea552ed3dd5d935f58ce8b56862a038e432cd9a7da8af0111ffb47f83c00094ef6435
zdbffee1a5498223e8e0aeae79bab06804689dd6efc37dfa35213ed6f6db46a99e99c870757a6c6
z1ac2702d8def125d034ca4c3a5843be3aa8d6187009d3582d9b00397ac4318a4c7dad3879ac1c9
z18679711b3a46f781915a0da6c591efc3089f82777fea335c96a25781d0b9a25be781cf1903398
z4b3e163717ff230007c59fd78a29106552b33d8a0b047d4b390928586e51fd56858b3baa8ca9e8
zcfe76c112176fc8572e1a9ecee9ca192cbc7da230c8972a28113c08dae633fc4f7cc5872d8fcb7
zf07fae94e348ed88c0bf219e96edf158f77222147ef1472fd55b8ec5cc994dbf7c7fc937715f8e
z6c4746cb5a89d1de6435f54002604d49db084bd3771d22f4385bc454fbd593df263587598424bd
z1af77aae5b36b797d070f7073dfd9851c1a8ba64c333f99121dcd24ee8078dc9c05409e277167f
zddfccdf7c810803ac5bd5a81a9d5773bdd15332abdccc0407dd6fa37c771157d9d3a629cd0ae51
z96bedabbcbdcfd6e875dc7a38a33c382df697114f0b3e319f699604ab1bb3cb502d83f3e5167eb
ze5ad5cb3bc36274e1cba7b2c5c0ae562a6e046d7b93ea92538263372b72b2591b6df5e13e39cae
z0c9c7b0a4de5ff2ed87f2f28e8792d8f3c14192009347c05316a3a1cdddae951e08819db5d12b1
z0808d858f3de50b4d1f287032d1422c0b9188fec94bdc5a5a33c477e0ce408101c3e9cab114cd8
z7ef9777ea6295ffd270b93e36ec8cb6d838d7c30df8a985b2fa3c843421bccb65bf7bae9d0b21e
zf2be1ffaa710fc48bf0c41faa2344523cd1c91e8df50e27056d6538163fc58df38dc902c54b005
z18ef2bdd05bea74e7a2fd8ec31ea195c536e83a188a8f7216db26de2237ae4cf24ed1c84f7bbde
z53f7f9417dcf3370c29ab7c85bcfe610dd15f2ed84b270bf41ae9cc00edf6b2e5218796fb05178
ze61987f33b6e582fe9de02774f83175f4b854dcadf33b56397bfab91d75d412aa05629005519b5
z0bda5813419c1d89f14f2983a53da563962a794d1685b88869a1555295170d46ce28f5f2821fb5
z29f6a86777cc9f2c6b83c91c805c58a616c65de5f674b109cf661feb09dfe7e597802c75dcfd35
z880f9a875a4f2fc8a24d7d45397e2f2f3b1b534f4a4d3c6ead3f2f01f5fa831c5a7ad55d4a5dac
z16bd74dc33dee7c5b7960c871a9be0e786849d9377498be3f5b8cf827ca935a8f98d57902f04b3
z3e3013167b564241e344890ca45b6b8149a9dcaae22453dfe31f039b02ea00f77edcdbeae56273
zd74a391fa19a3ac94f6adebf6ad3076890eac7dd91822c1f96c1fa306dcee9b2b6f7cb65afc126
zb0ffce27d1e50132c596b7047a1fc2cba66b3c957bcaa4a0e0298cc6010f00494dd97e63bb4c26
zb1ef142c28876ee8f924d0ab94e257e5b28bbce577e64925fdf2e267929e5b38dcf54e41998728
za6db11b1c08bb82646909c25f66db3998883af0fbd5b17e455e88e539145f704ae6808d4593045
z89035f2785a936036797fa41545561d46e820bde0c88f07f3d29e945b2eb7df277aed1e15f1306
z5fdee5405d23837335f2f98b574deae643c5e0dc531dec793859511a7d882e7e6197a45cee9ec3
ze6fd9205612edd0a8043d0704f4ffab617ce45e1973ebe51d11aed31ad99069d529d54ec7e3ce9
z7e362ac09e1a051ed22cb09eb10823468bd485b514f11d84011b2a2d66dec0f9fc842cca0e8d80
zab1b56d498cd2a5f3b5f2f0844807b79cb0fbbb9b8a44ebf9ef4d826394a40c732ddf5b5592b20
z92182bea108c4624f50512b7577aa388f636c61c251daac49766f41bb4c4f27a5d4cac0096c7a8
z847cd2250d967468435182083c5089d3b713fed92d56470c58e9a150cea88b2e083fc74507d4c6
ze30a6de440921bc29e015cf388abe72f83f151f2f3c32015589c94928f3c4003e4560feb49706d
z9a4d106b5468db8c2b91fb6112b9f4034365111f590c754f16a65d38a05ca55a5606ee18e170db
z42cb7cb228ecc36be8828ea2dfc294aa8f0aa8d22d634652fcba2feed61d7a7769f16aa318c4f1
ze83e6130accd15c33c4d39d0410cadde15faf958fc68cdfae1247712fc0d9174901ddf6deb52ea
z1831fdd59564716035b4bf4dca7f7dc73efa1e073d7a3c5b07de7050dcd0237499d77562f973c1
z9177a3d98d84ecaf82cfd7950e6f97f7a3b523cf1fbeb5977670de3c43773a271106992efca676
zba6a4dbc039e3521128e0c089cd75ab1744ef5c0c31580bac01d9a1c91033e203ca94e6e37a4c2
z09debdab688e6acdb3c8df2a77f3921f1cb209d789a083678f98c454206ab041778b5d7acedaad
ze3a30d1da9ff64c173115afba4d151029e17139deb73c5121f6c7368666a10e0a90ead84c087bd
z15a224b848d9d05accc57cd7f140072cc448e07056f3f1cd1b21d9b30409cca7dd8dba09d448fc
z2694284d91d610dd1450feb50d13ec6c474bd99d1cb93cecf17decd199ac67f53b81514243a0d9
zd0f144087917be072158df1f7a5ad083c0a151a7549e2919acd56bc5b9e93695c0128ff282dec4
z7e8b2890a1504f1535c0cb87e4f32091a06865585b9b7217e328689fffe6cbcbc0e27cecd70bd0
zebc1a765532d98acb70c158ab6f94a5a8e25e5dc08c8a29e72350a4c727fc922f765fd446c9b0d
z9292fdba8e5cd5f3b4b3c96bc4b94b46d0e9f33d4ae37cb0f9f8dab784ee5e2252e9a61e60bd7e
z0332fe41b77fd055630a656230052b40992ee79fa74d67a0e0749a33c490fcb6c0b370f4c5b195
z1468d9b7342f0d85ff07b312614f9a92e76175f294baad2aa259a41d79a3f567f2823eaed166cd
z527fe82fe0beec854a0f88648de09b7ec83e1698413cc3c6b282023ff4726412b7717079e22233
zc22b0170c9847c56ad65d80c3ff47c87f2881c256eb507c403805b9b889090ad702b1e4d25a2b1
zf2a7ed3c7cf7017a99b0691d3eaf1f0a83f5fe1f600df27bafac2ac5dc7fc118add243aee1dd13
zedd12899799e61fb00348051c0e4c75fd0d4850e28bb09a6900726efc2bd0762903a546b67d396
ze48750d51ab2d1894ea48d9741ced8f9d32094a2f79d57294e212e4316f0cbce9bf4154b797e25
z1b6ce610a16fb24f4ac13359460451c5d1e62d4a2384c5de2eebe7d6f13bc7b282fae9d7511fa4
z65564d63ea27eae31fa70c65c7fc0fc2eb0e62a682db918e5e778624c2db88d67223d76b9089f4
z4dd95ae695a53da1c9bb8269c1aeab8f3713d669ec22e6340f3ed541b0fdc1a24ed2c322df331e
z0c01ec9ae3fb0011ae3334d50c4b51d0b02383b512187aa50cf3a41f59f480ec14ebb34c3ee86a
za7921da985d54ea3fdad000d7f2fba073cbd3d780e06941277bd678fcbb62142bb79b0ef97aa0b
z2c0905174e4e1250237545022014a1e4997e363f84beb7e7fa7f6f539736827575a892963cf73c
z1a4b20581fe68a3320e2c27fdb38d51d8d9e01da7d12917bf45e3425b28c82d911f38031d0f1e6
zdc9ed70beb8ae83f62bbbcdaeb505faa2943fd3ff8521622836a75ccd9c9744ca17b2af47902d4
z729044ed31804c24383152fce2304ea6ddf01110723398b3969098805794c3209785bcdc893870
z2679187a84b1e724b0da2f3fa8eb98be1453a240d665ab77a665c4729e6a699def74d2c7015314
z5249e16e4859e4fce820abdb3e56e8c30551c98cb3fd81bb497876f3a9f9a7efcc266f60b0bf87
ze13c61a009f342f53203d52b03eabd6a4b0ac15a2331f2368408f7409cd28255a910ad1c069435
z4a3da6c8e50368fb3e27bc0924b3d061fb0185fdcf5d05a7274c52315f6ab18bde15ff49831ab3
z4a985fdd9984552352386efd2c11e87fd1c035021a4cb08e21a25c0df6a93eb15c09de858bd5bd
zdfdadf167cb058f503ae0b8dea32b83831edaa15d0a592535df22662acc306ae5fa7f7cb23b2b2
z8288ca2ff6824cc6c9881f090f7466814f97236a41313d3699c87ba17b05f2a1d8251b73182a44
zfc9ff3c9c4335434d79c5d20cb48acd1bddbf932763ebc008852410126dacbb27a182b1f448f41
z2107fab86772e6c5fa3d56307730dd3548fd7ed929e990d393f29c27d8bea5d8b7fa689e74a876
zca87fcc487f74ebe4b7fb3aee81fcaed50ea21026f85e394c5762ef6047df1cb0256b23d37fc1e
z14e95c27e733fde3135a71e5bec4165f0c1b96242c62c5d834a1db2a11542ad7f621fa9c92c047
z0f4cbe6ccaa62d0c84788fe320a372086a94b127033cfd924ee771f0c998bc9f9990f28727500b
z4f1378b22ece03b8c614c945146a2f7a906d2584453a5dfa78de0c17ec476a094b1da59412e1dc
ze00aa6f238cd2afeca64eb2d56191bf85c327ed1fced53d89907c7b85a02b18a5d1fb12d0cecc8
z0f6184557ecb6ba85cb3d37d466618491c0f3d6f6bca4019dc9436702bfe13060f06664d6025da
zd38dd61841dd3b8653616fa986da2ec63b751d94835c7488c693d2a5c80d13e92b76bd67fe5c45
zc430a841fe7e59a67ef850934e164b1aa6983603da5f475764211aec220fc5745bf3418585b808
zd93961942aba90a6a0a2837a45456a444c57cb307451e507f6dd405aac454fea9a21fc17016af1
z8d5ac55325ecc641901cf300bc8c31c46737679c09d7a42af5af6168ea08b264731405476dfc18
z11eaccf0743f1452f4fdd9469fc4bff44e83a835337567be329906069375ed9aa291e31de6b224
ze2e3a71fdf17ca549b35578a70d5838a90d38dad884a174a08ceec880d453fb8c285523bc140e2
z6015fa967ab72172cf4acb7679fc9eaf8656c86fd49234d8bcbb5d33e56fc77f3a09dcd66b6eec
z34154f2a0f39e8c785206c58b48629bcf44312e8f25a2248086157d20448835232f6383e6ace0a
z8393e4dffe4953cf939f668aeba3b787975f04ac4b5e2bcbac67705cecf63000da3aaf9c0f29b3
z260b46c3ba7c13a15ebd62ca58c9f9a0473c79758d0389ae3b32c41ef582edce8d0e2c5b31112d
z3c432f1c2a91a6ece0d22e708d3ae6b073c15cdd3393d3d149f2eb51662423bf4b635649d03a98
zd06eb95091450862c27c69256d61f0f9f62e697f25f8c56bd216de61823dfd706ca9110bbc3d56
z5c1d4e8dc071b6f1e765557bc69c2ef49eaf6fb19e01dedf37333d62bbc1bc696af3d26d17607b
z25e0d073f0fd7518517c1fadfe8fdab7245b2ae71a5a35380159d60771e1ede8710364951e3e9e
zed688d86df41782cd4ea7687082656ab7a49228c82ac6655d4ea532533ede8ec9e29aa207e7c5b
zf909d4de1c6e7d03b3b2c8ef7d08f5aaaa92c7876f04c8ecab0c42e91c16aa6ef930dd2ca41d9b
zc8a72e732d1e1892d0fbc0bb97c60ab74931a0427a1da79bded3bcea1022743b3fb4bde7eb2ae9
zd151f169a29c2bcb3e63a2cfabfe8e62e2143d9dd157b980e0ee6bb39f4740c64ab33526deb874
z0715729ce16bd23afffdb470e59b8ad06145fee87543b597d452df26d8ddad9c11047d1372f60e
z6a236b5a29dcceb42aea38aa28617050d52c6a98a388e6c3b64179c70fd85c7e7be95677aec515
z2dfb1ad0e44694875438c4349b202ddcd49a43df1a89eb5e6c963517f2e26aa550701ffcc364f7
ze64c5a23ded78d5c1bfc941a58951eef1fe48f73b5cd7d43dd6629ee77160e09cc68e5143cc7a1
zc9bb0e0829760997b6fbc08a5d391c144226bad929c2db300822cbdbce8494a1c2e4900633f6c2
z13d40b0456d17bf8175988a96906ec2be49bfd5ac7e2383f157da22339ba82f5fcfe07d3a6a632
z776acea1fde15fc077d5c2790256b7bd0aed1666506644eb228ab9c1f91c448b3064dfddcbc88c
z8da6a085d2b80ffd8aa4c222e05706ba384f656e881ed289bbc5acd3ea0ad5f40cbd852734a63f
z9ab3738576b8e3a4dd35042348e74145d40b537d2b74531fa9a457c3544239f9a5a748b959b74e
zf25f2773f4ad78185dab9d3c40ead20b3395c087c03ece99def00fc5bd824b7abe4909644bcdbd
zbbe841e145b0698253ddb1d515206e53d63c54b9931d6d48fbe9f7c14fde3ee5d4ce6cff1cb081
z156dc08ed30af853019bc4e82b30c36541791fc7f0fa3a78be203f06254325316de5c40b594796
z485ec1c2ff790490d0589e9bd9b1c8c3d8178e6e8c761cb42bdd8ca99c9e0d894d26730cac8f45
zddf8eb9281d49f5f57d1287a7c83cca5829f886b467a8b0713c3cbc9f50a306804ce1d8416911f
zbf559717331604515637e1144df1903fbf7eecad1ff02596fa091893bf8f830d988b4a1953ea92
z3f22cdb8989ad6c54a358de5b319d090db7796ea000f2f9b146b24850b0dcb113f14c06b246861
zba27dd79895fdad19885cc6a5cbf78104b085f4accaaa84e7f7450423661baed0cc9e7713795b7
zaaf68b974f46f5551f21f4af7a17aa424f0d82fade195406757c3a80428d241f2ed40977771850
z22121dc2d9311ad6b9d9adb30b4f55d60fc6da7c9b0525ea80d17e24e2b399fd7832398d577386
z1b1934add832d3f72059018268ce14d8b4ae9f9c236340004448971bbbf2155d63071475c442d1
zf0ec29843374f6b8d776a851d9b29ed584cda2a28a2aaebacd69858349fb70bfc04faf306dbbf8
z5df9384dfe38523d1f034c4a64c0e2e1c466a294b4051639c7dd9490a88dbcb7c6c2d4b096d648
z5974dc0c7b6ce20c6ff8dea19c5f54437e84f1861d092041ab31d37e7a39070653d8b9f5021490
z27d97a58ed37afb6cef025422d8135171a56fc2fc0d1b51d12fe06fae576bde2952d8eb0f0b8f4
zffe3662aeeb75f0fa8ee85bceb712675369cfc184e8a0421c811711d72b5f90964f993788d133d
z146267f5c9dd99c336dcb94e7cb777b59fd335efe544e91f88f74d00cfd3c2176947a55a7fce60
zafa29b2577054f188faabab2f0cc747caf35751efc271a2fd2c46160f1cd397f89f28b4821556e
z6a1b024b5c92a66788f5865d0b32dc714cf68bb23b4d7d2ed3509990ff599a08623be44e4f8ab5
z48d88ee42cc30025ad1cdb1c35f6d8cf4f7d632d28eecd038f0cb9e41423296e498139913ea79e
z419e7587691fea86800d43a1864916139fcb87cefd77c965db085632374fe3d8ffbce2687817fb
z6d0efb100502e7359fbc39b830d9df7dc79944c30d95945f9283282d638a8378f699af9cf89183
zf5900e6a6b8956e12dc5cb6665be52a2a812cd018c196f2f48977aa14167194ac547b376aa53d0
z300efffd1f2f5df333a1f584b5366c705555abaf9881fd1ef7899af45d56769d15002c7a21ffa2
z9469d00311e88ed4d7eb61d6f22254e006e06a6845e7f1180e0752c0b9e5501d3b1967d2a93ce5
zd939fdc6be7a9b3a307d9db205ff477aac4ea22135b320c8e3dfe7a58eed808f21fa822803a038
zf0060847b2c828c164471a7e4192b4779d7b23148defa7984283bd3e890858aa113617e9b0dac7
z324f4b0a40ddaf8c79549a9e6a1183a50ab9020a225ee3dc39c6c01dc33b2fe93c9d178c52c938
zf05fbea69ffd3226172070bc4e37f1174b7279002aadd5f6f4ad68633d0a51e88b8842bf0dd827
z73793178531b847e552a0a37f365858329cf4877b99ede669edc9d76c39772e751f5bc0a620189
z795b4cb8383671f186fdd597196a2630f91a6307ae753b0b6c9b33c85663e5086aa7cc15748d5b
z9982fb4a0d97502960a3e838a6ab31a8eba684c6b06c049da9abe18490b5c0ffddcb9fc0e2ef36
z8edff853fbea43fb6b4b0abb127e2f179bfe9f904781bb1791d0538fd9042a1bd4283d03006d7c
z2ec228ae1f61ab74350255038501250d7e22447a98c88806fc28deda0dd877fd7e2db53bb8cf66
z65903dda90cdf0d5cac0e318bfbd00befc1b48a7f26b653f26d7d550b0ddac6b30f392257a142e
zbc5753d32b0fb5775b7defc5d77250b93836fca81b4add8a4f01caf8e6b4eafa7f26411b9676f6
z8abb8822395fc498aed4fb4c9dcbfa6c7946ff05abfcb2396e3cef153539027b3d08d5a72d0b50
z16f8721d4506a68ecbba1efa5b6482c42c0055ab6d0e52b3ccab432a14e55e3005faf58ce8ec82
z663b442c5240c8727fd0710c39e4d92072e6a1bf314b44f15c6cac4793c820750a6859efb51bb9
z9a3a3360946169bb4a469b60983fcce05036de7e685c7a780d1f18b09be821d08b72c0f7273d07
z075c3002e9d59c923348f5eb0bbdd0f06f83dcec285db6d4a307fa0166da82689a546a7a3d7170
zc0efa32aa57572a1a668dda474ae6c50cc5e7f1a78abb97b880e996c2ade7eb3ebb78f89f8bace
z2663bb55ef8f964f0b6a0fec7bd2fd3065dea163286864369792c6c49d514d242888b2793ae525
zc18098e48126e8e509af87ec8acba03c473a3d1cc40650320d510e56a8d4d31498dd5cb040e369
z6a5ba199843ef73076b45190697c3559253d730b5a344bc1a9c5882ce593ee847a7512bdfa9438
z391ffabf652e418b09828f1f168e7f09d8c8e4275f588ab6bfc6b460a448cc79fb93bc54c5f1e4
z4c9f79a0dfbd4be3706a5adebb0320b5045746713e56f38fb6648325bf2b5b1d511b1cacae655b
za69afec2259082968f8844d5e7db8feb7b07cf6ca9072140af00e090db56386f55bb31f923bc9f
z71434b37c996ad0d2f59efbfc7bf936fdb52fe6f783343a5fc363a9b7aa04f17d87912c9b597b1
z56bcb796c0431cd3a2f4c2bd3a2aecf4acdf4974124c2ec6cbae8738580bd851f8474ea532407e
z044b6a0e026bf3f3e153f4df6b635810cae9f786ab68817ecf84612e712c29bf8a466a616a2c59
z3cfe22e1af9c67ccfdc3ee76a3e113c227f9499e11ec6e00dbd739c6f00eb60c57ddd4176d2f0d
z38fd90090e12e31dbbdef4b1472f10302030a1b5d31643ef4a98cfdacc85c46bc811a137bd76d6
z0278570d32d236ae6ec566bfa0caab4246a732d342a6e1924429fcb50264aa617dce6bab06b9eb
z075a08c42a3a5ca8d246990a00d64b2678e35934d67c2c0a125dab06234289c156a2df14ab2a1a
z27871fc91461a9da1c54a7ab0bdbeb7e68d625dac4cff0eafa1e2598eab9e6560db84d840e3f7e
z41682229b883a8a9575c1317f9c826bab544c7adfbba360413853d18cdc168ea81a44751fc0141
z4571e655afed0618620e3a889f0da8cc6b0415d7a89158ea501c0171b5bb3041b8887df83d7a2a
z25a35ac397612c8ab262b095d9d6487e287d7dbdf78de9d7cde3a297142f7a35ccf0131eb814cc
z4be958b8d44c5e33a692397dd411a754b78f08e3143e33fd10166e3221ba1b2825a7e0d3232f78
z33bce1daae1e4acd2e2a2d231c62c5de846c56a538d29013cb9ceb6e593c7359dc12fac71c0da7
z4101f3d5c255d3765002b8692844a98ae664120e9f92e934cd224d87710852e5abf51fafc0a564
z1c7d0670d4d05c61f90b3bacd2fc21b3bad4b473c741151fef99a999bd4cd71b744c26f00eefea
ze0eb2d0f7f81d2c42cd201fd9be0ece4a153de7d59cf5fc00890b5f6475ee8d5ed93f14c31b2ed
z3d9fe3d02c1438ac0287341b509d8587ff8ef56c3af5f7dde1440c0e970b9cce4465e5b98441c1
z89a1b716b59504906234a60f5e9c77bc3fce444bf91519957f13a7e1cdd35e8f106c0dfd27fe9c
zba9d65f75eceee05d5802a794879dc3cdaf6041866552e7249639f6728be9632be6223b04fb17d
z421d2e3ff4bd474f8d1d06cabad4018ffcf11cb551bc066e5f8072bb12bcbe7bfd538363e8bb30
z9fdb0fa890f3b3656f72ad2d50d08b0ce8a6bda4f57408536faeeb0b8df2299d3fe8bdd99985fb
z459b329912fdb371133978f7c0756cfa0a8fbdcb81c902ade7f9ec6cb15f309ddef18d147e90ca
z1877294e099a26ea758ee47f8be37d4c12c7b3b729937000199de00f1fb05d1440fbc7eb91912b
zbe6efe978259347848b9fc287df9ef06016d03f023197a2abed42ff7d30125cbded81185e0982d
z5af6df0031efe1f26d601b68634d34354fecce7b624b0d51c3088ccabe69cec0303b5d54fedaa3
z46426d36ddc03d311d3960b8cd30d78e790a41b8108e202cffc7052831dfc764850b4839ce2aae
z9d221e19bd752d4d573c1abf56cf7cc83ea9ef60328f2206377e51d0357d0b1049902118423c62
z4a2f528980e1601e98e1c9ed8ea1ed35fba38ddda08dba54c1025b3388b0ee21ad3c78ecfa3fe6
z3ddd73c967988c9d2b97de223fb7b70a97a908868f52e0ab3f3053176afc735ed2e16f779425e0
z141e70a21ec9bc5b69abfd19745be240f0574d0dd7a49d0c3424b97ed1d796e3b2bbf324882810
z766b59ef98cb94a9f1009d0f13ac761e82b50d6c0ce95671d7864f9b75705b260993a44ace1021
z253817630ed775142683514615691472edc6f3beb1bb7d1a05bbe49602fc677de1ec084c5160db
z3391d2d17e40485dd3164c4ef38a6acd570986172036460bcaedc1284cd136d7bd1494b28160d3
z3988868bc3f781a9faaa49439b5274393aca33204be4f4c281493006e2c35b0d43242fd135de0e
z2899266901786d6a85b82971f08006fd63fbdd4486af8fa3edff6156a7e4872d32a804979e08b9
zb37b6f15e9625bc4f7cfd4d279b54724fa2551ae5e2ed6fd605ea1f33e304d100b63d495df06f5
z2a880e5867f4b2dd1e9e72275e47e789c729d99d06ebdf70f3bfddae1d738d87e46ef3c7883d2b
za335c5b19dcdfce77ed283eef2d15d49afd1409f6871c1a8f47b08be3eda79590da4c7c0dc324e
zc5d611ff1394126f33f8209bd484a631ab9c54d0ee7f3136cbe936018883b3896b80763ea3eace
z45e74b33ae1cf63c1994c3b72635ba561894c4d50b35b709614124e1305eec1b894472a3b8208a
zf5b3f636302b95839bda1c1731522d3f18a92a7830702d7450655fe0848fc476404875378093a7
zeded27171360ff840ffd6fa4f535071f44df5b058c5f8e382efc05233d9769035e3f5cdfa29c74
zf8f8df35a1c0b2b1df7f8833d6729764a9f9a2094ca3f162b402499ce63030fb13906bf87aae37
z6383e7e6857220041c12958947b92fb3411abd443dfd3c6bce79fa2719c2017a5aaf41b7d06b93
z586157851a46fdc9c0bfd2f6b715f5e034ef48d9e4a10b0742a1ac78524670247607a72973b1be
z4c261463b8de4a8b703e7e7fdc33da967eff1e37c6a7e89f99cd71a589fd27911781514e2d1ef7
z955a94474e5a3a9325fa97489d3feddf9afff834e4d8da89dae6efd70bed68d6f3e4ae538d7e99
z29380f357c4335daf3c06b5310771b4cc5056838d4e0c11a33db0014d418612069b9680c8a41fa
zb548d37f882734da9fcb40f98e04f7f5365fa26bd90824340e5386ca281a7f67e80d844c859bd3
z1647c7fcb9ed5d04372174981c75b41121217a402d2ac05640e2092b1e9e28ecc7f29280cd7b0d
z7318edba17c9a0d6fb886ed0a3e48738a5969558559b457f30e72beb311b79f12e34950883b42f
z1f02196b5eca488a50f3e93319b7603b8e1ffba93e4b1860850beffa158469bdeb47db4f604e53
z03a6e1467b2c01df6d6b2421f4331a6a4e7a12fc77086d2afd65ef2e203c31098aa76200787d17
zb086157ff9c490ef4e947401c5d49563b5c3b2ca2e1b8af8b6469bb1b13fafae90c872eb1f8a92
zb8e2e123a735328c1bae415536db415321a61a615b7cec638735a5f2651f9ff9e176945885a717
zd015b5241874f9742a0483f3fc23298c95e1a31adf2996a34a81d0cd2ab8a137b99d664d097b04
z02618f38ed73f84531b723ca996bdedec37f98020fbebbe2bbb2b583b68939b823550ce769c842
ze61a336e258eadd3c82c45ab73dd1743aa2731f8220364d362e6c23695317749694ad8fa6ba126
z45a2d899eb853d5e17cb8c5914ac136ce433b51f46dbeef7eded9370441cd60762bde01ca0a58b
z7d907bb117bea81b24c87c21c8a84792a9b551f3bcb83602167f8f94960d44f2c901f2d54590f6
z51f6509ea20af5a7c54590979bee0abb0f6d4cdc695d4f8cfdb52f1288929d33597d346a798470
z574d8987b638cd058fb5656878fa7ea02ed51dadd3496ca105f3b8b3408e55bfc0760abad48135
ze8ddd1992c70fe3f7fc1299ef1769df51065879bc71fdab9546b4779a9120eadb341ed40a29c48
zb15891bca8d1e73168b7497cf0415ff8e8cb132e724ca3d4ba7d93996646bfe3f2728edb1f3452
zeb7f1cc722537bbdf3bdc44385b5da3801e0289ec008443d45132d8970f4b1685813b60dcbbf98
z6ece87f0559124270f3b68a861b4ec2c35020e64ee2c91fe5b9e69de7a55ad4e32cd5a154b2cd0
za5f5a34af5d2fd4fe42a5285f9cbef8eb9f158e10cb720d3b3ba5d34337f3d40dce3e4ee340ea6
z18c56a41923c556f8d8462a3d47043a3b092f41dd1ed18d712ff035d08d15cfecffe1399061212
zc61891a437c84498520f8be3bbc8546be5e5949d333580f3d70ecc94cccbc9af9907493321fdab
z8c5df9066e846f638b32e194246fbe43b58b1977d7a9e272cadc37f23b66a615bf7c0bdcfe2ba5
zaf40a0cc0ac30ea9059aea3c3572e901e289083d59741b2afde2ae8265cf4f0b9decbddbae07f0
zd0beda005882066b4af6fb489b9bc7ba17d9e8f388f1f0bcbfaf7c3b0bee397876a1f630a3beb9
z94cd2ee9026acfcb58291b3b40b0667ca9ccce67cb3da7450873d76026b4d33c65d322617d494c
z8152215fe0dcaa3678da8d191455c39aca9eba35e6ae0ac2e35be9ddc1ada58e3fe13b650007e0
zb51f3c67c7c118b7e80bdba11146068bdef24c67a9eb0e2bf7cda139740b73f7ee2f4d4456b992
za50ca1b40dfb76511b406446057cabeb8e319498cf4cc8906c85cccd08fd26411887837843ec33
z5e224aaa718530e7b96be9d400bc739449b3bcea47d4effd6b748d0053183544fbb3ba398a1c7b
z25e470d6ce039e6a4b5821e2e47289c1157ed03be2fd0974133ee2f564ee3893861d42367dcef2
zee06c3a4612336f6d11317c722908cb14c15154b293dde97ada672e34d7f813928c3a2600cbf99
zc4e72098451d99dc4634a688657b41ce0cb620510e8bb94c8814d11810c6b8e4faa37b61af65b6
zfefcfad4bb10ae3063b16c0e155eae4e4bf48091d55363c4e9ef61275ff3ecdad7e369d5508c21
z0f687f45aa05872f8a0a226a429e9d69dff854d0a2119cdcddef9e4b3bfa539cd4ae54c6e9b139
z54dc07db55a41d0a4f5c057ac4811d610209a3cd9c3f167e146d4d49f61e65aa561c8f917f4a04
z4612b1c30eebf61fff8a1430acb592569fbcc9ae4491ed4272f9117c9a4ed42a51b079f61c5f0f
z527e65c48219d62022bb146e8c8e26728788adc77e3e3985461ab2049861baeb425e61393c4edf
z299520d6128c76ec852bee4e1e125afce3282a1781abb60e04130765317e391a582cf5e5471ecb
zfe502be1976274207b0ed53c7659fd85a469251ca26ac4eb023c67d96ffe144d1b6dbdbb866c6c
z81c81eb8b40094031076ecaa2b840f68729c5510785722c1f69c00da0c4fc04971e8532f74a58b
z667bbe87470f00e8b39847f86df03e5e8190bc49ac4a6e68ea3d7bf6d09425a4e7b342ccb0d227
z5d490ad85a123853f502b53fe72fefb31ea0d6b813655a2b06e2a63aba18d6981a229a003183ba
zf78d47f91767753134366a28debd3d20b78eb0804aca49497ce84c342b2ead982ce68e89579101
z7162cfe80911da3409f1f51f55caff5ea45bde2f2662f84abc84f96bb4cfbdfda22008a0db741f
z103a7e04ccf9604ab5dad097de886f85cbb247c5f08d17e4c94472f7454b3831ef1789df09aec9
z3b0232401055850a453ca7d6f3089c3af074b74d2276ed6e48cc76f9546b42ea109f4684dc2f75
z3791a545caed5e13920c46755dcfad6134e5f839a22f61352bf219d40337910093726f25831e76
za82fb4cf97b165f2a1c2ccdd005732cd279315ecafef16f51c35517c4f562497048641b199df7a
z7cfb876282d74124a0afde67645964b978d77155652c2d3551f92a1fc74cad65852b3c85d89d89
zc63344f87e7b8635bd141e178b4f807f07e1d1c397eb891039bc02ca1ea25746d4de98491c516a
z323e2771e4f7971b3b7a2c2a2fe49c9baeafeeffe2b39ce9f5c05aaf33fa8788649c87cd6d6c22
z4333a4a27404c24464f9a2005034cef9b833d41463bfc8b9f46c3775c3118af19b27d97f5bd3e4
z0136a2be7008fe4794f163711bfb2f69128e3c6c0eac064eef276ff10d21113523c7abcee2f2d6
zd523b251769f36bbaddc2ead3c4f0b06ebbb5247ceabe42f6d38fa507f2d59558453cfdbfcdb3f
z99bcad8aed72f7c2cc84c8176df9cdf025ab702f344e1a72f0b6d564a99c06f03db118e8ed1b7e
ze377d9dfcaafe77f44525a656b093e819ab249dba0756e1823ec70e534a2b526b017dc7142aaea
z642ace7aaed16465d476bf7389d1955105c778a9b45f16d0f0b2532d11ecf5a423ab442a74ecfe
z8259416e4f98312bb5d27b6a73fc6dd718c4cfac59e2ea27f4e4856e41a645657b56ae643f2cf1
z3e51589a117072dd58307ea5efe826da950c8f39bc20e3a074d3141a04c2eee5bfaa0f744cc543
z97d040e3b7cf26bbbc8a2b32c03c9a5b2ceec0e56e7ba367a1f30ccd9b44024aaa8151ddfbc5ae
zfa46e0586f9bff11160631012f2b35039db5a5c7521ad4fa06ea5ab0afa6202de52b45b4873f18
zcfaef1b68b0d9681d529a98101fab7c17c5407a008513d91f9398e1c3e2a8c5afef0d9f4204a4d
z860e2179be0a499f70c1eb3af19599bedc23b3062ef0def9397fc4defe472a54c63e6b6656bd46
zc758a4376ad66622c4735a29ba4e45906d1ce431bebce8ddfcc476a0056c621528e543190f3796
zb8759da0c11ca19cb4c7b53a7f0fcaef84eb7b9f6ffa38986e137cede7ecef5850cfc69cbe2dc6
z09843ff1959c0c98f8e67b584b1e029836fc40f57c71232e8cdedf523ddde6bb42ab0e9552bc5f
z177c094d4f4e57dc9bd30aa4e92b76c3b430b87c2c25178f8f3c38baea4a38bf1d6963aba76fbd
z7393547bd54e76e629537f8ad7594219f840912690ea77a204f4cc7e7f3d50afa1efef18d2a546
z5bbdf11cdcce58848a14826562354bfe7e7d05da3cca51431fd3c978d04df473164f7b94aa2822
z8e3713900871dedb5f7f75dd746576c930b08fa759b734077901b45e84fb6cc266bc220de3be7d
z7704d35a952a9bc9ff463db1a44f9ecdb7a6d2b2f8050c5d4b90397f59c547c0e68dd758aef4c9
z8224453a12d66f02c3ce67a5a160bb93d25d6df8d273f6a0125c027353bb44a2600b7ced22b9f2
z40606c0f5d09905b05bff2fc4c2f649d1cf1cd23938dc28a58afa21bd13196d40c1d49e9b63aca
z15bc11fa2786b86435baf553488bb320d84a9ec3759ec97f4463555143101c7d38d1a6d3325719
z43f46596505d2c69349996e487a379fc1133e7aba67c901e5c9ae59cc0c90d3e2aa61cb487d063
z055014e539defbb86354e9200183d60b3cc5c5f71caffc0aa9eab604a684df76be7137c8b0677b
zf6c910d7bcbbbcbfd5a260d50b9ac32a15e9debe7bb6a9647a99910df029fd97c5e2bf7719e1d9
z28ab3778b13e1c90d2aebf0f8ac579ffae07397c43e77a823b24b7a47915d82b50f996aba6715c
z4e7dcf07e12d277c14085bc4ec152ca04b9226e4e71d31fc6bc413ce6ed0200c91b0b1d1b85600
z96efd95320b6ed9bbe1735925931c016f72d6714e839b2b789aabc0ce575fb274cb97eddfaf53c
zdc68b625e25b407bee965957729dc6564f3ba03e426f5ae24eb3a18e1ae0de900bde502520d8b7
z00f1bb8d8915cc7dcfad8af524ad66ba9b7f254e69fef88a8e2f7ba96fa59812faa4766098597e
z2d038e511750bee629c76a9951dfa8f2d17ef3cac8ca03ceefdef7af1784e22f71b0fdb4a395ea
z9408dfb6776d55c6bc9a7503fc03d63948d7aa6e68ca9cd53cbc91d6dcab4bf391f571002eaa06
zdb44c59fc9108fedcefa41a5f96daba6d6e3f059e9a39aac1265a5fee693d86d62c23e19e28dea
z64389899b68a007fabfc3953dddbbab0aa484db6c951d702c209ba2912a602f677e1d36605b131
zba22e29942e1698b7c260eda4f3e748ae5d273b0283b7446ed933c161eaab35ca280c8434b1df0
z781ef3b4af15d8d19368fe2f31d1cf6c4ba4ce5e6c7d1bb7da496d697969e10ddbb630c5919fc2
z85941a0b0c1970b45d824a4b4f30144b24b74d3778a3046fb65aa40ee567c8a670d13d27e99bde
zd0651ab6d5e903ac6a3b31d06266ea455db8f1eff05992b88dac200e7dbec1137f4d6779f0a94a
z858f5480bd9c5b5e6736792e73f555f01dc531d10ed5c50c992e1d095cc80eb9da92234cedfd5b
z12180158266b0e6c9a48e16c890d9f116c32e7bb9227d00661272b5b812009cd6048b7c6d713ee
zf0fcf241b3a61be10d7c0fccd4ae300948750b8ff0b818b24166270c58eda5e061cca79a91a43c
z13922b88564083f392bc34dfdee2871e1fd2288935cea7aa51529fcb42e8c32763fdb2058f2316
z8a66ed0c72525bb017b075d0cb3b196b503f56a810dd1465c88399493c4500d42863a796caf94b
z57d341c9d1e6ebf4977b11e8e990733031e59721b541793b732d20befb09eab65e8645346b2343
z3c83f443eff6171538ddc452082f9b2c1421d7e9f5524460b7eac7ed56a2b4006cc845acbe709b
zfffaaf81fcb0475468d8232b271d69e9bfed2bb40d8bc15fe73ecc86606651773e5671357b0d32
zc926e2aadaca6fd93305e525be3ca35df748586a4156ec051a1289d33d3729274098288aae9d1a
z40c218282fcbee6d01925148197d99dcbca0bf9e887fb74c758305ba185807bef5129356cf0517
z73e9ccedb7fc4952b3e903497a077d2c5f3639cac32b569624b95d720dd510334377a50e093e4a
ze1b886f40980a0b08674e28da346c3210b3edfa073ca99272af38bf4957d630be05835944af4be
z567942d1592f7063dd322bcf8c56ba9acc324038c8b0b2d90fe6c78fad00bfbe169199a209179f
z730d342fd39925380ab87f94e778e53caf5747dc8aa94ddae13422a6fcce54733c88f5e346a9f0
z26543ae19a0ee7476a2aec2debe8508595b41650eb2b77d2c8b6eece32f2917264b0e3e51b9c5e
z02d574b72ca690be9811190f1266c375ff7bae3abe1b9ba55cd09884c93223cd494f64b4466b6b
z498cfc5f2820cd0882f3689a2a5e96cdf38c07927f5eda09045aae23b91bd9e7de4fec2b89873b
zb122cfb7abc30441972a88ac87c80c561ca4e73843902aafd42461f5f8d3507b069b6fe050fbfa
zeedcda1e6e6a912ce79ec60938ab16449bb5595594b7869aebf2f38b8a4e45eec02deacf40d3ae
z7a81fba93368bd7d10576e5c921acbe8817f0a92e8984ed01f597c455e3c309cc655136293ee0c
zda71c8c902eeed83bca22a9705753ee17305c98d57de097c0ead4ed5587518b4d583cce3447c62
z7e7c7c712ad90e47998e47cc7ef7eec68c6aa37eb24ec5544ec5ad07db0d224f203b34b22c5ff2
zd41bc245aaa6dab6471a014b91326263b501fe48d553a4c3e1dbeff24792a94161ac2222af38a9
z81fcb374902db2b68f00537cc178e311f99a305f582b255ae3d550a4a91e4fc5bca7a9570e4f4c
z7e3082004a75f976fae36098cac1f11d34643c8c2cdf89beb428fae20cabda4e39a38e6054d945
z3cb3731c5b5128c63fb45f736bfa5c7a7eb9b19f6d3ab043ea59f9f322ea72f1a010a7d2bf4057
z5b2820b84283bfd7539959971e5e4190e341ea5b57b908a89969f2fbb62c9694ad065954ae2921
z7bd1c06bb06ea4beeb05e742c71023a9e1fdbc1bc82adc232f207b124561ffaaa90ef75cec63fe
z267daac11a30a9f32cf743376846d089a60f3eccaf4909335d24a07be8142eef40fe09df449dc2
ze9b970f43ad4e55a52267ad3a904f29e6aa6c4bd7167120fd1a2b33ceb39f20a61d52dc32feb6b
z2015d3fd48d55452bbf41063003bcf45efdd284529787981487c65b15371b03d046511b0696b88
z42feffbc93d43536a1d52aea0bc3be1bf0851ba0a2c3e28d61754323098838e25c65bebe23d466
z15d05204f861989df8f9746156cf2d29cd01dc270bdbdf20d6b9c2c032ba904c95f7f3e6571740
zad783699aedf1f879259726fec18cd9b7ee1495d6fb46f7a4bdd8db4468e65dd5df5f1a77fb9e4
z700d8f1d3cf9636fdbcef9511f7591b3f01ddcc6517e68f6069e04d1ea966773be5e1b11672388
ze9b58a91bf6fa7d19235c2660bc71cd67bc23a11a04812ce9bc1ef51bf227828d772ee40a5b8db
zbaacaa736ee908490bb01b90099ce98aed24e5691b89813c70cd12753dea526faaf2f0c313a2c5
zd8a42cfca7202c747145d2e1761f882381c98f8257bce93f351739fede630c32792f508670eef1
z533c525793b7d33e15f6ae26563daf0bb3bcbbbc983119178df0ecf8c3214503f05bf99d168d69
z41f573e3b41fcb29c3ca5497803fcf9c73ba6ba8c858a582cf6847d6e5a3393a053af8c0811fb5
z0756cc9ba96c73a47af9bc55faeb37af85ade706805e6270d649f1156d731ee7f129e1e1c817df
zc97dfa09172cfca8aeb626388ff8f4bb783af3ca0499bbdabc263731dee563fea95e1031639bf6
z81f8d3379e5e586c8f4b1927b82777284bf7dfa039db126e75624ec2ad0b8463ec81a871340e78
zbb2e24278ce659a558e0ff2c57b0d5392e3cecad5470c6d013f39845eabd60248d2702a190cb9c
z0db9656cec05ad5b9044b17ef2cf25d0a6f7c23281cccd04dc975d7acef0c06545843b05852788
zd92cb09c46fdd66548ffe75c25862d10ce5850ad33a4ed8b6c8e173ce63a5d48569d18e837c13a
z835b7b95a07858428722db5ceae2ee02af0ee8111c24e882613d1f1321bdd663e49b2de18264cd
z9b4466932bd68b988a02a9ce0f83beffc09e670cc05158e7a992e2aaec3728b70c0c96e21e5841
z92df00c271f38e1c050b69ba3e2d16d9244802f7202405a94c11b2ea7a24dd5cb9b160778415f6
z469cbdf84d074d4db7fad4b6f8c6a7a7f101a2f91cef1290fff9427c8f6322cd3fba5a8dcf89cb
z4ac2f94ccccb519a6e7e31c3967012285d17d937ea2f8b897e7237016776bcdd94b0d868ea6b25
z8054773f752c4b52d2ecc1ec0049e08b8be25b0475370cd784ff88b83f7378a240b4eae83f12e9
z41f8260d4db65f96390312e20e740f20f12a5e0ca5a92a46de76e76135bbcb857d81296eb3d690
z49f480b44098bcba1de5094c153c568df580c792ec46e39d162eb6494e7b857c43600d3d971fc2
z100cc9778c354d5acb5e68ed60def6be694e608d8010f31adf2492fba52da316d8e0c945a5c9f8
z63dbae672ad1ef1df447046e26b88287cc23663fcf49eef4f5a824e45297b891301123ac2d5acd
z833b8f9575251d82be620eee801c89e2cd9bea3d43a643137e5e88dcb6aa56898242add47e0350
z3765eaf7f20b848f11ec7c57596e3da93dce1ca8ef155f69e7a1ce78ad9ba99ed22bc43cedb846
zc6740359d12dc9ccae0e1936a0f3538e3aa002b3e66b213f54f1175f8c66486cf4a55420cbfca4
z611a0f99307b2ed6bdcec3ac5f7adaf850c461e9b8ad94e16c58124518b07e499f4d3dc15d096f
z34ef1720c2d9fa3f8eefe886dec614dd70fe4a9baedaac5cff5d1c81582e1777e654d2b384b6c0
z776be825ab71379136a65e0105866f9c09d88fe5c1e2bdba3b8897064f594cee20b2ee5af69ba2
z49ffde956649f0f59ce0ee935d21e5fb2a1f2154c2b8c5c963d423482344216f3e8a2112078f8d
z7d0c58c2c47f292890ad2ce1872230871b40b0866545b13ea373f8a0956f7c05d5aadfd5fa8306
z05ba0c46f7ebdc9496f732734e690820dede3b9c8196d936f08cd6dc8238b6f113db1a8ce6faaa
z8e1a20369986a611fe8be184f8f7a2899a19d1e3403075ba49a7b69e4166420990f946dad0a075
z66486e2e3ef3171184c10fbad7dd1bd4f26ee705984f0c529e26b02bb4680ed2fa9a59db432441
z9c5ce4b4e5f06099dbc2a4c939ab7915ada5708c33ec9da2d904ef343dfae6125fb737246b20f1
zcef0be6bb789311df97fdc766b0dc840f7e0c4fef9bb41736a601b8d7eb6f69e1b5e6805ddedca
z1f3f6965001c9fe6815f60455b182619588baf478763916d8999cedf3917ac9306f59e21b446e9
zd039c6777597569bcc4512536f6b165d5c26d86a17ce1e571b84885266d123a6b3444f6648730e
z20a10afa770d50a48a37c53697e9884b1dd42570fe7290a8e07caeee2d93be05b2cd118bcf7e17
z63f28eb91221c7911829ed1416f798a6e6bd7924631eea8870022b5a3126cb06f365803a95db57
z396abfc2af62c091016042aaad9d34c3527a34086f9247ca6f9e786db4163127452b2799eb6c31
z46ea1db913d2664779380031ab33e4b99ad4c66b70ba367d7b054db0e30ff68fde35f154f2a975
z3cf701385688f424acc95c79ea67d0f2f4b2c26a17c1d5f4c52b70ab3416993552042eb895ec97
z47f2ba9d9a72cf23f63bf06f6e7e9fc903b36f2a86243daa9b9a95362d9999270794ce165df6df
zee8880ebeb94c1fd4f642c6c2bad7427823dfb97fe5ba69cb76cd30f7817229a0bbbed63d3bf12
z7b12e92fe1a86107464cca8ddc40c2496d910b01726cf2b023e18fa3fc3ecbc5ec461c48bc9969
z905adad514375e170ed6baf68b443211638b92914acf975a0085244bc3d6319f51fedf9fe29362
z6980670433dcba1086af5e80509add9121425e311ceb9f6fbe4177d9852334637140a2f40124d9
z7c5c96e414f59f00c09f1be74b833cb8f368a5cc85b14c872e4592763b7dd311edafdf9e1a7a7f
zacae7c2b0fd8b43642072044f69a36e73a3349f118d8b38fdb820388c9302ab208adc99633331e
z7ee61a3143e7ffec0d8fa9567b75e4a0526df6b42b7af532fa1ab3aedbf8c331f55310d7878c32
za4f1d4f3ca6065c164813a2b898fa2b47d375a5069e59f152fb2e8efbcf4c16f701c53c05a9507
z7265d90e80651bb02e198837c896105c0a5f7d4d48dce0e620174626fca67f75efcebcaf66ede0
z6bff824584e3186e29ace6d0431708e295f086896a539140d8b1766aaf5bc04e9f778c407e24c3
z4db57c41b3fcb7570f9d59809cfb6efe0ecf5efe29f162705c26e48b8e171869a1f1b61a2b593c
z93d6b9cb2e611cc67afe3434c2e7129c8452b26b1f942166f6273bee83c12dbcdc6e416649891f
zeef4c74c2a58635cbff83c41a47323f6236d6a8226423d4e3fa78252944ca43f0f4151193602b7
z9089938ab8d6f220b57aaa4392244210ae6b4aecf8de6ca3522101772dfdadef30443f71afce79
zb24261505cdc28fa6f7739614cb6bb5d697b53921c1645af36711c1f703c7f37b521286500d4c9
z2ca4273e538aeb87166f31758b8af63c7b453766c31dea55fa193be77ad785fbbf9d777b3337e2
z56e6e31be88b9d27ded317f1daa8234e543943375fd94294867b1180521227dcddc045a122deea
z8e5ae061790c3ac6ad48430e023452916f5f4d90cfe86ea2f6b208eb45fe0462ec95c8de16dc2a
z402e187657bd66abc7f3c26db1efc2bfa4420fa6ae56b107aeceeb27d54f98dd5dc8ab6ca49cc2
zc23488b85314295159fd67d12188361301629c6cdabbce82832a7d2521ae187e7676b8dc0e2f47
z16be9fb3b6e66631f059d728729793881e0b6a52e46a9b4df2a6f2d89cdbb9cdb74540c47be4ea
z06fed2c89290cbbb7c17ff2647fa002b431762f3ba887217fa33c981d76e8ac51453892cfdb2f4
zed911186c7ace79e1d4373020f2f83fdd64dfd4db37d27bce95cbed739ade3acc46fde58b00944
ze1ee3e1f081065d18359a1a4e80d343ba495a0b7d918e5f474923f70d554c703e53859ae2d0ba8
zf7493b93875da9961210bf075bfa0ce080720e9cf22d69ed976e6996705e5e3180c57a3864c87e
z8f2f7c4ee13ca1c47ef82cb7ceae20501bb709665f7060b487da875ab29bfc41b5c1c1d7010699
zf26ce1d1276e76df85b5523d61501f5897b886dbd2ba8cfce07c3658dbdb7c76af6a4d5d7a4d29
z63f84be27d9cd016144b6a9b01b1c047d1037d2db3f66843dc6855d13ed8805c07d03b70679821
z75d0a97a431d3b33dcac98e2bd2f87f4e8d9c0a807bce5fee32d384f22e6e4b45e7057043d5f92
z79d4743d318639fff266273ceb1bf472147bc40e54bf0fe776ae3402502fb444f0014fc8439eda
z0c090ae5bd6d87e56adc3939be7880e62afa849a8b99b750692a1f1b69d69064e01948668517ee
z1d9eed2ff68abd6e9ba5e2bceac792ba51e9eb668cc895aa93b52ab981a5690412ca65f71dafd4
z17a1a833b697465d4d2d2f6f761d6e92e10bb39240cc68f00d057f72dcf8ee02a991b421dcf613
za81f1b0a882e169b566539101c95628750ddd33fdf243b27640bb1c0512e96b1f6d39abbdb5e8c
zcafb75d38737d772a33ae34378d1602bcf3586cb50bcd37cad475917f3a3b27fcf8e2257b6c435
z4848acdabcc49e4cc074f1fea408e602fb7f997f4fb7a9816a12d761cc5b5b23cc0073edead46a
ze8da4525a6aeefd5f69272200179367c753a2eeba29b22a55840e219c82ee0e70f29985a57379d
zfbc56478d11482c472e4acfc73cf3d399886c80212e2dcf49adca8315b8f4fe6541bcc02b4090c
zbe28e74bf5ffda626a408ce6f7ed863f3d8ce01bfa71b9b0aaa4d7cca437a1f89020987ff08211
zdba49b27d4e11621ae97494c742ad3ba8a5403827f551806eb7baa5e0d95bbde9d4965e22e27ad
za17ab3f8d91b52dd588191b974f3c0664ce9f7f8555f7e958e3b75b958a8ce77a4f74dba4b7513
z884c0bcce143011785601b2e406eddc63246733dd592f2108ebe9d99b3f35282a0a5810fd1691c
zf5f20060fba98ba36e108ecf4d67bdc17f5d8316190a1020d9b83be1d289d2a41d280f0c532416
z59655b346d88fc14c369ebe891b2e00046f2563fe7f79d03461f4cbfd7e7305382176c7f775c2a
zd4bd990e2496dd11f9a5ad44f7d590edbd82506b0dd431c8e4bccb3b323e9abbdf9487629b4d77
z9b3d042ae0187c59331dc6e58a392a178621cd9c2196be2ba7192f99b349d5f2de464d77677ac3
z84463a859980cf1d29a7eb8a27f9b9e5416d2d2044bde96c2bf0a468f500a0dc076746451c31db
z71ec1681ccba4aaf21b35c9db1c5f3152ec89312552715cf7c3cc2ccfda075541a89d53a95f4a4
zb6da8028e8b499701716d34ad0d65d41ee5de7b0d065b16e5cee546f2dccd0cf1a278538375972
ze74e5414192ee0828b43b1e11dac273fc57bb2e81fd72db44c10110710f1ad12528823fa636e13
zef14d57c9c5cbe8bb423f6e4a51ecc091669cf369fa14a61656598e97c024580af075b0f03ea8a
z6eca0b591eeaa3dc191aeb3877950219f180768159af3f2efcdb47e452bf12b590d435275d72fa
z8aba4fe56ec3541e6ecd137dbbd260c301803098637b93bb0fa20ed97b5db81ac697329b8d69c5
ze1c8d3349866d8bf1d77fe30440690d19749fb4397af69399be27ca4d1b4897bbcce52a7ed3ece
z751585b8c2bf5a5d1ba32f5ab4553c06fa88321f5f9aa2e6685d01bcbe573e49e51236eeb2a768
zae21d318f7b22b787273e40e3ce129c3c6f4e55977eb52c3e9608a5b57315e86d96c3337695309
zad225c7c41e1b3d2d9589cfbf1c63481a8dbcb4e82f7612866fa6b33d73e87696db2e4cb20f906
za93436c6ec94d5856cceeb8991ddf01d2c004a77221cfb6523a200a2795c34adb01f12440b4fc8
za3741684f264ea6a0e862f97683f7066ec482500f574aceb8c5622c6e82c4176be0126c5641fcf
zcf95202a10bcdad4c4f29832eedf159155d2c037a76e02d1f6f3d84cfa923a519f7f76f5ccae80
z6f889074765f91dd6f4a389d90b08c4d02c7d1388db071b1e88c7163a2eab2228c2c0416606d07
z4202f59ce0d69c095fa5a9cd3c3d89d8ff69190a6a5d60fb95694d15f158b8e21f6f86a7de9fe9
z9e2e691d48d70cc9cf6067d26e1fc15bbdaac868e9f890746d54e620092b36668d50231a917a1b
ze91b160eea41830a5aca040b5ec1d01f73a952e1825af99434289ccb7c410190cb589120e3d475
zca422c04246f6a0aa7fdbd2750860f91c99324a383caf7350c8102fba2c47ff93632fa2252230a
z6e02cc56a3ab86ab1a959374b792bba45d98f05a131338bb50c6540d087d4c027d0a3a6d6821c7
z7bd5e2adc36432582019945052537ea79f521a549a8e8bd38dbd0a9f0520dd4a7c5a3d71091f77
za4cf9bb71b063eb78db8b3de2f3b34875ef4265ca6677670ef5fa2de72ba0eff014edac2773518
zff3cd85bc86fd55b24c154eb0353e496975fcbf1b76608a4ddef19410a3b00f08934cf6273dd4e
za14cb4af3b10e7108b182c1baf85f22ee89abfb8441732069a857bbeadec504bb13b2115295448
zd86d6ed5666ef477b1f9afbd4f420f4c71f49e5c5bc8e74a0cb74cbe0f46f302687a9ac871d7e9
z7ac291900bc910760dafbff46c1a972cd6313192c4971a4026a8cf39bd489a08df81dc21c40d3f
z8b7fcc2d314cc7d19ab5b34f0e907a12be1a1ef7679dcd49ba7f4f977543b321e793647bc17332
zeac10f8ecfa4d5a2fcf13181e415ae7417788ccdb5d36bc83cc97229ab2824ca8ef139b87d1a3b
z719a0d0cafee28d89b336a9547166237cfea0099fc1b287cbb59a4708871973c878770592b4d79
z24993ff713fc86eef1d6f48fd8e5c3be5a9b7aa84ca12f2813f00a8cfa0a2173ac8bf5e4072de1
za1ed91930f8fc4866efe5db6f6586ee7fc6728292de2b4c5ee5a77d8a1d5a9979ccf4ca542b4f7
za618b286e75f1ab48bcaa817b82686550ba505587c679d64193030da276d1690b337e79a098364
z94c184d03b8209ca9da7ddeb3bfe3dcceaf6fd79753de07e6b60c01200fcc139a24b9f9f9af44b
z3b9c26245a3a6de1bcf309d1f0afaa952623fc4d3955d8ae40d909f995b24ef11b8ae6c6105d5e
zfdb91b659707ce164456e34f797b855525b06f77cb3646282c7e8676539fd8b49f6108c205f443
z7382bb44e2cfeb48e6dd5717370d904a62647f571fb51db50da5698f324c425326fd5e802d5a5d
z1cba4721620397c695b68631c2b113d8d21e4355fddf3561879ea9384b59d50791ed45d77b44d2
z9ffb56f76e3e90bccf2465a84fddf14235e2530d76818ab2b8b1c5cd3c68fa154c8e327fe58fa3
zd49eca16453d870a8d9f31dd5a8e4e77f6431edc19567175e5008cd8f6beb7d334ad3c8e9d5d73
zbe7ca1ae6f843bd335d00a48e431373e0234695be0ecc5c76bff6848ce190dc4c739c382a6ce8e
zae039eb2d2f61b9f92a2019b863c3f4cc4aa0e7e4c2e76722b9a6b2941b64456feb2feeaa67395
z8f18682d08fb378fabb9b2c8889e2f42af0f8602ae78725a7008be05fd48ff9397793009dd87fa
z78d130d92075ee916578dab1155ff443530cc420f028e4b63d0bb12657227e24e3862509319301
zaa1880b92c53eb4bf56fd1bdeaa841f4b7c0963718d9425fbf1e714f40ace9aa2e20a12e7e0dc8
z66e97eb380719a8663ba546eb1f2a478903d25305331f7667f11c1b4327a9748ef0926554b1456
z1f072b5d78543f0d359ee7fa5e1240efc15cef25e5ab59aa9acd1fcd3055c4e4e4922f0a8824a0
zcee2c61b84a9fa33bfb828f273716e023fb73ae2cf4ed179487f7110cd08cf2a950ae382071381
zc71cbb703ac1733adc222916459dcf2437dfffaea04ab62017e34d192fa33844126f16e47734a5
z8e9092f9df51a667af8ffba4d0a284a484ecf047eb91445577204645f5b340b79fbea5f2903ede
zac126128b6f376cd9ca02e305471482c1165bd40861d0d2e81b712f0caa9bf7a90b4b08e5f7031
z258e6763ccaeb9b1c9ccb6fe747cfe1d9d58a1360dcfa3450adcf2d23bfc7622eb3737f4317ae9
zd73bb3d23cabf7473125e387a56149fa479dc1fab310461aa8b0da75daee382af07988f6267007
z2985cd2fc8c9d91e90c098eafc02abb235aec142e1c13bca4be3436d130e5148d972a386879791
z9fcf80799d1385741421bea2de2b19a4bb5899417af1e57f691e051be75534cd2c775b1d318aa4
zc6c4bbbefcf2841f08f67f72834b7ab7dda89bf309803d8fbdb708bd35bfe1bd679efff7411cd4
z5d0f63617f91cb378e8953330d72bd365f1a79edeeb6f70b62427bbd3622195b4f6cb23ff60b71
zcdfa99e3ad85f1811b5efb74ff649820b94e27e96fc6d68b3bea49bd8c12cf2197bc6b46a30271
z31edbabc3d150d329a47150a5641fd633cd577ea9f7fd2f5652f61dfe6848879962ca6c99d4543
zacd391c93061323869863852bd544fd3378089601649ca21e6e1fdc7154f61fc7efcc03a6e7b88
z7aa963070aadb4e1201d7394972c5e2eaa6b93a75d03cccdabb686af348c51dfece27264d7baad
zf9845e56aa633c3369537b32d8a744a907aa9ed51097de9c4bd35b95443d8a7cafbfdfdea019e5
zfbb0ffb6ae53aa283f1c45e1f9b13148d9132189543a8daec428d56efe5c747df6a27d1de80e71
z4867669b944cadfd0b5d455ea70fce621ec14a1287262e6bb24db0c02eadf3be90ee29c76b6f1b
z3e0e5c4a7a532358ec9dde54d8c7fffc894065754d0b3354e2b1c7c7268ea72136c248c751e029
z8234f998ef236ade40bfb32d2a2e292c98749c6c6af3da625e582fa66b9afb9323130911d4508e
zeebab6d9eda5c38837b566cfb29a0944ca3bc906ff9e10a66f3d669fbf1d5a4071e8660e6ae6b4
zde4dbb983dc4c1002029348acd2954183989c26d7f31f093ab581291cc7e590d268c0da8da04ab
z82d66ba511081eafce090c68d8616eb241eca85d518b76cb169f861ccd3c3459c271b094b47c64
z06c1185f0d6e1e71a849baa43b2583396796eb1b880daa9a29a58498aa0b34586badc6af1bc181
z21442a06649b528a50a2dd43337d23ded525935971b5c6ab21975ac47cbda3f29b4daaa47d7342
z209c97cde80228fc4928f4e0d61309d2df0b4e5b7de676bfcf33a5e58006ad2bb9519b09a1eacb
z427ba936c8747932f45362ae79b290eebac12c075f54f4fb6b0e85f114253fb21424b8188494f3
z81f85e89183dd9cb0dec083baf5b670dbf520fc4d669339c12d542fb25782892b9cce4364acaa8
zc1a555eba588be1820058f36b21140fd05d007e47e371c39ce107e8cdb2a64116028815ba072d2
zb88b777f5af28eda02bd392477a758578bef56e4c2285acfff35b071872b4e17731ea64f59d83c
z8e65cf00fdc5a94e8f5e40ec26acfa24b7b8b3ed033b4a47f75e48b20fc88b87a75927ec55da5d
zd8f660b787802bfa0eebe56fa005662544e0b102f72e611e477fa056028d8172145851fed21a90
zbdc4294bd4761c60b783d6aa12958bd754979b87bb8e75c74e1043f8d1642816a8684e62298382
za700c47159da916bf0454b80849136aba7e7acd6e312b23f7f29b1378c51a8a7181061d7443739
z6d50cc4aa190407343e6ce37ad18ed4266f223d2a3c6931eddcfd76858541edd5644e09fb00492
zd1a11e8bc5ca4fb2657607564ac25c0032c134b76b0fd5b55b4b0c3ce31c01fd4465a32c39dba7
zd8efa9fc3ae8be0ceea61fcaddbc1549eb8d7f2766c3f98f748926ee0792e6a690207dc82e8a2e
zb719f271dcb6b339afa4cf298898e1cf673176e2c2fd79d4876eee7e846985d0023710d4519858
z946163cc44e8dac3378d446806661f58a20e0d5d1ecfa576414acea2a149b9ced60fa29d2c8626
z4df4c65b32c28f555de05f3d30abcb5bc11d6a3fbfc0a0cda0327af8f55489421caea879b810b2
zc2ca6e2212b1c6bcf652e748fc9c7759cc0842b347e75a1e9c8472db66d75ec871cfdb61e6de4f
z12069896166d963f6ec9309978a77c03526d473a388eca7b54667e57590afa7787fe9d8c0a34e2
zac2f313920f0412a2b92a9ec7aa4a045960c5667c6dfadb7f8d16636c85db0b284b86c38c6adc8
z58a7c0accee92fbabb7b08c77c0a76702b8f16eea33bab45cd58402df5a1a380bf724dfbbb40b2
z2db2bc23c1f6134f3e3054573e1b51d93316051df7364ed185bfcaf769136829ec6bfd294e8940
z475f6bff44eb34753c3d4b8c48fc3e642cd2953538c56747482bcdecd08eb5bc02e5e5632b1ee1
z28fb454e41962a333f460e36646aaea8de23175190434bf8c458d70e2e001a3d69cdd90b0b6738
zf9bde4a55216ddb3ec30ed360d261a63ac98759602844f2589fc591c79641ca4fcde62a73e6380
z45f99ddca4a15978e2523fe7cc97705243a4326e0f9688f5393239618d8cae1ad92a88e2305c43
za190a0d4d2ea05be5a6370bbb97eb686b9470e2b497ec01278d431cab006358a3ba79e3ffd74fb
z36d48d1282560ca5a72b8efcdbd6c6f7e2427d1601eafcf9cf64ca44b02bf9ff1c3deb5417d06b
z5455c7f88168cf87ee29fdaa01431cfb320d6db97b005595ce02ce0c6ac870d2a1fa7ff83367d2
z4ad55370b6de895270498d4d563665b3bad70c877e42724667cb03cb5696c9d31535ccaf99d21f
za61f63c7ec1ac7713bcd664804fe6b330ea06b7dad729770acfcb5e5bce7653bc79281ee99e5e5
zca8de33cd5696ccbc1094e89367a5fcdb319c8ae2a6b7dfdeb9670136f2274d17af837555b4bbe
zb072a84eb45f8a482dfed742053942b79ef6846c4430b5119556d7d4b0f0a4647ec2172576412d
z088b25edb8baa54ce5bc26eb9d06d354c083a470b69aca66b2fa1c8a81198e512ecc5f205e9242
zaff55a01f13dcb7f15ca767e90b24807174dd6ab4ccc9748ea6863fcf2496d0fba440449f89ca9
zca595ab7e1fc4429ea76bac9df536cf3244e3f97407f0d3937dedc04073b0e66847c557dbe5095
zb9bbe997c918ea1c194ae561470dc94f35946458e77389d56e995f18c5fc9f0aeecfe33a62f811
z6992f9f1b99259fdb964743ef05d0ed4c25c471fa194efa900b2861a523c1b1fea38c52c0d6249
z1c016aa0ee1af380b4c333dec264bfb9cc5016a01ae533f61a90d0c78f40e27cf72ff55b81b465
zebc5e134c2668e0d1055f608a7bd717d030d8d4760678f013c55ba846c14f3894e63f272106927
zbba94bb1c6c1f2bdb42de8ef1987d262963192fbcc5767ed6a6eed1b4a6a946ebc92a9f65afef8
zd14a01e95569addb398178f703830c236dbc693449843cfd1e145bc178cf29ea1efdc084611567
zdbba3e34bdf0dc1b3f8b397ff0e7aeb2fb0a1f8ea5f99cae630f2e9d784fc5e677fc34e8606984
za9c2eac644940989cde07125341a8504161628c92ea914efa1a04127132ec4ec5a79b2c1f1d516
zc6d7b2f0a2b4050cead2d1167fb5853cd1e26790a4fcd145aaa7bfed6cf02e4267412e1b09ca50
za1d086263dae6d5bd5c44c749194fafdbdb5e05bf42bc8ffaafdb945bec63306ad4eb1914079e8
z630e2c6d5748d1b5d397c135cc8a9d344704444eee575d6bef01d7e547b50bd5a190774c8e8943
z58c5940c7034f13f86aa1908b85d87e9abe9634cdaa788ae2d161b15abae06d04b8e11cac1e38b
zcd8f55652ecb6fbc534021704fde1a301916ec05378e595ea50a369dd37fd13c56e7794520e842
zb8a63c1b4f4ab1fb5b9abbce6d75d32119adcb03cd5c625d45b5e569ee4d44d8420cb4f5d2f240
z5da07499627ef0427cb66d80c24abcd56dfba362fd79f3d53062c68bc64655e96be612a299d42f
ze274da926e4f246c56c286559fd10c2d89838942c2471cd6cc3bdcfd28dacbc10154494387e8d5
zca578f492b2f3f4ba793da7ce865fab901948d7098eb23a306abc7e11da1b3a9f066788adea88a
z6b1cd3be7d4fbde7be20318d2150ed8677b4ef592510ce809ac8ecd8dfc4e1edfdf2afa8f1d08c
z0a9db40833e2af402d425026b08ed7995e36c5c49107e30e689a469beff27c6a906353e4f43545
z36ddd64edb8de93986ce20d0744c04ab903c97413fc3db2e8ea12226605ed19c687b669af16275
z60dcfe51ee115bad4d4e270976255b10d08d77b8878d95b9131938ec1183b9c177bf34dfcac355
ze3883a97aeef626bac862f5177dbe46e31becc263568a2263ccc5a933db1568b216c16ab893608
z6cbe1131f8e567d81679b67f58bacf455dc14d4116db4b842b21276fbc3a99e5fd06e265c1db7f
z1bfd7f459fc940376e5c9b66ddadf6a9ae8e67c7017295c568c296702b34b9384eefb2208036da
z09a7cb9c303f5083d5ba2055781deb06cf35d1592ef0bd006571faa337c9ad2e35029406ccf0b7
z3728aad7dbb5b3850b45d377ec47d16296c5174e3a51ca4e5e8f4ffe255f2b7372d38f00dc25ea
z0299c36286692d4af2424dae26ca487bb6ad6956f2c1c4ee43acb962ae9fb78d363df829c35d3e
z0d3d2081794d5defdf1ed4ca9a0798e26b824bd01ffe7bad6e1fd731df636bd58946c5602ec70c
z9813a651b169d0995571cd38ac48bdc534532d4be7a051109252256aec353b702b8aa287cd5072
z008cff05ff33817fc0540fbe88c8f54f57ba724556ff07077d0defe4d4d3e8a4678dc0cedfd262
z9cfbe967404da12f3ff4dfb1ffc5af72524cbb61b17c2a30bb472dbcd79e5e66dc2d436160495c
zb327a1cce6b87dc9a5521957a7d0d4d8dc2baa4cbbe3a38167aed96f3583329c53d99c83a322bf
z2d4b7ce2f723fb3efc76f1429f1dd3d9c3cb43e1da5e66a198b7d68f4ae0a9be637d0b943197eb
z0c5c178c78f32c31ee6824b7c5ca03281989ead6312631bb785f6db7a974a1bb05b55d1ff2149d
zfb21f5b9200302a0f7f82aa0cb432ec4fdb4a163ab24a71f6452b1fc83a33d7512c6984e112753
z36038d7d602aac897010362cf87e5790ee25e939db30d95d88d6984d11fa862bd9b0073aa2b8fb
z4668952d2217daff4b9bb6867180a2964f490054feb2dadf283be36b4e25bfb2e43abddd965ade
z0eb4143c00cc577ad082356eabce6da4b8ea4cb562c43328b6fde53ee19e5c187036f3cfd7eeee
za4079082f3c84d5ec971e109687deb62d33d12ce2ff9f43e064bfc61886992aeef12355d21b086
zf327dcbcfebb6412a06e00a2043e2fe2758da7f84b4bad876eddb162cba093109f91eff3f08100
zb294fdb358401e47bd200f6a6b4e4298023b11bbdc5078fea7bc51488a5d909219050f4dba3009
zfb342e480ba6dfd88f6c518b678e276ca112787f5f0236f450a85166d168d0b426c33f64460791
zb4adf7e8b0b035aa48abce173ef54b3c922ccec63f00ac8bf02bea83a134f807ba9217ea0ddc38
z1b19975e2f03deda8ad5c7df9999a501d32d27774ce218f38081609feb745141125b98283b6aca
z66912044952d8abeb3397afd22abbedb1bea8be96f513f4738815319514ded180cee61d160c7e0
zca67cbed35f762eb909a347da53f8c16e17ad2a48722ca6778313f70c7a8e4c9848cf6821e53b3
z83a81cbf58968c6e20a4fb69c630149f9216dd09ee526d40a720730ed97f4d8f763772e1dfc7b0
z72abb5f757baf31ad03f49f7e09f0417c86e0c34d848f07b61a9a045ee9d625b2b4db15bfefba3
z58c8e94349c9c3b201047a0cde68c87ceb661946d946607d11c721f56797e119f4b0ecd2f25e74
z7a93db781985cf1631218066a0c2ec41a45df1b58b91d85915a72ea23d1db69cf8699f4641af08
z5ef401e8a7be83805d70011350d764a1094b806d74e2494570c1ebbe9498a807ccd667d2b278dd
zcfca28e890b5ac5ee89d647eaeedda323198a55c7244cdcbd0404a21fc73e0a3c707fa24a67bd4
z4dd11b53adee1f7924acc90cd23256a13f9083e50ddb86d994002777e3896a9fe10ae89260267f
z5e64c859b30d05a209ddaa5f51d27094b3c478d0226c48105ba8d3144be6c9f6f9dba9da75b1c4
zd697f489925be17fce63632a5a00b4ab3343e2ffdad55f8099c81c9f0b2867885bad459d823b5a
z78ef24786c5df490a1b179a36b04837bb49f58e166d3b07de2bc52f38b364a15d8878b2b3c12e8
z080cea6837fb48ceb5daeef3dcf2e921eedf5381af75f971b2390266a4c8bf0a0b966b6465d408
z5c377955770af368274ff70d76dd356caaf7c884289dbc9681083504201e9215bf7eba590c1e9a
ze910b51fb4df6438c740955ae10665354e303b51d8f9360a39e86704a3b7a39c0215eb24946646
z93dd46f426689b80867911a3b99d02cf60254b7faf5d34d649190878f6cee6aeb7634ad9254907
zb11ae40f8a1eef0b1edad81257a504dd4b917627cd96a2c20cc583054568fe8841902663756042
z9e4b5d7291374640642933728809bed81659e90165e713c0b4380eb1d2b79a88735d91489e02bc
za818cbafa84e9d4223d4748065417da4f64c6632ab6dec8682d25f9d61884fa41d5a8fa3c9328d
z02d5ef6ae524e6c81f8e5318e3d3484a02a7de34763a7570941b766f8e3ae14440d48668efaf88
zb5464045c3b2a94ac533c527072818dbde9fe7ef28ec96fd958c2a53676a2433d4a016ea11a69a
z390f71fa05910f84b2c4ab143096d25a9540331b3627c33ff9650f4d921058aa562b0c66682d79
zfa8915e2307dff18afdfb15cfeda820690d9e7fd557894bb7a7b518520d13300ab234611980472
za06ddb9dbb004cb276445065fd7c1596c06b27f73708abb17294b74c959e6dc453981da4b6dbba
z5137003893b42c104fffbb23b14515a01e7a9846ddcea8602de7e63b8e625ad5dfbb01ecf17a0d
zdd1eddc48718091ebeb06f01900e4a37b5578cf6cea8fa2165bfa839fca028b410915297f943a2
zffbaf883e16487709b6e97dff35e5f05b4e5a2435a09634ab4c4b3b2a103f38080fdc21e4912c3
z42effc7c0a800cc80775b92606b48c304aa87a0604ba1a77eaba8c141b6b6b6b4dda8b9bedc73f
z3465cdaa2194f62f417ed3f8f569c7a5401a480a30ff6a095cd16d818ad82deed2963ca9bac2a4
zd8ea73b5b00baff1b30d96cf0dd694453684093798d5f738ecfd664ea49e0cdc9227d24ee1c1be
zea611c92c0e83352853cfb399584582e3aa2d9a777bf183d7015585c56510fa296224cc7887ade
z4a4481afa7ffe01fbf0b69d53812c073d241d8aab1b889cc36903212282a2803b68e9d442d065a
zb0e99a79f5a14185d00f2793749c2c3c78cdce0eb5b0ea8f05cd458b379bf7ef0673c7aaf3a11d
z8fdc807a5b81b85b7ae4d44135b2bea18c933cf7a27660d5d3a3b8584edb06224c2814a34a544c
zb9993708feb922a9cf67661933c4b86f31a039f4c57a381401bfd4d47821c39aef8b538e25d20b
z4377ec214292ce6cc26cfd0c0c87ed80283ce70457b787a6a2505b3ac9f20fa718f7ddce3fe463
zf963acb2d96905b33c06a1c17287606eaccdf5d12a33bed5b19298894f671e45e3ca88d77cc5f9
zaf79bbf5b0b08adaf991621aa3792e4a1612e98eed3f93b8945ebc9e9d8810af17cc2071b5b98c
z9bb690ce60f255ebf80a9944b1ef73d3db1e74d0b7683e17d37ab4670ff49290298d2b81ea5257
zfaa9292cfb125ca15c4fd77ad046c9364de44510526f7ec204f9a3812fca3c7694f38272894d41
zac8ec2d81cc2438f71afb2ef94bce3f12b58d673d991a18acd1ba5fdf20a454adbe9778189bc94
zbfcf5afef77e364488c2c170c8867d919c29bd68c5affb59270ebf59e17599d94cb572edd19acb
zf9b5cdad655b92a4cf16ef2628353866fd5798e207d89806aa8a3b378c46408be4cd8f7ff41d07
z08e9d891f3411a58549a00dd6d9d8ba927a0fee488431ca9ff11e9a17533b4b8e558ae6c0be4a4
z815136d23953af8e1859f215c7ac3035b548f743b3b6f6169bb598c2fb659d347568cfe7fde4f0
z417a12e8c21e22f0cf5ab3b8fe8084ec2c204a4520586ced4354bafb1eae6d8fda714697fdf49a
zd788b1d5836af645a6c59ae1a8a4e1d1efd6975657eabfbf236cc322a4fcd06f5704cdcf967033
z5d9d395ad41bd1b4b2022759de7d5504d7c4fbbeb2f578cdf7187b9ec277ae66f2e4ce995de662
zd0834843e5d6250c1dba4b2fa95160f18b7e63c31e9b4fd931ec63859790322af1707135b4f594
z466d849e820d341575ef131d84a21e260846bc419171e41848868f13f073434618ae62f74d0301
zd9b6a500750aefea4451d7fa9432da47892ed1fffe593dc3f4e6f79876bbc29944bb7bbc814b6d
ze5eb5f7a5a15bcbb25edefb848601f96ea18f110f470018d99ff499db88f354b573a393711eb93
z54b04dd8c4980b9236c716ef7530c381ec58baf6c42abb4442198cd14ee39e93c1c64b904da86f
ze9e20a7f7e2d0cbc258cb1dcc5b0c18fab69fef869b8d38266d5236b8158f0557567d3e35d76c0
z49efd4fab04a7baf8209d90570c27b774a08e54c583b737cf00539f0169e9a18c15b8c46bcde26
z502846c588d0c70adb3ae2cf776ee7748d6cd527fff831af0da517b74ab0b3af72e032a68c512a
z0e5124b3d295a2a3f14fd12a3520cbeceb93262281765d01a21f79f17a164a2d8633f10b0c48da
z1319b28558f76e1ebd92b7bdf54b202211495b25ff064745148745da32b55deb7b726510ca2e5c
z94bb4a9cc14b91796a07312a5fe6d2eeded45be67c9a0647ca6579632d08a35d82ae37efba91a4
z688b9d160b506c2c6c30ba78aa6b3b05201199586c7adc0d0ebb833b5013259096d4539b798ca3
z734977353ffb500bae19a21d42b222e7601b1936b4d3c798cc0a464d0ff2b7e6ecca29a283b6a6
z9e9131cc4eb2aef9968a250477bcd499932a97c631ebaa6222ac1bcdca9325a8c8ac5bce7f0b8b
z9f9eff82278d60735f4781d3176908cb744f93f2f00ec604f4a6282db2f6d8c665dd947c1dbf70
zae124a1f2e69e61e2b8b28c525fe557400285a7d31ede8a0243ca7cb58ac740594c21a49c0ac00
z266a865016fa2e0d7117cf65a38ffa25d2a941bf5726cdf04695b8e9cdf9a28b4a5715e09be7ae
z4ae7571b2c593969d8bca6e3447c7706ad4c6ed64498041b4dd6c539ad7cd8bcc48b98bb527327
z909921fecb8f6dd5d167a6ca62474a7599d10ce34ff61db9ed4579c3f96327b5eff75018310a9c
z38d57a58a1c0ed2d13047c31e198fbff85621de9aef34b6ac7083c70cfba62b7c47f26a7c1a54b
z2c8efa7fd6fc026c7a6c6ea43b0d8f79fb87e858f9ce438fba8e392603ee24c150e2d43a3db4f5
z4428d369d712f61248cace0840bc8a555dac35783653f9aa7435554e13d9857cab77dd668933fd
z278858f5f7bfa76707fe1d68b8c67576318e2dacdecac38028975e6b82d83da10a40e0552b4889
zab737444f0bed393fbd4a8c86506654d06ceca30f4ec9dbb39b4d943c0e3270180594e48233c33
z02884ecbc2740002b5167b49da65f783ae5667355d7da0b8ccb7cd65031241edd73c18e2124521
z4232201cc15b3f86001d292b57771bd7a600306a61c6b8321583a8875c3debb4c37e1abc17db99
z98395d3a131612678085070564e47ab52e14949fee75a5f1d2fb1ed59c810674b56836b0257ecb
z1792a0b0c9d05a13372df70d0ea0846b2ebed91cda318264129e1193c1454886dc76ae6b630c9b
z0a5b683a576c90e5808aaf4cf98c6f0c395a29ae44fafafe6560659ebf8e270ec6eb93e357c25e
z04343956b639930281bdff6269c8ba09a497eec525ffd7574f422f420946fcf7982721d0959140
za6b40682a678e3778e37cf44e06edfe1a143ad5f01ce22f7fc8ed5986275163a18be33c4844347
zf3c262523c414f273ac474c83d208ebc1b108465816742860f6246933a9c227f61a81e9fa406ef
z5ac6ca677b42084a4f177c86f1cf18ec1b3aa85009904ab87f3ecfb3a1f0e3ae6ae367127c25be
z29801f517e400deb13f78c3bededc5be52df5ac426103a6ec4d17d6566dea3afb54335f902de60
z8c877fb32e2375aff31a155e188cf1bce4a36c58db2646176923ed8eacd8ce577a087acaeddeb9
z449fe8513793e6b797f32cbc962c63c448235bc3cf5e5bccce203b3cca5c094ec9f147d7553af3
z549414a5496f03eddda4677bdd5f27442bf08d1fe233fae4b4ba67f827d7b2a52163f690a4a386
z1a94f98470ec8da8477d34af418e8283b00f113970eb420497d0bec602dd0e74e744a9e1dc2263
z6159c433bacb470636619b78aea0c961b27ae20022faad3a1f22304a8b4f9c95c7e1c4e2095b85
z9bdf500923303b5e3c218d66c40d4e3960de8cea5f6cd2eec604d433dcf91b3d165f3dac930d1a
zfdd54ec79ba0fb9f99df813e6ba72949d121888cbdca0dcaba927edb099a356f03dae8bd8d9b28
zea60eca2ca9284b0c03cac8e09711853798edcdeab8faa63b8fe5440deba57a12832b25e0880d8
z1279835234b76c61ef31d910ab14e114917720f78feff2e32b6ff53279f5b7ef34010806c075b7
z7a8382d053d6437930ff306b7bba133a52cf93240e6cfc1734faaa8fd097e01bfee9b7462014b0
z0cb303ee597dc5cbbb2359ddcc03edb5a65e488120bd49042d251b552e00d8d68688af8671b989
z99fa67468bd74f985416889e40f792703837b3656b41c852bfa0a87c5ff1bd1691ca57c33fcfc7
ze3d9870c292ddbff7c900046b3ebeb6a9a456b84cb035a2c5318db511f28bee49323655631077f
z3643aeda95009d6784d5fd6cfe2d3c494b860ee26e5eeb308ce22b45092d55cd2d548da8bd0bc7
z15817a449ee977adf7db54cb11fdc64b3dad4fc420586c6a295fca06e0399f1128ba77dfbaa9ea
z71e17b194c090f8b72683cf5f90ee3df8a28520044ace49c391ca4b312a26e31e22a69917f96a5
zcd1632a65e58023f461bb474f1273657edeb3e00bf979411c8ec6544303c1f0dcb4bea587777bb
z375cf67f7e92f39fad97e9258440e1b4fa54f38169ed3c1278da54ec667a82a48521af3c10b9ca
z32bb890265b50b7b1843168087caffa0667fdadeacc33f53e2aaeaca5beba940887228f0a0eed1
z5fadfdbdb84f81f4a63f7ea8cc97060ccc5e0c0635c736975c12b328ed5432829cd9556cdd772e
zc05481ca3862370c156a6605c855329ea000ca9e9ea2dd2b7da840d36f3c2538971340a97daa22
zb79724f440269e7739d396f1ea2f310813847387fbd6b58017402021fdf0ef1e6cd407f51b4722
zfef1214ae557ec4a5f391b563a4b48d4ff185c2ea18c9dd7e25393ec510199116e6cd763697fa7
z16f4475010cdb3324d1ebd5240ce181e8d3d6bdf3635a9247ba93bd1abaaa6a6661229734235a7
zca9ad0060708ab1484b531b99cc8ae6c768ee51a7ab6f77c1a39544994f1c4955378e8291a5848
zfc6f07efeaf5c9f1db279a815fb942208173e7126664a2faf934902a2c74ffe9f48f63a15cc193
zde13b8c35186d178099787d31b0a1a061b76e2ba5c6247cc0dcb39ef58930d130c96e4ab6c820c
ze651798079025b5ba69e0e78a77af854e5300ae0faf2dfcc3c957f771f28a53eae8698eb4aec8d
zf93b2600e307bc64d3b11066def9a4867812ae108e224193ccc0c0899369520c4dcd3856277dff
za161bf8484a464c180eb2c0ffd3f8adde70d856c2d572995f5426821ed95a5e7fb6a01158f119c
z18c026da45a282813fea7adb6a5fa49439e346b4915ccd5d93f084fe4e24a1dac4d63260c0276c
z4606c70e1ecd0c872476dab6f436e95a41010c198a42f3438680c7bca8bf4bcfaf39e1e14f8f83
ze5c75dcd45fa738a129f4ccc8f823f24937b01cbe6ee66a4bc7a84e881a2b6347906a6d3ef60d8
zbe81fc86590be4466329ab6154075af51db5fb5625c3da3545a0859f21cb9de2f5892f8eca2df7
z2a64460c2540868d22b5d78f43e9d3ecebf60f797ef1f2f8220fbc7a7d209be585085369d4a6cc
z136c5339b38281c9ae3118516f5a51c09bcd5781b7b07f9fdd966804ded4c0443fc6e1fa46dfaf
z3a04f6f7430373910bcaa61553389fce80c0466f78c9411dd675900cdcb4f521c35ab17a8a6e00
zcf310748f988bc6603006d6fde3d66744245fccd3184091ccf73186b6cbf9b4b940099089c5cb2
zfa856c70db448e540b31927138e5c957ee2928db9c5456758777c0d6c43656300aab9d11724ff7
zb7c2549b2c11b770139374fc8e7e8e5bb2809a43f11d728b88ce3fb9ad40050bb98b939bcd0786
z664e5fd4cb44ea89a071cd25ef18fab6510e8604554aa4023e4ad6d72c7451dc94cb61270326be
z52eefd098e5d05eb5a95a6e8066d9228e89e01bd8c83a9c6021c1f0e867f212d652451bbc64adb
za5ddb1a84145f4c8cdc57d90df3aef091a2819b439119667f9d67140f20dc581a8b1951c4865e0
z0a0ac88ec93884a7c770a96ed3eeb0a7ae2e1d6737c40f8632c4a25dd3c07433cba8c3bc954bdd
za588e7a02b2432bd9029ffa131bae403036c577532af5d9feecc892e9c62b92e977a8acefc5d2d
zab84582b0d309cbb4f367918266f4adce418616aaa6554e38dfe0d3d8be2282c48d6c1c3c9df21
z9c8cf6f43147fb93822b09034ccb185b33f11eb14969e503722659b7bd01e35244c866f1fc8f3b
zdbff929d4dddad5d685597e22f007c535932bcb9dcbe675a4a4e5029bea5f64a9876d34724eb3f
z79cc683a6d19fbb968d933d4d1b8e7512e1b7dbce18b6bbfb0176701057d42163ddad0fe26012a
z62a5a4f76a529d717cb0a9a90ef53452258f37691aebb1deb1c66d4495f682a31d4bd1a50d5d47
z04df1d6de87dd785fb8515ac9eac9f30d2c5d4b61df0d62b9b577b8e4c06dce86d738e7dd7b1fb
zde3fe2be6db1b02ab9fec55810ecf9f8cc27c4abeb40b666d731fbb21613de5f28f17adca8a659
z3f01ffbdc6eb18196416178016e6305891d5254a9fdab19d04e6c049a1e231260c0fbff357f24d
z84f354e0a560ac2d67f0fdb4e9d22fa55eda8cd46f92061b14853c7f0ccb66ea0b78a7a9857e0e
z2b0b18ce1abe44f4ec727efa1fe0daa51fb1bbdd072914526112757b38b28b5fcca9a373ba6e5a
z1eaa25390928d7af49f5ee918b618546c21054d33e5a19284fd752fc3a59efee61a23ef7b3d2da
z1e3a8b078e53484f41a889f2de4b87d497aef1749ad1acdfd9a4d4966f5d36372d043d9ef5b4f7
z0c36440bd664af739d082d53594d14ea24649b932fd09e6b3c807c9a732b966c5045e2ce7545e6
z2359e2364d9d707faa89837bd3f30e0a67953a079b43cab74c9805bb1a42b3d7f2140cb304b7e3
ze93093f8d0c32f58f552d48ba02ed4cb4f606f410405d7573a936fabd899a3c0c54fda509dfafb
z4c1878aff3c3e91772fa789983a0501fc720f2e7490eef1394eb9376e09233d5b184be97b8d02e
zb6ca19ec8e98aad3f67829cd444ae03fff0d5fef654d30c330c691a555a459024962d2cf4cdfda
zd7e02bf7d68501b96fe38dc7ca7c06274cd529ed552fadaa06c2e515c26252493df41a8b1d103b
z8c218d8e862f9070a071babefd1f5cde0fe90326b62acc188c9949ed3c367a1074001d6fa2faa7
z620dc3c39fcf4981042283c6abd5096c3b8db63d49815895132aeb4056cbf71d53d613e93ecc56
z46ee2afffaf7ea99972df17dcdad36c1361b132654adc9da422bcb4c6afb95385fe740d996baf2
z27c64330aa78183d7e3ebaaf534726c5a379e362309a6d5306e72fcf42bdd43a091808b6fe4499
z499566aa0acb0de5873a1308183c759c5b0b29f875b3c7f6c09ba16c5533f5792a349616ad1d79
zd8b829323b518429e937be8f55be39d98942ce8f506070be37e2de2e2071db0881bf6dce6baf83
z727181220320c06045ca410ab9878b3190e17844d158c705e38c989ba69886013e903aa213fc6a
zddaaa353d3be6c3891d65b849b8c265cfaba0e9c25b90dd8de1c243ce84c1742313faab3722166
zdb5c4afeb6a0160c360b2647ec11e922bead5f65b14b4f869f6e6bf9d7d2e9f728776029fd40da
z1fe17a63d6b4f31d61ce9e304486b0108033bd27b5898a879a6aa7f12bc1d9d745389a3a41f4aa
z96c9eaeda386cdc9d3245b74ce1bc681b240b9a8d6ead928db9250d5ef197520ee22cd2cee76a0
zc8c6ceebf33e6ec1b451089d7aeee2cbd96a2d3ec8440fafb4c17c283288ee7f101ef05493f2c3
z20b3ddd1d721fbcc566534bd0b7badefffa2b686f5e77fa0626c26ed110382d9f54e4261aff158
zba4e8abbb17bea4409da931d27741e41aff35d07c3c5d1b92aadd986ded4fa42ff5122555fad02
z12318c62c70dd87e2d6111c37fd85fe9a2cacab0ec11ea93289fe12808917e370ff194529f8f40
z6ac0763ad377d758a4862ab6af81286929bd598516a917d7f709b7f9a6f85b283960a336bce0d3
z03c50abaebc58e637037e2a3d04dc0925e2933f5dcedf0fbac855a03995eb9bff6854633ec8ac6
z674da9e09335768e3afa5299b920a669a4e2528eade1a272bc42268468efb5162ceb76858fd705
z9902871a0c4d048c143d5f721d1a2ebf16a9ff60773250d0d3a87732d5b932a7d5eeab8d1b5edc
zb3b8fec76eec85a1055d46c863d9194b75da20124bc4de2bb512d52e1a376fc92c7a9548848782
z4f743bc2d6ccf962a386fe4e88aa69155961bed604ba645e1b41482232ef6e693d2049579c954f
z707b0dcbba07a40102bf4f8e7a507e3afb378faff24604327a3bec74bed5c2a3f14078137cd54e
z3349503694f98521987478ab4831d5ab0baa57ba54a319008beba1cacfe1effc25c7fe1b17b99d
z28a3d671ab08614f9bbe2ddb0649e9130d20c146b8d65d063ca21eae0b632de27617fc5fc67490
za97da21f395f2deccf3d73b1b4a04e15bacbb3824ae2f84ba1e684c253ff095b8e5334ab15771b
z08987b21bc09c0e344e58d229f9e4967b63bb774077adf46ec5295f9f8bb8dbe0c9570bd5768c2
z61fbed27386c08fbb622ee38fc97a2b23e8640969a74d89b19e8e2d3a6ce7ecd916fc34c5fd601
z02e911730bcd132f3e7a10a81c911a1f899bd702da90c068c06a1d4c20b0a7504f2e534c33aea2
z84aa6a0496cf8a5b8b61f859d3a1c1eaba29cc96b9071609315d2529e17a51adb4a9df3c8aaafc
z27a3366989dbd4d1e83ada6c68814d5a41e1653cbb796962d67b66b7ce87169de050ae0fd0e01e
z861828c2661786bf95b4206414a5580243d3093b5cc9764d6e5ded29f3ffc3f534b1d2db8af02f
z269ade8c8da2e27baa76eed12e3773e095ae399e096d0d1c48f209658f49a3a4dbac9154ab0e8c
z23281f1bee970182ed4c560d024dcf26fa9e8d7a60dfa3cd74c48d4e4a599cb6eaf95463ef4a16
z3c5e1174f246472504c962a1389916d668567a41f8f7dc0db71ddcb2aee0979f504c02000a18dc
z57ee33f41ed0f4c43ee84703892dd807fdeb4b310adc5e9adb2c2c9e44f76b8ea83a5683de7db2
z81acf6f37d00acf754a2745e4c3daa7250c14720c5deb10d625bf0fd667538048e5b907aa9af51
zfc6f658769d05bd0265b01bb57f3998fa4bf6bc63a60833cf94cceaec5fcf0f747a1b6036b4721
ze73e32d693186c414c34961782af0cb9a02c3a3bd037de96930ad4c1470d7144633a68b087dea6
z2307830bc61c3295cd02adaa5bbb8e46848f54df9d1d93d7ce579144f7afcb0e336514a5095e33
ze4fc2f36fa8a9e92de45ec7018dff717d9e953e3e5558b80abc8e9da25557a2bed4b3899f44c26
zba391d0a5ead087babf46d7ee698c0324511d44b5f21b1ab9b04f21632063f039a6c489926ebcf
zabbd5b47f4350ca85d526a19147a4b8b7441eb0126a8c8cd89ef85ab21e113666b727b637b599d
z9ecd04b80a43c08842b8b3722003beb586fd5cae32338f5131cce1094ce4685c1f4c919f0d6eaf
z0e34c7b96b2a944dee13c18ce998bc684a28411de5420320445d3741edf4e7bf6e2ef9d72b315c
za89d5578956effc1f84a4ecdbcc500db80bd9c22fc9eb24e4d9c32782b412b6523e4283b1e546d
z982d1ada067284faaeb3d77211c66f0842d3182c82d6b8493a4e2669380d318fd6f6a476c52934
z91d8f224c360186d5bf317bca5398318a79ca71e2178506a0774506ea200972fa378dabd03ab52
z246422848457edf6b3bd158c519aa9cca6a9398e33643dd37370a9d62fa6b4476813ba40c5a297
z5b9e62095a2f75bc8f58c3d24a0ce705188e6f31a1ff2edb50446c6c60cefd3ade4342bb315e38
zcd9d468c833e211a9f3d46dd1b69d62813caa70eafae4abf30f40c43526170d395580b299aaed8
zb93a9a08f57ccca4c0977465e064443f4c5d8ac1ea4775439002b562b1cb19205233d5d02929a6
za14ce4b87acd23a97942db57561b878b778f2345655ad7a5e3c755bb16799f9cf5ddd5ca47d68e
zd1840dc2051497b95fe59c8f526123554a6a6fcf460373b999c27ebdf03752315ff75a3fd06736
zce18a2b273c1c48d5a1ad8b4100347b19a2d5114652881ca1a2ed496add67f765959bc29c14ff7
z5aad2055b8153ffe7a2364bf59f836d6f0abc6fd9e5172a44d151aa272e5c24fb0939b7ecdbf68
zc6e7d573fa7f491cd0bbcb9268a9f9bda1c009ba9e144d36d68335246274a77e0cf56114e0006b
z73f571b76b87976cb0992ea3039848c84bdafa6af7bbfaa713059040a3e88abe16c95708463492
zeb555ac9f5e41b79358ffc95e8a8565ab05e7471e5b42dd4cd8ee47efc7755fccf33575683cfe9
z75782a553a67fd4464336451ea405b26f8b149ca8eaef8180b96d16f1f72aa31c7f9ca0bbf53b1
z7c46c988a5cc4e2331fb1720bc7485ffccedd0560da64ed6d1744ee66ac3789354ee619ff518c6
zeb2f15e1e6547e36510062e6eb3b5b3b5ae7bdfd38daedc6efc3b8dc32435431aa56814e179955
z37907e856b95ff69266aedae448638b0abdf2678655c2542780d74dc8db2725ab2bc847f65648b
z24e4649650ed467cb56c8bf23ae19a18a7f3531928a69dfe03d30823e0c77c1f8760f5411adc48
z307e50a42f0865e5f024b57c979dc1c1e114e3d0f15339b486321fe158ac41d047abbd88a03aba
zb7be9843232a03551bcf0e15908d892f82c227213eb7934cac2ca7633f5bde6374daeaf9cc7903
z03a9de1ec7324ab64afb2d22a5a1c149361c98bcf387c695e5ed335108f00968266cf6c123f384
z5bb942370a9f3d016027e24ec8a09271191e47e986a71c25d88c9064d40efb679d3c745bf3036d
z2d4cb2af3ff917fcb4c1d0e3e1b61d49acf7293013b7943b66f789016621e24a780e8dbc03d210
zd470fe660a842c4358bbbd166cd733e497be92191b1cd15360c060c5e5b0dab9adf8d05eabc81a
zbe3acf0612158e1092e2a0d1eca3c0587c44262529506502be36551994220b7ea6485e7f8c2ca2
z9544198e8b7a3bc12a0e51799ede9002214912a3bbcbf0809488a770f66032885692b5c2c964ec
z3d36b9a6327bba825c8d3dae8120696463f76b5513128325b0aab3067f107ab258c8122b276aad
z7a6772ccac7c7350fc024df1782ce937ec5228a7a435638cffb700be51da92476ac09adeef2a1b
z451aa7caa96c31552b28cc6a585b73052d160b8400767423d595bb8dd3b1bf47bfc6ffa3fea826
z3a2e6626594d8f8ae83e668ae0043acfd9d9a221264f3c0881700985ce4deb655ec5295d02f318
zd45cc24d7d2386cec154f557acbafaba2ed43c23056a57ed7297d7cd215955d159a7cf8be42251
z279500c8dfcf979fb6193431e8b970a40765864dbc3fd8ede3bef89a0669055e24522b6622f2a4
z4a5d5f3bf8653131f83bf9d4835eb46252062b4e7544d54b97eb57a63b08bb38b39752d9c0d370
z78c6a44917ef7f8ffb03e8e5c1c4301bc096dc1a0dc5c545817dc6a4f6b995ad5a70b2f5e7b0b0
z0abbe3a04bf84b3f3eb880a2d77c21600675a9402d3a2d6d868bf861d842322971425d8357376a
z6f169cc119e73630172006a7bfe00d1353b1d34fd01b8228c8219e44359fddaf4871eeb450d1fb
z14117af3df75c0f263965bc4d9de36329a06d601d814114cfc0de951b101643ff00a04bce4bb39
z83ed262ae3bc1076042a66768592e3191862ed453397b9e48661aec860f6ea318234e08fd97c50
z3f3e81f837d2b333cf348a0a198feae8fb73176915a1f9f0b04b57e9710f67e3aa60546b48a46a
zb336b2e0700ad11d4406d7c1f866f8cc54467f971c3e3a4d6a59758a746be0a7b3f9149a7bb2a9
za4c4aab537bc5deb3b888fd75a449d32c1364a1388a29922ba9d435fac86e9a4b2533fe1e6e7b7
zad8f06743a9c1f00003499194afa3694feff546fca4868208a7a8f5ab459ff7430b6cbdfd9ce0c
z19de06429931dff6e408bd2e6da08f71b2e6bec161ef6af933cfe13cc3641ba3798812757c5c78
zc7d5f7d9d2d76c140e0a74eced309c06b70ba12ee42caf556a0bca3c27cb9c4b8784b5143d0821
zd56a35b52ba9ccf939942edf701c08666a7fc8901c12bff43d6f9cef1067a35bb3a8954fe8eb9a
z79d21ac0014dd3a92dcaa664ae0a9037a7118395f1e9d738b4b8873b00c8c1af2582b57ef52533
z5de4bfb8435eb4936345ee24a1f93ffe57c5b2ec6561f5059fe46eba6b90d83ac6cf3f797fad00
z3265f450e069d71e1d7e59aa274703cff9b45d5732da1a197c23892ff20b81f081de5ec4819054
zb650bc3d87bff5af32b8b903233337ee5323646b90892b11c4446630cbdcb1649ea404c41fc0cf
z95459ecd04e78a0e44cca8043dfaf08290b76760fe2b1c2d5565f23f31ebd5e6762949f0d903c8
zd3de38bcb00b86feb161a1c9620cf3924bcc3c9cc856c8780b7545143365b4a80a803d55dcc9b8
zd9fe4ddb50c7c8034fc58f58be80e3222905d57c23d643bebb5ed73551e5e84c2404f2a6bead87
z590b3af4b295607362ab0e215c32520a2c7077ec213523014d3a9dc29ab88e616665607ee9b9e7
zbecdb7792f14a7a8437c7bd62f6400bbd72decfb13e70c840b1bc022581cf7faf8d38021d4dba8
zc2d059ebfff9ea8969aa49256485f0c8bd3c38c38afb1f6ed5d830ab800bf3a071c838705db5e2
z16d76a7b3400d7afbe2621003909b76e925cd59e6592da5cca2b026d5fd8661d8f365351b2008c
z9de10082f06744e827361a98efbe04803a4fd8f18bbc2f7ba6acf53c888852db7b9cf78fba7ec1
z07a246ae5fe18dfcb693223fed0c725607c66083a9b4a42f3c886d144a30c404f6fa5a91b6baf6
z13c14fcbebac94e93f2ea9672e2f6178f383355a2ddf485334c8e2631b790cedd3c473333b44a6
za95ce59a0156a8d76ec687f50d5fb27f9535f03f98902ba6994dd7f7d4f85c695d921f867bead2
zb955fb0baee193e9dd6e56b40bfe7ae2c0294ec57782f72ca69b6fd62f893e6d286c5e3d37eab3
zc51d17e2f1ee827c763afd29017e113caed43a9bfd65696252112e4c52face8c245f3d0eb9b79e
zfbaaf84644a24aa9af31056fb13eef577ed84f1f9e4b80b00e2750db23e19a0f1b0e90333ca4da
zc32c0ef97deecee95b3d5fb30ac355d033a7b829dda901626fdba2e033488c9293ce0d9086ad8e
z993cea7891ed33186d9d4c532b36ec3deff16afae6a8c50420c8d99f1e4883f835623b6803c903
zdc5b761d59d216b8801c35557f7db8771f05365333d6c73fae18cfa0021fd169cd80d082d80ae3
z007ffcf845fad8d1ba4fbf1d8759bf7ab622c8ca1868f91f3395e6a3cff19a415b32ead3595c59
zed9f62cf8555a34f2e8368dc7d7bd9a3a9a34151e80b39ea7e00c68b06cb9db1e0e7869493afdb
zecb744991e24dd926848f7314ee4f04f638c7841c525d05604dec40bee76c8ae5ff6defed8d060
z375a8a8617268b12baf255adf307e6299c92f830404aa782136b3177ffbb92a97dde4322b89fe6
ze95b5222baf03e10ba6421050977f4b83f89340865bb14a4c03331f070c297f30b19acf507ca10
zfb3c0dddea4ce3d63c449ee22913a0f242705ad5229e1836b3977f46761f62023bb3d1f0e697a0
z41571bee7f0cb7d41c5908d1cf4a6494c026efd2de49e3d0a872fdb6c7db1a33ad95819a85b85e
za2f36d913460c3671158a771b8b5f5c7796a1ce1d4ff72df4109f35fc7e29195be19e6268b63f4
z6f7094e3e4ba69abba53f87cfe05feb8bd1804d75c4590198aa582030bfe732c529e4f01cdc9aa
zde6bcf581f63ca845ef90294bbe70bee075b8fbd1129fdb1b937ed98a7d944a1b792d84a0554fc
z69b34e3b6a81891781cf967ffce1b6d510d9724bfc7eb29cf54324f2ced7e0c9b9758261c742bd
z7277829b57c1203c2cd46dd1c2427ae5e39fd9b339020cb57926d9e1feac0c0acbd8e4bde2f68c
z356fcb08cce439cc62aa6d86987d1d33cf905f3ded70f1903390c3fa0464947d9ead42b405752d
z37af367ba433beded782d4ecb830d53e48be59a9e0a1d03762e7947585eb2ea21258c01c9b397a
zf046571e82ed58f8b96ce5c02ef683c2c0ca9ae6acfddcb24d997f1a11bfc4fc216b9bb5c3ada4
z02802d6ce912883d8766085cfa57f6d16335c53c87d05331ba25b67eca84df562136a21dfaffe9
z745760769fa36df6fb063e3d574658f65a718bca85e59c884af875e00893877d79a2e58eb7c969
z51d46420373fed56124f691aebbe0c29b0d99080c5025240a269d76fed0522b7345c9a48431c8b
z38331bcdacaeb0ce42f681ce405e0993908c49858a434d0d0d8a334d4866682a9a8f772bc2e052
z6ad981d823001db1784202c1b564d5ce689ce38c42429a8f918b3cbbf65d0a2aad791d479fa5ec
zc920a5477bf117417d09966d1035dec3900726fda00306cc957d86cea996a189ee640913cdf76e
z5512e790f1e38e6910a9fd2081cce9cc4927731b37e2f30b2b0400c36df507177f72b1404a09d0
z2aab55dfa2c608bcb171131af8557a34e79982744eb726f9f4bf4bebd431587b16937033d4ce67
ze296f6c6e6939bb1af38aebe3810a1229e83abaa2a1fa5a1e5801e325c329929b88fa9940fd075
z975b39b65e4ef6dec60e16a84880321b9efdc271128c96eb636cd5f964868426e999b452eab774
z0c4dc7b699e2ab05d892e9b4e80fc6863cd6c25606fce2a00126966b460afb7973462f035abfe9
z74aa90708fcc2d18f497ba83d4fb70a58ab9cea34471212232e00bb3fdc58dfbc1a9cb9deb79c2
z8d571070312bc3607bd2f6f55d71818d315f983a2d3f0d3c40b6f4ae8704e1d8cdbcdae14f75e6
z1d524135c32b7df238daf146119f40f0664836d4073595fe170192f1530c1ed1a2f4e5037a5b75
zc2913819ace77f9eb2cb428d0cea3e1cb5fb3964224506f61018b188ff7c47f3903eea9f276331
z69749a65eeac0b808b7f4ce875edb09d256cdbaac9d0574aa9ccf8ba2abdce54701e6e5135a1c5
z7db3cdcd6d78fcbb6312c6b0685df5505a7c13628471a31b5f95136924fff1f404787dbc4a7154
z7a23cc87b7ff97a464e9a302057210ac4b8a0040215fe6f716c862e687b4e27babb24aafc30f4c
z61550a5ed6c84e88fed5102e1e8d7ad18c365fa6d48da67dfa8895e9d0be676b6407e5a3f7d7b5
z13c364c47d8fa509ed3372f9df88ed23a31b37a2ab57dd590ef871efb484eaff5cec47ce96f3b7
z9b7929b8345f1d51e5b17c735fd7de2b0235e4740f674ae3106d69ba4816e358e7f712dd01f42a
z706d4fc125eea37f4b0d5779931df0378e0847b8c741319c30a2f752cbd7f47db1fc46d87083c9
z7121a2dbdee8559242667ee72e56b5c0ca519eca0c27e5926ba43e5f89ad5bd0c4d84e35299216
z8923b43191f9936b3a399b5dd751a5e8712657c31a190be81f380375f63f8f0fc6b7612320981e
zcb199f912d1d99232d2a3c610470b8812508b3dc1ba05068f3b40da8cdfe58e75b3140fcecff1e
z05acf8f5fb892362eef0547469a435459a287dd6f150b2c33362f7bd6b754ef6d6dde7addcda79
ze366d4efe93125d3063b15d30f0f94ba511b04ab1891282fca45b42eec42867e69d378091b0cc7
za8b05d447567eaad38de275e30a4204961bf080b6f61edf28df2afb30882379bac717de6ec4f83
z2b2e072033f375ea1284fb356b5007d9527a02b962c7c7f0dbc3ce3ae08c78a50b17e466ea6657
z9e139d469bf2c6cf5ece3cb9e19f97d531055261cd8f0295b94d5094fc24e50fd6d2545d082e80
z1b7d90cbad0709f1a7e06a9d67981cc6cd75d7f0666d722041f6544aa7386d992a98be9a5b26a0
zfa7eea99571b1d12f568c08998493a526a11708d8febce76cd746dc032d0fbe15432ddac0324a0
z5bf17ec00cdb0e88920c95d6dbb4d11137f9a09a3eb9360c754e9ff146302bb51a7b535e15fedd
ze5db7d0cc378dde67712666051f67e13bd3b5818e230ee7c5466019e61225f251801c5225cb92e
ze3d9ba1330867953c6539c70d8633de1aef0e5a19690c6de67e6717ea0e008bdcc55db21ccf7fa
zdcf3d7d56c489571cc025abe7a48fcca0128c80c5e44b5f9aabba1d12d37c5c90ffdc98650b63f
z15665321663a1c06c6bc837c4ea6c3ce2d9384e956324c366eb405899b38ee9d16c1929d69348c
za5db16581264c66393c5995c34c4e9ae7cafd14310ce1d7924262e8316ac73d85030eded73182f
z5b2721de323aaa808858ca2077da8728b7715adfa5b162ee2a4f0fd05e08790e8c46b040136a7a
ze4d753568a3e3be6313d2eb239b187c307976c2cc18be2255d02c9eac2ee358f2ba1d67738945d
zcab325d32789cbf8285642c84bff883acff4451bf451132156ba81c39a8e59fb4709b55e042b94
zaa6a7afe81fc501bf1c7adf0643203c2e0a207c00eab0e48f31c90a4ddfce22bb056fb320205cf
zb7dcca6761249e5164c95de1f2e773c1fe26b0a305d98778d5d698db3b6a78ec2c5bb8aa938f02
ze0e0e323356db658689fe22fc4ca57a19085b420af8f4157ec28018c864a390766a891d753bca1
z6512be0894bfe977c9606f8721da3201605500f551cc72a5d9b1afc9129bc2de7b9644ca341b05
z7e63d429ea5c7f72589eee219c0c9782f96968154ffba93a7feaf546ec20d047811d8ae131a743
za04207e413fab7d74ebacf186b23b0c20f12b675d3152d2eefe553932ff1615f8a23ae123d1190
z1eb8931f23e410bef8f9407f5210ae355d9e881eacb5959b35948bfd090f2572624dee64af7901
zae9deeacf2b3bbd38148b8be2a7f6882621746459e0a9237ec833ba2732d28350f7201c71e2abe
zcdd1c699349b518a7c10bb10abc2f701045f780379aa23fc3f53abae3022058be048d56cc7206c
z0f33a21975d31f925ed78d1b985f10b33a31bd8f5bcce871980d03734c4888259730952229f9cf
z421990422924b4f0b15957f1080ba70cf8868484cf2b4d94bf56507e5114636def553a2667e2b9
zc5c6c6122d958629fbfaa07cc1622644e3b99c2d74e8bc48ece041c78928b80c9fcb99ccb79da6
zfe9c19160d938a6ae59040ed5e763fa118a37d81d45e7ea091fe048910164fab09bcc233ef6ee0
z232648b8b0e5856c380e7f991c6e059fb921b4a986a16fe33ce58fc2e242a98666428815ab629b
zb4894e5e8fcfbdc665416492b8f452d58627b7f00c5630c64368ec21243cd04f909c79e80ef701
ze91a034993c2ff8072766d3febcbf4760bc397900264e55013de5badad7d7fbbdd35c2b4e9bd35
z34c6f9c46e2177ca76dfc8023e74fe8ee822c410b1b68f9d9043574741e7a5e75e8464774c7894
z6bc6d00074482f26df9149beb4789ec790cbc5c38828f1c70f2d54e5208a9fcf19acbe70451a6d
z0d511cfb90d883793e60eef37fcf83ab928d232306ecf0022920d6385a07a1dfd4c3cac8874333
z0987f7e248a6f7e9d2ea2fb942dcf7403f5e23680389cfddeb9116fcdad66636a68efbbd54de93
z0e4c108f76a7b9c91ebd25de80fa56ec7cf19d73141b3eb359172b969735fe5a14f3bae97c874e
zf9f0612922e0060cde28a4e0099f3557852729e844641554eadf9942fafcab5fb15124f21aecad
zd6e7498f0db39114024c2b6bff40c2cc366ce45a3d4bede0eb76d48a41b723f767c2297fba01b1
zee4212d06803480cde31c398811034a7b2ac67ee04f8895d1635131aa2562a8801b859deeb6139
zdebc2252ed039363aa20d08f7e6c7c2e2b3959f7c901c8314ce7c6d60df04a7f7f7f337694aa85
z929426ed99dea0397986866c8899b334fc66bd0e0a69d6e53f64951800191af120d6303f14007d
z3a5d720cd1e95dc105c4b398e944bd7b662bbed8a62bcb5464fde31abffec14b66e5145a2db2f8
z924a78576d9563ce9277f5e864bb2517d46434c70df19378b89e9a174ebc304065764094dae7ba
z2b9e2283846c0c7cc45787993f7cf56f607a1a71174f741e03587945c2a965d76036d4492681ce
z887637c378324828992ca489174a9d2ae841ae25ded0ed1f851901e101ec4df1b314518967095c
zf3d8af5dcd1f60e743ecc67fd546a445918318ea4435c94caf75fee0c4c6563185443be7d8dec1
z8c7687c5d0d258c1eefe9a22999ff0feafc01b12042c647bdf932baa41839d6b6499c01eeafade
z1a67ddd9edaa668a715cffdf59125cd787ab5f17b7812a3ffddc693580ad0d28c52de28f528e13
z34c483b56daed45b949f44f63b9fa7bfe25465be28e759902ca74cc1062de7f9b53df8546eef80
z1f9c4e743f0bf7c611e9b48a3788cb146c447b117db2113c08d3b496060a7ca176337d67d3fb93
z0f74defd7eba12fb2b9de5307f78b9670c1db74d8bd7a769e442ddbad7c6ecaebbe4a2d0331bda
z99542f9ef7bcf1b25da9712eb0e824c5f1bea0796e9c1cbd501dafe97cdf7ac48c9d33e1a38311
zda5d8861495dba404986e7ab42250fecaef5575b33cb274054184b326e3d45603a6bd06229bcf0
za0d807126a5ef32ebff4ee6cc0ab5a35df4c79baeed9ec13b5757ed1fdc317aecb4c17f615e0d2
za6a585ffeabfb53a7e2e51d42a41d5b27d7e3b12128872a04e26a81dd9ab9ffff95dd297a3e644
zac7d9ce8482ae656ad843bd528d1900abccb03d3d23eb9eac77831b3c5a962bb9cd8888f94c4d1
z837daf5a522e5356bec087582e3ca00f43d9b6847b474fc734105348d7f850cd615d22e194040f
ze76ba174897110d4c618acbd06c4867e959bd0d5eb1b90eafc13f4a69b49e9af12aedd56efd4db
z25ec0af6cbc5fe9cce811803b5c9620b23decc17eac5a595cd327c977deccb00f3730c78015825
z558daf08c982a9329fc6c9dfae713985de8116d533402fe08cbb7d483d979ff728d1d56acac869
z3951e382dde206644b9b8a721d581bb849b0597eac476dbe324f5906a0ae34cbef226fc90a5e8d
zc7e44deecac61b1f2c8f33073c905c31de2a94d117ddc6ca8329b3bc9e893400845f8494692826
z92e7979752c4dd46298fc15fe6e8a0696c39e5445337b7e5f0ca748a52b951ea35f44386a567e0
z6fc8a1d329ff81d26699909941c7f6039b244cce5bc3d6e25c72f4ec3f43993a35b2c95cd78705
ze2208433d6dd7ab4ece059da6511371602db8a66d4843a1ebbb5724ae77e8287b55546ac7b63f3
z093656495f4d999d9a44c2196c2f8378ae362d47f51068d11a0464d11102c4c38aadd3cad013b7
zae96b8073335496af34e71f5585b79d602e91631d60aff268a8a0cda5f05696a426e48c91ec078
z23314f8324e996f3c4f2a2cc6a39ddafeac9f94ff375c347aca2745b046f4e2df103d10774edb1
z6d690bc1dd4eb20af66a5d746fb264322ffb90c7bea5d4b55baaf8b7d267d447eb21431ca095fa
zc8ccb8d38f0f53856dc5af653de1f0d51f33ba5e7beab14ed0237e4f047c35d05eb6c0dd514b84
zb2076db8e857161c2812abbe1e17dcaade533c4299dc381c64348760c2fedde8a077ce6c915abf
zd38b70371eb1e4ca7423d6b44bcd6cdef9c2ed6f6321401d855e4409d102ea7d7b7560c1cdb226
za3441ad2182dbe1e8468ab4eaa88a5556d0291a32fefbe36e7bc269f30c10a3c01d65858c3a8fe
zf3bcb933bc1d25732d8b83bf748642ddf3e52facee22446ad8cb7a1eef9005bbdd2ce8acadc0bb
z9d7affe6369f7034833aebec5ed8948e208f1f831012d95aca7785047adc8a2aab5c0dcf6f6a7f
z959ec25993c4e0cc85142c4107a8b2a8b7a1bfd2c002d55b4253586dd5c02f9044e30d70c9bd75
z3044c97eb586e9ea0728071b7623216965c9275e5509a1863793c2ab8ab03722409682e660fbcb
zb5326999df3ffcc6d85a112ae85e8854fbddc459be6da658635c18b4f8c9a53e04f7f3fa135eb6
zc16ecff8ec1bbd1213951e4ed70458fd3d116753188bee1105218a43de9d6e34d12a417c11f5c8
z69eed00725f2388a8d4e2f7fe2f47f11cfa623fd74690b15ef9b3fd259a5b5344c2fd54fc47552
z4efff6cf71281d54eec6de311b47f0c103a3b32b4fb1f0f6ed5e871b0007bd33f6a16b2a96cfc4
z20e43df4753b45ac13df04ead05b6f65e9820e02d87445df0ee8455709e2b40cd0830da8bb900f
z0e9b2bb27d80b52eb7067b71ac96e5505f2870a5c960eed606482509e56e46752426f47b337fd9
zc474061a629c2c565ad5f81fe80b9a4e0b0636635dd51288ab96354a5576e8f67e0ba49fbdc22e
zf2c723ec37d272af2713b34243da27e302ad92b5253e5748387090c2a9135fc1cc659e4b1b317a
z5b94aa7a5d58a91d7a1eadab43aecf432ca8cf105c472ff8d64335b354d265f0e31693b6bf2862
zf5ce50148d57e8e741e6915c5c2afa5d91af89ce7e5b142236e2814ce99115ffce4b857e687059
z13870276c87a9afde8573dc21232c145e497c577d1a28e34a091491f58605a71152473de6f238d
z80bd7766718ea9bc286c2e6544c608f8bd5a9f7de63f0e2541da8f3eb93a96bc928900f86eedb9
z6fdc290d235e0f2a82da850736dc03522ea64002f7affed8f56f9c64855ae20c20c40668385df8
z89a4dc9a702851a201335593be802ef4f08ed812cfe2b97532977b509996d87751939be6f30309
z4e18151d50b0fbdccf58f4a3241f969e763caedd9ae781c2887c5d22e093a54ea51883b6145b43
zdd89d3d7851e11eb2ec56dd026f8dcf13d83d918f359950d28200429dcd947745f1ac0d1ee98a9
zac82898ba97cd1ac9dbad6a90ea80a373b981a2789c2592470337cec23d6b12078fcc9e0d34503
z8014a49612081386b1f48fa32c84956963292d8e6763f17432e7aaa1d67df8eba5c4ce6641186b
zc345cf72a12dba06bd95f4e138e271caeb38f3d5550b391708dfa2f695ccc2cf94891e155d9140
zfa91ff84a09ee9c14171a95229c7f5d3757d27dc59deefb1d75625d92398a25c8261d0818de863
z477a87e85874ab7f4023967e153d65300cdd18baff0179f36d15746e91be046459b554d9dae56e
z54eb070ecf7c55de377fc01c614b8885b056b28d79d3d1dffad8ab6a8af78d869ba9d0ea9efe8e
zfd39793cc8b53dc0dbeb6360a7304a4355ce383b021f3051f0112e0c22e5fb39872dab64e5b951
z234c37c83f275f01de605e7f8e2b73dfd146bd52d742bc8fc0e6c9a792cab8768ad2fbd988581e
z86ca4538b79f9edd014cef65e6d3b29bcec40c5b675564385e11e492b5fa3774409253c4aa4511
z444847660037e2f899e31b2727339c70e2de4b71c86f9f3089c861faa71196da72f64bb33cfb9c
z7c4868ef5538de6631c2e32ba562bcfc1067109e75d2915cfbf46005a26c6ca57a306f0e9c9b7b
z82e76cc426d5edbae5578e53ed6fefb6c6533fec0faafc0e589feb6b0a6a3822fdd625ee042928
zcc309d3d0b962345270151ce2dd07b7f0f0bf6328cc7f69f8d1f023fc73797a45895d508c2275c
zf66d541aabd240fe0e4763826eae41b932ee56fde9b284b9b091ac7019c7d64cbd579c7b287775
z40b87e89b70c1f8d7d2d1b4352845d4cf199344c06e7a14dafa8cb8469f5b4cf9720f41d7e4169
za36d6bea6490c125fe40d344501af1ed660fdf7827c2f55b038b14c965f655a25bc448f4ffb13b
z145d966d049757db87b30be0f77caca71add09375059dc79a06fdd051674f7393c375c31342d70
zca6db53138f743b230b7436a1f63f1ab351b3c0b19e79d73115dec08af392a93d3a8c0772fadb8
zde63519b61f13cc38bb0dc6f3b613aa09966070784c002397fb73ebecac2543216c301c69385b3
zc227fced48d89a7ba55edbec7863a54f2a69d7f6e8265b3fc5aa72fb784d33b4e834d4ca5a97c3
zd9a450fb8934caa388c5f166b599dcc9d51f92919528a326a010c1e50f9af76b65090c590db780
z7024930e34138e177ab96db3f11f6137001ed03cba7c55bfe12a6ea99f641346834e047e4f120d
z146e59e4e47034e999dec9b8054e79eadf7303b07e585d38b1ff453f1f237166841b9272723624
z85754efa6e530c203a1337116a028596203de1c1b75b91a16898ea597c8e8582c1f9e3bbeb83f7
z3c6a2c8bdde75198408e534a59ff6b32905ab0402f7fd85f507d3ef2c11c338d55de1fafa4f7ae
z7dc04e405d4ada7c7dd3d7c0c586b5b831ed6c6e5269c830e6a10bc625f3db539f6a6e1587e905
zc07e4e0e82f12f0ac831291dfb40c99903055cbec882ee467e031b163b858d0c87d7233eb397ae
z4f9192fec9c9251c5f2c0591eff128610f80eef28c1c2f69c03bd8f85d38a048ce5630c61ca740
zbff510159a96c8b16b8c4c4ac9c08d5fbe8ca593cd436d8e39847f094d648264aa277809a04c5d
z2554b1a2a069d99eb2e66dfae10928fe4490f39621f1aab43e52faddfd9444f7460cf16cb7ee56
zc8b9e8a630fcd308cf5baa29f1548b2850d14d65f09a476df45dc1704518507d919414798b382c
zf72791a0bc7617d8aab1cb36e2263834644fc5aa2bfd9612af6149f622ab9b2e37e792deef7665
zd23bf6a5b02b9cbae933311ad276c7c491fc66992e5f640506bec0621cd511a5c57da8f4021d3c
za9d1fa109e2a9f8b769b6b2fb08e44458f9283919862981ec4361000bde7be321222d970f2e00c
z265b6aba1f98dd7b035663a658a43006feb799d0734500edc4020937fdb5932c2359637ada327d
za250556b6170ba2fc2b4e8577d97d4c9084e19ca5f99154788c40ed46e72bd76ed9b377399a810
z0e8479cb189a99963174372258df7cbc41ddbee5e29d9241934332198023dc3467f439010ae0ec
z1955936dcbb5fe6f66a558fdca0108d612117e76d8ff4f85c56b0f2cefa2d6a6b719565d408705
zb4789d7570e12ca71f5ebee8b497d35325ad411b76a60cb7239f93f1f947a76727eacaffb7cbb4
z04bbafb6c21f5be0d307ed819b60d3dc9bffed1558ea5f6ee3fa790625d45951cb2805d842ffd7
z6259ddcff8c77401c1b4f8f68e9aedb7c2b43a3336a310355052894ffc1bc64926ec17bf9b3d05
zdaebbb7ae9d5c9a3647516e54630c58251a7aefa5d8cf07e27d10244c0c14e2b2a57d69979299c
z3a2148a1f655cf76c9ab34e4e80c42871f18b99a951934184f3df60c3153c30eb74c4733658da4
z1d84d038d01570a407f21efa5d84619040340ca73d6fcf83cf6027f854654e4f39e8f379613d0a
z22880c941b9b281b3c84223107ed7563b820485b4a259eef59aafaca82d9bff22bdb6319330e17
zb8c43b03796f055c745beb0825b11cf3d4f467e469614cf188d3ff90ed7d8c66bec453965e3b5b
z90f9cf087db1045a37b8672ae32ef69daaa17b28ea68897607aba16a4f27fa06bc7823b0201906
zef14e7d83b6f3e0666136d8e99447035c3d0962314d5360bf4ada3043abc1e0024d5733ddcf57e
z8139d82299f88dd29c3f8e6e0371aff3a2e26a22361b2e00f59aa95e39c13d6b40be7c41e2c35d
zf24357c38a08eafb2aa1b360fe128f49cc2fbb25b854b55ef5a36f9cd6387b3948c368fd397b8f
zd6a5da24aa51b59926c1136cbafd445e0fa638b0fefd1772c6c56fb39debf700129e64dec67e57
zf57472fd69a9b0f172bab3c39da8ff6de0df2d67aeac161a60256faac16ea53a0d7abd279fa855
z6aebf5f874ed08bbc2ef426f6dc5bfcbda96c14fd40f6362ec95faa6472076ad4807af81b10178
z4a7bb1b40f997e2ad4ad88a9af246869971a5b190a7309ac161f0fe82c5f66abeea9f29c05e96e
zbc7175893f873b6eada94add2e7966b0f8e0eb0343d66cc8bcaf1aacff2fe573f875ac1efc9557
z5075a202c8fd1397a1f4554e0aab9867a7c97b9e07351a9c4372f1d9544c435f40d3cf7c6f45e4
z29926c554228bfa9cc491cf095614bc25be0b2490de2f79a72406dde7ee9ed3f7698fcf281eaa5
z2cf38cdafbf163f220d77cc7174fa3e817adff68f1ac856d59bf6505d67477e244955a23e9e4ae
zd19f0f3a2abb9f4cd868ba65acc7f42ac5ae112f779172fb4b07122c4d6c7a393da9dc6487babe
z48dad732a3c64cfbe4c2dd2c598fe71b624b41ca23fa2db664591ac7e413701e09845397f6e0b9
z8c96e60a4b11178e85ea5fe3a111d25d4e338a32ecf4e3b30adf882c1e0a1e70f735a36f56a66a
zad90e9edf2d47c39c7571952bb644d6be0b3852883f508ee6794b9983193c9af75c7df7019dacc
z1b9f4ab7ede4a5f703fa22154c1d3b8278bc42b99b96883ded7abb34817e627c879bd0d846c17c
z3a3d29f800ea68c3da238fedd32b7926b12983dfd862f5b4465f45fdc7cd45b61829c7b304b5b5
z5fca3c869086674bd8ccd67834c18f6e73d09bacd3373aef05647713300807f5a0470c89a7b05c
z4d8b39794d9da0288beb4628405e2d7d5bcd2a13a4f3f5ee28120c829a637f0479a7eb862d6b60
zfef848bed71f88b9e6051013e87f2d3b5d11f70406e322a127d536f652811495e43948e0337aff
z470daf416893bba089902f0a32d786dcd12c142db174bb1fe4c9ed3105fb873ca6fc131c41ad47
zb7757e6f251b4e1aab3c4189d8809bed67a3fad67bb12b27ff6eaeb6757d5ec71efbab583c0899
z02414eca8f7c8cc81971151588862e665e659e687ebcb2edead2907bc32882db8752af835153d6
z2ed768322e3ad5df7ca6cfc73b017ddbfdc4dcbd4a3a8eb4dcfb94244dd964a9f8bd8e9ada6d66
zaf8a19cce8967bebe2234f329445be6c58e6a390c18d250dc86c353301618d71d953ef34ac4253
z67e1e6d844faac76daed1de0fde0960cdd7b5000c1c284dfca4d5de857534982d812a65a9d7c7f
z7f691c241ced7651aa47620ab7c0a29dc09f94437233ea53bb23283e02f2b5bcc933b19676f278
z48187e00698fdec4957a4d734964cb588ea5123eb9564bd2ed1f66fa9f70e78aa94b91ceff5864
z175dc68bbfcf70205e79e53a4d7d6cc94de98bb9af1cd53803f4382fb4beb27401b7966a4755d1
z53a5d3076395d34cd170c17f960de18a37c6aa212aa13721835b31a7cfd215c84b089f94637ce7
zdf34c74f714f436729e45c5999b7c7f2f802f31b9407bad50627a2fc9287b8e612174cac47841e
z85512a382c52f3e8edab8fae252c0f55a93d17ef145187c246d065f934cca275fd43d8e9121fa4
z97eee0c6a7f9fc138984181a44ec39fdc663063aa48066ce1685a836493b1a9d6f78347bfc5fc9
z00d2dc742d0d2bc8ae6df2ad4857145a57853d79fa4f819c52519a791353e3e69aa456e0da7f34
z84c4c1ed7d4433f4571822253d355c11d6e3d0ce7e7d718760fe4ace35191d5d576046bb159714
zb1507b40de29c8e0766be925e4d71afd6c5ad4424243eb84ddf66d7f4087cc4aa347da0ca708a0
z4612d950954569924917ae839b875f7a499290f246aad95ddbd8985efaae436d881819ede6c901
zc86cc6bc92f7615e7e999e6069193b5dec4b3a71f45eb7149b6d74e874ac3b02ebf28860fcc2a2
zd96b1138364af4ef943e9361b952331ec2d4e9bec6bc19152793f7c48b0cb0ae9fe682d19ca427
z82e7ff0c07b8e729e8a8805d7c58f0d23b5504e2b480c7fcf199bef18c909e39b53098b084f020
zedcf8f103dcef8dd49220d5d92f305c9c90afe0b99ed0676d4b49aa3a1e6fc904ad11a8b95703d
z44a7b0a3d5c09f201d696b7e4cdf7cd910c73d1641d65f062c04ef460eb99a005edd53e8bdbcd0
zcf592aa329e1d1cd84c119efcfa4b7716b5494f5900d13cbd03c3995fad21798d9084388f2a3a0
z8b9d32548cebf031cf2b7f549d4e0c4f25f08ec4c8cc7ea6814c6d2b1846ebe4cea657ca5d5423
zcdc6882b538a619a6e10426d35e73eedff6a6be452abf01d4a9764843455a4e444e240b43150c6
z3f4765501d6846063039e125d803cd9adedaf03cd057ad817176034f6f590121c5043263996e18
z68471ef62e426ed79d171026e388a26b4472cacdf69f762d4f49701b269a801f29dba4d75d31f9
ze5ade69b6f5d4a97df602d717fe0ed4e01366d3f012848453d231536e6077e1a5934fb0a1c3a22
zbbe713967582274f82490b071a94719743a1b68fc85906abf1653ab7e85c064af593daeeb42510
zae061b8d473cff54b8c0ee1954a03e2b800841769c43eba1201e0f8ff2ab4a7ff1628b88b736c2
z54f2df5e617c69bdf0997c166b632955a1cdf83b6005647ce859a84627b28f4bb9507fdf79f044
zeb8fbf12efcc86e1ba1ad50d17ff83a5ee248f21eaa3aa28959d631acdeb42887f30b2f58077ed
z7051784ca5d301a8af6090464872b2e4e2bf50f01c79c53f9dc9d676c7e667cd821606857b7e04
zcec4fd5b981e6891312ff86d4c440d9fc233356a9ba6c5af4401287b43dcef5da1d0979e9d218f
z7c93b0af5b269b6551f27474a5fa18c9b10dcc2871d0dd8d061f52b5eb8e66f55bea3b430a468b
ze947cc1a592519054e62fd04779adc5ea1105c8d3c32fbaf557a8f9c07cb1f2238ef2aa7c2fc26
z4e2e008074a44be6ad58cc0f9d08288034eef30f67ab933b769cef8e36bc922386d6094f795e2d
ze7e9a8174b9f8cc0f7aaf851a066fffa03816f850606d212b09c2bd3f8b72db488e63c2b62d50a
zb15a8bf595a12b5228ce469d70c973c9208d7b64ac4793f7a5db274b8b36c2fdf92f5bbd54a405
za415a4dfadb488bbb617ebaa58d182c7a5d8d540b789318a5f3aae8c11b847ddae3115d946fa1f
z87b27df8ef942b5cd9e3d2f850980f79f2c6027eb4c66c42da8bb7da5ea2796cdb913b8f16e470
z815fc016a3d55627af31ed5fbee418f99a321ff972739b295872afc1f9604fa8286707f20b8edc
z0047473662a69cfb5169612d5fd459c61b604cbe4af4f3c9f70e4c0cc3e163db9d0c2887bb7978
z225cea20815adc057d2414a8aca4c72b618aa02ab3f9d3596606e9438a285a01de0cd3d90a59e0
z219e2ad835cfc5cbffd0642b0bc8e774e248c60429eb183f4f4dcedd3b0e286804fa4fcdf1310d
z8d89f0551fa60b05298486fe5cf7bb6fcd05d369b1c6f30de25bea46e4f4fe3f1d682185c7c807
z9f46c9f7b08f67a696a72bcc7a2cc11cc7abef883e5f468295f8c3ea6869a63d311eb3f24615c8
z3fe2f200bc57372a1491886ca8fe5b84d3cce8b30744f3bf695f2c446f764797183ff358514e18
zf0f2fae1da74ecdc26dca7e65646d9009f8c2d2eb89823a2e8acc7e41f9b10f91181093939532b
z3ba3edc0176635d516af2ad8c3699263daccea9d3fd38116fb446fb131b2feb8dac4b016dcdc50
z114cac6ec5fb35d47f0d5d439a9e83484df1a22d2d31d4904aa728a100ad0ed1730f47e1a8ea44
z1930cac4ef90b2f58e489891bae381390e88781b29a8797bd4a38e9efde235ee06dbbb7afcb1e8
z86014cf99c71180c86d8efee060ef35d841ebb98070df18e6341a6796653ef11143fa79d95f3cc
z0c448865289c4e7ff1e534badb2adbb2c59cda34e071977e38b06da584986cf825f8b5397edc58
z95766f5de7b0231ec494aa7ea881e0a1b0125ac9410feb664d31b0119ef71d41caca43803fbdbd
z0a0d1ba42500e768e8ee1b9ca3b4f79b9bab3e5a4f8ce6d984d1eff2d2ca193e088d0e3bf7ffec
z2ac6957221e04f41d795047e81c9822cc6a5e8f121c9d4e65c76a0df570ee3d41815738f1e2350
zec0be07f325f43aeaaee69910d68a17285f51d0498864ae980a070dbf2b43f41ee81458671c58a
zd52f6bb3cfc29f3caa51f76bf9138d17a1d191a059ad095e89804ffb9609712e759d2542b66821
z9fc0cc9a8e5a090509e4ab670e150b89244c8a5df39198386067a1a58493fe1f210b220136c4c8
z667eb6006422976cd41282bc76d3e0b19aaa57e650be118ee987c9e6ac65de498a9b53be492cb2
z5c7a750b9f1c7b4d66e404d9bcc6a2e396e2653f15c0012f71fff84a981d92fc44ba56b4447a3f
z478ed600ddaba13fb0b96421f45792236f224d067d3374381a6d8676e9b64304675f3c308338f2
zc52b0ba101828c294f8b31539e483f9611f026fa304b81ee51ee75b02814dbbfa1c7b9cc64e94a
zc81cd5ef1a6e399a5d3382c167c97c66e810284dce1373b766c1db477ceeec8d7cd7374b860c71
z3d3f3ff897820c359770882768b38f2fe7ecd33e7d0965f0dce7fedd8ce1b245e0c06fdf665bcd
z25de2498de2f5c1f805b18c81a61a584763b560dd1c422f68381c7c8d12a83bc1e55eaef38abcd
za8d183a5b661b6c788108e4ba808c49f2e4a963d8edeb2535da6cc4be698acdfa83784b3c6991f
z7af4ae4ebbee74c416244e8a84811d66357980d5e83a45a715f4a3b5f23a316024ec6a8562c19a
z4ee83b345138fb0685c65765e2058a2836fd6f6f0efd696181ea9fe46d2d863dcab95be8292587
z93e42edb8b539fbf2ceeb70ecafc768e31addd9eb5189e23b7ce14700dbfacb437e18cfce43607
z7f6bdb77531c5b717a9ca5da1fe002a4f78164ba85347a02f97408a42eceada56343d9e04108f2
zc0e59e31d3ee0c0b74ebdeef3c7490e6b6211b9e2d3ada4e113c771905516ccaf3c6edaf4353fa
z915771bcdce81d7a01ae539d3e5dd510c74c0c190b8bfcaad0a2baed280b95434a39cc3453dfa4
zb8494e7d9cb768950c7a5b3df06cbcfdeca7bbfdefdd4022b79e6543a6a692b17a4d4fa0391d40
z37e0096435c7cb30994546f8b54486336406f04b54c2b4d2ba97dd5e0e772c648f1cdf1d81fbba
z6120804d8fafd51a32585088212ef2001f00aeec3d3fe2ba01b87842b95371d51f06039696be98
z03b6ff3b5581f30d10b79ce8fa64b0b53de6174aae92570d08a49f2cc321d38eb609804cf1a9b0
zb67c71db1e8cc71f10f02ee5d6b582eedbc36b39160ff67e7300b4869ff2351b19b3b3f5260ca5
zf091f7c0ba4ca150e4d6a2dd262fa8c8d89629cac68b04d90a81c4535910b8beaa492001c468d5
z0bca5f5a435b9f24d61efe8f3efcc12db19e4f571b29ae65653655584448cadbff7089fe4bed60
z0a9ddf777f73442fb45a148e312bc344c483f2a695f92fd4f48f8841efa526f73bd7239dba2af0
z919e5063b5fa30b6f26872dc01c35893968ec8a264f8c9dab97019116e936a695ff916ccaecb2f
ze632a274e1f51f94b8e1ec24dcc5e5ea8eda9050f1496f4a8f4ce77e9629cd243f20934570dabd
z01dd9319b3661ba4c81a6be36f5a9f8c86f59fb662c257eee36bfcb0bf102b180dbb7fea1fbbc0
z0482b6232fb7162945a55917015c17697efc48be92595341b4ccef843cbe4d6898a2ff8b1ab232
z1c0abd024ef10563fe7d0b6ed84617c5e189c08af84c27872975eb17cb269ec614f4f51603e2a4
z9f52ed6f8fe13fd9c4ed684002b565b4f6dbf6662f685147d515790693a1db4cf4efc818aa8e52
z4b72fc90172fdb884669f56c82ccc01bad65dfb31811aecd9774967b5552b9ecf2ba6a7739d021
z806a050dd4b1761996a8827f96b317001cf8383c628386524fe475c344a99031a5ab8a7672cbf3
zb35ad4f47bec1e3ac636b4dc377ca9e2611cbbfabd621cc1de14ea54c8ce24a71c68b25f1eb10b
z9017467eeaa7e91389c540c5bfff610f0c1d98e483cda8510380269be6ff92a03a0e627734432a
z0b8ea630385a01871c8467dc67351a80f1a2a8a70f8e7c1f50d140deb5b835460899353afa7521
z0c836c29c910691d6978393e94690988daf6be15be94d5f1224151efda057384d0c80142fea404
z87d8b35f5a9966ab80069f86034e9f42d4ad8e315f9461bee92b444710981b177bd3fce63574b8
z9a8b484f3ce4f3f765f6c52b5af6d231587ed70269d4bd9e658337cc757dea160e2eef8b0f6735
z5ce77ba589ffcd589fbd4ff669d431c5150720c4e677c32be089a8854bc3b5e1f67090bfdf49ae
z76857288f2d2eb3e34b1831271421cb1ce948f3aad109f4258c61e00591ef9c327ff960395f166
zfc80837304b549572ca27108df853e8ddb69bd92575a860328773433f38e1d267b0c4ce84406b5
zfdb052fce6881ffbe56c39c66700116431c78d085d9be1cf242714def997f9e1bed77430f9e811
z9206ef05a24a8d19fde6490acb3b1b6fa3d80ff4b1d7cb08efaab8396c03453c56dc6be0ac5568
z6e20cac1b0ea5be7adf6fa4b03808fdd889f7f20db5d47fed88c9ca1f756a8a9cb72608cbe7efc
z25efffb11c0039bbc43ce14eb84365f47d49e3f132677f7c4fbc30afea6f810bdf2886839ca4e9
z82c4487a1015b30212a7921098e18a94a01912cfa5280aaf6fae52af5189d0f3f7bd0872fb6d29
z27b60341a9d58eaf90ef00c3c9fba1817998ac650ba122438a97a941fb75eacb0d44b37360deec
z3c7e6df1121a6502ae63d0edab4a95dc6c225ec074f18d8db84bc6cd530c7c493fd48bb1542c54
z1808d5ca825d116603f28a6fde3f45b316fc0224a60a3a09b48834de9a4417b17e861e5ddf5fc2
z77eb20bde1731c6340d695cb7522cc20574310ec14f45798e440ba77f02e9e342aca8875fe3d7e
z28ba4a763c8f70c637d1fba3ab7f4732668c72f14b24c0e4d2e8c3f658cdece54272fa9f5991d4
zfe8b4ebb334187aae2fe9e083ffe5b6900a9aab96f25fb31977a910719f092e3b9b9be676b1111
z574ab96bcfdbb7a211af8f11359ae0aa0c481e1085eaf2c8bea125d38e6c8dec5be12dd9581a04
zedf3103e76d728980aaaa106504806a3252041243905f8c137fe3d5484d7a41e645533f57ab32d
zf26ea01162d524a8b016c69a50a42533db06a4a5f91c520d28dc58e357ebfddf1458836048e1e0
zdf15af755844653a4fb609f558eab44bb69776995f65f23d0fab4a5a67071cd661f27ebf58c7ae
z116cb6ede9d308334bf5e62c63e06542dba921c476afeceb7f2410e60ac20e88ebcf3bc4952e8d
z6e8ad185eda9b962c9644425c4ab10eae3ffd0c8e9775d740462579c9735945eabc7f552de1b32
zfa5a15457e76a0af3a61f5d6197acd5a3aeef51009c94d633f50c15abcaac8d190b36173966e30
z07301742648678f44167925a9b1678857ca18f43ee960a8656d03e5ac8a460d5600133fc61d6ea
z099dbc025078034e8be4589c5c21a84cf66220a03db15daf97778fda090612e0fc70c08c082148
ze18a5e47c06515aa04ec3ed4d2bb7f1fd82f807ab606833c927baedb5311a6e4ba11b0cc1d1007
ze526c694a99fa005aec1576a7264a6a9342b7d61049716ee2c8cd17676b1633f9c79f0d07e757e
z9a5e0c8bc77e304e6c5fed160cbe751cbb417767df90ff0bae7df4a67165d0f45404b94f7ef243
z1b224164c6fd9f63ae4b6c9d46e353bd3a89dbe70167b050c20475ea23fc6ddf8c8fd96bd1d077
zbc7666b9a45c7489a43d26517a1791050d1a09a9b220d61bc09b4165ed1edbaba6c96bb65fe33a
z8ef59a123d99c3c3ab878a5bbe05bc33f89e45564408f216800be3f81a4200760e7206ad59d9e6
zc77fb08ba7e3c10138b8589f71451d5189f72ac02e85876e4a48fa2ecfaec93ea5325486579bcd
zc41423f58f9e925da8ffef2c032fe2fc75d24c7e16ad65220722e35c49889784d27e6b214601bd
z65aacc4971d108043002f6c66bf24de9e3f2a8fd94662c2c5cda275bf3b8bcd2193156240198e4
z7d76af6b003b2af865d26b94d2580aea13642dd6d965b69dab5d8e591e3e5f9524441c935d589b
z37a59d71c7deb00dc550bfc95a6903491da0b55ef35f4827ae2d4b43a5a8c278350ed4b00aefc8
z1d7cef55f317763b7be191cdba8ee2e08126703b7ece209716d5c5c081e2e11e2eec205516688c
z50f4f0ede074ced9f58f3256446f58f2987705b56148c78f5293dda25686b3a9eb520094b1d4cf
z61835a40ddee052ef17d89a0b46c998585a7d4c4c2f2b35ea98d699c4c285dc076a7398768fb91
z71a8f6512a32a23b584d504e861bd77b6779d52291e8af4c5866caa2eaa9ad1b6a283b2b351e2a
zd7764cd38d1e50afd500216fe55513fe9f72f449e4ca549e5679365ad0d3aff043de43a1c2a849
zfe3aadae511242aabedc9524674e6e2228d0a648410496eddd14867437c2d3281d05ed25d344f4
zf2a55d512649a4856f0012ce82ef21bb474e1f42ed72086486b45047e7acef90eb7c5e37193fdc
z8285a02a445b890e28b7a3fcddd7bc7cb5bbf33c119abe21da40e17b13c6d1b12d1688be653c6d
z48bd9dc8ae6ab179ef4ad188d58a0a360d46d1bf2e5f7b5b27a019b2c43206497dc144488c7fc3
z0eb494dd174c276096e045fa1dbaf2a97a88c0ddcabcd33736632690adb63674cc0a3d535a8a92
z4ef889ee3514f98c0b64f68ec80dd3f66d9764fb572ece05dfc92be6b2c2d25deb25c8e8e827a6
zd1ab05464bb02cf3df45eb153f1b54b00f8109c7b96d9329a9b6551e6c3b507179e06d7f955a79
z4d11b5ab2ea659af7c296eb332d501a03bd871c8f5c1c943ba9df53cb49f5b1283a91f8712a2d5
z0c2f058bf65512f8a989fb858706c0a77c494ca0f81ab639b6995b53d4b1cc4686c9ead8061116
z569e2319a6783af888384de912a4b2ae558ab7b771a6747e59deb01ca683c870d325bb840c24de
zdda663125fbc181c15a6b6363a362344a22837d12be773aa69bc9354d97e75548f91fd8faa5fdc
z0195ff12919e6ee3c0f945c674010c1919e901f3e165699582b74aecb11a0e2a71a94075fa5116
z67d39e4c655315c5deb250b28b3fe88d6a441aff3ddc40f86d43253ef5d1072151a8b99de2d2e7
za92ea9b32cb1c81c9c06a70cb493fe3169f2ad130171f88f506dfe50d610c4b964378086324c89
z8ab7374f4b5dc5f406aff998fdf83e768505e887760735071a8cf6054b4a4a219f83e6ac1d791e
z3e60e24f4724d3f01584a420e26ad565f30b1ec46d774e581b89e08855974abeaeb60c376d6206
za35300607239c2bfc170cf13c535e7ffde3028206f1a4c90a0b391490deb6b8d3df598e8cd89e4
z291a627853230474ef63643913bc694e43039a5112254e916a9c10412e7449c5b8072d63039340
z811336b6883ad5f71370aa6baa3c23be00f3f79ed7d43f586f68379f4a842366c6ede23119e84c
z8d53d4510c94ac20dd2f2adb94061d5c4b46bfbfb7b43612f8fe3dcf715589859a5c33e0396aad
z460d75e05c3ef16aaf7fdba6e2fc971ab16c0c1d58e5dc6875aad8e1e8641d3d830207af882bb7
z444b65a7e3ac49e11af341766e33994397908d61ce722f1b00d7dadd1e8c64e70bbcd3d3e48f7b
z55a6633394039a4b6a18a1f029cc78872872cda9590f77102e218b0e0ef4f6aded81ac7c0091ef
z3bf066dd6f5f3d4f696737095303053f757030b87aab1843a05cdf9aabe3bd55145c2c30ad3e58
z403d976476cb837010f3daf09f99570902df87286b8018485b0614ad68f477915618ecdd50af98
zb674099c6b81667eb734fb095ae1acaa19f7423c889d8a58acb0952dc2f62ea6cd6cb32dcd8ec6
z9f12fab7db1726781e3a83bf1c80ff6ab7e3d9df273487cbb997ddea9f5bc84b4c3d05d096b5ed
z691a871280cea7cab8c636979bebb4ae9a9d4ab31051f5627dba9a4980ea19166d90cdd2b6688a
z7ed60cac1602ea00a5391621240f51cba7c9d51e76c6e7cf6c8de8911080b5225923747a6eadfd
zf7988deeb57f021136a15bb9269cbf9174eaa6fd2aa70888e76964cadcce451c2b443b4e5167fa
z3abdef37af9973f5066665afcc497747d38971d6b7c85a0b0006b8c75edfc0c3ba5bfb83f890f8
z930d29434c809207f51b6ae27653f036554d201df8ac12b670ce7f0209ca13a1820758c6e9522f
zc46521e8236df3cbce3323aedbd43a1908a371ec84674e5427d112ba19f06d1f59235edae150e0
zcb9df3994ee9ba78e6c1161302fa2e752472179b3d36ad233bd1cb3bdb4d2697d9c4e939ecf192
z909e0117dbb1d9c6c5577264e958fa62b09b9bf907c16129b8327e6e4c6d103656d90a04ec3ee7
z342f5203684e4385e352b1e31b4feedf8bca0464ddad7e9a6b6c314ce1e93e2e86163fbc7827a6
z02518606cf3419f9e0c5abacd6b481f3fe14ba607aa232d16adc87396d26c533bf8771ce666f1f
z5a32110e72250b14d28383c3b14395aca86ba6e46ad958a3bf74c0871fd9eb98b276b90627589e
z043db8d673c54e777d8ed20725c95e110b17f07114c478d2c22d786e14cd258f377df86e50a1be
z54e910fd47525906015da7b08915d563cd6259b544d09dee3af13be49f1b4063e880fc70ceae7e
za9c4b205f9991a148db1399b99d0f6ede0d63bb0846409d9e893f3af9f59071012ee38e44a3bf6
zbfb1adb09862a93a781da8e9d4b098d75c4ee6b08e75f09dabd9349eaed952c34267b5bd624793
z820a1158a68dfd2f634f6ba068e5f5e9f7b224a6b30aa487911021f986eae3d7c5cd7cd2729c1f
z9e9c9ea440f188db3c408da982c859caff76b8d4530215b8e1fe6ba5c661922ca03bd07b14a602
z2f22774bf6320598484ff6ded2fbc5e382de3ba4c2e104c1e68c97f16e58d2bd7aa2fc2e6b0af6
z9bd2899123297cd88a17835e2cd5db83156966e3e5a54fb9d0fcdf559c09d2dc380cfee2468bd5
ze7d13d10f176e36e18d3d014ac142ab07969a075d30b24a4d9839164003b99e0e51aa3495824a1
z21aaf8afc668f2b6df03036b4d19524c0bd397d054ea14ee6f0392ae2a66461929b79aea8a6346
zd14e7e5b06439defc3e8d2d2b2d3e8a95b710575fdce3ff8a37c0d1c5f72515f00b88a7f1c00de
z3f051e34d79cbdba62aa6bd2d68cd004f3e040958e10af97fcedcee496cb5c944cf9444e7eb642
zf7f9543588ad3664d1f141e3c817e923660ae5637153337fb4ff10ff54a9f0de366c8fa639b9b7
zd9ae9ca0f0f9c835b1ff2e09c440f9e2e26feae80504625f8227c2e2c244fcd9d43f6efab84fea
z283f0aef6e94ea819820da5c3e9d65e2e03556738f7a08a7d031550ca3d97a6e0a22bb0aea5196
za685ab967fe2cb91888041bc1dd2afc6e7667c55cc669961d23978935106b3d0a7a75256e3d88f
z161cf75217cc08d2383165a4ad8d0597364c9416fb27cc3288c64908393691b88c533a1043b6e3
zf17f6e7205a0a8c13ca4f7534801d2260b75840ae6f26ef675f999a61e0cd24df6023d94cc45ef
z24a89ae2e2020d37f69455d33885567f054197b3347f69b7718bb35bbf08784a9c8d1a2602a86e
z6f349185f35da65547e1711dbe501e19cff02c25942423514a0443d15e84c72d7626e64967e904
zf4f68c6e3f987c6d1bd2baa7bf2979824f38a6ac5f1caa247f57196001eed6f81ab2b754521054
z905e87eb2c291c69571bf0751219fa2c742c69e66c5692d9562fd900363cf669cc5c37267f7460
zd941e3af6544d62214b46e5daa8e1c64e800b27016d607ee2227be99902e4fdc216ce05fa619bf
zc2045b9f704327d8bbe0be95ec58762daa7473dd126a2a079a078588c6d65ce5ec1c67b9c65c12
zc13b54affb0e73523a51e1949c73ddcd6f2845191ef784b35ab208cd288f003318c6eaf628ef0a
zd86e555f1217a957c9f31df1cb8cad4c2d5363577af8fe26ce557686814c94727ad1d21fb77e9f
z267d04f68b31cd9586df79b5e387d837e8bbeb8d3b3c86c9083499fad775b6c086d3f341a403b6
zfba84436086e7376f49d1e51de9cc105af85eb984d3758b5bbd8c3293b1cb0c8e157445ddef33d
z4f2bd8e27e21ebbdda4e7fb8674acf1d147ba864b149d0f30a389a8ca517d88076a7f2ded61b03
z124fa793e92c8c1209619234308f7ded427540b5e94fab4ef638a5452a5241bde3a96c0da89592
z30ac2d70cedfefca6cde4ad6ccf50d0e059835d4cde80e93dbcef3c2e2e4ad67a2ead90b3ac603
zcb53baefff30bab12b5f19b608d5e4bf438a3c574a16d42229032757c4d49d5dadcbf417ae2aee
z4a63911edac185d810aa74a1514ea7b7034d0ba232bc6d750cc00e94f7910fbf5e3393a5b31488
z91b8279ac4a756070e4856eaf31ce3e5c591a297ca0ca72bef15ac90de8c92a0ba6d3cf7eafa05
z55e4807ef979e9a1b2cc7fe485fb6b890e09d68d3cb658aaf77b1a9241535806b1a59d3b2405a7
ze96629f4cab264410b4c4d1de913ef43239afa6f1c303d0143c56f123ac3c9e60beac7a19077a8
zfb83f0eee9464b2519df90517aa3db4605bd899675136f0159254d8c34a7415cf440f3db78a5eb
zfd13a3f518607315d438008ee9fba866a97a3fb150eb1008c3d46d998c95ada24e0464a81f0f56
zbbc5e158d234622335360abc0074a79acea8e6ab725b874e296c718b038ddbde56d7090cd2a22b
z0c9c225c440f103ef926145bd2d881b922a6636b7d3546c69d38150dc47446ab9e997483ecbe92
z7380954c9a9569a953faedae877dc88f6590d8506c6e7a6e490f6e07b7551058a3758751b71995
z467568a7efbc937305aae8ce37a7bf6f770b55a3bbd4f22080570714b61785ad58dfc384117018
z8134ec7fb269d65692abea87b408fff55a71dcf414718a867df6a6915bf94bc58e49b189e2cd0c
z867910f9720fe93868336b5b8a64e0bc822b3ae5b9ddb323f51e8de608d4b522e56ca2220446d4
zc87161af5900e5fe3fc7c679b236b0f83f2f243a5ec9c46944827c788e0f095a3ae6267e89fc43
zd8799fc2464ae5927dd5b6153b039af38b659ed1a18faaf75da1a4aaf00ba776e099065a08bf05
zcf5f37860e085016ec239f1c0246d5a1250ec17c42e71b42f551f5dc8db3efd197f46f7881cd00
z69108297a21b0f06dda7b16d2c08863c19bddcec6cac63e10772a7bc690384804cb3d75f03bac4
z44e639c0e0b3d70b3f9412b2ca00c1ec80b2061978b58326cfd2b914325fc60846f820fa9646b8
z1079ce0638ea7d7b32ccdf81dbe722fdecd975f8e5124e27c03ebf50ea615f70b0a4e804adb717
z29848bc1e45180fc83fa68617bd37bf8526b03da13bede69eb4c8e0fbbe4f72d73fe9f807c1b23
z25393e7eef308750ae9b489a8db744d518d37dcd52f7d9e97f13d89035cedcdea05ccb4ede4873
zd631dd17cc2e8bc6578e65f00ee9843c05a317d0a04b51efa57db9a8dc1ba8c3746fd22d90a20f
z196bbabcac53081848d211b56309c49670d78b8d81da936cb65402b5d3d669ddaa149d6d019b23
z25b48863b1c5b1e8ba0af6d991ad00801ab33db195a89b824c8f51e59b659902575c5aaab693eb
z093d37237a1e60b297194e0cd7285615b561cc729442584576a50b9f7d5f35f68d3c8897759890
zea96039cc2b7a5e53db286fd406d151c584050e340e95bbc21600eccd2c9612408cb4a64907619
zbc5b089ac87e7f1186f28f6679751fcf3535e78f6cbbcaf9ed9d441b35e1ce08c64d90152c03c9
z26d30a7c2cfdf91f25f795d554c747aac668cefe08135825808f36cbd4d8ccaef51564d36bdaaf
z8559e07acd9d3a83c8f20bd7a2cadf55d1ab9c3250508ae2fe5afc26f287b76bb708dedc98db7b
z249618cb7574a1088ab30de87cd9f8fd26dfe106bbf8ad728a295d6d9eec744c93e79353769176
z40a28b21ffac1c3e48b786e26c8cc47f9fe5a3aef37245295352c53fa5d1086a0e224b12c7d58a
z5cefd16e194b5086dbf31c5b729c358e882be6c1fda25a84bc583148da06137b5d561fe1ef2ceb
z2d69b6617b03b0b6ae181056ead5059322700c074997665f9b32c31d9413e9c1372d31554f5149
z487ea831995fde7d602678cb65bde6a8aad2ce11a1cab42bf953f35cba12a0c903e68d98a0f538
z46a7e60281afc4b4e0bab4f8cd2beea892c6e302a63c156a1c0c60d64755ca52da542458db03b2
zb7316470680847e06c24a350ead51192967691966d8b0d21e29c532076455d6f36147696ec6fd5
zc1d32b22100a022aaa0f40764893350ffeba9a97f237a12bf475bbe13e928d9299e71c04ec0ba4
z8674f7c785a13f9aa4f61fe9ea2c7920153e009d94e9fc20a091f09aacfd43aa76c6e64995f439
z15b87a7167dfc3c3f0ec28a918070488d612a93f0b9570ee93822d03a07fca3cd6afb75e462cae
z666dc2507c56b1e382703a4e0696bf6a871f972fed65dad2caf8d46fd7897fa101397783c62de6
z2936269c7d7020bf4a5f0fec03f23a020244814ab5b06fa80369a30508d958aa615c31275ceba6
z5cdf75ff633a1123ca59206b62c0326aec4b7a497567a60d6e79931dfd31a0028c5f37df0ce8be
z292b19e43f7ded92f58f67773cfcd3f5b76846dafa50e1d467f2967bc5d7f7af13b80e09573f6b
zf03f06b2c726543cd5efe97adf3fd980aab54ea4a6e23eab3ea19d744d535980c248b397bb6eda
z58e553cd67509a39bac17fe311dca34538916451adbd59b6837baafe2e64c8a2a7ef149d71c960
zb60856aff05f04502a41baffb05edd10a95ce3f7a1dff1184361c00d58b8856754f42c1fa50167
z2fb8194b2f3e8c9c1fe07ffccb1dc0d765f703f44ed72387bf5b21a65197c50e640b9417d60478
z07809a2f1f9c239338cefa564fbf33a742b3eaee2d57872ff29c323190cd50433cce885f72fb12
ze15bc7feb6829c568d192269674aa1b22c5a7689ee21decf3bf65e42097e5204fa538317f9f006
zd332b616efb1cd4314cde4fee0c9c6cdb1197789a5fafd8754dd8dfd685f2dfe96d567a8b14d81
z0d46cba5a51e804ed8e9632a9c88e3574514e50045482679ab836eea7c863988b1f13df633438d
za04e9d14475a50a3c041d43698df94f470cf1a5e332c951d49389d2efdc1f248920037187c166c
z44a211645917279e6bac5f2329bd84e50ace372c183dac64776a9e8f4f76fe517497e9814fcaee
zdf125774eeef5615776743cbeb7dcf9b817c343305e537850f62bbc05db7acef7c75440e4ead9f
z687d377f0e187023e197a3aaf9745934e34ffc5e8dc7941a90dfad17af23939bdbdd351b6b985a
zd89d6852e98181712bbdda9f0ac75e352eb26b47be3466e68df92ce3b0031d21147848e9a66a48
z1b1f0976bb887ccb65b3e5a016bf70d33e41c6532651af1c5e67a0545dd981223321c4b8e016ff
z51043505bf4c604604733f797fd88b6f0b0ec13192d65b6cb0ed9225f773eb6bb9c59a2a8dac70
za6b4f5e7228e5251551937ea050555dd744e27da4f95b3089f57c638eab1a02e4f8741d7453d20
zf978be9916e42df8829ec2ed3cdbcaa132db9204db7cc68e971bbbbada40f93f40907ae684ce16
z6232d532aa5f1ffa03057181e6e113c6c56a4e325683ce70c84910e183f1188fbd714860759fdd
z1ac41b66bb7b24f43d11923fca811cbde4966ad905d21f527637fa24924eb04351b7c3a5b32a98
zf36572dd4e559a58584344d32d027bf015697e7ebe86f10b14a73e6a02ee8cf2a6f8fcafbaa299
z965ba63999376c5b7182217d2b5bcffeb935549c49fdc7a5f8add82153fdbb186984a624487125
zf75d26de377d033eb97ef2a1d886c57ca038d57654db299ea49bf01a0cbc8d58221d8c96cfa4fd
z13dc585b3f2cfd37e6fc19e926696ec411e4925ea417ac8122c1c082d63fa194b1ce986388d28c
za8f09e0548506ea0719beb98e105579e15f07adf85ee3b2fe8d1e517bc3de8fd0810fb9a55f840
z80466570a6a1255e8d7ad4549dc17c70174f2523b2ce74a4260ae43dd94755f867887f8ac33933
z0f738993f20311dc32491d21a4a3350222d3e8428f9d640e0eb336d4c17857d449cda9553dd214
ze6a6c61e8bff39b54c53e1403eaf5c4dab6d280e10489fe425352e60669030ed2dd2f06c06dd8b
zb62c088d2ab069d1e37e14f06709647788de36e9b8b40e0654b56bc0a2229557e6ccae1f722f17
za3ce9c10adcbd47f5d265b0f263c793e370df68701944eddae33da4c0ff1d07d5baf9f64fe7c0d
ze85cba8e1aa75d2382dcff3f5daeb63f29e83f10e6beb1b2ad381474ad72a68b83301089fc4492
z656e5ac009ccb78b520f3bc45f2a62844e1c92b9086faa03dcebba06dd731836fc2d7a5fb298b8
z48f338120178455818ee1e350f70608dc77bd3217a2f2cf7e820b50dd61092fdba51281e9919a5
z7f69ae8adead351a46e814bf0e9110e6f69a06970120081bc5766052f8922aa4c2b6343c3742c7
z72f62ad632f35ef79ce15a3c0adf8ebd85bba34ba3b5bed57e7005a1cb552cd4645f284657b6bd
z7e500f8c9ebcdbfbfc127a702e9c48863c5c137a60f78b533748ca52180ecae4a7f1229d443ef3
zb05f693510a0a0cbaed218c21273c551e2bbb1b7f7a4e5fe3a5d18f979ee4c0d9a6729c1fab60c
zbff776491f639466b9d014fb91455ab38f33f04985e1023e711f7e60c4a80931bf7381ee374182
zc1b9f02ff699927c0207b69a4a692602f9fdd122040e52b7eb3c2277d96d2017050e6b9ddd3e74
z570b0463123851248d9544f0ff52af47d086e941a6c31f52b826257019c98e4874f0e54d76b003
z1a24dad8b4da1e07bbb3ec4534041469c22316bab9e8d22751e9c9866b2c3d3687b1b2e9221a50
zebd69b7bc7cfa43cc6fcd70bd30130b3e0af1be8b46e3d07370081e35cdf05241bcc1f16ef7a78
z543f43bea24e28b5ef5946f6daf8cc84aa538b78f68614b3d639c528c9239d0f6522ef63564e3b
zd791ec753e685bd4e7d825ce1e2f05c532f069cf6a3dd8c4ca44baa80fc5c803be3aee34df5849
z925c7d01c7f194e1b99251301e082962088eb400b09d730f7c915d40cbb89c502d845f03c62c94
z96c50b8624820a10066a515263398a42fac104125a62029872113240947a3afebfe8b2a3d821f3
z3fd802c872a940b92c74ed8dd03c4c1c91173f793fed8c55bb94cdd3130803b00453628e4455c3
z326c10668d5cba7ac82df7aef52edab6e592b334fe90ec0a4997f9f0518875780b2785a8a2fefb
ze6e1dc76b7782dcb5315c1120367b2bd7e5302c1a4fa0d787af7598303989fbd9544396ccad0c6
z1df846e852eb88612f44aa19f35ad7970c3b42af8d7e370d6aac699a82732a616fa5d75e668030
z0ae673b8620d9aaef31da81d6823f4980078432114c964268bd2f8bab1d5d9fa5cd617f3d979b9
z8f61fcfacaa2428563cccc655bf53efb893f746c82969862d4c441060525f43bd1cb7a0e0610d5
zc9f73ea8e6ed17e80c27702ecc8b1877503e8bf619efa9860382fe10a198832b0f52033d65907a
z258a4a497dbc4efb7b683959d2dd3cc09e05cc8d24066cc9f0281b23b74a5ccb557d3fe221c0b6
z713a8e0dffd17e8aef0ae09337af92b600d40cd8cc7d723c198a6d22b9c7abf48d5d28ff9c9316
z3e2557ec47da68d2de8a15defa709ac1f47315ddde169e36ef4a5b95591c087be684a9d8d84cf0
z7258ebbb9079b3a324a817c5fe3295bb90f981dad02e5e71c1e66881ab9971283b830614bebb11
z52473b8122561da11183cf65e003ff04701e181b58d2bba58c9767660e12b0af6ac625e17d2697
z90fa9bf2fcd61506e0dedad22dd17f20e2f0c34cceaa706a7a12e549759d5e2c6fde1d7c221392
z15636975a00ede734d62f254678b4d03317a1a5b3c635e5f2b635d888720db6285f45675460e47
z3167d35028de98cc7309659801fe1bf6c8396e5369f1f987d0658505402487d7550b5f4d2efcfe
zff760a3ffa8825f5ba55de2767104653980db93df142db26e62003248074609322ca96bba4aa32
za2efdadc3288ff1dd304a156c5f3b15ecfd064fb64e4f807dd625cd586ce97e1cb5848d7214717
zfa601adccb7592bb0d175c9f5d0fff14ad374a91e8f81e02317c523e002bd33dc752757cac3226
z9dff72687dea615f33a87afb36c7d087a7802b98260630bab5d1407a4779f9d1d9c0d957a6bfd4
zcc7bb923f7ea965d0228a6ab85e62cee06e427e516a7f3eeca650331e7eb5be3d07bd039939f18
z4793f11e75775394b58208385768bc78e4efd34abf4a7c7c9cbcacafc92257aa1f4ee542ce3db6
zb3f17c27eaf0e4c8fc964d6555899aa87e7b317fcf5bc488c1b96cec3c64b8ddb6abaa20940d9f
z2b1cb10265d3e17ca5645d2b9b0016956532379fb8aa25ad019719bd930fad2064de8ac09809fc
zc2e95d6841619e37cef8fc0b547eb71aa6f7452e1b8a2e21a3631d01fad6fce23595b32e8737b7
zff3b5e54e775bb6e36625814522cb3e05c7ce2e86685d987657dcfc386bfdffa276b0489520eb3
z91433af26e9d0bda81a2daadb42cf56e70e93d7eaa32349a9b3ca92d32f7891899d268e626cfef
z3cd28e6d21ee6ba61fb816c6a623d4c40cb40a64ebff4f239eded8c5472ebcddcadfbc99cb358f
z697cc80d11697c7917699784ff2ee30ca160d8506c21b2059c778c089903c6e5634882130b6790
za0592efc226885e9435577402728b92aac4e6000608ffd4c5a4cf3900a503a622fc8cf12e4d566
z3be0ea8bfe810c236a1a85592fc4b20e3aad40108a2377c5bc24ba2deaf49f374ee7a59abf2e23
z1b50dae0f7e70da25246c0af4d2b09c81ad7314fe7596203901ba8353d42d456907bf09f66edda
z941f5487364aa2673ee899b4246c89bb2c40a560228e319df881f71f6ecf913cdf82038c727d48
z1c9a1536ab5c382993001c4fb6145d5552c4b1ea1da3dc5a6f64fd112d7f37b12d78448a969a55
zd495cede053c94f47d6986f1f2d571bf12938312110dc6f858a4ac0dc4c722d97026ca4ef217e5
zc9f3d099c3460b8d748b0e202ae24f832cedee5025ca900b469d916f3fd0fc18b66656de86cf37
z73195d64d8f1a0c4d5b68afa34ee8bd427a3a5577b75c05f93722dba609552054911a8f5016c40
z7dbb275ae6dc5a98fd21a2b31733b9c679216a9368948cbeb5f2a010affe315a42443cf22ed9a9
z2576af2274688e02ff92f3c7de907372e1f0ee9f2f70385e0196a2b4c1b7c0ca2138f1f0459b17
z183bb4abeed9682b4b1332cc98f90c26dfeb0b893593531254ad482f0fc213ada0a9f5a4687df3
zce1254037f0d8f8585b16d3d456f23f750c9083148bd46348f8ca6ad5fa870fdd2c13bbe03d811
zb040b558ac130e37afaf3bc883709d5e80f343a47f308013d92e3decee5ddee53e7b4acbbaabf3
zc996905a2659a12ab46c8c3485535232ce34e009914dba2f20b9883ba705dbbc7e2e95c7013ac8
zd3ad997abfab02cc46f4022f4fc0e02a65af9147aa0ee089615042f11f067f9d2fd5dde64406d7
z936cb23a4a83d3d1536269d7e19f2554af223372b189c3c5d542f1f6e1383ce9ffba66ad25f441
ze69c5c81c6c8deee37d7d70a68f31ff5f189ef5614d7835255523fde420730001e151b73243663
z92bde20b81671e8961059264644afe0e1006e426f57bb5a74a6b23c4b20c07fecb31933bd1cf8d
z099d333dfeae68726a1787bbf7511c9aaa7ebdc82c468f7e69f9a24b626fa13ea46a6fa39a968b
z3a25a44abe9b030972af4bf213e802356bfb70330814afe1e3b90c2f08f3b426632c589352cabf
ze766ababb5f2999dadaae2a8280abb94636ec80f2803ceaaf8a38dfab7beb46de5e6cb8830d223
zda95fe94b6ef00cb0eb12c9b727332bd78bb08d7288ad08b92b7fe0c7e975f5a759c89c7a1c461
zff957e87071909400b21005b5c8ef3c043653a0f5107b89b263d2ec0153a902745e53be3236be8
z2e46f3ddec4bca69ffcde688262d49d904f5d05d9bcc68f0fed227a47fd4e407368609359ea1d4
z227613dcf4469461006490519a4bf9480709154a08e34a0d667425b62bcbf4c33912083b486d6c
zef04ea8d049adb2fd0f16effb0f22b23b684cfd3b513b3975ae76fce360ab3d23f6d2c01483cf1
z28293a75e0609410471a82baecd047c96cc05197b1534ff5b96f32c1cf4d836f41c13d265c7d78
z6247e4eb3af1968a5d83895463e10cb533df727c61c3cb7f4fd7bdc6271fb2e7d8274b7590be1e
z9c78ae7e281cc495a51345da711ebbc1511d5b958b79e1f03ef2f560f31a13ec02f3600cdcd980
z6fe69ae02d01d9b6bbb7f4dfd7a3cbda0738319830fcff96fd70aaecd6847b18ce90017b8f8067
zebf6deeb75cb9c15e09825c3193794e20be4d2041b8a6ae681e3fbe59c183d267c81dfbbe55993
z529b1965688d0affb38075572012491ffe62e1d9cd31e1e2e91bc54cb69251a93dbde0f60064d6
z28b0c4849b96ed9dd3c49ad3e598ac2b886048f650d92a19f101bc00f3d2aea07883bca8af1dd3
z14b191d364a00b635edbde518c542566cfe660580d6f99eccfbf646864117c05b82af3c5973bc7
z81717e8fd0579a29e6ae0be47bce542ef00d67f38d3bfa80cd788b5ab876568e4922966cd9c7ef
zf37a6375366a486d04ea139f9619b58e5f90bf320a06c8bb45aa203347a34249cef6bad7e9892c
zb8a0df99f31030ff576bcb6debcade5472a8455792ed86966464e8142f2e5e4d07301736c4d61a
z77299874a3d2017be51d8b9bd5d7692c09d8d085eeae48e400bd0c68596a6aea9baf71115880c6
zb349b646e8ce82dce51c54b73dae6896218ec26d03574c1f32a522cbd5a1062dc65dcccd504b10
z542e249735d13cdaa616ba229ad9ea8b5c487ee33606e593ef576051b79563faa102c2584b5758
z37b7029aa09ae4ecb797bff4983274befb9777d0b888b2829c25dd3a1c9981d44c21ef90142d6c
z8295a5e706b312d1828d97636c28198701816736d2516efa19958b27d2817c1072e315aef4bd24
zca8ce59c7d50a63879dace54656c2936332a25c8123e5c0cc2dff664163f4bc48e107dfa61dce1
zb55287219d562dc313fef3e7cc70fb62a687f1831fffe1e0c6d0ebab9e2312a547ab1af21032c0
z77b63f1b524584ee235d978ed104022ea020f694445b7e71d067c1f8eda9987d81febdf3be6294
z06619eb8a9c813eb02ca0fd9ff69579b57e9a157be6f23baf619a11a7c67325a1dae3b321ecc2f
z304772dae231dd1028985065e3b128bdf033fbfeb230b542f4383d9975aa0e66f0b01f1812c3cd
z102146aaa874b323acf9915e1db59a76be9ca24f1350789efe835fa44b6264b6ef87666cf8ae2c
z9d191688f6bdc913bfe029197a8cbfc7d8a4a7460d5ac086946d436e6ecf56994bf6eaac767829
z3ed4d689020104f68ebd2b7afeea5887fe6a47cf044d0e6f662ae6c729c5d3262981f1f362df22
z62db8904f48ce3bc7a127172436eb0fca42201f46843188e06e71a7fbcce13c5f4bce088bf3e3f
zacbde79af6026ba2073306b0c1672d12859cbf725e728a22ef26ff3a9a6cf620af228eeda507f0
z243de3204912cd5f1de81b6d41f1e8aee36d44604c6903018e3a9bf6507e52372795b87a78ffe2
z51c94ad66351b6ffe419c732b3e81d08dc166b5521bd7d7803d6bfbe94040822960934e56e1685
z101c876c61e5e23b8f44dea26b3dc2ec652b7eb11f5cad67b2117b6df40b033eec6a9302d435c5
z2c07c1b53daa8146351545f77e994644d4ff97d723ab8f656dbb120db712dad2a971ddfe28eb2b
z05c0b4425999ed7b4930535138cd829814e028560a3e5babcde91dff04c1b90cd8b3cfe79c9507
z59923819b0de0fbcc4b5a4e86faf71f6e7b0a5a3a384a08e8fea09e331c9096acb7318f63ce52b
z93ae8e9320e918d73f6106eb1bfb5f9757957b8e6aa3d9d88847c603b96f7319871b2a7938a87d
z8233f2c7ed078112456b93c2a7a4327db84aba45c8fe0af6152b23650707f9afef4beeb0067092
z9125f28071311e8b9d2a8535b951038cc6f3cc3439cbbe65fe1457f3be145b02f3f537c3a9b54f
z9fd21e6d284cc23311facee35b4e1ce4ff2c687891db6e52bc6a2f638ac62cb1315c6bacab1bef
z60708f0a742af6fb029a35050bde7d1d906626c5a983cd975c14fe5a35d6d586f9fa887521dcd9
z3f9eb509c5dc92938b94a978c40f5bc0a5b33ecc1be3413f0b27a1bdad4471f863e5601b3ce1f6
zac2598408e889091961a8a58debe3533e8ef04b87b80558a8b418e2de1cacd63906f5c3d6dba33
z7a3eb7d3c8734234bd90c283da63217ddf2dbc9d3ef3f9520e584380fe0f21d0192631764b2a0a
za0485b8bb5236ca273b31430eb2f07a24661d6bd75488da75504d0e70f40203a277ccd67d02ed0
zd01c026c6c9e3eb8a1f8982fc01e656aaefaf79f7aff565e42344d205b416f121cbf247d82a9b9
ze19cadaa93590328e8962668c1e273181e084ec75815acf23d53752a7deeb3a99306f76dd19cd4
z4b991d994d1a5dc5a212a56d539fed1680aa4ca7e80c0b9826c55b891f4a674a9454062095b4b5
z483135dd648a5f13cd1fa98b00fb275a21aa85e6674542c7de4d14146be2176f46ac95459cd6fa
zd86edf33a99036b1420ca6b1bdb2418e4f3391d5729546a66f3cf8f3a82ad7c26f7fa80d1b2427
zd3b7e941ab9b04940d4cc7b8a2a089f0003f6bd12c3e54ed9a37b5954324a6d38ee8597bf2b80f
za7dbb7a6c475a268e4e9b8f65864c036ced9812da57d4c0e18e47fccc8965ecc977ce809abd0ff
zb8ad76230d661091b3f926e4d590d05c46070b9320394868d9e8dfbd7477622280ee790d6e8bd5
zb3c4cac07245f71081b645129b25301b3ec869522ea1ace177037c6800bcdc5bfdf265c2bc61c4
zb9eafaaaf91cffdbc182d6ccad3474b0b5dec105b7707f8a78186fc45b7b4bf0631e3c6468effc
zef13649381eea10dc20cccc6e8048487725e32e829e4c22e462964bda79cd2109ed6049d450993
zea454f0211ae9ce7f205f76b917d61a233a1a7a5d4436ace6abc38b354508a034aed39238a4c78
z0ce250244eebf7f49b5ab711a533091420f0fec854b3a9eb3a8473384c31b7f0bf65d9a49e168d
z770b417ab70f21a68b8d32e73fce693cd087451f52fd76f374539ee0cb40163d44d7d0ca9f0d67
zc1dad1d8b41aa8cb353c12b45f8a6135eab3c2834d4153e1bf0c7e7a521f347d69c213945d2f14
z01a6f0b5d29d2444af1bd1db392751c142142d70d6cd8b6cd2c96b153404d339ae603eb8842ed1
za4ddefb7dfde131f1a0b8a2119bef9501520b6baf4cc94ec400f541a76cbd5eba18e3419ad9d64
zc68941f4d29bbea3d6c0aca2f008af2e08dd9a215579b59ce41eaa3c1b5f011b0f95c0b59caf2b
z753ebdee1071ab4a0a132615d9c70b446171fd3109d08bdb62633bc92a493a27947e39292ff896
z54887e164989dd337095230b7076138e7831d9eb5dd879290b1eac9c930aaf24e4c938cab85115
z8919a9855a5191604324f92a46f0b1bbb92ec5834f292eb40ec9c0f82d0a6c4403a196e5e77705
z0818e0e776abc9e22791e63f31e291f84adb5ab88c6b23fda5c879e65982fd92c0265be1226646
z48d073f78853c64a13c95675d189b5fb52ef2e66caa66280cc6dbcbbaf1ed31d11c5ff9b608ae7
z8d541d9f9ad44048227f07abd490a829390790b0c3d96f898ef6e3b60afb4fe47836b13dab52a3
z3edf4064b4f6cfbe024910fcd197b8e6fdade4a926c57b4d25fcf180d8cac6d82ab6ac8a28d70c
z01a2e3c71a46a538850c9bf1fc06401f354a41942b6957e1559de93628eb951a8f00bbcf0d50f0
z87aab586e4d5878743164232884c6d464523e82847eb64dc5b326728fc5affd6ba312a0ffbc1ac
z454f690c7b89e334d8eb35b1850325a1fdbdbe75f2717092b4151f8fce1cb3a37e5d0f7790dabf
z6fc9cf521a2f35fb04042905282c297e45a836f526af3a866a842e69cfa5e8f0f76c9981ba7d9b
zb8069611b98fa9f5cd25b82e32a80e2cfc3bc38042b64c3f46ec7642a190ce5c0e634cbabf6045
z9feee49e63f4dffd89e9366a32d7497621ba0dd9e9f5b4c03a16861fb0b89935ba33a48e457109
z2350b194ebeff6de9399201affafcb32823b10753d90ae6d472cde2ce1a082dc73ea10f7b5eea9
z90fd17d2ac4c210821ac67f772cebfccaff3dd79ced7da52376b619bd861c9868fea57afee1010
z209840f8a08381d3f3ab1bcbb660cff34adac4ce7c424bcb65e713a4f74f5a85ed03ab352725d8
z214b53ae3035ebfe1261f5c4e0ad3640a20d0d4ef3702a750bfa243a46ccb68b3eb2943ed1b705
z9df428696d88f6c583c4c3b752007443872630ace89ee2146b0acd00d13f1781826b4872b7fe11
z6221c980c81d88a356e0fb146eda29f644a83f969bc256372836685380bd93a8faa1be94915798
z54a8e7759fe2e315ace2144a216d0571d1b4fd64b099a654624be4f2b31a8c052b47ab8986b1fd
z297420864b2232102ccf0170d7b1690aece947a5af747fe7fc29b4eef6b39a27c7cd1ecefd54ce
zc48ff381809ea4ecfc3ff70e0e06e23ee2e3460d7ace040be545c000a8f343c4f6ee982d83d73d
zd9e5410eaf51e80a4ba6a1ca009b6dddf3551eeff0b69fc952dfb4876b45e891ef1f134861abce
zd77e4d330d3f39c0d193b03328f52024706304dcf39d64265e478130ce4685d08ddc1c790a9cca
z98aa187cd5f0272c8f9abc6b92dfbf35857d653d310346a92882c009c462518183b2b6828ae93f
z9320f54985639bd2725596e0ac78d2e211e628f7f46cb8e34abe8e0cf6a964eb2ba95b81811a7e
z0475124325049ee7f20a1734f7eeb019c6bb36479210ba4a4322aa5e3df83f5c466dc96d855bfd
z0374a6aae54f8f22a2d5c2d8c6e13a80e82297ad4bf35804419d5a20e26eaec3c0bcd40103a2a4
z91908831f3b4d636d2730270fac8696280fe514510d93e99215e4a47d736fad6b95437535affd1
z3f6dd4d9a4620671545a982bbf9f9948fbdc72e437380aa7c9e8f966de5e769f05545d3e3e5459
z230e3e367dd01f3d11f788aae93aed6b42bbaff8ca5017468ebc38ff2ea8227211439ff25058ee
zd73f32a810810e1c06209e49f8e0bc3334525b81fc3b0a3b17d47b2a0fa54883b23b13e8f5573b
zec4d08e8a2814b636eb175936fc1b22ef73d4e13c38faf43808bdae2faef4f61ca25b2c4f3a34f
z6ce05dc4ae32f239680032829f4b6aa06480e0cf00adb5110292662b43354fceef417b322a785b
z78b5e6a0fd10319293fe9828fd915166748d43ab20eef9bf5498f06dda6647fad22b12da07f040
z74d1802e2cfc4ca673d0b5ad0a0d0de9ce4c8dff7122e638948313ca9e7adf7d46888bdac20cd0
za8eb7021b8bf16d3a3825076c7949c4a9689451a26a6bab4d8c0819cdf8b7e93d857246f6785aa
zb0c14d533512d1d787e150b8615b8c8a39095d5729fe85645830851f832d6ffcd857c39658d9a3
ze5000e2f64c9d5e83a2cd0d83dcc53a3c3f03d7255c11ac5f2be6906afdc7e89d87aea53e6b945
z3499bdf32400627a877b024f557d3fd25b45fb856cd8e79f59aba063675b8b31870d445e096159
z26c3ef580b62b92d2910e20cf417da0961f38b983bed6969c32a8e21169e40913fa76a6754f77a
zdf50c0e2adac301627ed7944c42a4325fa98f5f62167c7cc750335db7eced8ee73cfe005affab3
z2dbc16acebb7ad866bdc463dc0584cee96e0f4cc3154f281f7b7caad57b9d5717899c29ca7cf40
z9b8923d804b23e69db56cb9fe4e5403208ab225802e4e63196203bfb99056b79dd58fa88f4870b
z53968ffad0bdecfb2a6911f14a57a2f1bbca22abc85c408f7da69d46a0c3806888b8eaa7b3f2b1
z08282fb4cf10836d76708db63926d10caeba83581045ee347f6ae8495525b14d35cdf93a1ab9bc
zf32b015ae03bdf847771b98ddaa5eb8368a54632082f85ce4c5d0291999274e4f9983bbb96e67b
z12d4bf184f9ae98df613a45e5ecdbaa98d2f385f954df357a691c7be5f3dd2f80509d79ea8c931
z87862a916111ab1a1fe8e4f9d51e54eb3772ab2eb8956043739e9436cc2b6355967271e7636749
z9643d9f6eae4e0c32b3039738bf8120a4e130d30737cd8361fd7f40cd7ebba367901c7d66df522
z7bde94f0a80eafa80272c44f8ddf4c45ac4be71139923a8319e343d0cef7cfe6a0c44721a2de14
z8a958807e7f9be0d4caf7809dc70ae6bef8e73f97af252623c6e7d53e830117017d265db88230f
zf0cce34dd6cf2f0c728c21c2d6987d5d18345a355a20342c8878da6813052827020f881c5576c9
z106e61989f3ab702621733cd6d6624f035a146604fef134ade131e4e442c3aa5566d19a2588b41
z3787c91990923126649ecb5832ead702b5e047ffbfdf6942bfa77d8c6fbed7da9d93c5447c3bdf
z2dce6b9a0482142a432bff248784b9b4604ca3c6cb5fa2c2995578a8ac674a2a68e9bdb34b7e05
zad99faf0c31a8f8cbe6bf9d2a1d4ddc9ee0cd962e3049484a9d0be0616475bc31f0b7dd87962df
z2bd8875635e7c4c6a98afd5a0e100f4ae882cbd94b750b88da826963d97664f3c83774c4596196
z156ff33070c3871b29bf7d615fd94116a9fe56c2f0b5d751fc7ef188d4b63837ce02b6d4ea4f34
z318261802733a816e414903f34c6e51e6e55cb0a7cc1516957fc875006c5e4b22af3174fb9bcc4
ze6511b6bcc1b8672f6e2c35f934c805167069aacb7cb46335a81b3c91fc42a73b794c3f0aacd81
z70dc5bc19f708e809126d6b00e3d488a940d43b31b697c32d05185ecf4aed78e7c9676328ab635
zb1423df947de4ac65819c5f061bed19739581068ebae44a5b10c61f81f2977a471f704415e412d
z94ad785df2be9970b4e294d44b08faa17bc1218ce4fa1b5a4b67b2084d3d466375c18131bc0369
zf4676023fab8913cbdf4aba866b2cb0caf650eb600f08129a011ae91480285354d41901b3fc9d3
z441596437abd8f1475e6e3a5de3dabbfd489756130c4fdb6a2d292801fbf6a69060eedaaa8a4ce
zc78a9808e045a11d2f5c61113ad017d591414c57cc6c1f74941344ca4fa9a943e4ba00d70fb6de
z68ecfe94affcc2a675de0ec1d47cccd1a5e00a1925435976223f1ee7304f19e0994adfb04c8f41
zfea3228b75a11f6e17270faba07e0a975ae1b91e273a4e7e2473f29978db195d223b23f8a9b3aa
zdc3f524ad001722998ad71305db1ebbdbfd947a03346affb90472beb186e5686e7ae532a87a1d3
z06d78b70f41ffaaec569ad1ad746b5ec100af59e2fa4c2cf2f47e56f7bb7f55198ce7246316257
z3811ae2f22cd27d776e2d77d9d01d5b8c537ecaec94c9175d43f5e854307269fd6bce57c6ceeaf
z42322135a8602016641d9266c91b6352aff778f81efef7ea563250658042e9177ef63c498a4693
z4cd6aa02651905158afc5ba49f4a588feb7d4275edeff8a4f2ba57755f139a40f0afe33f77a4f3
z515663770019114fd2312ded892024dc597e4bb082fdcfd1efa4c4c7258da8b08f8e27332b82f0
zfdf6f6fe56415549e43119515b52673599aab1609b57074894060885dc92adf3c0af3d9a0f5689
z28918b434d6836d203e3bfe4cbbe1741e7cd575d3fb1aa4c157c1e42787a20b5abacd22f8090ec
z0b419532e63c9eaa3dac6dd5ae3fc24a6716098f4e81550a34886604917179510163c9dc10070b
zc15cbce4b5c350d43b926721dbcdc1a750204f101f463663d08d8761d8a23ba41f928df63138d3
z0d76ffc343f701669c8d5a1e9e40743d9cffa47e5dbcfdaa6f40a01e14b192280cd976ac25d6e0
z225c36e6c4ad5097786547a31e6f1ff2e09a17b455004a4bc4594bd0b49f74847c473680e653cc
z7b89378a43688d839a72849a3f525ac143829ff427052fd056b83485b978bb3f837689ac016b0b
z74b7f9b064ac49268e99b7bbff513f032bd14b9252240a82bd30b5b8da83a7dc4cfbeed9e10507
z607fbc9a79e24e6c8489f86af54265fd15726837173d55d77f28d67246342c3c7e01b18b5f1e2f
z315b0aff46b5482384303731ada6e8fe2f421e13127758b0a693b6b02f2b329578065e79b145df
zeb70dc97dcfbbb45e8d02a6e52eefc92a72523f0715a9b8ebb976a5c911435413da16a5c688b7b
z1d1aa3da44146a72822fb68c1e463c46605e4c95d9fae2f727779afe2ac7dabbb12ca35761b0f5
z30a8cc5d2f4441a7b82ee762480cb5578123a440ae01a875c66c7b9410743dbe01f4d5045a697a
z3f5244afb0d61a8ecc349c0cc0581b9367b4eb38bf51e19a46f6c8e810cfa13e03c6949cde0176
zda92c1d05c6440bcb5a0cab5e84916a7f6c54f1801b5a0bf0d68319e312e5e188a094f62190f73
zd27a9bc758d46c8e647814506d8d0132a3aee9abfd68dd6ad635202c287591276245b93e88cfa6
z6290276087e25d0cbbb0d9de404489ea12198614ceb6032108638dd9267dc73420821300a5e862
zbbcbcdff1ddd83aa68be9ac23f27acd0ae642a00aa7076df39c569f3a562be19a05c764c2bb578
z01006cfd7830135122d6a64876d3ad364667eb75dba07d860efa734175676398f5d0f875736443
zf1b1563faec68d7392ad4ecf8526d9d4b8746733b068c14694784568e269d8dd68bd388225fe93
zeef34dccc7e75dbee37234d32a7c9d1e38d392c44c476f60af6c468f2be94a5d3bf053b57d3258
zde156156f362f7ecc0bf83f8cf454eec32aba9081cc61c69400833bf6c87aca12c3ccd44878dd2
zfe5a9ea9cfbe4f555f097c642bab8f31da9ef549e09c2561ad05b5153463d63df805bfd728c788
za493fa2f1c1cb5611aff2edaf4a97a53b91ca2d854ef16c662cec46a581a382b5457194b578cbc
zd1df1b0244d0cac3ca8c018e27c468f516b9ea9d92dc07ff1b3417bd6d2adde377d08d8234279e
zaa9fd15a45642d5251cc3832ebb6718af7741ec4db797775d9ce0d5a43d6c3ad44addfb0d8bf3c
zc30f956fc1d5a77d4e2945f28d096aa90879e1f2d64982e6a94919b2898f32b580898fceacd3e1
zf2282ce63a26314b7b4a874961fb1ab3643e38a97c2cdb48632dff8c513047a5e7226ffd45aebb
z0b8154b5db174ade8e11190a398d574fd6164b5a078197114dd17e598ae7ac21d04555fa2ede12
zc3a693d789c6c418a7497bfa2a821a6d88f51625e69bfa260a9529b9c52bb0b1f794f08051003f
zf59d47e5f3eed877af668a31b40fbcd50d850d118e5f1628f8b46eb9f27fc7ed5e64aee1e2dc45
zf0e039a96452c4a1d5e3a5f1b7542bc5d9eaf257fa98138a6fd8f1e5f52b3f7dcefbf7e695cf49
z86481954f2e485401f62d6c5ac582ea6cf701af424c47b09a0bdbed48f94dfe0773b9ab44eb706
z4ac533c51929bf47bbe586dcf0ec3f28e01aac7278950283c082ec82954011e17d34725060b956
z32ec32cc48f615b921689cd29331fbf71eb246b1f9734f30c054eb105bb41f8fa8e687dc64cb57
z3332485920ab5a620b83e55fb0a4cd94872ba6057101030428f58867da925c8f09be1c41fe9fac
z67132cdf4d5fe53c90e7cfde7d7d13d41e1f598785f89514fa15c00b29232300958e9c15450085
z89a1d6b5ad31b5c5d32841a1b75b9799a39ad5907da1d6ee8446b15df7d9b0da403b8772190849
z69f9a7a174afa0640c5716c1a4f70cda12a4ba8d52d1093a2bad75f269ec25afd21b749015aeff
z89f42856b82dc208868557f1ba2631a325890d7d82b158df88544693fd24f7aac360d515dfc8bd
z234b4d21e37ee3dcf13c9f25a3018219fdebe14456a8c63d6a7f681034f11ef20339dd1104fd01
ze7dc980b865ea1782e1fa95c53360ab12cc050d200e7772044d84d041563457de68620df4bfd0f
z1bea5b804d2e1fe1ed92cca18a3362433641966a175c3aa9607898ea67da110ba5fe8471c5cb99
z60b5ebaf16f836a1f3b92f93b2f3b62892f83dc285002dde1f3227a06e5147cfc6a56ef4d8235b
z3cc7fe0a0e017ba3e2fa6b48f7474fb5092b1ea0479db35446d70c9aa34ecd2219eb09d7a18b68
z173807bb559609d2bbabe486d5cb13cc35d7ac16bfacb4065a027b6968e4f1bb627ba09da24a9b
z9ac040a9486bb8e23aa74243f51646bfe00d99d04f25f4e1afc9628e59dcb4eabaa4ebeb01c623
z3c2200fa61cb36f98d85028b400e23e4abbbacd9cfffe6e30cc2b87877f5249710e71d44bf61ef
z3ad1f9fa83cd8aa367d6c524be13d031f64b3b7bec7b760ed854a3aa3cf9f32d413ae172042321
z63a4990ec29e4e8ac003e595464f0549b8aee0e45deb1e339ff231f014e0f5ace2847f17eb0196
zcfcc339ac5c7255f1a65666ed35eb3ef9a1dd31bcaccbb8ac0be815e089ffae5fc11c3a8f9f81d
z9588d79da0481afd2e85aa7371a3279813be49d3de927676402b55aaedcc722f775e7e762ef386
z9e842cbc93b54e49be6076729bd361a0e9ff2eb2e819a0d64764840b9b5ca827d2d2b6e71528ab
zcbe298b8ed7364f29d54978be8b2baad7b83d37e8c73ffaa3ba3611318c39c8614ca50bb5ce8de
z890b9cacea2503d95d1b63cf4495da9a3fc23b35a193c79dca31e27d19ef3a684e68ad8b3e74e4
z49a636f119ca32fab2a3188337b423aeefe7794f9d7a4f107f64aa2790c3d731a45b4a397b2dd0
zcc1e679468d58ff999fc766fc564ff4ea63a46bd6d76bdb2ff09019cd8492639b5cc71552217af
z8ec1cd6a10be28c10253e6c60128e6a1ff0fca4a68863bf731dbdc51ba018ddd49b3cea6a6aa85
z57af4a55760a28aad9067f5a8e54582ef8bbc5aa9f87ca95288f8a8a67cef8814b84e4759d1091
z97bc203da4a2c686d50bfe62563c7f91793147bb0c0a875522fe9f6cb2ff47ec7c4f02c343c4a0
z3750863531261c46982f6937e2ab0b1b465a6ac68b777a2f41743c15bdc7af00af78c161c6acf5
z872635092f9e391262bc3307692b947c37f7205232c39dd142d8a43797ced66d704bc76ce61e5c
ze902e675325b0eb03ffc6b3b587ba5a694cd592cab8bfc8b48c3dbc13b8029f15055a748a24d7f
zbf6961d8819fcbe39be5bc40d29c24db5d0db1ce8a8e0587355aac41c2a00784a464803fed5fee
z5353c122740d78781505aef2521d2b61acd71e17272be5cea233332f60e6e91dea0550c25e3939
zbc654edda438a038e6ea272c12c54fdb3a575708564847c3156d6bb83db8b39d7c66b9a11f97a5
z0c0b8b4713e3fce479ec94a3d2546db85d25c7893b4abba9f48be28d93c69adad85d7e85e8509d
zf1335cf399f775f559561023dba6cc6cf14948ce50effa864c32527c614b5e1c9ed41c1dcbbe61
z3de2eee2f8c62943995f152e7fe135e7d1aa25231afd88ecbc1ca9d00eb6149df89b6ea58a10dc
z208aea17e0e538339e9f053cbfeef6bcbcde33d43904d5e06eca2ad09b213e3920bc2e93d58d76
zc2d257b85822df1d4e16037f7cd78f84e652ab4e6f73783433c90a63a26866ce0bc9b317ea29f3
z13adb35ed9fa17558e61323888a5d41fb532a7d3be56783b6e529e08540851d86698a64749c152
zfb1636c3b66b807e55a930d6859134196de239915b6ebaa9bac7aa9de4f38d25b70bc4302cb7b9
zb32d81f0726fca06a9c5ef7a577dbb7a2e574455dfaeef9824b6ed899134608b0ee2d429bbce65
zc3f9149f584f37a5957162f6226f6b8d6f7aca0317e6682d8e473b0dfa56d50ae5a6fce37850ac
zdc111513a7ad50724a91165bd376e80c220d54ace1cbee46a8bf577caefcfe10d085442391eb4d
z58e7c9e009d30304ead4497596036afc679de159ce847e7909b8b6d9885856ed693fc1395795e5
zed04cd037db2f5657f933e4d14172141e9bc8f486ce847d2d674846915863575f382d22cd32acf
z8529a6fbbfb03b5fddf282b1d050ddd5710cffd169bc0106bbab591b34b93696a9dfaa5b6eaed9
z80ef379f627f3d768b806abf5dd2ea481d078c7b97f3083f257f3f0c1d41019be66bbab258238b
zc13ce611e0e875a345b7a725c05bb7b16bbee03fe7d30b62d8f1c18ae5aa2a0344317965ed3a13
z7c349fc86321c34853a11afd28c26c195bda770da171bc2eac67d84cc4b45b654b7d854bbc7018
zc22de1c7eafe2424bb3bbc19e09877e1daeb22d472356b690061e67c4dc6728432847a2a551232
zf37df5dd5472257f709cd61bb22da9da5e244627495ee81837a83a3207fb0b9e9394a41116ce79
zf5a3f086ee9a3ddfe24144296dbece39eb768ebde9d21cbff3a8050376b3bd6e0a2820057b3f77
z905c340c06a205a6d4901f944e683572de3ef5352bce789e4808445a5c43fd17fe21958bd076b7
z094190e0a64e8ffc2804499c10cbc3877dba9d2be54d3c6f396cabb29072b69043efb65fce461c
z2158bb6821e96d5060f4713369fa18e6dd68830cc05a64ce3bc1316875ca6cbd821458fd6702b9
z87d9dacf6e7ebc33e8eb5f5f68360b12a8f9ee8f4b8e8be67cfacd9bd877f90c615ac25b63ce4c
zdeb0b872265b8c737bab7412aa717f83b32fcb92498581e8d819890215b2ca24b286ad39c5f768
zd7176fd4ab9d2da854f2130408cfadd63532a1acecc2e0176667eee2d3eb18ecf2ae561eb7f432
z9301ee6e096efa45ec1c31809f9657abddd158835a62e56f9f65f9c74625d76962177b753a9dfd
z65c691535b407ed64bb71e58561e3bec6e0f8f220b8e6af4c3e041c1e5583f09f753098d6b0df7
zac91bdb6b4943e77671bdc690499180c2a81de36dffd3d0c170abe43789c542b41691d1cd4f5d5
z013e764dd6e5e71d27e511cc3921ac4c43aeea860f49831259ccc4f7ed85837395ef550e836704
zb19d6a819c7480da2806bfb8aedad1c910cb6e2225e58ef74aa9cfae3adcb8eda4a7293ef15592
ze088fe708dcb44b9abbe40bcc2ba9bb7cf7c9453b583bb646fc057643322059051d6f8be44e066
z518a8ca66cddb6cbbeb8445f3dc650bb9582fafe9f10599180d19c4153a2514a7c9504a68f812e
z0d7ed88f4c04b342e4cfcf824464f4f4db931b91b0c206c316d8ce6bcee755259f61bbd56f3079
z520eb66bb7e8a6e95cbab5e868aea0d36b94d92089213bf5397daf4c9a66adbd2c54583d3f0597
z970bc5d7019d6331c9cffb9bc270ecd74d8e7b0b7008e1d9ddd3324bccd7492d9e72cd878a190c
z7832da9f3f4e8de94b574ab158c355bd832c053928159a69e1bc38cacaf251f6c9f1af7095ae24
zf0bd84b16cb0ebda1f533ade40fce393fe6f72bd67a4ca7fbd511645937380b741df9588da6cea
z664b97b865a63d604651cc050ba096a4c21948864b625460bf426bd860b54360f11e743c926947
zc21b132cb17dae407b76f63117d670b716e0217a0896f21b50bd8e71cc0fd6483349b96c603e23
z1f5bc34fe461b685ff3dd1b62ad1f652effee1ca2fce4a0062b3e092d2828036055c38cc5e2aa6
z81cf9d26c4e8aaa35499821e3f39f55d2e4be8ba32c0f92f30baf24e04bac5622ce3c67896691b
z76a54b096249532d9240950a80e4f654136b748978c58307d2a15e85718a98b490736eb781dad4
z78bbd9f3ee056d7877e0c16c0b979a2a2dba8e33b16b2eda28720913ab9f7cb668e96b4b917d07
zc21517a4dc28e7d1aea06208ee467a67d3cbe32373fb2bc3347791240a7e0f499f05b0aa635b3d
zb3b8500889470524e3720eb0d41d5642d5a018473ba0cdd0819c8bd12316a283140200e91f64c3
zb4bc2c5926f4a0008f5ca945369da8ae162e511ab370dc3e62a22985a3a35a4e6fd3004d688756
z8c2d49110b54e639c1869f29a17849f9045d53701a317389c41a41ea5619e699f2a19e9919aa42
z968fd3ab9b766f4b41cde4a28e20853d66922a3c1e0bb211fa6c4680213b7051d67df370e061de
zbeac2050fdeb36cf07cf26381c64699eb7d9e52afd7bd143a5497cca98ac5a4b397846923a61a5
z1dabf9766a6a3520e21f7f6a3dbaac40385f5aa9dbf839932b0863c8146be9967520189bfec254
z83fdefd38703706ec86cb61aa20b0d20f60f3dc22307a5357003310331457aa6d6017ba0303982
zfca336deca36b8f333b07d2118ecb0695a88d5b0b6ddca519917f6915f4005fdba3abd82b8458c
ze279834ee38a84145674ac48dccb5e4c5e4048dcbcd352b2933e47d64c8f9621b2615bc8532de0
z50ebae22b1e601e4ac24461b9bc3a5af1cc10a6c555c89eb2b7c9e13378f99a252eda99ef99b3d
zf3dc665bbe566bb4fac6b11fa45a8bf8f5701681102e53941cc382e6b709b749e1b85c71eb6bfd
z799c24dc27fd2b308b5b41c15bc0c2ec257c93f1eeecd892368b86f9397acef93825be3f3a2e21
ze75c2e3be5eeb720c632d6637c1e213c38a1869e9842f6bfb815992eec02fc2b1a3da9529667b1
za835cb8092f215785f8949e9917816878b67822f608a8440df45067bf5459065d9ba733ec75639
zc852b2b7b4ded66d5e220d0ca34fdd91e164268f45767b02cc2cdcda7ec934b39fbd4de91c1f02
z4da44a98013d0c9fc2c4a4ff185ab31915d66d757076d567655a190842e20bd9e46f570754db75
z76723a5127e4fd4e91ee835af1558368bfd6b1ea1cd7a883717c2d9f77309e192744c843d86f95
z37a693812de9e538ac20eb2dc6119cefb48035de496e7aa9328e176ae9444b5f2bb99edfb8d92c
z96cc5ae09f99760bb7f5272cd94f80ef6bb0fc747ef4b49c8cb5894800d37034883da1f330362e
zc63c1350dab47e07b0b88ebb1757afc0b15ae5eb9d45df4c2f7d677da4d50abfd81586b6a6ce25
z577ac9cd84e99a8af029b9fa77dfe22b42ebaeddf366845685133f0d18e1a23ce27d788402acd9
z16540ad32fddd23cbcd9a9ec477a8009dff269325d824d3d0d6a4e4f72c1711c458e63b1102699
z9a09b3c1ade6486be623330487309ec70bb7c49ebcffd0998f7d227f56f0cf53da7d2e685f407a
z6b03a763afd58c10f0d47b4dee054cdb49fec702d5bc5c3f662c587a63539900335699db9bd22f
ze7af14b124d82783bcc513188dbd02d1821a51f13d46bb9c6e310bdb1ed33777f0a97479f4c5dd
zbd8b8d64a89d941f72ec60db4f7c9aa1a66d15a6fde9d85b7a373670ecb602b285c55219d88ef2
zbc0bf1dea496ea2840fdfebc0761a30a2e6107ede128b3d40fb90eabb6a5bf6ee68861449287fd
zacd51eda386f163ff4375bd58690a5bc195b86f9f37657ebcc668c68e6e1ea92f5188630eb1f4a
zb348c84e8e0dfafe18355462187e4e1f19b34e1d24b59bcc6a6cdf72c6bf5e416986f9821b50f5
zd04664ae0e8cce79d302552a51f7ac28cf2f393f5b1ada8daa69ccf43ab3a931644c2767c0b6c6
zb616f344d745de87d2c1f10132930ce8bc07a76cbfb1fc6982090235dee54600bd22419cc5b5f8
z02420fc03033de728705dd1a6f126949ba03bc40087f592c0b497d6d1b66e680ee8f84e62f390d
zce5cfd878f41c92d358fc54f9bb1c5ba5d1651b18a8f77819bf2de7e5ec0f4dbe84e5334c7bb5c
zeee2bc21d8d70215f4852f8d096c51be0713f7093aed8ffdab481ce9fc0d71669ccde95c2b19ed
z7f9c9d0ad699b2943c8f7b4e7b5259a26020f44ca18d26939c1a0909542bb133b94ce7d19fceda
z7ca27d4796ba019459b31b81e6e11ec8290c2fe40f8669442f5e41245b9213dfdb3164755b7cb7
za89fd4944c9ef2a3608418c15551b263705fa03d93344b5477c1162da9607f1b884b494a136463
zb5d15238e7c56ab341a122c885c0b90ebfa6dcbf6b38ad1db1020dcc28dd251a2d4abb5aa1006d
z13320f62bbf499d4ffacd334b93853b99dd272e9c52291f409ed605ec1f25dbc35394df25e430b
z3380d5b398461d2d254706541300c72bb897950403c78de312be78da4ef5e48f4cda331baa40ef
zba171c0f1fee42800864ea9c4b6422f65f9080777035611c42f4e087196fe8a10a72d4cf580d1e
zf25307b0973ca5d9de9087f342a0e767a01b6f70f9c6ca71619959cb6ce06eafc60ccae64a24b4
zef8752832c3884a1c5536aaa11e910947401bfb66149c3a0d2f5cee56eb93a66dc73746980c158
z8a1e6c82e5af92d69361a2e1c5aea93331be55c53792845e5887c28a11cef7de2e1f237d7817ee
z7aebb72a437fb0974ffe1492f47e2f8f395c355e6c8638e53b347a216d71a176035388a440afbf
z501cd47ded6ab13ba2689025519744d88003d0eeb43fa2073f6d287c58ac8728607a7ea015f55e
z9d6aa31b5ebcb9fe08c364627fe6e75a2d35189e854fb2f2af52572b46eabc8f8e96313e58e862
z0fc26241c52bf6b5f46e56d7bada8e40032e8e4a23fbc09e3dcb36523774a2b4516420ec527552
zced702269ba7cfef4d7dab70577697553edf08ab2d20ac392e541d3a222f5cbdbab916900b1eca
z65e2498769f8a31dbdb886bb5b819c7ac70ca3ac3d8499551d7f222a9eca881bd3a67a09f1a95c
zed67d4b8c1174943bbb3b0f85c50dd74cf8fedf6eb0ae0453e5b51ceab2a5cd4586ed072b7f957
z3b12b1c63ffa2e653c7087affa330c45b5f3faf014046cbad78c0979807bfac291298d315c51e1
z5ceb395f026bd45bfb4c78eaaac92ce33a229f2f99bfdb6a9ffb5fcb1dfa6f0095ee61cd926ea4
z2cebe4354d9362ee3cd233dcb339a7e8e6d931f0662e9ed8075115af465779f4b652396e76a88d
z0ff900a9e24c2832217a037f1660fff6ce070b08f873fd7489d09a39fec70f3ef2eae8d2144249
z2a92a8741978e502d2878046649e82adc4cc7395c03111240de1f655c38821f1add304161f3d54
zd6211ddf79c48f7f73bb6ed8a47622a992e3de60def23edbbf043d26f0f185a8ef31ae2103509f
ze336a0230d88c62bb21a5546eba71763ec2a8b10f726ca4656b9cfda00150c755e3905c0373bda
z4661962caab5c81d0c337905a95ad673d1648c30dc6c164734380d48d77f25a584f3116f394fef
zbae67d54b1d6defdc1dad395c6de6c6122f3eee7ef1cf7234502230ef5ef6ef5b63e780c374f3f
z03317ac988efad8c8bee67605eb1e129b312f6b655590d727cc34939f6094899996e58368f4e5d
z598511f848723d30997e5836cd28113d110107dc8c22d0131c8aac702c3b0781d9b7780294f77f
z9cf20e2668c548b093209f32236d44664b3dd2feb2a199c05b34687e5c071b411996873a2b853b
z7d02c2cee83c882a8f2481ac48e1cbeaa6111a1509942f291d2893b9d6c562958e96dd89e59a73
zabd0cc108c825b42e6965b200dfb99a58238adc28d0772a21f933054d6b472684b0ac299f307a4
zb75ff0065fcfaa6c881fcb91a6cb4210c21a48e1918b108951aa1688aacb44497bbdcdec99fc05
z068ec17cf52014a1aa88929489b3ee6e0c4c29e1a1d075b46da97a8a56202824f274d7acee6279
zb614fe5fe229fd2f474d18e97e2b5f7f8291d22198cde8b42b2b6057b62c73aa40185dcbba7774
zf754c54dfbef4deb25ba2077e8c0a8e583308fbc3e447e2a9260476e1cefe9b64c4b6d2384f626
z558ad7e9c3c41ba2d75493960593cffef94460050e9aa5b0ca1e55bfa8a8303c25c92fbda4646c
z9099203d12b10b83dc55056f22afebf22d8ebca1d6fe069148ccc9cd15d00e8a13e41c40311d63
z2ee4cee7d0cc01b070a6a34de51fe42c444d189fe21374615b8d38238c73ed063d960de4420b84
zb347bfb3e9d6458e4050bb0e44dce278172845aa641d8cc1d0436edc53d5432ff43cb1e3a98062
z21019ba43d57035057036413c105f9c9cf4e93c5b45d26cdd5a7f567e0246866a10cd8833ee426
z5813bcba04c26d4fa7375871f524b29c89f383aceecadb5e097262d2fbe5bde82ac2b5825a41b2
zeb64c87fd19560116d18b66ef2c7b913049bd60d34727392f144bd84823d7a9a4e4faa90e1c72c
z429890f03e3c4feaa2d07ae2012b5fd9cc87f5c9c56082ca055b664c01dacdd50c1015d6380cc1
z75f26bc4226b959a8e57482b1d74d16d5d70af0932fadb026c08233f8e47901b23111ed375d018
z17848e6d6266eba3fee05651b09789adc626bda368464c9785f0cf2c20fb3fea2720c766ad9e78
zbbc8041a8f7b2e5ec7a0ef8125cb16750d3638a34ece23404c358e1b235b7e7d0aa2d0881827d4
z14ec5557cc4c457182cbe9f14677bab8a03c325f18934a1cdf511a5b60d01737c0783cd6c92bc5
ze79fd52cd50d05a458a7a2ce29bfce22fb53e9d43912e7c66070c417d3ffbce8fae2142de1d039
z448d4c513e43d827a723658a831cdb04a3146d041d6609b747838ba06cbae88c44c3c3fe89eec4
zda228c4e758b2e0d374e8ae60e769951224e750ea564be74841b2710b8aa20a4550078228170ff
z9cce07ddcecfd0f77b6d73e17d002e3562c5efd844cf6d7e32b61079901980324109caca43fa02
z7857cebc7ce6614c30f182aa03608cdbd442b13a8c8aa68ffe4a510e9b27cbeb3f15cffb1d6295
z8ea7eeb9fa00fc5e5368dc6e01957b0de9767b29820141dbffc4fd604f88fb1393d6ca0c749e8a
z6d941a6b6c387b7c505610f291fc963a945c80ceb14a10fe1961edc3e147003c374fdd710a0f7c
z4d21d184395d15afce01ba1bd4dc1e6975c3d513e14480f45b3a1b32ee26f6c2932b7e6632af1f
zee865c7d3ad5df4b1abc375cfa3084b70322ad5428cfb4b5257ebd897411826318684282566c36
zc981b9e2409a10eab4d2d3c8b8f1f22aab6fb54324ddc5f57d9dfceae9e4e5670d5302781d3dd1
z79c0fe88e584634a1cc1bdf4680b08ba727bc816f1668bebdb7501ed69695ff6d3d59446c1fdca
zab6bb8277c54b5259461e27bb19aebf52005b0214cea856a87704d05c67e76a6c2a7e5dffe4fcf
za6ee10d612c80ad4671e7527bccf68c50a19dcdcbd1bb37f400abdc62eb3ae83b9b148564bc250
z47f57f69fa18f3cefdd704fa4967a9370365a6e0caafa3c13e122d2c5a267cea4f9eb7a0f55e90
zde664953869324747ad76cd95de2c51766570b5ddb3b2074ed8c481eeaba5024dfbf1bcad8082c
zdf48d03052ba75eb2280e2b74b3d80ce7ed01382e5f5429755a263084587a0e062e93987fd785c
z2f8073bface74d36723221933f127288ce6abcfdb0fff8d372af662456a5c76d698439b28aa6cc
zd8dbb4c650f3c74a70d2c5f98e31d9b151e6aeb1725a59f5645fbd6ec9d58f6a7e86b8e296a228
zc261295c512586d9ea84aa71a618b355e067a5a6e1d1050e37c21be0c7f5ead0a9bc75c9171cf5
ze83baab7533735b29990fce6af261408f85e79bbcd63fc0666a045da6591c08d1512e4ba9a909a
z5dc781c02c6bf7b9b6df3916a904438e38915bacc3097b39effc77a881f0c575debb9192bb46a4
z6db8b655af3b88bf51084bb71fd9f4207584001057d611c6b4e4f4d1632ca90ceaf02973c25d58
z83485ea30741d258ff8a37ca928e29359e795d90d6f5afc2750cb9bf7e154c6e6c827f0a3ef94f
z05009db70d1078dfd41d3ada485dd0659f2c73c7acd7c2536072a8376ffdccacfe1d3b41258c67
z4c0c240f13335d224dbf62a82c9162c1fc6b5a0aff805c411888195d3fb6b47d7bead7ec6df0a2
z68f7e00328cb56cb1e5f88a25d6250777da20737bd954e112a81653642cfa5d7b0d0828e22ffae
zb920ab4e6caa7010b6736977e78d08a91d83a78133053494e18573b70f38af7fc90a60d88e85d8
z643cc250b9a836f4af62a3806418774555cc528595d492064aa54da86cf8f578d072a50a07f36a
zddb7fe1710df3b116bf1eb8d0bd6a74c16b950eb2d5dc7829638d08c473316815acf5e8f52211a
z3263a839342ec945417edbf1271f0f3f1955b3c9d76c893ecdefae346c29f743a35d82bd4de180
z117434c070421c4017827403ec3eda687ece4da8f0aff6741dfb6ca57110ccd7ee96314096f953
z01ad8b03756de4b8751b9ccbc96b6a8596def2133a2a6c0c2b19ae34865d5347ae07c49f6c6555
z093c7053c053c6f8fe979f2b3bac5d7fffdea33c309d48731da71860372727af12d42734dabdfe
z0d66f02aec458d8b8c2c342da324a4d6de00e32df4bc12019050c60d9606929a182ab497e69e24
z1bd4624a2912580340e1cadd0b8569dad10e4f16ede4c80d42d0dcbadbc41ccc1e92b1acc85d7e
zae6251dca87cb60bfb910ce77d51e4d1c19d726ee99f985f1cbf7b795c87fd5f2192f14d986190
z41d60124e069bbc7e9329eb790a6de6f7fbfc3d5b615fade3b24ed94954a2565aba992fd726000
ze35c0924135ded8a16d9a38a6d597b5d3e6cdc79dd4c94317cdedf708f182c2d219a11641d650d
zb89383ece9d1d41635af709e38ff5fc01b4d035164f8754548e120a2ae5631d6f86260a4eb9768
zbdb0c2a849e9d808fea88fae77a92484fff9289feb925881b255158a717fc50c3e66e7e50493b5
z908a9d74184e12bdecf9d0432a51eaa43e8fd77892ae243ada64adb9d9a6c6f1f3f656b330215d
zf792fa84b61d21bbc7d1a82030b851ff8d68e7890753deef753b91287281a932dc00c4edcaba34
z446a024b3e3c210fa0f38d3a36a8869b5dc1b8e05740ddb5978d801a5ed339ff2b929c05b18d95
z11da46e03aeb3b225157f2a04128c403d2fb26add4a999dc6cefc5c6df6c07f0bd992f9eabee36
z84596feb55d6118a0f4aa95aa5113ea18243138f46cf46ff03ee1954f018709a9194f3369a2df3
z6f7d25df5eef3bf1235144c7b050fde4e1f9c30d2d2c1cee251cc93b744dd3baf51e3b8673f029
zb773c7bf2f929acb6549773d56b3e2ce4d55bbab725e0b8381bcb10570fbd40929b4c16fec0fc9
za546807b9246a5610d1d289df29373f58845ad70f2d75ba9f985b195a475b83f3572c1d6f0f534
zc299c73db828ad68c2d8b992a53ffe0bb254e180388653740ccee48131fad00a715a0a883afce3
zc665cf3b682ac0abb504e071ac3da744eb1e59c80f17f9d49cf456afe1e088fa94e5c7fb057a02
z4225c9dd0902a4fe4ec269c823ee97f9c519ecf678d71c4c9599e3c14dd2971be1c381b140cd6d
z80677b199dd85ac57cb7a548615d8bf145668c3367a1b0a365847ebe4c4484f7c19cfc414f131c
z58d1decb52b3833ea1bc04fef4469bfdf2ce2e7d628b1653cdd897883c58c1ba4ca0c1074a09bf
z7a8abdc19844977cfcb7a54ef2c5e691596a4f8c169f5b2745927bc5c49eab3f00757090e623fc
z2d14d950648c0abc8717286ef4d889eb0fc81dc4e9234e11cb4c31d33c835ee7c3bd1d41482e44
z7a58360ad05e983a0c9e6797653f9cf2859db77b390fbe3799eab6a5899c771ff02c0ac5d6467c
z5aa7210be060a0293d8645b5298d8d3d2231d34f0c4e51b41d7dac59ca5d064fd7687d70d273d5
zc8a9db1a44d293dcf0f31e793a9c4308c7d5651825bca01ae51bd35b4cacea33f3191858ab58c8
z932580e09ee326358e421f909fb35498f83a1346b5e61f884c692a064c02869c559432b8e43c36
zc47867b3e6c6e787be7e7803310add7aa173fcc318a76a1d69b484ef4d2c99c0e7d5ecca3132fd
zac78652acc6c6be378bed668224ed443eea8788a7b92309e51e08004188c2042d83586863afc25
z28b6ca11a976af9de1714afca4fd35abde0d9dd5e259fd7f5e72ed29eb968056f4ea88a15e5419
zb98392e91f59f4fd7658bccfc9dcf235dee3002b0e6b9dc48da29771406ae7d9dbeb54a8aac6e9
zfc38542629bc79a4d891036c6e317b6a702223f32d4d03fe1981a5240c3b08085baa324a79d935
ze08ff5158405a22c9505079998a54892dded682f14ed5073759f996a610835753629db9e5b85f4
zc74a91ed2290f184952438091cc64cad8dbd8d36ab2a428585c7b112e27d4c712cccb2f49ef444
z2db70f9f714e3ed50afe32553cac11ad87cc0056920a1eb3eb0b41eb3118cc7dc23c5093008826
z2501f803728f393e942fae3f33f03d838537783d42e721f9ae4f588b3571d0c115a0abda1172cd
z6746b60c54ac77345108badcdb3184a91b6d9bb6b8fd14f554cfe5ce4de4c0dace6c0d63d4c4d6
z55f56f07973698441f18e62ac0321b718b0868c209e3589c8c8da18b739e069af8f69401f8fb45
z48edfc3b0d10c20cf8fcf51d8f4dd9124f2117d2c9b7df60196f76ee1e0e4ceb593466e487e6fe
z40de62ff1ff84fc32484a58a31f089623389320d829adbd78906b7042dcd4093eccc110d7aa8e3
z2cd814e3a8d967da9ae7c6c5f54305ecf53fb6dc85f56e4782bf75c40d37edd7eed10cedc84fd5
z4c671a2242099627afd57036f9f0edacf1b11b8a8ca25ad63e3a8755cc132be45aa8f6a8a58e86
z436b9998354b26fec5b5eea22f02fab6bab7bcd35950f24d7eed3d58ac0dcc5e14916da37f99e0
zbff3d177c706986664783e3e710671777feb19e49270fb8e5a3fd6ccfe4c961c398b1080bf4bbb
z5798b89b5b2e359948053b7e68918b0ab2be231faa34e3ea06f14a7fc1ec175d4ccdde15667b93
zf5b209e487cb8b8cda3c09bac4502e13bb412d2d0f08816196f52c8c11172a69101ba70ea86e56
zfbcbf0e277f1870fe080b05d42f5d64e956b2cef320a4c59129f6691bc8aae49942080c7db1f7e
zdcc03aefbc6197bbfc765fb611a93d61ff3953395a33d936782dfb631a8e7dd86eb748a8499d10
zf04196cfc7a737607fdc6abec6e64d0c80c90f3ed24e3ae46bd4e9a93343cc5b3fd3f7327b2d0d
z36c80870babb2e91925809c4efebd7525bbd4444693b6271425029b4e44f6a4576cc06b1b14fb2
z870b89f1633f8a1bbf4a9445e4b2f18bac6c860f4d1f343ef5dccca7335551b6d168fc076278e2
z7e5fa6a05baa1b5623c5307b768ba3e5c3529a52c259bb4ea90363187999e45f451ab4ddfcfa11
z6cd6dd6d1764d4f77a59e8e270dd8a2cd1f0e35a5ab5c489609652b7a67ff98f7c61d900f97efe
z8834209d2b13d20475d043fd4d60236ccd3f8849ad6ea59f4b44bb3e203e56f1511d5fbb595973
z6f69c0c93cd094ad322081a6ab967bbd9075c332ae23b0ca748689c9a679212fc16c374f77a4d4
z46ace1a0bf62fa831c6ff7f14c9ca6c8cf966256c419f7a83a8b6e0ec2a4068c755c361132c79a
z9663ad91f6eecccc23c921d55538ecfdc27384bd246eddcd9f849ff3ba91cb1de36ead1bf34cf5
z1b9ffba2d5f8f8d5503795031487b4a15958b0b201ac93e6de88df29568a451e783278c4f3908e
z7fcf0e978342008b6fa1e900c634e4c6533c114a6f4a64c51a06c2a73b6c4ffb96a766328d154a
z6d832aa698857e1fd9874e28bed3514b9006a237657060531a3350e5fabcd9952a57a56901e1a9
z8ef7c83f3eba9bcbe01f55c53624fab48b0d800f27d6f941b6b92590a2380701e0b9afc227fc9e
za3df1aab0c85a68cd766aa2d0261f0732035deb172f104103bc3128b92d267785d7b81569c4a37
z45bcc9bbd9ba044857890c13161ae66be81a0ed427f72cd75d53246b57e690a9286fb3cb6a139a
z7d1cc70d034261e4a3fd6b94f6d40e2200b8e87ef3069e30601ea2cfc3833457b77bfbcd7d9602
z6ea851dff22e6ced0e52c52fc7cd31e0db649112c60f4910d934edac19ae56adfcf4755ca84cfb
z5d0bd30e06cc53e5eccb3a7fa2aa3fbe05b2dd0793c31ed384876bca3365bc2564bfa15bec9fd6
z1590348887b69dacd52ad89e0e0503f87360c9d20ec96136b6af9a69684b99d9f5dd2d29ee993b
zd6bce161ff9a3bad3a4527a98ba227179223293fdc8cf8f3e64719db94bddf49952a99943163f3
zd7ce60b746eba36175c39510e40b1c45c63d258d489196f1e50e4c3c7643a903a1c5a0e9e1cc33
zed4294e9769693262f8995612133c7f54e9794eae2e8f8e242445470b3006900612d30e821eb00
z54ed572cdd04f90346209be9b1b28b3d94ca1d8199ff393a3fbd43275d7cb338cb1c432b51c6f3
z23e193e847f0255d4dfc5fbd870795dfc60cff18a3adf70714853ede1641a43fa6bd12dc3a1dd5
z9d98747a3b426eb3872c1fdbb38fc934f1e997629443ee671e443a84338a0949ac56c5d032a347
z2654592ef0b9f61328a3718bdcfa2afc8f65bee79edfaac8426cdd8e419b21e69e64dd23995065
zbd29c6a3b637c2caca7237afe98b27a074d6ea43e38f047a64ddd3ffa7b2deb2fbace85124795c
z5c735bf4acd990ba993b39595bfcdaacb68afae4d07e92e1b93803497c84725107d02e2a2d8997
z0d2b8693626b2c4169ef95eeac06ef4899b84dead4e68ea29a1f42b1c02fa1bc625fdfffb7e8c3
z710fdf59a991acfeaad839b3b8e374b4ea326b5113ea4d1c7dd32d07ba45e9ba0ccf35f3c4633f
zc3fcc2c68d9fbb7d86ab2f4af1a38273ae2d1c9e07c8f6a87b0353de71bc4df1640e524e3ced1e
zda351cfbb74ca96e7b84924616a77967c8c5cb708ad43ba211498a879ea7f46a68008bd4f24254
z9a62845daad71105e94ac14799466cefd78a0a96637099979d16a0349b216f012fda3f81da7ce9
zfdb7e97e6aef06e729c49e832f13fd8eacf6e4e0ec754b6b00db1a1d629d9e80b6b836a542c578
z506862b19324343b4b9adfa3e341dd36e9b572af6c6d57788369756d8b89cb79578340c88905c8
z34b4687a00ba4e8de0951e2a131bd3c5e1c25052dae1bb17b5c4e25a61058afc0515258252a8e1
z3045752f39d453edadf39a3b3e9ba5c7036bbb50886ff0436fa001438132bbde53a42590cad082
zc0de8a361461ea6a1f48b684f953a746d76582885bbed92984e811034e45372b2e270178db6c7c
za03e6a8cf6a699d9a5c2327899920c59029c12a204bc00dc6b3a9b599ac9ebb65c404b5a67bc9c
z8dee2d3430f747f2f32790b80e5311bb385792084248a4dd5f5a136d5d451aaf3f19fb30edb4dc
zd5f8afbbc73398414a5ef833ce0301e4d9d3228bf12a93a1c4a92c3487f9203696311e985624cd
ze1585cc8a2754dc107f9ba07230256d0ce8d8efa17b122a6352013cabf090d96e79d88420ccfa0
z4fc6491acc4a123a2a8e5743a97ed5016901e1881b4797f75177593373c53b64d867f430997d31
z28af1855efe033e4150d144edb8ef6887fa3baea89d97102fa4fdaca720fada9cd231fe46a02c1
za0a9fe1961f0ef808a81129208dc79b59d29f1de5d8a8203d6f6c804c81cc0bd812e38849aee78
z510b4e4a449e76f826e80471fdadd9a5f686ac44490cefe8a3f7f5b229594749bfd483ea16eb90
z65d3063d281044ea9fbecae7ae463474599b897fb775bf38033e6657ff4af786e042429e5f5e12
z9250e3ccda02755302e76f443250a56314ce41182475e122670cf7a2a8c680b46be6700f830638
z53cd6340d2cbbe099b74a35ce8b796541f2c053c84864e2854b918fc17a0cd956aa4616bdd373d
zddea6c865f18a1b970eb4f7be3741eec35ad5cb8998a0ae98db1f63ce2f4116ca7761cb8c7e296
z8b21191dfef8c0638093dfc34f44480b7b5e740916a4ec8ba65a61a4edd0f24bfcabec960b1908
z81ff803e8f5d4ec21270fba91e6783638febc1a3d5429a588be04216c168ce932889cedef666cb
z7d8f75a6b607e10f7d58b34f89f6b5bbd61d637628c226d998c354861658ba558a9f8922880111
z5b9db7b4dfea905edf8132cc6be5c6de6a1bfe630204838c0dbf6897ec2ae89f32ababf3b10d31
z3530d6b6f1096881795772cbf8a7d9e66d636dffacfee43205916c728f6d2d490f86452db97cbd
zeaaf653c925c5a3e97a9d34f415d165019885ec88c03071a9807fc666381ede0e45fac70ca68a5
zc358f39d6bddd68be9f736f25d090bd4dab941244a93c317c8ae76a3c49bcc59c07d58f2e5efa0
z7c240d6bb9470f8422a81f107d009579189ab4e950eef33b826d5c289e88096cd584dae52a3044
z3042217f321a4a77838b4fe22811956edfd2d24dbc4321cab9b00f5e95c6ffde0c4af5156d6184
zb226c45d16b674d39d2ae0903b0a3cf82c4d52bb51a6333b96dce90490776c606d88e0fb6f86ce
z87665bddb2d47601bd867d5b19f05070d5916e0b393e895e305e97bed841ae3c43aab426d89637
z0fe65efdab4490aeced28b8c1525a061d358e3133885ebc07ac14c0a65587f954de62acee77aa3
z7d0f968372b610e8bf47b7ac06ed61827cb7da31078111a526707143695add0cbff6d01238221d
z7fd2dabc3b73189a1e0c58e7b8803b3575cb6bab244bc51df5e8d0b58696f068d79f06e0b13208
z36875ba5bc3b2c6388e094fc89a95f849892815ad534cd72e48f10a000345be00791c0547a4330
ze05a53f653d03aa70ec0a8f925122a37233c0aadc3a5a9705e3480dfb3f6576d362005070abb96
z95f42cf7c57f44bead28394e46b6cb9635039e336dfd360b907ab557d180556da09e662aefdebb
zc7cf7cdcd30bdfbb903ce1781d3396565424f8859f16bc675d369fa2c42b7a906cd72918a95599
z26975b2062a8db18ce1d48358ff16294bcb4239eeb55bdd7998c87fa5f909b2fcd5baf6ff818f7
zc91864f3b12f4b7dc95fed7aca1790572668621ee1c335c95fe2d4c2ae6dcaf654396ac16f1098
z65ffa1af5875d40feda5bf25ba07a8efb112dc8ed278dd7cb2780e4dbb81dc87cd7f3b383aae9c
z8f2278eb602e32261ef88fbcbda73db6cd4a8b491af28fbb00e1afb426d63b69cc545fea03caeb
z265061823d23d360aefe45e8ddcc753b163f720720be21abe6fb5ada5c7148474b24fb71c29235
z9741a3e64d44fc112ee9d8abbaed2413d940c6693b6da7ee6e6953825f52e29fb8b7293f36ba3f
z0e87de527304a610d035701b8b18c8263132ff835d020ac58d0fc11c4189d4645874105b8fb375
z51a714498e10fc301a134bb93ee0dfbc765d56f7c35cb41070e8429b434dbacee717e6a07305dd
zb7d1ba72de8244293128a29c8172ff909d41504a5dd76506b222166994fa01d366a42a89f496a8
z36623fb62b9db9a4069271bfa7581773d8c2e55f26533fe72c12532244e0927efc7b62cbe31f35
z8d0b9379423069584b63ae9da952dbcb766ad373bdcbbfd9a3be9271198dc950d94548e4bea5bb
z60a99758655e283e9926a7d466bdbb6f14610a948ffdbb9650f12698781d4da120e4de560b8813
z6a5107fa29b52665e42c6c36d7714a9f61f21bcea05b71d5a6daad90f33e2017d6befc90bca2dc
z3636f67f0f0c1420248497144fcf9bc312e9155b6b52f05382105baf8a81c317629521a6f9a1b2
z21d920e8ca256aece7eb423825aef1d8797ac7c069e519a6cc5ce5be45cf92d491ef7c4db6eb69
z1e3c56bdbd2a64da11c375bb4f9302e7153714bbdb79a1e7dea11b11da60c9ba727f267a5b1822
z910c8c8ca631c815d9a6ef663633bc417407f2c74cc32fdbbaea1c1e6e60a0049d02004895d08f
zbae9a581f9d7c4517f4656930ef31917ed88cfffae62b7cc56e6d35673b25402a6a340d75c8bd1
z68c65c4827fde314406ba6d06d3a71892cf628a6bdd9573c144db39e6d2f0c3b422a556f967573
ze99fe7b07c5df78a97246482c0fd942141e9f2c201cb65c1ea5c610a02514c2c90f4856bf2626c
z930671f1f6fabb605dcca0ad86a5eb9544c60d18d967e25810a5216f5fc9a2d9d79ee6b0d169e5
z4181d6c1491f8959066bbf4f2981b978dd6cfe78a4b2110b00161633538e15a443154bf4fd9a78
za176aeae87271f84f2efa3e5ac6d8d48b3bb607e7750c06ec948802a957d00a93b53b23c728720
z7aebd5da7a8a24231496447f3d4ee16655b565c37d7fe014481e9e349dbaff70dc6509695f356c
za5f4e1177a54014bbb02e3723922754ac5e39df1d3d298707d5f8bd01ee641401c2c4991714124
zdf2ba637d147a000a436313ff651edb6a6c60d1ee8df24238f187592e1438e7ec3802cd8fff321
z1b220994d9aa492ba90bb315222c285dd8bfe27c0e686c09ebb712762bba0112b62adaccf118c8
z6848496e55f6f2a9d5d3752aadf2e40c23bc3d613bccb61b49b9e004308a39a08e0cf3ad0c70a9
za3daffee6947df70b6b64b8dc2fa31c6b5aa3d3eb18c1e5f68defe2b7ce4dd6914f2a1032f1811
z8a1556be967f39d38085b6cafe58408cd18957f0c1ef0ae674345a3b6f2b296d81d6b2d85497e8
zc1f71b53ffac864d5a962a0771d30f4b033a1bbba1a7c5ad1196d9563b2117a75680db69c85c7b
z817ad7d6563ed3ca9b2445359cb14bbcc408bc10a3562a13a292395f483febad662c0a6d11acce
zecea963aa05508498b65abedc64242524beaa6674e574e69b2328f73eb20f792f95fa9a5bc0db1
zbf39f0538b29a575ee36fce542191a5964c8db0949ba384d35f4b5294c838928a87fe23dac9c8e
z56138e340a3a631a79930eaef8089d65353ee897b1dfa39a4a4e755a6aaaa2a192565561d836ba
za0b6940863b719543f343eeafa31b62ee4597b31ac8bb8f5b72681967f0f4c1dce52a014b02f3b
ze5abf7db5a09ce00fc59757d5fa3dfbeae05d708b33030fb1bfc4966b34fd3b5ae625ce8096751
zdf9ac009f6ff82b0dcb76a73a59c8b0ba9bfe1e941690f2d760cee715f9141ff0469bb7c1fa40d
zdaf75c971f93f4b020f7d53bb5f720c2d7c77b4c2dfd0b44b23461669653cf20e4511f087ff27f
zd1335c6ba03ef894bc5c5c346435056f604a9299dfe2016bc373054663c9d61d14e13083d3b526
z9cf3fd416f6159c4bbf6ff2fb3faa5420dd3d6eea8bdaebf081d90522d64ac8a69be79d62bf894
zb54ad49a56e3b85abbc0e3db0fafb3099ed75cc1897c8a81af6c2c36b16d995ad4b0ec34cc6bbf
zbccc90688ee8032beb218a7ca089da2985963cd178bedba8021cee488d9bd702d726b7fa9b9e77
z3c3fb9b1d5d832e5af118abf67e25c6261cebcfcf983419cf376f12174666fdf308a14e532f316
z23e5bfbbbc21de28d716abb4e583405c7fe82167f06936e4d10e8aca22c75581b5b6ecf7ff4118
zb3b4fc5bfd140971d24dce6f703cb2b1344f1725298e452d9b29b0c4a0c12ce5618576b13da203
zcdc099aa46ec282bb8aed032f14fe44a18927a7714f5e07b3c725a559ad658f06ecdc5e6e0e884
zc43410d8930a53efc547fa6621ab8c8e97c19f7c3760a4bfc6c578fe7829b26406746dbb95c857
z04bfab9ef5d583ca4fee27a2bc47ede2bc951a29c2689518c54a48a4275092264a7a10b13b3f42
zec8068b7a9eb8f71f13b17bc883b1f548b1648583abeb1262804585af33322172e5e7357185ede
ze39f57faa70813fc7ce03b490caef6a8c11f0dde54f30f4127978dc419bcc0df096e9a0f7c6f0a
z2f946d46f7e660a91b1005cc59d1a874cc31bb0d31bc176bd0e722ce0c2ff071147445e1ef16a0
z817eed94a2ef17e8b441d6d97edb18618e42694d50cdc5d896f2d725160669b336919cc0ea614f
zbc8407ee3a298b95f6149626c47abd0ae6a55d1ab67b362f1ee44f58bf47e34508f9e6df089fd1
z10ae6e1bb1445d09226bd1633210da7606affd267318c7810c04558979ac5feb3c22cfb0d90a93
z1a80ec996254fc875e7d82d7f0dd1a1b1f2f8b80a6fa92880dff51ca07130c3c83d2ec177148bf
zada849e9a4e0cc05fcfbe5a2798c08ebed0f1613263108d3dc4106bc19a3033b15992e61e6fff2
z8fcc3c87d1e6286a014a4b90a04f11ead479ed9b3474594566870c01a2dcd61041a3658b86b165
z590df50b42250e5a244be5b75479b979d2b78a128ab7fa87ca2a7faf75e03b8392b32279f44af5
ze9584e940af314bca5a3902ced15b3ae4c9fb23fb85fd3950cc8321c2e88c3d04f08e84530c6c9
ze1eb9f14dcf398e0a70044a6168dee9b281c199fa85a59b5e2f737ac7c60f6b00427a28897fd69
z72280151d72a81c203b1d7bf7badcc563f7171b3cef090a68fd4b7a8f28e6bc24c7ea38d63ae19
z9039993d9fc02504f3fe1c73f00a1c2df03d7b208bb6f4d1aa0d2bac20c2e30999f5724c7d6c28
z11a71e086518fde21dbaca4b412db33088ef12ff11401b5584c4b98fd03614fa1c6e9543c54b35
za245b61aefd848ed5fe9fe14d0df53e9e3dafd602a70e4f9c401f0bbc2936bb57268ddd5cdc28c
zbd7072e991e10598d81288401ed2c8abecd42f5ea32ae13c3fb30ac30f2c213d0c3277eef252b4
zb17b1217d77d9c0037dbe8b8cafb20b77eb27005b891f56e0fbadd98fad8d50890ecd0109bbacb
z1b750da37bdf1d036aa119961b27d1ea3eb7fceae7e5d34bf04060ee13bbf0d2c8344b0061acf8
z81ee2b7510fca075a81e132f85c73426d42d972eef2c666ec3828fe36457242afe4e2c4757bd96
zc949a376e7f4905adfc7cbf79984d5268a66dec0c6e2ec932a2a940787b485487a1813f0012d1f
z5b3a009d29284f8eef070e46889a438a09e85c04d6d15ded5c082b00d840081215926f9f429926
za1c68a0ddfc48e9fbea825ab0f20e0058e1a123e5e78f47e173dd3b574307d00c61d4cdde81be4
z704f72fa8bcd02f90ab444cfd4826dd2c2935af7f9977a9bedb6e8249fc2758ec173adf0afc7f1
ze4d57d3f5dae4243a994139ba66085dcbed3b52dfe44e4b5d8b28c1295f6f4ad1cfafe640fb32e
z9bbd438f7e92c56b96e564f5c68af514e58a8cff0be23adee54513d71a79061682d42060c30fc8
z661f53a75fd50eb6ba023b23c62fa507da67e480bb97e74b2691a0bb08f167d505afa2ca0ff1a3
z9984caa22b0c3ea9e15510a716c026699dbb2f81eb33b483e39eb323f075ffd914534c802a5b92
z7ded1d5c7d5e666d81639347e6ce18b6a83e2f3cd418310f78d38d8bffef80beee710cbafc2e81
z8f8fe88913b22819c00df2302a96fdd14888a70ac544f470991c33333d7e1a9969f16493c42d34
z70f6a4e9b35db4a2974da0227ff54a4cd7433c2ad59d9bbd4b3ae233f0974fa89ac94ca3397273
zcacd90977b87db6843de0a7e2b551d3936d8bfa897469eaeb0f3fb68774a822e76244d935d624c
ze3cbd3475ce7ce22faa733717c0c2ad1ba0ec732734ba55adf4f7477772bfe22a186e570ef95e7
zb4a98fac96aed88cdffc17a1988d2c19bdc69d8397073f3118ead4e0e7a56070274a63ad0d2186
zf4d3086bebe44f55ad966b2c17f4eb149a2d64005152050258fd8aebff17e6e170ad1db9e2d7b6
z601e522a4bdba8a9923560d96f468f8c62245f46b83f04a6e0e386762c1f50f1d8831588b258b5
z348e80144a110b1f1e26a1c87e37f7ce02ce53bbbae19522a68573a233ca65851939acc4ee1c7c
ze4f80800bd567cc740a1a289440d4f3c8fe7969384d348a9bd4ae02df50b2f0dd438e48c3f07c9
z2af58ee58db38ac3e7d56af52cb3e6c085bcf43667fed738864be36a075eb93959f4988dd16c30
z5fcad1d6aad2283576b54323e0c261c3c8ee4ee69e1aa61d76f681354c4bd369b786fe188b9dfe
z4df612953f3dc24f75695364d49eda5ff71d28877f851196923743456299e869be2bbed1b54f71
z958ea5d48b880c8c48c84c43a79ba5ece1f30143b6b747e80311656ffb5e700be1d9767378faeb
z45a735a04d391fd066772b0bdb6f384cc1b67541c52a6491684ffcae81a5229f0549797022f08e
z51404df33764cd60302700ea6f44cb59488dc8c5d86f857358c1cc0bd86033991d65a510dd34ec
zf68931c1473729444dd6bcbd77f11827136428569bcb33dc50175eee548302cdeea88471e9f04c
z6c97b483efca681d79b5c93bfa7284045d92bd727da620d311fbeaf6935e5ea1873fe7ed9638e2
z05e1fc1ed10b5ceffe39c1c997b0c348ae832ae2ceaeac22c8c0d14451820fcae18e37cbae268b
zf5c2326153ddf854383b079b6b3c038fe4a41dc312920fd0bbd3ac13b9e85918538184604f7193
zfc4a2b58ee6a16301657f965bd2fde1ac22df9c410a8310f7abf3ed9c64bc737a1ffe2d38c9f5a
z01cbb6b92a13d95dec4cf75d11dd51b88c716a8149455d5021cdea0dee750253e885e3780db41f
z0e3e2f50f034dbfb557ec5c59a71e2cc652fb2bde26f6ff8e99b9898ce0f0c1b36d7b71922ab97
zd04e08e9e96db87474db62f67b6cc8af8dcc3d08712369e899a93309b03c61b53a8bf241f20742
z321e071fc34831c83b49f9918046d87104d27e1ac74b2dbd87eaaff835067d6e847624a8252462
zc3c25b0abe6d09d6631672f4cb04f463e863251fa9a2c0a267025be3e7da3cbbb782f798d2a714
zad03f2b894ce26ef2b2a494af86f9abfba185f5552172c7a09890abad70a4bd806cbfa9a305d6b
zabd98498e5e44828da0fa00e2dd5374a860b31838a0b7fdd3a4274b41a82254061791e64116c3b
za64199de9cde1e1e99a818a96a5ca151e608f946629597b21736061864b14dd0cff19cb2f366f6
zfe8a25f9a4d643d79f0e0e64525c92ffdc0c042ba81bafdbf201f8b2734fa029ab1dbd7d2ebb0b
ze20f18d4fa12b6b7e43dd1fa12aceef0dcb0c8264d8e2ff76ced234b4473e534135051e6e7753a
zb2e8bb288b4908336cf766df96663b9ca715ee1f9c07bcc9949b2f0c53b314dc0f3ab74aa7765f
zf4c403f0af31b1575a78b56f33310875fb14ed1ce9c76ceea1aaaa32c8d42397c00b60e9bde77e
z7a66172a9c66dfabba8b9dabbdd69dbf0c42f8d9133c9dbb8a919ab551cd3d2d14b46902de7973
zabeab0cf1b7e3ef5825fff6c44dcb8e4a32f131e349934dfe83ee9c01a78be68d74a0269c687c0
z75a638b57dbd571078cfd4877d4027b0864c5181a988ceb257a6ac58ff494a3ee0b7c2bb21e03f
z382283f6234f6fd2c4e120f0d23292ad027b5e96e8bbc2d883af0572beb6ad4d3cb5ba8791c681
z9bcb463c4c176272a1cdb85b28ac83a0e2b2d3a3793f12bec8a52949ea4a744edcf359339f271a
z00cdd03b3f505148b61c9e6fd811d98cc5bbede3cd25f09be5803ddcbb7f53f6f33d90c7471339
zf895b8b8bfc76fcd5e2c7780e71462fdd56d32e2dbebdc8e1804424e29e24ef83f22a5939ac757
za13720d5c37a740fc8f00c4837da971f2c5b64b1590b66cdf68ad4801aec0e3b778d6b38933065
z362fad60d01042e48b976c15d52ea2f51d18f1963f6255d80c4f8fc61984bfe8f86543f85c3bfb
z67eacfc77c177305fd23f6f77e4b1646465e4652e36bb7dad457e0b3d07a66d85276f987ac8a6a
z985fd4789fcadbdcd2a114f5bd1a704c745291c2bfceca406f4c7b0afe6e755d07615289e7793f
zdfe552c58a3b02cbeb9a91f1974fb7efb7aac9b7f04ed2e6cff713aaba4f2373899125046c68d7
ze6874cfac7845d537d4781b9204b4d0c36715aee2f0cd6ca0e7b05449371d8fa72ba14b2bd2eed
z8ff4114f1a2746ef961ea5dd9ce307aace5f49457d3d2cca788d59b12dc34f45321108e9020ba6
z7c1e733673e467d5203cdf3c928484fdb12e51098b677fa654be41e5d1928eb26852e30aeb1ebf
ze76c6affc4694795b4f5e80350139c7adb8f3553bd2cee9027566f02cf89650ec2a5928a5afea6
zd802d75f08c442a0eb6afc3d2a8d5efcec985e4337848dc436b71b82bb3f480bbe1ed724b8c534
z24cbb53bd5082c81ba2ff5587195e28e7b9deccca4fc42cbe08c086b874574970338620b67fe24
z9d8b0706cc95dd6f8e49004acf471959ffb37847d98c24c381a38d7795f8bc9193d868a4c861b3
zcf1e75a43d8abb76752b84c368294948e8df55d0b411f8041e339c876968ae027be7ff565adbd1
z30cbfb7e1b37eda1a23590f5f540e2799ea67ff5309a1d1f53ad01e4c1bd87714a6ac22f92ebbf
zf7f6025bc149b4cf804b583a4ffead5e588e629615863064892ef4ede55016edafb97dea3b4a86
z4b2375626eecab8d1e4d9341aec7086a52d1982263f926daa905a60ac682bf58aad9d9ce4d4eab
zd10c00559c6def4b278f1df9aefd794b9e3ee27318f69c15c2f8595137849d2d2252555b0513de
zcf57e5d98717cbe2377dd7b7acd09515def2e9e86feda29ffbc69a949fe03522b51ba3892cbe06
z84f210b67cd6de3c8ee4322b928a40cc87330c9cc7fe702575b4166c61e8dc1528f3907ac97b45
z5392eb7a669f7b8bb8fac34cc79c936fce86432007be912713e63d09f1de8d819c429012016784
zfd0d7a9e767d56a9c281df705c2d604fa4da3fc083cb6321a563b575facbb0912b191147d3aabf
z5ac3b288783810b6ff9b2b6cc07313caa5763d5e6405187a4d6452c50fd34a03a946664c1be101
z7a10477b5756e7ed1de14ddedccbd692fecef94b11cb24046d67fcc60c63c1111b6b3fc5fc47a1
z22b1cfc0fc73ece38c46d987a4fd2d145c9362a40f5a56f36252d30142c263f3523d0d91ef26e2
z6a4367dca69f1b6788d8d73b6a487297255166cef49920febcae4b15d66f7187579e015d39ba61
z6a3356ea1098d7a9369b6ef99da29e2f6649a92163431c82d411aecf119596965e021cd038c55c
z0eba4759569fc12a176b0d4daf16b72f10dcaf2cc72dfb17952e9e8d698dbe58d48654abdf6c97
z53de563f4e04cc55367e8bf9548e8273b0c49472b95ac211fb3da18f0b88f8b4f92d81a5ea57e4
zfd5ba333a12cc2b4995b4e3714151d799cd97aadb7460a9176b49e722957cdfb2636759dfbaaa6
z3227e868005961769b7629bcecc1c9a11633aff5517b84151ddbb29c4130059aebafada778cf46
ze4ca05772849f1b8bb70da68242deab7ffd51038a9b1be7ef0b81c1af2c1a8708d8d5b5b75f89e
z3a60684a3bc359ef5021041d9c87494e96a16639095f81dfc6778567f2267e4a951cdb7e6da0bd
zfd849a1f72630aa8dc1e9e7f9fcbca88a07344965b56cef0cb6511754fa1aa54f2e92230101ad6
zfd3400efa2b453e7f94a0802689acb4221d412a4fe5cd6d0484503170f9edf7b66d8eb7834bb3d
zdec4245f9889e39676685f7405fa0c70b30c5a28f5ca6a010c984a280a5e4933355f74c534461d
zdc4e3085338c30e3ab50d9bf75f82657edaf75aaf3d23bfc4cfa3268dc87db2d9fb65615dd2869
ze2ebe9dae7a71262773938017695f8e3bc3f161af8dc1527f6c36ed6bfad13b1941fcfd423c8e4
zf58f3158e30c299aef4e477a3afc1a4bfc323d37ef0dda5865615103bc47a5dce5f38aed6fdc3c
z93371e04dff8f9326c12dc435772de8824e85fbf82b2659d099a490223f366cfaf035469632250
z7d693908ff932e1f21998a9807f3394d9308f74a0f8adb9af442f324487c2e5c8224440acb3d72
z0661b5db3ed84323fb9fb8509dcf420d57371d53e51a8ce422832beacfc922f61f0fa2ae1d328a
zdf582ec97381a1cbeb1a4847087a649acfa1a779d175033ed1ce3dd698bc1b01c14f5e57109509
ze9089ade6b239da75c5be799530d77fcbf2859d63470c4eb789de56e2ecacff371e30442d675f9
z5ecc4a88d1a14b42d0c98b86861a5371b82a598512fcb290957c5936fff1b821cbe0fbe39ed2c3
z0d4d02ecb58dc2daa81d4e3398c764d3b8e4a5c5847ff1c10568fa206d38364dbfa2c6cbf7d3b9
zf4f44e3b4f33ebb8d2237ce205bf80d30688b69bc7d248729b8ce060bf724e79afbca90cd1d06d
zf4341583a434bddb2dc91dc56f61787d1227bea1095509f3b72ebf55fd201b53c7d1c03c1da6b8
z184e757933b1ec3cbc05cfd6be9233c4b3376931b5aa76dba726a5f5c5aff8586d2c3e750af903
z6cca5147a3582d9e83bee17418dd443706c44f0dd2fbfa1738cfe1c30bbb798976c533a6f88822
zf163b97b83669665513d35e8030d82ccb3b1103cb965fdbdeb9a27c67e0b5ffaca16dc78dab804
z48993db56a62fadba6f523af2e44ea7825e4ffcdd93756ae394b176753d6ace7860d5826d4dd40
z13ff84c54ec77939aea4953babbc9fd569f0711e22541c7f04664c9853f5869685cc49ced76a28
z9f0dc088d26bd75c7d77ea527b9fddf23b7a06f903e56f3b53ae23ffc0bfcce0a597a48a1d6a22
z92c7c6cc52d6ea7d8ccee4611cddea47fa5d8c5f6906887647c4cc7357799b1b6b14bdbac90591
zf1a8aff7211733ab91de49430c1088c37d9e2bc360713b43f5a2021a250ddfa3b82e638bfdc6c4
zab2a7220f291f58b5a0129399fc5ce91266d14d79ff2bdd1bac68f42f5f931ce9143876433109f
z9405e50ebfee3a951b0334d57a6fd7753f5263fe8858fb47acb91ee4dd31670d738aa6accefb36
z44d1f70473894f541d284d791591b87325b4635ef794331291f8af54c9c2933533ca74287cef70
z455107a3893fbff507874da4d7b87aa0c60733d8a60e2a441244b01eddf4441da0ba434bbdc232
z3307fb42cd4294028b8d12934c8240ae74f57b3a6acdbf15411e46822e661d917f6c4a20912578
z0842f1f234d223e134609767324a17e30222d3aafb910354ef069c5d2cbbc00fc48c46e8fc4d46
z3aaba37d6a9d7c0468207c12de2bfabac04022f618932d97662031849f11d72a9d1fa0b434effb
z2e432244e046b6c3f1f063cc4cfbdd305af0c812ee608ea2e0adf007a40ea1be31f564e033a659
z22fc5cb843880d67080a20c747fda6cefdc810bfc266c1f06f39577deed59da05f63d3e2bda534
z4171c8bbb4fc4a9a80053b873a447aa5e08f7a174fda49c03df641af651f3d1767fdc4e9cd49b7
z0eb80286afc492788cfda5c1cbe55e9ec98ac5729ba3922bdbf3e6fbb86ef647e2f7c0e4d430b8
zf4cb90719896761f39537ce332d01eeefb2e5975f9a18f76d8a4559dd68353a7d24660c003a65d
zbebe4a543d36b8648364c92dff9657cd69fe446eb575f56b59773bdcc57c1832b4ad7fe549b982
za4196b5444abd017cd7b5cf0a46fb7ef0f5260380da6336d20c11263570a955464e6d9883b627f
zaa7c9bbd6f6ebf0d9a47bd2e3faf407a6f7bf8c2e53ca873c068baf9b6929161658c8b59a93367
zc91ab43a688704d2e5a14658fb707406f6c44e56da4dc16119db489eeef837bec509f510566646
z783167c7ad160ced8c3e95d444955f4c77085b6cf549aba5a7345462a7d9c027f83071182ffdfd
z06a9277cfe8b772ae0ee3b092d107dac1600afb0afa124d5ee3f9835ad5bbf540254e80cdf9b1b
ze8cade951c9fb1b8cc1e121ff374d5310cf415b41ec4d7e36771989d9b67713ac134732cad6981
z5fbd755be086cf3db025ef72ccd1474ec058eff5e704d0c3d59394e3f61d58bc8fe267066e06b8
zade10966163d3906052328ee6549fb074efb092925e6e4bdc5de37868c89d31c62010e0d5918aa
zd7f5b2e2d295f0d271213ec95d22306791b661170c7c5c68248d1c344cd14dd99e5b1f12d2da72
z7cc0116177e10c8837d540b1a442871fcd9ed54006355e9ed5a040017e0da8603592d975717e6e
z110123c271ca4ba9df44a49f60903b12f622da448b6c05ea5541aa901c587d6f6054110dd06a6a
zf92789bcc5905b59ab719d6b721d0bcff3fe1cf839527ab5a46cb561880ed3b62d3eaf1e29162e
za0b1943ef4a7e5f0086dcdc2b9a0f7ec1536a610d9e56f535ce0430a67fff48f87ff50bda0e22d
z7f2c42e2a4c0cf38b4eb77a4e577fbdd8015ce1cd587bf20f4e62206de2d8e3e4c9c7df2928529
z3d2884a7556e0f3df0b53fa4c50d4d2e65dadfae7f80c51bf06c3271737b6b18a064f4baf5f492
z0efcdfce30625246c60924105d7235d58a5664a897416ff21410d7cbe6404442744cc1835c6a31
zce3961729e5626238df102fcc16aadfd7a5866274bf9ed9cdeb7a62276a1bc20933a6ca548344f
z1c3e98934b481d1437459b9c9ac615344a180c99156b30840cd36bc9ff595a4edea8b50265839a
zd202568f5cd03dc55d0a124a6204cad64ab2db8389a057700446de11d5cc5c2360ee99fd86ddb5
zbaa29f0da19d4271dc0133ec29904c50a6b707fd51958670b01147e75f156feb62c256752143dd
z0552ad181f1f8482fa5f801dc3896617efa5353af21f4d7af932bf346c6b67f1b43a0d0c0ba62c
z7358dce61dc6b973e5484e79e9588846f454dc74d021886c890bdd8baaf6c6e9baaf3bc4fef0f6
zf612cda3f33ba92a9e7a40bcf137293befdd37c5288c0705183e31f146a792141359c609dfbe53
z1ed2935c15ad36a84e219f4988c9dcfeb1a3938f625975e9a680a4a41ea5d9a261860f725c4ec6
z30d5178d4c2e46a3a390bba9e3a10cd8ad686f59ed7d8320c5127e1661579b8549d640f583f6f4
z5e50c59ca40123d11677585fa839213b0ed897c366fbd6f1d209974e90e8cd0bb2f78e9320bae7
zd08071d2d37814c2ace626b89a22bcb8a4d165884045568ed075c9cc38af93680fd25001ec2ce5
zd62fe6a149c6bce1353acce5a3132c6d2b1e1771d6d38e13d9412a0ebc046e6c4b87e58ad7d25a
zbb5af773e4959aef7ff4bb95152b198d4e03333d29a3cd300eec04105002c64b20340d5983049d
zc36c5cc82c10ab1da78ad46a08bbcfc3419976147a0d07cc9c2a3a00807f20019d3e24bc988872
zb50bc5f5e2fbb805a87e3a6a22d9c70586296cdf03c12dcfb6f6a5bc001cb7cca8c548dd450500
zc7d82d0c0102f92b4126fd0e4a5d17d78613f91a4d162371170ea98c83dc38417dd29e66db46c9
z600326b226ccb03b868851e6313315210d602787cedc11a457e85533adef82536e2ac2b72e2414
zf5e2157fcf036f6b282974108ba0376faadf35e333b65c24dab5542a2a9c649466d866a16e07a7
za1b42ab226e7d28716028006bd4228f40550d160623b55871f3064395e3e89a381b1fc0e7a16a1
z6e621160cfc14f97d8ab816ba230cf3a237a5249cf01398fc99bf69839ef8e16294715a173f8ea
z8b34b1539cb4ede1cba7c904d4e0f4061a7681e355f88d60fd145c0efb6c872352c130c85247e2
z8d0e540cac71467c3a374ca0f19a9c04a45a2edb64fe2895c510454b60adee90852c8743812439
z19870d189a4a870b6228d2f571e0dbdd24baa78d35f198393e9d6e3561a379f30c8abb68b7c96a
zf3775b866da8710f6a5246b5b619ba998a7d973235760ca4afc814f1ae237174821985ff815309
z11464e26fbffff0b40a2e2e0f96d513dde3dc7088daeaced5c43a7d1a5d299704e0919e0c5e1aa
zf25d9b50bba0b4ff07fb9cab00f82087c5244f3e72ad0c0a685c092d0f329e066f259f524f7af1
z18806639557eb1e7230c8e2fc7a83264f07e78d759ca76c0756c6ff5958cbeffdf0cfaf57f68c9
zc4030a1a4367e55d349b02f077d7daf86576c7acc2170231a86b77926254724180b9a3c7175f27
z19c6ed704cc39e616de23fb2290b31ea0b8c0e83d117c42505ef899885fd29255570a3f894efe8
z9d446d0858caf7badadfe5b2bc3b84f995b4bf5de17e6f61f3a9229a0d9523ffdbb2c81c7352b2
z777eec3ee986058762d6e7d0294b0740710fdc578db6966fbc02ab9ff2453735eca164f86fc1ec
z8fff8c565dd2855af11c46aa2cd14a774dea16c1daec43b4b8d68872a7d6a08fb2287697402f0d
zb3454f614aadecda73f57e1989c2d1a525e265b23da047156f1a5a402c4fee822f2aff31750388
z338234dbfb562ca59376a122dbeb3d51ac908fb8063790e8e192bd369514063d0f985fb44d0fd5
ze414460bad925532e090d59e1f79235b019b009e8ae892fd09c5c10eab74c0972ecd3b33fcac7e
zfc78c15e7891f8f70686f58e3bf914e4e0b7059cb9f44195792c6e0edc414cde5c607fb953f2cc
zae7952b3aec6bb837eb4130320e371f6341e57a7fa326b0e457fef7ea335d39fa973d536e54821
z8d72cece5d6f01b8885b75391f6ea806ec8054f9ded784822eedc3f4276c0caea2f1e43242bf12
z2fc59a9c1f9e4ae5738e65aada55811801779665cd0b3975ffcb5789ebf65954f4c2abc821d4d2
z7738a3909826a3a6223c24e36f9d4643aa5e9a9455eb22df86ff605a7cbbc176de5d0edaadb8b3
z407b4d54364b779898a303ee32b70059c1e0261614bf9951af77c21815a99627338bb8b0805401
z0e1ed9052c92a5606beb5db3e0661f328d0d234fa21c79b8c9419b759bf7cca498b6497d3b29cd
ze1738978539b711003f36681b5b1d292344644035b49bb68b489aeb5cbc84a73ab4629ddb57e41
zbb450dd0769796a2bb178ed1f7941f1715ef91e901a4a21f60e0a6682c0d1e567c9a42fdda2e7c
z7bd086a252c436741b7bcc39ac07f08e3d399c12b88b9bda8aaa579aa7f905911cf3a0c6f17974
z915c9107c3cd7442aa4c44b9245dfa267fb6bd4cbc1e32d6a05f826a7503a1d43eb00e64dcedde
z9f111da61d5a8a68f254bb1a1bfb0d0e5cce31c1320f4ee1d43a776659a4fcda67f2ce6142bc2b
z21f024fbe602d996103dd2e6ca4dd26bc3182fd575ce1bbbd3756b452ea23f22baf002e5075cfa
z27ef351b60c9b08593d59518ac9bbe32c7f78f0eaa8332b7bb689480964ea223943c9110f2e36b
z5ba31c99c156b5a4db0e4ece41f9a7595d429ff91b93b1c4c244455ed837ce28f6d33c341f0911
z45a216b44af694c0c45bb37c7e7d3d331841d0b73fe64217a591a495a0287874934e7f513e805f
z6112226e1af86716ff2a5708111171c36a86575147eca3bdb75276ae2ab7aecacdde23b6993d9e
z49712e580178e4e24dddc4991672dd23df4a1f30b2c09b48e196f4caec1c0259ff16806b5ac442
z91b44901b50511039940b19b26e50013829d8d7ca0f2187e87454b59e54378f9a91cdb4e4f28f3
zb8d05cb4aef202b917342863493769b1a4aefc9a8b937baee41e71c6680be627225c3ed0fc905c
z9d446473a7c886a32c98a09357222b15417a2fea124e4701adb3879b584cf45be98a91160ef7a4
z6a4dd97aed125aee2215a64ef48bd6fea54bbce206ebb03bde90203b85790a25612683cf004649
z2e3baa5ac1c722a2db9e3dad87bd9209e8f326819f9217c33b46bb5774d7686ce27b68b6af3326
zfd329020f9bcbf3281b32bc048e4670073ee28b304a8861585160873f6b04b9c604501431cc6b3
z16512f1796f9e459f55d5453492154b05b957c72fc928d69cfb055edc98cccc8880fc548ce2bdb
zefccc58059739b4902ef47731ad840e03f9b9656a4e848e0f1ccc382be98a5596f362a11efba0c
z57e6ba41f4c87f27804efc0f49e7868d8fc5309afc3455e8afd3a0e7c41cca0af808eb45d306dd
z82ea31a29222d2e819ef9d2d2ca0e217dd76ed1cdb9bee49e0631011cd04d148ea6b82d32d17e1
zbadbbd822ef31bf3029f107561404a44d42ae3de12b559d2f63df89bd6ca10f382a7303d019a81
z616de10847c14187c3186a2e0d05c79d005ec05b424de0df9539faa356f1057500ccbc94a22e17
z1c632072a12c925d368c96993073c11385b8140aae805f37cda645c7b17e2a4ee9038986459123
zd320affa6d400332d9dc1b68a080fb9bc971c12241f49796992377108b7f68525487ddee3c9566
z5b9097dae5dbab0a188c639ffac5c83a9992f19fe859646ac5a8838fa1398e70ecbecbd6e216a1
z0d7d45b4e371014786e12b1384fe61d304bf9678838310177f1d33d41df8fcd88ac8feeb6ee3b0
z5d6449a152cf278199112b7044524ab3872934a209c4aa9d2e9e9f970d4753f2a8c0b07c235a39
z3d0f9d3037974bf4a212908172458038a18da02cc0d869acd3313b347e780a6849a14b359b5595
ze66fd24085ceaea12466f118f67a53e7e71f7bb69da881dd88e5267f430f64041b4910d2e39760
zec96780a0fc11f23a9c17c4a23af9cd70ea00a309909a3a3d8e699882e9e4c26f67b237ee44385
z64ade325258395e7b41cc9ea99ac0a4c98254e357c5b86a8b6f5711e830bd28d353f82f8a44cf3
z03c387dff1f18272d86dbe55951faf9d5f7b3fca372ab0e3f92b3137e4f0337772c981b6d59680
z64348775525dd361ed24d665fea30e6aac6da401c72ed1f32afbd7bcf809bdae23fb5a5847a869
z477e859a58bef8ff4f57733605fd9223b8781968c59c27c8ccc64397768f8bd41944ccc1001e8b
z429dfb708530c8c34e5cc9f4e2d0d2ae6f67a03df15c3f9659c4717d0a54ca6a5227d58f451c2e
zb6644a3c9591c345da75d9fed9e3751f1a84b9ec9d09548fa10af3e635571c6b22d58d920eb973
z09980c3468d758a0075086659b2c2b87f60c42d23164abf7cf9542db5ce505e521a55af3f61fef
z95e86ec229b2d45b171538d39958a3d00ea2c527b194cbfe905f602ee9060a2583edaa03cbbe0b
z3481938052f0f73f8041aadfcb569b41ad4f9799350c5c57038bdf294e93602fbafa15bb6598d3
zdfbd1bad9460ca210f878ff466551e41806bca0ff1032851e6db9e8009e607a12500cdaa8d218d
zf0f54e86fbeddaac589dc2de9d6699a3adbad077013b1de2506c586196e246cbb5bc783687d102
z20f9d52415eeb39c2920fb20cf80ed7ab6cd6772fd098df5a4d9feb4575bd1f857b1f127bec660
zba8c143df945e2df6e309e40e31b5969b97016df70312119f366917816e30e7539574f874bc358
z1d4af04a6fdced746c27b8cb615e11c0bdf7b8509e4f7f489951f70ca454eaf64662d06725a623
z6cb7875084192db00bb356d4d9320ccbc85112c631cefae68203d366843851b0a0bd806f66821f
z247dd363727cbd1754cac46c091e778b154d1679d5f1550ff0647e03ffe04278895f51f9c37f21
z1ee0d78c216bd39dbb4995807784df65fe778089f8e39f87d8fc88818e6bb683e79969f7389db8
zc31bc096937e39b7b0df38ff42d987c58034550b23f34c98bdbf0502dc7217a4a4dc8d529ca562
z559185f3e7332ef169b87b8f2abdf908d28a76ae7f17929436d6c2e5fabd27c6b8d81098824a26
z3cab9bb44f521aa8085c901c2d8fa3fa4371b096bfba6b4bfbfdf180d9a7c1ebc81934f49e8ddd
z9f9a132c2a4b2442ab00557cda3015488905c5fa0430eccdff4dfd20458446a97a76e1da0bf044
z024de208683bec8d31c2e25fae05445d51accde2dfd190b670368972e85d9b7f28da896ba3941c
z185f4ad04f9516b562b65b826cf16561fba3a30d7f44fdfae9752f0a3054deaa8eed1d55eaf3e5
z127531b07d4ee24dd5c1954fb10ad6ac8fbf87b5b62df98713aad881a3edc1347117aaa20314ed
zc1f308548274498e71aad9c00c5f42731a5986b7713e9dd13090aff875e8ef5cb2a203b5ce09ac
z4603c10c32c2164c1a5a8ab924c042e181fd369df748c559274e9ec5c6093f5c972c71e13fe061
ze7c1d4710e876188ec7f55950afad573a92d006e214f574e3872d49f301ddeac78ec828b7e377f
z9f4c061c01821a11bc84e4fe20b23e4b678d3cbac4991c133b634afae9d427cbefb21f3f933399
za07acc2bebc9da28ba4851281d884a59e246f44f722cbf65c56e934867bcac43ccfd23412b71b6
zae6521f97c4c1859c4c1756860892a9fd8c588ead1cf6ddb53bc3336cbd387822acc8d22da8a9c
z7de1da5863f25eb191aece547f911f0ecbe7dc96a399676c106225a9a1875fecd836d28c36037f
z26c88ad0fd64b70a83e4b6e51625c55ac2d60d75be19cd8ade195734c07e9f359001306e502826
za2fe2eaf7226ab82268e95bb50c34dce19a9a91f2481b738e7d9068a440619a2ffac44887334a9
z823fa216f08dbc333fbf9fb16cc6e9af92116fdc913604bf0ecc5b6442bd5e2151c625987f0e5d
z8d1866673a89a103c0aeb167ba2e14dd1c89a20eacfb8fbb3714ad26f09dd50e03b47b9b1d5a95
zb9f7fd19a38944e6668e5caa5743318d145aa8e7179157ead1dcbbdbcb100643c55a070ff73442
ze20d4e6bf932c248123c4b9b59f8913099e3655b806b90816687b36a3dc7886d9e281c3819a950
ze8182108dc347542437779de57f00aa56c19bea93ff940799f8fc6a585fe24ac864924eec56b2a
za6315cb3ffca5f652cae3d11dc4c9c5f129c103cc02918d895cb7140dda0c44ab4af9a6c0f59f8
zb0afb0e341033d37a40e74e53b4e2e59ba83307bcc9b101bf5a2f3b394df922ab243009c76b02a
z4cdde22ed7a4658b839602c667de0736a6b038b09216f5cc4d81feff47424001cf2ce95d782dfb
ze5cb52456e923f340b41c1987ef8cc52f359ff11a9a2da451263856a6b99ab5bc307b9434c434a
z395a4ce31a12ebe937f711f2959705a7d761b575905f266059b95ff1e68ff5f8fbf5859fef1490
zc87b6a4c90fd6352e936a43a36b3f996ad1d10ab43b9d121d43ac231c236cb4129343889795159
z1697aee71dbb21cff65b5bdcca790037d09e34cf93c82e9ed6cd25a32dc3ee0e04b60199f5d846
z982a7abf24842e5b7c43729d0c497f343033aa0cc1f8831778f3c1da6630efc9a9c393d3f9d532
zf20a5b4261de07f2576c7dd899c615c603df56467bd0b88c5406c77a2e4f35a744c15aaaaca5e9
z71422c83ca16de8ba1823448aa0b59327c3bc400b6496297378e9e18a5dff423cf32812bbc5c05
z900fcc593c6ea0aca9e5a059252a3ccf872418cd5ab36040fe1b76bf974715b84b8de036d386bc
zd7d64219bc08bdd15e1ede526c592ddc413d6f8f79ba435d30bdc413ef54840161cccdcb45a891
z6095a9d0aa2ea10e617603fd97ff0ed8d81696ff94f1278264cf922417baeefa99a41a3163f89a
ze5a78dd4a94303856869cae455445d03d562ecab74c5a2b513c56b6db00bbe870c26458caa5c64
z991fdb603fbf13b294b32cf0ab4e1fb21cce29ad54e8a8f987307a7a8672a277eff0c53909359f
z7022cfdef20443f9bf8bf0ec903bdc91e2e1f5924c74440aace6d73749c07dfcc17d56eb26cf51
z45087c81af65a7473eefd87d3a16fe739c1148b734ef9e6e33a8a2ba6588349909fc0fb047d21c
z57e31c2c66c2d74e6636b6b728f7ab1b227ca69f429d6dc992c05b1e7052d69c62baf9fd4210fd
z2ee2fbf8f3d1a759fcd114992eaa060ab467b912c3a061cc6a24503ae58be746ebcaae5e1c7050
z767a9da64c853ef01a4ae5e3350633ea37bc5100182dd7303e54f1ea66295b2e3c153f2089b4cd
z6c6173846abc03e2efd23c6acd6224139cb9469d1463a02be5ce5ce24c856ee8a3f0964da3bf3b
z14da0ce9d8fe8c2e8a008d1537f96c7b28ea45ac683c853ac0142742261a97174c06a7dba6f509
z7b0974fc9214db1998432ce3491adacc6f563b482d03c72ac54e4cbe9dc45684cb61a0a4f87161
z9ee55a167a2e5762b30cbd97665d4d7c20c88fab405fa18ceefdb2d11b73896001613280b6a2ff
z4a13fc48ff997bfac9363a4e1dfa7e931e2d52824b4e38a88528f9914c9c4f12e1cebba34f97d4
zfd6fc5630f53742ca59eb72edcf887952e88ca87b2d4beaaf738853797d4db38a3636e2439e606
zf8537080123acee5d08147a05891a25f9a490db6d824493f0999396ae3abc31aaa906e869ae7b4
zd07e2c07f895adeffd25080f6665af0b28fec7708184c3dab835cf2e484504b137fc7f9a34e89c
zad94cf147c50ac2e5470e2c9abefcd7dde3de6fc2979fe4b3c44fb86870c9e0ff06898962a3f54
zea8e77abcec2ec816b173c7f23f8c313f7ad25867eee145e25dd1c7b25dcf0d69649edce17c91d
z7e160b3271192156c208bd4fc00adfac98dc3c4f4b5ddf30159156e7d94fa0c85e2e8e6cd81e1e
z347e796ee8cdfc1708c946d15be8da8b46651a49b4a384a8299bcd783efe59431fef4ba3fb273a
z64b9e99d380d62f175d0e3acbd04a9570c3e52d3dca238aaaad8962efb820cd6f3bd93eeb6ed03
zad8519ca1d7b8803ae4b4e8c72661e777168e415d657b5acceb29316f9cb02d9957d811ff07e21
z8a9bfc280e133aa1c401f962825830ea33567db186bbbe6ccde35aed8237e9becf607d8a83f28e
zbba9f1201752f758904a4aa2c34fcf4e8df112c7d8dd7c28c39e01be24247da403c048820633b2
z8a0ac6e17cf82ad4beac85d9ac82f6fa9b19d43181d4621e271b82d92783a3ca74c12b34ffa2d9
za2973818b04a9e4c198c9bdee83a412547aea860bdf7cc98c3e388679b30bd90ca74aef7a6765f
z91f278b495c288ff5822a786ea4c6e0236b1ab21794e25a18a116cd0b49d3e14c67fd78b4ee479
z05560e2022a75d63228ae8963cbba16eee66ba077c3adc4e54e3346bb598e1a552bb25ebd5dc33
z2898f0cbd6fb379e824817345b848f2e23cfd0def11e7bc76e7e4aa6b7c3dc7a46074c12e7339c
z50fa3bd9b7bb1173db4e9978feebd45596adc2098b8c215a158eeabb38207981be469b905b6b53
z9bb5f24d3ba1b9bfa61758ee98c9dc641cf8f71e4800a1ffba961ed035d77dc90eeeec180e1d2c
zc56ad1629a1f5e174ba6f6822b7d82e9b837b92a4edadecef2008f33e15b85d98635fc954d38ff
z2cd7176b1276844994f02b928165006fd067995988bd100d5ec888e5a70779f1632c3eac9ff935
z3ab9b7ab59738302ed31e0be6396c6f0147c9000a4c5d1368f3f45b4a98531a6193b067dd333f9
z69514c1f3d3687bd7baf2fc9be595e8576cdad52389febcf9000a105560b91135d1535801be346
zec1eaaab50038687f2b4fd50d3515b992e3534f5638c142d81f7edf8e6c96fdb34140111a709aa
z202bf2eb7cc3a0f90b2ea5b4c02bdf1e09cdc637db6ea599312e2ab306b73946ca9417adb59c36
z24e4768d4b60bc8b1426ab24ce378253aecd72612cd4ab90b52cf473ba15aa6ebae5877613f737
zdbc185b5931b40fe61a86e8662ef4a2ebf69fd0fdc17701f26ce4c994a55a07e6efd84dec4f771
z2cac73d5f242b15e3b39db47c18c03734aa7f7a31d22b7700279b244fa33269e547f912e1bc576
z4558bd0788714b4e994ebaeca9f27f3a7497823d0bd06aab5094d5bc8995f93a0281001c30a4ac
z7650a6be67179fb52ca912ce3f6c5aac860fffecadfe5af951315baa7e2475c1b6bd335889fa0a
z3f3da1e5e7056880d256e2c69ea465bfe09295f48a15967578b9e5a986049ccde742f6866b2ec3
zdaeffd89df0f574903b85c13683659a174a2b2e3acae045864a13fad2120a7ac7a4fb170ddc353
z9160a00873a682e1a1e7a1f2510e0edd4f9fe3125e0747e3a50a5538ae8808dc992939df8fe67e
z2e041ad3cec519c794d06478e0e5fc85e8d7c26507db6f8364e8f242771d9c4cd6975a8ebd539c
zdb92438a1737c3a211d8c4600deeb3527251acf557a328c62b4162aac77b6c3fc25be09c295659
zd0a667715d157d091c873a6e6591d2791bc5455441f3b4bcf275bfe1979c83eb5e790e828ad1f4
z6fe8c64aec6dcdc32aab96355ae04d45a6ad29374da96eaa7b549e07eb12712b6bb58a7efddc66
z3e8b51ea7264e272cf1dbd3dbac8017e4ef041f3485c77192b94e4898baa73fa28db61c7e3242b
z91e79b9e2b5499fb35eeae0be71ec7bd594d9715b3ebeb084e23928f6e51ac36d0aebd54135cf3
z34bfd28a4adf7270123f6bb859637189b1b3a7cadb725ab521ff6721f38a1663d24980a194cc0f
z5a289efa8d3a025120e4d5175ff90629663e2060a10f79a420446759c3f6fea563fc583c977a67
zfe662c27ece3bd412cc670ee6dadc97d59e705daa842e3ad77b26811f15ef755ab35afc9809819
ze2d1ea60727180924d6a0aaffa0a6ffe258bb95b5139c9f8f845be0085e3ceddd5e753bd97617c
z338ba92aef669eac307e5bd5232e62d339fed9ad52f75510fddb9c36570a77e993d12aadd540f4
zd04a2ae803bf9f2830249e5aa65dd04e471f2da60a58566d7f8826f5140ccc5d7b622a291efb9a
z7836bd4826c3cd77c4f3afbbfdd547e6a98b0c8d92ea63a6b6122222e48803439b04e9f25bcedd
z175cfe1f4c0b7eea18632edd657b6e121de4ec51950c123b2fb7a5d0729a47aafddca7a2dbc07d
z1fa56cb5dc77866b8c3905889bb4283c5512a42874d7ee56c1ce6e307a8f0be340adfe78b568d2
zdb7de4f55c01479dc77b6254539b943414ca18e3643a3b7802f50517c8425cc7f4a5bda80bd36a
za836e09363f1b8a8c18e65bea469f698d04e150de6593eed4f40b4f8986164a1300587b6188bd2
z3dabac6a001fb0e08db8f7a2d0d4352b805c4a199f2711d75738d9b1a9c84d5f2356356839fe06
zd17e34ad8c4a93b120bbc682b63d13ef7bf5ec7a692ad36234648638c7ae7a5a08fbfdc1b7e114
z40de7c81d14d1ea5c31ab34c17a0adbe10f0cbbb3984977354edef2bb932ab2080811e97fad87f
z09b6251be25b781e5a66bdb1ecc0f192be0eb61996aa697eb6dccf7e85ad586e6b93839f1cfa57
ze43debd5ba0664f4d7f5a7038ab61b8417ab559bc04d4f1c167915337a107c10b68631f91f854f
z047b87b43b8711bf3a25cf8aad687d681aba969a29bf3b5a2a20bff0ad2e80a4a3590225b9303c
zcd01508b05e3e1e3945f9ec4f2eff2303782bc2ea6ebd78335cad502ae51bcd53fdc2b4f08dc30
z48c98b2d7ea65cc0c083abe6cd6e4d877c7bf20c5e01651a24af45943b3333502be7750b74f804
zc816dc21ac7479b60e459a950331c6c807dd1044c7b30726fd16bcfdd11320b0e8cac8618f1b81
zf60abc623b33b817495237da65d743f2bea08ffc1d6a231b186ce9bc830cee6f0472a10cb4d5c6
z3d5c77836e9a311565adfdd53a71b2ddc720f5a17ca95f7dd851323ad98076051e6cbe575c999f
z27268775fea8b2c7d1a22ca41da5c2ba64a54c2390ee6cfb5c3568f637e0081cd5d8cca44e6ce3
z3fa4b5e3563d7a9d64839afc5dd8ed402c0d843b87a68b5593fc539217cfb0f663c4644e0e86e0
z5c88bfccc1c160589383717bc60c19b1f5dba248bb3fc0753a71c2f01d56a9866416d437757ff3
zc48a0670fd2f00ee38c41e47f49b77cf640a227c1a6dd1220df25ba5750c6a73dc4a6f256d5f37
z1e7e690d317bc0038cbe06c6f5ed9c492a822ab649a6287767d247876f76d4a3a08c6a867ea6a0
z5f1558d6b50ee2f80e3007a34fcd0cb48e9ed484ebc6148f40720e211e332fd95af3fd4b7c03f7
z5d77d2ffd8a9ce0db291cb5dae39ab81fb7d0fa9371a4538f6aac6a9e6919c139af7f900db4dcc
z18021979b4daef6480c9939a57daa1265bf91e513a3a69c40ef30baea14d65010c8899f81cb9de
z09e8f317673d940f4e28b51b688f4030070670d8cdf6305fdedcf886b540072181a2ed3e255360
z92ad676197679f9372ed7709854dee9d30b1497269c322ab9270b918077a5de1320567ba61b351
z34d6b78ff938aaece93e4745d342b9ee8743ba4a652455ff56f344a47e9efaf2bad379be78512d
z3558275d85c503b1b72d652f812d97cb642d75b4b91bc8376d502e8085a20b3e0d3902cc4b8aae
zd9e6846ca308ca94cdd09b23cf7a9280004d1df7d19f7ee435efd7e14efc65fdae368e02f31414
zcbc5e552a312fa74b4bf88b084d3f67a40bbbf0a4479d58ae91ef195dd4ab795302e965bad879c
z2d4cdf74603d3ddf6f4d1ca5587985d19522c65a7152cf2a87bbc440be6a57e0b9107e7e32ef89
zaf439e4b7d151a2347a5f67a45bb541749bdd8fa6a607be4be15832ee3e34d78e578f1821f3d4b
z005168c1968156569f96f213c4da49ea26565780a26d6ed2764b172b5fd7958fe9e3020af429ef
zf025a6045125b3a70d7c77c8cb4cae9215a69a6adc5ff7607bf8055d05c7a882b8c1ebe436adc7
zbc1d1a5dba106e6b7bbb9305a4472c007e9ef00a62b7e8a32ee79882d50942c70ebf8590e3626d
zcec81f2e694da566373d2bfa61a2653223e47ebea062ecef694d6cdd0a70e419a8170ec7d776fb
zdebfeeed5e402fdbcba128f2b10257b3dd2a0b25e2cd6485c0d8b52747a06792f02df5b6ad3aa6
z798dffd446a7c3b1b6096019b668bfdb110fd907c1d4ee13e69e7e785c1864aa838e8912126cce
zb95783c45c14910ebbe5c7cc5ca2ae24254f9fa672757e8bacfa1a56a860cd157768ae76692b0d
ze1bb53296f13a7bd749a8bf22447f49440a8567f3456894bbc406d1bfb7186f8ddd43dbe465941
z40aa02e6275e8cb39978bbcdd8e9d56f17fb902fd0533bf1c8467f153f2e34c3a87845a0a25302
z45c3bef9d353c1e196591480b069ee97d98dd0ec4cdaa86184fd1850058b242f2793125378fab6
zad49990e5dd750d8bb05fcd1f9a9ac34e479943efd3533f00cc90b9856e8ac0b144366c3eaa6c8
z5c9705c4dc04adfc679ff9ec4f05892898f39ef915385412354e7eb449a995e97dfee6192eb063
zbad9b567f1ccb6b4746f87f66ed909940fa63d9f8d3b7e7ea22671a2e51f5f3449c0e69bbdd1bc
ze4fd404bd1abe545776db6b154df9d5a6b3bcfe53ecadfaccffc742766f51d82fbc4e527e83283
z08fe375ce6f031bb761088aa88a92edc441f64c915078160c6040f6b416e7fd2f9ce7e5f8e75be
z3e915fc0f67f7a236a2f1735d95d4bfdd3a0e6a03a38e6876096d95a5b776fc298de6d6e3c3d1f
z3f43b8c441c9e47b221bfefc8f880cec19ab0b0b8ef39cb00c051578ffa8c290a87c77a692f219
z22b6ce9d6a22b11f9620f7da436ead33cd5c6d8e2b4eb2151ecc74b873bae6604cc67ec3731f57
ze4536d798d7a4858e657215f5d5bc4d4d8e447670fcdd2255c0dd7d919df5a2f92fbc25c6bff86
z73595aa8e47bcbead83a3422589429722899ee246134038a4ff32f0ed915d7da1b93fcf26eb323
z026362340fc006b354229e10edddb2b986e769ce521b00c6ffd5a31f3f83146cdaf7f25f8c937a
z6e683421310d5a3f5cabe7920ce2c0fecf32c36497cc34ad261ea843a209dbd9114461c543de8e
ze1464268c802240c40d7b9bacfb1d87d9d9ea966472d36bcf778a2e4d5b18ca07932040b1716b8
zacdc730afa38f5d58aa14cbafce2dc4555144e4c8cb6054153bfb8db86a6bfeea1d5de6d69e314
za5059eec3b91ff1d673ba7082f0bfcf9c3b15192bacd98c7605b5d3e190600d3718f8d69552f0d
zd4ec6732fa4bb6287079ccd526e31f356b08b0022336d5f849b59bc772588e7e96f141b9f8bbc5
zfe2bb8967dab882fb548f4434dd14d74307fcbc107a014d676fb406e0e863ad033bdccd59e7165
zdcb5d23bba8aea10c2289c6c854acfcc5103c72cda0e53c53e158730823ad912bfc9b7c63012e7
z325381c6df6527c6d6b6052515e1ee506d0cbf50e5866cf949c68429525826ad38a1af2e72293d
zeb0929321107268bed7b477043525efd148f2a5e07667383a52b035f00228b4484dd1167052c96
ze1226e53bf4940e2b3bdebc11b61a6c1bb17d54af75c892393152407daa17feba45ad7bf46fdbd
z5e01060fc9010b17c8beb562683e002c0d9d5984c6efab6730074f75cc8412caf91dfd7732159b
zb8363aa7d09da459340764076fbbad98c9635353c3a2a7e209929cecbabf51604a85dbdfe48262
z7151a3609a052dc2d77b11e01e3322751e6b3421ef14af3789114c64a38dd933d0599adf98a478
zd066b5130560f2fd91b9d133adec35cbddcfe7fa7fe1ee4a3d40477c5b82d75cb78f3dc85761fe
z7db65ac9c04f88650092217a5853d0f732cd5e4102bca60b225234a8139ce4df60eeb2d2da151e
z02ca163d87405b55c058e03a3be8b3bea9f2d2dbead804160dadf721348be18c83f14688e3f64d
z49164371d8521366e534c9bdbc449ac04047eb87020f36e46eb2d3fc963964ad3d0899694a1bb8
z23bf2ad127d717aa4139083399f7e20458ba9292496fc2e1735c77a23248a57cc827f948f74a47
z2e0c9a251caac8c8fd9770f0171551aa792dc3f0fe557e30a3d5a8200029aab36ac2e01a43b6a6
zb779412955976ae8f02518d8e4830588773ef09cecda55027a45432e1f323da98dbd53835c47aa
zd5773c8fb0c4394db4ab46549d04b85af35f0670b35c732c35b5b0facbf0e78d20fa94c7c329aa
zef8b5239ec7bfe46d045453cdbf292887650099437e53145583efdee2aa964ca211cdf83a83e33
z85c79f7225083d53f7b89742830a0d36725f53b64a961ce535e3043c00d5e473ae3681c4cf0be9
zb253141226cf64c3a93de574ab66d1205282af5eefc06f7b80808ba7ff11d3bd44ca6bb76d7d48
z41e9b23681a13bfd1b0038d005aa28c9913ca17812d1768c67a79e8b1e0b01c3715269d9c4ef5f
zeaa5f59635082f985393bd88bfc7e5e903a47642b0abb249484604a840f07efad287668254d0c6
z39562511cc56ae6cc08c6a2ac72b10634269bf7dc8b02328ea8d2679e22d2df860e92d35304f99
z0db38c99435b3fdb9bd4afcd55b5f607f6ba2c3d2a69dabe8adf32100394db5d3444dd175b7718
z1cda2fce001d21081fd08351835fce7b5c96261a32840f9581a8c420f5967a758847ddc39088f2
z3101d39b8f58f6760aa2d7258a69d96596f5a440eb0e5bfde00408d82d9a9c78ac7f6d0585fe0d
z11af34dd6adc1a4f0b48ee401b9968e89bfef631a606f7a8b6c937d236ac06642f380cae9f9867
z131db692cd68b3509ad72d5d21f9ec61e381647025528630783bc05911404988af4a3682dd4457
zabe838ab0d7c99b2ee8ea5b6fb253a58e22064522ef3a6e664648e6b1830ea1f719379c6583309
z4e7c080f8548584e8701e0614f75d1edaaed511e3533f31c15c3368b8ed5824aa63ab2aa072418
zbc7f5a89d2007604c2e9599f14034bda261b3ee76e196df691dece5a154c9d77cb8e4dd0eced91
zd5394de082d61d025cc3d34b88286190d2494cacdb04158556e9d477a58f3e96346369233c955a
zd0126c43cb0cb81fe7654b2e62b21c67f1de8e065f5b4023e6edfc54e6da0738e540b55c79261a
z45befceb028fc623510fc84f172fb27aadf0a33c6f5ea11d201233ea925f27790aa33cf9a01329
zfe365a8f6410b51791930faf1689d41e6ce499b86b41c16cec6bd82ed5df8bd26c220af81167e8
z3f5c2e63ef32bf5f2431979af5d138ddf885ae296ee9402af51dbcf582c4e248da0da3d19b9585
za169922da0dab8be874dd53021cd3acc50e933dc7bffa27e3dfea3bc5ddbfcbdc382520b0ce0ee
zf311b866e5c6bb5167553c53e3c040aef2fbd42020b602d1bd3e8a8078437442f34781824f50d7
zd61da9e4e69ac610326c16a319a72a4e6e61243be63e9ec282c3050f80739178a6021fe01ef05f
z16bc24a599301ce1bb0ffc6aa3ee2add5054b85d800f26e7342345a49e3ec43a4e1afcc433a841
z9c5564facf10b15fa8230145196eef8e8763ebc8660ded5cefae4ce0061e26f70f10828c0f2f9b
z50f785bda95d00a02b96d3f802c19b7f8ab7349bacef583ab40fd791a045009465f9735f1a2d07
zb29bbbd9705f7e34b9c5a0789f41c3ea0f66e90424f7d0ef74270f6ef875d2550a9f1dbacd19cc
zd0c8d47b1fc7def02d751083e680e1c8d53e25023ef120adab9324c5fd5337ad43bfafaa8cc807
z3b5f22439eea5d282a20af2ce74f0bbae93c8a588e11a1cf6217acbb9e4394c27817101618756b
z9817fc4f003d8234995801310919358afe78ba8e01c19f389ce7b457b19e9146528898c175549a
z97ecf8c1f2bcf74d791e80f4c3d68293899e2423b72883c1084c08daa8c507d06859b0cbd6f0f3
z5f8fedff3e6148898dbc37f9b5285af132691133723cdb8e46e6d8e6cf4e4161ac8fc8f7faf103
zf833a3494edf68bc3789e17df0ca090763c203ceee3e43d3883204ba8d28588fd39158eb02dd83
z31c4f9b4d2a8175795596170c2733b855a50990feb0d2fbe1af219143c0d5fa6e198d4ebc7dbf3
ze4922839541fbff2b1d4569d2d44f695c4a1f1bed031567da26683a9b0de19970a58180992cb12
z1b6739d58e132e53b75ecbe700acf003f33b1b70da0a79d234bbde4200f2af3d26b949e167e949
z491450fc796a0088dc587ea778ff337959870bc0dccb2adf5f1f6c7566afca03ae18a17a0c164d
z75c475f1b1dcb967211827ad2766f7599739b2a8c9c80dc84d1257cc474679b630e6f500a0c045
ze5b910174295476c7c1a7ab71ff12278f62f7425263591ce13a5eab06263cb7c15059b29e05df9
z1fa31e5315b9d7d9948916437a73f56093dd197ff6863a83690cb0ad10de630b529decd3750603
zd4bb7087b778b88d2c9689c731696fa090ecd96f0b9f7672683cb9799f88a88bcd10e35ff98e66
zf2096bdb544173abd833b8e4f43da7ce3fd76af3501a3f2ffd66470ba866bdb4d77dbf3ce8e269
z353421a8fef11bb5593eb978f64edf42e5408ad3ab2392604e8ec647a8ae205c0df26ac6878719
z1ce5455a94f613f3b5241b619ad21719b5831c771a4c53c439432a7f5aa2ae399f6c4b2a158fd2
z62026a4a65e8f8ed321ba82eae2aa20349b554e65427b6e9dae0f5034e000faea2141562ceb58b
zc1f5c35fc75a72c895ece34be754c35af5fe032f586be677e14ea6cb4d8e9af79a9a8a11fd1e53
z4786361e94f0539a2fa9cb41cc7c5933c5eb3ae60dd098a89ed8e1b644a6232079f9df2aa74df3
z81500fba532128fd8d8a526451479030a8cca3a4177155dd79f02a43d93b6016f2c3d98e961a17
z2d9d9dffb198249bd53ff7fe913271f08ea80ce2f20ec0aec995d67f578d05077f5b847a8a6a78
z7e9036f29016d07c0e23ec4fb9078a090ddd240f0566de9f3e2693475f4a4e965f8b06003536a7
z535249e7a1ef482e58de75b742d00554130abcbb6b15c2bc03e05211acde01da052f0fc68ebec5
z97ef776eaa48333b0dedafecb473ffd736bcfe5b7a20a3ab3df1582d7dd2c9e0f21bf715800665
z7718075fa96e445cd969be839a7dabb4caf56dcdc59a3355118b71a859fdcff1774dd17e8125da
z38039983998ab1bd25117c9d7d4a7dec016797484a3bf1379bf03d69b070b4532d361f413b0a6a
z13bd04b6a1db859e47bbb7f532c9b0ec9b1f449fa771f73fa0cc09a8d67dab74662fa67b69dbba
zb961a001f49c47d096f9a70741b97d5442e382d79e7e565f247392ab28920a72f91f551aad3d96
zcfa205af937c971f4bb9eebe2225d83989c17fd92d2e51abee2b44ed337a6ac6bef6c70c43303f
zc70215cfa27a65e29b68b4090da15a655213f019a605c508dd48a8d019b129d0356b4102a50046
z6e9a58e4033c821da40c068ee0e6678074bec0b19bc0c6b563c03ef758dc7391a13572ec477a81
z4ce97d40bc2a576104840556a0354b1145cfdb19522357411a560287e6fc9810b821ef9efee01d
z897f212e9ded976d9a7eb30c9d401a03a43d7fea486cd5d3ecfae7408c7be95483018ba862d586
z23721532008a9a65e62f8ce0130a03fcec3745cf9ffce5523c620f72b66da4f902a2d6f3f0392f
z8ec986d10afd3478840f61f23b3bf8535fb4e8d7ef41bee4da9e1353feb5665dec75257005c61a
zea0ab5dffc7225f1a9c14a8cc6bd0bce82890ee9e1781b80a518ad780559a3393ba163fe6cd046
z63afb4aaa6d6c33166abe4eb8dcd70968b22f10dd3821ccdcb89cd893d575053f5f17fd08b1cc7
za9e29788afcd4daea008376bed228fe14e70d8d15bad42a327d98f16dea28d30634a90cf3f1ca5
z984d1720b3bc6ad3f163cae2277e9e18b5df2cc83f79f562d901cff930f77cdca3226fcd2d050b
z2088b5bc559a735b54a4c43775180202130606916fe0f1e53260f9e6c89d2eba7b7f5706675df5
z6ed89446ff383a4412c86bbb7b287b0b922ed94ec42585f5a91f97ff6cfc4ec0ff618310efe0a5
zce021823b22556516fa88bf565ebabfdbe4f7d53caf7ec6e7877f2d10e29848f191e559f693df3
z68a164dbb67a1eb529cb25860543106c5c7d939c678387998b2afe389b2c7609bd19e725e95f9b
z83c15bc3e29146dc886128dee2a8fcd597d06dcd23d80b305eb55d03aaa6d1870c062561b54af3
z71a24d2b13da7e46a3799c94c65f7308ff39e73f5ce6f3eb16f9afeeff5b24fc142e2b76f3e455
z3e41d66f3dace2dbb99aa55f70a7a3bab68442fdb5818d6bc32972a1eaa340b40872fbb1c4f4f3
z5974b5d7c537a5b8532d05e5d58308b67fe8f943ac3c86125b09eb11bf85d2fd7f11a237a54f0d
z0b6a1c282e725ec2594986d3e95ef324b0dc16388d051615fb68a22156a55d7ac5be5e2512555b
zdc4a8690c40b4623be7e8d1c9845b67928e7af2a9c6e5013606430161ce72b9b1e9eab7d0398c4
z02eacceeee5ee93300eeabe675a44e85696a19d7bcd4c11ec646df6d2a5df2ed8c2ef293e722f4
zc18776be49960a8ba87f46acb5bd4aed9b6b5f3a464473f4040f4a7be80f0ede15314bc2286955
zec83ee827fc497277cf7e93db9647193eb5108eea6a78750f682fd10536ca6a9d8e6276ad1defe
z4c3b89b19f038bd151129bf00c9f099c8794fc5f85706c1303b7a70ef5c0a5c9e35749b7785407
ze3ff4b146182ea35cbc88965908e05e21c218d34e5fab66d9d15f57f6b95e2153478c1da321d65
za0d07f2d7bfd5949d79fb63e166c83f19bab1c6c0c7f0e6006d0a2389c5afd7841314231cb9a4d
z02ed2cabf9592935bb1f5ae7292deaa619d97efedfddc270c673a8f56b02d27c21c9acaf53857f
z6a0f29daa6c0c76a12b5d4e9925f4d96544f4a5413fa18561fe1a7939d68ec823be8b687a6e24c
z6b235da9482d7f7f5899af7d04e7d975ec54fc6951a2e2fe1cb4f2341e4309dfbd3c1a85b9b435
z8b646131029711640a9dd3aa457684cafbcb54dc69af7579cb02e4e5e57c7b7c3142194f16e8fc
zd40f004872eb318d53ff8c0b5229218f9e1599d638d89576320d7f74dc5091df1451ee1d85183c
z0ea892122708c6d6450e76a2aed03ea30c6e04b565e5034c73b0019cb5f36d52d890e3444ec034
z0b669c00388316b9a83bc1dfff67ffea631fdc8eb841c88ed40b54a63ce2611ecaa1d051fbf896
z2a260ebe122f507ae012042fff38f1f375634e9f7bb74fb513281611368fed59080cdd4e35a0bd
ze9da0b34f6bcd7bec7fb1a9930643ad42cc3c3d0db2c0e97efa9e69c0a7c4da425f25b7238e5d1
zbef26a4abe28b1d853ae3c40b8cf106ecb9285c93fb1288709d3c10dcf9a41dcb042b9025c8c15
z249fd957900dbb0c9dea2ce4558ef2dae5f09f3d138f3d2103f5ce44d703e7fde1b56365a6b70e
z8602e9f77f54edbf04371a17dc1613f69cd9038a18f2ae77befc8cb8d6032ea36b0d6b0522f2f9
ze0883b3c91de9f2073dff44ea911b41fec6340e0b7fb82945d0b127f69678a53605d19286f8d9a
zda728ae175435f80859a94e1b0d5342c90ee7018201fcc6ca998973c63d611a6b6597d11890627
z71624ceba01f37331b8bbc562f171327f80e5037b955bd96127d441e36fbb725496a7b9012b274
z4c49df39128553f5908fa747e360a4238c7575dce529c4fe2cbd6394a4c5f7873f2ec352d691ba
zb0638a6e96829bb8494349d5b61eecf169ac7ff698dc086ddc78c70d997473428a761ed63d430f
z8a3d6a204f71b90448a4e8dbcb1b57d191225b7687679bb0b9ab5fd7f4f899d5680dd281364c77
z2798467559f6fd8f04c91087e8f02cf1ca83e29340bd89eae9a98bbcbdcc2d762e23ed308fccce
z2932ab0b24876085ec9279712cc4a6b5bff63fa8be905041f744fd903b8e01d8d39db84e5d961c
zb8ddaefca1bd8aa845831adb18e00ad4792419da553c6f295cb4db6613dc4477942b39b0b05773
zc077e36ce3982e768aad6be8f673b860139cc18b52c697caa714839dccb0a5cce83034ea11e4e6
z7fb033024d374004ddaa2cf0cefd95430faadd398bf26f076b3c7359c97f3154c305425e4b25ac
zaed303dac40c57bff75025d9da55fbbe094d043cd5c7ae1b45f9e4cd8b239ae46dfee2deb30186
z528cdc0947f4115ca3c398a23ea3dab01484436e786ba477065b18e532eb49d94400bdffce9cb9
zaa9e1d52ea8f5119f58d8601d1aa8dc4253222ef7f79552623f34537632174fa69bc2623786a9b
z77e637b436b7c63443ffe304724bff36c69e5476e3f779932ff0ff19882fe1a6e52e2c15e972f4
z4c9476eabba8a77d2ef3a73743cab8cb5710650ebc83c5beded34d727cb9559af91afa67e0c135
zf0a59ce1c69de557e6cc4bc25354528527e561633c9b5cb0cde8e7e08db6b2835acc420860742a
z07b3021633ec3e5bd428a85c0a578cb65de149e72269988161a1fad3a3e6e9ee3ac07ad91cb9be
z7c0b3b5a390f4bda90b8d96b5765bdb0e26425f37254baf940cd859eb3e4f6558ea6a1ff7da6e2
z965e46b8f2f4fa2986ee1358122a5ba9f349397169aeb998c03040353373fca78aef36b91ee893
z7ab3f0eca58964bfb1124305945272b5bc6a132b0987f7c43a9f479ca0c57e109c96b4d92a1c90
z3a9dbd16d92caa2d2b813673a78d590848f1c5a330f33701ea469cff2140eea0bd09ae132082e7
za58bab4b578535de304a670c1d82f14b91a53ce2415c79bbd631ff3cd0624eb9c1f63f973f2a21
z4e69c05e863c1761c95c4f858e2147ff6e8ef931407dffb49f6a20fb2a6061c4428b2162593095
zb87f54c76b271d5549dc240e38829a45084b95f482ea0b0f69bbbeae5ce4b8f8c10ff7fade9396
z0662b77c18c9f0c3223b3c17702e97426a55f416256dc63ea6806d380f14d40c2cb43bdb6711a7
z792b7d25ebd54c612e3325af07c0b0df2d9aeebdc4a5f33a7212cf3029f6028ae3d48667583c16
z2f757032b176a21348ab6f3d367298ad78d938bf91e3b833b0d33523343e5642fc70623c923e6e
z539ae3dad95c7428fdb39ff586071a1060d92c3a30eaa901ec9296f7449ce008dae42ef20a76b7
zb0f84146259012a86936fb47f76b40277367784599d37a37127b11974f400de6bdabf127927a1a
z0ead6cd63a7e8992d8d4792ab281c777034ba6b283340451c14534473c547753d7068bb691e80f
zf51fc3bc982fc5ce261afa9226477cbb15b1dbd468a4c6faea4caae6e7313490a80d1b53340f62
zb8eeafddbc48e19d03bccabbcac13542b9f948dbcf652dc3a89eb4cc8564d4a8974229bacbdae1
z7224c2be8bd99ccfd53c85bf7d378fb36fa8003d4467dff6c3fc42a8f488e3a11041de0e809a8d
z2e63cb7b8430d7eb5f3535b5ddbc82da97a0195b9a0598af2130b20e54a6db87019e306a881433
zbea925318dfa99ab214e1c71e14c94173a15c69e9e1339d78f72c8851b963c09337eeec37da703
z9e8fb64660930e5786a153ded0b98b21fe4bf9859e8b1a26672ee276cc2f2e2d3ffa140a9f498e
zac377b715041169c2900c0b809940ed9dc0dcf6c3093c7dace41b04891dc32f69e0ee1b8a38a7b
z8a137b97a54e14672e4fe7cc31700ae68cddd370717bd911d96b0cae4a8a4f7957ac3b09fa41c1
zd9deb2dddac6ae2af19d10668c4a410763c78211006dcde31833548e9596f76469c7789591ce89
zc514ed3b5b9e909a75e56cdc2a574b76e9b3076e9fb9e88e46860b0977df259933c59beb009d40
z43c4b1c3f71b1c9dee5c4416261a97b620f799178c22bc13cd860951417fa004b74f95a3053743
z04a59500a9c1156af94133e89d8ba4fb51cbafccd740c756bccfe28ba9f7e1a432f7ec91e9c551
z0b3772f859c512e38599818e971c65a7dea6c2bdcedf3196b0ad0a1d5b261215c6965730954ede
z7ba7aca5201bc5a62c12ce0008cdca8939a3dc837a20b7e52f5db33d55c4091a068e2f58c1cab8
z86b075ca39823110728dc46512ba5481dfdbf03b0bddcc901d757e4dd1c18293fc2872ea8facab
zacb4680b9f9b2d28fb1b0825789fb21cb087a5adb695e35c3814efee2cc6a22c8753f0e979a94d
z6ec88201339432f1a260a8034cacaa36303003b1a27af25089162d082bc4622cd45cc9557ade35
z6c577188ce131ba231bfbe96bc323cc61d09a0d3bec33ce27a881053d905cf841b9fb026a08d0e
z6275ca111995d0879d8bdb69ef15bb38666e83304b29f5993af8c4592592eec32cac8c9a22552e
z5339bbf6d5d1e82e16d06552f900179221ab14aaab938eb8684bacf00e3602808ce742dd851810
z7406da4d07abb40509809824d2e6097d102f4f61a5fda676808932c9d43dec8123d2bedda1d4f3
z3827326964ec8dd6b883e20305bd5256223d2e12ca4cf844b7e108e0756d34f4f0acb0709e9630
z62230649129dea91e81340901fd1a6e2371ddbe073227a0d96848c8f671d8cac7684928709128b
z640e9aa741b6fc383248dee2b2b3068578802ed9ec4015f38d7a06baf4bb8596256bea5f6db01d
z11cd690a5b9e270f483380c9fd36e4f65eeba6417219fbe3d6e874325686eddceb747d98a35c0e
z0958864b7597c766ea945463893e116cdcbc72bc244314f32bbedfb289cafa88158ad6c5566a8c
z093b9df4a35f36428e67f3bc4ced24ebd192066eb70867682c0c405671e4dcc64108b59729960d
zac936a66a004143b04761d8b785a730b5ef0d9fcca0593b993a19111f947b9788c545678b56185
z0b4c799b0aadebeac4d1c92c90a0eafca20c72d2bb758b38c2458af052e0ba8067c6e5fd790d11
z30f86cd892550fee0227f6b5350286b4f4368b455a7e33eb34bece7be7949974b7bef2a97b5c0f
z4e9d20be5309760a0e49a87154831e89bfc75404c3ce49d6e9da65946ee52655b70559caa0f905
zde6bbc1aaefdab3a4a6cba49433f0834dc4a2ae0df05e01113f6ec52ed5a677277c53a2ab0671f
z382252fb4c829544d09bde873e6a490f9db1599b4439c957baaa644e6e264c820467c8b882cbfb
zf326e04715c96f35eb750d212c8f3f4c0aca4d68964bcb2e89e433856a5a1f216e72f8f60ffdb3
zdea993526123ebc793494d547bd8f1bc09b95b58fa766433623c9e87e74d7996255cb1c0be34bd
z9cdc8ef7ae2506dd05128651b2b2c3c3609396ad51e1845c7668bc19d371d9032a5e56b5aac011
zeae98ce93e60bc02396a0a6ee2db66212c0731560a30b271dece9f510aed88cafd4578ddedc689
z3ddfa1c740210887666cd983b0709257ac675ca894a06add1457323551e01302b6c73f2f2944c7
z3510eec1fab0c330a0171650c3ebb533ffd6699ba80aef7b7bebc660c09c7dbaa094a5f833293b
z64a87624c35cbcad9e4ea0979aa0edb6eb29b978a86ec39e706fbd3b825a85f0bc140957250c5c
za3a1c23e9090b17f1ad2ac6bc6fd546f87d88706f20cde4b21860025a3008714c4751e4347e771
z0b5a4e06d7bd460412969944ddd76414381a3edb4bf1482cef414f1174e37153eaec3f7177fe0e
z88ea9f3a068a8db56c20ecfc08fc8c3ab77e3f96cf7c3033a0586abebd4139fd99430bd05175b0
z43c8923d8807024e61d43ac7c8d0f020b912be180305757cd6be91750c22777244047b9cd473a6
z800e20df88f5185bf33ef2017c83eaa6240b3d668ea8ca32ac33ced494ab53397f62d3ae65c9d4
z7ef84824acb7f1d14cf75ed6f7dd9cd0b202c4b2c2c73ed644a2e3b880b221b86c0959d51a26a7
z43e669aa636ec6f202f2006fa1ca2e8c96394c16b18d3df475592043c3232339fa09226bcfa57c
zc5f2fb6b4a814f2940f9df5ac5e4d7f6886efc4ed295750c36890c83f607c4db49deaa70f59886
z5ae905f4907bd46cebcb8ce7410c64d4cdc6da80055f2f210c0e0e475bb5947e9c1c73b410fb18
z49cdbd1a70ec7269ce096229ca9649d03bfa9e88d5608700183c2514716636770b7f7444b9a97f
ze28a9741fac5c3c5774fe2fadd354e3ad96ecd73a6ad4f2595abdf42bc41b19e3d3ec7fca8f00a
zcd152cf96a0bc567c5fd4e6c5f3d8b60ede65336a9fe055bf53d0207ecc875ee29befea925cb3b
z987acfa96e59bf7b8adfe6d79ab9b5158bcb2bd95b25f05a5b008f87aec1c8dee87ba547ebf9c7
z11e74c83068a1afc009336bd7d34ea32451eabc357c0be541f7a3c08bfb2390c442a55ce10676b
zcee75690129ef1fe15ad6d68f7c51a147d214bccf44d9745332b8e2d9d223fe968bcd92e26219a
z1133a3ee27fd89a49bccbe578a11e24e22449dba77d3daa5879425688169eb27b67a373d138e25
z26d1881927f2a6c998ac1e1be480b6921b69bca76b6df8ef6fca942816a433e8086bbe636d8226
z31e48b57434f0e3f4a9e12cce718a9f6e0d2d0b743cff660e9e91cbc87b6f64630dd9472a0e807
zdd90066eea3c842c96b69ad92202454491c5bfeca5056b7ced458475fa2b774b56e0b76833ef29
z82801559132a7d60741fb59c28ffca9d2930bbabb41576514a364e0f5ac08422ee702b58594301
zc39a13865e4d7281dc35b30effa7c653d72a0fab8ed300d59f2b25146bac3e9d12a5adfda3858f
z4d42ffecb9bbda0fb5b6993805d520ed5d305bbc4f0be283f64a6c703ef54f32ff17dc40c8cfac
z88a41d3313324dd8395c20a69806a2e0b5f7d3b3070578ed2399d8559ed444f8a65937845c5671
z940fdcb4210df42781339f16bafd9d7b88eae8ec68b21fccd66035acdd14c3285a1039b466575d
zfc7f73d82cd815e48dc5fe7e8f70a15ceccbf533637176b49cedcb3c794aada0091ceb38941bb8
ze28d4c4d82ddc47da5fa5366ffb44c1108dbf0fb7129f9bf3ee3671e01054e49dc5dd091d1065f
z7dcf2759b00239df9af2287641f22e2f13cc2d9c612f2156572c70c75e888daedc36a67cad8941
z0fac2d08c8f0b6b71d2f2a55c87c3ab85638e63793f0c13f331a216d7c19eae6fec08bd7681617
z9d6b3420c64f2ee1ae01cea3ba6ba56c747a7c404add66fd26c5af619d2782fcde07eee57ba1f6
z4d9da5c38de21cfff0a7400652e31b48aba7a5c9bbe0e5776b62eccc282ac516d41625000e68db
zb2c3d1dc051a6ae43bc711a12a6d665b67ccfc6323b6dbfb3e1f1414139156c0b61e969ac3b514
za78d3bd7cc9ecbcd16bccacbbf870a3a5fc3ecc6e30805c0fbfc602ef6a9b18cebc2bec312e891
z429df11b4493c344707d6c3272876b747bce8f6f8fa71a4846461a586e348f38c698df5cc01609
ze0f00ab79931a86da71ab62fd4e2f0ef283677c07355c35aa8403359b7347713ae4157762ca610
z03173402de1609743ca4a058af03eef642c1bd4bba82bc4f8d09ceae0c9d45c27d6ebc698d78de
zba416a7355ba10a6c453cbba09bf0f0f090164ed78828a18c24c775324df868040f7ba75919eab
z9e29dd93e6ba0de349e87896832bdd58cce29c5bf7c55e86359dca260f071ba1d76c571b2fc936
z85d693e229f03d6f7ed2a91902f7938bbc825c7f6700c371fe7e26a7057564d3dda1e8354f29e9
zbd1cf33342b067ca4f9f115d0eed73fd5c37682d45204251a653d8ace11368f88f4f21f7677ea5
zcff33fb53dea1642403c1cefe8f14a6b1e66a55c4681ac1ed2a67411678ddebe9b8c0fb4219f52
z1ce4c7389ccb56fab93b499ccd9f7b4937c54acef0ada02ac602fbede4856df85e1d0867405d41
z0ecb3da102cf879d58718efabf44d719295a3c504237f0a6c7c87d627ec698a0670f998cb55064
z0f4b26477952bf867b31256e58f4d2ba19cf6b55d437a3cd455e3d5879257123a931ff3a5141ed
zc0eb57ca368f2386120fd7f15425cd4b4228f62afbb207d67298de8a747533983a5c82f6c981b9
z08fd3f5d8a64ccda653b77b32a44dcf97fabdd866de77362e4066330fbba85def42d011c495cfd
z9ad23d32ec750a019d822e76972b05113b212e0dbb3bbf1d457237f648da316e4222f4f161a902
zb9017a7779d04e31213abaf8ba93ddcb2cc32d93ab22af21e246a613bf0e850a95b3f44f704568
z462f2c207bb35e559255193bf24b0d8b503371e6e62293edfffc17c68d954ecb96a538a1e4aa07
ze183908e42f9625ae1d6d3a6b91b30110cbc9558e3be5b35179da0f0eee01b709066380900ebe4
zc90fc483ba230cc1ad10402bfd581513e322a221b418258269efdfc4a8a113035caed67562b449
z46e9a149ce0f30e27efa97739bfcb6fae60e68042c366c547d931c9cb234eca5af36e13652560e
z20b6a149ba023b514dde2512f82541a40b3bfb34587e2c44287e1b137678a4535ed7a954bff854
z0fccd1e5b41b7f73a577fa2b50a31118061793c786e562e2eb99d655cb779abfe56c5c1a832c9c
z004ef5cc386dcb2020dedbbff091a75208dc7ed3c30fb001acf3edeba70f2f92f3d57d758ef5c1
zf105d26f701b405418ad8a45dcec60f42322577c31d58896230748c2ba0cf977c203eced488d37
z497500c77fc3bde8d4891981bde254ef21f3a757758b3ada46028b9e8b552b95d74b4b65672aa5
z288f2a9c2143f95fb8672376ecc27ace2bf0102352553d94a9ba7fc3924c43db50491fc4ca392c
z4c5e04080b641e4f1328bee86905080e4cb2ca8d0e13fbe6aadfe9a717af231dc1e55996872470
zb5d3fb48d0ef83c88b87440ccb1c128e80c4c371a04efa6389f4c7b5baa9b753981372ad2c6f79
zb50b73b20024d8c84b8588aaa492847807d30aba218d35c36e2dd4944a3ff283794192005985f0
z4b0aaaa8e922973472afa356c149e287dde4ac35f1a23b4525c085ead840509ce31bb086e9b064
zeb243fcf50a219cd21248026e858245ff73dbe860bc95b14a3f34c33a621a6738874fc7de1f19d
z915f71c08443e2293e29ea1db6830cf20e5f57cf37571560ec2f8bcb21a963b6aac8a44c13ff7f
z25c0e42aee006a93ab6a77ac65044dbd908b02ef713e500a7165c9164d0fdf4e4d1602c1f2787c
z461dbaaca49da2d463e8b5afb9cc328849da595e3dd3d07b440ef67186a1126596a2015f0c7c03
z64c416be4b8bea8ef2b0cde3d9b0969c4e9b8e46b2d2f3e3a1315630b124fd2e042a4f304c2b03
zb99ff22dc910a728c2c76219f586d00b8a405f6d4b7aedec4cff82c5e39f83eac01ed7b4ef643b
z128ec761c37ef4a72266ebb7fd78a899d65664dfe1e07a682bba168b495d0d2fb6872ed01b9bd7
zdeaa33c82a450e98b36d529f7c256a75ebb0142fb53620aa659c9e7adb4145a19e4ba430c9fcc0
z068f73ff4091e46223d148cb32bd8f8c46406b89d74eb985f9f74a7c8ba00a28e8ab6733ead694
z07179afe7b7f1cb99a321542fbd915e64f96ad26d52a6b99ca8e019b2f0462fa845a4a65968870
z9c8646da73653862ef3fcef73bcb467bf1df5278fc3e62b0c687ad6d56f7eac1f1c627c61fdbf1
z8790b22c46f732c14117870ac7628b445e6d8f7e45f90f800036603c02e3b38d9ee54e1e392107
z196628bc615222fe0a98fc3444bc5b041ff8f55746a9d614584f02a23ba5fa876deff3fed99512
z5f50cbbdae043c74fb7727f2ae32529b935254d7d5e7b062629e0771d61b005589f0fdaf1ac7c0
z1dde3b3f27bb696be564408401ae4c0a309818c0829a7e38d4fb0d76a48ab0fb503741e636575a
z924af822290197c654e53a87b8219440490c387413853464ab79cbed6279e671d430ad2fc5a894
z899400e1b79e58b9379a6647c535b940060409a4efecac9a893b66bd6c6c5c134f0a10966d1673
z8f91f3b24095d6beb5d961e724cc3bd327f7ed1945e70de89409ec2252c750a994b5febd83f3b2
zba2e5be8cba2fef78884d098844b4d1d34553bd2a1f6a47426d17c13ee1afaeaf9cc2e4d3ec47c
z5e8babc983b1adabd76cd4dbe783f96d7d1735ac5f74995ba7922ef4374ad3a3bcda570a5b0bac
z76c4775c7a7022cfb8d1a3de73a93857fcb0b6ad9f93055f34e1fa7a3b5fd93de062ed0e7166d8
z9a03ad1fb6d216023d0b0893201059734fe055a017346dcbb07fdfea2173ba777ab1cfc9903b79
z2a3736dccc41ed3443efe5bbfe1f1bfca0f6d3709e79c3ff69d9f23e9bad7b76de31724ad1daf6
z15759778529019c81a3a4673b43793f97c713b5e4c803c34f5a148788fbfc45f347aeb1a7a4c87
ze3c1decf845a2ce25fdb3c488c84cecb50dcf8bd6fdc6e82a257dc6b7dc8805a36516f06e080d1
z62ce0506a29665bbaeda92889ecc3ffefd692341ca51c89d7b38d2581120704e468260cfe36b1f
zea6aa5baf86ce2b2129361d86c77c71bb5e5da07adb9bd165e6e8ad023715918359a076509ff37
z04f987b6b259613f5d43e06cf74b4c1e2da66db0daf0d709e693c081cf61c353c9da74c110a85e
z251f7ad709c5b80804d90f799cb037c8e614ea10f3165365df7cd8a154f6504375956affe63edc
zbf994e92314e271910acc451edd5c0a5ea2bda4cc2f3bf2957ab1a290706ee7abe8cf608d10d42
z2d6d18bf11007c247824758dd9f37e9c56cd3eed1f091b50aa3b38ec30432868b518a10a105348
zc74d4c374f0d604dee427721d6ba1ce16daec3027abe086953291733ab5b8610b595e84c9c0b7a
z640ef4a72cbfa6f8d4b31799349ffb27d2a23347af851c3b773b3fbc26d273c3e98e0be269b934
ze610ad9533bd5de00f332fb27a1b065dd733148ca78c675cbd1d0918639fab43937f37183eaae6
z262f0273306c519a1f20527488c5aa236adc421651380de7d2b48da6761369aa4301b6544cd12e
z487e2c28cbb64e5f1247888deba00de62622026f740dd849f390a851b2606b5de0b6d44664adcd
z1a3947f2ec33aff850df92419db194142222d1238117226c56b38e91985fce41801eaaaba5fa48
z55c29295694aadcecca4457dafb380ba63e185fd5a825f7b1b27afe1386b459d00d47bd9493d36
z21fc9c709075f6486b46417e53ad90b984ac6c6bf09e8d98ac2f47c914aed0b34220324b950a36
zb024d46b0bb6447c41b3073dc303e89d5d195f3ea1ee854f1c96909f5e0224c2253608f46b26c9
zc5b8f9739dd040d2222b4c60da2ae0eaca5b1cdf325ba6e93720adb269bda83ce1902c73fc91a3
z896d6be43eae56c12102ebd57b0ca245e798fb1b3ca8ce07997a488d46da6255d9c9d80200fb79
z1e77fe18908a66a1cf24b17d1d1ae3b5fda9a2b03440622ad2ba43ff7b491565a0c41e6fd1fa45
z2da977658bbde3ce67abc37fd90403705657ca81d4d8756ea9de9a0279f312d291c2fcf3ef443b
z97989916040afec8ade72d857d8ead99ddd1752fa3171ca3a0b73f659317593fb7c664b29a292d
z44885c90a66336366780691d8b5c87a4f329f8b09f63f26530ff58c02b79d60e92ae293c2e08ff
zbbb913cd17be06bf64f44fb6274b7c033c8cee99fa9be605fe22df71f851314870f72ba95cff42
zd897acbd4eb939e1f5a817d009aef78cc00378c12440c605fcbc060343cde2f3375131a426b41e
zf378b6aef71de1c10189063212c128d284df9a2254fdd2735eb1b27bad01bb12d6762a3dac7101
z05c9ea31bee4911b4c4dd9b94178d1c51040a9b39ce836e07a45f7d3c66d945f009348e21325b1
zcdbf9ae408fec034a63d075a326146f6191f567ae1429bcff56e07fbd77b5e82e22cf49812b533
z6ba0c81a5fd40503aa87697014e12466aa6118271633c52d98422bb62abf3942ed48bc90f77668
zefbbc1c35459a41151f93f13450e887810d8829eed5cac5c4019b7f675c916b1600cf7b3a5114f
z8828a51ead653c1eb42a8b9d7021b98f137454722367ec24e0757bc729cac94cff652de21ba73e
z3a222e53990d75f30f7edae87e64d25695b717d629887197b09ab00e15c8abacd2656bcc8f77e0
zefefd2bfb30be0023d1ac8652020cdd9c2f61a5613d74fe7c59b8fd058004445d05af9b200d89a
z037443005d9d7560b9b3e8feadc739101d9fd712cea0bc8b115b07a66d25778ef7f067a2d7f266
zedf47116c9034184547ed7acdfdb6a4794d4339c8c7033af9be6bb64ddd95b6138370ddec46043
z03cdd0ebeb89ac271fc4565fcd21453b553f6927ad54e54bec67002ace4eb2e941fc3cd2016e13
z7da51ca3007cc9076a387582ccfa12cea57e4dcf37c0b86284802cbe9b69537e0bd06a21990467
ze521976a67623c5ac0e6ac2dc57dc4d6e169f481f48858cda5be520d4546a852281952d26e8fe0
zf80857eedde7b62a3aee9d8d7da25aa63c0c89b1158144f7d0e6d6328d0e2c43b566c936bb927f
zc60d1f49ba088d0655560f3060167516d2a1a417e2424645a1c33fd61302c3f7a2a83257cd5091
z6b7cf9060bcb260bb5c31269e58f8d594e50354aab0572bbff61cc091747e50fdd786a04f24fa7
z3ca7e0f8d77c841aef6236349405716d224264c337debe232fab43071c2ba8e4f6f543a3bc7b2e
z2a01c79a1b90416c69d67919da581b5ab7994391ba613bb1cb3b686746fe7de8420e1ae07e0698
zbc70f549aa2f0f398882b108efbe2a3e81351234f5f7ad118d6dc42698b8c8bcba7aaa23e58986
zae765403cecd073be1e131f410244a4ee1b871ed7d23d0096c970ae7b7a40c87a0f498ac60ca4b
zc7e343952d082f1202f017f05e786f426cd0584b9d765c33543f4e69611456a298cb2ca8593cff
zb9521e2d1228d24aa9f4c3aa2d7ef24fc592c62a0c3dbca173e2c6ecd340e9bb232a3afca48c85
z9fae6768dc7766fa02bf70a07540bd512ec715ad050b4f45b74ae7e44fef74c8a229be820230cd
zfdf2b8b3a4244f055b273a2d7d8f570409fee6346f2d3a236b134a2ab582cb26f3dda26f691240
z67c5d731a91a5851a307af1a2acb30d7f951a742e47a635b435f67f3ddc10eace6f905fc94cf96
z0837fa1d4239caa9936073c0d86f1728145834dc2907a3eff1380d148c84355a605c994ff2b9c4
z368972347479342e2bacb60d77ed2331ac217dc6023bd4678650f966039057ad1508eb8a5d74ea
ze325e3fb46c8a4236ff5d0a2d4734600fec923d96d46ce1b95aea298b8334cb71f8d7ba81f0133
zae9db166f2da2203e0273362d62cf3d57d60dc03f4c147a386bbe2d088a097463eaea73d661b2f
z4a6e17fd1376a99f54fceef062a41df0a3ac88fae6d48e3dba76c4ce2f9689a730d8f0bb1dc69c
zd19bc448e880145329e2463ad8b129d54e93ebb0c9fe0e4c0e113da242bf6ed39b3f12b4017348
zded7a5a4973743fbffe84ebaab6c212909b7e11e73464facdb1767714b2e917b1e3baa07e53463
z5c81223b2283d004b098fac6588370d70fc1c58fcde81a8645ae2b35cdf1147116b0469391307a
z5c716d4d371c5db5125b5073717d5bdf878ca308ab20922aa5b0c41388aa0876b5eaa3e50916bd
zb83a6a858bfa8e40bc78764f23b86604b45560b2c45a1bc9a0f183ac49089d460ed556cbc729df
zf15960f49a2d7cba8cea11c77161c37c5148dc9f9a3efee2b14048e343b7f8b37bc36d0318031c
z0ae1aec40af2fc38d1ab5d52fad5f108c27f11d90340b91ee71a91d1863faef1716cd8056c95bd
z0742d78badb76efc534f068653448accc4465d2535b8de871ae9dbc958040161aaa6ad4458cabe
z84919bc7eba0da9bd83b7391a4e33cb5aedea4f9829aabe8f323666a25002cca0e422c0d1f6230
z50ae633f34c5cbe1229c873dd858dac938fa9e6e4946f3a78d6186a2ea42f4bc123fee1b997030
z156fc39f396ec5048e96c8d35a5146365c02130964f93b5eb2dab74d8e4298bebb8032037d3245
ze77afcb2ebeb27d7d24356adee414f7f6bc8949fd1f9ad63d1172206b16c9923ded6cd8f1cd609
ze0f0db19e7297be1d90e588b2b48057a03e9d14dd3f49be9a851aa7769ae2e0a1613a8bfb8d551
zbc0d789ded622ee3b52dba26a8cda35a857b952a569a1ca919d6f6f19a690a4fa837acfc994d7b
z116e2e6e34b5cb400517c8876f53e63ef9ebe2b6944ada9a4ae76758e2e0248aa41a4e5d372bfd
z7ee661fb6125734c04d6cd729343640c6d16fb86dbb772528fff553fd21020bf01d3772457a4b0
zf775f4b71feec9b0658c8e65776fdf6fcd77dc9a6cc05259fe2c153a2e7be37d3cf699ac508ce9
za91d1d5e44944c396c73276201d5993db8c6519d89e0c846e4365c9c5f48e9355b8d8e9e1e0b1b
z078978d2ad67db140207559b06b0db6bcbb5289d63a8c1f531768981b3431eab1be199affd98d5
zd7134ff37226a5a47b01d6858c992a2ba7be8780a939b9c0770ed5b72114004527ac9778992cf6
z73763101b0fa264b17e56fb356043d4bc0da8a93a18351958a4255aef4bc4260b8803cff9efbd7
ze10fc3bfc265f277f3296e0b55e5a011ae6acc74aeb992520e83ef8732630a4339cc5a22259264
zb59e175b2bb42997ec811d2e2236f6681553c35ff8a66b13e4a917f4699c5f5daf37e9cb2fb4a5
z3a78eec026bd1dc14a4a0f9114221dbb3e8f16f33abe4f6d06de1f8dc73952c9abb7802407aed0
z004ef2ce2d034733ec5fc61d9c9f220ca95bb3fa7e74ebc202f6b4900974bb8cd7674cad714618
zf15fd8fb3fffbe2a46d32419cc53e5c548430ff908af5c22f40f8c95040b022771bf7c762df41e
z691c3127fc8e1647fcc4f49b9f4d0cd92462b82c963a63c9eaffbd0aa70557971d82e4b65cfe20
zc45b1f4e8c14baeac9d01fd8825c55ef720de119cf130d9c78adc060852cffd887fbf8ce5564b5
z4f6d1e086bf99534c98082ada0e5209469246882c39c8b049f95a7a0bcfb0655801871e2a89479
zebda927015777604417fdc02aea2385a62c693725223dec54e9462c6eafb5c56cde29b367aa50d
zb6912d04cf992d931615b782e2c07eb6bce9c61e2c5d4ef13e894dc50bdda05f9817a54583ef00
z5d372440200985fdf98e8f82b4f1f9c3362c6caa3a6e21cebf8494d14cbdc5f325c2efa9f87abc
zf1b1937ef11c56341be676612f4b135362840396881fdc15fbd687fb1b43e00bd40715c3b8bb7a
z30e1f6f92d017aa9f9076480d07ae0a99840d870d3defcf7383616ff6ba9fb23f1f9e3a4ab1baa
z944c45bd48f266dac9e3cb9e2af3cec7e3fbaa1573285882fa623abb77b217ed2d413bf940f8c4
z6653834d43f428a041e14a92d702084d767d9dccb48b8500b59c0eb68c07d819268133203cbd5f
z3bfda8d1d7c78316f09fd0c4edbb6afc886584cc72498a7449b05e54941486cf198e1340c6ad0e
zddeffa94a49070ea2aa124cca15b59520971673d32415df0e3f87c9a8b5316fcee5601211d5f84
za8715589caaee164a1517fed25b3069cbaf78b787a58e0f54ed93a4385576653f5e9518b30f64c
za1b5207d814d606ca34b8c666989a21e2e58ce1eaecfe2d278ec5b7aa64c6f43e320e633efeafa
z311220dde5ec0434d0a3977228667f42ba84ab95236c3a47dda86f6393b2ce7e8880e23a5cdf90
z01c0b42b1bfe1d65d586414a481eb38dc9740c473782408f04f45c9da344c12f39abdd34d44d16
z0b988bf4aa036bcf686cba024e5b95948c0615efc9d7c47d46114152013ad87112babedb8437ee
z6e9416da6739672c71e75e3a100992f92d094e33f2bf0cfc11f5ddc1f8ad92902c7ec1f45967a0
zf69f1adf0b9d3abd3ba253a2aa4dffd7de2c927ef6ba9ab430db86cc33e7af0a678d785cfcf78a
zdb05c5ed753baaa752c485aa278de3cf134e3c8278d2d3869d0d4f7520c4a19c1c1df21c84e5b5
z9f8d0a16128417845d09f4bce63f3e42c19e7239bb372fd092f7d528c0384d7ccca1b689d68969
zbb2527510cea4cd1fcda972c0da06e36f50613e51e7e2a9c03c49843ac6f09b448430f8689f306
zfd211e87ac3765f2041033e76b86a3907e6514fed02d48e46e5ef59b4ff7a2db3161abcba5b9c4
z06b378d3b45c2e538c26662fe4026b37c90664e6dbfb72f36db4ce9556af1b0e4f00ba9811563d
z95c9c25211355ba56e00ff422291ba893c0eb730c3904d33e03a1cf0a63fb2e5c7a7eb7ff53786
z2efb105ab9dd981266beb9d906c57612457bbbbff2df69d319f856bed3c9381cd845edcc721cd9
z6dd5b7f7e670a87e1b5ae858d54137bd8ab6aca78834cd85a0fae20dd104c6b919f4a8f5198b61
z3dee1603b2afe4b916b66704cac2a7ec11142b7cf8a6f0eb96cfeb36a926bd09ac34c638c05372
z69dd7dbdd67248feba1ba3ae2d19cc1be967d768d025a1618a4e031d986d46859d571136d52abd
z4e55b3b421b0b5e989db6660393fc1b9faeb1974f575e8ee064e4767745be36b6cd33d54349e5a
z8c8d3d7a5313af2a7f521e2fba6eec3e48ae1d7d683ef61d3a4ff8c2dc496acd73fed0560c03b0
zd57ccc09c1f15ca4b516ebc4a800b64c0bae7978a70f7bb1076c0d9218f8cd78de146f6dcde83a
z0b5ea97303a713e89c6854c134929002892424dff435173d5fb0dca50394d2244ca2adeb4cd39b
zd3a12f3c1c5ffa5aaf2320a80b61d7e464386e5e0fe080916f7acd48a8a18bc2c4578ed5151bc2
z652ab13d833bf0594690387788f9818c14d8e57207a1664cc501bbd9a89443f48a7afe63856b57
za7a4587c262234b14d225b0e0a5fd5bd5cdf8620ffdbca9a863f6b64480d59dcb8f281723e74fe
z402dc2d28e3d8b2986ef6fd96064b74b72877a970c64087e79a523a066d539ceeb3b7fda146b48
z61d89fed56a17599dd2c320233cddf0ed8516c6de72687d9f93fea48036000d4a689b50360e20d
zf01491e942de7094ec0a72eedf901ff9e1655f8c9b0227840be51940576c0adf7ad741a53708d5
zc355734929f3e9413979e6d54912e07684d7b4a95b4b41e22952ea3fc6ac1393cf5b4686ead811
z6fb016a81358c1589fa27c9f9d4ac94e893105cbbb5af7de77de9d2c0889c65b265a403bc94eb8
z48d639da349b3b157cd75dc9a903b25514d922bb5a56e4263b87d088ab380d632c4d14b249d3a8
ze638b0f66245cbf2f9c04e7090af556f110c6f252f91e3c04c02b471443c2fe655aff76d0070c9
za49aefe7c1c2d9485656aefd1f52920ff052d28e48feecf06f98b249c64f09a01faeaf02d855ec
z970f26aedfd12f98bf2206354effa616a5955ebf589e8066755735bb3d3ae987be63ef2359ccd6
zeae4519eb685f61f3169115342177a240f8ed749dc532aacc94042a4be4a0f4ce0cdf05e9c8cad
zb4365b0610d1266dbdf31ce8218ee46984f4fa7831cacc534b22bdd8ccdc0ab15eb271f2ec1482
z88d588ed49cffadaa5063691be4bfcb79bf7d010babfc7351872ba35b935d4904df6b25997497e
z4947ecef616e2782d8773f3d6d56b375154e4b8f6d8e28d71f7ec254fd695360878037c92ba4e8
za1af0635cb4566b9670ac0b64ecae86076faf36b1d8797ccab8547c3a706fe0def978edc309a19
z5d63faf2b3de397902d253be8d6599a3327112977e40b03360b48ffcaf92301872113e3599bd20
z9b463c874be95ba83f351ff1c6fd39f19b5b6283e7aaae1f9bc060041fe0c471f2be6405ff9bd6
z93fce6e94fc7cd32b0011dbd6c6a0edf43bc7808f99f9063f823dad675569c06a414052915d978
z9c0df0b147ba782383974619f9f267bbfb5951a2376c6088ab5cdde19ee93629d845ac8ed061b6
zbc16100fc5f14fc64cd2a8fc4ce000b0f4795962cd8bd286ae3eeb9f7014de29e51acdcf800771
z50cad08f798c8e4435505708403f0ba57f3e9c5b12938b6839f49c2d8b0e006f4ae3f2ef2c2c27
z78f9aab1fe1b0632c693b0e9217d726f5d98d3af0c8d2522387ee87b4c123395e6cb9e94409f61
z66f86c850d0fb7e58028892513ae82b4d1f00bc61b2091a600be1f0b1da703be08d1ad43b2e0ab
z0f8c3a08aa256eea201baa26873aa91a32d4d8b8c247a30510b60b8e4369e1df8cdf1d0f9ddc63
zc0261379831d90a77c1dd10cc1628baab29d49cc668cd41d0d026f325ade71f27ebb54d106319c
zfab04a6141cf4a21ff0ba61607b830662de9a51a5664138acb54d8f40c43c8c0d60cb50cbe88ad
zfa7b5358d43c30eea1b1f98697323d2a4fe5d0f76e62cdd5b8ca6a12c6fd8d10f5368b8fba6643
zbbca6dd7d93d23fadacf54910158ae2fbd078f0d8d8bf591c8991371c86177049b37a45f9500dc
zc8b3cc5c226d83263c0b02be0f6b47c35fc2aaee78a3b7133e9a544520a6555b25c3fc334dbda6
z332558803186bca29c37d8baff646acac97c707cf4d025863faa9f62e817835e6e10f39d519237
z90cffefcebec19c10fe6352f35b3d843eb951662ba620d9da7a4cd216f98d9512267cf539f8864
zcdfb4a9f2ba2291ad854fe9f4e4ed52104dadd9c90765840287f4e10ad49b23ba05328bd613f96
z41213c44e14f6488362824b0121a836608730c7a9725d4689f0c05c535cfb4cd755b061c3ed2b1
zd2134b944a5a60c67fc0e2a98c5b85305e4a4ae9a955a7e9f8815ecc5773b57ac44619fe75a033
z35f8c52cd67ccdc57bb4f523190637521eff45f7580118719ccef665389fe54206693916402dc7
z3a892cb8e4ccd155a0764f6d4a8ca981cbb5b472a13c4e3419f9c5f2fbe2ea0dbc84aaca6f0ff9
z4be9c7902d0e5d12c07c6ad9438ff250d52f5f9df68de415aa45072f6a6ace1a0da9975d6784b1
z8c63c24d78f4fb541bed1d828e419ec4abc0b657c38d7e6a19f23a29c48e4475f1ee03bde02c81
z404036350fece5c98d9cd3fe7163076ea64fc0a59bf2fb5e13da7b6077504e1c112d03c33e3ec1
z25a8888a5db3adca57614ec42ba7ae7c376f5e805d89e653ed9899ce73ac0d6b35aad48607923f
z11e864273f355c0c060d18ea10dac625da32e37262c2483ddacdc25adbf20036dad8b70d1244ea
z5c0290b579db725dbcec2319915772cdcb19c1a7eda144b0c54f45fda56146b004647fa6ed73b1
z0cf31539cf16ceed011d1b71ee15fff3d3d3b82d3d9e3937609900b989e6465b96edc98d72a389
z79b7992401f00d487b6433209543b6a456ec48b3a9e6e7fe1ca8066c9ad7f31ce6117e83c475b8
zf1e77a91739e05dd9e4957115f74919539f83593d22fb6c120a2d4738342e106b5d980b872e20d
zbf92b914a6006e1c84cb25e7c3f324cb9b6c8ff1f0dfec80011a2bd9aed221bad36c6bbbe8604b
z2853f5956b2a8abd54cc6bc887879bf0cd845770f80fafb3128ae44dfe3217d4567c7e794e84ce
z7b70562d1b75bd83383241e830f8af3e01e2e0a9505eb350b2233469349a66e6bafafa307123fa
ze2f4aa27f0559a81a48182b9e2e5a4855f48989e63b04cce3b124bcbfcd4d5d214ae7be43692c4
zfaac42316cd72a8f6d101dce207b3508deffd40664aeac8008842d9950ed201be984831ce8cb7b
z78015ff1ad658b5a89c7407fff30ece7a2855506d8ca3e82726e1eec3f99d7ff0fcc82ebbeb30c
z9aea02ae72611308b9ae51ef3f8fe8679b40d8efcef0f059cd2161f3654eb6a9b843923a3763b2
z90399012427f14f500349210db245fbb58afe6129aee1c7842ce3ead110acc17a1834c493bf26d
ze8a474bbda237dcbed14d8d528320426b63ad46f34065c8f37ea2c1792ed96f5f6e1fb6ec8d308
z5fda588f42421d251a5fbb0e7571e0c835d770537d606515205080e1d4ad316d2ef04358f3d493
z4f74d690bc10f82cdf8ba0a12cc45461475a2bce2fb82ec636c552e292bd760b835d1b182a7b60
z8f77adf07a0c3779858cd235c9a036d4193cb9d4b225809ad17195554833d44701a709bf6d8bf9
z2654f4ead6d8e639361d78793766b7cb3ae4337f4ee916759662c888059d0e44146a5c8e92d99a
z9aede8ec3a0f9214e646c813ca21ffc5a7b9e08bb24c304a197cd16f2f6ac50da4df925e49c0dc
z41cb1c9bfbe27f922911b264691b39f467780c661b86d4b23f2141c711979eb5101704ee4b4ba3
z13cb4034f6e123313febced2e40ae3d95905439086e6fe652e47527dc0fbacd2f93db1c22a7bee
zb00028360f6e429699da4175cc6cc9f0827956f12fe94c096eaeec019f2054159f0bf73ea28c6b
z34a9d4eb51c6245a18b37e7118fff130eebf3bf007de9e2def7a79e170b5f60be058072974ca4f
zf38d8d3e8718c10f06e65dd4fda38232f876807505938d97daa70662ff2c12fd3a7535437a122e
z530219d03786b2d1e4b58c7be7260fa11065bb5a2adebb73f5e8383e56e65a5451860ce79494d4
z4d1bc03a4bedfda536ca4ba5baa0c90b076ab14855f931dfb8dc58b54852db4e68fa5a74608b83
z9aae7c855286ef455f723e296363a170646f53d6591083f276a7638dda044266b0bc304bf7d99b
zf320eb3193499161e6f29e21173b27452ef1209aefa8aaef15fbc22420e944740f1719f66a53bd
z5583528d9b982c40b92fe0f566eed0c9dcc73d8bd62f00e17b8ff34341ebbd15f30143fc5eeded
z285f9003ee1653761588a463f690da58b3721a220f99ab0b043b3c0860f226764395aa8b221aa5
z437d0e5945e0efff10a8146c92d9e6e42dbbec7f02a3b06ee7dc3230a3f0bd6856fafc3dbc71d4
z732cb3602e72dfa38d280689ee6537eb6d595fc530ec8642aec9d05452f82fa20a18ff917321aa
z4adea9f8ed3fe09fc5793570875049c43c755abf1975d42a6552d9d771394dd31a39a743e90f0b
z36b1804896a11e364caf1ffdf3e626d151e8717bb1c0b9f3faef8c1c99adf4c9efc8c3c3a0e782
z4ce35f3f135feac356a8cdafac91bd8edaf0eb8c4d34851add21a1c36b4bff9a6f197a3b8ad492
z6e0abfea1db473dc2cbfc69b51d1fa955901b8edc4dc3d00f81c906c8600774bdfcb9bf6cf6239
z9f504cf87b74ecea33e443820dd78c133df8e3ef252fcbfb947b202a6505bcd3dca977601743e7
z4cb1685968d9523d46cdd4838f6a32bff08b3daeef1c98a62380511ff63c73e17440a123b5af3b
zbcc366f0a926372105b3ecad270e2c8dbbaae2aa98356452baa21d37c002899f8fef9634166f91
zc7e030ab76d1b33a673bf346594ae1e2661a13dcacac630f12e1dfe20abdd57dc40dee14f827c8
z1a1f4d0b3e5326158a9e6f40b86aaf545dcc9743155cdf08787e87ca63592c38dc1bb7bc88475f
za753d2448319bab34f19b0a370dc831c9d597da1d23cd5d01739ebd3d3b340d03bcda800eeb9fd
z9df222323014fdf2d68d12fb95772d8e312335913ffbb6790256a37690cd4ef4fccda23660f901
z464bd21fea822d32adbc04a9ba2ea16854eba76fb6d0e28f71504ddf5f200526b872c402fb1e1a
za90cc170f43f22bf5a09cc201d284f301e2213762a4f238c05a02803dac6c484683afb8c8ff77f
z402ed8c9a3693de637b3e50018b5c4b82b39ca8bbc5dc5c2ef7b543fdad357784cff6b04cb65af
zd8a2e4d94e0cdd2dc21b465549e1cd675907402ac9fe584d675f318a94dffd9d5d0a08d4cddb49
zca35d6b7b5c1114496ef4071af7adb4a4a419d877879df69810dbc0a891ba976253c9cc4072d64
z4708b2a4a78eada5fe3567c7c877ba4d972e10a2dc0aac499e655147615c74f1c85a7a1a608503
zb8f4372d41404bb1315b8fdde6dd14dadca8d42b60967ebfa805909f94da00a054f711637162ca
z37646b478e02165e8a40116660adaf2c0858c510e85aeaede4875c75d34e9e4281c926c7dadcf1
z433bdfe9a6f192e514b1bb4bdf0cd4f2fd3651f180641831db5355ee720fbc09732bfae28a2b79
za93ef7ed85049aa6ede3918872741e682f457727ba93c3b9bf4655947b1154fa8bbaf96e8b459b
z2d32e6a78abbadc504ebd4d794add0ae221583e5cabc6844fab26d8dc13c8b7d403fe04fd19464
z987f95d3e39445568bbb26e246676e4a61ba125a6e13d3cddca8408af1decd9e380389f4a7e678
z86511a554b708e0252516bc3f1755483b56938956cda61163611bae5d75c785ea44b6098dfbf7f
z830a83e58e1daaf4fc79644b232b67955bf78c5f433a72f821a2c8790fb4b456cef3a651d8a02d
z095ea6d1fc18e7f0b5fc15a01631d1facf61f1634ceee0ea27373d1078c10bfb5dce5e7d9c411c
zcf94da8fea2ddf491b3b57513e0fdf39db14f4a78b9de32c0851a35d1e6e83acbbf298d19d8a47
z2bc5920f43142a8639384cf8fc458ae2d8852064eec71ed162045817adfcd4983a374d7d6d1bd2
zeb567b0eba4206f88ebbd3276a72391aeb35ce613e191a07d943d7ccf19d1b6130ee583c110750
z37fb8394a1c7d2b65741cd8413d9508c714d3587f38a9a6398290f9b4efdb7711053a298706ed3
z917aab96fe60f0e8fc5e46b22262a90c99ace61f10d5d52d56e00ca6bb9b0ef280500b6dec226d
z71ed052564e32081d8228cc667a62e2c7612051931311b841d5f1e8008479e939425071450fb7e
ze0d4981c57ef97f4c5ace3b14a754410c7fe56ac907df85e05d7aa009ae19a835c0bf5f21e6be8
zc5d6875b7c46cc018328e2996929e96c124a90a888fb37bcc545cffd008a31f025441cd1816654
z7ee2f09f7e0bdc0c386382522d80479104d48ff5f1bb615b56e160b2e4a1f56fab1e17af021648
zaf7cb9879229a86a0a5def486737ea7f5ac7fbf9d6c5e457dcd15b2eead798f590d01510314c43
z43380acf7637223982fcaad1fd05475a3a9abe46d7118327223aa143d6f14843deec4be0a6d285
z3f9e8adab21936b0e9609461b18c5051eaab51e3d80e135dd2f2ae68795fa9281faa83604d9f4b
z2e9204d4baca504d4e48b084292b0887d7ed0ee82a94d42773d7292b50c6738a3108015789199b
zae80f30ae64bc777850cab7facdfda83d2f0085a5b01ce914f9bd5643b9362f9941b3599c6b6d9
z4e71d428aff05bd4bec4aced13239c4c2bdc74da2bf4c59cd601755e5a418d789aac467ada5c45
z37002b9a48baba9a8b65601a2abc2247c3779c3ec6e72ce7c1af068f3cb8a05bd68cd5367d96c6
z87316d17c9e02e8290d7b9afb8e0b69c4d9bf3e008240691c31632615ee486cd6298d4902b84e4
zb585a564cefb890f176d17afcb6b8f1a46434e5d0c257dd86875d05197c6060920520c724989c3
z5663f9b859bd2452af2db3d3ba7facbd69f3ad479af307fd6bb78d1ea0b3f2d6093695e9dbdc3b
z6a6025afbeb8b64c7b476084865960c6686904b9142744d3377fa9fd6241102b516af92cd38c0d
z26e6709b8cebc12542af989d7ad483c9d16d368c50faeafd561d665e4a0594fecb8ade907b80eb
z1162d6f1789446e9cca239186d24939810c99e7d8814a2ad0dfe86e1903f07f79f9a9758fd718b
z388c5872668b8b090ba7fb7c0997293a7ca922b9ea1925f6b6e0d1f4ae2b34ab1e0cf9f7175535
z86a44953d5d7be6bf24fd71b46fa35f08193771da3067d9227c8fbcb191499d546e1482c1f781c
ze732af3c648cfbaeb3de1ebadbbfe431cbf75bea35c890020cc5ecf63b34dd201e41906d47c269
zdc7caa55120539490aaec2e7c89e4f2fa5ef472281a10f8f7cc5d5af562715db5162ab15ae756a
z6b98e96c13442fa62fff50e6aeddbf095d6c156eaef8ecf546317c63f07d795a7a69f11321496f
z794f8a9d4c6bd8798fbf6b243f12b0cf562d1cffdcd4cdcdf452dd2d9566cc094f3a07d637f83e
z64548b17fa0c1ed348f2392ed5f758d22abb431f12b12d4a23c9e072ca7c3f6a148b6131375688
z69fce2c5c7a1fae511974f26e7993a39602cb515f2ef7d81c52a3c824043b373213ce8f51005e9
z900858b38d0917db579c1d944bdd1e40f9a40b93e565c45f24f937dd7995f07e9c5b4e01ce2763
z89f073131599faa6d26902bf4ff5f37a95483554e6976ade7e4ea5afacaae2a65ec016e090c0f5
z503baf558a97f6097411d2db790c95329f97611a1d110b22b78336c827d44377fe7220b8804bba
zb824fa591e0acb1c64c7fa2463623c9796588c39d38508f0b7d15048c681d59271738be7fe1220
z236f6c99f0b182718e63c0f4934c774ac67d13043506af5f30cbed08745ed4110f97699b7b5d45
z098cb76fa063afd0c58cc65f791ba921c7e982a5c3fa3be6b29e4776d52306c054ed8f990e4973
zcfb23a93e78271c6f1dc19348effb8d948c4b20a1179afcd649ec86d2778cc29145bec4ac5e948
z12172b275fa93d74e39c4430df629b41041cd2c4133e89434be3deb99d69a9ca4131ca7f3a8c15
z3e5b84414579813f3e6b52430f88cc67e26c7d999106e4fbde1631e1c017b643371e6e7df8c881
zf506451357d457f4c1e7adf79f4883bf6044ab0ae9ae5c7c2998b95ef955d1829d063a51ec6692
zacbced222f07a80dac2e483607a9a13a581cd0496b5a45317118a683447c2c2143aa7f6d26885a
z8eb7c842cfa4771d956f77b77f335511d2e2cb1b546df7079099b916b5629ac4669f48bbccc70e
ze8b57fcf1c3776af5aeb247a2c9cfb1cc38f17e4a4e31e52843c0f0ef0d043a5e5d8a13115cb7e
z03a3002db9827f0caa0e46429be7009844973a5a3776f767108cbab280fb06cd0d5fdd59e6dd2f
zf0a75594ef3e1501674509d8f26dfe1c0e55149b4ea4df001530c2c6e91f6a7d3336f41dc45533
zd8fc1c67f9a07c78d6b8f1bf7335b3c9a9ce9694ab182da678228416634306828b9b93caa6f11e
ze078d3e522c4d62cefdde9a398c4bf6d353d32b5a43316e636c8c47f809fea37ebe3c1886614b3
z6ebbe21ae8c15542736391c602854a7508889175f436f518c9e7d41b2bc57183b9cb99350dfce3
zf89d6ac552d8444f7ff9c68d9c24ee78b287b27bc291f85da89476a3ff136894e5d8e308a0c117
z5932ce4c791925f49ae7a66b3a1b9a30143024f19cd52534bad4f0ad309b6d519a1b210f48db6c
z8b2751496abbafcad418ca19fda9e1e186c80502fd58ae2889ff8a45d5723aaad56ee1c6c6eedf
z208d3ceda5fafbbd833f0e581d8b974068e01d607e4727e843694b75ea494688e340b73e5e4e1e
z1ccde4945977f26e01e79b5e184c2a6e2f67313551ef623b8c5d758ff5eb16080c48f997bc2823
z48725d26fbead619a451329b108af9751cc29107071b54fa3b03d950e796cbd65437b20790215c
z808761f4cf94f166ce673c70e24a18b893abc57fb71de1395585ee7cc6b8719cd8a0b9bb834b0d
zf31cdf288cd25dc3d7996d640e4f986ef3c43edf5e9d040e7e8af3ea124ba44a7c9e8ff52bc0ff
z9a4ae80c62944122812bbd26c599d3c28679076981d629a6c1c5f3ede7de31d9c48da399ed5f4d
zc6d8a15b54798bacd8dd75e89ddf457dc408a0b1deb6f00ccb809a7474634c7ace0b3f1ecbadab
z69625f611dc632be9238a922990ea016855d16e2c45cc75da5070a63bdb7e939036cd3841adddc
zae1cc911c2c93de5b1f39cda76270b95f51d31134694e04cf5defbd6ca294245c2f3620b514403
ze918cfafcb2d89115e30d46f3707e84c53755db229c0f84f2fa1dee6e610b43a0455c74986f270
z0b18cf910cd19ac64172c0d6e32760396055d8b83d117743587898b4e468a4b8bafa9c49b65c8c
zaa7195d5513c76e78442c48f046ad66135e903414b15689f3288701cc4d57d1e6b5f445ac9d4c3
z33314c2b23f67e12e0577956348e0cc5596fbe70c4a62316465f74400ac6e77d0a0a2d4e02ea9b
z690ef4869daac9fe38c849c51bcfc8590efdf0754760e6a0add106687d1d5bb2ff14d909711bb2
z97835791f8bca047029b66839d461a6855f5e6b4744bb4f2fee43c0c98fbd789104a09cc5d1374
z209090a986252ba55cbd4995896706b3041973f256c2784ff5de0a5a2daec3ce88ca9d2262c021
z553e610b6ef8568367cf6d0f68f83a79c357070b060aedb718d5a8af5462abde14cd425b34793b
z40ddbe58bdbce0bbecc9fc6b26ac5f7ef81df0d7b80c24bbe082de63af5c728706e32f25966bbb
z1cbb8fb3df43d9d4014adcc533083404bb08a9d80576201e7ad32400a1b413b8b50fe217c29604
z78be8f70f93c41c74e31d5bbf44cba307df399bb325c0f6f61f4777bf6eb4b2bd9a1dfc9c6c81f
zecf8750fecc4083f6f0cb2a4cde0dd958ee01ee390d7810999812040fefa7fb8000a824cc02a03
z894612b7523f2547140d6a67676040faeaa9305de301447b1d25bc6c9e6f886c30a18b20a6f4b2
ze8fcc83dccd5e1d94f4929e6f2a2c0d03339947cdedb1df936f222352ae6d3018e763d394a1cd1
z85fc796542ee1db74ae598114555310a240ff785e823244f7155035683352a2ba1b8e344320c5f
z528c9ae70b69db5f6164e0b567b2f0f94607b96cc8387f7f5a52fc5dfdfb29ac63d1e95b9b9609
z748ec3d83076985e5ecafe53095810e015b3a5aa866a764a3ec5dd4d653324907bf59ff6f01123
zfa95d6718a97ac7d98065d2cd8790dd38d4e9f80d8599eb0fc383ef099bd382926c2df645da738
z4a44cdc5341c8f00c0edf7a78f2e64b35a2167099cf7203e83882e57e5d372e406df586ac24836
z8bc204c3e0dadebbaaa7e984ca1182d68b6bdf5e59569893918de4cdcad4f790b7f3b6cfe53607
zf25f1923eb86a588dfacccbf5c3fb6a2b49f6053c7985634b1801dbefbadef5dd3a155dfd7c2bd
z59fbf582c26a033f910e630df3984cac5c9aa977510c853da4348ac4bb41bc2df4f6d0ad28dbe3
zaaa45b01f57edb6081ae98035dc5489bb1d2bbe5558030ea03abf855df0cec0dd16c49b681607a
z7698623fb2a87b637b6cf4f8318b1382eb2a6c74652488052e0bea2d0955097434cbc69e79858c
ze5656896b4d4e59b8b14add88206453ade0a74d5b7d15c93e54040506d395422373c89801c0f87
z5dfcc06ac149be9e80748648bc14366de03fce41a8c3cdf7bfc6045341efba00d9ebc17478a5f8
z4ac127ce57e3bf4d612d80878cee06d3dc8b572c5780396797893a8079f454833a7f4fc8093d7e
z5c10f9f19332b94bffbb39894b9651b6f87f4b9c38f71c814843de2d17a54cc25d29e94fa8ca32
z5df27e465607945801f58682552670ef643be0287115c7d910189e6089caa1c7cab8246a086500
z979ddeeec045ae0cd29faf2126e25b0158024c96c26578e05e071807d76ef03e167b672da66731
z5318b6ff156f60cb7e76194aa69b794c12d83631adf1826f07c852e9683ba79fbedc522b20d385
z29537be8abab3161c0d7b55992109489d7bb78acbfe8d4ffba95cc9333289e7b9732ae009fdad2
z3b1867f2878070f61c4e35c165bb1f0ecff93ebbb00423f18e12a5fcbf8f7f3db8b80796624d81
zcd8a97e874f8fe4e82a94b41377bc2fbabf93f84b498bd28decc4db56c61c55b335cbadfbcd625
z04fc9f9d4929e17c81590046ec3c40dffa5b662352aa90594bc431bf78e405a26960f1444f8eb7
ze507fdc6e24bf1a60a827848b70e696941a1801d48ca51cfdfe2cd18502b30107488c11070d6eb
z796e7d653ac9c620452ad15a513a64e3a31d04b04a7c6585fe06494521f001db1d55f36979a0b8
zf2bd90327707a77810c96dba48389badba6b3246eadcd0ad1b9544a9e4a05d6f92163d2dc208bf
zb284930634eca38814c482f602a7b16f5632bdd5d679a0ba4221a61d7e8e373c3cb67da7cd06ed
za95d058d774b658abc503c201c0129bad3da38f4d4e1647935835970e621383e24a19f698daacc
zcbbf3c807bf7ded89ff279afec0c6db18dc3a6d69ef6e24ba38e122e8d4eb89a074e19a219ac8a
zec91a00ea029a9ca8fac644309b2dda49dccbc4ebcc0824847c8b8332063e761b54b8a874001c5
z651c8d654979329e5a83035139ae1ccf93d51d8daab02bacbdec19ceacd2035c517414c9f4d316
zbcf7a275f9154ee4220c312e611083b4e7d71cbe26a8900394350275fc0b53056d6e0006cc95eb
z718e979b229438399d631844f8cad5fadc4991347318b45d1447c693ea32cd310dbabf41d4818d
zb584d20155e722a320ff6443c6ad4980f3b36a355d683fa4c018e459be3c88463b6b1658b61c5c
z0dcd31a07a0aabc42005156c7c17a751a3baac8fa88ffb1a33871b7e5594cd59e697109bf3f9d5
ze64a820549fe1fba1fa34e3e2847dd937fa339ab073acaf3c294be74414618536504431dbcb034
z241ec7a82b1ad68adeaca2ee2d885055405ad1f436fcb01ace050e9f6bec621091b286a6dd28b2
zf331b9c0089868cd38503a89141c688b57b46e3218dacd0c83b2d5d8d7ca1a157fbb5ba27942e0
zd70467bf362858654504b97a388a3965b709db2b0bbb0530c1f0d1ca268b109e89ebeb70972609
z08f53d64a81469f724a57266061748f2f3792071188d68e11f425044b23461dd39360c137642bd
z3586bf19f9f86677090855cca4cfa5666f8e2055a7bd6d5f852fa7961bc9fd85c86050f10b1a9b
z281e3d123281289cc247b4d1383be08d6efd56534593fe1dc6c7bd1baaee69c36188c9666fb0c3
z3feb27a58e60d09c7fe4dce125689771f7edd5f0f1b5fbeb3ec360dd2e9e230d41fe3a8336f3f9
z445e386a27bdbe9fb9b60a1196a581e5e2e3f34ec6bba8b821eb4198f1868c78c509dad7a14ee7
z837c13b0aa98a569c6c233a853c0489d1701bd76e324ea45daf5fdd09ecf8a6a7278c2ea9d7e21
z65cfc3dd11004e25d9432a6cfaf9ede25d268c78adf7b194b307cf4b3c64808287de2d56237417
z26cc605670591222f43b198c2e724796042a2918f8f852954add29214103358145ba20f80a770d
z523c9e1e7083dfd3f8c7e6639627074f31aa132970b7ee2f51285d3065481aea390d13f61c01aa
z922341a4c9f51b351fbc65c62c9006eabcd15012402e829aebd8af753b9a3435ceabda6c9f813d
z3e6c538e811af2f6b2676bfe6910e1134d4aa823b1b9371dd433b293c313e43ac9a86d0f1b9a63
z03e4fd8ff41c982f0a74b64348f9c3f4fffcf79964a8207d5facd1ad3c494cd1c34e1b33d5e009
zb772c2a2ce21fcba59e761ff3a0e54752370ccf6e203b8f453e5362b669f6c79784ef2ccf0264e
zad123327100d43036081c14ce3b87318800271417ea16eb947a2a9c1c5db548425966e659a0603
z609a79cd59e45c72abe3f4f7ba886073147b70d3420e67f28a3dd338bab375c7f738df5b0d061a
zbcb7d4b71376723bb07c6618ad2d355f41afb4ee35de3e4a4385d7ea5881b4a0a7623c465277c8
zcfaa73f465275b10500247563628dfde038c7f50420e473ab49f27aa1ccbf314bce4e8dc56f42d
z0b7bdc2e6cc2d84094cf08f0c1f8bf83ab44b4db4716da97404d01ae2b701cdd5dcd26e920f2ba
z38eb36b578b5e1830e5ebef0cf9d742361afb11a919e485b2bfcc1ed790d7757aa2b71512c68cf
zb26d13efd3a4e4e78b63084b87b3e99c71d40451a96da9d7e8810145c9f8ac6a87f688271b895f
z95f844cf2dd1571c4b21941ae91c286781cd6124efd6eb9348b70f6a5b12a9bf06932d3e6656e9
z8ed83d23d107cbb216c10bcf25d76e5b2581ada5e67bd4a76cd0db204f3c72a47d4e8fa510d4da
z0959a0723571c7d8be4b67683a8d5112ae4e2aa38ba5cc314be905390e8e26883e1e163596b05b
zdd6d67de38381b2ac557556a0736acf29c706e25dadd5a300ec11b6c01bc2aa2bc9afdc9bea1d3
zd370a55c87953d3cfbedebf9f512671b2884547c67649853b27438785ab3524443ad7dc8eeadb1
z8e1e8e213d2674f3ff2af211d2d186188239eab7014fe770b11a034657f99be35b55258f105a50
zc1d6a7fcfa185d52dc9cb7d46a5060bb798edc12c081e475a1cc755ce481b906846508172f8dc5
z8e38b961031dcfcf09579949c0b2052bb80e334304b817ebe4c2991b066f2e6e6b88175984b69d
z777a22da4dad36655d5b13698385a371a006949d5fdfd8ec7823278ff9d97331649fea7ee8408d
z9f41162ee4fb68b3330a3da11ac47bdbf9966b52be88ef97c66656c06ae27e7246529dd84142dc
z3710ef4d62827da67774609715787c6913a9d20d5db1350820f9bf90920d32d7d15ece43d19632
z9ba9e8afbc73f60a586e6b8be6aa16a95917210dd9d2fd024e0f2baa970ebb28612899088ed80e
zb5e9ca150a99f98897cf8641cf79e82c3deb204f1f44b9e1ffd2bbc72bdc1ce7479fa9c393cd52
z8789d16bf908b99900f5220f67bf7a833ffefa7404b4192570c6b063dbaef4ec6de0ebdb07cc16
zdbac81432f2bbd7a1cb1e7d7fddb0a59f1ad0bc58696c23cce87ecc4a7450a745c0cee12734036
z7d93cb0ec0022587ae874f4131e89ad692e93a352b4e37852d1854739cb71d1fc82813be70f18b
zfbdc5ffcb57ee7f2405672a9807950836d28d5fdb075ccf81068fd3259087120ece0d87c2edc06
zbeaf1125997f871d91401072cff24d8c79eda4f302043a4f26dd0c120026721bc80a838f8ec450
z9eebb802fb5dbad0c96f3d20fefcd9ca0c0eb5d649c15c00f8be7610a2d6ee5f03d484e7bf51d6
zeaee696cf7d358cd0f68c62d1e0dbef02be9fa648ba1ca005eb524e54bc35f5d30ab167c738f75
z6ba539a055805fabdac99b78674655a8a4da1bb02cde0fc15ff8afd456b4274d63f4e1bd6a2dda
z0dcf0579c214f18f7695afea13117bb606c347e40a3dd5d02237d2c4430040e6877091817ea564
zcf291f6d72667c448d749c866b8b797e8f06dc53e7ba36bbd6dddb97fc112e70d79cf18c30637b
z5387044956cb4ad851dc8e0aa07ce2d2e9ff2f60eb3300391cc9aa07779b91fc8b4dfa0a54dcc1
z33e826d1247d4bce9a718b83f33b96005ed4508ad0981f836cf0dca76a4be8757a735b0f156833
z8312eb4cb7c646e0d6056fc9fcea4721e18eb1fc0bc4db73bc05ff5f27fc0ae797462bfec03f24
za7c35f5e33772e90c5854ac18e77da735db396b923dd95a91b88a505a0d5fd9d653a8aff3c4ada
z56a47ca733a12f40c952796bbcb5c135eed1f863d7ce7e491f357175ca801d2b5cbdf487baa2ba
z3987b1645346a9fa2a04da7bba119550ec857ceb82581eb398237da8b212d32054f4a90fe51ea2
zf8edc2d311f60d0826fe5071135577cf62d3f5c65b981528dd38860ace06df24449269d9e52c76
z42421718590a6bad7085366185cc6dcfbcddf1626839f440cca0b817a7f5681e2267773feba603
ze487c2e09ce3f59969723387dbf118c6365e75b48a691a37a0a4aa43b22e9c6ca9ae6179bf7691
z5ff0153599d5daf312f14200ebb6e483c75bb0b1b85843ae07c919b092de6354080231a676bc29
z5faeae0390c363ca3375e97b76321a6fd543a573c6bcb00bf55130233603bd0b67fcab0fd5e80a
zc9fe6891d28868f4697726d3341aa9d9c8e7dcaed7779775888b6e73c2851a16ef5e3c1c8c0fa3
z2d8d3810203f85b36426b6bc614210b2c996daebe1db230826b68c8338da3db10f2b6100f823fd
z12f04adfa8e0ef5f966f8eccb11593cbda3eeb0dfb8782e4155e686b633d356214f13e3c230801
z064da94f848a6be74d179c9408cb4848e0f6959e4a7757780be0fb301bc857d7a2f1a2bb150862
z5d177cd3ab59e1b10a617c0a45cbd24c5f701191488e3718590e99f1669dac8cd3bc58ba523f6c
z0f7ce9762296724932b30c05cdb53512f1ed2f55df05ace1cbb6ffedd9019facfe501cd717490b
zb87737c73ebe738bf0847df6a406021e05e0fb5e1d5ea7cd64ce28e50660489a79699845359fca
z2df51bf9d67790403bc20453c6521a669bce0fce15594a089c4e4a9615608909611f4f02e37a6d
ze9563238f816ec108c807a8a8d8b4e1f0fd1541f4c13a4795fe90dcba3d37679359276bde1a216
z4b9cd90146bbca65c9ebe5dc596e750d6a3c23b8d091dfe4737456267cd7f39c888a676f5357b2
z6e481ed7212bc5de890b242d62c6d42daf0eb0dc482b31880fd54a5e2f938e1c86f506b3ad97a7
z9877d2032d89974075407fb7b6dfa256b5dd4dfe064ec0ad56feec22018982f3f4bbd886991af9
zaa4e5f7966f7dc9ccc09e5274ab04b1cfb9ab8190fce582cc14393551a85cefed1cc68e71e5bc7
z6c8ae33d89b180b5f358f45d31e25a9b36ae55c449a543fb2955b4440ec79f057d4bd7de7b2554
z4fb89e46ab564757b3bc6cc959302c6db40f5c2d6edf075b215bb0795e948b3e0f16d8f7803e71
z5e0c38b0cb1dd9ee1f36551c156af05de429753894da43af98245cd06c5ee7c8b1e34b4f8cec68
z7a97f6d22b6c8ebd2cd265650a62f553b3430e2e6ee11e635af1511e45b13c7a50fd851d3dca85
zb1ef4459da55a68b5712860a4a8d1a3339692bfaf0b80244ba7b4a84df0f43898f9b0e84217507
ze0e9c5ca9ea5ca58e9998f13045298c7cc98cb41f1639e53266b4d885669cd8316c5d0f3754958
z0de3a3708331870c75b8b45d349052e74d1780a5eb79642d888c798c85f3fbbf1e2a878e0d3c6e
zd653b55d76b9f0e841e9088563c8bbe22b4dee729f82effe2e9dc5e37d29231d4c05c8777e8cd2
z6f1392d8c55411725a37b44319ebeb28d745f2f4f19c9688d321f47be9a2913b6537d05bb29c1d
z5a56d1a141780edce52edf51098eebf5a7edbb1ff55519ab0f63a68d1537004e2df832f77cce3f
z0c8282263646af9c926805a8c8560edd723b0a7c33354e8e29a7e3f2778ac09808518f127fdda9
zc1fcf5a08bf9f1ae9af9ba90879dfe37d51d4b5cf6490257dda53fe228cb6d19e939601ee7f615
z4758c163ee0d7b272ae3f314a73d8db58a1007864d6c92a59a7a31ce9f992bb7b1d42411f2b6a9
z3514da9eb604208e189912d71c90164b91dbbae838abaee47ba6f41579da1369b73f249df595aa
zfef03fb9735ff8f7f9d3efa91ef85c34a52d6007f09b54451c5c0e14c92da655208228ae387fc1
zb7180fac46726492296fa787f08b2ae3de1a9384776169124816a2b6eec196be3a54d7832f69e9
zdd645bca68c0e99f07bf6517ad42c14160eb54ce03bb3125cb2380b2e570c3eeac274cb07f8b3d
z2f605c85cda87ea443b3d5e2a75d1a23e470cff54e52c21a62e018759a2799637fe7447b08acb8
z10485b438c289525b79c5e835c7872e2dd7556b9c489f905acd9fb6a997fe5e4f739c4f3c34943
z2ef2e545f46bf0731c4188f952aab9d7eebffe757290cd9ab2ccdca017396ee94d0e55457049af
z29d91f549776dcc95cdd8172b787671b51b838724846f4c38df50c60c86b1a4f1496c34c3eed6f
zd95c1e1ce4a0bc4321ccdd3492c1e63cc18c36273003dc10819471c8ecd0c31a87418980800f16
z81130efd331542e9a49523caf786a221406f0c1f664767ba17e1a82ecbba50bc9dd6b467bc7bf2
z45c8e7c6cccf06c481b2a0e44f311753293613a8d768cebb509f7afba6f83e0d0576828a6515e1
z71edc0f2533307d8928b88efa67dc6c561438658e4bf7e8e3939f3f9551d638a8ac8ac1031671a
z756d63ea0d676ed74d3b745326afd1cee4919f6a834b29843b6d19648f0f284c48842eddb6d080
z1238c60dd8f49ba942d69ec80bb3ace50bbf1ef193f8ea7ba44aba509cfd80e34e3d3633d437f3
z528114dad345703eaaea265b247a5186dc79e962216919e3660513d25111204bdf563b5712345f
ze27bcb47d2b1bf04a88ac5406d69d94f4bb8b7a01f85ce5cf0e420390b4238da00e885410baf9b
z7607612d77c57d2cf428f1effdedc0ac880c65e89b4b2f9b60f3b147e774265891c26e952b84b8
zf51c86eb39402d7686e7fc602a5de9f946e21a291828cb7d0b2a9b5ef9186fb690e0784a959293
z5d5620994b505097a4a4904aadbbd77f2efa85e9bac97b886c579f157dbdaad029addafe5d500f
zaa20c1215d96dea49c6398e6ffbb34cd68f1fc80fdce9a702f8a469f710d911f7842afc330b6aa
zca23341d06ad04c539dd6d514530ac59573489a621823103989dd4f3b3843891741a0a986b21aa
z2e09a330d023500e27d56b62f629d3649ccadbea4ba0c3bcda8788756779643a4dff2f12de319e
z2041732670b7d45e376c803e1a6809cb0e51261768bbd9f3fb9b008b588e12c0e7470d6d05ebde
zf6023e2b7e345315176ee88e344b6b59edd0be251a02ad91972d30290c284d4990d96c49aae0d2
z131f0564c5bb18505be328a2ea3f66963f370d2f30bf3a1b1872dcdddf9f98b5a893f918eceb4a
zc58fa41fdcd02817b2c36b46b0f675d73d560e4cfac5d8c4184992e72588987ee29690aa2caf84
z711bb5937fc728fa33dd75dac4d60050be954e9bf504f2e36e0b5b7c4f2d7e2e769015cbc67560
z243c9800e2d09bd11d5bbb22445a92696d8eab513c5253dce1926f3bbcf56abd90bcb13bbb0016
z4243a54c35c65a1781ae4b03a1476fdc15b33b5b904e5699179beaabdda61d9757541bdedfbd5f
ze509c0e2dcc1528d31e46e328e0dee90d7204d8239cb402075d209139ef6acd270cfdcba753209
zbf939ee8b96f6b01abee3a572b8e9cc87ac62b43d4073f8338113c8f49274cef10d32896cee942
zefb73b855b57504a8a42aad45225f8575e75a190f0f2a46c48ec54646464113fa995fcc3398231
z49c2fa7629e0bb21b228d21ebe3c26ba35ba701cbf26d223546abcb56c9ced103067e7ebc8be95
z2b7596981d3b575f94dd79c50626a6e94db0e7126935fcb60ddfddd4bb04b1903abb47cec1a52f
za6cf95fbc7991d5cc6effa054340278769d0fb3fcf0879834781538a50a5467155b4d1182bb776
zcb3d6169034b27ca25d7efdca1a90694a640da843a673aa9697053399dcc746a1659feaedc6d9a
z4fc5c128e0ec695ce17710e743267a13c452d02da7c904c8ced8b36ede25a0df9275f8b86a33a4
z9a2b373c3a052d9f3c3e28da6ae064add664be22c008b3c42ff854fb3fde18b4bce44d8809f5b0
zb22e54eec45304c1d8eeb5953573a3c7bb582951318210bd602533695d9d402c408e875f386fe8
z9fca617d0556d2e5404146d2826b4c94190bdbc7c47964f3fea1b6d5c1fc483add3587d6d2b9e5
zd0349d74fd4fcd9cb8fdd9c5f4fce4d3aba1f93aa1f66611c7dfdfc679ee60a159d48e9e183894
z5bf4f18e4ff69ec162aa511630fd6f4c4d2d966347cf6324e51fb8771d1dca3dce00cfd63b1237
ze215a85ede3926788e95519dd37b1c8c0a0b4288ad9abac0de119e3c66be487b6911f599bcb1b1
ze8d8fafeff54157909d6f996e08c5af4e95f86ea03201f90b4bf82734e1854e0e65b531747fe1c
z7d014a1f3e7247146ede451bf049bb97d05564e3ed5c47a28e63950d97d54ef976865bd3da09b2
z4371b5f9ccec8139ed4f0b28ec12a5c679f34ce58f9b0827ae09a0241f10257bbba35f36b05515
z7ae7674797aab5f351167f0a21949398ae6e63601f5d145242136cba7a77620bbc3eaa130f2900
z04546fa73d5c9781202df97d31afbbdbf1956fae59e18c6fd6d64c26597772a457f1d74a791883
zcfce0e590450c86ee0946428c9958000d0aa90e642725a1ec32f28c822617c1edec7fd66112f92
zccfc8692a7d6c3670eb1318d328ab1545ceceae03b7c77d255d7b47f0d5f228fd0330ae6bed773
z5e4c9fffb31692ae25c097723abcc2e91a8c7a738186c94cec46046dee834a99616375c832df54
zd7f913d2c1ffe578f9f5ec6b984bb7848016e2013fbcfae07a8941c288756a11c82cf3bcfb1d2e
ze26ab7c4482522915a0fade3f8168b8167efd991b94bacdf10872649b350741c21d06e16633683
z249ca51373bd958f262817ad8611d6fe275fd53778e0b64b6bd232a66371adc4321da8c1b7285f
z65212ed234021668332ca23cb13a5d365a09b92e7006e563a893dab618cd1efc5277036ca7f337
z63ecf0184660cdfda963c24af9831ccafd1c02224dc49561d04bdea2a46c4060a6a4bf58e3462c
zeecbaee52dcbf5448083c741a7b28982fcc95e20225cfd5c0decaaf21e4abdcd5560ba96c88902
z621f06bbef43bc7991dc26a3229039e6f2e9355ace552c1f9e360dc050f9f8653fa75e33bac6b7
z56c359a84a4233feaba636fe87cfffe3fcb18bd2087b8aa52c0b0621f7dec4820ae62ea96bb3a2
z78e705b2654c9f8b95dd8b166e147e21a5cb2c2b065fabe5b7dab3117b559e4e4dadfd068ec140
z26b5a15b8cff847438de5f710e51f6d5446a06df16a0334cb17b82d339bf582603787b5c199a01
z08019f0f57e8d2e042b307d66e4718add41d1ff1ffb50f0657c99a140f2604e4cf162fe568bd09
z2a1e125bd356a57ce3d4796979eb82e8d822abc1f9884dfb9501ef7d80c50275f613cc304407a7
z82b95d6ccb08378fcba5ffbca6952db5b0964fd9f4298611473d711f912940f9a1ed855982de97
ze440d58a23684f94754db359bf43596776153d78a7c579a3674f6deca8dddc644676f72235a4fa
z0906cfbf58297e80409179b5647378fa3e23b3aa29e097e41d3c366d2c8729233f848007103c0e
zc451e34c489c085e8a71bdf07bd9b9d8cc799298d41e01c2dc78c4e5dd3bc860d8e4cc73b19fac
z2f2a448b07b4f80fb62b278aaf24b640e5e76e59050e1733a950db845734083e6d3a3971375e5d
z558838b5f9ca4ca2d681f9f87756cbe3e3ac5981316b19b0bba871e91373ff1a5bc04ab96c7d1b
ze8a6533090923aceb562a60222a03e17712c2686d35d4fef3e792a4cd112d72948a4ea1e97f3fb
z52afbd0e02906c97098c676cc59defaf9d91fca900e5973c9bae1bceedc8a7e306e3d3b218e400
z68880f50e02f54bb862531d6e7a89ab48eb7e24cfd5360c9652e6956fc6b67ce0652242ba17f1e
z71a2831423dc17300bc56ecebea0fbedb676afa7e06084afc6ed22fd952f00523b40c4542d4ae6
zc88028c383ed4c402d9c6903a88a29ba39c6b6bf7cd22a866ba400d07b6594c5adbaf8110a6d91
zb858ec6af723e754add07a4fa3017d324471f0bc631ab4cae9615b0668d2ea8cbf4e9c1d5b6fca
z0f754cb97e7b6f02c77a2fd21d871350e2c92e460dcf6b42a150997e79a3328720093dfcef861a
zeb9e1b4e5d6ce28b6d5768339f35d072c79f2ecb6c69480ba20e4c8ab506204228dbfe9745863d
zd09730ed30854c0be45e5c0912dee274c72e46d8333a30c3e5f7a8abda6e88d2dc911952114a09
z4bf269aad286d691240e2fd326681b05adeecc1e9f55b92b48878b920cb89b164a404614d8ecc8
zf1fb65ef847075e16e0e22c7c04626fc89ffc20827820500ca6cf2641338bb8dee7263ee319245
z34aefaad811eff939ae5be41632e0757025fb3b5e8cb27984108f437a33e632ca0f3d68e3ba839
z974278e3b892093a30be8532dd2f6ef3f953bcf4c39e70780863e7552ecff9da37e16ff08491b6
z1a7062cb05e65037eb947ab4443df9cd9581704bd4fb4e508c18b83dcc504e1c948ccd1e26fe14
zdf0360ae21075c7740d25ff8cafc79b79d0282383270982a2a968299c6d45bb586dd817b2dd401
zf4d10c7341129514eaef900d6ba3973fa9bab6ea2ba1d99e61da93a476e98768713044ea6945d1
ze3cb0f128c73fdf082d4a6eb40d4c7b838cae172416bbe2370b5d2b2ca6a96533335d955d28d79
z19c51ae030943521d99cfdabbe823e55f7be22923aeed9071aedf3c58ae45b1757dea2dda88474
z516141ebb94880129cfdc7a4b1cf0227cf2f00a24a552c43a0490a9e1c1d48cb4a6d39db0dec0f
z5ce7da0813845094c30c134eecf3a07cbd1f3337a8420f6af7e66bc1cbd860080efeeb1b8a1150
z1aeabccc6970028df22a64eef26e768c3f7d670faf53247952e25a470cd080dd59e532e07e13e5
z5f058569efd7a0bae42ca4872b52c714c0f7e3e429bd937b3c198222ed7d473a39d0ee952c80e9
zcd80e6f2a2038498a0e50b8abf564779981a6cd57c1784212e5d12e0c0495ed6ba943593343b9b
ze57c21ace22f48ca13db5716812f6cf02cc4f619b73d374432f8e7e5888b6bf42b89e2a7b12d74
z7378e2d616614350e22f3a5dd8d97167a4b48ef89838fe650b4eba4f5164a66dbb5d3f2f545a7d
zf2d9c2a306e444f5729210209164813b631a4392cf9232826db720c6495a35e7eadd695f29e46b
z226cb71929af186f3bb1de2b23748a3de22404883a35063b74b7f5586e56cd6e6c6a2bb99c47fd
z5cec106350d61005fbed2421ccb7235c9bc70af43c53b057c13ffad0f4e1d58fbaa261f3b63563
zb4851989c75143ac8f11c7458ba2f7708871646b75bcc4dd7b87bde97600b720f1ea4dc7a4bf05
z2f3ab6aad4106556ad9c3d51d1a590d5c2422b48f6489e8a0483719939fa50bf0545a3ef78f7c3
za4beb0fec8c73310962dca5b6928d2aa0a32251290286cd136275328467ba8069228b0da6167d0
z4144925a3c1e9f2f294550534e2533d832a044e375cc4fdd6a165769d75dba6d2b66a99c6c88ae
zcf9315a1335bf0f153f31f7b27d9ccfd012518e2c59dcf44b51f2908f088f943e034a2af57d147
z7ada41479c644844639fa4b75f9100ad88e88ca11a7bf5e93059b0a3c4cb13818042d7b2872d1d
z513e69a8cd2d01af4293bc307003d0036195985e81994ec718a2e95fedda58ab30947f8e428598
z2d0be16d2f664bebb716cd512c8fc3306995e3dc18e1fe59334f969c732c04ad6087b2b35a4522
zd99ce7ec39d06cedcb6727c5090b09321d58710082d0c7e4736eb16b4f5ef3d4a1cad51a6818ad
z726c56c915cdebe614aefff50ea3e3e9c804b0280346d370edd6bffc4d17262067f9d194546dfa
zddce9744dff29cdacb987c5d5448804d80b276310115511dfda76078be87afce9af8575cc4c2fe
z5e91f360b106c9c6257661e65bd63ec7984dfc2b510e7b26242c70f72fa2b9f2491ebbee5f68f2
z0a1c9cc05d9a10829c22961abe4f4b7446553ded55a652a6181f373f2f976ccf8f0815a761d3fc
z9a23f749eaa6c863be787d0d158c7e5e8c65ca571f91bb2255fcf8f627f2c1eef5406ad9b39f32
z75687061972ea1bae6ee53575f8bf610ddae278f731de98141dc9a12fc66da1ccb2638d7aec6d9
z30efa9cc29799330ec1a745a2672497efe95a0673b2f0b30f8afa7e072d7b99b9e020fc2d66f24
zf64d835326da1f21bc1c20ea981c70a096f2671944ed44233b2561d5edd0d8adc8b7891e6b11b5
z2c1266befa177bdf603cee42b76ddd4d04d569d9524180665dd6dfce44e8035ef8e25338273616
zdd28899d6b90614b210181e18820b1569fc293629ff06af49b6d50cbfb80737943a50a3d4ac575
z7980094a262aecca91189f0bc85a96372d5c2c699311e213261fd4fe4225dcaa7cd4ef353cd1f9
zfc0bdbe68df59a43d0eee1cddd86abe1da065985b4ec515cc4b66cfe7c773eb2771f2bcd81fcf4
zbb102c2066059c6fa6d61537933128d9b5849a93866588d32fe4dbe631e947ed8f13d802d7ab1d
z418366e8bff8637509f9fb0dd0fccddef574a03266360d699192509e262a272593cc172dc39d35
z3743671627efb7dc21c225639d24cb452e2bd3b5d596933aeb53db4d67e204461f49243b3e71cd
zf36a1ff999dd1d00f089c9692fac0a7d0c1f23224a4dddbb03322a75bdb0760b9642ba28a7b46f
z441128522c144bbab48ec3e126c9e47ddccb9b21d1a397b94eb8b2a0b8f4447c756e5d5d231b21
z838e3563edc083e97f90673b17e392a6e8c4af599fbd9e26d4cd1a9a9ec00ad9521bbfb6b3d939
z0379afab32b71df4d92215361c880f51f62f5591023636d7c3e8b6d7ab46214f37f3e4cb374eac
zf8413008e6517a8fdc3dd0dbba841d02a1abe533369aed1408f65f3bb28fed547eb8cef02b5be2
z0200fac224485a9927a1d85af73968e3253a08dae25a4134c6808a7f292b788f6f327a11c94dae
zf3c0f295d142576cd60c0dc942528a95608b7c87537118ba1d132a1a365ad8726cada440c8bdb7
z6e6830c874950d42a6081d66491f6c9337752de9ad0ecb9d284b38fe2fd750eead1f0c0d46d9f3
z4278916337f8e78e39bdc08427f3ff4a053e6af3b1fc04867c624556ebe738286b1de83c612a90
z276b83cd726e41b264fc30ef96aa236cf1ccd66b12429b3fcca8c57785b341e530a62b6351c4d7
zf4b8378f5a32097f1b26d1d730df7ff8a1e7cd383ac84d0baa185faff8475be33340443872ae79
z55bb7d157bfc77cb30f6ed8847eec0b71915189dc07cd95f6610edf0b5592d9b70885972e0cde4
z6f589c5a51ca51f88ad36e109974f58d0409593b70921f0c625b3e4f193b371a74c68e1154c6b3
z338d4f8d08138479a0ceae02467d58bd62d2a290de071142cd5959b37d5011138c0363a5ed4243
z050f5644f46f07874d154950f2d5fc5ce987668fa37388451d4b3256e52ea6bb553fc9487fbd85
z3896319f8453aa20d5f6bc50fbb1667c320db778c8ead5df08a745e5a1b32003d4810ab52c4713
z9c5b043e7a153d87e5edc54504990d326ffd4da1be0caa4042a85fd34063f7f61ba1b83c401e40
z75757b85d47e1fc2f439884c1357b9fd39c7cc2ff532b9a3fc50c375c0bfd8bdff562271c0d251
z8465190dc77ce3fd9273911c849339599615dbdbcb6119ea36f4768d3b1186a2093d4485f33e5a
z170a800ff5aee5960ed6d624b4c2200763a1ca876d18ec2942224c1e093a23b3f25dc2ee676f34
za404a68209c4cf0da2cdc9c7ef541a725468ac3a7e5aeb81fc5894e758d223f2debb43dfa1b009
z35b177654637a3928f5a2f62a9f7f3f9757e68620efbef6231e11ffbe9ca4a998befc1e2d0dc7f
z8c6261d558410665dac4db7cd4b7eaf45c5baa2ebd820314d1a0354219c7f758a74b06e46e9298
z9b3d07f3b98430cc956cd6c04c83f7c98c0c9d7bb5ee7c62eaf0f2975b640afb0780b39e0a1be7
z2a400f5cdd723393b58902f69aaea54792add595db6bad79ad5f036d10e2e65fdcef6dd3c1aa35
z9100d1f51c4c79feef5c4b0dca202aca2aab0d9ace72c5f6bdee90cefc30d7b93ba1cae58a7aae
zb6f62f0bd31d90ebcd360b19cbfdf550e83e2b6cc146c649dda1353818a71d18a2671d0ac1024e
zb3765182ff5d8b861af6ecba026a2ce875a512716dd8de72554d9ffb42171dc2d41a5d9c04383d
z4dc3e380437f49b6451dc1ebaa082bc2f4cc7d889d79b55ab1b5f1f513477b3f63e8c7701fa83d
z7a1665f26a7503baf85baac52db2321d4b5108b2e0f6a4f985580537220e733572aaf36eccecbe
z7dc9d90bd09f94e83e2219f38bc9adb7ac6202f5be30bbebf17465234599924a1abc7f59026cf7
zdf243442e559cbcd470f80b31a19606df14c9d3619bc05a2ade2fba6882d503994dab5523b005f
z3f897a49c9661cf7449520c9ba28cd59dfbc877419fff28ab97e576cd0c65c2d7760227db61f6c
zcf61c7c8831f8dd246bff00af133cf752cd2a4ee1277fc0336db8d7afb09b2de5544bcb3c27688
ze09f161069a33f04244ae98a12697b0db4852e6892103db844479345ae925cb5d387d9fa23af26
z9e97a9996d50459ff703510c868eef1159d2f3959956d4ca74bd7d24449e3d9f057f499acbe96d
z76eab0aa0ccd4c08328127dd8862afe715b42daf547c5d1f6f96776c80e33e3ce1e0405bebd1ac
za999b8d11807f2e770e7c9d13ba438e6edd1ee8d987e285b1606d3681824cecae72d18a5702560
z9ecc0a6041ac1240f5bd6a7ac8d0602031c944ab996fa6c810f0d798ba4f8aeecfc5a037fe5905
ze5c0f660173c2e0d10521f93a2ae0edb86e78bccf7e79159e93affee168dfb510115f5c655f4ae
z1acf5e9aa2d43ccf3c2b056a5250e971c857ec3b30330e56caae5e132b5c952b3a8e42e159931b
zaf44221eabfc07444331f50ff6e56605180ca4720e12e66991e7d323f13292d945cf532295ebb0
z235c995529be832e3579bae94e34243b662351a1ad3e527dcc28142fbdf4236b37601304fbe7e8
z889a49f8a5359655ec3fb2a2dcce5f5b4ce9a9b488bbbdc53d3af30675d78f023ac0b9253d5d4f
zd7b64e31c1233776477b40fc7397f0100aab7b1f82ec96bbf61ee7581298603cdb5415e9ad2e75
z9704d413145bc819da6899f65d96994e4ef352cd0353466f539153548e0e3b5052cf8e28ec96f0
z20e4bd816075d26026a8570c3bbdcc473b98f0bb5018057381064c57276e0ccadcf2e3aa31641c
z8ca96487fb0396f1a4101ba3e2cbd214555babf3cdf1951fe1c2b9f23a432d606b6f80a0b848ab
z99b10b7da9e2394b0ba23c9f5a23c0eddf27e8473370b1c74eab8a25f70a36e6f575287a5fdc9c
z4a36b314d5f89986fe21d7bcb8af0989f5ba7dd55174fd9af2a2e59804fe14e0ea1e9b66721206
z589080d862c7c8ead982ea8613b38415ca3fa7eb075a32f55cc32592de8292578512949db75190
zb5a0af5be88361455ce78216e9365f2b5a77e47faec0d3d402a757be93ff5a6eebfc92a86ca0f9
zcd0eb84bced63b3f8a0ff967c4fe0b4b1a0db3b98384f2a3602a5817f544e002738a74a490a2fb
zaaf68154cd165ff771f3d161dbf3f17146dc94bdc7e61d6d49f61ddc74e624365c1ddd7f5cdcfd
z71d1b4709032f489295bc6b69f44d5d5c14b5b294b0a4fb9c57bf4a8cb8403c771f0882d919ad0
za093b768d81da6dfd2afa2d2bd3a72aabf064b8cb1ab11101e6f9a31aff31af7df5a79ab4a688e
z6d3f0073bd626ef4323efa564fe4d2768a93d4c081ce0aedbfaff96cfef33d524e9d3f4237f6e6
za9bb9383ef12df9b62013df8637192a22dfc3953c8070aba6bd70ec26e026380c36dc79a1733b0
z75929771451797b25f301f2d390121efab930c137a024f262c829234b0b05aa3b1d2c848e6dae8
z952432b575e844a3bcc31577739940436970472c8a5fc5ebc0592548e21dcdd3dedea13111aad2
z26cc401f1c16cc51e5cb20a15aadb3d99fa3406259822180c3780885025dd712caab8fd2984dd3
z1d4a632604fe564f0d478778052d07e43a4678b619c09066e17b7f209688c08b8c225be4b7e617
z20ee0e2435db9b7e82c31204caa975c9efc6046af6b630d82acb1787dc2a71c49e36af5ecd338d
z4c5f041b6dc3df5d5d29f79c0201efbd6e7a2073ec4c5b378acdf385cfc6ba0e124a5b5d10a089
z17247cc9d3281b3cf7c6d018a568c8f357b80c27402962792cf3ed571f4c72fb177d39594f5f6b
z5c3a9cf291f8f9fe67e65b8cb944492f20371767d5f292c1f68e12ed87fa7fd075cb755e4e58cf
z2585d71d4bfea4d6342f7f1f31816c53043e365adc008f001ed74fa21e062ea8582bdf97bc9689
z1a2b2d4a01de1e231bca96794e3e31d8ee2f2202f89577d05ba6b22aed42f461e4ce2d79570e41
z53d140e45a310be9ed9b0e3122f71615bb09623b143073470690864930d0884ed002515541a3d8
zbd3bab1b33c55e9808f8e07bb52a265cfc2ddc609296e882f57bb13615eced96d7503dee1a8c2a
z054b5b9c812652b68584f356bebdfffe47234cc88b86cd6b21fb313ae6634b6d64b981943d44bf
z768cbfbb80af9f125128842408ee51fe844af8963ee9c4da28f48af13ab9c7919f7d6a9b26d59a
z39b7088f9a93c17fa0f78970548e0f471d900bbc715577ec96e594179de5784d24cd3bd0165ad2
z268bcc6e251264df9afc0f3eae343da34889b5f0bef0d1f211b286d2ee128124875a48066a17e8
zc165c0d6f76a02d1c0cbac96d72ac43b1f5331277009e7e9ff97c58d97b016786747dd8335faea
z112ce80f839213bc4e1878698799e7ae79500baa676f2d5c85326295cfb5a24b8771b024508b58
z3ef99a17c2d9f9623610044bff51f43d77a1f3e53f37e1e27107869ce6993c435774e7326c79da
z54cb8091bd3f3dff70e4302be23a2bd0fae805335fd230fe4973dc1b016e08b78479c5c25cad68
z345df745eeb7f3e02b65e51810814cbd4f7392da9b5d7ceaf2a003e462b7115c426db4157073d4
ze6e8ff417ae04df8f6d01c2555115d1fd45eb1cd08be4e9f2797848131d86450329558dc7fd43a
z69bf02033ac47909f3c048df68b158406cfa724bb4acac08c4bba66460db6dc951e288d8637879
z826d495a8da21ba33422d46e0d6c37fc6a0492128dc61b1bf412f4e38eb61d492644b01686de66
z54dd145c5f7b76756a64a5953d9bf6307328a2c34f7cd24fff9db2cfd97ee88faa5de2ec3ee9f5
z0940da75e983e3dfbceff55da89027035ea2078e362c6dc773769dc80808c1751978d67e930ef9
z66521eb2500598e9d5c9f76d2c24d1e5a5b80fe378bdf90f7013f1893591ba5c0d46e74350c75a
zb8014f513cf6262d3e1cfbf6d40a73e2913f196755280bc7a89a7222e85bbfb33501365354b51c
z599f0d369017bff6bb41422d8f9c532874f6a3360da175b954893d03e6d501355ce722c2a5ee9f
z341bab3bc90fc5810921f5a66837fb15c1147f386895b294fcd6d44bbd40153c004bffc1a68684
zfd5e211b48f5bef1789697bae07ed5a7e43e5af3a47dea4b8629373238d9e82882ab685623162e
ze7faeaafbbf5a9077c6502b1e69f2f79d0b413d7bc7f582c39edd838e51db39e0cfaa34e1c51e6
z37b92a8ee2bcff2b14520d575e8ca62086ec23affc74d1ea65c16b111814549698f891b1248e8c
z561c520139062b607ca959de55c3350f5a83a8b40018f9f83c089884ebc911285b9bb60b0cdd96
z3a281938a48d05c75935a4509dc51a42863b55802e36a170c4986f928354e932c93d8d47f5566e
za4579425003b75eda0f57171da3530cc53a66fd38ef157c51a127aeed23f37a682abfa882cb434
zccd26d79b3f2974b6e2e8fea19d983115db217c96ada50358d197467c59ea08fbb2dc3d44aa11e
zb68154b6f9df256fe04984f782076d12e3079d38ef14ab086b126269d88143d728c61a7f0f5303
z42bc17f49b314c6ce93b30068393231abee3d694483a59f99fafc449a2476df4ccca0e52ca25ee
z4dc16984499d040dfb9fbadb536de58491d6f3807612bcbe33a211c324003d4a695629acd060bf
z018178c2b1567344ca8bd904939a081820bf1e33c15db650249007252fb8d75e39b0c54a47d1e5
ze41b2f4c828df7adceb9157f4e1df7ac160b28cffb5a307f78c521e25e69926f5fb2af479b0b8c
za8a71aaf93422cfd2294743dc0745135f7be6de068979afc238c3ad8597565a6dd004dca5d6bf1
z48ca027cd1728e501d18502b4da07938259de90074a6ec1f478b50de98af8af41ae8c7a97b60bc
zb73e51ae8160a5e9e6b1120971869512b20fba6206f44582851fab86eb7f7463492949349b0745
z412f788d02880a59a7dbedc08661e16dc261c462aaa419f2a16c2248afa90b8432c362ffc6ed16
zdb4d697e22a59aa01f0c416b6646189815ec3f88f32bb012953a8c07755099bca15d7a1bffc40a
z2aceb3ee6bb773c811c0126998bc5a9c0b21a7e6f37d251543afdeb02b856bc740cc79567a3c0b
z624df71244738e9b9ace421ac7cc4d997171eb307968b6f681d4dc8d0fadccc4ce4bf5bb52dc7b
z4b8e4bf1201ce90509d84b07ba7c4c558cb11d7ed8fa47e404a7e1c037a555634892836dd131bc
zc542de565fb1dabb479bd1e9eb8e97280533b1501486152cea7ce59ee85efd57dd4b62f72e0338
ze999c6f0fd148e49d96edb22eb2549a9185a91dc72c19d137e2b085fba914e8d02a823a5716128
z62a0914d79ca4a36100ebb0f17fb5fcc398754b2df04a2591c925451e691f867abf5d9cb2735ba
z1292bae52f37534980f69b4cef17bd86ad8658f7dc31578acf057bf79d26f5359b9499f44e49e1
z9e65998d45265faac02442350f62954aacf0f281aef460756a0717843da99b047f9d7bfe46a93a
zcd915d447b562f82f63416cd4f20b82ec2de5ea674073b194761765c192d1decb40d6c3c0d1aa2
z9dc3596d12aab45c664a4d7fc85eceab569858363d12a24bedafaec40d0339faf69d5dfe34f6ad
zb985c742759f4e87d5f2925b383bf5c251effc47809c5322521c5e9e5362af090765663f8a0e4f
z031d68c454bc5c88659d4aa2bd36b26293f017e42af703d05d6f2709c89be609916e2be5fb81ec
z03dd307004029d4f08f08c467c34b551d84d8f43a97459b773fd77507ea49b8e9aa13c2d088c05
z67b2df34d0bb9d01839ab90f69e6546be06e96bef1759dbe0c140960f62d44dcf84b2a85ec78ce
zea8ee982df800fb037ed11cea2fd8847100418989e808fd443befe76a2f9a59d1559310fa2de6c
z0dcdf9d3bf7632cc59068b500c01116db9a78ef3bbc9f50e200f09ae2d127e4d28b50b97347573
z64ff6f9ee26d3c8c54a15174c2c76906d4051897df337974d9a955fd3cd95ff485ca31647704b7
z189d37bd92feba59574ae284821a465fc33335f5cd4944a0d3d981658b65b23466ce4f9dea795b
zf806f8e8d55211e1b224ce30c047e7fd9ffb46da64fff8d6dce36a06f2a9ffcefa94d1c270ba9c
z3651fd9c3ddecce539c5ed25128af31f08d73df17c32ac89739adcafca1fb5821e780fdd173f5d
zd9058353e31a0485c23e7728bd2d088ce9ce3099354d0090a82b3ba3840ecc643b8102e34c7e9a
z0331d27a49c754396da4af482d532c62b3bce397f2ba1974e63a6ef96949539ba93bd5a8d18174
z42bfb58ba8f9d7b462e9aec0aef791ffe5fb57cb8b43ad6d1ab3980b5e91fe170de029d8ee8e7f
z1b7e30641829244180eea063410a2c57574008a2265e47c69affa2e2227f5875ab1bc151dc0b8e
z3671502b820271d18ff17638e2155b7dc147ba6f890a376991c10812ae160cc4ea2bbf5c645d5f
z0d9a8494bc34497697ddeea0a314e2683614a4049b63da86c6dce627b8fe8eefa00908d8058711
z8282de501b26b15ca08263ea6b879cda64e978bb2337eba6408fd8274c88bbd34bb43cb7580d85
z18a8a4a55b4de1a29fb0d7e6be19b9bae9e36727c4b5fb63ba92fe3c1dbadbbdc3070d91dfc1b7
z2312fef0d6ecb04c875554f7aa03d7a20ce1a43a410bdb7658b0889478e77efa5f804042b74994
zc8095abd084663fb97aff40f925b5fb535356a7d01b943943262717783a093735a8961673d7fe0
z9bc844887a3613d44c79b97926b49a7eadd3eb9ef2cfc2604fda4f9b14a46e202b079b96adc851
z2700fd4e8730bfde878a1250cc9b5a353282248310256ef7bf521697cc2b27b135da5c8d6ab562
z249f1bcc204bf7fb4d216893796e5287d61bdaaea5f791e33c475d146d14f612970eae89c8ee9b
z8770973ba3dd1958306282863f6e9bc31b702b804e832dd258b9fca824d66d26ac0cb2cb447e0b
zb43bb0a943d9e6f28e57a74f4b9778715a08631d34a0cbea2c51849a12c4a2f1a4027dc638a911
z40dbf254dff7967bd8e2fcb554168b99e28e432edcdda6bd988e20031b44c43c86aaa710956160
z6df9d750a75185dcd0b8ce5ad9ea5ea991d08e2cbd45c6b9dd633ab60b82665a385a864260902f
z981e003dfba8b89e7149ce06ddbc00475e512d8bb873c2fdd10f0c048466287747f0b6b7c45374
zf3d4bff46d94c674be8830fbde2dc1ff9acd66c13174f5a17500a3b5f529789c93e3d16c1c3522
z28945ef0aacb3ef26f3b687b68211ff5e855bcd5efa6ea5d0a72a64e937afd1e2217dd554c8f34
zeb5c17fa1946f9eddc7a41dc57827fd3b6ffcc8023ad4c09d7c438ba28ea508d588f13af4f3d87
zdd60778f57c057c38089dd0043e0c61a84ad13e40ebe4b47ae401e5d82d2c6aea8bd9b7e657d21
z8d1c6474f6dc35b0fa53424530c66495e9e55cba12876d88762407c16fd4c6fcf01bd5cd8110e8
zd697b9b4e116af1bc2d76f550e59e048ece7c97b97c468fcaad9b1cfd6435d133db96cb7ab89e2
z635c4170faa6be5748e827bacd1961b13b3132372c775c22c92e578ef67e252098c4a6e1b81e5d
ze93cc0938e7fce371ae97027d7d78a39bdc68fd6c6c2e266da3f400de0f176856e3568e2630a73
z9b1df5a23beeea613b58b4c9f0f00f7bb2faa0ae14c5ae5765560127f1915ca44b8150dd033504
zd0479b26f013a7b6212f1494580c13ef7135a2439a8c054c62131b5764a0064e8fcc91c1b4d276
zb63a48be362ecbc8ebac41d49f95460e1f52921695533599a259c523e4a55b588cca05a8f4fca8
zd5f9ff8576054020bd9f0a6fd211f47a6e6fe6b226ee78e3e42a2e2a63013a0c0215ada3eeffb7
z9f4426b0fa8f3136da22dee194dd9e363bb3e0e67306f846d29ab5b4a25ac63c397922287de564
z0c25680d7a1f934860b73a68b6524f938d97f504ec720b2b1f2ead2b6d9dd56a4b606f0e311f81
z2804385e4dc408820d7ab86e67bdcf820e11d948fa66798b1dcc62c02255c8e281afecda3d0ad6
zf7f9af1ff7ff41124a5ace0f948ecceedefc11001b5afaaaace594430647bae0e6fd1d5847ddb0
z7485d87ed31729ff0a181bb0486b7701b7a3976396dc4205eb43c38cebd3b6729dc426e52613f9
zb374e23e4b80602184e1e381122dc05f48c7c41e68914d0b98f1eba4bfc3cc61173507a2a384c7
z6ce8692c9b80fdf755dcde983a7d7a439b3d456ec822c9bf2a15f1ac29040f5bf9ed03f5688a97
zeb7d6411f800198c46c58b0081c216e3f2195f79c0a8dadccaec1a7a2f7ed4ffc7ba201f42090f
z35f525145ba5eaee8fd5317e2265ed2fe39dc1d4b7ed2b64d3b2d3119af0dd48532a12be8d434d
z23dd50eb9d847c8f579a0c668793a536cf5654bd7dee8325ecfd9b85af3b32ba4baff9f6944294
zfb5184651e1714a982dc6306b733012dcb36c3534692168e91c2290e978a1c4b7b9b8d336cc0b7
z2552a34c5b9343984c8db0a52c16a90129f8af5937c75086996eafe175da9fe69d059cecd9eb45
zcb810bcba101f94563600c89dfff49342001f67a8542da724213154b15d4cdff04a3494cea3774
z207d36a2912ffcc70a6eb87dec6c1527a2ea32ebea50fee51dbde3eb7af344a0d73d25d8478d11
z0515742607889aaad34d02be7085ec423b9af41d9ad2e20dafebf9c64db5408e288007b2df37b7
z1c3cbc88dca332dec4e8810bb05789719cdcea6b87b8439b05b8d4e660fbcc668123f80f251122
zc5ac41aa0da44792062013e4a3eb3466824b4c845f4f6c39347a5d1a44d488604eda5393e7dbed
zad2d61568c30be569a3d314a43e0f29a6518174276af7f94f3cc9a64200ae0f2203a8423dc2000
zb6fb679d9af65eadc7449c36c73e4cf31d08aa438236c4c9158a5c7492f9333bc46166cef1f406
z8db33c55e379e8c1d223358f042eaef4de95d8e49cb159f2b124136e127042bad9a6b3eb130acb
za57f8ebc81fc94ae7f0be31d8602bd1360428f0d7b10fa39b66a66ed4b27f7734505095a133b1b
ze4ca078a919339380d2fbc8bb3893162fb99782dc4f4268c7b237c056ed21108c0721c8b0f6a30
ze6368ccb89ab06f4d71a63e8c21c72f5a21a648983e74213d7266226130915ef83e6837cc08e5e
z4ffbb5f0f63caf82636b195cfc0faaf1d47a23c1ff287cc54d63473adde6d177809ce142153056
zb9b6df0c03d0c2d28dc67cb11247b4a01155aaf832d86231389fc3c863b42cda2923c0d79decf0
ze6835c279b430845597f261abede4545197266944e609fb45ad37cbe5c317e07160b32a1202593
zae372636cacf9b3217db997411353768e6ffdd6213ec530e8f44f381f6c98a8ffac4a17213683b
z249c234bd8e4fc545044a73ffab50c83c28888b7f2ecced70b77c920c434b40d654f0cef1b4ca8
z662a9797a3360481ecdeae847b638c8d98e783667f680b95cb0d01d3fddc97781effa8364a0f68
z678156fc974fd471720618fff3b4b6df7f7a0c904e4639cca73bc9c566f455edb060961324cfd3
zad4a899e221a14c3f0762d604f8216d21885e9419632ba593574aca1a678728daea44c42afce6a
z5ce7e91a5db85da9733f60b917f849a68f5849e40bb628aefcb25049b5c9937945023412745194
z70ec8f6612035e44f41102922c8ab7ce1562b4efe11575a78d2ebc5a6057d0ee8f7e2c6c52e06a
zaf5f52a8cdcc306eb64fb388f840052593fa03a40cf04060a835d0290c3687a4c349f4074878aa
z9a7f33f32811fcc3af243dbfb800593e48ca50a096c99cf5f59ab22486b3c77c4c0257352b20a6
z2175f9224c9eb28313708e0c45aaf699da62cf8f3c885f5edc87a17e00e5f3180236c6b9be3ed0
z36c0899b8f926bd25dad96050756ecb9ecc45c3043914c52e35e74e360bbe63fe9738afc61aa91
zbc6b3a32704077cba4bd07f5e47d88502e81fbb6aeb2d7e56509cfcad5ac46284e6f554c0c2a64
z0f37410309f79544d5a102d8ac8a494f61dcb04464db776a8f8a0a8188df222b0c09b555ed80d3
zf6e234643423712a89e7bbd3b7e61112cfc5ffac12cfc5027810b78c552ce4a023a34597450fb7
z723a3651fceeb4db486cce54b259fd76086d35e312e4c93aa35260bec1e33b5a935cd4a2cc2c59
z8bb090523ca25e68b7b7fd407dc724c359f60deb18946de344340baa43ee2b87b6fc1235f130ac
z7bea0b8edaa25578f56d57a3d1c39dfd7be0625c084e50d5894109d8bdc26946826b5bea0d98fb
z49c8d54861e3cffd6a1ad183ff27577942027b5fa6dc53790ac19f0f93a6b6af5559b907a87059
zbb673987a5d45a91a86c4bedbface28ee80865aa4701bd7d38c9e73e19527f31d891c58b81d94f
z7e5bbd3370616c8e86b417ede5fd8ec1bef9bd927f45691407c4a7c1d4776b4aa8d704ef9a1f85
zd91f4916ea3c9b835f80ba0c66c599a50c2c7f91fe9c7dc55c116e5e9767e0765c361e7b53b674
zc938be5e8133fe7313056902963d1e56d8222fb29cd5b6e11e7d9acbe7414add3ffda9610ca145
z8fd7a574cbe1448b9d44aebc9c25131683a0aaa3732fa37414e98496a0b95f8eb435726c98363c
z2090548b0f6e7c9fcb4334a1da0c5fd6f13ba7f26b263ce6a349274e1454672a2598dff530abee
zf4a1cdc182e9431898a684b3f2f93c6e32c659ddd9d5e3f2578f5fac850267581b9ddeaff936ef
ze55d378aa7b1ce4cfdbc7315f47e35f6ce01af783b617b678668d5a0cd102a3e6455631d5a7992
z9f690cff74f45147608701a281d9aaa13cd88f98a46697400f590af01cd7eea3e000e8969ac600
z7149491126e7525582fa7000569789aa67e5b136de11d023e6ddbf086af934b4bcafe2b894fdc8
z8e202604939d96b640f7bc638f82353d65bd21100adee408fdc9ecf2b2d16abe6c91263d5213a1
zb70588ec5634fee9c91ab0d8b053c20bdd6539c66baac2ccc5fa0b6fdad30d1a4ad6da734f8463
z21ad17adf8a824a8962aa9121f70308514987d90460b12949e5129ee5206a23bc2303456b0a723
z573bf3f7215d1dfafe544fc3c9112359a8470a1b5c81f36a8a7d5d6485467f4df1ca8c61801483
z5199d68c7cf6af8eca5298e65f97ec993d0e9304a59596f7f02cb769d351b43746794fe1c33e73
z193039635bf7257aa62e7f998179cfca4ef350d88a12de7d0cb142fdb8d2c61cee26ad44cc7324
za5145fc86820f588f81b3990450e80c92893e7108098726c0148479201cdd11352a9ee2eab08bd
z3fc5f02d22fa9c2a5d596a5d382d00ae7670c8cece226f416052296f38f485ad845c799b98d9ba
z72d2613c8f8d394f8d4ff2ca54e34bacdb9d20e6e00e3fb82ca2fa8caeb0dd9cc143b40afccc16
z8048039572eaf3b81991a060e0d95898666630671af455883dd6d5b895c7d362279fdbe60bc572
z31409c8f084aba20be5b8e8517468970da8071e0dfe0a0ddb3f918e19e32cb15c6d5cb5964fa9c
zd033227bd00027b61ddadceca38ba1687e702834ca1b93e6ebda52eeb6235a42df08bb0ee43424
zc2bcff00fe5716371cffe04e07a766686fcf697ad87f7e895f900fc230aef0bc6f3356cb231811
za548ad431a820e8072338fedd4eb39ac886ce4288a82e1206fa9a3cb5cd39ec58cba8493c72b49
z43d828e8795fb132ce10a22144dec0c2e9fe1dd9acd0f1d1790b3096249fb62b08f3726bc30c3e
z0dae58dea2680c22d2e06ec95153ef0abe997608d800fd0685e36f3ecde57a10c60bde073df79a
z518d37738ac9ad8bd34982c8396b3ec261207cccc750ddc3105cc38aac1f93807c9ff7195c2aa1
ze66864fc4e2079458db92e1a62ec9dca8164a38bd0bdf314e0fe9d9f0579acbcb78bec991e921f
z9dd0645c666f186de71ab914ba3ca4fd1f73f75df6d79de3c73c73a8091fd516733a1fec755e58
z7aeb6d41562aeb1ad557cefcb1d6981f86bdbf525f8256cdf74a7f5e81502896e0dd647f1ba520
z997534c252cbbe5c6c569a21a1959f667267d1a217d4f5868baf61a119d880c319da841c2b2502
z0a6d2c3ad50a20c0e17528cfa4bf3ce7bc36d6f799c7c5ad92c9ce79beb55a7befeae92a0f7fa3
zd8fb968700ace5dccece6a78beb6305da608697d49b189f53f99cf2910cc91f08e1d6b2b8d1e24
z7a99a25c13ba468649a0eb8519a213482f6b49af92cac1decd6b98ab0527bcf02ae04a6803e1d8
z4edf839e6e022a87e131c6af132a551571fdbb7beeb525ef0537bd4b0c98531f4fc4701f1db97e
zc199e398331f97c8a98d04fca45121777864ffd278b5f00918cb13f12b5e66d5dbc44d87f50f54
z170cc10faa710cf27d233dee48e4c9bc20bd56fd8dec2dd09abb913628438807e1f85d069060e4
za455749de47cf1234e6d341e5b3bb2d88593bb35af5cb4ca3b5ac528d7f181a61220188acae417
zf4d43353c989d294dc9d081a4cfa9953a82ceb0bbb14c622ddbf1fdb39cb9faf792f9620173511
z9af6f1ed783042b62fe1642299bc726867fa48fd85c5cce7e03e7706bf961b5b9515e287ab153f
za581afab8924997e7a666b697f1cb9eed72afcf5d405c2526d75076401f45daf07bf0890880875
ze252cc4fb1c46e2b86589ce306ebae7dcc50752eebc13efe35a8cecb4def675a13221c552267f1
zb6bd2dbef414f510baa5169d6ba2dfc9f64831fca9d6595a50d4b77db975e591563d8373c589d9
z262f6f9ffdb0537cb53bc491b901eba41b31c16a61ac99328e7219a78dea283b0b75f1a431b291
z4821a1c2c6824d31a45d606942050a482871b458ec352a28c9764c6f82b444d84a3d25c2cf7268
z3bac5c0655f23c960a6aaea50536f5a81f62944a02855f541fb5f6ce2e8192fac81eb0d194db85
z809e23a7b24bb8d181909290df8c07d23dc21ac4af4b6664809f0fbc63659443fa1f76fdb0548e
z24f1d60c46f4f7abb563d42cd9bcaf4b48cc7c431ce30bd59fdd86dee25d974e1a0de61b095cae
za7d194832b3edd6f9f98726cd42e86e0e595e1bb05153737a12d72e6b906d0f371d2f7a58b7c46
zab6a9565d0249442ae4599dcb7b86633d6d9b426ea99221536a3b89b87896e22f041bce2c5c130
z0258426d03572969bc8ef004e61698ff6f44a2ed289b902717b831f5976a682141ef2936b99c29
zdbdcf2a161a511a73053b13da1c6f17fb35cf987eef4fbd6b235cfbbded9d707edafb1a18cfb98
z62a2e1fb5336d3034b87bd89eb52d3ff5eff94d33d244ca1ee447b44de6477f8405e48f42b257a
zc6d7e3ef43fa7ffde3b9e8a3e4f3c85b1f0e7a53c40340ac2464574419a998bb9f6b39a707eaed
z708899876bc754bb195328807ef5cd4c76a8a7d651d5c5f43c7648971e9ad93f3d177a456f3e44
z870747966d5272cadb802eb0e544dc59ed9acc5b3b44abd2d20d808843227e3a0be8f194d76337
z85e7c210c84f2f7558ab188e36422da9f2ff76169a4d1629bec07975d31a6deadc29e2dcf6c2e4
z4306780662d06a615f588e26ea4c833f739faed422afadbff70ab43ebccbc27e8c8a1c3caf04df
zc1683ddf7b308cef561f01bd50f45214eecb3c2146cada5eee43fe0dddb85a5b6464b4ee367bdc
z8af1587ad9e02feca31851a4ff38b9fcd449915dc3efb67681f241b4a9d582ba6ea24f1c88c82a
z62b3d183a898a7aed829d838af3ea49a43350e19d7b48b44e50f80dddc5d9c24b6962f73d8e94a
z4ef640bfe9445d399afa8085363e67058543763b580f9c9d8de0a43e5e517ba14882e7ca8d2c6c
z60b577746c1b06e94fc5dee4a9ae58792d906ad4daa4d8142561c31dcb8000d8329f873edf5974
z688cb2b7c8729d0610a44ad21ab5332180043c796465b1b635ed2baa729f2c8cb691b5b6edede4
zca641b0d5c6ff175a3801d0c2abb14eded0ed4adf1ed21590e084ff9156caaf40b4684d18c0b78
z512d3bb20142ee217c10a5b6345919ef2d18f72a95138a9fcdc73b074298eabbcd8e70e5f29d90
z91359a192170859a6e7563b933b87a691cc2e5d68db24d799ae76f5b85693a2d3a7c59a47e19da
z72c562d494458fd4b034a86438867087ab54cfaec4a94f39112dbb2e10f4b9990a165358fc4335
zcbada96d3397d487006aeae9aa3b848357d47c67896aba28a2a7ebdfcabe09c7915a549a63bcfa
z82af3137c1fe4c2d731222676d2b595a935925e238628fbe127fef2a4244adce0f1e7599403c5f
zde6477ea70e121ff159e0089af6061d962009b82509a546d41553755c4697d80aba0dbb27f3950
zc2a2bc2a092f4febb64177e75a5c3cbe98d54538fe5d4e275a65bed8990466cc13ecc212223cce
zb7e8ee18beee1d4f1cbbffd02e8b55875038d6f7cf9d742d5ae30a1b4820bef46b0d718a66a658
zd1e70b229d628d5ec4e14924021283c8cf1ac98cb0a8a00d97f499bca0364bf2dc9b27e2f05748
z454715af38163670c7e1c27f253e814485859b3ee9ab7ac33bc1c9749cb08faacad7a95d59a265
zaa047c470416c76b41d606125c3a507aa9c9f3989983b9698c720d1652eaa82d2f6bb2366d2a91
zae17f8dbdf67ebaa5d023f90bb461bcb727dd199806d1f2ecf9268c711371f866de51e886e48ec
z9619365a5bfaf5e03162339adfd83a5dac49379ddb2f0e85e16ea29a1e2797a2cb75f6ffa3f85e
ze1c1e48807f10dd868830537b89043a534cceecf6bcf8b7155e7aa79497856228a263bbac3a6a5
z26217bd42230696ab9c5913f5d4591e6ff23a3cb1b2a02cfd4b120db60b26b82286293fc6599fc
zc99c2cf09ca0cf9cf9755aea54909301303d9ee443d5944d58dea67af8e26ff04ad6808e4b8cef
zac762aed0b39f44928d3c316cadaaf891e93709a2e84e6b9abccba0b95e88d051dc597690c50e2
za089b176e16fdda6cdf11e1d08bc48f2d3f2acf3a5bba78ff5f833e7833042f90aed3826dc053b
z5d2b409450997a1903d55bfc1d195dad54d3450f88b08d3138e60ee12c36f599784e2ef5e9d745
z12da5ff8b9017d7381c73743a99d24d5db60a5ca651fb6e6a591afe8f8ce893386110e08b824d9
z59df5e407e5f1a1f2f70b05ee63b6dacf751b20e300244c47a5d370b5bfb3eacc25b1bc0f5874f
z3b57db14519b30ef5b91e0b4ee034964da0df63d2fdcaea0c73cae7abeb0412c908e7ff0016831
z439ff7076fb4257afa28600e0922a5465e4356a28a140a7f83f1ee99a859bc2ef7d9f1d215041b
z2a06ea74d23e56ef05dfff4d8e99a959c2b203ac4975e9fd846c05251f42c6e9e33e1cf5627d29
z28a0dfde25c0da466a6fb7a33dd148253bdbdb267fb469d771641b96115712731c70913f27e9b9
z71c2cbb5096ec5b945934bd0491eaff5970430c6f42ed16e417ebf5e71d4e8c0ad7579469361db
z4b3738bd2da8d29253db751b24a1b723ab81252698444836826e8167c01d02524fb56bec279d6b
z018e8b611e7d6748eaa448177e9933e165011731d579de63c79556b2332e90062b9273bafc0e07
z38a938565dd799356d27c2b041b6d09da6821757a256046fabe6cfc69f980c3051578e2780f9ea
z986740adc9eaebeb0f75d40ddcdd09a58a4e57143635780d45b18107109264abc514a7f1786768
z2f437d86b517a1988df98e984b58aeb45525fa6bfc51d4083bc6fba76b956b475cd0b772a72f0b
z5969632c47aba9accf3c15188ca58891497e86d2e64452b8384ba3381f82ca2dd1cd5e623e02b5
z0837003e0d957848fee30ee3dc8e353865b3200ff105fe13bb0470cc0c1c3dd8f81aa1dedf8301
z37f47a6f0e8a8234ee1058e1a2469dedb1932b7079a3cf318a3973a0dd0443b6d10c8f411ae838
zd5740bdda8fe75c5edb86edf4c62feabae2d6ba1c1b23e0936fba2b64145d8c961e077e250b941
zc539ec90d72751fd6f6fdeda4b7a13e34e3bd2e7ce0818925fb57df9ddacfe1b29ba792c7f5734
ze861b7493cd910dc56f0f396e21208a2d623b9a9a4f657d4b107a76fdd490f172ad9526b269494
z71865570154e80a210c219eae4bcbcc56adc9e3cbb412d059b4295fe2602815b070bee5aed1e00
z5112285c359cf7aa16efa40ac990f433a3eafc15da0fe912162d78030ecdb9f510a1c3b6ab530c
z1b374bd648163940014ceae01936b9706cbed3b83892cdc133f3e0580744af0f272133227dc820
zd6342876d5050d25fc91f5a6c802da141383eb3ccc36687840428aeff766136ef4b8d675164f73
z6e3c3d571774747d74323f14a646fdd1956431d66b4d2189116d78b6fae3bec042279eac32fe80
z0ad617c1742d3bea450ef28d5b1013b678efa4b28add86b611cc6f2664d4c03766f7b9047afb3e
ze81ca18c7bf7dc6b1fe4f1754ee81571b775d2dd67259ec3c1f67ca01865286d0a8bac241c2ef7
z5983975133be1a7738d3913b72d81bc35c35489f7dc6059e1f7e4bddf7efcd05df2dbbd24a1a33
z58084b791397608119a60830bd265f43adb9b4a70427ff2e978fce15fbb5fc8bab9559071156aa
z7a6b8c5e52bf58908cb1925882be9485f720f78faea1347a4c5c6584b147b13d94aab5d054ca8f
ze1233139077ca5e08abea20aae7a01056fd792b0bbc99fd548737f7bdb9262fd980ab0bb6b0f47
z869d17a254fe931452c2b53fca7d2cd1b266092af4b880e5d28c0d17bdc9b3a21f36f44fe96b0a
zf1f8551ce645b859e554e354157c5fba38d420bf921fd716aaeb1afa015888744d0f63ec60622f
z8644fcd499565f4e9046fba554ae65d6e75738ebf89105361f24cdd9957a412ddd02a2c7ee8363
zc83d8d740660ab0e8965b989ff05f20745b22a261a50a675117c06785a262f3beda0abbb95e74c
z26f7b14cdebdf95eb2db45c26cd561870822aa454b2a12ba234d95f7ebe73ef6f39ba3c0fdcf75
ze665750e3df530eaf104a8f77fffb36b4d4a8c71187489d87846a2abd444ad7557d6119ea56a7b
z9138f5df1ea50891e4ae4b921c1656c5d4ebaa4de506ab7e61eb39969eaf9dfaf6b75421a4c071
z7a16daa6c8e542776395ee87e3532c73564513a27bfe130a02e3dd145357a61a20822915db8a01
z03747dba08185eeb5bce87d924b1739682e57e7ec96e8c0cb996468b951fb0e3dbf7a505e98ab0
zb8e46208d37ecff8ded4edba3519ba5a4e1f5587885f8979a24bfb08473b95fe5d37bdd593b7e8
z51a3c1538b5be912faac0b7f6a7faf24cd51bac130becee783d9a93d9e40ae0d16b8ec6e805e00
z38c37b2d8d92527fdcf8e142138ddd5837b3bf625b2e83172520b60f2aad82718ea58a8020e955
z0eddd62071afe4633e4852a58678894103b8b29ff0dc9d0a0b0c8cb2f854395b3c28020114e7a5
z5e3c27c6c91fc9794e8ff46372dd0e0c4af5285eef236c9c7aea38737e0fc9a4500d874324c9ce
z317f5923c73a044d370df98418814e56a03c28d3b9f0107fffc4a99d2c160fbd9a1e14cec3e92e
z793088afa500948f60f1439b3f90fbafb1c49659b40b8238acfaac1f4109bed2f57d427c7e4f6a
z97584cca74d45eb6bf477f3047959458fbefedf86237163c499719ef5805321075245001e61d36
z65f5a4594200bebd8717ef2010e547e4b19444e885e60bcc458ddb7126f9434a4f31d1b493f96e
z58735ce50cda76deee02d861ddc45411b7020d6517b66f08a4fc0ab6915e36a3efe226fb881490
z4731a0b7105fac5700fad97077556e9da174ef7c223c2817bc3549e0b1eb49bb15e6ec083ed10f
zc3e298fdb94a2cce6f4a30a35f61d9d821528d6849043a64816e6d20cb127368f221d2905a2cac
z176f1bc87414ff766054eb67986dca1b8df08815684d126b1227bce0a3beed2d94e225c4918d05
zda8bd91c2d5d04968fd3225d6d7044b65c2e0dba418df09e88242ddea7c3e5321edeb2ece56733
z37cd155cc28e5a1ba3162aebf2938825af684882f32038c7e637a2eb579fd92556107769792eb7
zb958a0f81afa1770c85b5b589bc867cb91379d47c33520f31793caeb6f12d7c9eca65476a3462b
z21f8e09ad6500376246c2117978b42bee42292029686dbf79cf794a04e2aae7d458ef4254a3360
za2364f8c5b847fa8feb2c1ac969ba2bf41e46d13a4f128f4b14c08d6c3e7fe56fc6a761cdcf1fc
z0d8044e360330d4ab0af65cc93e6be272566fe269ae30a92a67754db46e1bb2de56cb44af04625
z62d5c9a0b2cfbd4436e044584fd82db0ae833f714dfbc2f05bc975cc00d9816d93f0845150ef42
zee3844c70bb89664d8a2a0795be547d02567a3bdf5e680343756816ab51bef783dd422e0d61869
z902ede840e2bfdba5e08ef0c0dd97276882e9cc120c01307668db75f469a40ad20e222938a588d
z0f57c0180a7325ba98524501c5805dba80a476451d5abe26c82f634e677acf8ac5f305338086ab
zbfaa1b69f77a63ce0087daf4d865e62eb53768149619ef749f762db62518b0a4ab0548c4cdfc10
zeddf251888bc26f87940a359248081f7639a55e5e14500b4a0be76299cd2b88fbe20007992eee3
zd43352edbcccd4b731edc5aebfad6e05c6d33b39747e1d1c1ea897e483abac46e084c93057c951
z0947a64aee30736f50572b0d18b7ddd8514f213824849464ac80cc679974a04b537d55c559d1a7
z651591f21e8399c6366ee1b8c5c17c4a01cb30e212807268739edaddb05170595be3201314d186
za8840bfefbe5abd85caea50e42c14c9120e3ed7dfb91676be474fb8476e8b5a66480719dcece07
z2a65eccf5f559314cc41a2ae01f282873ed533ecef18eebe25d979ef70d47d653345ca4648c796
z439c1476833ab9880b0cb47bf99db278f50a7abf913a6c6ffd6682bec2216e83c8ea9211414803
zea0ed22b2f9f165ab65c38c89801701f1ebe24b7a220833c0a1def5d1193e21868ccae420a727e
z20ea7ffc29c95e0e5c6c4c35e3820e7836ba02c7c548766a7ad30c5a8e937897ac8984b2d4a05c
zf15b7ae38cad40a33e2540bd3de1f8a704aea46963363c67379de5a2d28041d45dcb9d9868946f
z6a802a4f37f4944223e4221e9afa7c1f6f980d4c5a34b7264b8e5d31aad520bd7eaa13678b5028
z95989d0281bb2251c5756606dbd4ec6c2267c5d73710c23a20c0a7f1ee901ca7d7c282126ecfd4
zca34bd2bc1715169d8b8bd37f96231ed8954a26f60ebc975bf50ff1a595f138df40cab5e057d8f
z741d0ccbc08358e03b4dffac81148f388d64374dd3f1aa0dd94a23efb65d742fadaea504cc2660
zc4eeee1869e6abca38dbf754cd0b284d902b0fabb8a06e77fff10ba0d60e0660755cb9b5ee11f9
z76f1b73a4c313dfdc0c61a875912c9f59bf9abe4b2f729f9332b806c1a96d37a143b464d85c3fb
z76f5f3869d40b61a076b94b460e15a26349618d603fb91b60fde72b9e5be623a86ef9f90f27d67
zcbf6c752e6f09990bb0e9d83d44ff3b1cb2abf79366b0a3e6eebe8d6ce0a2fbc7d438d1f122b90
z69d100da2fa790b11dbeb8db8b34db56b013ba5408edc8c9891b16f16fedc518531f141a933608
z7bed011f288336e7a65e1997ccc01ae718cf09d4470f741742b624916559a7112c1ebfa19b8935
z62870f0a8e1f500926c815bb16217cec51f65e7f0eda637cbf211d9127c68cd80438011afa0d9c
z6056af33efaa9ea1cad8bbd7ae4e1caa9cc8065746d86b416a15082df00e5cdf7da42fdf70dfc6
z6366958bd7e20a407658238a94b5b779bbeb1b8c3fe483aee59540f2e521f8d1609923efe47144
z4272275c1a48380d97c7da5922bd92fa9577faf65535412c63426dacb9972f278ee4545f41dde5
z309410acd473b48c82717dc031ec6f96181bdfc5ff876bcd2d3a98f50eb83b535f51499a3aab12
z24758c9183102b787ee39e7462fd9a7436d0057afb1bc887d64bed7fd2423ab66ea579523b07b4
z78698a8c1e6a131ae14f12bccfdf74c6cf4ecc4b55c6639b1d1fc198ea7ae6230c539685f278fa
zeba02515acf320e3dd953791136e425a3de92fdcebac6c4c45f9ce8bcc9d5f3b7a52874fa33296
z7d31eb4785c2588ddea33034d75e8a7106ea36672bbd82aab173c9bc8cd88abc50471739b705ff
zbaf668ed2bba0d2fb3faaf11e3d484eafdc843586fae5edf36f0eeb39ced58a59566e9abfd0901
z34295c5e4fc0f3d8cba1bc2df1a74795a06bfe475e9e3225148ed3ce28ac0c6707ec0ca31fafc2
z57597f62b56cc2c0a8fab92899d8759328bf4cbcb58ab97a4fbff411e09a22b252642d91387f9b
z3987f858b3dff5e233d3dbed076a903963405b4036a8d2d74814286a41b794265465f04507bad5
zb24a321c000e78102ddcb21c2496a60eb428a1cdeedac565e8c7aecce0e2cdcea7fe4891f0c4ec
ze29db63f1233c75e569ae52d3e6e5c012ca3347a34cbc741ddd0c1a79931f18381e47fc7bc2128
z4a1cfc144d7be7f81ac1212d1d1380a446c94cbf737315cdb16c0a57497a82bb2201559ae6b79c
z48a82e82289ed134174165f045c59ee4676b770594046211ea7eb37e58d877e97681085d5e31fe
z0dc60af4b6b4cdb439f5bd8e4f6f1f1f70a7b6fd5b843a88c446203da4670a4ffdfe0cea8a085a
z52c037fc2baa0ca6c3c57e5e8a3fbdc5f0f5a8023ac8f75b5b401756efbe5c8c117b3207570679
z3cf72ba5754e8562939d90be412647857d2c52eaadaea5f85925d18de9ee4053c186e518627a72
z0aeae1fbf58ca6aa495ea5b96bd0b052aa6f64f2a03493b53801181def5b7e1e750174f5c789a5
z63988ce6fc4229c3c969ae812f01a77113ff97471716e8c0bc049760c9f1477ad58d184881e7ec
zae9d7f845320e2e1eb54e0818ca0b801e5ce01c1c975d6b8fb51f887105b8d74180748b8052d75
z9117cbb4b0e2e610fa144ff56940edde2f8213083d90974f05ca6adcabedfcc0cc678ad7cc4823
z0d862a544d07d375cbe479e30b9f2be8262443fe29c5a4ba513958297a57b03b33193338c20120
zbcde9eea32295f43025ebb339b147a9446f529b02df32de735783a88bc921f9b5a9102af6bd47d
zc6899c24f65058eda02b775a562cc37353bd671c446a0e4e61fc7fb101292f9891514661f1c8e9
z5a4f1722b506ada9acd52736f20333d051f947f240cd66a44d80a17c8de8722d2537b9b53cd0c1
zdc29943f8cd29c3d50bf132509c306529952d20c873346ca6aab3c78a17dabdddc816d13a3cd8d
zc3e9184ce17edfda504bd8f5a1cc4393b557fd35fa07fe18905317b4664c484fc4ac10179b9822
z5988e97a99f2dae3b3b1cb06dd52f3f7cb33fdf5c0db000d049439e9efa645aed88c7f5eb74d18
z64176cb6a8bbb812bc0c4d3185fee69e1470e021bd2fd84bb89d56d7c49b6a1da6ff4c64691346
z3e3e44e0f8ad9623406aef69747ebac1509428536c19b948cdba7803e3633120010cd96d9c1124
z85836cdc8f28155e929725ec41d80a846c89b0ff944128bc8c207343aabd898d8b43ca9e3a77f2
z7c76ab94f9f870753066055676fdb1b469b3c97510d66bfcee3c018fec18836260b6991ac13589
z1e57516b4a86bf970795443f8ab6bf9f018b2ac93d80ba1e9a8b4b9d89df3f848f47e1e328bd1e
zdd26234e40a0cb74affddf74cec61104cfe626bb7d093b61a115ef0f8d3574ba8c7f9da619cdfd
z4bd5cb54149f44566e0a197de3d614413fae860147ab729bc6ae116fc51ad328925531589077f0
zffdb190288a6c241d2da1eb51c89ce07c8d1e0909c01775db8cd6c3d4de7dd8c5030df8a3c885f
z7bb576a87d583053f6c358ceea464a82e9d2b68dae03a23fb15994e36da430f3d9205d9bcf77c6
z51dd0b0c544c1493527593604fe971083697f13dbf6f8ebe7aef00bd4a33a3ab5805eb6e1c4eb3
zc53f55c9a2824c7ad1950e30f45aa7d50919a6e5e90c34491692c86276d51a33681822f9cb980c
z09ff684a60a88b6a5eca14e3bb08d3772c7818dfb2b20067f83194e42cadf662f541c0166e1643
ze65ab968e66e885f2464cc3861fd9e61e37833e181da54c3664f14912858908b354e1d3d6a422e
zc59600bc4e0ef9c3a38cb28b005eac9a0e28dafba952e7696e6330fe5cf452f402e7058fc25287
z5700250e86aa3dc339fdba41abdd7dc575f4e48872169ef1b4b6c3d121285eec1b2d379580fe81
ze60a1351ae35c6a37448de180a0fc343da6b33c11e66d3d3e8e9f7de2c542ad0b6e094ab30d614
z8395d4376dd3393dc90770a364e1d93a62ed41247305d0ae8a196ea0d8028bdb95612a28edcbb7
zd0b1ca99f5c896ca3d2791b15dadf6e5440df417455ace561c042839551c04839a39421e318e0f
z70fb21306cef5e116d55fd5156963b0e675d6905cc5186e58458e77b753acc15a7b8a11cee3cec
z47331ea62083a368bf3a28362eb3d6f60fa5751799d99ada87b8c0bcaf04b9e7a15412735405e1
zf3024d63e71e5b2c50c984cda94155413a206adc90c4201341cfebbcf9d9a71641b6bcf36ae3ec
z73a7561c9024050b9a851731d841ed2c6a13a6219fe0fe619459c67bc38b4bfafe67c47142a18e
za2848ab6929e4008b4a8d157895e616b454835027c2109cf6509e071c0c26c45ee8d70fa20cfa9
z88d006ece489e641eba5b48435ecae20ab5163d96e2a71cfe376890f2e4dca4e2f46a06b7f6e54
z9249e04986a61becb92f08133a3fe6d7282abd59541b8a5d7ebd90ce2d750247fe879e7d2e70f7
zbcd2266368aa2c6b09b8e22510ce97d62d5a560644a694f4fcc1d5bd740316e624be31dafad5cf
zf1b37fe702ca86c985f43d965a13ea237f97402f68804840882d587bad6667554741e3979ac27e
ze848481e0f42a8c709ae5ffb9e3a70be1539b1c3b20922f5c329181870024b1b9810c1c8474d03
z1b3b208a14d768f91791bb7b7ef00e205a86a7f17d6094456df17d2e67a1a13bf179ac65e61b51
z4a3492ece0fc8938c7618045060d26b6fa7f138ed5023f8ec228e9625cf384de0fba411521b40d
z4047c847ccce28642718cf4a4e88d7283cc6c057f3ced1186a3f3299f1b8b8b26a234e175137e4
za7ae4f1ccf7cf270f1f976b118f90ac335db53e6c7c414db09d92b0bbcb4e9b0d9f053a148d1ca
z60c52fa474c993d43888306597e261af5857ece45f9be440a1be3a0d442ce90a3bbc86ccd9809a
z6b72cdcae587a7d1dd1952045322d1375654a0ec69411c84e6532c7a79d1fa1efb17374b7ca5ee
z538501b68b62fe8a72d197e86fca397e3ea93c9b3039b18b68ac727d220e0e06e83e559045c844
zee3ce472dfbbc9ec495ef92b7bc74fd6a80d2cfa624d5a3475a5f65e222a8e5fbf600b97e77cd4
z31f87cd8b5bd506cdd6582417571ba2fdadb18bba695c72c480269b250cfc04909907204db72f8
z9926c7ebf862b46afeaecab9cb272ac65e77dda3ed548d8f51c58cfe0ed4d39f301f95a1afc7c0
z7bb01e8ddb4cb42faca95e85357f7267d3963c7f4159750511a20e4256b4b577d1afb4fd364813
z2e6afbce964aa00691f98944bed66eb4334f32c01b2d3617e20cd1ec28a626873aea716e7fda54
z15419a63bda843ed3b834177794cefacaad0068658f741c811ead4252afe165f3ddfaf1545a1cf
z1c079c7cc42b56ca777b7e16e84846d6e0545f9df81ca3fb3236578ebcd1090f5b0ffb51f06b83
zf29c3d017fb9debb235f7d5a79948faa62e8bd089918e70feb9f6df5ef77e734488048335195bb
zad8a059d6a874cd36e0ba1eb29080ecf88e0d4ceb93e7abd70726758678d01106a2e476a9e3dba
z3fdc35b6f529ef610029e13317d05f2404b99056ee38a4979121c53eaaf8b5945c60e6dcd3b06b
z1cc5eae6a8fdcfffdcea42ff4e4fe8fa2d776a0f46511b917bf228312d4f8b21e48bf5746a30df
z56d74d46bbbdfa9ccfe3fe1fb6a728e56ed78318290a529ba312e440ad2a0fb7bd523d68030912
zdb78187e72cd4c59f803a537115d728ad799f874b6e7f20cf13f99037bca2e6cc20d75d4a5f565
z2f3b3d6602aa90953ecccf73db4377080276f3e8c5990237c208ed11712ec556f94eaf368c7e0d
z7089fa308e37d1451da720dc6a00c1d7dd7fb8045341a70d564bbdc17cc6ada92b3c56d8daff3a
z65909d91e0282fe9dfdee730d88c710a320aee178cdff08b3a31da75705ae0dea7c3633915c42d
z257294a8ba9d8bf021d1b1be259044bfac6ac92e4d8791c5a378f401a53094843f70b72a463066
z197951322dd4c4420e464966643aa0e62ecbebdec7b42b8358e7fb6aef30140ed0c8c40702d9d3
zb3b8ce0332efad4af9c7f1d19d763942ea641125411cf0dec7f1eb84797eebc699b97010b225ac
z9bff4927eb80075e6469d106250367cf38f18b104f5ffdbe568e58b9ca777642ad78cd3d4fb4be
z27473b997c4847d03fb2b2f986a3f6edb5099f17775bba66d31b2d08f5eaeccf46bb64b940a70f
z17db6f16d8d08bbb2c31090b118bf5b7eec46b8d47784770cb13a60bb4f6a0b764ce78cb6f906e
z0b793ff6287fdb497901cf8f3c492e3f12d5e823f8053676b21ce73795574867db324e281d8687
z325aafcf7e500da076177ddf18c97b69a387e5f0f12d5ea1f9857947155a944d017546827a6660
zd8cb23878cd69f1ef6490ea7ed41d8266b7889f4849d6ae315bc6cdbb3c5d2b77eb01f70bb2900
z925859d5eeae756994a265dc632b5c03872a52209fb2e702b1dc7287187cc73d0ad4d2db7d8e5b
z5e2928bfea1a9b79603c082029fb69baaf53579ff6fb8f196dc991c5bc92607a7d347b367c86c9
z24094d6d7d149751e01d5e59b381576e829945f4f30330811afa0b82ccb56a2bdc8556b6043e14
z6f8f385ecb6e063116d6611df2999abf7a32654309524fb2493fb96613adcadd65e48295f4d039
z5ebb28fca6ccb282db62cd02fd47de41b45b4f13604ad785c5dff2121bf5f155abe45bdf4c957a
z6a4caee86121c5ea347e04b6c2e228befcd19f57e4598c7545d4e5446a97387a07733d4a7b377e
z019725e00ce450ceca37886eedba316545ae50c3559e3faaf6e6e2e7b9b3d955193395c23aabe2
z79309398d9c73b0a340df7684c36b15a29e61e4e97b917e6bd45abab6f10c8c2b54ccd2e9a919e
zbec41f41ff2835fe4a50a300e2b2560e4f8de4a56b23d32f903a265b629ce066031f92ce3ec8f2
z53bcfaf4657caabe88bb408692daa2009eff41c3918e324d272063a11d6d9017a8190a25e62107
ze3262098a4083df11d0a4812fd101264c54174e7026ff87f084ad217178a1ecff80d4cf06cf74d
zd801b63ca87227e2fd19b073129f82b933237175e162feddd53fdb2372a999d42d653298dd4377
z23cc2803713e26af57fe703673abf274bb539da597846dbc778d3cdf27e076c43da9786014a198
za8d6286af74d9e9c3b23c3823ad66d5228dce85716c55e1f8700d7045c04b19aa69dcfcc805d6f
z075d0f81d1519e0001ba86a21c25108d1556fdd4509bb83e4a8acaf22988741e802d8e1769c3e2
z40e212800161ba719082b70ef2283730fddbc7ca5732ed02430b8f85dbe9fd23911c3cd85eb7e1
zfc291af54237fa0f095c032c1b4c4f7774ae4e9523b2f3d50d2f996a49cb3404653b6b8178b2bb
ze79ff7f11d38b3c3e9b2c98de6eca1ce1e7fee8c55c87990b377a531586b1a1081f099c6badcf5
z59e080f4abb33270ffe84defe6970e3972b71016d82aa0482c2b73f9464d3a15ddccf8b910f31e
z97bbd61976c61af75fb78ff3b35cc5d29635721098701b779cf2367d820c48153e3e9d6690515a
zc9ea3d8bb788eaad490648ccbac3354c8fc6f974aeb9908f2b037dc0dfa27355b00c79b2a2ebda
zda4a53b1bc6633ab34416f5989e28e344b2dc7b2acee0513aed9683ba37e4afedee33171d429b1
z084c186c84c4f517a0016f81ae3dedc49c839464848ea51325374f251e245bc067a563f2ed374f
z0784876bc2255a6461c98eec232e209a60c9bb3569adbbb54cc8a0a4b3e30e8b61b67adb0b1765
zefcee7848218610bc90da244a3bc1000489434ad1fbb960c177b5f891c23592f0ed44c71a24065
zedc56f23996b448c7770ea71f186cda13c71b90b0bc0442a5aec3d2136fe1732d4a82f93642418
zf8d525213ed80709fc4903c4a736941fe2362e798918b8323cd75fcf1dc2dd5de22c473fe1a25c
z4b802d2638ce0b2e053d0ee9b044d2372c09e20a9ef9f76813b6ab68f79c703dcd7944a0d62b28
z1a130dce06c7f099ed0c1f4475c885145f89f035055a55b46ff00dcfa0b0d86196acf24cf23558
z4bf878cf5d15e22e5f1772a63ea2045a69f5f2235ad33554af9a37b9f91cff9e50c53b2dd73350
z21370f2f183c36c349afaec6f9705e1ab55b86afae3908c5dc679dfff7cddbd6f267c1e1248ad0
z630194a75abc0e7c93d384989d4f1526a9ada96863cff4e074ab2f7d8de1f87ad0430e0471694c
zcc33891be467ab69650e4730b937b5b8ed733cfa9a578437d5758edc3f9ccd35b672bd55c131b6
zcf263f38819305448e716dedd329573b6612b4848e458110d51109afa9c5ffbe523f45198b56f8
z76893155992bb6922ac98839278ede55994397234293837fa8d511fa05654a5463e9bcbe004221
zea1fcc04876b8dc0f4ed9c4a223bcb41831518c0dac1b0c2d02d1816646d1ff1fd5ef1382bca8e
zf4ed0365cac843732777376b6475cc62fccf3a7a02bde9764fc468448dc970634b185fcdcf0f5a
z98429c32766eb1a48b56e30f54cba3eb9b961ff6cebc3a125a48279f9061bc6e403440f2a38bd0
z2d0fd99fb41d16469a622cea010e0650e39ce1545d970fbcd08bf50b9cbdb011f0e77b6667382a
zb126d9b7685eb44ac6322a3e9748f61b36cfc60b513e16f6a246c4f8164563d68ed2fda2d7de66
z9808d431f5ddaa569b2f63be5ae363eacf9bd11fa9100c6a3aaf40be3b69994eda3846129998b6
zd12370ded54b44351a22e45f57bbe6ce8c9390ebf47c1ab62ad3224ea22037fcafbdee7c582d2d
z903924c38ad78724b9a466c42550b0e30357fbf214df526b97052dffbc7b385aeaa79a734a125d
z11d384bd5238a060115fcc01745b3519ccdfa6ee54d994129866e7266a5bdfe14e34906cc6bb08
z433f70539c12eaab64f24d77fcf6351d7476882ada3b09d9840facbda04c48822b0cf936261209
z02aef5546e68ae34bb24ef0bc31e9ed42a900dd47017b40e7417d18e9921a85f1a8ede9edcab41
zfc860c8d6844af39cc4eadf4f48fbdfacb8d988dcaa05d3cfe24128e8dfbdd02c0ebfd48ab0349
z140cf7fb05ca96129fc575c0c2741d6c18a4d1ad6cbd49841e1d3da2672072f7480b9bbbb27356
z1f44b4b7edce7a50db20e6f1a1e36eb4cd624f3d03d517664372f0f4e248fc0fd8bba7f1249e42
zf9027f019600fb9d8722d2d8f442bee1649aeac280b184006401ed9124ee21d86ffafd03807c4f
z8de23bc7404d28c028e5979bfc5d770b732534127faf7d411bc5ed1ccafe0f1516d21f86a93ed0
z7d90f0a92b627148d1b2d2f917a119e1b52cfa51d6b2669425a214acd2d32b291316f7aa26e946
z3ee0b220de4100600f3c892b84b1621d56be4078a527cef7ad745715aabc5a9b0b9f202605388a
zb919f469ecafd577a6cebf8c0a626419c38e6bdbdee680fc77dc623053d67e09f7c0576a0a6b2f
zc89090336d367c17f232b43189cb3637f91ea7f7efd8f1fb5afc626d92faec238472623afb7842
za37af1e0bfdbfa6df4d4592e3f31bc2f2d18e9a54bacda684b50c7bf3686c2df0d71fe6f1af845
z79fb590bd52a25167373d2b8809badb31c6916a8ab82894be0aad87cf6c0b8e5de803c01d847ab
zb82b1105c748b81d848656c526103a6c50f55dee31e28a150ce61787ffa57c8678f80259c0e2e5
zf93c87289da83c6ebd9082bdbb750b14c43ba2bce3ec5b4983822d4a953581aac7ace0a6f881ed
zb5be620063e9bd1985e6eafa9018c1fa896580154f7955f883f2cad207d53d5cd6d12fa29fd709
z5512d91610eff4b20d9dbdf3b65c990ab6a83a29b3272a2fecf5c70391d78eef67155f1d28179c
z6166bcfeea54546012f18c4e598a52c829ea263b1c966aa8966b9ae17728693b41cea0290246d9
za6e356fb1d1cef35dc145647244f75a70fa467e8fc9efca7f31e9d47a17dac0b729fb54d31bb85
z4fc0c26716ef5567f55065cda14faffc19acc8e4be29158583dace91855405babba526ae0b97e0
z7ced66c2c2445847cb84e96f528987e60e71f7766790ca477eed45b9cbd05f47d18ff887e9ef73
zd97d12c9ac226c155c0af13ea5ae74ba3690b4180236576d2bc54fa9a5eaea22d5e6746f3d3e05
zc1e69a21ff2b125f9aac81a6369b30a0e7693fa9d874659757133074b0b27f2a8000f9db7d247f
z5bbda078abd4b40d12f5c0a80acb1984b96cd981a1614e3f72f3fc22fd9fb1c79e11a349f9c501
z6a641f182454aff6c49dd422ba831ac2f59445a715f57e8ae88afda3badfd3265d6c145e16b490
ze3525b75d011f42d7e4784dfb4041bcc3ba7cb176599099666a39c6390ae7def9b8eaf74aa1530
z48c3acd25957774eb0147c924430641e9b363bd12b63371861dd650ac2dae4656d853902dec878
z5b5ca739b3c34c44f21e6bda361d94248ac4a435bbd4168e1740ca342632a867d0bca1cf126207
z7c7dcd7996fd29f00226656435322543f4b7ba45a3c92373403013c42bf1332590c937918b7f58
zbef91cfd4324200da8a3084b5a140b6f7154885ec9de1c07b9fd1b78a7e0ee16c3b4451d2ad3b3
z6b1652e0381e040a79904e1c00c3f30e155e7adc2b219280ef8672113c712a734230049c6cd8b7
z55df97655b263b304ddd89f4a945127062d8e75f0a684e599de1c92b70b15a481d505273dfbfb8
z1b88b9a29f4e4c35617e06b0ffd64015263184cd0e17c94c4060df8386844d0726a26d1766e814
z79137f8db8e7f00d2ce1c9e29f10df0a70e46a028f5d4b2d308e7d69af65cc6858a7301b6355be
zad08f7a6cf05b9ccb5784c2eae7f74805ac06a6455a205590246b30cea8e2491dd51197fb9e4bc
zf9c3a0ae4d3ea9d032fd21433559a7ac17e52153ed5ae90f654a9afee3ac340eaafefd5da6a648
z0e31529cb412d06f61bc6671600626f8f933f71c0eab5b1ae71c24321d657f6ee693429fab252c
z9ab4ff1dd3726107412f5aa130b9f1790434322358d93f82fd0b46e6b6d9772f70d3b99477118b
z27964800e6339ee5fcede3206799aaa11c2e6e70bf1bfe1298fb9ea776dbb3c1d741b075cf902f
zdfc77aa96992d9ed0f7328124400ac6d68305eed2e937248d29fb4c13f2d68560c23532d66f7e9
z7d9fb33765ffe4cea7dcd8ea971b52fb4a300981dee764ed7cea0621205af4384ed44917c4610d
z2e7e39df605c6c1ebbfb7292ef48184b6663c446331c95ca2a07496133c82acd927655b507b998
z36f28c5e854c828423daf3b2e7f909fcba22ac3e0790d095e26e68abf2b58c943ef781038666cb
ze970e5532b5707f5374169efc8028601c510f97b6c68d44c73e60ed781f599030a3ef372b79974
z11f442c6f876b1ddc746ccff991be76a17b4f6af6ccfa9a329727d395700c733d8b3b33a06cd8a
z97c8a5bff493fde48dc267357403ef78df8536813def6cc79b223f8b1583299827c6f65b2277c8
z9c43a9c58beeb9d530df804902ac464adce7a68e3a2db4b5a4a98bd793a829e3ce8905d354ca2d
z275e71b16cae67445a3e20390407b555a0202a6ac7fc20819ffa1142d7d3d2c6413ca76d0a421e
zb736b9c1a09e03db910483122b6e8def1ce5466b24626179587b6fc51c5c9d08e3b2576f0947d9
z3e79834876e2466338287796b3f94b87117e4f712e176cec99bed8fc642d98c2efc85e5519e0f7
zfcadb138a6b908902172853797b4f0c225e7b9af71a1147df19d2d70dd0513acb51b4ab8203c9c
z16febb14bd1407b060f38821ad4ef148d8871c0447603dbdf14362a4cab9413bf24c5cc841bea1
zfb0db6069c116e60c46bce69adbf796d49c9897757c38c63cc96cd9cfa5f8f34ed1a71cddad29e
z450cbb6b52a5dd5f442f05e1567e26af2fbc0c9c1e170581214cb1535bd03cb6bbc4e8fce444e7
ze82738d03af1e2545a753f47693e47f1bdbf7d3106e74d7749cf2c800a29d8c19644eb93ff694c
z9b7a325318e16261b804b6dcca9319372f67cf642778077c72b4181fe64331057afa3e52577766
z9284ac56b5fce2ed6854be12476c6328d71cefc44b266c4b21a28b94cf4cc0abf452586454d63e
z605a05659744648b2b7682f8950927d324a9fc2456f577153b7f9610ab752e0d374fdcaf5a79da
zc6e0704e529b5d6eb8f4ee1c8cc02764334f5feccf4a3b4fa7d3ebba76cff8570b034d140229b0
z1ead79e81481baff038b2cca2fee68f4c19576d808dd2cb923d399812beec303f2879ae84bfc12
z1a46055036689c4556cab3282cdd6b91f0b42ca295a7cf1f75b4908b3e724e175b3180dbbe6835
z68f5178a86830f445d64127825573ec4176625473e50fd761df7cdb6a27dce353ae9a6c05b0de4
z2102aa565322f3aa85fee7adef5d8acdc00074a50c625a15877b81568d9c40cd8ee20f4ad68b93
z2d90a04a5253ed027d16f89f7d90a64d743b6a1e55757482893a8105916d9087bcb0103c76cc12
z9446ef03e23553dd6931cf372307cfa53b24e4cac292009b792e430084074fb00738a4f27cbc0c
z6dd57f3d61c63ee00333d868ccee45abcf4870a3bb7c5ffc31f29d75e467fa364e2dea1b0308d2
ze21bcf863280c75cb0a5300e33d63ab98b2ffd82f4775fd0326f154393f61b55536d55cf352614
zfac0cce64e69a41eeb614d7e41d4e61c6d99a1b36130ccbf6857086e225612014d8ecb44e8aafc
zb0a924a1f590d803211f1f03786964986b09cdc32c15751f907301aade17191684c579b4dd10e6
z44a96572b413e3a0f02d2c075337b3f2bbd696de144ee173b5d30c444b70674986b3adafd6c6db
z1a8b22ebf9816d7d211b4c4b9f40f4fdb66fc3518a101ae7401c6d53651111d85c75893753c07b
z37c7b7621540839d03ba4bbfb921bd1fecfde2f3cb4239bcb0e559bf67d45c10b16d3c4ec63f42
z6fa79d204238ad2242fcb8de8e230513cff1fd7e906474b8bdeb49cbd664468e03d79209a179af
z1a2add9851b4e9966c884fea23b48cf223733fb7157d8275a2ba1b1d10cf7c75c254fa8df26e30
zc1e419d514600f041e3ce3877a7b3281436aa71be29b8e30dc6d9da92868b2bf128e0506cff2b3
z92a6d3eb455a858d35c946646125446c95bcb98666da036910b56f7a7e4456457fe57238c96f3d
zbe5b9062a57ee1560e661504808622959ecefe81f3132fbd6b09d5940fa57954f0d04c06e998ab
zb943f3139107cbd2df206e6e27cd4d27ee6559c986031dd095a84ecdcafa9e4c11094ad1e3d442
z94011e4cbf287d8921a274036bd73d11490267a95fd2601cc744d8179fe63afb32840fba08dd0d
z9fd133613198d0182fe63374b63b1334c9cd8947cc7f348aff10acbd71843d5ac992cf70145dc8
zae2d615e7d50d2fd4253b9d3badca1681e90caeb9d7bac939ab12fa56b6863e5982cbb775be07e
z7edf9e493c0e77e3f30c2c7f5a2c318bc0904105c2495d893faeed3e938c74ec874d39aa86916b
z9d6473f3de298693c88d7c5b4a792df199ceb1624fd595cccea5d402386e9b6381f095145a76f8
z73db020711f38ddee80f8d9e739a7ffbf60a8e33be7c20c0b1f5a4a9024ac5e8646333636323dc
zdf209621833539efa5e3474d59c0fd32eac6a2701602d0371a6abc1212b78603a0537501b1593d
z2fa0ee09dcd5930561e4b7c5341eb995b900ec59dc6800785647d2d68b11570abc8612c9d44598
z79a770e6e7bb9caa26be878bb77e7fd6c653a669d8a91aed01877fc9ce5530c4d2a1f6e9da7ffb
z4e2c2ff5487b33d22fe5f19611bed26256704e23743e6887b72dff25cbdec3b3aa3225b6001491
z1f31fcc5a36fc1391d85f99ec3acea71cf01aef5e0c156ab9515d1704f2b7df59e1822e65af71e
zfba8cd1d651540bdebe4baf96489baadd4bcfafec47644c8b7d99bbecddf7bd9465a4fd32a6066
zb7b483ba7731d250f4b870fbe71d7a3576463117c7a36c332b058822d8579b75ea1c4166068242
zbf7fa44108e659290e8ddb480d6864089735893cd74bf71ed2323a28ee4cb6323a8241a0dc3cf7
zbdfd1a4236dd4fc50b39a317dfbda4b6582c2743a0e9f04826674f1249dd192c0fb91e4d4d88d7
zbdbc75df816561381bd6831f0f64529c922dab618e6aaf18be7eccb088bd9fdd7d31cf2882065f
zdaec2ab3c1508fadcdcf060c47603dc6ff237cb3a150678a91981b4ab1439b284d498f1ee73f0e
zcba3120b55ca76d42494881ef4e5efc778df3bf7a9f0a5fb9765d961488d31132cd82302c08365
z43389b7366da41f2a84831bc2a0a785252e963fc1812cf0e5671051bdc76be5265681108c46a43
z72136f28404a2eeea06eba59922e76f35a16514d0cad63933dde1cd3a0f0ab5d82da956246bf5a
zb9cfdeacea38310baac18f4f6ac10f07268f77f17d1fe40c2e2b025a940f2751bfbfb4d10f6138
z393402727d43bfffad562c4764751196ff46ecb83d2d241cece54380900f7d7a60430990f3ed9d
z89c65e5055cdf7b256fdd7617f16f30740410ebc9dc16e9f0a16ee1a2d356392794905e3a36884
z9f83d4fc5fb57de41a07ce3131c1b0c67bb21e15b02050d5068b5575e5dacfd86a47fc4ebe9ba6
z863458b1669ded4800c2c7d92aaefa0cf4af13c673def8cbe2fbbeced8096f820a1a72f8260135
ze8da4c166e10b30a7118c0c9fdf01d65f53dcf412a039016b136d91ef77ec7e8aca183e2626517
z911e38441ea7aca7edc8e794b77b7b9025695f8ca6f2687ac0d97386ba950584ec9ab0efda89b7
z4366e1a05e20f4a5775e8a9e5dd95ac5393919feef88b630dd8b6652aa3e6b1e2bfbb8cc96dd41
z7eaff76eece80716a50e08b734540e2c9e2ad1e8097e06c74d84999bd3e3513980e081330e58f1
zb7b66882523dfad04482cc8b207d1f9be8e80f3be22970eacde9704177a041209cd21b97b01633
z84045597268d2a41cad95ec573bb3315e02f731279000a83f31cc5679e756485df00a9d2d1610b
z20fd2fd28f64d7e0ade72bab85da3e38d2de8bb9d72578f3941c59f7f95321ba94754553390b93
z848ffc2efc3bf606d3afc245195b208a5ef29708aa30102227c75715c39a9a57e85c78a5e6e5d7
z473744236c2a8566005c07957d263a028dc0d6ebe46e85919a55bddbdbe8c8967fa20b8d2a327b
z022160eaf35f29571394fa40911e7e6680798efe55bea9338d75f5350385c611ce9d18adfca092
z567f7aefe39bc3be40ff6b32feea02b89e4dbca627dc6da01f4cdf91d53252d805578a2728902b
ze2ca106644d903e145ce4346eca1cdd46714b20076c2f109c1a06b0d4374eae2d5cb18c4adb339
z9ab3f7f30e2eb0d406fd40fa588bfb3355ab66f301da883574c2c95e617cfd3b78d217890a9178
zf29893bee71473b12ce228bbd29a91892cb86db20daf02b0d7ebca6a36bb04f30aa39b185aa488
z7d9b8ccddd9ade103b4b8fef2ce80163a7fd8dd91541dd5311ff397668a9303919f53bac7f31b1
z88d7b4ceb84f92e63736f89c8e7e79b721915a1f7561ef64da9cca3e6bef63af236665fd05323a
z0dfd7fa8d82b7b4eeb3fe4a3e3bc08c789cec94925331dd965aaaad5400a01e38ab04a8c50276c
za6bbbe9ccbaebe3227179ce4d5730ec7f8cbd162affc0940ac7019ccf6ec3522dd730e36d43a5a
zba6b7acd0b217e7640c73da554ce12230b50b99a07788a16e67c0d4184bf0da4080d45099f0ea7
zaa3ee46fef1f69e9e9963a84ed7589ea8c976b48693fb20ecef7288ee9e0e8ac900edac366c62f
z28994b9cc2a2fb77156ff4f27231709425f7665e9db8efbe629841aab374a3a711477b93c80de5
zea243759920511d72637966ebba456f2b4b34404fda5caa01d092171eaafd2b254d975bd49eb4c
zf96fe8dbebf3daf4ca240753a592bd8da1f2ccd6f7956ea1a6661a8df85a73f5bda9aafa22fef1
z619af7fdf0e881341f0894a750490020a8b1b64c2022a2ccb8aaa109490edf797a9b3736c8c0e1
z736cad922acdbf96f5537cfc48e81199866ec1e55c0f7fcd3dc136b3828d007900140e32806217
z6fd5fac4563d3fc3e12e9741734ba7e7fc7b702907d835ed47e04b1aa31ff4dbacf823cb913356
z70e9c1613f7f349255ab0eec0b1b6d1e3d121d70b126c4ce568b60bd08a91f43c8e24776182e04
zf8ed6c4c8cbfce628e1cfef53821636f51094d960d98df8ab5c1f0ba5d4b51a60a4f3a4fe62ac3
zba0a2ab2f1059ac7884ad28709c6de5a80e9e000e688985e654519858a7054b130e385f0b06f98
z89cb42b61b0511540298af4758832dadeb13de4dcc14d47f20ddc96e3572f8213987af1c221ebc
z5bd1f2aeb7e640f57f9e93021661da703ac0a95f47cd64da16a736bba6944c03f3bd88477a687e
z133f1d8f63c2d5934200d88e9c91c4d845daab94eb7e8ccf1f593512eb368e4aaccf6083541705
z5d62a2c8c1568574f76341e1eae3fc24349609e07959ff36a47f935fc4fca94b0b0ce77986342e
zad989356d2c6ab4ed74559b7029f5ac4d9849ecbcc00c792b6babf477f71e4d9658cca17eceaaf
z32e36f194e8c6fe8ffed83c603d2e3287c16cf88745b9e7f1f74fa4d66048668bf7b79dbae873f
z47ba0b7e352790c167d39727b64fa68c1d1b09a6774e27eb473d676b68fa7e7adaa067ad60c977
z567a709e0d5257978dfa229ab4d850eaae1e5df8f5d62643207e36cb72758d2e3e9c800d5693ec
z4f39f58309c8459f66c535739772e28ffbb7db4eb960a82c14fb3158655551ac2ad03994443e4a
z58ee62fb160952c9a0c038591599ca98db9a2c90cd628d1a88aeffec58398bbf688083a466d4c1
z38f0d4fb8c54b28ac79753c03c82011c0154bd67191754af42d0516b49cbdf412bd46ebd181ed4
z2ab44af052614d2b60d87c2cc35acd28576ba72d9c4904b60bf8aff0c2ca09be9a8824b9e3c8c6
zee1d57b1f9e6862e3f745b541f220400ed6b31e9f298822d5beb863992abd6b1db1f917a2e8512
z232bb48433981ae26907c03c73db8fe148f43f87c3b240d44170837a709b0189dd8fd73bd0ac2d
z71b968e9dc7d233c6469504206fd5574eefa2f3ae7f08ac76352c18f1d9da2836084c06c40b242
z537e5ada14125892345f99056b151a61cc7ff7801315ff7991d1b565d3ae02d6796e8c9923ad42
za5928fd7c1743294b03b322e3e550b0225df33dcf7fc15eef4d4edbf939028314a80c70008a909
zd1f6a7a774200adc2fdf5df745175848cb792b39c0d2305ef66117aeea6c2e48d83a1397237084
z3ef27ade92fb797d104498ea8ece8e118207a1fe2d1ed3740d17017a12dc3c5a870950c44e5dc2
z61a2d9b40e7a9da7fc72b8d123c78394c3cf2fb877fb052204b7bdf4d44b439e5c975459585f79
z9b9a6466812669c5706d6e13955bfb982c2df7b301c3f82aa55c3d21c59d14d62ea15da2ba3b0c
z763d8c24482d62ddd66363adf66aead8f07807a02a4ce9342365fb88b500cad4443942cb72c921
z9732de9e71288cfb5e3e25f090a9e536546aa361857c979ae12846e1e3540991c3a9ac0b1d10c6
z329bc118386139419c689621331c742ef7955114617bc4d3879a5d11df016166d471a4dc05f300
zf398b294d5126a73099ee1fe63c47cf910aad66dfafae257874ba15380c22778162e7dbb0e5534
z04541241e4b15f2bbb19e7b95d74fa1b82fa8648763e5971add8e87fe929fe4670539c0b8add5e
z3dcc774ab78c9b2a82e5b1cd305d05b72b916cbb65aa4adc29abf3b0568ba43b875eedc53c2383
zb380fdb786c3e8e66f61d8aac252ea3fdf3dd6bea4d398135027b244c3455a9d72338a12278719
z5d1e4c0c88fedd5de90c9e759e4d90f62dae52622ef56baebd4fd5bae1797f7cfe9b8a62cb4b12
z7207fe8b4792e0f06f14eb03294e459e3c678329cfa3b6a04b25768ad47292a8a3b482ac93e23f
z92ef1af9e42014eefc318f3b689c0727ef09a6eae1abcb20e71649c91e72530eb3b45db3e87528
z38878d8f87ec701fc6b2c7ebb1092110a5ba7b97eff30b054997aed6ea537bb468b7c35d55fb8c
z107ba17ca9a13be0e9250a9e7e9f695f41d295c42e0408c28f877e39c817b0303b0723188bc18a
za7a747b9b6c0c844231e33a2461ad911ff4227e8b283244bbaaac6838ce19c371208bd9c5801b5
z9cc4b80a88e6d222b46eedffda1f4d97ac94812aabede71d992604529194c0e5bd061de27f579a
z910e4b182619dfe7e28684591412e08fb3227a729d506f921ef2defa59432562b43d5a75bb9c59
z26b0dbddf6028a685a06efe6d8d9a61433eed41b5ca680368982c2f5a1b45beb8f90fd0ecec1b7
z8b63fe5a0efe75705b230a18917090f5a1dba98b63e9959f1569b8b67952e56b6672c06d88ac7b
z30fa4f7e83e18e1790020e62e66e33eec270a6d1004f8af48033f24fce4e74c855ec4007718add
z2feeeafabc0ae72f247324c0349a14c5022999043f8110094a96bc786c64b5d22840fd69c45d0b
zc15ceacf21735055d4c68f24eebab6714a2558d30127f2c4d1476660d29bdbf9a5e8296d305195
z985a4b4aa41db3f8c5dbcf25b5ccecb0567e367ba65932da07c92b23382a43b4fe211ef416e77e
z684a2e116e9fe1a40ab9622f223416f63c0a9df78be88edd2845b7710a162d64a84a4ca4164485
zd0c58cb294c7e44df564ac66b79305b25bd540c8a2c09470c72f5a1f178503b993f50f8f21dd82
zd094efab5cb81256a2dca68b305363c10d2438bec3d64d9543d76c22d281efb8b11135f4686361
z87cf92bead5171edf3da7703f3c49c1649fdabde978c3898b6cc6c68a2011f002d083543402786
z312930b524ad0e0c34608f0c036ce85dd431a1ee10b6b1b5e2066612804aaead3ba3145a8f8636
z00068c7a6e17672ee434735c32b481c133bb93dc94d28d487d4c417de762c54fe764bf4cd81dfc
zf34cd2257d9a5b17fa960ab82c3dbffdab3d5341627619b3b3d1de911c6a92e52a7e7be31f8626
z1154a1bc13b8d67fe12123ad839f14f1763cc93b67f9112f3edca6f77a78c1d8dae965a8672189
z463367691c899e4379c208dfd184de05d0a84d84e233e27091e3270ed882e02e4e2a3abf536812
z6a0867bccb6c816671546d69ef73472fc42060fe711af2b153e625573da15f4889f649486f54f4
z9d845bc65e300c88925c98500a8bf1d2c7283ea523938ce4a247a0b55925a85bc5818d321b2557
z0948786b4c3eabc6e70a45ef44ece409855e1066631246e8028afec396a5afef2fa26d36e7bffc
z4544ba03a6822bd0a4be98ab8cd96917fccc62126d41731e9ea0d04f77733fa727918a23a9dce2
z0d6a0d8c317f8300911ccbd6383fa57707f1fba57cf2333937cb2b0efffdc4d0336344bdf7af3e
zdb7b52b602ceb1cea3f44ed5371301370803a02158961cf94e38e82138bd29f5015c507ce85f8c
zd12e467c6bd8b501cbe1dd89362b358389dfa1a679d46342decd61f7c2a9e3fdd656edb285d529
z110dccfa87adf99fd708aecea6a1af59cd55d54d907e5f5eb45972ebf2723f849aa3c75b798480
z04fcc98a65bcf8ce37559e4470386edfa2ee6c5d3359a3a2d96d7f2b79c06462652bd3f7d27928
z1f2f3ddf99c87ac3a8145fa878d4d85f4b3c016688715294d4939f856d31c7699670f1ac66e8b6
z6a5f4792ad43354ca4ced9cb5303e16e600ea273ef4790c49e6407fe2fb89fa7a36a01bd61a15d
z001f6154230b17c218fcbd52d504ea3ed833ecd531aa23477819cd1837c9360bc8ef3b81b63e6f
z88633b337480463dabddfddd8746610921cff1881dbf07a5b2119c4f025178fabbd0b11b193704
z32263dcf4d13c9b2fb6f59643d3d9db29ff977fc3ffcca37152a24af79a2a2a7ad87fd0d95960e
z6456730dd37281cc928196731b266848c8bab3abf174cd1da6057bbfd1712e4bf9ef21a55b0afe
z875324a140a5b770e2a2a7c2dfc6cc836777a6d8fbf1ce51a378bcdaaefe666eb3aa2206352a12
z8bc4619ec45dda1a8719fa012b215aaafd56b4ede15207b4e1fe8903ea248c078ae4a83b5caff5
zbbc495530fb4c9d25644a89fb1eff234ce4d420656e18ba062c1524f2dfefc675499cd3b3dda1a
z13715a2bf02234e721d511db67cd3a4307e060e7ca7bdb98c3cbf3066b5ff25c58bb535185b142
za2d147754c5fc29794f2c190a78727b166f2b308310df1e5fce15057bcb7695ff93523004e29c2
z269bd06c3199d302712aabecea6d4b118cae7bad79f6128b56c77cb9bb1fc6ea330de95ca961d9
zc372660d3f9500131cfb3886e7c7295f7b475f615a72beed13a7e75bda952484e4a8fcc11af71a
z4b9d2219f0ee2d4ee71daee7ed839784aa59c0ae03818c254228388fe8e27a4b211ef40b1fd996
z1f8e42b050eef841e9a56ead7e71ca7f72649f184e27969e1d38edb0ea71bb9243f98743117459
zd23bc6b8b36ef64a426bace738ebe9bf8780c6440d4127c46d1926c47d35bf82062b1116a3d241
z90a0ec6e5ddaf5320d8adb9e4de6c821662773d9e30d41e305648966f263541141c158a8aeb762
z740a9557c610438830aa6779128a6a2ca67d55df105ccdfb854bf6688f59cf2381ea3527589791
zfd29dbe6de13a0fb7a38df45734c6dba0c56e4704b6ee09fe0797a2b9958c189ab949837da0a1d
z329e77eb0b21bba5e625e5eb0324180e5765a49e073b1eb4e700a8983fe85c96a52a441ff6440d
z7fb67c00b19cb9f9837da2df63cdc01f4e5d68d126f8f2b9f611cc1a8d28ff21b0db43dc9f51c3
za77c4ca478b644ddff5fbc8b14acdb3dc0186aaca9d813daafae0cf289442aacb31148f07adffe
zbc4b4fb81364686f3bb18255cd4e9fd85a6ce568103292676f01d3810f41300ba103cd54593726
z04293c2fcc13b1c48064c1a3df399360b9d3d5259f18ce530c399ec1a8e97ab7f527b4df7340ec
z4078d12a016edd1c20f444958f3acdb4856ed834e23585623b9618f80ca76436afb7673676f56a
z62c5efacfc4cbd600b2711854bd045159fe4b0273b12e96714a002fec2d4ba1ac796d7d0d5e6b3
z10741f304c3a854a1a2e14ab8b6cb5efb196a2001667e49fd2604043da8e96449772585241ed49
z96aff36c5bbb6ace112b96498da3a74c36531fc2da80dffd105f5fbff21d398d637f99739bc6ac
z118a88752923ee0af93e1aaad06cb1bd58da7aae6da00b08adc9194d4209fe13754881e7f78019
z257723248acaa9eb939cd77cacc946eb85ffd40864480e65ed93f7b439306c907836dc51dc2f0d
zef62f1734d54c49868d4dc6d53c4e9f2b75cdbaec9239faf9f91182476e56ee42d344f3e39fccf
z08b789ea0baae49453146d36f0aeb1b61410ddd1ca761ff99692bbb733e1b214ff0588f1116481
zaa5505b981fb184061f6728fa44d5e69e848b4975ae71d73d83f1ce6eb4c761e8b77db6f5d6f81
z0852c162663a36ac54fb16bb6f32326810ab0b40e92e8307245f0c381fe1bfca16c3d32f22bc92
z5fb07cf9ed5cc74ea09bffbf8dea2fd6f435747f09824a9b7bed1d847c26c58cb2410dc9234eba
z366b01dab78491dfebce6fd904b8b3e4eb9d3466dcd047b1e4d581f8b52a456be7e5a01ff1f895
z3ac82b018863cff380194edc162f7ada0df5568074cacc0157b95a0f70cd3fbb7bbf8adfab6b94
ze01712fe4e9ca991ac0b7685fd6f1642476bee70ea235e31a29f5b0e5f6e2405bdb3509e52a07e
zc26e46bf6f98150decaa998b8d50a1bce900b0b5e61641783517c205bd0ed2312b0207cbacb2e2
zd712c9330ee6b871de25f6343008fb5e416b970f6f65dd65d72f4bffca69766842087a73263016
zfb1fc657b0d1a278af713aeb2bb3b8a2a80d7e0fe1dbadca1e94865412c55f47d911dd23bff92f
z658407cf96619608f4c0e2316b89d8287a8052dc62f0f1212c394fb39b8edf093ff79c20257ffb
z37484bf956da8205b4ee6b7e628ce44db1c608213a0a55ed9b627f0e5ec0484989370e0635db9e
zb38f8f60b99b8cc0e166f5583ceb6ba8776b1d99748dd737d4f3e6d6e46904f5beb025dc82c68c
z85424d853a38304e9cc4c7a014c6142c74fb2fb3d2e41fec088a1a3ec180388bec32e986c1947b
zb9e7df6221dd1de11961ce5c73f8f5d227774b4ff1655c2ba0bd475941f14d8186b0dd06c2dc86
z2da148b3b883f9840836634b83582a291bb9f9a772249a6021923162027dbbdd108e52f93cd32f
z06320400ac6daea83248bb275bda98f53ec1a46d86f9cd3ea013814c35b3f34c84daaa1780a51c
z4d1b9e176ccff59a130ccbc7a36e3c837e5a4c24aaa9486de92f840a2d8eb2e4f462062f7dd84e
z9fa81486ac57056bb80468d848e4e928cd737f867537b18ec29432a8dc95bd75d59dfcc0dc6f5d
z9096c81a0735d56361df5916085116e2c2d0eb2d6612f60d33dffc6b52999e15d17522c8625907
z446e4acd5361e108d32a8e153def05d69eb12a06f32b6b13ceb65941d4de65b270af2dd1bb3922
z7541daff8a59a2c8d734170e1929c23a057a6e038d80899992aafdb91063891b59cbfd7cd04637
zea800dec309bf79d1e5fb32cc1d8467b0b47b7fb789213ce50769c0a2e4e6ca6a3fdf25a32ba1b
z7d77e95daab4f5dac51e638c14eb16cc6f0d0e27435a89712b5dbda455643c4a56398d57b39ca8
zaad55992052de8cb04074b17fbd828c020db42edaf4edfc55ba81216d3e6f6689e9aa563a2148c
za2dedad8b682d778c58a4d23702b37c7022dbcdf51493035baa52b4955dd8b52e1c2e32dc6010f
ze5bb952652c0b5f13f1266bbe64a5cab7422cac143d716171c2561a76d2869c42b807364869d0f
z02881bb98cf31845bc185c3a5763370653e4c91586770234844910e854884d5ac643fde43e924f
z0c1bd0065b8c28f543a12223437c40c779df1d1948c45a1c85436496691e8f424277b25a6b8ac9
z233e5d65f4fa3083aec9b251ff90461b59ba489b051acda02b700075d0cf060308a6f2181d9565
zcf6bd1b558cb06b6203c5a38d8840372a2b7b3617cbbcbf2d7966abd1915b2a0a85921da862776
zbd8bfa96c2fc3f8b4c46b2ef77548d4d6d85a9e0f46e7257ed1db6efdc0c7eaed0499b40cd0576
zaa374e1af4b98df3d02ab7379a89cf1db333231ca33f31b8f4b54fcb735e7297a0461439d08290
z0acd2b45662854452287ede5e162e6aaab355c2c7b7017fbf491deeb3da957e5cc16ca4b93929c
zaa0c0a80a0031db973e63317ae24faefa9026c37703a44ae6954d88bab005457b73c05b3664402
zd29b100436ebcdf4b24aef3ce74a3aa8b0f18b3696698a23dddd8c12c7b0786317a38c9674ff74
z19a342736bbd93326ebb2ddd2551951acd89c7ec4c3ad1cd2052ea19406a6d4cc7693151a22330
z69fd01f6293c824914962effe180451192a10cce2a4a030ae7b87e971904e84ceb34e7b08ab663
zd240a3e8e25e488b03712f87be7975b291691bca4c4511a547097ac14caf24ee9b73ab93e66056
zc4942d289da4ae2cb186502d90f49f139e1a30f86159843cd81df8af265067d63ff867d2dc2361
zc3203403bab3ba19571020a2a76f93a8d287e83ada5b2f4dde8dacc8e47e63ee7d8b75487d278a
zb86de5a026d132e5d7c1826f442be5acec8d04bf02390e416682e15e89ccd351d6c759d5d63f2e
z262d9aa1d28819297c1963ff9ffa0cdfb0d7fa222b2a6b43303bf1e89f724ab2b3ad61c3ac4c57
z4509090d5d62368c842f90a19e0e54e19617f2355d25b110ab5c8cc641eea880511c75bbff9095
zc9f29b22c03baf057dbd86dc87ffe8dc085c3ee3fe50a2cc3623b7a1ae1d39e5775dc31f7feed5
z96d91e31d55401fe783623f6352bf714eedb7e6908f16d0e636f0d02604a5726180de9a1beeb58
zb96315ecf7b8a78620d898733839edf0451e2b4a600ce01b8a6e268f8e183e7595833173e31668
z6ef705a28a8a027adc76114015ae8197054ae1cf1f32c870466de1a0baf0a3360f461381e159ed
z3598c3ed7fb4badf9055ec55ccf25166384c32ba347e592db5949ccaeb594eeaeef945431a4681
z6ba5e2e2a1d7f80cf5c504c2b66aca6818b52f8305c1135209e09f799d7d49720aba81ea6883aa
z08c00810e2bafb057984d3b22d40b2b13a0071441ca1f1c32275749f4315c7f4f96bb3427ff3be
z4ecb34cd56896b1ad68eaa05b34e228e5bff56759516e8bcf4619cd64534b8a50cc4abcd7decf8
ze99692f5e2dc1e7977eadf29428a4f7c65bec2694424bfd7259350dfcd8c30374a054d77d3837f
z8fb034a2dea2cda8671844190583cebe48438b076c32ab0da6a155f6d1e6e6e1c6982066204226
z2c52e5d8ff0df1af2ddc5ca842870ce78504a52699165a567eaef4bfed6df5967fcec602938014
z56fa2326d9354aae665a4290470061922b71f1b5b6455d268b8e5ac529c7ec314bca3e297e9d5a
z20aecebd620b739acd0bbba9814aac587000cbc1db4e1b6337b3012e7473bf4eb3447f8543fd3f
za07b2485a819ce6fcb4d8687634fa655da7b18fb776a3ba276f0bb6e561451516412cacf6dc300
z2846b6b5a834f9be8ff454e4487f8693712e636045c98d3f5c6c4237fa2a52f83c4cd8d51914de
zeab28a26a5b5f8ae1063098cd2f342435992fe547cad99b124704f61310ae699640796828b6140
z38d1f024a1f616eb62ec36da6bbda0d62eb1059f36f76e14db409c7c8b86c79af949b89647c6a7
z0aa0ddce90a56a2e71f00e9539c0ebcd455626c69923e8ef72c5f61afa612c1fe76d28f3bb501e
ze14c93891513bb85c219ff7fe23ab39390e07537b8affad8cbe3662b0359e76a0c2b6633a057ac
zb401f412f73f57d54cccb335bcfa4ef84228eef228b87889d0e0f2e6c610d6304d61c9886577cc
z1338eceaa96049b75b919258dcbf50136e7eacb32e81024528fccd2be43474d7750214d54d465a
z86743f5b4d09d9b3100a6bda2e2adc2fb5d0443c49c7ea83ce302a75e5e87ce4d4d20a723c0db7
z72b22cb26f032281ae2335c8d21945c4a81f07f276d06f54c2b1f23c8d02f5647106fdb772fd48
zdb9f93b3c7b6008599dbf493102a5759586940fff67d26599143dd89397e355ecd332644948200
z436eb7c666e46eb8c3ddfafe04a2689d6875f65387ab9b3d72a297472269de6819b9b10ac90179
zfd72746add7d0dcd4b1b0206105c32d718e13c74de47a768662a231ebc2b9042998f66d83eb3c9
zcc85c745e39fe3355a58697965d6b1c8a0fa60b4048faaee5f284b8699c53452aabcfc81893f69
z33a9815daab9444b164681bda498d5dd945b622a131c23611d357b8c7c68360b663341ed1a11ec
z057e4c397eb100989264726bf42580718efe6e59e2032386fb2429bc641f212751cfdf3228da19
z269ec76f215a730f81fb7eca9acbeec5556396442d9cfbedfdd02770fc7424365fb7ae9bcc5d79
ze59c58f9fb28a5b67c010a9ca4ce6f04aa178be2cda0e59cf8de2346f1ad8ac8263dfd18a5af99
z0e9992ff8ec0c6ac230be3a74aae09f1a1dc6007771a0756520f75d75ee7c9441b60a0d37a2986
z5a0e7e5aa88dbd15eac0f78045d26886cb6e2475136808df96d124d04c98cdf3666d01ea1f467e
z9db8781d8b8bb94cd03558590df7a84573158005480e582056cd04c9285b7a421c7c792c945f59
z2a80dcc1ab4854a9b7e35b91c6277c0e6c1a33e58813fbc428cc75e8539a84e66c5d866c1950ea
zf8a573f2c49283147e4065d35d9b721761126e2032d59af0a37f4f76cd96c51c10ab857ce05dce
z31f334bc23c2af1131ad109959b4c01437c84e986e5b7f5dd011869c8fc9b7020f018e1d3cbe7e
z85e4d42d1fbbf247d143f31b97fed9b3a45b5a4154465a7b5f2e15db1548512e9f7e80a04ab2ba
za7a8333c81a761167d9eeb867b4d61e47d061f16517cdd6ebb58914c496c4f18deb477d7c2abd3
z78b8177bb6fef95a34c88f7ba22cf6cccf6ed32ca9dd97809efc3e47acf82ceedf6dcfcd43506d
z1e0642d1acc5e9657f510fa898dc71d422b02971d17d25dc440c8c5b0187ec06f02b2976fc5f1e
z4c78b768a09bb70f7706b3adfa63ecce2111fb0b87152f7e1bd34466f14d924246e9710a73f312
z6333beb25043b69fbebec459bf7b0335a21d6858be2e3e82d02803e30174b0dc70181117881704
zadc33ed8a8eb3d1f436f6bb9cf9b7b02907ce56c98aa514f55166c6b663f19df1e973ec8194710
z9790b66ea3ea90820e45274329cc655532c6eb580c6564a01e3e47a9935a5df591d686e7b240b0
zae4b3cba3cba62af1da8fb4b8ca9b684afaf812dc7d5ac7b43f5ab2e6b358e82792a55708cca90
zd2f026d1a44a0d74ded56ae4bb6a6f25008f823d6c9ef2d02a82235d1b0aa15324bf632ece777f
z53acb7215bebc8a51bf7f98ef3d2924cef27247244b472e32a8e39cff12e1f9836824bf2589a88
z32eb5d06087bd6564b5b3bce6bb1fa47d51ef71bcd157c926a6b292b507505ec06d9883c31c3d2
zef819a5af336ac55da0f0358a83f63976784d6e072fa78b72290383df44d7e2a5b666995c1d02d
za5b67a878c6cad87151b4571a35e7e360b67af970bc1662f51a949cf053e2cf55c11fe8b8edea1
z719040dda6062a90132b169b7aa22a5dac94d2982cecc1619a0e1d37bdbfa380a03fb73ef18bff
z75d0e78963575151dd149024b81d6ae970a5a8096c119aa882f5e43eca525c652ebe3693790c10
z19691ac7d1de2643a785c63911e01c5ddc5e75bddcd6e943d8ace1be495b439baba4684f6479a9
z162851dcc584bb940c1fea81fc91ae3ded9bd374a05dbaa7c6a7afb34caf33a2e3b482fe2331aa
z54231ec84b1f09b85406638d6652c8a18b77165ca7cdf3e70106cf5539b85f5fc05381ba1c4924
z76a4ba2731c1b302752a93e81123079926cf749ac9889b2712d2f0409878952fc8f3227c7dee91
z49efcd7c81a7422f41ce3e2badc394b26496618f1c95cc8a1120e4634b21f7ad20c1d0393f6aaa
z792bb453698b8e68b0b9dbb6f41a85b78348451f320b840529e87003f38e347385cd9ac7721141
zf6e16c9a00bd9aa4bce47616ea20069b5f88f20f4751b768f2cdcd40f76a3969d68d3c1edb5afe
zced97723ac78529eaaef65d8636dffa2f9d3948c957302ee5ce6bae75a2c490f44c37282f88d3c
ze650df8c0dc198b31854fe6c3a4b4b52992a6894578060ea9857ef9131edf8f91b88cb41c65134
zc3aab3be5637db53f9d087850c734d1db313674dc4f14949cff38d423eff854e38dce5f701cb20
z307c30f14836953bd3422638dc8b56339a5034a8c009b50bce89e243b0ef953ff11a92cdbf4312
zf6541e72d02e7c01765e757f0452fbd5ddcda29b3a779c5f6a911a9bd6a88a923188ab01d440ad
z88a2dd539251f73214901cdd6838ebe4efe5232a4cce499b6a0bec1fc478db28fe5307177c080a
ze9d18e3f76797eb9c00fb104713847e1036c175cd6d802b196ab359446ceafc7c9175e51b60a78
z8f4139817856cf9081265b82fe1d7f135081cf9cc09c85499d0eaecbe122dd1e53830dc28b6206
z281659823d5bd4f38342e33ff381ecb637f516911b641e7e154655925614c1c0a9ad01a10c47ae
z36eceb7f7b0837c9e4c35d938309a7c7c719b6926b92626cdc50d13bd4a0d71349e6b18bcea71c
z98f866d23e6275e100fd82fd78177c594d2f833417bcec331dbff059f37dfd61e587cb9f03edf8
zd3f46499ca0622dcab50de20dd87fd1e72f427c4dfc0d7914fe56d617920387c77ba4be8d2a97b
zf50ff0178e24a0b4943bdbe70bc047564f7823dbba603795f2e783fe10aa3112dd9699d4434416
zb268a9b97dde03eeea52dde712f34a37245ba77b6b5f7e2c52a0a7b5f05c029944458be9fa593a
zee8d5dc3925fe1fe228fe68137fc07ef5995ee0da1f9a596499c2567a7139ebf1c242ef0ca4b23
zb0c68a313d4373070ca9e7946b14a4a70b3f572fc8ac001180e3651956b135b32bb005d194fb71
z1e0c353df96c0bda4283cdb33c24acbcc9dfb29f8c7661318a2f5f96fe92e1df89bfb8990ff03e
z976d42b8e9b2fff957e3de14e4bf24043f122833f2a87bd901e5b24b2ff0cd39a04ecc1bf482ed
z5c76ff08d93f601d48242964144e3be354b2fe4ef1658a6941632d7435a2e60cadc0c5cb8267b1
za03c6c5b7520618e9086467ec2cf8256f7a938e1ca284d3775f181d01b71f8a82cc327567b4030
zcfc5af30f61dd1a2a36852c7b30728f52f3c3ecdb96acc8ec34064c3430ceeb436725cb8f1e68f
z81551c338f87b16afc748fa38a3df93e4a0b2fa7b9b9e30cbf9cb52a1ce2d448bec320b1f2c3e4
zcc0b7eed5b76a12cb4403df072c9e604ea12d820537b55a005e2903d0689e0f31e7b0797cb969f
zfdf93e3522611b6cfce138b8aefdd381060b513d49394c32f7683c01cc3d9382c77136116d5ba4
zeaa203de8065a778154994331202e60310e92fc06d5bedc7345be846f7523b5f45fd82f59a16f3
z7dd0c82ce498638adc71b49b803dcdf1f84bb84fe76e5261e9b7683ddeea35a7ccb83cc25d9699
za0249dfba1da62e849ca7079fae1ef31884d63cf091af94edf7f6220cd1b787670a8684e1b1408
z4db9c417b009df30b414c9d69da5a592058cafd986e54cf2a9ac0bb448cd776e382688d66f6806
z9fe390973febfa490d296c6f92d762ff50060e06690d4d7522c925eda2b35400f27aba6fc71aaa
z07bd00a13b85022b616961930929adbfc32ab99095d0cfbbb8ff2aebd4db99d8440e3d19d301ce
zf2c9c43f3172843d2a74a4996d6a5dc7f111f53bc2e4267802efcf71a6cdaed9212fe904bac8f9
z5024a56cacca246b8c8c85b9c995e0e17c7ee6f2dbfa0eadcb2601a4d70629742e9b4320bd2c79
z4c728a0c79906343302d57a29ad0d02e96f60602211ade21c67f797b5d894f4ee224120bdf7ccf
z642d1c754e0b839113585cab98c0e77f3a5b819c745085e87dac2b8158f2b5ac6eb1483142f43f
zd5d8b5e8680bbd3c69e719ada8ce7155498d4c547647a76c0508889c9f0d67f36111a6967a87b6
z55bd7fb02c282430ec96d2a272bcf75bc4cad47e4755908ce0adad3283e99092cae0b106efafbd
z453d4763999d73834f875a34cb394fdaa10b8fff2a6b73261acdac64c16840beb8e47282fb5ca8
z88481b0535f0ffee5d851fdcbffc7e5f562a615f5bae9dd765c1a97a3de03b8db0294464208b07
zda3c39b293ae4ce2ac96951214be909ba2ae049885aba9de2c6308777f03ff54fa358708dfc3fa
z8a46a4ca849b5cf463752cd38a0a0eefa835db573629ecd74f12bda6cfd64ad4020f4e32915f04
z8951f672cd1c0c2aa18c58186e12fefe340a60a7206751a2df10fa50070ca8abc2897a1bf6443c
z78a6adc9862509d76de7948b9c51dfb418c452c935637437dd5cd009292164471865ecdca5cac9
z7426a85ef4e43c8a7455f73f210f5b7de7f800c781efe9174ad15a4d641e39f72ee55a57f53123
z46bd14b9470b934db9a886db86d731d276cdd701fc5afbfec779dd0d5496d89c7c8f1809f845aa
zb7e710822832121c5321e511db76b02565b2093e8d8ec6f45c880e7571c3f0bda327347444e1b3
z1b99697fa04cfb711392560b1c11cd63d6adbfda05694bbd23328f7f3dd5ddf872c1fb4fddb747
z12bc504fbc401a1dc2fbd7656d2b8107f84b49fdaf89eae1980203f075cd153fc473f4152d0895
zcf773be906884ecfe5cf777d0944522e329ecee4dd66f3e019c234faa83b772ee11d2c8e97fcae
z4b019bb9cb2758c2029cd1cb029d6d600bea1d0473575f8646825a967912e7102bda46707f4b10
z4520e7caf5c8268badae79bb1e344b9695f4afef30a010d7d36e19029297a5b0c07f67f31bc973
z43421f60a2572c4004a7882bd1d5b7b5f634bca5e278f9bc300e75f0fd7130166b261225d7234f
zef81839a27156474424889adc43de725b1f8b317f3b41c8494b2bde31b682036356f6f23b8c917
zb47085114268f513086eb4b8814124cc034e8fc6a3bea0f85caf0285b83aad7b43f2a67cf042b5
z40e6f9db8ed935cb5db601c2b25df4a5c890b4c74d5ee9eba18ff7d0206ef654186ca878b12fe2
z288d8fbd3d56d98d860fd008f7fa88005129a19e06157281d056d77862393c365eb2830a599095
ze797684cf6126d6011034a7bfc10c7597419ba57d2c13c699add2da38441d5adc69a72e0588329
zd436042e714476a2236fd4e3fe746c4e8fbe1a3cb800cb768319ada664749ec2d4569442d6e974
z59c695dfbfb8e7f6d117382e784b7bd276cb08c6119fb452604a1d2f51a0ffe67ed1abbe064b78
z870cdc861e9c08d8b22b32ba609d0c007e091d047a02e70989dc52e77935a446e4ebd7f6b06ea3
z3198548d9636f158c427e0388ae2305c86b750d09d0bc13e645c08ba9f90ffb26dc7221c3d715f
z721c39156153d4653512dd1899c345f4576f4d28a53982c881694e3258ecdff5711f32b8edd495
z4bc8e455e540441504e94749253191b0e0e0ba38b6d0172d09cc291c4bc00b51b6ef861d9e87e0
zbe979329258223917cf5e2940fa392ef754ccec5e85727c9035455a40946eb6fe6ca0260867fc7
z5dc03286595c21affcc55d92177ada90abb3ec178f5666cc2c1aa3d2f1956262bc717340a77179
zff3ee8a164579a895b7fc440f1b3131f36aa23b39ab41fec750ad667bfaf91e8c3e13b25f1c13e
z1be11706b2cd3b8bc6511087dce3758ee369d103fe97311fad825544565704c7e46ad5c9c6bd7c
zea0970e27b8a486f584d3ac12ddb533b1e392501af2876642c504fe72cc281da5f939468860ca3
z47e11faebee48ddf3955e67487ae4cdfa0ebfaff172bcb5bc3401232c7da586f638c2422f4d1db
z99d656d9ad7b11cd16521bb4c84d23feb24805e5bbcaa76058c42853ef1e1b3d65eed97b79652b
z1b1e3a88993f309115ec6e2dc4fd282ed333e275e74cf96cb1eccf7ad9e6cb1dadb1c9eef3eeda
z64ceef986f95715e97a25f43cffa4d34de23b16e8bcac4c23061b5bb0901018cce509ebbb01e75
zf7bc85ebeae4c79eb7ffe5560f563805b9c1639c645799ea4570fbc71d6082977ebf350e713bd4
z50c54665b0055924661b073db242ea6c1c7b9030c423e0f2ec65ec0788fd7905e06e6ceb46481f
z56cd45e9df207d57f9232d6658dcbe5ef97a2f245cc56a781da9f963bdbccf4b00ceb44c3d7726
ze6ab87f4b96e3106f98b869950c1d3c5d200d295ef8841406bb18427401a0a0a56f88a382461dc
z1fb1cb07ad5fa71b85127ae9b4d9f5422c8f3aac1711de480f7953a5018326847b927dec962850
zc2f078bd23f890e30611db80abf4a544ceb771739ce25f8dae66bf2c2daa072bea8e7f31c3d8d1
zc73eb6d278e4bdd452056f34bc1aa6e86c90c906a31da05b8d7a3f8602ef05e3c19ff110e6e937
zaae4582b4ccbd5085d6b967fd154c20b5d6bad48c512dd5380898ab986660720b96ae580b0716d
ze6a94be7081d39763da61c243c58cb624476ca1c78a3547a4fe13953b2b15a87f478a2784eccc5
ze674812860accc2546b5e1dab36c832605b0c58e8c59642485ebacba609b6e7b67a8b64025c5c6
z6f7a9593892372e8621c1039e5b6d7cc4616526f748ab31014eb0d892d357edc79ccd50ffb8aee
z6e4e584ca0486f7983c6e7ef74058ef1188b82b1ddccfcb43e03151ad8eae4123a44ebf56b0a3c
z123af574b5705cfad005db20eec94b7894884a5570d27c17a09b0901e0c1db11ef0fece2b9d417
z41fdf288d8ce24d58431379edc6f4e8807d4dc599b7c27c060d97c8fdb99fb1574cddeb3182b6e
zf1c069fa89eca746dbe5b65a4df635c740c0d4d35a6fabe16a080314c2788e81a4517327f8a762
z0083ffd474043c6d2ec2f0775b5f309d83c7f70c870a0f71ed6f4fead211fc4bba7acf24961c02
z6955a5245c096ca8779eab61d8329fa4d2c6d7813646ad715ddc3682599a5cb885fabdfee23e42
z8a3caf03670b25182c353b3b4d38270518592a9eed637bd464cc7696dd8d31485cedadd228e379
z3ed979cee9f0539794383da79b0338143be0cc36bc693af717661ddc5258291379f943aa89eb14
z2cf30b28e73a0a1f11a1ccfd1002fe75488edbc39228704400929f9d6c47a13b087bad32799700
z4a82d2b7483ca01d4fd68983dcdf9e0e9a74f6118a4d0db86a5b1cd5f0a492e272f521e21f73b7
z2b22c589a347f5f495698528d115fd051d4b5cd4623f157ac8a35ca276e0ce0b5e1abc6431672e
za27274eec415921e11d92cab138740627a15eef900e9fe64d89d10d3cb29f2b19da879bfa8e6ef
z3fcc8538edb607fdb5ffedf75b28a53619e0c3a5adb2ef120eb3ec2fb7ffa08e41ab2135bfc499
zb24d755482d1e52e9ea6ae6c48311f54e712fbd52b8e5b6eda99e0aca6b1e28a6a683558c774a5
z19804b61767b776dae28af7a344f6a0d82a2152c540ec64b44974aa365e13361dba94e841ed977
z8242c6f22de938cffd64c871f9d647dcb1e1cda286246628ad6ff4fec8bd7d0ffb4e914e37d8fd
zfae3b69333a37af84041fbf261b41aa47762ee0dbb690b572544d448624cbe68cafb265814eab3
z42112893fd094664701b87676982532f647fb20e32a19194fffcf100e22744577da9f55596a500
z8e4c169943250daa2f820d94ac407ba61bfffafb319d95104eff5acddab9ade9ed7550dd510b15
z5e9d38f78f6f6c053f41ee581fd3b03c94a8624430f115f8673425b2753ca69782fc85dc7395a7
zff93ba0d40d5316eab5cefb6fdcff19d941bfa0cb6308e23b381a0038aee41a3aed834264b26bf
z49005ab27f0b1cb80fc7c69273a2be228fc7362efd14267aacb7cacdd863d262e49f493e265a74
zacc47cb2a5a8a72fad907ad7e03c8e447c6746b6521ebbd27d904a2bca22f0a7dde632d9d1d3ce
z50780f24ff58d92f618078cb5c3b4ffc3b3605c5df5ebfe337ed2cbe00b037530ce8f58ecc6cd9
z942712a77928f83f14567e414dbb91afabf9979dd16b37d7cc826cd395b6ec938699f3075c2005
zf0e80e0e76ade5ac40342ae9f9ae05dca724b516d9ffb5271494d6ac2eb99dfb9f9697bd366cfd
z576527cc08f739adea0e72bb1172ff3eb856d883f09d2677f8fd66cc6145401dcd5e469c94e7e7
zc94416a85bb3b95fffbca5e374272dffb949ad22a873a677aa31417ffc6037ea352e8f322eeac1
z6bc6834110db3089d72f9c18730c4cfc88d11609bcd86ecbd00fdf268e5fc985b70eee395d129d
za9ec936f6852a2d110af6ccf6802f4c0d327717d6aab10517c53709c0db4ab8b6b7c1c63ecc712
z52c593c0e963a197907a311ba0fd2e47a39e5fc279588eb9f5360f244167d83bdfa6fc24e78e84
z751cb08dfd143a862428be15017ff2f8a35716ea3f2d79ebe1ea8d7c4b469d1a0dc983b0142389
z803e2cdc8b6deb67e3d7e194806c153fcabc10f9b5040f469a8801e0cc309b9ac46604d4cb9a7e
z4f28e8ac44f89b4c142d4956282416ab47556c3e3252a88135b09bf37bfc7387ba704bf8d46ee9
zdaa7ae7d5a13696d1843610463af7083eb131eacef84413892664a4493f9ea82fd971316c1951d
z4d415a51233bada2c9146ec45568ee8e0f3ac7ea2e7e64f1ecfe5b281eb90e134f00e32b101ed8
zd017722071f337dc7ada0a5db587877533056cc04901fa97e9769724636ebbd2fc23f2f4842e54
z9288a4deb43665b4422620d4a42e69a8f946721a0298db1829de697be75e0172199a9474794c78
z0cc5d062f536a9ef1d64f6b6b322528708ede70eb4ebf81d244936654177598072725e026dd831
z2e85f1b94cc5d7a9555dfdd9693c976195c4f2a486e43f2f3e0c4d8a93da5fd1e6f1e3392f1414
zf4a44c719770450fa0f5ef122ae2ef1a8018b95206f622a121ed65b8f8d1a395b27b0f007c3888
zacb7ee10bd0753caaee328819bf8270e359c9a8bdc6ba2071bbd2c36bf4fde7d3d55a50079c960
z98649584cdc597b468703205bcb025f88fc3cfaf4aff0cac3bd9fa777f1af8b546386ef362907b
zbf26d645ba572e61f6b2fecd768f21e5bbcfbd60a98f5d582ef5af03457f861f2cfd5f3ec1116d
z0208d20de1291d33fc2b807461f9691113afd8144949aace1f471c345d9563a9e38f2b822a96fb
z94c8410292b06c9c8d57bd5645428073426633de244a8807445e50d6178e51cd54f344c8378b54
zfde8e760a7e3065590d68d5660013e269087fef69afdcdae815ce9ce7fbd2bd99f40ffe59814c4
z3c9adccb29ac52e57a51d80c5310b786eadecf7978b317232ccbfdd99832d589307807855e3544
z4f10597aede84fcc9a9588f59cd9b271b76f8d1514b5dfbc5f6576d7141fbb27e8407bb289be23
zfd3eeee46eb944f3ef7c99a8ef38706ed35aca384500e4717b644b6c1eeb4f910eda1cf6232f1d
zc73b22ac181b787fd7f336def0c707f7651514caa708fde8334145dd3f8cae4c857a4b5e809a38
za5da84faac5366a82c3783c5a12e1714c29100b015c6d158a75c668ec0d31c362fd00637befd7a
z0002114d4a4da690e3229f0047068ee8606c245419275fb07864cf3ead170f1c70ae5b5507c085
z3d6eb340c83f87c18db183fe9a2acaf84e6883f08b614b344281508782be24ff42c2575cbc88d2
zd12fb7712ea0429ed1c6d9222e18b204e697028de9f85a24438702b0681ea9c17a02f45159ea2d
z6f4827cc2ca5b8ac06fcb79f967ac5ab2ccfac14dfa184a4b27054e0af22963e290d19d25c87e9
zf683dee86ea227b7fec400b2d4ebe83d9521eb6eba7c5c9ecbafab5a638d3041f43f15535fefee
zb82e830c36b637815163aff03a3a71ed217ce9a97246a6c33d295193f7387c1aba061a042bee04
zbe1e1e1a1f08d0bfb1b6ebdd0ba400b83690014dedf8204353c2db497c0374ea5ace267ff0ef83
z22ebaa45e10484a3ff1f23fa9ec2f4e9eddbc61ee112141a614502df4239f7c03d1e3bd2fb7e58
zf4ea1a05261672f40249effe79c13fa802a0d95bc384503fb7514179566c8adea8b9b84117ebd8
zea076c9cb3c68ddd9216aaae3e80400485f546aba0621b31dcece189167454064025f5e4826459
z658712adac604779b7395d2bb0fa2dd987429a0f3066e309672d6cd772d617eedee86d9024593f
zfd4a5ee4237ff7b9bf1c87596686bcb03914f4592e7758a2c96db16e2a2d8031f52938cf02eb60
z984963e24625f4e8363ab8a81676899688b1b875f019a1937281be956010812e07df1f9335fd17
z6170eb4d0f21bce3080d9aca0dbf69256ff35e742abe5056029d2fc01eafe629947a420fbe91e1
z24202aa79f6ce39c22fd46f3fb54fc0a8ba2fae86b21ea04a6fb98eae741f7dbdb20b224ae0129
z6d3ea84e4c3f7a640b6d7eaa48282bee4b2c190a1f490feae6f450a0ac58ee762b0e2c308825cd
zaf89dad1de5bf3b613039b716e92737fb1a78cdf4e65a1f9f8b7ef4d5abf1971316ce04442e295
z49465b53e6dd98ad32232fb7bc146a840bc117752216c5e9904a77fc9fe9158faf1aa4215ac525
zb66191744572d7c912f2097d43b46fed30be3b2c3def84ebe852c2aae26805bdf9bf8e543a4912
z0ad1f8b2e584fdf777608414acd9325ef18017f280b49e52311ea7fb5c54e9afa505fe5c8022e5
z5556f58532bd5cc4b72fffa47d3a15c47408a36761ce4630049a50ac40c8934f63462142c28ea6
z3d53f350b51e13fb6f2483ba33e16cde09845e76cd632fbdd4341260809b10825dce7703fa663d
z61ae047c0710d531dff9fe352887459990059399205ea1fee506378a62352edaddac6f0131d105
z88e8582e9af8c83882cafde03fc6b5d4cc9738e927474eb2194c5c011c1674a52df181713e5789
z89d66cde746c3b547fb850adea2e5969e234507b8fca82373dee37769c1ffb13bbfa2a5dcf0730
z7e252e7308a9889596992614db9ea63f466dca29a170b58e987689209446cc341a3571580b18e8
z5d67b718f850d423db868a253691b0f15c0f442068a647e8a53fa8ab9f3a0640b33658cef82957
z517f8a603fafb0d297006bc8d2f3a54041248cca1ed16ec1e010151c5920b3a129802eadc240f3
z1adaf61d235c0526adc7bad01ef170bab69b19f9284d5249106c92f3335a089c76ed555ef336d3
z5e227571d08230bee3996b8d1da1792a6607e3ca0bf59410d20ac54eba0dd76f2a6be5775ef671
zc046a9a3bfb3529bc2dcc26e228ef1747422e2f1571d03a09670c5242e6068ceba9be84b0002dc
z6f3d079efa1f2b4c58aac2d7e980a0c4d0277a619b0695f45cf78222c225b6b294078618370a00
z547f27e65262f4bec738801b3322e6882c57ed482d22d04760ef6ef46d3c94f32ea9dff1c42002
zc5f9eb835f5579803afc9f2bd279828cefed23de6e4ba2ed4eb823c647d4db3f6fac3e11d332b8
z4ef962c8095162cf769900e534bbbff85b3907891247be981a7129bb576c2af3f2a91659bf408c
z0ea334d0e63f59dea63439b224e9fa96650dd21382f11cdabec8e984aba45f6d4adb0dc1ff7e45
z91b55681240af4b7c3ae249e46212e033498be81974f5e033abcd662a8509fc4406d45007f8b24
ze9a45e3f6b5048e067a0d2240c2eea3849a9a721139e70dff53371e346406a083f859fefd1789f
zd283c9551ff199b9eb2f080423ee92db9d10375bc8b299635d63ce3eade1b5249cf63b628b7392
z730dca10ea19a6cf8b4051f57eb2ac533d75a14f6f177ceaf3b5db447839e046a5d36b78e06b05
z5142c706f2e0d9bdfa6108476008bda593d3d43e68c972360077f0eca2a77ec40095703b9807d9
z9d5d00f93c3428e67eea1118b4ed65ca31d8405d894d5c7a1051a8bcc474859dec9252b152cbdc
z21f5176c9fdccc526b15f16c1e6c3e6a23159298f1cdeb5ef502b1f8b245a40b846980c530a5e9
z8aec867a46a786cfd3b50b68d9c7a286382f07facaa679033acca9734fec30209735f12fc12d9e
zd66f476af0149d7cc23360bbf898f04ef8a313f3d812b2a2425b5445cadcdd98ae7b87e29d31fb
zfd9e71749e9cb5bc030733c1503447fd1fdb8636a7a98a112356cddfd8e6ca1a13e5a818a0343b
z13a5d3cdb8ed3ffc3e6ce306dda04a0f2eedd6607ffdd0dc045a252a2b7c60a90e5fd535bf3562
z2feecad3ec9fabe8b49196cc30db3d2c59cd4a892eeb3c51db04dcc1ac0013ff9229e14d2eefe0
z49bec850335a4e73e4de5faf11b98b77be76c31bf29e487b22d4d67d53255e55b44e6527f5938e
z2ff7a769347d5bd5978aa4f2397192511f0fbac80f6311cb5dfa54325843c775fa67055d0db193
z446641ac7ddbc53748c08c2100886e146c6f017dbe75e40c959218cb6927825105bc9f5d37ff83
z679b896936bef91cf0b99c475307638917482ed437d57ff632fd2e9e362c66b83d863119fbc71b
zb87d2e537e69d84c300fb2d2e73a3cc4ca28ae9af2fc08c24e30fe483a0e82ed7f8f947dd220d6
ze6a3fe8f944d8709450235d9de2d381012c6d97c16edb8e3ac7716abf94b7f38f30863519719b1
z3ab4b86d4a99d675ccd8e41bb696a1d7e56c97c455f29cd4c28e9280aa23fb4edde3e540a7d65d
z08fde5a306c966226c857216729bc8bcb9cb7356d1aa61f62c1266eb25990a802e92ffef25e793
z94273df4a6876ebaa4bf0a0e5cd4e9200f853fcc7a1cb6e3ecc26c57f0776fd527ac2f41c85859
zbe0f042e3e4fe389abf2f64c402fc73ad60f44ea13d20ac412b03d079e4fa47ce7ad2c3e5b5d9e
z08648f59c9c14a82063c4b0af9a879c68231ae907a34f9bdc8e298a61e06fabef6aeb14db97f9a
z4704d5616593e93402b4d1beba3ae57717a04ab0cde4b7da6fb6b05b76b50feb8649d3560cf875
z3bb2500cef123a2515c5747b14af015893133af6b5fdeda902815ddc488c3506cb452ceab07e57
za0093d10086ff344235fccdbbea0fc7e826863884cabe3a8c9b4e19775476e40420e464135991a
za9879a997e5a454ffb7d3f1a4a7a12cf6bc9e7c15d91a4e29b297d151aeed9cf1bcfe93ce4790e
z8307a2efa0663fecf77b6937a463ab18a066e5489ff6ae29ed3ded5ecbde894b16c9922b660ac0
z39b99caed41aa78dae2774c2ee856e1e6b30c7ad4c3a971142f193a9a03cd65d236aeee28b6c29
zeaf9a1fa751d2c252c54b80c6b8489a670ea785502d59c24fe28a5a8c9ca0cf32776d785884ce7
z326033fa4ab02a569bda949393ba61d6bf69f5df62a57623be32815bbdc84edf9fa9b0d11f12d5
zca379ddbeff1bcdc4631927646c327a66f412745b774794aa316eccd46130055b226a586046b42
z2338ae92aefaaebd55d700178489f7b907702d4845daa67e74f339902a43121d8701dbe8848d07
zf71841df30d3d30c37f7f5e6b0a1567f7e130a1190651b60caca1af3b08353027d0af65e3551c4
zd71ed63fc75d957533d5f149ec4152a30beb0dc755c2273a188849c9408c24a645934ce16f1ae7
za8d94da0670ca9b5185cdf5407b6605d8dc32355fcef6c942e839d40ca7a60cbd17927e6f246a7
z856347fce4cc0067b1fcc33bf2927ae2cd5b9dfa4b8e2996d61a7d0532aeb562678414c77e8be2
z5dd79f9395a8ede2f64dddc1af496327550edcdbd5a5749feac7b1b0477f1093d027c3ab17dc73
zc60cfbbf7fc1ee0ec6496662b043f716dd37170cb99e1290931d48c0a5da5d5780fcb42bed05a0
z2d83c447c96fd397a2ed02ef70c56b3120392d4e5553080a9ef227cc5939299596a877965e00a8
zbdd96965c454fb2dda4ba5793a1d44bb1a3f059b9c484a843eb002bd82559d0479bebba9c9c59b
z3d7127962bd435bed0f7bebef72272ea867c5fc9a77ebb0130793ba1197e4ae78074aa29fee055
zc4891862a7916a38879dcd9db9a376d8ff47c6e5623e6f08bbd19155513e4004f8ce2d82716467
z24698fc3d3084903332f5cf5bc9ab0c27042f83f15a8399d3a08ec856dcc867740c2a50ded2382
z51052100f2f96118c9e9733765fbfbc73507cceb9f90b86f9d8119da5da8be1d0ea5e037567af7
z0e86197f932e74e3b17654cf58e81b4ab694627aa52b84e530ba2cc7afce6300afef86d79dcb80
z185a63c16681c19a8a392bca8db899e770caab90638ff4289c0357e4007df93c6b807024b3f2dc
z1ff7086d29149d1382c8f8ceaf46933098cc3718a71bcf437df6bef6612220d1bd83d1a3a0da7b
z19dec74681670020c07a03e4cf591f8471391a151d031107eb0b1b84b5ecdc20c5430ffebdef74
zf5cbba3eb4718eb80488da71ddafe0117c3abeb7fcd5425b2fb296d0357055b87887cf662349d9
z0d326ead052bd1ee58b48e322b6158b9858c6114082b35cc6a6b961d2779519819da8dcb410d27
z6e377a52214d6cc68026df30f6a683cd6039e70cbe281d19a81f84fe4394157abb192da8782678
z2778c151c2166c444323c2d17aca89ab65e76e61477543aff80b61effa5306f4e5b0063b37525e
z4b33b313276a7700f128d2951cbf00120422e97726aa598c80715368cb891907dcaef37f376e41
z84a997c7f223af856510cfd34ef1913337538a8dafa8342dacdf7aa12a59815b81b0420307d1b4
ze4e548e34bc8a3e3561d55c07c8be034c9524f4c110304b38a7310fde03fca8ac232ec57b63c82
zd05ab7845ad3d07e8a5f0190fd12f780a96c283657349a77119080268544036c140f066ea31c16
z61010ff74425d36858231dfded050afa31408439d26f4f9bb364d14f27821b424e6b008a7abcf7
zcf2859d3c38365bed5df2a637c3cb9261f1a63341c30f82dc80261eace0d617079c9928dd3f057
z93538eb1a9bed755dc2519f57c44b995b9bed9c5eefa1ab85019487eb1d257fee14f52300e2969
z1492eed96a861c1962788a18db20128a50d434bf908c35e50c3ec8e7d977d781bff3eb9c356581
za10006fee90ae0cb7bf352e5c804e4d63537c8fcff5363c578b818bb8e537a61f9e00e28de1a8a
z37c80cb146705c7e0ec20e0e21da80b1916ac8ac173ae991aac033a681532594f2c014b6baf553
z295529878b0fc8682818ff2bd44c9114632189a221e1c58adb1fa487006f729be4d7ad76feca15
z5cfaf5068bba671cd4493973f8fbc168a9deeff75269ae60089c7251936fdf4d2f1a4d32fe2d8a
z882171f131976f64f4a727ed11fea0811f216e804a95fd766361831fb07d61ab1535466dfcc615
z67e47184d92fb87fd6749f931f0b4abd28b61951c298558e4406c7150b1c0771bef209090dfcc7
z769378eb57c87352f7b7e4aab5f8f048f2a70276ecd752179ba5c29ddc603b73872c8d12c31dec
z506fd5154c1ccd7a7096dc4bd589826a6fb4c3854156f2f4da81823c98ade9632bb34c019b04e5
z675d621d985eeb7e80a53a1873b6945aa1873fdde7e875e79307d3ab29c3bdac121fc4f8fff9db
za57149fedcfc48592a8df416df0494c8548dee77147e8a024ea975eec4813127f5efa3c9823033
z90d337b1c47b4708907762b7d74d106d177e678463c1770eb76315957d088e330b5f6b942f9064
z119b06290389b1ef9121b59ca2fc63cd08b7a74e067b943f5a0f9f2ad354ec783c2494771dc265
z7892952f927e42256a7dc8fad241ca94d8ea4137d294d7635cd08c7a1570f783da243ec8af8e29
zba29f52f644a7d42203661a04198a1c99cff7d9e91b088c7498f43cd327331868f42fa24e29b31
z0718c5f03d45776daf2bd839335e0c2e4441b722956a6eaca4dc242a9949719aab2d5fa0631f6a
z59d3d077bf853380dc7cd15f365bd9b95e9279c5dcb593ed7ccdaf4637842f0332889d143accb3
ze82319bd0e4ce22251b7174bb8a1627e8b35719b006a3901a8b0262dc07068164a507d1ac27f83
za586f55331d46aba77df291f647530570b603c825c5fb59c2aec1f458c75363a9524244cee1d41
z32ef10f791b5e6c39a374862269e40603468097be6d37e18e4cfd1cfdeb8ca2535b16fb7f11cb8
z0c528bb4d7897ea77534368e9b1bfff0f8abef99970df11f37bf60cfd85bdf77770ee1115dedd6
zc41ce652d7142e40d9b11620cd98d12b73be634078d652d51746800192b11968613148fb1c9d79
z83f80503722e773080f19cfecb515a16c9a6c43e7824d01d3f8a6fef02aeac6276919be7dbdfc4
z82af69c231b6d33427116b752f895ad2c879146bc7d2b28be30ffea267312b5fce042b1432748b
zb6c4be142e4d1289c1e4fffe28c8aace8d8879737c29b5f58df3e457d5b4d1eddfcad02fd69a8a
z825e345cf43d7ae5070d9bd8c48ca04e6c143ea737590d04559184a2766c3182dd4eae0ecdc620
z8f1f73fbe203d4682b93d19ea53bad1c31443c7c693802791c906eb184a5fd38a33a2637184031
z3f486fd2778eb8b24a4a9e48d1ca57fa631d9485402d5b6e79118fb75dd62152398acf183c278d
z9486e849a4f0c18997899a8cd342d226d135c967c593ea7d62e23956d1289bbf04e485a062a592
z54fa95d8d2155650c30707f5bd281feace8146ad05aca88ce6afdba69065f7deb3ed6cb937dfe6
z79f002652bb4328c7d4cc30fe33c82964dcc9fc098bdfa205968ecdbd30c9436574a1c784f8276
zfb8d7fadcfdc1ebccc2540ec0041eb48517d89e43e2ddd40138dad037dbb3719686cf461f99ef6
z5c5b38d8cf9b7cb2024eeac5bf616cec2c7a11b69285195887d6ebe48b2c428831e6ee6d41f845
z40a144ee704ac8590a2ee871f9c27f6d09d00ac6b7d7677a1fd46b09592e2dd10f01df379a9ba5
z4f32c7c6323f0cfccd4deff1a519eacd169389c53f8c9d9a02b4c07321fdd6e7751d515a0be9cb
zf7f5498a54955631d976cffaa0d199e09f3181696d2228f7761f261fc61b51f3ef61236c7f8893
zad463b44dabcbb48d8304dd6298b0ab4954a6191b323585a90cc8bebd2b49429764423d56c5299
z22c9042994210d05ad34f0eafb938a418484e6fef1889b1f67dfc4aad1d40c1dc5ea67541a3038
z9a618b54c0a92b51d6a99029b86826e9c8077c8ced95d0f3c28a0d8658ca62af32adcb0b496c4b
z74b493ccfe2262b7fc8173a7d4edd684d1e01350408611baf9a42eb46edf4ceec33486178ce6b7
z86dd03faf657c3f5ef72f2bb8b38c0765a5f2a00e491652fc540d272c38549467e35d99ab03416
ze449c3a80fde2f70b2e941fcdff20095504d6ae39f99103654847c287e89a6924665e356c10219
z62aecd4f8639871989cb603162f0bb1c75568ba1783ecefd62ac73b7eb2088e45e985717a2f936
z094aeef4793490a46d0236a003baa676cc29a2f0733677110467790a7c1c13bcaf89ee8d9b1d79
za93c95d309d6d63e23f36c01119e9e80c5e94057dcf2fe464297b882e75c17bbe9140c5e13ca2d
za1fd168c8b83d9bceb8e1f418c9c8a1412b10059ab2e82272ad12c3b2916524eb7153206f3e288
z0adb22f394beaeaa56444ceb9ab784ca80a3c2f0d0636cb77c7d6655e6f4d1887bd0e35bd0bc4e
z1e77630d10b0cafbe6c3e3b4e03847da4890da94c75a7c97059f04e6772ec9a1734367b679d8e6
z6252b80f07dd56c6a6703d5dc36a8d207473c800e63bf83a16816abe16b2537e89900329ca7542
z4944da74fce086e5a1bcb1b5c65eb5c5be9c2f37db3791057987a352b99bd5c0f3b5d939e573b5
z2942397dc94d93dc75448837383d51c7d50ed28f33ffcf5d6bf8e13ededbac6227db5210cca01b
z695825adfccb0ae01f8b3d342989e7cc4669ecb116943962dc5ed9b4c69017ef652d7742512beb
z3b569484705867e5efbd8443882c8edc7c962d47f4c45e4740349c526029b89ead6fb4eefb38bc
z512d8756bfc0bf79fa3bc81ff7161ad6793bc489934b098b104859418771219243cb2112ca41f3
z2bba76fd206fb7b72554c4f671b50ed8fc39efec22f94bb565b757a9fdcd3de808c414c35bd58c
z187a7473f4e4fec730f49c5b1277d7e715b9d4362ac32f5750060ae86ed74fc7101e72994ff5b0
zba969e202a04df883e7b854e693640e26563e037ccefaa67e0cfb249c216e361a4887d496ae11b
z542ede7b34aaa1207d09c043a718a1b0c77c91b52d015ced9619194e7e952d1f8f2c4590d77888
zdccb079187dc384354436fcd4b0f5e1356275295534d35053c01ef4123500ee791fa54d0b2416e
z844fcb52bc49e20519f4d5a04dcd39679132ee086887400362b07bf82ce55ee92cb2c099454520
zf985ae9f9a3541e36f604e8e855dafd4edb76ef71ffd4c3349c5b91b17f474c355f579cb4f5c10
z0e39adb9b7e49c544eb207f21040d7fd3f72898d6eb365489e2d1f6f6ab1bd398f8d01b131a5bf
za127d611d0fc8a01104441d921a592f932d6fbb9340a6365d6569535d2b94900f02e757aac00ef
z686f47cb1f7ce1b14fbd0fb46faba9270bca294a9fa91511af1a9d33221793b74361e3a8eba553
z3d54429b0911d838c62c2fd9d63ef7ec3d0f7f4de747dcdab9eb0094834ec460f7db20edf14fef
ze5f6aa2fe7c849b5604d6a335dd0ff992492e3e7613bcfa4ecff43d16c2d0c2ce5e5f8d9c2e004
z6c7ce06d9200e6a30106ceffdb351267b5943dfa8ed0c5ef7a82da4661a36694eda8640a99b526
zca0976572aaa1826b12a1dafba9f489f3369c541cb7aff7399d93a9e8453870050991ad1c5edba
zaf39debf69cfd159ed9d0f6f2e3166db126f32caee67131acf1f86b1a95bb7d13ea9fd6cf1cb0f
z57f446ec504967e28c0a0301067af02bfd8cfd7abbc400b9e6df507253faae67da4033c518c981
zca10ff4eeb3491fd6b993fb1c993d88fc3b0af06d3b8fd257ab99cad422f401e21610ab01f88f9
z73754b043716d98e66a4304e8463985156ef60b2568b3fb11e3561da4fda638518be7312fe330a
zb31d099fb894d24e516c21688e0f80275d4ce6b779c2a6cf1e75a4e9323bc1197349d1605d9f0a
z49998c2f640badbf574c0b8d586904a47e3cad6f936d0610619cf49cc147fa66adbedd21cde590
z43edf0f0b548df864e7ed667148316cfac313e13d059c86b3232360178dfac40b9842f212b6f5c
z1c032b77c5e74ef72a24fe2b895ad8a8dc0369b3216b34183ed9b7d2444da86027fac10ead4ac6
z5781a3e161dfab091d9ad87e4ace8e2d8339f9d4eb1de368db62b36e8736401e4a54d490284b81
z8a33ded512742b91ea7bed6c3982c54a8a6271d27e8a2b919321c5063893ad8a84857663febb1b
zaf434ef9aa7c412d8a0de86249a30a9b475bfdbd9e80ee6a9c0e9d68070cb42ceefc5f534c356f
zda572582754d06c26ad2a0cc0984afe7c996fa2413e5e87ceec8b8c8593e63d8402ff4cb69616e
z9764c408a366e7867e6b0ac9337cbd481e702cd3372fabb4951ae80d646cadad8e162c1f86e3a5
zf87a0c5203979773f54abe710f663a46d70eb1d1bae6e0f038ee4eb866870a481866693b94829f
zaa2fa03939ad804054ce9b08488059557956767d8ee707c955059cdcdc199ac32508fc2288596b
zbbea0ed359fd78f8a9e7826440e73f4703e44e7693907bbb51d3e18a04c964e9e664acdf80ae2f
zd31c65e74bd056aee6cbd944204d0d48ede8ff5ede5863d75b4c29c37c5fa5107a09b26b1b4fe3
ze2348f1674234db647b19d8e7ddeeac173b77ca88e9524b04c02a25097decf69cb4133bd0df217
zbbc83268b158fde3b6a685fee3f54c5e38da88d68b91508380c05fde9ff2c84bb349edd3523737
za7734215cfbf8ed386b25d3f54ef01263c604221d17f35efb5887711e9f7fc06856a010c2d068f
zdc62af4d9037da9e53a1a7006b1670ed7488e704dd4690a7d03285d0d49a7a33f429961b4fe2ab
z530789b5c5d600fc4221ad51b9f2446c864abb2c9571e95b22d19649fb12695a7642572c1933cf
z6d58e1f36f6f3895f64813346581749d78e9b74865f538b7f39fdb5a8ad6559696c9f5a471431b
z68aa61c3ee5b0b735c744b418599f1b8b0e10da3dd93a525d1ba6ed05ea6c3e6d48b57d5285e62
z7f11b4648f6564eb29c2ba12dd105e21372907414a1c870a95c22dece0157db2c4b3506b845a34
zcc1ec18e3ec9c1867fd6c8709e27349a67a56f78276958dccbb5e28993d2724b4ffd1e73300788
zaf278324cad3e25ac77f24512665afa258219e16f6e34dadfe03672c2dbeefb5de0cf34a13aa4e
z52b2eb961f4323a91863104f26e08256d4ace618bbfd341b58caf236c4e7bcad85d38b353f7f00
zdfa1621b8ae3716472bdb045468e059de8b79f1c90e9f2e9c1af97639dacc7e553e5eb7d2bfeba
z152d5f88c70b58ddb204a328b26cfa016bf6eb94e296a5053a66db3043f5033c3f73186e3fcfcd
ze0eb0bbdf151a66535db493c90bf171cf248b378d16b27fa52252b2fe0712b82695e5ec33bd01d
z93564c4594a1ebace7867ccab8a7f9357b54a585bd3d9834841c53911f00d6e59c681f5bad9707
zbd874e15a752da3c025fffc6392e5a61c89a11b898330327b4a2808d15ef1c7f48205d09b4f673
z69b0f4702572282b3a08baeeffc128f737a8df543e043a242d477a999693f9bd0ab371ec7f309e
z519af3b001868b0d111b0de55ce824cc46b669bb6b837d10f7a1c6cea6e47b9e4798b9ea359b3e
zf28424d37ab8b2a3fe60e4f29dc88a2f13cfa0bf0f5981da7f1308b096daf238458bbb63e1aff5
z9f2d5c3385963fb8dc949ed3c5a0e1a6add4b116070aceaeaf773f30d384f67a910cb97f50e0d0
z88653b3ee8c14b887941799a4e4da56d21c0a3a6d30b800bb050a10d2854afee3f302254a7657b
z0b5354c90e44f4cc89321c5f468b920e0735a1f276362c3c3a4892733a6c44b681e76eb392c8e3
z4f9398a08f36a0dfe58004ee176e6ee6cb40be877905ac4440246482a34a1ee76fccc2d05405e3
zc612fc25192dbd7cfcdfde585c07fc66de1edf97bc02673f5e64d27ace93e99186d5b2067129a1
z2d1f966d9736b8d3a46b2acadbfeaa8d41d2ccd4a95df4815e1fb6d128fbc49635fc3d73121343
zad2a14890b1f8844ca2eb357f9d10b2e96ad40fd1697f44c6bf54ba7a95c07be5d6789149acf9d
z9e97cc4e807a0d198e1f3d92bbc6cd634ebfc2f618fef99e99e1463b1544d585174999f151d4d4
z564aaf8fc0b6a3fb4f98fe651d973a90ccad666d46221c238d31b183d7b66b4de27e0795472b33
z7b78fcaa8bc37d82bcaf4509c59fa21d378b3e1e73410bad092b691d02fb0e6cafce095782cc97
z4b56c885877d4c3fa8c15d5839652c742a20ecfd74a922ac93c9cc6d4d43f3bdeb96dcfc799fcf
zd6dbdff9292f4fe5bb12e8fb0ec774ef343ca77df2093e7b6b7adbcdae35dccbffe21cce859ab6
zb98c08f750d44dd628aaa0fb9a5afc1ceb709a987d6da370b111ef3ee4b6b087ed1dd86a5724e4
za0c5c3f105da9cd767a29d72e6db430a37cb5777a864f1df897d14a1953e8e3d8293aace55dad7
zefbb60b6f2112cf27fb750ed05d3f4c620be12766317af47348025eda2ebd85f4acc3bb4fa706e
zfe11a0de1c3bf6d4e512839943020d218cc887442c5908e36bf4daca9c5d323851baeebbd83cd0
z81e344acb37ae9551a82c1752d517fdd072e81b7cf569d0bf3d933095ad25ef4b5b57386754873
z989f713b06bc4444c71bfb90052158ecc2df5c265a7cd8b06dbe6c21672535f59a799f11f8269a
zc8ed83b9ea90b21330afba1249f71216c9c9c70aa65cf049ba384ecc94dc50a57169582443411f
z3a842698a953d87ab8da7b444c8f0686572d7bb0acbfba69fce585cc31ba86e6cd4f39f7666589
zd6f2ba53474205f2bc84ecabf612ca0c3430ebc15895a0ac14a862919aca8096d5005e268e1aeb
zfc2aa127ca506aef2ddd026e14a947454d932ead70560a5ee317e09107917cce46ebe7bc665e35
z547478c3aab25c7264974187bd993aa2772d13eaf106e0f671e84942cb5f66601b17e23d411474
zd61dcac1269fe8301ff89b369f0a77ceba12b019994aa79bedb52c24878c80716751a4cd283d0c
za1d00b1963ebbb07a24527ef4b3aef402c3c9bf67f9d6ebc04bcf33fdb3e99a915d4fbb05d2511
zc6366871c5a72e60bd30cfdaaa8dd738b636b1b6865601c9db7d23e560043eb4450c32442d322f
z0707239a44bacf8af30044d2f099e28aa856e1a9668ffdc23f4963b86ec91db943e127259e2b56
z9dbb8fb7d6f813176fa308d558dfa7062da5992e2a3808ed0d0469ae02dc98f7a2eee18efd1b91
ze177dc79ec423297ccd43f46f338a4c7bf356529a9e4eef3a513168d82685ff1bc8f08c03a9a31
z3600784d3ffee311eb4f28167688f9fbc2df63be5fa0ec5a58ddcc297ef28358279971f783d21d
z264c8c355d4095f83db777de3053f01eb6fe150fe8543084b2e10e8bd25a5f8be4ee3b521a4ab2
z6d14c509e95e38daeadf12c9be7f6bde13befa702800119ea706ab5a81e88c131b2af2141634e7
z536bef103a848b0d5903bdc841ceefe48f761ef8156e51f773f3624ca09119e98a310714c98f88
z6113eb2dca017ff19bb0ce6ff5d2a6ac572b97cba50b3175cbeb0ff8eaa7db7d508bce3bffa202
z7730400322172872396840b40c06301ec7cf222bcafcf10d29ee39ae5897654e9675c61cec4db4
z49e156a0e02fe1e1d7336b704c5a554478141860105aa4ed4ac3a0aa8a813e8f17076c0db705d6
zffebea81a06a1e1210cf348f995ba3e7abff6cfa72b8b86ee7116d926ed1aaa33042e5105fab54
z69bc7f2bba4d0dd28de818e5b109504687681fe1c0ddf123c25992e905783d038789e8de177db5
z190b77f53ffffd449d5c357811672bae17666565b477b6c458860ae5fe326be7a6168824a0dbfb
z932a6447309c9510f68d97be1308a7556c55b49b982314709d1e42d48b0d173e310e818829fe5b
zd6cea7d7fe9c549f61016c5b4beb8aea949ae87c6a3629849e91c936fdc43e3735c89700e11a50
z38e18f7852efa5561a580e0c460e0aa6986a5e3524d31b4864782492238c5e31b4bc3de89b616f
z06d2a309036c571bb658b82432e8acf342b721e10c3a9d25a6bc51c7504d575962e849ca3181e5
zb4ecc3184f0b526220ae1eafae5a3dff883229386089c155257ec4f2694dd4989eaa83b12f130d
zbc14a641d309185a3f9b49b1f67d86aaa529a866b0eb2752100d22a61a65fc90e537eeafbc27a0
z801ed34d787591f4337c791ac3fe88b82f27671d3dde986678a076df256fb6853872d12421d614
z5e06ed0ffe9c836a229425a7a23e2e3fe09afda886bbc8e95bfc9ddef7e07e50497a9558fc29f5
z52d83159769e4d2f64dbc39f469d45be2a75db1f40099ffd5db372129e0d806ebd117784577d75
z8177da8201388b714b0097fbc63b3bd2dacf694c03dbafedaa539d0df6995ff72a30692ef545e1
z73f6bc48d781f3dcec17f9cef1b8de4b8e122857e28ff0c234361431c4355ebaf87be2c94f2b7e
zb8252cb631d292144d772c27190ac5558d2b7ddaa616548142331063164551c9e8d9604e7cb5ea
z950cd3709a8b5d2e6ff854d8d8edf35489737bd0fa7bd519b32c9b29e2cb9515e6f1ac7c84a314
z5059fd261607f6d54ae176ac7a1004cf14ce914cc02c2cd407961407944afbe54d4f756adc7c96
zcbe98e533c8530e0c62c6a3b9c4be3e1a8a640f252f411f94e03fee95aeaeb78cc6b2e02bef864
z252403294f097d8abcbf7ee9153d9c7869768e68c99eea271fd34562b8bee97ea60d79636b951e
za5cdbee66c3020c7a3837ce4266f2980dc66bece2f73089d82dd3fa308d643bd381697b6257ea4
z19f94c1bfd55075ece3e5bd03197b3c6f251d545a656b2c3ae1dc3a838be54b5632bf6f2dc6e1d
zee1039e8ee65ccdb8055d7758ea1846ecbdd18e5d49b2d288a22db189e618fed80f284adc14f3a
za31f07bb07194133fc216f4574402aaa772b39fbca0885a9fce54350fe3709af57e47d36f0e7cf
z97b50654f04e68b884bd3dd58fe38d76fe0d7185902fc6f2945262bd322a00538debbdfa89a3f9
z95db67f26c4be79d47d6b63cecba6556c863cbe0e3d83804901db67f7bfc573afff7cba1be4028
zf5a5767090eceeb1762b874fdf1f36ec93a74d1c201afa18ea7d4a9b12e30bc0ea97f02f9656d4
zc5268f08b414528a939970a27b02fdce0f238cd1d7d80ac2ff3b80e2f1df6315326024c5916ba3
z0ee24c08149e7b5156c2a08d0fefec111a924c65c4fb974c4b6531e9311f6da208445662ecb740
zc635f0c18a6508429914111919f509fc72c4479ea5308561e9c913608e1105c5f7c2b5995280ef
z5904b4f631e53c9a294c50d07fa35918378d5fee1b47f5578c51b5f3c8f49bc3d98e8c77d63c50
z8806d416b8383a10f5c6f874df47ceb97ed4dfc338e1dd1beab56f6e4440b7161858f4022e91f1
zc687c9ee46d54a273f4d5e899d56dacf12eb403b0880dc53b88de3a3cce26ed9aeaa67e09e1f00
za371646354ad3627e66cba1d7d25cc42d00c21b04f2a81a4699927bb84c28d4d0ab6b4b6fc4e9a
zc6207fd8200e92894667063de475051850077c1d19b05ce797abce51c56ee3f1577aed9d38b995
ze8ec29ba84df0a000c9b5526109fb58d50b91dff1c2d74b98f04514a4c7d5f8db0e13e3ebec7e1
z55b064982a6450a62ce1dbac9659c72386b00bed515997726182e162527f1ee511e3fd188d6183
z709974a4a35754ef46e1ff86aa096af03b0648662bb32ae44d6083ebd2a21a7aea44be29e26908
z78cc13b78966ee71b519d1119a8baa62eaf7a9fa4bcd7e8aed0c2a1aba511566cd25854f8e3404
zc2066069c1ba7e4552cd5484c5ae4d2c1f5a64da094eb79b93f121c6a8d84d0f8a696de8d80944
z0b2bbc2a8601d60c11e4d3512f2ede4e16edf0995bf1d0778aa0795cf3ca6f1bbc57f4bfcc56e9
zfeb813e3379f68e93ab776fb999efc369be717ba0b36fabca9d9724b822dd5f0da545034f58f4f
z0bca7dbfb26d62dddd5ab0d1cfe73e47a0e0c173fdff5e0aae33c52808e7b75ec9290ee19bae87
z96c269d8c8be913717994602769c51882f0c201357008d917c211fea913459982ffe2c43b683c1
z743f1f3ec9f2cbf6a735ff4f550bfcd6e1c827cd22949ebb40b26670b234f1b02a396cfd48d4ce
z7f381ebbca102d8aeea221a9779bcb0ab997a95478e006a2fece768c7853ac08f118b206ed93f9
zf6e671cec65f28f383897d43a285efb72644368d77b394dec5d4849854090c2187db603d83a130
z599f5e67b854e48012e73f576c6691d9e8e5c0bb75a1cc1d35a8ccc94af44d9dfa7e11a0df99d7
z6e3159b9251f225f50f1e49762548068678ed3da4e506b49901d7420f10c0be5e7c5e70bf2e5b6
z807ea17e204093ec7308d3d9b3bace623305d263882656946de3e5304ee0e99f33bba3dd0ee6ac
z733a1ffb46286565150e44bd9d20f15be1b7f6e5db4eff1498f93132b3343ee61f6a1a3ed49d72
z7539eba4b165bb30916f59507366a6f86a01f2ac730d7a811a03226d2ff0f8b1d23c3b1300fdc3
zc8549e2c81e8b6505b42b15f057df117194f56916acce6b15feafe0eae174ea56cf6e85481dbb2
z4f8e95b3efa35442f0d5e4922ace42f274b050813243961e7860060073093c253c34cb99e106f2
z19f4f3e73ed5b103682772f9759943509c1fc7ebe0926340c32d0f4521bf4d94847acfd18a23d9
z67e78e3b46ff9afbe87b4c9dd69105f9f7c1b8bf802217c5e3d99213cb609a33012aaf5f075d33
z8fd63998564dcbe0c05ecceece704406a1c6733d38623672b014aa8429488654e958c9e07de4b6
z539195d132dde94424f31b5ef43af0f634fbf146bd47c5dd87cb87b1594227f47a6d6dabc270a6
zf0f66d478c4cc6ce31365a6ece83db123fb878ed1ace236332d5c61d6db2f53a972b3ef97653ab
z1c26b13f64375b960780a151f604d33c5f0b1f1f284daebd4e47a1b3fca5ac6b883e4f2c12da5a
z55628e249fab07dae552256515737854cb63b942fb42da2d75d223f93bb56eccd9e0cb1756904a
z90f874d7c940fafaff16266ea909a71b99e9dae8499ffed5b95e08a431d60a8761370113153486
z8a7e27a2ef1366f12665620166a060f88d701cd3c0cc550315c850eab80ac1569244f4b9a71f90
zd833f82a15c5037ce4146c7fceee704fb589bc7461c6fc716f578711b2f2f51e7833fc333a03d7
zb471e45d5ea2f1b6f5a73639a96d15ba1012c36d1ef38eabe6ab2223171c8ca206359dabc0fc1b
zb31922ec43a7a74a72ca4cbc1ed8aded398fba9b5d8487bafae7b0bfd27b091fe04013487981da
zb3da7e2d4e4403d97c17c072ff33f80de781a68eb61dcb7bf1568a4fc1ffcdc2a38471e23c1b4e
z27c7619abe3c1b37e1ec86441200e506a86f8b6f5a32e5aadbdf7bdcbcc7e8f6fbd2da1df8416f
z380c8576d46420aac8b4e4ff919e526538df741dbe6ad1ef49ff26fa8042f2e855581bb3b9544c
z7551758cac4e1e73ef09ab114cf6b31739fc0ba5f9157f44b81b21086ebc8368d4d6c633664fa7
zcd9f051ceff02aa54b95715c3f0a83717d05a3608200cb83482597353190eb7cfe6c692d8fa90b
z189ccb79fc2fbf26bd8857c334a47989adad91bcc42df936c2b84b2fa4b0d16672306088cb4c9c
z83b5206528fb0d59fc646db35a64fc627b8024844523399dbf510ad3dc934c967cd3f98599cff3
zdce651de41e0377394966f3eb26ed137ac9f4df1c0229004130919e0d7be630b7344a7e1c10e31
zb08bf11ae898a17c58ab2fe41dc65cab0b73a0d01468ef26775303709907d562f2cb474654ee01
zcfb5af8dac2d0197f73d9f2a257f2df73ad87cc6ea197e9de79d0f4c5b2ab4c2d4b8cd132a6c0d
z072c2b037e43cff30fd0636fdfd80aeb0b3c3dadd57d995898a5be43e4b2c74df89adf6eb978da
z686ddc34eb9958a70b6566102295f30da1d4f5a2bd43623addc47244fac09ac7a6800349f39636
z63cd5803b2767b2dc49c5be84d6cf5505254bfa72bfbaff1d2a32b2aac253fe6ff15ccf88f8f2d
z36ecdc04d4892db58aae2094c048304c9c6c57ee224d3cce624e01393244d96a9e2d1e908ef9f4
z74b528672cb5113b6e3e772f8bf5d3271d36b3924a5e3bbf7509fa41347c0cab9b1668d2770193
zbd078b0f67bfc1caa4d2b2e2f3cb24c35b8bc7490e9f2e2a506d286190d01d1184ae0682b74201
zd4147a54f1762b2369be81ca95e7e003b9c852b7f18560ab7ce49ed106fffc8535779762a7cee7
z1731906de06e134f9b8e9edb37637251f56dba070715c3de5f2a1db8642e6b7808899c56105441
zab6c550913023471c49b52e774cf6679fabeacd386a70d7366300eef9f548998f59c87f4440149
z6adcba2d1504ec00e1c1835dfe37ab1ccec9631df10d58edb4e8b253604cf17e816c184bfe07a4
z041e9d3caa32dd45665b5ace8645b6bd83bde001cc02087997f6a0e59cdbc64613592e40a4cc66
zdc73b40fd2964b5c1d28171f916ac2cf808e00500abf29547a7d113502f268dc5ae4627e8d0886
z0281a475dfcf198f49d096570971718e227175be6532f572efecc9f9b64f1831cf7f4de6cdcc4e
z8dbdc38789ccf03b3b847b220d5ac864cc159ace7e311e5838b77a7ad154badf34c9ed97ddbcf8
za0ab34d73381e87bc00edd36260bd39fae3b441b325edbe0a51329b21b1c7527b950639ad87d41
z1529c780999ceb1a2b14965f0b9e093b16d350336aa1f96579e4fc8d6a5a3b2aa2eb57594c3b19
z7e1bc511fcde9a9c22edb1f91d6137f91674c5fd6947780f71b8b1e9d1213f24dc0bcd08d0c075
z39e2df42583cdc4c5086882ef7c5ed9f5ee83f821f838dcf76da720603915a7169308724c4c551
zbaafc4362faa9f9d5f4a4eb4936798c67c4857c8c76c555fefa50cbe30d078954ac67891383fc3
zae065acc427af48e9c4e2ec2a20cdc5ed05023ea00b7c777c2bf6b1c5c49b7b5adf77fb0cf9b68
zc47d6d3008c36ba8a904f974a746a9ac1060681d08434d3a9e95aec7bc0aa089e46c68c3cf4a20
z754be49fbb9311b88955fde07acf797e6daa2dd774ef637b8bf541328ac16b45dc7f897a88d4f9
z0e3237ba8a1b265ba16040c44ce8358b8dd0d2e48fca6bdc8e704e1297a41ccd1d8c2ce9e5384b
z7dda5ef157b9569393fc1ee2e774030ad25602fd72638be9d05793d2e318463be9c9f7ef811598
zc39a255d1994ec9022fa7be4e6e6785497ec9687f30025e01ecae02292bd1921d2c7d1ceaead86
z9cd6b681f19935ea81877df216e0ae253c36d6efe0ef211ba06de7332831569892d154dc16f7c2
ze8ff8eb1ea235afafb508bedca9a1e6eb606eea68a8a915751e1517ddb0e8cc0b3593b0f8ecfd6
z24b2b71d01a11454d406ea471adfdd72606c1739b1d5552dc05eeac08e0fd352867033b8cad88e
z9959e2aeb6882e7263d0939ee2f80d1ab1eb55797c541943f886e93003cc98abebe35788287402
zdc96f12dc839bfd426c3a3dee66d9e74cca86a2838faafc35c44fbadb2db9a1d42fa551cdadfd1
z1c4375dfd53cc83f1af28ddada223dc926645bb109e6e873c8e7a28395fcfd1e05e5960da8a1d6
z40884d19f8250d7a27921f99b46197d99347e71dd2e8ec33f283b0a1f45cf141df342120d62940
z296abd5728fba13d5fe908bac55d4c6187576ea12f1c3fbd71392240cb9144d28fd6b901da145f
z3039c036c707da2377bcb93d66f7f5d898b1ae91c56a8003251ec8e24fe22d02745ed0f89f4853
z0d2362a097a9648214cc03bfa0c43bd9fe9f6513f6030be9fdb474f223d413ce2285114a31afc6
zd7dbbd112ae02534ae8ad3155157e50229f1c20a1fe1a3bf046054c046cf440cb7c49a9763e2e2
z428ff9750298223d5535d0d44c698aae10a9bef8babc3e00e492ad3ef70d0d230db234819dd74e
ze4d8994cd9fcb0f4526d7d22f8ee54a47d7f5533b1b4e51194181207210afa1b6169f05802e66f
z48612fe9a4f40b1db6f1e9db021025b8c5c5867987fec68bbab8a3a82475c1143963938d23c270
z3c6f6612aef7a6ff1b16b01233764f25d82f503423a66e4e631ecff8307eb7dcde6265e7d79fc6
z36748dc4196c303a06b524a8b4330fdda282aaa46cc5dd748a6f552199c9957d1c3a5ddff3166f
z28ef7bd0562a99c57ed48da6f3dff3af356e35014c2729571224aa4e0a91fb69f3327308b2369b
zf277fc39657427fedbbec01cd8708494bc5ab1c6a9455b170dc7451589878e00de07593284bf9a
zdfd8b0e3d40a118047c53361abb15c3d2e1df78d2616324d370fdb8515231865241ebe84f5318a
z83a2c629a8810f2f2824fa98415b2d9773281c4620ee6d87ccb48cfef09b5be615a2080a8ba084
z6b75e679c71bda0b4b131c2c6f2af5ba670796a5f14784eec7dacd3ceab8d3cd463ac4b1bb3db2
z9e0d85c1e98b4652e1c277f2dbfcbd870fc0adaeeabb2c4a5875f161b875c6c44c36e37b21ab69
z7ff5097d8349ec3bd8e862536e41ef3924c50e1e195b251ba42e5d86053a1930df1ccacaa38672
zabbc7ba9240ab47d2fc3500157bd144026a00301bf7905d9b646dd063c06cbdddf573cde727a14
z3bc001722af7c913670b367b58c3c764d852c7c2afa819209afb09b66b1987b95d6c8c1331ea4a
zcb114f92d7ac4aebe7a09dad740b14e20c9aff122d305d12e829a194e51a833e45d7a589b35cfa
zcfe31b0ae5048b2cebbc33b167dffe51afdcacae820aa999eceab93055bed90d2dcfb19551eaa4
z8ae35c23b3adb3b59a1587edacb351e428e4fd674bec8c8553a930086efe5b2ddca21de837fdd8
z0fa265697dfa57bf34ac3bae3c712bfe9e644644cffb89b1935abc56a99cd31e40eb8f309e1643
z8785d7b90ae3df5b064cefe5e694ffa664870636735281db81c9cd3df94039a6285dd2d7ab0479
zb59dbff8fe6b6bb7dbaf63eb7a97427623060a42107698da4dd9571d542b8743f49a3c9d49eb6f
zbde547c1447fd815b0f29eedbf0b08087cea2e55aba42c062872b1c74a2e9a693b2f025701d0e3
z45b4ec522876c78159a6b9a2624a246a817203faa1e2f931b193d2b7f8b580ae63181c11a083f2
ze4d6d41b2d3fa1e6f3cb8b9cd15d7b9313197240a3e4eac4da5094f709106d7095ff96291a6f9e
z47f3d8d03f7aa1e47c266af9f8389815aad1ed54103faf0d7893ee4229b8e69dda4be55c5f2d9c
z827daa522bf964b41f0eeb735f52e8c0b62efdf65badf52e1bfbeaeaadd96e74f2fd20a10bd6b8
zaf57a2571254c0e0ef86fee9de097a939fffeab4ac3662f237fa7d1a400be538dee15c791438b8
z7ecd7d63b7fc7fb207e1c7f3e885d46674e781372ab01035dca7b917806bb5182c7b8180982f2f
z4d19790f2ad1b7b2005f1c8670db7caf8dc6188709754d3f4b76e42bea87e6a7aae55419c1fc8d
z9243ef6acecf49b622c3beb8619c92b4282556f805c27f933c064a441b7cdabcdb7f26abd5a516
zccb0282d988f63e46fa88d02581bb123276d9f96d12d4b75468eca602fba39f53d30428b7445c4
z3016a159bdaa203abccdfcf9276c06df318f746361f5c9159975191956c2dfb51765f9fc1a0fed
z8ffdbce25160a359c27be32685669cf4d25c8d954a0fadf4bf1e3a81a7fe28c8200adedfe3ed68
z219616aff44389e556b563e52ed918314939fe0284d4215381b0c0a03500c96c9a1eca3a743c4f
zdfec4b48de5264bb228b58a9df64313811c0b72c8cb7c76c2d79ca3b5b8123a1934861eefd5a24
z61c3c97ab161eefdfa09bc5a8c3bb800237a61690d7686f8031aebc106f483c881abcde33ebfd0
ze7626159fc92f9e9915c2243ac8a91aa10e781d3efc5d01b00d12817a547ff3dfc3a151d23b46f
zb7e996fbe56f408a20692de15a98f1021020523a0d17d9fa710d5a0d5abb80a43088bb7d21f03e
z205f797c61e722b75c9c5e2b98bb5bbef43e2e54e81e432c9b345e702f5604db7d15a862e7ee15
za4300af633914dee72a8f3e99c8cc24e6e7c7bec81f62d9be084931b6c27ba46a63950a9bdbf22
z0214ccaf6f23e7739cfce94ce85628d0719d89f1a143c6e750d4528e078078d037368f4dbf5b46
z583407d52c2c13716fa81b7ea472beb51c0a002778db0c49cff10b8dab5a798db53005b809dfaf
z5680cbe589628f18765163ceeefee701d1fd03a92e6f41a8df72b01e25df7210d6a40aff868a5d
z155690e2fe8b8d44716a68e83ef4a7030635aa0d39dd21acb4b1b6f805c3adc1b7b49c9d1091e9
z17b41f5b3bd620ed461c5010010f4b28fb5c9cad9ab5e82998d1b417ea8f7c9325d23272652682
z4810fc4d5f90e23df506a1e0f237803a92734a679f46fc25cd5de1faabfc3315be7ac5a3779190
z2a4d0511d8f9a1aabf5b163a321c04746cdd666a9c5472e9fd828d1e02f476785182e81d5cbd53
za53e8eb67c3ae478d1e4f67742e65638c5ec6f892b55f602244dc795c7fad3439b98a6b9153029
zf2631fd052d54925120ad5133643b763a92ccc463381e1c31b4fd0b22f09114ea6c500f2414abf
z79f926d42b928008f485c41794dfffac7c2c6a651fc0b1ac8dd886b27f1114fb63790b7553a833
z32607d66222c0285bed23b28aaac7967370a0237410d38785c5f7be42d9beda22b23ef954895d5
z637e8346c97fbe4e700517f3d1b9b9a06d9ae9aeecdc590f1b5bf2af3bb8950a07541ef72476a0
z97658bd1dd5cc5e28351ba4699d09b311240df1dbde4973a37dc07c694a93c0767f5df56414674
zc64273ead87bda85ee28b2168081d6f96f31cab4ea753d8b2e8e4526490745ca876c0698484d96
zcc30daa80a688783a48297787daf583a7ed2d30a13ddf24cf99763dc25d08d000a8acba2c2d1c9
zfb42a058a6b72f2cdd127342d9c44533732528f2baf661f9ff04de74f014ebcac55c2cba12092b
zaa25a41566543fe0d4bb803ab7dd0cb738c63a9ad008654ec8412a84f98d5e041cbdee9c6ee076
z93f4b9fcf2af3b136c6f0f00111896760bfba6b876b0a289c6f4445f69eb0e171e500c05e55d54
za13e6e3efd23c3b66ac099bf3d6e4398b143520524636515b048767c37c0ce35749f977dd06a39
z4ee2a6786153ca6d5ff694c5a29d3bb2aeab1ebf039843cd8ed2e5d7f09abb9e03d4b95c21cab5
zeaa025dcb12d80fff6b4a7ad5f4a2c5a49b9ff6d35ac60c69f4858fe86693ff1fbeb450ba8c4e4
z6e3a4dbe6bba5298d857deafe026132d0673d66ac5343df12da3b36d58fc4856ba6ac96bf644f0
ze8c40baeb740511a85e0154ca4b90485de6f8a11cddee67340ad9ca71aedc28327fdcb3d0bd651
z2228f2d9337ddb627a7e36f7d7130e0f97f5a86b62b731100cfbb37753d77ad48ed7c74607c1fe
z99fa73c215d5c9879608964629d018436f276b7eeaaa5a6f1fb77675a122afe09014eb1e442dcc
z95e09102a0bfcf93bf5ba4de1820f0d2f3278bc43724573ff815c86911a0a9ffc48a119417e8fe
z96a8ff6296481470df4a2f3a5bc992beb87fa0090cfba0c13a2b0aa878f344fc5ced158ece2fd1
z7cbc523bd2c5e22e7be91a6bd4dcf886c65a4de7cce92b5a52d50db39ce6eaa00b198bce1713be
zd131f5b61c4a8e744977b7772879d36f0cd1cf8ccc3ed08d25d43e7afa1b012265488d01e90dfa
zc4967c3ecffe7d7d8d0a592a89ab54a7db591a11a043e9672fb3e3ac6a4a4778f10a9e79d55da3
z3b2a7dc98138fa146b725b5da192661ef0f0ba886ce4abd3c1a97a447ca2a2101ca5449d0f8acb
zfa1621bbcb3909b686f4b0840b4b25ebe10946081d19b938a3c92aebab5335818e2d220ef5e30a
z06993784779735f13e4ee4e20c4d469beacd5940628f5aaa5648aa94e71c1f17b07a7d4c4b5f50
zb922f3be20e15098fa1f6e7baa0d42e4d835f522337fbbe7271817dc9621ebc01e3c7c25f87790
zdc4ef0f0e62affdc3b4f89cf1bd8f6d6c69151735366455d5038da15e0b3de005b11d22c7bf000
z6de84cf5aef395a0c5fa9c64f7e40ba9ac8b3c6a7adc509219b50a119bcd7504701386862fead8
zac8bd50adac54089b842ea38169d5f0a207e8473230e6190f984bdd91956e302ef029b0647ba71
z28e7f82cb6f741599dc8b80494720fdc35f5ca6abf2f838647c294460aad0de06ca59b126f26f5
z5e45bb7a9eb59fbc467a0f084c0655dfb7da62baeaeda57fd3fd0271e409dc3f01070dfd17da31
z5f607dd6f4a9d7a93bacaf9732a9e713a046ef2293f45ff27c5f506e61143e1c3b1808c54544bb
zd523d6202ad9638243539b57749b5d79cd9ae0b8fd127a500675eee777f7fb52ce17759125768e
z7f405547491ec65c8b105ac428659c0c5353643f106931ef9faa5a79af19626a9d181365fa4b56
z415fdfa778d605d9fd7e9fea362a641423554f9d5aaa6a1bf8a68e7d4b35358b4baf08efb7acea
z70aebb3cc2bbca03388d6c06714af2ace48c1fa6357b042054149e94875249bed1bf7f4ce646cf
z904960f4ed13b79da5345178df2a559e4cf7b4a78d41036d9cf966c2b70edd2a37446a74626aa0
ze4cfef1c314df6e0d038c994c33ca9fa2aee01820a1ec9d93c8aacaceb22c01c3a921e79562594
zc5eb4425cfb0bb7fdc5cfc65db7c3012d582f5784a86c25f140f9bbc8e4a5b36d9f95c1ae7b5ba
z4087ffa76b3f24b7ca367b70a293c4991444d5ce62b7329cfddd7d1c4051425ceaeca28e555c64
z366988e966de020e028cfb686e5fe969149d7b62057882a389e611f81cae3438c4315d00e5c763
zb5760c933c1eaf5a63177fcc42c1a02e24894a9c8ecef44d2ef26da903d87d8af40e438a106762
zd6a5ad902e820cdacb37dcf06c1087502e99ac88a5231f3808713ff5ab4cd0a3aa2b92d3e72fde
z1f014cf6e948090fe548643ed954e8b7f28b665add227c6177951678a7c009326b51341b88507b
z345b4719ebedaccae4d02b23ffb4fe285ab4edcddc6e444bc352f79f8a374ea4a7ddd9827ba8a7
za8f3ff813090f60f6beda8ce4a4526fe308a2bcca82eab1de747a502fcff5fa50701802cd360dd
z8d2613d7657ac8177bef6d577f7bc8102212e1b35053e9710f1b0555a2950545fdcbd16a4d74d2
z9331bb3831af5683f62b3c28d3ee73647d5978af5a4f76c744bf0f43def725eb09c361ccc24f06
zbda1b8e73d4a6a73ec218e1d21589fb200d0a779931e79dc694c0c06d4cf755871a01f9afa98a9
z99b6b0b04521edcf1b18372c2e2d13485ec646510e210d46afa2ebbb16b0d0fe90aab0411e7712
z026fae6186513ae42cfe9b770c6cd27521068d42b25b7b8e518b1bcbd1f3bbdcf1ad7a32edfefb
z1a11048e83b451c9254d30d317532e76ac25058625af37bddadb6149fa026cf7868b8fb1e1046b
z9e6201b2b7bd6804f1535df89a982c5fdd5339e6ab64ef7b025b770ee143c5eefa28b3b291eb25
zac16aa9edee3f9f6b1fdb4e0ff69a456cb9911250f30e78a6d13eb6c2a9f67d8a93480cc55d8b1
z6fb56ff26113b9ace7bf0bcc67ca979670a977f233a4a5f3682bd373e779fa9cc3a70ed10410f5
z359dd38194ecc044ed18b69e4c2a6497917acd35493b7c9a0aa2bf13be05a15af3cc00dbd2d0d4
z07a15a58fd4c43ee900b8d1a53f7c74279ffb631ffd3a28feb219d1b39b1e6d22fd2a5ea5003b6
zaa7955d1570face26f71293111c4485c03723f3264baf147233a3d3dbf751cc52a080894cf66e0
zc6da94d9fe8b6cbc6d6bff604064278890f71bfdfd5bbdcbf5dbb6089d83b33129f4e5f2033bb5
z93116bc12e6ba8e7bfa4b0329cf6be963ba591baa5d4927314d730b9bd189bcbf6c6531ee6478a
z20defb79aa94c6b5c7bd1a272054c4793539cfcc9b0111aa1b159e0c32f98fa97e3293bbb3b13a
ze1a9ccc380391aed1d3619242cbb286cd2d78befc1aa61850f664595b5785be18668e8fd52c5c4
z12111f3996b17eb6a3fca410a2a746c78ce9c4da59cbfd53105e7802554be248569b93b02b91e3
zd3f14b0574590ee9fd3f45108c3d059b6c148b61e806a35fb00aaf5c5bfa6a9e597e7f6c8bf499
z1ea10a6dbea1945b834eee8220d369a2976951e54a53cd01108e0ae95e7f44fb1bc04eb0db7d05
zaa24ce11b6d87dd678fce9e99d6093083988adb05da66bb1c67c8b83eb900e227c6c335f7e4ace
z4ede995c02236fea976c7237b00ca35d67d7e2cd60fc00693104fdc4f6531b170fa1e1d7ec08fe
z12eddb6d6db527438e5baef41f09d85a8c7c04ace79015664b02189f457b8b8522f9a29093201c
z156ee74d22d626274df3d590d828b72afce985671abb211245bac9fb68a68366da4ebad863f4d8
zd5fe0113055c74db0f8fd4c4de0a7ce99ffbcdffdab6501f0c241a9f7c3a2f3ccb7cb79f1f39d1
zbce2c100e719c469ff26729351d7bf3a0be070c7cc0dbf21816eed6cf12a645056a87007aa8d89
z37732e05589d7ffaed13b9286e5a4e30cc23fb5e588fa014254725f6a10b931d7fea6bdff9232f
z66d2792f519366fd8db067ef60c8897926e347d45d155b9cf5af9787ded160441e2bc987d22a20
zc53f64b4f7c5fdbf3f4f85d32987194021270d2106a9b5e9a60ca19b27ef49d8647579da9bb2e8
z54a74f3fed8b7e89e9d00a790934a31dfeb2f41916898b20f884bd5f6926ebf9479f157d16d69b
z61bb7fcb031e499051e5c7b3a0b26334ca6800e8c9eef94994ce42de774d2da65ab684f26ccacf
z3126ec306bc73774b131d571d9ef22fe7494603d8d0d539141bf1337d4657d26a938a50b1d6076
z9175a2ac49bb45cd36b299aacb503bb8af052843d09a58dcc74df84d9473506ffa08d365ebefc4
z81918563e7c74d41c8401b38979869fec957547d78dd254b1437393026cefa4bd17a747b68df58
z70a6c57715ce2fddc09f2147cb840fcee58bfbbc592d9ea183c68ac212289a86334e76cba49bfa
z3934b166f27b61fdfbacce7fb34d49bc75bf93572280a71180a61e54931db5bd331a5d9d8e5b03
z126cf42e465aafcde5dc0d7d69906e64514a9bb278761d6420f9c0ac2dd1e2fde8dc457cb4b78c
zc1fc4ee7a25cad978d3473c949d08add24b76be5d37b66edbf8b12694f86ae8f80119a875179db
z2236a8f5294500cf068e12037774752577532fd12a89aec8bd90a0b163efa09a18fbb1bbc31610
z3760ffdc6c896b69656e4b82d51b0ae26b99098deabb9b8bf27b9d2789ca9522cb6cbf5c9326f0
z9353c10f724eedcec27a7f83564637a3aefbee38f50ddab2d4e1ca53181d4de5deeb735fbe794f
z216ff72c06e32f69d1eca26d03c03b3844f1632afc8397e0da012b11adf857d012492987609d99
z351ecd2c4e4e29045951b954dfd1ca58a1d3700f3061a117014fc05a72a600eb739721d76c863d
zd1c6af84f4540a902e5767fbc1d690162ceb36bc9e1dd6aac2f1c5b02af69e4c56aac7fd329736
z8d03712ff67776b6bd35bdd3520b10fa50108f390abc392c216e183849c50a8ea10b16fa5e891e
zf4b9261b47f8a9214344e12f792268cbd3578546dc4d5f687ec6f922acc2f348cfb3bdbd4c0ab1
zddbd08f5c6645b532cb6c5b4ec6a4de0d30d67def017463abd9b3bd82bae1b3c6831f51bbada0e
z90143f35b980ac0c18fe4c21b66cd8e7e3f888321ab0c3944381a4f3ee32118f0bb569104598a0
z9075f25e287e06b49060a9674594642cc57a8a751e7c66779898ad82ded5165824c72926ff01ac
zd75d388b8514b93e9db97c0466510fe0447392720b2be7bbdeaa9c2fbc9cda0560bc38eeaea49f
zda8af50b7484dfef1d56f7ca78796c9d46c088cd9834c29be231c62a540f465efb17d28ded67cc
zfcdcb09ace050b6153c61222612b0cfe56bfe060ccf2127e35f5d02e4427938b6dfae18558c5bc
zc1d467ea13838ba0aca6fb5319c7cf524ffe59be0ac8ba3692e47cf6b4e0f167f70b35d835f3b8
zbda599f2ef57a1f209614cf1e81c2f5d14a1de62b65171068f2529332c833a781dd32ee8f7d601
z14511834351f5e578e6595757ef6c607e85b0400a6d832ff5d7489cb06efd9797b0c513c2de748
z932dfec80fef109b1eb0a30ace5bcb430c2f585b06d97680d9789da16b6bbda188d071a3886dc7
z6c06a3bb397d4145b28f6f5810fc3b3a9e56620d6955f6ea32cdba62574dfb9817240864687e46
z863a1a4a01253e8481a502139a2771e3b4bb6584933d28acb4ebcac227583b6875f9b5c4952a2d
z81499245604e5d1b9881bb8de1025a048bfaa68002786ec0e7a33e33f260cfaf5646b41ef3efc7
z5aa40774a38de4700730abf33f77072ccc17e6da935f9e33e25346f5b441e51aed6ed6c3c9dd1d
z61d60d35a1384aab71d100d402efafb2ca03a9d4662ebf1c21f6be5c8c4cd0c4de58089c0664f1
z44c573df7f020318c01dda64d44859e129a37871ccdff897d4b9615fbb4d06d835b85504979bb2
z2ead6f87b175cac47d74c08001503ccd1f183da76d4eb59cfa2a8fe5aecc29cd3f48a905269008
z1a9ce2a2d9654ffe7dd9826051dc0734a9fd7e5617f823104640417a9e520e037b8941424e0398
za40744343fe9e6971e8d28f28e0d3361f8d9ce63b5b068673aed2649afa076fd82ab88a0929bab
zcb4e926f8c4138f9becb2a4c6a1eea288717e0f0351490172eb38a39343bd2fb3d63607f8750de
z0f78e195921d0c4818f73bdce9b5e79f6ee7a527b5e4b6920dbde2dcb5ff430e74eec65f04d41d
z4636b1ca024b1643b79e4886ab3a9525b3b65f7a7384f3aeddd47b3b200e5727c93414e4cfbe3a
z47105de133c09fbe668611f2b383c6b339c52ae66feca98e7944105ca69570580f0735f64c89d9
zff39cf34adc5004b8cb2d6faf0b3772577672ee94fe41143da9c8ef7671eec49586d4efe69a743
za1032700ba5a4ba4fa59238753512db7c5b8222213e3e4c1b191d2e6c6b2e53d6f6b2e890149aa
z376f244c4afafeeeeb0ad7627f47b280926091fce1aae03a51ebd04c0661597376c4e7d8aacaeb
z2983fb6b6f3e3632ccc70e6843f421c094311cea3df9a6a2fc07ff06c1ed156bb559565ab922e0
z02c0a8cde674a11a057a702f8beead4bbfd1b07e41478f61ea80090febc87251ff2069fa9717cd
zb24d8d91d30412a6f9dd5bba4a412c92ee811341295becdc7c0cf5dd16f8773124ccae63fe7bac
z2d0aec48271a7b4eec0d28d7bc5c791b920cf9f12fe249758a9d51b086d0eb19a5dca518a54ee7
z275cfc143e97fe10058fbf857a43dbaf40037279dc64c154a33236cffe96c83d5799ab6d747e32
z71ac7885d6c6357a61ac8a46f0d4a958799b7ef21ab8f6f24168d60a809a2006bcc163308b1d65
ze0d64c26be56bd5b223c75683b9d4af92701ba1c459777f98c55143d8b86b059ee9556fba1be16
z913b8413ecb75d585069754eb6c8cbad84651524f146a3ae5065c6773e2310f8facecfceb8b255
zdd8b8d6327e660a9c7dcde7cb2a836e3c2f997f96999edc647580a6324ae721c851822a22ad399
zed6e25043ed220100b3a4a66c3970b3a87b8e55065d0622a6ae58a73b9ac557d128dcd68dd7424
z12d1c577aa249df3fd301c38a5e3b39c44ba4940e640b725f1e5108c68cd1b271bb02ec6f7b351
zd73f00c2f44f7114c7bd5353cee5b0e7afdb004e86077f5af101e04ae8ff36f98bc2f4b7b4b78f
z0a276624be63fea9fb14ca0386e5224b77c9cbea2a403d113f41b9afcc067d284c314e2a2a5b2c
z28a48d31df8e07d1aa1450cec5af4bdf0843d6d7166616cbfd2b4b95c4d193467478f375ac3a7a
zf391859de63b3a0ddf9d6e9ab415fb2abb7c3d12e252f7f7047c2e726b8d20242741c4723425d2
z92afa272a95c11c76d296536974a988dcbd2d47d5f152ba79938eec7b7bc1e9b11a0a29c36d468
z6633ece9a96a951c6b8f55100555474185ace791e081bc01c4fda97e3998016b5ab03262a90ace
za9047b30b2783363d6cc596d450e58343e4eb9817a9482cac3722982efaecbf8ede82bb4ce28f3
z35b19f053de84d8a0e6d3c104c945928dc93e313101002982dcf847a550475b8769f53d773011e
zc8faf527da1ec65468c0b230dac3800c7d8d020cdfbc61094136cdcec8b446fe15a1f096d282de
z95c190781b364eaf7bc2bdd4045e4b9005a2f2d8e2b5a217e6abdccedba7fe084c7ef1cf8d8ac0
z78941a5f12eb3024a618818a8d77404d2b3719a48be482a7fc8dc89f8b4b4b802522b097939f24
zc9c370f40c1afbcf99c928e1edb45989a718b693424788b6c90fd087f0830c2dceefbbf2b4682c
z8643cc8ec96c1523653299b39d5f60f751970cf34f68196c54ae624be6c904545eb476b18ed1a7
zbb0febac77fb91893dec4541f8d4c871cc628fd5a7c7788caee376d0e1b55a4f260c53e9c3c7aa
ze8560d38349998be893f3c8afdde5da56bd5f2f6bbfd35082aeba83551a85769bbd05fbbcc9974
zc11f72854ff61c2073aa63fd0ace53f1d49b6a972c29bb2408c46077a3af21ddecbcb1aadc5ded
z233745aa4a8b683592987ce1aba3716df50dca3dfc9a2f3e8a20bd82adf08eb2267c68fa66b3db
z85deda4399b17663bd2f2bceaf8f6df46989ac37d3050a91e43e112ccd88aa8422d17b55575d51
ze56eaa31f151f642a2e382b404d096aaa04c3229a77aa856247468b8d652268bc4fd29b2dc4343
zca2871191c5b98b84471430d5991718f8758aa4f035bd3abe0593cd2e120b8b105b14411c23498
z4d2d00c0e42c2114d8aea3e49ad67bc3de566813aaffd7e898d3ce24a83f92b3f7b64ed94743b5
z1c0dd63bb4dee068871a17177cd5bccc3cd2e045e2583acd0f25fcd5374ee8d597d3ea4a8260d6
z8bc359b1012ce0e3afb6491dc457eb91578e51eceb2763b62c960ac315a45f1eb9aaa863e24512
zfc7521fa7ecfa738edf816c4e1e6378e7cea6cd0dc293b0a897d14d8a0e4c1b54920676525d13f
z6edcf6d3378e9a4b832575436eddd0865fe3eda499d8b1c9736faa2d1d2723cbf40be3073f0759
zb27be0f401c1103d7b44846d902da28af8f5bd98f2f960d4d53a3f79cd3b1dd0d576a15a620a37
z213ba3a8957fc49e38823d49718dc796c5c4871c09cb88d4061d135d7dfc494b0a39d35e6d59cf
z67e3c213f0061ae2e2b7e15a0cd01a16d4eda891902e49eab703acd0e8433b545b255e9ec327b6
z0861d5b544edfa28f9656111e2fa96bda22c91d9457a2b85fdaa051555cb883af525cd21b554f4
zb85d4744af552e775a508232c22c4368d915f7840c2858f4c8d826a571121094eee394ebef9c55
zbe61a61fbf8bb8da39cc148694008fbbc053cb8609fa111b863a1306c8c064aac1fc0409932343
z0d9f71786e147c16130f80b2aa65f57212083d8c7e4f316ca03c5ef04ddc8ad850d132e23309f7
z665dd1d31c84ce1de5867c3a7d545ccb278024676e7f31565f060bc74351cc174691373686d118
z5367898a49526dffa4dd1434e172aff869f8229725ea36f2cf94614a3e41856767a5ebaadd6b16
z4e73bda881b1d4766135568dcc72639e51ae2af8df934f9bd1500ee6a0743b5d56eaebc09bece5
za8de81275745069d8cdedae4c9834ef49ebcbfce1810a513b6c701f1dd42bf571e14ffdedc7f36
z62e25e931232b6063c7c98141813ea68e3d1666ff471951930fd85fcd400193bb552c40e1a6935
zf1ebb87e79b51e4c18621988e2de0055e916dbbb442b1652ec4a0bc135d06b64dfbed556336f72
z700819f9c6f038e99ee40f97ef9a439315ddd3c736ec5d04073cf1c987cf4cf5cd1a2f2c4020f3
z60eff15c82c6e53a08f0c3883b7c85d8d06b8a8a6e3f6b3e14b9cd0ff9ad58d5ff86905e891faf
z2b08a6ce22e629b8f5f6500efd6fb688ad0a288489764b8c92588129c9bb5ecf67d00ddb1f1a20
zcf3d3a2598d196d018c5e52a04ccfda0e27902c69a3afefd268d68002d17552c1f11d31280e836
z860c658a288242ab8c0a1ad3f5ae188e05baa62aceb1e312954cf42eab6a0985f1957ed84ce0d6
z9babbb35ce790cf07e0cf2ac34f1826c95ac516a41ea97a9c32afd5f2b2b01c2b4438904858423
zec5076426df73a35eee676501318220b4792bbbfcb0f3835fe365f62c03af7776cd9afda07a0e7
z320de53b81a4f461dcfb5339254e6ca891d626c24f02b12e59f68600cf054049e2efc6e8908ad7
z6692fe3033a144cd9b38baf6cc592695b4484d59e262b1459130620ddaa94766236a2f2ca95f4b
z915f22e2cda16c3ee52f6401f3117351fae6e07e260283b17657eb1f62a90b2c7aabb0189f5125
z176a6fc2110b6de5acb08ebfcba002257533f37c1d41c3263d23db7645b2457c1a92863d89fdb4
zec05606fe108f33d04d493469eb80f206e2df1fb5be588bc32ada16479b0a53ddc41e7f32eafc7
zf9cb697878e6c25598ff4335d5b0a06c003151a982ea341da8ba78b86aa143b1906bc41ad63d6f
z24e96fc27d7839c0e072e7871a255d21f10c487dd4202564066f21bc539340fd84a08db67fad09
z94521f45da7fc460ee3235d6fc1f8c1b020d111a68667e78798159f7850b72169cca283146c0bf
zf6ff3925344a396438897a23279b77e522c1a6873db7de15c78fd3a1dd07185c1865b1a019f78d
z2427fc0ce9490655e20baf32b15162ddb6ab8f00f7b8df580fa3cf62f61cce1295ff3adf20026e
za029e3cf099d675db15a07c53b581c75913f56851da1df131610f556b5c039b6bcf575ba4cdb7e
z26f05e58fa87c63ca3207b6b578074e505e0805464abeed1799a8d6480082cc960b6699f03673d
ze3e20ade08a2e2650e5d769e51675678c4f221ac74d2cc40abd68d9ae8024f7ced475d81d62a9c
zd69c27e93e0987f1d82ae3977a98629521aa559cb8b97bbd964414c9cdc308e6a5216d0efef147
z89a4da63bf9c851fa45041f88d5da7d286cf750313828500bbf05b5531f426afe779bb02aebf5e
z1b809c32c49d7446a56db91000321064602cce820d9780b42c0f95ae8e3c15546f041cf37bb943
ze8685158c7267aabbb327c036ba34324786c9aa7ee0dc6c57a93fc0708f28f195d2950f372464b
z1681784e4edee6b386ad7354c140349fb9f72a85ce028c9ed8b430d43a8661f1fb13563fd58583
ze90ed65941c52b987e70c146d99e26f56fc23368700fb6e59e35cd80f657f47596ebb701fa5fc7
z2e4424ddf70cdcb329cb5970301a32f7c33271a999baf91b997638f3c7ed08fd1ee289aa120121
z95871033696f9afcf2e44310f7ffdb41dfa66d55beb29427f1c206f0c162ff9c7df3bb47e77152
z6dc3b3aa9b6591f27f08988c4668f883a514253ed1594d1f7d76db79da2929b1ab1569adcbdb54
z67bcd2fea8de6adbd99087c26f8f79152d24e1ae16dd5c647969c6a71846debaf6b4a7e07355a7
z92ed4f74db138d47093e9001eabed1d3d63d32cd1d7f7d04285a1805dceb39184b14a9268a6c9a
z9431a81ea4fbc6b4aeb09904477063699a4fa112a1cd1dd0d66503605b6ecc42938b982c41081d
zc8af12bd839e4498be6978b20814db0c4913153e9c2e0a711a4ee9a4e177d5068656f1fa928ec0
zda35db536149bfd8d5608ca816482b0cd9f637b1e698bce5f260e026b3bd1c387b47a19fd36542
z7612c2348f5e065ac34c5297cdb8a931bb8b76fa317f1260c10e1356adbbea49d8df32e1fc4791
zd22aea9061a2a29bdc43815231016c466efd2581c5075ca0d33245d784ffb7afb47b690b68c92a
zc260580af3f0beb0306d030b3fed80625842b89a4e807183c437613b25dd72102fab4caa6f0ca9
z44d926d15b2240328168dc2f99a701b3a311cb91eebc0ebd99c6c9a69cc2c6ca2eb4702e7477fb
z0b5243e57497b0acc04a55c01b76e7683c3b3ffc635aa27e030d93566ceb53873e96cef8837e29
z9cd3b49eb6bac35e5a13cb8542a728c70ae61b4d3da65874086ad401db94471096174547869f5a
z61c7e42d6a16a5932ab2b9e1e4b6ae145862a3b9e0d3984845e7c1d4700b101cdc8c530c6d2581
z1aec51c3ebb0926300f89defd4e016c012d1dacc2a92c7e42477ef1e60e2369da143e48af4749e
z49ebc2d6ee4f3afd6877e1650d871486bc97d6424761fea6f9d067b9ebd5335f3932783c1b4000
z2a9700c9a5081de685a34d4085e84c1de442304723917339701c492bf570bb2686f015fd897c4d
zae3d28935251164286a504fe2094aeddf3ad65e84ae34577cd28b9b7dec70083eb59d0a89e297a
z28a419c781c90accda0dce5f35d1a72a9eec871de697db85447852f9a1524ddde9c89b4040dbbc
z5ec140cbb52199dd6e9f5b167c6a4b6569fa3f8878eeba618d885b358a83fc10816edea4de8a53
z7e422234cfe7ae43c6d5f386e59c70d07acc566c548b6e3024670903f906c4d48909af82dd82a0
zb462bd87732817333947f5393b7133de2f3aa5bf785c33a6082837e9f21f11e3842c3004047446
za2692a1b2a55949ca4a0b3b027f4cac2b27b7460f6dce5f82154648ad4321d7f2b9e9d801c6f42
z87629eab3f4b3d42781d1900d428a9b5cf46448b16f9d6f350bbd9434ba05ac535e510099e57d2
za0e88bc206596ecd1a3c00b4a900e3f6bf84b65bc1931d9dd281e4d4ed45b2a7e865c3588e6160
ze5a04e32ed01e9e37e0d9966241414b47353bd2a81a7780e2ce51b4a68b04c7cdfb2a7a956fdf9
z6d6d94227a2c4a5bc9f88b5637933a702e4877f3c1358fc545459185589bb949ef6319c1b1e2ee
z9ad906bd36ccd77929ade0e9172953b0f5b795ab2674f8330887db386407d0a850367eaa5e0b42
zd72f07881dd7f61a6755aea38aaff862d673a14699fd950fff2da7c03983b41b50e776cd91b3cb
z44903a753e684bff26de3d28a3659e2daa487cd27411bbfba9998bbda716945be4ceaea27d1cfe
z9322b0648b25e304d550448b5474a7cbd52a1617028acd5799ec91d76896c65d01fa662e006260
zcf93a1a11126afddd58f3a5428bc259c08215e68513531b2dcb1ee2ddc5be12d0febe68ecb5f59
zb9f1343c2fec84d0e9df1d306ffaeb4118c94cc00ba29ffa949bb9b85bc342c607a6a04bb34246
z9ddd7d1bb93c57bb892c750245dc7712812251a8a4a2acc0710f660ea1bf6816a47b95fea5f851
z418ffb03a8290305d91c245f41ed72e07443433d71e756705057938309b8733ab3a08c9afe9c7d
zbf40dd916af1b776c9ac47124ee04c18f1983257f49c7263b8b8ece47b79733279683eb76d6779
z121b30f11e1cc7515e87612bc1d9ec21c63eb4ae45d92c1ad547ce005895cd776999bb3d24f628
z7e3e20017c5a271be1ae2b0ce2cd2b651ac33c599c9b2098807be93dbc81a48b6f3576df7ecd0f
z3a66fbc927eae34d132c74446814c57015c870ca9de7aba47222068eec45a3ed6e94d40d9880a3
z9e1c0b158843293e62cd42480dbcc439c50776ad7095415bb8fbbcc4ba7300da61e192fcb43661
z2c6b694e1f2a8bc61e7e43f6f05f4e88344e80ab1c12ebaf1525730df0143e4efa0cfb820f9932
z95be18078f0c87498336793e4dbf287bdc5f2bd6aaed4bc251d4113e26c4cab5b0e6513a8fc71c
ze7d1f8ce6ca6afcb8669e50f577fbdfb1f572f4e8ab31c58b99d4ec845baf26caa2cb08d7f13b9
z50fd448dbde6ccdec2ab3ce5cc7d685ac1b0529cc90ea30f0fab97f84f4c6456b235c3c12a1315
ze528439d219c96a5f29d8a262cbc6694562252f52b2acf346e8c4e7664b4c49513c8e98ab2eb1e
zf0936144201fc6e984b56d0471b672b12bf898a6ec2c0ac57e2198eb8c88bf5fe29dc900ec6c78
z036c727eb78e2e18d375c8e1fde30a6b262b7f42afd0215199a12b6d90456acae66f0dc4c5534f
z1557ae778e5fd5cfee37990f731a0d31e170b2710016f3be978908c4da2fcd04ba41c8cd6d0548
z7637f8a3eb36219dbbbcd9d98466d43379463de392ea08195604c5c55c8fd3ff8c036c4f877207
z2efdcb5f72dd57f148a07e064133d5f3cfd7a7ffa76f7ce78f40b54d10b2fb8376ae116682509c
z1e900bae7a3e61c55bda0e71665d52dffba6d8109fdcdb614ecd923add5b12708d774a2a9b4cd1
zb8691debbb088b054dc811d3395720f130b2969c0c20235381553b944a2555852a2c17f2847b54
zb8d0d2c7df785a203ebc65d66236776103d37b72d15c44ce3a427affef16ad7a4f0732c5ca62bb
z36e00c6eb002e0679c7a409a66f4b18d1752fd11ab63fb9f2bad25977c70600aad463d6f61caa3
z84cfbfc364cb66a9400692a80346e5f73f11edc015a798ad1ce4a5e1ff82b093de74c9649351cd
z16d96a6080386c73346fc1b418fba67792de10d5d0ad4aa64cd091347f5b143b86fcbcf95be6e8
za6b45473afd72c59b5614194e585bc95deaff591d192d6eb0959d0b19aec6932225b63706232b5
z1a96c5f23f9a06064f5030fc7a75904094d5de318478eb4a15c19d082767e7a4a61e567b003113
z8c187fc3bf7d5ae5286df9c26b0e0c514d4c5240d63138e88edac44d13063901c44628923373c0
z38c79755d1506509bde33957927ee883d5f21d1a05af546eb553aa8e607f20eddb7a294fff39c1
z2bb18e31fde0fd62d458b9f40d2ed1ba2fd697bbaecc41cad5c86db076bf5c181b1f49c5a9e716
zc4a2c91f14294986ccf27065d36d2468a8eb58911a5a361d37fadafa010b75af53261cf118c009
z46d340e773b4176dd43d06576f590b07cacb448752288dd8b33aa5e792c1eeb161a494ca7f51c6
z85079478240636df2b2f1e747d626bfdfa904ea8597ec262222e5e026fee276fab72a66f3cd19c
zf65c49bc4518e038e3b779727e14716860444df2532eaad3994073e90890b3f7ba0b8fdeab29e2
z0d02f64afff1e28248d78e6698dbf2b731a82e0679e9f73f8ba69ff82c0b0473b9bb8b3055fcab
z8b4292ea8efb75f034444ab64a2e9a24c2e1ea9195c537a418e76a71a1b81fa645d4cb3abecec8
ze0ae6b905b86440cbc8a841701ed2b898d452dfdcb2cb8ba725f57568e94dfac1c4cfb77a92c43
z5e32aafde0d351e3768ce4da10f8fa6c017968908a5045afb7cc227ffacb1bafb5c28f02ac65f6
z2c78a737c2ce4c989e75c9d3777dc94bf6aaa894b6bac2b91313e25054c8436690b2615477e50c
z3fd1b0f6d9d93c630fc567c66bc215d82a3a30229efb3ae272fc67836014c557a7450b1c0c6524
z6b9a93970ee1eb06cff756d7cb582b981b79a080207d9a56165f07c937660ac7989f9f88314d76
zd8e2ca3bc5cdb243f6b483e5c2c9c3d6c2f19589b23a49e5db444d96201969d714b480d557f8b8
zaed6becbda134a056445a77b9ec6ef89555f59584b77a6d2c923245af07cab6711b052012c350e
zb24ad2f9790d423876f6a041709146793c5cc44ed2ed59ce0ec5e8fb77f51f65e4e6d2f7b60eec
z7aefff74d4bf7d105f64dc761be07845a4616e3300c869db56d905d6ef89a2a00ae5928f1f4c28
z16b21903b18b6fcb9de9572aaad4b2d0779a18e9743c2cc706c407c758c83996d2e1ecf4c1aaab
z1a29d7704ee7a09b3e598ebd1ae06e2c0d60dd078c928679b0ef981055fc7c945907c55c9f41a4
zfda2618a735507ff703e95b7327397f7dde152af06ff29c8314a2c687e7151c0d5f94c30c72662
z2d27fd1ef5eabe04a8f3c49d2fe76fa1a7b45b08c938ffdf6db89a3c90dc247bf2a9ec6f7277ee
z391bc54deac319fdc5ce3d6b6e69afd8ceab55b6dfe0bed816af08563961f6d5404291cb20eabe
z4c06dcb88f8ef37986ecede9a39d09fe05d8dfa3da732a16f27b74dc7624fa1ea3cb6e93188f55
zb57b7f04db202db38ba9cf7257e28ca26a756800ed8f613e713f3d8dbb910952758bd8fc75c751
z660eabaa1d93da992fcf772ab1075d1d019f87df50ebb6d897244c1e6caf6883f5db7c9056c43a
za661fa2772c99d67c60fcc114458d1286cf2ab4569a608a5ffd594488e2873c54731c0e5d9007d
z3a3e1dac7c6f692f267162195003ba68adcc35642e4d59043cbe864e9acc0a9cc38376757855c2
z19e0b577f6b0f5fd13ec6e1039a6a37988a519ee1e3dfeaed0cfbf4819df67d6bbe4659f773236
zaa57796126355be2d32b273057bab9f77c6cb40518c5a1f8b5348af5e4c06ec8abd2fde9ddeb0d
z2b99bc9c456c4e901fa1e9ac9f47e77cceb455dfa35646602fc22f441fd181fbfa4cc540870fc6
zf7655116ca1eec68f138cac0c720b5cd483521916e731482363b028a716653c7e18e248615ffd1
z93e56805ed6cf36200f18efc7511436a03966520cb3263326fae3bfc2127eeee4279216e5cafb2
z64d721c40511284ba38bda55bec1ed7a0f058d44662bdad87d80d10a4e240c41d0b0d0e1bd57cf
z069e9f047dff88c33f45e825be6a3956150888fa1906d276c85d056736a798ef33539f5c213dd6
z0e9dbe3aa58b51499ab05c6c079bb3862407f76e117719ede2230b1460fdbad99ac44ca3eae679
za2b7c100103691dfff6a94c06d9f3a0a35e825a3f7409b9adce7fda988e2509e31a3b0504d6ab2
z0d1fe5295b51038d58b03b30e7a4cc4157d197f8af76e151fc5e2f100284953e85fc2ba5a8df9d
zb406d47a0c1be1e9cae7b63c1db971a5d94bddab9d86da220ceb1fcfca0ae5953d0cfa45560c29
zf4d68938e2a18cf9b67b630e874ea9f8b8253f46140cc5dcc003d79be342f9062ce04cfaf7a280
z7e8b289191cc24b522ed4073b280681990fd42e72f6ca737ebd73ef455c46fbceca6a7515ce5b3
z8d77d6648718fb643f25add0d7e69d28142ac57155436b770505d83ef20c65783c9480c46c8140
z0471fbd339b087c103758548f92225d10fa538c01e65fcd4a9c34cead4be3a0c5f7a3a834c2756
z6dd8db68220668f5fa91da20196fbb66fbd789f55f5b2c798ccb19e96dd0fe8092d8706dbc16de
zddfcdf169eda1ffa053daf7e26e3d8925baca5efab2db784dc32e4fcd973fc73df33a9a393ef33
z2e1560fc4af3c7ce11361b8cc09cb3b8d8ae8c440ee4f9e495ffc69d26685f1948b7d5f492023c
ze4a6d65e8803287b2e67ddc2a08d72c271699cf885d2fe443f9ebd8c6e50339ca906aa60d8477e
zc27008ebde322dc6719fdc346601a86d1d5c927286d23f58ccc74b6df156fb8a4f3e7b16d6fbc2
z065597775d5a522c8d253cf30b7ec848593a13ca4284f900844886b2f5e8a6a8af94bae548aa1c
z8594eb31304a658b20edc809e584c94c89b79fd7a1d2a74ebe86f7eb9355985106aa6d35a4cb60
z9863682e46217a5f6b1098aab03fa1252041044cf6ec6132fa92006f4b950e5de24a3b28b78a51
za4b478a665e827e6fb193308139104e023229ff853fd9f46d466da78c770439dc75061f8908ccd
zc40b2f47c0532a541bebe8ea36aeadeeaf5a841a8151e6475677af5cd294b2616b416a9bf8ea34
z37a5894f9a7607e6eb70f938d6fb93c8632767403a1f3f240133b2f66938c727b77ae11881ce5f
z74f12412fbddc366e4e63719d08b86936bb4bb59b60bf2a55bf8c526f4e80e9fadf05601972cbc
z791f29fae97c3e096144b7fda3dfed552ed62d8c98c44cc10f638313c3f9c8b4ae0718c318124d
z18988716fbf4751f80223434543f960211199ba84a2e0c0dd896ab17d699d56273c5fde6a0d1f5
zb5595bf56bd54fceefe398693ac424ab7fc3ec7c03996fa967b4ca414771ee94c086c4d1ff1af0
zd757ac986ad571d1b8bf02d91b99d6c57d260632ba90a87bfaf4fd0cc04b9e8df679667c82f4c5
z8611c9b006a2737a65d733997790680a65b502bae1a3e9493459c63d2a83d3a2d4ab55d85d97b8
zad498431c1a8bd0f6ebbfa0c55fb5b79dbde6094d7debedec76b0100c09f2d4ae253457075a4b5
z7b9205b1b0ae94c85aa50dafe6d684d240430aaa644be1e83f735c1c6ddba259ffb89dea98a2a0
za4898c70b9e90188a21e81b8984a8b1587ca115206468577e72d60888340e6cabae46800041abe
z0b2d330a4d46c0d1c456288dbbd4ec53a81202d8dbca4fceae08996404f0c300c0544775a99975
z9bae3d9b6d5e39a73763815192bd9558661e1f4faa718ca1a007cf9826c4f241d28cf484ba6172
z2d0c055414573f635773215f8290b3839be9f938b58a318f913f3a4079e6d6dd8bfddd46483b5e
z6bb4fda8748913d99bcbd1a6332805993d308b141f3de6538f3bc39f455a1768c12caca643bac9
z4906188b2ae76ec8c92b3486a6acee20a7675830941a12a1b345ef4b77a031df594dbd93aaf699
z802ca5cc827adac0ac887cb124deb9f2cf323be3c741b9b08fdc32ba3b20b29844586c3447af5e
ze0a029ed452864eea78efe78c6da3f4c692b88857fe9471c568cb796fc31f547c1850dee9fbc8f
zf34e123f6543f9629fbca2b79fe9eabb39eb28c878c15ec562ebdd32453f6e4b14ddfd77cbc276
z2cf77b1ccaca1bb20a91f01c77d4080ffdb667bf7088c989a62bd205949d190acf73054bf8434e
z85e7bef136f78345d1021dc13f32c081eb99bc9e29c4a66630f1ec86c44d5b6122ae8e4dc4d7ec
zd221a9c9ceaf94e7d19e9f6315b415c8cf82602eadf645880b46419a1a60ca240ea77b457c3f4c
zbc6706292906aac6dcddf4f304ca5fe88a63d7f2c7ec7332a23c6376a929debe0ca89898003a4f
z12d471056dec1dffb5705e55e6348be7b2ce0be7d9e7c15dd44c8484e3f5b917c695d065f1bcac
zc2c1727c57463bcca05951d8fe68faddcee7889239b12b33246d84be8ec4b301b28dfcb4230f1e
z6e0414957fdb614b2ba42a8384a21aa90334c88f01dc1c809eeb24c5b18bba021ff34264ece2f0
zbe8510d8c7ca29415f9cc8764cc5715b85a4cb3e4f6516f855adee91e19570b50ce20f7062c70c
ze9ff3e97380070568e6a51f26cdd1f189b192f176a44a5c65c4e0153c360712a4e91d7c1ff8041
zaed5ed0585af9a45d0213228523e1f8a6e835f433697eadeac72f666283698eb6e66d260d39636
z67317640fb152fdc2303e845a7d9832bb7909ee1e0a860d1c60c2389c4f63b8e923ed37ee7028e
zb516bd29f6a551ef51dd150050fde7006f53a3cedd87ba6758677fa7709200b7bcbe469e8fbd2f
ze505e6aba2bf48a67ccd8ed16d45b5ff63f65466f7ebd773c1fd3f914aa09d1f6cded5054baa28
z17744346baeca1aa714d97bad2f0274c041cd9bd38b8b7a0b099c77be7f3caf2d6311b2e41658a
zc1ba8409c4ed9597fbab44d0709279304caa2acc8afc660e1aca933170e4a191f5123ff49edf02
z23398a0e758f9c5998901bcd72cba83cf22877b15a6d71f0095dce65a5222fb30f1de7512f36bc
z290f8fbf0f77a9fccdb3a238ded00a3b2927fefe32cb241d110f74a36fb66588a984d3f09ec3d2
z1f3b9aa8d2767dfc3a8befd92bf024c6734892f30ead43beda23e4054b23937942c2343ce0d4c2
z325acecc00e5f5f5120a5401582d8fd073e78a8bed161a1f241b34f29ef2dcc00b7a65886ebf5d
zd097eb5bd962bcce19acf7b774c17938d114e291d3bf6e5acf39f80def76463cb1048e33b69c5a
z482388bdebc488c47e9bf8c28318846aedea0fa4038bd53bc75b792da55cf2160c2687d54f4f51
z68f43cddf875742c9e4f455e2b29901bedd529cb315e0de345f462d91fb1954d29452ef06ae7fa
za7887887ec102ac8bce7243e95295d0f1bc13a974df7f5ec03ba1d3177fe82c7388b64f267386b
zf57ae2721cea6fb2769f00d33036537a1f101dc2bc58a59e919d827d8cab8186f1fa28f3202f7f
z9a86740c315a21ba09f42163d15d872eba0cfce46528d25d8cb7906c8ac413f21c44dbed1e999a
zfd49f1c4ef72eb3cdf7c86e859374f5d1a4530231936e5c8a4912cfc7a0b2bfb9e94cac91a0109
z16c1fb21ac5634cc01f2658716d93b12f70177cbb3ccfda5742244c5ed8559396dafef15710740
z0d6c335db11a1e293691019a05288d1e1eaeb74f1e3d0202f59027d5fbfc9fce4bb3145380b735
zf39ff239fb4a68fa8fc0cfed21dd9733170edaa674b0bf4c7f25327736951188283ad40677eb23
z3b13c141b229c415be09788d39264a5e0da172bbd3a3ab669608dcf8f8ede66ce422b30cbd6430
z6c19bb39fd235bd2cbeb36315af4415c24fe38b60a9ef741086f68b7ae3d33088a09df1645b2c0
z261ada6dfedbf9ea2d23f37c861bb9310909a2500a6cdb0600114260bfa296051c93c1e481db84
zf92e0629cf4851f7970360f0980eb6d8f672454504809567c13d56ab1f2d4c6d7b238bd12da22c
z7e90bb6b31ba687ca1a2f740582dfa1f5d11ad3fde17463db9c4a0b9e4c0e60720ac54fc9dce29
zb77d5620f3282351fa5b26f0a9cca2eaae20f27f32e9775e273d8459beca2bc85502335ef87629
z95beff8611fc16bf1f629f9911e840c768fd003325542584029140e9d7d093ed58f9d2a6cbb314
z31a5ca057442ecb270f21ce3ca50a3ee67aa4c7fc9b2db79f1bc0bb866d0d31ca7cf399087aa7c
z9d3f122726b4ebbee7cf26d6e48e13baf21195404f63af29fa7859881b8ad84107dbff4d3f353f
z0aab03573e989f8dc9a75fb917ff91b0ebdb90c28779ddf21ea1ce5b1bfcc97181feab60ec62e7
zbefa3e18fb9de2af3ebcb327f87ad96ed8f8c551f2caf5d41f9f95b39c10ed3f4d4f47db5bf6dc
zc86ddc0cf2f45d1beebb809ab1c9a577a116d3394b075f9b7b4340ea497110b2dff11d5c411291
z9f50dfd46cf5558e2789eaacbce8d05210b4ed62ef1c23b26cddfe2db479c9d2ad11bfe2605bba
z2cd75a44bfb01ff66e9cdba0210ee8e3af50fc8b2efcc74223d86b384767b504bc21a83d884865
zbb86e8557eac2d16f0177ec1d364cd412e76640b0c3426a39ef1cedb40d12e40633e04de3f9cc3
za9b97bc9d7d3d1dc684e1b9d39ca4fc40a06e083bb2322e66bf7085c951793ba002b9ce940c38a
z6949e6d4a238d7f146658c288813635ead27af285cc7de4a5400f91b1ff4d0cbf734fc6df2b0d0
z4455e39585ef479a75d2a14b8527ac239c950b6ce77c6bdb7e649fd7be1161a1029668d623d331
zadf0ce88545084dfe3cba2f5d524132d1661a42acec76a3b2867fb0d2a3f1c53a62c2201b3febb
z546a615abfe33a6024daf56b84c7737a37227dd199d693afef236ab84e1f8ae0ae1e787fe89a30
zd4539423810b27c1678e2a06883dd8435b07551b1e9ad0a7178aeb43f26c9bcb48599c9cc38a3f
zcec22bf8052d21bf4df072801d977ff427cb1f132eca5abe5af99235152ad0737570b84fedc219
z3786485ff0fb722b7ee99cf944ca8c739a0a07f483d1d7e5e5c827a1833e14783322a9e7608455
zc87d2c1566d4abd7a70f81415cbc0b523e8bba41a5886c54f8faabf9be4a4dd062b8201b6b083c
z1aa9f0e81ad355a9dfbbe9d89f2e390f491cc8c7d946bd9379263534a852fd38b7d104864aa6d2
z7d166314606c253197dbff6045a01753e073bcd0392ecdf512967b6561d5493424436262283880
z699846770bc4c6d010e2170c51983eb45a615466ea9eda36209f7dd933952324ed19accb4c0ab4
z17a12456c9968dcb0a7647e78038300f9c5cca24b023ddd3e58c3eceded5e9594a777904541040
z22970bac778a3a8d38f30e37adb3b536a48e39a9f65544f32202fab8818ebf220fc66b7f8e9843
zb4273fa1fd99173a466716cc35664c69a987daa162f56b6d9a708da970eefb0ce160f337c3d107
z4e1980eaf97cfdde0eae50caa63ae4b5991cab7e57906729b27fdbe31d187747a28b022afd5d0c
z361040a3d692ae557c355036c407b1220b61d9206ff2fbf2a9722a4b760d609812c2f6ed809c6b
zb0a1bf10c8a0684a2149df8bf17b5c50c4ee81ce7165bc98f222254b1fdaa7709c4f55b6d5bcab
z4077133437c76723215386a07fdc17275dabcb89f20d4de5cf8aeefef8989efe4e24b0f734d337
z12b03a06d588ea1ba98482abf8d048482e9b3b9c8b16dc407fa45a2ec8906778eb825124d66952
z0d035d23b4004523bb3892de7178880e01199e49f6211ec3a9aab72695cdf4f0c1bba96e8bd064
z2d0ddf14aa9e8c68afaa972f785328decbaa2e413cedf561f55b8e4f4da848fefa3cba413716e0
zff73c949a232e3563c8674db1b78235576c1bde60993d2ba3addd1f397a7fdc247eaec87f546ba
z2fa32cb711c2ae78a59e65297ac8a4f3ad4f22c7ead6b26730f764554748efef88265e690f82b3
z05522a5a36924bb6a66c4b404b6d9432f4ce82142fb6279af30d05174c052061e6242a69ce2882
z942dee8089c6bc20fd1c3092af73a8f8ff570ce3001e0e6dffae09599183a0d5f13383cbdef332
zeb5bb673cf53ac7e991abda6e0467c54c512c920f34d2ec3d8f4e86d702fa6ca5754627a059a72
za1ae847540ee33769247b18bc501379072ee174a0b21934349870fd0184934c4a52755e3732c8e
z98dcf1ef3ae2c1939eb6b98fbb3c40ed6282c7fd59f43aad3f510fc2ca660547953e96805888ec
z418ce9e57efdfc4c8b13ab43027006ebd3c4faa1087f62d8ccf0efe98174bb27850c65881426d7
zdf0ebc6de1076c705e6b7fffcc6a365a5c9afd6db507cb32f1e54ce95434c303d897dcea238038
zb3aaca59dd492d8860f8c6a0a4f9273b1a38385f3289873090ea3363a5439eba922e295c48da9b
z508da95fda09cef3f7ac77624e972d57d74253d41217bcfd3844a9ff9814ec2c4bb154f0b0af4b
z6afcd4d03100d9618e607cb2047601c40877a6f614944d5fae401d5d6711ff425e1639e16bfb7e
zc57b025f7e5c178eb72e27d1d53565d1bfa0dd15d27a8de9c27d1255e61af05c3cf147f93a2533
zb314f41051c1018cf107731fc574b4d03db68fb6ea097c7fab280aad427643422f7f8df97a6cba
z883a9c3b7041bb55115ee515221caaf443c89274882d6d4c5940b1553cb5b6ae883450297b5331
z6d3a596c034674ee429c9071fbb6c065d23b9510fca1ee80c543e296534f546a369b11b81a88e0
zf38ca8119ef8face294e2ac53fdea136075e7b4ac5767f13288d2b2a357a8fc1bfc3c922b91e09
z3ce9f0d2bec09f9dfda4dfc8c7fb82ece329f1e0000af314c9e5cc81a35c94704e194c758dcdeb
zd58388286c9baa949e780f1fa204fddcc80097f46f28b090c769ae7558eba4def9241465ca4ef0
zec6fd61984529889f4a56be6105ca4d5b204ffd79cabd6a14ce03085262e1ddf798d945477f389
z10107b4b13b25968d91b898672c7431ceb65f684f9993f261476ac8d9f1dbed097c4f0f711d34a
z53b7ecbcbfc2f0be2b91330acf4598a820b7d1641a3b41933631480b6cabfa1435a9a0260ec6e0
zc1f68f556358f9e6897f4b7df74467b7d08b373a7c9eeee5cef1f3794653c317d19722c58a8799
zfb515c22f622e9581df7bc5c9efa0057eef02377bc8f5b8ef1b641b96d16ae75716b1474cf987c
z49b97187554e140a0ac4e344e5b9c426bd820a44f4e405659022eb1d15ba7292f02e46da6b32c6
zb32e7bb7ac7c2fcb3b87bf0942ecf220ec6fe251a13635f1cd5025147141e228ab3d99c34355a3
zdf32d512f96f6219be60ee5a3cbe69bf1f87ef03029acceaadf86e7c06eaf6b830ed4446e7e29d
z59314cc038c1c660f21e394bdb1d7835c11122c1b3781f8e71dbe2be58dd32cefb6bf05289a14c
z644e3b30bb5a6059874cf5db276ef8830d26bf52b999e30e6a2606b9c7cf2ec61c66a5c82bf4d4
z5d7f1b849b9f4d6e970864b2afd408d13a1b0403170f4d09110677707d52bc38316008f20f4d79
z01ebe807af7054f440e21f180600d1d097a7c14e713a9dd195b9b7e205b3d6959be79e185091b9
za13e0a5e8acd2d38ab698845293e4082625b4d6b3e341d852f416ad452d9a0fea3a3d1fd470864
za99da9f30abd857df63b1a6700dc6a9d959c79da4ba2d3fa73fe034f8fbaee164b3d10848f868b
z857813fa9f55e0fc62a101bca1fbaf178f0630d22f9f384482ae2ddbdc22047e8779a5bed5688e
z9cb22d8ee3995764c5d32ccddae8c9b6357d79deac8d2e8312bc371499fbf5417349342d4c43e1
z7173ec899cbad396971cecffbd6e3e1d82caf879ae33828be04acf951d812d550828bcfcc215d9
ze50fe2d6a04f6a7fcf02caf064c0373d0761a13c3a649b95d981b808f3596a34d7323a1190963a
z8e4cd7fe006118e384f2210d0c73dd23090d5881067eacad88db31993e8e5ec0c3333f5c7c4478
z08bfd380f7e61af5ec7823598e3796981ba017a07a21077f32ff351333ede3482a9a8578240dac
z3d4660bb172a75cef0db48530e8842c35800e07c5e3dc8a6b3cb97d7500ee4eb1c1529fac145b2
z06c5e1e896d49e7968b6bb0c40f515f969db302c09dea84446567e072aad020227199351fd6620
z35c07e7efcff4a87a033594b34f15512b768d9c5b1b3bdbdbb35b482307175cd1b5bddb7912644
z0507bf07d469767adb241e58009975de0a827148227e1a328e2eb6de4fe12630b6cf1ec96c517d
za02ab8449b8ea65ffa7115dcf74e9c4ace56bc1b7f8fd293c425c9ac54e1b8f9b289ff24d4b73c
zffa681f6ebd028c2b67f0af86d376d2966342aa39336cd0b01a3446e18718d0a17738edef0145b
zff62208d7acf86fb4d112f72f92f8013e8bcc66139a8090bfe7e2e57f9cd5b2bd77ce2e62453bb
ze5e2e6baf09bff55095b6ab67804159fed22df4a8968ebac4ba6d5453bb08442e35838ca4df829
z14eab1f0ba96a59153744afa0b50cd458d3adbd261f01dc50930fb815bc169575a9e7b610da149
zc0da5c60e90b7215f1f2f3acfa6bcc6c44a874df483044161aebcc3be5ad54ceac21b599ded887
z7fafc8f0752c9688635fc2e703a0def8301e6fb8f2aa77b952f95ef2c75b41304a8aac961d00c5
zdc8b008395401d841df8aa374135b62fa06e0898b2694d8137ae77d61d75eba21b18386135a598
zde521dff9a41cffb06ffcb7bbacc549082995869fdd204e095fc1d2e4058f18e15f516b07e0ad8
z04d5e655fd05fa679055899e6a41e97ff28ca7e73788462023d1149f58c3ccac5f3b3a54cd98b6
z636ba6d091f67832abaa61a9acffb1c4d2314f581afde2dc9cdf38a4169dae9c7d28c3af51fee1
z3c6943ad8db47b415127ab67e5bc72cefb34834f2d7f8a5c05f636e8a7371ddf0c898afb9fcdbd
za0ca6b5cb48a7087564a0d90bb73e593c7f04fc64c7b6361f7bfdfde78267164f20b7d1b7a32b1
z2365901279290081ea21c70400959de9165867faaf434a3afe96b8c8a2605f32276f3235c6833a
z5fb534f0326dddcd62e12c958be3f8b3edf356ccb57f120e156f68081ec9124ce1a48f6aff8d69
z9d0ed25af5bcec1e320f5d1edf08b24da5459383b6da5ba779ab4dfe66e5c8d4d8fecd97e2d2d1
z1fb7d993ab2079021a3f77eb6f105bb83f134259e39b934984954b408cc382c6048e6249c44b38
z20194486d1a943a7d0d647eef961f55d1528aeda87b5f44a467f6dd2a6fa0e1e2d189f0195352b
z493db8007c1318ca5f2a17011f049ffa66272ba3b4ae928ca6e4d35d19b56d4c04312a94dc4647
z5f139ec5d6691e585f17c27cca26228ea10ca0d22ee3cf492de087317caed23e9363cc3be428d1
z01ed83b866260a0e5342cc02554d932d9df4686744738aac01fc0adc4d7bdb6067f11ee1d94712
z7a06ae1dedf10415067ae46e1d1db72618c2b1de8c83986c76173ab83afab42ef09d56f67ddd45
z4277d04cbb573cc738dbf1b290a02c6af6413ec3334f1178a35529e83d1ca122520ee6f1e12597
z4983df9d79bc6c8a51a2c98910565510f84625456ea266a18e101fa5cc750e9f242f5effe12ff1
z869f297222a1ece2604bb56f3ada1b7839e1baabba14e94768c7e3179fe5c5f2eb1fe10a689c44
za57108fa2c1e533b3e92952b04722dfa165e64641439d9c2c7123acba5b818a3ba6582f8268067
z846e8b8227d786c88cc44d87c43b1bd1dc261ce47ce440a7dac68d36f6f3a2a709e938bbd8184f
zd0a4be76b07c6829fbee37a243a66d6923a637d30ab23693ed276a7d881c4c0c32dae4c0627a2f
z9626c0d290104333226386c69a3a1d18bd2ea5e18352e4c4bcbf7b8a0f2fd686bfc07398982ea2
z3112de5bc0ec0f047c42715a5f6a47b94085eab3b0f43e793e70b4c01b7c70333271d23e5673c5
zc2fd5744a72797b49ce73eb2d29505849ab0049433d343c4777654c26bbe4f78bbe9a3d6e4871f
z02b0b3179ac7009cfc62ad6420f51fc6adcb0b1023793cadc14d0a519e5876533b1055892a06ff
zb76abea2c86600a0f4c3b6069e004478b38b47ad809261b7f0e7cd13892caf99fa179aa8bd4941
z091c05da54c862322ee5bc64d91861bed66eece773a50be4a7ed4e0675c995b46030492b289a64
z4b2ad5c0dcec9bcb9b36783d66e0d9223b40c358f5be9a5ec0bcc87ad705ca414881eea22a3ec6
zb1cb36292c4dc0768b15cf9568ee3aecb266407699fd57a65f9ea3ff00e97a9819055613a3a0bd
z212f8ff84fb2e17b4e8ff93a133ef8596dbeee537e77337fc796b8523ef2a6018637db444527c8
z3c509825b335e087e8483c28a0baab6f5d3afdcdc5f63cdd5c96d9e1a4e7f46a49dae467743d5a
z3c62a4495d2a1e05ebf17f519b689314d080e19f5910df0e9f2f3b4dbcb064a80c2ceb9c119ef3
zb66c756268e3f18d5561cf4c6de96e0970097be393c198adbc81bf0b76f2909cd12c61a2912afb
zefbcff514bb4372ae9d04d4d67fe45475e27e3ff26c971abcac16391cfbe6571f61756d3596513
z079a76d7673c158606147a8fba1b99814d681005c556d31fbc28764bcc4d23cd4a873a42cea519
za4e900081b6850d72cd8abb01bca31adbbab34b526e49507e8d0f6ba6f9009bcbe18d06c77298f
z12081b157904e874184da42481bfda8993d98f948118485d24cc3fbd28be16db7c357900f06f65
z54ede0db7c67b5b7f5fc971dfa5479900964913569f42ab0664d0d18fdc4a76f9c50c534c3b1e1
zd2996e1acabc0951c67a2492084f9e42423f54543cb38a143f3d99f1feaedfbed2c5fd375b649c
z1d9b47ee16cd1d173cf80df5ec83268cff6ee3474819a83724f679baefb1f7ebe1dbb2368fe6a3
z596ce1afad6dee35c5a814160cf7fd75e3449ad50ef9b43eced64304953192bacf53a4dee02b47
za44af17bee57d78a1cd2836ae2e4ae13a950b4ef01492b6bf8d18f0dfaf1dfaaf00d59eb1b8eaa
z82f6303aee2e612563d00c700915ba5ee0606c7fda06d4c4fe7dfcb3ec954c78e94719e9e64e4c
z522a6c17ac85e969d25d6769286360becd62adebc00b11bfc02a6642cf6c98cfdbdea642d4d343
z937bf1132dc63e44d8c3a143b80e002272519be5945c8d0e3d99a129ae99c24b3418ef8cd8d93a
z4e5c0d2b2d1a565304245db40ea5b94852373a43d4f57ca2965d1e3355bf92f4097b660164f5ce
z60c912564e253bb455b21e3ec738037002746506e6394251bd6aa800773300a15db490d7d38a76
z740b5db08a247ffb2efb1e232226893b338871db0159987d72e555dbac3947861a9414690e1380
z1b41fd684ef852d89a862f49bfe030389e85b0555d5ade651c54bc945b05c7dddb7b0becfda4ec
z691ce79349ea69ff41c085e0cade5b460d061125b89a08bf36e3bcbb34d96d33fb131eb8d29953
zc6aac789163fd49292d031939af29208859dc2462b892e6b36669a2b233650a0627d42d301ef2f
zba9afd30281a3c7db09396f296f0eda1823997b47f670ee56cde5c9e81d068fe5f78cf02d506cb
z2f00a6afc270e8c2389cf53ec05cf0464a225cc5d7bd3dc529f3dc218a69d537f50ccf070cc5a1
z2114ed329d8cd645798ddb17e2720daf6be8065802c0a0e0411e7c9c45b716659dcc92e45814ce
zcaea5df431060291a80eabc7700b03ecc6f4c5b786b3a1f3959cc64ef2b12e44fc2c2c9d5f9453
z5b425a2ca3e0fbbf9f9de8e1b74053a8f6bfe73bee77b1e6ec9c0123adaa28545f1a12f9f275cf
ze904ab83878572bd983ab526218e5c62e685419a2f6e67e39f5be48d68636e7133e9bc5acf0638
z3c5d0a8cb8c6145d68f91619e34ad4b79e30a509eaaf3484fc840853af93ce9ff445ccf2309db5
zcd14df774c3eafe6d3ca04e8e488708bfb97ee61c600854f067e59e04731d3ec2bf4f61fe0f037
z2681730fb4ba7b419a1f40cd11a27f292ff6d3a56228fd0a101bcf51324ea9b37968a288820d99
zb0c751dd9c8a74509a71bab4d8688a131dde6f5c3d01a15001085b2e7bffd233d00848dcabeaa3
z6b4e05eb924e71d8184ab56fc6d581e83003d85dd264ab769afb36e6584c76e9318d7cbe3a22b0
z10e5132044402b40205c8e0a310613005ef0f1036609866c860d088ea5e98c3e56d82f396d48da
zff5f627c4a43209b7730972767b5fffb8bea222eb1ed87ca4ff028982a960ff020163e44b5bed0
z76d19fa90d48c2f5f654f57c8ed71534261ebdccf26e4b4033a97584e04aff7769e41a2f238818
z1f55c76dd6b222a6de6cf4569886c3e668fe7bf708a05bfafb3eaa51a51976e20cff9d686dd19b
z8b0713987a75c67bd2fc5e1bf9a1b208147777bf3731dc55ffc3ac8c448fc3c4770fa7290f9c1c
z8dd7e27b10a4f3db4157acc12ab9996460df27f62a0c48501e8a32386615d2ffd79062c964d45d
z6c04d53cc5ab60290fe5e60b1b96915c45e31826981b11e06fa2e1cb65973910f2333df9fcb8e9
zbc27c813d9888117a4eb7cc7aa8fa1a8e35a22d841693bb26c88c4d9695f2f5fa08b3b9f0f39d0
z5df88cc62e5651c86332732c140b0db86ff4ee94a993dc90934d2e733aa400f73ba102a9ba4aa4
z281bef6e4f0351723b36756b8b656914a10ab0cf5f69d68de7d49992905b74e2b076a73656ad7d
z4d0ac8fb5877cf34c352e5ebdb6084062df58febc493f5337f9d519ecfc8131035256b382a0cb5
z497148b34d720c51fe0e5f99028a7172e2765d35bc8c7feb64c0dc245ce64c63523a5815be06c2
zb2630357ac18bbb8b820bb2b9610f23d4c899ddc69cc4532de693af47855ce2f202d68d26885ef
zb444ba3c2256572bd0280510bab66923b6cc98e8cb6e949facbd2eca97dd5d675a58e5768cbcfd
z2284cfb4d31a2daa5880fae225b70d27d9f96078b738025613f95a22e26744c09895b7a416c8ce
zb52f1196a54294c7d1999a8967443012672c2898551e57da0fba6fa6e442a45da7ebd14cfbd085
zcf7f53d2aedb3ee6bb0b20f8bc841a84396d30d50b22cc4e477cc8e4973c2c9bbce072b3e3dab5
z204f360d69468a24d88f593104b099f9a3a29f941e1adbfc36d2be1395c6749c62e24ac58fd287
zdfa55c069e2d40b6b62bc584f269f5764abd4c40bc10927265fd27aaea4f8ae08871af0df3f505
ze47b7c9270216eccbc1376b748d5f94b440943f388e88c050935bd4ffdea29275eedf297ce1f1f
z802d34c2d3c031355e7a71c26dac7ccb2c572c5c13d526f20645ae0a1bf9500c56a3de60f48500
zcfebd4e37b2f822210e4f9ecdad10c66adb4dad57cfdab3fb5a94e0783d8dd59f25fbda1a68eb7
z76aad676480dd7e72dd323a5e95132c4c1f3132925c0848d81ce16d864062b59879757c1f159af
z57e64be3653c6d749cfee15f06c2ff62f7fc8ac82b501c05af442e3e19288ca76c80cfa0295e81
z1f5432d3e7a45ae78490e2205ed118606ed7a31c1ca46a579f7916b8ff7b18bddb9bf4af0d505f
zf1b2612e50364eae3334ab9058770c6a0d680d126bea3009812bbf7a6e9a091150742e35d2c19f
zc8d0fc099d62cfdfe91c847f630f1d1a4d522ea60927235a01f0a352838082732560889fc285ee
z8b59a077ecdd7427b7aafb4490e981bf68668ad8b208818c51236a3e22ecfe6449712c93826a41
z75adc22603f242b17e98a38e397bc66043911ab05d31bcc477686d399e341318b106edc057bea7
z8fb65ebd7b8b218d6b73ab401417d0568135568d7244e8f912fc9d97ce27fac8a71852a1829aa1
z32cd60b819518e0cf2213c311bbc09b44f7fb1ee29040d93bf74cb3082f6d1ba49ebadfb5736e9
z8aca8adc9a117910aee897e5f10e2ff271d8fa9a297b5f362a40bd9b832a46667b75f1b741d1af
z8470ce3488812b92c0f2747674aab90ebc0c9b4c512bfbe85d487b203458813b34432727c5758f
z27f15dd4922ac421307133c144e0a1837c01c07d3317052f8ec768e51e84e09ab98a524ef00449
zb4c9d7acb582a2f00e6eff07005ab0d89c58489f670c9b0eb4a02785101bc7844e375a6320ce6a
zd1e7beb5c7797a08289f231b29dfc28c367c99e18a10c7c9c81d94711e20da2d793e21dacbe4cc
z369a6452e3baaf315016d316caeccd104a3f9f0a20e1b7894d5e1bd755e0542476dd4af6c60486
zbc6803ba42a57d61199f1a53b715a278a4b25e41d298cbe64dac56ba35947931a9a0174b718ce8
z7941519421a82ba3a7cbe3a1905c36f1a35a8569fcbaead9d7c3aea087d2170bb17a377d36fe20
z849175e7228cfccd6a86072f0a79191a78974aa1039e488bf07e8e0b4b5e0d3f8914cdae145f62
z16d686f83d7d7dd37e18665cccd7f5758aae4319e27500059e78d0b9855225d3aeddd73c8ebbfb
z8120cccacd669d56888913b1e28dff158ef5d83b664cb94b16ce853eb829375e3aaf9651afb0d8
z27fffcb92984e007b5815fda552837f31ec8420f83edd38a56d36a5aaa82504621437503794521
z7963f27310d9a155be281c3b86a11a83e267f0d79c4272def97effdbcc242c9a38ca3e1f02db7f
zf6a2629ae7162f3d38d6014b3472eb6e8358eeb75e5ef69cbfd61eab97c9c928e8885d86684428
z72efcf9712d94468395c6a0e35b13c01f0e243c76e59a87a3e6318f85b0ac51f538aacec944bbc
z31a621037fad4e8b5a7e603dd7be1d8d5bd5dac29e418e6f1d45212853cc31d9aafc61cd69e6d9
zc2afd4ed5f5dc5562f68cdebb52fe69e67a5bcb207bf0d91437af9af9836996b1941f523725896
z2dc9fbd246297c77c97fc4043b824e4cc3bb637c63b4585e94f94dd2851dd59fd0d485c41691c1
z7a3d83e3b7df5beae90d632b8fd1c6b4eb3060191c9ab40cadbd3a018119ea189a119289624afc
zf9b7c332674fee9a11cce3b77790a5f31df8e99aad5a16d85c6071b61d7f3872060723477c39c9
z0872912be55cd09546b09cb3a46b8ef3684ee62a18c989fc9c4a82aa2acc5d6435512da8dcbe70
zd88048bd176a796344f2e4b9e21dee1ae3469c68c746b78fab2b5254daf950246d5cb205a5778b
z240f7a13b3208c30011299d564345b96fa91d890edb107ae6555e92b19b60a2421b0a5f86a13e0
z093c0967d79af9515fa363d0a7bedd45d395e9fe35524274ab33d6565fe1638fe22877aad3374d
z1c4644f1d5ccb47c97849f4909fc105daf783b96796e7294498dd57d5164a0df0e4918a4a41e61
z3d7369b501d89074ff835513ecfc46fff506926c3ecdb1bf51d8c069004a18e078fc3cc3ff28a5
z2db1e3f050301cf20feca0a42c5eef4b84ee8d7e000f17f052bac438b0d4d24a7961e8ad4950b6
z41f0702036931a24437ac6334e5844a190a658a6ebf18943bc16a56e53012c6c86fcca1937a8a4
zd166c21cb8a10d7c84bb388cdf188c767ba9316db478d9793502ec1fdddffd67570770a504c1f5
z4b1bf0b5055954f986528c0923b458a4e5d92bcf13ae1ef683364fa36850e8a67ac6d85cac5588
z2a891289a966118c9d8d8272e68822f3026528cfcccc418fd087facb25e21cfed68c4be3e137b9
z412eb5c60eafc22baa80ba6779a712048794c8f095d6cab8cdf1ec0757365c00eb3fb724cb2270
z23b442df77b2366ae782ffb9e64fc3bbe7c23b8fc738d45ede531d1ef15a9b0be297e076764821
zd26da5b2b69c028bfb73eaa3bd64280b26367b41d7bc5baa090d33005a4db041a65c6a78d6b0d1
z0fb1ae2e9c511cf1fee1b5d594dce555069cc4bdb34bcf8a676c0151f95db18f16de6c3ccb78cf
zc8abe25f4577f0c6d1236d460196469a9e8c3345f1da01a0fe30df574f449eefe722c5d6f4bed5
zf4f7442d0ef7456f4a673db60a2fa9a078cc92d6dd4e2e529e3924e710ffe87c57e7e246a4eae9
z45dbb2d7efe11530b1bb2f1e8b68f001f078812f19bf0fbd9db8d70890c44653cb35f28ccbdc6f
z065cfa6d81d01047aba375c106691442344b9f3ea93d929d751f930c3c3cb4cd4524051d25b91d
z132c96adee10e0eb01192eb51d5a143344cedf16daf8c3ed1b2c49d4943a57f4a04c471738cbdb
z69fdd3e028409617f02fe434d5d72896c57ee43ed00af1380255ad5505a9e408f5618695e59455
z012b621564fccd4b517c1c2623b430469373cac9372ea50286e31f3d0475561a307c71802b1291
zfba9f33449cbb8edbdc109314ffdfeb53b9913d27feec7410abf52987d58431d4a426bc2d41c7e
zb23efb229af7d2aa9182da74a19f4f592bb291390855e2fede88616a62b24a9565ba6e803352b6
z521a43e54433cd9b3aa42ac9ff709cf18d10a873a8913acb8678eb5e95ebc18eeeb648717f2e1b
z7b917484f710076bb0ccf38e85af7e10f34df37b7518523c2e45721f1d4071ea7ce2521581a1ad
z18cf83f29702351987b7bad1f164efc90dd2217fd3da0c4d5bfadaa77995e196e4907a938dd4b4
z5a77b26954b5cacafab5295531b3ba7a196919af5a6d83d5ffaf25eff7312a443fdd3422275df6
z7888684734132f17bb3cd999de2e532179ffe30a6c4a6b727e13c443f79d7f2bf25808b896dbe7
z0f9d7822fa0c4f76fcfccecc98b6fc0eec7fdbc088d4acd2da8ec391363ed47cc005393f0eb0af
zee1eb94d9d97ec2f3aedc602ab09d6d5b2099a60b27909e5d766d1a456ca82918542cf29aaa687
zbffd2a9d87eb85359fde500cecf6e9109f995c0b2180066854ca64daf193ece4c6e19bc4a1de29
z692a074baa600465ad6e2168fd938a0b645d2ad02c5ca9afa63722b6172f490b0e4ca9e383def4
za560c10410e5d756d02bc87f01c4d1cce6ccb95e714f1dd2da0500490cad7d998dce867163368c
ze2e8569efd827137d0099682084062e009329fe86c43fcdb05f8335b3c1f3c0ed568c12412efe8
zefcaa24675a18c1c92f69369c8d511d16ca924445ebe4bd3b182093c56d63fff44478a83048a2d
zad289f984d5027acfb9a5f6f255b19fe4bdc080a0af7fbbeef05814e028890d848dfa106644250
z2563d86cf45067de831a6aa7e31fb22c9d1d5b011bdd2201796231b36db35c5d79b3c02b13f842
z49e0df1356d5729145c09572daaca97d57fd268ae7259146c15209c019cd74a1024654ce6c6218
z186b9cacffa193400252bc37a7e7b5de3dad3a41cb3a6c1f2898304d63f76e375535ce0b3455e5
ze8af0bf100513e43ca1346311c4fa9032722ca325efd0755ace7888ed95e1a324e6fac797bf883
z419d3a7fae289a5cfbf1eef9786dad9bdbb2a4e1672c162af2dec08d32154156ca4fb0fdcdb733
z22601eac4bb7606b380cbac18f11e8972ce35b4abd3d0a1c29d23eeda0b8a2c8be2e73c499f4bd
z082343131d94d95e9b31895dd33d04919799fade72a223775db3240465128b7d966543d2dd8d03
zad8aedbc76ae081a6d37861eefcc712b374cbb43d59889393ff14a0b321308d6d58280e2861f22
z1da98e910f2b5eadd810e86d23e044d56bccd656f7f8d9ad1618455e20f69d7cc4c405aa5b3124
z6c6707aad6910b44f01bb1dc6be7171dff219a1247d1b0da58025634902ea2622d01c8e1b36c18
ze76acfc3afe8fefc18fd04e6e162fcb24b765f07a99828033c178160c81b6a4ace8d9b2f71517f
z5627386cfd8a147085d0e8c20d3e09bafda85323a8be78e6f07fc1c3304038b78bd3fa4943dd73
z22f1bbf04e97e9abe149e6d05794808e8bf3a5becc0e3e6fd2b718b824c6b4adbcf38048de1d65
z824c6086f96852ee320a113459eb246e379f54f79652ac0142769dc2f0cd89963e4645458526a3
z4284d607ab56ccdd33359b988d28c77c1ae87d90aa19086d613273e176505195c0765295613a03
zdb71cfba6280c21389b516598510480a003562b1cf0a7a2a8bb65ace574b99dc2c37093074322e
z4ffd676eb7fe0524b38697271a429e32261e4b1a6a7d35560c598f9d0c0811470834941ad9a915
z07625fb21aac6d1178fa4dfa9e3878628a1a962838580774d152e94858890dd337515426f124ae
zc00c13b5f88c206ae9f69f9f0dbebbeda9af8b12df2ea594a7d7eb0717e14e21fc776be45bcdc0
zca7bfd1c6e5a82abed0e4c25aa2208c92f7a552fa199aebdd580ad66502058d2f0091b48edea50
zcc4f2fce4f17d77e4b0545a758dd269c1b5583a36f7d1cc292396fd94f0a6a39e38b359a9e2c32
z9ac2e8ee29fb5eca08603730e9323eba37ad706a1027f18d0d2980e02cd4556acfc51f3dae2055
z41a29c50f582b29c8da36a190e2d6d0818b1a906bf00e436acb2dc511bac865f9c7728c2589033
zbb26b08bc7705ad7e9452da55c2db2c488ed9e328e95ed655fb7b79856c23928a9d88ff137c218
zb3cadb63c3c9bb44580c371c335e67f79fee13082cc27a2025c401c88c8fca99e3fa1cb9208e23
z58b71269dbc25f698e6946a768a35c836d55699b4acf242420e83f2c76039e77c528af4278fa64
z37150ed240482255745209e49a6271ea06e0567046f555b8b85214eab284f8667a9b61fd582083
zbb3530f150969a15d952fa495a3513b6f443c0f258fbfa6758fd9014092c0a9d61651c39fe93b4
z11faafb1bba1e2583f2fdb9be8c45d396f4a76ef6ffd4d66abefb73d4271c6c76de7cac6ee8ca3
z337a1fd6431711875792f2dafe98e3363e49b8e55e2a698e5dc8d939a89cc7c7d42e8e27b2c3f1
z99a579f821a5581df2ceee361bf97b7a8c8cbc45f4af69e3b3a5914998781b0c87d6b53f561676
z7e4974bfde7f6e6ef2d9f8ba87b735f1a79ca713f7fcbb834e85a9280b1b4ed44b3d3786ed8539
zf297dc0a78ce02685a036c21951c297bbbc7f9309974968979307429a8e780384b3997bef16739
z02b16316ac88ce52f6d4225beb6e112b52242ed63aa586e86f919b890ed0126ea525ca60c25486
zb98a519354db4c68253ca453af7c07b63a34d157c374e8f798fa2d79a00bf8a1c6ef5de99691b3
zb40aa46c8279af4f0cbf05ee928fc671246c432b51b120b1ea5710b6c602e9249d0344e5d79a29
z6194af0b2c71abe2cbabd0a391396a2b94eeb24264bb2f52342a5a3116d1d6abf8cccd5d1f7bf2
z66d77b9056ee83148a19877e68608b0803fc84c47218515d924f125be9637a6b7c25b54b643574
zc8f7231306269d7d70ea96d3f8901ebbe8826667ad8d8757dd2a3130442340f49810ba69a08996
z22d796509f8fc4a608237d057488c8417a53449396af6b30481b224def955e04c753b04fcbb63d
z0349afefdb61b18ce22840f53a6517d31b6659d897764fd540267f2f3420ec1c2c232bf2307813
z712a509b7279e777a4f5a2f4c1b5cd95877cdbccfdd58fda79c8b9d4cc60a775bbe0e8a85e4e71
z257cdc5faa7541e4f8a7cf3bcad47921673a9072c725e9fa464dd7bf3ba832f87507319773e67f
zcdb7ab1bceb1dcd2d761e1dd8a1b0af39a7cd32b123c40411b4540ac98983586e210ac376b8cbd
z6ff2c11a3c849588319531d0a908c3ec478a9eefe7b86f81ae50a868a7ba839207c3b709747edc
z323c8769196de8c081a1e14fde26a96cee03f844a88a50f05fa3c89046d18bf3340f8926132157
ze41d52212f33e6c08b2f7c4027f3cb6699371e5c81e1a25682ff14ecdb901a76dcee23bf4c4b26
zcbc9f6207004993281999b3479ed5d1f1da81bbfb19645058033970c071189bcba2c3fca3f7ed9
zef3813005eb81be0a77ef8b135f4dfc9eb4f74e3620fe42f9915513bad0b4cc0b535b497bfe68d
z93e5a557e4fd2ed7084dc1b609caa6c7e98f97427fdcd9055c65f4ebb0c61005268a84be8c9f2c
z8c1c0ffd829d5bce2d6141bda4767640818e83dc4723804698deb2df655123ab9c5e77397e103d
zdf98327b61bad5f3e6c910e25f3061783fddc59f385c42f3e8ad9af9f79c902409f17c8a552b13
z4cfadd5fe434fe674f0a4afe903410c4c1b5b1ae63a0745ef58413555e02434c33df5baacc34ad
zf91be5e88fe59b6b4941601458d8e03002810c15a6f1aea74a87e46bd22339b796484397171b0d
zc191811da73c66e512b6c9cd4cbf8c1845c2930a38a2019f8b52afcf110300f9baf25cdd09b6a6
z6de9fb9bd417b95709b1d5733880184c061c49054a5e3c33ee03348873271c431437690ba869f4
z1a2c97647c2cae949219076ec56d64fb79925bcdc64a509c9a71f347cb52e9087267c46e90e0f7
zfbf01ea3dd488ceaa89e96fa746a49fd2718e27540c3d04f088be9eab1d86ec551dd50be8f9824
z117c416772fb89fedc73169546f377d1488b052567435577d0ff67ffae26070d244068bc00923e
zf55c0cb0c20e47af78a449826935be4b860ccdf8c3e9aa742ee45f160c26dc37cd1f49bee83a4e
z55bdfc42474b24dcfcdc7bfb535175b516ed38da1af6b2506b816f6c25177f22de30a3c3773810
z9709d7d932853e959c79d62ce0889a2ed45c88bf8a194ee295da33dd90377e2d179d6718c677c4
z913b975262dd3f4abf2c4dcda5f9474cc63e8b0cb93893d81409ce1fbb0d48c11e506db5910a86
z11cafbffec0b931a905367ed34399afdf821ccc6eee55c560cf3ec470e303dbb19dea9a9a93443
z23dcb26df69e1093a020be13b4d0393d8d2e5e04e3a8938836feb20f0ffa9b548f6fc6aa4bef85
z79249f00cf8061014905b0440dcb158635ddbbd946fab3e6a5975b17f73253e4b713e58c45f77d
z3c480925493bfc80a7eaea99cc848f79f2cc1aeef6fe768233fe29eb461451be6a2abda8740a87
za669ebebe560b6390e458ba87225287bb98a9b917e205140f00b0efd7c7b2ecacfbc2bb2583a5b
z8fd689064cf7eb5c43712a6faa6597b533f682f7b3a58fab20432cc03cdc88800c43b45c52485e
z6b0aee7b0648e60e118057afd83fbaa1be1e5c5a49d8a1e76569752d1614f58b5d7c0d17a8c442
z958bfdf00fa3fc55a092a78523a4fd590e0fd73af81d8e2a59ed7127a33722d184d849a09f3711
ze8e4ffdca8cf32110cd4001c88aec231916dc84b8305bd1fbe23a71a4b9be0f4e64642a06cb1c0
zcfecbc275848a98bfcfd2b15e4b6a7b995240d6611690007229d94920b925c61217a76f33bd1c9
zd61791c24c6ce34a9a830ae1d5ae6c482d7600cf34bb2cb88239b063505a346eb6efb42a967d81
z96b11aac4078a3943a7e3f383161595312fb8598e1f4565af5def50940beaa90d15b965336340b
z727042e75032772239ce083409a0008cc1461838a2488034cb2f0ef86534cc39b6c139c1fbf597
z4a9025be1fd2ff41191529989ec32e76c93858bc98d86c61d135d83267652c974d2b6ff52b5929
z4e52fa55285ec415781e701a406e0ec78472e379909a6ca347b605e0491a5ea4ef5d7bf17e4e28
z4c4ac1e615369ea9c309a12b7fa24010e6750e41e77fa9883f682cb6e4f8dc5e032d62000c59bb
z4e37e7b948243a984cf08166363eaca866753118a89400380d46c88e2da95476a5b44085560d8f
z5bbad10708afe4427e6956ebf6bbcab951d48ed851ff1986d2a9c416bd134ae4a70111bbde132f
z125ce1e3804bf575392a287dd0415d478b2857547297e1be44617caf4912973db735d2352e0268
z81becb6082714f8751b9ae0029ea6596669808644bb9e3e325646ee45fe714f8f9a2e102d49836
ze2b5b037b9f233c84d93b61a4b0941b1c30f965deb1bfa097da44982d58f4579f8a94859c41cbc
za2360ade8c7d84d26f42dd01750c805d13d2716b268c5383f3130281fa2bc7b80b67ad6679e079
z1c322da99491fe18ab26ab1f1207406a3e268cdeda4e3e8f851bdd3b327e7c26c0915010481621
zf2bf1522ce3752d9e2ac19344eec527e611428f045004b69d8d22e93d7768f110182e729ec49f4
z54c664c53bc4791b4f6ff9075274d1b21e107ee838cb105e9872a398ee7fb7e3f03f1d99541384
zcd77b01291860d31f8ef581f3ea7776cf22599d87c0c9e236e52ecddca740b86bb6399adefc5f8
zde6228775e233fc799ff3088995c71b8dc8a0f2346f27843cd251c379222574d2a4e6c5a4d8075
ze09e9407b11f82035c6c25573f338fdf30385c1442e9ba5b668a2c4974162dd592d817543e9b65
z12f722bcd39e418f0a6e59f036f451e90916110820ae257df04c78f6c0d1bfb372c028bcbf8dbf
z8a521b0721ea7aa6f89f8db489cb3d90f212f28b83bc80b6345fd309f0f356fc346b9cb99eb1ed
z55ce31bd5d2ddd54dce7d49158fb1491230c57b33234ad34d24f7c61ea75e68eeecc2c198f7d44
z2d112135a6b12b7445d7504d33feeb57b8ec3707fc0fc8e7154616f2f2c9a17ecd8199d8da5d02
z4f9cd103337f12f2b47511c49eee5b2700bf8e59cf0fe1ccaeb908d811f0126bf18d6854aeb3b9
ze4044102f73be37a7588a7b329afd163fc1bed54174fca41fed7cfca434197cd960bb822b984ae
zcb62d550ca523d14d0a6ef2cc251db74843664fff4ad18ecb000f5aabdeda8533a554b2aef44ae
zaaca3465b13c80c2f80f675c3c25c1e69549c7c771c565afb63dea82e2f27ccf24f43d0ac4913c
z53c5074488ba9c794a3259804e4cbe3681b4bddadf96fcf65bfb4135c2731d449826de07845950
z4ee3c76192bed51afd20858c52b2f01302dae0f72fa886a14b46fac62d3902a7adc8e47d2ec9f7
zb037216ce13d5d33a7530b077b3a9cbfc67675f09138c5720a55b8cbf660c8fcb64b1092b5e554
zda98201032c151e2ebee8d3a6b22b4bbeb6c86710b07cb706f43be4c8558bc9fd7333cc379a553
za2a44496c5612815fbce9378fb715a06ffb6ecf280dc8d3dda4bec0c2b8c59092a4d0a3789c466
zeef04b0d56405b2f75f7a7c5ebb3fafca4cda3ddf28c95a1d8843e95300a30def2c550b7d4af9d
z69d6fa389584c0dabe7d9d30a0c86620fb96f933767992f4ddfd916433daf33e9c77ff53aa647a
z57fe911160e3b1c19b59eeb547da3bd38e77f38a05e9baee17f634b8912ce2bf1f67ee1ec27177
zfb8ca7f7bc08f6631b56798925e0a7470f2274e75f78280f453ce8f3742d2b00f3155a90d17838
z2f9f2c2183dd4e8ad7398346e91900aaf31ba749e993f5c0e0247ab889bea63ee1b77bc4adfc4b
z4163d04711b17a4f97fd4e93caa44a9d5c380284c1525ba8942cd70ccee54f4668b4d9101ab57a
z3ebca617dc5b9a88be3647e540fdb448ce87e79ebcaa966c7acb0d61b442a706affb0313ffbf7e
z7339580f2d3bcbbf43505741ca7133417a2d44e1cc03498a1f511877adf23d7d224c537d599f65
z588e85d49845df9d47eaf4e4365521982f0451b20619b3ccec103226e2131353a832d8ec06b51c
zca3de2279c649e73cb7c5f49417b3bc9b7189233a3bb40ef5de49be97aa0ca987a80cecfacd3b0
z130e8005a716cb3f1c9b1100e322533d89aa978d79c45f63cb8abb76c775cb05752029bfddcd4f
za8a4a962dcc402d248f0f6a35ff22968450fe37f483a6a757168803d817fa9682b98febf7ecc50
zb5d529ab212d9e367ced113ec0b4be25491efa1ce604c364c46c43a35b60d50a50300a66532b34
z10984a166f8200917779cdb8bdd893e1ea6d8727b185793d26c0fb7771820629eed5c2abef38d0
z129c7868364c9ca9407ee3f30e104e2b2d23d0be7afa59fd21705760f1c17e53723466910f249f
zc68375ff1b18607b29186dfdd793167255f91e741a59adfac8d8c95cc6259c108c81a822a601c4
z338142987bbabf9cb88d05970ef09b1c77314457b7ebc7562d038ba2ab833ed4cca75203877efe
za6bbe3d7bc2b1a4343e220f2c226ebb26fdbe515b02a8d60ff2a7ca08bf2dad4d6fc29c4102e5e
z56aa604e5bcf6bedaa5dcb65541ab3e07255839cb25507335c5606c1e6d50b95a93e00b1eb7aa0
z5bc6866306118af11a0186904f827b3526d8691b6360951e9a33b09e42b5fdbbc6d10bf6e5bcaa
zff9fd4b72d8545ea229de41a8d24915f00f5de330f3a2144a166abd681f2ecd5caac48e764f048
zc16e237979c25a5430758d01d3371ce2aebacd9058f216e3a431e42bb4b106fb807cf138972cbf
z88bf3ea12e4899d4bc8bed33cb02caeef0cf8050b1190094a4299f56ac25dab1a22095ac20681f
z1baaf19466f004002587b6776d9aee6adfa49f7dd5e739a40776320b97e3972d9830c1619ca382
z17c985c231d6e260b6d948ecc42559d4b9bbafb24f200a07cbfac3e36e0784c6027a6103fc8678
z49277d25e0f63e0a9812a77c727627b3228b13be6c9288804568d5cd45cd5b43740b6c51298e3d
z4a490c0ec3f178deaee2212c6730425e325f2a4abdaa5c5b6cac831429c4f94d140634d6c989d7
zcf9890de654548c66417c08a27d327fd2833289e06cfb15903578b85fee0cf2a4da9edf2da8aa5
z87a84f13ed14deaac7ad62aa341435e0a32f8e4043ff96ea250fc20769bad0492b4c49058a2d0e
zaad8ff067f22003b2e71114f552fb5627819713088949eb63bc651b93dc70b1218c1832c83c1aa
zf7ef85ac38026522c4573f89f84e3ea96def1fef8edb5190c7e5d81e623d3daed7c2bee3af5943
z976488961769376afc36372ff10085baabf9b6f7f6c4f2ac06919a63edf974df1c760c56e51f2a
z4acd64f3fb9c9579931f38c0064462390a0de58cfdef745656f4eb6c152af17ea8980a24f8fab3
z0b24390e110931b1cd73100dbb5d6310a3c7f759909cac1700efed68df9876662570036ba97864
z0293f0f1d4163c8739822b741537d7fe49cb5d8a7170306d5074d8f2232e060c44da4b4f6abf10
z7a1cf1cebb64e9a127bc3f60819095cd8dc6cef6712265f9def4b65a2376da96f9669b302b2a05
z4fdce264d74e48c0af36f6a14c3711de730ad28dc0fa177ce25e0abb6642edd8aadccef3090d51
z36295d95b9b25574cd62c5e8de1cd418ffc5e9e48f31d39b13d4522bacb82aedb88980215a048e
z62646de7e4b5396778ef60ed535474b0ded1f75ee40a5a72724d34414f3452c45c0abb04c61f95
ze44844eed075406c0a01d921bbe35ba8e0c21b9152d64a025f3d3facac6fedd15b9734a4e52dd8
z81f8b81d11b25d83b00e5d096de2dead2780bef4657e06934828e36a4e0f977713081c04942229
z6294dac8a884371b8833a9cfc51f21a2b010a30334b762cfa63b565bd2f6b91f6526293e3af17f
zc1c3859a2597a95188e74422fc6fcad5cf7155487dbb8c3236dbe470a7256947d728ccf7f02c6e
z0163dbb10ce7d1b64da0962c96b762110237535145a20b331a3aa77159f379dffd51ab7dc837dc
z10d950e160cddc009cbbf7b67a30d7dbbeadacf90b4a87b4b49def32da74d1b1d85e842e9b579f
z9e9ecb3a78859c3a5d906e2997f41c974dc6cc5fcfb0b9e9db055e4c7571f065007dbf2974cb01
z02fd7f5db9584ce00859af5d17570f07825be29659a1bdd280f4aac3fdc993452fe87d5d01708c
zd635b932c2ebf0646b25d7094a95433fd88bec3fcc7f68032de98d095dd331b1bc5e52e03f8de9
z9f0e09f545b90895bfae4ad973494aa2f4ffcff446e3dff9d1c25879c65ef5786c0074c3d41540
z3b4fb64c29e50d904295f72600252abbf47fd3bfc79c33d66d780e436c2f50680d77e63dcc6bff
zc3c28de2fdbb7ab7c91d633b87a178e7cc9510837a95f5c4ae260e83264dd51e4f3eb83da4e266
z7e81b311ecfd6723dce8f62b3dda3d31e282d7d0eee417a3971005a7841cbb8ef1ae6fc3dab825
zc8a78561e43e179b23b8e10b05581305eeeeab48522df9c4592116f3a70e177f0a45c26e691ae2
z223578245a387e62b906c6c999ca9a01476e2735ab3348fc032f9517502bcfb5101829ee8b4db5
zce24cef6050ef1d7f51c9d5d977442e15f9edf417729b97dcf1eda2764fcddbd6fb69c65ad8cd6
zb0371ec4da0161bf3fb6a8d26696e3edf579995938f2b8a5104b002715f3b0a4eba3af83da01f9
z5cbf14c56c0fba881b0a27b6260c4d0e47899a7a231d27eb7667024ca4733d30078370985b69fc
z7b8018a2b20966821f8f5dc37f1dbbfad580cc2dec38c1e3afd3bc2ca5c33262b0cf88039156eb
ze89e50524d9c3df6031f4f29bbba0cf5d209525ccb76141fa809ea1410cb660a512b0dbe102151
zeb6d47d10b312f9912b322e2abe69138630c4888562fe83a142231fa21bec5ba8524f189dfdfef
z01ab6b5091b95371d0de2e9614eb13c3592edb165c9d95c71602b6ecedac504b7bb8fea95c8eeb
za1f571de68bb80ae3b2c6024b142a022a9e2df55288fbde858642123a157d8bffd961eadf2606f
zfb4ba52221c63e21f9d11947591ff2a34f1515ad9d1779ca076c181752f3620e0cab979b118f00
zdc171624da07b0acb09761466352aa60bb16173b565a976847327a20a64970ac3fc0b14fb969bf
z6af63137b6cb83ad5d6cfac861661cacb8cbe60b0bbf2368409387cc2f21fcc0890d6766bd3878
z42d40835ff7e9fc1be07ef1e3cc037ceac19e408dfbbbb60b62723144c142fd54eb7e4d2bba7b5
z6f7b950990654a471292c6e216929d580c8ab9700cc6480f1d11f09e0975e929700fb5e2097b51
za8e0913ec1e49329dfad58a6579f2b8c541e6d50ad8523cbce74f85a77cab06e3fdbfed3dd7d3e
zcc12b73208ff9310b95a775d4e36afad1ec08e664132464e9d32d0cf41976c419c6c853a913fb1
z1269cf76664fda775e15c82f84df86d632036c106cb98ac6c0e373387e89034af583594ba8e75b
z2d16e239423b0f2062863fb47c918431e3c0cfc39d12790776d372c0032462cd47a0377038ae3b
z2c3a14c2a474714ff54cedc087c996e20167196784fab4b796820a2504227597f11aa50c254a59
zb60347857cd359338e37f1db567688177a64fb04cd607f64e412923e96e76cb29304ea25765173
ze2399e064b508b7247656ee0a8f57e83aa6a043226575baacc73e6d9718a03d294b1899969c1a7
z4f1c4a8398413388179c20772bfd52a0218477ca5c867efbc69c6e4702ba1a92e4d23adbfa96f2
z4939fd738566caf72fffc755081dbd5eab7bd0344d61d16aa423be8b429c75e62b5b3f9c94fa88
z9b51d43a6ab7c0fc8651ede2c267e06374842e50263f9c65916d8b3148630972dacc7b3c495911
z49768e834be519ac47f0dfe849d97d8d127e814fd668f390fdbcdfc27f0839fcd3b09139a105e6
z07a1915289fff68cc9f42da55e4eee9ba100c4e1edbd085fcb25261268c901e73f71637d7253a0
z491eab45f0c21139c71b6e9a8d248a4aed1cf23246aa0e2c437b118b908a143b287d4da112b138
za63fe70ed3a4336678f9241f4696c5ec5e9a816a0fc537684757e9be7d083bda91b93410e0ea47
zbf15b22bcf8c54342735e92b862ea6f0414a9013f2b003710212c5e4b35746aff7eb91912ff8ad
z7212cf013fb9f15f831228103a56da17e5d3ade015c03eed5bcdd3c73a0f678e4fdb9f78f094f3
z5cd42f8f20ee4f485270f1355d29625f0003f23f98b0c13af92238136aeaea598dc9c168eb5fdc
z05685a5c2cd5c637769b6866de0e322c5af3d5c9fb7c72d99e54e597d69b692ddc5fc810566067
z9afc2049b0fab4d20331fb9893d1a6fb5929081c83d45e12d208ee097f2e89775f304584493bfe
zcad368ccdf1d7affebbd8ae44b5bffa741893622d7c30b3aa09464cbd20d04380efc366172ddd5
zbf679805fef8a73a8ba6597c2d35c1e7821dc452ba99a2b5124334395d7cea374986fff54c1fbe
zf63e0cdbf5b457db31dec9d5641566ad03a4514782db7761ffaa72473571befa448dab7a02cd4e
za810e34dbe8fe655eb5e04927bd579948392fb0d50d5adfe99e3d34941fdfaad96d01683e9465d
z61ebb494758d65573d91d56d9f7f93576e7fa99bbbeaa221a57817564adbfb00003d64867f3364
z036f8d2b5a43ad6418a78586129d92c62a2aba16de521ea5c293f058cb05ab89dcc7c2112f2a92
z20af8f09e5988138436ec6d42fcf4fc5b31cea6753e52fd6cae4f0afc2ec3c9fb8f17f803217b2
ze003949938c84add536105fb3237f9deb59e9c1709d00f48f663ce53071f9e96a154a7f5a178e2
zf0ab712bcc8b3322fdc21b79209b40dfb4d7315a7aefa04565581e9cdcc1ac71bd9b3a3d107aef
zfee00edc829e15b866d8a7c92469d6e4eda89edaac8dd488cffe0e0ee3b87fa5bc03ff84bdaaee
z397ca45367468c85667e21fd9f9154c1996f9f3c7b40b8b3af591916fbcc687b393616452f67d2
zbb991c5291fbad33e93fbd59b3a3457f7419b37712a08fa17358a2101e70354d8c8e299d5a80b4
z97a0b6884bef279ca45f590207c9d65febf727d8dba7704bd07a16f67e4d9cfa6a76695bf2cee2
z6ee580ff69d020ed7e723619230562060e894b345faad1b07191d8e670c97c9b989526d6c4f161
zddc5c0fca5a951f54877c2adf294abe0ebbe0fdf6cfbdc6e8ed7163698fff7bb8408a76002070c
zd0c8a928c626f1be61d94ee0dbb07c0d2a46e389fb37524e6eb9d9a58e8269ee491c610f6fd4a9
z36f177f286e2058de75bb7c054e538e7fda940748ae0aacea60b8d59b1ba535256aae3000acf28
z6212ae34a3351a2ef521c543332d808c26b84a1d038e46e605778cfae784ea9378ad57020c56ad
z05785a499f93697c5f4a7cad94e603612656467a0a806ff50c7bb2dad40a438ca7a445c927b256
z6c9a9beb9a00877f1f98fd972c12d47f1a6ef472027b910b3f3bd5c177788535dc8543321533b6
zd8160e2a302ec6f7b8d82aa1214fed10ec75ea170092cfade9ac189b21541a04dc5f2e5d85ed87
zc7e7cc5a3a77bb445ad892d76b759b09880d85bc77af101e4bf0dc46c9d4f098f60aba62388252
zf91238d13a31b9d8ad1aef366e335f3b52046a6d9799a6d45f8c6edc94abe3b0755365f1850a88
z9a4151bd335fa9dc9c7a85f50bb962b58aac90d29104dac85d1f09e9dcc9d7321bce7f68e0e53d
zbd5ac3deeb1f46440f27e11058c9ba98691f5c9b1ec0e27e0387d514ddebc104439e5eea30657e
z4006e6749c997921bb6fbbc052b63f34ec74576d88f6e3e3d19808f24703e94b08401a71e05dec
z1348e849b97ff5019d56fecd80534e14c61837e656d26804b5135144a46c21e5ff6daeedec35c3
zf2e7d501626baa2dce9b159cc874609254bd759fbef76f708dc95c8dd7027086119f8f552e7b98
z6fab8cd5c02a075a797d3af34f64681007da570be4477119e1ba49a721aea552a5d8dc17793f33
z0982a5858c5bfe01951328eac328ee05bcaef810dab5dadc5ae2153790477dbb6c378e82c9f622
z026f132a2c5cc1a32c60f4358be1d7f0b6ba578f78cef8ac0496082c8964a58ada722320c1faae
zd0fe13c5c9890fbc9cfa8ff83fc9777df3d425a844ecebab1e25efd2a7cc6817e579d56f5ae467
z070221c8297ba3b8d89bf9a89ab5ce08b8c708aa9c0e239a17e92679f089f180d2701acf7ba076
za7df58a9777e7a7b8101a1ea070f620035bd6179bf33b4fe760ba51bde52bd78ff7e7889a3bced
z55ff5f7936152be5d22167e5698b6019eed49d94de1f70d2b82da68a18355d0df1f6d15bd8ffcb
z2676281453aed0e5c3b8dc81166d136f62439c6e2f977c9965416970492d53d5211599ab33f4e6
z86329e0fcc85d1009ee73932017fda81e92088786a99d78a7f3ab21d6f72329a58df02230b1020
z61e560a4e3f16d8d7ea613ee87c9bad72b2adb76bd3dd513eb776ca0f161b13f8b80154106c1d3
z3a57a7a7638c7cdabcf0462a661f8ed729140c3d24b72e4510e78c3702c574d36f1d6eb3066f74
z074b5782b4d0c94bcc19c020f555576b3f273b0c225eddaf4b038e1939f5c68b007d90b68b7c82
zf6c715c53e689e457793f45f9ab50049610215980460040ebd7cb459cdcba4c9776538b9c3b6ba
za3d56078860c2010251b4cbdffc0162c6a6a24a0c68940afac2f8c179efc1829565cd008e10aa7
zc269a6cbd9e4a6a0eea37a26530226ba171169576b4da5a325f143a3687b491f9e86bf17af8541
zc8a2273c4a702c7e33888a647fe587f291c00123e5b863b09132db3d9a2d7ed931adfbd49d57c1
z5bd7c323c2740c0cda8861c126de98f4ebcf0790933e0e0c9ca49575b8824847ad6dd29f6b88c0
z1f885052e654a23a7eb32214115365cf6d131e45e659c200d1a03901d7707a1f174a69e8624ff1
z8d0e0ea9b0486e7ae2cfe2c747c3d391fd18f96e483d563ffccd2ec903d0c283b869be2a0aa46f
zba04907f1ff82681cb5ed7d9703091ea422e8e03086f3258cf54fd4f696568b2b5894d10acee4d
z5d55e2595f43b87f810152b34921dbd527e29b6e9fd03e60ec2e8b6e25ec969b21b6630f2b9ced
z649152ab52012e17376469f328c60bfd1175f304f5bfe987fdf4e6edbcef601ba6b8a99528e7ce
z4fa652b8caca2e24986b1675d056d749b2b53b2bada648abb6a60cb0d3f23566816c0ca03b59f1
z016ef3d84e0891b674f76bc2a6941dc962873db0c87939a143dafe8b43974ed26d1bd16ebee77a
z2449a019c1d51a64254b230841402f51f3c1f3e8cab32bc4ff2d4e3b38f2cdb8469c49c8cf9e2b
z52756b3c28bd1f8388938dfbf64204ef7d40ad83366daac7925b70888a3ae7509e18dcdc96c391
zc522fcdb8048eada482578d7d7c68837b9018adaf462a8ed6ee0f21690fe80c9b3a0e2a2ec6915
zde8a0de1a6043980711e0607342a5386e7dcee10cc3059f49bc6ac55b173d14d56c776658712db
z3fdca7c3fabb984a2c971a1bab7a2930e13345e3cb951ab2beeb63f5b850635b6df34a52ac1115
zb6b507b4a3d04aa5585237bfb48f6fd2eeac3454850f8243cf46e8fe2134f072dcd1430004491b
ze1dd7c47ee76ce7224c2b3595821c45dee5081917168157d66ad0a8163383bffd8bd87065e9b7b
z4644a94e91493593090460114792581295c3db51b953696a167f4ad933414a8ad29d60c9ff2ffe
zaa8cc250e9609a0aa99a1caa2daa094b34e8f1af873ab2fa25a96c95f99ef9d99f9bc9f0615f38
z663c5089c1dd1e1edc3a7d08c1c9c57f11f83169392bd50017db0fbaf73c307a359d9a9e165207
z9cd8041b101a94f24cfa8a9eecc6be36a498410d065ec0f8aee47fa1ae38dc214bad2dcc10a8ba
z828638e7060db0950f6a61a9f381b450cbee747677c913c76de428191a08e6015e862f9839eb6e
za1dc4f883b4fe94fadb10a1ec9faf19c9566f0d303e6d740e1d60dca06f4aa30596ba8bc44c7b4
z13c40db2ece05171eb9f11de1353b1b1d11173e9147b1aef7b4738643cab01d1b77739674bbbb8
ze6e3b6904a3e388b876dc8733fdc31be58409cd807f80762514e1adeb543d16a58e10b7b369bf3
zb0b955aefada61feedf807e74aac7995b61e82800cd22f596b531430e9e44d8670123a2de25a03
z48026627baf33acbf69c8d20b1e2255509605187a25bacd530faf6ff366ce8d22fab1614bd0aa1
z5792c1c9d4ae5f9f2ee9c55ba6fc74b4c9dfe45962309a3bb5e0af95612dfa3c9177dcd1151c92
zf9fdc1a6fb99e61e384f5badb6f0df459031ec3361aa3119cc009c9f0ef6cc996d6b0e0eac2cb1
z2393718726d62db48206d0ca01acf96e183fe9d9f4fdfcc3c6e2059390224dcd93094f54fc4318
zb199f900dfc1d525e9e108df1cb008d161ae2d766c6ad88309d1f0b11ccb47207d57234222af5d
zde163db32bcdfff9a27e31f426bfda10d0714c67129f84980095f58406dfc9ff028578d05b3d54
zdade971e36da506b5b3a8a0469559c92894734439203a39caa23733fd2cfee7784152e7f74c46a
z81d00f6c67df1b6e4401baac49c997dee19850233607cb8af9f27d2a938384b5c900fb5a407c42
z84b109a30021f0e4d7329212c18428f5ad5bb21e6f4cdc46b52a9d8f2a394e6222d9db40a17d83
z478b362e0344700b7eeb1f65156f3c8d76c87961ff6e1f97f1a753dec07a17df659982f67937b9
z12ebceb7b9f968a7e40b1eabcec830af87a02b20f338f0d000ddad0856e5d56250bead23382122
zc017c74f936316e47bf86b7af504387e4ffad989fb286cb75508b60206c3459aaeda14c34f5a11
z479f80caf342c662a868ad27b7a089b1aae5bf0ecd84b7335ccf6813bfee95f8fd8a63ba3bd277
za9e30f1df9ad9b8c57bbc98d9e0244c1c64a1e02fee04d5c0f4e876d4268f5769b448846b73bc0
z8b5351adb1881bb163c89bf1cb2828764fcd74f1c224b54ff7465dde4e1d3c4f2153437ab72e52
zd7105a417d3299f18700d6e479e00c77b71de3236e3dc908a66d1fd81eefd02ad423418d4f8ac9
z0c896493ab5002ec6a5d22849ce6eb5c21c589c7a4c95fc0b2dbfbb4b6b90887745ebb4a2f2d83
za739dfa62485fc071e55c610bdee7219001fbf96a6d9e958af44befa50ed1af6404f02a541c67d
z5a58888e4972939acb95add6f641854c3792fa56fd06714d402237962911ddedb04526ea18192f
z569ec3dc7d90c58ee502b30107e69562355e2be7c8a83b35a2292544845e3f52ce440712fa5ad5
z54ed13d4b49eb1784475a55b5f7b7a8f40527f751f1e1655b54e15b8d4ee1fd2ba07953610198a
z41b66aa69a22f78fc11bfda451e9ac191e3a4401422364b553ed77c4051621d4d392244447e548
zab3e471d8b2aa0b9c95aef3ac5c41b18689376f907c55b8dd277dd2c9ad0cde3813491ce789ac0
z8e0ee77f4a0f20bba493adc774078f398b1add176fe0a5f917d6f87dc0cf4caa3801d65ab619cb
z278c3fa3a89e565ac37b3594268b04c8fedd1cb01ec393c4a52d1b9e8975ad4685daaa140fd090
z33b55d516b96807be091a90b8b36cf6b188a33e8cea6ea2dc2252566d44f66ea81c85a39cebb55
z968cebb9c73f964d3bef10c58ee9ce5b163126dc2895a13e16620cede53c8631b3958a6a635946
z54229c32cbe2384b038a5b3709abb31d2fd310c7778eb358cebc9f9098d7c0139d1c701f684493
z67e4c3ef9816f1cf0a5d707d1e4937e07ec6f2c71e5cabcece9a403c496f7a21cc97d7cfb07ffc
z4d9d3278c537188b433133cfd78a350de8fbfc2d91c7d5917a76e4cf39a59663bfe30ea88e99be
z35a426a21525db862afc46345e4e1d8e94c9d9d76a014724caceae4af394bc7e3f09e5248b1d5e
z0d971d034c682464975d16b18a90af832c654d75706644ab6c664a4c22cb05556b6428685adba8
z46be732a8efbf36a6aa09156162bce95ec8a1c22904d79df90d6ab73e36bf04c9a5c9131163c28
z7c82b6f6491d486de8b5f99db915483e4c339ad540d0bb73ec06cc75212233d3b5a659aae75d93
zb6dc610f7ea98c576970469e5b4547bd03b760eb12ce0215cf782a656eeb80de44d3e3b468787b
zd752a9247b3ab17c4fd27964aa4f1ea2027e7973088de4158764a7728fd73e69beb82dc523f4ca
z4a9f1f1091355eb1c5c1743ac1e5c2112f73ecc17f4499024e8963e9918eacc97744a4974b4356
z81f22a19a486ac461298f0998edca4f2f1af65aa85c75cbcd7dcaa14d0de407b667195f61bcb64
zfc41d8331f4afaff590107ea5e5610028c88f6fc10a4f33d5ac2d3910eb839089f8a918ad3d43d
z499ff6d362095e9604388d9ae68daf658f5046a3c8c987a6ccd471521eddac7f5267d588562451
zbad37dc4e89565b3c623f4e4f2b31713e9c201c09c4ae0ec5036ea5e3d3e98d894200c7be0ae94
z9cc2f996381bc03af1a34b975903067a7151c5b508259a23344c315f335b3d19deef11ddd97487
ze45318a9148504a3fedcd8e622e620f2dd54bd0c6e8197535c676ac9122d9ef6815b0b9d46a244
zc04246d58ff1eac0f88c9609cecd94ddc27fc735db53c2902f1b7149cdf1b8d403e70196d20751
za8b512250ea66a47e3a3d15d2f8cf6cabf2a848972672b139694124d671e53a7ce69b417643d56
zb74ab777596c901c2e846b5ba54be6066b30de22be7f95a692babdcfcbe83e7eab36bac1b8ec6f
z349e86ce7c240c8f545fe3eaee17b310b58e4c1c955da31d8261796ec84ce498f795df5b998258
z43c0da458a2ffae845df683ec4c8ddc4c29d5b13d2f96edacd630a83ecb304543c83e27ca4c8a4
z42eb0b6e6042eb4663635b30600078143ffa421a5d74f9165526bbeaabd941bb20032764718bd6
zd117881cd6a0981198320f8566e4134505309708e95fa15bac7b2ceda4c259463f75ebffdd3254
z1b86e908bd2e5200295b2e89d65fe0b7e4ec97cb57692959cece6c3b7ddf92c7d7d6a81c66554b
z63f22fe6dff162448c8ef0e4bfb8efe88304141fcbf2cc7bae0d4789e489acfdd19c63c41fe68d
z76d6eb1a50a3d3ae73f4279ed7170ea4f1baa0acc8b02777ea0dc806f386e1c09ce965f05e50e1
z82d71b5bf2859491019296d1c94e9357cbf0b6b6b3674ee9d25866783c2f5ee2a0595104690ceb
z57b555dd3493101d59f6c78ef6f9d4b73194e53f033b63796b67ad3f0e6e60d169e2be7a8c4377
z0bd64abe8e4c8409ca6cc5b73c0dec883a2825b92d7539f12f44016b3d7634782592db8682ff8f
z3e79203f55b85cdc3d9952a5d6e399631d521908fab87835d4f1e3de35d18a1c60a5acadd59d92
zd640847620ef133055b5bd4ee7eda07d62efdf736201823a5565fd599ff4d261acb6ddfb99f67d
z634f62a8af41d8862774a5561a5d3cee7b25f0a1a481b1217a9fd4c64154c28531dd12df1847af
z66c42bff9f8ca57d21430bee92cbd195c86d2167269ded6eea2911691c8899396a44b9c84f25a7
z57fbc8c51c3ddd58c62cfecc94e7a03744009c0f58d56e9643d7327b5dce20bd73e431b384c604
z90b065d36a23a88181ca9f11e6369e452ff6d2b1eefda4023537661c692f551ff1ef8fe3d9f4f3
zeee9ac6eed0b1e2da33904673ec2f08e416301174d3c1545298b83ce0bd7554461c0415bbdf290
ze50d55c61853da79267c1b45b4c493b2b6db4ea3d396cc802a8bcbd30ce3f1b7316c8d8daaf452
z37ddbab388e4cbecc7a65a69567a09367a283bb4edcb318411bf8a2b3df774609d2e47a23cc75b
z9772facfa1ae70bf5801799284f4d23fbc09434e48494488e99ef62683289cfc8e216665006ff2
z3bc9995c18728562fa9ecf1e8ec4ab3e479a3f1aa0f34d1f05175c457f4ec981050fdf2e3cb6c5
z36aa8dd3257e0c1f67f1e4f5d31c26c645cec05e796bb508b1b0a31e4896e7a7d803ebb34d04df
zadea46b2077abcca9b59d205600ec3e0c8c9ef18d55bbad44eb88d9a6450505bd6aa0df64cac0f
z0bf23bba2cb1c501ac74075c540a9e8d12ee86ee6868b00cf0ba9aadbe42c16959e766c49350a3
z0156911be9686b0f530651edc0c9ceff3ba3432399a0ce2420f0f5750ce0d06c23b2c8886dda51
zb1f5f4328302ce130a8890d0a7d8fd0a55dfde850b781b4404f6035d9048cc7b2e13c5a1b8d8f3
z8e478f36491d72e32b1e0447a81eed925729b355139d9a85f8013bc9908843707ff8eb8f24cd79
za76ce41de225548b95542a307ba6f7281656deea5593456f543fba195e7558231cfd221a9053ae
z0c64333577529b114b3eeb2a5851e76bb5956531b751da4746971c249ca6aeca3fff544cbf5769
z4a955faa418e905ecdc9f222b19141f176576f75c046179abe3951e693a4e3afc476e94bb596cc
z6976fe44c93fb99e9e9e432cb989bd332ad4bf22959c763ac73ad53cebd1ee3be444de11fb0cf2
zd0cef44c4e091a395a9ee69aa6ae7ba07bdd38371424c1a72ab6311790db8d8871e9659955f5d8
zeab3d803713e24d16405ff39219508a5584c37089c7840887c04907ed53df052ef45235c40963b
zae62373cfcd4064dd93182e435cbcecefe266df800fd88c3ab406f042ad5d5d8cba321b3f5f41b
za990de00ed3f010f90d7fa2bc9fc8958a346b92992301d708489a460b4d33d7a3f7420a5b69aa0
z5639ef5c199d31efed1f8179db64057c1575a0a6d3aa6925db92283fff5601c78498ed661a863b
z00696517e7e1b7e1edf09cc38f20300c174e4482e9b1575952608e27e035740180bf0469c790da
ze91d53a12ee1b36b834bddb4b8df84d66050cb3ca662040cd9a0532069dc4a1d8f20ec5de20211
z2424b1846952e04915ef1d9e51ae4c565fc70ed557bc1c88f4c456bd6c39ef50853b8f09831e18
zb01ff72aa0d838ed88f67da8ce5e999ca277f31b503702d1fe710d9261f76ad6246f735ab58091
z2cccf2547a96acea13d4241bf2375721e853cfc8f38a211ce54c226f9fbe6bdc3cc10eb57e7265
z788a7d7536916a4ce9529f42ced8ce880531d0c81534fb2401b2ea2ac7b45088c50ca4ea1098c1
z475d2863833c3716ca9656d2e26537b3c8a54c736eb3ecb35f15c9ae24ef45cdc0c3a28aa8a0b3
z9eaec454ec713c2c15b53d2761bbc5f35008449fdaa3981f3be97b7b01aff52941197b355733ab
z869968a660e5591d5fddf26bf03bacc292c682651a4d22b1cc3baf134e3bde88cfd60a5c63a383
z5a6691614d9abc1e2f18e92eaa484cd5d98b4c5648b6fa0e8e476514815e846334fc02480db91a
z09512a19aa928a885963b9f859b43ea2f60bb60d21734248fd114ec2a0c2c78a9332d36aafbd0e
z6da7d3b28c4126ba694ca5c6e9d20ea670e36e0d54f7dd19cf8e6f0654218a348a9c5982171516
z61800f5581683a54a25590551a0c7d87add8542005e767716063e4d8ec9b25a7fdbca2ddc26d5d
zae62231a1f4112f41b0cf5604c8e93b58483d2afc3f04706122c23a81879a58fbbdd0bda2a6e95
z3b8ac99ab3d62260ef275aa795a401ff2bcda105b84903dbc44201a2f1574b33f53ec240a837c0
z4a882b255270d4a0d54c177d33735f4e541349e9c9b4da3f5506510a179937685b9ade50e35c83
z6e07bfeb4f15d77be1d0de0f64b34859273dee73da36ed84335c42a44a5f60bbfdc40c9f3bf2d8
z2992509799b2a4a91f3a66c827d9c7b2db6927012889c6edfafdfaad289c0f737d21dafa1846ab
z4aa283efb8cc6ee8cc47ab79674a498e2c141d03cf2cbe53d7c5b17e001f3c70127fe41bfae49d
z8428d4c5e829fb7579cf5f56510de978af5fc3578f4ec30369087a35d0cdd31eeda20568d0ae21
ze321a93aaf681a819a87b970c898f6d894d3379e9ac3dfb58dcbadbbb1438acc533c0458777107
zaf54ff6e05391851341b1abc323c85c91f841e7147ab646ec70fd6231ada06c35f7a12e3443f03
z786bdc3f81655b3350a71c2aff34b081b987711aafb87b7d9240453a0351b95a5659ce3d9b84ba
z5495d4bc2147d77dc8c768e22f54a319e363831470ae8c3b5429fae5e998a69d31894a2e8f404b
z8a91daa5adeb1916dec88779c2bfcde4a5f39f64d135fad1d82a5aaef5d4413234102a757e8244
z52bf8eee071bb7097f88de3d2baa6e03126e330bcf55a36d8836119ce2a5d43126b793c4829146
z4c192ae0f8a93e0595c2d117398a8bc0d061b00add8fc803ebe635ba225813abdb51572b54fd53
z916f20e3e0cc3bd426aa4f419a248008e9170aa0ef623f9b418566ca69b66ea2fc7fe555097ac4
z205bdb363f3bde5b2370e36b120c3a69c2b33033c957fe62ad2fc467038553455be0fe4018975f
z24eafaf77d53400e2725c03108b9aac5c2840ea2e84990762cb9e08c0310b965ae4d06fbadf924
z07f058a25bf697bb0f03fc027de6bca8f77b9d818e9469f8c10760faf733a1f0aa5ff9b75a601c
z5094618bbfd81dd305ed323696def7a258c7a8958ab5dcee6d926ca871c45515548b261dcbd40b
z9ff4983611d67ebe0a920b0e8b36114dbac2b2742af32bf3670d52d4c44b25d052bef305e55bb4
zf92c724686f9f0773859936f6f13b964e8c28a8104c8a26368befc00cb911dddc4fe413a8899bf
z30caf6f4927455bfc50d627b160d7ffbe0d934943305cd1f74d1ca00e3ce4a9a87abcead5ebb25
zb987fdde59e54b3c4736c5af02d12ba64418aa230df00440e4ab99ebd0eb1ad39e6e01e7408b63
zd8bc6970c67363c83f6d0e7e656fa0dba879d954aeb60f2257f2d9b3617546c6f2de51c5c1f3a9
z0789c46661fa2b4ad99dfea196ba5f964aa0f3a5d9444e269e7c901bb530059457fc8c8237dc0e
z08349cd9d709818cdef61809566cdce98d17d7959225309af8c17eb2c40881e2d55384eaa43349
za948aba9a4be3f9aa69f80b963c06d862aa190135ad1873973e12d7fa3d43e1899ef7ee31b57cb
zfb706865681fb5f6a02248cbb0b1ff2c98afbbb40daccf970bf6750e40ce7f9e97d73cdffdcefe
za0a812cc47c9391164dc1c9ce438a6c574dcef6a932c73a8af21ff06fc13e863cadf475cfcc8a4
z274b866e287405c50dbbbae6f44807d8c4c997d76c97379a4a8e330ce7f2711348580db8edbddd
z808e88312a703a31d30429b29d4ec745416159c309f3f011e58215915a80c1363f53e8e1784456
ze690a47973cb18ee8153aa6824978fc7752add86faec095c4c298303d219a9862ff8999a9bdbd7
zd1ddf756403cb90f49fb9d837027129f429cd65eae1e25cd2b5d872295e507d034ca7ecd13398d
zd3c53f38dfe7166e05849f817aa00e303f52405f2df99bb276bed7fd07c796185626dbb19cd816
z87d7a35c3e79da093df2484baa084cd68543e4d7b89ffd4679be4c2e4318654fd82271c310d7ad
z6d5af9a22a72b869f1eb8f8fbaa20eec4a2e33b271d61e3a9aaa633a789cdf5032e3a651829ff1
z4d48eb5b458b2a64e9d4ab061b8434dfbcaf5affe5df2256a5c4aeeb484725a7fbbe91fc85bf73
zb21a7447514a82953da77b04f3748d74a8eb025ec964f393a38d9e61b19242184a140888c208d1
zb20fff8dfdd698f9320d7ae4c902cadab0cb2cca1a3b624ce4168f14b1fa902fd7746910a05c99
zab115c669ec6272fb43072ce50a3c3c5ae21dc8b7caec0bc3c6200404450cbf2d5fe319055b90f
zffde7d8034651e4ed320ebbff0cc7bb42c28976a190d590f698f40206a7b365f8098a2d6620e2a
z840659c513e920d1d72d7e83806c784344d64e01cc1a78785fb9b1c57dc0ad06908c658c03e7d8
zf25274fe924b5c4577ee1d5d224152329cc13ee84abfda72f17126cd9aa195bfa875562161ddfb
z24a28f16375112abf91999b17c946e4ee94143d7bd334c879109ab72a58f5cb785b8b8390f1f2f
z24a468b37810f3590e5e63e84a687ae37b765de253da5ce74c5359826895adbf446d33e95ca98a
zceda818161bf111437bc9225551cd59e013e4ca2ad4a86b88059760aea867854314c3c48eeb919
zaad5acc090daab11c0ff365f0416deb5bb1c36c57c8fd18ab04551a29fa9da2f9991e21f7c5b3e
zb37e2921e2c616e3a2ead7b64f16f1e00ec0e3ce3b4b074c4c5037dc4efe52413ed49dbf8f1043
zc3cc7b60b02cef264e27b1d4d7cc803654355619b881867de9d3c0b8c82bde15323e4f1258182c
z9375fd34a53c2a8d9641d0400d7b882fe6a11eb3879f9c18daebf9e0098d9e7923ea383d5d3182
zcecfdc10d6abbd4238a47da6462d66231f405adec3bb47bd0fff99a90d6a6f4c9bf93e063dd75e
z234b5506aa828e2e7d351867ccd172c80fe325a5d98747ca696b944e05ee190f88cf3c06e1fa3d
z770188993d90376085f6c01201565a375e21a569014dae44da7dd4fc63e455255ec088e1ce74da
zf81953a0c9a6e20b0fc8d2aa232167be64da89b2218a4f7fb091d0ba59f8e8037957b6c51273dc
zd9fdcab20feef64abb6911924ab7204457532508f44ae8d1abf751a0cc230c998207b68f58c3f2
zcc52d46f30e0c579ff635b26fcd70959e4d5cad5cbd8f3092bc997ac835d00aae0bdb5a865e870
z79026eef881753a425a1545a344de60cfe1be8b8d87f643a91bd3d77d767138ac8dbae30ad75e2
zbb87ca657701a894f9e21aefe08921475d6e8c3676372c8e5a17dfdecd74bc85da14a8ac55c8c0
zdef675c2af0adbc8a5a0994c5ce8c4032b308480c36592b6efd4326a612365369e3be5a2a293c0
z1bf1b1f63e7f27e45ba2011849fafd4e53f580bfe3cd740a4dafa2f96d077d68b32907e78355e7
zbed30ca5ee8824e872541c8594132f5df2f53d23d02f85a5c3fd41c9b7066f3763a2e1a86977bb
zed6b41517c1bf2b53c2a4ef05ec23c85cb67ef4b12972b2dd539d7ce6d9b11fec836464f4f1a40
z69fe91aecc693f816da479d185724201bb18ac8c6567c7bf79f3b520d883ec4be6b96a47b08bda
zb32773bc2b2081547d238fcd3368a5d4f7744b45c5298ebfa4aa1618c4105a12c00f6d55aa5dcf
ze5914191b64e90b255953573490a84c3780ed9b1f77a902dae54bbc4247cbbb2b724d22f8134c8
z46b830fea7b2bebdc9868aeccb998894f337da54a44eb3abdeb1181db7803f95713e8df017ebc4
zdac08402ae99640bc8af2965300647254d43298e6c70254f551bd12fb37d7a7513d6e76a15a89d
z3521c0517419ca66455c30c44dbc3ab8d999c830e1872d712542ebb28539482cd73d4f2ed700b3
z318e57f0a6d7d395182680ec5d5bb4f73575e981e0d942a4260bb0e8860bdcdf8625d1fdc31afe
zc698e38a9c701d915e5b9b37e92235e787d8bb23c4503bc40f122336cbdd96a40b733ad8b31d9f
z93a828c90ebf4743a61899843f13ff98b11f66ad5e5f856eaf44e9a9e0812fd62982fa4ee03d39
zec157c03187f74762929d4666f5cd71b4903dfb31c9e2870d8633b529da74af0a1d34af1904c95
zee3cd65304af388501979a0b2ff898fedec2affa9201cbd9ced67cc60103a11827ae90f056116a
zc72e4a61af0acb0149ff1468b04db85f99c440e74facb616baff42f2bc46cda995d7cb215b5dca
z502212e6c98bcd7983e589ecfcc90cfc5405d410c42b7180b11f18245970a8e56573ed8a21a089
z3d84eb90042abf3ad7dc4eb740a70b27a2410f95696d62a7a0478ac97e5f727d7381514c2f35ed
zb9fe6e867874525927901a236d2d6ecfcf523262c4cdc036797853907dabbe4b8745d7310b2e44
zeac0b7ff9fc30a9c0dea6a5bf331ad123045e94b8c086cb0324d9c6d5ce13f9c0bd821def399ef
z77e6636f697f9130e800819f2c8bdb183df2099585389b2a1c7c899ad3f885f0567273f2271cf2
zacf3652aa196f1215a37e7293e2ccee56fa5aade7be5c917a5cdfdc4da12e237e26f71c2ce92f2
z925bdcb49892aa605fa968b2d864bac040a625b0f64f0a62c8830ce760cb736eefc14a74894e09
z13c4660be4d836a403170ad0deec6dda4731670796c87437973e1db65c92f8cd08b886435ff4f3
z5ff4bae2ac9348a06dde20450789ca76eb3ed8ab12e5ecc639d3653b1548f04f6a0108768a0b19
z84ecd8be51ea8e1db32564ff21b9ec2c80856fb875d3e5e2a33109f87116ded0d38b38bed79802
z4f661fdb9c07db901de1797da251c849a14615042806e27ad51e3bb6783e920b22fc0652de5d51
zea975abc28b2ec0318e74f9dda9377cd0c9504def3b94b6c92ddf4747035e76e18ae51473ce643
zc17f0f96ffb54915d02787b77a785d4b862d192455eb6fdaffcba1aa412b4ca2ef0cc1e7e75b7e
z31f39fffb56b90096ad44d70c318ada95de09d14b173423fa8d56661da6966ad63eb02e81a3b1d
za5a2ae0de4dd53e3e617bdc2b1c9594f05def57d01e42c5780674c6071bf5b801b8b4858afec31
zbfb4348089327c9fb36c127bba686118a39c00fe4d500dce0383943ca31895932b0ab4a01067de
za996361cd00ff5e4bc2e97ee7ccda01987679506a4af70ca03f95622c7d84c7cf77f6b52e048be
zdfe4bdfc87eb3e00697cbe82143d96b28afe2a5dd4d58aa5b99b3b9169a5babce06fae6c685cf8
z94c228b60e1e26306542a476a776bee39f52a224e640289e722ed59c9f60dfb617bd195c9b2331
zcba46e19116f5cd8458deb3bdc892f57aff0e9cdd68a87e3ecc2c58ffa22555bd087b1e0030007
zfa00853722cfbc28d9fd50867f2c1a7c3ae2dbe7d546b00a67dfa5a1eba6a414acd2f4ded45b9f
z3047576a6b339d088ddd7e6c8c34dfd9a00d8c83d6ae8728f8a82f84c86134a6e277863df6ce63
z64fa8dbd190feffe4951e06021f267408c7b4c179bc0a9d09753f557f4a115f3dd5fd624fd3f14
z68ecaa74c10ce949da3fe66f61b3430244c6a80bcf5d0cfcf5b6e84c782218cccbf873b0fb6c2b
z2dd99d5603132bad7be689fb443eedc55651ce2fc86eeb4aa4712c047718dcad47d4eddc40cefe
z7dfeb1c7e1b3dc4de44cc9c450164ebb4d64b1e27178688dd09f07b16dda53d9fad99aa89ac28a
z9e82ffeba85dc3defdb58680c7087b7d88ede8e8d1e3b9338df8e89708b3c93baf882f57088c62
z6ac40eafc6c119afc54f840b7bf22f1151454a2e62e7ad14aec672825dc030cbf567ab8da2506a
z2c693f2d36d1e906292dea313e116e99eaf4b8dd9e353c95818b038a94e44689a6df91a855cffc
z5a6c73c138326cdc370531cc91f7b3abdf87c11bab58d879ece11f6a728b4e1c9ae69c7b2c38a8
z1e21a79471eb3d7fd9a1ae79cd4943b61ae0672f2ac2d5bc47dcab46a6d8093f47a3280668245c
zee99235a72657cc88ab67f892afba64e492f8c196822056747741c228016a712b0889748ad1b63
z34b4543b3b4b86da183081c10c80028562041849414c92acc3765aecd1563e5862008778d73fcd
z1db3da97df8ba7854eccf8f1d249271f44073c1e4a6e2b94a3b1bb6213317745317e4efee807e1
z65130e82e2efe3a4bf563dbb4e7d419632803ba45400c7f3ed1ef35ab6c5b8455c079ddfca7b5d
z90aad5a54ec641e6a9c4ab4cde9f12a5ae0e1da33fd6f7d6375b439a9d331a15656fc5e53be294
z8fb877ae893030e2d20e2607e3130659d7011ab9cb376ac9c721223dbb0a549eeb9c12f4c7b1c9
z4ac1deba2135901ec76f75597630878067b2ab9c80fcc6977317a95ecb67b8e643d2ff75125376
z2cc8de02b37cb8139cd96fcdfdb508913251864e477f7868d14bcf819c08581e074e96d626f09b
z88ca96794e606b3d6fd1c301bfdbe2fc0924e21b76517c9d1f9cb4d5a66d28d702ddc4cf341f22
z44b0f2cf554cc3861c0e0f6ea4e5b0a1c6799cba70c2e6be9b0e7580225d38f17a4ec9a49306e9
z9aac9d98f7bf5d26b00e594fbe7d11e8e3388fe4e891cbe9e57d2dd272c660edc0d65ecfa2523f
zbfddb1a30509a8067bd300f65e674c54ab8c7a10913ecec7e8bceec239901a3d3a3bc22586e071
z0772bb352691c322076c054d9b1c090bcc10e927180e4ce561702117fd7a7d560aac40c960714f
z43dc53427e436b2dd19acf087c528f8e3fd232736adac26b3f8774e61494d206ea323b9f6fa148
zb7595489b3ba472ac8f1a22f06ccd680fd2f04c30733a1fbd24aeaa72cabe64b66326f8b4e102a
z36418885d40b45ae50d213c95f854136b96cf30b176a4941e347c513d8705533a7c7627308d233
z9f263e6b99a22aa7cdd8a5928fb2171302c60632c5de3b43a91162bd3cd8cc1fd2078aff31942f
zcadc2c0dfc834626bd5d1b065af80b554dee4bdaf40879b42b448d2f04a8495ee3199406061d76
za0b25a4ac75a699741f6eb13072d9f53ce3f78d36b519ce75e26a6c24251d34203b9fad1165317
z9294c845caa542d5414349548f3595735137ff404500966a789a7ebc2b4824e6f402ee6215daef
zccec9682c37bc337b50599a07d9c3e98fe8b7a9bfd07483b74058470fd77890c8dca41531cf83f
z22137f99edafc4ffde653283f34a2dfe82de779ad90bb81102304fe58cf0511399595112e91e6b
zdc39c701dfdd8c3adb9d57b01976919577c3dd828b451ebcaa2edf9597ec1ec1b03cf96eeac78f
z2e9b83c89fe7f9cd9014bacd16c0b09224a3c86ce8eccdc3d9836d3cec60226e3df90446ba487a
z7ac943254ab35e4ac904f196e5683e39187402dae95ecbd9e5dba94310aa049bad8c7fe6b63523
z31506d757fca5440fd3d6b861a1b849fbff34a7c2b18c19daf43e6035fdeee4cb20da81885f3ff
zab6195c8552520e46276ba48e69a5b2bd2c8c3cc691544d2eaeee73a60e35fb3e59320431af72c
z2b1433f5da85ef8fc4499c1d0ecc6687e248e43573d56c310a8a093c9fee541f3737124f1ede8b
z71e6ba7e39eefba3cfd0df733b133552685f290f437ab957c591b9b85725ef4e7ebd36132e4c70
zca6e4baaea7a7b7980950f19616af595c8a5197d61cd4d33f89224eab2a0b0f77a38c33a5ae2f7
zf33dbdc43257d2ad842b482d2ec9696405e55801bfa5a518daa2616dc766e9524040498036e1d0
z4636f9be44d58fbdffc7b41db597dc840c430ce120b1b25c60c3d2febf78a873afbf5d86a8dd9a
zc67740203c609faa2a7faa496274cd4f68cd8f1e4c7b5bd3c57aafd18b96614c8de7f83d5e1be6
zfbdc19512ecc733dbad4061264ce012346628c4f4dd0ea0a610ce5880552cfd4483216e17b506e
z01e459fd4032c6860564a62bf4539f84e35a23daec35ab6ebb8d7eebd034e69f1dfefdbd13e094
z0361612f257541f5359ce20bd58ea2a8c9ed4a88c5c373d8ebaf4601e641e026ae214bbd9e046f
z75c72a5a3adc1f481a48037a603c0828797a1c8e1198a37a42195a5d5af2d8d5f12d97845a4a25
z65d5dec1947de729e36daeb7e72d66631747ab147929af99b41e81e03f09c9f26af8217639b490
z003e98ea7d5024f34a6773bba09cfadc33878b82cb9a1690f72a5230744677c6dd6ca651eaa05e
z9c25fc798a8a2817cb69c04318bf148cdcfe23ee4e25f8bafebb2232a6c7c3ba921eba6e4b5df0
zc6532f785bb119739318dbbe7f7a737254894980406e8b6bc96b7e503303418ccdac7ad5353667
za55688f70b7f6c3c10302b7e16949bd1e23b852e2535b1e8c8c0604e071d38d72ead644d56b951
z992e182bb499d6cc869a25b390690534423d9ef1b6b564edec5712217d1494593d7f10e4938538
z4d30c8c4111fcd9d9e34f2c9f32a858933a68a51b3a76248d4a2327b6600c5412e1b55b4c8f4ca
z9312bb41954dbaeb3424596510fad57070462c057c7c7b68e32fa1a80a9282aafee190c452e4af
z14fef97a17b843e105757689cfc7fcf219f4bc9fa9bd1289dd38d9aa9899d2adec881ce106be71
zcea863cddc0a1d97c978e2f2727e4b9dc4616655d5ecf0b54a3d6666a93e79d6bbbb20ba0c2a97
z1397d957d1d7f10970786812af9b6c826846773919056d654e0c4d9339317d2d1b9454cc64e7d7
zbe52e7e641e4601b500f5cea2cfd0aad15be7c3260f159e8d68bfb011e864c2c06b817bc5b9408
z859e38a91a981060c137bd96d9cc83e18cf603262fe7a64638e323950d303bcecc265f698313bb
zfd63fb614664dacd6f37057f643da4671084f10dd95d762f20657e60d88095889b71f6a9d33c05
z18c68b4f3dcd3b2a62b93a41b47878dede5d174dd535978a7d88cdce82e31b37098411084d0e23
z3c39a12392c34c75cc0faa4ab1e43475831aa8013b5186bd7ea7605c6d30edc36572892099f53a
zb7f50fb1505ff3dc41a2a9179780f6c369e5696cdbd7199e171db835edac3562ac38d7bb76fb6f
zb37ee63dbd9834c2d23c2495db180312ef009bac62dfbdd55812d2d8aa51b931f54568b92a0a85
zb1132dc22dd97c9de69a928bebe122a2d6e68a5d9e9840d1f9d8fcb3b35046fdf156cae8f81376
z32f98153aa1c8aaf4a65538b6d50059004b613559a7224d4aeca12b15655461c3200107fc4f967
z3dbfba055b33b7ba1253914e50953d61cb0727b495833c033b0f2cba6db040092c09b65f243c55
zaf3352dec52db61ff124f19ad935b5a2c014cf5e751b2b482539e86a879ed5cecc081db51e9e35
z5d7484d77888d80663a9f4fc9d853fc6369411bf2db1b774f5774fe37b85639ab34cf9fb40d496
zfbd08a5034e1ce28b2e96952ccd5c078fd42c27fb68ab2768325e6c72c462b0fbcb6746d7d12ea
z730088602b4d72944dd437253292499d80b9806ca41a56bb1d410462c9847756e28c8e8cbd1255
z8ce3162cd5709d0cfd4682c06c2344a824b9c0f14dcd9fdbc92743b62c5920458c425451995f0f
ze63d2c7f4e7397a95ad4b4460271ce28990aaa0a313ec80e2e6a0f526d6dc8d43600e07ff4bc05
z75620f3df996b23fe8831dda5b20eb3671e44d0ab3f5981569db6bf999871e66a230f79cea7baf
ze7ba299d796a4b148de1950add13a7cbfd34ca03f6d615cb87ed9e32c34c0aeb089a545df6dfb8
z9aa210f372778288efb1962217c36b21b145a87cb81839db3016076c092115e6c03538b5a814e4
z48c8b2e104c601dd0df2f090cbdf3094923ba7bcf6b1afc54c3bfc2d62d81b3cc0d3fbac42941e
z593af940e71feeee913b79c27d9e1a815deca734c6da20eeb8293edb941060e97a034e1ddd402b
z27506d2afff37d5ba59b84d3dcf61b06ab7bd1777f0713e4a6ef614c0199bde6a41501ff47a338
z14d9a06e9ccb7f2757412003719e9f16108495d1c5810b2240a66b5381097b85ef8c661c54a52e
zae041a25b6146a8a125f3e24c8e0ae9d67b2acfafa2d1ba56041e4e0acb48fb655e9a632e9b3c4
z8a29952a34d97af75622cd87085086ee1e1ff739b063ef5b174a4b9576fb2bb7d334f1c8e39dad
z38950a3a1a9c3520a5284f7235cd99119855a39534fe4c7b0298c43a0716718bd13f3b110d8827
zf85169c39b27dbe3d71c0ad7b28527a31ae3a604f6fbbc6f3046d37ba1a8466c5333e86aa3a629
zb5ac6efbb9552fdb423bf6466d93d8dcb8d79f4dda9ff68a3b6c91db752a9a1caf23b821cfaa00
z4c0ed3893c4564ef2d783f6de8139b54a0807b1efb37d6925e377caa4869edc9c87f6c6d4a4b5a
z9fa0c353730960768dfe5867ea3ee6fbc14edec9ea58bf313ae1162a2a58a39e5bab17f94fceb9
za28a21d49f30ecfabdca09d057b1f0c7c67b967c3a79d37d527a544a6c9435bac0505d13d42581
z85dcb31fd2bdf96b8a8454288fd8bd19c10ae80f738a5ac2deca0f4662a52d9cbcc0b22f9f4c5b
za2ce1cf82709272568810e35ae55f472cd4342e29c66a1ad3a54364ba10c4bf912d1a9db4deb03
z1ee7f377fb2818acb42995c4a9ec18d1fb5a0a3818b0b5f1377e80f185a7968dc125fafa71d1dd
z14249393ea5123b0fe6af01eaa2ddc22eb71fb1422759d0718df913996836c19280d1d27fb851c
za08b817c54d8cd398fdb27e398f7b5ac14e2a850faffc09fadff809a9042ea5e23eb265d82ab98
z941fdbaa3105ebf1dd81b5f9aeef40e3a2807cbef30ab35ba96ea355a529f15e9e2fc9bcce74b1
zbab0b9114f4d8586e187b11b51002878c0c4eeca0205b655c1c0c4f0a73ab660fa7de870c6a6f6
zae19b29af2714f1a13eb02a3633ed62891ef3d8ec55c7df67cb1e618ca35f07fb09d5ecb2f467f
zc4828cbe680687f01d3de3bb973a9e6f70202e8aa7f4679cc74f5bf30d980c6f840cb025deaab4
zfac0d58c976f76da385e02729647a95a35cf34ce28ec81007ee7d1f9ecb8b8c9a9aee76677be89
z6bd53aa4a93739de0d1af44cfc5d28b98ae4e9b5da69aa3987b4717739e844bf6e1ebb1e46ecab
zbbe3fdbf530e865acdc9ff4a3fa54bf156fd0cee06a18325b496d5f3b62b6aac35b41d4a97fefa
zf9a188c2cc524543e695c41f88a1995d66640909cdeb929b40a75987802120a289b2785c26605a
z45b87422888a924b7a5359da1a2ba83515f131cc2cb547b2d5c728d66fe331b9396ca73532910b
z04a9e87f5f8f320bbe4cc74d113db3ffac80a9407c800af752c74ee9c8bf320a0ab15e77e915e0
z08f1f7652f70da9cef8e57e44cccbe1e4aef214faedfeb88fc2ea9d4e840b79a203845ca815c68
z3888d3630d6a3d44f388c2a94f5e39e06c88b1924e3f7db13425a4aec48a5cbca69a4b580367ef
zd99cc75799c476b647d92e2bbc6cdccf1558b79c74eb585ad083cf35f852e24dd43b270d8c1194
z6f125cb91fb0726bc3aa067d23d218584446a999a0b14ba4eb76e1b15247d6bb1fe575eb62ae1e
zccc0986ee7c126c0aa3c8234fc35ece782960d5ffd831c5045e9c0819312c56972db85a01eaee4
z699deefbf61e8c3f7338d2488d2e454b50918354fa6825918079ce18540ed961afebaf514e2f70
z84845ba457346af243ac31b81f06a8da25f495ff7e4002e9275157df7065cee9308fdde6006d6b
zc1d90cfdb1390b04f5dbe069638950ce06b5155f311b98e0360a67e7c0f020f2299e1651114b70
z9a99e0bf30f3d03961e4226c680845ba67a70afa6f51471f24e4af09da74064db71e0dbb65ee4b
z97f05356e1e854c00eb84d5872a6459433b57c961f2567d9971b707b9a1177bc6d6f240068b106
z074c8231c8d8ef269c01bb13c0cf568c4921d96fb8c382b1e31eaabdeaeeb290b3b05401bc38b8
z2d63a8928c7f92c4bcc5dfd621a7c3cdfe1db271c91fdc382480b06a047beb3679002124b02875
zebcdd2e4424a3485af71a98921814e3ed8b25048b8bce6fcb7166eea2287e502ef5866b4db6ee2
ze5bb321aa5e298fa1ebb8328358006eae5411a9807aaea785baf1ef6612417699698d3a8bd6d99
z4271e279cc948dfebccb56eab0dafe339dc5dd52e527dec3272f5b1ffccd2f74797740a2a85e9a
zd2d38dc6d6383c19a31bd3cf6fd8333ab893062c7ce290ff778e5faec6725de8a94ce6f7a00879
z9c0a2d6c3bb26ef13461836a84303fe38ae4f8800a9b47cb3a039e49e6f122c6e85295cff13002
z97372766d7623d2d63749ce9d50970c8f23e0cd94f232afb582a04dbecfb78b676c442945ee631
zc13c6c8f5416f530c764308aaffa365191fcf92472e95aec7f8d9186ca9428deef28c4f2a10379
z82c8d55134b84ecc7103e10c2dc9c8d0fb0392b95cb700352c9540351e2aa834990be75d54fbca
zf17492c371fce2dfb3f3fb93dcda21766df4aaee7359a73cf5e40a67cb16a7fe5901c846c9c2ea
z1e538bebbae2117f59685d0416e4892524f04b21ce12e41c700da605d05258693d0bd518e5f649
zeff392263ebe72fb73e88ba7f1a57cfd4039adc5c75101e6faf6159cd14f0a5fa078a65e45575e
z13d2d18981de9ee056d0265b0cf1307e7418e8c8f30eb82745b35af044b708581bc98bb9b1ce12
z1c6ac85b71295416f6f154ec158119cd8a911ccdae858a301752a15a318847cadf0a86c21348e2
z8d3a992e2503c11a2deaf667afce9a05b21490208d29cdfc91d30e9d35d217d04e397b5c5520a8
zf09e81b4d96f7a35415f11b238d0027fb4901a4d6d06f13e4eb6c915b3dc1441dc5a1462f07ccb
za63962e607adc1a547f1eab4c989af7813991c77bee73305487180f9b4057596b8f0dcbcffaa47
zd63f627e4be0eeb9bfede8935084f2ff5fe9bc0d0567e7a7ea5ce37d53bb3d38eea37f30770ec0
z64ac435c13647e34d390b8049e538307bb66a4204370d53b6007d8732f2fb223db811af3f83d13
zf453a7ef51dd6f2b0cef6b87fc762031433fd99ecde812a88f7b342a9e7c7dabadf68889346f08
z00e1b881afc5fe95df7b80c1c5a2102babe504e9e8d3eead0aa517b83c8b8a50be4837cf28441e
z03b9166c82887118dadd3d2210580aa6eb9895c7cfe2a33e4b1c06a8411cb09b5116b822534949
z4a497f49d2bb0759b3ff21b150d164e4068622cb327bc926193b98c576fa743236c6de49166aee
z31aa37d137c526b2928443287a0f3accb3bed1eb7b4da10d5023a5dc72dfc0aea02497c04740c5
z113e70863c6c555b53a4a471aa2af7764b206e3841baa503a8d18b46f8c0cb7de545f22f511408
z1bc0640db2f5c1d3ff919a7cf65f15d531723e59774bf4cba06bfe3e7dd2bb35264c10cc1f43f2
z47d1433d5128e70f798e41b7cb03d7c6e1d80b3da78c9bdadbbd70ed15ef31fd0cab07ec13b42f
z746ff10edda7ec7ad8827139e953ad7f706fe0bf041c326f966cf9f98079cee98d8d4464a5af22
z8f38528209c714834f66b4d43d0c983e0fdd525cbb19f00fc030ed4658199d7bb943507f5e0300
z1404c082ee7838c882405ad9b1446ea3c3ef70529cdc40c6a3116b7f3568c461c64cf6d65d5c99
z9a398d5a64ef61e779f43e0e3592bcb08beb5f49c707be71a18f39b0fe1c3218764e4cd6b08269
zc8f8b544dd7acce43853be814fe205658de18e75e7de15e6898b7446c8587fccf4ea1889f657a8
z4fc3bd79388c764e1376da385d1b7ee31ca6dad1d22ab1abc6c70652d5dbc1e282df28fd83130a
z5940308551371a05e1365810aaf23e7d2efb00f774b850a37b5e272ed1f594eb4109b2e7d4c414
zf3b9cc0e9bad23220c295ed27eed083216b99c21da5a73b7a23b46980fca70626f51c357e4d363
zb3db3e913aba9c2ce1a5426ddfe942ac066c2e88608b423b563754dd9a4614b6d4e5334ddb1b45
z83a789e07778bff7edcda562d529e202ab2865a03476fac71afa094d9f05b079112451143e4d62
zb10ae2d6374f1157f0a6a52cd421166a47a63e7ff386e1e3941c5aad43a2dedc49489bf0631f6e
z43005aa99e15706f1cdcf3254bbdefac72738047fb12ccd999d0d5df1474b7ccc5d0fa23ef4779
z95518145ef09c41caf20b91d615dfc11c3529a85397a1eca083eeeba902edb2ecff4b22d697811
z9f8e93f9758842f6ccc4c5a92a2249395dd10f3898cdd0a3d33b9423b2078b21ab8b29ce522ab6
zfbd72b7183eeddddb2e65587308311cf3361a30b7ce83fcf12b4822fb686025a3e527f7cec6f26
zca49ab9e43633673a94cf3c0174f25168a595864ee77f1f439caba6822c723bf7c2b33d8b441b2
zc8f09a88de8fde8450ea1060861a1113d66cc53234176f8b95ccb434d7fbf268b30d126786f37c
z5c9024163f85e26ae75395c1dca93c77e67dce421305b8947be716a3ab8c68ff7825d4aee71dcc
zd9ae38a6a636422e2735ccbcc8fbe4120a0bd22af46d00cca721f2024b3be0931d2645e7abf853
z3c33a78427f650e86c0e76d7eb0dd8452e0092c918e81d3fd4ed06e67f6d2c9d651cb8e84054f9
z9ed3b17d320d29ad077d0ab5a4a0305a3a15d8017e42e51b38cdfc7ad07f6687baf246f4d72feb
z71cf4f2f76bbfeaa1b3d82dbfbee049bf0551b81b76d279d4d75fbc6e1e142e6823c381fc78715
zdc038a10930a41b8ce782002dc9099854630a9f937972165d6d5530f133cea7582a9b1712dbb1c
z600b14feff323d3c19edf5c46d5a6781ded03ce522548e1aef19b22834e4f131099f4665b14d2c
z465eeda756f796aae036ad4e27d77a552e5cad797fac17d47e9b1d801285c15fe27ded68326c1d
za3366d1b36e722096a29fbb3f8936d6ba191a60f6744a863bfd80ebc6f36f16a83656370917e67
zd0d198284d448400662ae81eab2b3821f48f8786d641f7abd1508da68e3f27a9c532b47c784294
z450609288b4b50277a7dede89d6489d942aa96d519f3cacfd7e9cb34670d04b3ade87e5f251300
z90bae9d414582c3a3085b5486a2da3ce00f2906e16781dd9a7508b7e1c068f7663f07a91bb2b32
zf50349c625539744ec35c90728eb6aca86ad0835fe95ecc404e1d1f16b18a20f4b3056ba551b35
za18b650784c9034f0efe836f4d8c033885491749fb4abb03dcb6c8815f43cafa274fbe45e42b38
za1972151f4498a7e372b938195e44f7dda5f69791f525e862fcf3ce7b3612fa51cfdb9ca92a69c
zcbb0fb98ce0fd0c733b6930ab8742a23db83240f023cea79d66d7e21b3e6fde8730e2e843835b4
z7a0a66165cfed3502118d0c6e0f7adde580230fab15021d90f55977c4b217b077393a2d6c06cf5
zed15b90666b547d4edcb6649a5bafd80809a22c973bd6ac3cc676ec99693be02d943ea3d48a8ef
zebb1a00d704b9e65e579f877bf56d3879dd45da1db8d487e20a816c532a4930178527b3eb008eb
z8779e0df5ba0c12ed848651ebf60363b840c5fb377c78e1e11822299560329831afd8ebb2e6bac
z9a50b9e9d1f10cf0dde875322d9ccc8700ad162aac73eb34b7ee185836b15cf6b86c4df5a3878f
z35c0b9c57687e8520813ffc5bf42386298b1bdbb418cb1de908e6e00914e00a8c6a528ab5ebd6f
zb122cdbfae5b422602942c2ab4a00000c81db84edae57e709504cb524f2c903364aec88f252abd
z15ed6a0154125900182f93dfe3106ab7aca9c463db85cdbca44c70b73c80603389c6b32c17e030
z2f16137885ae1e5cf54cdcb609a7b0777907419fb45528db98a5865479cbde6eae12b37f6f3abb
zcf0b3f735a564d162b0e9090ac08797a5efffeabb7be006bc73cfa94e5de515e97552043ce05a7
zda73e8547d8c100d7e0d15a871ff12d267504244d36d63c1f9bb39b3ac856e587d91b3afabd3d5
z93a32276ba37da63977eb6b07f06a6f0028e63cdf32408501606ce9b4039985a8e9471969ed2dd
z0b12b7ca15a37e679c3997d14032ff437cce89eb5fb41ab12286f58c46accd2f6fc00d96af6baa
zed80132364b6a036b3e823f7dc9d093b9663c83706dbca2de07d54f6693f53c3b7dad31d55c164
za3573487865bb7b45c4f7e813a8e42a9595c2ba201fcd387381e0e0518be99ba10120d211ec60a
z28decc604d818aa31457830ceda975dfc950f98093256a2f24f9bdd12bc853c6fd3412b9eb3afc
ze6f1ad0752228cbfa29729bd25a05ff8039cce7a2620feadb53864d658a0dc80d20b5b0540b21e
z9a5786c4dc0919b9585d034dd39b95ff20d14f2c07e581eb3dafcd4571d1c54f4750e49aadfe28
zb583e41471cf3dc30644361b835467393772c8a05e2e4cb5e0e0a15e0440431b79a5bc64f92f33
z48460d38527de6b456dd561bedd56daded693505d10cffcf68080b9b2d8dc67f2be0627b86ef8a
z04c9daab64b1baa0b854454418ffcd259ded3d246ac5a19d609fa8155d0bd5ffc0dd99d5f331fe
zbf8927e51c3626b16439e935f5af68aa890ca67f6438170abb939c9c9683e6048cc029b030bb18
z75fc7d9c84db04ee4d1ecc508fe16309b37b517d6eb77a63c0745bcfe36b7dd4550c666e362b84
zc19cadead1cf769f7d41a91504e3028d79baf3098aca519d2ac0fc630ded7bf7c953a71e48954b
z5302f2ad3bccb96c63b4aed939a7759830d0427f769da3c61842aba90024b298a6da8b9f65fda0
z92020217d702ed0fbc30d0fa4cdd80993f2eb0baae929b9616b7eeaa59d37a673550eb4d60f1af
z3596c009f51ac844ca65395b741c9f3f70a193d7629b47b648f52efb80bcc43f4837f2caef76b6
z1165c25902974204c36601ba8f6143935daeaf9745c8c5513b2204d4b84b8af3438e4ff0a13eaf
z3871647e6ffb97eaec295ea7d134ebbdac9d82d699a96cb83e6e91211524b70c0bf5bd44e15e99
za3a686099a4ed26cd40ed1c9cd530ecf34966a6708f0e1f0d3a51507232778c1a047358f2ae857
z407c061c6a530a0ef0f5593d25c5f85b15968a66bc8df89bfbb3c468787be627291f3c98d33ec6
zd09f58ed3c9d4b196c5e4207903db53f94f21f75b2af91bf5b3e80a6476b79ea3e2f265dbc6841
z45777969a9a00a6894f072b2c6238b8061f7c46fbecabb5585d7c64b5f0d3edca8a83a49c92e28
zd88fd344263e4f312d5b0cbd17b314fb2ee201a34cb7d356635ad4a504d22ba7622f0831976ceb
zb1bdf42b4d50221e2ffdb6ab67f749d727ba95adbf6156e1b2c67e5e178416f380a3d2fff11970
z928249b977c13bf7110d371df92d620b0779360c076cdf6479783429fe3725508780a290bdb3c4
zcdc7a21bf6063035052c05780db042416cd2aa0418b3a8fa05391f20a28f78b9218ad80b1af511
z8147a41d153876d33c5507fd457ea5da21076b53548f64913ed8bf513598d5c969fd692aca4b83
z8479791dcc24285c95fabb3b9dee10f09e19eba1053dd77e3ee355edc9190fc5dcaa91336cb32a
z8511032b823f45389d405d6d85b62599806012bd8ec597e24194d888886114f9dd18b209866fdd
zb0d4952040db87d13e63de2020a401cc04137e1b23783e216198c8206f30949eb3b2410d1e462e
z733deb78d619397bba936fa7861e30a1dcc143df13b3762d47e654b15b43cc3ba25e67128f7758
z1bd3fbf9350d64337eb10245644268c5761c2c636078a036dce517fa237c24f40f80dabe59fa32
zf5f703e477d84bc68925635d566e1ab91be2f4227d3710267aa282e1e3c7b86baa5f5e3f66d1d9
zf38ef7b7a706592acb9e89b7650cf75bb70e8ea977ee07a6b7454f0d591e5cfda07e76ef358192
z467919cee30d5aa63da80c2d46a76f6bf642dd53864b005861ebf1fa87f8c0d71053eb4e17e9dc
z8f64e26cea89701a5ad31600f4e0a887ba9ea66104fe3f6092432717bc7245c4210bc17d16e289
z1b17c5bd12158bd4830369921731f09c18b33d235ba42fb89b1250d19c555c05ba0402480f321f
zf9549bd8beb5cc9316d571c4c3e11b090d1a885c488f553be72cb77498d9d2ddbe2ca328d94196
z8dbf15e23cf54a6beff31a224630de3ac534be8f816afb77f8187a1f7b5f0e03dfc8e6419aaa20
z827ab9c2fa07fe19b0b427ef299475a415df0924095fcabe690c75694c24f6d0200f6eb097f752
zb05bc76232fb2aace0df9a73ba9a638942737825c9dd96f0dcd8fcae6003640c29975a91d74315
z39a0d19423bc6238521163a8b369a0829eb6737c1548afffd8ae0a5f50a1a88f019b22e3890026
z2ff3b1c1f0d847ef7890ad8db8c3cb00ac601b3a9be4d90c766fe765b2cc1c2343a7c2efd0e6f5
zc77b912dd65dc8d0c03684c3bdd55e4a57f647726dd53641da7a627f5f465d12e3cdb98d26059f
z583113bf703e6bb8155becf07f23e9103923d23916f79bee39beb966564ce918681a28695469d5
zc6af342400cc6a6f4992a464803b76d96f411cb29d702d7d42372dc5b52530e292272d9277f4a5
z330a421ca106cbd121860b03add4d4c31d94dc93078e07b906e9b641fad64ad0fc2734b4b1d1f1
z119a4528991a1758d111d8e0a60b8611debde17921813f167196a9da7f78551e7693405648f06e
zb18f4f5b2b384d3a14746769438b651301e3c725c57e4c59e37e58b60f16ab1278b2902b8aef99
ze5d6b96443c1af05a7399e2fa0e1054961e076a8e7371d65b6c785c99bea4efa5c82bd72816df8
zac48d2e931bfa3b688e0d5e8c0c85550a75aeeb4f4d6651e700bddd141a693c4d697dddf307f05
z221e8f7ab592cc4aeaa8d47bd627c00faa68315f442ecf182069c90e830f8e0714028ec403f82b
zf8be711452afb9a25cb6182afdb00a4a67f7a1f1418919d780f2eafb25d1d60be4b4d801a85661
zbc84ebc70aef81c4bb07067e5449cc4328d79699d0de5bb5433ff6aab99ef976dee2a33b82d49f
zcd4de754060d2458800c468d5df330ee5b2cb20e0184c6c29d4455a3824cddc78a15ee17caa6f2
zbd609b221e4e8b7c3a019204152a43ef4b609bb082e3cbfb901b170b72b5d27025f785c77aff1c
z1878b438a515c0a937117bd4f6e75a3d0553a6fdf66cd4c8981ad2a13290630c6432b1a7a6bf72
z6850ce160eddc5fb6ed066658e65eb1d2a3c272b7b3fbc38399bd4c6aff7c28744d9acdb683afd
za95ce73a1bf98c2fef256151849df9fb196ece2fec1f1c65053b0df13ac7c35d4d4d0050bf8e22
z7ad77496d77c92c015d89ac219dfaae843b15a76de4299e46beb8bbb3d9028b4689d0d27891eae
z495515a14e9db861396438c884e4ad59372401992d78c9e56fdef2a04097ff1a93f93f170d70b1
z546340e65a93d2cad9d5725c659c752d49c708b9f91718783b4fba34aca339c9ae4977c5d73429
zecea36a839ba2a770220f2c2eba4486891bc5a89777c16a83b793576b761ee4df4db3f56451ebc
z157bafa709541db042a6cd0813ec0c978dea552041761ea3cbf492ebadfc4980c5be4409d71403
zb71d39d204d04758a3731753280e61400a49d9a6525d46e73e27e7adb2281b3c19267d2f0f86fe
z64be49690fe2112d2d174c46d1ed9ab665f6f6d080e5e89264f11100ff6c27ae414937aaf42ac3
zbaad6f5d29d98ff8e23eb057916387830bcaa063d31e59bf5b79eb636b1cb12e1af4553fcbf526
zc807ce5925b28e602115add029f347b02318077432234c21345672e6b9a52dd4f8e028dde7c716
z5d0929d8392511fad2e33382678bc37f32f98a62c0e29aef1a6d465dce849dd00343a5ee076f31
z53920ea76c4e704e097e9f01efe14b496cad3a1e54ee60ca504a40a9e92188e97108aee0a9f768
zb6f0c80d8ecfd92b3407afcfed57555666104c54fb50ad8c10bf1a2ecadef09a6f5d21c5dc06c7
zb1e8aa4b10b81b821bef04b3a8c1e77e2afba9b13bcdd5e948caf1312ea45d9f8f4f70f19bb79b
z30a9c3c913f266edef5f0dde21b7627c3c07d0045840811a26c4b11bc8bfe7a89a07db0b8306a9
z278865c1c6fcda941a51669ad032417aa937b93929a0b4ed29a8b13038082f142dc3ba9ca71df9
z98f867bb365e31c5384ab365e89224ffc8777da92021a82bf3f5c81f5d4495c63d106d9fc56267
ze39954bbf16ee495e9d5ed57997ec4d2ee76678a47bbf3ac92684dc7deda112856472302662944
zf5861431e02abf65aef1a5fdecf96924ceef4d2bf9b3918b1f62abb6e6a17b9efea8ccfb131361
z3f9c5010dd57cb1100fef4c57c99d956183b271d5dd75dc6e278d8eb2c489cb9ab3536abfd8b27
za00811614077a557b9e4d718e7ee14a3fcc866c3f09cc3fa54dd11e2ad426708c6191bb8291161
za6de9146b5f6793bb359166070ab48fff37ecdd56c864c62094fa7b00c462ed6e51bcdaca843f9
zedb21496b811b79d46bf0f008df6bf567072ca54af56280f06de4c71f460c544a0186a855df016
zbf988751db936d4d4ed736b8ba0f64b939d57941daf0bbaa85de26c2450b056db5dd59582d994e
z0f954824b60953694d383d3a14fc77cb33eb12f8a1e3554395186c8dacb1bd6feae114b4be893c
z41365005478eece7f5151a88188728d7a5af1dd81b3876974b92271d328125618dcdffec593707
z8871b4d7a8b221b7b1f0b9b7c754f4d73c2b786514413ba956c1355bfb5529d1332149b639b67e
zd29c4571ee870a71d47031574b4e14dc69ad9c3eb668e8743e47b9a25a40268a4a48721027aa80
ze98d3e64f8656f95fd8186c169fbf2c42fe520b47485d90230786ba569a774ae38aea04a2114c2
z87749d3bbdb940c3ff15ffc23aa153e9370912ba98fab439fe5c751a1e34f74158c1a9668b5106
z71e81179fbfff90517e084da8d1ca9a7e6710acb3e52cf09765274363a417a4c1ac07ac8000e12
z2ba979809823928a5ef50ca8a5ec1c78e4230a32b7128a123ac3ff01dee4417d7b459a560544cc
z6cf6e62235fb47d05a52bca28d411d2412ac53957fc7407b7b9e9980aa6139b05b3d1bb814805d
z224c3dd58110d4aa1811eea493e7e68d061ee2c3b1e7acf38c02bcbe293ab63edb2d676a740194
zc41d2fb5f2890d1040da60ee10033cd1659a6fd5c950f36c9f37add72d30441cb880056034fb10
z73daef47ddacb3805b3e8849b718bc9ff3c02edd78d505c5815c5c5dd16f9f19106bfbe00f90a8
za1d0a7937c903cb47d2a281dd923be54a4691ba00d179807a6e30ea06d3d1d36b6725420a3abb2
z53c29fdc35369eb452b600a36abf5fa8e8a8a10b9bb8608c091702eb07cdaeac084c28e5e130c7
zec0cb9383f0482eab3ec0c4ce62075c20e78877383b84660b51fad5cb3b995c8431594132970c6
z73a2f2fb2149b0f592239114cc7e6e34d40ad2c058e08e182f92581f15cac83fd6983cbe414ec7
z2a00bb0a49ce66995471517b96d0814f546d63a63f7dc1422a90a448658ff97fee88009920d569
z5e241e191bacf67235fe51c3e2ec959183ed1a411af51db36cf4832cae4e517471f763b7cf9272
z3080eaee863f5f03f8580a6b6a7c6a9deae6223de067d0fe43216ecfcc3bc39c05c4f8050555ad
z7a36b6b86f3e6b020a43217a110ab64b0e4d9fdb57bb883c5ebc250b760b7674c717ffe96babbe
zcb5c2f3a87e811da86c5c5b197fc945e47f3332222fffabf802d246cbd9439e3dfc4855e3a9cc7
z094c904ec58c8628e8f3117e2f804144784004c44212c754dd489285ef04a8ee855c308cc21f12
z5042df236d05116fcc26f9f7bcd9fd5777204f4e20f7699381d2495e0dd87ebd2b964db97ca875
za2db7dd58d5054be6ee53aa19723b50bdfd47fb9cb3df3a66925fe7f27a07c57b283db1ff8b0be
z57a813326a10c5f68afa5d368e79d20a7cccd31cad0154098d6508cf821463a50b12c5f350cf45
z423eef0299da65afe80e766ac9998c57eada643351a4d7398827ba5317d24dcc3c5984e582e195
z751efdd1ec366d492564338eee1062107b7cac101fcbe10329436665a63cdabc5e5be50b1cec73
z58586aa245277cc653d03f2132154c7e324dab420a37537a54d94355d7beafd3e5d824787d36e7
z6ac000467770c1e3c29c26c241dc0c101560c8b0c53b5d78b6fbdc3115a7d77af5ba1199bb93c6
zef10a8a22ac7fb050db426bd7b367c3d37d0ba33a75b3b65690f8ee5c8dd6f2cc80e5e86d1a683
zbe4aaf05b12fa70ce7be93d77c909205a278783fd638dd16577cd7615633cb72fce313b48e116b
z86b3682347710135812f421d6e2dfd012700093e3a97ed92c2d742faec193322a5e9f96d52ad75
z9496f8fed84bff3e2611c82827383e569f5b215dfd01227c00b5342140203c77516aedbf529d37
zd5cc28ea45472d86fd84c670883b4c372c835704d846b801760d5fa9a41dd2535a4178f8e1528b
zd245173b574728a152393588eff935a12d11e5825cba4b4fe871605cf1d43ad0c8412338887d17
z742bbd395c6574c5e95dc0dc88030ff1241e0c4211deb6271ced4b11cd55509a4e04954f2c5110
zcc1270f1fe30c9742dfc06c0625fa54e928fa0a6d4d4882b19c3893639445c50cbd54062652f64
z8fccbb248428cac7b8bf954f144327378f972584c04f7d94569f475db1f1aa366fbc27c9b64e63
z753178af815b284c7eac32985dd3369a846c2cd3c80cfb0d88c8189604c399e0989b415538f38a
z219713bf696e8f5926cfcdf515b50a4cc7e358d6a195ff5965520489c7cab4ec5f5f1bbfac6e6a
z52100570f95eb99b262e2495eacba44de989f1ac79ac11185b20f0eda8316c807385f845c3f63b
z64fa4682cdd2fdf4fba5a324f9a7cb47c35715068fa90dd5b17a132fd372ee28892df8405ca53b
zb18f26c4e187655e00e645924298e0082e45ec9aa9d12a3f3d2f1d98959f0df4eb715934735343
zb9f0e5f24997b846faec038e60aec5536fcb622ceb16c4469470d5b407db69683ce54842eea2d8
zb864fb294d671344f9bc8a9e8755d1d443557d3fe405e350f6a65bb865e60950b72d81eb0de375
zaffb3b63b47d6bc423f1a395a8cd2998f873281136ab15d725471a2ad986c44492eb05ccf5d529
z388c82cfd8ce57511666f456bddbe1428967a8e5ab3d721c1562d4b40aa5b402ce57deeabc378f
zf0c0b31c3dc39aec2992edce9c005af9263604b5b0a85ca7d2c5bb3075ea2edf473a4344aed07b
ze36b8913540b0d205448024c52b0bd1ef392748f8c8ff6292f5ae8ab568ebe921820bf7356ea80
z70ec077323f9ad573680d0874784aa06ec5e1b237865f577bb16ce4f4d6e26ee1f01aa6f331e13
z0b0448d5f64f90e1eb95f34925a04d153cb2244989e7796db6e08465f0c1552ea530d9351196f9
z045d5f76c3c16e0d8a1d800681414457aafd41a54460cddeafcd7d1f2992c3f3fa308e511a9fc8
z0836691df13a87541d0e2f0ab28cc75ec287c4890955fa34ebb014b11d30132e2c41b01cabc9eb
zbf3aaafba260c6a3560a6d6f6aac4f2d5840f198ba54ba7e7a84effa006be0b89fcffbf07e2e22
zc9c1af4072b1befe100d9267cbdfc2eb152500508868263500248c78bd930c00a428ad3e6dce3f
zaa8fed7a5fed5b5438e895e0e8e9a25254d189e9521e0729f46296dfff00cec34c612f1ea4c9c9
z3febd4ed99f9e55f6f2cef27de069713cfc44754c2addfd8dbf23cf60e7578c612cab1f666e3d6
z1e3779b306ee4b8c6e28506f444399388214c353420b2bc89163618641d0dcff341f462df539a1
z2ada530ca1cc38f99e503ee92b53fcb8c3dba67196673aa000eda47fb45a77ae77f79480fa5b1d
zc50bcd661b51a44bd5d4bbcc763dca5b87be64f900f831a603c7fa10df61ba025353a1a068dd67
ze152855ce7dd0aecc62e3e05e953fe2340476a1a2edc7f75cbd16e3d95b9a4d60ba5a34bafeba6
z3ee1e3105c3c3efe2c4159b7f6237ab85a8c125f5ded30685beb1863cd02323aa60259494926ed
z9b54ce6f6081277a6939c57a69dcc30a3205c583c9a5f59e4f749654422d945e8c6e0672bf5b02
zf5eae65cc8b6307746211e5c5860c770f94333654c576fa640b87e52344ccf8927e635b0c82b72
z7ffc98b4169dccbb1ec6e814d6ab3a7e0d04ce91a1f62a7938cc73c6194fdb510280ae45201161
z3d0d1626b6d3da4934800b9696e7341cdf20fea7873c80b1e0ee9ae0f15dfdf65ece08399d7f20
z3c9d3faf04b18a36798663731ec2a66723089040eb1477b56e0b96c9f5f2dad2f5fae4f93cc529
ze33c52a2b276764812941b16fb4e202cd36f84a36543ddef8fa252dd55da402feea83a0fbac746
z0af9cb5b281c0f1995b5fbefbf7a2d1594de7345e7151eae52e4ceef6938d49a814818309554a2
z36e0b8d4fff686e2154b1bf51a5bd6eb1de968cd6b0dafc0f03753bcd69d354014de0e3327ef93
z783d631bd4c6f404f61a88c5ed07e83cfaa88c3c7f93f356a532c306e6fe0490f0d32ba9cff968
z181a0f101a3ae2b02fc45c52357b9ec1dc2f892d16a66b7af8b91ce9e8ff6294042090d98e6d0b
z9a5cf00c387d242630abedc5c17b279e37733aa17df5e650e6fdbd3fbee4a763ee694de23ffae5
z994543c119b7c42ff5d2a96676f434ae256dad5f12e24df7bad323a6df3fdd82795062138aa491
z9143a01dca7eca80cbbbb29acb4ab4b62ad446fad0eaf4600c9718497d224a95ed31d4131c6e29
z22c0b34f0af27dcc6b758001369d94f6d4170eb25632ee3b7e28038e850312ee0409d9b7b40462
zdbd9d7582239a0047f34e2a3339e76630f0fe38ec6121fb423c1cbe156ef4ffc0ebad0d7981b86
zce22d1929de51df538e52d742e3cbecc948201cd251d8e133e5b4bb8bcce442d9b9cd64b56441a
zff1692a66bf68e609de95dc198ea67861c52af4f44fd4768f876ae08e17a07f19d5dacb97eb893
z01b22798f4f9b7805806e55eecacf5de452b2b3fb8044d74d93831e6bfeee96430ce99023e9523
zdb5275938b6aa171a14ce4349dc2c42a1420991c7ae390263e6a4be199bb1642b944f997a81904
z41fd93b9d9d795c87923e07da9d5b6a70e16c6ddc75ce4ecefb18fc959dddd426f5d767de9c50c
z919482db4a2d18eb6cca5f885cb3d99f5cc62f3329c151cc7947e8e9c74d58b8bf9b9e6722e2f5
zea8250cf15f5e2aa55d29c2d3b29ea298eca1e72f4aa64644b55bbde84a347f4e85d37b121a94c
zeddfe9ca4e04b634e2fed135f0272a1c2872718db466b5335b465627e2cfe5db56601dce60de36
z7339d3ba8f976719b2aaebe22d217301b928065651719353708baae349ab550c9d6c152e35672b
zc71cd58468284d919b1c2a0faaa3520b652357acc5717bd560a8b1be2fa8a4d37086a3af7a7d89
zcf24b41164120291b2ff90b3df6c790ff17c9956af7ab832e592ab0c3b35c90d49bdf513a6c03c
zf15ef9f96f73c5fd761a18f53ba5a861f9abdca7774a5e99ee160c41355f4b9489e51d2947b141
zf4ed863a7698c97ffd52a0d81f862582956d92bac73f30e392b8a8d7a129e8a10ccb4241b91556
zfbb5958059b9d173142b8e9a65233312535a7a4376e188ec7d0bdc3c2bab8ef614a3dd22de3f81
zae7147adac07eb72d3252fa817128d655b46ce2024eb8da03729935a2616aed76e84618f394bdd
z41176b59404d289dddff89d873ce665a9e9ca3f6600fc815b3bbb937cc45b05ff6ae53fcf907d4
z7931f9f3c035fcf5707c112947c9100b0215a736582c669958618d665c5a9bcde7f50da34a129f
z8424b704d091159ffd338457edc3d9201479e4960bb0face5d64de22d95fa187bf837c40a931c7
z6aad640bf05af53cd7702c9704221e4d25557f7f9b87b22f5919febcd24d650d21ae3f6b214ef4
ze4fc5345e0d2a594373b4bb9869f033d45345930015de34d70c1286d3f8bdd7e2e5d76aedf0cb4
z6d8a3c96f105fb12b613adce9be198bd3f1a1373c4d58f7ebd2f4facc9f9e5d3282a1274c29c37
z5f1616276c4d9b969e71824e224d2d88ab7dabb9a92eddac18d2454080555d42c5e4dc6332a561
zd286c58a40f70aea238053ca5164f1a36da263a12a34e195da3e9bd503f52f8ea8dbc046b4eba3
z45f9b3f0d76abf5e6fe6bf31fcf33e49857f1f0e9b3a2bbf82c4b3f0f49b7f96a23428b2a01e6f
z757e399b99de30ed08db2f417a7f4006f0f2083a01fa2d65b3f94c5c87c3bfb50cd4a44583a7e8
z113d51053e471d1fdb011beeab9d4a465fdfb1774d305e18bf891975f1d1bba1fd5804ffafa85e
z3c6e983efbd6e966dbac4770e99591bccfca085858e995064e7c1f640b289b37e224cbc18d9d4f
z7ceb788cc9f5c4cbc15b0324788c92f035ccbf8286dc542d667cd18fab62263d11d2d250993534
ze54a77e4c737c48769eca6c7841f086ae9a95ed789bcf6f968f604bd586f152275d422662c1c87
z42d694e3102b3e0e7b8f979ff6c5c69a1e0942e1883459cf2003d78674b8c47bb31f05ee47d7b6
zc3b208000979b7275770701bede12ba45a0b96bf63fdb889d6745decd71f541a7efbfcdd9d9e59
z35f45fe7f56f1d9b07e54fec270058ccf07c39e1400f03f765815337290c2364892f07934502d0
z915b151a1d9a76278a6d254c5e056d14d9f9a328d0bacbebb8832f4fa5f5c7bd54b4f6b6e94777
z99b9b62bc6f4f24d8e8e1373bcab75e3e67fcea1870327b4a046e4f8d12cbe2abaef429e600c69
z3cb93c6ee271feb468f63afef412cd3c5289fce358b9b24fb1a8c173ce2cf394be2814198d04c5
z62934e096f2465219e5127f24f3fd62a00861ca251e7fcf412453559b9c5ecfa315c162ca6c450
z5ddd1e3f7629ea7c3453446ec303ee2213db4c95f5e91f41ded7a2cb1fa8f294b408e250a65098
z10db7354ace3423555cd877b60e5a2907c95aef96bd9b720abc1abc8cbd84452151c4af0e99495
z852ecfad297e092146587beb257937045ee972a77ac03f6b362452f866f03b43b1e493a2e4bd33
zf81c68a21a57960847bf71fbb9d44edeeeb7409c74d3439b368fc59c81b9dd3d0d2b68b6697d73
z5beb864a511a8cb8c4bdf50ab29e8fccbf5f190ff5ec63e42001e9c9c6e4aea964264f8608d84c
zf42bacfbd35a6bf09a2d37079c6dddd5e562a35f0092f0307ce6d335de7f73a44cb00d6f54b95d
z2e366af601b7b247425aa5ff1b25cb2c9057228e7b3aa732a46d5ada29976a3823bfa65eebf784
za794534ff3fccbc1a52ff7cdc0adc55781f476742921c8d251aa02bcc4c8a815f279f3d12e5947
zdf7f69e794d92c21cd996ca09c6f4dc9c0566a1d7b48e88076e7b628b3827ddab848c4b820d542
za6eb553e623c921424c75d97da7bdf3d23dce61ff41a366850f5a6e4c34b49fcc0e65902ed0d66
zbad3191bf5aaa134b99dd698017cb59b7e6219ba394e595eaa62ce3cf8686f1e5793cb2143d151
z751b29e3208c275ac29cc30fb59795afad72cdf5e2be037585502b80960c53fb888ae4f8d0e326
z1eee10eec614363f862c5f89ad73c4ff31721c908946768bae79c9dc12a9f648cf1c3408cfddf2
z2f74d029b6b89468071b0a448e3d96071bb18184f2cb13d8cadb460a19e363219e5dc162673ec7
zac5b1699541f8bba00f494a20d240ad426dac672a4f36c26ef5753218578dd79f7b4c972005fe8
z541c6c9900766f1b8718d21a8fad13f41a016fb2a037ffe3476997d422492144489c294d4e66cc
z126d705e19f9c0b838fd79e43b97110bf256fe45f0ea0b1e3f2f9671fb32c116b35c7017a0c35a
zc8b9754262c830f4e6ba0ba6eaa92af218569e538a9efe2f8552049c06e5e525f505618e5a54bf
z6f730b10a1e039987a18c1e5d1f3c85ce6dbad65d21f93bf94e377855e109374a9c07f2fa13b50
z34e6795fe68f8bc202c5ce933d828ecdbc4b182fd238c16ee71648000e1b5a4fd60cc8be70e57c
za5dc9473e2ba1b6d8cffbcb75f9c4ceec61e2600c1ccefa635bcb0b5635e3c64733349b93fbb82
z4ec6ade896727f23be2713a54e36b1cd2ce2e82cc61383113f3f5b65cf744df8dc7fa72ed9e6f9
z3951e89f9d44801a954476410cd2b61648ee4277a7e507e6f3a2da1a181558c8b35aad8beff9f3
zec553a28be21acc4292d6bced01c599b9e9a44cfdf1f08eaf21798c1bb6afc1ca875794143ca83
z79a0c91d5d9c64a1865bf6d8ec11dbd2bd60bda2b2f2498d9f3b3946d68f2e0c5bab77fa37d7ef
za4c4ac8b3feaf9263dcafad94ed8a475394790324a2343f72a4f88e5f32bd331b1b246fc9f5a63
z25fa990b71079439de5e54b76bec23eb8f8772561534a7fbd9e64dbc8dc2ecdcbdb975336e1143
z51c5f21e7aa1c019cf79821a9b1c628d3b38323b5a276a924798c1c83cabf8e6f84a5d5ab7a0cb
z877621be32501aeddc3bad12f65d24da5b5087f8f9129d081ca4d853625f2ab6e6cc1c33bddf30
z6f6d4f97c4c61474a8ed76710073960fd7e1c696c90046c19caf1b5293326d622087bd49073099
zb46b14c53bed2b0041f925ce2b9d5ee417ff5863e89cc22b5708035b070f7f483f511e964db0ee
z2c0c1335834702c8300b69d168ac202338fa63da9e69b696bc9e59b6ae5a658d811a0ab317fe6a
zf068656d0259bf471b484477d26e883ad3f10bc1098a8d36bbf15e8ba465440868f786515bafa5
z2f4606ff9488b82e8bb2dd93091a33dc77a4117828cf32c479ca032035d53b78410627322161fe
z37169fc84004e884d318572a65d48f6ce44ea37f4e77d126dae92c330ee3e1bffbc4fb84a987fa
zd67e272626b7ceb271e2f83eb30b1d90479544fa6af46a2c77a9eb8bdfad908a2234a47ce9008b
z381f3fe776f30ba0d0c4867aaa1e1808664defc5977cb7bfcde92696a84057bb378c06a4ca559d
z4956669f2c6df2690f48ef1b6b7ecef565c93a7fd02a720c62552123bade564ab5ae1b3e03799b
z511fd64d43f5d78a94ceaac38e7f8ebf939da6e0ced6968dbf67bb5318f54a366c9e64711b8d35
z62ff12f569dc46b2eef3c024e4a670903020984f1b19306d97e19bfd94d69a959d83f31715fa20
z3ab9eb12873818e018d6c55a10924fd201eba5adc5d644134729a0a05a9fe3dd055d7ad1fb9353
zcf3537a338c1a7188cabd1df86ca1c07b93201e21138e19b870f65bfc4ac132cc90730dffff3cc
z4f1d1bf42cfd46d1d4b6e74ea35dcc3144890e4ea05b96f78213ca466c21caa7ce5670a4daf0b0
zb9309f105ca2f33f2752ccef4d05a1bc807207490d5a4fa72379b6a21e21144bebde121b73df4f
ze655881db7a8e9abce828997b8c65fdc351c68b90cbc397cf915d97c61f848957cdd89fe11c1fa
zad1f6e57ab48dc9e8b1582f088357bdd0c8b0cf6e2fbb9f88e91356c2c0573c00f183901b1dcc3
z2a4b584738d0abce58921160765f5834b0fa8c77c4d48c9fbdc32a02d54a857ec7c0afaa0d77c5
ze3b1e234ea59ae24617fb1b69ab1817e7cfa2f0c1a69decddde8712857b6597c825bb80dd5c186
zb0eec3db16d10c75d339416d5916bb7077ddf35b8643427aaa4c51ed1894901e871ea402eb8b3c
zfc29a78be197b885b29280d054850ef46f63a9c2cc601b8c48c78ccf3d64c426da1127f905c81c
zff49b3228bd7168829b2aa12f50ca9639fe905b14377ea87afd1923a7b8f8c8c27021aecd5b818
z2aa55a79517708856a8b2f9b9141a5ab42bf56f732af685486bf0f004fc1760769051e4e4b6e23
z8ff4e9fd04f0ee21976d76f4d99caa6e47dd50401b8453d03d87c90ae38406e268b5ca3b5477e7
zc2c691d7fbd55bd8d515a6ff0c46f50f11f0535f3fb082652522a5d304b2099ded4afb5503cbf8
z3edc95e6e4dd937c35172d139ddc160c484b255e23461dded434df53d8742ec1759aaceb87fd36
z0b7bcd8a867f45c454b65e4a1ee9beabd383ddbe109aa7c6bbdd01c6277662f436fa7055b66a51
z95b60f221b46b71f85e617db2b99d106ea084145e413929ed91261e1e356ea6613c6c469b94d67
z76727bb40e3da2314fdd5e08a540129377eaa10dca4180b8bed1a9e1cecbd11a6f0df86939bf9f
z8cc52e8aa729e1a94b7ecd6e38792182b19ff2c8ad7fa9010ac32b198718132fac21e4d0947814
z015f03ff4dd9f25bea8a7fc68e9f04fd17f898fe17c813e832490dc7a6619f997ec0e12eb6bbc8
ze4b8d0c9e6a67573b710432ab0f26275abc2e7885c7420360effd2df6b12bcaa04cb9965f0aaa0
z2fde98baccea501ce5ec03d4bf8ccbbb05da0401d1d8f75370b4fbc35a78998473dc0fe8ca41a9
zdc0112f65018390a00cc6c2f970ee6ad8abfc3943d8e4c5f47df0bdeecfb8f22d95106b980b10a
ze842016f3eb6770b492f2d77bf0c15486492743d4dc36fbd74e561e56d615913ee8cb689cef0cd
za07f9aecfc7b9c8486b17dfc74be99e987edbb1942b5e76b0f0c45bab2993f766daa9a450057f5
z2410c87cff2817ab4d66bc8f43e5cf478bccc4d0fcea1b71b8c77c29497d3c00732fea537100b4
zb889ea2504c52b49e9ab7b5db6a87940417c0731feade039619c566b123ca3336a04d1c4adfb5b
z30500542d429b9d61b53c4d87c1ce6a775d72489add2bee504488b3660ad200e621351fd81d710
zde84185576c1af522369d87aace5cd653e7df172687c1a05d66198a3ebe8766977725091f548d2
z1b91ba9d22a5575d2706788d7ad2bfc69e93c6a0a7caafe9ea214902466086ff01a158dacdf6a5
z949810d23a7e99ab3157d88c35c61650f9a2fd67a2e9eba998d3acfb7bb2e2efaff57c3490f94b
zca5d786f731eaf4d9ebd797a9551fe21962601cb9fc4f97c8c4279350453e4d220204b083ab5bc
z809814e53d0a03ec72e82d151529aee82283ded1c2a09cc9d4517c3681f6a21ddf63b2dc340b85
z78c98014e62c12843c295bab0951011030c2aee80cdf7d9282115d89b8d92a783e1c82bbae24d9
zcdca66f6cfbc3f01bb3c35787897f06b84f002c7082faa53c078ad0b259d81faf8370b9797e3f9
z9f22e8f4f617933b0be01798631861adfbd30bb833c10df205a4f6023fc9dbf6983f2ebbaf95b9
z88d2e6bff6134e2a9fc3830959564687a69bda6b0efe3dbb964fef21cef7a02d8fc6f20f0eefb3
z19d845cb10904ff6943b76bf0ba20f66e087d25b05ac1653659e960923776ded23cd94bb924e4d
zeeffbae32dccefcfb889cae93f013a84b408c6aa0a929cfa556c119d53ddb8f0c85379975d1a67
z953ee423cce8c47ae3847396e8dec38e081efc063d07ac782ae7da55fc6d5ea0733c9cfcc23511
z5f17157f6715cbbe37a58676a33b5f7414bf7ca383a26abd7b59cbfe597a8e22c24a8a37510b51
z58c406172aed5d5f6b1ea2b3ce7313bf762e51521f30e3e27a56c25b27b05726ceb7588e762db5
z51229ffdf49a87735b74f479b7fb54d833f4889c4328b6e9bc8a64b75e2260b207eaa82bf93ab5
zfb3b2e805fb6b9287ddd0a6090409023bab1a99a7cd8f19263d2b16f25375db200383ed68fe850
z16f507f0e39e9e6dcd653a920812db5cf0450c9f55167c82450d11b57b8cebd14b50a4ce90130c
z6b3e7df4b482a14dc0a664a3de384ebbdce853a5fff01497b6fa989344813359d5feabddb5ad35
zd9552f6bb314f4a19dd092a1c8b8bc3df9d1cb760fdc2c4b60de0503fa9c54825905f9a047054e
za3a65dca360433daf73f095d0c3d4709c6d31e1d188b4fbe9e9fd4feef8cb232659e4913ed4b0b
zb4797caf73a6269b3bdc36cdd62f46c15ae13de001893c3f072402fd1b985eb362b9cba3f3fd3c
z9550bc4477e53fd4ea2a0cff43a7f948556b662032b0e3f9954347eca93bf425f7109d9569faa9
z9eea571ac00342dba6d0488a31051c653b49539e649e1cf3b2ae4c2a40842debb3fb481836084f
zcda6e5d7d76bd783245982d4e902ec8ad0b6fd2783ca9b1bbdf6a05fafbb6044851162628ed1d7
zd033e4a0c14c0f37d1b7bada2fb41cef823fcea063ab677144fb2742cafa57a761a1bd01e86f52
zd87b6e560bffda91befd0a1726992ffde542e58692b582a191a32493bc0e11a0dede3bcdc6fe00
z709575a334ae281c126976fcafb25323fce6ba9a4486011a39fbd57991c62e6cb268024f1fbb56
zaccbcbe635e9ecd2d0c344575e968d84a8a5f773abbb1306da43b993ed250c1b082b4e46627ea1
zdfb18ea55ad85068f8f645c860b71bc159512c29686110e3c3998f3995dbf0f8fa5e78abaed1e4
z9750d47fed0ad7810d2e346b126f8180ab3150e514209b87d399e3df8c4617ddb7d4fd81812f12
ze3343990c17fa19ef1ca8b7092ff267ffaf9a89f4c3625b56d9736e9e52bd0742a0afa06269a6a
z1c6a9b8592595e67e373ce6f3e606eca14df61a57f6bf011d9e05c53befcbb8456d3f8a645ec2b
zc6d50d88f23cea4006308da68fc080142234860b03849d83f363e8ffec543f9b5f5b6e8d46a767
z02b90c9c0eace7711783aff62e1aafa68b721469d0615c238ec0412afa7d8e9b8287c620eeeddf
z128106a21766d4f53f23af3345be55d0b00b211e25eddbabe4eeb81189ca5ac3b896f345542c43
z4e06241500a85caa4874ef40db87e7020bf44552f0e37e2cca1cfcd15a6c41efad407a33452ba9
zc160fa0923cfdd3b5ca1db004391d3975a389480331d082d2b3fdd4ccac1ba284eb3125f16521b
zd5e431203e1254c474690ed422b421b205e033469304126ec85f94cc0acea15e03fff1df44e344
z1bd9445586e33ddc047c3bc2f06714114834fc0af395459697cb4d28801151a97905c69efab92d
z2100868f9af8700d5b1e45611d6067a1e679ab7ed8e5e42b9fc9c9954bfd0c87166f4f350c183f
zc81ed3a161312a4b6341383fea38b6048f47adc3311099402bd4ab3a8d8241db3c8a290b68762e
zf6d2465208f72e4ce98a387aa4012d6483d89654b55d987f2e4d424e5b2d5a46ce659942b5475b
z98bac1487053241b51144d1d84a32db31e087646f1951e8b2c5552d5cc194f2a2dac287a0b2e55
z76a98459465c5dbb0a516042cb0ce01a5dac1e3539594959989a5f82a5a5d44cdebc8ebfe25f26
ze4e64d8fcb18e092ea721f538eea5362c09d02f922db727acd92f1d0083fea26b3015c29f93335
z7a7b22432049251e0e4f102b5453c307212f02b371803fae5b68485a8d3b330322f12a2f4b50d2
z5ac8f63ad05346c4aefd89f7ac41e908170d91597a2f3edf1c60360cc0e2fd92b62123f1182661
zaec38001a7763bc85da2e14478434cf4e3182161004a5e4bd3b07e9ba643469b86d43f549d874b
z3a3223f5e7de66d7ab4aa83bb8b896a4280123a67f92703dc08a01e1f4be8254888c92216eafe3
z0cdf73755e2662eff52844edeafcdc79d99b6c92c3648348ca5f41b7ccdd6952021b771090a6e5
z6f90920df9968b8a69ac866940e50e77389a3115ccfcf9e8694368389cf7a196b52a209e783ad8
ze0484157c8601b3dcafe2998e8a55a8af8699583a062c992759e6b46805b645512209a37068318
zea6048b7ef10c9107a5fb1e693ee285f52d87f260173d7cec525cc7bcec7d47b3752431a4246ac
z6920708e0b4630d494d9d73fc537aafbcd56f4e984b178a762ce87b6c2a6f689bdc88b344a7010
z0d8e1b73b60cae27d41e7e5296dc9d06d7f21839c0627aa05a003ffd94efb770934d5a3afecfbb
zd7f511ea7f0e4b9472bab2e1aa74031b377cc96084b35611debaea498a4d95e80ba9409d24091e
z298c7caba4a3ee6f774e28c4a23d02a29f305fcb2988e97d550513a087998e8fb605814539dc85
zcc4e85b90b0ea9abfec6cdf531c4f7ce4d13ce29023fe769b8e9f979222dbc0146b51abb8b2189
z45c8c2ed2d5d27a69d989adc5cc5265df932c99f48261cf9eb5216a2bf28cfa47f68c4056fff48
z9dc1c4b4f910d7e37f6be11495a97f4e40831c450aaa178488a74234cb24c64d024044c306bc50
z004c5bf14955ed4fa175f0dfa0171d8790dd1a336e1fd5964067ea3fc409e06c6aec42c2633aec
zb43b796b74a07c05763ec110cf48ab0d6833aaab698ff527f9faa510dd7b42afb1b5a1f803f4d7
z4c6c9c283acb08c5838e7d9395f2b17612168752a5663d01856be985355b7d564f1718d5d63f2c
z70579e15299a14ea0847b10b95d2d98a2819162c9f4fcc85e4f3eb1fc950e152c70f1f807d6092
zeb8a709dea07f3354bd1a2a6f914a591de3de755a836e36538b7870f47952231a35a3ec9182540
zc4753fc7e8c81bbbec2c5361cf071456a0c545b686c21108e3deb9a6b2396f082b329c2cf668c9
z7b52161404598d517489c13fc7b41c5326148cbee52346cfa029cac13dcb958a4306c99121d2c9
z2c6417052a348de68b82b6f5efaea5ea9233a1d6c490843276198b9ff8c02c071e2c71e8f41a50
z4d0fd7389518dee0eb1c93c109d0601c5440a60cff6e1a168e983d6458c05ae226ea1d813ef4e7
zd4acffb61c8c89b09459ef6a3d572216da37bd3df9e4f468a8f063e5f60dde118f33a6b5e4af2f
z5e60db4f996eed5a4bc54f16d90f0f894a4f42ee7fdaf57fd9ac96ac07c11303f956b95acff9be
z61bf6a0967880b51837db4888711fa1d802f666db70f57194eaf4813c2a3edc38785985c2366d7
zee0d6982fb9157086fccc1a2cc7604d4817afa3e52f6c1bb90803d4cc9b6881fb676162e96c5dc
z440df4af77ba432790a46ee5779384bba3a640cc026b45681cb73cc2118b78588cd6ec66f4f42e
zc93b7fa298198eb2f226ec6ec4bb9e9c868bee89bdfe375f136993ac9723c1243b9d01a4e275d7
z927c7beda3923388c302915fcf7ea385e6151b7596e97db10430243e2a35a1e3716eab2d60c90c
ze5158ed5464473c3bf7accb7d0072d14b4f77c3babab2cc3280aaa1d956743cf308992a421a9a4
z9fa808ea83c53f2dc58330bdadbdf63e1cfcd4f6099fed4a72b05cfb412f19101058c768369178
z3a3ba37c08ccd94b10640370e03a30708a751219b40b9b2ed57e05c9c879f9b655040cb2077abe
z4c3b6914b1bde494d42a50372fba2f3c7f5636c5d424385bc39baf68aac7e55cfd90cdacbf5c02
z7e709158cd6d39455afa4c4a0e156c9cfae987a3e9f662b00ee3062678831f7ec6a8feb229a439
z6fab50c23d37378844cc8adb141837512768797bf0d4abbe4d068d15316a191aa8a2062054d49d
zcf738fc986ce8b14f18779538aeaa106731050755936e43f4132637a79d856d9031adcafb29cb1
z45ed6af1676d97063024ea3d54d55616a5581e9d99f0dadc9b95116a3e040a2b4be8f200b99336
z16eba29a152c39a5e2413e764e6c0dcb6d5581c92b16e6dfc38173669bf5e7192e5e2ce6f9e46a
z5bba098061bd680c4a0814d4f346371526c6ac68fdbaf7754f6ee03f0bfea840ceab127e6f9d88
z5004230fb51cbb4390ed57db07e9cc8c687f8fc5b0085564dce4baa7fad9d83ab27a4f422b8240
zafd5191fa850136add62c803fdefa71108334592d59d1fc2e2ce66d42cab1eeadc353d8b03f5aa
z9ccd5935f1655909dc7e20f405427d0462559118961fe88274c4099ef1e3b44317706a7a40d82b
za6f5269a3744066a1ba8b4c61a3450f315387d330355a9716d28c50ebad065bf2fe1421bdaffb3
z879b196f3135a9ec56de5bed98b5d4e5f2fd4eed684652561a7ddc9e503f6adabb18ef5259bbc0
zed697801e7f5082a52346a7b249a4757b55f31baaef4b8b38d2ea00cfc400d9b19f5297218e398
z524460b38e384c9e55880bd3ffb432112f60684b5bc4223a81e58bb5f6f3a8683630266ee39219
z235d41742275e072bde36eca8a7c5d3d540b5ce727731dbc4de7e57ba66022f2025b98d2d0670e
zd6a43ad7beb4d2672c893539cadaa965b36a8510d3da06179eaca322209151e4051a608d3b0fdb
z0084196c5cf9c61c0aaef303530d00f4d1646d1f60e03f57955bd63701b05b94cded1900a8ba14
zc7ff6466e3df718ed142689aebc509cb7c1f18d0da6290944c4dda90cdb50dc0a1b9a49da46232
zf6ffe41e8a1a1ad7a9f3097452af7063a966932ef8ea027a747bc87b9b0c1c113cf48848ff565f
ze7f501ef86113108d47b3068ede48e6894a8001b079676e1804c309a418033bdf6a4a97bc32b2d
zbd6730e7195436c2fd2dc47972b7e79c4cdc5f858e465eda22bb214d8018e91e0e03c4a1362af4
z2776217e759226b1b86a7aaf1f693f6c9a42e81c497be3fab9e047bf04c4ebf166b46e8a3eaadc
z50e67272c2161d3c2ffa9fd2f6aa85c171d4f791e35215aa3f9a80d205f3b413241c158087abfc
zc4ae8c9e86c15111d1bf30819a0897b1b4c541e8008eb14514994161bb8514f07bf4378463be63
z137ebb38dfe37ca1ee274971978219455e711d3cbb9a72748507715e8981b0386b0cfd5339f7b4
zcb6cb9de87d92502cd7c04798801dc818aa7a5a500e365764c7af7b365a0c2b5cf8cd445e122ea
zbbc47e7bc12dbe5c12f88c280cf8dd2edf4a395307e21e383cb7fc7b3953e384902ca756173d8f
z3dc760bdb6d2ed02f1624801868d298e037653ceade06f198eb47a6f194802cfdadce1c6078534
z736976465b9ebeaa8deb8ccf310c066403c14e47c3fdded88cd71beb99e457d96ba4ea0c846222
z2a5a1b39c55a2a24e726db2e085ff4b77d540caae1e8b1d3b675a08c05881cb391970b90f748eb
z20aa32c0d5b20fbd4b41f1320cefb0dfa918261d8e65c4b1a00404950c9f5d192451f50a474f9a
ze1104bb392aac7a92e1e1e4c507bf9b9dae5d17dbb9bc36df42365a239238dc5b5fb8bef1ba097
z79b6ef1eed02c7ac3bcc5e5a601dab1cdf61307ec6f2d4ba519d0086e5db273cb7121447952ba4
z89544ca91fe5172a388669eea6e1ceec44a1f012365bb03ad7896cda20ec0c61aee464eafd080d
zd7b19595f8adba9c9626eb43653b93d435dd8de8f4eab4f53027b7d59deb61df54b6826d186312
zf22a5d571f8856dfa8eeec0056142a6a3400761493eef0432d2d07c5df84d7a2d8544121589dea
zef85eeab9de43ad65189dbcb7c816ef6f82c97025e4a879267b51e912aca411dc5b94c98bed547
z5a989c49d85df346a1f8ee908437d975a08f5b40404798a9bb0aa7bd460d829b8add3059492d2f
zbc853f0afdc1a65a82f08fc962744ec67e7972d3aba0394e3a33251984b26c39ee6c1cddf9a321
z93cbb20de78dbff5c64068d613055375c69f78b2efa6da747a8183c3508a2050b8c86bff78ca88
zad172bc8c3823374c58236dbf5701494d921a4c795b57b0217c1a98e9dfa650f7dd3b215e7fcca
z0c31ae55a8ee62d369de290251ed77f0b7caa6130de67901e077f286b3d9a5bfde7d3124846bca
z4f92301874ba11745eabb9aba5570fbb2dec3cd28469122f9a3864faf7617e2e552515ddb6dde8
zd5be88527ac0249f7488aa98ab3cb6a535ef28ceba44e7c1d3026b90758be9d3bc1456783d11fd
zdf164a2fd7b867a36a35efd6ac779e49527e87ba0b4dfab9bed46ab2a40ac0bce4bc1284ba03b6
z1f2a8f042f4284282e29eb7f3ada2fe652074d5cbb8c4f89bfcfa66abd47776496a0102a610136
z071b76ac56f3134d20a9483bb7ad37c9066f048aa59488bda6c90b3e0950d66548c94d9899ef00
ze63e62bac43b5bc043ff67284ba2a055cb1c5210fad588316b1725754153941555ff04fe03521e
ze1d230491913339c7e4f540e65e228a3beb05ccb112d38d52e840fa8c88091a49b1c8793854885
zf7a2b13c0beba0e46bed8dcc39e808f6ede75e05eeab131fd3434923cbe070664f32e7c0a89bf1
z76d0839c5436ef8794d41cc9156757f6c192dfbbf9fb076699cfd432fecb3578b5e8069ff8f802
z7c3749ef9d5ebae8164980be82f93d2c981b3ef498953dfd00cd8a3bd6d06f47f15ebbbee14843
zcdfaf85352f716914322d24fc3b31b6c41ca9d8c4bc05b7902eef3f6ca78ad1cb6d968960597fc
zd2e04b6177f7ee9fcea9f957f3ed45f90d3974a6cd49a03ae84717fee22477404747778ccdbff6
z418cfab0eeaa44edccb14be590db22f30c48de5c659193359df978ca33e3ff57792ae5282a45bd
zec060fc71f79814bb26b408eb5107ebaff9a5308ebca5ebf61f89a983a39d06f29041d203c7e03
zdaf31581e49382ab9d02d39ee6750de2f8d25bacbc056f7d1a695f19065fa38ff17473d0e4e5bc
z1eee595aa6f796ebc17cb5394f6e3654b99c1ddf12a13c6c6c7b2db1a78c5471d52a11b692de79
z0fc66e89423b9e95da603a8c2f18656d21a8e8744af687678b8641ee823e2cf22266846c4ce6c6
zbf925b82517781b41e5f80132c73cca5ae4e1576b0fcb1e4dc5657ef3097f23a11fbefda9233bc
z6da84565389d5f4c113e59df65b8e512a6bb64c3e40c122c8ce447a036c8560bfbb571576d9a8a
z0d2f6f530342827ea6af2ac23bcbac6c23712ae0d292ab680fb47904a0e2233eaeca3962b9394c
z7198176aa0741b62824576d951dbbdfa1a5214ac3b8140ef05c6a324b181fd2ac972b8e8dfc449
z8e151368a9405a07e68d10ec939469a98e8ffa446a100e01e47f47d37548238e95c2252112b07c
z4c7df70b397f6395888ccfc533deca1275b382bdab48dc4614c7756a9554836571f80e13206fd2
z1bf7c3fc24c4c7ac4c0bbd7d05392abd56731dd33bdbc86745fe757ce1a1d69c33409b6c817883
z87f43c1c68753b0e81f788cd24574e149945ab6c54365c5cdb24fccea126a137430f4f2468d913
z7e76fabf47750e0e4f08933a400a254dd41f8839356efd6b7d23ac5b796b6842d10796c4f36e73
zea136bdf5dc084a13c399d293341b81bf4be469b5f848706c3a24e65249b0a173594a2da875a26
zf9c62db28e1a7cc94a0f7a12a3ba12b87eddfad1d48d3c564135eb97ca0818cc26beec4b888d2b
ze15c64f90666f88dceb8e6738216d7fb02ee5f83a4435c6a2275026b8e143454504a10e15c5237
z2e6e1899ad09ee0b23dddb557f791db72d72e044d7560693116691cd4184ed251902ffad071701
z7cad2e375fcca9961be5320ca2c8fe1a796bc396d8b17b6b98948af1a3988efea35476e80cb305
zba792d8e924948142e26001097d68c69167132c4e2a30a42dfaf352279175fe9d7946e15ac4962
z6224c2274ec94b23ae8a1f72746f8a4468484da3c09d6888590e9718aed0984b93c1b54a010a16
zdccbd569543cc39d74363e4dac37ce83cb5267e6f73480a583267168f1a97ca42b393e38f183df
zcb19dfb4e8878e13c374369dfd6b49fca4701a4d03cd37cb0f876df8273ab345597df3e785a59d
zbe74f29e1b0fec21225a7d67cdc5c96b7050b22fe48f1b0314f68fe97d399a02b03de750049ccb
za1990bb799287669876b0c94ac2a63f432c3ef8cb22e6fa6ea0965092ef1e5afc98e9d952c432a
z69ef2248acc1bb4b81d317b276cad247e0b88097ebb186bdf83bf75a0b5c8e919d4ca6d868935d
zf5f78664d5ddd725771a904d0d0e2246ba69cdfc32c8c97c9ea8b5331642299352690972cbb9b9
z1008794f28ab5e5e9fad29e91b7a9df106719e697f5be8f450ca673d5b176e66a970baf226c13a
ze66584a168958d05e7aff24e4ff13b75a31589c9b0c5b7979fe52f8c55b773ceecadb0797f5f89
z2ad825871d53bc5dd764c05297986478f28ba4454ad3453e68e654c20a5f7e95cef5afb4ec3aec
z3da1bf949b5fc288a2f3e810bb44998ef3010d54082d33900a58b55abf2cd266fd8da8f6aa9e59
z180ad1af7098dd1351d5e4cc73b01e532a9c7e110a61cc567760a4d8a3529f43905e88e5da8524
z8bb2c4e110d9a7eeb207c9df881b5c7e367090714730a987a82281c1a11f01f0d60de8ead8da8f
z9e729c4cd39b1cdaccf3eb7f89c14c954ebc1352cc0d8578004433ae7e5052718c8bcc7b55af15
z5945e7976236c0fcb2aa4eff38b393ceb3f84a4df30c9692299642c3628fa23ac03489ad357511
za1fc00a4050ee1dd0a25ab41851c4bb4f504bee5ddb3c57281dfefde41bcb57a473fa96b6c793a
z37bcc3631873d26893158f2f24ddb43bf736b53c529a2957276b1c6d47a806021cea5d4297585d
z4e92f32a1f0cbf989509d5f7ab6f4aa9851918b7307f9650069e596d8c130396553305ff8080ae
z51fb172f22c0aa082473e974b4cf74c675f610cd458a5e7270710d9668113c7a4cfbd7af155fd4
z1c0b5d2e8d102d582b4cb3e688c9ccfe2d31cd6a7bfa48d42a61da2e78113cd543faccb125943a
z660fe824bf01a56bf324026249a0adcfa1ae2297a1fbb7d07c9f9dc956fae3c1c1968f977acffe
z41924385d4a3b18de6da6b9207088b140ae2d04911a44475c4f6a11719f45dda8d9345c746ba71
z8aec162e3dd81c4dbe3f118aabf56456d407a1d907a4c43d4052fac019dc89ab4b528c7c3fc0e6
zc539850806b4a795260d994e3d66d43f224db2934f32a650c5caa1dc971f115fc89873c479f60d
z81a276fc28d7253bf1ac6dc699d72fd7586f9ce94ddbce44c1768732e29155ffcaf2798a074312
zede3f333964363f1ae9d52bcb947c074abcec0ac30b966d54600197b17c71e844f1ac3f596ecb2
z00232b34b2f55e4e6133024b4478af67f298f96bc49cfd5a9139b70499813924fdf27e5f813a2e
z7c2efc89f5c0b6ee6aa8131e4dc9559204d513db48eb948fa1987c8e33252b852603e8339b6bdf
zef6d1a93bf49b1b8acd96106861bded176447672f625b2821241a718a7fe8b076a5dbf93f50419
zbc4fa59cd6b4d858a2f467f89bf2b247c8ad82d5ee707ec1b5488ccf7d0801c511d8f6030af4d6
z9225b288d30b521574fd5d487e11605f9d020fece9d3bbd3d55b7297f768a7c1b54173e19468e7
z7043392903196e354b30f2522f2443bd30692ece7bd8007e1926134ab73f7346fdd5ab35d9b64b
za0c28032ce04caa0a0c470fc44a8163e200ec133a33c5bb660f690a16b447a7720da690fefa81b
z415b3b000e16cf401f8c67c805cb4fb9bc0432e68917b19629c3de324cf9e31debd940b84c60ec
z90c140800dbe71f4e833544773d61c1e6bcf24486a6e0f3ecb47c23b053a1f36bd0e2d6c07c342
z14bd31a6de8646febad00830fe360bbfdadb3476a9982bc12c7a9fdacc280c91765854a40ef626
z685efd9c7866860dcd0b369f7aa8ad9945d0e42af4c6d0356fb668ea3172e124f02fa9b613d9f6
z95ed45e3de2b74fb2c4e59ad481d359df31ede1c9cac0c9c77f445dcfbc237031152f3183c72b3
zbe1f4b78ef0864fb1dc97d09c28ca2c76524dcb177be839f93f98d60bec40d6e8cd26853e66660
zc7ab15b361296b970155404f63add3c3a81348e4a299a46adadcdf2df69624c9e5106b2ae5d006
z94f651618998f4db0abd04f703c5266348060fbf9a1d5f27b457c263a1a74045680d3b03c7b134
zc97cdd398f95b7337811a15f708f7da92f9ba1dfbbdcef3c0d16627472e19370587c8feced4084
z4fd271842e354a80141aa569e10418ac9944a39d80125bf13db0a005212c2898558a670afede17
z189c37b415b517ac14a060f7feffe31c325285d1e76ff12c31afe5df8fc06b72fc109ef1b94c2f
z5bbff73cd98ccc05994d223441fb617ac86ffe4b5a0c07e8607dfcf8342f54b87676cd9f47d44e
zfa0d216ae2e1ed99b5b512ab3e069151511fe27dc42d7b71c803d542a66cf89d0af9e370df8388
zcf62bbdfbdc781aef01565926eb238de2cd37e34ec2f0589beec83d4011a8ee680adfeb4083090
z49d0b80ec6be376f0f2ac6c9048270ba71bbe253f94cc8c0e009d9f0ea928a6685b15494a2b7e4
z2fd56f4eb8be6f2902da474037e7544e1973f4c8f179f8637a8c8b39775e7c539973b7c0606618
zfd7b3bea52c9dffa201b2c1b7621d96617f532bffcb24a5c59bd832b3003ca4e24e3aebe56fa8b
zef6ed54ca6e7b62682c5cd33e73b4f71b7a493bedc2347f7753b674d433aa99300ddc49d98d091
ze343373f2f5f18aba609b9b7ca77bfec264402816705ed24312f8f9c2019f32cbf5564fe66fdea
z12a84b608bdf810f53a1b1fd4845dff52e1f4173912ae8b2ddb21e32abb0563e908aaa6cbb243f
z2ba845cc10f0d656adfdcc015e5283c70851646f5b3f2ec2d61b42d13b4f9e1f4d64faddada5c7
z161e927008ec337f991709882d12c4973808797499097d1a51702b2f17bffcf7496643168081c0
z5f2edb8e9d13d5a0c6c2f1e4fd1f2b6a33dd21e4db1f5725225af41f7fdd3e8b73b65e0aa915ed
zbda0b18f37c72c600be7878de64af631e774cf4f2bfe7babf46be24b6fed2c2c469c31cebfe9c1
z40ba3d61e23289bc28be722cd08eeeef6e329f33620b29d44f6764d495b1a219245e89b00ba416
z4b09c068defd320c1660acbe44f7ec7a5e377e96308c0d8a6b568afd0e2dcbac69503ee571b735
zf15d82705481ec4341911e6db3dcfeb1c9eaebe8647018fbd2d1108bde1052b48508f6200f1bb6
z00065997a5b02f9b7b28140d68b6dbb53252d03e488236c53d1192d1d108bd7eaf197a62ca9c17
za33d33c5e5c1aa9423ce47536844a27038596b0baa3eb0deb82a964ac01615f3ee3bc9d30ddeba
zccb6c43915ea0e5d4e7e57a42e3eb4325faca28261379c7d7ac2e55c72cf00e8688ce1d4788c86
z69aa5fe24b347419146549458bc6c9a94cfa14b23b6adae82affae19ce4c3071475678e18f6253
z3222cd1dcee85105fa9fe0c4340266a249736296a76d27d16d9e537f737e9f4d8a74cce39d4f58
zb702851b3de143ef7d02b93c469dbefa3766128a5204947b3b9a70a5f00a1c967a27f9e107f4c3
z93dd6e363d55742b9ef0de0a0e61e91c52489c5244674b762e7f6d251cfde1739341d20ef95c12
z0d44616b9ca9466e0e5e47e43b2c8e2b9148c0fe23fde0808785d526597869647b2e0ca6d177bd
z5c86e0739b82f99d8d2ebd8f44f08aee76cce5b7ae99d3f0a6f05aa23d2249891110e68b55bc30
z432397f01adc29fbdca11c9db422b59a9c1d5c0b765f5779269f899b6783664b74c58bcedb90c3
z5240f798c97142b43b84c94b9ce43544223a61cb74377887c7cea0bc274ca8c9bd069f72713ff0
z25abca206706986168bed77fe36e2b1be56d13d5dcb212aad15a3a79984d936af55a4ba421ef0e
zcdfeb63ea8d45562e79728760fdec15958b8906c68999bc554bfbfd6c2c1bbdd7c03576060031e
z885cec9b2c0f29660855dcd2b84e8c6450a5555433302ec69b943e10b2c07d0616aec023e87930
zf79f908e9712f6fb1dd0114e05193124c40448d80ef409a0edb4ba36fdf5ffa5e0ed13edd5dde7
z4191c93aa098c3c950817653b388fbdc04de8ddaecfda5931b7ca523787607b6fd0eb0744df9a3
z65e45475da1994ab7cdc77fc0dc3971125243ea3bca8d050b85c4618357fb2322616e95fd9f72e
zaf9b1ef290672b6031124669a7d299049cbbbff09488bdf3e2d55a29b068e29a9640930f623eb2
z69ff24916443aeb23d41f36fde9f83e46979c5645572c8d0b4418a7ec59d621e9642546d17cf66
z20c5b187cc0413dd9819d2e19b341968d7c320de2b8752edaacfebe0a377b5640d334bace98039
z80b0c4d6a97198cddf6686738e16db5c8d247fd6db1dfc636134d2c7c7cebfbf20341be9986a56
ze3bca9ffef06ae9acea10b7c9828e2f503f3368d2a207d4d69ef57cfb3c329d6d0565fc50bdd0d
z333fd1863a139b541cb29c4c7ec88b0e3e1f756afbb04390fea1cc6022efdfd9f5de4eadee1be5
z9e09658a1927e24c323112074c0eb5eb8216334368f980dabdf0d1d28840ccdf36e004887b88d2
z7667d547b7a16732770bb255a8e9992eb853d6cf2b40d51d8243e01bb0c728752f81c245c6ce9c
z3866adf82d9c2e0eaa873e2c426ecc699ea7d1a789a5130780846fb1b71fed29caedb303c27a11
z5270aabce4a5c3bb9d046ca8db75487991ce746ed347a28ddce6fb0cd92d7f7fcda409a0d06ff2
z9dadd86b99da2a915a6f27896c3533897097487ca2349b02a02688cdfe8c391e85ce3eaea513d3
zbbf83d10f86e19e243da70ce3d9a61904b39851b1b55e088f8a71d5dc3509ab7de2c48597d8eeb
z6da02e625aadb98ba46c56e31c207253ab377be298d1b9e627b702a31321eb6ca66b9d3921c839
z13fac4b6c89c621f0d60c2815bcf356b80c595a11b8f36eb5680be32e105af078e1bf58b2443ae
z03d5b6d325eaea9877988297b1746f1d29f402ab61bdd8ab61b2d665f4460c3041b4eff347f3cc
zf2b9a02994d77ba3a295555d235ff505c083811828912ea31b1453bf01e1c11ed8a8738e547dcb
zf98235558e8091f7e17a59025c3f4fda45c396fe5d84bc4bf48b95a44f92836cbade175f765835
zbc0a7b7b0e8787c1cdae2238faa92127a2f3d4242ee4545fba1d00816b27eb9c4382cc8c97f9bd
z7b3ef535fb6e3e18761d46ee449843c79d4c276e5a92ab08fd506d496fb39149d253ae06034bf0
z3577c5a7f34d776f3b7d2d603f17b5c9e8fd9084a1590fe3e3135b7515103fe1fa5f069928bfb1
z18187c040a3842782f2ee47949462131f935cb4e08b77114dd5fb617571899cc0bc4f3a166ba4e
z0ed4224f290a4e5b7c38eb00116e8bf15dd8cb3da50f4831e734cd1ba9f3d9e8c29801dae8a8dd
zc0fec5ea11489fed02b63296aa6f4635f3e1ed60ec41705e8b50bb7a705471dfd46cd04a2d04d6
zc51b7688c53dbab42ba77bc02f96c4ec1458cc3edba91553da06767dabcda85a3e153817fcd7cc
zb055ee75408dab0bac722ca8dbb84ab03dd6165414a2f5d885b2b04b0c7b151a1c9c8271732bbb
zafb4215de82e562b2293b44ef45c3643885fd0319bf79edf561131c0953a15c02aeaa000c6daa3
z3ad14faa650ca7af863a9dc877107a96aa7064d1e56adc8716bc56641276ac296b86583ee11923
z419e5e90005c6f7ca404a0dbf785c86139c957055fd56fcdf1d86c07f404d0285cf40a68ff0dee
ze67f9316b5438f31a1fa21b63448439db4f82d1b54a4f633f905abf9899089a2c4ea5103c40b60
za29d6218bcd2942d4ba3d9ba4aea9fa69fa656a2f75ea85a668793f81530127bc29a5e258baa04
z4e9eae70d413f32dfe02e5a8e68d3928f370dc799e664c57653a815e22738b9bc60e4d5b498fb5
zd6e85fdf4f3d21b77fe642045d852b88b8711e05aa53232497163b0bef89a4576bf2c72c669020
z0bb0239b2956b245de07fd8feaedcb6b0b116492c907d5371755a9568e6954cd8b749d32853096
zfc7320012985d6b4c7d96b68f95296766bbc27f7d10f5375b730027ba98131c88ed31340b0a78c
z838b792c104efbf7ca0668741eaa4d9f4cc346187fb55e14df6453b61d83eb2d403ea80c1b0535
z422ab8a7708cdd2b51e4314e4a949c503b816e4af6027c91e6587463d57260f490763ce3cde5c2
z6d3fa49d6046664afbf6b155d32c806f9e974642418086b356720d88a65cb4ad9e5ed4971c860c
z5e2a15dda9eb249e9145821dba3b7ac1f108de38ba60714ac945ff1fa6a16e310033a73836f399
z41ff2c6864961d4377b3a407d182257df53a0863484eca4c766c6d4d9bf26f894d5731b4afbee7
z1d20ab6eee71654f66c4914e1eb54caa875b96cf0cb2fd9b49e02ce73dc86f72e4f6179b7d18fc
z04018e8953ea4c2e9da29261a6fbaf177c0716b25455160aaeab8989c32c3d8864d535acb1f431
z27c8b97723997a1e10bf2c899a8e996572692770dd99a88db29425d98402682aed44aa29acfa5b
z6b32f56e04dbb4a014af44ebb27abbf776454bfcb1048bfac1589deba4f547ab4c783c6922abbd
z0dad539923df4088f24a03bc9b389bfe8f2faa5cb227043aa30651525dfeb3cb85b7877623c862
zdd9fb8413b4e44097e549b051ede7dc3843dae24538d9cb7c66210a7905e2260a5150f1749b85b
z6af1b710f6fe5c30d00e7cc82188dcdded566b4bf275e28055eca8c79fc7231dff4fc85f186732
za920151af04818d938ffd7aff08cc80f2a3a03b7479d8740bff1e20c24cd251f2838ca8292c2ac
ze5374ea220b3f56a4d04eb5f01e6090461f40e2c202d4e3e4265e045c8ac97ceec7b76e6aeadc3
zc4372106625fc7a749ad7ae788c8fedf40fbda17cfae6ce5f5c73104a86c85baf397e770d88304
zbdb9e301a499edc0c3a1c638ba1aa71c6ff9b4a82fdd81d813748ca0f3ea9daeb90f78ad36defa
zae36c7c52c03f1d0e1451e10ee3f76d34e8131f260ca1f1ba8d5b4d75afd7de62c8e36909e097a
z0c77c62326f8d171feb713fbaf7a2ecde7507fb796011859871834c50a27e288725987ac495fc2
z93e5564494b23011a28069a0f7dee46e2dac97cc9ef602d13a49d0a27ee30cf8fb0c436e382ae8
z5515683c1874d9e0ba6e851e1893f3f4ece2abc1264b11f4348e8eea58dc0fac095093ac2099b0
z43b90680c760f7d8f2d91d41ce8174c1c7764832e67d3f036cffb69946413a57fdea242343b86a
z5cc3e2f1baa12203de3323e39ceec665b2b9d6e998975b502a55ffb1bacb3e45695fd079995bec
ze03d893b26206b53b3caaba28fcb5d1a602a2edda55b3cc2182125cfcfaee8a8f0e5de55449c22
z605fe5c410ca11954c9a07ad8d887147bfd7144438631be8bb7fafe1912910b0be4b6ffb8f18af
z2b7dfda5039c1f8d98121769b9470b5c81af366d67e32076e4f89871a3e10679d1ee016c84f471
z0a2914cad4f542205a7a96f7508de60343e79ba9fcec9458967479cbc2401654baae5d2ce5b1b8
zf72fd460ff05bced1587d25205dbc81aa188ed848ed6ab7ad0f2aaa76194480698faab295035e8
zd5344945a1d9ebe40cc5f0d94c39ca82b178c286d4ed5cbdd52bdf0a1737975b07cf4419a6c0aa
zbe2ff120df3cc2ed981b0f144050bab251e9acd025433c1fddc10ddeca1f395ef2e87c010e8435
z81912986af07e63be0bc01c355ef4969dc79f567b2cd72129f36d55d0925b1bbf2973dc2bf5c33
z2439e0b14a112916ab9f923af14870b4cc9c36c6b9416f5fe36317fdaf80b95e653593786df0dc
za6978de1dc7338b0d19c044cbab87ef7d21395e8fcd4a7f7c7980dc2b6a8d593d61b2d033acedb
z057b8f3bffe41e30220d67489e405ef1c661db09d6c5a52bb06f3fa6c135c60adb15e9e4b4ec10
zf6c2d57374ca6fcfa771a7762d5c627ef9af5422e6f893d36b3e82b70020b2f8a4949fe3d23369
zf07a4b9ae785b2f033e05ab18f6e5ec41fa137851553921eea89b2c9891bec813f4c965e01698f
z61f6d10c6712dff8c013d0c8b64c984650dd0fadedf477460059af26c04f23455d4d00680a602b
z4c625fe506d207b75ebd8c7089077010156fe348076c0a27a2241fdcc23402537173b589748402
z4ae4a61c157eb69d295a84249dc065b8ada6cfe9eb1fbab37346bd37715fe43451f96ad37acac1
z759804e9d2a01bcdcda4306b8cf863489c526d9597604406c19342254ae50f25cc9d3dac258f07
zbf17e38b3693af0fc886137349a23d68e425f218f48db863e430ecc827b31fc5c60df9ccae1907
ze71eb8857f7ce6257e15a610a726dbd8e38c1d13ce605da57d306ef53d9649669482a25d580af8
zedc64b122e00f8edcc8a35e256346afeaa583a73d95b551ca68dcc2eabd19523e93f1d833a3cce
z267aec85fbb82a433fdba43a64734883705f7bc30add63e4280b472719eb9298545e84d8d6ae7e
z714ddd537c9bb8ef01f0a2ca639631c13e8e270483f5ef7ea08a4e2eb1c4103f6a8a86906b00cd
zcc82de1758722eee83c70e91f0955dc2728ef8f6cab0ae60fa3d05d27f1a0f4d2141faa45db692
z8b8a1c630410c5f568cdccd67e4faf31907a52754d2ec104ce8006fc30aba00cb922ad8295c404
z0e8093472be440b64ba4ddce37d18e60942b8849685f0e52ca8fa7923bc5cf48b1a65f554a284e
zed660c55a99541773f8c1c70ec5e069e68c6540e099143cd3e4b4365bd313e15256a510418afb8
z037ae7a947eb2df18b7e7bafa139330b9edb4f1a6b715df0a116909bb088ce575780c1e12524ac
z64cc8e71c3ed634bb055b7c23b45fa0577009c983cdc113dd8cdcf8cd71a4ed41bc22f7049ba01
z3b893691f725cd54816076c7b143cd9972b72bd5af006c3b9b67276b6b19bbb8207f5814ba94b0
z44ee43ffe7bf2f9ebf8dd20ce83da346506bb2bcc316d2b5b12b67e6843bab7b12bf2ac67ef602
z46d0764af2e5b43e5ec3e7e4b6d82c001a9e28656cb480275f85fc33f2e4a2149d0ee86bc047ad
za323b62d81064810b5f48a7e0db9c543f312bad667307f7ccfcd0c372e4c368fbf0467947388b9
z15012fd267b6f25cbcbbe5c7d9d9d7c9afd5ee58b1ed57fb354995662594a6e7df06555e112727
zabf595f3cdc79c9ae3ce4caa58801dd5b84533761829d5a3247433086ceb7a580a9abd2f6d6943
z0fa168ef99f9d3ca0cf51057225c0d08d243e3b73fc15db700a53933092ff355d844cf7bc07d40
z11afc69b1286f91abbc060781b0e9e272ea4ec5748b55c7bb156552ffccb1c833dd24697d2b300
z7392e202ef530559527b822373e7c895f76fc3a87f0fcec6a72272c135e3a91966e4a5ec057f39
z1377388166abf98d40365cd10c060c9602de033316752dd04c223d0ea5848c1eebea7d33bbf889
zb734a28c7320b325b326734a844c846551d82be53a269d5e1f1010b74f3966e4fa90c1378c2749
z1d6423a58e2e31ceee29daf5152ee7c601539fba03dae49285c4ddf9d89e9772dc57a4ec3d9876
za7b2fc31fb12e16895d10176d1cf3cf5a2a0bd6b98a349983fb8c9b2b1993a95b9298f808ed710
z22e377bd0792f0b9581fd519bcde721b9497912ca5b2caf8444b910ef1eb67376ce53ab2660dda
z4ec3be7646c926c73d97860bfa4d08da1882baf502453a1d02faa963e55e3491c0aba208a9edee
zc3cc40be0e3947a20ccd384b753d6afc2ef17cc463e7576eea142c62213a3dc725048106a74f2f
z0bcdce76784e58e1d9e3265b93a3a1e9a032ccb54678c6c976dd5adbbc0c52f10ae145eb8da0ff
zbe96766a02461dbdaa8e0e78d8389b43bcdb52a2ba8c962ad89ba654718865174896b9cd240bfc
zd79e745ccc3d3a7c6c0bb92e2b9268916719eb0203da4b115dc805236d649ad9b7ecd1ac409948
z623c9c6fe259c40045215b420bf7cd6ce649cb824047c01912dda721dfb4fdf1bb9a06bdc1b0dc
zb830d6bfd1887d0ef3f937dcd77314e656a2b9d13ec028d05a3332f36ffb8e51ff09cc514296fd
z4181a3d66b459caa6eeb93254f9da35b5b5c4b66af10cb90b928bc343d4c384259043314e25782
z0eba23292ad87da435b3b4083f8903e1ec796f17384f450e40fc831b3f29579973afbf6bb291f2
zfeb3507f7dfa99337a0aa9511457e2f4ffb12de42739cbbb56847bd61ea8c50c266631778a5bea
zac828690a21f35f41746d7e4504614bf46aef016d831f7b25ecd4d0147b9eb28f097e054a1cb32
z99c4141a61cee50104048f5f183e81d32185ea8bbcb979a0b805124690281642561bb8d78d7b47
zdd66cc6d08f3d13b6a61de396b5cbc7edb45f88407e3585311a7831e4bd98827a00d47d560d8af
z71cc1b35cfa4d87cb2c941574675121dc90db965b608a10d0d6b0b28affb192fc6d82466814130
zb3bb3b0d8a4cf4b45cd4ca4c0124c3931cf4cc227108fd8fbf1c0ca2c08e604f0dd2f42a03dbad
z288f4e4a40386ff9fd1ee9e1c29e3fc8d910076cac1e6c764801117009329716c5b9bd4e349ede
zf60ea26b5baa480982d304830e8999222e700f2f3f15dd963a83cfb7b7fc5fe696527783a07e86
zb35f63115933c049eef067a6412a7d47f4781a426bf7403ab53c8272cf2e12e71e8b28d5fcec84
zfbbeae84036935078ae4539f7fd7b0cecc1c15552d70c3cf7aafcb37d28be1aa1192f51b52e127
z9237dbed01010c60329a13177e3c5232c1e693d19be301f7bdc76292117b1df31f189b913d2df8
z7744f4aee26bad0794fb242202441804a77b25442578dec899b84d0585ee91b7e05d8661a92306
z15669e419bc1e9a66abc00ce6a311a553f8296ec44b6a24b18c33b8ca038b002050a14b12d461e
ze2da7e08ef4ada3a0561a10a716168ffbe7c483e7c80061c003738b66538003ef0b7efeabd6a68
zebe19ba0b2b7db1ead2bd028c639e6a35b84792f813129b1508ee657e8bcbaae02e78bc5994dc0
zab981d4f21fe58735a36f48d35e1a54aa9ab912a650e7c26e6c5dc388967ce5067c684ab3e2cf9
z3a2c5c9131dfe4b0c171de883ddbe29d05a14f4ac93d0111d40085c93714ee88ece34ae5242135
z53d2dbd9e29f47524c77e9ce1d31be85634bc51b8cd1356c2fc91234770d70066770cdac340f63
z8bb28d12cd64e3f6d6ac43549da4ee61b3bbd7c67553bc07f3e59f1732146ea5ba90ab1d36d881
ze1ffee094f392457d3099ee77826144a05dd6774e2dd42b8bcf0ecdcc5cd9ddc98ec075b1e1c18
zed1493e48769db018c1428384268fb956054cd7a2e1b536912b7bfddc66e0b77db90fb46789201
z0dd63e7c0273cfeb036523b99e1d40e40ff570756d88341570c8efe08c6b41b965c60fbf9960d8
z9bd21bc427d595057f253277d3d40959b97ad31fa3edddc37c09e1bdf64c1270b79c1010a4a488
z1af3641e93a6d9edf0347484d148a95f14981ecbc57e332aedc080ac7ae09cf4a2d5df308516ed
z6654f387ad9143bc8fbc67ef1b7e3628d9b26733e6d1316df6aefcf979430527d2b5e4e16c0519
zcffb6321d45f99b766354a985f4d61ffeb3fd6d9686a19135e0990ab8e6ad372954b00eb40c171
za9754b052b9ffb60ed66e1a80bbab51f470b05241ed28ec1de5a67a87691cb9d31a546412a07f3
z58acc5ef498299ef341ca012d28d7ea37a31ac524d0f9634f893532c0ce181804e61c59086a4e3
z4f6f9257c1562cd109be1347415aa13d8cd3243994118117578be74d85bf6359e07c6e31e4dce8
za25b838a2aca3027e2b6d93c36eb2e2afa0e19250f10223e2909072f957a9b67d70d65f9000a05
z1c5dd748bbd19b43e9cc138b16f166d55964faa65ba29b9516a86723b466e501763e951bd208ca
zd0d1bad31269b4277d8d312beff736cbdb272f10233d9eac0306e1f330dcdc79621f63073d48e8
z81bbe22a419d404b35f370f801388d25e6c5994b2be07f8b003d07b65c2508c665789fa1dd1d98
z97fd66819f0e17017b2efe91fddc68e3c77045dabb6df94f83855598eadff41c2295c734a74fed
zc3b6565351ef3863a3bb6ea7685c28a9b2519a8839b942cdd9eda5da106c619f55aadb9242b79b
z204bb949a651ca9bf5d736e948fe95e8abf4c1046ce9e53f3269a031f514100cff0d89c8c02bca
zc6fc2a0045344eab5605a4046d41b2339828a32e112e6a07311f264b79149ade684f034724835c
zd600d34471d725162bc76b3e6dd33147088dcff2d73b610f431ba60bce8b625cece245e544c018
z827d20bbb5219a431a1e206dbd3ce5ee62d32b147f51b36af048f18ffcd46f8a91ae0e8ac8e725
zbbd338f6ba49958f938b88a6e49c97be14e72fa8073d863ccc57681d9fd3061e410b15ac865db1
z36119dbee73680c6e491fe58234eadef26554b010f643dfc36dd0d120cf1d3e4b6fb8bef6d1810
z68e133edb274ce72cc76a0c9a60fdef60f93dc61ebed8d8a9671264ac366cf0b4f17503b4eb017
zece9b0c49b9c4edf1b1ee8f0361407ad49feeac8aeea13878c396f4381159753e2039d3b02065b
z397c616c15f492fcdd95f087b78984370bfb367eea7fdc811aeb23978a12a8c3018d2b76c9854c
z04b62b53f699991bda0ca381331acd80c0094f32dd157ec187945f7cd583052b8c08e54c36cddd
za329fb83744fa4a8979326f2fa29987104d65af94ae9c4140269ea19b5c606c5f2d49463f1497c
z5d9f51eccdbe3bc732df19ab6da49d38aa82e002c85c8acf0cf31f004c7969fc534ad2a4c261a6
ze014b2b4f02621025d58888926dc7cd53f9bec42ea835603c4e1c3f71b34df356b87c458c02e07
z132abff0b4b50e15ebe06a2e7017249883c653615fae6b1351184ff6e8a142dae947ce50e217bf
z89304d01e398a5ebbfb74b3bbea9ba129bb6e0b431b965955aae7eb096dbe310584cffa73f730d
zd666d74b749390c4eff81d850bae4b5f8f38a24cc4c8da697a7fa9fe8208f69039602c5763e282
zdca3c890dc804b6a037968386ba36a35fd79f620aafec212ccc35414077df20ce0b680e11438f6
z82869f45f9ec178dc38d45215076c25feeb0a1449ac407c14e0be220230344a0b2b2a08738391a
z84ee0129fb2bc96e0224a512df6f25b0a391bdb10e63a8484d4a967806b88538242047438ab865
z8587abace44089271bfab111c0780b98ed2d2f930c7595af13f135902bbd5ecff1d70a68622045
ze902a2c6a2a398bcb3321bbeed9e83b4c4806c9340f73faf9dde1dd1c5f380e266194ec9513e92
zdd489ca27ad2562bb4c880aedf9e776edce3c2983ed820ff1745c95c7c77988f2ca6b8f45c7255
z2a7dce3c907422879c2ef53c9cac09825a5120ef14340c522f7c5b6debbc24b86cf4209f294da8
z53ef78b64ec68de3d0f44e8989f3081223d4c18cd9c425681e5c303f6e7a0ce341b2a1ac73ea56
z210ffc5359f66b0e26200a425b2f9435fa57702c2a6d228a5af8812e8639c7db7874e6942e31dc
z8b3bdd240fe26d49d7c3b23e5600cfaea6704771407ad13a3e00d4fef961da6c4a1a1a530ab2f7
zf7187d6c4638564aa7faf8db1616abb6a89e26e76188bcbf6e914ad88c6ec7693b5d0075d1695b
z83ec717a4894e67d8dbc1f36dd2236679b2bdd7425cc7548d8cec6a47f558adb48332eb3d15a0a
z156ebdf2872c23eb1c367919cb7fb83ce8a4d8c8a4ddd84619e15a8c42e81ce95700d2ae859292
zaec3cf3b616a4c4ae79c3a021844b7755e457edcbf7cf9e78d839c251ea3597042dca0754c9727
zf75a621d8b7686836ae3444724213bb6948c1248ac62fe5fc262592a18ec66c945c3b55fdde99d
z61f85ac250368826021402710b273baa5e540b70240dff1af67a3100d4b93ad70acbe7453c7aee
z42a3e540cfdcabc6a8a839e86962d1d1789b47a96ad96a93d528286252066c9de52fef2601b761
ze1553fc89d64fa24670760f36309db2ef3f0c77994c22856c27447b1ed4e6f23d809b7e39d2c86
zdd7ab4a84d194738617afad733221c6c834a61dcf206e72b957528048445ebb8a8e9c8cc63fa43
za2c15ab7f06a1caf9904b1932ff1676c9f8e3f098ab5a51b396fef1a94fe4199d30aa4d5b99de3
z9ec9c1e4780387997503cb99d14c74bca7bc20662d41b533ec1bacb0c057d7f2aee5f081b4d436
ze757d2ef8bfa6515debead8277f432ad529c17f058a0d8fb6b988a494f8d8cd86ecf8eabe6c095
z9cd663717117ecbef1a8dea19de84303608f76bdb1c284e0c06872f74c39001e4b5b9d734f5fa4
z180098b0cdd1336570014c3413bcadc900d3c947a8607ce4ad4ee2e13f22b14956ca1fb6978728
z196f4db270a15cea6fbf0d610bf19fd441791a2e5aaa67c52f5d01f22f1556289113ef0869e126
z89bea20f595c83f8ec34eb1d0ae93a9ccbb3234270e0503886daef17961bf23bbc398cb4fee4ce
zc895f9031e67af749def525ab30bc74214175cc89c2cedac2d61d2991f691dbfb3777d9ada558a
zcc8da659795539f7cfd800eff46b3ddcba6ab2d358f79d6812ec9810b5141b80786b37467a5704
zc41cd1fbf4796e60b1323ea9fee9e8c1d7eea15c20f3202d107554d3faf00417eb2366d79bb5c0
za04bba74f0b34497c95a046a75fb5b954e384720f1083ae75ee5762121bccc0259d1d1bac0faab
z31ce892271c7c89208cb1aa09f0462d86dd266badbf43c9ea1aba030db5a9d2200e74570ab632e
za0373ec6b3b7bfd944c9ebd213ae640d90b5ebfac24eab54b344eb7fc13a1994aded808cf24be7
z84ab8655c2e1b9c8d26e5e4743d4841fe3d5b1ba77ca56b61608844c4fea07bab121f8fdb2a733
zed857aa64f7bc020c215f4dcf7aa92412a160d770e1ed11a764b3d12f82bd385822950ed83dafd
z523080cbf984c3533259a78fa7e15de90a7437f3d5bdfb458b4774aab2860866959309de23f0ae
zbddffdb0777b8033210db2913b14deb4dba40360f45c97ad22d8a8ad53e77e89d746cd86eccd9a
z96ffa709320b97400df97e7ade2dc68a840e0f520dc8c087eaa2ffb3b12141baf8edfe9e44b9f7
z44b6e614fbaa1d0dfc71f72b4d4cdf96f8323d590637cf79eb18b409f44ec2110a2b06ca9645a8
zf0c5f7e75622785426fdefdc2eb39f09fbe0beb192a695541a38ab481a80190c16c72401bdbbbf
z454f5000b3dae84177577fc10be98cd5b386e2e08f89392ab76b7f78e15e4fd7fcf6ba81581941
z1fd6b0a9428e50f7928137ae56ad6937e940ff553cca3132e1dfc504f9852a23a68d3e75d5eab1
z6b92700c77ca28833fe381c27895cbc186541346ba46ceac89956e3ac7c32e212a18bafc3b2173
z1501e8eb0cb0d1ae3cfc400af406f03e0ab1c212f18edaca010a79969ce81e535eb1bf8129a8cf
za084d937ddeedd54db7b6b64f6c00c981aea502d174b7c3c224ea52e198009efbd2e250da31bdd
z2bc6234947ef347fbb60506167302cf582da15d18dc057d842f8b79a50bc23f217e8e91c8dd414
z24f84bb28334de49cb0be1259203409948f2f4f87cf09d53c8efc004e0663bf9a4935375f22b09
z2cb05d00995f51e8d657f3d4a1c1b352270ac2d6f7b4062218e5ef52c8e0156fee0b9687ffd983
z3efe946fbb5633c1be034768d8a9953cf0fb9c1d3f8bf7a66cfcc1d606f78addcc0ce3086afcf1
z32109f4d0fb66a7a1bd543ffd9d205902ff8c48e68d85a879030254d45918ba5f04ec7c7dc0049
z602c0e9583be6bd92d8b6076a627977a892b31fd13de499e1fd376accae9e2724e878646ae52dd
zffdda45db03c1daace6e8a4025a63225037d20c2173803ae5426207953018dcebea59b8c97f71a
zf107ccac73959c5a91147455797403c429382d266ea9ba407652d7d89391189ed793688a687f81
z8402be2c87639fbb75229ac95bfa02a9cc8a79ab3ad7e655c2ddc6d08b6928f21c5bfa2ea3e10a
z08b240f08f12605cdf0c05b3ebfdf4906ba8e2434ab983435564537932545991f629aef95f27d6
z37e1990c40d805bee9bb19cb8a0a85e75a9f5102e85e08882ec0021ec748dca9b48e0f0208ee90
z28e3564df87cdb3c36c65b9961e5b09b3d353b3d0d1c9a5d58940eea85d4de42c2535a8a7dfaac
ze5ffce885e0082d2ae12ddde51599e1072ce4015694477f6b840b005b4589860e62a8987b1ec10
za91711aeb562e29fb81c666f5bde4a2ead06bf74d80456cb7c002e7604bbf30ba15fa1512b87e1
z7f7a9f7e40806689f846e72a4c6a1892dfd6f097debf7d3b17d9f244f48d6c8224ba65e28a7449
z33a3894e9f081831c917143f2835744d693102e446195202772ef23997cf33b0c7769f74449724
z1e24bbf09b82b90c520fe934c149d6c092bd5c2772ef3a3b371bd5485928e798ed092b58e3f603
z4bb9ffa606ccf5ae0108356ee546525237654ea01b54e1f595e2a73d58f4953ba44cecaac528d4
zc64a2b4ce70055f91e9f9666bf5fdec10b3abdcc5bf737cbe45cdb0864ce3cf48866fcae9e6d10
z2cc851a7cb84f2931c5ef2ca36bf0f9211d63635a390fd6d39659abe8e0039ab0c88f3d93d7583
zaebb23c200bf7966ae252a1ec23e1ac93decfc63813af55c9061870c4485b71a047810fccd384b
z236e38e1b5dcb21b954bd64c4741ab3d3f09c5bb70cddc314b9339e7998880fa17b87777c5152b
zbd29cece94b14b5244e0ece2165ed957c00606961ac624c97de56dde0201532b12494e318ff7c4
zbcb0a33c6aaf35afc939a947184fa62555760e7aa1e4578556cf8a53d7438ad5afa5a7c3082f0b
z430d70821a9459ed7d500cc3ccc4f5cc3a0b4a070d120f7c90efb4d4a5dbbb226b2d67aace5491
zfac92a096e40bb6d487c5761bd268b5bc7a4435b800e5cf2581122803cbd8f28a5d001d4bfefa3
zf79d149396a45721b00dcee3c483054854a438f8e1fc5c32972f5f03308c6a2a1c5defdcbf4051
zd2d9efa0a41e856ffc9bc19e4ce3e01ed90e993bd1757f246528e80f6aa23ab469677e5407356e
z148c2da8d1939047f3d08b1ba72dcc334212085be2cc96cee3929a224930e0a279ade071f18946
za7a9a6c762cb48ab2c2182cb7bfb538606f6543bc47a245d6835b6b009a8dbcc4329790a66e765
z75775207831c5bcf258aa16e2a61d6582005d82bc30f6c0373146c53202aab3662ee5e93cb549f
z3511f4230d6daa8c3a49573033f2177f3a7e14c828e3cbdba54c63648272e10adfd11ec79fdb97
z5dd47307a02a227b06be09c362d858d5e48e21f589c0ebe5938c281de2a99a8343564378633a66
zfb788ec2a162ae84c0e04b70024ff7bd0e84b4b5e8c0342530fb046fb9fd90e7c07db494b2bbfd
z0bd5667af35cdd32973b67639b24dbf82f9f426ff55b6c158be8a464a2f52ac8d8cbe772a9f755
z0c7e14a99d4a3f3ec915c3eeb4d40e3b8e0b6b03165a9f3b6e45c072c90a4b23f7af5be91ea31f
z7038a62ed9c03695baa64cb44e2102d1e2cd3be9278c5fef4411432e045dfa38064746d8256d86
zeec6e0e736c8d967f9276320364c9d9c79e0f2c2053ddb9e828c8c8453530e04dad78ea266d91d
z59db71613cdd2e41c47786ac1a31a4513c9f41dd0a3ba325ae59029b3079864233123ecb4d2c2b
zf204ed5f41f631a0e8f38db259e82fad32a86e53ed95cb42b398ca36bb32dd1411c1b79b45d0f3
z365eb772b579eabfee38af8cc6eeca6f73673cdc078c515d9c4ae359ccc00c2b211d693d615470
zd77485ccd640bd0b1c02e891949e696442f66774c268e9532de4a3f6168677e30a00e8e66e2e0b
z8de40b1807dbc9caed47a3530ec0c98d92499ab6247b2920af0f4e679d459de0e4f4af6adfec42
zda3c118b4d41776ed95ecac96effad585a197d626d016ae4a616be4a85b73c3bd78513c271b60d
zb246f348ba71c4e4f6d9b74680824cdc5ca7db8cec57c3bb6bfecf09cf8061d61be40bdabf544e
za805fe967109fb1a7b3e8f50496fd4bfa5650e63f2cfcea6ae07aea75e1188d7250b822f49b71f
z8f5ff0ad182b1d43193f69b0209a9b9e985afb72c058f0833b9462b0a3d4d4ef2bd0a6fefb45cd
z3fd976e2aa0267212c1c3682c2bc6e081aa2d33a2da27ea132a67fe01127ca7fafe3f6285c78f6
z9a45c77dbaaa30e1af37dbdc50bc38638b4f8262afc842e26b81700748a5a9a6e5f4411814af80
z6890b08a946edabccb790ea2fee85c785dc55a2889aeaba7896f1c1cf7b856b3001cb5a7a5abb3
zea177dbc8cfbd666a4402090e132f627a138eab87696b382a3385ffcf66f42ccf57064012fdf68
zeddda6b92000b195d3cbe4bf86fa23f826c3504c5ee0cf813d08c64a5fa284d53ada4fa8efdb93
z11e24bbb88b1a9cd3bb5642eb768c6666e8c9f7eca55164484dcdd493e8105fc87c288f7d0f194
zf17e4c98cb19608e466118ceb4a387843c027beafaef3b674f0b0751aa5563723de1311ddd40b1
zf8971ab38294a0c440b11d1fed5e0ea8609f52daf2d47dac900185b16fa98b1c221e17ad961a28
z228c535ef272d0c95ac70bac72038d35876deeb64aafaf8ab5b0e0f04e5e21c348c1fcda264409
ze71bc9af1c850fe01d560e5a6f788643342b9b71cedea2a7f868e1e183f0a0d9681620df8875d2
zb9ff335a6445adbef85bc2fc1b2e74a9b69f2fa22d713ca4b8774ec1467625ed3b728d3bba36dc
zc8613f15a9f8763b5fced582c9dedb65d971e754e37e053d15e24a71b79147220ff00f0a07b320
za1dad4b5913eb4d8e8fb156cd559974e26e9fc90ee19f29a6e660d1fbba709c14ac6907a3e1b88
z76547920e3b1d505a24250d3b553e18059cb8be4104281ccad7fb14a3c8ab696863e00a902c804
z6dd1fc73f86ce2b86c01aea5b8d5899dad55e2ca08aadc0c56ac66f3144377865c2edc5fdf5bfe
ze4c4bb621c7563a0697bc9d56ace87626d916003b3bcf446121779704ec9b6358a90136d5fe302
zde49218d30e7747ad93ff6a76cf0fb7b78610f9ba5537a4572bfff1e4f50756a96dc605459b24a
z2725187e48254d2ffba748a6fcb3f6c93546aebd99df9bc87d5be585322c0e2d1760d5d98985ef
zf8dc308fd5d26cdaf22176c303a90968ceca64d027eaf5b9d5d2987c6c095caf05edbcac620202
z3ab4321399cbdc7aaeca17b64fb20e8bf1cccea2efaf8137e3946cc462baab82ba3c4ab458f3db
zd6af7a2ec1127b2a70ce63de84548e7cb28ab0c1641018c37f73241055474ec26e9995570f7fbf
z473b31060b61dc5d5d5e132bca86004d098f44b4326a70a5a91adbf137bc7fdf7898187b6bdd4b
z04c862d1205765b319617d33a2ddf15468f84b06983fb710e83643b672d003ca460e53ae5f0ed4
zb70d5dbfa8543857bbf50bf0459193a83649ae2f13ba254b28da0d91b764716d9e9aa617ff9722
z2b331c7cf74e1787eb557115a5e38748f928f8512f01727b4708338adba7a5862f7cc4ce8b3485
z1085becdf41924bdf166c69b79ace9759a368b9c4af4448e669585565cb6f92e15c15dd2f9a994
z3f8b294494188453227dae5b46a0985516c61878ade784d1fa64ee34d519f35f541e08c1e7f5f3
z246377a82bc4ab207ef9db1416ce83a271774a49432ba28c80f86c33c59b9716e674a70907912c
zad5c5b97b12e30bbab5f73a4aaa33bb9ddd74b04f62f26a7864a0dac3b2d0eb19404ea3528daf3
zaa4ab684c2285571ff7b7caedb9b05eea14094b0505f7e8ff52c6f6de3b40cf260ac0c8243f4d6
zace3d09ed51b5a4f35768721434a605cb79e1277b3fcdcded1414ba5effd12e6520809b576feca
z3757037c00ffada0a33e9c500102056108e9e6e31c434fae1984d7a4a7ba3322c21bdbbddd6baa
z3c1535bdc9a8bcd0ce7531eaf4c69d9033a3cd23cff2bf0d421a3fb1595254b35223dce2bb72b4
z160ed5bdc9c7a6eb1b93e6d6fbe01d78be6e4140c7a9b8e8dc2e44dcda734eb543245b5c7ae7a7
z8482e5bd946af0ee8aef72b4e14717bfdfd54f34f2c8cc85cd99d0dc764008b871e15655e6d644
z6301edb38d60b7c8027fcb5989666bcf11a86916f584390c93a4310ab38557b66f5629da22a22e
zc57ef85e59024e68ec08680e758b74a702ffd4012b510f68f285045304754b58c6135ef6f58e18
z5d739d6ca2314b68589781d9315808ae8f8bae1a29d248117437daa44238507d66bc323a528768
z34d52f6943f0fdf3e196b1acf464f12f6d0fc9dc29473bbc69feccf8d22a662f9c632ce6363e1c
z35c7ee9ac7828895941513510abf0a5cf90203d64573e1aa30ba51c61817575b6dc49a739e8048
zf496c5e0fb52e5adef8d206e01f59f3536bd4e1b4dadf5b7af078567c1097710c07c89e0f1b49b
z7ec9fd2cd87b1410ffd25ee78a58deef704cb81c7a04911a2ac045a23cae291c39317ca1dbd2f8
z1bd7d3eb752033c1c824b012557b2e2ef1ce26c9eae18f7562b667b3d2fabbd56104aa92b8941b
ze23c6d34a36ae3ce70414cc7f902076197ad7d02b986f42ca6511f7d42ee94d197c71d38379e3d
z681d0d7f7ff59dd3017b1ffbfef0eeca7f2418cb1d90510a44b28e824c0225485eaa79c339d62b
z2da63aec6cd208775d8f0a7441d601afe26a5a051df27bd0c9888a3f86834e95602bba2a5ec51d
z06ed524a0e96d1ffb47387b24bda54a082232fffa1387e0a854757ea5d2f1417426b9a5be6e360
z8dcd359ce935d78b476762b32f58ffa4d81aa7a2861e2547ebf7d06266f2c97e8f54eab771bf7f
za902fdfb96dca5295bec061197ede71fa129c4d50de533d389d18105e440a6e744e7768606537b
z7618d63c562cf0bc17374fb7052e5958f39520c8ee460ebdd05f757f9322488c988f74580bdfe9
z9413c5dbfeb114e0b6461b74a3a133a9c0c53222e1b4e750231b744c7d308d554ce854c364aff0
z20fb4d6e170e9e58ccc8e37594ff782c0a8ec615fdd2854b1cde830d07f8b550357bffb2c89674
z2e08b167fee909e0fc249ec2f42ebc5ebb4efbb30a65a5c777a3f723a318af7e1cd0f6451fedf4
z3679b493e485db871fa8c945299b67cc93d99cef4b16d97404c638532b84d04f7c9a6a971e7e7d
z6b01a46db8c9b1a14a80861ced964d88fd323aa9d1c53c2bb2b5f74599edaf200311ef2dd748cd
z98138dc35cf9d60b2d8bff117250bfbb644beb110ada659cb8ecf7b62790a8b18f17856686747c
zcce021fde9bdaa1249c0a7b1460132baec609a4eda683cbdf4042302b787d7cfb2d487905b7b9a
zb890446c56d8844c85fc9c90eb5ac6776d05d42653c0fdd624d5d9a11e9ed3be99b547f00b5723
z2aa93a16f717e080f0a201798b0ed6eaa50deacd67800e49f0194c76babccbec9f742222200994
z5c88d25f722ab27ce4c6a08c0a98dae29d98df8b2abd0b607f13f2bc0671cbfabbce57c7275392
z6f305190ab6fb6a05efcea0e3ad002704ef4134ce1d4d7f3f7404030320f43e5801fd17e811fb6
z156bdfb58896c1f907329f0d234ae27468e2b88d730871bde08605d5d3c3173149b4b6829689bf
ze5f6b3a87e4c043e8aadb7e4c77bf13531d4f2722f72d990f16b2877d0ff29295d4fe39d4c3e5f
zb215dd12c61b93e91d928ca52c07bc80e8be9e5c3d85a0a6722eceab25ec09203304c823b09df9
zf4b55eecfdfd11ed69c4851e04efc778b26326da47a00f1faeca2f2f9e979b6f497026af7776e9
zf4363dd4511fd628ccadaff6d60059a08a6792ced3b8c1e97bed5ccb386c65059e87956dee502e
z196c30f62367dabe8c92e676effcffa01a67898196c263ad07c961a86e35d74fa44ab06edc7f58
z28fdc416e0cd1ccd331d0251738750b242689e3efadbcecfbeccb11b060d64d88095339e5e905d
zd65b5267e95383cef3b07f3e970848d7d4b26ad6af3d45a4fc894d992f202309e9ea0e18dee712
zb57ac4fd6c87f411f347d0250bafcdd9cb03d155a8f73c07d3797242f8943ef0634eb11da71bd7
zb788ea7e7fdd7d51746ef4955b5eea3af2ebca148fc0144a2e6c0dddaffea591bd6a5e76d4fa23
z3be4cc8b0ed828ea32dd23d701d3d0cd09405b06009c1651f07c7beb555e46b747fa8185af1993
z601aef48a531ce7af8f3a1333011ae99605483d9f2e8815ab585fbd6f4b5201e6f49795c1e62aa
z807956d0f3a43ac126f6370e23f5e95f1de6835d5484e774530a38e325a77a7938887b62b23f7a
z36ca442642e453d5225b84aaf7f9608c7a32d323b1b5b2e997e5332fda63936acf0e64e494e5ca
z0d95c99bf230b4ea6629dd4f5bde353f5fe7086dc700958017fb06dea45c83394a841e9faa7c1e
z2b271cdf8e1966b584987e37cb32e43b055c5d573946c11a9d5dc8e847697ad7a6f07501f33fd8
z40a1f4f71ba9c9187d9094aac6cbfbf8e9cd67225ccf2dc2e028f038acd6f3a18e3025333d0ec8
z1d9cfadeaf536cd66fbacbb8053accfdb4a174520761a05f3a447aff79bc35736b15338851f447
z8073b7df98f819976f452c00b9546b51e2a6b40b28b2d45c35c24cec540a623469215c1bfac148
z8869adfdc899c8651d8f5110550c13fdd1f500e9b7c6c01360a0a1140a5d86777de2ee2ff139ef
z3f8df53232152d11bc35a667b73e240f47175009d20f8346f4b885900a7bb0adc7758231fbce6d
z69981c3d768d80e952bc4a3755b5b8786df532f28c6ea3c848412a844baeb3558f36490f4e02c6
z91cdfdf8ecc147f1335dd5ce74b446a1b1937c91229c8b8c56240610af4b76f1d12ef3a3267ebf
z446adaf4b02af826fffe495ad5cc00bddc3e59d30f288a5cf3da42afc22cdecbe313aaf435aa4b
z0b1771c5217baf1b462ca467c5961d6270337377944086989d1f889ccda688047bb0bff5d35c56
z05dc50a93bd31b9b01c0a6d835ee73aafd52fb12ec8cdaea258a50881fe49df701bdd44774bceb
z207264824d9a0822935c8734d6710f12cb9f0b3a4eb3a74f968efb4163e8eac644dad68ec5c116
z85b9ebf6c42e9bc675d72dc3ec3699f811838ccd0113785c80579c1965454766c73db54c53d772
z0485db8a8ba807d432e894f278515fe102b13b965c624a505d4d60d11a66269329fcc59ff30fcb
z4d20b0d422249d39aa76bb1810a187ede1c00487730f9fdfb3173ebe7d87d63c46809801dfa021
z6e92357aa6441fadebc9b54b5ca9e6626585d8b0e16f3e465222b9207e72fc35f67f13dfdb82a7
z1fdd43416504945d51123149f4b5f917c0a3cd6aaf6561ee5e77b55238e689500c292acff16605
z29122d9f3e528310d2a412732e2440177aedfcf3e7b1596c7aa4038f19b6c7ac70a08b93a87d85
zdac12eba113922b966c5a454cb8c49848a2af59a87cc5fb6a2e490869f5cbbea0a3b8af3938872
z49d79132dc3ab3db2070aa7dda7974043442a4114c8a521972738567bd7e49458c36b676283a1f
zf45747bfe9a5535238095841960d3174e95b11381258a0efac470be4db95871170f588a3e59891
ze5a89ab96f010ca2970a49d6fe251223b2f7212caae36598f5711cee7c99f459f3efe07df71dfd
z3251fdc74a479dc0a158bff2df1ea966726d29c4eecde20b7511ea9c561462ffd88d6fb5995ad6
z0469b88a42072ad7904f4c54e39197e58501ff27d00339e25671793c8e89728c6052d13942e660
zf287207ff7b62519ffce98123747f332fbc09c1a0568d64e82696f1fe8d227f4a8ae0e5541034d
z8317b926b47c6d7a66d44c511ee8889558f51705bc22b4b0ebe356e63e7d1265b79bb5944c1bc0
zbea973dd570266759f0ff21160c5203dc641266d902115a5b2f10ba2da135754321f923e284d80
z2979a0255e1c9df6ae40c8c72d0495acf6fc52f86574313420f19fa686f9a82aa40b510a1652b3
z8e732d7c2434a28eb2b150752275f1760a5e4a8ef4a76e1eeb96555f27a3611af2c392a0af17fb
zd0bb7135e6bceb1e5afc1a28ad23752c4d02354e09374cc646145911364b20cf293a47b04986bd
z29e503dfb6e1e677238b31b76719bf214103c4e7ea9a4d0deb5bc97f95a9b723799a3b86bc39af
zc436508d59bcd16cd90aa1a2ab8eb25960efeaf2dd5b085d30a0b3413fa7946d9e980eaccda721
z43b6b3b3a8efd2847577fdd9a3f7d52f98b969596984b9482f34dd4c25b08f45c74b6d06903a52
zb4d3c861a013fe0e6420c00dc5aa5226cc2f35ff4f239fb8eabc2170a5ef3e3107c3e125847425
z0e7c1071c81fa1eeb3ef3cf6074fbc38134ab6922abf3e8418c41a4458b69faee70ac76ce12d83
z554f7bb0fb25009ab3c00c60e54c8b13530c0c8de7c9bf616d06037dcd95ffae3d53da10256e88
z4b69c3fa21ccb32681ba7381ce0e676f7c8521e65128d2ce950860b52192985559ca9cf540abd9
z1ea01e550030ec645d5949ba3d3a8580c8a799cbd3946c00de2327e5d9c527494b9ef337a5c970
z6c0ee5e85adff1a7704236673c6b9166d008e3c971c3f343d1b6bcb3d6f2e14cecdc5c9ebe729e
za3bf1c3009e6385719ca2a3c12b0b94cd4f5e6eaa6aaaf93e7a30654f8cd7a90508ec7cfcf2c96
z56272cddddcd43d8a38902072bbe45b25e4a979b10bd36a77b14f874c3239d9e678aa134272513
z714c084c3fc39bdcf797392afa4be76b14b4372521eb5e60755a612732bb67b18cd9a7d8c38e65
ze49c4ea12ab0186f21d765c4c3b59e7bbcafbd9ac1945f4be8a0374251def4b5f5cdc92aad71d6
z03d0d0e6de047c47d69bea40b6415d470ca63cfdd788fdddec6801ad3676ea8a312c45881260b2
z9a8cd379f28ced833d9c5c5954b5c099695824bdbfed53dc318bd6b3921a0e18dd1ac4665348af
z65f34f7ee930446287938945fb1931b4530c0599298db1a6c9b5b3bfd41a773ef112ee84e262c3
z688406cbe7225d6bc57fe0b33b13e67c4d7279df71160c7cae96d0f47a79a49f9827548ece5d9c
z2e61edd04bee37c3c6c93d961abc4a150ebb52af02c69156b1edc5c4ec866fa974bc1d8c5d1b8d
zf89cc6f473212b8109d0373ff71cb8c4c532b3400f2a51c4d7c8dc251ff6ac2527176f41dbcbec
z7a4c0bf9535e1a3a797b07682b76c04ebf915b447290ded357971bcfb2f76344f8bd90ed9ce22e
z872ac973fcaf080904df5730d3748b9594f6a4027cbaead8a7c378c9d34df6c6e252587387e790
z198568df687afc3647928e65d35da5be7bba18ac8a9a1f1ce93d36a469872fbcab213c255a5ea9
zd51c4a1f4a7a27d743624d5f6217ee3d8b9ee42714e44c05228a7a95fe6c981a2737105794fb90
z359cd232287ff3941248c0d0d8aaf3246cf5dd67f77213cebbef14980cf881494c32c4ba344c7a
z8ddd4a4c97d02fa9343e59417bb868b8b1c6a08c64f904995027f8a8c4e65c2ac920b7108ef5ab
zba74c98fd740bed4405faf4b421fb10aa6b4cbb51ddb176d422cc69069986c5b5704cbbbb9bcb1
z72900fc2a218aab78e149a9df621da616bef8bf19d2c80dda962ccc71d5aaa7f0a79e246d72f91
z338045da9b9450ba7bfd28c116a09086005730a12f6ba3ff44723b9a026b14e9b29da5cdd537e4
z7c090869764d5a6e1c8efa43746f966cd590899ab7bc32ea2ae276006891365f43d2dc06dc8833
z8253b1622d5dec4cf8c862da38d39e769cacf11a8bcf104c4b2ce310eaaf4dc13f2d8b5e7ef15c
z3cf941a41d26638fb9f286f053a59f1726afdda91e18f47060176a368a41dd2f6889a3888a7e31
z73b4505f0db3a7188d95da1dda3e740f6308a53b27a827c00f2b5222c1ca626daa6c97ffcde669
z6a9065de16287d1c75dd17a1d253a2b288440c02da990f52abed1dac062cba6f8a2b9c578632d5
zbd0ed8b07268b81f790f51fed62dc7f4f865ee4474a28b2227e6e4a6f434f6654475f29b5e9457
z4963257c90054f01bd2c80ff32f2010a16cbb71c5a6630c895f20004f9d04f7cb5db10315877ba
zb48ffec4d29a728b6cd517d371b3d3fd3d729088134eb2aaaeb61c3bbc54112ebe5b9c9272b216
zbaf6e14f84ce9ea3977da3ef75f9360afd9b512b9b1c8ac788e96e45f16096327204965fb44b5b
z982df8376d4480abd639ca16a40ab24473698b22f9bb04ecb7f74b9d0077d66f85ed1f0c4e3809
zc6536efdde6d5926dcf203c119da0960c6b2d1dcc441b8c129aa830bd313074ccdbcde78cc93fe
zd7fd85d3247c4a8a8b071b3fcf2d6f1e5985bf9477eeed679ac1c913a47e3ec151a2eadecdff6b
z0f50049b92d9be37f8639a7603678e4ed6e9ea088a85a0ee9378b25114a9d1eb9bee24b02ec26f
za6308dc55e746862098c2f5e69b1d9a0e6f76e343de18440179d7ad3f60441cb190492b797942d
z38d5c32516c0080aef750fa733f645530c9fccc0574231d468c6f0cedcc76ef02b10def04fa21b
z32f6fd76fa1a6a76293633ff90c94ca690f1a0e4211d25ec68a7702ccbdfc4a0d26955bc5805ec
z32d6321bdd4b206048fa4d1bcc05c2aa5d23f6237ce813ca5db56f460ad52fefe555e63bf745d7
zf19ce1565e69fb843e64b068f3f5abee6aa3bba5b2ae1b4fa042b28dfc1110ca772b8030f65306
z9c343f5cbae5f19d9d2517a80a66c281e9471451a670915c343c828d3742acda9427f231491bb2
z48d8e81b06b789228363d2f4083e12ad354f38a10fac3d9e56468c7dfc1db60727a303f332d668
z587b3a63010c1bed541ce42362c62124b2ac088f2b6b89565ea7868b200770735e732b255a40cd
zf10ea282617d01c4c21d371c52523d969e230b90c3b2f37f3fe8e7eccea0611a3d6f64f3a205ac
z7516824634d32f0cd96876821a42a2351a48ad94a1b6cd974e4e616157a912191faeea2ab5d201
z68aacde3fb6234bab2e931c5615dd01281623645bc748d10618a5ba25bf1c8c3d5d48a7b173560
zf9a2e5f2c810f4442f3d457443c3b9a7a74c3d0c75a6f66dfbce38a8ec9ec75cc81a28c42b2e28
z3a0f091a232687c11e43a9a7bdee53b52bfeb06343e93aca8adc10ec335dd362f1f87d40be6caf
ze5faef1acd00cc9610cfa1b158d04498c1686749db9ee86bf1580692d039210b8ae903af7add9f
z42e9b60eb688546cae6395fbf9238bb861a1b462040e3311356f5b0e8a6b4e54b471e60a9699d1
z7ccf2d6596e0b41bda25850646c7c5f9ececb2b2275d3d4b7eb49eafdc1e50ef9b8038a0496872
zc9aa772b88b4f7591432236d068289a82b8b15535745ab1872806bcc4ebad9fb447bec2e6a5a25
zf61498527f0d7c656c87542657d6adda69178ef6b8ec0602f9e9fe5a517cdc73d95d0977c787ca
z20e8ad20f69980b258d23b2ce07eb923e4b4bef9a6f78db832041da414a9f1595548719fdce7a1
z5c09b08c50fbf59e8842284c5d5be51c11d1640ca0d446d68d89c186153b2a4ba4e884f0f56fcd
z293f2f175449562fd72eb43d282a0fa177e0086ab0a9c5701b4f7287a2ca33cf507b2d0f80aae1
za3d65e43f879546a45765fc186b6abd86fe4cf88cbe253b21fff14ced82d24cb168bfcad6a5e04
z94cc29946d7aa79eb3bbe3649d1395c8f1ad40ad83ead66adfb98a0ae446aca7d7e5b1b0fd54d1
z5e329594b8dff29a98e7c25051d806499dd78852e7283e3849e3ebc0b112566b18a8bef004179c
z0a09cb483eb82f2454bd23f8e13f2a84a42312f2eacf09de4c90396153fed2e283a756c9492936
z9efe1697c70c7dd0e352154c3050d3ea323f6b4a965bce17ab2622fc586a2fcaf730849f14860a
z50e5064cc6e4b75507c0049c76a195b1b9cb9cf1dca6641a50c06c58cf9dc5254b274e9898d9ca
z44a2b2daecbbdb6cd6dc09d3bfa1fc8746f96bcd0823e2aa83de8f33c8d1c9acc455c2c5c160d7
zede1d60ad79f1fb3b140d5c91e8d9d76f984dcc5ef1179efaef5a6e13500f2f56c10ebb6de3755
z2893aa78befb1d0124e0e6c5a6c9f0222aa23273f4aa5be55b17b808492092cee7c476fb15dcbe
zda9058bf39feb2d24dfd2261699e23f71b888ce8ae12ab957fa620cf4af525f603e3bd5b582e92
z14547625dd1b0944749f3abcc77d323afcc6b15573627fda2f3645f082a71ef7530665df3d6bcb
zb1fe82b033acba820c3d706bf7394af38babd543c716a708082877e84fd242636ef25c88a938d5
zb7b1ec811211e1463b861b296ea957d050860a70b4439e3cd69e88fcf88596abc1fb98629866c6
zeef1e414132c4b6b9c1e6c72e0ea5acea9d1651a2398a034550c6e61311edfb9c212544d905d5c
zedd7cb5a393531059ec883bf4a47d75442c0c78864eea8c00ee1a06235948c0ac12857f65f8b52
zf75f5d58cc90aba2cca5f96422aed08066cfe0fe1c11fd9532d164fc3a7d34b4dea598f7abf1e9
z4dba2cb30e19370828a20be34b1865089918864e725a3cac38ea74138e2be68f83fe7d7d40d444
z869d4df1282ab8975b266528148db2c936a8adb6d38af42aeb3cfced5013c9e63235996663cd14
z45771dae883e54dace2a1c2e5c77751f19ea63c6d3f25f122eaa4ecd97c30dcf50f9e05e703dc7
z20dde5708f1992f5add96b118e0022c8196dac0c52a2c7225612f7af24e8699635cef55c6fe645
z3214a39e249485992df5ca0bbb7927a84378395cb8a02ff3cd5ca29b9daacb9444ce8dda5eae2b
zc6ba52fc8bf8e77351dc84e274b4571c8535efdd9b6238858d72a8d71000c55778b3529ada7b5c
z15758e96389017ccf1ab7a05c7bea1e30c588a366cc5083173fed11b0888ddb32d3c8c4999f22c
z47871f48bea3088479afe20ce774ca90fcbe9402ea80f4111c2f75cd355e8273a0868e78bddb46
z14c578e4fcb7b4e8ccd24a349977ff4eb9c26aa96eaf62df718ad5a848630239b125e558a29b71
zd5f96008c174bcd73871c738c4acadbea88ad0d73e4c5189fd354098ff15111ba7a8adf695b2fa
zb867ae1d8c55feff0e5d9b458a301de3b0f31acd7ed0704690c07adf0ac47de1fba100204c8a31
z500e8abed080a7a48c3cab7b473df4c739a454e11f78965bca7eef022b7932f89e82abb7d24959
z45001e6d6c8ba2f592b56991793e25a2aaca191564bc21ad55472ede2a5ff2b1255bac1f1ebe7b
za329848040c69479b4e1a9b0a09f4ccd1514fa0dcebbeb175fc8c4d37f9cc8cf12a58d2bd37941
z205568a0a4d0dfca26ff414027608808afd978805888f2ba06164fe1ae0aec619c276398ff3ca5
z28acd6bc92b23a61d5aebe84c9c2c18593fc1d9649ddeec3ed75436d01a40b351ac25e6be37aea
zb5b3d084ec5b738c23fe4733090a510827b79b0333b9c9dea5d0ac76a8274301589ebb77e404ef
z92c9902fddd0748eefd37222cde54e89c01ba0461d67544c655b6fb577d252c7d529f93ce01729
zc3505da767ee6fc8806f8bb01f4686dee9babf002fd18a1486323d24a8602cabd28575737f18a4
z4f2b1206fd9480e50de41b01c3a964655890425ac399527cd16393c9ae99b14480811d02f0d6c7
z88b8508ff5b9f0a6a87173d899e7d8347de4b7d41535d33a2d698d1d9ec9ad97e046d350c8bd88
z7e2e716d9a67fb60d9579dba6090f5b5d6ffa2d6256a8faf9e75b5f3eba7c33ffd26a843122dae
z67f0f0916565dd6ebe5b412717c34dc25b49913e41fbe48b6275e9afdae41b2a9667d102c91678
z4af0c55fd6ab8b12dda0c8255710a6d779d8b1da2f3fce7bee3e2ae5837af358186cdeaa43ec0f
z5b4b130038abe5231d2e02a69c02b5600a2a0d3617f9176cbbf4ce54e90d3f5623b4e495ff3430
za689c07a060588faa26a98effbf782841a36470d90aaa77fb0cd372982fc3bd9f51ab17256f21b
z6b77117f434015e112f31f7dc745d4e397d5551509fae245aaa299182161bc7180584502a619dd
z96d68266f0ef236ed5599e74420b76be1293aba01c54b7ade8dadb2d2d218ca44eecb7792c8a96
zfe625f049d491d0476eb888c74f3b9d5d8207100b81e7daf6df8c2eca7743f41afdd98d46120ab
zbae6745c35aa265382c27997412f823178877a77046bf31dbe0d87fa9b89fb05d103599fd1b38d
zb08131be67a9051a6c80add6ad9ba937a4c0a38a4d2c40108b368ff2a6254cd050730b7d8eee5d
z61599cedd7cebd4610d594df3e28bf2193b2bf40ab66ba98f436da1b6e15bed19a8f1f89ed897c
z11691a9029e1d23a17f3c4ae43d0cc4edb117a5d51fd78143fcd28e5b0f406be98fa0c505d1b74
z90158e0ea2f56f4e366c2cbde129cb256676b846a1cb7dd29d4b6daeccf16cef2ec99e6f74d666
zc5878fc026a52b2ab6a3b99a1dd01ffed7feb17a86976a4575a8d2f5704177b93f13d09d27d34b
z148a6dc3572290955f3eb430b8e889f20f9baa8bd8973296d9e0f0aca7b53cf484cbacbacfe51d
z065c35078ffcc96ef449f964039fedf048ecd4245970b563ed62ab409288f69ba23b143df614fd
z007905260bc005ed695355d5d5c056de5dfdc1aba8e3f5fd2cafba196e09e250928983e88b32d5
ze104781a4eec677f3860a90916c55582b687cb414253b89e57a82bce95df850fe8e1530d455f24
z945438cbcc37cecbda5fb6349db514d962501942aff9311b7572680e7628c6cb731083fd8a5243
z560fd63ca83706fd43c99734cb2b2d9561f463abd81ec331b20d6be041c1b99be56639fdd7fbe4
zf05b04c4f37520049577923764a4d46ab2ee6ae6ff327a19d6e4706c847ea088f5f89c46caf8ad
z63d1a6a93ac7bec87b64860f0e2735e8f97c476942c10bdda4ea8b463e64f96426a3a0a2c9a090
zfe0eb236df274ec59ccc990a5842047dd85619ff882d96642493660fc1423f794333618bf5b66f
z68bca283015d4be1a6ec7202b0e074ef31a32c011e1178a2b23e56a3aff72fdf3ddc709d3b682e
z29fb1f4ed61d72a5003770972b976c207e052ded29bf7ea8840eca6d0b7190b4177bfe5bc66ec9
zac4913e450adc273d5e4b8bfc93df851497118ccabb23756c865679b7db03dd02c02aa5eedad44
z97662c8bd8f0663f307d53e3992c61a458e0c5a465a79eefb4c2a8c5e354af89e3790f49fc1fbb
zd1317b9b62bd66f3b95c1893ca7e9e37a31ba4aea398a4a0a4f9c80c9463317ad9e9ad1d7e9613
zc3663b82c599be60adec631eb4b9cdb678eae4179612035b832c67e4684d5ce4d55fb07472d8d0
zf6ad832596c57bdae651065e13b72b2f2c12f402e05dc89b5e9732b0256cbb7c5bab8b01d950d7
zcd5d2372c470987f180212cf25d72f649f7d6f417158965ebd42fb2840c0bce95808da0e4788ce
z6f36bef4fd918e9e4de97129cab5087213a845c0327a9100bf687dd00c6d5e042c1c15bfeda844
z0fb2ead55c5c69ef951bf41a90b6dfb352924492df9edbf8648ccec18903bc8b275ea068ea7b32
z4998fc1882ae3fe80026769464f9826a12a640346961aa54509acc21f8ab6c4c59f8a9ca982d80
z4123fa72711ecca70be2c0197bc20e37504bdf3d2e42345025edb85ae1cf05bc8e211241cc22f2
z5f20519c8f105cf58332c6c421a6a32ae63bb0ffa96c176d2d53b3d5e738c22a63f08dc381fafc
zd53f160ed0f0525f0d133ca7886825943b1ffa7c191d22b000849cf4f4b1f01fbc182b6bd3ba00
z6e969657dd5a080ffac4c4f33f570d349d06428c471d726ad5f6695d65724de2d519b250b9107e
z4f1ba3c9cb9ace0ceea14b7126978b91cd7a53aed4b78bd789c689df7e93fd49c3368794245473
za69f40b81570c243b30ee65b5c33a1bfef64d82f4fe58ef79bf3e845b37a3cf2ae39b926ab2430
z20a920c881ea7934b4d78715a8a9648b300352f71cdf8a701a89739b3098097b8b82f65c947f03
zbeebf334f908562ef03c4ae02d379e64184aa5d1e4a07a2bbe4c1709137b75aa4db8c23999b143
z9e6e7e0572fb0a959ead8250b0a8ea509b8b265f77ff77252e759cb1c5511850a45456f09cf382
z3e1016a53763ff3512d6b0fafd48d4024ff6b4e32906ff8835902b5b522dda8eb8968457bc8206
z8059ac82118d3f5d3737648ddf05f130923ea4d822de811c8007b6cd00fb1627cc205bbb2d4402
zf9837ac799c65050c338cdc2e1d896fb699bba5187b84857905b3772e9f265561d1141d2999b1a
za3c0fec64aeaaaa76669ba2d182d127b89eefac5570dc4fbeae9337a0f8a3fc8341ebfc69a6b4d
zf2227292d128b5cca14e0414ccd456174acaae667ad567b04d66d13e9c81d21162f15374743010
ze584d337499e56028e3439de5db87b158fa63141e3ec8911d0f1ed2624065cfb89a074fff90b87
z9a416711def1e79db381b8d1c974d74b24a9e71e9535357f20e8498a14546f4b1383f6b57ddf36
zc9ec74bf7d89dc6a6d152a98778199639a9cd2b697d660767d57df6d8e5c31eed51f2d93ba94e6
z377646df951f74f4e85bd2ee8d46e0211e961b121776c6fe42f14f883f737eb13e873617b7c971
z32fc4a69cf9e69d36176a197350ee1a597f02360acda2435f4106c181d32374f80304b841c4ffc
z391e53077b9b4772de1d5485a37a93301c0313ac454b018ec03032725c240d5b5c6fd2598462dd
zb02a274d648e2f464eb329c7fdc3d1d9cdf1a8b0e509c4d6a1bd8de33148a9b72f0f04906d01c2
za582555e6b1e95916758b90cb62ef6256c0f9d95db41159b6c0aaa3931c89da279ad7ce6cdc331
z98337044a2e3d7451f8a759ede07c54a17673fb3d9f3e53dce63010de9c6d3eb125d9069ec63d3
zbb1823d34acf7dd9e9c5aee8f43ca0f9a82993d1625d9565b8ef27a4b35e79639e7f488fdc4175
ze580bdb468dacc42ce4709ff5baa9c7f96d83f5d9e9042f0914ba05e701348472eeab0438c9418
z5db38821d843d4702497553897e74b04781d43aa85d195828e09405e14e26ef271b338986bef27
z3c17685d7420b7b6ec67b3b9cea60d3dbe8f763fcd39bedf99abffa2b131b13bfad9d66a0d26cb
zf84ab10d0e773cf30d0bd376d29107a474001b4998e14c32c9b8e2f68130e22214fa2bf5fa8de5
ze1fcfa7b411f99ca8ca20863201372ab483e35ca2f07bdb17b1ec27bac1b47686292fd62587eef
ze47e3d4cb2044a49d76510eb67fd1c4973fbf9472049c347c7b5f8702027c6a83c13655f501360
z615b41c0bb389a56850b40ee58a36c0871dc56b41e826726d9efae44f7681b3925667d84524e89
zb595f00a8a099b5307af748ce464b191ec9894ca4658a56f3dd1ce9e8fc742934078a5ee2cabf9
zee9f5c92e72fe285024109be9a27eccc70079928a1a0d3f712d3c65899961d81db5bd1ef279dc1
zb240320bb8678022c86eb09f1cd1523df12ff39a46264553afc4b1325d9f6aab3cc2dbf591439c
ze94fab52fb4882073f0f78175b57585ce99da6f9690a09165f6f21591db7629257d8be39320868
z8939895dd9ec4b098178084e16708f422fd6746ca0ba57e49ad2ef55b5156db71c17a099505776
z21b42628ded09f339b1e3067cbf51a4e891b608ca8f6c653141d74cacb6248c655dc559d6baf19
z879a7f9e8ad28bde582412eb82a143bf49f0be48aa22372e869e4fb300b306c3dec2d100c4006f
ze04b2a0b8914c5e29e600c569940d8ba0fb40f62cdb7f615fe0fa0bb48838bfce865271a08464d
za878f0b302356a37fb22fc1747a70f2b29e99afa5b5cd24e934786569676bff9bf861e35fa3176
z0cb06506c870556bd5a73c448cbe6c81bf65871900ec92df663d6869d9ea6e6065b9cb475d01b1
zbd7c5384f16627383d31a23e4e96ef82f5af385eb6ac9feb74f8becbb08d00fd22ca3f5f21a2a5
z9a17854a64594514189571da126dc3f20cbfac514ba10b50269fed7f58a852457dd28e05ea8b94
z9bd742be99fc63fb7e2b9a6eae7ac737e80de41fa5474e839ea06dd1d137bbf3fe9fdce7f70811
z3ffa62985b3561d08fad09133c8267e503c4dad140694af827ccf37d9d660e785ce78a4056bbfa
za51eedbd3bac4f8e521b77fa38d9ef9d012c3fa7259c3331b530317b28ac7576e8a893dca0ee7b
z5429504f6b5ebbf678e875435af764065e1f05b45423d8c292e368c549f5dbb9de3907bbf9b1f0
z2d6e693033fb8d6a9f45eda73a8dd17b6ce80377f2974464880b42075bf2f291c685a019c30563
z5572e4630ede25eaec1ac28d7d0d7bf13f8d220608a6a96f50da38b6001003b87d673a5d9ba48c
za9c30dd4d01e2887551bd93f1319b4755b90adff2a0cfafcbb2ca9426567595e9e9e200c82aef4
z17ff20367bbfcba999ec23520d24d24d8e0ac71b48c368e94ac97a17faee6141d6e59f55460734
z59143fe5e536fc9fc2df36f0cb6f06c928e17a02c2edf2031972a4d2a1f1f41d357d9d466b40db
z5939ef039672749266ae582a95f8298840eb0b76c9d314f5cbdae097681f75a907ae18353e4adf
zc5dca31652c349c59d4157dc24bb45b4fca37cb8d1c1f47aa92a5e2afaeb8e9ab1333aee6f4029
zd05a556fcdfa7eeab0a8b2d5b4210ac813c59873b8826f936d285af512005e77b5f98a2724d293
z678078376820fce4d267ff49dcc51ac765cb25b3e41bd1de45a5a10704e45df91a6c11fed6c9bd
zaa311a385698ee1d673ef6fde7044c18f089512dec90aca4a51e76377fa7137d2398b5a9363126
z41233f2546d992f7df5d4b596bfb809202dea66025744637f7d14da78927f4e4af2789953f11ac
z38101fef69add56216f06de88af7e7fa87a7eac695273e6926d8abf60075003d2b319c0c239c79
z39d5c49d5d8e9fbad9e4ccf6556c1a634acbd7f8097d9abaa712d12628dae40fe0657f81cf9cfb
z98076b5d026d25de6d11651c83a114c3b4d5beb746084ae2ccef165afe29991a7e5c3cf910faf1
zb9264969cd9cfb2dfbfaa0692ae8f04cdd61c90331f88808c59c4acd4c0f720e41f85cd2aeefd5
z28008cc133d9691176b82087f48af601dbe0e9a557e2d197a9436d92ea5e72ef2129bcd286532e
z8e04157529b514e65f68d5e48dd76a2755d10fd3e7830d6022f4d14fa08216625954eab5a7ec78
z2d2e0ffa45a0f68adff944456449d8ad0804063f23aee35ef0088cb2c391ddf72b95a11bfba759
zc1a127188a40dd42f4a02bb9bf689c3f6d7cf0cfe8972f99d568664b581602d861340ab2f49214
zb07398f362024fff871ad142a33e640cdf9634bab1ea30d2fcfd4eebc3ab51a809051554ac4f30
z72d011e93e5f3ee30df62adbac485c3f001a3f2c9470b3a39a9bff15f4d576543214aa6cdd6109
z70a83ee9c0fbf29bf344fde104052ab51e2da9c362248be747a0303491020f2bf4f1b286a62c24
z96fbe5dd81f145a358959f3298858655718beaf2eba0ebca0128767c24caf40705dc5365b378bc
z58070a482e6a11374a7a5bdbce2a63ff951a7e6d3046d876aa20a2c13905bdd587bbe51d75e5da
z5d80e4ae584df9d75188feed0624ea90355c1f1b799d070736398ec003185cdcb820a9af01b1fc
zb42114cfc675860112b634840e99a4c600e2607947adc6b83da005f6cefbf87c7794a7679f5ad0
z517954bfbffc2e193f4adf491a95defd1d84760a8fee8298b6e9f781598fc04131d5efb270afaa
z90f302fce2828994cee046d287272651d7a7b3f6fec573fcdb19f16fe7bf024b338163d5b53a82
z6e03152e13e30cd830ab50813c216ced9ab4e505122dd2082c18d62c060752de6de2cd1cf82090
z575c5a5992af144338df6dcdb0036f93d33f12356e5762247c10f2010768d85e4fab656b2bd430
zee88cdbf8ed718926bd3a8a38cfb7735511d0c5cb17d3402410bfcef838435b9ed619270fff626
zdeb3fd75f361961735a9817fd51985d0fb122d414f719da3535c0ca06127147da8528480f82122
ze420914e33c2614596db0544eaee85de1084a93e580c33fb080b9bf75576f4e3dd3da53e5ff9e7
zad8f8600bb498cc13bc909b515eb8b6eb5a5d101c0505b7993c5ddd38d9ef175e18bd3b14ed997
z9daca2c73d6bf86f3feacf70fa562fc98d3021b71590c5e49d5ba4bafbf611cfc559d4d3f9127c
z9a864513978a36f03c2a5bd25213c0fe93c351e39c6e73fe39fb1a553319df5da0cd2bfff719cc
z762c8adc9b64b42dee418fa4261d6b68a4232e2d63b6d9e9ad6125b3fb0f7c62389cd8c24263b5
zdb8affbf5545feefaf7b267fdc9171824235515046ecf9aa858d6608321aeefbd840f8e2be74bc
zecaab1202e2ebcb4b6e69d489604e5cba47d737dbe992caa968ae305b50dba2d72ab2ecd7f5313
zfd2f0f15c57a8058b3e870bb1ea3a73c7e1c803a14594de0f3c9345a36c95792f226f1b2207def
z19c1d9d59b7abf002482cb36159c9b5b59f4b5a7b78ba26baeef7f00c55ff95f22694660e4c747
z768154982aa97ef9a3729eaae598042283f868f5c45c83fd5129af38686465b544280eec315723
z653ea09ea0b44e51052f58e60b3e63fe04bc2b679aa69fb7317cdaa146cb91df5682dbed12c460
z269d5c97b041cd6cffc4d3607e8504a2f5b02b2defe499b6469cfb29fe1cc7039365948abdfdcd
zcb56da7f23828fcec669355910084c6725bf45f01ec8671f5e6a2901a5492be2d125f14d0cf591
zc947acbfa36f2b63d195ba7e216736e3be6f7a7b26b09cb10a28c8d749cc3c02b49aad110e9976
z12b5ad6a04cafa2ce27aa93266b1b4b210e2f380caca9d544299b817beb10a6b6805ac404b659f
za0e71017653903c666c7ba3095561fda5a3b4aa29e447a1d55fc3f667dc95267e5a15b28ed3fa7
z9ef121c4ec314895afdf9c8a6c2ecc92c64e642cf44b18ea3fec13f871cc7669ee79ddf5610272
z033caafb0b0d766df6c2b1ea9897e53c64b04f4ccea7055c1ab2da3b0eecd6d264ffc8d61b20ae
z074359c699ef439288984dff90974e071e1bddb92038d77fdebb79c69fb291e8ed1fadeecd90be
z9b5232e56fd728c5e5c7a7b83873df4931cb02053a5d4a1c505550862e61dcc24364ddc418869c
z53103c356ac3a4b88baf384a18bb1b8cfbc2c3463a9ba44975926303736393a482403bdf6a3043
zd94d4c22249906f6af432a60d4d082f3c26d3ab66ba14872fd80a1d9091c6357fb36fd5a371758
zb5ebd5bd8f2b4efff6b13959d84c280cb4932a0526c26808a4b6247bdc4876417af0ea222cb5ee
zebf658faeaf5cdf0c653fb10b3daaa2789f1c965703cbd695d6c52b16793a5aa17d767131f6ccd
z8fabc3306c3637a69eae861a2c67cd005d972242c72fca5c6f8863b5d95973eb012c92e5dc8ed5
zbc800c59e62787bf945f692f18ca8a5d7cc1254c1ee3e0cb78cb703eeca9bbbb5394238c86f5c2
z0380f75cb9952169b2a53d666908042505c8d5bdef25aaf3eb6413da201e817e07249602d6653f
z9fb258c49ec2a3c06439ceff6b71f01d076435e408294d2262c8cc8552d909c3d8cd6401053875
z819a4192963d0f6f98705dfb92eb38b29ca9beb2d8c912a20bf6b651e11c119b16af03d86be488
zd47d8ec7916f0e56c8b27cb7812b288b7a49073e0565cc1429bd8188c19e1c10c64766df0b209b
z5ba06a56addf7863de334ee5b0becf535373ac97db062ac3f7e866d88af5f0fc7c15ddf01afef5
zc283e4bdd944340278710be5ccfb90378e60919f16797191dbcb3f86f4cfeeb3f6cb68bede8d18
zc713e68b86e0fcb8cf25d07332a7e93733fb28af48eb5f996c05f62b5bed1afae284f450d4b4ce
z51c822f6b80959e1c8ec8fa33af46a6b60f9e1241bff0b4f1e3f46053bbc7b1a0751f305eb1a29
z9c6c71523b3604ecb408f9585d3af1972d0662e35c9e11ff4d3acdaaf289ec9c51d379d3a9a497
za7b4d46dacc5d9ae3e6279a3dd9da9217177e2b32597476609415073c0636846d3ea00aa8ef35c
zb9543495751dc1ddf9c80a4a5a65bd8d009a0053ce216bd7904d6c023f943cde1b8cf7f31dc843
z38b0044be231ea96a2791f9d38d2dbc498d7ce074f6e0dc9a3c84e15541bb3ee5ed474f75f2200
za637aa3ff907214aea5ca26362af645459bf911e069caef989dadba837c34a8692f5b84a6b7385
z77332e4bef3ed6262ea28c1f65c8a929098f74e63a64c9827327df7f2063d9c5939e2b856b9ea4
z186fa2b7cd43f3a64d4b28c55cd5e6eedfeda7286938187e3c5e0a610a5177b2e872031f0858cc
zffc70a825d6d1c65ee95d79c1ad5b40d3d5506b8945e7bf0e05cb2f9aa03f15e91ed556de3662d
z84cc3313a23805054c25b73352b6245b03e052d40ad6be4348a235bdfc2ce9c194dcf3e4b32bbb
z6e906fe689d865810f2c5becfec822a72898fd61fd9313a15e8daa67129011e6c78b6047e1edee
z23cf71eaf1f75caeff588a295b6e14d637f64dfc5a1ba8b14c956b3f266e7fe24a0102e442c245
z5fd7b23becaf4f031e29ec554263de645a0f71f8baf9d3d88b69f113e768e8acd065e1105e073b
zd0be28a887f7774cb7c3f552881738bf200bf657e2a28f6f49f935dd4c14c3fbdf4f90d31ee2a6
z7f374a6ad027247da76e641609da521352021bf507da4cfb7ad8aee2903b646d11f959006fddbe
z8cdf4fa76292c84e8af267e24733556185b4be8f9f055b16908fbd7a7a090461a02ae61a2e62c0
zac1e47a53b431b98858e031170514810083aa823db11cc2516e323f92442b2b591e657b0e4747b
z2028ecb09e95608752486403328ed1c8b16efdd6cfcc7ba44e611d6a7893772748870576883f60
zc5f1885da6098d5d146330ab3d930290a3f5255f757d9a044763fdfb331440ed4f438c729f3f10
z6590b34b1387d04e2590438e43dda0b3516a2cb0ac61c3a3239265b51de6262c0da762ff1a0850
z002c3905089d13e3d4919446a3f88d94bda4f825770d617a99aebc791a01d0441c63b4ceec3f0b
z6215ed9fcb447c40c3e35fad18c96c9fd03d88e5daca8c471280164b293acc0d6ef881ae6da82f
z480e9155aa0167696490ca1b4dd33bff28346ad7090a41653d39a9a5d445f1514c7d2eb0bb1ec6
z3927b9019922376c5037836e58bf1e2ed76a85983cb7c892f6b1a8da776bc88048f2dedb04cf76
zd7ec96b8dee127dcdcd4d6febe595a96443f8107d82b94684884fd07f4d9a03b8c3386b4ff8777
z0479d7791eb1e1b8316b33ea0e040133c66c80415ea92ebefd9a281bf704f85ff5d4f7b7ecb251
z44ad70c03249f7656b6a341eededbbce545bec26aa5d9eafb1f2881a466a320bdbee474b1d8bf7
z8a3058e2224e3a577dd29a0d226846c061611bed751c3bfad78514bbce7aba74c50b3a07b2efec
z7f43a49cd0176d0a541ab98309eafdaee8ac8ea62c3ddcdf7f0ef7fd3234348b27762207d169de
z5eaaac44e87edfd12ced72b63c5cb5a8a89187b63011793843b0c9a0d6fbb3b6320de45454681d
zf4972b11e24da76269b9595ad179bfaa2fa1962fa5f294c816f3ac7ec7087f4a37a23979484aec
zbc238f809f454f545cbbb868fad7d1f8227be4aab7ac43bfbed3b5c5db74feb921c165c1bd44bf
z0e17988fc631a842e8b3e8e49a27c2d076720729c703aab43a045300f927422b83a60cb203dee8
z81d1044e9ac5dd7a49488df799e119a9f3bc37d8132223e20eb30a26d066c838d1f9940bda59bf
zfc26d2e45a7dcaefe0441690d2b31aae6143fddddb2c2098196dfb6095663378940de69c43990d
z177c5287f427863a773406ea82d5949e56422c1279c3d8f0c83299854060415f95c75a35ed101e
z86584abc9b9377f4865c800216991d84bf1b48d6a199029bc67356f3f7b9c9f68f8675a7010d6b
zd2ad5c6b76c2ee5795707e2e40e28e76f7cac6c4afd75c4cacb88e98b3781e980a265f181e82e5
z4db46bd175a5c16e1d416d6e098756d05a0cf43d5819537168380dfbd0f871dcb89f9a8eb97078
z21892c73d2dc4df83cedd014df328fe175d563532524287140873f35ba825a3630635a48956599
z19dd470647b95e63d65291657ed4ac944e63c307b03a52ca35ab58c3b79835b181ce6e102226ed
z20364dd7a6a93f5ace0a968c1c3630a3e91b117ddcf184ae51869e2f11dc7f82485b84d96b8753
z95be3889c367df011269105befa67abcaec8eecc61d9f5cc9980af7d360feefa706c67da668974
zb307b8c2a7a405a11d0dfa3f73702019eecad96bbceffe1a92cdcda86508760b40525b9003833b
z0ca90f42dd5c501a18ced0235dd1317a51f33a3cf84639244a74b63fdf260c7a992846df2132d8
zd899ae40ce08aa6ea0adff8f8578d0f228824701fdf4ae9022194d5f42950b146b763b6d9ba349
z191286492287c01eb610139e1143a20d241b775c35fcef12fb6221c966d16c34bc0334614398b8
zdfaa9463b3ddb43e502a2d438f47741a80e11b4d6125a211e0329ba0500e8c21552f46e0654728
z75405e719907b6c6b9bad698da224cbd3f059adcf54a72feb1c1dd1d69dee0257eb19750334485
z6070f13ed57a693c876bb479aae48fcc9799c2401480493820b6872ec1421d45b593363273a07f
z0582bbd0b069c7b250d17d20dd3c825be9fd937d46a4e28333d8143aa8895653bea4266c3af6fa
zb3d9797bae6e708357f821867ac2d00c9582096b65574bf5ea6af4f6d0169fac7fcfc5fadb675c
z29a6172697e304bdeca4d18a63d730d1a17183f9d805ce4ee42258b4968387b655fba99707dfc8
z9aaa2fb82d67da06f6c779a050688fa48a68721977c74eb99cbb89a2c7cbe8b37e7b59186379d3
z43b314badd7d50590b811f17f90453ce9c00db05cafa9b2952d95cafc034688a62fe251134218b
z569cef43c0a0b2fc2bde802c508e742ea3eada8549ee76b345a7f6b7641878c06e076d26481122
zae1f43854dad17e23012ad40315b1b1c63874d989e0b6f3aa43b7644762a715e48e1343b8b2016
z5634c6441ba600c4e7192bae7531f5b8696c0b2b5b8ca7f386fccc4098dbc247f37564e075873c
zb2efb582673483ab5daafc55fa4055f753ff945389bb9656eef7bf9ad4cd5de8ce0d56a1610f9b
z539a61a5b77eeb6a609c3f698c7fbf23540510cde110165ccd9fafc215501896a9b405a270956b
z628d49b155227841eecd6aafad59c67139e81dc743115cad28bf657ce677fe50712c5e6df79c2d
ze81a4e4942095cab57e6485fa86809cfb2333cf55cd08e2f7f3bc2c698546214f4bcf28b2f9ed1
z3a08aa6af4dbb4d80622b3cb8ffe2d476f8b1bbfd7669e2c288aa04efe3ce50be6845470c497fc
zdde6332cc84540f115ec66f4273ada5bcf6f314d94265ddf429c6f96b49a01e32ab8fbc23c0282
z8877ecb3651d0edeab58d66b42d0b9897343f591f8431c5368d1a529a288ab2f62a683228a796d
z55b5fbfcfb8dac195eb18450bc94cfd0d7e341cc5703ff11e5b25416e0a9be782776ea8046a92e
zbdaff91f4b463787e1f2d0c8432ef4b44e6edf0775133c7a601b293f8a803a5a8baf65df7e92b5
zd3b7a574082417e337cd8acb8d26f232520aaf64907ed85b377da0f30fb793eeceb8c6d72161d3
z600c4f8d4553b57e8648886c95d995a750a9bac61b271da16eec2e1f6efacf49f3da68aa41a250
za38252f098e92eed5d1dd300e23a18f08823aa78de5422f6d77ec6bc5d014c8651161dbbf0418b
zd56c4d935ceab3456f5aa1839c0c63680354950969629a0c0b190a97c31d5ba514b0a661f7cd27
z218ae1323843e9b7dfb39bcabfdabfa4564cb0e33a7fd0e5362d9666b42b033fd3e200ad676132
zbff067843d3b1de6770548d9a3cb8849a5ee247fb33d750cd6218cd14df9021f48a341828335fb
zc23c484b9d91ebb295933236187f0b4db9f069f995f1842cde21c3a2b7d5e5534bff3752550312
z46458fbe2ff4bb9f60bb7a0239f4dd3648c37036c4a687395641f94548235a0ddc8f31716f8ec9
z65e2e121ea11ba32310381241333d47309b997a0ad16e84525b0111683596ba962c31c79f50271
z0c7a25fba01c72e72a587ca1dd941ce462dc9c84c90a431b50cc5fa2c29f6aa073f121107a29a9
za2f8974c21c8dc5e4cb8237f572bdebefec7fe02b7b299c4a913ea6e1a2661ac4026f13522e8c4
zb6273c5a6fe2f048713593240993084e351172d04db2d590ae8cce4addc29a54ce7497f9dea429
z1b74efd3b139f2c3411badddf1871640c8148c1a39b73afc7b60b9538bef54c001825576d7b388
zebe89bac95137a6293ec797a3dc0847215774cc4b9acf53f32c096dc7cafa2faec3f26cf6b0761
z84df86e5fec72dcc170445b4f9b470bb65d6b037310a161c9ee10ab440c6e8ceca9ec48d367572
zbf22a210924a29696fdddd9257fe3997195f92e815430f86d257104b576df3cf976a7f4dc32960
z21de98d84f9e4f60caaa136354dd6a523695db70523e682d82c1a8af5f16844679bccf07293643
za18ea3a886967ec908f33d3ad2f1b3e94ad9fc0ad50008888fa9e1913895f2d781b8704a602627
z2323f81840c8eb75e7323619f5fb0a315499cd20a106a1df3817cafde93dea33a279ead05af9eb
z89c6b43f9d138881b2a8f0b23ce8fd1925edd5936bf654dd806862efcd7fe74311b6ab75d2388b
zf445add19feba7ebb1de717081853c867026e796712be942c93838e7a0f42b935b81777cdf64fb
zb27f3ebf6e94016c21d3d1a642f151c28e3daaaa48d437b22ed800b92f2e5eb92b9f79bc377c65
ze97fe82be706d5dd48e3220d99e652084db9626512e19b5cbb87dfe0d2ba502e93f568da7f79b0
z29ad65694c0b451565a9e8c9f03fea55f85785aa96cc307011edb880963516d6e6b408e94ac18f
z083c32673e8fe9bf3651db7fba5997fc8504c1d2f8ae57ed52725b396395fdc9a5afbcc48209ba
z8561cee83e636e3b0c0e7d24151c308f05ae88e2838f28717b8bdfb092715d4ec4ff716f6683fc
zb65b88cc9301363a4eaad39fb840972ed15957db2a9124afaed17704eb551d10e795d76ecc0f1f
zca3ffcf78fc8a28bd86441ff55a27b51fe3e2e177aa8e912474a6b076abc4067b7484a6d7a7ef9
z0beb78455256cc01637084df39c229b83d630f6b0f7a2fbf8d58c4e65f6d4adbfaaf8562e40e66
z476eb01df2f06a68729d50dc64252fd85b2f28a8e42d1b60d5577588415d81174b2ab3ae89f55c
z983d03bac4dde314e7da720b793c4e2020b05db796894d78cf0f5f868e31ac9598ad30a598073e
z63094f4ae79f76356ba51fa464ebfb6f1ccae1847ebc04bf39111a7e2c9ab949cbf22112ae57a3
z7ad0392b4f10a84bd164f98925af1811030118ac7fbf6411ef32658ce4c74ea9a6371e0b9f9789
z098e06522533bd6348422cfcbdaa8ff19848557b06352e491eeb3594d9caef873a036e86e07559
z8495dd89df8d7c22b2b672db87aeb22bd237fc45fb39d416a85c20cd441a362d5233e8de56deda
zee5015a269c13e959e8639fd981346cf29c2471e192219ddc79ad678e6b1edc1854e8043147725
zc42df6555a68c1aefac8c02c70bdc2d9119f14305352723b50c6dff3903ac94bd841fed6f5ca08
z090e215b4bceb2b3206efade9f5b87c1f515056dd8eefd758ef603c4593ec5bc252fb0985d3466
z55ccacbeddaf7a7dbd1791c3377a771848c2b4fe0645c641179768d5d510c4ff035f0d42b84b46
zddaac83b69e7128b9103f5cb773d224f6157fc85bd9fa5c547b0b8053b9dee1a96074a8a6ce549
zebddc0c7fdb2e2bb4be07f8042dc98de295891c86aae06d3b80660b549498f823f69b4399c0498
za6c6d6807a5e149f53a551965f4732e61d6cc2423de27db5cec0dccafd8be81d0a205bb2c6e141
za91efcb47d5b42c7bad6a040ea6d31dde74675744830c01ac87d85912e7c56951aba4de0cbe3c4
zd4d1fceb089f0527ae803c60c667139de53b0aa7d02ddc5eadf5b5aded0db0c198878f7911117c
zf9c8f40d4c8bd05a6165aa63fc82fb753fa14c6d0abcbefbbc2988b422d2e9f4c833fbb2a0f442
z670fcf6083ae22742c528dac2f0a23a45be48ccde67748cea6e33e473986a94939705d418a3eec
z12e41de441f55cb9191851ca0110f177229df48cfe52e9cc748dda35977030307367367ad0c48a
z97bccab048de8a9f8b43573cafd2d2473ac6d555d38da9bb8a4e1f03d7636f0490f9567c2cd4de
ze743d8526a55845140e8d89ad9bfa2f0fffe9209e17195105e290486656985b7e535d5a8f78d34
zda2278fc04ddcc4de6adfb02dc396d7f892805f5e0c6cc84f1c96a915725aae3d3d052a5483e4c
z96ba20c678781ea3caf46a62f6f57c28fe8fb6b253f22db32f601fefb786585f7a0d07b93e6db2
ze1d3316695496bf62a6252d4741dad5b4932f871555b48e17b3185ccebb8954bb64c16ddd33166
zfba9becc95ccd3fd4e4e48096525d403b5413b7ce2714f3d2f9009777d40d1f6c15da320e5d827
z11977c770913e78d781def0f6940c9bb8ec25a77593ef257ab610eeab3a6d76d8458d8109e2ba6
zb8e5c966ec15584ff833cf361b6c6d4a843669aa161c8c95624850dbd963b2ff32608e5a423704
z9b78d38d6f8dc00fae95d551e4c0c61c78dceb7f1731b2820204d4f1f9e1c5d11489d73953b4d5
zbcfeb43029ff8263e18759779f307010868daab5ccd6fbf0e6374e808bd690aa9d03930cb89fee
zb966676f361a8d94a6a566d6a0ca8cae9178fc816b854c5b26eddfb94742b0737b5eba263b25a3
z0649453878a24779a310cbbaca1ba82433818441894ac0bed54df16f57d2325b73a3b99087e8eb
zffa5de78ea1d6e6b750132ba37d9062a744c0606d9befea48909865be713e2ab980f584b9b898d
z2eb086481049a784cfc3ddc1616736fbc77bc650934e08f9c0052ba1b7ebfe8c55be5c7930bbaf
z63dbd88bf96b5361f29974d52a005ca051b710115428f1f9dcace224cf32ee1750f028074ca711
zd831ff9d52885eb5eae6cc41074ef0d2658e747d962ba22643bff0250758623fab3c8684146f61
z56ddf886d80b93b5fc6dd83a5f4541da7b8dca07c6455b253725e356bbc1f504c3263795acff4e
zca30dd8a940b34b2c2c266e8c1d020811e7e06d613b476e8455b86b9ad687b651308076a9d14aa
zf5d43ef1090925741d095af87eb087f9302a1d37c6d75264cec7f8b2f9c7b2e063e95211c77499
zc070c812a9a6b79270cbdc98269f110f34336228acd11fdf3271b2a341f3065cf6c577cfed5f7a
z1f4847be196f516fc9bd8bac29cd6cb16ed1bcb842656e066f188bebf8c2055d13f8479bd8b88b
z96ce1df39c6ae8122b986bea1a75fd3fee4ac0b2dddbb4f7e8ff0e8d69cc12f80470517678d149
z97e179057209b9012c1adb3764758423c572f69d1af6bd0175ac2680d93267346ce3f448c735a0
z27d2047126c04f3f2092c73cfcb724d088559720ca1b592f4ef917366522d682062bcaeda8be3f
zd4b78c3511a0ca1e2289971d76972e95e32e051b89829f614eb4c5b68d564ae25884987497a996
z99dede101abf8d859e722b33ec8e6bfe4dacbc258a3b87e50fae46193316985ce4ff8dcfc1f49d
z46906dcc82611d43eb67b7c84136bc8e2c8b4645a2d77122123b7a2f6525b3f8ba38376b2b07b5
z1f5b2bd26748024d7b9ec5c4064f513e494f6197a142f88aa87fdef7ef21ae00a63201318deb69
za32c8ae96cbcebf1ef0e06c67cf7a657514485dcdb8251731ac4792a9e15955b5a58a9c879a347
z42cee8ea6c5175c845ff623b1566da6d3f6848fef9a63b71aae152f4099afc6edd08f2c316aa71
z0553d01ccbbf9d9a16e8449a8e132be39248515491a55828f273257720be7ca24f3210b2ffc1f5
z35b37ac8568658fc2287d89c6a989a6a9416a24ea2bdc050c36151d4bb04550e092019b9763bcc
z7c3b8db5d292e1ea56ef5e74a823881e254787aefc710a9de3c02bf679af6dc9352454fa546a68
zddb06af67c4c21d4aeb8e482929d4c8918a7b167b9902a44986264f1b09c180780f6aaf276d635
z0ff658c380739a4b7c2e52f709d59a9e371bb6f41e672cbdc7fc8b637c930a09ab73d0a78e5c28
zc7ecf0fbaa393775bdc7dc6f6dc51469e1d70ce83c223780f7de3e2cb22e2e33cf1ac87203ee7d
z8898f07fc81579f6030a282d5cec5416e287fa3dfcc916d1bb0287ba3d6f81e0f26f607d435aa7
z08bc53b532bc34634bb17443ad3be7105759196f43529ff950415ccaca3ca55ac624e94c62b5c6
z34df6220a1f4fbcbfc54d5e17be83fc7890c160ae1f4b9456704723ac78bc72b6eed3481d359c0
z6ec472ccb5533c53d2b817be5eef910eba4c79d091ab9e7efb368707a4a21eac684e4c1c177316
z360c72e132c558cfd41f4a7cc45ddd0d385e68bc70e51537b6fa74ab641817ba27543cc741e4f7
zb4ba68047e9e4e4dc4f8e6e287fd9177cd6197df4f09ce1063bcbef8d0493ca364a4c2e47015cc
z3f369dc2b8194119ca857134049d9e3d1dbd52f9f2fe8d62cd8a3c26e90abd108c3ab146e9c0fa
za0f53972b01095481a72f79c33f8feb61980cc808088175c6d0f7e3a170a51742d789683c39f59
zd22049b46394d82908cb6a00640e67cf9332eb18c9b3383a5755dbc246e7680a3ab711ff7d21e2
z850e84a9380e5af8c62fb5ec1af50a5ba3977fde0e28ec573c8efc8f2ee989f5064006dddc0157
z7c26f838b32df89a5a15254277912c5503469255ce424b28c81a3b39dfd87df97079db458ec284
z175397b59aaef211d98fa329cf01ebabe152028fc6b98899482a670fd51db8abb0da3ddde8657e
ze1493a07ac6fe18a1c4b01761bddb7ee6ef59e701ffa6487df8c13599944d928c118914a862b2d
zb75590e2d198132cea9088ca9455a143a4a4e02d9b4e3b53bec89cb806f354c9e82498c555734d
ze907c9d50c1fb83f9f26c46f7dba35df593a7d9c0c958166b0cf1b2c10f080ea9ec7553cd66654
zdb0f9e3547dc8c81d3434ab5320d8b7563a2a90aaca754ee12faca7443638d604fcc17cbdf04ea
z9a73bb0bc7338b2398ad574af93c68e33f74408b16c9806ea5f1b23c225fbca3a1d94e781e75bc
zfd049871d89de0abc1529d397b20bf4553a703fa8409074c6565ace1d519f9bd381fbced8db590
z78a8bca3ae61c2510ccb160dec926893ddd8e42e379b8de077ed065e0551315ae997c7dbdde80a
za29d386eef49fd80d0de821636ed8ea320236ecdb779237c6215459789f2d6bc87055e3810369b
z54f3e19f08f3b79179ead12bf17256c014b944ff1e58b9a3fe7ce160cca20a9929b682e1b0748c
z73cfa028d562bd5574d096997212c70574efb793a9668b1ecc564bfd1f9610ab015b1f7116f042
z919c4242c1c1162952e3e4db20b41dc1816a605c4b0dc1f5a3eb795c14ea795f503f5617d6a780
z8d1e94315afe755bbe918cdcf77f1f64f221ce95d90c7c287275c3f8fb6a5fe3afad79e06a173e
z4e4646a803211eb623b28d130ff3027abeb2d0c14d6b55eb3363e96f5515c7ef52bd662f47f695
zdcaace6e9fb1119fef39ce0d8a68dc329932fe59f5fdff7d91c0ee1eaf6b3c43613997151ef26e
z4d97676f17991d75e569b4cf7b84794509f590e626a89fad5832c91951a9cf7375c5c1568479c8
z150289c1dd42cb2fc8d4d31583ca67ac2c11c8635508865ca54b252e99f0105edcc51a950d1b8f
z56d2c8f299a53c5a3a6a54c9b965ae540f21994a4b160bcec87ee395a8bcf3601fdf7704937f46
z8179e2a069e1daaaab7ec2208e5b1334c125a2b04a1d76e025f3dfb74bf7d3ebbee48152ecb782
z25f8193929ee0578a3c9f4acb4f38197e7da3ecb539553fe3cd7badfb2123197ac0b61b92816af
zc31864f9329463d1e1850f8ef28b2718732946d7c0b660f0f6d4c974a32712b8687902cc78419e
z37c73ef7c02236ec0e9a053c9e742db5ebbb50318354e24bbc5ea4fe65fc77572c4a91bd31ec8f
z22ec91d78f8745d87a72efcb96a4e14158fc9fe8c091d4a5ecdb550f785a4812a37bc1db9d78a0
z64dc10a7178a41c7593b8f18e706f9250928729641a3671f189099456c0b6496f0b8031e8b4fcd
zb28a3075e3e50334cf2dfeba8d0bb7cc8357e2246572ec2908bdf368c37bc8e00649f57c6255b0
z1c726563bd07c3358c92fd8a9965805f6b32fbf9c74fcdcb0231e8cc33cba480d757249f7ab36f
z44ba42c87347d8f0840879c2c31c7fdba6db44e25a857cc9a7e24d3189f850f801ae968a27f346
z8f58cec0bbab891627a42c0d3094896b326654cbdd526b6b6975727c53710a20e219d0567ba843
zf9b203dfe7f27b2dc6748f415a57983c789a7755bd28407e1b5a8195d4d0514c05ad00edd2d8bb
z4b9c3a148a0e26d25240aa0676873ae696e80ca0278cfd3a39688fb1fd584d551493026b292e68
zbbac5738ea06bdadc1e67a77e0595516297b3d1e69b1bcc18ea7c508d75121527916a4f173ebd1
zbd93ee50f4168b0b5db97d838bcf5f03dfb5d4355fdfeee00bae9d48a03b5b9ef75a545f996297
ze539ea0e9417d37a1cf8a050cc5a2f753aa09381fbb65fd2ea25fcb9ba5d61156e5c4ef154fa26
z0a2223aa4f245c42af173aaecdf4fbce9ff04c45ed7e07ccba75548152b2c9fc92b44b50bbea43
zb83218b70f42d27595f196d6d6c54e2388c326bed8e01c491a6c0c4dacbc04e33bb06a1dd30055
z19a2d7d60c8604ab8d58c861640d904189bf5867389f15f5c7d3a0c83c814e48ebd35a42514b3b
z5ae166f369695032dd37fd178189fc943ea5362252a81e022b1310e8b19c9f8c82bb2096b08e30
z3bfd74e71438c20caa24fa6271a707945ad925175cf35d7cc9454d4688c4068044f7d2c2722252
z2ea659040b7d508d6b484277e956432d89d8f3f5d5a24dea499a86718488191e7c718d45fa8b4c
za5e9a152e4a3356556b9cac2c225377c0a44344898c165563920b2ec1cec1ac8d4c380d0e37c5a
z00b72fc2a0a747691683718a9c3c653988d9a3492655a48047d09437a1450930fef5a56f922c99
z19a111316f6b518398a03b53777aad38e885b18997212a91d04976cbdfeb72b1397781984a9f24
z87646011cf81b074cf4783b342ba0394b7af95b69e17213020b0fe4623e18ec5b020c4c9d37655
zec62f98e15bfee1aad00be3731ab5d2e4b4f85a1880ee13f1c7ca6fac99ffe25584611028f55f7
zaeaf56bff934324ab000ef965ee971e0672a0fcc8b8a0792e796ac73fc09dd2d27712f2bffe551
z41f417a35e9f933bcb14247223e83b53ca2818393f1031ea4cfea476f8124d80d2fb817d49c2b3
zdc4493b661a22e4b8c28f804a2eddad8b2c073be55cbf0d1b8d18d77e7b065a15f0e0f8dfa0288
zf51e2eed412575f58f06e061b4f84616968038a511ef13cf7660b8a4fa7637820673544f0ec1a3
zae2e546d8b7e351a32b199ffa86f827068901750d85432b69c9a070ccebf4f498b82833d5061a5
z3ab500708274b2cf62611dd76be72e8138bacc782857d4efa76a43b1b9c7a232cfe8ab76bc9bf9
zc7e21325bcae6b39b79807ba14f04c2baf1841a273e9d5b664c241358323ebe0ef9eb4b60ef3bf
z75d819cb3da4fec0718158b34c497f12f736cca3e9a95be88f467e66ad66ddbeb7bef79bdefe7c
z8e520ebf39ec46bb5f815540544073394cdb15b82092f6048cf80643063271dbebc6db8cf19ddb
z35932b800a90aeec0a535d968adef19a9505a6f540bed3208aa288679cc2442052a19290b02b69
z9ea10d1c316080188a125dec57cacf5dd8439aa15a9c39663588af64fbaf046c4f5548e5c9da29
z1c86568988ee61cafd614ae49a22ab095e1a57f702538d2167533b8e796b9b75e6105bf0bdaa10
z0d8f04ade3a71f9913045482c410016e1fbed0d3e19c8dd894fb3dce35c406505ce52072bb02e3
z93c1d792d334207d37254465ec1e391ab4baaccd0ecc669895c1a21815d8786905693bd7ecd7c7
z0d551c1570746fd3ad28271865355c6fe311a720a940b972f1f4e50abf68a835e9b5bf3f275068
za1c38a864463728f007496868f8a9935367b19c6aceb5f6c67c5c0f9978bec6add44653135a2c2
z30aba7ad77a74e4963615e54429f5a9c2859f9e86ee2426f2fcbafe0fa18685d943158778c2560
zaa5ffdd01184266a72a76c5cf9bb9108ae393ee3919964145a2c0263bf2f8dcd1f37274f945050
z6b20376f40deb47531784da3285f73602da190641f418dac3f378a486468fb368465ff257f41f0
zf7a9d7c46195abeca459188c52a745d40e6f55ce65bdc5579dc1389eda1de233d0d256f3622124
z4bb67a3c5f86981dc55ad22db0045b116ed1765aee2bd38c9308fcf12d6793f821a0b39214c13f
zf25eaf3848a96e1877f261aaaf0286b9068cc737e648f3b366b4f7315a7f5f5165ff14a7bd286a
zb10411df9b1ea88bad35e1b2c42f85a534d1374fb69c50df9ab35b161038d46a4c77f157cbc740
z53dffdda6da8afb45f059c4ad4fc866586b0ae34561d54d9e24373a2116eebaef2faf0b8b8da69
z470b5fd05df0dd7b54756c09c3eccbc51d6cb9524e2632639cc29cdc554f4598aa7cb9e68127b2
z41cc44deb1c6d5e05b2b652a6aff6409033972b2150424173a9139fd5a848c8936614ce2e1a967
zdba12be79dafcb58fa50a3201e9570898b45617c456ba7fb78e21dfab6d5efaa48b0f8140f8cdb
zed1610eb770a45a2edcffd3366fed13baf73af0f245aa37b7acc1378cbbc3cd90086fca70d934c
z224cc3f0de72a51307c2c9c9b6219a0eb853f810941343919d49e8dbb705e5c9c6eacf12dadc37
zf9858d0b55970bc4c82dca396b55d1e07d5570df1aada9e1d34ea671650ca06262d787755acd2f
zea0b114aaedda983953f24ef74acba051634389285c4ace17f51270feb46d320c555bf26cb4d3f
zd530d7930bdc89dd2fee8e75c376411d86f011d933a4b60323d3a97ca3831eabe3964334b7b2a7
z6bc0e411c0b02ff12273fbc812259359a2a05364a43a302723c8bd48fcec6603d8ae970a18dacd
z30988a7bfa5bda6b8513979693e2ab6479eb2a6734274492a0be9d489a5fab930b984b47913d8f
z4404046519303767690d3c3b4d36b6b66867853b50af26db21c844f6959cf0dd4cf5d65ee26fa1
z8129e0444518ea942aad08a5241142fdebb3cc742db1a63002ef4b3c599e0720a8a3d549c4fc57
zf9f9e5973fb60a1871403ef169c3600feab8df823305d0b46558b757050193fcf9560d471dbcfe
zc92986ed19061c6f610edec412d2eb87ebc665538f5faa15971160536655357b0632b5c6e31af7
z99bf0c18de20adb577b2056b33ee4e2ff55602c24ff054416cb3d1f0c7595ff28ae6ae500a6b35
z1da186e994c4a22d4e03594e2a9a789af63b22123dd5e99b0bf4bf63fa4454163210e818865362
zd3be94c2e0fe5c3eb244813079e085e98d9c04acac26a26cab00961e7c65ded31b33a6a639c8c2
z87a9e40a28445950bd76ac0fd9f4a013206e31f7fd6c4b14e714e5eea2141912d007e64322bb12
ze3fc5a91965f631b783526104e97a255544a6cd506f88f1bc6db24ffcd5c0b63de50265b49a76b
z734b6b477f27ca4b5237625d27daeaf72436620331d9aa6e7711e29f49b3314039aa7cc49a2947
zb6d3124e4ac02acec53165dbc658be4b635176c4951b4e2670543d97a315b665abcc570155b26d
z4a286c9092ce213fcb4d3d49d365ec43c3aaed9a099f23e953b917ce056c62e7aed16ab6671071
z14370887dc1b891c848a9f81f05a726d579ff6340d9b44a31ff32401ea7f0bc1d87db22f320d1d
zdab487e3f1ec5e79bc9cb8c4f14ffa45dccfb75c2075472f162bea96e4f2daa6c746a6587aecb4
zdd48661ef4951a0a9443467e073a4803a58739a3eddd4688d7f52b460cea856e3d2c4d8b2c2def
z865161650a690cf93a72f5203b64f4e7a53906e28e9e0c12b26600911274d82c2702134c027eaf
za497223c26980a12a93676f6df01e1e7b2f8a7c0289983c5e76f79fec80a08a606f1fbd323faeb
za669c5494fbd10aab0c17512b9afc219b0f643d5ee3a6cf528fbd8cb12ad2c2840ae78ab037439
z2cec129b32b515a904cce9b3a927f0094f709c57f1c1f613327365f98a3e64b0c4767fa4804813
z5ed451c34afe0610506ebd5ebfbb5a6e3151003b5025d692e1876feddf525f31463f3c5bc624d5
z213feb4833b141614ad3a81617548dec6ab1c3649bdf8f5c9d9fd5092ffd2ddadd01c08b94507b
zcce8d5f0bfacc65cc8dc899568b5840a6900b61846a0e5f466d3fc10707d774c213e0aeaa83abf
z202e82937cb1ca80f22089d60b0e5bd2bda7255a6d3b5a3d4668ae39b73b8c599d41a95592dfed
z5c86cfd79cd2f28ae093846f68cb79e2c4953229baaf9a70d0206e28fbecc734015dfdc3296e6c
zb936b7bde1de006d992af577dd418f4656e9191c6b95396d01bc9023bde7592808dc0c94661db8
z32a8f2ab73001b7b1185c58099f9a13495b4bdb33bed4aa11b23c552d58905b80eda2366a4f6d4
zeb8c43ea6808e386e36286b56e1db794ea58a1487447e0eae9bd91ba2ac7614f2960276f5c5a72
z93d946ace3409c542143f392c50194d9b644798dd6c8c108406b96c4eb12493c80c7b5d2457fff
z5ba6c722a743dd48274aa5385ba19a858ed8f7ebfd51cae4f9b0ef63204509d4458ab54c7937fa
z315f53c057b76390dac7f5e43f95506e3c2184fa4863f3a61fdc5eb65c4349de5addfda532aa36
z2aac263a4b1463b584387f5d532cfef20a3f282023759c7d95276cac4188c4f0f3abe0efce8ec5
zaa4d13fd4af1552da6e784663108d9dd98fff4a06ec0d64c9e6632fc8d80a6da8b60d19f6f900e
zd8db082ef902604fcde1a9ff7ed05245c08f3bc31dbb0a3bd8074ecc2e4355b3022a90b33c291c
z82fc458d5640be3651db2917afe9cc6d14aed8228d931e9b65e50732405818592122edaa323f25
za069638f9357d1cfb41b079eb2594e0b1cbe8bc3a4bc92c929831c8f46fdb9230189ff6d62c262
z20b1e11ebc9d19f57c26986cc37787ac5f8de83d561a3c11de0be7b00f82127d3b2ff64f096cba
ze1a76b277fe82eee204675a37a0b8897416cbaa04925626ba996a26dd81e2c00d9f24efb1dfe1c
z5f57fafac90b998ec3aa6a2a3bc16d2f4eec27d7249cbc183ac89f83eb5cd157f01e337dcd7c38
z21c4364cabe387542c5a86383406e20f1db26f9f90df997e8bc1355cd2b86f857f024fa418ad76
zaf4c02d0b2554bd119cc1e99b8bb87736e85271a6b39a89d8fb726984dafbc0bda44843c59be7f
zca115128772668763caa5e07336da831e2a5c58acef4903efd5d7392b48b83092521c3b090e15c
ze8e85413ad4afcd918fa863fc2e026342f8f0a65ced03ff589ef120e7215e86743c13ef3b6a720
z8bc53e3221d00584cd9d45c2ea6f5aa854c5b3d7d20681f736d2908b3ece4fe9bcc054549d0d9a
zf2f45ffb885b59fe3606b03358e21606546d0e767c13410b94c6e837caa5599c5fd75e2315204e
z510532fc12412ee777938ce5175a157447f13cb35d5fb0d1bb791421396684a0885432eb3b7a15
z59b3710822727fd3912170faa5bc5647649db8dea331b5e9a920eacb161db62edcd307983899b8
zf998846da8c8aa272111b009a40a28810487bab41f175e7d7ef9fa21f7a321832fd82b44f8973a
zec2469d53fa1fb5c5a2d8c216931e72a4104f71a404d255233bc469303eb2fad1abafe09900926
zbb4f7a5214ec357ce6fc424ef34eeac6b2139d4ff4a18d0d262814b2aba2b17ecc7b2ebf05614d
zb95299d2a8152ef506afc8f9d6cf990fd73e8a9fe280ae799d37c7d94f4abed84656f3358930b4
z0ee416435c5d2b2f01250f4837c72617f465a3cb594153417f8cb314bf902ab4931a6415e7146f
z5363d3f8f9594ea246ca21e34d05c55d1ec473e28223e453aa78be88b7c962a62e5eaac7db60cf
zc66532544422295759e96c498734aa8a1aadf7e2ccf5590b4ab1636e670a0730ae0c73841c0d0d
z940183421370f5f31e5c60754559cc874221f59a8a3652a20ee77e50ebaac82556f074c2ad9c68
z199f6a4939d153fb07d86053236af703d6edb9abb2ac2b6fb1c1b55ba83c3377274a8636401c08
z03a9d468432adb37cc0a4d849df607cc2be28c5c76fc6e99027905805e62ef96f43f73f9c5b96d
z1c94d932f477500d8ff1a52ac976d9c74c6fb902facb6dc187831ebc65b51270a7e9caa89c8d99
zab6b1b5f16d2b34ce287a5507c2485f80067f8fd54de9dde3f0fe390254c4dfd77d4b74d2ce754
zcc7c928254956f436aadcf429dec518ffadf835813fef75f5d5e41e2c5feb7c89fd85a8d869b81
zca940e6d16dc3286716f355aba1d2a66ff34cbacc24dec02a9fde1a43f6f89a065f16e03274dcb
z8c97caa04f4e85d1351a52946446fd48d34d183dfda1fa2814f4368707af46723fccdce8c699be
zd49e66dddafbea76dfc6ce5c42029706d4ee1917148455dedb3439ac744ac050745e2e90421afa
zb1e93201d06040ae2535a4d397145d4e9025d4030b477d7aad2b300d4668f4b0d5f0c2a3f206c1
z18f51f0634f78d8bd796aa4d01d98da5b04dbf890b86049efbc8e8c294f501a9cd90ff63377496
z2f90ad08a134d29498b70e5f620b3a75c2032c0cfdc0c36b0e69352066b8bde20225f71d212b86
z5c3d5bdb99c1ead9eccc6581af3932124218b4a69984d0d0d1ab0c0e1267bc5ed86b0d8cc1404c
z6c30c3e9252d50dba101e9a40c4cb8c4588234e65a919468978ba2d2e9dd8407cadce8eef8809e
z9a2b09a647b87b02cdf806d61137118e1091c0ea9c1ddb35f4a8324b3de68acb8e8035c794178b
zade354f2016bc265d96d21f94e5b9111093a0cf78c9b24af29d0f4d0ce2c464dda08c73a66ac9d
z6aa9f137ae955be2e195f965c0deebd6d736b026dcb00edde139cb89fc35861cbb931bd91d04a3
z58c1365d130a832ac8688ecd55879cf36f92363ce30714440226ebc919c839e6574e5eca9906c5
z0ededdac57e76c2c4f80b5944b5e7044834ce62d43343628eff3095a9f2fc7f4c51b55d6a60a17
zb4c0c7d869e75ef173a4b0d9293538b7925c7aa99a1e340a9acae8646e7554c43e54a75afd4179
zc34861dd0aff9d049f6faf2b53d18a617da62028e0a6b8485d6e823b479f443b705b10d297ed97
zac68c65ee4209328735915fc97d55ce60e815e03cb2c3e87fa9c9d7a803da2659d486a1d6732fb
z894438ed3094a323c5e8506383b199f1064b018de9e6962ccbf0b5ff3c34b6a5c72cef6ca49b8c
ze28fed53524d9e350ad24f962391b84462274d35b9b76577fa5c57f77cdcfb034407b838b12d1c
z92443a4d17e22ba46a8a5e6bee5ce1d6fae98b97778254cd5eb19b1e5a5aa8f1d341f7b15aae7c
z52620a73e8c3d73c5c8cc17e2b52a9c627d0b4fbb9aa7f9ea6a7e77e0694a1aa5a28fbb0f5da63
z334627cbcc7a1fdbb2ebe248b012f0dd09587613241c9ff86fcb31bcf2707524d4353f2e2720e5
zf3cca0d0b1732e4e72eced883d8c24a0df6b9c2523c75a0963e4a7bdc21b3ba43a2ecec5864840
z4a77a1d997a3028e51bf14e4cbb928221d6fbd019a25c466554baf981efcaf41866039669e2743
ze274d1659aa26a63f852c4cd27d6afe1b0c1fcf202740b50522218b74da1bd3676b851408e076e
zc0c31dcbd9526060f70ac429ceb5ebd062de8cbed5abf461b55f519c7c4d2bb0e1a271b1a743d9
zcb3927576f69f7048c1be5dfa3d63fe8e78bc58c18c797ff6f1e985a311aaad59601df82ceaab6
zb7d4230af4ae5b23048b20cda3bb04fdc8edb0e611c1885751fbaf917294cf0dae159236e58f9b
za82a0ef9710cadda56a77dfdd06a612de90045717a5160a0a9a4f4173f3649ad6004b7eab09c6e
z197a011c02b20b428c6eb4d07f7a845dadcbe6a3b8e0227ae934f6f2d1d79eb040e84f6dfe8328
z704c4afbdb03b6d822f9cc5e13cafa40582a321d7f28c28ee0785238991020bcdc19fce059a253
zf27db5f9215f4ad660ce95b97aedfd81ac5fa59173d9a1b970d3867387f49b559ee909a7dfe4f2
zbb00ad6d96b524b3e089de840450b74ebf8bb65afa621dd6e0358725d402112638738d68df23ec
z56ae7ae8bdc3410339f93a4ddd376a29f03886fdd4728faed00a03564fd5daefe8211423ef6c91
z085e54158c80b050b4b5029e8264c77872008ba61136b4ebf6b0aee759a45e9ffa4a9ac945a775
zfdea76a83893a18ec8279ad0e87f18cdb481aab3dc06e6408acc120f46d13ea7e56bf9964d78e9
z0fe57316afe02fea9842ad347059f4dd8741c3a3064f407a373562203ed1ee8d4647ca309157cb
z4e53a1a8a451dbce570666f53d8fee4aa44c56494e9563bc56da613884fbdbaf50fee88cd58171
za80147dacf19bfaf09e704c65d8dd10391c9f3357b9a97b363ad6c3ec03a557b1e987d1433a09d
zf4f6335eb7a54e3025418b4756c58859c0e6348e501afdf4a1b48d63945c58c62176c0ff8dabee
z35f7391dbf79752a34ab832276adfe59589e519285e350546a4274242bf62715f3e243dd05f4dc
z689950b0bcd103c8313c4cb2379f8124e97523ebf226e92311fbaf90a2cd7312e4508de718b1ab
ze5b66a9a1875bac13c990d8748b208e6706762112b1363649e91ead3e21b422d1700dddd335078
z4d02e613116aa9bac756e52dc5b3cb82831d6a37c7d633f3ff2872a051f0c3350aa7855e4bbeb9
z00aa4c22a165fd9e819618793820067ff20869c95a9a89d236d1f8363ae4e9e9330f8da41f6f0a
z04061aced401c39a9c6d84ac1a23edb875f88c7f514fc26c1627f06b0c77a160d3fc64bb3020af
z3803f80c5698c73b6a19fac18e4bb9a4ffcba884951e611656d0a7ed7d3de0ae952aaf2358bc62
z59a012150917d025628c6132319a6b9405a9a984ba0063489b6e2610e2a919dbee4bc3cee58036
z06dd7e6f4eb209fc282e97b8155af34c9ecee8914e115c4e3154a7fd6889389920e19821380631
z4a4f0ca2deb48260f47562afb1105548c17c2a6d7701b24886208a317ce0895776a2a61ec3a689
ze3110bd49e8d8edcbeb587e215389d5f2667e325c3fd94e9d84b6ad27b5d5d52bfb164308135da
z4beb88f449f06ca2f401c2b53f3fa127b9018450141052729941f648298e82d9cceddacf63ded7
zc31a2169ab3a68dae9262464231280a7150d4a5ad6968f8fa4eb23e692f00438905a33a13a9650
z91b3a5a7e26f9b3acad1bcc2aea7313e13940eaca2c860dcaa35a06e359550f41393271913dbdc
zfbdd544fc90335cdf9b4029335655d5b01f7d04be4e14151edc5103d551447ff4eaeabf20ff3e7
z002c2345b5a104f15df58dbee4b2e21c7d49bd53f23b80f9e7c41d9ee79ab0d4a3b9abf36682bd
z9ad10323f7ece7258849081c1f9d483ec39c3523b1dfc5f086ca0327e2fa145f96b1a3a961944d
z160874528691bd59d80680278b93dc7f7c2d16d32775495bc51580d96c599cc086f6eee48d3c92
z2744c8c7ac3c64240abab1cc9736138faaa5d539004d57833e491bc0bfc6626d037feede211d29
zc72f271c46e5a6d47a845a29e7f51c30438b1710d3782d68bf3b554280fa13f6f68dad984724d9
z4177612e85aff57ebdb3230730bf75a501183feeba52f212e6baf2f3b2b3ce5954cba126f0dfa5
z52627edb2d55f7cc383c39e1dd9860abf120c31d6e42d6cd98ee7b71b73d8475867b01980e8bfe
z0bd467d6b67d2f6a8d2c47957a24ae8019fd5a98fbd18268750bc781da2108b3c578207ae2d15c
zb3855781ab390b5d5e8a41bbd55a027a1f33c2fe48d375edd0aee2e51fdc79ee70f8fdff4771a6
zb8225ffe6a878b1508713cbd60dff13512bf93b244816038682ae81fba2e233f989e91611f06c4
z3c9ad3cfc6a29b38856ba33176da15822e9e3990443afd43fbf0c1cef8f0540fa8746304de242e
z657e2eabe1c7bd4b974b4ea121b74d8096ad06c33d4127448e37bed0aa77f66ce8d7d103f1182a
z6b85c8dcaef21b036c3f922113a3c2da7095b47286d820ad90c208203e1cab1895093c097b7b64
z987807c27c36fa4e05f34cd1aeb096952d063eabe5870625541c7d66c6d7218054e551c9fbcdc5
z29f59bc320f6c85b94ae30fd1a1c844ddb28e40b71f719e8b73eaf1f515dce9f0d48f5ec1ce4ef
zd2a5f4124fc6538055cbc5c22a58f9f5718aeaa79dda25ef2bf51e575f5e1ea277b5df703b12ea
z41b239783d4c3e436f1e49850a1bf70756cedefa8d0213dc783ef92834fa37bfd4de2c01cdf090
z0a69417046612b3a70725e66530d1b9b7df3940e0ddb88fcdc427312930b4e0c4e470e16f5b232
zd8ab69b777b70a5653cfc13a7b79b5ed591a59b5543b7bca42ff2737aaec6c2d193413929ac82c
z95c7f671d59d47f218ad722f9de77a14813779d9c42aa119b6b2d28b6ac5b3b418ffadf0672632
z939bf34b11250dec32d2f30aaac5cd2de97f5e7a5e51094dd14dea5ed2d0d4922b85c538c44cb3
z0002027dea63a1a413abe9d076044b74365d4fda99947cfc3e9e890938d799896e2a59ed730113
zc2f41801a60baa131086940161eb51e1e6f6068842fd29eafcead0f029b85d1b514eb18dc8f7c8
z2ac59f67607ff22ae20299efdf07f4a947197b58ec94c4c5fa005162c1d9d426e242b73881f930
z4dcd64923f375867b70b083806e8a712e492119e901c250bd9045b727ab94ef2ebadc05decd212
z118b983bcb700cb4d17f54c3345411d4791acd538e9c1d385c8ef9be070cac2d8d363d8a674556
z0b869afcc4192d323a97bb5f417a3eba8b36cbdfd0bd19d0e097d70109912bdcc3509c825fc0ab
z07143f00ca3173e1bb534837363de6b3f9dd5e54de39550bef6b364e7c3901b21a90b9b81f3a25
zfe931cfcc22c3f528131b05bc658e16231a07c1d97d23ff79a4f57d1f774b1b8e20c25bc519446
z6920b208a84d893b5650e883fa62b220cc6ef39a647b40eaace12a7e5a3d3de7edcbccd704b9d4
z25ae728464434c7af2e25191a47690015a21f3eb9c03bff8bd4824209f374c4f67f45dc44f83b5
z65709c900a3c986b0038766f4290b04585ec65b2d3e80d5188ba5d105720a2b99445326fb615fb
zd2fac5741ab07ca16ca6cb158c5f332f02c8a9561622aeaa3545f2bebcc476066648fbd6ac3cc1
z43cf1d4e930e380f259e939f7f9a92c12ae2e35531ad8d2356101fe70bc931df576e195bb9720b
zba84269437dbfa39e13e7b7b3b105c691f3011bd8abdc6f016ec3e1845413ea6764fcbd81d45c2
zb0e172c446fcb0dc45fb83ae2d7a982bdc86155aadeedb622731ee27e23740e248c2e2e8ef8e09
z58919359e80b3f820ebb496a208efec3a52c1203fada9697b10b41497350923a367dcc1858c917
z08d8b4551e17751e30a8f9c1b091f8987b5ee3a5d74617ba90d1810f6c4c5a24351bdecc00b613
zd9694026af8518309193bf5024cc7472065e32668f08911a29f06a664b34ba62c43c32636903eb
z046ef613c99147be6d5a67e40c1f4b09b56485afaaf674d773027b50c52fb332629c3a114523c1
z4554af1f3a5ba2bfaeaaae0866d5dc27229ddff9db83c80beeebd58800504488141bf4f5cd0b6b
z64bbcfeacd438383b2a2025dfb216c023eed32757beef4c5c4d459f7222607158c53032d254659
z0415315b63481bca5169cda9f8fdc013b1ffe2cf813353480bb0c22e6fb6c4deba9a51d290b68b
zf8ee991b83858a4d7aecf0e5310710166cb440cc12b4d8e773ab74531ec7885be989ad46375b04
zeeb5d0bf5f281375d5388e3c0b0ed3d0fd7be102f6091a63ba90acd53590e3765a249ba3a84a31
z4e70406791bf1ef8479bcfa192a1cde5c7450b07814a24a76ce6ebd756e9a60416fcfd68526224
zb56e59ca94967d8007550c6aeb07fed204e465452c9044dbedd1816429897c0c8f20644dbad22e
z6b33bbf1247effef20277cdf69ddb89fa7c028db5acda81e7eb0e4912a085ca8135a06b5926883
z67f4f62d4e0269f0928b272fccb1198dccf6b2789b2983d7102e7348551f627c5c2f27ed521600
z2cb9eb5cecddf3700fb54be1338ffac997e723354857aa3d94ab7366645ab7d650de29feade5be
z8fb73d7d8a18ecf3946b7d3ef8fe9beb353651741928f36958039ea7cd6f3fb66005328886fca0
z97c671c4da69e3b88cfbbf661a4b6cc21e3d5edb5038473f111b0d452573f87fc17a0d9359b0c3
z91dc675935cf3a0913ccd2ea7a157b6029e51c167dd9f7baf353813d876e9d3f4226f4929da139
z87421405e0e35dfdcda849f503a5a4bd41726ca297e46433bb73e2f913c3c8eced42a4a8e697e9
za1cd98031a654538f819e8818bca333e0b3572bfe1d11fccf65f0e9051bb80e2df0f17ff90f7dd
zd34d5fa1bd843106578a62e51efceb7308fecc5e6cb75b853c2377e40f11450ab20fe409e9a43f
z0d8964392b92280ef25591a9d1d12c0eb5cba910c59abbcd509f67d6d2c5ce36c003a614078954
z662ced4a2bed861f827c503772d9fdecc2ad2844be80d8a065c67f22dd913fc12160258800f0b4
z8040a7122f1378f59353a0038baffb0aedd99c444c8ef9b362762c64d3d14269d6b66c44152443
zcdb177fe73778f70a0093ac788b844dfa8d329180d034cf180761410ddc6bb650b978224ff153e
za3152549b0c5d07ec22d3ed046593f343faebd38aabde1f7470646d68b19387d2d59a7edc67ab1
z6911ca101d8910200729cf01b71ae2d6d8f1683c34d5755de15328c7db3f36abeff0483218c3d2
z074af364afd55e3139c7a1ae123e0864aa7a1f3aa50a92718e1f357b8e67d607ee813d03b02c48
z73fb7afa508ce0831f7c80f9527b54367d4185c0cc6c0e1daba37becdb840cf569662a3e986316
z14667b098e00c64a1d9d3bacb71a2e30ac0f00232b0449e06468f5a64d7a5d7f820001037a521f
zb82e001bb52d56b01ffbe0d6bbbdc7f4a15e3abc1c312c8011c6b61a17e4459a643d5b2a66d866
zbc99c1cfa980174d76e6f9030fcd7c38563ebff4f8d336f587cc7d7351ae4e6810953ddcd76193
zef2d5f7ee4f5ca14e93e1ff3a4fcf5e3de0504248537a922ea3a9a8450bac379b7adeaf5fd33ed
z13069bc2013baaa3f1266ccc73e7060a3e8127fac8b6e576e2c2a3e29aef63a184daff5d869d7d
z4ebcf800b4495943a3ac63943d340bd47c94c66fb7e64629f29417f8f9f387dd7fb7346d7ed944
zda20299acc13e0e73f477f76b2dd470bcbe10a5e0ead525645ee5e782ebadd0599c59e007b0367
z653c73b5d8d414d28a464bfd43378ca3ae43b188caf0e2e81397d539094e10ad9faa7b89f219ed
z09639201c2b34eb1515013156a30ae4261ba707d75a4269632bd7bf4f0ef2efe853a2cdf6f2323
zc57a61659a8ce1784d567f01df939e5a2099d8416889351141f4f4105dd8e37056c616edc3f1fe
z3d0e5bfe0a269affb048d2ee59ce631a127f4fbad95070314ced87f4c4408de8a8e2493a1dee03
z6837913b64463b955476ef45b0bbf20d67fe1d283d13840cc80074f055c5ed462df350a95558d1
za40d1a4fad1a13016cf6eeb7a963e80658abd7af147bcd58b04c4dba887f712335a355d574b041
z1dc58a33573a81787ba93c6034faf5a56750befe49b206677e37ebffe1713712304316be433515
zd3e22dd96f3b5d511ba7c42ffd43eb1fdaa9a3e8a8a1264c94ae75db4f087aed4e990fa807d282
za5e603a28566149ea9d49fb06487d47c8d3c5a927932d06f45fcba167774fab7d16a5bc905dc51
zdeeafa0ca159c8d493199ac20a06ec5e9a5d36cac07bcf23e3e1beee81f085b5eb7bb8f2a634de
zde97dbff0fd1be3fa802afe30ab020f41fd1c56b413bdecccb9231c35e85121f76c8f676150724
z7a6e11ee8e510e12500e74eea51c40790dd82570793813f881f45dcb6d8b73699c02eb96943ade
z35cd674b24912d4c31158c4d06c835e8d808ffacf5adab8d39da1d43720ca2c3360f3e6c6084dd
zc256fea6e98ba309d08d24e0c0bf86adeaf16952984814c8b38e2cf9aa1fcecdd7dc7b69869773
z7901c9bbd1e2bc6c353877bd3d155c8799cbd6fbab0ad2f69bb65ca1176bc13a4f9e71607628a4
za2c5e8c75eb1d344e3373a8708d1057584598ce90d5919560f3705ba23a8fe7d194b027389d055
zf9ca4eb6abf442e52096ad7a240d1aa05b266d78ca32f8ef0a21c31049e61157b9576e3d7f14c6
z264c5bb85d979193a9200593e07af3199d085d8a26dfa3dcc7fdd8a54f05a811a3e7914e2a8615
z6962d7e852972c92ac0565d188c3a756b0e3d42bed58d1f3cbf58d26d05576b6330cb5176457a9
z8fc8b61a225af1c89b5590b713dd464740954051190e3f1d45c5b5fca555b11ab0c36eb88587ad
zed58039d37b1d4305ff9e153b4cc454416c77a112e1cf2812b2ab7aafd397229596e8daf371f1c
z8de876c1beb0eba650ea57ca541497bb98bbdfa93851f1456627c19affeff5a0ecf0d08f8f123a
z915bb1b437c59b4f616f094de339e1982ab5c7d0dab6af78d9de625e9496db9622421fcdb3faae
z255055488ae43d5578f645cb646034c5aafc78d1a9739eff90f3e72b71d0fa361f40dc2800a6c1
za64ee7b51a9a22a25537f2b2b6b33000d60b7447725901f1914a04c910267f8310dab7d43a6ac8
zfed8d1ffd3546d342ae0cbaf09b5d58cbc3ad9e994183d5638c7bdcadfcc90cb6a1d69f47df5d7
z2bba0c550f885ce647e38af1d9839eb1dc0eb93a1e7d94c1656ddb257019d3905b256a5f449d04
z12b09820842edff1e2d67922217c3a9eca3663344183c673b3f2ceed8aa4c13f119970d5d55e38
z901a1ba88e8ef979286058fa1dd64a0917d9a21c0498ccbecda56dacd255c94f03df446f2f4520
z670139015951624d218ebd06b57e8e80e334bd6980ebb829cd0e70c638dad74129b3e5e98e7196
z964fd977427a2149746bec32d6db7f433adee1ccaf5a7c4ea7b01a9bbdaead9a0b6e9139fc3d5d
ze321c6e890ad1d6fcff4f0f52a8300eb29addeaa0dc9ef58ca36232ff1bbaa51027961ba283731
zf3acd401c46fa5e252c85d641d436e59b05aff95db2c3024fe9c043b6c006e105f3952b4bb4237
zf413610cc9a072b6218c1b14a9ee57c5712f54de8bf6c6efa8fc6deb1aa39dbb164908ce52e18e
zec6b320205c36c9106ecbd0c80534561a7bb69c61cf660f577c10ddb08523680d4e550fb9c4f38
zcc3e6b91cfe9f058796ecaea0306d4a492906e1a82c988b6eb802c581a64802d4ad4db42c3e417
zf2df5e34a6cbee710d0ca305cce7695745f5d85a9d7fc9d15573ff49457771230059e8d00df717
zbafa9f4931332d1a053943a25d7781f66e3f68c4e03efcc27a8052339c2cfc6342308a48985196
zcb2c331c8b910e77f9c03b44e3130b46fc957a5d8abedfeb16583540d8f6b63c447d9ef8ee645a
z623e5cc7659d01aff4ca62bd6e25a4d20c260982a70eb303be2fb2942ed079b0aa970d28f37edd
z78508220747919d4003cfddc7dd3e17ac4af70c75baac2290ec524226a4689c3282acb7b15f070
z89d8f583847e7506a1bb19c2e5cca094dd9bf1c8acdedb4b65a155d4da438b1f5816eab7f98ad1
z83fc040c9a982e9e34f84d81ae29696b57027b4cdd88c010b82f1fdc67450f07c300409c9d6f6e
zd8f7c3cd903e4b6aee47929d0583ba5f26ce49826c579b919f7f2d4f399f9710b4519589b7212c
z39983369c95876610495b1176bfaac43867bcfff709ae1b81dfafdfd2e976c5c23b2951c7ffd3d
z6db12f70ce8bf11ad73600e95ebd5b40911cd6e94c7de431ff194b62e134497fae138ccd093c2d
z842b66611b4adbca5fd19b988d0a5b3e567c82d8e9457e25bdd0d799edd0ebce6a5fb8f54a0a46
zb5b0068667459a49f5f0a41c877ab67f87a4aa47014030d31bb9c9e2a01100413b0ee912fb869a
zee8a1b76cd0357cb4570abd517c5109149ac562e93d1c385d2e6301fe8fc7ace84d8e9cb7100ca
z1403ff34ff2b662a296907fbb59a17fb35a9ec8ce16395142818b00d0e3ba0ff93c5717e90bc6a
zc5efcede3130c1a026ad0a2d766a34b6890e30fdb56f91d0ce27f9d05383e53535b3c15903c890
z20a9da17e433673363e0dbed9c92b4d87dec81cbbe4edc2d1026144e7393399c5e4bcadd9aba4a
z4d1c55cc4dd1623e374e483266a5c43234e5cae3d01ea00ecb6e8822256a7bcf3d8bc0f0ceb240
zddd32c5459aa7e62a15b27f6dd9bd957752836fe690bd82992403f931d7613eddac5177fd868c6
z5308f53d776db1eac6a9c69219f46e54ef27f313a8f3eaad384f657cf5d54da3935f097ac2deec
zb675d22c287cac16d0ed0d234043d5cfaa8acee14c17659b51deca763c47b936dd70b623546c17
z3d8036d3855163ba3bf06e36e2cbf88cf330445c8141785c67ac8ca1bd93ed2cf59621b95e2fa2
zba6a224d1ce4132a407a2a3c010539b16cf111935677a00d7c030ccd99638440a9cf429e493769
zcf00e4c90b87b5064a778a08ba7b6aba181765f9fa4c16f769ecaf164bdbec9847d1cbf901d80f
zec4c30b766330d353e979237047bc628814d01668ba319d8fc421256130c1dbf0c0c1b74afd221
zf1ad283e994634670d72a14efa999acb5231d79a7fd118ccfa940066ced50a2fe0c298ebdf6e98
zaa8374dc93dfed27216cd3b2237f3f18e7c6aa84247e53c72585eef722844f9cd31f32054764f9
z63a255d70638d0af05d0505cb7c737a05ebec86ef9325e7f1b883d3560b03ee1c1364da15d6b0e
z98f82741622029cb27f96f4780831fa34eaa352ca0d7091a120584a6b8f8ce51879a10bfb445d8
zb57fcc41f8d9daab83e2d7c4673fac35b117ef43744a8f8bf5fed1b5d8faa29a7aaf143e7df11e
z40d58e92f60fead0c51badd904ba52348c2510fced180be347e847fb9ad010bb46f47e28d58f09
z07f0cfb898cfef64785a6d5ce5c06efc00e08bd9e7bd217aff361df1750da8f52c25569ae7469d
za04f6ddb3f713019d97b54b7b9aa03b5813d1c92b8ca36b039df2b1fbd393b9f0febfea17adf40
z09ec6f2c4f68a6615630d75c01b71314b206e8a5fcbdac8957efa5bc54cd2e1434946cd40f669c
zf0a87696844c7e728d190ba74cf797654b058722d3aa2a17a1ba344672e499ced68cb94d246ab0
z5435c99d24e4a4c9670254580eafdba2122c53ba27e382aaf918113caa0edb27e1cdcb7e4174b0
z9cd937cf5f6d7f32c4bf3685a2f24dc6a41982c03b97697a9d780c20ba47a69a503754b91c4b11
zc7ae2529f59034d74a572ff12afd38dbe1928545a37298bdc12ccefdfde16686f084324da96657
z2ba38a659966b71a09bf9e2beae330298abb0e331407d051cd167fbc7be5e593754100a5ef08e1
zcdc11f8ec0fff3f0a9f30df4f8cb694774cf72d3a65f7e0a18b7edf4d3ccf8d74ac575c343a3ab
z59c98eba47a7dec7d40fb328929096f77581e2ded02921df62869fb0738c0ec30a1e7ca3cc93a5
z2c9ed7934136011e28dbcc10359983e879992f741dc8edd7f19f5e8f37c282e255e03b07aa2098
zd40dd1d9c17df6965e19cd7126181283032434c4db5f44b015514b440432b6d313f4be1bfbe9c5
z26edab25e466521e031a68d886cab247bd31ab08d665d5b54f3aadbe17ae42b71ec05d38db1091
za9a6f85abf25e5a5c7f6bd02958e8f66f2290d3acbe81babb7f98817f099aaf18743b1f91e82eb
z66706f4da85dcf416e01241d5f5d5bae90d7d67fb1710e64ef8897e07b6568e018c554edc3e581
zf0f71ff778c58de303d3f69c3feb3d763d7371c9774d4409c6b1812e6c23ed78334b7b718bff89
zd7cd1a4b966244f8f74db431c0b9a79bf75aea3d70998d1db59bab34fb40976d4684f61345243c
zfce32dc9c80363762fecb8d862f849a695de566ea35574a33965aa1cf8cafd7395fdceff27fad9
z9bbc3b277bbf6adcc8b2608ba6d03008a868f960f8149e05e01e62e3a6207907d2bf134d060fc8
z3d51296a1a45ac849eb07348631b795c4605420311494742671e1d6f71161262dc857fe51c7280
z32d9806dc7485ce221f5d69ce146d43ab68cd321be97290554f7fa3ed32262cd016c99e5801db5
z9fae0e29ab7bd0610294ded689952adfdc80902dfd0cdc0786210bac7f4020cb040ea79969f253
z02bf2573be94259241463b96a9ff57b41c46a9f41fdd7abf9ad11effba46a05f89fe3cd0af1470
z130e2fd0f6446f6cb1c32e9c79c48b7cd586a83756b7dea7a3524edd844815543b7cb47de12c5c
z8f60567dee49b95ed62787b6ac13edafbe601ac80935a9ce2cd25cd80395433d841bf597431730
za06c87dce8840f9e97755f38069ee932d0806af93948bf085044d125b4e04b3f9b9bd6512f0ef6
ze2d2d78fb343a2bc02503ba30093e5b24943815448c7b026d5c3a5af9a8dada3e0419528516e14
z9527821819db4e8bbc0a65a6848453da751220adfc03e4ecd480dafdad07a10cc7ed13f2ab8e7a
z4160a94bf2aff6026cedeaeb3f389741396e46abbc945f88098e6091f027865fd5145776d8118e
z66e6e5b635e3ba49a76fb028caffe1796eeaf0d50ab1a7951a106be509a9653971c5abcd66d81b
z350c6f82ed0aef66c8603dbd1f8632ca7a3c87b25860c79ddd17510efbf62d90dce83380343eef
z00885d388b998d32608e5d25d1cc08882a964c95e68df778d29a274ed39a33035267da575c17b4
z5233f72c84febf8db11b6955ec5c209ddfab8059859b6c2e2cb773180ea2cf1e34be85fb24af74
z1d1fb5d7250f6d801a99634b8e2aeefb810ffc966cdf9b9895ae4657d602e83032e1f15dfd833d
zd40ca9c83404946767472110288f79e6a9861afa0d0a477a3d563d87d9999fe73088533c3b4d99
z974130fcb020817d7eff4ebd40ac335d387496c6bba7222c5f8f8a163d4538f675ad871ec9b2c1
z358d975c5c2e9093e92ea742814c550ffd8cd332012b4fd739ce2bffdabb782094f205480da9f9
zaf9c810e134d930a7dffecbe351da7d7fb21d25f908a1862e4f9ccf3856ac4b6932e8aa723271d
za73b1e83ed1758e1e7ff570bb66395e24d4943905285babd65a7a472579e3f84cafbca99293dc9
za1978a84c83b3d608bfbf086983ceed27d233937476746cee50a2eccd135c86692802fe3355302
z5b918abde27390a8204c84ef24339bb4d8b6b90a874932cfefc12cc457bc76047f238b827b41f4
z0cd15da87b280b8afeb8d1fff62036647a35b87ec864a2e4701f4d47647c83928a3e2d72a43220
zc79aedf7522404a17a70016293911cca07201f7194c22fec04a11c3f38b54f123f04c44d5c4075
z6429d994c2a3a3a03dca0437c3d3cd9a8f6bd0282c36c05cbe3e246d32a54af22f9ac1d9797ca2
z8592db8a3e2aabf35814b42b791c0294d1231419f712d1bd6399c43bc579f4eb5933e5aa330066
z056f088fbc0f86e7e637c3c0d7e06aa2f895b14d3a9728daa30843381650cf4360c948097b8675
z52f2c3481f50157397cbcd783ce748a41d5beeae950efadfe615a1b65e6b69dbad593ffb811538
z98faf0f21c166e578469a86553905ddf89ebcf26c78c84728b7819c8ec7c1905060f9ab975a693
z01172b2ac89bde082093a8e8ab0da2cbbe1ff6214fa2921c1f5af862c7c66335df50c03c5006c7
zaa6003140db2d419edf9f877566aa0ab12e674e3c7dcc6189b885ce97be73af92cd08f4a5c487e
z2233e3a758c7300992503c29455ae49a9eadd3e2573e3e41f12037811c04cb575f4d1fb4a1f91d
z6dbdd44c202aeaab2d7a66253bc220aea517f208ddfc9a3e37f1f92dec7aafeed3f998722b2f7e
z0d5c52042738b0449db53ac4339017ae43832b627317ff4dcdd71c13fa0270c41016d3bafaf1ff
zc8eeb0bc9983b6f475127ae1ffdf6be892d1f964015a4cc9478094b7c35338f5940825443a2477
zf8547105e90fa80d8231b763d7208fe43aca1d8c538c36ef43cb25dc6eb809f76564e0432c5474
zd6521516d00f26bf033e0c2796f26268abacb3310768262c9bd9af2d05aedc5e93cb11745e115f
zc91985e6b1a0874025c76383c7167d1c221bbab1950bec34d03f1bae3951c4032029d15b888df1
zce6371c9e135c893a58411bbd89cddeb7661c2fb75a1b4da91d141c9d8e1e2c93eb414f2fcf9e0
z21ad1a171639a6de2b118f858ef86dca553522bb63a7556f0414eaa3057d58881b84fe23c004ff
zdbd44efcb50707307e4fd5336b5748e55aadc178b68035c6cef0d02cec513d9606d3df0a7d246d
zca4559bb08d60f508fb7a27480294511599f569be79a7700458aa6223c3ba8e941850b0e1aec15
z77a2b630e66ddaa824c4b54a3d61bf4eba8d6772cef08b93d6e19ac8c36271d7fb20f4d81af34a
z01f7fec3bbc17058640486a0eac7261192a13c61ec853ae4f19873baa99afb1114282f24c521fe
z262223448b55f13339b549204a7ebe4f1943e83c85728bea295ece1b0c95f0c998018b9316d2b8
z49b70d650f5f593dd86e3dfa8952bc9673cfefd70a5795f386a9d0e986515681d5add803e84f5d
z77123e25bf75728736a89ae8e6a4f25b010074f85a6f795ece35b68ee985888c06e7d8277c6ef9
z97ff0ea0977a7c5191f1c01500a9be512e51d7930d61c45f0e69e5d2d8821b91a3ff1468854475
z7fca0b9239a4b88001407fadceb3e69d85b705d245aed7e5524b4d7669fffe7003b2b797663be4
ze6a88f6e1f8ee031c599acfcabdce22263f96892fc47dd34640e1124e58e4d4a3f86f9bc4f3ad0
zf07be9292c0700c256ec7f208ff851a7568c47c3c7e2854dd3f0768003bdaebd9b2e7b084955c5
zea1e0f8fe318bb52c72455a5883412bf5b6af01de364f85df98d0e4de55f39947caa25fe656187
z8ebb73f09e79ca8c1c22ef4b9f698ce38b424ad8f0090f68754e86f4caa41610ef36d9744232cc
z02af6af8216f0b1f4b4a36c9f3d053cf3469b71c04b0cc5f180e711b373c680e784d90354c6bb1
ze0bd257cb22d95f41a3acdfa7a76aa86f4d157c1af65994cc468f36349ec15034571378558058a
ze7719e81f7939b9db6e1d896f2cf7edf6d1112070c4c1e0bb828b18f293e613e69eca37ec452c5
z5ea9ee36e327e64bea15ccbd17946e4249ed25fd8a7b2bb6cb98b3a6d7878661bbb96bc6492e90
zb74ea12e8df845d383c9c2e19e503f4559bef28aa087f3fd157e1404a5e3c86cb8f995de7e3754
zbe55d550c4dc94a1d485d04cb552bee5ae02533fddde39e6c456e206f297a198fa470ec186c5fc
z1d624bdbba0802bba3bdf507e2de61d38e13c16b287339f8a5fc91717646eafab4ce1feb85d006
z5527d42d4be71beec296ce42b3fd91f6bb6f31e8983ac45ee1a7a519b8e5d69421bf65038514cd
zac9fba9787559f64ce7ddb8477c345febc6b1f8817e97ec0094a5cf85eb787ce52c4231ee945c5
z7e88d3bb2a79224f2487a59f59d39c5f91e4063a4192aaf520bc72bdcc00cf5106ad4c2dc30c10
zfb85b17697a8b0f3ed6f2f2280117f14805ab021d3ce643e4e9c424c65c580084dee7877a20b75
za6ba2382c25b3556538b1364b0179ee23acec4ba31ce0210ee563b867899b5326007e747a0bfc7
z18f0a78a962c7d42e701890ae9c30740870680051727a27d1991b077b0921f1f89535b1cd07d50
ze3f5969a664c8a13172da4a77485ff13d8f6ec8d4110a5673c9f65ac091244eb49fe5eebcfa8fd
z9741098cf50c27df0f7b9e1bdc6ebabcee975f9dfaa9eb7526e8df4c98fcbc437efc157655cbe5
z3c8349df8c296b0a587a8cf166099d124384c594cc8959c2008168e49c8f6dad90777b585d26b3
z6d1719fe9955a8ccf88ae5cc3eea6a414257d1d01ace7ab7448592ea7e9c6561df9f2be2b79309
z8bfc8cad69432ef589c3a2e8a9de0b79f2dc494169277a83c2ac0a038ad535cd81b4b882088d33
z1e8ffdf562d5557823f96b35dbb0d61d1dcb6931c49acfacb2020f8341288288c45e9cd6b18219
z0de879f7fdc2856b7e9de267209511bf1bd8b3c2d72e5867aea3358c25c0b6764c0474e47193c5
zfde5966954c007fe1bd1e6336aebd49342da993dcc56b01c43179c59f7709b72f05a6c56ef308f
z4085d5e2305b3e69dac033b782897476e8fa731ba24578398e729cec0851f8bcd80d5187b923f9
z309e64e80b63672ff60d5c86187087a1e136d0565a66eb4fda1a174aad32f01bb629101837d18d
z67cac3fe2724b827f48dad7c50ecdbc4b1ff735d5a24ffff5aac047c2ba437ee453090ef753a24
z1b96701f0027b12499bdffb4c74a373967c5146cb1444a16df6568713bbabf703bd841c8f77990
zbf9156500c19581feeebeacf811b3bd5f2371f675a6c27fb3e8303a796cf873dc83c596396ce37
z6b378e6630890d350616dffb504bae18b7aa8bb33accfaa13597aa0c0ada321c0b146cd1da23d9
zcf46ac7f73d0365db506c87b8c41733c660c76f50cd908413acc3787c417c59213ca8fad330e1f
z3c623f3a8019dc03d03c2039acab0c66c18396c32cb6d2ec7fa1c0bbd6648ad768d98ac5e6898f
z25f792472ac275777f553add7a9aa291d8828a9e4168e8bd0287ce1ee074deaac37ebb02ec8859
zaaa07bc0dd4b88662f550554058afa9a1015dd320f23da0821d96c52569f550414cfd8ef7e1f9e
zbe1172f32dcd9ce5afaf88828176d319801f78775d438986048f2d66b765272fc535f60f40c921
z9aeda53fd19ef93e61558510dcd7f6949bb8da2cc1bc67f06b8d4d97dc56006d22e95e80363be2
z36da32a25184665ff5da22dad4aead7cc2b10a9bfac899cc9e0b0f88426c432fcc54bcf19d9814
z5c511612a5e11adaffed997b6d0fc04867702db409bd08dccf64f89d527ccc97d2649940687f2f
z70ac7a16b6d85c8c358935aff787cdcce6ca74aae9662fa3c83a578457208e42df4f4af7542c74
z34ef7f6e11ac06de639964c970f19167f79ef412ea39fbe535e47f15353d02f22be7759c553a61
z067c221ba72561d6af842cbf5911eea8be0c9fb5bef6b2b6c64651939db8a9658eaf15416e35bd
zfb0485b7f6fe07da6cb1a857861ab80a1a621641b25ca49aecdce964c3e2ad9df13618c47ff43f
z16037a3ddac116143c623ebf7bb10a921c234215c105467e389c9bc2f990f4cd6c70ef0a47bb0d
zba6665f819a794f9a96051c105a571d252a41d56533037ea88671e24aba676835bbdedea15f448
z607af1345d9f8ee72c03e5aea8cd1a4955f856819fb475cab7beff5db7af8d7f498d80042e52af
z95d7ffe4ae02a46f0b038899e46dbeb87b629ec9c12c3a0a9804f1bef728580a8b36d55baad2b9
zbfb83e32544f5393862e72da7438dd5f31d9214b63befb61862456023f89245a8011bab62872fa
z81672faa6d9466bc0829ad1ef98c42951ba8571482731420a330379b0caeaaff9017e3d30791a5
z4d9f1b80b026971eba044387ac1be27ecd6df9f83b9f1ce19ccdffe37ad1b956925a9ea8c786ce
z8ec3cb367c5c12064fefe6521e9950971a985de7bf89ea523c8925a54a01a01b56b6a36e84c2c8
z356167575993c7114dd3e4b32ca47e2f5be40b9a4aadec0ccddbc47f59db46412e1b69d9bba9bf
z5dba5a155d60b5f031f2bf2e025d1ad528f7dcdb8e047e76514a0be2ce8f0f61c3d65943ba9899
z05fda6e27e7d80a5bd9f99695bbf5093ce79f9152088247e477b124639647ca654069f2bfad357
za04c5f10eec4b2e5f1cbf42f7de60ec2d90bf934530af0c7d1639c53e82d34ccf1034cd217e4dd
zdea6f7ddf75657f17f4b91296abf0e282352d36aa74aac768741d2932bb9b6dbba730a95486576
z782095b14fc179c074ea082b5a3a2229c3290a14bc9bc487dbfcbe4c9ebc59126a3668efd0c9d1
ze39bf7ae0530ac3edd4554daeffaff81d3752af4a41227b832b314908ac0b55bca77cd9c8bb06c
z3b3a716b751071e1739dd670ff7cc5477b117b65bccf04ccfb476ffc5da18b12bdab26c4cc0715
zb9a3b3511829713933e259bef529c451f6b285e1e9cb5a84591020a3f25e16b8f4411f55e196c3
z0c854aef640ff590698fdeda18e3594cff2b51a4b3b96b3b5963aca927270d802594d07353d874
z3b7881d9138497b7102073dd4ad03ee69a8aaa7c0d9e6f2080e522c4cc85d412da4d67bec73022
z839bd1fff90df9887091c2fb9a308fb833da6d85d4ad926baff86d3ef182c9c4ef40beed8dcead
z128b64c136bb5282cf231f2ad0292bcfa415e8395c85064f011456055866fa961bf56b78219d30
z0d478933e79691ba0ed5400fac6990363b637f568af4b03115218eda9a0ee629d50a130c932361
z0c90547a91fce84072add45ffb9d690616bbdc8134a4919779c7a019708a8128a4b4169ded630d
z97f4b70546f334ea2e44ab2926b9740b0fe7261b4d5c5258877f2df936abfb9e917e8e8cd30a56
z632b9b155402bb1855325b306ea19e99c14f2d8cd34167a04d958520ca6f67c9da2cbb134a204b
z241643ddc2886eb8f530ecce2943486f845f0ebac98c9720586a4d924935e4cc4d65645edeb318
z446b6da4fdb118c02e0d117d9c5ac2a1f5f80185694933a5ea98a06afe97d9ce7924f9d45e196a
za9da9f5890251d27e423dd329a86afa6cf3a4cdc8671c9f27dbf3abee77bb595be53f356151d8f
z8fd73d9a816b11a24a7fa31f97f9d201449f1c0b2b3586896059d549c2b79aa312eec564060cff
z4c8f0fcf59c02af657b2cab74914366845ff849f864936ab1ee9be11807b472fdb3f36bb31272b
zaad9995cdbfb86da6b27e0673830884d996fb0a0e3f326047d5ca6b6b5840c182b88d67d57a4a6
zd5cdd9d28c8e987d522ed9cda17085c832b5f664d2a8e1a506419be077daaadad970aa8ccfcd7a
zba40a0c8f5a7554aca1fcf0dc303bf8f71532ac872273db17b2b78ef05dccfd22ea023494f49e4
z3035bb2781215c54a7a2bdc39d4862779bf428980e96dc7e1384f8ea781f8973934bfd46106b79
zf288a1e20e8a6432cba12ed69fcee7a32420b6063498284e21b51559c4682e31e5dfe92b5f9dcb
za8fad984a2881f1dafb2cd7a704034b6989ed33285206e4fab0b2b9f502fd38e73bdc6e0d33994
z91a80dd93ef077ed8f60e1a3a35ff6a2472dd6270a537e0887c3f8a98070d8255ab0b883fa7be9
zc992c0106161ac3ed50325f1f5029ddecc39b1d31e2fe0b925c79a971d7e06c575a4ecd8d24ba7
z2037f8736b875ee62411b388e9e19a8912843db8de883b5f0b5382387b5309cb924c8457451458
z85fa261aed2d03e9415adf9b9a22a5f43cdb633992307bbf920e39be83c9a2825d722f239d568f
z54912d4e85ef98f59d4ee2308fe9bca1b62858aaa791a3f5697fa3173e252cc1642febdd7e034c
zd444b30c0d674bd094bc3939a80540b879bba850bc69b278165390e8d1105fd25ed7cd695aa4bf
z92a39e64716b72a857e6ccf55c26f9ab422fed79b05ca39a211315789dd73d55b028cb3891dcd0
zd04566add92fdff201c01af9118b32f3ba8349e3df9c8a134f04c8d53a904a402139c1da46347a
za6f75632862c2f4136b98da0b9f095d20f83238d8b6f89989ab6fdbeb6d6dbfd7d54272fd86385
zc3a3c444aa8e2de8d505284aeeb303931e6acae34c9c09476727d16efb4b6ca277695f9438912c
z0abfe37503d7cc5cefb2ef72f5c4315d1fe91dbc5b64d3cb68156972881860816aa0e72f2400c2
z43848d9fc5248365a87ff506337dc5042e39a9a63709368d04793343a4538721684613ac03770d
z6168ab4d2c01d51676185599d92fc0231046f070f7298cf2b620fe7d82ffc2a6cb897663f2ea74
zc725cad40b09166b0e5ab55ad3d6920aa29f2ecf66dba863100d82d2808558e9ac679ea42e4136
z4ab1af07110f4d3f7fa2d8bfaf7e4a1fb4c3df4f29933012dcda0a898b57ecbc1edbdb6bd917c7
z276000205e059a298e1af64564b243faa869819a6889b429c88d21eab662aeaf9fde41dc153371
z0a9def48a15ff155bac34157160e21df8d0b3f1602632d71545b4223f04f4be1345b931346de54
z75d603fd9e727ef06e4c0572799c61478a7590152583dd7b677e040fe3006822e7748c9eab0d1e
zf63a01c2467b5a2f666568d99921716aca6444b5cc0dafa44e068becefc441dfb33f3ec3732565
zda512b6b0ceb6ef37d07e47cd6d36dbcf7e4211ef55fcc38c2e2dcd0ab480efcc2b9d82c34b306
z740c837e334ef696f3295fed55cec96115516b6806a63814c7d9138498919a16a3f6e841bda11d
z201a95abc6a0958ff7cff1c27072b4c4e6e7dbeb324e4303a50816399f4f5fff4f116a9aecd285
z72340c40f9250b92e10371e26c29c0f1bda88b75fdb68806900dc77895e89f74255eb1aa88d8a3
z3fc0bfbe5af12003b22798af60a48479b481c6caa41a6118df5d5b71b14d62de56d0f319e52cec
zfe8cbc2f8f72d61b5a626a9d0c7e8d2ddddd275c0395c4a0797b53c6d4e346626634fd2e1a5230
z20bf3b057e58bb4b1b00e731b84beb7c5c3864d8d91424ac37b262dbd6405dd1a27d5dab026d1b
z1c4149b48fc40e6e25aa16ea49dfd70c62e143761a3d301b740c0cdb9c38a74a00988079d9131d
z90c23c0814811cf344f0b6790d9a81c86559129620b45d664b4d5b6ee8971a501b67af0f5d092f
z2a321758b723d1581617892528372c3a7c8a63233e33e17abf69063266e33621b4c0985adc5a5d
z11a1a1f550d29ede44af0798961ee9ce7552a4b0d162ce6427e9ed0faf9ce57f16ece41720e504
zca12024822be982a06c0181eba97c9861d6eb6fb5e911caccbbede8a13c42272b109e907e4464e
z408a4464de76219481f5b239b79be1ad2f170b0079f39de32209194004c238abc1d442d18b64b4
z136909c462eef57aa154234fdf681f8b9d69ad0331ac1dd38389d00a096e1c58035d9a63485900
z7a5ae3ae61f69b68d42abddc9c564e953f8450716d367a5a991781f2663bb25e3cab60140f344f
z103b5d5d5bdf56554348e7a42a3843c38010d74cd83ebbc427b06994e527c2383cb3a73547175a
z3858f97de4bd6341a7b51b114a775edbf989117a6a672d544d9ee7bfa9964ec35ced83d526b582
z277ddda3440271a75822761ddb7f3f3a97049bfb34482381233d3750d3a06178783229bf8c0a41
zc8c6eb91879b8ad7e2051d182970c4f4013f1ce49ad018710ea338dba0c4c6a20df676630563af
z5a06020965a05dd0c410cf902261bd4f8ee8182af70cd464a67ad603c87ae36a1a568fcc952b27
zf8d4074e088cbee32489f1259503142ad7f2d04e3ffdc5b661aaa49baf71db5c66415f91402756
za2e5f194f250b77c5af55284d01cf8ff0503a3110a5755a4aaf7c991d9ce6d56b9307e152c79d6
z08552f3c64694cd25e812d9c1f7c37b5ba166dbbaae260180f368b751706733747b162b21da573
zd019c25ada27f7bd98f57cee7bdee71392b46055289e977867272ed3423b4d9b5db1c3e8a891a1
zf247e408e33e56c8a9e3b15032312dc932cacf2ac92df528d1851d89642c24f2b2267f9eca1dcb
z56af79ba23636c9ea1120b86b849c321971b158b5de5fdd66f270fd9cc9b7bf007cfd3a3215398
z9cea11b2afcc5dc44821be722a7ee9d23b558ae93a597b96d50a211816342227b6b45365bad312
zee5e77929cfd4e08f68abdb65cefd3cfed5934cd563ab2d7aa8252c1d7f954c28e9c914c95d2d6
zb62c0c694518d1e798e0b9b63df60d1270e4c856e47b401b4588fbff73db104f69b4bad2db26dc
zb835734fe36690cc094d1c04f9694f4101cec974d46e0d4eac9d24c24d39c546b2582c42076970
z3d8cd1f5e446d2ce762dea43b0b1ee76c51bd919a5ad1282737d424c112d6d75e257bc4d15b5b3
z236eab38dab09b24346dcb26245917a8547074478cf2e51979745b7023c32b636afd8867185bd4
zb6077401a8a1839c7454b2ee0e80f5d47e83a42afe0a5255475f204b2898321769613eacf893d3
z6fa0dfac536cfe4fbd90dc696415e3bd3244409a89f3ddc1757ee381f6b9578ceac64708439154
zadc431dda8aec486d098304e25cfa30b1c7d9276cc2be71137cd0a6ac929a38811443cea3f5c99
z3e9a11a916506cc700bbd074e6df86d72e76fb3046bf443a1ee9db76e46690945f7bf4815635a0
zf64bc5c4b98cfcc05f675f460170ec5aa4a17b6be2b49e7bc4d8d4b21c0007fde35743a5c56bc0
z7c0c7f9d68548abe5b01cbb81711198bada2e9ffb68584b8efe9f362eee005daacf6e8211dbc3d
z0cf2886a6647cd0e0d6480e6963e811190fef80c7a4a140b6bdc1e357108264f1dc07c3ef61c21
z9135e4b2f2b45f4966e1e408f6fb36fd92c104c4f1c834dec672de2c63ecac71cc54f6e5c7827e
z3ddb1acdaeafabd2c4e116687773f8e44c055b2d604b00c42d69d1ada3cf983cfc32470d39c723
z0e68b50840afe297ae92f60e86090e69e76a53fe0099f30005b3048878af3f99828d374345d7e7
z838fd19eb2b6d811c95c95017ed16e71918477e3ce924919cb72bcc9b131f81b42c0fae6cd856e
zeb80ea370392f77249e0594c0f7281149d75b55a264c6e708aa1e994c525f3cb26ae1a9270674a
z68134d2b4ef8a7f2d18f185a5ac2757ce0ebd4004eae1ee31beadeaa0d26f570a18548e96fe5cc
zadc27c3abedf3c98f03c192e2937732a017baa083086ba53044ee557191590c17adff78f46bce4
z0d5d345b53ae7936e35f4764c6fd245e3df1c2fa041b86cca280716f03d3c458ff0f7c72fe7712
za6fe0e18c8f23d417d8ec896cb9a3e47fbf0c84c95b966b7fab5d73dcba95dacf6154006eb2ea6
z722c53c4c786b17821bba542786c7c6439b92b55fd4904df4bb298a652f5af1252453ea33bdf16
z39561f65df318cbbd2d9c838d980f520f839e2d838118a77567e1584ecaed5981084a47c119181
z271b187f4bea29add9354387491bcd316a4aa9aabd937578ed2a4aa9cb1a4bc186d8ebea9e5df3
z00cfe90ba7711b513f66b674eebce0095f1d1ba9a177c4ceb8caf7dd3545d8f4c1e8ec68b4d7ee
z2e1a2dfa7df69324a65d98bcd611be0ee900e7c45729733727a3730b4a0757ee7033430379f326
zb5a3ed22eb813eaa77e17bed8cb4cd0a086246342a75dd38918ccfa4e42b1989ce6fd91d3f4722
z21992fa224e62e7997bfb28ac107834f2c5b44903a04140081fb98b153dacc179db32b209340f9
z120c049d778a583bf73835384ca8ba4d875f33a70ad7c766463bc08ab371f96a6389f67976dec8
z7da7b6950ff2ca784ed2100740fef09bc42fa4f8d8a3c4e30b508881033b63c2eff2030ed750b2
zac2601bdcd284e21c0218975218cf5f49bdce0f6a37654bd4d29a87578a574c36cd1db54b13da5
za46ef9a2e3921a432263b44b047da460a1803e5f327d29465ab86513a4210476aa547b3948f4bb
zdfde2587a26f8ae5c6fa5aa272316fb9ae220de964fd606a19d17d4daa338114695cc549f63c3f
z23ecefdc2b54c54636d4aaa08159a2977275bb1cb4c9ce8a1dce8c94afc5c55b3367c6c5ca7984
z1d7a265e30f413aea4376de44bcc8cf0425a3db23ae906af0b9627d6cb64f2e0e7eace33dd6df8
z0a15a28c3bde1fcd99e01d13fb3ecad4e45424fea8f65eec7f99569cc066cc27d41cf97187a705
z920c35d73bcd31e3bd648caaf9e0a27b141d654e51704d26f622621b97bf68fb50df53fe86a287
zcc8056e74eb56908d4180f130847da53acc9308ad069b86a211605484cff36be50ad70682ec74a
z2c89feda439f01ef36a9ad8d7e6b964096e2eca47061b4e01f4be33f0ae1bf57dad0439273e5a3
z208ea76b50f53669830890ca3b54903dcfa43e78411d5e267cbb1dc4f1ea6f11cd5fe1a64d7419
ze7f2749a1d94143ee572f19ae796af67de1e445b0e390da1103944ea6f9bd7da6046618945a5cb
z17f6b7dc0d435120347894fa5b624d7e0af966e7e2ec2d53a2339a760ce8ad380d8a0b43997204
zfc31c2cb6f1a9454252b2c38d724ebe99e8952e72052c393c35953ad7747e8b8140360fdc39746
z4805781d305cd58cbe44a2e46e4c601cc91487b5bf2c8c319e3994557f7d83fb2d4081a2448a48
za3a3776d14c1425141662720042b5a8930253d2dca8b09b92c5af59041415e72b4173b4cdaa5eb
z5d180d4a608c021047a139a01000d6e301bfbd4b1e6c3b8afe55b2b1e506624003b4da78c42e67
z0877e4f64a0f803c0fbf0fc8634db7e75152da732ff6e1a3f229bdec1320d072bdad15ba1ec3cd
zcc490cb306564c82ff024e90972e21e73e6753e85abe47d79983e264e9173556e39c43cb0d1686
z01b58a7615c86c52e98614671ae3a2f157baa4755ce4680b25b256b77ff820834268721c1a6a7f
z6889acdcbe2b10c086e84f283492a076ad4d0e8a624ae9fb5c880fc738381babd2a6324062c68e
z1990456deeab2cd01cc62fc931e9f833657cdef54da05580650401698b0d7202da375ea9d87bec
zae0e2920cb097fa88e41c1e4f23b05b0455b8ad30c908bc0fa338b5f7566c3b3016d63369b8d3a
z20be4dfc4d84baea613619543796fe9a6b93968193a33b9e7611bc6d6cf970731ebf150efb43e7
z8f54dd7b3e55f1224760ae9fc40e42aeb15e4257f1202e3ff96ea335d49ea57a30c497d502afee
z70aab9a756d9274538062e17f565bb3716aed850c27e5c0d5847e6b950867843cf70a117b37ee2
z86b30d5194de929f7221528c44b65fa2c9e5ff410819f98e76ba9080ca5a3d1f75e16007d0c3b6
zfec5d488b4e857b7cadb4b1ed8641c410c19f6d413ad6aedb41d7a243d34860dfbfb707d6ab75b
z4bf31b69484b1b2b7629327bc5df07a959adf512c2c2c6b78d86a467e0dcd0c5a7486f8ab55652
z57eff0ad936a5c164fa772072a42f5adba8dca54a5b38a89be00373a84bbb3c2e35f8421bd457b
z2e323ff398177db9fa3bdabced43b23206647440ec5b1f8d75d2cebd8f3586f2368ef32051ff55
ze9d481da13c96a291293306738f8c0e0dabd438feb41257064592a140af0c58546b768ac660a1b
z2331fc41deab0263b69c7812c038d80ef6357b618713e12f7010fe2ffe9c7c7ba427a234d9e415
z6b24ae3ff8f38241ab86312dd33c55374e332a3de63394bcd5151bd06a4ff07290b3b179892552
z9129e02fedce4444dc8e613ef6e24214016c00aabc13e41cf91708fb650333ceb65582ae3126bf
zf4352fa680ecfef2435b5fbf3a668aa8704b592d9d9844548e299dc8798c8dc560c660baf4aa44
zad795f3e66e67330a7042f14788903ff9ca1b7a4da07f61c9e87bcb25b3bc9ae2fb3547a96ee81
zac52df7f46e6368e7560db519286e5cec9081d094bd0b3af236f7d50e56e89c1e78d7bd90f4de6
z78307a2137d3342d7ddda2b0bc89ee58c880f1b372021291a9666c9c52ee13072b1973931015e3
z96cac6f259820b986fb7e147acc39a0ca76ab3d08c1f6bb81ba685b1dfafe62a223b8c2bd611fc
z480bd38e128018c57b8a6a08dafdcbefb12aeb7f8f5b52db11ef98c8ec63f202928503194433d3
z2b00cfe48d5e60d46e01cf20138f481713a5f38228234721a42b7b951f54b9b53984d0b849cf73
zd63324661f432d4c5e665ccbcaf21d64f31324d00eb9d5220aedd57f77cca82bed84cb7bddb676
zb3646b130d3ff7cafd601b3f18310a657ab29985517da3e7b1edc7fe999d4e11f9df33e5270134
z3d2b9cb125c5302aefdc4315efb50180adf1364b9465b411134e0ad5f239bf55cd23ebbfd3563a
z99579ddedb07d381ce769d3bc7c1b00c0213ca36a0bb75fbf5d4e72e6d1f0202de360740edb81c
zcb0431758d7e7e95e039552ae800d6de5e176a422f5d96c5f13c537e199de13a51dc0c3a94d938
z18bd7fe318e2abb540d8b219e9987e81a24a68dac320e2a92e48335289b66b1f61ae5c8199d7ee
z896d3e664578e1e5460ffd4714bfbb56aab0b6e7a31970a954c04b125bf718018fa55965a24b28
z7d83f132906652e6a2b7cb76843482884169c6b41032791aa314a5c8aa6c8dc46eb19024bb9529
z822dd6df98cd5c6f6f36061c8106b5c4a4001cad7c96b964d67f49d4ea40f216eab549e12e5d2e
zc7e40e99bbdbd9f7240ef045d509e24c3d6c7bca2bbe6ba1a838f259d0958c757f9eb60612afc7
zcf210a754bbe4d3982fee1865f153108d569ef2f552ad81b99968f93052aa50fb16a81d937dd22
zbd1af12b8079e7cbea7751d90f534da96f4573e5bbbc697f23567e00b4741e127e410d24f030ab
zee4a3dc0db767e1820c95f9bc1ce12c5263998417f25ecf9897c29cb760c701184195013f6d0ba
z1ebcd5b67aa628c51c6c5c6c7abf9794ccaa88421f7c5ed74675af3429c3fe9e6162e331abeb48
z561294be607628f7204fee77f36e8ed2b087c689dcad577facde6a069de7933e4212c927c0c9dd
z1bb52ce7f8bd02136eb416cd1641a972b9ea3b14468d79e7ba10ca4b04afb976bee3949385dcb0
z00adbca0f152b5a024823e7c3257a0101355de287cb71a778e6a19dc9067fc6041e6159a18482d
z461b8465640cac11db732de5c743159033baf084986d4213943527be212f350db30a5ddd3fbff2
zc75f83e8596107824e9e572f9eb992b3caac36def929dc9cdb5729218601633d70c508c1488154
zb4ed1640cbcf544f8b2787b12c42dfa3d11d18bfd8046db55732c2805848f9b2c6e977289b1d59
z9d248010cac33a7b86a4b907cdda2a299bcdd57d33508b436c2bdabf795e943695c93f2ceb96da
ze7ec5d816b7bc8a143ffae395f986d45e14e5c0ab7b4ce0251226592e7e0a554eb7d650a6f6654
zc3a7de806a9770a0795429334ca1ff8570bd98f3d4c06da8aec16fb22210dcf2defb1dea187e1d
z5a8db62bd3191654c891ae72eb260a0529b1ce7a89e3b489278bd987d05534031dae64264acafd
zea541819a48fff2f6002a4711c0e24f74c823185dcfd89c4292c5d71a40a80da847ddcd33cc570
ze718cf5815ce32ee9b21a845cbc82b9a311243f88164ae866ccf8bb34eaf8b352044c5e60b16e2
z435ba4d152f8fb55277ea13a60beb9036fb2398be12f90a1c66e2db59187d62aad7c0ac60259de
z96679ca5e1657c50e02a4ab5acc713616fd7790a89caed306c3b7fd1799a2498986c92f714b3c0
z6a3f697f9066fa3aa1840339e1ff34dd3d4df56ecbe650a5dba850e7d1ce74571a10626d3bbb6e
zeb7cef3a61b467430b745fcbfc92b589088cfa8fcda85e0e961a1b22ca51663a9167c6c6877d82
z710f78135416dbadfc38c2ca523495177f2d7419929fccd3d4d0ce5417d0e711c7575333749369
z95b34cf3f9302336dbc673dc475d3b215ef9e60c026d876b9ad3e8c32a5426c7f5281ce9763102
zfcd26f1ca2d0489fa9a4a6ca2507af6c0ce815f4e090d13b54138630a48aeb5d1b1463daa42f16
z5a27fa13e1037b5256f9c7b8faf0cd3b3b334e0e175ee286c3b7a864b561130feae884a27b1835
z85a5a950600b234b7b499aefb0197dc33aa268c0afdddc87e0d02fd6cf2c741667c8f975ead67b
zca1b27e8199d5277848d4ff7079fb9a3b2ada048f364e68cf0399857ae62fa9b8a7af1b78ea0b5
zc88873acbca6e5eb4228f27ca7664e2a5b5f54cea6a804f506d9f1be50c1a1899c49f9f5634a18
zfacaba1d8eefe9b70c1bb60c16e0757cd4954dfbbe5f3f69a873762d51d06281cfb3b1d0616528
z30c4c1e939c96ff99d5ec9a636ec5a03c8a6e02920577f332dc840ca9ae303e94764db89bf41a6
zb0f7ef99a69b765ba09add5fe452943b2873a554d92bbe974270e68f39f5fad66d9ceab62b1072
z9a551f7baf4b75e52215261434c8f19024c03d3ade28fa721b73c6f07f93f8c1b1d5593fc6a317
z48f03b1b5933c4c0e19e84d5b3c546162fe25e6f4b3ee7f7cc353d7ea632e8ff0754932fb094e4
z9a84e2171957aafc1d01490fa0c1fd49a9bc34a47a7ce5bfd0e04afff9b409ab5fcb0d2c7580e4
z1dbd0c3980fe5208afe339ed367bfd00a67211114b5402578ae31bfd05452e083530fc4b068e20
zc815e510c6206a9c5c618520d8bcf154040a7b8384a4b9c7abcb82c904df5eaa2361d90a6e2a2a
ze668ea0ee58612f0e37b12bd86b1857ef5f38ca0223e304cb0c6964908563a1e2bed6fa21542f7
zbc7451dd2d99d37ccc4ca4e9232c826dd26100a19a304e94efb8f95252ac109d132a6d8a1d278a
z5a8e9db66c82a242055b42735440c51a66c4201f9947d6e20199ed5640458ba78b9359f5fb10bc
z9bfe9cc989dfe1788eadeeb9e13ee35c65810b07c11bdb6695de48d215149be81b08ba8e4c9674
z4bed2cc165a1d853abfeee19c16c9f6c383a7d123527ee3acc3994b7bcd9373f57da7d91bb8912
z4d82d12adda11fc8573a76db811447df872aafac843915562f8b867ee53074e84411e0c3ece394
zded26e6dbe1e2e4d1254b2696f30dc8faf56ba9fb195263e015a5131178c8df94326894dacfc62
zd99caaad8f178fe488f68da7028b40675b21106cc06882eb8df4e4916c2c7e494cb1f4f747165e
z9a3bef5a33892b8f3a6a300a1dbde8fb1255ab6e7b33d8533c56ca0a742f1cb949a44d96b69fb5
z24248b67f934f7a18bfc9d29bf49da3becf2aefc5757dfb6d7a2de4d72fe19f33846594ee197b5
z3647ba758d3d4f781cdf5b130379c6c6bf6da0b12f74472d5f7da5c0cfab8fcf01c54b4f20ffce
z196401aff1e01bd83ce1178bbd9abbd442f99e81ad6f28b6ca7270a2d307c69d8b34664d902303
zfb5e0e42c04f7e22585aefe579395eb0cb93ca6cb9ba69308c9376cade284c79e8ff3fb619fd7c
zf98735bdd4014f1ff2dcfaa83bbabed4f3c98af715c8bea18d18fc26ccae237a3b9c0823fd7d68
z19d54b803257fad51d7c88294b9d7be0350578820e2d19e55c2173ffa5ba59319deb399668810e
z277b8a56ed696c1fb196cc2693281f95e95a8f49f6bd403671f5725df310f4b78f74f523c4ebd5
z0c14e34f930d6e6806315e5ed9ef6717792e929374bba8905a9b452c9ac15759d7b73f8f283a6c
z414efc604133b1191c53d1c3e844e65a872a8da1c21f2663d04bc77851a04dccce37153b41615a
zb8a0013ae99fc49d971cc5578bd09fb484f137c62a4d0b7d9000fd551a4244fb577eb92a647638
ze0436741def1672f7cba7de089c103e7c22bfee50c1178b4221f05f77fb6d64eb61d0f2a1305ab
zc5e3801feed7ad1a3ecd8d275949abb11de7aba38a762a8d49d6fa95c8eff993fac3116b3e2b41
zcac1e26917c9aa39336ccfa74c5b48ff53b9b47e6fa38e19b3156ccf04576926c8b82c866b7e08
zf11a4aa193452a7c00ba1c688eb701a5afde3ae7687c679eb531c9cd497d42d3493b701904db1a
z142e7b58e1078671f42508d2c232b7761e88dd54c7e7831abee9a12fa88bcbad93722030a6ce8c
z0745215cf1a7f18d067f470aecc540b845196e1fe3a8790185e6012686e222a1ced8455b832272
zd2e4e9d003e6e945fb6d21e90ee78c9bf18df4e85e419d225aab4ae0e3db08b84731324d744ec8
zc960342e031e6fd25b6030dbdbcc1b8e91b58123fb039171b1e8322c80f74d6e3bbf14390178e8
z95c0eae0738bb151e7e69445a9a59a11c67476d4d8ee7a2373239cc0b7da7955387ecdd2fa431d
za437936b046d7afe8cede8c2d6cef67cc0d329a4cd503bd20291e883257c85f545854896a0e979
z1c2276fd733d42e40b3d8f6da2a5635079722f87662081d411fb48d2c2eb2b31b0bc0302c7b411
zbd6d9b2ef9682bdfde767bd3a28b39073e5bc5ffd56ce7fc8eb4ad50b2e657d9e1b1c0953ed048
z8d38b8900846ddcecd1830d1f4511301b255c6d065303cd2f52537c7df0bf65660753905319d3b
z6669dd85229c4b74188a2808aa7803bb0f591e440b2677b50ac68c95d954b6c81f4a6c077587c9
zd297e93ab21fc25046ea4d5843f4b9545dc393e2aedb045fd13bb3038de81c7227f6c5dfc322e2
z396c3894626dd6cad0795fb5556cbd93707deb63d87a91f4cbf46da50c3c319c1cc98c46f5a2f6
z185e65fefca60eaa3d679e97a341e99b1ab5b51b429fad9dc47adacaace22ee2be985c7775f551
zb18e1feb79cc296b3f0e567c8747dfcc6a2776b3dc0960b6a5a3cd917b18ff8a0ce18623a79dd3
z7b33086c724955fa0b0116a433dc9028b79e407d53f13e713e3aa6e1c7cafc119bc0e65ed95fcb
z554f0b6a66bf04b0174b0820ba447729e5e353f61481d4b1014de645a18ae46feeb7ad8bf148e5
zbe6ffaf6ab24008f07f3600e97f4a58bce311fe50b2c1237f8649068323f64231edc25db46922d
za4da90e2ae34db05ba759e352542d21ad0a5078887de7d17bf2a8c3c5559e78f835b410cac299f
z78a20dbfdbec2428efd6d7e76513a6e35356abc450fc4b1dfb74b08edc7073e09928d654f5c020
ze7ccbce4d70145e2d5cce3884adeb02d5f8f93ce1a162a6adf0f89b61d60d2c4610ec26dbeffdf
zd87b486279569cf427970f3ab088fb7eae4b58432ee169aa958b0ecfd40674104153b405ad0804
z377401991f8694f899b471ef611bd07ee548d7fb1c860e4aa9e94497aa2bd2cb0836badbc4050f
z4bb29051f320d25c4d7e344cf01813704bc02d6353f1a7bac10d4a1b7b39aeffa78f7a2295f924
ze612ad4cb367ca4f75d4b558ea2fb8fbdab49c1d51da77d0131130cab79af5ae5583e05812c46e
zc4357b9204eaf7462b1957e6059715122a9e987ff57c587318141046dc06a47bd0657dc0fc6b43
zb140bc7f3aa83d905a5ebbf7511de8e69ce26aef9e720452755b2c35eb949fcffd9269e2878417
zb256ee4840f7f31800239d0568b7932fb97edc6caf7cecbd7b4406fd48e001dcb10117505627bf
z77aeab8f46d569fb91f5bb70b2c271a3ac957e69b05064b76dbbc0f55094e5ed5806f78b5ff0a1
z7d18e28dd892990fd02b6fbbf34a5b0033c364b09be72b41a81169102bf49244e3df96091af95b
z592dab50f4afab67c3c819ece0ecafc4a77014956d9286af49be8acd665830eb482422b867e844
z6297c814f271d5644ed033b6f18cc92731e142921af88e8d330702ca273d2a29a5a18b98ab8529
z21e2754356ef86a3dbabf24d9afd995f7e1b0e636bdde0223f5ca3e3ee2417fcdd7adb3ec1bb13
ze7359eb0d2155b525ef5eb785dc3028f2564379a29a1746338dc561f7814cbfc1f5464291e2533
zc13f08e57b9d89048bcf4f09ec3cb6546e2648e05e5b5dcb6ecf3571570df4060a47480dd914de
zfffb1d722e7ceff9282ea783231c9658f64e68c2b2d8e12a3b383bc2915f950d62454ef47150e9
zafcdbabf067b5dd0e302a327a9ed89909c33be4f8bd5165f2229d63ab61ccc25f3bb6c79d70768
zffebeb570e1211848d641db5da1ab68e5dc1b4924f4ec88cf00c23c4b9c61e59e4822421026366
z15e9c48339e00894b5e06a01e769fa6555b49ce7b706ad23edfb0067e86333d572c2fac8b089e0
zaec5abb227771b77ee724eb034c61a6f0b67f151fbe3addfae1c18eae7c75a8aec8c328eccaf7c
z9a6bd455066421cc1ea9845d6513bc45f25971e188de58ba71a4e5ce6a7e32ef093bebeedd2eb9
z786772e6c30b1a9ec24f5b21d5c071e0786d96579b0a67836f6c7099782ec58d42af8aa45fcef3
zf86a0155c9bebac173a53b1b5da29b7460f11f3030af18d58df456ba6c2b9648a17469f1735228
zad05af642888f65cd2af2796b32314418918a2ac951c98ed28c375e3029bbc19968ac5584db197
zc55fcb05735cc2ec24d276265808ea5d49841f6749c73a9fc4c7b22fc404ba9d4dd7616a596fea
z8321df2cecd8d4652cc7ce22d1c8858e6fca4aa15405a004d1182a62213b6ca917ba91fdb98bdc
z5cd1ee77f55da50b30a676a9f384702cda01a8fc4ea2eb2b7fbfd443ce5540eaeebad42e64460d
z07be4782cf5d0038b088c04038eecf7fec385a84e6d65a91f8da2c7b8f36eb04e82dba80139d82
z7212ddbecae96a7e7a03eb0b4bb37e91f4415ccba60de2beff098ccf67e12d7ae4c70052c6cb44
z6a0f2f833d555d3a3afbf2ece9d7b434d829cac50dd14063766629b2d0c039697a75f40af892f3
zfa7bf210ec545ec12f0b98efecac02312e53295cb7fb9ee746c3674481aa8125de229becb33ad7
z868cb4cd78374ab79da86b042fe89cf534d76690dc2682a1d4c16aa97da8677d1cf97b24cd859b
z975cdc0ab885b9d0d4827c1a86cb6ae3c1608080c7764c2926c8701943118dfd6e762d47534994
za4cf89c1524f5c835e808557a2ff5ba40f6795248a4cd2308f42b8e29cda9effcbec930ae78ed0
z1615ba434fad873356b4655ef792b68b1c303b80f7e813aab850943dd37a595063a9f156d79525
z0f22b3f5b0910997821d148e64fe0652db671bb1a0f5e4106942d83da5682ce128182deb14127a
z7a5295cf5284878c5a28abababd8a30e2aaa0c84c31daed143f0742215b4791596124fc0e944a4
ze5d05772854d21696d7c8a9578bfc62d743083b84c26cb50d9c236af2123d52a6144bb74ef7a18
z7a02430802ff6eeb025fd6a84513fce2596ecf84baa4370f54304e23c9aece1249810e7e84639b
z349424aab44bd59b623f200f0ccc1e8b496e5975de1cf2892a383060e3bce0b689e12ddf8e2571
z873043cdeff6e1cad2fb46e0937dd0771abdd11d4b0f36c31b88e389a1b3022b6c9a63e54faac0
zaf9fd5daa04a60dd890faee9e8dff6f52827b09f67d6f26d07a25b82a35c873086e090d873d2c4
z5c5f6cf1e8022309183c4ffba135c46c8b2d575eff0e61fd10ac839e97038340ab50f12ebe510f
z4850b941bc68391fffd742a1213d09a2b851ad3330c9ee5f6c5433d88f34f146da10499f5a6157
z7d791b69ac531bdab59d02c8a76acc9f87efb4e48a07d81707411a7046c82eb9d1602313b4e994
zdaaa09b589a5421cbb860327744c445c1808a67aba45834c72e99b5e1227de28fa54ea267be741
ze621d6d974e1bfd64355bcd437a320ba7d6a4da8b3e4760ef12b91e8a6a82a5dd28b6a5420adce
z9f73b03ac06bf6c295357b7ed1bf9b585d64a04f7517f27f40b2f136cb810d340bf2ce84a1cbba
z08a5b92ba4d6aa844ebe7b229f2658d1a2a4995fd5db8201aff9b38611a69681a13927195085fb
z209fa5e57f94f660a307b9593b665b9ce69f389053c6daf3af30af758a500e8a03f00592bbbfc0
z4857a07284ebab99b59c3dcdfe65dffd36188d9cfc8967e35e125590e93c9dd02a6f14bafd4c85
z84c9a86d9bb4f739ce0b7a96f158448316a7f043123e50d93ea882e7c024853db9bd3c110ec3a1
z3ff8a946989dd5d94ae24943f58058dd309587af98b7dc1479451d03f88f0df0271ce0c14616c2
zb8fb1b15bda6129b7e0f4e94edbb4e34342f21bfd33d0769a1cf7516e58bbe4eb0b220aac4539b
zb60a5ec2ffb0615ac25c26914130ed8d777734474b02267000f5a035d50e39658a95485fcf8352
z11a3e85fc03f8ea8cfff95edc164abcfeca942dc5c2c9454dcf2e26c10955984376f80ac24c78e
z48e4a2145cf715fd26a276291dc6421d7d6179de66dff2171d6e9740ea58680d1b8ef54660038c
z18c0fd4ed6ea17281bdcb72f277624b02b0fdb0341b573f3928dc1b9647b6a4cd65c65055ad334
zc5435fb21d105c529e1b2b89fae5ee1cef8f0fbdabf3ecbde7b97807861de8a8f9b0a9c2853a7b
zb2d49737d471e672808aefe1021d0f37ac729ceae3375cb54e2f64686be86e518dd341a6a65156
z316b6c009dae28e2954f6736adeca9937a7d5100d5864a881d2dc2b5b7ca4b2badbbeef4948321
ze15613b5e51aa3c60e45d2504325df16d380bd4481c4fd13940e73055029b953e7b5d390948340
z08e9522429b3ae7417cb727b315ccd0b382c7079a18d09c8e960fea7ad68b797744909836c82f1
z9b3bc8f3d853548dd7aec95fd23581447fdfc5153d75cef9fe4c664f6fd98f1c75dc16676b362a
z5ce3fe49c202a7d0961e4355356246a1c510e0978382970e4941e4fb668b85d00b27a526351f23
z1de8e9780957ba362a7df7accaae069ebdf7d80085b4695ab0d2bf3c907a75424f078d9c76d34a
zf287b83619c740d221e96492116f95d67629828f46ae1c8329a9b38d7eb841831fec42f56d1079
z39883d65d257658fd5f17e455a37677fccdbdec77256f8a57b5d3e7e709708b56217c88698f6fc
zd5abbe10197a3bea9a9a7a848a95b6b6588189c3213f85745b386e9242863b15194e846244877d
z6f81d538535505e37727a52f8c645b9953b91639272ccf9bdd8d8e86053c5a824dc31e41ede3ad
zf1bf979619d22ba000e82123039c32a079a5a5e911943c0dd329060d85042f0f762b76ccbf59d9
z7b23848059f4bff6995954fb98b8e765e1130104d40824925782a513a9491d17ef781193f7f48d
zbc11161c7e593340f5b1961fc440f133e73272464ae45e98aee4015988dc2c4c1ebac22730421c
z7ed8c016b4d4a7973bba9998810dcfff8e53fe8e276588a725abc186fb27a812fe162da58750e2
z605942f50fe290add83b3e2fc5392d6930d136ee77d1dc2d35d27027b6cb2cbfe5e16e2f38454a
zac5d7187775749f13c6631d386f8bc5f33ff2e99ec4ee47415309b986fe18521bf5aa96304b32d
z5bd454da6ff0d7ba7d4c3df708322c6cee035eb915f36d9d60633af3a7bf82c77de8a2eca46148
z47edfc6ee6947fd6dad90ff8db23b5dcd06143a386a4d7f2931402a58f2a7cd8f4c78352ac3251
zb97ad8a581fb7a20a9e51b90bdf212967d5ebbd8a96ef303595c49b9e6bc935f2188dd984090d3
za119052f1cc70d9de755f0f2a97d731a7098c4c29227fc9bb19dd4da5f66df975daaf390571b9c
zc20f9c799abc2197bbd5a39e0a67014ad5e6f95ee57ba285842e6cc4894c3ec2dbea8cba23f02c
z28c95ffa8f51f92cea0c2adbd6b1b07a33fb92fa19ce7db763d108c902ca5a46cb9cbcf2997a6f
z73224fe7f3dd6d60430beca1105209c55ce0f3359998be7bdcae3f5ee34ee55b0201f623f57b35
z342361656a0f767f4d9d8a4b1adae1ead8926c9129a4f48443f4f1cde46a69fc4e2d2488f82740
z602ebab52128330b89253f58dd2df0efea06948bbded31942a99b524bafa0022798ab0d8ba24e0
z6d683531739228de4e72a729c1b1da6890f0f77055567f298a9cda333039c04326efd96ad120fe
z5f0276821ee58608c3fbdcfda8440ac42ece1392a52ab031fed7d5e011bc61bbe8583866c50daf
zeda634a8c551e2a2fc72c3c38664f9eb2f9de015642643532d2ab63f088984d7f97342badaa0d1
z4343c5365ca19d2fe9d463cc612bca4316a64cef79fbf7b206a0449cf64f8260540b0683889cfb
ze8946213d2831cf94fd4993258b0d62b755f6dac044960b1d33ba8ae8f35dfd503f83c22521575
z85fb6531ea0e026610c4cdab6b8f1233c7a026feb3b56854dc1cfe6ce58b23e43f6df68b12bae7
zd0f813f59c4808d4c69335120b9f05ae4830d10ea93cc50121bf26ba88e521876a5fd5c1361421
z415acab06689f6a1ec30d80802d2681d5d4874f998a197cbe860113356b111f4145cd9796a1156
z932874db2437ae2d1778d621d4efb5f17f2cbfb6ff03285ceaf9fe4bd9eca801cfa772fde1b4df
zbeaf2119f27c74c5e7ee90b13a0f776b2db7528695b699390195030fc73ab59380b63142920303
z5ec0e01bf06e14b92ef55d312cc331a8fe8c012286d89df04ce549ae6a3b473ad2040525ab7f7c
z8137a61cd80980ae8ee6e8dfaf5aa6773e823e2a4617305333e94a3d37c4bcfa38af2ca14f36e6
z1297cbea8777afe0799420ec0bdb83ea101cf608deec9c8355b3ef6689b215dd5bcd2a2be14871
z0756950463fbb2769bd25e6390f0b4854a282d2b717297857046c734f4bb8cff833986a8ec6fa8
z35149d4e2ef537f9eaed90b8559f6309dad0e21296cc4f3b89a6cd0bf22cb47de269d770d9823f
z4b0ac5f311f153d2d71446226bb193c1dfb92729fad88acc9aee9a316e265727fcf59b440a7446
z4288f34a8ebc1e4b7d25c2a7627e364b53a2a216e95370a26ac436cae4ce2341efc12bf75530c5
z43e4a619262b92cbb2f6daa3126c1d48d3c7cdac01e675f611a2f470ac55491a48486b88548936
zcfc56f3b212eb9984cb6a01c9a4ebba655ae59dbed394763ab13ddc952e14aeffe2e57a0230aa4
z1dba639b294c2fb0f1023cf9291a04b4cbf3c3651223c3ff535881ff76af1bfbd26845e279f124
ze525c9b08c16c249f85545f95f0a62831c823f7bea607e9ffe5efed31d7fe8c1b773eaf4aef176
zdbd1e1aceee4bd42772b9de82f5717733352b9b02f59182d87e967584b52b1b9279d4a6a74e315
z9cd1a2292d7c6026dfbbb2b07913002f7f8d1f7f9d9f63e77b11f7c21114752557c37fbba75839
z9bda4ac27eceaf887225bb15d37f4e09e527458e1da6f5d9c713c3b90ad9a8893a4e79b58295e4
zb8194132d00cf69d0666aaa3dd2cd20f515df1348b6040eeba90c7ea99ab15cce253782055af46
zc1d2f0bf27ddd2f34471b7700fa2bdf73deb85e1e8c84c96dc5256a9b6aa74e4d9a301761ff71e
z558bf1faece424c9094bd7d4e3752d2848da056000aa72d590b6d79fe3ff9bdc17292f9479d446
zc3093b22c01f89349bba26749da1a53c136a56f1b44c8af480afab70723b7dd6bdf313233f6e9a
zbfcaaf2f96398bb5107ea0b599d23e3303e7c0368bc3ee814d524e85a611caac95a5bb1a72d362
z1e0138e4b30309277298c86ef1fd30e0c69291f981f761b4d3a16ac39b54d02916fc877ad7e2db
z578d8ffe11c878d86850d73f8dcbea8e54c3b72c82619ec92acee70c423d222b582f6f73e44ab7
zf3a3ea60091b84e624d007f034d9dbb7d505ef3cb596f3229ca01ccaa9b4f099bca1c55e43257e
z96375929abc19b33fdae9febc35c332e384b183d55549f150f66ca562a5219bea29e189e1bb9ee
z83f8e22d5b5daef3f827d03751159cb5e386375660d4e6ec9aa28b90c8cdd6a3b1bdb39ea143e5
z69c83a2fa81280402c775b30e941060858b2fe4053c0468829ea20c88da182fbde4dcc8935891e
zf04287aa662833fbdb9aeb0eeffc0883b251849604d54b4287984918fbea02ab23e6eb2fd19240
zb9f9f14bff3427ce59a5fc7b433ddf53e1883bcfaa3f5d25535100a7f93e265e17de3ae7dbc2ab
zc4cacc064c1877b1655cb3cd9d059875672a3ea2b340eafbfc3c4d039b506c7b611b23f01cf798
z5d5f6d2f36bc0db04fee26265603fb20db25e34585dd8aa87c14ca4623aaa52202b5e5dcbb7e7b
ze0c52c508fedf1746cdb5420ca7bb3861f1bdd70cdc68cae301f0029c373112480624ee1d87eb9
z3594a0a72f76a760882d176d1a7171322fba091b8a1db8ffc6017d6d754f106fd24e5e8854a6d3
z51b53850ea042398d5e3d7436c27b38a0f790500152ade80fdb165523f700238ad72ccbc3922b6
za6eb9835d2c50e26c9431f45814e1e6b09d280a5107e07d95fd28241a7d492f152644aa3fe8a53
z6b3178b385e2652d6c56d80c5f73248708dafc8361776789cf1c45fb9f00164f7812615b8996c6
z1940ed8eac435768b7c48d55c3cd3dd4a38a6071149149b67c2edb09807158b89485ad293171b8
zb54dcd4d0bfbdb058dc33f1a764341fafe6cc9407a590976fd0de94373454f623305285a7836c6
zb0dd7d51f7b820bae96962b5c8005dbcea1989d2246f22c83f4db6f68fda19ac45089e9425aa06
z9b3ada68cb4f338c0ed511c2fef1a0952c91600de4e6a328de340e605d9e4992e40696f1f8a62f
za9881c8902a778151e4ae79ee17b293f1b2013b20f1fa210bed60c5816b9f427ab8bc7d8011616
z064018e8aeebd4c1869a20d6ca0dd206fd952c6316c51e1196d036fb828bd27a167ee9d04f64f5
zbaabf1bfd5c65c4c7003a98240c912d5b801fdc4aa8ba49b4be978ba1448024815ac0a150bcb10
z50b48d0b864e874267fb0233d6475442d0367c8037c2aa49b3b27aef4dfc13d356ad7ead492c8b
ze65d75a94c8f3ea0cbf01815711cde13900502cc67180942235fa00d4a2d805f767fe734c66d0b
zd910f117dbc9663559038634b3bbbdb5548f1d6157b0f7059ae7b3f26a7309165bf57d23a2b300
z51f25d88bd2a3f22014601d5412f9a7061bae25df21ae91c62c3236539252fc7618622ce611fd7
z6e0e2f556d5147e3180baefb01c44edd0abac1b05e9f746917fe309225676a58a71941fc68d764
z3bed22c7c333ab75dc82a99fd38fe7fc835f40300f24b0e67627c4efcfefbc0be15fc46f0fa955
zf8f2dc9a2c0832a8e1d365cc9893e2c68df84a65c4dad6b449ccbb22ba63c17977d6f09e1d8b43
zbc81c44ac31b54a6d882fd1adbe012eee784b9e18a61a65555c7df8e93d1fa0d8ea76593366719
z01a498de55a352c9e3f790bec8d7f4c59c55efe658900b2e1d56e3ce3434122a1768892bb66223
z88c641f26115ae1eadd39d9c5a5fd083571a51aaf4b2ef7ef3d9d91a1a9fa3101c778383a235bb
z8e8db3b31360720207e4a437954070e451c50564b9ade7db553dde2408e8b2549b2405173dbf86
z7d7a8479da441560d51d2af19c0cb46e54467d27c1335428bfe0d6a2dbba142e877960b94bba66
z0e40a8dfe4f3a4c016f6741437d71d48cbf100f769c3f0cb7b63da343af6811d23f5948a7983fb
ze6f11e0b07a5c7b5079996f62865de6b273670906d36206c28032bb7f2965c7ef0c2ba498a173d
z8e82a44ef252004e122acdd4169aabc4ee3e9fc7185e1bbb02c28cdaace2b50e7e2806ee1fa48f
z3188759bdfdcc099148107f3c4051fbea3604ef55061604c53292d661f2e3e95e86a548c880357
z1c6a2c08efe26e9ad6ae76dc0e6e824c17325877a0d3a596f2ebb6bc33244d41013c60c54c43d8
z9e4c400c2ad408a625e355b7f9b120ad18f1ccc0c52b0ab501f79edf29e66009259592e60d2335
zb5b5e28a806495322d144880f23885c82d733b59f4b071c4f969c7228cbf483dc8c10ee61ef2c7
z1a25fa42ddb58287e1d2fe0bbec47c4eef72e85f7785389e0da6181fb3d69b3fdb469dd52c2f86
z31662bc535e951c3ac638ec4bbbf3676584a0a6e558a6ebee7a57e309874dec00d006189898d8b
zfaf8c5bcd8f3f6db3b253ee5344eb5b0595087dd056c653dd598a4fd11efc5ea0930bc5e81883b
zf5723d1da8ae285d6403f21b46f3158a22f1a872909a2e1a559b5dbe72a139fb9c95bb13e7d9fc
z25952493f9c3b6ee1dbf5589da15f9366156cb136dfb2c17caf99a0adb7d9f976fb961474da5e0
z3d17b21f361b38552f2181299a45f97e54fd15c1bdd76905eeb675b47d9ccead9fc0dfc1cd3e90
z71fb87ce60852aad97cb8cba3b648e6c62801a0c35111f7b096439388a78da45d3098af18c3119
z1d74cead613f3b5ec1e15ad128e40055f2db1a076fbbaef775f5c1134c6df0a8740861d8d376bb
z1c2356bb07411c7f5f865c60699e26e444827d8a29c14477add4bf28f0edf4eb9eaf9b46613a7a
z773c012e645431de2d7144f6d75f46ab2a60415d444e8643a1ce82c707afa4b4e376aa105f10f9
z7e3bfc98a5c0c5228dcb99b18c49f1fe475515fc309a9ccc1b312b9941c9604e797a4fe4fcf642
zbbd560fe9c31a1982d8c5d09379c1a337a0e03d5aeef78799b4631034eee7365b154f32aa538d5
z468e7165c72997af97a0fca43e390634d240f02f0a29548f926aa920122cf2f1c45a1615ab9816
z6cbf05fed6476ec91ce46d4c4efa371fef5285351fe43bb6e4f8f5a2da9fcf240fee3076b4028d
z70592f169788cff5a24a37ee50954182ecaf81798f3b409e17a97b58c22899f2bc8d79c3b64c21
z00c465b37a0379771de2ef054d20c58e244c001155f6701f0f16f6352047572ea4f1670dbfe6e9
z8032465e9ff5997973730b9fb20c127f23768854696452e4c139a1ab82aa25f511ef2aeece8205
z96d338f30f0c134c78ff9020c3757f57646e304edb5b67003771757b8443e6fddfb9ec1322ab53
zd6c760d7ef7ac7cc8199750f1775205e34ec9af1add69dc5b14a675ab58a97faa3524596a7a9cf
zb7015985d92d35834e41a68445855012f075565d62dc191d9258a44cc9f9690769b7cfa33fb7ab
z94912d9b9ac9bce5d58cdb183e9ca5737f42f81319e162258e863df8ebea0d761349fec6fd2d10
z4db47930dd2a44d3c9145c7eeb8ab047460080ab3829c34573323af3aa5793c2119333b2d66c0b
zf09d860f52c1f01da5078a72586f683841e2a42b17400aa8077e080771c371b00b1c06ccaa548c
z1a7bd867f650ee7fd40a7fa8730b71c620bfd02fdb9638eb79d0798a018f99cc8c011a26650b63
zd4842d09475aaf6120a25b41b8eae5bcc898e2d19350aef6f890ac65d068a023b162a93ffd4add
zfdc2acbd3506c2ccfcebed61b3412717a53ee76e5dd29c6ff8c2be894392b624d81f1967189be6
za1c2371a1393d02d6fd96ddebd1c962ae6058500af992418bc677b04ee57580367a9a2aa2a7470
zd00919d24aa2b82978dc0dcb20ef29fcaac747459827adac4aea232d1caea183096a27781dc798
z2f89f130982bcc855a513d293445283915a01b123be6f67da67847437f46e6e628f60d1c3261ac
zb0b8a7640b9d0714faf37291c0e52198da0f2fd6a193142e49303ae0fa5dc137a4770714141708
z4e8169e7a95bff57599a81d143c039a251af481339fbdc31a158596c5b1a126e42eb05dfaf8e60
z45d4d1a3a22a89848420fe1d251082a3d623339a897542f60c01b329b4a3bd9405a4ac20ad18dd
ze6a65b93081ec4775d1ef0ab4174a8f369143130431dd01110461b9c41f87188d3b79ff2288114
za2d5cce64baed3376befdb70edef7b3e617ef69c104b8dcd8e344b98dd7e509b0eef1697c25e97
z993557b63e08d22c0ce52acc993ca9504fa99ca5e9252f8dfbc4988e1713c555a1f7e0fd3bd6e7
zbf867d0ecc4d98d5caf0a440d1241f90a70720ab365abe93fc0d5baa00229dd5fa215359996a20
zf673ee9b67fe4ec9ea32d3a358be5c544866458d60f91c25c18b8a5f2fe75e9e937d3cb399399e
zc1aacbae261836fed9c8e74b19e1f99b4ce5cd055cb79933fe26c32436cff125a0ec6e48a477fe
z4c561d5898fd5eb6bfb6b98471d76189ef80f9ccdcf18929c5d73893f22f88d40927536adcebf4
z7d8dc213cd6d76f6a1f74dd567dab8402a895b3f6c1bb67cf06650f3cb9472c5fa5cb66d840963
za3e2c08a7c86ccdcfc1f610fd874bd1de6f4093acc52ed4a01bb629299a2941bc0727e72dcfdf4
z849306a5dc0628885d5bbd3ae3fca06caa18d78b65eaef1bcb5dbd7e7e9c56fb2d9ac35804c0ad
z879b83fb8e3dede00c19b8a1888ab3dcb8da2f573988030b3c0d09de4e641dbf5c7bea7b4a590e
zef056d0d20221b33609237ac423a1d926888a94550f810ebd496440f1b54f7b71e6458b4abb964
zb7d66981492236fbbdf4ef171d2d8e3b7199b946debf8cf9ab1ea0e335a9a2780ed829dea93ef9
z0272e265e43440271c11e5e286ecaf589263c4b5debcc1882ce0142d65e537185cabfb24a6a8fe
z00f514b332e3a2aad55b00822f1adef9709643a3c284298efd1420667a67758bd5c747744cba77
z9b99d10bb0791a74a5f1ae3f5290f5c9dd1e86faee218fd61e3d4d93ada16d551f12eb12f0377f
z29d3535191ce39c3878e61452aad22c17ce75c0e2c8e6f05c5d8e4c0fca517cc569cfed82af105
z778754d70fe3c69aa216a6dc9288dcd300b85da3ccdc173ab4e0da4330b71ab54218499af73291
z5f4a1c366823be913af28bd73cf30f2d1f536bf60c6d9734b78d1f3e027eb5f10bfcf059daa075
z41e38a6ecb896a71fe1d53a08951d93958ac9f9a2b369b65646143e863ca5ec1779216f883b9c2
z32b17fabdbfff9ae33bbbee3a02a15ead136a7bc72fda26be39b5c4fd60e3033933377b5425ec2
z84ad84a277bcf70347c2b8dd0d544a9dcd9e423588fd878e77763faec1f3b529f9953fdebef9bc
z0d89f8fe3eece58d15d4d96ff3587acfcf18b6903af87c3205b3c01029ee87cd9120490d6a8545
zbde8f114293e8e66697bfc6dbc753ed575e54a5fc602bad730bc15b609ffbf4a2ad081ce4a9c43
ze0d2d8fcb6e1b2aa25afc988d9951c58a740ce51b0dd76de9acf68b02312c206a7244aae0e3ccf
z542da4f9b4e8f5d6d03b91304de2d9d2057a4fe020b1c8922ccc045fe971620a638846fb79ff30
z189b1564c319ac49e4d9087a1beac3930e175fd9353e4cbfad6a5a3c55a273f6ef27789f493d03
z6bd254f0c836500d4518962ff0e45bc72b10b6373382d9b4e9f1061a2d2e01cf7f00b9a022b65d
zbb9d0696f867a77301b84f9e1cdcc8e8d2abfcebd03cf71cfa607772a7229d1ad59c6212279d52
za88716843964b52fd972f420d7e49ebd8b8a93f56bccdf322b4499afbefa138acc6322e82ccdcc
z1516dd526d9c29189cf0a2c81117bef9da9bb1f0c9ff302cceffc9d3014bb40b6ec387ca242322
zb6b252168294e54cac5ec056bf7af69bc78a5b22caae120ba68609f34b38fe143eb6ec8622c142
z0186a9f6941e71d7615af86a6d334b66d545809df8d9ca639fed62b4e47792c9af9769dccedb9d
z35930ec4c332449db6001fb3ed595976731c650f547cbff0b2a3e54e37ad111c178e7095ca5ca5
z5f6679bb1333cc95279afd8c03c0583a78222db168cfa3f3abd446e8f2926cbd3cf493f8224482
z2d29c6cdffcc33486aeba2d3efd5a8ef2b861f7b7081ca2b8cbed8a597ff0eae7f39be889d61f8
z9d2b4678d15ca2010ea3bd3cda21e88267dd8b65746a996c89f2b83947836ce617e6ca05f56a45
za40acebf1c6d34f3c268caef74222431e9350651c3782d1a6f9d7240eaf3403d067b3958747138
z27aee7faae6b197614557f35edc445890344606f912ae34bf22717e68b9aad197a228298a5e7c5
z7faf52b64f4c11822301f5025f6c61109e7d09d5e4a6ad051e900fe98c9ad1cdbbd7e3455b6857
za75da7f0898acd1f4e07aa8cec7cc8b3f68d288059ad23e2a011a11e8ee26484005f846c2c2ab6
z0633bfa439ff2958c358036c3b5f8aa229abef8c61936617e40e9a6b33f9417df6a14d63e8d7b5
z4815e8e44321c5e868be6058c486dbfcb76697b718499246349e37cc3fa82107b7b5e8c9ad15b4
ze6cfa6af2ba11e46cbb623176f909e28d4cf077661b48a6089bbb1083b437b63d561bee7d3af8c
z4f07826676703ff53f703278b39c123bb6f15f398868f7588a99f9021d091c2b9f6dd7372a695f
z1edd59a6f387d3bb0d2321eff0337e200f2a3cd2f59c217c6acf84c30befd779a2cf802098e471
z9f83b08f7bd40359c913f326a2d64513d5127c7eae639c42df12834d16d3989287e5d714bf1d94
z5d32bf8aeabca585d49c4dffa2e9d29eaa300eded833cc2e9994951f59f9e5579e0986c91d2cb7
za7cd0de3c6cff97f3e68e8ce91f0d45d4ec891349595d6d9142ebb00547b55ee72ee48dfe541b3
z114a6a2a3a37e213e4581cf46dcfd6e00a34b524fc71cde6f8e508bd99ab7b631b9af0f267186b
z5a631d9ea08dfde0f118e3a068832342755d3e7e115a529b87af2006363df013923a0425d965a4
z68defe74831ca2937e15e2aa23992c399768a5b3c7466cef32fb1d411151fa0b24d4e5d2ab6b18
ze555a080809277e4d6ebe48d0ec4046404f1b5b5f593af824ea9fdb7a4f2c6f8ee3fb22d73c61e
zf9938eb90d004bcf450154afee78c4298c990f5233ea6f3c5f2c0ca39a33b364ad0381d87b6b61
z1b8ddbeddd7c55bc806dad4b780ade347a8eab4285a0c2d417bb2af19e3842d411d3defa4bf949
zb64c68fcbcd8f86f87189f2bae8b2bdfe62ab1b1570990218742b218bdf7b790b6e4ac2a696648
z25dedd2bdc9ffd95968725823a5605d2c5518971f349936c9691ec5a2ca2d7c31e0278abccc91c
z49e331410425858c67fa28938d0dba5cda6587ecc9349adeef6ecef762da71ebefaf7c8ab75445
z0c578eee35a7baddb604ffeac41588f7de59130f9f05c9067afdbffbee91399b383d876050d473
za44f86fc37e0165cb4b9f9c8cd99fc637f58691759dee9790fcaeb30609489f3b64641b37d3d8e
z7d14af2407bc58124c854e10595ec3394df97b453a8474b34241135df72af75f80d0270db710e4
zaa0584d84fc0dadd1ca16e61311bc2140e29862ffb4bc014d6897836aca1b75f2a0d85e578a3d9
z8aa2add05665996565f974406cbac0143ac025fc0f6dd5144dccd90be9b93807f32ad023444789
zf273ace3d9abe29012dc0a1c76e8c99ad5b0d83fae654ff3736e154db2d04d1ea4a6c24c29d97c
z959043199660bc8673d23b1e944ae1597609d87156a205951d0c0759ae1ad80aa885c6a43fd4a3
zd84a5a5af0b2b6f7b1275a4c023693043358b3a570fcabe6f98e50c44656d4819c213e814932c9
z634076cba0b9356710a46edec0d0757f0f77e223bc8b7abc946c88faed1f6f5ba8e5264e2766c3
z8a02bb2e8d35160d2620c607b0ff69779dc5c8c548cbaf77954a20279497a63b17f2870cad3005
z5028a70b6416bfe63fd7984f61b24d7d64a07cf72b0ea495ac64610eed36abfaf99fa335ab516c
z7b64f1fa3ed92d512eb723e0b07c4d556132cad18131e3a4f38682e7db3eecd3acc8c21b6dec01
z2c75bbe4fe4ee81c92770349924ebeabc2bf2924a27b31c7cb545b3a1631d8ae654e73ac20f2c4
zb643cb82c71d7ee5036269a227412394213e7348e93a4cbab8030aa5b0ed8aa9cdb312900251ab
zfe91262a80e36ce712b3ff46c090a794f2e7ac9dd457b24d384d9de17844dd8a4df8b7cc2152e3
zddcaf362504133415013193c19f6214fcdcadb7946e54b6e76629e2561ede9169f8a788ef67556
zd2ead5949fc049fc38b331f233418d8e4669153d50ce4dbecf81fd83f274ecf553a7000e209d0c
z242f3735bed84f6a1ead7290a1dc21b99c3474dd8acf47b6293afdad3c0c8950c4018eb20ff52b
z95baf42f0f2d058794ea95bba50641883744911abd6a8f9f19f5c247d82d2963750db65a45b049
zfcc52b88f726f58fc091b390183c73c4f79a81b60c156852ca15217699e0d55aae9438dce676aa
zf3072d13c18c34b7e37255d4d2bf58d7a3d05f5a6b56a5a335d644e82b2d5d9873177f468147a3
za1e77730198c7efb585d89ccb5ae13421cd340fd4582b6cefd89720b16ce20694bf5beef2272c3
z5970ee9c83a0f06d908b56cc21fac99c4d4132027c1572b6dc440d5a869d6f7260978fa629d0f4
z3faf4c1a9e3d4e94f0adc951e99acb5e1e32cf50c13c1eef2fa25aa966cbdad5edb1ae3446b40e
z9e176fbb4395d19faebacc5814633feecfc101662ae9affe4602402d3bef114a69fe1a74b31384
zdc1511e6ecb9a529d0b4ab7dfc6be50d500c3b7a3545db589749793a38626a7be8557ddbbff611
z48e4f4194d12044b6dcab1fc95e90d6132faabc95471d366b2672c7f23ecc8fac009882f5c32d0
z29bebeeaae69e7e7c668ef09671682afbed5358b251c95e74f2e2e065b56847b323dea6d04cba0
zc1b7329a4656e98c5d50e1c7b846361e8c7206fa1f0ce1a1c0008497582fda4befba1d3ae0e8b7
zd0404d2681a8cd46dcb270595b5dc4edcba804cd5262a1f1e7f0141295fdeccf3ae3675791022d
z37716f4deff33fa46228379056853a200d237a3e3df70616c6019d369b6f2a195a063defaee4ac
zb3b8a8a67b7e190e46ce8990eea96a1aa9313b72317b0832d2316ff28384b219f18b85eede8f9e
zf74eb18783da3468b2977c61f8e04e7e28dcb4c076d47f16b242acebe68ccabb91afa0d98104f4
z1b973cc03afde0a0b3b4dbf34c37ff293f932430bb28e7005447220f7df6f30def0bc0ee3912c9
zb88dd78e6db7ee06af9a22e0ac536b7deace6cd5dc4d0fd6da90f83d902eebf8a183bef46373ee
z4d26ee671999912cf74ecce62d0abe12b2e6dc360917ea6eb3b2233fc1b67c52ac9103c15f1780
z7ef4359e2cf557f216edf033146f82b9494190837dbf122bbbe14e2f6c511107c3f18e2c8937dd
z48f2c5cc4986571e844c6aabd3b599f2920d9607b87ec289333e8f817a678654d105d199dc19fb
z0d29fab6de05af374c6610a3e8b91fec6f0c6605c031063fab9c31ccf52902ce03466a2ad0a2d5
zaa894c4a0b99d18c12902c53eca99d902c40f4fcfa05b8c3f4583120fd69dd40137fb5f99746c1
z3a9162ffc2f39bcb75e013cb23d0bfaaec714c66934f933abf3eed770f02f5b8c3cc260f771f09
z30f9cc3838d223e51b45e826e729c433cee63e63cd5c9ee202861dc340b19c5fbf466f75eff1d9
ze01d2d50187c3ea2715dfa4d61f323b44953ecbb195963e87e3c7dd0bf5694612e36755b76c250
z1424b9abb4d6ec2238efdf44cee5a92d1935e4a146302f26113bc1e0e893b626de0d024ac7decc
z366c7ed3aba1ebecbf4af291a9ceab0d0a4093f3225dc953ea069fbf1c18dacefbd1b0d814adac
z476220798fe3ced1d504842034079885714abbb852e5c2911f9b7cb71165e8acbb8f18d3469c0b
zc7821e43926a1dce11be33c629ef55184a5da7bdb76e7f5c6578452f2d9073bef477c037f5bd5d
z587d7f5d2598d1a30e7c80d497943e67050e9fa56cb839623f27d522a05256495f76465ec67290
z81e7457a94c9c361d872f489462b8a38b4b83aaca9830a42b95a8d6c0423b8515a15d74c54f995
z2e21ccbc2753e9de3e9e08820f331309820b7f1102d4a51210a539aff11391aede0214ef7e5c40
z94ed86f18be464987a272dd1e843b091d85e8577f9ab2060c22f6e53e16a8e3a1443abfe47621b
z1b451a1823055d87904e63bcb26df0c28447da3a18cd2c573d2cd8e710e083874e7832105038d1
z6f43f9dfaee35c1e9743d2a5978b04578000c047b8dc769d4b684bb2dbec673cdec7a34bf2ca8d
zb47e0989389ef124b5e1bd61d1357722cb2c9071681235212650c1bf852eb2e5744a6b1f74cf62
zff83b0dee2aae8228fd637106e71755439ee7b5f5ef36790facc303c15b47612fb4f40781763fd
z0b8382a2945f51fe0cc57d3c529ff7f1ff11c77813854af0727c634c34ca62e4bf0872ba25a01d
z1c08114fc6ceb5542802fb89e870d8e2202c4ded35e79d31ff9a2fd43901011ec1e6327e720fa9
z7fed8f3aac2a5a762a77156760a52840d39c85f0277dcf8e92d98feb58b269edb7a8740b75b7aa
zc4f0f68211e69df1954cf9937a56efda90ee7ae8f70c36f076c51dd6e6fa412a5bfaf56aed3e8b
z971b17cd08e5dfce26be7bd6e3193c1edbbad081567741645a437282ad9d2774a150525460f97c
zdd084ff91022562b2ff607afbb5b30ea4ef67cfd881a330442673a90445913add23d663e64d411
zbae3913937ba5b78ed6abc64d8f8dac0c920fc72481be52d4308f1b3df01e219b6f6881bb221ce
ze1b2dfce5fe9d2b940c3986e4417de4098c87aaba05f356ca0f8c598e73d249a5074226de45b18
z60f2abe055cd5a4c43c88296f48937bdffe0dcacad7d32697cceebb20b212ee20b2cd406688b92
z37090757a5042578990288726b013ab526eb2c346819703d5aca55d9f4274816de50ec81ec16cf
zedeb5fe92f13ad7b7e3acb05b24ad57c4c7e8009a1ad325eea515d3c380bc97b1b847a44ad1bf6
z93dfaaa570b8a3a45aad0949fc1c3a2571073f79d03654bc9990e088a7c1cc98141a547a17dc0c
z69e902d00c49976a0c920e163d0aafcfa229914ecdec4ebc40bf86fbc9ebc078eeab3749e0650e
zc919620ae97c9ff078ff5d56fcc51aa3a830f3fe25ea056d93b8c6b097cdda6dfd793384d74581
zf99cc23b730299d56a9096dcbe5b227c116f27e3bc897bf9395bb34563b09e4c8664635a6a2b6c
za72c3c67e79934da4e24a43c8d4f3f609bf49e4fc40a566a8f681042d81ed1ec00f5e6d1af037b
zb6b6a8ced519a64fcb3320b186437afd83e8d2288b83abd73036379c1a94a9e02dd4a9d80392ba
zc79d454a867f1cee35c50b6d68044eeeb1e1d1cbff0aa52c0f04e87fe33c1fd253eeb6d3156a83
ze8680c6bbfba1b90d6baab9b5fbe373e3a184d773e8850fa30630ccebfb1d655351b724d3872c0
z4b2e97f4f15da535e75c14faa4c79bba68f1a49093e8c6ba1f251bc2e6d34a2e2c390c8f4a17f7
ze82498afdb555475445c27a42c3e671d20e23f8d0ff033ceca47e9ef3dc7a96651e2af7976f885
z6c77bbcf3c3bf2bb8240cd3b63d4d3c56a9bba3d14e20370f2dcfeac73018fd5aa2a2a64c3885b
z5cb16fae337e84e8070a791f5ea5abb07cca8b82e8b4f57cbf9771f1c13c4374c89a0c7b0f5ed2
zc61e49110fd267220558c7984d1977964cb02de8f22254e10238e43760689e4f84fab58e3337e0
z5b35615681d40a0c651ba6290f6a9b5b627b2929f5bd6c7d97cfaf204bd7ed4af8b76b88e1ed3d
z41a1776c7ab052c4d7528e9674d7dda4449a5d3bb26d1c38540066adc290468e283962a13bb724
z8991c87208286c79f1ee738b3e46f7a109d1f5d8ce019a44b3aa40e886b27f06fdce7b6e48521c
z39c97c4f8e854b07e2c7a6f675b450fb3a15a5ad3610b118b14678eac2e08f6f1c5ccc5db3f79e
z4236e214b96fd2f46a744bbccb7cdd5aee166f93c9ceef8aadea8633870a1a50c16396fe7268d6
zbd6bb9b9d9c9e8e4f8ce5f3cd1d3fd4319042bd6cc9ac3ee2319765df931e527f5f3d179db5b41
z3565c09e57574a640b88115a31c4a63cd196e3a97ff1970cddedb1325894d9d17c3cf37fed0e47
z88fd69ecaff82eb9d33aac3cb54289d5202a633b607a46322355a89fa9212836951c1dbe92820b
z93dd251ecc752ce5da117c9a4bbae0ecfbf17a5257d30f4dc8d66717fb4e38bd58dbdfc7fe2fdb
ze21afe1f88c28c886df2fe89aa29120a31cd0b64ac6208e31564ea60860160441847dc8f053e27
z5451caa37149eef29e3eb556fd8031c5f84d250ba4fa22e349e4b53b2695ef417a12227b2b0f27
z8b542400f4054aa8412a1c0342e33d60fd4065950cb1addcabe41b68578a31d1e1226d0aeb3598
z6cba3fe1b074e90317ecfc64376916ef5d3eb59bcf50bdbcccf6cdeb096842df361eec6510a39a
za1f6da1bdc21f273f484029d43b53ece04434147044fd651298762104a013959bae76a619d2077
zed68db34d7e21b244a8dc82b56e05b60ea6128ef7bffa0275874edb6043f71910172138769a421
zcfe90b59cc40e8be90f086bad550e193371452d1293028525c92f30bbf21125999abba88fba232
z68876f3a14667c696868f0d454b90169cda44ce6da7f572f3fb8e662457c5ee455f8d9b42414c0
z0bf32a997331d0846bb448fbcd04c4afd4a755c9518b13b9875ea7d928b7ea8d0a565c4434ff77
zb3896e4c5bdbdf88531b106e9a3bb5349bc03f8ba9f401389c8751ec1993b617aad581b68d3415
z03b6b9728d036ac1e0efb854f32d4e289026cd4c2e906eedbd2a632625cd370d0675d47a53c978
zfbb50549c21a47e22a41e1060995c2c3dae44877bbf8780ef49bb6f66481713995c57acb382dd6
z629a6dc0b7661a091b711c821b0f0991b8a089987cdba12df2b6dd09ce8284d586d6dc31af7e05
zb73991c8dd2e0381e6bbf21f08b31733261ebb3abc10ad866d388c2be686fcf0a3eca9698526f7
z3d16546d00092021ba6db9576a3e43ea3ca405f347400896b94ccff176f87817e795317f608481
zd98bbca58da35919507799e83a80b0910307f807335cb85b3805330de3bae0f4672d49e87fefb5
z31656b40b5603a212d69cb0f348691806e7f6153fc4374bb1f9db7554ef3eeb0c120e7976702ba
ze1d17c9b81f9bf4a23b1157e76ddb08575e4bf0798f28c4d5a837cf9b28206e1b359fc1f155568
z3f48ce4ad14c474ea0047a3f5e601836be5e08a6855826c1a3797d916747ed7e5838f7c0d44102
zd8f1ab2a982c234221d092f2646fc880123cb97f50c951f5f1c48252607c836834da20478345a5
zb7d046b88178d3c26f6ec8101ad7e8fe5f8a02ba249c2fbb23f4c35dbaa53e1c2f9d2df3c1752c
z9d4c4599352b85bc3572899a6c2028c7a5c2a0826ec03850aa71adf9ffb05fc42b23050b61bb7e
z102d309d2f05a90d0a6243b627f7462f5dc82bcaa997bf76929ae159e923daf41b9fb0c0dbf6fc
z29ce6c36bfbf9b45b97fbeca8803dad31ffcee42e2bb65688e53a1d7d85ae77536c5a054515fda
z69f491de9177756abf750b050e284573ca3b24cad9d0686bff93dbee628526ae96cd1b2e37ebc4
z1738c813f8dc7245c136834980a189de0cbb61a13df2da490e2dae21192c3de730a7f51c37e701
z69fb2b1aaa0003382e3a4872b66de139146949d6214b9c945dd4a24c0739f350f78b6d2c41c2a4
zc911bf710a7a46d8bdb56d7ca3f3790579b383d2cdbba045c7dcf613a945a6a41b5323cbe2ad9a
z215b168f2f8f756ab41a9f09c3322c857887395637322c66d7e0a67b24ba47a0a2f32c790dba4f
z55b6d19e4e00b49d47101e5407937ae25bce25a609b843809e8f8f667adcc7cc9b75cff91f9701
z154edfbb07d1b7e1da0734e0c259293deac098257e2d1de0ca6d93ba80e0c79594a276d08ceb2f
z0db47c9272dee25ca8be58504dc369ae8ec38196dcfcba93d0600a7fe82a48cd6362c6d57d1139
z54bd084fb1c1f8f9a1b11bb421113ed07343bad8d7aa8cdfc221bf13615d57af8ca606febd1e11
ze28562cfe4ecd7018c9c8683e2c4074d39ac87043dae57aad2e4313a39233628368c1c6f5564b6
z441e9a04aeb7ad43b99946edb0a888700bceb19c901e72a5e2c05e2f409868575a99d21418f1e5
z098da96429cd570e4758e58af727be2a6efd6012f731cf0027ea100478139543baf85ffa80e206
zca2cd7587ef3ba5209d92b8c0e76b17c5eb06c730ebd4ffa4f7de8cc82a983d7c3ca569985beaa
za787a6be62593d8bc8a08862f5b44077eb7b15e3348bbdbd57c09a9a485cc8feabb40fe106f203
z1cc32a77bdabe9422510774343456104189f50a73445c80c35b76c510224f05fea13f36f20bd9b
z6ee2cfe786d5a2e9bf64316eba1b13ed1d0253d87294b16567d1c2719b46b1a6ca5f7640ae540b
z0b68276f28c6cda95dcc1969a8ab80ba6bd8a32c77a3eeed3afdcacac413420fb9fa7dbec0aa71
z5bc2fed53836793fad631408037478de937349897f870b348f37e1d272e7a57eabefabbe6427de
z1f96aa747cfacc5997e3e9c220a7d3484e3a06eb8e8ae434b0de8fe8ad929e4ad0e9ea51cc35d6
z30dbf12efe8f94be9c70e2eaaa6a09c90cda57dc53b3c319ac37f81d7ba7532c24db17f52cf712
zd001d82852c3d692778032fd31fe4013a4d485838d8e96fdbe8d882f8338d71754d6b170eed487
z9450814b5f2cdcdff58f76154193ed770147eaa3cd21e74ba01da244b5924906858c100e08c799
z88b35a9ee0e6ca9471d1c1ba6eb401a93ec7b54ba3593bca5029a049b8afd601b8df3c16fc3769
zb6639f35766a59b30110c4c9237278574a49b4d5613eac576c36d742abbc69dd7468ca5d5e288e
z76926a7dc4cfdcbdb131570627e7916ea4449c0b5c74382d38bf218d90f1b6ccf9fb7ec6de9cc7
z7caf8c5ea025fc80e75a4046deab44adaddabb3199260c5c38a9f52e07d05159920ed9e21f3bd8
zfb4d773ee4c991c147f5e6101e68b4d348782c92cf96cda90c35dc9d3e119d90ab4fb8aabe8779
z5403ea1f21b97e64bee18c3d0fa6e0cbd889f61670e2dcd777eb8e0aaaa61233b36c95b12f63c5
zb75becdfa12fbd4b811b582ec8045260290bef7c88604dce164a1cc646e76f5f55e98fcff3e9c1
z7e15e547162c79eaa5a2bf4f203b3bd1d124610caaad21f31f7f619b66ed35c8ccbdf1db8923e5
zbfa0363e644e27627cb5b80b1a1472bba35aa06d477ab641c8a07c5013550267306e4e54ad0790
z81b2febd6fd9af2bb36d4d94e1454e266911aa1f4185718cd729f69d80ef1c6c67c03404dba5a8
z56fa2c30dd6d98daaf7141515aff8d4574490e148f3e407bf221168fb1dcd09f9e8afc1e621eb5
z2034785b13db44b56894b1e701e369a32e7a6a278f0f7e65aeac6dc9f96b5eb945c6123860429c
zbb2939df4216796a6fb3925e128faebddcc01fbf1ae9ddd6d7d60d7989aae353697051f3fc1e5e
z677630c7e1c1fce8872384b1a9d81acebe4b3ee9ff2d7c46c48b855f2610457cd611ea803860d8
z21f5e5b3749767fb7815d7d387054dfe3c25322ca422156f90f35bdec8655a8f5b44ddc2103824
z97b5700adbffe24115863466c24e5af4764627e6fdf9e65d9456f13e3dad2080486671dd1e683a
zc94355641a339cca29110a5f177892f4fae2da2fa08607b009a8081cb2f3eba93e2ccce25453f4
z7fff72613d99015bf8bc11a6f45621e80cd158258b24a13b250e6e93ca06a6eedffa2e90109250
z202729eef7a11f57396fe52c86166965be958eed64858edaa443a64bb3d04e62753ccbd87aecaf
zb5d6ce8b045f9fc04cb4f0e7cf31790de5ec6df72d4e66045b90bd74b197716f19669f74f94399
z8a81308026a80d06dda448ec1bdf07e115857a01a888d236c488e16e3fded6a26227b2a73efce9
zea4ee9023490223d11e2775b04ce6e15c84cd2c829c1f8adb9d89678996f8cb7c5a1118c461e9c
z157050e2e87515354f7a3f7b1b35c384d3c07be3b5fec2c4482390a65abce10829e79a55b7bf0f
ze073d49973c17039276a9ad67acf37ea0ff7e33a514f9746a45d905d89e5e9d5aeb0a688c558a3
z8e6b1951f79b94ff180b7e404ba733cbe2d95c7c212fbb50cc821e093f01ba1bc26f3a5d802293
zabdc565b784a87350e0d7a3743aa27c523d9a9f33c0f08466e613a35fefb30cd97d04009a0ca14
zfd8c176239ae5c57f5c269c9fe8065a78de9b288a2ad3c75ee0e056e9084dbcff17f0bf65bb15e
z150ddcf652a1032c92410415b01a29c9e506d55a6cdfd016bb101f7191855d1bf8b5192c4b2cde
ze4359232a22e9e657f64faa86c1f37c2d46841c5c9877f428a7319748e02b20b529544785dbf44
ze11fc07620de8d8f5a2276604f2f544c08a89c0fb481351f2def85895174aa1c418aa5e2a64ac4
zb9eddbd74e337ad46904409a010767a782c1c572e8b439eed6219bd009e650015ff9f44ee581c3
z67c69f381ddfdf4dde26cab2c9831b8b9b6b8ff2c8a874b3be77c08cf7ee156c66cd24c38adc22
ze05fd21bf415288216cbeb872ba83310ab1f00e9b06d0314e73ab5ce302851d726e864a39d1ae9
zcdb595f1f460b030c00719be24e57d239451ed37771aa8b89dfadb7abb620844b94df2ce32caa9
z0855e5dd1aee8fcc655a7fb4652d163470cbd284db20e4f7f466a6abd3e6cc59f3c16503838ebd
za4edf01cf600f4e64afac9a4ebd20f854a7c9ff61015be6eb310324ec33e22db0f56255bdbcb98
zee0dd6fd097698ce747cdd8e843337961a034947cdef654b5d196e3629400e12ec97dcfe76a5a3
zdf9398c312bf593bebc72d4bb57fcfd113fcacbfeee98cadf69259fd99449e793ecba86332eae9
z20c12a3cdaa97bf22ac29729d0b39b9ec55ecfab2c0dfc89cc68d303a95bd88ead0711e1a0fd39
z7786609235898b3266048518915ace3f83e7afe7cc927c739eb0dcf8ee075611cd146857db46bc
ze512d1d6c0126246b0a39bc8dd21c6769915e1e6918f5a805ee809bae23c05270fb12fb33c05c7
z3e4d7b960ae2aceed32e5b1c6c2eeccc416385f074fa49fcac5addfc0f3acad4fc15d8553726c1
z8c244b80ef5b5db64fe363fe5b87bcec9729a15a9e8f892cc51d04d664e4d4f17ec09c245a686c
z0c46d418fc5be3317f797229f737cd54929bc8ec9a2f273c64bec589af5def250696bbd23d5b2a
zdf6a16f6e7349b8ded8496ad69b2a6d4585faca36839ed0ff8e798b36d9ee9d0098829e7ea1733
z340ea7f8d151cfc822431821fdf5f0a478de9f5e05d10b1e8e772094ab42d735315fab8c767a59
z1b16773ee9f596813a58baf044a96ea4e88939d2c47d4bc40d337f7a568feb18e8d19bb51b9069
z3e5822f435d3b66bcd9c6b33a9500100f4083d4a67ee4db419cc3787523c9287b03868f1f7bf59
z6e77dd73174d37ea77fb311826981f1f938a8c230772148a8eeff4f35898f029b303f806858232
zf8d54b78aa030e10f12da6e7b1bfc59e4b888adfb8eb51de445a463cedaef0a1c1a3c464f359c5
z1342ace160a5f17d84090a6e879cf325aa52321a3bd049571d2b4ecf7e4981dd6a6e0fc24cd466
z054b65a61f62206520fb7a48ca7e4f026733da02e22c4928b951e9fc5eed250c8ac378843e3702
zde50f6af0e20ed09c79e70041934edad6e27467a53860917c375d6925952d2c4ae3e3b42d776e8
z93f064ccf0b78c45748deabf5e9d0634ae9b28b0ffec06f611c03a5d9c7d79793586716b6ce538
z67e0dcbb942a11b65408d390c39cfbbe9c70d89173ba2409e1bfcba7940c3eabca4964a20c8b9c
za60391c97621547961c2c7e288665d9596f9c8674e2715e744631d26b9d153fb5ad80d8d7d345a
z48adae7d869e7d98f041d7b526fe42cd31313a0e880431e9d16bc52ebbc1002f2b1a8ee3414eae
z8f88a374163902d29f6b49943d1321e4a8c5bb847ad56c713eccdf3bf9ddff7a261a24b82687d7
z14cb4e9b6536f986ebbd62cbdf74a4b813f4a4bce49c69c33ce4321ef648fb54d298bd43c6bf04
zb8bf10f4ce6e69d386e847414cda8517ef79232bfde085e5db3b7bf46261156640163412912e94
z28ff2cc8b929b390a451993ebfd75f172b6376caf22d68307e002aca666b77e2ceacd8eef77829
zfda8c150bb57ae03ef1620cfb85909a463af9b99b99c20154a14bf2e58937a01f7bf8c4b402f31
zd0f5976d338ac07243ac69b41485f0194166770edaa53c4212344cf56d491993bebf7c750d59a8
zf6828160354a0d750919a77283027fa7af5abb353c1f7061b8bac1b3d0e2d2768ba87e80c66a14
zda6b88ff581c26d11efed947eb008a377ae35b94da3ec43872449963ce059d0a980483dfe25795
z069a8f433c0eb89284eda689f9c2d58a96dc6829b85c33b92e6addc215977f95ccfaf95b43ec5c
z08bc68ea0ee8e79a279d69317f1f3b344f098e9cf979453350155e41c61320af979bf308cd67dc
z56089e0ee9e72b506d3e7b08baa485d833927b62dfccfe74a7a23e821dc2fae223327f1a13a2cb
zd0270958dc319a26e47f834d6d8a18588a552081e9482c5f4d6609a8b8294e474563ba917ec0ef
zfc7a565e8ca2356c355b81eb265c2da026ade01ebfc05530bad8dbc69334ebd2a9e1fd1e068fa5
zc06e54e626c112745f06a834e1620fe23d13e6263b550fd07f1a89cfb259e319f835bcf8ddb2a6
z98e4727b46579c320774e2985aa596527609d00a4fbd5bc98282b40e79023ccac5f008c7a24345
z05373a24d7e5f372b24ddaf29631332bae639b79bae063a5fdee71e4bd6bf73354b8ea5b3eb1ad
z03fc7eb0c968216c34c3a26c687a5a30c326811d0dc7d3a9cc63d6454eb5f0ba9b23dd275cd860
zc83084b55f4a2d7f2dcab27d762e567460808351e4c88f84a15d6e3d73fbf12d060571b2547d6b
ze8bc2193574a96669768e7492dfbab327aff9a48e18e7da051e8ef51d667d703c823af7f136115
z0d7379990515771f4a5441c4c28d61b747f2757d5847244947d33c17cb2dbf695133c8e08e875b
zcae2c2fd049435bdc17730059cb905e07d0c9c286ce261a9142308efa3a96f88a4770b04d2016e
zb14cadddcb7c739a8ce59165cec0329f6af5d68b760f67bfb5a9dc68fa117eb72e2351b21a12ec
zec7e002786b9a6fe8fa81c366eebb8a0bfae1aec14bcb4806d1fb0becbbff0bff20b8286dfb88b
z38a1848457a4a049e0c5cf746b9e145f5d739f76b06f3c63138478db3d6bd7d4ae8a7ba37b905c
zbd07b5f8ac775f5e23621db36173ea2cd0731f80a125b0c1b4ac29b76caff4e5623a056f243c59
zbeec9f7155c15311fd03ed262082b1c1bd0888b8615b682ac686c6e05dc4529a5ae41c17dc0842
zd13460cbd6aa654b5b415e7e22152309f4312a3cfce0d8e8037b28d90dbae9fbf68d245a1cadbb
z2a79bb1e74055701f163f948ffd2ac7f811ee12df1ed2504e2f6f0e5e835932ca203e53bc471e5
zd581bb22770dd342544c84d271ef7e8cf78597b4c5ca04588a6957047d178dcf13a04871ee4813
zab54c10c8e867798212d10f248082ab024cee87dc5711fe726a25be5f64d7cef015d91b123842b
za518e7f65902bc832a04380d9f9e66c25dd59f0da6d9a7cd12271a3f155a51a84005e7eb368f67
z4f51798320b5687e240df9a00e4a6ff303e55aa371222febdbac3c4545cbed9c2b3768edf9f8c5
z84c6cb4d7d8b3f25edfc3c1440f681298f8ab1be75528171f25f2edda563036364ec93db3b3a89
z30efae5aaa7221899ffb0d2d10c31d7f60618dc373650a30c8124e5bae26e3b5a566d5087cb172
zb813f0edbfd6e42151f7bf1cdc3e4d0f3df2e197aa69c157cafdf117bcbd7a4dc70ae614a3432f
zc2633ffbcc4498feda8d5115a68500f3cc63503689dc18455520d0af2303f42daadf451ec135d7
za9ac83faea11847e8f98c5531c9eca766ac6ff4724edd60423e8838e31cc855c61a0b16f55fecd
zbf1a3dd11defe0dfebcbd888feac4e22a05fba40e59fa6f9c205e66d6f4e569fae4077785f2974
z61b80c6eed6638216c13127c2e1736b6226ba62f294db5abb58284b86c7fb1e16d0a9f4d9a471c
z4844441011cdfe683d2b4353f2d44c7678d12c42d6bdd3f80cf1754bf6211b59f721145de84002
z22ea972a534d5b3cf3b7572a5007d9f1fb753f08d20e424eb2cd68e8bac7dd3f2334195ca12c39
z2ba513f81f0685c3db5bdb6a055559c36b4d6ff65c5041cec984a058ddbe95d267ea93dd89810a
z1828cee9549154f4830b6d6521e5e3ef965bb4e85e93cd563d4f542b6b980a85ae2573ef768e8d
zfcc255ecd06f540c7d7ca6b068ae67a843ac421601a8de1d1137fee80e73809b6545d1bfa2b972
zcf319addd3cdccfebd629e58f904b2576e29c66b0af02fa971f47b791646921d742f0ef2d11204
zf0ddecc77e90816e10c8989f8a0ea8ce79e9d74fbdc2be117d416bb81a37fe316db6b876fffa18
z5c83c9fbe3bf1dc6dcd69d154717dae0b138d76b132dd2cc4c283c731323978baa20c996f72fe6
z9ac987390955f0e02f70c0d5e1e0291396a2755d115a650ec6270dc325d36043ac84fb1af0a669
z18f066fda4a85a1a406edccbd993d2938d9957a2b222ffa0f760154f02df92e38da5f0aa04fa8a
zbde704be2fba3b101fa720d35a13f1486febde79bc2dfd1d10d4f9f07c20d38ff42b366d8993f9
z605c3f4ab65ed7ce8952658e9dfcff241e8b311aa9e005e24b230e4f203f2e27bd3db0636d169f
z400bf25ba5f50799729a06bd8e18859410a697f44fd2238d4e4a4d83503344da87f79febf22d03
zb4d521e3c4aa637fea70229db3ae7d8c94e22f5e821bc44b9d8769e2afa3fba070190b6ca5f094
z94cb32469d3b44e81342e21fa0d32fd59c21b6e125e42d73c4963e07be4226ea2b178aa76cfe72
z789d2fa40a7d265421bd1a1b48561ebba4f33fd8c325d13f5693f9c470669c92569618dd0eca64
z892f48ba65a746b3239aa505ff3eedf7bf7d7fc8ff85c4fefd5807dbc09d60d3eaa86dd2f37c17
z5e97f035897f77d6b83c408958dbc146c6412729f89617951d68532072a57f97bc9594eb324613
z25de18ef56b84005d8a35a298398875011d50f845fad21baef5d513c56bf8253335aa077a353fa
z8b8855941ef544c1f8f143a98396913e46ab204e6f7e58dcf0fc53494d48d7b6876e53bc9ea191
zbc4c1f1a8a81de214c270ac0ffa9c375cb36b3f02655f0ddccc328b6c9b22e10d0fc8c088f0401
zf8c112ca8608e402c1d23c6aac9b85354ab47d181ae389daff7cf5fae108d94c252a25c90d82fc
z687533121af69a7ecd620a856268d08b01cd94f10bd49049b95308d87f21774692b7312bd843bf
z66ddc690057ae42c83491637d627cae656ef1bd2e29afb30a21596ec65f43452bac108da585354
ze0a96c40486873c816e938eee3098b4467d10330c6ca15fe01f11e5d4fa1cace55d41b67a07e86
z66e9f2061a978135106683f8d791227b9724b8abf7b0f4e77a8a9fba21fc7d01a06aaaca3040e3
z90eaec7af93b5caeede7292136336a1440ae13afc6e8f84f70ee76839677189c5bc927f1db7d20
z5680fef484bd2a0fbbbf01017f2f00221cf69c9a341e12f621b7f6cef89c7a95b6b27155e16f3b
z221cd59b9709d74b1cc72019c2fb035c0b01292cf0ae604b965846213f61fbb23d6f9b6aa1d788
z1368eb8b916e4a787692162d95ba72fe89c9101284d1afd57d17eb3033d1a556da5179fd1fec71
z63cf8a7e8b880967eca6a08475946198c1e17294e28d9c36533d9fd40285550cf4a7ed874f0409
z5df3be414849718c8ae595fa698e562d5b60b438aeacd486b45dc1ba32457993a7e1bc439613ed
z07bdbc04eef11152376801ce3dce1f36c2d49c6165c55890a151d671f7d27cedf4e8aa6f3a630e
zb437dd1cc9a409be09055add2ba97935299ec6c41104223fc0063e1a7642fbfe404bb7803617de
z1db0d4742600d31faf2601ba29d346ad6202e78a453506ffa5c32c00a6dd89cbdc39e7445001e5
z71586c67a9c6de66a59edea98f88c73d6230abc685b30847d8422869c1c728f91f69bc41ff7329
z8260063539ab7e4083a936846b0fdd6def65067c2d15b6b2e9502d5380c8816f23a87eb238e100
z666aca484389d8eb2400486101f56f0e517d4291a130a18eb94f55ddb6ccfbf3ab0eeda44af869
zd0a12d3ae57ba717971d36112aa79645dbd4446937e40b02133e2a0e0ad033fa1807a060210215
zb00c44ec3ab2ba333fa336960ad39cf98dc049d43af6e4c6564ab9ad30dae5663c38e88f511bb9
zb02a7b46af5bbed3988a4e7f4a9ff9c324dad28fe5215ada5d00bfad475fc161b1312789a9bf0f
z71fb6e4e864e9c2fac10fb8774d9146e5bae8b7709da893d8fad3938accfbd72feaf3ffd9f89fd
z18e5d7cbff363676c9b4b374f51391c7733792f7ad836b46cd78b073a373f379efd2472b1b21c9
zb204a245ceebaf4ea3f27dfe3320bf304ca221b52ddbc7e958e4fac3433d194cdbaf61ccd9c155
z77531abeba11a1f7f0f242e696caf4180bdae954bd2e288cfeadea09c7d907f2171551920d8663
z11a618c49ba27e316132a9b84beda61b3f46a8e1bf5b8068b2f5ad424ba2203be65f804f09e88e
z8abaee078d9e09c836cbc416273f78bc9bb03c4f6a78005334b54b931c8dd3f3039e1e96e2a870
z42aec3000f8f1f1f48bed08d56c8f2afd7c98b24387ce9d68c1a6d7de126ec21f0e1861ae6f4cb
z04b53a80cce613df85887f54665d3abe6c8b12ed008c16a1bfab1ca5c8f9c0db96eb54dd1be6b5
z598bc07ba90be66e933fdf2833b1a3bd50bc14d733a8ec13a0e524efee4302601182f143274c12
z955194de4d171460b65b1ee433c1ad63709904d464e483f920ceb53c5676d282b7e89e11f67b9a
zf1484cc52a5394df751ee8198c0f5d0f716c6785912c107c45b7956865e4ca6fe6343de983ecbd
ze1cebc4cc59ba48d66bc1b66f341b732314172994322ed2877789be59de1310d788241df64fc10
zc8c0e0f7eb888f8731e9fa188c8ca236e3d10fa6bc5b788099ffbfb1f72e54169fd2a1d54baf11
z648bf73fb365281b5d6840cf257f9bc9597e90a0ab9f62c34808025dd88ce56c7e5db622dcc1bb
zfd7d5b585e02722cd5518ecb7ebe0668225f2896b0f6326d2619185d178b7062799b508791cee8
zec6194a3795ee42df2f0f93c54b42fd899a13d71ad51c54d974005fba38f8fce70b911eb8ab17d
za24250275f793bbffe07a2fd1d75debfae0d4b98100e7cfd0c3a78b875edebcf3e6e4321be35f9
z6d3771775e27b7df41afd95e8ff967c823ad3d25ec21e118a76a0292578a111da1549826b6bf37
z36885e87ffe48504faa2d673c3bce9af8f393826799cfd2e59f73d0e063ecca626aff0c71f54f0
z848dc483dca677c8a425b38627b9db994069ff707326a0861c458664895b0d49b446226afd4ed8
z25704783f4f9dad1598bfd21abf2b56926607bd06497b4eab73534b19efb9ba13a6608c32c07c1
zd7123fc22315309717f091ae306e7c24af641523c7cb69821f5460fb6816a0d4aa4080b0cd83da
ze50ab575182952d2ac753636ce31431f4d2b15b93050c9cbb398240113789d314fe71030e7add7
zc7c26bf9cfadd576e4a8f156da9eabd2b7bc97ddfd945c802bed564477755c6d26cd20daaacd9b
z1d43b3cc6ca07e28a0f0ceea9e2d10a3ec3f312a393d2d3be3c1008a3922d35b1e57c5dc05f178
zfe731b267064d837a684ae2c97f5822286795c0cca07bcfdb88b87a601827980190ff98ddb2626
z1b09ac66f7a42ff52751f97fe9354115498483e387c87db73f883b0ee628323111ec63d16673db
z6e8f03001a87208fd0188b92c0be3bc220192c704f231fe875b21c8cf9755bdcb0393bb8618568
zbae75bee31ece261f0fc28a149b928c22668d8ea51114518600bb5970eb6eb16ecccfcafddff7e
z6cd43da5da8ed2d280a9909fc8b49ea16f213690dbd57bbdfa8b37fad254ab87d912e2dc8c1b51
z560382b0b767f663c27445e01cc1cbe8d50aed97466e805e001b436fe423b21a3171df3953aa30
ze01d8574d3463e4aff40e4dee0ae98612b921e8fc782e5813d4f65bcff7f037f65a19ca9f132aa
z192e020093476be7ef2366144ba1a168e893ef4adebb6cd1401d63cd8983696a48b31c2b4b7969
z8accb7fad1193247befee454a96508a04e2ed1a510add65b02ae4bce1ea8d6b3083c64b984365e
z68fcba48bc5aa45dba3bc0cb82d6c24a280077fd5839053a0aca5f58997c65d02c7df1f074f49f
zb7908d53e161267f4461d0e4b3b3e248a06b2891aec1edd46fde35333f906bc9eaada20883f3a2
z5bbdf20d1910f6954ca3a6e79965d72f41f8bc666574006f40d6080809571a7dbc3641f0c19cb9
ze9f946d5b9c59490be98cd81863c2bfc23c4b7312361ad893bb2973a0d8ef414af1f4cf71fe309
z80f2e85d3b059cd7e5ab89f5a7ae3d10c9e1fe0b7d4193494072ef09d9d9dade39ec5b5f374545
z2b5c32638764f4259bed2547746810c42fca48055e10bc5fbd3095837b6292b1cad6d0c707a3e7
zf273a7e365e86a41695de161e6939682487f91944dfb135ebf3b47248ab428c808e515216592b2
z7f1cb7717945f94f7b3d80002638e57ae2477ea5efbd5dc35b557cebeb4d0d4cf795c0ba9b2a70
za47ce4f2a0fc31d780eef9f1afac3f7f48992f6e17a71c07ebd9e8aea0404eb844451c0a328f24
zd1e59d27665e2918269846d6b8b1c1d5d32ed77ce4ae13663de90b345e27184e77c5014dba7960
z617d51dd4ae1472e2fb1db37184ba7cd4c8349962de6858f2097d93a051d5dcdd31f79aa6d0cac
z1e204008e56f167f4f634d4b45a0ffbdb26604e96b2ea050116953efe0f687f0095e31a31fdad7
z66f6e398570c759a8b205367e24f3550a9e198cd02fb5ab74740953289c5ae0b9e52f1678f67ce
z3bc8faffd7d68131308e0a9426795d404d0d5e8737e029556ec91c6ee3266f25b1ea9910c6ddd6
z4404965cb3f03dc36191304b8fef30618584b64d869d5a9e42bc5be21d9ab7d2c4642ad4da21a5
z06fe52fe5a3dade23a7e30898bb2b6c98905378526af9fb5db5abf9a1e93d017e917602609efff
z9aa8de5a642510cf4ccf92a65b22bd486547f544d75f7c33673a63effc17f02212826d4fc2b176
ze34b1ab2f67c024dbf3fc21983014e97b54a7410debcc82c759de7d283349fe193999ddbe17c1a
z4634b28f1fd7b686e9bb7249fcda8030da12ad931b688e52148ebe26481ddfa5677eca45913c11
z9b8c9ba461d5b04d614992788d32cb2eb5746e352497a7b982105c5cb975bbb805d8df7cff96b6
z8c4a354ae07beac1066158a7295fabab534af1692eb02e8f189b51a2a6783a12ce362a8314dab8
z756911fd0665d94ab830a571efb729c5eb7e935fa132abead57a169d98513b5a887c11f2d98806
z7d2f41a1709b8122013cc20fcc0af42ff1d80c71b3a8b4677e49560ea4f46b1f11a386c36b6a9d
zad7bc094a7882d56554a64ca413054fae5cd9cf409b239e67a59f872cb7bdb282e0202042bac91
zda5f324711a29e5fced24b6f7326aeba3b2b586ddeb0f881a72765028a9b7fef2a4edc4580613f
ze3c414df24272381c3560aac899aa9539dd6a23bd3a590411687479cba6defb00646eac9a4b9eb
zb75beda48f85deacdcbefd75f65a5ef23d3ac0db90c455fdba154550373236694d240e5d07e902
zdc714624721fdabe175940102bb66e2ccc44c52ef1c1d32214ec350c6c48c01e6d9ef88bb045c4
z5df080093698b83f18c1fbca93b1bb0fac59a628a7797b8effa6bd360994d41d9e7dc80839f874
z4f2e03e894ba1a919b6aa0e2b42dc6afcc0eaedc1d07a6c3383ced4b1737becb8d3bf1b0c0da2d
z1660716d0de5f826735f39ffb9daa6313f8a93f44faf4d6da0045643a9eb527774454e45ba1f59
zdfd637c4bff0b33a21c3472aca5ea96c6879548afae1faf5d9b1dd8a5cf4317328f9f602ca4c51
z3b4f28c8be40ca0308e33936719d65cc37c71eb56af9fbfa7151d64f9bed71a30b119f977e3f31
z2696546fed0dfe351c39b6a0ed8c235ffafdc8bae2eeb7536096b14e04afe377f17d5b0b06b25d
za8f612c485afeb4a401191de680ad2c6d552ceef992ee9aafa971941f2f886a3231656533ed7b0
z9225c709c75a9f065ad52d407117f6f55be9f814d440c630917e860a20998e414fd3d863e58af4
z551ca457548ee84c74ac6741b1d6bb71682b1c21f2305629f919c9782f93303d48dcdd71e58cf7
z14fc6680e7aafda39e59e69b1f080e2e2c34326f31845ab379ec8c0641591b6b0072b678538280
z310f32894a8b8e3491a706772509e2615ea71f55c9acac5f956212b7a3edca5bb4926f0c105daa
z33c048a59fb21053effef5710f0c059015b46e4da40c0366817ef25c0889b89040ac34af7a4cd8
z1a2b024baacdc70c7e5b8cc0d9ad65db01883dd3daacbed6a06b47ba6519df468dfa3844c27cfd
z2dc0c762e54b6df5d9bedb09f96bb9d9d06a19314ca343e964bf18c094a1b1c62e3ccccdbccd09
z1ca4ae4bc41b14efe1db53cf03a157153ba09cafae0aa72de5edb33867b5c7e6ae352ec954ec41
z64ef4c3fc8e44c92989092eddc4507cc386ed924f929fbbba1c115ac116799df88dd9f8ba3fb78
z17378456b1fbf7eadbd33ae1fcd8921a5928d4af6796a9a9935d52ad6ce782a47e69aa4291c984
z90805fd3c295ac252923f0344e419b345a660892b8121ea4d8e5b896a01109590a2d06e7d2d3be
zf586a3646b5e8d673bbb2a53203d1f434ba0211d02b8c4ddd71ea45ba9efcd956d7a3fd0cfbaaf
zf8b1672f7a8c14a8abbfb94cacdaad0ff5a562ec8d6b27dfcbc3d3c22df657e234035676533b7b
z1ecc87ee345a38a2e41423d549afc55f86c69e2cdec616dd429fa60ba01e9447809c822426d690
z7c6920c94288a07cb70cd12ae90cd64ede527ca245fea61ad0ba085af5ea08e757ab241a56a36d
za2a35eb4cdef821c265bb0711588f8bdfdc08478582afda9972b4c381872b34f3acb8bfd4f6560
zfeb3cf581c93c24ba12b7fb958e3112cc22423154af09b70d9c2708c8494af6dfae37fe18fa80f
z3d22285deaf73f96c280822eda8e7507409c65117a3ac88323b7d1822cc0a629245d4bd574d255
z9752ca958ae4a0a0be2cf8ee9544ae04486582c1b1fbce73a88538e332dfb8cf2faa7630c8716b
zbafb5fa784167c4bdba0568183ed7decdb8be1da1ae8f2ff125d7317e250de0b3113ec67512532
z34bbbf91e12736bdfabbb9b6e00bac616bb1b99a4db5d76bd87868dce9434a929fc2007eb20ce7
z5ee4f5720ebaa22863f64c08a8dc44c48944629e07b30007e2fbc6ce8aaf12303ff33cd178bc36
z3a012cf7e789522816d96633232a1f3b798ac08a866f3952930c1096a8a9326cb89885caf9772c
z535351cf04e87c60ea4076e1fdf6ceaae12b242bdff7e87bf88f6314fbaf48d95038afba9ba918
zffeb7ad8ebd35c99ad16361c65f3016e5875eec3c6291040772073dcf667e1e7c902771e33d5b2
zdef40c8a3be5229bfd57c6accaae2a7eb57cf54da47180134c83d57ef9c646ab701e7ae25cc8e5
zf9c7478307a21dd421d148223943b338a81e39d4111e95f9e3a3f1d0cd46657d206eb89eea89a5
z8489b689cd0398c1fd0c5e0d714a872dc3196e9f24e705e538ecbfc7a24dab0c10552c58c92844
z83d8faccdba26d53d6a72deb056b816dd634c258932a904c7b7d7d13aba38a667210ff5a357be9
z38441741fe73a8026ad1b72c8ddf4ca415a4b4d1933694b56f0503c2dfbed5657513de4a7ca742
z0e89e24ded6ead5d334fb67d32014fd28db79985581fae2028a3092319b61ad093ccd649471012
z60387ab0c91ea208bec0a19efddea735d2e01fd3db446240a96e64cc8d612b45b33f588572a520
z628621210f0164063c6a2b753daaeabef699ace0f01649aebd35a9f9a72fb8809359e71d6aeae9
z44e4a04cd37bf167123e3e7b569e541519c67376b2a0636dbf450ae4f45b91582abadf9c6b7dbf
z1f8c239880130e65a88f903fc0751cfade16a8c1da66fe5e8f808366f26f4430b91162d23da02e
za2cd73fd23bf0c8a1cf3a8460298471a8eebeecf37d4c55f01c118e3fc4a45e60380fa8c7bee36
z77545fe0c2d8d7ba4548f31439f9a7b105f5b1a012d5979a9452b797cf0ab48513e006672ad78f
z3e945855b68625cc1cf274ed724894e9ad4b86f54a7cb2a9fb98d5fc8f56ad2912b14f441fd4e9
z9d8abc4a1b5f3ed9e79a18169c235758f87bf4b9a6f6f2fa94bcb623547a6f85a80c8a3da24e83
z95544496c1011a4657f9f106a7ba1ee29070908238b801b690f256feee0c10c278f16f89ce370e
z4aa0e865089a016fd930a214efb774075f50ad2fd320096a62e11026239cb8fdbea90494cb4c53
z469ce46b789e91f04c3f0ac1c7ad407c322e10ae69ff45cb405dd220059d1b888c7b6f9338f157
z53994195696ab87f6e519a5456e5fa2f12f95b120b85df1fc000b2834033158f8a353884387c35
z4fd9e1847052d9c16b150ae59860eca7bde287cf077836d525500888328cf3e1f5f93d4b742f66
z08f8484b8559019d27cba3ed0f110853da93cad052e468e123179082472fd670adf902f272820c
zc50dd690808af1c457634fb8f386698a20bed242c1c2fe5887a75d33925e122bbdd60151412128
z0be1076cadb60fad3f50579d768b9a179088c999ebf11b954337ddf54a3f63e3098bb1ce584aaa
zfe93ee502ad1b4d46ed9bccc702400061e3e6e8b701d9b41dafd477fe143d29bad44fc4656f369
z0e3d2e379a1366f22ad60922cba76200323c6c8d0d7410c57f36b5ca8d0f57bd9749d48b6da28d
z4ad9a4ebb52a9abf47062bc4600909989625208ffa495ae176bf7709eae93022011c5ad05c928e
zb5f0632d5d4d120e97a04e971e8d19d253b8f70dabcaaa88bbfd9e792d486fc8c1ea702cfad7d5
zfa4a10aa0aa07366ceec6f00fa531e730337fbd23d165bf0979b0ee8b428fc3e7554e0376835e3
z93b7754df6e0c73d4e41e4cfcf51dac8b49990c4f086f628f256863feb38959a1ee92aea2d3673
zb1f4f11db027e8bc28b4ba4cdcd6c3c4a0f4e243dc22d3cbe694e68b5feb560b2b1f652449a1b4
z72423bbda1eb9c16df7e342a14c69e3bdac8112fd8ced12651779d7415113372af88d4e11b85a1
z3f8c03ed065ddc34b347225b869dc4064e9cae8728d8f7fbcba77c463c7dd91bdc626fb4f0d5af
zc935881d78cba47594d3421d3c77d04e8336f30c35717f90a12866d0756e43c8db104e68a66a22
z994e3c8fb6967dab2778dd2d4cfe45172a3d9dcd23a298993186ae7a18e687b68bd53ace98b4ce
z982529687f2e35d42f09449f83c3666438e8e1134d4eb1654852663dd155e3f24c07cab7c9c3af
z55231a05d7bc8551ed4aa273ee54a33b3e9f65b4862de4fb6d97906c816c5098942b680a0465f7
z5154289c49a39b38fa01a6b5ae49edc8712062ef4ef39decbf135ee1c3dac60f3ae61e0132a408
zc05e1ae935e584f007c09639309a4d9c10e2df66aec7b6868ab4a2655f2fcffce9053be242dc29
z2377360a0e6806d61b087d89615ed52e55b313cb820d74926f63cbe21695f1df8a89de3f5a3b8f
z31ff671ff92fcace664ba36bbbfbc29eb11e46c5925a81b59f7ed6bc14734a2bc3bfd0311dff7d
zffa06064f820da3b9f449a4165603a9c73d05728ee958d85658aac39321efef62ccc639333b765
z72e3efb5b25e3601ef7d87bd9d033dc4d23783a466a22c956f4b141a102328354892d8dcef3813
z25990dce07ccc07ffff43b30a23c75674e1ff40e66aed0edafd59e649014a00da4beaa8d2d1de8
z5d5110f2681a2efac6fef69384bd8ca63c5f24eea8c5ee797d6bf1eeec3e32bbb637118d857da3
zd2ddc58dea8170952b232c06abb36145912ef887296fdf98d7065438f67f5179e433beb72a1d58
zb48675bb32741775cbb98fe5fbaec402f02068064f91722afe15a96da7ac20a95fc2d7d71fd70e
z48c4f0735dddae96d3802bceef587b59a5b1bbd5218af050108df56a8d6d6bb7c69314ff53d571
zb7b027a424bb5fa16aad9c33c6e07bbf071fc0c5834a023a7b1015bfc9473dcc9eb1f6a8016745
za6a06ab46125a3ea50c11c7bcd8fc4c733d86e8ed541e10d2da8f85b2355f377d02e6606ded71d
z3bb77d427b68f029667faf686d174f67828ef6ace8ea7c35d78d5c1bb30409b6c5b87eccdb75fc
z4d1ccecabe8cc64971695defc8e153902b65eaa456ced85eb64868ab9c401e7ac0edd43b20a119
z295064e00d1cb0c798addaa742c3d86572efad5185bc6dec235b1d67d87e1f61e04fa8b99e2608
z02786eb04b0437812de158404dea096f424c289ade466f2996dc3f91d0dc5abcca863352e7e463
z95aa10541f3f322b68b9e0df50e807a7871270ded1c9a0a03a9616a1b3bc5293579b58b455a0bc
z38065219d3e6129810b6d26058bca6f414565b9b88a048fc4cef563227c413a41e2c6ba9151658
z970d9c4404422feebd02ca4081d4217b009abda17add3213e0187680c170d6ccddb30ea9af33e5
z445e406df95704fb31642963d6dcca5ced818f1779b209c689ce13fd300edc7743417267a67d58
z0d8e9d4829f5cb77a02ffdf78dd11e751e98046ee223746685d76c8ff165d58b770cd3a85ed344
zc4fc494d8e12e2dc2ab1cd964b3fbed3c27516722ef4830a6008760fb4b8dfb30c52d414175684
ze1f646de1da536b6e47870f49f17ad53154f176315e60d3d9341ece7e808ff9ed37a49633c10f4
z77b3fb9dc533701cf0d8cbae3ca3a0fcdd1839e32f3add87b3ee573a43e2f56dcc9abcdfaec85f
zc4bb70af4131bd8fd203e3b03a5347989cc4ea2629147373e2ea69760f635dbca9c45aa0e3de06
z9b359799fd4346e7d58f4ae1e2b60340ea874d9ca3d3790b012fe683b00b4d99d199e1a4c6852c
ze268f80a48c9f35cff8e26b9360ed33ff234d8efa8cdcbe8d3f631d1a4832c1df1a9338b4585e4
za58f4c1b00dd9d3b7a6e5df673e849f411a7b05d0917d7023569f146334fe2f7477cee961dfbe3
z396747ab113da81764880099e220d87604ffc97608d0a79d5040f68f3aac40706bc4270373c630
z0f2f40c6456ee5c65ae9bb3ce34f970d2e381b13393f0ca9dd9b475d2a925e69a5048abff939e1
zd1fcc9993592e8ed72543837786c41b8846d29d3091bdc709dc016b55993ece40d025e2b882010
z9d8f4b05ea7239bba1e50b0583ead0178eedfdf66471e3f7a5ae3e4c485a47f0e9f13a75010755
z760c04b616968dbff65bedb735b9d90a434c61263909200f0b7d3db72fa42772596d2cbd974611
z7f1bfcee2e584d0176884b64a88db653e473f249e24faf12ef332238b84d406507dd457095731b
z47f76e405a75ea2bf4392fefaa178b88848c353d0cb565e63d34867534d925c2f1d7fe8ed1ccdf
za7590b431e57381e3a41818f97d9a8545bacfb56f072c3baaed82ce3cdef07e2885486fc438bcc
zcec23e380cfe01302dd4ff12d3c83cb63740a395dcded38e752478d913d1421ef18c24eff3c5e8
ze45f28e4993a1e51e3a0eef6917f57fb73de4b685f4e8c25dff62b25ee010ead70e6aac24f9e22
z7cc3641b531e38b47b382ee4f2970f660649e606042e2fb2073cd81cbfaf647d21c7e19702147c
zc8168099647ed918de99c3565af14c143cb828a475fe18a124a6ed25702c83edf04173d2ebca58
zaa31510d41b35a348bc4c7ce3b4dd453a4668f5e5bb839877caa055e06ecb9a4adb76796032eaa
z186df007a5fdba07cd4f8b8f90db34263520c59009791edf9a6bb8835fdf4985e6f3dd7cc64ec3
z0e13f93747ec8386da57ba67c7e551c0fdd430aa554c7e3df54f4a8194f5f7080e26f9f710e733
zb313603ba09fe1d404fd55c40b75bf566d05ff5bff3d3640c7f023ed2313741971512658751f28
zc0f549fe6498c900b4f8cf0b55c2a99fa4a88d84a2a4a8ef1b0b8f595af5a3d7c5dc48c220f0c0
z262118fbf395c1ea871e17f991301d0c2f0e91cde05955fa82c97971a76a53dc2dc6e9d11be0ef
ze8fbf1ed3c125a4a67602c79294eed564fa840372adfaa760d3d50bb0e5783bb8c4e0b37c3c30f
z9cb7ccefff63462288d4923138f9107a27891e07eecc54019d12c3164743ce3ba07a0ac27af296
ze6b37c528650a47297bd1c339797d68c7c7d95ce4fd70b75d3104fb0e6f4a1a08397827c303d93
z772e16cb16509d73641aa53538b09cda163a74e69ddbb3a8a45a0d481beab5e4526bcbc196d725
z02e7e3f1f1291d83864dcd08e9a33bc15662da97c6258193f8947120f136b11c16dfb908228e87
z71fa165b9e78423609096df8ca055d228d9bf626eefe3f0f855f6ad11db1b123d7c4c6cb370df2
z822a51504f28f5855765e7ade3d2353560dfc4fc7eeb936662006b337caa7507adfabc82c6da67
zfbd14bddae2daceacbc04e14399e21353269e02d18533c452df3de7cfa203ee4b8b370beba58ae
ze3ccd31a026831ac4e51015c74d2d7fb1f83b62605aa53f6d8d5935a808c47b702f74486e59bb5
z8d9c15cd89e1687b44ecb9f9aaac9b834ce7af8e0ff98207dccb163162bc85011f9ce4167739f0
zfca1db8255de5939b7987660d2190f3079acb3ee370d375fecaaf792f962fccdc13c9543661a27
zc26d5c2af1a0f030f841e35fcff19a240ecf983ed440782a1dacafe8a205279b8b186f6d44e136
z56cf6457ad396da6b6e168ce1cefdd05d882b7d78ae3fd7084a529f3b0028790ab8f0a2b66d9cb
z8a6a9bb1465c3315ae397575e0e3b1b904732d26252b984d5574fdabdd2ba0e29b23aaa1b91eff
z2ebeef3e21076d0befba900ad90dbe21a7cafe54cc6c777eb883396ea755a0b0bfa98e8636f989
z8049db7df57649a91023a645ec7242351b2959c4a8f4a8403818cf41dcbfd961f47600416af838
z74858f9e5c4ba20a7d4437d129401c98fc8dabe8136df6d96c72b9f7f6f9840df7573aed192465
z0cbef16a0494195d854b0b744f15c556b93a0fcfb11aacc3e541c2e1c870574d62bb0bbde580a3
zb254c95521c456d626ea79191484da521e1baf144865bdd4300529a12a3c6452fe7960f698c862
zb2a89a08ba6751b4687654a3e141c03bf7bd12f095565430f0110ccc524aba814b9e4741ac00f9
z352e028357c62ee025f360918e7ab82cf24070593598d040f036a487ec72aa0d70e5b35fa12252
z0d987df4540a325a8d54f5a2980c11536f36b93b866fd500549fbea6107be7724509f9b731539f
z425990b9ab4dc7811538acdc68ab39e1ded48aa53e24e14366c9a829188debb7228403d8524ee4
z73f7b2f48de11a619a800ff9ec8d727b65b582fafff0a608674786f588e84350aaeeb2f564bd04
z60c2d08d61842e437d2340c14d77e26f43d3f644fa99ec4dbbfa6ce0828d9e0e700d4e31ff0aef
za93be4d42dc8298566f1fbce5f2182bc5dda5446dee5d4537f0a1d55efbd5be586699e95fef308
z97d6f0c8fed56a5a617019089bc3aa684d3e442647e51850302e2d7c6b7a3a9cd30ebdffa49dd0
ze28f07808731236f742551712c3562f01d0ca98535b068fb8491c2e20f7920df57c24d0b066d1f
z3e60743a58b7fc11e5531bac2d63279efc02f7763eceb4491b6fc33971e8f41a123add43ab1ba7
z7cfb117239361fb0eb0534eaa48f9cf99d072d7b8a6df52408d74d1fd6533114cd320c5e563b6f
z22ffe88a032a3f22c0c61861271a8880a627cbc5fddd8b8515d1e90a52ff82adb39c150868c3e0
z209430cd3ab34e9270d2f774d3019e2c091ba50f4a4b19783460d9e010f47c11f21120a434c272
zd3848a98403ff8f78f1dcbc8e8f8e4d01f01a12276223c6a2bd0cab9f068a010f2e6bd410d1d73
zf0cce288cce019451620901c1ad374877412f0b46c45a213f43c6319cc82dc0a5f0ab537ce25d6
z70bbd3752458a18932a56abe6e6acf2ce9fc7b3ac817492f722fca0a3e9b48536e551a2d4345ac
zb5ec6f28978458c8fe91c1a45e7e8cd1024ff1dfb5576a34131b92b9602550a265ba333e56a8f5
z97f6c8bd442617e5bbea8095891e3b223162bd96b885139e9be17ee197d345ba8ba817a2c7525d
zaabe52642c3a30637f5840c29e479ea04126c7a019ca45473d321de9009ea2647fd4d0900a2454
z28e0498d1762f19e1e626bfe78c35b2c68dd4da3f2116711284c552daf2d90c752e727114d80b4
z3f9ee721ed277f2827426dedd3b865e1293351e4ac28825cd4a27ff9fa2894c06c313a894a7648
zfe6f837291645efb11cb9737a9f81dc433967d59920c0e3821c9583d0f66643f8d0c3da3eb075a
za5109066914997c411ea54fd95650229ee52ff9e89324762837080f7a8accdb0c20bcc7d26860a
z9f4414a34fd2e4c7d11ec136997b51cc0fe68b3244cb46f210d8c3cbb6f652d21d5a2655140406
z85c69d2c40cdf3aa1408a79c31f3932e5a8b9d20a93d3acbdb463e9a9440040620ad7ab260f0b4
zda68d7591c8e4383999e052588a506cad96266ffbd30047b530d0313dc1680571a8abe6f361b7b
z88f8c61e4e20402ea0a54fef6108e501fe79f99b7e6eb3aa483efede0addc9af83314971fc9cb5
z903d5ec511718fcbd20bb557224814fcf03e1e6cb025360c07c98e460b4f991c6766f8d233986d
z055041dadeb2914227086bfe9e55598aa72af1e00ca565991314bb902df60297d6f320897e42de
z1bc6a6dfb300054e5595bc5253afdcf54065dbe3a53266c357a14a96a5dcd34c3f848dbeb12f9e
z1e58a6bfd956b316cf50c4d0613c90ef24682f0825918a108ce0c6dfdc514d78e5b6e51f973c77
z625b02f826afd2f383ba7707b639080ea9230091b84eaa7c04079a94f564ca68b64a9682fcb69d
z4db3f41645a9df40ee95991fb2dc09d795682fc9afa1c300fb051bbb860f4f9237cf16b5ad0ece
z0e19e1a7db8fd5b9e4179fc05d2527aa13aa2896a68e5434983937f64fccffa7d084ab20a5198b
zeea436942866a646009e381f1733e9508722a7a2a32379d8a9af523456f7edd73a13b9538456c6
z1ca7ba0a607707ed7208401061b7163a606fb19c3616f89edf1e67a9fbefc6d736f9752685ad42
zcc52bef3d33ed7c0394edf4fc798a52a9e94308e9443a78e88ac6d942e3510e22c6e132359d985
z4733b0c54c1c0a1ba7e4d2b43928663f710a87b7f30f4beb9a44dc453bb389b559756d2fc85ca5
z986617bfa5d0b7c5e1cdec3d74659838a2f8ed7397f86b830232bf06641db940d30bb2b58d3f90
z65a54b2b3d78647cff0652fbbd3eaa9678ad2f6152b139733d72c904441e42b622d9cc40530390
z32843c880b114694513196c74686d2a1eac51f78155daffa183c01b7e90d76e44f3eb00c199190
z2c6bd664b2726911373d98d17e8ffd574766b05888050c303e96d9aada3e38c7ec6dedde7e3f04
z354592efe51cd25aa617172e531f44d81fe177e6020bb0aae94c942e6cab15561e295b17ba3e1e
zca449dac03d31d63a794749b845f4db2be1657449fb134106e5ee091e0ac91522444d5ec127af7
zcd782db8c683e83ec90b01f79a7136605a33d7a9439ef9928793462589ed662f3b405e137ccbb7
z75c21a9d7f2cf75b7f748714befe4ba4b20cae713b618f35c828b7e17dd41129b4d26d6b6087b0
z8472897ecf254533c13cbde71d9433da9e63e258114eec2bd6aba5943731fa44cb46f4ef71e9b0
z154ecf8819c4cdf32f0d70781b08db80332e1add509e4060d90e79edb47f05136ecc2e8e646e66
z0794adb352b88c93fe3e498d741f6caff096eb60f276c7e8a5b309e47c69a7fcc326c9a64708ac
z92fde0d4483eea777861185d22a6f4300a21ad2f7adedd1873111c382c8fcb777e9b8c1aa180d3
z7b9b64c0bf04cb08d095cb217e77dff8c0b4e350fa2ea70f9c21a325026ff8de508c5bea916ecd
z9c79d37dc13a6986745488964d0e177c00fb85ea1d5092b100897c9797b4fae6bdeb20f06c7384
z895c243557e5f9df3f7cfed5352c608a2b60758347c5f0e5d20ceb06364c3294ff43db0f780830
zd54bf0a714a9fd6ede2c6b5fa16b253333501b20e30352a7f3ed049402727197752b8fbc02a358
z62c65c2b611b528b12843caf4051da039602d8beb4ed5726f6fc25b7ced07577c56ffadc9dca9e
z0614080f7a5fa0e72f2a61e33f0f68139d0b330532bda0c47db7ee412101018fc84ba4d4366e5c
z427777cd1ca67abd3e9713a68bf69374516f2a4d7cd577d6f96f1f8cb01a56e8ab18ca38b1ae2a
z75acabcb5af9a760987d33cdd383ad0289ab3357d23a7a353211343737872cc2b190f43e2c9a56
z66ace8abeee5caf668dc2c50a0b162fa14fd5c9186d0d12cae14f3f0942589d660f80dc1f1933c
z204a7a560dc5bc8bfda59812c4e972dd7e005a05822550195680b1db0040f24587350235b72d8b
zd1cc932feb2b2f6749da68035adb2d804001ed4f92e4b7b4e92f24b4932b0ffc43f2066fdd51a6
z3d152ca758f91f893a8f57a81717809536fdb5ecc0e7694b7f8df8986deb1fb4dcbbd01c83a063
zfa6e33b60a3ba9fccc0b3276e7d09d4e8abe292858be7d792a0b886bcfd7bca87e11ddd0612370
z25b3fe7889bb3f9faef529eef152757ea07eeec467f692e4b5df5d7f9ee1d2a9ddbe703fcd9731
z8e70c23360dc3576465e89fdb69ec7fa622d4326c87af18596a9eeec3b7e0975dcc6e4492e093e
zcd06104f4b773c98749e45ac484ce9c251795ef9ab199243885b943c429e9ce7141064340c5e2a
z4ed407d0592f268091c0c9ab4a03337e246a92a45b76efe35bc4fceffd514937de157a4934806a
z79bbfd86003432bef32764eb9526cf1deb76ee5327da25a6be358f7eee4ca84d9b1918facf3da8
z68752c26df351902e4dcbc72e7dbe9c682368927e39dd32f7bae59905022c2a6d6ea7c3614d3aa
z826a17a0fcb59f001ce1848542873f3a211703067075bda648ffd26427e805883b7697370a49f5
z1f13adf4910fd5cb73b55b99df86072b4ea1662519ade59cf98ac82bc658e7b797f2fdf3cfcea8
zc0559197f47fd6d3e5e7087092c254d67a6f127954d5b1387723d465a69076915a5153750e108c
z04c03bc9470703b426c233d21282be7d213c21bb4b052a267239b27c22c125034a6a6279c34820
zadc3c8c0f0df2ba4b54a5f6cf926d9c9bf8cc71041290e09c311ac21f0ed803c38725d7f7f3f09
z31adf566f48c2091fcc0ad3795f9c7d1fdd2683c8c0772fb156704208701d6883367ccbaa30068
z30804820ca76552373c4d00e3877470510fc91aa02748d43c654624252a19d3baefe87c3e17ddc
ze0562272698c1edea36de7648554947b2ac1a7d4722f79ded79c1e6fd6610b8a3b1ecb319f0bd8
z600188bf6b59075dd28902b6bf8337ba760d0d17a5d5f1ccb4d13048db7670c1c0d4d682b82618
z095385a094cf1305a71778351a1653c7bef4e43e59be3b4d6f86dd3c567f1efec414c49204576c
zb2d1ed2c3d24b37af9a27bb88da2d4b8695f5e8d67664a4966fcddd5f3245bd71246be34abf2a9
zd9bb08013baefe40ff22aa8640280b49ae49decd745892489c440782560f9dd598ccd13ae29d54
z14d24615e1831458771ae422fceb0445b3faafcf867b77c2c09c61a16bf9daba0510f9fad47516
zfbb446e1dded1cffc88ff45bfcdf8c500548aac29f365c9ebc3b207229630e2fefd4f9929740e4
za6500fd78386f9d527414375d83abb43a1add4365bb81475515827f5de447ce51378921ebffc2d
z19085c2b0ff62263b25fd120237b9538e44c7763f1203284387162780c653cd3a7940df0bbd949
z88cd74101e0b9cd1f787f3550fb21251fd2d833451e1aacf2f0a0e3c2d34bab784aac155b296b6
ze5aa44f9fafc2c840ce3de4695e0f1440eb46391c7a05061ae7c058785575d0c3cc3b6e8dc9402
zf5122918d97163866b312d6a0d250522ac0930e75c22b2dd9ba2601668b45c03c1a642dc560676
z05143dcb148e2794ad149d744a83f2421a19ed25c3131329eceacaa2398a6feee79cc53746faa5
zd92f6eb556b4aaa5daa3b7205005327e01595701442305f6a4e600d408569e7d33fed53ed445a8
z02d8c6cdaa4abb9e08b0c7285300e922bbe7a17f1fed61957e7720894abd7fd1ef6f8b454216d1
z375cbd4c18bf37345ab8a1e3e09b1693fa8a85aac02601cc6022a4e721036839a0174497a407c6
z4cd35622a5b91d11949ec15cc9af6b30909b26df68c62af7811f169757d4e89c617dae920666fd
zaa55db34bf51d919a32fb3ab18e8e12e50286f2dd2aff720ac774055beb39e5384d758896268dc
z7bcfb5ab95e275e3a3c289da66e11128dda54869ea8d860b96f973ba7aca20e3a4d4b16d39c761
zfc228d6b58e49a2d6acea70b51d352d04e3909b5e4fb11c9e4ed4968494dc664d372e70821a2a3
zd53381bb852fe2f0984c93240a1a3eb14ae59d0449f09db912379fb5653e4300c6bbb46ba11b78
z32417c505b78f072466d88e959fc384fd0c3ad2225979d5efebdfe6c0a8bc28325134b32147986
z85f4b423db299407615097afdbc6bc764f407c5b4be02bc13533def5c26dfe6502a8d1021751cf
z774e4cd44f93aca61c073721032a7e4e22394c44cbf16e6e6aa7af029179cc1a17fe4635a2bd50
z7ba1d9e1f59d9f6f0e97954753e9971858b3a881c569ebb014d731e36f358643cd7b5aee4ae938
zea1ad90a34dd65302e09f58b0097e81199e324bd14d081ecef47bf144ab3e60f485376a566653b
z4995fa04291a2781206b76a5dec5f920149f5659b8dc5b50883b0d19b15225295bd34c0ea12b8b
z9006a9707a7242064590c3fd6efb48c8e9c4345ff3ebf9fbc3aa10ec61eecb236f30fbacb37514
z8a3a4d24f5df73d7482203aedc9ef1b6fa6e4f62be3a49f99dbd8be6bb566ca5e371465284fa08
z15cc36ab28b976ea0c570ffe6334c8dac5382dd3abd8fab0f998df655fe1c977f3f17990cf51bb
zd7c5bd1bcd5660eca3a153d943e12a1aa1b4dcd61a02f05cbccec1929a14c99357cf0dac403c33
z75c91ea8a55a7c4b891bb1a58f76394cef7ae78e8ecb07392101db0b46877ccfde80b04184f670
zefd2378b65906440db90be736f4667907287b8ee901e47004be45c07cf21bde9c6c599a1ea0b89
z5d0616b43230f8dcefc6fdd608e2c91e3ca664c7c027722184a85932ce4b7eddedeccb007f2d81
z91fa80aa9c7e47cf3e76f44b91312623ec04bd8155d146d3525292747462cc8a14583dd6c29ab4
z2aa98db985492dc7e2159d7acb480b747230d8d659dd5189eef357d56699c54afee14d82b8ca32
zbfc5280b0480f41d9ebdd8a312d0897225fb8edb9330d74d8ed1e4f092cff8f163d44c2cbb67f6
z8524e85205800195e121461b96ef4060b1884ba006c6b437886f5b09b226925f933d09388ac302
z55182785130d7f8de1541f0ae289d2d6ad5593d0a2c8631e8d3fa8e00e962ba1d4a91ac38878bc
zf07ee2e4cbb5c87dc7ea6e170c7b7ed43ba697fb14eae81b37a942600616f02123b3441d890a35
z9225bd2417ee07ae9a657ed397799379e9c2fd49d44cb28521861515579791e4c0bd5417f54628
ze517035a708eedfcee1b97b9bb1a7f6284d399c3609dbfd4698d925796587c80a732b517c6ea8c
zc242da57b9ed3b302e4703e867ae5cd33ff8163367c7fcb3b900899e274cf71691e1011da0976c
z5786072bf56227bbdccd636567b52658ad7d77eefb2549cb37ee66389550043a762f753fd418d4
z03b4f9f1ace8117adccd004811880498574e9f327e8cfc01472f1f40b143017cac4b75e67640fc
z198a9131d9cec5164040c10bf6f5d64956cf8f84893d7e000c3f551251140b344a130979690947
z3f851a4365e47539cd21ebb530916d04d2e96b83dc5e8378d5f051adb7a24a56d64ced0dd08eff
zaf7050b15a85449bbe0d733c428c893b8df0e763ea91c217847ebdca76b42e748e6e37b4ca5804
z9d09bf30e82e3c18670962712f46d784b2f619c0b8969d942567859f55ab185c1e0884186715f7
z422c47a0f4cf0d2c9aaed120462f8d20b45f25f6d87e48ced7eb20bc1d6d977bba3ce50dcb6a5c
zd749d02079e856ae225a8c40c39fd84dd2a389f545ded98acf7ea47f43609940313600acab32df
z64787b8706b2398f0cd37b8c1e203591597d784ac2497946ad184acbdba544b07927204af8d381
zf647e0bc17703eccbec54b83d40b87db835361b97630990487c2760ebc49d6f3702f28e84031e5
zc2a701359ddcf14bc13c8b0772cf5a710d56cc6d633d7972d5958821e66589df1349b579995519
z509f20fe1fb314a923907bc7c3152dbfa37422b4553c115e9fc3f0d8a7bbcbceef07919e1d33a4
z0002d433491b78177402278a3a36e478a9be2f44805a59669ccecd2dfa1da9800e05954db75c42
ze57a646955a65b27e4e21b90410eca14733c34d7093f0f530d7659ca1c6a387e244eb401217de4
za87652acb2e0aa358715a00e0fe980fe81ed35eb0a223f37a2cb21645ff35ed8ebb76d767938c4
zc98a03a9d7015bec93fd312a1e731158834376e135f5b80721a48537bade543bb0a41ebd4092e4
z2eb084776fdc25c9c591c4ae05f861a6234f4639b53223ea633c71926fa59d207503e6a4097026
z7adcbf8fefc276a521b7830b17a48fcbd15201c182bff35063173961812c4c56c8f55edf607387
z3625b3f52c33dbce889143308737ec52917ecdf4f41cd7462f69d5a47ccf5dfb2a08195075726f
z65b1bbcc97e2f2e5cef265d3a0e83faa37e2f9b4501015f6880dc46794b7a9cc002edd61140d13
zeb2cc24cbb066c6622d0a9cf186c87f9b439b25cae1dc8cd79a223118c09bc407c91eca99c7903
zc8def2083f2ae7715459079593694043cd75321b3b5db99b60aabae22bd079f55f6e8981b72480
z9711e54f36fdcca0631d91dab2993d7c9a1b4f2990706e3b653f7f9eae1c6073e698d8b8ce81be
z8c32b8c5451477a4171962e423c7476599e45fce8654da5ec50150a6a54134f1b7d4a9054aafe1
zc030ffcba40bbe309e0f38af162125a187e3f4d61ea498f3811b40d0dd0f0c5f57301ba4f6791b
z6024df94e20d25fd93255b11cd4d64c7140a4915cca24289cf448f8dc9ba44fe460312b5388700
z68ba128f69031551436807cd5b091a9359615f4c2325bff965418fb9476c2070ea5e3abdf73bfd
zfa5e3efc67ab78f31aebc11913d8b32c11f1670e0c22fba94d7b4ec1d287fc24da21ab24aa833f
zdd6183efd959210a8eae83ba952be6ebaa54085f1099331cf6e91453f0f947d1aafa9e797b2412
z23cf40f4fb2024343d37535ddc2f0faf3026a36d2f80b12f658700c2adf6c900c2aad36fd438de
z9aff59f7a127f403be25ff9dd34d87b3fdbbba3e8f79e07a84900b5f399142468b7bdf16e67363
z2187e3cf1ddc25f69e5a45facdde135bb41b1b1467228f109fc7f00612c36fd03c1d8e68a4b2cb
z0690ff2d09eac5b0100cacf43aed8783420ae146dca55a262168d7a47f0382627847d2b0b78c40
z8e838c9ba847a7bd67cb7a9d703ec6d810341ef24a1b4dd3f698f4fda11ea035e03981b23fa592
z10088938f6042484d329cef8083a895a78ea91330e20bde310b8f3cd227e47bd1ecbb2d587284b
z6070b2903c5e8746d5bd6d82edf5c945b224d57d47d7a8dac00a9b8ef03f6900063e5498e50dbb
z0ff41d3a8882f18ec19197a61551dc80e8b586637054ebeb959f49f11e44793c7c0b0c4faff7b1
z95153493521c682d4cfbcdda4a63175a74670348052d6cc07dc57f3e8c45d16c42f147adfb635b
ze46b605e6da5983ab141f1641bb0c0ec71f5d2bba6627b8619ff7b6611cffcc12545e7ea5648fa
zf3f49e75cf850bf7620c76bf1edbef7bef7406b4934bdeede768313ecde16b5872d6914e5cfb15
z639c5a01227859c3d88a1efe308fd1b4630bf34d8b20b8b677a347858dfd6d0341d904bd7eafa8
z8129ea7487868ade7882782a9dfb3bfcac541a25abe70190907d6098190ca6789f9af0a5d9d234
z207dc78c7bbffa94c6d9af857420dbb81df766602da20e7295ebf603728829eedc1d432fb42374
zf56f29de59e9e8db9d10609a7584223a3ff34d7aa075797ff48eef30b9e2f62f3e9e5a99a32475
zd37250b159f1b51c6769979473a85aabadcce3d08ca66d1860ebf97ab204deae99c1f8cbf96dc8
z40ba1cc14f57a3527c96f9f736d53129d45a1b72cc1a262b1aca9e0dc3f9b329bbef1c55b16ecd
z1d2a5aadcdbdfc5a8d2cb81de94f91872acbf5219fe2644c6121087d4f7fbb14a01cdff80be00c
zf73623b52fd10497169b04e96c606eae7106ca0ad144b25761876b6644b45ff5f6adcdd58721b3
za9f55391e6e0b43997994fb9292c4e966321ed5cf7a5b8c386a816cad5cb5d8140ddf55e1a7748
z5ddbc235f8df846a594ecb521a344d87af6502b3f823f9afbd0b7294b7056f83571b785ae31ae1
z3f7352dc527f3cdaf808667d24f38f947aa6b2e1df83a1826071633b8b82067790203ff11a0772
z511533919bb8c50f345dcc1928243283cdd0e2d6f1ade3ada038230e6ec36111940699ff6b1f5a
z6a7139cc666cae49f2d14abe40714ebcae9a7ca8b5b3fd2ae4f5b49b5bce227477fab86ef5af21
z439507458f090e9415826651e0ba5bd4abee0a75dd42a6030dfe5c3f5fc0691e2928541ad6f124
z31e0de1168e05f892b20b216f8880c375912df5db9607993f3c60377f016dbdbac5b6e64f7d345
z4f0af8c7b7052d66d84c997e755a89cc05b6e4f0eb32afbe381c24b6d467697f414048c22623b9
ze1688dae8e2347ec3ce2b7fae78b32cb7c2e8f49219a56e7929102a64c4f08b2f5be99f15f5c3c
z74a312a093c402d38b25ece19362daaa6a070144d89286a95599ef1f529f64d18520d69f1fab5b
z061efcfaf2877dcfbe88d93f1caa232e545528541ab18be0b015af3196fcfe6974eaffcdf4be92
ze983e06b7eb535acf55dd8f330a39b30b4116dd9dd93b33216574b79d5d285cbd9b8b4d6ab7f5d
za175bfe6e16c64c327e248fe8e48d31e3b3e708a45c1931acf129142d79c90c9a6ffa3ccdf64dd
z147093869e2ed328d71db8fd32f9a64a52abb14291014b76d65b2441e378099610822521955854
z575c28b619d87ef6d53c208092e192eeea216a81a81051de3b67f67d218f27f2c637896d45c4c3
za3ad319833d0ca85b0f8e42f09ac13d362621fa83c3036cc562b40afab27a52a53362aa15eb671
z58cf1d0f2f17637adf8b7f7fe18d96a660b9703a950c625fb8b1b9adaf2f3542b5cffde94715d2
z4da0705874eaca258f02a32fe742668c0ee997444b754aac3653a2b0e4bcbcd2f13f97257ce6f2
z8422e746dce9cb51dbe05b5e81bc9b7ae0709be44b84b4fade97c713929018641147a9514085b0
z4d05a483e7752f5e8366d7309fa19f0d23640ea3e41a4d704cd99388bd555232cde88b0015bcca
z35fcc5e9e05716c54fc10c5ee93de58d668bb413bb0cd372d8cc878088f812204933ce1bbe5111
ze1d5e1dab06c9ada6426247d0d98d61ddd7ecf33cdfbcf7ff0c780a900c71b4662d2d51653b002
zefc5a0c098f53d9692f80b331da6cb0be36f4f371e0c7b92324d8734f15cfe0178dae241f108fb
z01b7acc0b3d3b02564dd4d990c4da9eb84da1c639f6cdcdda7b4dc96f8f47b668a189671f51378
z634b5441f994dbeca622ba97e2f3aba33bded5d0c09650bf43967a5833184e23e060f1a30e2e3c
zfdec282ec9c3dab49f39bb33285f8869390a62e90adf2527b5c048119f61ad8f979da0dcd8478d
zea7509a773c21acb3755b28e88c008a2394afdad298bbcf85bb7c46b9c89702dc96c0406e1e41c
z3c41cb2db6d861958c2d6ff9ceb407a31d20480956f21f81b9a438506cf26754d3babdbdaf6794
zc42b5ee99b9c8dd3d1afa280b2c1b9c57afbf87e70cb93311f48732b0234e5e5c950853002e35a
z2f689aded7fc0a389a722238b62dd6693e53daac22f3e7953106d7b552ab0699f2040f41055b0f
z439d8d3f084a98eaf698b0d844e5ee439582fa71dba83c2a40b67547b7d7af83dfeeab4cd71b60
zdb9c140b7eaa50bfd06094633f5600c931fc4715cc6be0595858374e86754dcd3f53ba98e13b8f
z8d590d032f2b49213d0c04302bf21d453bcf99920428a478d2de245966c9166699cd2b1c0a00b6
z88a0aba64cdd0584ddb3189033961c86c0cf65dc3cc29e58c90d85be988a5d23d1522f343cb1d8
za704e77ef482e33217fc93b5244e6af510aab1075b7a20470b7bf7c492fb2dd79970ed4de695d2
zda05aae93d342e112b99486d190835eee5b37c42d38fe390eecbeec77bfb2f6b7d3111e0eb0fd2
z6c944ab4174a47aa1e9297c96c880f5c736bafba9ddda39e691706963c5c00aa64fa4248db55a6
z392d1b82e1ac8eab69a2a2193d23ec3ec1673034fff356d8d209fb83c6f5ac6a603d484eaad93a
z5e89b3a6ddf58f06c3884d643e321aefd4499845b432ba825d8c1f2906957a481dc5597c41d2ff
z1e52cb46a4645cc919dd1149aad2998c465589caeeab3e02d6d799775c3c153279c63fd234855c
zb387711954d0c0ba9776d86a148b5fc1a2bc568f8640c468e20c7ffeb8c9043e6c77b0627cedb8
z73277270dbc99e8f938e68d1bcd6a529ab55996f18a1079ba8644bd3e98566ee1a4b41bbe29918
za718baac2d3d4f461031e55f486a1e85aa06579764737331bf59bd7f73dac4e150f2c06cacb097
zd6b3b5a35a0ebc47d1eb09e2bb3d9c1d5ed250d4a569e986946bfe657cde0ce2e78b4ba5e1b72a
z1b89fbb30ebc4a792cda6fd875c36ced0f8b5f223382f52da5fb8cc5b8d8d08aa6998a1b3052c1
z793d9d9b2435e594e0dddc1809e76ac77d08b0fe8a4b997fa172b549369e586151149ab2ddec3d
z8076dfa3dd9dcc6faab6fd72f36d5317288a760e87b9882b9de2019591ba41557088e2dfd596f3
zc72d7bc6b2c5bc986c57fad39640854fb403ee0af1009b66e4fa1968bf72431ddd41061f3cdf82
zc606d6caf0e8ac165eca6034c19c1d82d8eb69f2d81a77c7a891ed95ebd154583986155210507d
z670974d21fcf6cad1aacae1387777be73858c5f9983a1099cfa04e5a84b4138a4c5c2c704bb48c
za8889555008ad3e364d5dc0a74d009169ad00197c8e8adef745ec475d00975d75d4a59d39e4f23
z52ce458f25d2d416ab6b62974eae5b421fad724b063e3492670e7fc3b03f46e7437de14950b4cf
zed1446d124f181dcc55f980774fded259d28021bc219b055438b6a3f9cd073b42d9e72a876b0c4
zd4623ad1cde2bfc45593c76506b1db1cc5a14c4bee00bcec219a702222e2698cc53d9d4b6ccffb
zbc820d5b38cd77508ae8dad5c008190692b3d4c911369699271abc92ef796912d06228808c578f
ze8f8f0e1ad02d5a8cf3ab047fa23466382c05a0824cce6ee6b798cf2157af9e6cc1c012ca1d70b
z524e3e01911ada4cc94f24686be580684d96ca3b4c320d825c466c762e9e7f6e6ed0efe8e73a1f
z72472d059faea5497dfa0fee87d915896ed6488db310d65ed65806fc6f4a38bec9c6ee29f30549
z72d020541e2bb4d53c02fdd3b6bf3bd2c1f275a831b0d7c565193d1d27a798e9cfb1c08f7243f7
z1e6df8432280eccf560a5f3f2258c3ea4af185e1737dfce0ca9abaf8eb558e8c8fec1d9bca5c71
z42144fcc677cb0c7c99bc9179c626b2c4a90e608195b50097c363d6eef6982b893c1ab1bccda55
ze021200418a920e0b3718d5b03c732e7479fd688e58489db2dc3941ca0aa6c53b2000b13597b39
z0c84892192e8cf2d69f3b624c2b454acdab5bd056ffa35fad26e97d5ecc1da9c6c7434ace54de1
zeccfeae192155efe4e981a41b2af80203fadd3abc277c34ed9a1403bf5856207ea1b1a83725858
z86db1d11019ed877e139085192867440f0bd083fcd32d2aec2c723633ec9edd72260d6b5bc11a8
z99c2e157e5b4bb2822188bbacb94047259332638d3ff6875d670b04a9223952bd606db82f80446
zfd78fa4bc69878c1348a13c1c99e334f36714477f6c8558d7b1fa96ac0e16c45524bdc6a543f74
zfdd24d01ca638b76273cdf2d36b30abec0f5b752b3feceb8e42cb5a449fa715975166a9b063112
z6eabb259ea5fd9e4ac5d041d194599b545a32895da8ed8efe455a6bbce003c76b8183ad5a09fda
z967fb1035599c6e0fe5ab08b0eb97619a35cab2a0a327c21516966fb3d92d5b85f6f9a3ae4a440
zff3c7eb1a1b1f5f0579de54dad8a6f7c8a9499fbacea1211970c0301bb38966dbf8902608b361a
zb356819e612510fbbccc5e37e05073069b4a07a7ae47a393ce776db52765e16954ef538df85d1a
zbdc33039259cf9761498f417d5b41c870b8fefc07ef767a0c2d379b8f2ac3189eba4bd8e957024
zeba95fc276c3ce69665df924e224d9e9670425c9d0d0975227ad053530d40668cc3d29e1726d4d
z24d28a69e241c5e92d2b15502cbe2d5e90f405d7383b257c217e706cedd90910d9320d562dde1e
z1e0daf2ad9c972b60da0612ea719ec1ebbdb54e24f68c1eb3649387a7fdf7e71e8c08f835b687c
z345659245e994acf0e2a8fbdf79174d427237410019beca1ec6d851f7770112c07abd3031b8392
zf0f37c2d43f4d4b894f049b54efeb3a5352af294a5b0b854c72e57ae072de7e8edbb844564adf7
ze5eddee5f16d73fa2f16ac689dddf6a18647d17799833ca60be12f740e9b98fae33b0eef64f189
za812876dab2b6082912df887b755c5ad4fbc84082c136dbaedec3401dceb30f9a8389c26d97258
zd36d9e14c3a7604b710899ad99f5e6a0f0585b25f755baf810431dec2488e092d41f3c63443fbb
ze36c5cc0c8020d78178ced6bc1a96e354c08de97d892b43cdda38e16d4e8df2805b3c9448d9ff4
z12ba45f14510336f75304da75025d10911d7c3f34b68dd099b5dda88c978a29b50201338d8517b
z23bc9faeb7f292588b9ffdb11d81671e16e0365373b13399b9954500e91b62855c848953b0a635
z10b823a8cc743a544c72796bf209956ab8c1faea1425910b472efbc276fc80fb338cb85ae35500
zc5b72d61ec467e30f6b3ef998156c8f5cca6a7f8a1730f15921caa0ee05846417403ae5ac38ed6
ze303d75f94fda8296134a8b1e1aa605cb1e14380b92a892d1671e9e32460c0e528bfcd76317424
zd279d83d26eb395679c74f38e2d556befead3cd431d019dfc6810ab4d9197e15d4824ae55d4843
z9135771d53215fa3fbe482808eb65dd151fdc0fd3f7c224cedb52a1056578cbe873db520dcd8a5
zee9999662a8b29da3844c013c0121e335990108fda67c778f5e720bc06a8bb4cd062e85a358943
z68baf5d56947dc396314b9db8db8dda64b3d1c50c3ad7e2471075589ac3f6cd0382c4e8157d4f5
z37ed19872303c2a69a44a12d19bf0c71728ad32e2d859b2b8d126e9fd141d2c9ab4f53fa5b4fa7
zb1f0a427c490df46763e21d2253a185871afeb1c55ebd11bb753a8af81db19ca1ec3b36cd632cd
z0e37edf219caf622fb36356c2deb230ca7d8a3c02fc624c34f8a2ae34f24d0381910f8cc51bddc
z9f830602f6e73995818f37305af158c9564c424840b85636080b34f046e2ceb69f4ae82beee778
z6815cc3abfa0bb946b229d2c9cba2c063c15cf34194a96814623a15017725057e079b41633a629
z36b0fce9e2773c5083bdfc468ad090d968c3e05af68a0b1382a4333655e09ba634a057a7944b61
z50cec1b3b1a5371617d20d496bf4694ba7a3cc2d12de4689f412d44459af33ae5bcfcbadcf4769
z7c55ce1d897651b40f9bafc8fb6ec0a6b27e9d4951b7e0c15caaef05c67df7eed2a4e52cf13e9f
z5a82a3d6a78534bdfb978153362cab292167af0fcf9c191429c7f1c09d542b2d1dd2e2040d415b
z13c45279b734a5b2ab4cb1249b8351d7e6b3337e73692f0d51bd70b79d5c821994a9335ea0d56f
zb40c4661635dc7b7a9daef3c89f28ee07e7d17c4f4fe67dd33a245833087197fa8776b4435a6b9
z52a7186408c7a6f64cfd538bb55a2818fc3091829a683bc428843ba5209ad87049e3a2c3a97d28
z6dfdd12877adf37dcdcf3f2a7289291268da636f982c48bac1cae640e85cdb606749cc484d0b3a
z45390bfc470ddbee49178088765db5c6f1e1308a196da789c7d0ace520cf847a6feed038702368
z816ccda4922d5ff3e76482c7182baf7ff512ff01e8aa1a1095d89bccce113fa981a068a7de8c99
z03d1ef695fb63e0dfe5a22a6ad72b6034b0e3cc056f06b2995c0b2be60529239830dd37cdaa7bb
zb9682377caad4d015caa49edc1f7144d6c049c73aae8e9ff94970b2674bc2448a3a3af29515425
z050b02c8251e83de7bac0d5e260e28241310dfb9634368cc00dd105591f57bd56ea409274f59ed
z08fce6804b73124235c421254bb16378f0439fa0e1a52aea35958dfd05e7b4643239a03dcbd553
z5947ab8208d7bd62732dcdef39396597a6431ae95797d493f690dbc02186401872043ef3b3f9d4
z2a3eb407f38311ea1ecea8128e91deca379f61b493bf828b414705fd9f8195713820c67ac0b97e
z905b02df9cfb978dad6addd1032828651881eb00036905468591146af0645c5da7d1585fe84f58
z3b7029e981aa1b5009db0db9a89db4dc24a9e14325eca34892e060c408b897b24904292104bd98
z113724db0886eef007f455da7318241d211b5678c58719357de56bb7fe3efb90c025899f79ad29
z78726f60ce3dd5c791a10db3e4bf8b7271e8412ded9c0e4e650e2f8082342bd3f533b2b99387da
z9a25d2822d88b022d446d1bd8a75ddf02dc858071a9d1453f6d7d3cd28dea07cfde69741c32802
z147f9de355489950e64ba4f672e000c01b1571ac199096c83530344ce316a4d180ee7a8ee73796
zb8d863ca0e60159d2997817cd5b95184c76c19eac7d17d5ff5fa529029ae04367478f6086734d8
z9d988c1993b81ab12c9658f79c8751cc384c3901fa3e865436dd55c7d15ab2baa429d9406971f6
z8c45bf5465eecbae8bba3a6de6bd64f5cf3667eaa398c818777aa5d7d37f9c6c91e72f63a3d9f3
za1228f40525b59f3ff702c2ff71ebe82882cd229081d91592e8842aaf4335211043674594b94b6
zed21ce617cda495b522806b06f7db8ee84f92128bbcb1c83cf5985f103e0916cfea02c99b3b4da
z936587298f2c4c6e881b5cdbd04e1dbf2de25e010d0fa3e4c3a1795fa0e8bcd3931c54eeda1bed
z65fce8661c7d53f568dea9026c29998a8cf795274a3917489e1a6cf53164ac45a2fe673fa47e0b
z9a144138498e48838a669fdeb6c5a1f0ecbe4392bce16469345411b1da87f21f142bb524da08cf
z0b6ed03c275e820089e63df58cc15f397ffb51886e72718d8f46f242965c6000412fb68ad8b92c
z0442de57ab6a352b36cdfecab7a036aa1ca24a8af1deddea850ea193d1c50c0452ffde11bfd8ab
zbb188917380aceaf85189dac69583df113d0e39b9f3bb49ae9d82a33b838cea97b40691102b6b0
z25e131124a1954772ee1afa44dce41fa49ff69033c66c0b59dcfc9f8334ccf488dc6f969d3a2f2
zeeb98ff0eb125346a1e1d4f543a74766be8442d72b8d72f2fc1a8b14ade9a8f47f09427fac1020
zac2960a7c6b96b09357d712d1e4998f760fbb820ea8d4f442efb11c9ca07afc8f9969433231943
z599e30a7b17ab2f263a36d625d6d7975b53be8d36944175e0b4459112f0b313c37fe4fd0f3f3de
z188d42ddce21ea8443f507a5a47c101f0e32cccde59ebb4aa5b2b17cb49e6b72c7679783bbe26e
z745ff2b74c2fa9e851d0d592d552502a217d581fef05b09cf036ceef021fe229de2fc8b5dbbe84
z4569fec2e7daca79cc2e53e21ec489b39e14a29248b8d58169dd1f313af98231850b6c42a3284c
z2779e973aa574f39c78a8204fa88ca6acb9cc32dcd3e50a01fe3705a7be6b8815c1a721583e825
zcf0f6372fef88e3caa743bfdf66bffcf25ace1faf0071de31020572372b385afd49bca3c8be58a
z6b40ba4c2289df01050f08d6af90997ad2bfbd153111a38f4cb0d0dec6dbc38dc0094d1b69be61
ze975ef43c1c390edec0c04d8779fdef1f2c3c4599f2838994e79ad1be730086bef712e1c36ffea
zc608c72f6a4162be422f1a8a2d649172b901a767fec46e813d77232f01ea1f478c07826e732364
zac77ecfe3e2c6ce132ade432c13058ecaa9c2c388f113bd46c8434c0939daae11a53d48dccf600
zb8e85cf2a93c708c9b9ecbef182280ee5250ce70192ae2e31e7d308e3cfd9fc957941afa21e863
z5d0671962aedf32d31a48501f5a051fe78fbda476e51e6327a72c60462008078f54a403597210d
z3829e554f769247701bea7403468f3f3848718be4b28fb3154407bf15e90abf41e9a9fb942b65a
zf3abeb0323874ac49bc0686f064522baec8842863801d5eeecca90a17f8e770d66c1c4eecdcea5
z948168cecafbf4be31dcf4a820efd114f8f3c579bc5a4f4f689204ade2d211fa590a40fe7dbfdf
zccc826052cdccd554624d05a0c21c7d5d71fa1cb6b6450e53d8a620d06038586e097544bfdedf6
z10a4b4960bb4918d7fdb3139bcdc169288ccd324e069368791e55a2ba4bde5503872591b78a02b
z7ea21708502f80b8cb9989d58dae6828de68288f8019eaf1f2bc137a50271fea12ed95bd3f7d80
z9626254eb0ef5d9c76223759fd99d981e1400153d3eaf4b214b417e219c107e4bd8f097d2b05c9
z73e920392bf6c717a6f821491e62b31ac92b3d9efcb7b5beabca99dbe0d8afaf66915ef17b92b6
zfa02ed108fe50795a536a7d2286344701b4d2a2c326af02a500bfd29ed71a5f99cfbceaffbb540
zee6656cc6c91849671e22d2d023b3c186d3cb30eea495be0ab1d126d8e4aaf42f59efa49564769
z18c6be0c98f0dbf2a4325dc291c7329b5844120f5bbd67a8ec9b2a5e7e85ec7b9f7a24bf3484c7
z21badf9f275dee44d9a51d05685605dbed3358362ada6b1064c2e042a67b5bc7e0f34d554d09a8
z48abacb201ef210b647b2ff3d49a0f1eafa1dc033872f694591fb30dc90748e81e467fcd293c0d
z824913d5e4103b74482b5aeb7fe3e7c92dbaf1818f127bd3303f8b23c252a0ea1d54c80e2588a4
zc7223b1f152f15bce6089592fd7716483e0bdb745bd2ab72cc9054f3bdbe5f40dd43112882d115
za3cc7bbbc11bab328e068eb7fae08e6e65d1bc598714f27b874226feee7669ac211edd7d0b1571
zdf4cfb9f81075b89aebd26e83da47984c39e03c53ea42fe90392f6fa7cd486d8ca5b6fe06ae442
z0a5fa0ed081b4f6710037c0801e60a315ef8cf299c966e01bb1849787193eb786034bd91fc8308
z29d2f34fe397399a5ea78d24992f3bc1263a4c2d4061e2dafdab17b34d2ce7e675dcb109f15122
z1169ab018bb3f8e9e056d8b757d3911eccac6d70bbbbb2d7b7f7260e87eb1a48be110fd1b5e6ef
zbab9655d06de70e6be2422be4426a69616b4b76f8996c6bb1dc8f147d93c4e581519071005ca91
z3a97c8da300a5e6540b82990a24b3e3f703490ef37455f57c1b2cd2c5ab0dba00e123108d42965
ze895911263261da00d062c7d9f2f8f0fca87bc164aea897189514e8efa2b09aa7fae6c2c88bbe3
z023826b4bdcb98d94c1c6d3e425397f9069d1375e919d058e13de5a92db904c561a7eaf0797e47
zf7fa765753c2daacd6c0537fce46a0f5a9bba7514ac83416e6250a3f508019c8a155ae53366f49
z0e807aadd42832f6a97631763315938842062f175555d0650365afa052f4ddc86b84519cbe4519
z0d50b00a3d1b2c97249e0c666cefd0ceeb1b5cef3d7003cbd477b7daf3c836a0b7b0afd904ed2e
z48b79f6f6a29ba5af8a2cad6c5bc464ded684cec1488494d192430c7ad545b0296d56d68513a00
z318189712e4bf304937b698bed07f8fedb31a7dc14c62d3bf8400eec9d748d7a7e3951b8b33c2b
z6e27294469f7f4931d20c0bbfd14095530b360d5b3aacaaff49eba2e77adab13acfe79feef12c0
z375a86cbc7b631893aae352ce51e6e9635a2d48f383d7d05f98e80df8d60f73b9817885fedc892
zaf66e7031eda7c4b149243c1bf164c7c2ec99d4b1e538927ceabfa328f8b335bfedf67d683228a
z41a47d96c89431b310fa9d0ed3d9e1abfdba88e3f86d30e7d72d8677f723cd575f14a73e9e401f
zf022bed0425cfca52ca3ffad50a62e54dacb593c1f95091289845da45aa79af8b35115934f2d0c
z53b559266981cb4adcf88b6fe7205a8f51f11718d5260d34b951b06e453e8d1e2b74e63b4d83e1
z85b65f1e1f5b46319fc19e9e95232d13f10695b26d8ceb3c6ecec6ba7b06c6f1bef4527c709d59
zd3cf6199bf5356892a4c2c7589309f1005cd9d086a9a56a35ebef4ed98a7fcb047778df78abbc2
zea7d9957c623523865ee57a0059e1264a5135f6d08e74b4a31867544257aee3ab306fef7a93204
z415369b39c678b07b4791604080d2158a76cfa3b4a1137d38ae90d497160876f1108293a87bfb3
zc27c62b92004c69432f918ea24f256d92b6e0d91d2eea6fa1f3c368ed6ef9e835411cfe5a56834
z31b711c1a91d3dd24a5fcb0e1f1af3208579f22527e79a5aa3c762a52ee7ff3bb3096b30e9cdf1
z3037858f2d85936dd954acac5fe6db8643a50c00cf28728671c9671e461760d3df6e1ddcdd3157
zd621b055251b0d1ae67da44fc5d5b9a2c803af51168493977538829511717fd4b975cde5a9ba19
z6ea12860fe7dd72ca5c3ce1f335576a85c9b36b52a333e23d88c35f97ced3bbdb2469373078840
z5057463b6f619e3b81d9961120126d6be9425c1fd64015618516a463283e56740be62e6552b45a
ze122cf8acf1f8f2cbc9bf7ad69034bbbc11b370e894a5a35cd1ec89e04ca7d9e3b254088c37da7
za267584cfa23539276ea6ae63347616a29ccfc9273406c10470ee1ca6b662f89a363634c126272
z23819771a1589af5ed6dafd80bd1cbfde93a0dad312bda10a2d9b4274eb46fb505000b2d12b296
z6b8cb79d4e2b960dec3c12ed783dad530153ab7fe75878951edef6f3990804fe4a025b66c152a2
z200f40733ca2698aefd4ab1b212ff549089d7432da1f564cea1314d4b89e68ac6492bce37f2322
z89f65b3a60744ed06a60a577b91164bbd907cde754cc77daffa6a172a3e316f702dda3b35722b0
z2d8a347621d31bf9f2455be51fa0d5cb4c74f129142cf656d035163ed42fca1eaf98fd040fec44
z05fba1a5ea1c7f4835c3d69924653c2418c3d91e31865e9267e85b9e2313e832340611fe872fe7
z447c961c87bce804e364367168f4599987437e50dc2aaa10b579fe54d6e8d03042e7e3d0a7259e
z26bae80198c6d34b42096c03f0691df53ce129fda8df0b07c704002a166ed2f91a78e703c83fa8
zd589239de64995ef55774cc35e0bdb76a0ac05bb32a7fd424b3a6dc91276be94eb2f489cb9d0f1
z0277e1c8a25a9b791730a9b1a40f6c46c9f7bb6e3175a377ecca6447a258ff51d1baebee19aee8
zb63e1578b2ea4acb570503e8de4e96c7343c07d87e5ab0b753f272cfa3d1695e4ce95137c90201
z15226071ced86789d67bcfdaa6f9f53a205f6bead8147465952a20ec2b3f7bcb3aabd5c843475a
z8e64559b5ecf44c257e3ef86d367e3b51d1d88a698d07da383d943f23d0df7cb9077877886d712
zfd13ccc77b058ad77a4e85e41128231e36211b84978cf0659563307045149a2675b36cefe5179c
z5dea61e07e7fd8cfeedd4d104cf9bce95607d810cb6966483121300d8197bf42e76f020022fb58
zf56235506df8046dfb01231a0299885967d05b8d2b9663522609f0306fe700fb99fb65971a13a6
z9c594cc88405f8a316394743fe2f7bf40902648d1fec17d4fcd0e43720760ab7412aef466343b9
ze244b922f5018d8af3c8a8f860ad28d67620068ae953ad9ded1efe92600c931c295310e4a18820
zf81075750f3bc605c42c3c14bcb2f2d57c42e9455c59c1ec569b0b377a4e85b7d8886eedfb7a6e
z1af888140daf6d8cff3a650920a5e00f04f6a25b63e7cf74930f242569f83afc7be3ed179cb8e5
zbfbfe5a189d4d05a06e091fd1c7dcce8cfcb401dd27b1b738a7d23c0b7439f75cc07fa2db51e63
zb2dfa8769d7300ab87f308af6cbf19616cb2fb6bfef046163067f3443fe55cac8eb24eb0b46594
z6624e7f6196e0b6935fd05f5f93745d5c3178942c6ecbe39cebdf692a1844e5f443892accadf5e
z42a629ecfd40470110b217f6856da973130999d3af52bd742b165defa4ee17d175d8bbfa7b5588
z687936294cab2ca5db98040db7037c60013b8e0ce0a8bfc068c53daf906a8422d8995a4b00e6f7
z265db215a3b110db2b24034c5b44fce4c09269f3f317d67b5639ad23a6a17182b404189eb0d8ec
z702a03d924338d0a8a01d37e5af1adb93dba8a0a9eb91b130cf4d0e94fc27bdff882a004682b43
z0eacaaa07e373c76e649fef5f9d1fd0ae3bec13497747750a94782860bda14d005b27007b35835
zae1e1286181b7f8116e1e82205c6c83d204d47bcf81c7e031be200f27905891b9fae4efe6ad5bf
z2271ece9bc02a488e964247c8db0fceb8398ff72925313ad3debf4fb3727769b3b5cf20406235e
zbb3c3e75cb613200b758fcd27e67db1531c789e0fcb5406cf5b81475bdeba6f4bea0f5221606e8
zf5bbe81a6f8c78d99d5f3c84c29b601616e7886c8b2afbab1822f24cb5dd97d38975480da30c86
zd7361293ed9e266e2d99857ac8ebe944f991e0ca31f597e4f196110d8eb8c521343b7ca4627916
z29f63dfe3d377a3e7a2bc77db78117e01567ce8d2c6670b0f687e6607f850af441fa61ada45409
zb4d547d72abd2cf3e3a61b61857375f890f038b701bc978970b10eadb129bcaa23a70734f9699e
z090626104978fadaf18bb8404d7cbc33158f02a41c98599439a8b84b7b33c7da8c78518e0fd6f6
z2bc9cc5c679e6e1bca32543d096ba18008be7479d32da7de6a08a8e7520e4001cd9e06713258ab
z7c5ab7c06b47e18e5f2ae74ce8c285f60c8e3d6887dd1919615266d046360aa4d90178aca47fb7
ze44b522dd8f3ec5c01fb0a316110d871b035ccc8f241c1df8f7f6d2a097d684860e5531bc68e7c
z39ea9e3093dc0e5c547452f10675be969c87037dd517f8bf81839ecc7c422acccdeeef639506e5
zff1235ac7678443cd57668a4202f3f65cf5c0b93c0752cd6cfe4f4f28d3ce98194e24d75c63312
z5bd064adce968344c32c5e8b122bb80f2245301a6262e98ba44c4747f04ac19471eaa1cbf74800
zc891926d7a1c31913b2ddf15dc0748692a4484176b9a045ffa68874963e59671bcc5f67792f121
z23feb45e3068e6366c0de8eb4b617c006c9aa1716d17bbda986eb63ef63ade84a68c1d152f02ed
zd403e9141ad23b483b2968a7b615458f5be59a8d5ce8a367eed25dd622058f879b7b97899c7625
z4a46c2fb61249715fc4ef3c60a03db089239efde1477b4e07090a6722d430ce3fd9eb9b40f86a7
zf875058814b3f76d83b31ab5ebc7592c87ef058e5ac7df8f71230243da9ece5d60e957c7f6cdb4
z338279679c2b4a74370d3c1e9cb32dceef7e9a0027038db78c13127658b3d0695663afaa30a316
zb77d53c6f3238c3d7432738eb424a11c0f53e0ea1c470730326f7a7df0e804ce8e2672fb21a1b3
zde12f5e1d2ca6cc79e21836805465c3487b959f0b363db7a2693b3290906781bf4a71fc30dbedd
zdb00892317afb42b53e90e6c1bd9b0be71eaae6f0ef84e21064c31290e19fdc6deb382c29e1eec
za32eae67bbc1bdcb2bf0a258641ce8d499c62fd8baaa752c63b84303903b60ef193156dd036025
zd1b60c009e1cbd504ef3cebde1dd2886de9b45da13af54a141c840dc9d417cc89645a1e0e32e80
zcc4b234e0aa682c7b87741c56b11fc65a90d2cf328009f7db0836632897ac640298aca8f5036b2
z30cf7a9102a6e4074f5627a422da1ca2d976e27831ee99868ed4517003d818a4faf74a44568d3e
z5ed1ad66d6da487a129c2ad582f20259c8e058be2e0fd244dd0b22e2c4cd8cec072129fe9bf118
z84d07e1080c4ad02fedbda9db86eb90cada5819ce81f280cfd138555a4cd1a49a5e82968d3dd1c
zdaef13458cedd671d5442ed979e35e01956eabaee5cb177410433e6650ce03a4188a873d82aa8a
z1f8b07f1bbc519c355d8676058ec3c2f15cea3e32d43f99caae7d3b1e53fa7fedc54b78791949a
zf911249549b52abf7358e17ed433ecbdf30114a3401b8861c8434965cd7b3c770b2a01a06ae3de
zd61418f73ccf730dcf4d5e966ca1fb10f0c8304df800bf5f2f9238ae9c37906171c0c30f45f906
zc0385f16885730bb935e89bac6f58c1357a4cdc0fd83d80f64cd22302b4f5bfc410a244efc21fe
ze96398beaf751dd2b69c919f3324c5af887c39d48ceba8f21c36682e039284ee3fc9ca7ce766e0
zacaef447585b11e72cf7e337712535669f5f0aec3816c1b6dd7c136ee24983165b30cf5a676a20
z058982a2e3471d593c57f9656342a64da2c2b41fb20a0128b463f8cc9a9269c7810d2a8935d3d3
zb758d67693cc30a7bce4c5ad889bc4a2a77e80b25f2c5bad078f4fae130114a7f01084a4337a67
zd3bb05133d11f25fb49c134e16e513481f3fe4bfc6cad9ac9e991a5d8719a166ca312a2ec4e093
z4564314cb31406e5a0299f86b5f104ae1f1a965ea68644d79b3edfd01b576b73975cf2fba9566e
za981c0f033ea4aa28bd9e56c2db725ef282424ea4aa72a5b3c0a14b1f053692e33b65487ee204c
z643281c66a1e9d56c06114a632e4c8a7c77fa271838355fabad839da594c8b33771939a2cee3f6
z6fa9b7a4d97b3b939911dac52f4c0e5e493b22b3375e434efdbd75a3c46b71b940c244410864a8
z6b2214cec70ffef998a95d2a4d8531cb60f5d4bf3ec01063e8be8c09133a0438d7c7fa09c22894
z1f52a22aceed97a83fb166d2e5bd04a03be8abe6a7f9cd2be221c2d7d5a0bfd987acb8e7d8159f
z695fbb6abe2782281b4a8baee298f1fc977c80128e8ed3474d455de81067fb5cf0756386621b1d
z7ef2d024f8ddc36aa6efcfbdb71ee5dc631f68ae08a3ced219b28fdfed9c8e4b10f4b21362ad8d
z467784e0c95e16bdc3e614f2d87f8a89cfb35275ce7fd9f779400b97334bc99960feee0192065f
za89496109cb8b5d335cff64c653856fb533930d3268d94ae299217e9ef187eb432313f5c66298c
z24d545b64feb8d7a0cf614d41c73dcdd81de7e26312909f01400f5de85cd01d33bb9096c41854f
z4100b92a8017ed7f042cea3c69dcde5e926a2f9ecf7fc836fd917cb0f76d1ff66ffe9cdaa1323b
z79a289933750fdb73113f2b67a4f76ae1dfae745bc41685b1975c9925c44b0612af92b9c43b5f0
z71d49260761eed1ac4d1bfeb142d1c8767b7eb34e30f0d47dad600e200ad0e3185eb8bcda8532f
zba662900b12e138d1536d289c16e3ae66decc5a3e12840b013fc0777597e1c6ada07aa0174a3bf
zae3ad5246827ea33c6e291a11af51ee5c2e3faab9e50bfff43669a0f31e6da4fa44dd038944ef3
z3f49b4747c7e9e352a59e24a88525ee5bc4b2ba4c2d88b4940e1abfc68ff122e8cba57554440c8
z9e5232e2bc8bf9c5bfc4e56c6321e5a75ca6677d2eadf48608f89fd34f13fe53b281fa7a98b2ae
z92568a1797ce14218d103e9944f4306d76fb4f9e0986eac161bc2a9f2d462d5c816aca7e050aaf
zfe64a3c8fa18dd93603ea3e6231d0131455407030c510ca5d2d9917c07628073b5b95631793246
z2e5e14707dae10d3f1c9d1b6d61aeb3771578e4464f62d107b115d7c99467285a7e703a2f7a77f
z5e7ddd0fac81f48d428c3a02e17f539fd61c3fac690aa2663e4b003a28e16be642d22a8b9de4b9
zecb00af80a4a1015d43bd0b2895205e45c5a79fb9c02fd23a0709e34486a4f5e80a504c2e2d5df
za687a237a90cf834e196f86036644acf71b594bc2f7af319b0a464c5e79fc60d390cc550e1bc45
z388ea8af60a938cb26da366c04a93738ecf9f2b1a584b0c65f401b8f3181bfedbabb592ddd17c9
z1edcfe2f4c5b6fe3c59f3024507ece74819281833f362853432d2ac9fa11b62e08f7cab5b37344
zdcae2674d53d4187933bae527766f3be9a420ec471dd9eaa2e556fb1c6c94c669444688b951e8e
zee9b61fcd48bca9cf7027345cbed22f82c26bcd8bbda7848d3d7ef03d1d6ec1d20703b60163d9f
z00745ea7c56fb1d98de00f3668927d118fd62a39cf83632eb58c687c63c8339a6c88eb793e7593
ze7650052dac55b8ade87f3d9b77c96271dabf29f1940a7b1bc2a29f955fc270b5141585c658507
z68165f6022530f24633e823c5aa5c34216e635e81d6a46257b8c0d9f04c5928d0e58655079bfb7
z6c6bf2172facafc7785a53c53bba9631a7d7b4cafc7ddb93543b7ff9ac0ce05ab940e523f35120
zc07f059b971be7eb81dda9c00d9d7979142aa6375967cf83616765ab4a206979640f93b354edb9
z18992983f417e87ebcabce9798b8cdefda3d9714cbff94d0d97ddef1cd751b8a98b4683dd17fd6
zb014f80671b0ffa1cbd0333e53564c116db8d14844db01e68039ed0e07c3397800f9253260ef4a
zd483d200ead762649d368382464c375d50f366ac05597ac18d4492a0d34504951f3ebf15c796ac
z7b1bd70f3afee721b71c41f8409280d84b860d52b3b5e8c4599ea8801df307ca0fb43064a748da
z9cf3ba0f2544eb684e3ffb11ea1369524acddefea5eb85c4a9c2a1d53d4f59244d51e5f5299509
za758aa2cb988f1a7513e48dd6af62ead5ab8a79ecca44a6d9eaf6e564e2eb67f379d3a981c24d5
z2660e60cc28407e3a32f14f8211402cab07bcd472cbfc917dbb2e317591ad41f92eb6b4c928544
z2b393634a075e4da48e3c09ed52ca464292cc904fbf7248201239a2d18bd153de1b3473a2a7433
z7301327238b490c777d79bcdb1949cf01fdaae9e8cea339fb6393ed30d5a45579eea44766a065a
z95bfac5010044d4a8e1688adeb9ba63fa069254c5e77fe124eff5fada768d4fc4e37697e712b85
zce15ea7b3c9947510d5812ea1d7674e779c994db369a36bc40db65fde4c1ab0ecbc4534dff0ee2
z64719162f5e60512a487f42e6b1d0ccdadb7567ed50fc183d160912d59de1de014e78fdbce60c3
z64fa60adbdb3dc7d6d0f71fc658558607d73b97cc074183738ec23ada6fa612774ac3109390274
zcd6a584b67b6305cb317e386b1706a9ac477ecad19d8a1df91160d5945bd6bcf2223b8e9e0b7ac
z2b1c809f6fc75040d25bf22cda1ec94982a08c3b46af81e23c097f333986fa2d943831340de27c
z22fcc25b57eb036efdd0ae4420c2943cb4a3ffa4ab4727a35abf5e80784bdbc8d2ed76abc566ca
z165c80f83ccdaae14e29bbd9057e7330fd3ef98414d8c67bbabb519524fc368fe70e614687dc2a
z07f5ba93444027dbafc147427f3044c5a3f23aee57646c33da9ba775caa92ff3ea93f6c158bcec
z54e6e2caf845b37df8fa73ce205ecd6ee64d8ed0910d541e60bce1622410a3548a242f606399f0
z580de827e8b1062f050cf2eb240d0cadcc2ce55f7e0e50ec175d0fd8f0e68f89efadc5ec31abd9
z0135a15a7977c8f913593475061f0d50b2a3988f85450feadd2db14c6da636e21dfc21a833cd6d
z63fc693390b9298a0cd3183e1074763deec79eb4ed0c14bff696c9e1715bb2ea1b3e5df07bbcae
za61cac0e91c7a2f27f5d908a15c363f55933a643851472c7859bb373ce045eba710584a3c2d1d1
ze65444fa53c178ac299c3256064b537f8521aa4c0848bdbe6242e60fb6a528e58e8f2b2b9810f7
z6be7596e8b642883ff1548038d796187f4aa421639dcd92c7e1072e928ee9af354c2411aa297bb
z6a3ad075e7bb5b15469b62a10c435225e54ff100b8898f22f4fe899a8707cc85e4452577e078f9
z2c01be0a5215aa705b6bbd75bc6e3e19b8faba215adf9a127df7ba310ae4437d160c791e14f6d6
z3c5dc2f2129b81a893e97153ba8f4891ff9feaf8b393c30d554429f6cdd3c85bc7b4bb158ff828
z57ab36e0fa8baf29fbee26c3f53388665d9fd0b92bcded2f57d2dc7ee33c888096b20ccf8fc4e6
z15a4c828f94dbfee935190f4ef03a58816476807f15a09478913a635db615a8f4bcd4c222d7f49
z19e9f3488b8efefbfdb22701e326550b063454f8c3f75db8efb4f5a601978b984b4dc2737bed91
zaca683c9c154cf9a6f6ceaeacb190414fc3d84a6e65b8c0d76b7bfc8a456c94fe8ba5c08a54234
z8cbaefda7bed2749664f41e52aeac1217c9478409d97bee7167c5fcc1f7927a015f3e4cbc8504c
zc92cf3b10e332df539e3250e1588cb4de62412c2036f804890a87f8bf1625f5b56cc5e3cb96f0a
zd51c1fc1d33bde9ea99d4e250aa5084fa9d1ffce2982cbcbb647d77205dc89af044361140a620a
z5bbc0b14da5b1aca94da569c839a962546e916ff71df494e8ea1e6fd681d95aaf406a9643fd620
z0356b38ed40a20f471eeb4501d2e29dc00b2cd242544a17eaeb951e94b46e72028452168be5d83
zbcefd20d4672b3a2a246655273b4913bc49afbf0cde4866aa434700dfeea31cc38c5a2d0b24612
z064da02189b0acda164ffd51fa80bfdb749449353e1335cffb778d9bf539640cfe078090fdfa95
zc7f7c4283e03118525379462604620bc4555990585894abf25ccb59bfa6eba1c4a194ac8c47432
z7c16d74394381d44e3be15ffd53c534b2724ecc400c471052167cd7d2d342ef24d8caf4cc845f4
z92e02fbb6f624c05f0fca0c2003b2baafe483968a0cfb918167a3912cc0280845ecf9c3c341cf6
z931a1e9b56ac874030f563c2474702fbd574c75c98fa15c1cbf5d85951a5b96c96dd7d151a77b6
z231a5cb6a9ae7d279c0cf0cad636257e944a4f4e5d1741298111336525a66feba488062757361d
zef3f7b8402676466785378f6a91055d02e6ce570bd65de4ee537f4b5f4a153fd56c89e7edb1837
z5ce7cc773bf78f132674a524eafaa8925017c4f05d32021a0c91953fee9f032f3219e14c403f0e
zd3968f5a1357c51b06ddd00994c53790331778c471e2a399d223738f652b91af6c21da884b1224
zad88f08e0a059b2249a21e0570b301014ad73fe4f091b39b3b55fe84499417c281d9eb4eb744fc
z29456ce46fe2435cdf1341d11c34f775017897991490da7d2e5bb01aefd9886593d1f44ba155c3
z9306cdc8af22b3ebe83e7006f8a81135bafd45371f0befb3a0cae9e6960008ecbac9b3fc0bead2
z1f957dc30aba5464255749df5e1464e8047f88eade0e3159557e8e234b8f2958e3697c1d337090
z989f296009f472f3ce788c62d48a89ef1713d10ae89973442eb2ff5337eb475d5ea008e6dd59cd
z72bcab0fa62ff1f498f1dcd2ccb35197c684dc30261df8c5a53a434591b522689a5eb386c7b1fc
z7f7eea401ca5d0d5be9db399c3bb6fda6d0feb678a77a784dffdce944a3d11f6c87f014ea84d04
z84cc5745a8cca9fb9944e1ab1eb6d5a86409abfb6c55cee6e474b3fb4977dff2f3d734a959d265
ze6f8bab5b849d6b3ab60f405e3aa5eb53238aba7b25eb94c5abd8cc2715639d270057b1a95cb6f
z6d29f430a4bc55081e5d97c830070dcdb2bfbbb220d184ec70e5677f67484ac2a3dcf4a1e0c8e2
z09328e1fa87f6a157f13c8e2f50461bcb3e5ec0da91ca06251a4346d2c5dd00f5b9ed2245db2a6
z79ba459a563414f9a0a04eb3cd1a135e8c87ff826fc4f1662f105e520b3df658275ae69309c9df
z8c3d3f0d358710d4113be41d9c61286c69ddae294573366e6e6955ab254d5a3d9e13ad4c0c0fd9
z5ee591c63597029c66751b87744aad15ff69afe9de67493ad2d28be3368f75d4f54f0b6008afdf
z7d8481890fc9f3f0308dc82978f4761a0abc5fe20e2adb588db339788cd2d78204f3815524a41c
zb906e00142cdcd58b40956367b14a73167bae2c0e23841623de094b75b45a7d973eab0587f04eb
z22c9c0eda4121bd53fc1da6a20a734e21e1627bb23db94063587595c54b70b09507c28b0b66819
zb75e944f17bda2f427f16032f3d4fd11e4a6669b6c08d35dbf6f555daefb555d3204954481a2a6
z1f2c98210f065f00a2ba813946e0ac30a6a4bf3687abebf85e9c5825fc789de05bc62afac759ce
z48ba89bf2a911f5eb8d64e3fc7a7c0823dcabccfb7e5e9ddb050b4379dbb42197c0ce8385fa751
zdb7667ee180709615162b43adf1d8dcfe3dd6e6a0e98a93b99b3d18297edc211cee4cf523bb171
z6d1a325237697960f2d03394b39c82ad56e9dd182d4390d10b52f94c781a639599bd18155524b6
z8406822206ecdfb3a009a152e1c1a343f82b389174479a5f0617935e6a9ac108135e30efad76b2
z719e678b0d55ece0be8a1b24cd3ab8f5dbfee2edee204d59cca3af8b0c69faf6961dd17a7626d7
za8a83b56a2ed1950031dad274d0f70c013fed1a8f476af1fff44207542fd9ca5f3c3a9b3ced098
z53aa84a1bfcc066ee4a599cfe52c89a58e641cde6cf0d087a5cea54841f3fddb9f21b5d01fcc17
zf59ebb8ee53f2c4f89a46be5a44a1c27a0328d5009274feb079851de4eac5cdeea39b7e53636b7
z628c01c3ebfbbc946d211bf9507926e72015c803edc2e6ce6caffdf0b593e1f71e56d0c255c4cf
zffcba1b780ada174db5b1fcc4f10a6bcc1b45c404f7808074687d2030c86eaec37c3d258357618
zc5336037eb5b1445715111030ad3eec2e0a9a7a3d7ec8f70abbfa26d661a3efa47f4dcff8a3bd0
z28de6404fed87c4d4d426bbda3cf63a55a5aace53f8ae502a58867430f43697bb8c9e941284a34
zd1928339d5f0e72cba07f974d6f9276487c9c052abf08c3af955baafe9123e839b4d2c5e0b1dfd
z168b5ee01d234989222f887ca0483ff06c06f7d984a16a8bd9b59e5caaec8cccd6c5678547c16f
z0c3c73d8e9c3178438ed7e955b8cbcce7be256d36501944cb72c977dc087e53326657adb8c814b
z9efff24dcaaa790e4765791494fc22715f6f9f361b3378e2240297121e87b374b2b72d8c41bf99
z87c294e8654699d7fa2d11f0135344ef49915dd27e2717ff24cc773795563eb0850957f992e162
zb4006bb5263bc93d0ce7de878323395c725a462efcbd759a06b5e6d0d7a7e09a7417dc851b1204
z869629918d1f6938727dae5f8154c9824cb360f9d02395988700d70ba3b90272399cbe72750e9a
zd715896b148064f94c8d68c25dabff1a9339d06bba839b8b088a14a241d082cf088321bbaa8721
z3156b48cbe6962199e55b5b5b7f85ec1f6f99035a8900d4ab868e1203982e07ac5708657ec6ccc
za1552c306dd09b2f485052df466b62bb81978adca8ac893ab81afcf0f6369a360935814bc2c2fe
z4faa296e2c51aa4d6ef92d1647e9dc65a5e6be099a231993ec81d93bc851fc41d4d19c14f0d548
zae37fe9f5edb9fdcbdbfae3b1dc167ea24ef326c46af17bffbf96e8dce4cff4c640d8892e7fdaf
za0c424c93aee6e61db7d637b83911cd2bcd3ef246ce1a555a72991446da6508bd590cf99302f60
z354c5797fc64fd488149d2066ae33b60cda35ed701a77f3c84d403b09f537727ce719c5db6c80a
zfe612f07545e8744b6b602751e20fe39fe7ac4c2269b7f4679469ed5be2a76cadfa2a1e30f16fe
zd994e50365969f2ec6d0bdd003eda3152f7ad83713ac69558d780d6606b16119ff31d14caece54
z0ccee988ea813690b44033d5b98dbaef36412012904295b9c20c7116becc9cd1abbce89367d02f
zfd5dba3859c907e4e14991b0aaacbb51ce922b52f0d2a4e5e9945262fb9a93ec9b375b52075b60
z0943b54141f38ce17817c9937b60203aebf1a60396ae02d6aea2258b037177c1a803a00cbab931
z6a64f1e4bf972a6f032b9cfc56dcbbeb1d677b8030a6738e6c06fc5e4017a62ef2c79b0432c80b
z5cd9aab6512aa89be267869238afe56e4e0811b74de2d49d7e5f609a13a85e21db3a1760e0e651
zc39a0be881f99f6e6670ed8e651cd1fdeea89021db3ac1ad0b6970d5e25b8aa9c8925cf27fa596
z4885624ccc5eb046c6aceeb1216c11bff42a3661997ef79809158efe01c8c504749bad80afda21
zb8fd24c4140ffb2a01c617ac131e7137e70ed7548d256a5e290b52f45eb0285728b953c3cf784b
z2f6a6f46440ecf83a8843cf18b0b7f245c6c9704bc14550703418462d6db4143b2307e2ce11eea
zc4001cd820191e34f9d5332dcb3db4d5dfa161645bbc334151c1dd05f4d37031dada689104060b
z26fdf66b665198fb0aacd7025f8c74eda51cc3c1d066651773a221a7db21bbcb1c5d1f92e10955
zcb9b2427a95aab535b109f6feb37b8438b1ab8cf4c64c95eb8bd2b7d36335c2e7eb2be61f2fc10
z3b1c1015f31f3a45c6430e375050bd5fa7794f18e94b080668d69b697631e3ea01e5e3fafb4b4a
za3d319871b9fea26a4530a8a6f77cae579c5bc83ce8661930f747421e7b7e2ab46729ace3d81ef
zcb5d9ba0f7956a2aa68a8f77c602b0bd7c44ce8b0492a5ac5f155c7706aca2eaaecd1b0977fe82
zf35acc444a720d69266c157870aacf761718bf04c628c29f9a57bd8320f2815fc92c7c96a99aa0
ze9a5fada1828d26401c22ea754d589bbb1a6e68064e5ee1bc2c271b48eaca57ad5f9e494677121
ze3a99160b42e169ac3bcdd6ba04e8fbfef3c687290541d0e035eca91f9fe01294d7f36ff6b037e
z3df8476c11ae611042df0d60d914442183e2360c0e853f9afa653072a9b3998a45d6ebbca32c91
zea51ced2852cb613ac4a808fdaa8ab09d0e5a85ce2d5f8a2d1826806fb0b2e6ab755f3a62430fd
z1207bb0911b6c0f72367abd206c133a6f1a90da9d4a1809c09fc37acc6bdb3356ce27ab912490b
z1a0451ff9de9474a4f59b847c3a97c6a3f79dde8aeec01f5b31e3c52f61da094d2d9c8c505b263
zd8aa36205a109ba90a8b0c641cce66dd07520970231a2e2846177690c8ee20c8c9deab830282c5
zbe144b500f26a123fe52fbbb2dd95d74ecc6b714e99886e5d95c23a5cb28c44fe418e4a8a8490b
zfb8a587d21255cff47b53c5bfec9174f4cfafbebc51f80562717a0f979310cd4e2388b031b3b26
ze4a8bfef3968e47cc187edd7b56ab526f9a4d28632e546dd9e69a790bb3ce65dc135153d297373
z4ee0c8a0e9c7444c5c76c704c237a26d7ca2b98e9665ba3f152793749165ed82eb4f811e78f8fb
z4637451f9e86e32b79fda66ba0b0a5b2b3337c5b27e83ccb48782af0a50309361c5f9607aea3e5
z17cc6278da87c8f850adcc3f260adf6e44cd602a2cd0473c9413277fda58e7739bfd5c89b7676c
z5942d3fb8be8dc6ffa60c28910beb82e4b151e3353bfa73fb18528524c50387f37154de7c46c4c
zca5553dc7b91e82d52d7d52e8360b00b2ede46aff6ac9e0613c734631032193fc04920d9a895d6
ze7a321bf0b58506a5eff6ea621478090598a5c6afd8c1d603352d61f6e983f4f0b61d9949e331a
ze2b43aad341dff9f7d8c821b51c09e58760327fb335d616195293b9497239dbeebfbde92ed8ff5
z5ff19e0dc3b31cb33e684457cf555ca357ed2c6b379064447c94897598c6b243e6a97b5f32c6d2
z268b71661298a93e3360a281e2836e5025946dfa7a9ca796671ca927a990076f3ed46e94bb343b
ze329d457fd658e77aa22ac59d037305a056c351bab2a61bf52cf6657ea1cce25c9b5ac2f0194c5
z83017b58a36b90d3df6e4d337c5467d351b5c8ba95d11fd43bcd2907497fd7717ad361fc1e44a8
z70d88d4fa9bf78ebb77334f73bcebe5b3f489472797727faf7a81d641d7705f0dc4de263e7d69a
zc6adbf7dad26ae8ce2bf0b189cacec4333e1f28cd731cbe4e02a99a3692d44df56daf47dd75931
z36e79a5e6b52dcb953985ac0a4e156203c8909033a2c2e114af7eb2b555f8b5d9777d9f7537858
z841cc590c84acb634fa83f5326b38b2df09cf4e52334ff269487af687201e73230c026533cae37
zbbfa3bb14d8333b050743ce363e0f3c0b2bec1ab3cac467a2930e45ef7eac7a624beaf714ab0cd
z3f25ba5d2309fe79e61226d4619d2b9a094dd3ab415a8f4a418acb0889e8aede7ab4beed197329
ze22e372987158812ca0ea7586a69690730f6a05353d10be75fe67e8b381609931d9ad1e2590daa
z6c6807c0dcd5e7e77cfa09cee0e3afc225da45f905aa929ab40603bd8e49799280ecfb6abeb368
z5a64727b92fd9715e52355daa6129230f0ed7a44ae249eace62cbc5e51d1988fc4520a01ece71f
z166d901079faa4f54d55a9ee20fd6c583b33ba5219cd02695dccbe57c3a9eff6ea7339b563f6b5
z9eae9b4fea000888bc34ef869cd3ef4267b7bebf224103864ae4611e011a6c20f2c20fb98c0391
ze49f7de8ce7ba585d9004a2551756a7c9f91938b014a9d8a5d8c47a204da9e0ff380fa57d32431
z0a78fef3924d4302bdc39c2664cc7dc7df7b1e2bacc7a664b7ea244841554bd4ef1509ed2a91ba
za9ac86af86c543778586ed93e995a8357c756559386fd43c20de12b43befbfdf17ef92f3d9664b
z2ff25cc23b075dc58776a057c5a0195946e9e956bb9c562a83b8dc237bfae204f0ffd32c927891
z60a746ed07735d0b76e80439b75963f50141f4db90d3a01e0c79fb0cb37b6608ccd8529785a7de
za22c37d96ead782eadc3929d9d5b06880e0e42f033d7a87428e669506677f37b6182f198cb3375
z36a7a98c62262cad0af0d163867f85fb76f39af3a5b3a1f56562d168d9145228be4fe8e251ec12
zb1d5cd0fc95d7f1f8c7b53f7f24a5bc21b29b0e2d72aa13add5f5bc38d28745c4f150d7f7a389a
zb2b320e1114d9520a3984475b05cc9a0e24be17e0a32b47c93701801d28376ca891e8a035d922d
zc894a9c6f22575b988693065d4c52fcb1cad01746293dbbcd1557ca343b9d9c572e591c35e0f61
z22ba9cb5ee90aead8a6858dc2bdd71b6f0d024103062c1079d3413344669257d7aaf96176791c5
z093a520fe1aa23e76c691ed2818fa54e2699667cea57900be1a865dcc0a01ef424ff208bfd247e
z980796c3ede8a77098c7137d54de29f69ad20a835ef278a6d4a2d479ee9d18a16be55f4313c274
z30f29a7a4968319c0c911d3964c10cc11b52f06f5f18502a693a995c70feeb78e0612ea10da72e
z5eaf73a171167f60110a3ec56f947061cdd67288a6949ed5e60fa57b0494cb14ba521129cdeed5
zafb027e5796f69fa0fe65f0e5dd6cd500502f576c2a4027bdc8fd9923480805e9d72a6365b2216
z8aedc16c56adf13d1b992e7d7d9e75ef5203a813cce05b9497cf4dbb729b2784e7ea44cacb527c
zc9c91922a7f48e0497f6f6c02b011439d1d899b3ec5bbac9535f9925bcdc5dc6d9d80f1c9a9ef0
ze744628956459e4551a2d013bbddc8495cb0d61c7a8f1eb8a003d5e76b531ed5f81d42721cd679
za6dbe067240155091a2a5125445798d090856cbb53dfec0a3ee21b4543197bfb7b3d0da1ae1173
za1e376c3e559b75163b1a8738891c6ca1457f00d832e086bfcf09d8f3279a53e3604119244d7ad
z7e4dcaef2e534fbf3577c77198fb1cd5ed99713bc9f5426b7459dd2e1b7c63af8c69c839d49a4c
zf424b988c117f365be0f9ec3b5f8052ea4f760dc912def9395721c8338d7bc821576084207ddf6
z3cb92ff179fad2337172f0fff7fcd6e4d019b765bca8a54dd70013eee1b34706b05cb48fc3c20d
z8172c4485f046117efe831b88e35f787a6139883e45dc6fd0149800ac5345fc89d0b8312ca67b6
zbc6a707fd35f6bb36cef124d4e1bbd675f028361f3b9641c8e8df00449436ea38811a361799af2
zc7532b833ea2cc70fb89af53701b28daa05e4287f3add93ba6e48c3018d04dc42788564878feac
z134586ad0bc6cdee3f476d6a5df37737d47e53a0fefcdb543fc7485faaaf20b6e1816495240bc9
z6b86766cb5ead17f702ff3105f5654c67e9cf827994fb8be95053176b4cdd9744050a4053e0f32
z4e679d22b1d150d2a0cd595949ae68164be56da8b155bffed46aa261f62721f2b51101941e3162
z41ca8f995cf36253ca0ac4f833802df68249b81f7813196888e6b400b0c7c41a12dfc60ea02191
z067907b3e6cc0763b301caf82783d17542dc935e7fc186c6d538163ede350c156517d2a5685d9b
z760634c5a1f3cad711e88ad4f168795dd6362221751659cb9a12a18233526715944ca5f55cc3db
zbf6b6f9e55c455fe251c6dd0bb86af1d3538bd7210999c33423ac8c77e904836a771240cffc15b
z8aff3fc351aadc35c8fdbd2621389b1c436d704c6aafefe5e132ce7ae80d0173b3bf08f68498ea
zc40920b543621634d512239ada4446857537179e1a48d63383d05af5b43c27b8ce29140e190d39
z8176d76557deb23379dbdb1eb677cc357163809d802fd49b5822e21f79a909e712594c5bcdf54a
zef2ee2d6786964381edfda1554567a295feb3d332cc5471b9bfe0cabbd19d714bd92c77cf340b7
z73e4d4451f8c842bfc347e9484924917edf2dab1ef5c3e98e8074d2778617d42990f625446e2ef
z8ce0c50a90834689eb5dac62a4d14757782254b2975d18c5b35c7adc527cdc2c84f2f8896d59ff
ze866238fb58238f81c88754033b633285e682f8cf8f9bbde38f429532bfad536305e729d45b20b
ze4e096507dd28274c5e21418c79f45860f0f67919be1b008dbd34e7507c38abe97967ea22a487c
zda6e235440147615670138782c7c43def0a00ea03407fec8ab3874d796daa00d2d55704061d193
z6dffb7ce7b6781beb080360be038666bd2af531a694a6d6974c159842b6fd899ebf93df4404d13
za16d2eb5ed1b4269d170e5dfa4b921cbe18deeeee0d4e36368130e6e93e9fa416309295a92bd31
z8f8e77c04e4f8c788794b50b97880785642b8d63b924501cd10cfb21b4fba1a0e2ae8dec7531d2
za46cf7d47d0761760e96144a46400ab88e49c58a760646c9a58978d5e62e381d1752cc95ffe64d
z351d9ab16660b415b0bd9fa057521cbc35a75c5eb36e36119d05d58aaadcd3eb9993a176815699
zcf222d98adcd7d04d00f1973b5d8041549f4c8eb6fb28881e43434f62e3a34808bcdc60117de9c
z8f09862d3dd4021ddfe92fc8e6656230e406b96aaccba1e192c33dc1c01dacc2ae8d362b5d3e9d
z3648debe3c5cfced75e318be3dd4f1f080463abddfae66a0289e4dffa6b179dafcf6cdde240daa
z1d27aa17b1dd8247f92ecd48f52a9f2635b96f94027f63e1e6e098f7605e80409ef9f547cc6021
z7a7bed7e18b72a882bae159ccb622ff569de3549352dce32349badbb315496631c7c5d6010d849
z15705487188331dcdfafc5cda60a8ee8ddb18069c0a4fbba2b67075edf6f83f3e65a554c600002
zc5fcd84d11c72a72a595353887759272f4d75e8f015b96f4e4b6e972dd536bb26dc300405cfa9b
z0c16107a4151a6414f2cd70d9386f931c52d7399f3e1429f058125f0a3bb0b38f90fa09b06248c
z82191319ee34624c78e5d842736cf1f3638f224becbe28f3c0b05b65d194c135b0d3a2a64db292
zec76930272e7602fc41e5a0ec67134fff467b53f3ae7d0336c9dbab13bc6ed35d8ee0fa65ec51b
z8c030ccf9e22356f106021fd927b5004b78d1741d39f98d9e64d4f4d93fdec4e86a7a37f48e8aa
z308d3ad9c5e0426733ac37224b619ac7009ddb3d5d67cf0005193c3ca8d32d4490f67d5ec9c3df
z2be2bdde1761ae6971a42e357a5af7aa3bc6d99e3020f675f92ca2f55f4be8a9ab78abcd6faa5a
z08123732e463ffdee6cbd211aff0eb54498dff9dbbc516912b4548e22ed6bd5e2fe0bed8535217
zf09944f27312745423e8714fca92c78e5b98bcd5cbe5d787d9bb2d56e1dde29eed9ca8c06bf5a5
z870641e2b48c3b3e95fff97f6b21a9b9983939279c5f9b2c32a174978f5585a15f54144df6485d
z4378d3d41eac52f3bd93218ca8375d85de8950fb7d12a2975a51c111ba6c0ee40000f67a1db223
zd005190b0a13f3b455ab8b7d9f1a489e3be02095f2d4f0962575cd48358d3c00a86321be0b13dd
za5339650b5f1f688834db7d4cfc5924543dea4cfed484bdcc180aef7bdb91990b8e087c338ba0a
zafdba7ac23240680d76b571d9a21ebdd74db00c59fb7b9f1ce53cf984094d47344ec38092fb887
z0864342d22a0e42186efd8819b218d1882ca0598a15e7f8506b929dff8eeff49dc4a7575bb7fe9
z2ade673fc49d2f8f4cbcd32aac14a870bfa97bcbd2df6e91e209fbfc198f4cdfcf1a1c416efdfb
z063152944f619749b6138e55a7b9743cc937431ae67b16e4ce0af9fec3af1b1d1b12eb362514d0
z469187772d9b1c4d9b43ee6df4c10f32019197af6a567d4d72a59ace17efd5957e1a6d93e6ac0c
z3e44f6ea33ad342ec1d1836003ba550f6c53052a58f4c69355b78ac454fb7bc65c6fd48a30c1b2
z58586899307ee1236b397446ff35e9a6bfff0fa77bed774d75967a7d1375aa5065f38c131a389e
z4aa24e263cd6c2fcd531f8735e756646932393bf4c60bb4e61fce00b0de9d08089d7bc09911436
z4457ebf1ef4d7f63e8350177ffd7c90f5d50a2dfbd26ee64f5e81ee14e167dc58da0209572e9bc
z083aefe754b8d9bbab6b11af7f013da2d17b656ba2b463beb35a05c836dbb44743910178ed5183
z1e92f95b85373b29cd90e52bc8cea785ad5de1b60fa8cb92c5ab83988079591ab8b351dbf60ea7
z2d2a4a0190ce7b5c63ff8073ea934e8a64fb2118ec825b0b1c34df25debf1f2245eefb7d0bada3
zb0810579a462d2b75a44047ae2cbfac78cf7119af6a2fd0e13001159e001ee3288a7576d66775f
zcb6225216fabe1d33c0927f703229dbbe4fce6181f4e687d29ba27896aefc471f1fc97338f1b1b
z93d5950b80f3b5af210270d3327b765ab753c8fd615f1733ae49d297a95ce85c2e2c37217baaf0
z60aedb2a8b1daf5527d97e8a36c9af4af7248c432e51697b136cd3947cfd786e54eb800c674c38
zc6181bf703b1a4fb6c71e440143d1d24e416a2f44a3537d07b002e957c2fbd578624211becb58f
zccda9e7f0aac6be4bb7703b30cb5bce630f1edb985b39baf602ce8529bb77d093dd9a51c43a8bf
ze6c983396ad745440dcde102753c53e93bca176c2e96933840527d4a719692ef2cf4d70c207a67
zd1e25ce7c99af6e8fc0457ec9a61d0e84e82831be45a3a4a437832f3ce4994caa5803d5e16ded6
ze896e2944ce903fa597ff7925f1752f3ad668952a8757fdb54e86c39446a69563b9e55652b1192
ze593933af06c67f021acd90a0b2fdcc974b914119f7dfd18ae44d2d76f94cc612cd3e30b5cf0c7
zc78dce2069ebab381661ec0a8cedb7f6494631bfb683273a8b4e8d22e8d8093a4a3494b24c313c
z43988ac1c8c7a3318da76478aa532758f3066d71c427f22d86a1c545a61c1f5e3893283c90620e
z60d7a1ad32731f74d0dd4d36754f6431f9708d98e4a2fb23d8f0727827d028134219f753efbdd1
zbc44a322a434f9a5a814fc7c93cf2297b86b845bff44aae04353fc27420a07a72ef57502da02cd
zb7feca3ef5e325fa6a37a24ac69bdc9c81fc3c68c17557f2799197a4160957c5279a093b63a537
zdd71e4d5f35fde1519da27acc1a8274a622efda903a3ab556944c62e11a893f8c673018733cb20
z46078aa944fc4713a38bf1c69ed83afb66ae2ab4797216394fe518911bfaac392563d0b6ce963c
ze92177c64ba14a2803592a862c960c6a473932f54615f6c4867d248ec76ff3414b62051240f50a
z1c916ab910f6fc5c019c28fad90ffcce01ed69389b23de0cd135bcf19e6fffed8e70cde89e6e0d
z9fe84ad5ef6cc1dce7cf6191c21297ad5a145e22573d1faa291b8c0676319dc06e3b4c6ddee079
z08615ed641ac7bc4b6fb67f309f4aac210bbaf7088a9016405b0a21f6a1d8c6c1d293d259632fb
z7fe49bc60d1bda2b8f2794c18b326f50c33ea28249f28c0916e801ee21ad8c2251298116dda435
za30d68996dead7e30887ececb53f82fdebb503fe2f30cc581a2b848572b6878def8d37a4570b6d
zdbfdd3581137ead4d4113f09d70777c84207b2042bbbf4adde3da03d6af2058d130514d2ca4792
z73fb4044ce11f6c8978c908a4ea9a95876500c68c04cfb3ef9d152b585ee3b55bd43541bf9457e
za68f7b2d3e5c8b04db265488d7e28d1cdacafc6076629f4416224b22a58ee7d50f86aa821f8299
z4a066cfa1ca04ffa180e9511ac7abd92b2aaf96fb96758ff41f13012c50157eb0dcd85c36fbe13
z370bb38d7b5e9ada2a569a98371656e72198dfb00d5616942e5ab3aa331b39b91a43344d077ada
z7e22d9ad9958272e93487389795c850c25d5d25816397cf570f349d77c1d81c863d6179e66ba2e
z95d689095d8712cddb372915f4776ef90c6bd29d936805519801e2170abfc5c5f4b416088f54f1
z100f377d83e80688dbb911d37ae939333b5004f02c3ff2f0537662cb56260b036db6d258a9840c
ze7eded2daec46f9173cac90fb36a1a81975e68fc4162238c61adeb167afb1f8da4812f7dcf38ea
zd8905f8d547fc54e1e723809ce7732d91aa15bab88f27dc5a4780f588acb4edb5f7ef935797fe5
zf415b7132df23e669ee449a315dc744ba08df51795cfa9e1fcf8a9e766a9ae94d2e953ed4c643f
z2eb199c61ed5fb2d75f9819cee625a10e89ee28e30f369ca45601974519bcad746661a75982c69
z1beced2d4768d5491353add5f55f3057cb653f3be17dacd74f1330765a38e685f4b46d405f7381
zf6852cb3b4031804baedee50e61889af1469e4fa19196b5947df4ce73f7f5fdb43a1dc2c8475e9
z51c2222f1f5eebc4fd6e444919870dfb5d8fb3cb3355006745021eb9728841693e10268e23176e
z40922923af034b6d95e103a2e1fb4ddfd82a611b9e762dce0e653d4e2491a204a59ca9b2a35231
zc3525738e8bdc854d39c45df9467b8bcf895a580f415bf6bb31b4b0d7411591a0c8924dd53e043
z266074bc1c2324c27f7552e7a729c0717f00087a9f0097359a0639270c125b0a8f0caa0004c981
z476b75a36c73d4bf8a95edbfce766decc38f6f8611f26a53c227a55c48403333dc2264277a14a8
z6f2f3371346354f9fd42ad417ec2e27fdb701208a576e84978b060e7bcb0a34672be24c6dbdcbd
z1ba35c4e7b5ddbb88954e808f9fe034fe4726436cc02e0ce444a09d010be8aa33fda224146145b
z6edd7ca19907da103cea576ba86ee205b94266d80a9c2474200de49b034c90185fea46fd412861
z694565dbbb22274903eac34a748cc0966a20859e4cccd40e6359629edcb3ed60a5708255847fb6
z82424b4b1b9c757ef6f0a8dd5aebddee80c11d8735775fe8afb285c53b1ff818e5e0e5fdce838b
z3b1a28ada8b15ac3b54d48b0b30a9e93b547549d0c0096f80fc19393b7f8a5a828616c968d361f
z5652e37b745db6f380664cad4a551631ca5891e9e8bce33f4a229c7a4a62d66a8690fb307424d6
z8511208c884e77ea968fa04d7ca101debba0d39e61d062a8475c2f67b61f940d57272c1291bf63
zbe586249970d3b917b497cd2df2aae630f88a78550c91677b4556eed174119800c135a47d47b39
zc390f9e0d95bd33a2b02521740bdbd21da94951120f2c36f852f34b36edb3721eaf010c95acb4e
zad39b82c9d6896e6fc710e3ad75bfe3279d1d86a724937c2072df788ac88e1db8a94c92c0a0f43
zd2ddf447b70c98249ec409bdf28fb14ee7be804ffb9c9058a3efa110f3c4d97b86de210a581fb9
z7e8b50c576ca90e6d395314f06069824f0a5496d87abdb3c0454d68869f529363bce30ec6ded47
z93b5a70ad135165e5dd6d518073c160a6791320fdcf8ddd72280a073a74512ea8d37deabb6f1e4
z98ea7411bc9dcb1ddc54da7a71d14b1e47c17428d24153fa7005c9ba6592a41ac0a498019511f2
z84e5b236608cbd1b7a0d7df2dffde9490a21c2fd70b92f7f8dd3650cd813504d2ff71ece41a84a
z18ae89228a753aa930506a94832b18ac221173a6f8e3df4c9a8ced56568d407a702ef23c80380b
za6c2469a5f500aa0dd2b6441fed5e856b049fcf70d90f8c10685aae6ac1beffd059dd9cf87518e
zc59853a728d7d263e42961c81abd46db3526106ce0d840699e2ed99f2b56b22ef59f5b0a209f2f
z1d8e78261500b4d917a7fc089faef7d7773568f7ffec1bd2289fe77b5ba9e8a77b2a3435faa9b8
zd84eea8f20fed8c2b77f26f76a88a63100e68ac592584a374c76412399ed9aef14928fc520f775
zc91a6fa0ddece0bc000869311c181a310bf3d41430f198b17bbe6b5b25a6b230d67f8d60cf64b0
zd00c182dc36b2b74109c1fd0b4c010cdad83b0256a3f517c9d906a8b33b47cec991a2d60f83cac
z5227d36a9fc631398e49a9743a4a46cd97c9a327143a1ea8c41a5b584a3d3d943f44fa616df24f
zac26417d8d36bf82ca85774774f89b8bac6b207917ef68c28af320b02f3e5666460bdb15a22f37
z81add33119c1e83c9d017d6c9cf5f53bbf7d572f5ecc9288acf76e530debe92c2ff1a7fd5d8ffb
zd9025ad36c3c2210fd3dee4c7107d097c5a27b26513c3b130a3914f0dbe44071feb1a7079d0445
zae1d12eece3a5e6ef49045ef9214cb14a06b1d393b051d6194684b4eec9f3c898a566ce6a3a11c
z30e870dd4684a6fe8c7394b96628295fb88e3b3b672b46abe946abd8ce03e9d6b568cd5b6b56df
zff7c8bbb5326fa34b82d6b6fbaa9ccd7b10a6df4ed49f7eb150f6dac62dfc9206b85e6bd13acaf
z8072a15798d22b60c048885850417148c857b9f443d83e70445dfef4babf9ac9ef785285b8ae0f
z56d00efdc23d3bb20de3248774d44f5af213630236d9fb1bcecf007a34b11f1dc0a5994ecabddf
z3de6e321198fa18d2c9c49ac71b57b629ec1b15c9f065aa3238ed69b936d45ef120e540435c6f4
ze6b47b8a5559be54e6eb4e4d903045426825481d131fe698f96ebfbb428266885df05478633cf2
zf030a6b2e8898a5416f84c8bdcc3298965f3be9c78295aadf2d5704300e4e1142a8499cb87793c
ze9edb0e459c8154e07b60650e44f9a6e77c27f1fdaa8110d92a0dfd482a4c363f24cb782796e17
ze931ad8d163d55ffc057cee17386f1cffd13da8aaa24d297f363c5455ed67838f3d7e963af3c76
ze96945e194b517d77196f8d4fac4541741d8e6804c12482ee38582325a991095e4cdd7f6ec9306
z2608512bfa13685a24f6501863e24a9060c5be98e209a936ad0d3143d574135c3ed53a27e76ac3
z2001893b21d14a5dc02aa75f6470869ad083e14ba5276e8a91f826e9c21ad6f6e2ac360f2baade
zfc5105af717814945990c6339728cf0f80b87715d7f6d959910dc3f71dd02a1f2ea2f4b4135757
z9f31338f4a9185cf0762a13f022661c588ed7ac68085b17a024d11643c87ba92b06eef9397a358
z3a753537488ab01362140123bca6c6a52d6e11e903de1b9e8011bc95bfd348a01650123e3f6801
z60324be80614674bc9024ec13965d299b0880af41692f9b096a02838c4e293779c1897d9b30fa7
z60456574367f353640151dce2c3bd35aaaa5397178ad1aeb47e330f051674a9113f1f414b163f5
z33c3b3e2b242287b760bea31fbc228f6822fcb710995f52244a129d9fc8e5d7bcc51036abe783c
z9053c3bc6a565ce3416a200ccf8a7042079984c57c69b5e211bfc4e2f45d3c333df0413abe38fe
zc0bfaf17c1a97fa6eaf8b418e323ff0bc34405d724deb76aa8c60f81994f58f9da4be1957e9f3f
zaebc3c0b9380a2ec5453fcc1fa488e75013245b0ea1b52263cdab27740a6d6a1b766b7d4d63038
zdf8e07226f389e3188e245457cadef3edcb8bc98e7589b40bdf82c93d308f7d6085e089bec8c15
z1e4e85371ca343f951a8b37868edae5db1e417a6cb81d4326eb29ac8a5d169166ca61207887613
zc62f000fd7d71b434a33c7e5fcd4d0a7684beac238d064b1e5cdfcfa12e4f1a4ca5bb1f12a182a
z7d7a82683fe0567875fa59da71b0295911ba958dd3e0933834e53282d92dd140180f8f3603de07
z89d67090028a709eb4c35293a8c2c87bd328c8fee74386c6af9d94939349f844e23027f3226aa6
ze4f9310f99cd5f23d7865d46a4560acad94abe8cdf256a2ef39441aa3fba9f58a8ed446cb795f1
ze0918e085005da40c9a7bea83897fa7d96254eb90d6fbc5c895d42d3f75cb991c0346521319ccf
ze67ed8f01845cd01dc53105163ca262ae8bc680aeed5c7648d09e10baa3c4fbcd4e9e655bdc07b
zf7ee594a75b9ceb148ad1fe3046ca7bcdcdfefbc25bd4304ff448f1144416e4014c600347288f1
z095fe6ed4a397f3455fce8851b7dbd9f170c2129b23a217d2f298e08e8d7da3e8844cf511bb84f
z3787a6407bfc65c6ccb14903052cbad9e11ef213560a8df379a56786d076a63cc7ae4f82aa0213
z3450bceae8fc44edb1bf9e0ed3b25aeb6cc7b4fd24efd558fbfaa334228deac780ee32d67528de
z53368fef4a959a156e605f86d5ad631f8ce48921d801c69ec3ec539bcb8230cb050b9552609d9e
z8618f68d2c95724d7cae04c5a0d4e4c862ac90bc873f2a00ade820556ec5884eea12dec3aa1e23
z08fc0f66d162b4f660c5101d38c27fc93bdbdeff409b7bd2e0ff93eeaa292f8888c71cbfd2c234
zf3f46886039844706c21595566aecf40e4ba1041ca73f1dd99389f04f21ce4ffce06f7a285154d
ze75e502155ec7e049b019d5529494c3e7d93df44606f39cdb43448e51ce8ee3bdaffb72ad27c46
zf2c3df2fa75e968d466e674cd4b4823a721c5b626a3d29bd520d26b1c9d619c814254261fa79cf
zafb5227937dee19fd1b4cd935f3f0c84c806c906685e90aee47fe48c8c06e8e575775feddc54f9
z06819f5c5d7cd090fc65ff369207b05ae0236a441c5fcf25c8c4302a4a9351bbe703cce3cfe193
z55c1c2e96151a7e631536ce04fca694297cf3e9fbe5301403e042d4ec3f2c6321383552fad1437
z5a62cf271c8d664f626d006fd9ae2523d5733887bee1cffb3ec2e31addcc39839eaa516a12fb92
z3c0278199079ce22f1326824087bd607fce30dcc109c6e8a52d63b7995e50a2af343ed99d2ea34
z387150cafd4584e2391c7ce4e6aefe6e3922a6014193c87fa4372c94d18d0841d66de71746808d
ze66881406b0046167f6ac63546723a1ae37d7fae88b5eb71a0deb2f1f74511af4a2c0dcaf02413
za4faff638e56dd319c1e890048cd3bf63e4aa65afe5a062e717c9b6dae0d77af387113ce5a8902
zc7ea04c9fae2b20df3ab769cd2ab5f781ce6ce733f34c2dd9e01aa0e15a033fff224dd0810a5cd
z53cf71fa65c4ac83c0e4e64ac67127ade31b5aaf9c16edad4f0ad65d0a8e64bdb0fcac3a905342
ze7d22975f9a6b50bcd534d2b574431640cb435d811135638beab31a37c9d93e867ff82e6e50b33
z82556f99b36a7e8793e95ab7e292a2af44997a239483cb76476acf64781f12b4f43c7d80625f13
za55cf41fd45d18c6a003db14373b53c95694e35a8037a5d92e238e15aed7b4b1aa3bf1455dabce
zfe76bf71d9adbb9855a1143aa0201ea2993ba464dcef048e45855909843788d4379a87f2110c3f
ze39a8272173524106017393faa70aec2f861b963a6c49fd940f1575c255e7eee963a31dbd66ba4
zf3b790328b565914d1410acf552121f82169de6bb568a56c60cfa8be582a23693ce3abea0381e4
za4783b9aea5915352ce66ba4b6fc73825e4f74a002f4edec99e712d9524969f18a5f104cf23cb0
zc2021fab98b7dafb53d8d743abbe15661dfaef1f0005d54abd5ea111aad0ab6a2054297b85cf93
z2f2577f6a1afeeeac29ddc807b4a41a69186e0f7b5126c711b74841511973d4ddecfe6bab8ab7b
z009e29890409587e78b343c2e34e277e7bde9240c5e22eb9c7f32488d9a5ac2bbebeacf0f8fda9
z30091c00ba0110a4b668a58335a1273f7da8e0c4e916f62793c03d6a57bdccf34563d93ebad2a7
zb85d57fe0c2d925581596b174db2972d38281013f78a8c624056fe9a77171e027c3d934822ef3c
z1076feb5712f1379138de375ef8ff399b6cb78838f27d97eff27b4a28c99c42abd5bd61e4f5b3f
z027202c6c77b6bc371d8a1ffdde74b136e1710738ac3b7c546986b5a06b2564b3ac758f06bbed1
zf66626a2cab3cf1aee73820a7b044aaef2acce5af4db8d3ec1bba969ee3c7c06497b1973d733d1
z21389359a91d0ced2e02f99425558b9acf70ad81d4800dd4b5b89a1e92a9d78b4e66549433e706
z40f10a65e6fa1d1ea3818ed9ee0d597b10ee43781ea6ad33abba7f8eefa3ba92693de1efa2ef99
z290d6f4c64f0c273f4441a9a24dce0bdfda76144615d34a17774efd909e9af7ca4ea147787fd98
z1cc35faa7c8e247dd35908d43105b65ca89e9618edbd370e45df3c19699aea758cf5564cc36309
z62c36df29ff0273fb2c55b1ecdd0e5dcf1ecb8ee36a157c56e533896fa73897e314a539af00c7b
ze245aa33009665e2f0f2496cd28cbc04282faf38746fe77f2451dedd49c3dff5f5b194e03cb97c
zd921820e39e88b0ed1654e68220e5011a8ddcda0ec5da610c39e904e0e81ed06b15d83596d41e3
z51abcc880cdfdd66d8af3ba53bc21928016c20aa79aa612e14f7247e499ca0d9f0f9dcf216ab0a
z091cbddd11874cc45a03309f49290a82cb6459d005630bbe686b1a75b4ffa5d6ccce2ec014dc2c
zdd832506d39c37366f0a7988797050e3d9ee5ab8349562624d4c699da74139ad60eb81cefd2947
z30b1d5689ca1d0a98d5250c5255cf85f8bad986fe1eb69ea6d0edf3dc3408ea0046698089b17ca
z11107be2821116734314433e6987722eadfd26710abcd80903588d354175e8ac0602ffc8335588
z2af8a1d76ede1078ca9207fb0b4e6b226b4688ad8302b1f2f501d829b445d9d4468182b415815d
z1c513d6ce11a581b9c90d2355a5112523a0e0bf28ac9d180e140c8a1251ef9a531fad7d0673bd9
z7f011ccb274b26507168bfab401dba2db2dde7a1e4e559ffba78afb5aad4cf6d9e6b9124d801cf
z97bb019657c868ef1e1d050fd47fedb96597d49faf04de66d96c0957a5f7d5526c850af91da9e7
z78a3312b9e5b6f0756aff2de3fde46e5810bd6b68edd806adad5eba23e383cf2645883c0ef4ac3
za517801ece17d04c86bf9434fdc7d1a34822aee59c2c6bbf11e6dd0878b4bc32d4f7632b43cb07
z8c52a133531e3e24b2d5a7e78f028227c97db4871fdce1e4ffd0a53b8c91bb327cea7e0511f9ac
zff1c55a531f7c70bb2464c803be689f22dc8a680724103c5706f9be28058508e41ea271b86fa85
z26755dfa3fbeb89d27cb222731fcbe004957f3e460cda342330e2edafd194e45e32fe5bfd62158
za4ceebde1687612c9fe26a217f413684eadefd4e64726cb2e1907a1fe9ec2420764ad27d639eb9
ze248435ea714706997d1bbacd9ec676f71a4bcd59d2e05a28832b486ed1e284bd15927e807387a
z8a3885510bf1c103651ba4f830e6587eb220fbbfddd96b5d1219c051e08eb1fd666011b58df364
z37bf890e7bdeb119c9365650140b6b651571b02f374453d19f031c6b33a7d1c9e1235ec3a552c6
zcc2f50979d6360ba1166557f8fab1d162032a8ec6e7188f42a9e2f7fab9e15deeaf76bedecc45a
z83eba421530dfed568831bdbb5d3ed481c376b81fb0877d0d04f1f4c124018316ddfe130c6d982
zcba14b612a20ae5deb5d3335e662b6904f5cb372167329a921dd4bb83b3fd3198c0530718531f1
zaf56151ab444982d4def07494fac6252aba70384cb44737cdf19bcad1f5957de9f0df8b930b135
zc4388ac8146ec84a01ba8fbd4c3946a4f253f738798dd633a98ab928704728b9e62b166b73cb20
zcfa0cdeb993833fb415058a5f8e4f35f2d69b470630f749aa260308b59f38f0f1aa1026055649b
zf880724261bb4c7ceb84b2701fcd0bd6340fa1e921d8390db38afa47fa8b1785634d2b3de6e7e5
zf20b33d8da6e771527dfc17e38ad2a2214d37b26fba49636eeefe4182b3becb7ca944ea278ccb8
zfd077f124533c24952fc59ce3554fa7845f329384b0fa2b07f703242133aafc496d65901b4a81c
z59bf2ef22412e903475dbe3e0e6fd017b6fd019efde8e712ab58ba804ad845407c49777eec0ea6
ze4e33f8754d6abfa3e8dd67533fbde6232036349373b0ba74d5248e2a8d4b92624395ed254b5d4
zf4b1a3edbb2814c6df1b4fcb816338f1a4adb1466a1da4b3c02c7441aff9ed094fb6d6f4b05cd8
zcb91f2a847a81626bd6a98685bf1f3f443289cacc03691fd3b8df39e32206103d9764f042784e4
z030075173d9cb3133cf803b7f80f49a0699a3d96e32aad0791205947f1ec969bce4d84148ef701
z8ed2002e3dde81142b62e04097f060a88ad3f1967df0d1f020d06631a05401d612d51d924612f0
zb5a06f2122f9866ff70667f0d098afc3a39ef2cd8a9b8afed62ce4b847b3bbf6959a60f7275bcd
z2ba3d2ea30a1b13e4a6527ab4591a9ed4d0242e2ffd7a1974d3364b06c6effc0e9ad4805d66ff2
ze92c1366ac17b9472605177a0b7934980fa0d0cb7d92bd090c5071507e7d1ed8af04498270c7eb
z64d5a56f56e12cb24019dd346a6722411b022e7328108070c5670fc753b531e72fbf0d535c1811
z414f8ac124b45d3991d0c0a9c713eaec9c5f75cea0befb9a8d1a40d3a99701e062512df5a39fb7
z54058fe88550de25d0079aad8ce8e2069237fb0dce0aa1ccdbf110f86a51df35c5ced986b5851f
ze2a43f381af933ce8ef88f983a243c14d59d2eaa3b2ce51cd0996c426cc9a304152374318bd0bc
z286327f248c1650fc2d3bcf30cfd15a27f36f2b2273dec203f22752b2056d23fd48a5a40ee6dc4
z75e9c2c6bd989ccda3e7cc9add58ce5ef79366acb4cc72cbf99fe554eca370568d176d44e47e0e
z89d329a388680ddcddc57eae18f76d726ac8e9e750d3967b08acdfb412e92db1f5afd0ec63435e
z448588f35923ab957a0cd15d13a094feae994987e12cd056ec203329a0fa342a85e2605a1df4ec
zd32537b87198fc5907955b986e1e3c2e020e4e3705f8bc19b889b01dd29a75f6539c320d128d00
z94ecdc20d5fb41b3ae62496e26854746ec1cec5fb14453c04f1b2507aa894817c20e45e771edcc
z3026488f57972a8e7234510007201ad73b856bc6cd92dcda4d492e3bb2c5d528891e6f09860737
z090aabb32b0adbf16e623bdc102848d523defa85462d7f15bfe4259c6d02978f4f9b10fd00120a
zb75b78538c4e728b986935da94bbd3598a25136b5620cddcd0e57d13aca5ad859d0b24fc7029bc
z50c52ba604063b63a548475ab57a7b6b60c13f81429bc08189c1609ac3f88b0a74b5ea7536112f
z75ba10e6e9046c607aa540dfb402fe115887377f98018e92ff63a612288971b437f1d139f65d1a
zba5a277e94c63b6f77116dba83b5e7d1b0f2b13a4afe5d19e952690b788b716a657292f25c4de6
z6d08e3f33307a37fe8e9d01bdffaaec38a67887071158c7bfa0179ce964dfec912ed5e52b491ea
z7450b586aca485c1e42fa85a8e2707b7901d07dbf6a337fe18a229e82dba0c075d253449d85a10
z871197e5841971e62abb5435832bed4a3e329defd3855fb6137b68aecf70168c3eeffe1add0d46
zc65d2ca980ae79b929277b2a93148782645d1ca59fc6ea32d937b4427017428f93dad05bd6ad00
z641c53dd1ee4acc0ac518e4c0efb23bd70a0fe599797d1a859394d2f91017d73c7b2d0326a085d
z04414c160d361d702ac81ed9b5412d01f77938894c7a266cfa8363eaa2fab995d2fced3ea38421
z1c2e6c2e32806970fbd8fd7d3569e1e5517e58c18c3f77a81f9314165f3a5101fad3fd9347aff0
z5e51a30a210211f4ce0426802966911408259ad18600a0e9bdcdcd0f4ca3a0087eb43750c3ce73
z1fdbc90db0c4620087e1ebcf312f584a5d1ebd7df85e347ff8f6120b44c4e19b19ba31be4eb360
z74a2a324bf5dfd1b89f86c7153c70ebf6230321b76dc8a879a6058b79eb5de90eb5e1ab718087e
z2430318a10d5e36b59ec547a965a3173bd1616034d36d3e15d63ced84ec3eb7b4be09270c9e8d8
za3b1a754d421b452f1ec358ebfac0239dca0b2cd95901e421495626fb1e12a2db3debe06f4f769
z1dbea63f835649d178cbc3cf9e1af304f648156b13663c32f72364c3a4d4665f2e30f6af9fb571
zfe439916034ce9eb3141434a622765b525ebf609370559068b29dfc05fe4e51ad78f23ef50ac92
z69b6761f1dc17e7233330da18027633a015868d8bde73f190a2a5cb2b6d44d33a97ae236d58290
z457414b2edd8a3a517cfb98a8915541f60f6431e5d6eea7512bb190ff3015889a81c7447bfd90b
ze8fb64eb61012e70f01c8aad2d4f70b4a643fd573c73e3483d9409838f149298a979801fb194d7
zcbcfe40b653b4db408f233d1ac1bb72b0a0c28467cb27387a5107a739fe49f12875d73c96c7fdf
z926028aa7a61d57d887a8e25ea71ce58ba9ceda980af2ca9b5f3f3b5da5bbd064763d6f44af91d
zdbcc465b222e246d7a54ab283a1b84a09813a1b6a1981114c520a49f4410adff85b7a8f4cac9a7
z1d51e6a021f06608baca066d5b8a8c2e0a93600b8d0898beed9515083b810298df222df26cd604
z6424aac644d485695eb3b2196f9a5be47b08a7453d002d1cccf0d7529626708ee5e2b1c0b48289
z7d881672be59a1f223f27583303a070b766b86cd1275223845e9ebe07418b1280557667162fda3
ze7d5175df0f2e396e220a08f08cb6c1f6028409320da353e5e6542fbb1fb0d778e27a84cf747b4
z4a53b4dd77f92e767b408396dfb060c0182bdde57f74e8c0193b86cea754dc25e26c3f4479ef05
z576390c083cc1ccc35acc6b5c99ba9beb3afae5a51dafd4690606a6905ab44e04eb932d701c320
z8b5359d4549bbb61a4a717c6c9850f57c499cb6969daeae46dfb55d6a0081822e1a370cd32aa63
z7fd5eb8f8feea8e486c7ee7d1f40416dc796fec9904b643030e9827a6eab5e6e97d58f27e682e4
zda93c8e74e40aab46a0487fff98314afd0c54e0c5ac7521f2dbc22825db2c2db263b0eed7b2aff
z5930bf72db4dfb9bf4f898c5c408c215d9825b4fe77be004c9bea55b79e14b22edbd839df38cb4
z2ab6fd79f451794a5d248b14bbfe9813aae4ac9a77bc6400e7f217f83f13a927b22c55caee0b3b
zbfe3d609583724ddf57f1d2b286e33568bc6552094ae31293256d9980484bc823709d269a51439
zffd373c4d6e441febcdd08650667e176c3f9034f6286de0c9ed449893895a4634994b46e822958
z3948c6aa1821bc6d8b7565626333743dcbd4b14a933d9ad3b1f782442896ed1739e8007dcf288f
zc8005fe1fe7d57cc649bbb696cbf92a6ddd3964b7bfc9ea98a4807899e196632bfe5cb45ca6f5b
zb49bbfcecc970f33b80e6ab39a30a5b44cf8354227dbae56a9dc20c5746a7b9a88831fc9ccc664
zd5df73edc5d930c083e053d67e24b86544efa308afd33e80f407f04774f926fdeca1df42e9cc22
z8322451e89315c70f9be6024c44b8730f9b239d319f3731daf4fa5007157fe6e9e433e4c7227d9
ze252da7449212a57d671b8cfc66e61c1934373941babd262440e0f8bc43517902bc965abdb9e6f
z39f11dc5bdeb36e6b64c19700253d0deea31bf2fabfa9b6362930aca9c3a80104f50a27ef1165d
z9c0dbb69bd0c1f0c5b2b2e6c46fcd353d52edf0603bbe6c62b3576ac083f102f79b12437c1d13d
z8e37ebfb53f274737d75f5d89a90acbcd30e0567e58368bd74ef0fc2ed39f335b96dc1d2dd86c7
z40d46313bc6a1bb8db8cfb79a69f3f610e6764121f2b4e86c5e97ea4a77c7ac0d399adb5cf9fd4
z1847bb66dde6f4198bd94ecc62ba028623e2b900aefdd4e046728be6b3297f9ff03a6fbeb77c7c
zea6870bb052c3e03d1fd844c7d0e5fa6c0438479ef3afc10294cb3664020019ba9a7608802df4f
z239018f27cf58a788ad74cd761e165248b840219901d50ab84f0fe13efe3575f05cc1896adf404
zfc93807e96cc1c78cff2e12064d77150dedb73398bffab048dd2cfc8faa8728e0e82ec55a963c1
z4179430ddcf405048d0bb8f4768dbdcb0685c8666d6ede99465fd3b1330275c6bb4ee495d1fcf1
z47301cca84d59d52539198066a3d5a19e647cd017c584921ad35fec74bc906cb4df0ca0cf67968
zf4c46e0f77a9ecaa66f237d752247d0d7137ce7354fc6dadc211cb4a143aa92d58804ea37f6802
zc6e997c4e8cf7e42c5448823edd86ea710e3ae5fd95c94e425bd79ad92ebc65be9502b1ac7af3b
zc08437f1d420831716786964c3cdf650c789c8ff0075a59fd37678885895d3988dabab249a1977
zc6cbd18f8c9cef7ff39506b6c6828ae1fdc2ba4aae0ffe1e06b79cff72900a6a1a396af67f3b79
z60f43ed0ce1542809876cf290211e0d2d498104796fa3d5739e4a68ddbe76a185898cf4eac1847
zc705ff3438a3cad4ad8ea4b37c2d8e14d5c5033be05821e7091c8d396cfe55bd0a7533632632c0
zbaa3cb37fe246cb7dfa72f40c3259e0704f5aa81e342cac6669604738cfe2139d4500bd1fe734f
zca868c0fb47f61743149b8bdcce1030f53b7897a0509aadc85569b1e0c66cf404ba0dcd0fef719
za182d299055d67d54da8ba9b0f8a0273d12de3e484dcaf5134d04f5cdd72577ecedce0567219ec
zee85b25ee8ac24dbaa9d301dc105b3d156da205758bb4f03de67ba89a7de09ac3293c81953c4ea
zbf5a3b7127ca1cae5c4ec75a923db5119427eacf4466e84fe3553a70e2177b58150de88580697f
ze4440e02aec28ee8ff97c8e6ce1af1469c9840a767c67f61dcd4e00ab8da8c2abb223e52eb1030
z239d43933904b2e939346bd4233def783e56b10b7bf09e7b0e3887ba68f33d2b29674c99639c01
z3dd6f0a28271d3b11b664727a9148b3e85d1f1d9f539e59a8dad3f87e37baff88443cdd45efdfb
zf061aa6669ee5684dc7172a7f9f06ba557b3b82b687553e13e66462eeb2a8c6840478a67de0a71
z0a6533a79eceac4b8efc78a448723300c4c63de1e1fd0399176c9a9bcffa1578dc719701c72389
zf709306971b5434adf08c675d1efe1ec90df360061cae9ebb2185da85454c28381faf830f29820
z15838fd5433caaae8e9d74ced376a6597ea5e6474524133f67143e8d10e64b6320312c250bf437
zaad93a99bce2626ed22c3ef101fbe6e9211edaca4234879c05c2911f0c792cf0e2453701c65dda
z87f7a7fb76037db2ba7187ff0ff46f2bed55fc55781ed2ab9ecb3e4229f12b033f72a3b98d19d8
za780ed9e998d5d5036ae7f02073d2f3cad2aec0309ad56918a6ceeda7eb108eaa262c68f16a52b
ze5bd60891a7c1c49cfad22b3eb8e782b3535312b1776e34b5963ef82c0371855512644eb0fad49
za6899ce02c8dfbc6f8c89ffd00d58836ff295a118fb90b9495e750fea8cb84af490fe22ab917ab
z235b361d0452d6f3320ffcdbe6384ef5619059b6b628a6d96487a9fccbaccfd3bb0e8023be6c0c
z0578e45dc87b484938bad06c98bc0bb24c547b76b683c8d4fb97543c00c126abe9b33086335306
z8ab7b951f6923b67ecbbc6f49bb3e7226be014f5533fd16eb3db2784681d04185fd56ab6841807
zb2732ef14225463d2362ba92b3f8e98e3151959add75fd5fb9bb5a9e5b008027812e1ab47dba62
z7b1cdecc86621a0ff7adaa3353b64e31f556fd6fd1a9b27e4ca218fc34029c2f83076f4deab09c
zc72d9041949208016a44e6de9961c4cc99dff56ff4543ebc9ddae0cba1e41241cbad59b6f90ab7
z63e8f18878a36e1a3a84bca89365f00e40f4d50294a6361d3661228365571e038dc44cff2c0226
z2ff5fb1139725dd23abe4c8c10c20fd45cc8d5bb7dca03c22135481a7ab8c4a3156aba667bc33e
ze057777fa9c7632a6b7bdfe488448e287217264dc00e3db31f8cc09d301c76e8afce01c713503f
z258c36942ee848995d2bfc28aa4e2d88b882c4ba6cff2d34fa69be3c565f5b38662b9b51e4de60
z4be1ea04a44fe466d2052a22012c8bbf8594cc248f4c39e60acc9576c73542d208892f78fb6b57
z6ff8acfc5dff5ddb50635c442ea4f2d456830954b7b18d7980c433ffb10bf370a3644d4b3df217
z1f43176a2a9efd8de2d0cb83e6f4cbe6874e0b43ad32686679bbb6e94530ac84da32d934e7097f
z53e496214e76a7e528177cbfad02142314974df3d07e4f5c45ce8e2e50e71909695e34078ac39a
z84f2529656debe5ca98b6abb8f831c6c57da0fa3aef3fc558b3b5256670a37a43b9ae25d5734a5
zb40dfc1ae7e29f600261011c2fc544a32502688ac018f5447ed8888957345e5798af363e346160
z725e41004f74f6398f160fa90bfcedc26dbbe0961313b51958c6595b4699c8ecb7bfb605e9fe35
z808d11885c240e4109a360c58047e992928078e4eac73f144fa4f4e744d80243a5c8e7098965e1
zb7826429dc94d76cf4f31848f2436138e203a64d65d39841069a478b7198d330205444cbb329e9
zad76150d0e7337812f8fe5ee67e9d8b672d1d27e84288b8c51d5c85a6148ab116abacf651406aa
z1d1c522f170586a156f4b998a6d5adc81ba938da0a4e8c02ca52f761f18cbbaae09dbb0b8a011c
z6efaed14d11522e854d7ed7425bfec77962a6ea97003dfbc99fc42718928d4e662e3e7c19d04b7
zb363708022efed7b25208453cce68ca4e7667215b17114d911e4c0ec0a59649bc299f1727f2c7e
z900561786a1c6adc1db25b19bdd4926f2073af1f24b807939c4c0d334ef29e11d2f0d43fac36cc
z6616671bed5590ea95752f0f208f3ef71fa83745d20935c6f5fce030189e92b926b540a2c7e2d9
z3cb442cba7f4daf52072c766beb4ceaaacd81bb6c6353abab31ef3bfaa45151d699c5118d15a22
z236152b9541f5093141ec29cd2384c69a9fe58e69a539caa67ede8613ba27456a1aae0d020994f
zb02431ee3e17c5df2aba64ccd7907c2c4f2f63c13af022c29387c0d49b7a677d808527e6832ec7
z94b61a6ee6cb24316d50cf867a6d3ce78b0c7a98d48437f7b9389af16844f82d01b56592d72f9c
z28b599b1e4074d8c90b6feb344a35009af4ec645d4d516bf3de6973e21036009251b181a14904e
z471f40c7342b451c6f2daa8783b6d4ef12f8d27a33fecb3e9dc2b5ee49621c9cbaba2b03e1a6ac
z95c97240bdcca71311b8a2e110b7f47a9fd9a411798cb210de15533324557925c874fb8be18841
zc027740156c6c5b66639a7e74918566f2a3236cd0f913ff853cf66c20f7ff5779e02ce60bf0c50
z907704a77e92e03ca61264a03655bd8a6e8d8b1ee9be208d89d8e3525b233713da36675cdda944
ze960c6aee4b747903ea6189cf9f00d38b4df12428ecc0002f4386e9dd6d49d6b7c4c173134efee
z5d681ad19e16381c71e20cbf16b8ddd6cdf373dace6c11cad55bd1f9ab81285369fa82f1bf7e78
z1bd2c6ae7e0fac45a917cae250ec5ea80ae307b9cecb0cf2843071791a49fdf143729f61b99a5d
z4c45f3ca64eaba6aaa0949d1d16bcab5c6ce2369140dbaf035cf418d46e2a009030c3f5ebe2b22
z5c9dceb3c56da803b16d1eb5ab41a9becc33a3c93ff5b74638d473ddd6d9b1f1114f66489bacbd
z55eaa68be4064deefaae3a52068a34004c5674df68fe152d397547dc29b0aed5aa59f8ad1e2059
z7f181a45b73549cc43aac377451666381a933f295d64c6529affd943c6f73887475e8289b3ee68
z7fc7395b07c6e6c2570df9ec7393bfeda1eab234058f67f476b016bf2794fe4fd1a0e171ac1dc6
zb8138a5269de4edc11c391eb1660037230971e5ecadcc7fd7d1dd8a21b2914af55f46c80b22bfb
z998efbcea553c301f8664b1e303512c09792ff9df5a7f03d67acb87dfaef169db2e199e357c19a
z899509e099ad23acc5229122782ad20563ea15bccbc45ec3cac198e0db5a27ed6c3ab00d5e7906
z3e7672e467c741a92962736b24a31703464cfad2ca0b28496b9ed338362ea8956119fc3641bdc9
z74e88f7168cd59f5c71869482b4ee172cc639df8f9bf5d29d7cf0ca685591f224db72c5428e1a5
z46d26bbebe394d5296221ebb99db3811a3dd73ac278a03a0cd7fd111d5a283f68b56a8e0af7733
zd92030f0f073bc71ac8fcd45b30738e2529fab80f8ad50ca512640321645e1fba55d999e9e43e9
zf6008d214c12fb5474834cf09533893eb42f570846e978b461ff078c8beeb9149478a9b73cfe70
z9e93d4a80c6ff45133fb25b41521d673746bc1b95c9aa8f094da1934a4fadfbf20375a6e5cb081
z634899fbed7dfe35a09e7320b067557341e3b2325219056e585b71dec9a7b03aa2bf064c66e06f
z310c90345eb9e6afe16009deada3c11fbf4ffa1aa576b6839f8912d37d299e1d9b67cf6cb0293b
za6fc6b4330ae257c8909388de686e7d32cf02d5ffe04491a49a063188aea642389c4331a0d8d8a
z6d85a7ea09c0199e30d18e5604d4f6a88a672af25ca9082b5451399be13c8c0334d19e47127f03
z735c9f6655a7d3f377877d60053855cc61c4c21cd59331fb75ece159a335cbf3f043e0cc20a23c
zf6076f647b96e586f7cb30bfe523ec1b6852b06839cfe64fd2cc317784379b18687a7ad5fe1fb7
z0ce3494f3b56b2512426442fb4a7429f5977384065e4cb77e39df9a2bb854cd6e026332cb0242e
z996c7772e6352008f5b555be55dd3e9bf785e3db32cf4d9e811d80697062b17f47ecd9e7a48948
z3262255cd242905e1dd2676c2c1c105738ef8ae63b09d52e0ab8f9cf95812595f917c0b820c63c
zbc9185c2fe8fd347f4bf0b394805c3314af1e7f7dc6f9b811e147ed014dd864a86657616b3e101
zd38356aa62d132ab8a95574b352877829ee6bd2b31c9bf2a393057408e18e996fd4505ad6e0efb
z5e36283bc8b8ff0398c7fcc2d0bdea8ae82014b2df885963dc7dfaeb6bd4eecb033886d0b1e332
zbf48c8f19e0dcf0a51730752fd2bc32124375d72de163962a2ea77c03a78f93526b7d93c69c7ff
z8f50d59ba7c0239c3585fa2aaee32da1a2037cd437c35a0b55f17b8a20fc896571257168022e24
z84cad0a099f45e88b609f5ed4f783e0421449be42da9c1fbb90de599707db96d6512b98c0f6662
zc7263c156ded7eee5fb0a011067a4b513beb79aebd7dcbf0e3b59053908a8458114fd02e3f9d75
z7b60923c9b0b652a89f5ed91d89051866439cfbffbdcb3d0f5e9f7ada1b9970d54c004a6bab685
z5a742b9b549eab6198b13eebc759a81e9a406dd3ade53ac75041fedfc7c669d8779843471844ee
zd4947738f12d8ff0d1259ede4413333aa0657c88298a913c72e40624183ef53936118e57a51710
z52fc2e9d6f72c242b31db425051c5a574126ca3152ceb3c649d24a0c07e6891478ebda80eb677d
z1b7956be53be71163346477e92889f0d3b018f628263b5d4e6158919b7b85165a0c0bae205a357
z9cd75ec4674fbcba3f8db61d749071bbb8b57f509f4fa6ca287a8c659b03515f3822c6e200c55a
z9705e737a08e5ea438b479f7d801deca807ca91dcd8d2e334bd3615144eb65014d1dc22ebb48b2
za44c3e607c11f3df0ef0bcea59966ed208f73c8238b3926b249ef7f9b6e227b4d1d03ab678a83f
zb0b025cf890a6de5c2bb9c653c85bc75807357cae21912c82d7a7ad2f0242c45a70a114f38486f
z69d53edfbf0aa00a24caeb307667b6855a1aadd331cba6a09136989ca8bbc7ef35cd122a58a95b
z1404999d0b0dd4df88eb9efaeff7f0fd9c6e9cef0a64c9810679104649c3cb60beb4c65076d3ac
ze1dfc331701e98d866b3488b2742f86850f55faed91506a8344709492e436adf637f3733214a1e
z4cf120bce3dbdac8a15b95e64e6d2f53c8e4a87241867426191ae5d884ee0c988366bca11fe4e6
z610521ff18e68dd45fbc724232d72a1f372756fff536b73bc7c5912df6739790f4ca63562ed572
z16566c3e7a41947a76715f902f9a0fea5672c1cf34e78c2790fa5d58891dc651a5fdb95b6a7ca4
zaa501cde52683bdae096ff6d347171b1b892e3a47e2c13faddbf03ad0bdccbd9f6fca4b5a7288b
z64662ce47aad90d4d49ae12b5f0708f51e3d490140c39632c697705a4ccd62ae47893e4d1b3600
zf9945b4d104d4243813c4d5d61c06728822e36ebc2732620198241d034d768dcfff47971cbde02
zd13a9a4093aed71a07c89948081d0b2ba98c08967892a917eb0434128bf40a078d7d7c653254e3
z7173d53c14a5474925f2a03e99ddc3893c4ad2c7e2d37705ad6c9ceb41b32e334fd99ee902892e
z7735dd03bb28795105e5d30122436a1af32877f6b5f6424aa3a6f1d4f8418a8a44bad0eaa583cf
z2897ae3a99bf39a33eab760c986bde24f35323f048c384997ecc487636c27a323de0c3aab81279
ze21752b25409ab3dffa6b7854069a75eb1ba3340579475af820ad134d5ec6b6ed1c04590831118
z90466af44f793ef4555785d719be02018d1dd80754c739d60e06325287d7c0cd796ad80b156f1c
zbca01144219b16da16ccd2c003ade23e6ec73987470c859fc63455c7debe2cf41efa8f24de7e74
z97c40d2acc9cade600b6f3384514c7343838c9ecea75896ecb365e9a8dec2797646a75c052861d
z9d325fbc966034dd51dc05cf7f06ce8350d41c99440870b963d53b342cf9f929bf1a7f8edfa9e2
z3a5d617d2f7b49e38aac04517239b53202de5a5197f6cbf9155dc38f6a0d59b5c7fd6c2229a133
z13b62e95801207d5ceac72d6aa77c03e16c3de26aee2899863341145808d95b064450e3b26c5c9
za13ba850ffe39197872913b9de64f32fc245b28173f33323fce42ad257a52b829320458655152d
zbe390a6677968a129df767edac69363a8b168ba75181fcb90bb6a90b46c6dd1d2cef686389d264
z0de04ebf20b532fb60a3454748dee018a45a79692bf5aafbfb603fa35f89ea5e4f7fa96d910e4b
zdc06224bbc8ec5329c09cd013f076a1888ec8ca947bcfd742934192a4c1a3f1f54ff3334d37164
zc13b0bde548d30b30c04450298fb2da1594943f3c1d61c13b071e9b33134a1f770e8a96493bff0
z6678e6ab325e0f6e8679672a266f01aea3870afae4d1f44965c99b365686c48a33947177a0f7b6
zc93b9b60795f321e40226b062fc351705cdf02e7c8e50387d6271d2ee1421b6adf1925f7b857b0
zb39ada7e1aa3f58f4150a18b4c76bedc4e723ce5ed02bbe39e20d7c6d92e354679f91684c6d8a9
z20c14d5f36ef02af72df6aba371044d69d5d086746d8fce310fda8a24d4678dc131292659e9adc
zafaecf048cb783e38e0f095540a4c80e637a98094ed1a4aded7c4cbf620960a59d3729ed2c7371
zb41588e0df2d9dbc941b890b26b4a800d32e59b1d77e02146d139a631b897bfa344bcf7d5c70cb
z0bf8abfe7c64e41d2b072a0efa3e69908b139fd3c66f8aed45721a52853f0fea3d671dad715801
z38559ad78440577e90d531a8568d7c9866c3b16353fc4335fd2125f402cdea31c61b482a7f2b5b
z233afdc5500fb5d2202341f3d852e0f7eeb3c694589ddd135739df667c9ddbbd9445bfd0b4eef7
z232f4535f113e86f9515f363a557418260f19307539f7e0a90296d3e3a96c386075200ea00cdcf
z65858246429103474b3bcde94d83bc58439e54eedebc421aad246113d69080bb1d76f9b25dcf21
z5f1fe5340fb1819b20c01372e8289ed0c368a5b350c271a5727f4266081656b853aad8c18db495
zabbb3134ca4ac08bbcc801d086cf20ed283e76f5a9cfce52ac6d0467f01ad006887694d4f0ba43
zbfe1e1aec88c993398dee7519c408a75fa6fea43e898d08de501bc566534265d6b91baf21ccaf0
z47c4f875ed09e527046f58d9a6537166479a30743197d616cab3d7c28aa52101b1d2d5561ad79a
za591cf0cadfdfc3f1b8a49907dea9c99ec4636fab9a810c50235b24fb3540e439f997f0c6b7b7a
z0afb449a0539bc3b01c1d4bea6bedddf4c7c399e68950914b596bee88c84112824c1927312d29f
z4d8d811a80468e8c488605d45837ad0a382808bf0f56797aa87fbbb220f0747faf5effbc291da4
z84f45b8068a168a49836f9a87b915220d3ce6cde5325921a7baf42d8c28183e4bc677f6c60e0e8
z7ab85fed5734777141070616bbac9e86faec903951804d9a55ac51c7a8342a99882a50138f4e95
zb8f32ca71d23051f4cb79abb32008f31e5c02c913fce163eb22ed903b746053f5ecafa900e1bcb
z41f8492675ab87f5b17b5d72f7387742dbbfbb7a23bf29b57cc4d162027e6b17059024cb877dac
zbfd69b09ed7507ff964f2a1d13d281e9e4b7dbd58fcb362b8bbfe80527d37df2ec94b06e237c5d
z7095b468989b19f307e000657b0a8c1046489ee069006c9e0249cb14ea321b6f2432260a35f05c
zed917c4f5457926fefed5d753848df432e359f5253557a192734bc2370fe66c58d86519684ab51
z2ec70b167d3f565f61cbe738c4b7b9aa23c5c79ae9c56ed423da94017966ebf692c6da0f8b7804
z158620c86945d71d95aadfc60729f86f72e56fdf3a96644e2b57af9a9c3cab2e6955dd55771b25
z5260c2812473950fdd60997187c500468781166b4be0b33b8a3179af8e897c18663e2116619184
za47a9b07a71bd7e58d7097c82d12c0a1e9ba0bc9e082952786d19d81a8b0df7632f46d3a4fc22a
z6ff5a83b97f31b900310f5478d05ea9e0ba281ef4a1060ad8fa78f6687977e3f0e3f72c1e89ea3
zfe7824db2d8f5fa4805200868c130cdbcc78edd96192fc749e7b8a0c5ee5ab2344b46d7cb6d0f4
z3669139f53aa8b666669340a4dc36bcda181e8d3cabfae61f6d878e1dd2ca2f9651a3772cd3a32
z50dd0053d9341e3ef9db4829537fe8caaa77977d972b93e40d002827239cf55cdc3cf7356d3d2a
z5ea45fd00719f965b5cfac33900f3fde67e5a8ae5eab16d89f0eb00d226afa45c3c0a7421ffc8f
ze69ba063a7a8769f3f306843220e7ef31040e99d6bc8401d839eaa937df13917e8ead9187c1532
z4633565aa69e896ddb03cb09e584987c09a80ce22c62983004d7bc1222f95da7358d8712bdf145
zda7706913000e1b5453cf1cbf83cd0b185cd73b03c3b9bab15c183e42197dab9ffb7051689d7f8
z0ea319cd564eb03cfd041a7d51febc944e99fea10cee2429104aa0230a58870a152e2fcf56cc82
z57d9e5b55773f3834b85d46dfd93f75ed7c916ef213ecf241c2e19f46e2731a0e265350669116e
zc8f3afb8b2db015ccefe268ac10e0ab8e0fb508a0e77298d454e246b1a1b03d12117bd7e36081a
z3100ebcb544b01d2ec86de76b20280eb526d2b02e36151c91bc51602f06001877d908a78d74ad1
z7fc343a6b7d341252049d9e02ccac98f647e143385f0cd2ccf7988c7e733435c6d5167242a05da
zdf9f414380dc57c01c155d1336a9d28f8538226d4c797c6d6910b247d5cc6fd5f439a019e1b5a4
ze8fc5d19adfa15b3d79fccb70e70e4abe758b91febca921ee82f656210a0fcf46cd3ffca383b03
zec9ed0f67d89d1f4df751bc25f753c5992cdf77a3c991d7ccf155ed66c0d051a315ab69629cb03
ze7b94eaa7dd412cd2d1e1241bc8b18788d2a0a9be0371dca95938ef64858f55a85e8373d04e5ed
z468bd166ed132875d9c328f74a0298ceae9514abe2f9017e5bf2db28592208df793aa3239f6cc7
z67fe411769768df5009c2698630afc180e8aab378fc6984ef1478af4fe7b84e17c20212a2382a4
z81b4768754589f70e01f478428747b06f894405ee52a8ca49f350e76e4ea9c64bfd70d26d6de2b
zbf4cf32d1184884496d7928e459e7b53efafdd9e3c2f4ebdc7d831f3ace70f9f058fc09e9f91ae
zdea9f01aa11ae3247e3164d62cba1b3883bbf6536be1a816f417bc23b4ff10da89356b06bd942e
z7fbd6b1550f54e8c758dcf8798bed15714ad017ec14ccc1533d72ee090c39cf2c798bc917f4b57
z5514426440998902f288c3e2bd29b15719e559326e54309d757f6eefc48e8309071f32ebcaf859
ze477e511e9032f0467b7c975c9f3b504bcad16257c3c94d07acd8d91fdb3984ac37d6a828ff501
ze4cba718af512845a8c62c5e04ea2d01eaefa4d49436fdd59465ad27456617cc7c22165c05aa69
zb5859183aef6ae4a95d2b3374131333e55f8e337b58506a9f7b6c9e3b6a7aa077679bd611470be
z6cce437b51f36d1fa671ee81fdeaa14216cac69f434839859b0dec8e9a449757a12e28b52a3f2f
zad2e6bb97cb718dd1e1b74f11713837835f1840c783b520777317c02a485cc0d20a3fd1ca4ce98
z1161750eeea4259b7d1dbb84163332b64ffcbc19ed8087fd8f3cfd8e8b623af33a0c8b9a7ae72f
zf11784e1dc914bbba93f9dc6f136ecd8089aaea5387757ccadb47d966c094b77df3ee9a652a31b
z43013d425fb02105906fbe3b62300e487bfa7a45fadcf50ddfd8e18e635a9ebb27c52bc12a0677
z9a0322258da2677ee875fe10873265e111698133cd85cf289f4f96d33ed24d703e3759d442a55d
zdc801727ecce924bc2f23fddcba21a66f4395333cda663de8e6650347adb65e713682b28cf9e7e
z2dac73a52030797c121a3abc580b5131336553c3fb97e9249e66a2193858368d334e49b5d7633e
z09d0a5c70a252533a821094437ebde9c4429ecb496806cf523d80deaf468d3f544cbcd46b0f53b
zc2f47087e4d7a57486238ff73ec6f181f65ecff8ff2c1c2ed6afd1356f4424ad9bce8792f23bb6
za131b655f21011e9e065e7106f1f20a8ede9e0aafe1b32728a546134021885b59c68796a74dcdb
zcd21483e679660bab3c88369165082094737c4f0fccfd4b9103c2dd3ea48ad49a4fa190dce51a7
z7e884f4db0519fc367d1afec9430d6b6b9e3d29751d4bd4d07f094032a57d6ef985c54ecf0e788
z3f21c615b76c4cc35be352e427576027ca0f4df8cddf121eb28981b31f5f3660048f2f60783232
z7c591826586efe497e4eeb42aa1a5d705955ec534650cd8f390ad2a56e765df23e91755ef60f6a
z66ac0709a233c7eb476d56cc6e9fda2dc5d7ec446bbfa037ba04f7047f4a07c88202c3fcb380aa
z026d32ef18ecfeccee01c4fad7bee79100a838750c62c59020382e5b38206890f201fbf2c41806
za9c26efeeba197fca821f38fa48f44888c97143f7204e11cae9e48fd856921ac1a1a1ddda3865a
za6fb463788dd79603f1c3a993e2b45feb2c6048cb8172e60a9cb65775153c1e7a59ed63ff57abe
z3838da3f9303205557103634c3c3fe1c70430f79c61b0e06436371b4af3e1e33a4342168d55d9e
z744b87f460a7fa7d0dd3155440b45b1891df779ebaf327759107bc9330ed5125d22aa02b78ba90
z45833eafd3308c70188d4710f75deee5f1e549bf5dca849e4654f40c88848c5165fc7458abf7f6
zb473f305fd362d3f87fd6a19491293ad7f98ca11ea12bd6c933216c9d71bfddd41d2355d33fa98
z5582056ad7b61e1c65c0519836a611b0b077a115b561618f48478d24e9057175cad7fd99bf983c
zaa33267398d4d0a7431dec08780f9ad343d3069d0a596fe09f5a91be20c4f04c3f5ba4ecd2a71e
z9b1b8f82e82d8942e4b6d6b6d030f814139069f48cb52a63e76f2074ede2a8ca32c43270dde995
z174c9d9cf4450e9e27ebc864dcdda5fde783d97418894a4514c7edb095eb8b4c6f48fcd1c9096d
zc5041c412e512ec8e81f6603008f75da446bf282ee186e8bf9b132ec3f16d0d15e407ff1b934ae
z02c17e522a134b46f642c1b2c54c89993478a302e4b5765e50b8fa1c1e0e9ad1b80b9293627073
z0629a823705e4a4e70ec86f51bc4abc142aac0544fe6030695d38a86173fba9ce3c07a9abb3a02
z27f495886084850fff5c49581d444124a397daa87514d60ed7bbe419f8d653d40e2c01dc75989c
zff633e9b06eb049e2e596689a7ec12fb76e87cf337d246f26677e63eca2543cc239fac946171d0
zaad7cc6fa7c25e01a8a7500d97f514a8f9779e6701cdfb05b524413b3f345ee5c7c6b26b9417ad
z954095539f24a6b3832081e098bf414e8a76779c1fbfbdebead8d7c91b3c2b69de0f416cfe0f16
z52a93f0a6e7df9ccec4eeb626f78991213f219af4ee4330184e578c77bf4c02a527759e9bc6967
zc8b1b3d00cce5f733a571205e6f0fbb9f4694b8bcb693f9e2519d0beb47a20ebcd1096c640c0c1
z1b25fc8678f2037d85d13b92db1c197edb90d37338cbb62a45cc56a44923ccd9419045680c06bd
z91682753bf62f943ffdfcbe02c379ac401de120c75c0189dc4d4b2859df3b75135356d82ee9d24
z2d879aa7831f9607b861a79badebfbc81cb46fed64f14bb61b07afbcbeffa2d247f6b535e39952
z6b9ec6920713e2be78a7ea99dbb3ebacd05a029c0d6ab312d398ccf38bf77a770bb5a4e30548c7
z7e439834812b9b62a190b30e5f95ee064e6d9414062de3c3d1abea26431c88eb97b1470974d848
z5dc8a9ce2edf96c592af364f9fa1b766e648e9e0b0238e5b938a225eaa8fddbe4d20c67b8a8d8a
z2bac9c65678910bf0adfa747f672be83a83b352133b89a130d729a66c1be2215436a796fa78cea
zeaa11b73db9440c246848a2f2a57ea4729c8e95ca3cf28c3b528ee34d44a5e0549716ca930144b
z28815c128bbffae37e19548e4da09234caacf3b7000855087da60d5af6c94fdcb1028cb2bf21f1
zcda185d7fff0829e248cc58bd95028997d1567c27ec8f2ab52495141f24f24372849ef40a5fca9
zdbf13e08d0d0985f5b2a706c2b6d4e3a959658800bb92650458d14a10df1b24558358e68b81010
zcc2110ad139aa3cb98c257b928f7bfda2c9f929b93bf4e62f4449468f89404cef63d036c938884
z3a126af7e1066a0a2085520b075c1f43ec0767ff2431094e03d3f1e60a1c359e03c66f9fe059ed
zd6bb1a22d89e33fb67072301401408ac8878ea9c23a00189b20080c6fc79b67aa41d67df8b807f
z69d03d61d96bafeab3ced2f22f2a33523684c45c445b20836bcf35463fc03cd4f61e23291f4b38
z9915f53f132cbbb4e3a6be6cd2e9dd2516534efbc3a06cfaa3873820f9795ece5014bb47f27c71
z70331fac08e0ef1f84c0eb9f9106ed2b4b40a68f83a61b7f4ea4c445a88bd202704fd6edc2e72f
z310e5aa868efd72e62a395a26e46017b0d3678ab62fe827d27879ccefa9992e1f463554500a6a1
za188dad1f177c2a90b7acf5cfbf3dce7d95a891b69ee636c6068f3ce46fdafc3c246b88c60bc59
zb000ce65a126cfd1a620b05a35524b2f195d558d4433b9c5d3add80a058fb7ea41c6b9c218fa65
z3e145a17dab15f1ce1f102956808dacf0e78c340deab3a03ee7cddf4788450e91f1fa4c0ab458a
zcebf3ce3cf84a46c3ceb0a90d0c1eb2459ca25f01072f2087347d380d322dc96fcb78912076fee
z1be812c4974bd0d1ca739ca4f87327b5b21f2ca122bab57ad25ab9cd1fae35452aa0a3097e7cd4
z02dbe864b1e09b0c5f742b875da73c94ce5c8a4fb745614a01e4f11f34a11ab10d643d3fbd830c
z9f3717e05d2b89bfb5f54943d4746cceb1c3f334ee449fa2f0d678a5bd190147753c094a9d5b80
zc014e27ba4d7e46c8de9518d7975b46a78ad0abe3996de66332401fe1f6310161813d61f3e77d6
z90c5c831c8ca681c35d28ca5ad70932c498969ecb3431d782f665ef4fd4d852b887bc98526a806
z927e96573a94a2eccf51b5dfa2521b880dd8815d07f6fafbfe739f4604eb3e57f872369c6736ce
z33a55179f0fc7a327ef0e620573a811fd16e89e69badebedc77405c40c8d9ce368dda48fcbf4ff
z19132f2d6f6b1b4ac58ae1fc9239e42f5f68daca7fa81b9cc1a0d0c3a46063a54b8590a9ec880e
z4a01b6657d70b660dbfa81e23c4c69a06cdd9bcf175da3436364083bf09dd260b792eaa2a5688c
za7204d51e54a6543c51ae88003d81b7594552ec78d5456e81f782c656d701c9ce5b594c59daf37
z2424af19dc6d1f8b6b7e4059265dad9fd637304ad756ea2134cc9e82c37f3a996dfec20828db24
z2d90525247d76bb20ab65b91acc5f76e87c42c80cd97cf8a9c01c762dffc8ccf4a3f6f4e5da153
zc4d0e5d9ac1730676c018430c069377b730010510fc9a2c2a94b5a752342dcf7ead254e7a986aa
z4dcc38bb48efba757c64b490fc716cd462ecdf44cd224e791630c1173d6eabb200b400ee643163
z022f548a2645072e529dcb67dbe80f21d73d8ab4bee51656b15fbc21bd3998a73dd280c8152b36
z1676c9ab59fb42b57f2fb2d0b4c8ca2aee0511b3ab1b2a7193a5baeb8cdf78507197598b548917
z3403229893babfb0647da389e7f757f3819bc2a126efd0f7c16397537fcaf899dcc8b87c4d88d9
z9f8667c35fa92c047e066b23fc25e48fe500c08a92f2b45fe17d25c4b17942bbe9178b87402338
za1e5fade2f8f970de397fc3ff1f71dce4b50bdfcc3b178a357a76070d2b549297408bbd11f610d
z6376c1cc6da6ce07c4d2297dcf6288fde097a31b30df1a94ebab86665835b925fd472021d931bd
z6f70c0650b757b5859fccd9a3474014542a31317bf2d0c66addab9ce61aef7d988987a3fbcb860
z57f09b6e4897b77e5cd351f2783cdf32d09800aa342eb6e40d0c7eb9ae5b50f63f762a98dae102
z53d8676f49d255a1312ccb38f1e0f93d0d3542387cdc386c310e0fd9367b8980ebbf52eedddfab
z2e2c13d107ecba32195ecb2eb3fa4e1cd1f74439a99a7e4d36dca704f9e935b4b4a107122154d6
z28660eac39862b22466227e5272b32e9bcb3bc7e0f0b551517384f3febb5153dc95d99114f9ca9
zfa76bd8de39d6e47c040ac393127ee81620f1d0619dd85266471cff49c7eea012ed07607afb247
zdab1522edd67923eeee905d8b5d695da566dd0b29e776fdf2ba77995a23c77483dd934d87f2f55
z69ab3c53cd2a7ed8426462c445e4f2f1b462c583dbc3d381aa46955dfe300ac9a5283643fd4611
z1e40b331604da653772ce6f19ff360004928ae7957690503fdcfc8273b57d16b5e4a04baab0277
za52189b7e6c64b6a7f0748e171a71659971613e5e9e4e62135d875b335c1515c993d7ac821770a
z5eedb9eaa3be381aae2167da9bcb6c6caf7a49c129f2b8b16ad47f14edf9b6f26dddf23af96dab
z22d021725114f8f8196105f8fda5c0d4bbee5f1db055dfcb4890ae6502277fb4dfebcc3d987fca
zeb352bfb849c48f5f081d00b601462cbc1bbf389f7a709212e6c24ff2b6a6be4eb170daaa55c25
z688b4f5ce954de410c71c26f3e6c4bac312f4838d8fab0402cb1661f80977fca1bac2d631d9751
z679d91e96035f1ae421647b263d81372b1f107d62ce60eea00413b04e5a8db408062d0a7bc3dd3
z13001819ba9375ba84cbb03d578720fc8770ed067dcfaeada8f6bee70873cfe262c503d7891f54
z48fdcb6949d5f8f7629db7a7843fd7898e99603899016e6a500d4e1df556c65452a58464e87be9
z7559cae7cf1b1b491a7127deeb0b852ead09860c9d6a6691adc207dea3c720aef90bb4600c97cd
z07db4fd15167dd15b98c7bdbbafbe5d1565425608bb66364785d6101aab0fb2fd258ab49f28543
z85e04f04df838b7fea84da44613168780d6a41f194a36297e0219fd2c5fbb02412f843f95f4977
zc9e1c6a10b175216b122a70d7adfd40f55328f563146597253449f728fb4f625fec6850245651e
z1a55a5e7e8fb89bbf58ef68c7de073244479735d2eb420491718a5c7243102c202192836196b0e
z2fe3d470a60f57af26c4523802f6b2d22b38bfc957d3c0e72de58c97fc586c7a19b524b46c4b0c
z37ad3fed6f25ef6d705660559d75fe024aff65c487332a7060738d0e3eacb43b9220641aae62bf
z9dd5bbbc0a9d1faed8de835edf2467b4c34deee2fe428f10132213ab1dc5edde18e66fcf189c9e
z818bad40df77cd553fd2c84f7aea1b9283757768700c39dd4adb897e44fabc361bd5e2fe44bd77
z00ff65dbd17ed41bb2a61160a181d211e86d5d99b8e416aa28da80d34205a9d2aebbb51d261ad7
z8b7b120282729e955b0cedf2fa90dac8fecfe8393d9617fd57ee4089a7583a0c539aaa2d2cad6c
z285170779bb2c188b02b2eff4497df474d94c506b90092e9fb9074a4aa92e3a3fec0358ef446ff
z1109ae8ea59f6c22fe05d2a3c66d42c506adf555e19642179608991364fed12c2648fa53a55553
z04ab64f83f54b1d17a6655a3ca0448c8174227b9ccd2915c2e2dff1ff4f477b0056b16e900e87f
z7c9e28b87e06be2a41f86f2e03ee59404b7dec70b342788168e5e6cf0e1c5798ca61490ac7a86c
z365dea1620914514bb4f601027786cd550127d136c396d16de9d0ae8871447e7c62b93cefa6d4f
z77924bc160db33c726662b7937a7ba983b2a6b46aa20a9e1e21a7bdb60885b9bafd61d309283ce
z6e149a9651886c8d7a70644ca6c972abc6bbb1ea33e5a00c23f01cc234110fe6c1d2e17ea0589b
ze68a6f49b3d1464f86f9939125b3a25a8b40b0316edb0fd23d1610de4d8b30679e3a7744939dc8
z2466f5b583fd682ec56fd0c2e8b0dc22244bb835d0887425e03e4bb6ed848e61b10de7d5455b96
zfb64e002dfd4ff4abe8c770d128aef169c58c653314c98d02b0118922eb23b49365aa9fc53d749
z8b48424edb3928e696a6ad319663db2bcd4411e22f4e9b76eebc29618974fad217c66be3d06013
z15246ab41e9d5bff864df3f57405365d861e1e94549cfc377e486247d74227b774af9790554775
z0ef21387be21515475d80d82fb9e44e97d6be3c4da9da9073ef0a6f5aced1c76097d0f9a302232
zf6df6b6382d976c1c01083e94e65dd8768b2c30a1488696d387844c2078409fbee190548f4cbd0
zf20ea2b0dc3bee7ce5a33876e0cb7ab2860829f0dadd546c8f363f3025571746ef465a8f413278
z7d9e4e50d6a33011ab705bd1f0bc775a36b41ea0bc06dbb922dac4464016fdadbdcc99a37a6c0c
z42475eaab355dab5178adc5f4f5acb39ceb344701521f560399dcbd9c64253eaa61caa3b2e6cfc
zb04ccf3b3faf728520930548df159388701a9c825bfdea30255c191a08ef20aa19e9bc0cb5688e
z1708eff04087a6acdd4de4a23702309bc11f67974feb90da70b25585d75df4407a3c873a361391
z0b818b53a90c7eec5c5e7f10dafdbed6d420428313470623c1e39b5e5efabda54c0dcca954e7e4
z56f99d825733d08f45cb87874f17303c01e9fb751e3bcb38cbdde568c74a0cc9204146351a7340
z845d053de4fbd4867b2e6d14125d7ffeb4493982cb7a2a4af49a172d141fddf96f3c5b2dc6bcc3
zdb9dc34a37a02f62d3dcc703ca2008ff2e653620ce00216e86256c2326d2338beef5348d40ea3d
zc75901d0cd6ab6d9545509884dc9e31369d87d2bbc4e63d6f68988c83cb1c150959650ab361ba0
zdb1fe3e034381306d624931f04340767bb5aecb79a4a2666bc22defb664f06823e24fff12f6336
z125a46b198a210593985723f3d52f2e7f3070bc6954dcf72756794c38fa343426bd8d48f3275d3
zdcc4a5cfa02148cd53378b67553e6bcd4aa2bf2be3f679ecd386f4c4fdc149cc77787791b868f9
z477cbd9a3965ec906c4a5a5f246609f75d89cd6462565339d287f48653100c34823a408a71f708
z306440766ddef6b727af6b88d8ae22248032da148a5c8e0ba5c3363b38d7b22c10db1c606982ca
z4194ffc4717d698dc165b691b27587430334e9eddd14868cc1e94b56bb326e534d0f1919684956
z102c196274ee6c9680f901dc689eb3f4eea53dd54a5a40d04b95cdb1b33cdd978ec9e902e53626
z922f4e3eb1bf418e8c550108a8089cac01beaf88a17613e5310774fd4d0668bc519880357c04c8
z96838bf645d0075adfc9e8a54cf592aa5ccb85034c1492136391fc707adec9bcced9399db59839
zdd9411fe799aa98766628d3d9e36833ed592383d66ae750628a64725873ba0f76426490eb876e5
zd7acb262a5e8cf813d57f8458b4556e03959ff83dafbbff6ba796288a29838393988c25ffca807
z61b9d39ea4c52e784abe324230449ce53fb270c2417504307ffba4a6bb5223472dae0f869b84ff
z9d46ee34d1144c98c5228b865f6c1ae81ac1d64b20df428e91bb22a695906b2fa4d7d20c3b2c87
z6a68710711661b5660917836d1e136d1ecb26b1cc99e65d8f0ef274f277eefcf92b966d3dca617
z8bed84c6b39a209044a0bc9f8526e0cc8bf84b7cb9c1b008a0acd21009e64f2ed3ea55579223bc
z4a5e8fbacd0e6ec4456158c32848ff16204262add9405f58cdd4bc1b593e414c6bbf11d346d9f1
za3e6cd40627b4630afe165a788cb6ec495472db1bdebd46e2aa627583ac6a8b2d85f72d9266253
zfbbabe5a601b4761add3728fe266cfac0c59c90353e1dedca767ba8e5d74f0adb3a4eaaf4e5598
z78c6a3a63fa1ac282f82d11731e141b9e0d1725b46b9d1ab5533c385e898b7c5b2bedef7a0254e
za3967c6a1889be3df3466b4a0f34a284729f48e8b3a50d05d3c47d3a3f487a4495a2aed0a64d41
z6419782d979fa81776c8807e42740d67dd651a7cd1a31eed39dfeaf5826493be294611a50f0ba7
ze675d8bfb77b3c539ea0360052e17e33de4388d15cdaa23959a5d1bdbaf6f422f13b0493f97046
zec6f0135e856a03978dfd3ecdbccec694e60ef784dae8f981a8f29b4cef7f006cb51b251f29ba0
z6e3a36fce42e306dd036125d09852b925dd37b19f4d769faa185001e48413b94028ebe8ec64e87
z8e42973d76d52342b02f7f8ae1f08c22dc4703ec3ae657a600d7fb9a8840a1d54213d99b814246
za9ee9060bc41ef2fdff133febc363672128dd76e3f63fe7d5fd600afc96b1fbb44439ce81fccc6
z613d83fe541e451cdc39969287d898f7635bcc7f17a62eae00cc766e19cb0dc1345b2133e0e4f9
zee202a4d2e9db7ae5c43705613a3f706a6efb9b8b5bf8ece93fe2534ee42966721bb56c403afea
z3af3b71c9977d38ee82d33ec09df994b5f1768ebf90d6bfdae2e321261c8350c9da8e90c9313f2
z75bd7f9140836fd91f4bab6e53b1963761ad3e1dea8b5cef9d4e0ca57f6b091ded756a464112e2
z30b0239d271174e7d4419fdf5215f9a2b0dd622b2d7fa93e6a56dec259c5497cfdadabe341a973
za3b957c88ba3de34a13eb58b0bfe81433ee53c228e0f2a5e3e466726df8f2c53684fd61234cdb3
zb35e017892c8f55954ebc7c89179f6cbe7c1aff1e74787b7f38c4feb6a376ece16e24dd4f5da55
z9467f0228f1df837ccfd18e5a6e727ee50d2c2c29a7f810cb650e49a0972d61e83d432e8086c63
za31b2f0fb976e59e4c6c00a97b96e1356c9ba367f25f454150487eef334069300725b4822faef6
z066273e0f2b3aa684017d4c982995369a5ccc5a0465a36c387edacb93eb3b8cee2c2f29753beac
z73e1b8591467ded4caff6c671d2845268705fd9e549664a109a5decdfe7b367723d826fcc5355b
z3e9f75027fe621945d9fc056b5b51cde31dbf225e48954374a20cf37b2707f55392ad705f64b00
zb4e99b0b7889195428c6550b0da1805c63761c2c355b59b550b97daad290782601753e5225a159
z3dd08cec0672bbb92689505646dc9a2c4a0c376a99f824857f2064e6bf46792684b3c681bfe037
z532997df1842b854fe8e0b9911aabe9e4fd478c586b40a0951c3904dd47c008821460b8592e29f
z6ee7f1341b45cd01da48985ee505ccf7e70c727395f4c580eb9d86a3dcea83ee855a2510d518ed
z0e5d7441c71e0083766aa386251c0595fbdd10df1baa7b1f9888093361186172dd9a015efc84c8
zb38b1a76f94d953590b3cc58b84963f18c2a0e897ff8f8731194e3e60691b4d54829c01a6e5e03
z8240ecfbd12bb6498e1806dd99f55df5f55ba9d4a9668a8f1e8be04896c759d46ea3a69384107b
z40b643f1ddc601bbf6ab7dcde59cb70fd5bde87f1e56accd5ed3c2146b56255dc35fed2162bd18
zb1822b72f24bead785406fe301cb1525b5a295af0f3f3e9a0e8a946575efc4ddf7f5288a87e449
z47e31eaca6e5cc9b411c91c8f8e7e9124161e921344e27614806317d9c3279d303cc42bc3d1dca
zb04bc8af6b605a29ee5df69ab517c136eac57dfe5938cf70ca78906bf408c878bacc5f40a559d3
zbcc5570740ce8cc3266596a62abae0887c4ff759c4955cb1e84c6e4151009ca1376441d01c59be
z5aff38387f48574e4f384342be9e236a8d0ff6083f4e93f36657d6f0f019dfd26fc9d182a9e269
z2de209f84c8124bcacd36c5c183e1824244ba48fbae41d3419816b5a59047ccd990be54503b7a9
z2b87be8efc34b62e47579353275e81ed57a1f7ee6cca1dfc463f107becfca5fc9b3b1134199f9a
z0c65f5ac492268ca07bea4fa65ec39a0ecf8433254745d5dddc87fb23375b4c6050dd32d32d211
zc707bbb900b78ade0e4768591be244a6a00a9bd13a434fe357175816672a7eb51038b782c2b69c
zcc80ffc84de13a71ecd30340b5f50ffb3a21b7fdcfd867c1d516e6271f436a3904ee4d42ae7b38
zbe6008c5e48e5c32fbdec1772a3d6ac282ab5b86267e9aa0ec3d160e02c80689ea34a5b689bf63
z1e0ddb37d2311b7c83362d37415b4d8ecfa39b5016a2aeabb68ea0e266cfec5b8f7a91ad9214d7
z84c822a7bfe7174441fc3c2039f9e1ef31138f4c452afcda8f658710835c1fb5cb9d1f0b2a212c
zef21ccddeef9f84611be8232f138578f43530bdea0c6b053ad75f96a48898df4e5e1a2b6701516
z423e5616c9c261d0f673ce66716e5a8996e91072165db78cb68edb825d860abbc765e7604450b9
z8f1d20aedf028a3ef27aa95209ea2d6e0a0e873e51942d252a7db950afe83b5009e677a547f070
z43d794dbd4b1dff27972ed7479a3c08f7aaefdd1e51e44a916d3e77a4d09944993c98f618c2005
zc02fc24c24da0d16846f5e1890e85259a399934d2d98849a4db3709f3240224e31046cecf44417
z6f33c861a82e549491bfe0a450256103acb856ec53c61b52ce384cee8c57e6c1fb9cf0944b1eba
z6bdcc3d052c14685b86efb32290f2dbef77fa3d404e66b037a29f651c332c94fc996f1e9989cbe
z2ddf330c11684d212d77b05a1bfdff7d7f8ed96851108dc8cb64ed56093d963d994d69b949b282
z555cb613726ed0176f144836f115f21e269600fde03ed0131d13aa9dabdc0499b8f8c125092c43
zf76a3ce03bda88aaf98e692cd5e3aa7d5071ea410af1d8f57dd45d69996b5867af90e719dd1272
z1ca6d6f5611233a53ea97d013d0c79d11937fdd9e963b7cf9c392aeaa0e9bedf6ac8a5e53b8814
z01632a4b85462884eb06f04e2cb24fbf9a1bbcf151fa76fe8af8f286d09ddeae60d038925b29cd
ze16902c932af3a1fb12569eb6e0e188d1eda0d4537fcc064b628a9575ef9d3836f2ec1bc9830bf
z2fbf9466c83628d8338d1300a55ad1afbdc91787057509429074f889b1a9f4d20ac7f33372ed82
zaeb7195b4ae6a779e42c67127315ee927b32eec529c81696ab5ba50a0162de6b68dbe7bb00deaf
zbc88c525454353b43cd331b5d44932b4596d56efc28c9935df957c111699a2848fb82957f591cd
z169c1f2376a07a1bb7240eeef54df03012abca6807c52d2869ea14d12ab3951491f79537b11060
z755d4b3ea496f7b92cb2bdb4d60ac2a7771037940a9d6610bf3092e45657e9b7aef4781e6be78d
z126fb1232634e24e0ceb01b22afd1930d305c576c35b4260ff347309294014bccaf494a61f5ea0
zc9405b74ac67c10ef1c9ce92da872e378ccf18253b49dc7dea95f66c818c41475c364fdb749e71
zc3767c14259a72aa3e918c1740bc830e8a3f2e7736e5b90b234c543bd5feae6feb7a9481a16c8f
z780f2faea9054de55c2b9961ba64b7dc3f4c1836ac02023bb8385c8805d551a023614f9e463d61
ze9bbca12b8e81db80b3d276cb6aa7817927eb0989d35e4e2f890a47d1ff0e2b9f67a0fe9c82704
zc8b2ce6a00cf3a7cff7cf1e6df4b4effcdbbe5f0e810e37d81da9aa600b41b842655a9e0e5c81f
z45609eb5331d289e121534d5adc9fd678ec61950cb93d6a23bec02927d9cc67af7975583190f57
z6117c4a94d19d349e8d36c869821a85a9c47c394802975dff2844a5daaf9431c12d70e006077ea
z6648b05b3bdc0b0b7c058961119a386b9e9f0b109970bcf4b1250506e14773a20b3a8a6579c3c6
z76bab038346a94696ab69b53b705406427a5e1ca22d62d66aec1d25860d7bb0b8a81ac6e7de62f
z22277ea7ee465e68e6e145a9be8ae2b15c8492cc0b75ae1f92aafd4e43ebf7e4c8d6b261c40521
zf4214780845f5ba45ef1f0be16686cd785bf0a34177a87119f9f6149aef2fb33f903dd9b89b24a
z7fab51288a3e4c003cd00ec876e3d63b1ab2849fecfdd888fdc8d03da53090969a50e587ebb7d9
z7444c7d9449fb3b1ad9ab304cbcf7a628f3e3824fc5eb3549809ea698d245605cc85f776499d06
z51ca45f66c610880080fff334e1a0271363cb4e7b83264299c29c98e38acbb5f9f3c04f1ca7f3b
zf21c79a648c1428302ad2882424dd31f75b6f39e16f252fdb85ea608890f021fe653c1ce96e134
z69a26ecc42c3316584f681aa5a41bbc7e2d2b730395216ec0f8d7e44dcd47df3220c47e9d1d8a9
z6186e8da13652f57eb85e4a3bc6eeea64f84ed4b5baeef4a4e09d7d8003948eec363711024352e
z0b62cb20da9aeed347ea03fdd381f8ed6b1a904ca561203be9277703195ff304ea52d5962f9ac6
zf8ed941784b3b66829eea16fe6b293110c5e32ad18e3d5ea75e67c252d4edac64257dc0a73caa2
z97b2f7fade69b5502048123e1bda42e6b73cfa9e79380bc5dde2e94b5d7cb6057f11d2aa6a1750
zd204fa06f50fa28fab0ce541862e5bf58a6e4999aa4415391d02ea3141433b4044200ac4ddefb8
z56eaf41a04ebf39c85af53845b78ea812a0b3856e50f7cefbeb264b1ab32139584aec0d4245087
zd6ee4fd2618c82fecd66b42fa235ab1e70ba867e3d2405344354800fcf28b3810e201315cae43a
z5e79b179d460803b4c7018d28f2943ad5471b59af02cebd87b47f4dc3876ffaca4ad5c462c5be6
z835576735213a5d98c521c231d001ef40ae69c7d3cc4523421d68bbc567b9d31a3434d0a030cf7
zc8abdb8c5e547a0cd31e5b41eab3c3079a890eb852104c1f001c5b1923e75175cbef2d522be518
z52caa04cb683e7b4a94f5008e5f0082d4a0bf2bd84279bb5a265ad6840354177f01ed74d36715f
z71f230015ee2313c09b1044ccc27d8c73c3fd51e5654722181d250e338f98cb85a684d30bc5280
zcee29ec18bcaf2ca6599015a5260a4ce1fd34f84544c78d285d626901f5f40257bdac3dc6f28e8
ze9bf80eedb4a4bf902206cdcee8543f9899f9d767efb07c0c3863225c49677ab8b516c53af4f27
z0e660dbac9ff481badc4f20f7e53bf30ccc4b55e22858214b9bd45c8fb243dfb69cd3171701b3b
z0234b67c920c6a77ec278f867bf33102b5d9ceb1e94daf0d25d6f8b5335d7e9e30a5cd018d3313
z9847d996f93f1c3e68266148a2516a41fbd196691eb1ca857346ff4d8991902fcfe8654f7d0ab2
z220070625240cbbdfe1f9879a625cd476801958b57ce460e0bdb44c1cc9d67916acad371ad35aa
zf6486d25ef1bd9ac29283ca77386e27fdfeee3f7d13145997b9f626509edac53e38300a66abec1
z8fabd7cb429da67f73144af973f8374ce6deca771bf32fc3c8bceb38ed05ef0a40a36cf397c390
zd87412c5a69494458856a7de07b6d492c7d52eba1909d59b4548ad1cf1411f5dfcb584e44532fd
zb3f42126557f4e4781805ad4cf433ad333fe0a93fb7ca297dab7b17c6aee3a0da69734ed0cd1a9
zff614ca9a8ebb6715ecf3f226b0cff766e44404a6d32271e5d9d2d318a90584622b8e3beb9ac25
za935b03bb0b4aa275390eb0c33396bdebacd146f8397bfef61176ff6458e0ef37c0412fbb09a18
z0c8a390113ccf14d62381897b10f75b7a59e26b5c2a5a1a14af42863e0b62d052505c2b6b540d0
z2f4aafa4d7e6b27e661573ff68d5b881046f702d1dcbc5a6544eae8b830c05f4a299759a2957dc
zd83cad023ef6d22548136700326c898c2f319c9034e400bfbba6a64f0b2e6de2a3a83ded648066
z0c1772aeffedf8c402708ce46ea4756d705c690a34f2f120a5bf41246a363944860f602b957d90
z0ec58041d8519bce51fe6943417f51a2796498e7d925e18b3ffd7d95661618431702aeb5f6721d
zd9f89c7cc5f37db668ed5cf595775dc423367de39badc5150c5df921d7249fa535fe829810641f
z6951ef30a96050cff7d55ecc51ac24a79b79b1b8d59c39be5e1a856ef48ef78c16034dce093bde
z74d687a83455d288a0e33b063ea62ccbb67f82455c277f50a7f0c91ca54aacfd91a06e5d14f0c0
z333d01d5a99840a3efc17c2b7d5d83eaa24fd278ae3fba6126ebb65bd5bd17b74031e939a3dce0
z093b73eca4686d9b40594b3c43fe37708397fb40f820a22cd73408cde22d877fbd499ad36e5211
zd3dadc9c530e7020064c4424544fd047262731fedc4eff5df4750bdf18edc8a526f84ff98395a8
z8826ad4cd86d4a24a7cfceb018e256a6d758a6873c46429e8f0c78dcce313e5659d798f71a5c54
zd9bd4225be2d667eae0829c6f65b0b201bf092c405b640d9fb25093133b527f206b06b6ab5edcf
zef1dd7bc16870dc858511e5eea303f8f6258660fbc03e4309db168af2b0874ba41df45e60c208b
zd91a805dad00db2e46c7a20200305a7a65e91269400d42f2211dce22bc742b2941f982ea6ad36f
z2ac0cfb7d050a610e19034cae0bc0a0aaab0ba5468a6674958e5ed92c980b0970f5bbed589993a
z0509b9d6f6394d01e3b374c58f04c87b23f0209b43712a9387611db103f9c088408476adbe27ab
zcded2e3d835f523229486ddff85c23cc288c07ee34c3aab9b96dbe74f7f6bffb9982e121eeacb7
ze6cc0f71b0c0b518c1ced5fe36429bc5181e7b0e0031e5a6c303420b399ee81a565c949fe00f57
zcbaca9854d277237b7eb58373e4271120bc49c99457de2b2ffb8f49685637d98da63ed5e41bb15
z5d7f6ebbe1bca314ea5925505c58093c02b030bf944d8e0f437a5d625923fa05496531faf6c56d
z3aa0eed66d3d52119abadacbe156e71144c4d94552ffc177cab0f36f193271fe1adadeb98d28d2
zbadab462e21435268d33900ce965db0b0742ed94ee40f963c90ec468ccf867d4e8214006603283
zdb67ec3df8c80ca512f659d1c8f5cfb78003ee89ef4571b767f735a34d6790ffc5dbedcc83b0ad
zb624661f6bab0599eb365ec85dd6539d4b38f7973b88b5af68faa5763648661ec6beaa5b34f507
z8adc848aa89e098593360542d7b528e3c8722a77d812487aba3fab103d4b717269fec59861a408
ze06492f14d037d6d38f36236122428086d3bc24339e67b4c9d355047c6b33483dbff958487c070
z148ce3367efe4346fc41ece7c5e2334df7be982e0fa1a26f895025b87708356390d06244ffc7e6
z25523c9222bfe65220b0cce75049bb35ffdaa41c29f4db355cc0a78136e56fa20800bcf59f96ff
zc1ee5a4cc3642f65e0973e9d932892885b89ab346888503fca87673fe3cee599f357e43980091e
zc849b21aea4b85c4d1afacb3bb5332ec375980756cad3c1c04253d026ac6a344574a729ffead69
ze9dbef3e90bce9394dcd0b05bd98db8d2e953f0313c826fc34fcc927e586ae612128daf019feae
z3e3bb0b9b7c38d2c5d873c176d67b21b70c4c97fdfa7ccf622f6635ee68e684b69fe8a191ac692
z768a380a55ce3daa6650eb1a1b2409a65a4db5bf28e780207e66e095c90b48e74e0924d11cf5a4
z0cf7b62b71d264755e7bb5f181cd73dafbda437bc9c8e8e91694e7121aa39ad6007555d3e95933
z02969d52e22ff17ff30a429aba7b81b95fa806ec0edb95fb37e13091810afa5852498cf60af728
z89814dab8f3e19aa068540a4d7ac761b8d48da6bd163a629d1f2c808566d512c69f855f2ccb348
z16ad3432fc7468828037283437e8108755511072f489700c66288f8a3fd3df45e490b5f8a4c665
zcac9934671fc4cc1be89af87b3af8f1bd5f58c2849a8707bbf91b23b86ff72a1766f2fbbe48c4c
z664397ed18d88fc739df8245fef32db118bc8a65eb36c9cf76bb94aa19fd008ef97c629c6682fe
ze7546b5ad148d56b44c1e9fcf052f04d717ffad57a297d340d693c9bdbf5078fa375d44fa6776c
zb4a302c096ed4379f066567cd919773a03e11bf7d9317f08b4c52137ef0f56eb0d2325bca2f35d
zd990cddc192e1a708fdfb90f07697cd33eba89960ef199921aee698ad63e679ab68f0088ae6023
z36ea4e446c0885dbafdb465f29772166071eaf40da54e1f4f6e8a1372a81ada59d4b5e7ec77e82
zbe0cac643e07b1985bd7d283265959681ec0f19e0ed36e88b5efd4413ab9493ac5b7363680e9d3
zdac367aa37251186cd6837519788baf36aa27914a5bbf8e7741d98eaffce7bf4d99be9add22fed
zfad802bc3d410511bfebdc05b1d1be61a495b011d41f45c4cf2ce8426f202adda913486a102cc9
zfee9bdba71aa5694838a67aa0eeabd8bd52b810b99c8a2f863f780e424db76ed71c2734606f6d4
z8036e270855032686b30701bddc6e870d4c53b4538ae8c361a310ff08d1f94171fb6290c607c8a
zdb8f1ceb5b34ad2d30d387a9db038bbe9099565e650cb418a3a374fc4104c5fad74c4adad1062a
z3cd547c8abe760a407b2bf73c5e13f77847e038c0fcffee93b6ea6b8048e23b9fb819685a06069
zb6d35fe867ffc9892cbc6b843ce0195efdb6752e9ac8c87819dcb50e9c98174c4bc5943ef8ba96
z95632286a4d5d92649a38afed3819102f78ac75affd6763806f3fcf9b2555e6b365df2ca2c9d3f
za5ec0e81b55158df1469f447ccd4a1c254d210b8f8a58baf74a8200a4f7bac340a905667b4f8e2
z5eb565f59f7769210da514d70585d32eeffda92242deb627d5ffb57ea1a2b837077bb4aeeb6613
z022ff27fc57f715b5230339fc04d2fba67c516c30f74c48ae7daa41a42411d33ab7ed15dc25d32
zc2093265e70ea5b697969ef067b7fdf9add1e73545f493b6fadfb7a6e7bb18b2bf287704b9722d
z7d9388d4b75582d7e1cf2dd0f91ac3bb3bdfc72b1ba10cd19756218285ba7950f05c3a79d41daf
z36cb2a57e945534f1667a14f7481ded92a691c6230cf5837b4292803deb99ad0f2384eefaba04e
z88a4dcb386a5a6244620082aa96ae435dda7f44026a3b285afcddbebeabdc584ceee5f473ba98d
z26a6083a030ee311cb18c34ee7f0d47c8d7e47a4688cb8589ae1ed755c403eadd84337d7553522
z45fdf1c3fc665376719ba3e8ee4ff51ec5b4b18cbd2ffb9a48e5336fe5ebaa9c89f8b449b682d2
zecd07fdde6c5fa8f6b3a72438bda14269cc656022a75403bd10ce4ce07214837590555495fba98
z4ceae5c33d5b1f8327808d7626a477be70d89b723713eb4126c7eabc7b4180d9309ebb0fac3807
z8105f56e621446969705c0787816f1876d993ef9c3b396543dde880f858adb96d3a8731bf3a73d
zdfa12fc6ba45b79d75fe2135c44eb6acae1b883496efbaa9e195fe72aa457246de6d088807075a
zc67b58fd8edc52544f3a0b60ada4ddb68c4f837f73c766c0bb00a58b9c5bdd2e2fd1d36aac3209
z3e9d7e01f2790fd46a4eb338d7ba4e297473616aca518a54275e23abcd0697f51bde70e6a990a4
z90e1b06ca2252e414326a791ccf93fbccbf518192bf8132943cea57ca7cd39ff6ab4b05d472bca
z2794a718c81403cdfc8ce297ec9074921291f3709dee5291025657bef978de561b745119f772cf
z3938818555a31dff8455aa48c7b8cde34d3857d20b1a95137bc99512d9aea8c38788d0b6fdc8fa
z99aeaa8d967cff22e6d73bd6ca4e77c5c2b3c7e4273108df9ddb8cfe6a19d5082675f8542eb172
z71013cb8854ce3c7855de464b6e45852987622839eb43ab77bfaeb4643b49937af16a2efc05880
z9319907206452e45026af8dae8fd40273c9fa670420695eddfbc66dc3e0b3ac6cab455e3bcbea9
z85e61dd26944774cea5cbcd0b670e0119dec650b47de86bac4063c6e0b4326e46dedc70a9a206c
zb9fb4b4a02e6cf3b989c0147316ed967a5adcb468d6edf54f92c2a6c9c6a0d82b4434de4f257f3
z12a1780cb905d195704114e8f491fa1c6693f9c49cf9460e00143c106ddee16fc146a259abbbf4
zcb8068cae38aebf8553caa3b382b46bf5d547e3399ff38812514e3533b42c163cb2bda8f2e0512
zc572a51d629d01cff7ea9f112f2b1fde2f6fd7a5bba744fb47d7aefbc37c39a00b72f7d6f871ac
z2b3e60fa34355d40eabdac978f0fe5f934f803cbfaa6d47c5a4763e86a21268f6e1a79e9cddbc8
zfce54dffa0a6ba4c4cf0993585f6734c0d7cccff33ccbd610c911a08a649f73be5ed795c51cc30
z73eb137147e40e0a5f8070449d4af0bfad03e1e13c62bb997d6eb211933785f4af80e1b1d7e7ef
zd08e09dd8435586bfa339625010790bbaff62c8d3e85cbb69ddc3f12e42fe6f00c09b6da6a5f34
z3b6d9bdadd61339d559bed2a5b8ee8486baa31cc82be8a17b3629dab6cacde49db136773ae6875
z603ce4ca8efd1aae7bd5dd213c31f150f31da25c549ba765a39b02296a5b5b68ad6fcfbb6de847
z1d020d4a12c5895e97362de2d480b608f6f7733f3d60bd16842d719d7d79a7340503bdc3e2e995
z5b671786014a95e3e4a24e1976ff1d7f7d4bf0851d08cd7fd626ba0f09e5f728ce2a4f33e17663
zf3a55176b9ac149e376d4f714610b072dc5920d8eb53c2484170f7a5b4db07e474d3b3312dbf44
ze5dca19db9954a15304c9f2b3bab15b18a6edfbc6fa07329542432b86d61fbe16a8205fef6f8e1
zff26851c45e7fe5ebbf3a9b943675c26994b0d8730cb8bbf1c85b9a5e460269dbc01730ddabd89
z645c1a347031ba2c3a5558cc4d1c5523be4ef80fe00dedbe421fdb3c56b709189f48828cc6c654
z796742666eb8c8291025f0c1bf928c16ff751920f018a211f7da3108a33ec256efe0e0e7a06b05
z7d0d893581df427b5c0111a27ca24a0a9b2d298e0a3e6ba26fb2aad7cdfd2537603472cd1d692b
z8f99f85a2506c83ee568647f7a5fa571aee78149cd5b0c6402983f02ac2b188a465e7f7b682617
zfc0e4131683e4400380e3cb7abaf4d61f0b3f5b3a35361c01d092e9f8726b872a0476c3f5a4f7c
z3dc68a18df3873f1b37f385d87d7433b75de4b6f1e8112b5ebe88664a7ec10d612e5c2659fb5cd
zbada02eef40afa580f563bf193ac9c8046712bbb0b18d87ff703bb7e6c35553c61a5eb140213fc
zedf319c20a7c640e4fdb2f006339dc488f46992dc15a413c03765ed91b68f547f8440f4c320e1f
zf215008fb321263e8e38fb4a68d189eaa33c382079dda5ee40ecec6eb7e581bda9c58684875736
z2806e243b2845057d3a2744de5b47807cdfe60a84cf13c51af4eb9e92567ed52396cfd0c221aa9
z6a44e09c748d04f0157e40f6d532221b1fb2065efe80441d917ae04f5c86bb622ef2685681d664
zec54d6972cff474a69c5acaec73ce8b96e67fcf8729591b816a9a4456fa3d314d4c4354934ac39
z94af9f195977d9bcff8539315ea38b6f875478e70d856882c57651bd613260044abad0b2a0f144
z119d50fbf98d9561f218f3df11a55c07c2d0d2726b4cefbfca9f6309e6537827a56bb1ba4e1653
za4ff52a3209cb16a81152ddca7ee27208346573030f02510dbadb2b52048ad029558f67ec45b95
z20ec28f4820b5dac5a1b8d813cc08ce614d6057f50029ea677ddffced1297af6bddc2cfb3396f0
z6a8769756599202a9de336430720ec55f2bce3fd3746aedb252d5ee7153f1d5c8b112114e12670
z3a80b6f7e20239f801fd9cd44986b1a3b397e69402c873043d08bca11e39a234c78e5f976d5984
z840acb8d684a2d1e6199ead20a0f0fd8ae576c80b13310785d8692bf849984103cd82b7472bbcc
zead9e7ebfa1a3ea3fa5f5627d319b509db0c2470071614ebcf1d6664be9e84ec55784bc6414a80
zdbc716bc759273770b67fe673daa7c8d4f2f9413b9ef18a14fb580ccfdd09be36c965bff1609a4
z2e27e46c5999e4eedde0fb322f9b4ae4a12f06b494a982fef54dcd5a8be1ef8fd136a3fb7451d3
z91306dc4b121501ea304412a453bc5914f09375b6e008b91358182125e8a447b29ee56a9afe5ff
zaad4190fbd9c8255a211ae93b9eab475d008f734284b2157fe39f9e7c138c22d698f1f637182e6
ze385960f0a168b51babf8a242766d72c11883ab635ab51bf8e3cd1710e156a351a1d0e439cf268
zce4f475b3c80deeb1d3af41a5644a153a58671bb4df3e6fb7aed077fe80e7f296194fe5f123441
z5ef1dfa5518b9f79b59b59935858c239f9fd018bdfa61b7b530e9f12720ee6dd369afbbef7bbbe
z2b855f319a1d14a86ada8d3172831ccbf43785c4deee10aa72f19a61766f2e838302c8740317a2
z1cc5ff1b85c12f143b7f103a08e668f2e67d46c2985e9374326ab53ad40baf62eb61eafc6ef6dd
ze9045f76bd48a476d9bac1396c89dbd9f9eced8138d83ca5a0d07cec2e9f5203d7539e98b5db83
zc8bd7f89e78b1a2cca95522b4fab0dfe581a8365ae60882377bf1c5f338593cae26cb4b9e7b0e4
z1f245f3309038b83aeaa1aa755d3e0976466a42533dd5facbd399a0023be9a8370acbd14fa2a0b
z37ae756efec83d7e082d6271cb9a65f6a6e9e01b7eccc2dbf510abff361c894c4cc6b06f631252
z9ecd59db7147a2346564f37079600e8a9b960d459fc8e1546066cbbc897845d2fd134d8562ad08
zc1705af7b221fdc332d727a4c578a6d966c8ca2a5205dba17c9761b7cfff043c7b7e5399ff8bbd
z9faf6e27d3ff240e113fe4394d40ebfbc14a3ed6ec13f0f9d075cc606d8b5a63e23a98f5eb9910
z1d8cc2f121d29ca332cbec390352aaf85f7dbf33cbf82f567d82505c78ef651178af410c094e46
z7db01fec7e29a14f3fc590767874d6e052c9fd90372cbb027d5714d031e10f3afb9036800f17eb
z81402566e2536b1f8a2f8f5c991ba414706cb3daa8e85dc82d1084faf6d5d54aa3ab5516b93276
zedaea6548aa0af65e82caeab4d033f4e5bbbfa81809e8fb3522af2447c9b1586228d0a3d3509e5
za188de38e82737a7ec095eadb4e15e510d623a00bde92cf34a912186cf9bed3908ce953881cac8
z6acdfd7e1e75ded386e79235c118e0c4a8020e9525709f3664494c335c25e1cf8fadb2ea532481
zd027cc0aeccad4ef1068e47e987bb1f6914668bd2986fc23f94da65a7db018833a1b6b547ab656
z910920838354b2d2d6d2a592cea7ad37b3ee4efb3dc6791949ad563168bf13f41648786d86e0b3
zced7f65e4463f7ac861ec5febdee19d5d0e7c95ae8f323c6f577252aa95e6709a7e4e9b4aefcfb
za91a2a5298f811573bddf72060b1c74d7609a05ff59618f591328c253e71e87e203f8d7ff005a3
zf0871b7f55b0d883f04a311d4b31588509ac7f7bb019e2d15ec17be466f401ebfd2660ef807525
z2b4b7a0e2cb793063ec551b09517a387e9111fbb4ccebe8160dd8d84e9debce99c259907e68228
z98ba786da42c601ad60d50038264d5b670f23852154c31077f85ce9eaad0351db538130a674958
zb1f55c0d66885c0694088329ff20b626e2e4a6ef8ebfe5b9d08bdc68c6b86cf1f2503fd3a12a8e
zd4c9a792822ccce713decbd4152f0092d936bbbc99b2281e2e26ab53abd6111f2734bde2c7074f
z34015b359b33c414a38fd9dffab740fa240c0575bc097138d2d72ef7630824922e759ccdf50066
za984c6a25e89b0b10113431a1eaa39a88cb700a9a533bbec8a685136f055f7b140be4df4dddc76
z987280461ba1383c81888938d06a5a7c36fd05a4e580697e50aeea1d04048e5e0ec3e770183161
za1e5742bb237f3801174b1017d7e53910c494ce4a485c3442861e4d0dab35c58f68ac1aa747a74
zf127fd9b812c2fad71efa102db87f3838ab96891756fefd9cb656344ee38b1e349d47686e75c3a
z3954697c4526d0001f49011ed63239036d77dd18cb461582ec0d7fedba7fc5cec7aa3401394e61
z38c842a9982db928876c0d360a594b46d16154456af5579ccdcb666c5e4a3461facea2355a9e88
zf6245096adf7ddbb23b1114cad176713674064e040dca68465a6ce7189076aa0ad0a56945dfb29
z842695cf148ddcb607526702df0143243cfe7be1faf317479a7235451b79a6e72034248f2ad25b
z16b9d6ef57e65fac07b8b2e0f78710c2bceb7f510f61a1a2ebc956c30ac423521df8159e744416
z9769de7a94de143d39065219ffb8c5d1226ad276773a901b20bd949c911988607e565bdc33a792
ze29a23ef369b25b9381f68f77de5caf2f7a8ffbdee2594466d26cb02eb32e55ffaed049a54df55
z529828542b69f06e1f811d3b51aee1879353ea1469688aa1d99f07d4ea3196bf5415cd03db7ae5
z80cb9cd93ce53559e0856aa813dcace057391e779eb3ee6f9c7a17ae0534ae9270fd654de828a3
z53819dd30a0b58fb9929a6ccdec93be1166c501ef98ed69b5381bfa35d82d1567f97fb4419a946
zd7e1d0aa23de02293a08c3cb15cbfec83d6d0c8a7b3261fa16b9becc14ad6c178e390dba3b42a7
z141e76114dad91e1e76a8662c7cd983b3a28cda9a1a784436134a1c16878405bfd790d7cdf084c
z218f49e3e8b5233b8cc4fc9fcb4e55a17444ff2a58b5f08835cccb219100f6ddd4c258eff158f7
z48d9ea31c41988bb88b4a33a5a283117f87f54ed3e7712a87b26f861fb03972fa2974a5df5b6c7
z1a52643b51fb8f0250f12380c9a0c92e279c1e53ee0b28e333dd17556b5c8a4be38674afaa2136
z7f7e7e33cdaf89a6c18d7c2011ddd4d61379b66d671fae37d3b21151e38a51db2470c085b689a7
zf808f538c88ac29fadababf6679d403c95971d645fc3a0502cd726cb278e29d5e73a21c2ff977c
za8c6c6fb5111047ea6d39a1e00ef7b174b2b3bd27bde091a87d00cc3367886b81be77eda733e4e
z9c61f25def6359f6b19645d44ef50ec88b8bc93146328d63a621e20b87b12e28b75240f28f49a1
z3f3a441833d319e008446dcc64741c9517d251be2d48f0cd40211030d0712bad822cba8e5648f6
zd3cfd660e5992b271e58d412871310105a56dadacaa41dbc1ddd0cd53f36cc499e497fd4391955
zb17e5b0979df416ebfdfc6d1fd2e5918f0003ac7721291eb30d76ce5fc754fbfa90a05c4d3328d
zc4eb3012f8eff607de0e5c27d4449dce96686415caadd096a38e99ef0a173b8e7f77a157bca551
z393de12c2f865ec185c7ff7119f11287ab56737c991a74f45956187ee2f0606a9905a4fdcb102c
z7b437e9d918fca2b3d0af60dc1ab189bd9c0786ca629ce669d00fe6b6289aafdd7dbbddb8056bb
z3041b54ebc710db1ac8e6cb440eb6b71596fc4458c9f42cb238356110e67051bc15cfe5cbe0f92
z17bb3c06364c0e0000c9e51ef189b424a9e97564b4ed18cef194cae10a40aad41664b82128fd41
z4cea284b5a9ee51e95a3591a8d767307841c09cd3137f8eeea984b353f6c6da0d5bbaa6d6f2629
z8f8caa26542c515afb53c5dfd16cad3a4cceef4047105f7b94e942ee2c6df996ce4d7ff9c36a92
zf361e5a8c97673d745246891cd3c912eb2baf747139aff805d6bf6f3cb18e525e0c318895dc014
zd3f42091a204832f0ec3e1f9ee4113182510eb875171e291257e2da68b63c3cf4ca4ee4d8e073d
ze6dc08c17553abee3398d8671ba2fb4d4718a994037d14efa3a8fc95d9d35c20190a8b35d214b5
z2e948bec7bd5697467d7c370f9d06fea3dd6d1b23a3c50e9bd75219d29111d5a989ddfb44e1826
zb9abcdb9bbe2f262fba5a803ffd5956114d2018942c0c7b8a5814f453cd237c14869722efd596d
zca76fcdaa0c2870902d3bc28091fd558d92ebe84e0d0bdf4598f01f2fec87f28221d69194d96dc
zecc06eb74d14c91fe2d719e8467291ac74bb72a7d5a80fe19857f380477f8ab6f18cc6c3a79247
z88deba326be62f4ab44b3a41930cff55a6892de26c45c67712e2b9ec2c8704f23f04c05d192ddd
za8f024f5a78389904e71aa19b4a132271169ac971f60371636a150b9be65133f7d7ab0e7d28fa3
z4ca89afa97a52b23863ede6cca6689a6041e388ce49ee54cbae7f42f49c794fa72aca6451b277f
ze98601f6eb786da5bf391468621213e896662acb130d1e37d1628b08bddbbff99c5d44ef176176
z703ac81524078743d10cbea4a726324ff03438e8746f2173feeb6ba34d314be5888a7f5c431a52
z0d13fb9e7fe2f62c68747bb74de80e3ac14c7c2b4b733ecd5699cc4f43c5577489c021f842af03
zb30e439d586095f42f5d2192413861b5becd104fcda401dfb076ce0995eebebb095dd95531b9cd
z764f7b4b306313c500a646fde618bce92e81e19aabbd043cf90c63e6c6428987e36e8d47b172a2
zbc73a53143402fe8dd961e575fc139669c9d4c7f10138a0e37467c0983e135e4a500b777e6f46b
z2489f9a3ced98ca40ebcfed84041d30b129c3d2e8430dbd69436d3a9efc065d3acb3f9b47891b0
zfd9166c6762911f8c92b5347f51832e1dfc0e2cb2432f13fb1f601923ae23c3bef7c135144869f
z3d01b842073e85228beb872d5463006e32d2baf6caf15e340d26171fd5a8e3f8240b66717034b8
z1fc66fa2cb7853d29c10ce847a809b270ab479f0a3795c4354d73aa998fa226b38ab057156c1bd
za9b7f125224c378172f432324e3debc17cafdf7c04a46f37c1e749f19bd661a1d5ad37e9c95109
z44a46e755972abca720032f85f41ed70c73e0a3c8cdefe66ba9526fd43b76b37dc4d5fdd76ba68
z7ded976a388f6759f84570dd8c5bb5a926ef6beb431de85c80c32622fe4e80f1e1ad14674a2e93
z81acd82eb5c399249bde5926eb76e5cfd89e870db56ec75aab8f433acec041971f87ae7dc46d44
z7fc4e1f11d27c5447f740b122064ada907496ddbf8981d6639e9004a922be01d8d6679f05f8661
zac565d05a3f54b27ea9dc696979d9cad7c5136c315f034dcd9f8eb1189e93014652ff3e798a5a6
z1202721ce7b0882fccd8202e52d5f6c27ccc2c6908c91fa5ef2a1c5147617bc515f26731c7d7d3
za671e12d4dee89b21f0255de08131a59405dd6b86249d4284fb284eda5d4c0270abb16649390f9
z279f0c411decdd3117fd9ac83f73c67097ca00ac8f1239e4d0c075ef85b7a33f4c2bb7907a20c9
zb1e9cba3f4aed517e1e151daa7f6d90adb8019b391ab000d74967d4959f179c4e150b76d2946e0
zf0bb915f15d1745da10bacf4b052856dd729e3f1453a2cc64ac2e61a8fb06c6a7f94064d51dfff
ze7c24ad51109a6ed5ded25592dafdbca5b551b79858e0c3b5dbbf7585db4f35df0fbf86c1fa5ab
z627d87be329cad3bd53cd6b800f1c9c2841c2e922a99a7e28a8af18494db59a0ca47ea2cadc0d8
z4250c4d38c3f3d483b91122a3529d269f646147e850e2c569e86bbc513a4882feee3050e7e2e8e
z96183084bcfc4b839dca95ffa19ae27bb7b9017ba30314fda8e0d2804b882bcf0562485458b5f4
zfa27fd3c62cf69c4bc67489e2c2395e909823a9e1e6f0d18513432f03ddd8a176c2f886a13c24d
z614e04718f7a121d31177e735a466ebe49ffe03e7e50137b4190f4448d6a18b061709a5959c0f9
z10000254f48a9cca69b9530006fc94bce4eb39ddf9fac1262ef63ebd8c8e0dbef7c119ff397b8e
z9f939906696b0b500ce850eb825b7edf7860ae652760192f4105f4281a67d244d175f4a173fc18
z07dd9e5082de7ad79caafa630644c5095ff5b82a39331b3bbfc62e1a1a044afa4b7855c2c4031f
za03f3b80724c3ded099d2c0a9d274e5665d74de74d2c5aa028d2e07c0e7c1dfce05c8eae339603
z449ccf1ee473f2c4d03e0c80342f0022333acc5403f67c6390ec1ac722d08c1337e5a148fc0304
zc2071679e8cb156ce05dfcf17c26326bb360fe27f58d1fe11d4b3d78162cb8f5cd8b25967f6509
z0fd2f0d7ad3a7cab9312db2c8a635bd6ff3f3c8f7071dbac90ae1a878f7fe8c937469cefe6224a
z16c8a4b33fe29e8c457b1817c8874a882448b3f8cb7de5c646b14c3b6dac7ed9d59cd41417019c
ze7fe86f35f1a384529bd2447fa7a0ec1a22f9a663dea92f985702841b64633121d87f12896b126
z8bbca43c3f59b40fee2ca08f937fb594814f2ea35c3d8c6e8a8701e854ce7d10bb884bc3473958
zff12c68d2623b46cdeb9ecbad40735fb3bd761eed7e3234f0a78b653143a2280095db77c131083
z811919bb6e099eaf3a869d667a881c4551492a8085d07e4529da41c1425620f45adc6c521960ff
ze34e696c4114eaf84eb43ea8d3284ff927d6b309c5c97b3dacb3cbc68a642d4ddd7bf2a8f3a968
z744307e88f88e43bdeb67212cc3e1918f88b65870f4977dbcaad162bc0c6ee00211e3ef2f7a3c5
z406295c9258396187ea4e404a83ef03e157d16745577012286415161f2080f9894a00590a7690c
z20635fa6137d0d95ee3a30121a36918debb309f097a37880491a94ff9f85863f568d7474ada641
z3f06f05b6528941cd4e45c8a862c33c7bdfc3c983a66714614feed5687085ce88007da607a1244
z73c9d00acc2493b9d36a11b72e20a8dac845813447259282f0b6f559d43ffcdb73eb555c8e1652
z61150a61ec40c7ca7841dcaedc3f6d5edc6c9ee4fb837a72e4cc76ca02f5d814fa0dbf9711648d
z6ab70b887373374f8f801e144111c4977983242678ede29e9923a2dd024bfe3f81eccb5c5d891e
zdb0b5586d8ceef0387202666f17285c0f344b9a0ec4e6b085fa2ab3fb47115bed3c23fc23a1ddd
zb5991fd60cd2a70e4c9abe699e6c91289e9c19e610d2d16e2ecb613dd3ac65608e82749edf1151
zd2f07300657a8032d23b70ab78f8932965da39e9b24f4f50ceaa110e58e8b5cbc2fe55f736fe29
zd8392f6fd01ff0831b1e74bb09859590994df427a38545d9c414c0ab973c30b5dc3a364feab831
z9300368d98d0de10564d1622ac864de3f3ee6b3437269ddbc0c0593a0fd865a061fe6c24d9c975
z2f41fb57ca9406295155588d97b153ff54e138f8835648944cf25e14cb7e2d467287ffef79e017
za7e1c1d56bb686917301de3623f2dd26c26a07784cb78acba88f2b4772465291fbb377411b4d3e
z0b2a525208e8effe082e665c84b9239ac070ba525f737d9797c6be4504bd3397e4dc0e0690e8a4
za89043d44ded890888ce2b7b69efdd73931163fbf6012965f4c5a82508ba6b09920694611b9585
z3105d6fbafaeecc25b3ca0c33512cca6d78d7c3e8abab186d9f8f4625204adda219151dae47452
z2ed9ba29900eeb0c5b94121ab75a2e9bbef9876bee7098da1ae7ce92c6c3dc90affb43cea664f8
z1b842f8bb2470e7bb18c7afebae6abd8ad3781064e5bbe5de1572c94f20781340654d5614e862e
z75a957913c3e3c06c1e7c0ce03df30f0c3b2f621ed87fca687210b8bacc2d4e5d0a8c321032d77
zb6d09751d3355837a3f122996bcbd686d56f2d0744f9bd34992ca48de4887d34652c2603c0d82f
z4e323e831d4f7d00b5ea6b4fa4951f3b177543e2589ddf92866103462d722bf2fe5a6f2381916a
zf3fbc92bf127fc9afc777b0bba1d61699652162a15d6639e5980e3505876c19771d72fe634b9ce
z037a7c358fac989dbdfaeb2a7618b80f86e1ba58f9b73987f68ef2b5bbc6bc44e9a3541bafec91
zb46db077ca53bcc893dd15ae9ab8254b49addf68c93b634a7f35a06f57b7bee43b4c26712f03d2
z291139eca21277394ccbc780e76b3289ba60cc97fd7e8d8c8370646fc53d709cbfd108a3c76284
z2d76600639d871e7127b949282be8683e3cfba02cea5a5bc6a75416b77d41f5fe2dd029494ca54
z268528b1f5902001c70e2870adfd68b67461836ac2cff19f595f66ae82d67586e4bee048095039
z9953294bc7f1df82364d43d0a2c42a49f889855f4d11575348eead0e21a0e79788eb916178919f
z6d83ce170c4788c4f32188841ff5a84ed35f2348f1bee6ee077097d6fd0bd3f54defe75bc2a5b5
z698dae07a656cb14acfb1d65d2d21f218bb61a0f05203e7b27119dbacadc7423a61ec910e94756
z08b73a30c781eb6f82f6c4e5edfd6c80669d758e8567669375c954098bd044f118332770da5982
zc44d1f06c9a0b025f3013a385ad5cbf59a075bff1574366d13b483204d7eea1b59222f0a920cbd
z2271e3b279f54fca1b388ed97c567a05954f3e88835d46ac93093eb4ce4d943fd4d4cd2220ced8
zd5073d18869da6171de4ce3d087dbdca4aa2edf656f3f016404723097eaedd6e53fa2dc7c6ac9a
zc64a5e74bef94b618f94c587f5824144baf557ae927d8ef7df0a72767083fe0bb75a90f22d8630
ze4bb9c5f0a321c189b5c2bb8b14f87aa9c7f82c7b17924e55d8f23abfca8bbf0b2c1fa5337cdaf
zb1d057583cd2ec0ccd9d4d8b537c636ae7c2a359b613c026749e71349634b6cecf0b7b30e593d4
z45510f684c447069b4f9982f7ad288ba842a88ae9e0152982ea9cb8b7e318824b597432546b698
zfe93598a4945515fd3c18d6fc8733a8500b0d8f140ecb0871f77604758506d3335a3ffe22c4fa8
z8f89d021e7e79318cf30ea143b0650fc57d6f5964671e1eb72520b4709f8a343eef1cca4863127
z8b84a8651531d2853a1e0635ea395b8734d6695ddedb42449ab3e459b60f3f06c1cd08265ac838
zdfe5f823aace5a312af72a166856e9b7261afb835c9b952fb01619cc0ac481bbfc230f43f0e016
zaa4fd5ed7680ee035643ab4f8fe0d77a471715100789df7810a8ea2793af6de6bed9f18121942e
z3415578af7d88b9e87dbc795465f8928bcf21d239ef15cb25a3f54e0166242c8f9e72a7d506d48
z0323a8f60139b5034d9b1186c4c5f3e52a0ce0affd80356b697be6ff48f22e414a251a3c92861b
zd783e38e3ad5343346b286f7d7fe2e0baa5abf6164ebc0b0af7dcb3e8a10531cad4579193fa303
z19fc12677280981174d6c9e1f746aa2c34c220b8a6f6366712a0fef4527430623754d4a8519197
z811764d0a2fe75a2c84229d0764e419fe8487484716daf3ebfa5c9c7097b320edb230be327dfbc
z1c15b33a8a2bea8ff3b4827dd205d99594cb2631fd37541734715b0b5f06e236bcf57d80bc0db6
zbc18acd1ec32add4912dc85117cb044e69c358768b723a043cf7c5bd12fed5a67e538271492049
zf0cd6776ce1b4b15214357a7d9a190b6725a8f5851c73714c6290426f040fbc4cdad564e751e2b
z6f2615e9120854ef4bbdb9da0ed0bc1d7bbca425d9505f40533240ae7d55221fc27ec25f4e3725
z78c3981d20d5568bb370e633f632bccb8a9367f501512910d38ef9b5c764dae2b3a84c8ab6b064
z0d7c408bbfb0ba978723fabfc7f91a83ec246ef4efda5b0c6fb806754452c123365cc392c126cc
z00ba367e66122812e35f99e4adc2ecff6523a205846c7efc57674b3a3391ffb671332f48ef85eb
zc2d0d7412f6c429c137ed05c185826c12b899ca2eb2ec6e88a634cf918565e119ca21d624d3f92
z2f411afa8034a8193cafe1d1cd4d142020f0679415a0542ee5f95b440468cea1b1745c67e11321
z71471d98f9677bd78c04c9e091759a5d740addd51040df56af6c212498cee8e50f7f86444330c5
zc8584e7c1e4848d47ed3b95579ddc5d6eb68d3decb8e787aa4c4579b3987d28a720c408a05c348
zf53b450c1ca7b3b00b804eb79e8ededc93d0504b4419e5206ba48a8c1e3c2ebf1027c0ef9b1a65
z1f93686b7b09ea077018bf69a861027614da10626521d839416bdbfe7cb7c7f8c4c1c03ce53c9b
z99030a46c0f03f2fce0e54d54127dee772755ac089f6a0811e7bfe43f36ef03487d8efcdcc8c6c
zf038dce910ef8064f2fd07334360139ae772d32ba4aada519ac9c534b8155ab044d58f605c5e94
zaacd7fbc3f10f7b4eb31621d5b027a66c591f45ed99e9d9ee643ac1304d98c57aafddc03393bae
zcf21b5b722a7d4d841b368c0dc599c4c9fc1af6d066d7d2eb0f9847376d9b4a2ad06a1e5cba371
z22d60223ab5a3f023620f8598eb653e75b541620dc589282e3b1ee17a2a0cd62a525972e2b53a1
z2fef1190d97e5b183ca733a3db725183ddefb43481ea1d9099b61d9abb0d92753728cb7cfdadaf
zbb1b24b0d9dba9f7bd13edebb6c514bb03a9627262e3098422b20b6f0573849c13afaa167fa0df
z6e71a321fdeeead3f66a70f30b9db92bc8e153e714d61c0e1d89e643cfc2b98208ff711d4b312f
z28c0fb847f9f4328d99d5210bf73d15f98fced170312c76bd057ecda5db6b070ba039f4f08f090
z4793b43b76513f89d17487582547be67a4c4a45c971fdadaf0fa1793453303beaedf0ebf4c3e28
zed6ea31c838e4d56dee68095e84057d0acd9ac24857d479bb106fd3bd7949ef4c491014873bb70
z362699f2b0afbf83b27e9ef26e8d6025164026193ebee7d072881ab15a954a98aa4d5a4b50ebf3
zdb7ca40c2861f9488443cf9607c5dc92110b3dc31e6134b1d5ed5ce89dabea20ca7bfa6df1d8bf
z1ce4df330ce061a850c67f648c6efa04858604fd588d1317d4abf678eda2f09fa2e723e41c5823
zded100ae3c02981773372f537d476e8f08a6952ca315b78041ce8614971843640dcb578d70bec6
zb93e7a3231d09ce34f982e077e74a62538f69d8fed7a29a6e65a67f5a6513c66cb111a64379d59
z5d0ca6f38dc7b9166a3b1bdc628a0a0cc5b7fbae7c665da7da426beaff431d27398370c144f3e7
zeba547626027c356879ccee7d3158d0cb15a32d2c92f615c73a30856466730507f6f47af0a20b0
z52dbf70b038be97ba66786ee5bf86effb4c495c943272d94485656895b30f63d3953bd2f36d408
z118c820e402329e5b81ba51feec1273a701371fb7d9e629f1d67b7f778659351715a826c2e8440
za114bdb589d0cbd3d4e65a9e18a46fcc01555e00a547312c283333f6a4ce3c1f0e225f8043b458
z41d64576c9e76ce31219420cb33fca272387e97cf90e022b03e8b553b412c8d2fa4b42a7d04661
ze54043e5405099ce9e7d1273b4bfcee2c1e4f679df8b637aa45a0f06af12974ea3b00a0ad4fdf5
zb87dddc4b6157cf739dba72ef65fe7352ccb37c2e515e38767770616b0f43afbbd350405f5157f
zf8f6ce777327de37e107c32bfec15819e2e3eb7a9b9b3a5f3c345d06d30a2f0d67fc36fcc95b24
zcc99c2e8f5027ccff2ce794515493d50c07ff77e530241651394b501e61b96d28ac2f055a6d40e
z137a710f55dfce2f9728c6617fdb2339d74808d65e55706348c91393bf5aec385fe152f34c6286
zfdb5093dae1768b213d09fc39a23871569a534143b9c09f95b8ba07e1c09aff8d56cb734528b11
zebcc3962c7781aa2faecd96366b307c85b4c2238e4cc365fe76d8f4601150a00591e78002f0018
z2b0a645edb44bd73b2e34d94a183a823ce9b86706644300d0db59d6b70dbf09cf0362f2a887a67
zc6d7546163dbdd793f79abbab068080abb1ed0a71cb492f980eeea44121e084d4289ed49b6be34
zbc49b3d2d083c04e188d91d1e2fac7cd9c3df684fd22a653a2d49e96dadee4cb578ec1992d64ec
zea0efa176ece418afdc2f9ab3cf57c5395cadd1929da35e185cff1f7c7721d11aefb7efe1d7658
z8308a7bbab38a1cfdcccc3963e469c165f2e78c13a10941f6af0ccba8e74d150cd017bc015fede
z1899b4c9047526ba29a6912abc146afeaae85e402cd78f82e309953a0a7ddcad59e9f5e3904cc3
zfc0890fdd02a6da76868a209fa451f24cacbc4e11fd534a0a52f296c1d68196f37c81bde4eabf2
z4063822e57287d05534a7f52b6fbd7c576198d63dcefa79a347608ab46700959f69212f64a4e35
z6378c58063f4f81f496cf015946740e5c8224f9edbff776732618b8674678cb16e6fd8160383bb
zffc883ae27cf192edf7ffd36c715a5c8840b722ba20cfd5bf0e6b1362ced988ec684c2b7e58ee2
z703cd70dbab77d3718d504b754f75e90c875eeabad8eb7ca17f17c4dcb4f6059d243a066dd2e32
z4ce32faab1f110eae83a2bd98e48396e1c9cf81ab1b371ec9c145733ba8ee07652d73297169c3e
z771c3a076915bf1f5ec6481f8520eddfe5de16dbd22ad25c393fe3ff889f50a949c3e23f6908de
z2a313ed4ebd0aef60369ea25cbd024964745840667563f5afaf3dc83be1320d6a0d29bfce89546
z155c5e0b2f7e2e4fff33df42c83231e0c2b59cfbca1b85d414aa805133665933b29b871c923601
zf75aab1645e9a48c14d223ede33ab2df3033aee4616c501e8feb6818809b338d88d791e34c0d95
z447ddab7b9b9fdfb119b748f1b4a409a9fbfadf0565c8db7c961fa5fd7ceaf6d8f19e8cb70aabb
z114a103ab7cb75e67983e96f0e438503633aabd6c3869c74f823f48649b892445b46c8d1cf165e
za85ec70a03908e1607c8949854e4903aeda5f4f90552745efd20798eb10661fcf21a0ea26ad9fa
z340f1af01bba20d32b957875cf3402f3512ec25e08b86f2e6af4ff19075cd74ff255be93396d95
z9c217685482fe5b072268876cc97be67523cea6fc4f36104dfd0ecae6ca213c0d57822891769bf
zd447ab68c91b2941e6f65fbcedf9a89228674afb0deb01dc5bcc41e764d64de29fa1cbc1a82e7e
z2a67f39bf4272f2cc80fd2f686becf0a748b0e57cf90acb8152185d81fe70f5270a5f3c4fa7ef7
z13f262a59bc496f5c71d2327a98c251d239a2817841431ff1546655fa2531f094fd309546f8b15
za89a79e1587bf1bd8f4f640b343164d3a639dc79a1a1a1d3e4306127df35daccc7106c89426754
za33ed0192b1fb5786297a74f61fb2231ab7de3afcc1d4bde5e70b6fd0edd2c62c5fa88a650808e
zb1034946593ce4d68c44c9b2f2fc5522a47ea29c088be51faa5eb3c5b9099232f97ea40265952a
zc30693279d5594607ea68c092e05bdc02b6cc5f5c81976a09caa71f018a6709e215d69141a7a2c
z068135e75f3609d9f779feea6f0036ca1d6b59baaebead0bb37b6d4da49b151a154d1896a84718
z804d98c58e05506d942aeefdf6d00bef24c1c407a2d88fd7f5d7c5e30f3ed39ceb0c25a2e16a39
z6dfdd80b0f6567c2abf885bb5296241d4c625e9838b67d909d20458265e087833646128570a931
z7953583073e10ca8d2df989a41ad1c5a4c537578c42f7498574a6cea47171e3bd01a8286ab12ba
z06da9a84ec86eeb95c08baeff209f1f495d3cde79519c6ebc094e5491e061aae45a5ad7e3d951e
z7eb734cb2200eda64caba5bd95dbff7e1bac31b2125cae641e3f9a44c29f9198ca04ab5e7bd85c
ze6b89aa972524dde0a4b19ac2497ef4ed0675d3c95e1a7007314ca562ccf5b849c9ffba57a433e
za176bc0d68bd914de988af616fea3a5c2e83a6898f9173aff43bbd3d24eddf79dadfc314b94ca7
z028d0b67986e8ffde22961217cc8117bf7ed01c35d59e88a544eb09ba538c233b1cfc8f7c68b01
z98091dd45f5392f8e6e8147a0bacb329382375e586a4786f0f40ca1bf61ca7e462e3028e58da52
zc6a7cb1e107ec32af252dfcc365bf0e1ad02c2a6cd9fbb2fd2c3d267a9ac0389518d66bf93d72f
z723504422bfda040a14744e2aa4ecec195fcf7ad7f9f1d1d5d947d00d2c9244d50696d1e5de47a
z67111be1a0f63ad41411cae5301ad3eac59fef1dc6fb8d3becddb86a39cd34b5eaaa175a1dfc73
z80975a52439806cfb55550d78bce6ecbf10842b2324452934aacf981aefa4327fcf7582eeebb5a
z589460352ae73225dad78bdd53e1c03f807c95fddb5725ad6a22b9cd49ec0c6526921e5f94bec6
z1d16236e1a7a74552fe32fa588d4507a2a0c4a001ee78617c1ffe1ea4fb013fc582159e84ce4a3
zd34da057f76727bf012ba6cff3120a3d5638f8a0a75d41dd243ff87a77343f38457f76b65c1501
z3bda71e675842be4f914777522276b83f158e9ddac53b6f90c8f0ab86f8085fd90ab9a878e9d87
z5b6ac701a59d0f830b722e0e28a8f5055b866816469b4affd6d17d12c8ab1e2dc2b29e4c2743db
z0adf10a642e00867857bc109c368b92ced7f441517eaca2a9e2239c27ef07c0812adfb18a2ba1f
z09ec41252c5cddde27de0cd33c4bb73ebc97c44f531c75661dafbaa606cd0cfcd1917e1e11096e
zb633573460e4cfabd11b72f70439dba3d283be12ed28d39dfcde9da430ebdf00538b8443149a73
zf97ee2feffdbcbfb4466ae3b8774453b9713199446cd3384bf1a1e4c2736f479a4b47db68811cb
z59c946059590665bfbba969c63e15e88d6dec326921595fc754c2f45c73269d29b806c84040762
za803bea0b92591cf4d7d8d2777f1f466b29bae1c1a31b876b052cd51b784e5de27552e4d09c9a8
zd70be93fdc85b2d4c3d352be5c648b142c0b455a0eeeadf63fa92c927c424d10cfc5716fc3dcb4
zb3867a307a94b25b278f0fda88c55727d0890cfb841b67deb0c66d66a082b65cc050fe18fc8b19
z8d7eac704d02873b9352199116a685bd110d899350b3a04182bfe3dfe4d3e74363800d25cd51b1
zf2ef225d3cd677b025cb68d88293e9ef1ec2512042b8a2866396b1033ff4bf5adda717efe8be27
z65e0efd18e14c4edf2f35e28ec0d9ddc2100f94b94585d325da540c1a2956d8422fd1d4e3508f2
za2bbd7edcafbf255451be46853d10a067b09541003054a2664aee71e0aca410b9277d29877bfcb
zd8b349ab1b1ee0286b9567ade2e44a1d9391b40f2c4c46392bd387ce7cc55c5c4ba223ac5edad9
z48e3d3b2cc177e7e455b7c1fb74ce33181510b6ccbd9738eef1af3b4b351acdb0f8c09fdefdbb2
zb97a6468ce980896b1fcaa2a64038fd13ea35c5f281b71a77f18a9762de55bd6e1ee8bee88dae1
z5e7453f53700bd4cccf495f2f500fdc835b805956b9fc5e6a2329cb14cfe0fcc163e28853145a3
zdb4d8a43eabbeb78e3c8cc4c1845aae439e4193442bcfe21ca38c69a791d6b265c3ab3993545d0
z56098be4a1bc562692977827a1a081d073d516bf0a564d8c2f2d820382e87278368f79eddacb81
z7abf22af289568388fedd8dd20c5d03e7a6493ef17fcb387d11a2e8cab4056e4c4aa21e8ab221f
ze8fb708b7aa6876da192d98c14eec032b82a2a6a8960fba86323c39bd73072b6f1345e9b76c486
zbf3f42ee0578bde1d1df10e59e1c552019c3200c28d155dc16392bd98b95e3bca26a75137f1970
zaa742e109e4ba98fecea0d52c4ce4aba237ba9df597c563866b27d0998dab29f2b40862eeaf9bc
z5216bc6787a74bf940984cf5894526df4fc365cd89da03a0ba3277667b962c5977a8f1a68abe02
z2251283954fe74212ae02a577181fb0b2e09f82baad349cb47daf3356811a472a6e4ee6068b2f0
z6aba1c5b79a16ade4caae32807a4c1309e7c86acd686a5cba8a047305d69b6b46bfaf6d0df635d
z79fa916f06c46db016050a46bb42e6764f51ba29f874edca9e7389f7d9607b926c35a371d81e7b
z5e
`end_protected_0in
`else
`ifdef MODEL_TECH
`include "qvl_sas_link_monitor.mti.svp"
`endif // MODEL_TECH
`endif // encrypted_0in
