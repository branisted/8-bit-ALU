library verilog;
use verilog.vl_types.all;
entity mti_cstdlib is
end mti_cstdlib;
