`ifdef encrypted_0in
`protected_0in
ze74c34e226135848fe16db9ffd31815111b6d7fb642c521a3f628cf6da949865580b22efd062a7
ze90adae0e65e66a2c36a587d0a790699161455169ed55a01f2084f11770a774ec4c588039b380f
z6de9c5084882a40b79a175f5c2114b2b6d78b070cb806e1c0aa9258297f4687ab308bc470f0040
zb0b1de382961eeeaf2e279e1462520fc31c119af8f2b214846f56c2b3cd2eadbe4099496abff18
z15cec83ec4a77b868344aa20ba7360908f5c0de2a79abf8b3534b883bb12180f68b5d4beb444cf
z3fba8f13afb0abfe8fcc4294810f75afe452434d2d0f1166236c82f76edf1e12979f04bc35693e
z32ae028996dd85737a8f5adc1ebb94f39c940246e887647b64782cd7ab429b0544c173176cede7
z01dfb26b1f73408344a52b7e1f117f12bb9c8077b34876c2e6fdc085981637012dc9754765e1a9
zc512ce062e0b8fb16a214591f5c81e1353b900a611fe1f4886b57940b41b7f2ce99a7b84b04b90
z916f717e73bd10589c81e207ed77ec660a8cbed5b487fa50acde1b055c8870bd8676023f21ddcf
z9c98cc47cfa2d654ff1365d1f45035a045a66c5dfa8279050262529d2cac9e64fd27d9c7de62a7
z731bc808811ded9016570962244887f98fe5440167bd0088f2f049df882af501358497c3b28776
zcdc5426c7f52a851c35106bb93e16fff984784050fc808fad15da3306022d17da80d857bd32a53
z2ebc5737d466752dcf94171cd2cf105efa9c502d8d409200a8150244f03fba3a90bc8d5cf172ea
zadcf57f1aaf8cacc562c30d11230bfd4b456201e0488a1919517c8f4390b2a7a4b4b904dea5234
zc5fabe55b24358240562a4a4c3748d32e0a62d645c1870af4a6e67e97350e8d4f09093855f19a8
z33a08e8fe6224c5ab4e33bcadee89448a3b6ff131307138ca3ca0a1c684c94a515d8acfe73706e
z9e50e1c95177c559f1a230700684027080d0cbceab8f7e5774be4cfa9209a04c5149a3de08339d
zd877880272e338d825f7d1020883386a16a61280af8ebd71e95c264c4e9beb7271845437415e05
zaee6067053d6d032f27276e328ec0c2ba07a8e9d807902b7e5fc0d3cdd9cb1bc5ad5932fb4cc1a
zf9acc393d90817d240a02ed66e2169408d7ca775fa71be58564c336be30fd523f7b0f015bab450
z12572a17a67583247b55f471c6ef6261077f22c34e24d61c1fa10095322b4d96dea2b5db808292
z7e759c09e1241ba78f5dcaffc0b3e9d1b59f0af01fd46b995c126ec9530cca2f63499d27500baa
z08f5bbd03bd308286faea8b6eff8ab00936b6ad363a8775ba2eb390e210f9edcfd53c18dbc7f9c
ze762b3e1bd67cae815e35a7d56e1323b162db5ca08d39774ad54676e6915701445456f2cc32500
zd59fffa2daf23e69c8bcec740cc53d8f1d43b4c758fa2c074ebcc2ffdb8d4123632cb719a7f1f4
z73e5aa34b72bf183ad8acf67faecbc78ca5ca87967032c27fcc9ae2c21c1db0f4dbcd5600ae3f7
z7cbe7763f06d14834a84a8bc7fbd797fbdc45156a234a33f13d6a306326e8222ec75aa55a8bbda
z08417da7c167da82ca7d13cbc2c3f5ac726edca8ce59c15fdb76a374b8e5abb7b227780284749d
ze9648021f4675e2f6933c54cd63206579ca453d21eb5f6b510d1463cc62fb3e5aa36119ace57d7
z357e7e022ba5ccc9b0e7b6ff3130b4c91f741f3de52554ebb01f71c4b97e832d5c6d3eb3afdae8
z9726ac898dbcece5f029aee852eb4c90d21580c3d855b90ce7692efb352629582d0572bb1814e2
za822df20933f1e0191bddc3d58afe85f883232b90b04a410c990016cec3e2e850e81214e81d7b7
za4eedbeeb0ae96f96c1172aa7162a7421316a2f3def7097c3293e71514454298ef0d19a75688d6
z13c3701cf484b4144af59ef1f04c782af1af9ac78ab153f0ae3f2855b6d26ddced18d2bac4ad49
z1b196276adada0fb727bb440ae9af0a132e47b613dc32d46bcead719ee05790173bd6c9952fc5a
z02ced3b4379519ff2faa1dfaa7313218c1357e7f67bc0d7ac856bd706dc45ce2a05dbe09dba7a8
zd1a98c79e01b7c975b21ae20b6ea5f7d1fbacf20e8a589b00de6632c5016931068b21628d7830e
z458e1c0bd6629eff104a675bf253efe762b2c1bc020e68fd34f1f8f5c71bf94551802e960b0f46
z72f27a623f978e198e2d84957a738aec01b1ac3bd859caf5fb46314903870d730beb2dd57597d9
z0029d733dd43aa32fb00c14259a62a3b7f7432e941091e0cec8bdb5234cd9069ff9f0dcd3be260
z1fcfd7ac052de9ddee448d9b06aa6f8d2b678e8e0902887ea4d87cd09e17fca14ad78c5bdb1fe3
z93bfdb1a39706cbf3301329f97fdf586ffa5f1c3b24397e1a381b1afd963d5b2f7dc216e29e323
z063e1502062a5503ed9f47034dbeb3db38540a4bc10c325c759cd2164fe65bc07dc6b678a2ec0f
za3bf1476bdfae0682ff819c77cd1f4a62b1bb555d0c50cc35fe5e2112c3650d3e8ed59291e8d03
zb3cc12603ed876fc360356e972057d08a091f1a9cb25324413d5ee020bcc389ac16c5f0d3ca30a
zeb68f965bafe47a797660c0aa3b08a13b40fd2d82338fe7762023e7f5dd6d42574c604fdbfac1c
z78136eb0cbf8061b4c878a71abdf9f02c6a2d1c077c070a56b2132876b587f963c768593540344
za9c912763aa60d3331db585e80c1b0afd4ba607241d839daf2f38ba17db0ceba39269db33967d0
z84780c26a8589487df844daf6f9103d6888ba7689f2e30ce81e369dd08388921f26ddc67dd38ec
zdf20142f9fb34965025d20b460923bee4017c197f3e20ee1ff0d04edc1e0e2f8b992a8cb89d8f4
zdc1683bca36db2e51aaf3b4b4bec3896fb62bbf80ebda5bbbb204b618a5de05e4fcc1c322ab709
z35cd855f9ac1cbe69f7da77304d3a46542d5db8cf159ef6f4e5127580d9f5e7555b17e8589f861
z00666ed048c06a3a6282cddb5e7fd9ae2134e28bdd7ef0b42f06d43b9b995ffc55b21d81c8ac74
zfeb52f983b0e8198081c21a8fc1186f0fbd8a11cedc5a938146508d366d9be0e0cfc76443e11fa
zf1c6cd2d12639786d25434a65bfa2fd0f293b4f020f1f70ad29c35250023e6463571313776b5e8
zd6fe0c40c1a2b60ebcacfd30ffb60d042f76dd7ac78991ef1800f17f98f91823123a0046a23537
zb83e60459b97cc3df0c841f7753b2f5006bbf14f43ab1e4ee65409120db43463081261ce23305f
zc2eeda998587132b855f5a620335bac529e2933b32be9313a3f153770e5953df1283ac374dc910
z6bd7cca577ab9ee2c297970e064b86efb3347e52c1c3b23fa27c8a995fb957d5131d32b85e2095
z3a86b01f527d13d69e2f2ed4decffd903e8f991afe50910e36ced7b85ae4f595b85e850009c4cc
z811727344c95410a55a8cecebc3d24f93564db159af7b52af76e4515fe01f836e06707871086c7
ze2a30b843e1be01425de49fc809e1845fffca14b25254f3f5fbccd46c674e3cd00607ae54e8cfc
ze5b5ef7e81edecdae3424cd0d44f264a3a047856961c822fe6787c19e73c644d29432ce2cd2e1d
z224bab55e84fac4cec79a3dcb74a1ac69504baa1a1b65b17b3d4809746b0a90c6cf84ccb481be2
z87901036bc4830525c7bc3e746798f18fd0f0e066e317ca46e82e48bf91a68b5547b7de8ad66b2
z22629c6bfad0c677a0cbfe3dbdc9dff3994a2f343fe9ec49dac5b6d351084d682c54acdb7844ca
zdc2d8383cf2b05394be1eb321ae43f3383385cf10a8fa10b7343624bc8ca70ec9459d52463232e
zdaeb9658ac502ea8ff0bc8c70529f488b6fd39daef59f2bb2d431e05a9d797e30e4bd0cbd1cb45
z5e7bf0fa923a27c7a2a760b79d2106ef10ef39d2b97db41b329c47483fd883d9c8aa406e37fa70
z172ec45a97c1580e82c31057a3c276bd4b792e3dab48edfb586e4559bcbed2f9c5c8a4ed9d70c1
z1b28a1ab3831e98099c8bdd4c3c1d5241c704bd8eaf9e87f3e3265190f65a9ee1bfa03c0de15a0
z245cea8792c76df1595b91e145b2686d409c7dac5ff2adbf492ae7d34df830e53135d5f687d6c9
zfaddd154c81b8108f25e71c9af0e4e53404109b95f3b8897e807a4ecd63ce6a990f18742ef79fb
zacf87e454dd02b2ff91404b742d08635caedad78ce13c815067fa1908c61cbc9c5b81650c4a047
ze15a299c00d8adad932be545f78414eac3d88320fece3c965f7d53d1e43d2e62379a68a58ae4ee
z6246355d81c30b6d6c96cfa3b5fb672e005936333306421c44c095f46abeaa6f46b5ec0a9edd3e
z0e662684045248ef73b5d42c15a9c02b3a538e7020df3f33ef544f5b76413a2f45909149392952
ze0379c9ef0e99ed8da46dfd6dc90452269776d2594d79d976c1b882ab4bc8e65e5fed8fd54f7f3
z99e3bac9df6c5a8dfdda2300fdf0e390bb23a7b0df57d1438f1c8fb7a53bea2a39e5c857b4eefd
z0762c8ba95638b5e7834d5de48b77415a1c36803f6c3df6e6c78a3973e4e1d482cbbf3be9ccf3d
zf02d8f4c36e83502f2fe9eacaab96c867f106fb89ef7407797508ad47c9af669fd83f182acc9e0
zbf6307924a4f4101c103cc94b1f97aff31c230e792d97b89a8bba05f503218c267e81ca2dddc64
ze1d636cae378dbc76d35d8479de7883d916862290a9bafc31b553fc583ddebb390d28cb52bea67
zbb1765ed1a7af8123fbaa0bb5e4b858359d715ddefed5f35535317b0e41aaf2ace9af3aaee6cce
zfb01f2c5296d9b5d7cb8edfb1bdc6f2cb17f38890724befdbcea92182a5891b443ccfdf3e64d19
z1d69f8af142fb370644232cfea634fbe7e1b1694323def01804c7c13d938368de4b869098a6f78
z4743502f5386af2197a172abd28af2d00e037165da0835498b5d0478a66612b616b64d57d3bc1b
zd6a4178f63ac16598adb67ee36bb5e14e2b188e9ad67bd5b5a58452c9f520839e0c800ac284462
zec4ad379cbd878268feea512f1a0fa74b70d53cd4773c3d57a8e4bba9907c468c87608bc4ef94f
zc8f917447e9ac542376744ed41f0d6a1481c03656f7664441c60073dfc5acba884bc0abacac20d
zcf31441e954dedd1494da7bd628dee7d394ccd6ff75f805a9916a3aa6cef231d4269cdf18535f8
z67f52b6bcd89e6d55e406340ef07c667fbdffabd84a0e9a55528aab06b0f9f1daedd1ee343e8ba
z86c0d48459c90ce1d079faa89c2d2fb4fd24e61a368f08607eb2119c3ef5d6a87d393d86b4c49f
z16d30292280892cf3922951248344e9149d70b54539fae52e0398494d00a1c582ed1eca24d761a
z20a0dc39212db669be771d99fcdd6c26e12e0d8441f2616b925812d625bab36fa0d97fd2ff61af
z916abe08787ae0af450c813e2f9d5c3693127c41355a0e91646416ffc1f447e8ae5c2cbe6e94a0
z15f9c3d46d8b99845f049dbbe89bbb98d5f45b0631296232a8e32ed2952c026a07e1c94731aa25
ze03bfd2bd0be599bc9d375ef493a8b5a638d63c3e16aca269a7ea3b21c6397d1905627d19107b5
z92156e36848a04c6cc453f5d2aa5c9e34f79c7d22e713dcc921c257c67545d9a1625868fd45ebe
zcce1d0cd9ee011470b88fdfa2d2d3c0c399a13d765d4551c1504932241b4b2ddf65ae580de9455
za9dc02c02023be92945a674f010e4c72ad2073c61f5d764a9b3e36dcb2301a7b92b2f3fa66744e
z0a22b9e382f9e71cc5919f2853a249e2092dd7abe302699604dd8ef857b221a8b60a09beca35b2
z58acb7fb3bbe82d34fbb76e3df9c20a605dd3d45193066f398e02c0817bbb4f0de1b307fc6415b
z5a6ef59eec30303aee6e129394e584ffd55b93e7bc848b90dc63ed0b76f58887d3a51f4222aaea
z063ad8696fe8f4bdafefee95d6a3a85927950efe7ab0eab12708d6ce6ed6aa3bf10b54a43e6e00
z997b6a3918e9471781bdfe02670c3924bcfd35993b888f34548fb4d59704908bd4ed3be9e96364
z20e2f9a9b8c42e6ca129b4d59849728cb09ada524aee21d9ede991f5960bfe107b28f7f2239c44
z863629056e1d4dfe73a8a361dd084f0bf0d125517595c5c9d4602b6e043347dc18ad944525e62e
z610750725917c08142340fc4a130bbede22baa1388fdad4794196a5a4f5a7233ebef707365a54b
zab76441caf2276c269e1ce8be94301a9eb7d9862be02c47967a3a07f4ceb956f5b0907b4f4815f
z73de7db22efbdff76f52b78b26a0b6aaf19832eafd2e7951c71b45f2b0dfbfb3fc4ff1d1955739
z6e41ac1d689d3c04123dfa3d8b3d75994dd95afe3d356717a56f0b22528efaa679ca6492344450
z534cec19f6e9983b38d2300c580b44caf402585b03a8277847b579f1e2037d14670b1438787614
z21f86ee6b691cf108a0b4ef108646138a5629bf33e568c3ce1c93213e73395a70b7db1e7f3fd5e
z665c4fc972a3a04dfa8ff5589450f5a79f1d5a092c87a58c5471b729746f9f89a471cc1d1c4b9b
z827d0548f1dea401756d02335419e26edbe5779e1544b07d9c0c4f175329bcea93bee28c28df97
z8c87f0ebc5c25d1a899b913709ee6e465b435bcdfd1456442cbd3080c50c680e6cf99989cae116
z73d9ff10f37316cf2fb6f335915345a04ad5e0db443f8c303d33e21becec41ba74996377615899
za046f86fd34d15328d6ee1005684a76691058b6780b6f6466333c640a18b5212cc8e9f9acded65
z6d22c0c3897b9a7c7b93e3852930a033cdb74c40865fd6ff6fd74646b200c7307f8782f2d26a7f
zb89be47c12ad85b7c7cff5130e6a1a62624ad4da8f0e0fabc4bc0a38b5aa5d0fba3f39142c5fce
z0340960c44fc9b7a12c93a98a03e4ec02874aeed1d482a32b94cb259ab90a4c4ec87ebe2bfc60b
z42daaeb4867c874a3993c52f762befc0fbe1c087479330d5f900fcfed85dc3ef20b623cadab85e
z46c0edf0498f5d7400a77cbe4c91d0db9ee3b45915502ebcfbced67f4eeeb1ee27c8baac7528ea
z050034c3b7177365e0119fa6c74952dfe73b9c873e7cdfafedade0cbb9e0b15030722205a4d763
z8f4b7ec8c21426fe363e0a6a8f67e67e5d8a4b6ce963dfc539b9cac7baab073d92be07015c1a39
z29ad020e7af3625069bca6a3cfe9c8d2d6ec5fcfdaecf9106f33149572a653cceb83b695944ca6
z41188b8ab6e1ef672d8b06ff527a700c306219d97b0269fe9ab288573bfa0b980ff0d727ba87fa
z1ed73497e8187c1e8a5f05d11765a3f70f2bcac73bbc3e8c35242a9d6c54e9f82539fbc5089ce2
z3475e34f0396808b54906ee17106c57ca72badd41a7e642e500d6e1ce80a13cb9649f8c42bccb2
z28c60a90ec23f0a53c267756125c8e4bd3e3b73f4c8a7036eaf436dd53c866af697c6661d5b91a
z3edfd3e3b8dd12b9d56f999f8015bb9cd8abcc1edd61aca2d8a0de2f43801301cef3cfa32dc133
z71bbe8d75eeec4910276c5e37f925143ebfccf9bf56e71669a80cf01027b9c095c0b1fc16cddb5
z8bec7b5b2a56a80a7908981d382d35ac53b65f7f731393f4d27f4d2c2f430e670dc8f90dad8b95
zf9a476a704e84c7db8ab7dc24d941e68f4947a89856dfa7f9dd5e617f6084f86e381f126a3c9eb
zb484b801c83bda914277fa90b4e3f006178bd7a2d1ff6529fefe6f304221ff8f21e10319e562e3
zb3cfd2cbeb3814858cb3ca9408236e873f52b4f24b5ec035da9029ec233cd2183480e0b6c558e7
z0a7721052026ae3f2150e0880a5a89ea3c6f04edfe038d47522a18d39770f083abf2e16fb28538
zdae3c593808a044d7ed33ce18cde197e54c57e2d8ba9923a38a0d42416b18051777b19b04dde5d
z97550371ad79b3d7a3df5e104bc4abaea266b4324e5574006c8170153ed1cdee9ceebcb0150f50
zb13781277666770fb365d9d6a40fbe73148bd059e740a3743962cf70ba5c26c4cd861f9dd80f88
zab0f478babb2bac8424dfcacd661c6661c95be4de530ddb1c9e9e011684806ff95f60f3c1340a8
z587d2cdc3394d96787f2649bc09d3f475e1de28257f8dd14153637aa641734df80ee2f1e03b059
zb6f956909635d71a94e273b7412c222640ef82c7bc05ae618ca2906ac57f5dd6c4c7ffc64c88d3
zb00a727e856e32e814862335f1fc83275ce2c939d5ea34efb9ac0d42e37a72fd73b4aea42414d0
zb4cb869510b70cc033760c054479a7d2bdf420b1556333d0285990f7b7c52758ab68313223319e
z72caea6dad52b4c213d23352d556c944dcfa64298da6d377f39d1e749f6c5698b9721a49a5227e
zfded658264e1487c4c154b58ed4e492dbafc9cafc321b8198d0dd878654f5ccbcc36cbcbacf557
zb58ef0fd1b904e060a6b2290e3827f637cc0435876636918d5209f10eb3c0b72d4389c7c7ee662
z648560b9b67e57f396caf61beebec473582b719dcdf67ee9b0da4bccc966304101f05a7ce687ff
zb68dbab24f1ea19a39c849d0500f6023c5f05af06ce6c00517456268a8ec5412113106a657ad9c
z3349c8e85a65e9932efb2645f613bec646a79c91164cdc053535fccecc6a957999f8c7da799ed1
z1a86e8c02af205455610c9b7b834c9ae56fc741dff1d90e20e7d098a379ddc3646d482c364417c
zdd8656bc24972fb842550062399f4a9cfa04ebbd1247dbcabbe93a5bebe1f9edb23597b366738e
z4497bc0147bb4bc19dae1bde7ac5f744e5188ef449b83f7fc5ae2d31168c51b35d14d669884092
z643f2bd2eff7afce62bd14cbc41beee7b29eedff9d580b430e13837c3e4173c44613cc2616c30c
ze1d6e721f803986e0d3a3a5a65a9a609e8ae6d5acc2be1bb3c90f649c407e6fa56d745330c3304
ze7010f99b0053ed6f4ecfc9633efadb796f4b60d234d170695e34bd49c8befa25f678a8d552e32
zdf7b5141e287f50ec06bf47988d099f8fd71608a5665236ab063de320b7e61cd444ac3e3bc108b
z5cb2e966f6c788997c966676a04fc2f3e71367da3c950bcc4c3197aef8e9fd90da9f14dd606b76
z61bb05f7b58ed2e8ded1fe903278be439301df57e0280efd2fb0ab325a33dea61394fea63180fe
z2361766eed5012676754103012f061ab2353a0dd47df529c94bdd7a019d1f7426bb809b8074ffc
z032d8211b52a3aa94dfd32e262460d3a4b1ffda89438ef3415047e5ff07c0a66a2795ecae5981a
z1dee7fd202f8523772d3a4af8e0b6ba8b39b118205dc8d250a984f8ab1af6e83efb3c6fbf0b0a6
zbd56b1e946bd9021185e45654dd07e06d6ca580c2a52d0f28ad3fb8bdd1f4153d62c37155c6705
zedac6b0727645abdd91919bd80cc90e3c92f88eb266a0c8973f6d132cdf2848222a36b45195a0c
z2c842df5d387ff10d52a225c012fd9500f03002861697309bca55612617747fa06d380aa924e03
z519d6660531614b259e2d0b3dfce76299665a22eaebd04d5f44b5f93969afbd226efe45319174c
zb951c90e1e83136262afaa2289ae24713c66add6674348ee18f195c2dea8228c68ca2517a3b28f
z29ff0aa3d6390305d280b32e2e43ef8f26c16828b7df6f5d9eaba6674b748fdc61b17fbd566719
zb16839d05b6ee8ef98da94127f8c2dd01b54f862d48a1ce597ed4ac6d3cade638996c6a570950e
ze2823f324c648513263fc0f91bfbba06986f24e7bacd0b0c0ea9abbc5f9c3ab9532a8868eff184
z96457bc8e9e5eb6701a78459a8d8fd293ce705929ee4a77f7b46d0cbd071264785c33a3239c5e7
zd81fdd81d3ed52ea4fda80b41b6761fba1261653b1f34a56da5c0c7ed485aef6f7f9bfe649e7c1
zc2c361c00c412d4e67c8fb00fce46dc0530ec97c1ca69d6762436c4c318a69b161d8f65eb00e4a
zaea8c6c4b5796c1e34e6d0cb6065a080bdd76475ffe4a7ab0cee72a800e61c643caef25886bed5
zd407d2ba0cb026a601719cb79193eef796fcb5f85f9ecd75b0db7149ff894f4c73c9f2445cbd7c
z46a86f22ea869f6111a335c22fedd9cb34eaf77ee24cf049b19ea590babc80aa3dd75459207c64
z0a81a20ad40081bcab43f76ff6a5b8b1acc9495e7d9a9a421cc8e1698030cc2918fd757675fd63
z85667f9b3edc454150884233e80f8c1e1c91021ae0b512356f94a14961e9259b0c93756c27f9c7
zfd1d0148e17ced9d887f943c5ec11fafa5ee888a896f1554c26a2d4490e1698b2e4d720b20b587
zc8956c375c23e8fb9ff384f5b16b0f33822a03ce3b12058accab23f5587969e1746d4fe3995fb2
z14e44514d9e4fbdb2d9b0e3a13b68fff971bfa861243e0e444e99d645c352880533632561e04c7
z528a8adfdfccf6a794976a041bb02df03a8bfb83bc636ae0fd6d979bb0b1b0c2d396ee44e23b36
ze55215fceac62918a0f190793b882c4e02c7944617948cc200f56617f8ef6335d98a579f95ff95
zae29baa5e7c7e0900ede2647fd7f5b8b905650ab914fb61f0134edcc6c1a263e0bcbe392935c40
z9f787f467db8a3dc3de6317741ff8ea7f5d78115317532119fe2fb30847bace7c5f9878cf3a2ae
ze40b950098ea7453f3d17588e82710b26353bd78d5153ba1152151c2755a3ef856c635a656825e
z08c95cd568745ffc4322ed9866cbb3ed19f44a9075c95d9db39379603cd7ab4126e6af8680febd
z173f24274a146abaf767c9fe7fd4d8667859f0653ca17d58e38128f609aa20d864509f70285a74
z40f41598eaa74bf5aa14ec291ab108d4b88645ffff6610cf5f9d052eea29bedb7b659d40e81098
z6ce8793996511b61dc9f43fdf5fc0d7d8c9534c87ddc1de56154270ef6522a2c4d153ca4e5711b
z5e8c070050d71ba85164c7143c3642b78b3d8bee437deff50de35be98c24087438d664ffec1802
z05c0556f7022b38f205c1cd115931f9ad8d88f2ee65863938840c8016317997457b1683e25762a
z064fa56edb1e4af59a4442aa7009bace039b8cfda96bf5fefb5eb17b58d07cb390d4da9252003b
z077261de42af0d111566d33e5e84f30601985fc5fd2b40e5968350f4b9b9c6eff2c4613ba5c874
z25817dbab3ef07585c3e9e9b00f591a1da6e52f15ca07db362104a636fe1f7f117e18eee6b706d
z7f8784e0db900a2889863c1d7f683940357b2e44adbca069ca3e2981f325ed623baa2289453c89
z9e7e135ce2137d9c6e136c5990001521701f22a88c1a0476904847bcdcdad9ac14e2544d9604dc
z4c8e7e5bd34bc9f506976c2fdb479139bd51b7da2f8089ba2c6165c896996e3bfe598e17163e7b
z4d8912373e8b0c1b0bf44b1a1d2996de1b0a89c32391443004c64f5b8d10adefd43aaef73e8dbf
z93ff1d79f43cb0fa9b44007a71e3d3037f62f0e7614cd3fea8038904507d1bd57d561c8d6bf1f3
z4cd4cacf5f2524da6e8e39da6c77199f949126dd2d36efb62cf99a0c40b216ff32c1cf47fd5530
z13d6dbe9c98cfc545205a80bf4daa07919bdb333969e0623b013165077cf72fede0c6dd0126114
zd562cf637b7ea1178a528922cac4d7f72e551255125f30f65b26c3a87f853b45529aa93804ec6a
za60949498bb962c96e08332890b7bb46583961d0e0237ad83bb9a042a46a3acb26efad73a1e37c
ze5a4905cd9b9ad9ab8537aa79174d211bb2085fbf1c8478846a4624378bbd8dd23d23b469604a6
z6613366334787b16fd5807fd7d535b09234c3eb0baa2ec8654100f2e7ffe4f0ce13bb94b47c16b
z2e10ef8881f9bc8d63786510d15350469285430f49b38afb83be5a8ca350311ecbe517098369db
z94e9d66d6b432db95eb142de7a665e3cddc5445387eaa592e69dde3ac45627ddeba5bd605271bf
z125f3a8fce8ba34d29bedf99c090b6117a6d7715fd0970d102e27de0be0a93043262afdd9aeaf3
zf7323650d7216df7a9296a4187ad1abb6518a0e8807ac0ba93f0a54c720652d2776b59a28507a6
z580818233b80b8ae6d0cf0f42c208eb24b31bec1e360a75c9c15fbbb30a521d1e841bd64451317
z614a8b6c55448bb7dc79cee6d91bdfd159ea5186e3b1f51cbbb5606e56ff396c3adc05d8194533
z931949c39aac1776a883b24dca9b706352186c71bd376330a796019cf87bf45a8304663492d236
z6bdd7d19e47d3243fdb1b772abcc574da8cf239e0ad55edaf117a931a1eabf45b2303810402c78
ze0bb94ae93ec15b303982de8e3a44092d82aef949e55691d84c36c8109f8b80f5347cec0ba44e8
z28429b55a8af06f6b505b270e535bb67382ef1970a37ffe9a8e725c8ab63cc46797683c839d735
z04ffb1b8f7b25b1a8f7aad83089ca452fee868122d20dd491a34596e6b317a02b38ea4aba84ac9
z03b1fecfe9219840738461c013aedd9938585aff38800ec5e94de0e222e471a163d74c534cd8f3
zed21f5ca64b78ece0e1879cf97cd46ae807044f3236ea4c5374cbd9debd9b5ced19c74419c7172
zb01e848a106d037e34fbda66f3f197f8c6cd54c23775f7c13e74c5f76a1b2d739bcee2f8b9fe98
z7001c9c9f736f89874f291e8b46aaeaf7516489dc7a12b6ee0172e90da82c9238afae91ca0816b
z78dd4b93a4cbd55593395dbeeed2a9d5eaf22d2c24ec8b8f15250237b816d019099c36bb470135
z894a9fd84b0e21f5d7e94857d2e1d573f5a150b7a0b8ef8a176cf0040aab736cebe920bf82f391
z936302c8888b7e8a06ad45aaea27a69b33d041155b385108c333fb4dc9701950a36bbc91e43a86
zb824812ddb5d9657bfa50300b7e7e333ec49005247d82a9683893ce76607bb1ba7b523b0e03476
ze9cf27cf7454324959772966f82ef2c3d03689265a9c8982f5f69051721b6cbba5815fb949fb4f
zccecafb6d56e97b7f7f17bab062ddec64396610e3f21dffbe83c7d3eb3ecfb4848fe55559bad6a
z18d73c3491acba5fc2042d8c793292dff777d4e58be3ea1b280fa193eba72285730c323ce17bf7
zf1572057b992db09531e5bc23fe3a44b2ca0688f9ec08b0365f56c1ce0a24520beecb6d4f4fec1
z3f6901bbfba2f07e2faaa081127d2ae456d361cd3357eb89abf5df9854448b37c841544af20d30
zf6917bd5f27de24a62ca1deb9b806c76aa22a3604992f745167ee8d70597461096762608ca3b28
zdf0b35bab5e936eefcedbc01e49488c0e994f20dc0daff24a40650820a1e5ccb3dae3bcc3fc18f
z0b8e6063afcc60a1d27c8a39a522ea1124bd90d3960d1a1be91296281fe4d69f9241a6feb180bb
z538e3988efbb32dcfafe32feadd0d4b3967cf6146dd2f3b279844c7d4c8609965623b84e677347
zbf38c02c55f4d8fcbe70272b8b0e4eca24a2400c9062d0bfafc2be19a70013f0aacf553a3af760
z2f5c01892359a7b05d69a9684b52af667bffd7d31d1d171e8159876ca87e458a154f52a1472f5f
z0d49687fd128b5d1c3f6aac549312a08b1ff1621223a4df7d85580db02d3b7d89d121f1170d80f
zf04c4a2f71d8234a272fd48ab6f0d4a03cb752beaf72d2b452a351979637c7483587d5c1faed37
zea97e9012fddba0c93cdada09c37ff2ace3a7539d6c4a3bf998fb6dbde7739253d8e859487fb25
zd5344e0c0c7256cc376b8e62bc5a5c3096480948c44f94fe0e4583fc35e463100523ec7e36a7a1
z43c0b3c92034709caff9a549122c4caed50659a317b44de84ffa0ec5eeadebe04b51a820cfec92
zdb2aae0fc0e50f5b35be612aef421c9b1af45013b950280d5c24e7ccf82775478a5a02dfce72c9
z810246bb139a8e6589e2dec036c1e5a8cbb5b8a8f5db4ba96c670edf0c00ffd59f9549cd7c6916
z1f66a0ced1e18854fa742659c5f0b9dac65ed7b1cdd35ff24a900a742f07c9b9bc5ee3bec96a93
zbe15da067e05c723af0231c9e555855ec41d1a47fc94adfe453e29e4f306536a125b8f6540e724
z020184c9709b0dac8ea03ffa47510a787d267a4dc8732ab5a07a2a925f63692967af87a2077ff9
zb3e92d86449d2f4bf3f345f37d9c0193af5423065e31849528585e48a5d288dfe32c58b1f32e97
z1e6796b6cc65437e25dcb72003364ce87ab7af48928c6fc69925fcca37a51a5375e14603b82ba8
z329344fd4735133a7897fa4d03fd56f0757230a5113606e9c33e2bfa2621a3db1af8b8a6172a98
z5a4e48292a97587d6d3e61ce0eac74bf65f778b93dd0a70b1df161abf975b23783e216bb6f23d8
zad977b43cd78dba56c13a81924636b00b0a9b63041665d2f2b9b61e07c53050b0f59c93a907130
zea1600773ec8cda04cff1cd7ed4899cf8807d3a15ffa50b35a26e68b8b8f961f933a5007e208be
z5ea43277726d2e54dd397e3488ba4c1df3dbe3269a1e1e39fcf6c828a80725e22bce08e4fff4cc
zf356335ca306b7e0da84c5122d61e2332a9c2086bc7cfc4f36ddc7febd76debef87e2d7a3c5588
z79a5fef98cdaf895ce8d0f6afaa34dc878ab92c394d569a32075627d5815b6b827ed027a0b8d21
zb579c13dfe5a46a25a9001bd4b7173da3a2a0dc33d31fa24c18c529b70e1f4a44426bd5af5039b
z01c915f3cea4b62c970823003feb730bd890f9d0850aabbf0bc46c2eb98f0b119358970d3b2202
zc736b966d9715d79fe40596f838174d845ef76696449c1369b0f9cdad59aae7cda254c0dc80c33
z2764a236a683c3ec9744088240b35656cf80474fe96e385068ccb6fc339ef43a9abf2549df67ba
zc4fde353164b6efa5419ebaa704e2431dc5fac0524173135f3f4dd0af25397c390b861e8a5d521
zd521fa34f552c1a7de3f903586aa6245fdcc893215edc7bee26bbf6d426ba6c69f81f79582180d
z656c6fd2c7d6dca01a03219f6fde30a3e4dde3d236eb834ef5fcddceddf78dfdc8a7cda978a681
zac8d8d7873216c2682830b1c2fb9bcf37b4d45caf09dc3e87515fee92ce67ba5a5e3213ff515ce
z65516e60394dd369c3078f93eeb535ada45e87335c307863c45dd059c16d36a6fdf7d5cd25a47c
ze7d8d100097288b278ddad95a31ab8c60f550fbd2232b54f98a62f877bcde2b82edc4f7e82278f
z4b7adec2c89cd04510cb1759827589194f73d2ee75390f13f7aae2e51c5d99743bc34b2b5b9325
z97f8c7e28993d09d0dbbc11184df12f5fe9bc11ceac10d958dfa77ff0a5b2ae8994c9da42627ad
zddd64600e835419ceb0c43b0452f9970dd379c8e2177b9125d6e9cfe2bbec9fd0296c457504218
z229056f28415e97a85b26e3e56dfa29e0f8817c0edac2fc18d0be7a1fbb767d61842fdf9f97d22
z827cd5aef24c9d5cc2e6af92fd09aec950b7ee4ddf6a33886f2484050f5f14751304cbb1276650
zc17dd55fbeea66d01ed43c926182626d77c1dcf3e701018f97bf0638f1671020341767127bd3d4
z6a1fa509117ba8673be537f617a6aa61d0014d5a355e0483af7b5d672fc84b18a491b17f0124d4
z88e463959d1e03e002d8e664cb32798c701b30c77a607773bc1df87daf132bee0938347b5c28a4
zcefaf118bb340c667ce0c9ec79d371091f3f2630c4074442b7d06cc1d493fa554b31281f70c6ba
z331a5c48f663af2261c4a8cbb5987f487cdda8f144ba92b73b3cc76192ca0d999a4e2353f4b972
z9109976a52b8241ce8e062a0f44a4d67685aa61fa3d27d76e3e4bef541ae8d323d4cf94b9d24fb
z73b892e637caaf1fd5fc3d6ddbc850c991696cbdab908d062e990d4c902e92bd971572f002c1ed
z2c4d8ad0576fa292ce4206f6783de70e73ecf26842775997aedd603d1ec1cc29fa392b593aedcf
z9f705c68d31b97591637c6ac9152530c0be064786044fdd65c8e41b0bc487d2605c3cfc21af6b9
zc5cf5864ce37caaa96000c49e355cdd3c65ef81a5419908b44a5ec6398ecc751e6777c58af0514
z90b763370c6690b37c77ae6512f74675040da5e615b3aa80598fbd7f4f77c8d1eb53e84a6e858a
z3947b9147625974d33db9120666027ad6a1b746f2bfaef5d4edf5622631086702683df5a0311d4
zc47c1ae9681b495bef4c49a4f11ab69b9ba11d6dec5be70e01e8f84393e0573d5ce363960a27d8
zbd8c9e5460936affe5bd5418ab64c7b0344b5880954ad35535364118a3f78aa37156cfebce2291
z2bd95875b5d8c309eafa5f2949f40e3304b94f7db51dff40f43e2bdf463ce6f384a483f1c5676b
z77bf5f07cd981dc42b26c7228e80c9aeb68454ed980f28f87cd3be94d245cbed23f0f6a25fa54a
z89e790900bd867f6824403886dd76793ba13ae96234d5baeda1d5145408a3395928b158127e085
z866fcfdd7a64863dc394882732a142615592e804640512b77d632955c3d3e48f92c9168f4ca368
zf220c40178b9466c0a0d9bc96e99d5cd170197015ead11178360b68120ab865fa5d5d6c8634232
z3bb3f9cc5049590b4d3f60077d2676f2b4bb779bddb1599cfb9159ca126ee77aaeff729b9edd45
z0ac3bba2874191f90974c2bc4978f6bbbe2a5aeaded21d536ecb78eb4e0caa01fa6372bae297b0
z2b15c77638130e72e9dc29fb902207489cbf79cb0dd9c43549831abd8585d11abe3aafb5eb32eb
z5d84e2a0a8cd28740d91ebf695fbd54dcba508355815841489a836b1d52341894d22f12d949e5a
za9ec1731d2d36da36bf64b6e9353e981d2f1b4d50b44de5924f7de5fdcc48909908d061ea522c4
z48746444933ba75abba470b5c21d166094e0afb3013ce58f5b3f4d7aaffc515cf14d693cad31c2
zc6dac4324a1896872379e83dc7904377948851e9ee858a2564466d3debba471d67497ebeb9b165
z9a79114036c80c27a23f41bb782a0fa96cd2d17f125f6c059d85cd2851b19b6fa963f377bfcf97
z55e72ba671cd210be0320d5df5f9b274fc038165282a248722e8b7b23c3701290d8c1007e8d06c
z5fa337ba639260e5b99e95c1131de15647a2c497048796dc97ac5541d9f64836cc22403543082a
z30a0c4e27b9c6286e761953b156f4d49c0d1719170f1c3298b605e9de58d3187cbb9b74f139a80
z2d6e8b30e5310d43cdf2def06efe617f114164b8a1624336c1bf0d707b7766b0d2c11dea29a56a
zf2f856337d39218ab2368a06a8a5b35a5b996e2dda6a9bc4d35a7692751020d74e831f4f4cb369
z7f2aa77af224c6739cf9b5a8024ec64981f42bb168705863881d5f377c3dadedb95d7ae183947a
zfca20709eee8d3ac540957286f68eb85c7a2519b2c4e0c6ab375a82e18ef32658816b06b176bcc
z22c6a3acc6ec7ef6f7f65f88bb297a1c758b3cef21cb35ab67ee25ac174fe25399d1fecac96607
zf9f36e4aeaa57cdb23d6730b8816b6726e08e81ed3cb47c205180e479740c5746a69460f045126
z9cefa1c67a8448f3b1062af9a6337ee03a7fec565699e91c50c21e28d229cd3263a1fce2593598
z8e22fb2c9b27f8ee5ba1bdc943bf268dce0466027db691ad40c74476dcac9d015640d60f949eb3
z6369febb3c15986a4ebce9156c82320b83493625d4e7c9f0e06070faa30bb72666e334ba198f81
z692e41341783e568e267efab1194c71f5c8b5e8ebf302062bb69c32974ab4837d60d0f74269b47
z1a740f8704dc8138a450a83b84a46dee5198e55a45eb6b0c92e1a538889b07ff6e435b1d0fe75f
z7813892363e7e931de7f34a494623624330751ffd74310bacc4224a79b9495b8d6c270142466ef
z29502a40b0985797ccdb879081547c08d3c690988ba4d009885f5b58711f7f0899d2796795d096
z1cfca1e2e403a93c079f5d0a4d4dd86b7fc52f3a5dd5e28395f3f7bd84b4b97b3e7813fe66560d
z1f5adddb54d91eb9ce8190a53e924b8705e3eb443073446e8ed3663fdb2318aea290f864938be5
z9aae1c1a0c560f260a3bd1696a253ec261c7fa0508a4d44f9f9bf7859122b2cd08527820819d15
ze78a0702c3a0fd08e774c91686eb05285e4fd403af3b483fc7c967f5a9aa8963a7f8a982c1d974
zb410b557225da83dc05981797d942ebcdcc3d441257dc8ba668837514b15ef6e8661c3698a6d61
zbc2ce7dde430984fef458c3d6059d4ad4e3d990143097f2928f22c719f491a88a62db735e5dde9
zf7dab5cd8786a741770c0e1a5e733890c00aaeac34b54616ed4e1e66ba2a669fc8c8c4140b0e3d
za716e481de3dc7a88ddcab8ffd91e9b5da68a216df25355ade092194bb3259d4fe71d43c4f0c37
z1459ad4fdec5a6257e71578c226def42e2d86163a48f9e12ab7eabd58947ded94735784ce211b7
zfee356335011648ca504fbb4d1541e1fcdf9b9f538e76f9e39989f0372f047d6e708807786c341
z4837f7fd5efe4711c234a42235d6366026e8ebbcb46f0c977a774bc875d6ef42f7a4cd69caad34
z4d98cf605b522bfa059b1e815cf70442885507951cccea1edd3b4ac1fef3b61278e8c9279c476d
zef90bd8bf383fa78447f8cf615aa81159e0d308fc15659c697eaf7f57491aa646f0fbac3810c78
z6d459c118130710042b79218cc1893d66461c4c3c9d89f371d29d31673c5eff4daa3b06da4545f
ze18bcf90fe3ffdbe7f815162df55e6cc86ad995cf0d20e620ada0d0d91991ca754d7f0ba2b4f76
z4756b8ebb373de89df6bf2d511d8fb0ec99755746afb9f77dbee550a12e64074820297badd5a62
zefd1236149fb842d4245d4b9870107c5ed393a9c44e0696dd2c9e43311b49953698713820b617c
z2f312e2f56d31916efff24a6b3ca061940745b9e3b13ef7a7c9f8a312588bf65df32ca8e807150
z6d97ac868658b5e55ca33b635d3fc687bcca88639d11071b3ea6a71545afde49414e4e076bcdc8
z9d6ea4b30e60d476bcb48f94c5e921b5d24c6999d545c3a44509bdc8bc7202b5c579f2072e8056
z0c6e17d09fadddf86807cbd7aa4790f372383e5c9c3e52da5992ec51240993cb3fd1b792ea22e8
z5f311ba03b4a869d64367d04fc8352b8eab5bc6e3c90622e477b93012cd79c65df70cd21e17492
z363507b5e49f33b5d301fd95ff9292a37e1e921f77ad016bd8979f0907f726e2dd67b40442dcc6
z27022553bb2b8ff045aa29c776521ba2672c964d009eab8770d1161968a1dbcad0c54f5972dd24
z05908752e1e14b25c6df6b66e6f9704c1ae40a361b061a847d5a7e9a6dec8aa17a69182e5777be
z14e0c8fcfc470cca50bd2758ebce1138cfd2e8339ae6200873d8fdac1a518d85dddbd554cbf21c
z1113723aae788eef57a3ecbc1cbd37ae9cf750ff8b99dcebe20fbaca0148bd522f380a6cfc4b22
z1f9ca64446216f9294af0a8ca2caf873dcd1d8dc5bebcc261ca7647637e880812bba665e338bae
zd3fa069f8504db3c3faf122725b525dfdf0f6fd80babbf175e4c4c29b9dede69e3d098630d704d
z40e593c61eeaa4ed7182e6f0025175d05dd79142fe9ed3085bbaa23a38d3ed2b135ab3546ffc32
ze06577cdc5ef4534980309fc7adba7d946a85e1fe24234e12201a41af9d1345d4f5631cd89dd6c
z77a3bf208b080250fdef4b063d8c30d1dec0ef05f9b755f0086eb6eefa50d9ef239fbbabc6a8c7
zc7fdf2d3956673f96ba7be02f50292dab19ef861e40aa95b04577dcce69d74582c56b2cfdd84f0
z4f50aaa2a017deb96a9dd70733c045ca4cafb1c24cce8ba3df99fa00a9dc4ac171a290695984ce
z7189cac401521673c514c1ff3afa320447e3028eaad6cdfd646b510927f4cfbe5f9c7c758ae894
z8db334c6c6d7e8673c53990caa742e894a0948bf341c7242fcbaac4dc14aafc21d4b903b65e2ba
z0a2fa9615108b7a4ee45ea8fb947286959119f2cd5b0d4ec0da2514344f0e3e6f0deebed4667b6
zf9dc6d09539e58f58258c6441c7e5d75181137227db78355d8d58a23b9c8514827f21fadc4cf74
zceab8b345484f21478fe3b59682ff68fe64331903fbc9d4703c2b427928575df38effefef2b177
zc53daaa935db5a46b0069ac2e77bd4be0448cb54217ed5bfcd59e396a6048d6d706826070636cf
z5a245b910e181f038bbc18ca96f10b414afa6d78662f3d7bb168d536e018761b7f6a8dced0d747
zbc7625c9a7e55f7f9180f6426c40ede8bdf170ffc802c9cc9795083df7acd04d3afeb52992103b
z47e890a87b88fd38a49a5bdae113214323396754352a961eefe9b53a70014ea6064617bfd7199a
zd0772430291d15ffa85e47ea924c308d1262b557431b708337ddf3454306094eb6820ec481ef25
zabb6c97d104f4f134d3b9187df1fe70f0c95a32687e961361232de3f4012e74f805c154ff214ab
z97ebfb82466fb104c42cc45514f9c03455825adce7687bffcc0b3b5702e859ba6376ad51bc52b5
z6d384d8195f9ee742872db2c4ae94ecc556a8d44d5413980e202f748eefcf4765df75441af1994
z8b311c6ae4f486f39dc16d879fbd4792a1f8ffe8635bd4ae8cd714c17f5313de2d298f54ca7938
zcf9bb8dc6ce8138073f30dad13582ec8aa11d0927219e0ae1250a49e72810959a9249480838403
z5c59c247a8f2bdb4f7d4ae9cbcd4feeb819ed314711bdd8695d45dfcfbd157a18db0d237c60cd9
zbeb0001bcfca924a6f7cb313e79c3ee27b86d5673b162c2bc405b816215b23aab09c8fc9e32011
z79509dd49046da23b6953e15892350a7249d5bc8d2e6e0dd487ca535f2fbd972cfceb2dab60d7f
zf722e3a8d47ef3b50b2e7334fe503f099e0c137c4ded601c45be2db1f71ef82ecb8f572af7d271
zd7d20fd7027d911b4f946dd1266bf36d8357372046fb548a38e9618a4cfcc83b33b0cd0395e78c
z1a9402aeb886c08fa40fde2d5e87715639f78ac6eae9ab2719247c3aa419f20daae6f2d3372f85
z3a1c191da70a741a85c86395fe3a5c91fcb236294cd40844e1c8597117cae67d71f70d22ff2d45
z237608fe71dc30bc6011bfe9a03737f65bcd0725736dcc11d49add8a7dadf0a8295b436ef0386e
z2c5ae3c97c9b1fbc525ba58c6e15fab30378e4af81afeb682b8af2321858a6aa078e57877e7539
ze690357bb26d6e26da0e8ff09dba6fac977468ae98d237c27bee0cd75d023da770e3156d5ee663
z335260e216d769f66761f3b919be8017e492bf6c4295008459c31c530dc5911b11b5fc4a420657
z3d8813fb98352a0d84b88d1312f47bab750d208ab4dd62ca81690391dbcea76ae64ad90c1917d2
zf1b0f193cd5c47d8ab1ebf8d30547eb6425f4b0ef0f202b944b9495f36bdbe55646c9f00847877
z4fd7ab85760918a0c3b5f84f6354360dfe9433b63d8372f10f5e373ba75cb59a9a042d094a486c
zeb77cd286966d6eb14c7104f2fdafdea536d41c320ac42f3c042e375e53239b31d11c46bd1edd5
zb7ff4a942cc2111ce56b6ad59984cb390d2a96a2435c5fa1087b108c469de4834f901314055a51
z29389ed3fcdd94b58e36c56b79938fcf7599581970ee2588e942e6800c7a0dc179500261a0b5b5
z56d598e63a6087003bacf0d71ee766b93e07341fb2e5dcf96e654c4285316def645ba579b60039
z17dbb3a6ce288deb78f1897348fc78a7f06bef86d30f12ba9bb375fb69daea27f8afd0ca9ef34b
z35244c05c0a81c2b5827605be61c335abdc51440cc9a281ae1636500f1feaa974b47fad0878dd3
z7ae5e936ddc0df925bbee2c2d226804c6df831ed3ace8c8d5ce29effde2fe4804ea2412c0b6c11
zd33ee5e81c022b174eb188bbb366a27f489cce0b22c6b3abbffde2328b2fdd0a3a427c4feff0d7
z92426913bac006ea71f3d17a9bd5a32ad4c7d8930b5c7f3fa439046557aac7618afe96f3f79768
z64019ad5811a8e160c589ca00a9df15c59deebb507c06ac53f4d4384bc58afccb0574366d64268
z25fae31713ebeaab30731cfc87e43ca13ba54fb53be0f3b06e901be9a43e9400a07df928f2f71b
z41172c949acf302e6f1c843d5bde18032238e79914069e694f15127cbd9c16f1fce6647c502e88
zc7aa1e55fb2161f2a4a22cd72c31050de4279978b513befc5f0a4647805168f88648d342d46ac5
z88af1292d18a40bb9e3bf2b4a7601767a27ff0e3f9f1fe1830f067440cadfc04c154540f60a838
zff94afbb1abbb9f1abe66dcba70d716f9ef5d72631f9c4a52c27d24898e1a0e8f01735730a7168
zd73bcfbec31668405f684a59e4b90d5eae160f01fc28b2414fba3e016b0e3ead48c7e2dcbc9041
zd32794d76d9b0eef872cdf346c3f5b9314462721766bacfd6b625a2d547b8ffe0dae70d1856d37
z725ec76d9e22ed06213998f2ff7aa632790055ac1a5d5a5a88d7a680d97305a699150faf654ad8
za6843944fe21ecbba38a9fe3a5ea017da86ee6b1b6889c47eaa010886cbe1e18c75486024469ed
zf0330ca55bcb10113fb70f530d1ad678ddfa5600fcb541fee7e457ff277c02a4bc274d859cbcaf
za19d58be5e02bd7076e3963a661d96b1f48f6ea798cab8cf9eae20749ff0b64e08b43c48acfaee
z446e4fa11c3344ff6d80af738b574a9f2897e4b8179715c48b2cc5cb3518d63bac1845efb52e26
zaf906c34ef019f821e09237ca88e7f710080d1e12eb028571891756acc1fa2e64736f1daba5f6c
z6483dda7c3eb2446439960baf01ed9cbda6473a34f0e312b14b3a2a1eae2c21d02d684ad7720a4
z3c30e69b15e116aeac9b13e831da0180dde8dc0253f1b7ae3bd7f6988f9d0f4aea9ae79e269fbc
z481d75482eeaec00b2f6c57830084f5ef6372e9c90d36b941b84b4a500fe022bc97f39f562faae
zfc802e78aa1cb3fd070dc8cdb3d77da656954849263060b68bcf2ae428a0bc8079adfe211f62b2
z36f16fd8e294ea73d43ad29caabdcd50346d8c58953de6d4f9ed60510e9a979625c4a957aa8453
z5c84080d767deffa5f8350bb9e934e8319068fb6c1d63724436953c49d90297cf3f30d6cc28574
zdfb6b16f3442f497b36f179fdfd9edf866d8a81feddea4ae471c3e4b2186e6b0ed51b80802807d
zc0f1bfb0bbcf04acc8c988799218f3d5ea69ed513cf50b615c9c8daacaa607cf90cb27ce7bd5e9
za7c4617a4f92c1c63a1652dc33ea848d6a35c63d29ea022eb9517d2b5880c7d317a292c2474c80
z367fbc0fc93343e66cf76ca624880883d70002e4ec839f832b1a963af0d5484a756ec72392999f
z630075f8dd789769cb3dd5232a03a549a15c68da39728947aabdba0d2972737705d66090f6f31b
z76267c94d1d495ceaf80783676f99ddd9f5e28081a0a8122082435da84594cd92188094d718a76
z9d71e1fd5b0465dffe3504e56e20f2e26fda8194d39107abd4aaa9eb740565e415db1a3fcd6f56
zd5d60a4faa808ab533030f22a61a0140539bf73c2e7821459f867776a7f02cb7ee26942fe39463
z8a8cad08dac3cb35a9d3f0fd7f34a26cb47d1e83bc01fa909befa82af6fe62f71f5e32ee4de4ae
z654697cc8fcbb13008a70709cd5c09bc7bffd666fdb63545d7d8a6648a1b25e984feb141c82c54
zfbe1232c215cbe2e77025674fcc5f4f08f9208adda7a07b0066885d0d5df40133bbfa99ae84988
z40b7e95c2ea99799d1c081b013a208bdb50f3fc803b182ff61cce0c8c855fb9d4f9f203e3151b8
z805e2f0f2d7a0c6a244f0ab1375f49c8b7a04a32e42e2f18994b1ca2e60c88d6caabd794fa6881
z626aee7205dcd4c547b1ed5293c25fc65fb14c21c7fe5cc1d9a80af8e4d94de5ad9f517e93e014
z5a21cad6e52935031456205ddf854cd250a4ac774423a8680d18dceb1e03ac998882725db64e1d
z4ed7da53e4f52eb67e04904fffd6202e7e658e3f807ad2377a165554ec689192d19b3ee474b284
zb07270bd7b6ca4af010957b0fefdf2b580363e9fcae5aa6b8fea527984a20a152b202f18b91b96
zdf63649658bd9e743cfd1846f0ab79638eaabcadaa0ac075be2fb9bd32bc61ee73276e80b0cb15
z05d7ca014b404db2213abb04ec6123d4bf5982febe6b6790eb16b518c583a7a9853a71f7bc2b4b
zf6fae14eba5dcde2c553e16fee66c9891451cfbf5a4314aeb2a27a8598e893e7a9a2483ecaa66b
z262b59ccc9a3a82c69dba087508056785c907df6d7ac6e639631f37e2fde1af2f792eb6ce86585
z253a1a5f189defbb96b2298f0a62db300887ccbfbac00f92ad7a65b8548410e046116edf9978bf
z0b83f875e0209d5b13b2e2f0f0f8742f44fbaa7519a04a2dc7878961c245d0e0d969c9ce55175b
z7bc00231ee0780f8f7d491f73d762fc67022bd13a350193d9a81b4587d098d2705a84cfcb270a5
z90f7eebb3dc0099b877e4f1ddf7b15c28dc69de1784c1e09e6757a509c71afb7d9e34db4e1beb0
zcd6fd7023a2d8094b4241dd26728429374dd0ae6cd4528247c92949e5af41ba41e45aa96def7c9
zb3eeb1bc420a3d4a9386ead8415eb00b665d71424e334961f89a12de99d0c717993d6aa0b0a430
z40dabbb6229ef5e1df02fd6b580400090ba3a74667abde40f0ff61f2a92e0e3316e52406a26f23
z42839d596b0ec091b1179ec769763842c4a54fe85511269347f41f64091b7f30bbf32c8e2bc34d
z20b09012ae05907c1ce124bf21593af4f345b563d99844f6af6975a87f91473fa53a2d9be6b093
z5a4da335cf29c52a490284296030426b0861a588cc1930e84776cda5c139c1621732621a79dd87
zcfbcfcadf97083f0aacdb5b2276adfa48032e57ed774367648fe91ce9578cbbb3d8fdc73e39fbc
z9640677bfa06b2c3e054727885306128261ca059dddd5c7ade2ea794a636d93a4d850eb5439830
z1185745c4cf9ce8380d8ea70042dfe2e866941869f4889cb2e80491935169da2c2f6652d7ef86a
z6b365e3319976a385372f2762a98576688d57fd6cacf32468680f6ee8c3c2c8c8d8953770b9dd4
z0c4d594a26d85ebfc9f7291ca3865bce4bd6089629abfe54f373ce70c38c5db7a8daae77146fb6
z93c3dbe6e0ab9edc7b5a5dd2890bd903bf230ccf5ffe757e273bc21173ff232c908a9c2bf99130
zc119cda2f273c1a4b4d6a91248cab1915e694b9f9bf002fce2c3726bb37168be7aca7c90b76180
z777cdc33316473db243efee2c928aa23a97080b9c41fee7532fcdf19c5504773156b417adee100
z1b12c039f32a28a1ebcd0ba1f9f09a6b74d2a6978bef516d78f170887486691458efd9be950382
z929eddb4cc601f3f9083c4daf61f51cfd930f5c7217ce735eee3daea90e8c114cf43d0d3dec973
zb4632dd755cdbee9dfdc0befa7898f9c085a65cb23d4357afea7f2ffb46cd3564d207ab20ca6b1
z2be223455bf90430c7fcb898680190123521cc36737d150a0a5d12f045e3e28fa56350f1db2cba
ze0a3466e3dc012a24e03a6171a876720e21992b170ad33952a5056066ddeb3bafde3f849c9294b
zf6991f1e2ecb077c1c697154c23cfb73dd24c897b1f230433caaaa1ec2883421a8b634488dbdf7
z85b154ed66478647b00a666158f355fa8ac4bd19609ead8caca5b012610302de2091bfce7473f1
zee9d80f75409b7a5e513b84b587759eb2f3914ace8bd1611997345ef32d6911fe3235fb377c4fc
z5cd5a51b474b0cbd0085722b394d1447e69b211a17bd2bd25b0185d2482eb018ab9a26d9328ae2
z5f6bc9b7af45aeee87ea5824c9ba138a12707c3f9c526a228e9430855908a5ec1decda31935f5a
z5904b5eda7be0ca7dd875b524bf4ed8f92eed5c6ea79f5a405ce6aec6c11f09fe4da61289d864f
zeafab7dd591e2a7b2d092d4d72ab940e0c371bb31eef9eec1f687707b3440e58dc722abdece4c5
z7e3debb394e604006dfb9fc2a355229a88352a461c5fa82c54aa5c57078c5e316581a95fbd28ae
z637d77c923c87935f8f459f12690bcf80bfe68b80a2916b7631a1755269cc99c45a5fa34ed9044
z7d95f1219ad6c72836b1cdfe9c091e5446533c9e2551d65704e4fb631883a9a61375404e129a2b
z6a8c9fbffbc93a5d5f38dbb7dbc2041d1f7368e11722941af97b8ef49b8cb3f7e09304fb5614da
zf9f14039fa08f1b40ed66e823c9e5e8c1f194169f2ba21c59af678eff860e98dd1a70af24e7a0b
z034aa516d7536f62078e476aa7bebc5cf76d7054f2b5e3ccab558aff6d36db94a912f7df3fccd1
zdc897aa51b7a1d22e860c64b2ec3e4e9831bf7fb775d4b0f58f8211bd19ef40d29fc2292f799df
zebd7f6c5ac68ceb3ada9db5295b2e7f7b57d8f59e803d9cb6970df0385b25a48479fc00cd11230
z06fd7e9338ed1e9a8685b5e7f8d1191ad7345ecc8cb6322254cd0de3880957da1259c95c3b135d
zd5f0b985ef78c3233c886e3b0e63b12a441ee102ea20c4c4685e5070a0d260ceaad31e585e7b8d
zbed3cbfbe9959afefabdc2dd1dd0d1a6865504a5457322f563f19d747913d50dfbc7320ce2e46b
zeb03b3671c728e6f45a0aeff4e4324661186c6fd67a5a82ef8692f24746b4f9e36e6a532447fab
z1bb8b1a91945ca3c2fd5f6b97e50bbf1159fb1840b1aec4764e8f7dc8947810ca50f4def1352b1
z4c9206f16fbd2f0d76738ab8e2452abca63b0f5d64314457f8e5e1cf67ea057aef05e076c12f7f
z4c412b43215ecb5a69cff4e3ffcf1f98325e7b47a8e1c58a49cff1fd4635018909125a77d4252e
z81d2e4ff0e4a07f4898251a42254ead0c3c5106cef678b2e7077e55d3f9dcb4724eef0feeeecf7
ze0f30ba419d27cd94b322d21daa5ce01cdb10f86728ecb92254c5cfc5e29a4df6d49c6be67638e
z2eb1580440356b0e9829d8b75c42dbe322b92aac6be88b5854db6e340aa6749ed70082486cb855
z4573d9588371dc8a60fff33a55645d5b42c8e4ffc33ce3d6b834fb0f8c998a6bc911e459f47bf2
z1a64431fe6446b93bc1ea6b80a962d96f25c2a3c4bd76b05cea5bd6f08c6f3b8fc0223dac12f01
z92039ae9297ef59d62e6c3c61920a2e3d540d45518deb24c4a40a9659d45d739c75bddbd92261f
z46b96ae1f986776a96eb4629e2fdbfcaa6539b797f3f3d6439b93e42f42f97bd1674aabce8e8c2
zda3cb679107c23c98773214d144632463fb67e57f5bf2acc5308977985e4d8e1f9e72189efbcdb
z6308e39baa86fccde5d65fd91d19eedb684ffce5893a449ce03e96411e6249285d0900a1b717f9
zaa0b45fc36a9dad74a71ea0c8adfbd94b47c8198c2976eab967119c3b587d69a9a5384b2847d79
z4e52da3ed77eebf2d968ab88c3abf6f67d8b05066897286752fb2376c11e703744a4b9120d689a
z48365c2ada7af2f8d1ac24cdf4fa14a6c3bce738fc7722b153857f59751d9534af2f7dd59c2ce7
z85ff7bd0b32fa908708a1a5e1efc7bdd2a87426412440e953742a1a7f64d170d33de097d9c809b
zcf1e9a248efa2867ffcecdc447524320eeea63f70288c7acb54da6c79ee4e4f29e318f4cf84d06
zcafa95116634176ee6ab31966ed74f9ed9a9ab7b2a7f4233432903393761b5b86eb18df47d3d2e
zed1aca41e4e928bb2db6f7aa5e839980e38be2d30e699601325cf5258522231c3b1b0494085f18
z367c668d122b92eb0c6cd35ebaa83e36724d47996002506e29bb057e4183134d9b69d22eab8db3
zc8c27babb57f261345fe05196379a3e9d4f6d0d811acea6183e8051cf208b11701735883e08c8a
zb3d7916a9b9d2d543357fa7e46d4671b17711875ebae7b923cf6f265bf057579b3270ce0e36c10
z0978d886e7345b407a1e7c9066048507f717024aad5c4df0d82f32806261341cd7b6d7137167fd
z7912073ef0bb17d5512aa3ad08778ab50332e122596a571eedf47c41a1e9b37e6a067f2ea429d5
zbe14ec742b8009a723509b7ad40855017e5b54c9ab4635b812ffc7d8259c249ed0c71ace5db0bd
z3ab437996a83f64a0b780a2317df1f91361c855431bd3eea91d470400d09a47b9ab12d056264a0
ze4d87d39801dfabb4cb169b587e5b8f0f330a68eb9d74c475ee8288d5391d27dfe38588856bf13
zfd5e5953248650b343ed53ebd3319355850f6aa2da463dd5cc98fb6924c76ef7e22905d107cc5f
z76b0d3b364b0f207a6445d262e23c71fe88ce4c34e45704853f5e3dce529b5704004c1fe312b21
z2276b0eeabed5f0d01920923d567b0960a1cd9e24ac6281b7b9f56e322e7f729a877547d44db99
z2adfaae7b238158541617753ddbab901284735484656cfdaa3aa8e1918629840f0f6e671f9ba31
zcd32d446b26b02c7a71085813690d4648de77e4ac167af93462b84727ab358d3cec3e39ec7b8fe
z0fcd07ae7b435c959815268a58cc6c13235f5b764b6d8bbba5f08a807ed9bbac16d142fa8f887d
za2b00183b1c0b008b121862809cb3a9609759b1cd63775513e9eff0cab86624ef2c77625b1ae78
z201b7f8d21413d7df097ca25281faec8fbbaa4effe9c18b7d7a4537affe0be00ac29902bdb437d
zfe66f93784bcff186af2350c47f936b04e5d38c02fe15ba21201e8241c7ff9184be7b2792530de
z512c306ea751232fc2743b93f8a2c4b167f5e4fef09fe3ba0d33c3267a5f205ad90577f3317ee4
zb4687b915336f9e733eb3ffb8ca44db1939001c35025828977984023d55a7c2126e4f234f63dde
zc223529a7e6f7176bbd8cfb60211ca4faa9cc444021974069b8503b1ab7c5ed25df2398664eaac
z0f540e16543b1c875e4b684f57dad40a930e3ed7ae552ed118a2efee1b25adfd93bdb532c933f2
zcb05558f3e6a81c6c0af6be33808075fab8a9d07a35c587d626fa2c27cba2e165a701709466ea5
z560fe7960dabb639652914eac25c6e3cc3a7c3ff091ef00c2f3d3fca85247c57acc4a60976fe13
z696d76fca5af5fb31e08644477a36d5545a5e292ece42e593ba27cf414278dfc1076fede707788
z586f7bd448909256029b287726b62ed91162153abab2ae0b485979ee1dbd84a78e18adb7f2bb00
z6dcc9cfd517099d073721aaa3c697cffc801591bc54a5d4949e801ac03c968237aa546b63be4ad
zb80371f6960eb54108c65d5280a595006ac006ef4809df1ea0b7a3b0496da01a21bd5e090ad977
zea7d1a55f99b6349b9f6a0ac46a94a8f5dc4a9ffd12672c3c1ad2d3bf63b41975aae3be5b9b2f1
z7c38c15b7356b70d16187a7172ec97edeea33cb4e40ecc1803b5dd2f48461590f863670fd930b1
z04ce78069390e83368d07df2dc6fb028122a39714461df678a5bf6f5ecbb43c8fa056b1565d1fa
za253b5f7abdd991de6467d49c8b0f19bff72c76b791cfdbc6789ad13197d3aff35087d4c021ead
z59aedad7d74405a3a1a61432a5bcd289e9feddf878a753569d3406d1838b4031e747433540389a
z4dfb310e6e2ae353237e8cfa7541038a423d0ea8d6b7af6bf7307f3efb1f4c4d110de262f479f5
ze247d32cb5b204831e5dfe5aa217a09a0e1979c15548de23c17f52a5748b32a68ab07c0d3b20f4
zeabddd60ab5257e15c1511b5b95fcb379d2b324fbd5fd8ca9d96f24343616bfffca390988c41c0
zc39cbad3c4d5b30ec403f072af4a31966b18eac314df84c2ce3c82d43732076de9386774d04807
z7251e7ca72b88bcd5012635bf76ad2f7572625cb35bd07a27a842873ae57ba03da00f2c64971ea
z96f97f8af5881d7f44d84f084175b6d854e03e716c9b89c41ae956779b5a322ccda95dd6503e04
z1285c5ade7370dcc2424cebe97fdca3d0932ca5b5d70c0b3512546b34492405a45d3ac8c079100
z4ac2e0c8b49b21de696993359fb43517e8cceb8431608ad9c0be98d44fd45ea63a9715b8d897c9
z248d5d987598af372d58728f0079453f8dac61f2b49df434705e7bb69dcb369a53bc90b9207796
zf88a884ffe58ef85469dc67600452618717fedb1cd07526b2f25a682106fa0caebd27dfbc2da89
z10908f28c36324b88fa8b2c6431d0b1897187e2dce9997d0a1aba508f0ca3d5c20d83fbc907f2d
z94dbb38e1f777eca2ec8e56984475521943cd20202eceeed18065750858fafb8ee25715b09ddb7
z338dfefb585134e3232ebb71e50bbe31f716d2159da2fc0f686dc3955ddde36f8efe25f6d18d50
z26f6d24c3b3e4840366c9fe09c6d5f17557a6702f3454317247b52f1eaf864811c8e9a3cb44512
zc11b2484432434fa1cc2a0c112eedf06e66e1ad15a62f392694be1b801d8da222a2f6235847471
z1a33f2fd72330eca1e92e1e6986a76eb71bfa948cc195afb95840196b263669fb2bbafdd80a20b
zdad26b69fefd5b715aee68fb6bef78a7699053ff242e612551e6d04417ee3baf075195ff1d525c
z16fd06d202a28fc88aeedd8eccfaaceaf9a81408eed1234309f5f7c818bae0ec79f1b51aca1852
z83da3a15310dc1267a189a4e7edb5898a748b842660ebf3e09997fc7fa4a2fc7f0543e28236aa9
zb62c81a7d52dbb9e36fd02479819889fbee97f144938bd0a002bf076150e47faec6937427fa0ce
ze745057cc466c15cf214d464624c2bae5fe857429c52384585d174449f984475c5e808610c230b
z267fb3c880aa5331edf1fc767d09784aec225dc27e9bceb615a520b38d35d0c5684f03851af9e1
z1bab7645a1f79a47308939bfffe0ded6bf04d6624dec0a5c15881b1f2c26dea870bd09dbf154bc
ze2c73bb4109e8f0a7ead4f96fd99a7865a99e5e962dcfba60a2551f0577b357a1134cb7deb00fb
z171e7a8f56175104c267c97a2e0ac87646a72f627b6a4e9ae0d7c2006ff17b1de202dd4583704b
z4d83c7e4881336e34bed15ffc088bd88c94ce3af595f7d473ec8084884ca9247bb7d1149ac315b
z64881c8b2227cf9080beeb9dc2c5f6bae8283b40c3e5ccb402d13422d0e298291c3fe946446259
z7c3af3f1d0829ea0252b58a8db20b50a350fdf257d2cd4cf8b60622fbb908b68ca8ae17fa83745
z019a9d9892fc492b3a836f16fa367e23bcb79668e4f5347b41f2c47a49af8df1abd03d3449a991
z52683911354c1382625ff4a89ed11ae83d8b4ef615c8723781241caaac8e0146676659eb0e9f76
za0dd5ed4a0ca95d4d887dcb1b9a87409d4af0013c8b9c146dd9a22b0f913e5261e8d4d15c40b19
z45ad66930543acccd1be1db3987b8221caf12a5d3426cd38520a97a88af9ed7a25ae1938645f48
z1182cd6adcae666d77cf30fbf0a94040b15b3ed8781e904e1c2589896784d3ac90450345f8387a
za4792a1b86eee10d167cf52ac282011896c37a8a0f3c95aca51f35dc1b80147bd888930cb01180
z478998dfd2f85c3a5fd31e7498525ff2457727eb0c0e1808c5c3e3dca49459e8ef960c00fbb91c
z4a28957e7c358dc4c25346c0ff8b21db5f83c65612433a5088ccd9bc18d72843aaa87cc1e75cce
z899c9a6041c17ea72c01d0b993eaabdd397f45c0feb7d40f161c88d53970d5c4144c7f4b6b8f65
zd97345c822bf7eacfe46dfcd4ae9beca26326c4743abe6eab6a4772f66bcb0f04fc6dfa2a26f45
ze5bb917523400a63aa01c20fea1903757c93d0ec3329432b92762f2019b0f1ef41bfcfc4e8b618
z4225f47acdc7d451d53c2bba11416bd21d48a8b35e4f54d8d6fd2f6db86529478a3b940109e275
ze511674c1ec66a37b6e23304a4e109b12e6aeafca3281c9c85416dff53079bc348062917680af8
z6175dd9377bcdbe4b351e5472cb12ce53f35ba235513a7496c5341cb9b93d459bd4e95098b7472
z98d44a7233178cc67f190b90430602a31a0dacce92e5628726493c7f71ccfc751e43dbd87c6458
zecd31918e75919e4f59bcd1de06218194415526af59a62267d0234a3982c5fcbb3f4f6edf501b5
z94059e2d40415c306f9950a4737dedd609b7fc0cf4be07f5a547ca31dda3a14de3f733266faeff
zc572e95bdf31cd8df632ac693b149515deca69abf291e02869e272a4aa565b7f42d68a124d4caf
z1a5ce9671198429bf5b68c5326a91fbdb700578dd7d317d7ab99720c1424e1c16c63a71fd2e456
za6360fe8e1c584113894b170ddfe137bb8f51fef63b56aacc62fdc208dc274faf10573b5fffa5d
z43f53a89376909593123ef09550a58ea0553640f1548c94b937fac852b6541c9018fb0d17c300f
z1282a568c2eab73b524f9598fea5f0648ee86174930ce1214879cc2d5ab79763ceb6e08a72df60
zb16caccb8452a8ab4fa6bfdc4cf81f64ca75fd64e1e3f68dcbb31df45cbfe82f0fa18f7473f375
zf6d926d3ac832e15fb474052a657b91a383fbbf36439c3f5ca4050a8ec175da7aa962d005f52b0
z2a284c38fde5442bb05624a4dfc12ff95b3184b42afff506bf7e3c1aa0cc67604364cda7fc503c
zb33c370f17842145c0575b261c0f0754daa8c9ca7b8e913bfccf897beaba8715336ab78af31d17
zdbef629b26a47e9b7ac16f69183b356b8c7115be5f0875cff583443d930872f250bb1d4767befb
z9156cb690f1a5b53a476df892791ae3a5e1efd4a1e23e7fb1be41a8c6252fe390d69b2406227be
z8cf304545bc0a58a92c26336119adce86ebf8fe232e0a71b2e17f677e58e971f15b4cc5293dab4
za731d3cf1ebb1ad1f40d560f8b76c3e5010bf01ca633a412932ac05a7b0821725b4f90685da3eb
z1587ce96edbc00fa8bc107869f07b0e3d668b2446ad6af086cd630723055a4541e478aa4ad901e
z4cf6d36ee2f2b14561e91fb2c4e4a30972f7d743bc63b518880746adf2b39fdebe70f923739729
z496a1c7f514f71b32678fce657d3e367faa4dee35a644f61b34a8fc8bd967221265bc1e410f090
zea68d6a643945008706d8e59dafd391e0f43f58fded97eecfadbbc39e37e214b5ae23412aea3a0
z04e823f1798a2d002e844598e92ab18719838aee04d9efdbc6b4d1a1890833e1c6503f3c72552d
z30af8ef92b8706b7e045a7ff01631aff719ce63d52d5ef2c365a59d20d5802cd30dd629f482481
zea5a6090f53c20f3965826510fd8a0bbed538d9999090db71dbd9d5f66107ce9ced0f669131a7a
z2ea2138eebda0163c82072d78f08c0ee661043fb19fead5ea93a57b31bf54587eda830abe43b8f
zb4ea81e965eb1918e63fc5379c11fdb9dc37132789b2ddc812f9921fd18309ad5b7991865f673a
zd3bf7c215b1a356af14e45b1ec41fe342226148d7a3bb86041d637198e03b2ac3c3ed8de5d2177
z1470ea362661b335a8983129decf564b2060602c60304b8da3d3eb57413a6c78db76129b1186e8
z05acfea6ed6274089a3727daf700c57db4da7ef2a67ad9020efb36cc89a3275336dce6c41342d6
zdf7d3689a0652bced89707d4e559f8cf9f510d2be4872e03a39b7738860bbf4a30383e91f35fc4
z522084bc11a22aab74b739dc6fbb7a2823169312ed750ecfc6854f15df76d765efe2954dbe859a
z5ad09e844a284d66120e3097a969de5ea0d818730e575edd853b035629d86aa39227447d195db9
zb5915ff9db2dec63a62cbf43b5c0417c4e207449c2da345517c95bc403a447c463e47baf2121a4
zc038aedb3e862f175ac2afc59438ab2710144b945c6da9ce32f8c92393353074892ef494562a2c
z24bda1059ecc2763be0efcab259b857bcfced955e81e8c6e9d410933853cbfe1a30b6cbb7dda3d
zc6f00aff5610d7422dd148ec176e53da6bca2759878a546128cbd0462cc5a02e68826de5b24438
z2cb95f94ba114365956c54791ab1772cb633dbe1672396d291c2b0e187e94ee3eddb49f4ef8b2a
zc5364c826ef56765b49201fd88c1ff43fdc75394f56e04519060256f260caa57dba8c1e4ebcb4c
za84a3a66f0f489628bd5bb3aa89131a00f1d48078901e591735e54f935524c19f4bb3ca2c20f2e
zde58ad1d79f5fe62233068d9b1f8254c6fc8cc22a3d10c8f95906cb23747a6378193f056a644b5
zdcf392f703538f22d6f3b1a9957c5a44f7d2022b846e16650776f1c70e1557851d3203d066cc9a
z9fc7c950922a5902c7f1024d7cc916080672a1f29f95e52f679160cb18360612c7d23a9adcf8dd
z7287aa30e566b20d7ddf7472b7f1905f6cf570e1b8dfbf3c3de1b4d5f11eddd1df0471f27a982d
za8bb992b1146e8998cbc505e4ee3c2ef0c9cf691ec6d15ed99906612aacdec5a0b269bdee35c8e
z2168b8ef205ccb3bc7cf223211ccafd31404be6872fa4f063650cf77f929b1ca4cdc555d1acd57
z929e56a536b0c7f33ea608d675b1081abfc6e9ca25c0cc518dbd08966578e88cbc23815672ea66
zccc38c1d9f2b7c660eaa60c6f823c23e9b55cc13ae68355d848affd71954d1407c80aad0e8318d
zfdcc02b5ad2d4f3d11964ca7419c1066ec38b9a2b79af51b9d3caecf98b58372c07d388abe4195
z8d460202fd22a19f415dc1f9263c904c4c07113d29fdbf4c66a234f6743f8b9045de7f42e6decf
zfb80661095e7bc63307bf3a06c4bc3f7099ee74579a8b9326063b6cfdba1e7860bef62ba467b96
ze0efff13ff282752540bce816459a221a7e4531be42239d98761ac51852203f8a597bcad442098
ze21daa8a766464e0b38a2525cf12e7e36ccce60d03658927e5886a5d9ef2068a02d0f1652a55ee
z7933bd4598fa548a8fdb551ecd708a12081c2fcc5125a37173fa66ea98cfafd38ac7dcf8dfd50b
zcf82c96d3b394e1f3f7e58d6f4563016cf9f15009834a725e652592850673f223c96c8ff369c57
z54a640e2d0651c563105f3d6d1854b989c10addab7d7bba1c8fd3e6b7e86c01621142c0415e972
za7dc65096a88611e66564b564e61f530c3167647947c9bb77c08e622b18df6f87d98ca24077892
zb97056aded256d6333c20adc38f877b208b4dfb8beeec032eb45ef41365e7da1585bdeb0a3680c
z4994448511df0f9451550a0d6f1004083c70599f2903a928130ba5dc542e87dd88d80668b5f033
z37d2883f96b944eeebbb38f08d3cd356f5f3432f44f1e7845ee0a173f124a222e228bdfaf4dd69
z7a081ae9532c284d782ac9967e753c8418caa286cf2db470e61c2e8b5ffc4f26cd45a9a9793f8b
zc66e48603ee354e456ea18319b9ad326a3c98488e4a99137ce33c845dd28d510f70a7b18f6d3ca
z1687c289808ee2a05f7ca6547760795cd6f2480e2dc828565f508a5603ddf19665cdce1a07e77a
z4d88a16e748956b75b1f3da16a5ee789b2a9b01d3741ebcf1bb94b918f5f05e9d5529a890615f0
z0d24906e0cc439f7c691d6369176cd8086ef940f2f2c65ee7a581043337f44099f653bae8014bf
z3e7b0b5173e4b6a80364f28f83ed0b6d62edc642be15373456e58252f68a04da4d8f9afefc9620
z51c749fcd4be5d33d92ce7b5ddf51433e60b975e91748a8adb9864bcb37089890bc04150a27291
z28eda0d59e7ae745edd8f1105b71273ea6d98581deb87dec38cf7c843a7426c5552ad8241b745f
z2fff30d8d60b840dbedd5fad5f7f67779406d70a441cb2d7ef3bac2ceff3b2ecf44fe488df0903
z7028244be75ea2ebef2183aa245a396e00ea658c355b3d1a9719adb916746fad1903f4a938e4dc
za1a649e6b9a8d04ff2f1cf37df901c4b989dcf6ce381d5d7f8a2700211185a642cbfdcded8c636
z133ba8e7b1e793c656cf218f50f9e40a5eb5aeca4f27a5eaa0d52de2c8e93e92358697f0e5ac2b
zea045b3b6df6c4624536971ac5c826826b3aa4d7a23329adf2258f02b949073816509c69428e71
z841226dfb7b4ab6ef97c6fd8a525cf813d0cb65152f546d587fb6761276dcffac0efd7a61f0054
zd51504da9a3168ac40779e0b2642440c1711e8610902d04e97b90f959303190179665135e20340
z6c4ecf03eb257d134563a89c6e64bb38b12561160e92fe6f01bc836a0aaaa430ac65190745f780
z90450ba5b2ca76f0a2646830d813dc9995227ae6615ece113e2acc0165895620a88da79ebe538c
z16c76db226e34f3d0ce36e96f04a112fb952a78975f1b12188673c7a0682a398dea557f30f167b
z88da516484e449776be59cdbe2c5c863e166441aeba0daf273cac6876df972cb1bf439f67d5e95
z3341fe23483f3c4d82f69f21b994dfa8e5402c0befdefb179e609701a64418b76384a7adc040c1
z2d046eeed073bdd941129aed477d74eb59d70a7d242adb2dcc65f2d6f7d4fafa701cb7bc67f880
zacbdd4a78cbb51ffc09e2493b363babcfdf4f3cdb5c597afcdcbcb32d508570882a6bb93c71f85
z0ff0ed8e2e12ade5ec0d54434ed86b95a1f4101cbf8d7584e48380a6b7b6c6c94f87452cbf5d08
z3d162df3a3f2169de0b160d5944382e2451a73097264e896e52e7879e4841b440f11e955c14cc6
za4e2c915a2b4629ff655e350abe431be6d1f68533770c2eb200b480e5a8f33611b3412cb6e6097
z2249e2d623264f4d16e152b93401535940fda307ff98ab27a69ce20e1faaf0694af256a34c910a
zf4e22d09071d943f101e7cbb822673ab94f847477c975cc197058b8349cfbabcb4ed224e6caea5
zab808e9bdf9c8fdfd8086e72d62e017e4366de2ff74221f49f788391e4e0d1a7dc88c1806bfbf8
z54d6c842a5bbb867d01c85fd363a93f5d6d7435a1927032c54d15292182cf9c7f94ce4fcc0586c
z205b7b1a70bc6387bfe3527db77bdb931807fbaed5668e19ab9262c21f1ebd78fb1c8e40c6c80b
zf54421c93f41186a6cfa73dfdfaf1cfbcf0262ad72b29b722886ede08edcecadffc70ab9e40d6b
z19b2c7f84f0d6dd507ac604dc0606f28341317e4fac3b1c71bdd574018e4071ee3a6620edea1d9
ze9762e626b0cb337fc137ba3819b4758419601459433aca6ac56448c5c368cea59b3c8bd535c86
z3c563833aac745406db479ae3b4b41b07941a2371f9dcc99c6f2dc513352500f47e8cf7e45b459
zf7adafc072d4e4e62b9358438e8b2147d6ce7fea714d9a4624c8a01d0fd5c91707c37cdc0e6edd
z1c4787ee529d73a2e6416c08862d3ef6dbe52022cfaf3da2edb6e0dff2c3a366e8177d00110826
zc1f60c219cca23c109654c0adfcfc0e352533f644c775933eb8f17ed7b0ada702d9964ea92201f
z96ed5bc64ff116026a8e395fbd65948b99f09a647020fea9fee81da2b1aaeac0d363bc800babd5
z8f5cd9f2c30838ad560207bc4eac187465d96bab9a72bcce790d1009fa7eba44d5ba84de19ef26
z6e1aa6625ea343f074cf704c9d0907a29351226e75ae79fd25a73cf204bd052bed4f0119e5c1b2
zd8e2c02e70287b0d77e8e06785dd9e098d5e840a6b5df61f0008955e6838b9e4cff66f9ba0adcf
z579646d426dd40843d5962926d13fda4e40f6860dcf5b1238da4173ce996fa657a5709d6eb0217
z00744936236d498468d55897a0492deb35608d6948300691b0d4bf0f23d7e7a23c4d892935c0f8
z58de29c97a953a99b246c46b7ff326fef2a1d90efcf3bac388935e380f720fba522ea5b4b8c46f
z9e6a92cfe3f802f2291fa08572160095f26178487a412298f2ad473ca509180664276a49f678c6
z31576a077f8d4fe875334834ac5e51182a2e8033a652511690f2709725832108b9af6e98897f9b
zcadb208383a5db7a49a46684321fdf938a1ffa43ef0b0ce8f1554f1908c02b7e1cbc1f7b253406
z7a5002de880a4ba10381e1bdb820ec1cdac54fcae2d410488257f298b8c31e5fb44a680282697a
z11bf8fc406a07c038fb24e868371bd1e5b5f71db822a086cf4bf715841baa892afb0fdff150fd3
z090b4a5395ddb12779b7e838b946115a7cc7bbc2b9e5e59fadf25670de5bdd66fd87214d507b88
zf815bb5354825179f89fb1b15dc6833c67931ae6ca996b464ce696e02d5688ad009551d8ecc808
z0408157cdd9f6a3e4d1b582bfaea512247d8b7c47acaea94200b730b4d268ce19f0e5f5acac9ae
zed3986cf6424bc91c3b2562459df55cc08055e1793dd69fd53d5a33fc3a8a931e97f73eaf44900
zc07c2cebec2d987a19ad176bc7fea5dac8646d22ddaa4ec0daea7f1bf5e602c8cfdf73ddefb370
z1319c2f84a8b9ef4dc068f3d950bfb4f0e4dd97765a1352710b60f3232f452d49eca80a2f7fc8e
zfedf968318a6c6380c2749e4e170bc73edbb0c0b774f8110be1413abda58586e942893ea4f6746
zb0b35b090eb6930a2108ff0f7000a8968c1fafcc01afeb74f77e2f43ce9b9d50d3c9907e79c241
z07f92da25c5f96a49c978f719824f8a60c61ebb3947f89635b8049275c53b676c0e47624b7ee04
z1dd36f7c1628c62a6a4843fef63d7f5b1b4811ae029246ed5afd3e248d9ee4244f1eedf02d6c6d
z68288d94c9e992ffb06f362713f3a531f7d7f17d12a8b1f7a886ad4d4dca7db0670db047df46d6
z8fe14f95d7af97f049af590bbacf6511f1951ad41a6dc1cebc3af71ee01d7aa3eceab3616ac397
z1abdce51f40bb3a6e329a84d0f9c9005ed7618a646c8c0a1bff35f49cf129f2e2d0c5559c92f6c
zbaf8ba8dc9e62c268eb6ca2009d69053cf2bcaab65a2358a43e1df9aa752ce231404a720a9d232
z40b3fb726e352d9aa6afd37448c02cb86719935244748d7c4c1a873fdaee19842a2cf11c841b24
z366e41f07f07cea83cbe2ccfcce94d9e8f7593b6a335776b287b1cdf749bcac69bfc7afeb18282
ze245ccb99b8ea4490ceed421494d57f13222c278b2cb4e631c78074afdb753175faf9785b0a7e9
z870fd2d6dd82890c9dc3c649afd3ba494902d3e6a1889c0b3befeb6131f55fb15972ed17a6b047
z89f107b686ccc59b60a986ab663cbada999abd87f64866160ad3af93c2c4ac253edca52dbc8c66
zaeae6e056b16fbc233d9ba4761a0b99edffb0ced6d8c2b4425075f838066a4c339c00232e13867
z20713bc0fdbe0031859021b2dacf142701cffcc60fde28c701025ee3e01cef3fb59fd8604e2dc1
z9d92d10d1420d701e6912bf0f5725d7095cdb4cc2fd15f007c78eb20d52282779a88690c4cd2d0
zaf058415f6d040c42912f791eb123d8abb792bf78c85dea29ab59307a7a2b7ed81710ba5844608
z97bf1755894de26b31363d0feb8e5ece00a21a66d031cf2219a4b7338ef7771d04a12faa33591c
zaf9b6761ac15fb1a14c6f11d409a5c45552dddeeb8bfffc9238789da03dcae83417ea671489358
z0208a4d735184f56c12e5ba31d746793b0375f10e4db7d34000fe731cb1267ef35c7217c06a0e0
ze48aa345d6197c6ee05812edeccfe28c995bb7e739a2fbe3077ad59e9bc3c0535e8ba3f7a6b545
zc73403123b9d62c9d2b38a322ea220c0f58d71dba22d7ec0c1f712f230a771ce2248be84a043b8
ze0c0e1187e3e114ec4a4c1c025bdef0bb58087a74d9b3d23a893d37027101c721b2040eaca4efb
z7120c64a31aab1be20dbe88a4b53d945649b16d2935bbfad96c95b6e1f7cddd512a662e7d7cf83
zb80794493dafb3cc7153a2318c2b10949da7dd4a84b1889de737b60e1e5589e73f1e0d2dce92ca
za43a31383e2adfc0b82e3ef7029ca5c803853856fb21c0fe677e51f764d428b4b467479dee0924
z547cf53758090b3c505126579f27c16216cf0c5a621861d36054f4f090ff95160c0559830a39c7
z2406c274487f3dcebb17029ce21727678b0aee221de275c62d91ebba5a2a433372f7c2d48cdc1e
z1434337b266478075092a977156f081d1ae272fc4f4d0284da3d7104e96bde7033c903add398af
z82b46857315d0c14771fd0d9c786ca1f5238f21279e7b09147bd5a6635dbfbd9c777286662df9e
z0517c92acf843797a0190f6f4b3faec03e64411ccda47d55a4d4fb0517be2ada3c39f5c8af7261
ze7464e7d0bdfcce7004bb443848ba40bd5d502507719a234a9f6ac6bfb8d7e173a670736afc650
z7a5987255016776fd340b273acbef4a25e7c6dad5d90f6575de34cd16710be06523055ac4d7b6b
zf9dcac664654ed13ebe2f5d0a47cbe80c41d33b00ab57b669f3ff006311f3c2bd6d78249153262
z3c544a22701e859db2b06bd462253d27e76413ee06d94b85fc992d333200607e4ced7e98747f92
zdbd2441d32fb840db6cf28fc6369706a2cb9652ba8056eddeda018a4c5856d87839f66fe0466b4
zaab89628a6c035a636ecaa1557a4370bdedc07fc414ecbab1518658184301f84668ac0cba755e6
zc31183f982e92a6272a3c950072de74aa8a1d1beb39a51ba4762db6577565b7548f4cc24f5c7ef
z17c56ab76f456244d02141fb6a315cd0b946f2c5794767f7270aced089a1feef18b6b689d9cc2e
za78e45f8c0763987ee0093a4f099c40c7d907176410ef2f472c3e4f49155c74d41c0a6c0a830d9
z428fb6f0876f954ff2de69d2d6eee7154729994443e0629e63f75f9e56d8c28abad42c52e75396
z49afcb7aa54e19b1ba9fb10602052de2463eb1de5345f5a8ee6e3db6f7e3604b386dfb490e7633
z5fa5d71fe9d421c552903c6080ca7ae39977f95bf8e51f981adcd3c9a606b211f534d1c748ec26
zdaeb2f439694703bd4376ee5d12c6c77a702ba3922207f5dd02164ff53f200abbc86aa74e6e088
z864fe0d6368afe8ac2714e42e784e5d14d93fe77eae27d9d742d55b5ef92339b1f88c34af36191
zde53e469f2f33cd645f62bb000081350df0b8a25b40fea5c667903e404d292811d0eb0b8980fe4
zeae651afce55bd7492bbbf49447b495740728891f61baf7c3fa16197cf01439faf1e1cfd0b86d0
z8f949f9cbde1855f3ba8fbc47e4509b3c54d59f7b9316fa406c06b7704f62f27df5787d3b10444
z7734ee02c9906018dd95d1ebe94fef8496f8a8743be802ae1eed911493f382c7c3ec90ef6d817d
z0d31a0352ab814fda84c13d67b0d50b72a3ab1ef532b6b10ff8741b5fca8d5be5eab172afb2ea9
z5afcdd5df15eaa4a73f606c0767f1cedab5215ba450e09a0cd1c9b8cc3e444284ca46e14ddb1bc
zd54c79fc9b88d16fd6ef532326b50ca5dd6cb72b1946fc931f0e29f453a9a96e13056ba29e6724
z9240e5c3cc336495f6580c2a0841e6249a95283b96461ae080efcf19e669d2e34ff2eb27ec0315
zc6e0f9d9ea7d958f70bfe20e37ebbbf9ef9c8b463e0d0e887569eecb752ac6876e0f3b894fd2a3
zdc09d3647a5a1911ac2d875b3885e39fc8268ffc9be6ed986297b053505f77db4e6773cf94aa81
z6106a893b3cbeedab02a8e22bd0a566fd6a5cbd394671564ba785a640733e7449d7698187399ea
z3a331a0aeb0f255017984081f0b2501cc0c5f3b000e330c032d74265e86c9994d44c303bc0ca3a
z833be54b89878fde1b6512a52b6abb7d241b6572af13397e2a5ce7da8177badb7ef08416571553
z50f1485d21c962cb16b6e7b8174c6ff94c288bc5347969ad019109e00935a62bb269737a060f7a
zdb3d2291493741e14a71e1677ff280a4ffb64345093eab654c49970dba7c3a3bed9b12787c4120
zadf9f79e3c8a70604dfb3ec319fae51afdd710fef662a28b641287a56546a4ec91d251376fb913
zc52b022965a747935d90ec973ead740a3ea0b836f077c58af33759c32e43ce20072588f44c0734
zf74fe88694f1e55e00c46f77a366c921299d43b7ec7b34991f677c2113b7ed56ffd58345d630b4
z657936d203a1e36819d80b2f777f695f86033a997737b6f2817288ba2cb541507231de70be3c51
zb204486bf8b34ec80fd9a90dec4e0fde5f0a87046af2bc5fb3ea5a54dbcb4088852a597c7d5f33
za9243941c252a9cd51f033e627d15fb509acc86e5e46031abef17a8e6850b46cb4bc58b9f6b5d6
zcb21322d17c87b50a0786c6ce8e0e2a11b126ac712dbb546cb971ae2fddb14b7645826ec22d856
zff2a96aa8b2d3d50caa29d9c3bb9fd6568a1223f4fe3adcb6a1e409aa3b2ce6551aa68ea18df88
zd78bf91ff25a41c878b964fa849d9a4f6e4849e34ce4c14c4ec3895c0f93015881a4521bb02b10
z3a2f57b01381829cf108b38f46430328bcdcd6fc4105ea41be06d777869f20916f6c6cb422b1ba
z9808ffec36c84e002c7406dd927413bd6bd070941827171cd7c943c5a4b5ca32b0a6b20187723f
zc302542b638d2ea8cc42ea7d7a9423dfe4ef56fc82e00de6ec6ff41181d803e84f0037c5d43320
z93ec7bd84841dc9629293cddee25bd7f3cddb798ede10aef2ea35754b68ee856ec12f2858584b5
z2d982aff5892ab06cb87878710d31e3695e094ae00121b25120561f5fe066a6da1ad4b6c06520b
z4f87137d086d4f3cf3320c4c517df596f71f0ea3c0269166fb0e537ba9897322a2733cf19dc09d
zad85e871345223e4fcac1e0161cbbd475ec00774d8e039f2587f26594003a06b25e99687701fc0
zd3f89e70f3312e962616e3cab4ab341705511756d5ad37f304cb96285bd3765e07c6ff72d6102f
z55c4148b76861365dc6520adf89bb114d651a20f8211b8ea06af76ce78b93508863675f09deae4
z31ca47c2600fc1c828f4a3407d38639de3e054cf2c3ab8c24bbbf1cf182d5839b5d0d02a22ad1d
zb3e73ae3def63f7fefb90918acc562379205bb8ea49bf24985179fa07bf907a348771ffa87dd0b
z74437dad9ac0c80c8df4ee45bd680c0eaf18b438fe62b0d0c43b734d2b3067721ae07932516fdf
z362f14e840afdf312b26a5af6602c964c67da837a8e62273d526a59c669236686d1875bc79ae47
z65c81b6a9ee87d80f0e6fc24081377a8d7498a3d4949aa5f81edb2153b89f6a910e54569018879
z46a4b354f4362615935d58e9e1b30f9a171c032dde834511615fd80baf86101cbf4d1f80dfaad7
z531a04727e01c88129aff41dbd80e643f878ef29af2938d1a44cc4c2837f9b63dcdb134db85d9b
zad01fb557ff7a10b679b908125f0b4409f97f7301bfc4d342dc855ff5924615005b0b180029107
z95e9152d551e2e0bce9ddbece2dbdcc09b8a7ecd097d9d2ef861351e52d99e6af0eacbb79100b2
z698e181f48d7cbbb1f79b60f453ca855488c29e9f1ee6167698fcc21a35a05a21267c4ea2ccc44
ze9d6b5d575c34a58fb87605e213bc7d8e0e67da1ecccb092d56c5c6df15040992dd15b19c55fac
z169c5c9fd0c8492b3c2e19b616b37a93b4841e32395f1264ec87e7269c1475d1837bc2804f34c9
zd9e28ae26be1d70f237dfc428af695150646932e52440a25a81b23857269f2318928c6848c6cae
z79e49c0c43667f9340c8d567c6e87b8f3256960e10c4b9626e5b631d1754dc7db2cac48293a4dc
ze29098ea22b6418b578acbaae418c0c0ba63eb00439fe393f7f3ae0134973be158144060dce275
z2cc93f3b35f9ef30a98f19b7b21e4b0835f1b68c8e1182412cab2efb8b1d6cdb9783e94ae62e70
ze960925eb151f835d89e1da2281b4e92447ac603b381f14f98ecdfdc6c33228a8f91adbc71d9bd
z594e476741117ac1f4cd85d0feab9cf4cb95632ea03c43c83b21a9587abc04fed3947ff57b3e69
z23d2bdc92ca699f96a0292150838c9018be445566256bcee248122b7a05044ecb9d61eefa1ea99
z962f0b76e9b8264da635a058dd9ea09a16a8bbf687b6a5051bdffdac8580d86f0894b6a3db61c6
zb12857aa6b5d1d24799f00c63f3aa898b47cd9ec10fe7bf4a16c67437b321f487639a4d045ffcc
z6905603c5d9546a71b3cbdfd9fce39ed940ab46fbfe2b2c8c120090120530b30156dba08d1419f
z1d6bd3cd486231d6dda02a2bb4896d09a03ba98b082666222049b9aad731b03b8d12db915f7176
z1229c92dafcbdcc558270ca7ec6607013bc842edd595c553a5b3880233e77dd6e393fde6246110
zdbf6b14dbb6b4635928984bd017572a86853b8df3844b38527099d7ae587708b624b9ef3c52106
z5e3f0d0b2b982dd7f24abec9c888bdd07727b48fdce36d8cdd5d86f2b759eba9964c7cf464a6ee
z9c6c2b3929eca55f1e185c4ea48c2c04dd2706a7d0dcea138a00dc676e9137fb1b606abfb2dd8a
z5fe394b69f27dd362f82c489440b4f8e0b5e1ed96a1ec3797d3cce5a075fc6830e5a227909159f
z42f1e5ddb3f8531f6f1f667cde0f9525f9708551f4e08f80c57079ceb3cba92554bd99718ba199
z1dcf0dcbd025225a3c4aba6e210c3f6a6d5d9551a1d865fb9de6cc333206845a290266b1cbaf5b
z8f0ac7085519aac5eacf35c00e1860f5037a2ad939280e34d413088a3d79c9ac60c90715a555c5
z47f8058a0a47395c421394c34c0b34136a6c15cd160ff6c4d731b2e6561a5d96b96aef6d021ab6
z12ded1fc7b6d326619d545d6cd9c54273ea9511ac3f2c2d3f5834627a1695d3ea2e9906fcdfee9
z245af5d07e673929c7a8404f70419a1a1a4b77a749bf1d5fb2a53a8417df65b6d73593f8704de5
ze58c7ba42506d829f65adcb9c722bf3a721898e3cf7240d96ea510d7aaf127f52b51dfda2dfe58
zcade13e18688afa3742121f8be441647e2c12c186a68e7a60fdcdb692e420267bed355e44d0d58
z0a8650fd02b5d68fbf87058809489bb0ad226bafd242196ac6c5f66348378c835ebc2f83c949a9
z8923734735000f6f5d57b2c1a42431a0aac5fcbcdb647d1166a434e998ddeed782eba7a0c6c058
z7f2d31b7dc20acee9b27e27639806dfc654176dc7c1d1b8f00b7a28edb72f6f9974ac9e759926c
zf0d4b97415bf05485e583189c640c786d671bd89ff7faf1532038256fd14eea4cddd2ac977b4d9
z7f41bf91fd1c9c9f57d7916742a1adae7fd2d0e793de93e3a43d5595a6fd888dbb0ab5a25f81ee
z450da11c02ee4f53ac82d9736e90371674fdf5c03b5424bc6b1f93790d6940470c3d02ec4eaf24
zfbe4319b600c20e9c5bf8943d0710228972b8096eb814574a9384c5abacc0912469926b3dac72b
z67e1e89d2c3d34a628a760f0fc58e2a8fb31dfbe9aca7da1ba7c2c30451fae2d218bb2b9522238
z9f859272cf47fc8f54025782bebb1fb25694ed72feb5da490e52307a60ae5d11bffe14e378482d
z90390c1f35318bfe667d72bf72f0d2e3d00e090ab7e576e0792e9be00427449ffd208d82a7a3ef
zc2c27e0a9b347dcf4162ea63cc0d329ccf5144659f2a521fb9faedb39b9913a811f6d20100121a
z84838c109496e7099e3c79c3681cce05e4c9da6eed8c700e899cb86a4007b9b68278e4600305f8
z367020e15fa7c19bf3a4473df5717c5bb8893b775507e01fc426c0ec3d948e198522f87dda7bed
z9cb3b7d202f7d12179c555f382220ff56c7b574dca9cc0d9cce793e808bef266ccfd59960fe971
z1ad1afc55d1f1a47685719c5ca59b04abd042ea38fa73c91383ca756d0669ce4402394c36f9f97
zc873eb4d2b34bb90ac66bdfadd05948c1bec70a94fa70c5d24f03221ea6f612b219607dd000827
zfdb708c5e3f6f767aebed49dacaef066b30bd6596cfc348e06eb29d77d942010752444688c917d
zf444bb9f58110f33298407ba34244d10064ba39ac3ca669df88ed81c9829cfc893af3bb7728ca4
z9676105c4fd12f1c6b4b0b27f958dd79f6e8748d6eae2853c90374a24314e5d16aae71e5a9b58d
z97a45789bd9fa5ef7fd63923e15d7e533f41a0a6008ec4e524a704c7525777ff2a36fd3e0ea4de
z093d43518372c0ac37731e508e0a05b70c3fa5fd8e95191783de4cf779c7c6f3e4228027c4a508
zcbab81bb716a78d3811c8b79dda6b4af5c0d85aaa7d72077051db19c8a25eed40c344d74a0f757
z6fd82679d242e391c41b6a0b51ae28f6aad60b77041e6daeb94c3ade17209d14da21bc41317b57
zc2949a2ee97aab68982d2dc6cb3779bafdf7cc92f62729670c688dd0b62982cc95629d723a74d1
z8a24b7140c83f4b93430ad1e68be80ba47979d15ce4a5ea33a286996c352dda2b9aa64791660e8
zfbe49e0de49fb28616b67395e9f46ba6d9ac2e3e6eea4bf4ce183630a3ed4d5f83b768ad9e002e
ze0b5eea46ddeefedcda59cf56e3a691cdacccbf4304e2c33e113ac862f5dc2a6c55d0bf0c85139
za1ff6e375e1434e9acb177198467d7ac476149cd4711ae70158acf3b0705cd08f300126288da37
zb14eeeb68019aabfb1884d2d036186ad325fe06c8449c493e3f7a0a768d77966c216e4521429d1
z02ba50f50225446c474014a7aab65695ce1ad1a50135e72f9bf4e46ca90350a7a8b93e13e6bcc1
zefb0e160e7e16f05e4edba6e8c1624a3f1ae32f1cc0795fce169cacd66c488955c928fb311a781
zdddef0e563318e16b20916009d90daaffd7f495dbda90cf37c580d3edac6ec2dc200de652b279f
z8fd910405bb3099e9200b5029210235ff5c6214c76f6e879305ebcfd0f6531556a4fb10d1fde74
z8aea3bba49c0b66d6e4f148e312b50997bfdc204df9eb258d4b36142c3e15672f88fb0ca2583f4
zac486da6ced902974453953da25e892c0ea3e7065a2114de6e9b380c39cfbb9a11184a837bfdcb
z0c39cee32a53642fe53fa77ce42bd090b7706458f8824605bda5976d0d70f13de9187765d5edd0
zb39b7a32df8798c5ef431d49387d4c9bfd813b5cebae6191b5f60ab6d93922600de8b201d9fa88
z70b849548ec83b3174fca2181fe006b0f03c85edea0f77ec49f9c67ce39896b82eabbcfb754013
z6ac80d0d50bd9890d771c0d1f3fab643805fbbaff51eed28e843f31add2b8aa3ff7c50df216120
z212c9d42ad3ddd124bbd7558cbf7103c5df556e81a0868dd324d55f8855fda814d19ec9df88304
z8e22425a2dcce31cc2ff61e314408020e5deae0dfa22f3d0641bb3edc1b2364d9eea62c3ee2e9c
zd6668910e50109c9ff3f24ab3cf1b0dfe3f0d6bd1ef1d1f3b264fbbcb0c3d661bdc53e533f29e0
zf57a7d4daef10d33b355901d34985c6c7a19dd4e38366b0d2264859ca8dc1a1829241b73c81286
z2670a0c6b078a2186ec81070eda8f014f585b72a67d2dd9a3474e4f1e6c68f74af07c3a2796e16
z829cb664de48518f599d1bd0d1e47ba6fa83740f8ef229f285989e169210eae18ffce7fa95d553
zd43e345967b722f9bca5b42c9fb7b1f6bd73e3415a2df3c423ab68e6c7c5c0f4a7bd7c823dba1d
zc92bc68d72274793a5a2b962fa4dc41c2ac0b6279a8799dfe5ad21fa2eb0381a3f3c485185f2ec
z04a113ed11358754eda274d6865f812802b76aae4ebd49d2df95b5fd67ba973e0eab32b77c8c77
zeb523179240499d9a90dc8f34f50674f0f68b5847f7f4104cb8d3e41276be0e4dec63a1f54d064
z4a64413f8691e3cacb959b70229cf96b271eee6c2b97bffee71b5c167308b1c50abce6f5c459ab
zc142815a159066bf32e0d776d52f7bebd1aa8291d568e3fb187b9ffb56672cc59043373e8c6ff7
z167d0a777c891acc06d9d9f1bd811705318aa05956f3862ce20c23b4fbcd25eff7d48f70608306
ze4f079bd41ebd55b5848a7ab5e3fdbf268c5746fb5d86d89198b8f096ef8c6b75d625c502db91c
z40fb3c6980028879d285721d844705ab025daed9871600a31a589650eeec91dabf3635e31f176f
z5c395d57c9d15b7742566849f8a106f06e45381a006cd2cbe562c70aa4da5b2f3858d15535350c
z591238a7a6ec42abdec23b25f5c09f76e7e7059cb97a0d408cdce9e34f9b12ba01066b7b118e40
z7b625f717fa755e790d617b8b47e688fd23f2ae1911e27fe979eb00358ad1ec3fb413cb5822c8f
z452fffc1f1b8c4c09c866114be511c9afcdf7df199c4efca3de4639e5ed9247047f4296d0d9926
z78008683fc93457f6fcffea52396a88610ab01339153a5e8c568e1e2b50b615cd2dc7f113ee77d
z5894f1f4145dfea23269eef6d14dedc6175a48246c91c7ed8dcea260fc3dbd470e629b50ec3a15
zd0c2af5ee71ded6773d0bad6215eab78348c6c1e0e00f1648dfc6a9816fc12b46f86d5aa27956f
z13db9734049edb2c22e9ca473149d6681dbce56a3796b8388017577f57358b548d3b23e5e5b26a
z8e0a588d15cdc154213db326b562b8144e59a58d5567ba27a0f5e7924b8ab221020db49cd1f56c
z00e42cfa0e54cc3f3133012e91b5c4f3481aaf21f5fea6cbe206e38439e6423feefa67a70bde5d
z7fd5bc5303217159dbeb3fb2ed60231c0da48f2c4c48e3e6a2a555719f6cdeaf37b177baa1311f
z43332d9fbced2429697084dc1d9dcb26c8b8f7d96bc3ee781a11ef412231adb4aa80d12f5c92b8
z4221bdc4a86f4ca5f7535eda09288c195d9b77041f4d945c851aa3aab2c33f3baefbe0b6ba9092
z7aabdceaac0310ffc3060ab6b1e448611ea91b10f8a03434b67ac787722d6c5babcfbdc7d0d3b2
z7eb2798f816e44e151ab0a1a8c01c1517f8df026235f6c3633aa6d9ce8594727f1f6984a6c728e
ze7d88d47c521df57bc20ae63433c303ea31927720ad197b8dd70594ef6d7b4c4d49f86083c7e7b
z1382a254fa7bbe72aca88491086d3ac837c7f35195c82df900bed80bbfae7f22010a559c00d1a9
za7e70b1000865f63b3fbcb429ac2e14373dafc51ae22a5978f7c698f1e3c1b07a9533e74ccb99a
z8594e27051ea2dbc27581e3d37df7e89cc8f5c3574bf4228d13ba86e2457fc0e9daaf62ebcc728
zcb8eb71b7913f5a1177b9813cadc0e9bc7135b05c807e450eaa1bf5b6cf96c0eba11c41356c7bf
zb804c298c5b8d1e739093b74ff61424a29ba65dd1297c0b91ba9e4154cf33acaa9369205254ab9
z323932f5af0e1aeca005476b05470fcd0833d305a39f887e2a6457e8797b5f251a7046aec5c250
z0a2da723ddb037e7c68369a026886792f38e0b43b2286ff2a8f685bab71a6f888eb5045c62e6d6
zc8358330827415b5c70179a63d62749ecd7fb9806118fa88920a61fcfac358eb8f134eb363c580
ze6eb1f55a5700c4a4b8273b7ff30df087ac508473b8e5ca501ced61b7b9f7892a3b8c02a3164ec
z9d10fe99ee100f5392dbf1af04c4b32a2d58cb9d0fc7a0bb63096706dc2c45c764e5dc01ef09af
z21c81fef6020245cd0ff40378811c30a9238f1a1a10428ad281323d8f6df14e48c662c401d56af
z478bdac094057beee335ab1d09d83fb2c7fd16402d9aaf55d7427e00aeee2bb459374b86fc8e7f
zfa3bb34eac519d47a93b3b1f0a473739ab3f468781a0e1a3202cfd10d469bff53769b709caa6ec
zeebd1609ad0cb914a902f8c8dbf331dbbbeafaa610e900d123483e797d2434d232beb39c95426c
ze69145b78a29256333e2f2efbe8257bf837b737545a9028f153a9414368b7abe9c4e37c095bfb3
z320d2f96449db7ea646708cd42786ab4656eeb7ba01058259fd4b4ab88213a5c606bac6d3e98bb
z1b831d40dd10850c49beba103ecc9b011f88afafe44160b67553552f133f2075954b37d57ef6df
zcbd07e1c2abe8ae1b6cfde0cd5a631d663754a4806612d8d76edf5701573a84e260204bf477047
z4d4d872d90eba6fef100f93be98c7e1bda24baa163c41e36a85cffa478793dc9f4aa6019ccf23c
z97c5925d3ab62b86025efe2f091b427fde4c64eb96238bb0b963058efa217c766c6275063b1626
z2c863d51887d69bed7bb5096d25b11b2a879a2f94fa204e4f2cf517982ea6b5042bc47d10ab27a
z0c154f4e556385470fda21b89c60e8009611ce4e5c67b59b91c911c8c92c1e69248bcb95876beb
z9249cf4fcdb48835015701402070569e03d927c1c801d00fbe0bce81d9ac82103fdabec144c35f
zb3eaef3a6d2669d0631897bc197cc67e1d1568c9b9019ecd8d1995124e2609d371a525eadcd359
z928aa96f8a6a6941836806fbfdf7ef170eec33f2712de4eef6e40e412ca3bfc20c563658ecc4d1
z091893df429f4bc3abe5080b8ee6bcda788c4a0d3c79b1ca8a918217126b28ac3c48962b229b1c
zefb3779f20a78ea3d597a32aaba2f75461356d92743d983db3edbcdbf486e55e80cef8d35980e1
zd1b2e976a3b975408b06f5abe7110778e19afd6c2845c71bdca1ce7e964d7b6541a6e263fb3015
z904b74354d868d60dde1ba9e04b0a416a73c41fed117e49e1a199cf290bd2401759b98b9dadc10
za8dfcd22ba94abe5b1c0cff8e40838e92af63b783c0ad98bdb85e84728a1dfc4fd6cc26470430e
z71a72191e4c3889b7522bbd2e6b9ef871b24eb83bcd124478a25c4ddad1b9cf6d005386a15f546
z0c867b2a4b2d890be8e9a1f1cfaf8fed758fba1174130357923d527ff1f0e99cd150c268ec03ff
zce1bfa448bdf49a4eb8fffd14ed817e21c5c1f07855a4e6c957844e17bcf0b2c59063ac8bf19c4
zcc596fcd6d5e6087d6dd51b0a1436f3e9276557ce2555edbe9fc232a219a56dac3add387f2e035
z28ca65699ddbb08ca23e2018c19ced5543c8f5054d803b02a426b67680a5a6ab245b12af841992
z6ef3a41dddf30298af2c867c13b1911e7f32d14bbb08628b014da86812b681d496cd4e2fc1160d
zbdeac37f9b5efd8ff67d3bd8f088d489158eaa7fa1122338029f1c574f0c0202d4a4642c5cefcf
z915ffbbc1345ed2a7944ea3e627b0c9b88a9a52d0d804cccfee0df6ce127b5efbf8b56c92e9528
z527a751a3e135633a1a1970228f7a7560b3914a24d27fd6fbee5cc449691dd5bb045fb490fea2c
zde7fdd5a19709fbb1ffe1f339a5b5aff50c19a047d90aff0c8c13191c6cbeaba3c2893de50b914
z9ba3a447dc0566c71db5d1dc5c673bf704e7b649f938486c1f5c65558df2281c974c9002b6e7e7
z4b8f3bd1515b0e9cee7b327eae9e374af4e2e39607e90e017873a5da0b3541767747232154197a
z791dc218523974bca282cf11c2bb9f6595bd681298860aa4896d7f6478863b233b1b63ef3eb0a5
z61071a84617214f391009dd196c6232cb2d9c50bba89927d4679a4cbfc14132446cb670a3303d8
ze971ed622e13d31aed9ff7dedd8cbf6713a7979fa485a3e3025d3343dbc0a931b864047d346dce
z1ddd507a155130ed971a843014b9838ef2ce929bf8c170b3ee848700013fbde8566d09e73d45b6
zee0e78c8eed6d103cc8cd2e570a56c2daa249e26fdcbb972c7d7d0bbe53c229e844148f7ab136b
z13fbc4e753353c270550f89fccfbc98197a35b65156ca44c19b80f9519eb97f4e11961c7d6ad5a
zd7b4c6bb19b57637d0b5538a4c01137c1719b24e36703d19ad52440845b9badf40984d9c34c258
ze9a1a0f14f28ac62701ca3c5ebc9b7f24e78596c901784a14cece0af22382151972692ca4785db
z1a663b111cdfd9614d9565af4f27775fdfcf3a28363d0ae58d2a998137eda8907224f291591ae4
z1e23ed0621dd1a5b5278a590b338d77c8ccc7098120425c00fd48f298cec88479db51b26547926
zd003468567391a7c2c646b5be6c068678b95a86543719cb18107c16fed731134e344bd2c9240ea
z3fd04a5babdfc66d7cb09a78fe29b1de75d73c88f4ce15e8eba381e74ec02e52ede1d0fdc2bc4a
ze07cd3d93d02a5aed91227ff0a86ca531f56fbde3e67abfe904ae4aba93d3b44afb6e5c488b5f5
z09609e8e9b3d98b9d2cb61dc9a7ac34039016501c6876cde04c0d3323fe6f1f4636e2901a30b47
z5a9028f21c036b27372917fb9618413f125f07fc17c1d6106c4b5f155e08e80db5d31b77729934
zb4a2c157c1d03e2fe53ac7d7f4a3ddd3740fdb5a8b098d06eb3ed06ae0ef06fb4e3b5b09ff9bea
zde8aee335ba323022e214441cc9128b17c292a0a0b8b423dc6c0294327e97288b437fa682aedb8
z74dbba85b5af22c8fb6078d7d076390c086a0a4b50b31fc77f9fead43fe18e83441ab404487e52
z53e353ac472651dc4d60560906771d0fbcfe381326417c27a78cdb523b8e5094261ff657796a82
z701068e49981275590e4d5ca9cab6545ae5918177b655d82308a0e412f749034a943f02c34ae64
ze0ba33f68e1896d1ea03dbf46a9fd3da4144ed4a2328b50dcfd0e96c8dec30c09c2d06b4a3ff75
zc2dc226cd804f02925188897d8928a90c28b276a0d3ea511247a2d498adbf47b288e59dd923795
z8d1174b83bad5b0d94f1babb02ba8944b4f96d715cac4080d2cb7c98f630d983955313e4f07b24
zafce7c62809a36c5953d3ea9d8d27654dbf23cdf3b6f4f2ccaa7819a9a095b8cd6629e7ab3a8a2
zd5a87202cf639d37b54de41f0f6843481e33e99ece2e50926801743e05897c12369634ee85ae5e
z30eb32e598f02bca1fc1a4fbb1c2741a76b79bcffc43ede5f340d45a58310e88413ccb34ad299f
zd29db05877fc255df736e6aa12d621933f7e8ea6f68564ea562dc6cfc6e9229d385b53f1543e6b
z982c514804d5d56854179bc2b5fb412d7f7471993c8854d7767a8920eda09899a68d2a1c3cebfe
z98e4d0bab3ba4d11bdcc7f672250248bd5366093479c7c9bc81a04a03bc61375b40e839bf7230f
zb96ec10417531bda3baeaf77159ec6a0a46651e9cb5ec3d8e6650a336fd740922c5aa14a979e4f
z544365c33bca429c397bdce743e699fd09ebc3705d17ce024f34eb9ce62fdc6f603e9d45a8f8a9
z32209169c89f3d0692cdedf322c8cadcd50b0763f023044951df035d1229b609c849ce51d983e9
z0c8eb463ffa69c9c5546cd5212617469798ae508b2fc0275847cade1fc2d293f3c172a4d08502f
z0076d7502bff441be11ff41d01bb9e72af4611724f15414ad7f7e044d9568347582a04212e37c3
zdb593c0ce0134b2b32bdae8fc747fc62d3645d29ea2aa06ce750acacafb535a9040a69fa464bd6
z948ff4b6a9bbb2e08fdc1d0b6eff52c5896122624faca4e21307990df442d5f0c1e1c3e878dc5d
z06c23dd147b6e3f29cbe45350ace431e198ff3d9bcb96f5082d39990f8d9dfde4d256503048c2d
z5d0402fac472e74eacb9dfc2e00a237449ffa4bdaadea26d350c2bf0b5addc474d606dfe113ce2
z6c4758443ea1e036cc045dbfbd5d06078dcab55a703d1e8da37e690291996ab5d6ee14f50db190
zeec68f4749f710e80242e3e015daf07e8929b8665a4aee1f9c770fd45a8e7ee4514005267c991c
z0be7b8532464edf76c53af719a78aca5ce628f0d5f4dba90ca09410e85e53df24ee5680f545204
zc3b87c9fde36f6f992375536e847eef6a626b7340291a839357dd83fb1ee0e977cd3bfa5291e90
z7d80af190b5daabcf1d2b9baf92fe34076f0f94403c94ff977618c24bb2dbd141234043cf3f579
z1f48455454d08fe900e0e59e2454a33067c77f109927916c2765f73b1824eac31e8c58ddcab26a
z2955835a8f46d031e65dbc63483c13928f10e763ebf2b90f963ea2a6f279972401284037ea5bc4
ze2f07dd170ab8cf3937253fff880d3fc65580030327bbc4bb32817e14a7d2fd6be03a968030c4c
ze02f09aa311cb7d4f7934db62988b99cfbfa30c7a5f0e2f342131063d8abe3327fb9557f6bde42
z441095a54ac7ae42070b5835c777dfe94efee01c6c5022f01db4cd9d6d5b67f23bbbd3968d82a1
z88abfc569485745c20697b2cbbe24f5638d90f637abfd4f1db93847fa8e3231de6f1f58744d7ff
z0ed5c7ff1fce9b4456b222de060986583bac0bb06dc8f8f9de4d9274068b14405022d9db2734d1
zc9ede1c3fd1f2fad0588a086c708a1cb39514ae7a540948bae14972699391f8eda4822b2527eb0
zf77d94e9cfc6836152479eb0b9b79d75a3aafc43f9d7da2f4eac5b6ed11f04f1cedc76a61eb724
z8e1352a19353017a967bcd116b36cb7b79adc839a09bff4222abdd62e3b65566dac7fa28f769de
z02b918994d988b8b5d12d9b921a3740ed31543b13520ddeb9e294e90559293686491ef1f2d6a66
zfa8a35f95a701ff8eab6fac4b6b512bba8943b1633bfbc594ae5b9511ddb1478d5e2cacd055f65
z6415a7c489505ad57a35829844358c4c9b5edbf55be1728704b82adb1ab590608c7db8813e8314
z099f807daa189fab419a3f98e82b6dd8803ca4732ed8eac075288cbd85c93f3689d7da4ce0e10f
z6264123ef08767a103d6caceafc3f2b7c357ca3badd8a9bd1de39820e7075902baf2c74cb53ea1
za5c2797e3ceafc78a19c70e13bc940dbf18ebad15c341d173ea3535400b845b364485d2c8e6814
z345cce849a92e81d164dfdd79ab2bf8e2fcdb41199ddb48045e7e21adf5c11115897d056e1f8d6
z1d4207aa364c0d584c5de71010fd302a78d79e2bdd4220d21eba06c50cb0393f21a886a14c7956
z5030f49f65db1394d5868c19408c76051f0b089523c6174635bd18e06c4bd28e1319e16e8abe69
zf55e2d122b07ff5d8ddb5eea46c18492d38ebe08f18bd3fda52e297e764861e5a4b821acecb6aa
z2996a9c2488a575497d0eb7f9f77338f843923322b1da6877dcede869b4a4a6f96dd63631af93b
zb6b8b9f712b21f8047117d8ce0cfa20bb3a754820556a78bfb9b5f66cec3a53a14f610564d3d06
z692efadac0d5354008479349821cf7c9d6f491a0d7577c08b11493ab3a752b748a424c43ea5fb3
z6764ae48e5237634218da9ac9b9208e1715daeff82c6b6c5238e2b3bcc3c49de9679504b68ea02
ze48a73dab36025f6ccb8491b3711f0bf159cb29fc7d517c89e6ff166afbb793fe04852d3ca47cf
zf359ed967858547a038cd2397812f3ca275a5f12d971378e5f83313bd522dc3f9aa92be9d9b415
z21db32cf54f4a4334fd7a7784f401ec5913b42d7f6fe2cbf362b1c1dc1f7ba851755f306930a30
z435ebba957536da7115c4a797cc457baf560c8859cf1fbacb1d831ddc78717852f5db86b0ac190
za11b805df1e81b0a3b18ffd6fc97a0a67fa6e8b7b19ec45889b787cd57b1b8a3457f94cb115868
zabfd358c508bb38857e08e3aef8948886566e5c140791bb208bee700dbfa4fde600e1c1e5154eb
z1927957284cc64de6d4f5c5e42d02bf9997f94fc83bd72f56754267ff18b9d481eb0a8ee9a6746
ze4648086a85c275f34ec38738b7508147d5da4c13b627bd46f224fe166e8c4a2a7969a128bb3cb
z17525e839a232e7b9a1edbe02624e8cad3d71d94d1a54530d5a274ad59f055c462e6d19480c98d
z4e75f0aecd87244c724fa5a0ab66f9e3f121732c7591f4b0500dd768cdb12582c44701d58e9452
z60a349ea5ca866605a5bf592a093a956e76c25d0894ca77edddc3928a4ea014178c2c870c3feed
z0854781b715935a9b5a9d6cad1e5f262d24e54525b6bd018186cf9e898f0b892b85c395d39f7ef
zdaf00ffd1989073d7dc47b8e6bcae5f02cdc59da14993df1eeebddebc216f5179bb66625878ce7
z1c4e2be87b584661f296fd69fc8e4bdb41bf280a0b9c4be1f7b4582960ca0d79b69353c958894f
z4cc843df10d14b6a3a83911b030c50f4ffb54451c47e1ea3dd3c4dbb1ffda833e0921c2f35e210
ze862acda8f4c8d0e9d393ba51168b40b6933384be60045b87aa5d55746196452ce20500cee70f1
zca0d1c34afa2642c4099af558f59c735895c344e17d5d07f76e8560eecbf2949d628547f570318
z9568d63c9c054eb9d1b0ef302c8629ef59906c455966c0175fa251f1bb4a6230ec283028099ef8
zf6a6da2e4eaf83ce48e3497650333031c037f09c0c961ec25410740502fe9bcb547bf91db78987
z436e21fd02a4b848cb82214369b68ea5963f4cdfbfeea9e7ef6087ea57f564e0ff31a7faaf71d0
z8b70e38ec625db2a88745514161363ae462842f5104e7e7cefc0d11a6130e3c27f5e7bb7f9e37d
zc9426a7eb9a98176b2e52f0e6e42b70bace6367143cde50fb6806a3575ba6e4e6bd06ae265d2c2
zca3c322f24042f59c2e832c28c15bb1e840cb5364870435c6904ef02bf149e0d10d138c35fe7b1
z5aadffd100ace91b1d3e6f93a57fc16c373d42561e060e5bcd0aa24311a6328cf36b009619f7c2
z530643af16555fca18cc7ea3a76c889b4e44c79ce512f70432302fea440a53e85cd89120ab57f0
z898ac6c33390e3b5720e591ae0c11e6e04194a3f6c051e6951165e8f1c2eedd725f74981d6b421
ze164956d0a8a89132fb6b0adb7be6f455370a85764c49de04f3726eed848c1e037d685c36832ac
zbf11218de7978a871212ff01a018d1910b60167b56db1bad44fdebc4a2ee22c15dcc42ce2b8b7c
zbaf9a9f6e666c8878a2cbf8a1b87e684fd8b80ea99e733d12b9b3dd72ff338d369b910b456fdc1
zb6495332763d8b84943596937442331ccc7ee97758563377f2adbe20781b215d5bd5f91c280284
z35b0d9a5ce8ada56b354b5a2331790513dd68627096be3f70ab928afa303a3f10e7215e132eea9
z7fd0c89f76718b664a72e45898c470d8c3f6a66ae700fa0d3c315c0db8d0813351a2487f26df7e
z1105e2b2de30d4d1f9793b3747f7a1293edfa1ffd456d6938f9993d06bdc0cb7b8a69dc9fb79b9
z0543878000663b4b67b6ddd1a5a791b2354b975bda6ea839e6afc38388a463ea8b035868f02bd5
z337c9269d8983bbaea6a0a17bb78d905df20721917b7032acc0d499f0cc3a73b6169708d52f6ef
ze771853a0a8ee065904c321d9b02f6fb8f87b5ae325a872fad275940f1fbbc204d6f70ecaac351
z8c5de3a8c48f26a846b97ff4d124131e02c2ae3f7df7c3044ea98dcf7e5091f55cb4e14d67680e
z308e34af3087a37f699e89aab1dd66b0f27c11d496271672ee404eee7fd341b99e9622565ebb4a
z382f535be4c1735fdda5d1a555793e7233639090b798585ff0b6e87bb2653c788da09241f57d08
zdad257234dc470de0e6a1ee664337d476b6df1e4020b7cfeda29719458ba13f4fa7fd7e3712cd7
z5d9b16fdeb759e7ee4ba88f1c42a8d1a029860a21460e6c85fd4541631ef10f92477b5c4a5d237
zbe8552a744f063a8f2c9719a5f2f0db4edefb692099664e15b6b826765c53f56ec2100585eb17b
z9597fc3137ffcaaf1ecaad2640bca245d62b331c9484b6a56a70ec969e8bc4b8e94ff8606980f4
z548b7c45736e6f3b69d6898658a392dbfd3475f74ae0647aa839504b4ef1bc17a00313cca8ef97
z1aa813df044e07f0947e342c7089dec174954b331f111fbce010bf736a2259cc8c38f13c9eca8c
z5d35e470eca3ddcfacb1efd50eebd2c0151ebbc645c0843057592af5cb9629be61d9561c1a2b12
z30353df9c8951b21991404f499a7cbf8c6c990c05c4f8cb3a51ecbf4831c46f032830b53d62c21
zd2606cf60b6467219d10e51e89c027a36f5d4c65ef5f8b9410a5bab1d9a6703a34643227e92fd2
z6c8660ee160fb23c5e03adb6a0878af35b55dcb056a4abeaed5a03a1e09f163dcc87f639cbbdc9
z8b2928acf87c839f7abb667b0c8716fdab6888c0db24c84bfe74786fc2f06c8be7560e4b7ee023
z50a28f95a9b736d1d19557206ef6fbc4ef6e6210479257adcae66499d8f5c0f187a19ce97dfd59
z6f94361f403f051ef555deffb8f500b38a1a89051690e356e0be58f6e4dd205aaec71497bc0f4c
z3b71ef12ac18f83ed3541ad724ad8a42431367b20e319b5d2805feae1d2d0bd1ba58067282cc01
z86b61d302fe203634ad5ab947e987dc05d8dab32ee2b7b21ec127f72162eb3ec02bd3f5345abe2
z3fc1ebeb5313fc27c1ac4644008e884f63043c9097034d930ec23325744bc0f7dec91e3b34e4d4
z64e61e1ebd8a00eed1cb16b2004987070dafcae9a14dd5d00eb65b45814b6d6b96118dac6c48bc
ze0660b75f5aa3084a0aff7433472f6525e8d0422d555a4630a8ab312fe40bbcfec2f26703712d2
zcd4f4a1a713484e552f025aa936f727aa529827728f14c83314151194aeb7ddfa8df73490cb69e
zf3d7da465e82884d8c9c299a780da44cf6cf6eea0213174e45f55e59b76dad9ffffb2c94e06d8a
z11f8fcf5f82f41d438523005c1f20aa0a62104aee548850723e78515daddada49f5c96374a2f5e
zb0e77ac6215fdde3b7ec54ff621ea0b86a561c1561acaae0a3f7bd2946127219595be6de6303ba
z6e142612285d4ba3e0df56753fb007432c42b88686bb13d812bfcd63962b0bb11b375233fb9dc4
z03c576fa1f31231b56b91ec394175cb7b0805ceab56589f8c726e36c7103f3d5699dd8624f751e
zec586cb7cbe638f59febe407127c7a1482952da5490c1d0f6f21fb34d25d63fdfee28d67502632
z1e2930d86f0a04791dc75d6e4d93f8c427262f1242584eea04a16031f8ca8d3ab6ca4845da90a3
zedec3315676d7d4be314e6f80ed5789e5724448468c56aa196e99fb795639796435012cad74364
z50d3ce7638db239b92083359ba91e9d282f1d638667ccac0a9d2a61cc4533e8960b92716494ab8
zcd1814148e66567aa9d59646986051f102d2b5b5a48595fecb0266996ea4199d9a011d2ea64f6c
z346db5d2d3d8f7ccb9b77dc5ab5da119412980c79a487c715bd757636079c6ef208c3a19a22095
z279c05778490b36103a033a818c0c4d154308db314fcc6f4fe607791fbd4fd4f7a4271a7b61c8b
z6185e19af53daba7c4d035d3ab29d24708733d5683ffa6bb1a40d2f5415299013b425d7acbfb38
z63fb28b4275df69d50d8054ff7f26bdc22edcad7397932d5ddec67eb966002fec555e2d278b23a
z910c98a9e3a1b4f71b9e21e3251e6934143f09bcba2e74e9e2a91bfa823d1be50e1f586adff4a4
zf3c0d8f3ca7febbdbb3022162df20ca33228f3e6ae8e1afc03de351814804113001259e7fcad7c
z56a9294c28f46f53078f3a1a3fff555b17b1299c46887025244a00a10f09c0693caa9867403b0c
z20db125ebc638a78ee9f6df3b3583a8edebef747795e6c292045f8ac3c6ca4d7a1fadcfbe4989a
z471f4bde5dfe4e5d86f52e3ea1228717d18291a707942b9ccc1210ade4c9affc47c2f30523eae0
z151abc4a5ad3b614306e970713cdfc36c2b78d21d59ec30a4e11a77e9d6979d27e0cc519a537f1
z7afbf07e89d11fe1e0453b4389e97aad884438b7770a76037f0647223b3325542b51becfc6b050
z9b7a113fd028d394b3817a8b2108b7575980bdfa3ea762f83afb2d4a0bfbbfd686dd96e122ce00
z1616f10043b88ab4c32cffbbc108dc46304c1c074c77845bee77ab010e285c6f1c1508e1a96212
za2803d4e07154e6d8585497ec589afa0a6b29beab737417601adc6bc24b2102c7a57d650468e1f
z7834ec4f6ec361f58a1e72d63eb763197a22d1576b495626ea05c42dae8c67550471d1c4b7654b
za51bfe93cd4c4e5c098c913ec2b1643c18bca3efc29b05fa6e778af2ed118c08294e373cdc0f9a
z744a44c7b039c05c2cfcbd10bbc8b3d476cfef475c39b7e8b64f1a949a7a4d15e4b2694eb60145
zbfba608f872eb69f2f22c8fd48e56bf28037ff21e81c1f6fd18f89a69abd2e7b3f5a259b52e713
z230c43182169e44463ca45db87899ff13999dad01f60c453f79737ba4bae6f2cb495c9d869780e
ze81b964a9315d1edeaa3e0b3602f65c227284f4b43492b23cbd74f016f5a3de7fa98c7c0037c95
z9f0b3f3978b0fea760046760a65c02375c373aeb5542546ecc9d5c322779e5692f8311c17e31b6
zadf60f0162186d306b29e3488077a2a57349f4e86d0fa43a7bc48e8d923c1258de0ecf0cec5240
zb02cb720b38ae4c298f390ce26338d4f3c5af7a089096addc262cde769fde433bc1322d3131aea
zb90e6401eba665b8308cc0c051363319ae97d726ed6bac4d7c4e42fbe18a3a33c3030ac0a0246e
z7421fca2b86b8f5656eec592f62eb1eac6b3118902ea1acdd787f627b51dda9137f8eaa3ff7dd3
zfada6db746681d17af476f362430713c1e9997e00f67ec6a91f823746e3dcc7ef11c2e6ffad984
za81f86763e9ed264236bec3ae38275d4cc70e1a3dbae21ed1dbf8c631409005517148599c1d861
z4cc4fd20906e905a3370633bf9d5034b4c4cedb14aa4cdfd040459c202966964f006d75d8f83ff
z5647cf707c07d6c1237a524980f0beabc77190ee5ef1dedba1a3972861ac9b2896eb646f276138
z3a2b438797c1fe4d53b1fc0fd36510a33f3b1a2fbb8bb5772c0abc5e1c81e3b1eb8f1519d0c714
z62ed9ab546d08de3a63e591ab2f991e3fa5cbdfbfcbf5d1b741c1dc1faebb3f5d89ca01c620e62
z2f8ddb30dcaca991493c6b5c74a095c6dd5fe1eaf90ab33f0c65bad10f7164aac7521923d9e2c0
z2f4128ef449a6591706f35ccc61646fcaf9cac3139c9185480fe8e49a671985cc070455a3f99bd
z8cea335089b4c6c0d2fb564bf4e35b61fba710652257317cbd1becbdfd998db1f48d9bf8d2dfb2
z18c3ebfc8bbaaa7d1d92e6b09498d0f38489af0f54d77321a1a96702c487fed9f33fe9e708c506
z9a70cb143a12fd5b8039e3d05d8a17ccab75a3900cd06e0c6d34f89232fb3a395aae49b51ec2b1
zf2c2d66867624b49353f51273670ee70ae4d68d198b164a6c3026ed689a94aa94d8f7617a36435
z6e0926dc501baf4b7f415d594317bd50edd1a8f192705497fbcd099a2084d17ddc224d49bd9e86
zfa0600d6ed263e0c377577579f0d2d032b324f66e0c9e8ed93aa052e4ebb3e1473f8919248c963
zc6414ad71901e674797a2f1505722c7a038e5bdbcbf435549c0c83742f88c4c1bbda45ae77bcff
z60b7562ddb6c38bb431bcdfa256b991c08363964016a6fbc042f8c2b96e6b88d47d853be2b935a
z44697c19cc7bf79e406870f423f29177e7ed5b280e388c7c4626fa415b1760a3b35a3634313aaa
z1532f989e1edd71b45ca789dd57cebb86ae5189131a9f7dc5db0164f077b5ef02067503230b7da
z59ec167381b2d6b90a570f10ba4954e670b5a9b7896e4e8451c4a4d48756617677f7f1b320d4c1
z4bf45f99d5f80cdf90ac0f67c07f9470e5093bad81870b13c5273685b18d1b67dd6baa2db74f4a
zb15c20884e870b4a5a3f07a2cf2e3899c7246cdfde236d7143b29edfff48dcf0f6de645f720a24
zd62aaa7fe9a282dc93247f735bc1a8708236967e1af25fd885c68351d780a1582a1314c3b45f51
zbeef60f56ebe1e94aefa9b148c296b5f3e02dfd22254a0f036f9b825fcfce8c1a46a2682bd9702
za81adbeeafb3bb4ee7c3363ecf780549604c1fb0b811ee08109a1447a1b9938bd6368fbd71d22f
z39f3f00319df3904e9eb044c9b3542418475be7702681b6c257ce8165b16506c048c7f69badcf1
z34d4d4f56dc2747ad9a71add0b8cbed2c5ae27f50fb2570a8a761d1d6ff162977e3dd2226b2e5f
zb0e14c00bf3c640f82761b97ee53fdb3eb2463e71abb672d50190d866695ba57b9d4e5ca3972ab
z8106ac1faf5b41d6bfcfa05cb15e24cb71bc348db333c5d9cffeb7b4a119b4dcfab6037ef740c2
z82710f8f79d5e7841e5329c56716bcdf80f3ec86b8a65934b319f085b0bc28fba40120e2591fd5
zdea112a15a1479b5d1456907ebb67dc511adad18de02620f67a9dd373ef05b5613144c814968d0
z58d92fa901b0f812d588fd7d96c5b59cf741a956fafbee8d9828006b67a766b0a164796a8206d2
z80ad31e5b3ce6dffc5f430807f652b4c411ecb7e924d9366b281f686d63c05d2edb7ed1b2f3bcf
z968d9cacdf478a2dc493632985e808a4590fc8d867bf777ebe05350fad6abe8fa7224e47cbae32
z44d6358dc65609c67fe3e8b22ef7d3723578a59268ff8297e542b2733ff2ccd3d612e550afa407
z6b7edf9140ab303931f95a0175ec352f5270934c9d1234927414f5604b23648ce40fb5dd058dff
z5b5248ea5ee447479de76df7560e7104ee22d46e7737e4104dab2a657838f73e21fa4c29862a21
za49a0069427cb7da41227d74ed8ab6529de456514b562893ef7792e9c441f6463a4663aa06ae2b
z9426f31c7813e2c14bb29bd9f8de6ced43248086cb13ec35efc9234465d56ae2cbe3be07a6efd8
zdcd885feb2b702957c082b54105ba31c691462a44c7ba5be3fcdcc998f3938c2375122868e69c5
ze496fbaaa22858a5426eaa7a33f72dfb46fc93ec5ea70903580c1e3ae880a01bcf02f18bb95e19
zd84af93ad15e7e8fcc5197cb32396b752f5360b7d62b053a71fb552a067fb8cd740195edd4d293
zb9272f34451fa7bcbec5f01094cffea954eb03ea09dab73856fccb3dbfeeb2bd3a6dd11a440fd1
zd8c2e1ec4e24dcba6066fefd5c95533ba6ec204dab0434b8ad4c85e4aa5a1655cd970c8212697b
zb80314ea8c9e235369436903ac26b804c6bfe32038c320845dac5bb7a93750143bca21047364be
z2701c8bf2490e837079e0272ac1239edfff2e758fc19bf2addfee3ac5386bb5637fecc93cb45e6
zcb0f492df499f347b785a7cf9ad97abe654636063f11d56d367a7a277841de28c944a3248bc074
zcf009d3e58f12c98edb5bd9beb1448bd520cfc287cae8a2e332a870efaab74ced0e86e2d1bec90
zb1ab01c560168dfd484ebf3569d20e2eaea381a6e730b4f841c50b3ef72c1d56792f8cf5cb140f
zdd2ad7a5d5ecfbbf0c0e99425d42ddc2a3c8899d331c431d613f027f4420eaa1f5f7a9f297e536
zc24877b3f13ece812d116eea6c1493488506a3e299131c9fc10898f6682abdc1b0699ce6509d63
z2ffe576038d983ddc8a602955b410d07e8cfa94c92a4fd5eae9ff152c9878e1e3a5b1c42c785ff
z4ccaed2dbbe1dd197278f7b7cb32d1ea3667fd9b2ace6746bd45e5b3cded9da301340160f6c7fd
za64169d543e16c4e0be7e8c6c4b3550fb180b70e02eeaef63a2f3faedc1dc6d901b34c422d38e8
z4870585170ec399533b42777069a498b27a5360503df83fba2850e018c754988dd37736644a5d2
za3a4b021c26acfabf26a0e975683e9f59b631ba4bcc8ec94b865dc9b75121ea31f9e89dab22f80
z8645f94fe433ab447799f6fd99d4ef9ee4807e86a4c254a5b039ed938817c13c2c06212493f2da
z95bdf47a602fe1982ca18a28507edc4bbcd653ad6d393162f5784a68dd8514983396ae8860a9f5
z33e0a0a0f307e2252485665f8d300e255783bb0d41e077ff3a3f8094857a03d844e4a45b76d860
z0cb5a4fabd6562068ca6809515339ddb22c9e01086e228040f5d7eb4831f75204709e51eb64265
z6250bcdb2655e4c83a2140d4b647c3bd63e158dc7c96158879beebd33f3ada780e0e37d09b7a17
ze50e7b56e4d10a77090659117d92fceb3ef4b33a718a39743c889965c9b3f9dad20c8e1f084fee
zbb061dca868dfdef57cbac6884fb5a1eedaacb0048a311bc550ac011cf46dbbe32aef1581a380c
zafef6f08dc54418346b6dd117f5ef39d46f37285ee484d258544cf37128478ea2b36c93e09fd4c
z8ba21788017f9fe621d59433bb2bb13f2c53a6d08a015369ff1a360610dbed0463b8a09b8cdc8f
zbce919628d4cde9b43dcd02a7a7edf4675283618665244b4d5c354b6a5b553ac282277b78b4852
z1bf544da5ffacf8ae6d16f9551eb137c75a14369ed0f48d9486bfc8acb45524b6269695096a6b8
z1d6da8401cc8eafa35431456b26db7788327b0310da8362bdda8081e0d3394775a07c07691cae7
zf02f2640b6e7cf2c36316aeb9ecf8fb839285e46e074d0a3a85fb0fca19fc4c9c8ee567301ef92
z6a0cfd0fc5d26699cf85056d6fd0407aa9b350e3907fce78dfc6b0267415be24bfa0b887827fa7
zc38bba64f1d56d35ad5fdebdcf2e2b865237ca069f58e63df6b073e9ea81aa2c2677648c58fd5f
ze20124566208c6541db88ae67794c89bffa022294b38c0d4a1b07d7f03dec056c727d66f009c3d
zdcc13440b457043bda3978dacbf9c4ad4ae761a94cb08bc0a661096cda112ef856bd7a80a5d2a6
z0ab2f0a429aff1e83bbf2b564cb6c44322a381f7a44fc8d7a75620b72f8e7f4f40bf218f8bd562
zc29538c196f80dc6b2fabf30c499b1e169b997f61b6859b3c3127ce526c2bfc31a0d5af68e29f2
z7d3ab5929e64f78a9ce3aa5c7fa3bc758ca52ce1e5013054b5fa69b5e599bed9c58e4ce37cf8a4
zf782df0cabfa9c91728031d6dcca27de4b0ff916eb76bb6e1d26c2feddcf37b62054c05aafa788
zaab0756966beb8a93c8c7427ad901c57fef5a3f290fe699f7afc44537326106bbac6921afc1b50
zffa944b8fda304a2cdfc07cbc9c1426b41cf8515445906a11378fb73452a01a5438511f894b95c
z305778b076421c40eb55a96d3dc21ec4530c6d8d033f9674f124665f66cd77a2109fdfac7eb1fa
z3fb311ada16f30fbc6fff28ed6b8531efa201b41cd3642665854c1eb9e2ff205da8cd2e5a0c06d
z656cb7609c876b03683b9b43022a2fedcf98d78805b0a586ac5e3e05dbc95ab2e6f3dabc4af357
zfdd98cadcc90bc1e5b79849c2a2acffa2b3b20b879feb34a69acc1cf0203eca1b83753d9ba951c
z4cd235a3b5bf878bd663a7aa68c5e26d9cb834e50eb494db20d182b7fa58ac19c5dae9fd10d0b1
z7bef59ecf21f42e579252ddcaffc47a1aee3a87cb8ea495ecbc178a3642d44f9bcbc3cf698f54c
z4e9f486ec6b4095ec3cbf9ed5ee631a579a3114d2a7930af522628ef99a1eb6b12aa81b3b4604a
z6558c933d72b6b4d70f0b0adbc40ddb07ba930c168a84b847308964219eb1d136396114de7f413
zbc23c0806bdb6e02cbb6ef8adc327593f38080f1bdbb01e0b0ecca44d580294d2482a42dc72a6c
z8b21df2839876267a07d74b2f7fd9ce5dc6111a43943e969ea6edcc60f4a0c2edfb98418c16597
zae3b6b35ad95ce719853b7276674e59929fa1aaa416cd581276b68b5f850dedb6f86d50ffcfca9
zde2a8bafc8473d7b31219bf62f2a949c73b15564381036b3d2421e900622c07cec84a3a43718ce
zfa0e41100dc1d928e608564f530f496c95e60ee774a844805b8deb7cf81ffeee47b917a699b6cc
zbeb32ce6526a6ac643485889dfc1384b25abdc5fdc491440b45c3d1e773622a6b4bc9c64d3cd9a
zf453da8aed7f728197af54bec30753bcfafb03dfd2457663d9f8dba357d7ffc4e883f1619506f6
z5b1ab536bb1d71681256f09b9d064f924203344388e48007885fdf018b4e5b1272b83436d6c81f
zd69345caca22134de365b67140f45fc4eed93de812efa216a024e93086d320100100131f0e9900
zc59c9416c7996747dd79dd86ee53f325d0682667e891790c867a8579b50ca42b8fb6d94fb42b73
z6893127eb9b3074822683eeb88f29ae27299562cf8bc2bc2459ae05b28a0c5e077b1dcc9a32d0d
z8507ba9c1d024a68db4c49bac7a5342a7da457ab62af9bf794443a009d0f3c8410d34d9fdcbf2d
za67be6f18c3a3272688400f50eaf454e3e19d211b8a1ab9054fd8119046c9c108818e51eb55a2f
z4774de899e1dfcc3f28296850b121c17e0575f485df298d7beaff9b494b882c1bcd7cbb95e1154
z5cc8d0d37dc479e9649cba9e5f94697fb68533c4c79f4b5961d75fccea4a7b18332341bcf79d99
z39df273e2a875a20e5ae26c5191c2016ca8614961ea3bf2718f3551adbe251201da67765feffa3
z8ef64d24b66f6f3f31ea185bfad9e65672e2425911b349d533bca8c379de9212e3887056e71b74
z8bd569743d55938bdf114d200f397df4c270cbff34f38af321ace51b699c2cdaa4f9f49f541ae4
z8b46112facc65673c885818cdbe21de25ea5630abfe418ef320ccaf78b9c0a1c02fab8f5b0eb68
zd3b17dc45b035e0e7af3a4e861aecfcc26d1dc5f1909a225cc98e46967e1efe4633f75507c3722
zb85de2a775852b1800f05a02b1270db9abf1f949a58ed6b9c7b1e4a23c063f29f4589381ec3c19
z846b31e905ba0cfadae0bf926712eed728fb1bfb5124aee6dd529a1f241ab9bbbb727f3725fb66
zb8202450eb3a0139e9f162f164a39d7d96015953a5449096f0448e9d09cd1a179a170ad81bfe74
zebaf8b2cf10388b709e4d88723caaeef92e6279088f1c30205ca77ed1915f93d7b51f473d17eac
z1054886c4313a99df84019d7ad77b470678d775451a1a2ec306948afcccf54a401d611dfbcbb2b
zc39e859424941cd7d5cf4275fd263c4e64d567eedd4a94d07283bdbbd450caa7ced41b53dd217c
z7f4ca7eb8529b0e35dbb8b541778c2d2d1de6ff35e256c6bd120c8900c576d73662984d4f64c9b
ze3dfcc4e31893c950fa85fb9527677eff7bab686cbe4709864ef82d849d568ba1e7170a241a2eb
zb45085ebcce2afd084ff08be18c84ade1e3c9453019c8b623f931ef85c62cde33ffd611192c46a
z73faa22b6966c60e2e3db556e3eb45a62e7803565b7cdbc125231db1b48f5eb7b404eab3c489b4
z537b32dd292e5a24b593a7af9328a45f08df71f243fdbedf5d19aadcd5cc73091c53408e7de718
z98e627c456f4b0004605395a98946b9a991c7dc2f3a9d56424ae79ad7a8485718c3705c653f78d
zc86cca3d7a8b7df5bd9bbe81a8dbcadf250e2015fdf1c3d3514ba16be1dad6d079a0a15bc437c8
z53b6ab2db9b04231f446c7f2051f4feb4c35d1a9cc812c7966bda6570081d50de0f9885e55d41c
zc4accb0c64ec0c9650e15b1724a10c62db1ccc6d1c77ff40af0b07355676741b44430cfe3782d5
z19af9ca43055ab5ba7aff1dbf3fa9db15be7578e7d80821fc3fba4a6e31c9b26ddbe93eb986e79
z4d64d97fe5b7f16f102365a3e53719e19ee3332508d751ceb18fc6ec793cdc5df6707d153dd9e1
zb1a18bdd6bc2023965d656166f9228a0def4c9c0d7a82a3b65ea6b14f88336dac664957af24d59
zd62676b563f2e31e0324a4e565a248a6e2f6cebbf05788a221dedc62c81946ebb871403dd58689
zb02a6dd124804929492460ef7f92f271285d2adafcabab678c1d295d3f926c1bd462ab13151edd
zfa86113f585cfd370516e658d81c6797048be1369f3fcfad849fee2032fe571e3dce3d940ff30c
z0d350833c3276b99398e8cc895c32e524f8ed05368345af65d6d326eb1cc8b0e46a88fd7148698
z6b1fbc93b27876ff523bc46658ebd5cca5fd03ad3d502dd7359565a63c0d476b40837ea7b437d8
zb112445225a45dd2c6ff938b74f7e76d67a51ab394d863bba7142b4d7eb29c9d0777b0624c0a0f
zd00e29002ec3f45a3a37ec698a40022d9cd58d9c7cf72ce07975f38557b5aa5e479d76193c166a
z4fc0dd05b995a86533763c9f86bc7e3f33bcc419cddd71c02fd725ed56678045c2afd2f8c0431b
z10282dc7ae93337a637dc2604a628bce057570f1532c393a78060e67f9ff5f53fbf2542b184ace
z123dc9e973036268e552386199dae01d7eba3d8fe904446b2648a4c988ea554b62e5efa6b47777
z495253508bfdb6ba69b49d9ce983bad50a0725b992178be9b895945e1828cd2fb1d454bd0884ef
z8ae10802c042b4e98cef176a634411e1f30a52f182afc51f77088b70c94104c91895a959bd1163
z62d04e7633640925811e0b7f219d34122673e7d6b6964369852897590379120f38a9eff383ada0
zc38e0576d06b28f9107063c1374c5f7d335754377e7bc82a9ff474b90467122186d4bcbb99a5de
zaae04bb29ab7d2332bce08e7d8c27473936a01ae9b8944318f8a58d7b4ea8ff01de5a4df5e4099
zacdb4d18125a6db8cf2f502010caea708b269a5756dd2b0ac05e6d1551477715b9b986bb1cc2df
z25bf7644d04f019842e4062afe514fad450712742e29d9c79d2cf4f78a9412922c4904d9fe77c0
zc690ee330f19a6879ac1103f55270988bac2dcce7e3b57e8a99e7e0406d652819a2db505d6cb8f
z8a3135566a4f8e05efff84575361465019d570028ae3c042c294964c2e2fa7325ff2523928577d
z0eda66d088e2ced13a8b871c2ae71f838b022b56e38ba8372f148373b86cef7b65de58a8a7c633
zbfc75bc8198449443ee18eb4e14da34cec4d218e1236d3056edd9af1a05637d87b088c8ce15de9
z75f24f0a85cc8fd11b58567da9ab5531d63b290c538efbeed1bc5aa2d8ca5cbd92620c3c123f4e
zef69e72b77d8f5e8799cc09c58a20d4b8551f93eadda8d20dbb0485536351c0edee48f2983f06f
z28ccb18c2a64bb40a030880d816e6436c181ef6a238e309e9cb82e1dde0439968b872c30ad5339
z6a4b9fe36683653e256009cac493f671e75a28b3b021d7be6a3074a6084fcc01e06f0c5d928131
z22e4b44aec33d8cf057ac91bd7db92fba9a02df10798bc60797d206517b37919c3c429c47563f1
zbda727f30d88da4a4fb6535b12cf464d8e495ecd4c1997f06611ec998f6a74b27cde3479592efd
z1d5df087c9836bf124cad8338fafc26d6d7517298d1a31a2cf36c3f6208a4ff93846851ea46ad6
z0ebaff453fec0e5e89df719afec56052351384a18fe3fc057ba062d183d3fb07460d1b3dba8fc9
zee72133d71a5c22866d5b87ff170dfe208853c3834e25b4630ae5a65b246a36dcf652438c2664f
z53581c47ba4233887ef2a65c3d6df2e86ac4bbecfd4829b086dabf19c1a4c19f666eddc9e1922f
z97c0a7010c2faac456c85795398617728dd33337083cf7b52efd986003b437a264fb6df76565a5
z7631b2f4c2116d32d17b439dbf7d7df9ada20040db90d2dfddcab18b3f2f6e2cbf68ae81a3cd3c
za5d843f49d4d0765e966b3fb78d84f4433f410cbe3adeb470cdf5509ef502202f358b10bf1086e
z9b5599670c565b9217e9ed352e68cbee7726660f52bd5c6528a5f0e90a3a9aa138321cb11c146b
zdc9dc09ed0bde538c9a862ad61ef667ec1dad46af85297b146f2e76f41e18311331499e3486b6c
z9d78a6ea32ad8bd9c376be79e538f77e861f8a63bfd50eb900e57e7aead984c2a2684d20ef0e12
zdeb7a3c49655406f20cc18315a9d634688c4b32c51b436920382f24a7a87bf1cbc90e25396406a
z05d731af6f03bb030ab248fa2c06947ee8d8eeba8b0282a1ec6dd54fcc03fd2c45a63e5c4e6bce
zf4144571aba413aa1d53c1b71b766aa7f69143e292d8f4061d58cb9391533683959e1c0eed7ffb
z40f8866f17289ada0d07e7522ec03e002c1ca44a490a8df7fe11ae04cc61cd032cccb0a07fd911
zbc44e27ee5764d6c7db65ba8ca60f3a7581970c19f6c46ce0911dae1d68aa6271c3d3fc9a6d594
z947751a686c72a3aaf80ad8315b265873a3e724b933c7eb86ee4c532f1d065ea969434aa396483
z685b300aa8ad68d1b795818e1f0bc1b705b936484d7740f79133d6d3aaa6e7dcfdc0d2a36bfde0
zfed3f5190f868ef1d4b4e683ab504cfad12efb45ca790271407a4bb722c4507df062fd48d6d956
zd1e4bc6772f14b57c056d5186053883aad70505529135265eaed0695ee66c46c04abe13ee9c2d2
z1016a337ccb82d200d8a74ac178a234f96523c553161b5b117e16328c91134d19071046dac43a5
z0db60690bc4ee9e125feede412fb09d40b92804d366c98ab6e82f8fe182498ce30f57725a2043d
ze10e6e1c83cdf8b3c78fc3b1ebea90cf272f3682880edfc3f9ec4933277544261f16c17c2724c3
za09f233fc4091025f7126ab486eaa8d4f1698670644e2adeb0cfc0638dbec4befd95f2e4c86397
ze9a6c5abe6332a297e5049e734b805076cbf68d40b73befb54daafd43294d694189e8238c97e6b
z16b58aee5e5ab11c204f6bfd36527a0be8e6b5b880d9c7cb8ae094412cd213de8e35cac47fe266
z92c544ed61e21846a02ff6b921b260eeb454660818407654109136c9abd686516ed6bc0fdebff2
z5315fccd2e56297403ff0ae6c739c176970adedd646e2b7df56ed1c4d83a0091524f4e5852bda2
z6cfb6bc5c7f26b5a2d854129ee24f144093041b623fd334c78b1a43cb4bc0b1b21eeb55f2ca189
z7611657f8575de32171ea883d14f5e848ec4d5ddca4a0fee67d0eb8488660aa976b0f8eb605349
z3612b02e2ff8b535466c7d25363ba4aa20c46d9af2571bc251d719428266ab77d59aa2af02a9b4
z13fa873d09753f051091b65b95fde73552de350e54a59dd77f7290bfbf5f4046a1c2bf56c41d11
zc4d27228232e7a760e8530af6998479900c365264f91e1adf4164d55069d209c6c7f1364a60014
z304baeede9ab9ec434c2573b096ce93ca099577741273e89a601aadf80f7fcad7b97d6b41c64c0
zbaa70af42625a5e820308f30b9b432d31a1c6a6a527284f41dbb6218c2f787c751fdb12d590892
z0b1f921fbc18c26a2d606aea2222f6efd900e5250c340dc619544b9df95994c86c7c5ab99b1ffc
zd72c4cf389f732720e5a155e8c84cbb52df9f51f045622dce01b8c06e86154ba50731d3f1e0103
z99b58b180b263ec39a37447f119662750f2aa3d9ad7efb5e1a49630f186cec07d5bbd68cbf1c27
z9fd9e109bb9f7c000aa082eaec0dd6bb323335f1788fc059c3208c981bfe70dbac2282de644d52
z901e473d93b68e62fcb54aa2611ef912ffc004c84e8381a474626d5c29a2fbfd6060b6fc35b3aa
za674ca15ec9da4a6257189e276b37a51597992bd4d5e96c85dcb8ec68cc063e231530e0b3ea18c
z7c4a7c26263d4b99eec6d7f6b36cf97e92995e44d4f32022fa104b26773de287f26d06d9d8a060
z264e135ae7e62c596e3af360daef3b92cb324010eff2ecae37bd7463b8c122a77d615ede18eb2c
z2e8df11479a8a2a12e019c92afd75e18062cf8d1f548bc28eddf447940c5686c4b74a7ec05af03
z9f71b2f6404f603c78f47ccb9a01ec7dc947c91474e7886d38f25ddb4aa31c649a5d7c8d10d6c3
z7d8160d2100a47dc477d01cb28c16802f0ab8ef3dfbb4e22f0c94e333293d19ee65d2b36d00416
z2d7dcfdb3651f1895766402e0def238ec340ec124cb15ce1a6d8e39b1e172fc193132aec7cd7f8
zc2d0e18aa9a9ad90f2408adc79bd1de2053aa27e9356b7c8662d23eddd1045dfecc00619ea44cd
ze7e21d74292367651e6777c1c8c3d0f967d75d4066b9fb01b2a35403c0a418d6787c67ef766a80
z6603c18f1409f441e583bab55b08cc062c3fd96fda977b9a86a56f0a88b44ad1c1d9fa6643e08e
zbb82467cd86e2739130a0de19497feb3e51897dcf9c502a7237d94c1b12bb3d285b9be7885939a
z63636851117718cfe916d067963beddb5a4d96e5bb8ebf87a0ed30d0102acbe11a6120a847c4aa
z9e7d7134632d29007fdb9d51bc2fb94df1bdcbe29e6f4b483d7e19dd9671612723f82ac9608b1e
z74cd83b4e6d17dc033352cc4e82066274c2ee96032f5668198018e32a1aa68383a1502576f4079
z25ce7243032f3770654e357779b6de2b0fd8daa3e17e8f66c5cb4f86087f64b653aec3c68b5601
zcc304ee712710d7c7a1202619ece506e3afbd21e392cbcb755b9d832de29210b89218f4f947a9f
z47eb40a4d6110b5843f74ee46604c7061fd7246e57fc1085492f1cc801cfcdd9fe374e30c5c801
zee9f2f2a412e754fe7e9b562fe5835059d19e7e6e87224142f77e60168fb643341c787c848e4a7
za02fd7c5ee6d0a39a5b1b747b046edc89f0af540bec56a0ff42bd37f7ce98c1cc91871357abb18
z87acc79eef48580b4d3c47046cb911e008b3bda35ed379203ef4d9dfeb3e0df2c61babd6ab61df
z9b8ccd6cadf1c295a822767283315736897b4d736319ca07050f1cfd1fc5a7e7779f0b1589bacd
z6cc6530558cc2ccdebf3aff9f1ff880ff89ce44cb2cb626c692d88c7e50155ac92b46042779dba
zb9bc0c087c66fcbc33bd3fbf9d86443d6b7cae714a3ae7dee77111e8c510459e985e0953341dff
za53ca67201e96f08ebdd5343c99f541691b740a8bb7f3dbee98c8f6c7f63d7c9ccb8800904e1e2
z5cebea146f59bdf7829b23bbf2a5b5ca3b5f5b70fb333c3c71f4351f961e866929af8b35a8108d
ze6fc900911aa373d6fde24a58804a459f611b69df8da196fd84e24b228ca64272be6d9f93bc49e
zfeb79093201054e82956d241bd58bf5de0d83fb1e837e14ad10b06a30dae73827bb7309d5fe392
zc6b27256be46a90faad9bfad68b536a1b034d45899fd2733f780ef76b8d6819816f2f0a620c89a
z9ef303094c8917296d7265357e90302fb61431a1dbe5b2af6b8448e21107dec5e43adb0ed8cf10
zf5318e14a176a78dc8b82956dae3d51915c1f4e26a8a0fa71f477950adf2b4062fa160aafa8570
z550731c9ae2e255a598f6967ab6f117d977d87defb075f4984e009e39d58e44e960cc11ea45301
z42f83d9e3fa37134a37560b53b7526a40cc2b30ed72fb4d4e2d9eed877d7a66a7a68a8a7e16a8b
z83c03cee0cc632de7f66f49e3ecd4f4c9f550e10e2b790b0d27e774fb6fdba05058c5d670b95a9
z3693d0c75d5d1817eca29df24fec8c8303413628ad869890c10a8aae5162772d3d9b39c4da3383
zb01cf0330d804dc77bd60409fb8ac21278d6196a690d4e121ab28b75656133580a157327a01a4e
z48dea2552caf17efd2ac21306d2bb0989f9e9a4b0db2d43acaba3b5c80b0b6bfe8cdb1615a6dc9
zd31cbf218c0a651bbba914c2cfd960800a70c13840ca552bbe1de5c0ae00bcf7667c3040155a33
za5b98f0c670d8e438fd2c1d397f9d06ce93ea0cf2eb5b45af93cffaa25c27eec2d2c55396f833e
z63847cc0d3866567d94a6cddab920f62535f3776ed9aab3d0c4a0c5b94d31c832c20775244765f
z3a8b8c2ce433841280b76fa7bf6cb011afb16789190eec20aeb22b2e6df47c21076ffbbad96997
z31e9915d7a307a5b31355b9a9ba99663f7865246ed1415b54a2891ed39e886d88345fbbd215e99
z74ed15ff91eb9a26ec2791aae1c34a7d3925924eecad0a0bd2bb99c5305f1b9f917478d5dc814f
zd53a505dd003095b1a979d3ceccd9d309f9306c105604ec2ef8f8e7bdf809aedae1227b70e1784
z2dd1f433c585c93de627de7871d119ac302016eaa17a42bd4f0918b193aa10dda1f9eed986ea52
z711a7db4facd5d69698fa4a427637a9dfdcac87a36e234a93a5ee444ecc9b4b56c73d536ba0a55
z2ceb09ff7d2330297b44231afc422b64f4182ea06fa6ec72fc7896ad64c2a31f4418d72ffb6d59
zdcac278194b2122603793bc4abb6196c9be180a8ef54a41847f61273ef748d46153ef3f32094d0
zad0c08ae640269178b46119e0a9a8016db039db2e7e61a3121a457dcc9a1c117619f95eb632ce8
z734fa748069105dbf19f86943c6d2e5f8a79cd4e4d39e2bd0ae05f45d9e5f9f990b47e8027c38d
zbe4e5986fa820f9edfecf9baf806aa2f73b99497dd98dcacf25ae15d8efabb2b6fd64c939557e8
z06e12b72ce5d5efc8cda4298c5934fd0f270e378b107000e848a57066669d89f8b9741497dd7c8
ze64e8e25b3b1acef3f8b7d27270ebab9e88453851d174d061c35d7d7271fd912e4346bc06b0643
z2677eb8549cb4cb16dba3b1fbc737e5b790a2070536964d64dd4a6361f7f424a9f8a5f358cb1e3
z4e0452a6dfe3f7c17762e13debaa1de729223990d23dfb675e39e7b034c9932015013d696fd434
z2af9bd39a638ccf8bc30107a31902071a1b04efc5bf0ad9229539b063736111c77a88c03668ecc
z6d7a89b78aabb8f38a9d6c24e6201a2885b1dd16fcf4b63ee5586e1051eec7cb020afa2778345e
zaf645516bf24c4c9a463d898504f0668db196c6c3015fe17472c049fbe71330aaad14c553a05c0
zec0d77fbe9bb722c0d70b518e409898a7f8ca26c9a952810466f456a463ca8fbda0c69bce1ce26
z421d854e565e97596a9f40a82f7164db2deaee527350567466e00d60bee04e258056ab95805ff4
z88005f50f4369f9e6254317346b2353a0cedb543a928bb070c2d5faa8ccc15e61b0dd5623ea34a
z49c1c752129d0bd73f3374aaaf6be84291a4dc1feabe311a79d6407d86438771520465e1c62376
z316297c339826dd6c37d9bc7e6c89efd115b8d24a16a740980c289c05c4d56208990acc2739ddf
z043b3109b28cb834e49fe913cd54ff1a364dfb0fcacd9262b7f1c65c25845ea247e7b54fe4bb88
z1cdeb19732b3ff1a5e3210af5315c5ba8d16696a198c651a13b8b7d3d43717aab42ba8e6b51769
z65a5ba82167d669ff29e52b7d43af05dea8ef6a9fa01776e00c961dcfeefbfadca44b56a9ec151
z7d1f636047d6756554881c411211d9f0a8e2f7857c28efd9486ecca793323525962dad70721506
zf180a0347a4035a65ed300be5cb991b582ddec58767df068630a58754dc98531792f604ffdec5e
ze8261d05283cc4f6fac01a7cacb77d2468c6ea6eecbf7362562a13b8c9f1e1ac3e01a8a56865dd
z523b403896c0c30ce89c5a7c613144e7c7252a5b7c1854cb7b4947a6aa0c8eb91af74a3465f12b
z95ea25fff3dc68a4395650a629a321a1774d8b1b1f4ec9839f7682d7179931190d0edfb44b94d2
z25e3b02de1f98a1dea10fd7ee46619cb7437f412fd6be8ed1d016a9329bffe3a569af86dbcfce5
z9a886b1d8430a4fe89c3b65eae84cc398797c1a6497e0cfa7a4ef6d2e6afb706008cfe0300daeb
z601c23749662f9a122adb4f1759e4d0ca342b8e162cff54e69e232e0d6cdf704e56662573a4545
z198200fc2bf78953e699366fb5690f599fd0e4f719e44023e74c0ff10a51e180b381db082fbc20
z38e549857729cea0868ae37b999492f40972864a86241878d2b9ce8d50e74c5e0e2138cc7a1da7
zbaabe8420db10415cb9648f0ce830fbb128440a3f1df8a8521ea4f19c7f17f4a4f0af985922e56
zfb6400224b78754189d279d2465b815f5b0f5190ba3bc3f6cb5eb3bb163d0243c6b8f61c22f900
z382a7390c26a960f0b2cf90cc77393b0e01950147d5d779ec432f2fbadc3c0547da21007bdcfda
z112de44b728db75f6e9b842a6af2c96f4ce844709b07860ea7f18a6278a7e7513e440b94635f32
z9721839f6da0ac1a58f307fad28c38fd9677ad72d67dba27a354f9385b69af2816a4fc61b6d9df
zc213822b5ad219b8b7dc481c99ff5b505c2e672fd943933600435e5335932440abad546aaee17b
zd2996fed7f79ccb9568f026c0f0cae4368d48ebb9a35abddd89084996064fd9cf3f09230bb16c9
zd1ea3708677433154a3db9d59987626aeaedb9e26d1d74015b7dc63bca5b8c38c36376f70d9fd2
z72ad27d0ffd19fcaf62a3476c50f5dfe65c52a06eeeb0e359c4d084b42dba785e6c11d71f4c6a2
zb6e4628b2056543ac57b5f5cc4133197f7bd33130b665fe9580044fdfabd203894224b1da0b7b0
z4df25937ec201ffe4e65721f6f15e088164724d842f6f12743aecdbd7b6c4076c572329811a345
z8df03857a335e94c6c7128471310b0cfd5521ce2fd8dfa73925080a21cfc57ee359610e3370c56
zf85eb708d832afc5fea8775c11b8365adaf120dfeb33d30416536e9d79bfe541272a3c84e08c83
z0a893875549ef87825836757ad82e0b5a0479862221718e0bbf4615d451c67d5b0b7d3270ea7e8
z4655b32ca3042d68838b138d24f32e9e8ff35d14f4160df4ab008fb0a21e048016519a1b6dadf4
zf8e8650d37a665d9c0ff650e81dc7ae27f6d7f7082d810fbb2260a30ebe65688f0390884015c55
z8c34aeac6cf9586b4ef5c9b6890e4743c0b63c2525bf28c09ebd6e8011c9a3f000a27d415dd6cc
z95fc589fddbf6ad0464b8547f0b49c49ed4b8613d528dca943cfe62c0a05fe5bb76b3379b71a74
z68211599f72c21f5087a703aeb0fa729922af3ae464bc49adcfa7fb478a851beb34920350b054b
z801a17fd33e47002ceeb8e5b9165bc8f4e1df9d3d52dec52981296d43a023b267b4a080763e8b0
zf9563b0ea322bae18ba9ef60dc61c2ca50e1214e2bade6139c6fa0b976dff0b574c7049699825f
z44d2798d3e7df2d3278b48c60e0065e4ffce5a97a6ce16d70bddeac27ead763b6dfc72f13fc969
z2e69068fb0576073c7900bac98b0119f482f762dd14d7e18ff75f75d8fd56a9b11e1ddbcc833a1
zaac0599dac25e0ac1bf3bde8376a777e717ef0dd1d3db9e85a4e31ec6a10745b5e8bfc1c5ef7e0
z9c43edcef2437c6a8ada48c7975a8e46625b284361c5f06f54c03eb7bcfc7928d7061a514c411d
za47f0e7d9264eb811048b1cba62026d51f6710f1713d7e1592da4d3151980da91d77ae8e6efecf
z1ccc90e263830de0d365166013902b5140df0c1191bfe64ef3b2fb6a5af7f70e72909be4029f14
z6a33be801403a6c5ea859822bffb4071d1e295c3fab47831b83b76b24c942bfb9ca6a1d7151e74
z762c637b4a60b100782f65bdb701d1ed25d8f3342717cc3fa464b0f5a08771a3fa6474fd3f6c8d
z5560349170d8a449f32f7718f99b7c4253aaa94a96bfee51396ca12d2265d5fd4e98b9af20135b
z8ebbe7ee9aeebb912bd713cd3c265324998f43c9f57485e6ebab353701511fd00f4d481fe72403
z628096129a06fd101bc03bf8b78537f200f340a66f8e672bae5876cdde4fff2ecda9525dbe1cff
z35207d33dd8eb39978af46fb1f61b686e12f3d6991995bf7fa5a6a5c9f0958ce5a1bcdc024863a
zeea96ac763f8115988e3c5aa4dc2ab9984cd13efe9c477aaa2849dd3c3ac7c726b73af31c2279f
zb1450eb22a00b3667ce64810e5d38ba3a9888af9f5da6ba358e3de676b5a74bca8d67233f31f88
zfe7d9c1f97792b336869660c47c167fd07b74fd6171549c15c3df5517effd94b23fc05fb71f89e
z5f0cf66883cef69ada0e16ef8910249f7c6b6abffd2b2f6d79efa3d0e53288750fd560bed4b8ae
z6ca5489291824b3e95e6716edacf1465da01f9564b35944b1405be78b8d6207792843f5cc47618
z2246bbf671bdeda1e08820bff737eabb306ca6bf88fb11189ac8aa19fe84de6277a591d7dd5a0c
zce9a4c1ad35b4c33e3856f4e230d28c35db62e82a05dde54320442d72f84c25fdd662f35f8c9a4
ze5e859852e622c88db6bdde8a7117857f66fd23fbdd4ed66e72d0d73704c0f83ff8219e40713f2
z782e719d22440f1042757cf8b33bc12cc2cb290db7d9ed8f91c34c2bc6b1f2b6cd09c5c1ffb976
zb94f71777a5e2d4f0e8bc2e9f89baf98db3609241f955513a601b63e82eb1e33881a892f7abcdf
zb692c516096b706b7751d329b3ff9fe2305aa27ea02cbe7f0c9a8267de1cf7435aed079d993619
z552e79faebc6eb10afba8b665dade24dc498f3a43d02cf69295abc178bf6dba9a461eec5246019
z3d89eec9a7e51e2502602d7971bb2ca1bd505698c0aba0128588550e4935185a198f4d67ccf328
z4b779d9082f3560af6b3861c0abfd710f307fed02e6373b8049949458d3a1981dda34c2d678488
zdb38ac8518ca49137fe838a53abeb603ae09018f2a8f4d371d6f0814ccb51e3555c4812c1b9a2e
zd95c5bf837176c4c2268d9c70b470da5793b7799f9d85b3abb8e4d33573e7d7cbec0f7200a9c55
z242a0792cabcb51dbf081d5ee24b83905f7b818dda739837e5efb332b67e0d3bae1790d6339f29
z3cedc36e4641c3d66f14d26ae4078f8285c64d8ed2173fa6781a27c80ba0ffd9e637eebf0e0e7b
z2f653fc078958288f717bc472457f569c4c79b23ff73b4454c51276df4a56b13dd62884be91a67
zd8f74fae48e5070460c8004eb64b733b96ffd9566dcb1370928af89814c2c4c34f1717ff4bd734
z7c1de7568d8d3969dd32986195142476fa20e9b25d07e15670b037893b4220fff6271d4bcc2d1f
zf6811a62611e5eb3fdad73299892f7e75265d09e2b90c0a571a9bcce7ae5e71deb7a375d79d8a3
z0a6c96bfdf466cf0f125b7cc3a4bb99c15a6a6db7c7dbd0e088cf586fd97f3ed64ae57771a8a6d
z5894f475cf9130c1f2188a41dd5f35921cd71205609dab41ae59f8c56fd92a4c22e5805efda38f
z37da2056251566b8a1467a47b63bfd881e1cb9b7e81a046a8dccadaeef933a810c39f0c010913c
zc4d34edf7b97a59f2cdee8bc842ad2a859d6ffc01f504b0bf64d117bfb463061226808e9b3a5b7
z8bb544cd56f4b9ce4de96d1e6cbf2183b4d208e25481923a60bc12965ed50887b2ddd61c13aa8c
z1e3a9a6857824f94154d70aaf906850ac55a68a15dfffbbd1cf7118cdde771be67ccc89917b4d6
z00656664923051cb2e872b78cdee192f880f894dee62e5f6c84927a3912cde88b5b099c1939157
zb3e4078dd1e272e601bdc5c3b7ebfdfacda0172eb3761c5ce422fc9d5720ac6a616c60472d83c6
zda86010c6b32ecdc6ed68421182f94d604c47fc1ec14ce522aef8809bee0caa9b2c4bb5b144cfc
z65dc087c8c06176d4220cbe99e920c0fd120a844a281a75963c13e5c301ea104745509863e7e0b
zcf506b458e47a89fe9e4ff5bfb2d6028419e087897e23c2251f228f9f29dda5448b4e41750d7b4
zc6e9d4f740461c17a2a59a518da434a3e289c072455f257ba8bb35db2011c8359681ad2f6814bb
zeb4ffff29d7c5ab47078c989fa72228b2554103f930dfb3c52c26bc9c236e01a7e93169471077b
z71e9a1be913441579ad3d15751da75dca8774387cf08ec6fbdac624a96684c495e99ef08fa6e38
z84baf489687a1bd7b59a535d5c81d027ee662aa51c84a912de4b9bec47f6ed0548b328df7b7a06
z61ae8914c8cb9bab636cb88402e7e3bcfb1db54fd9a2517c47a22de18689ed6de416d50954182f
z62d0c93b7f27658a842c05650aae11d1adec527361b10a529a6b7a0a63d511e02ef54e63ea833e
z227e631f0e76ad48822208a0247c4a54fa7e94e9386e9d4216ed26292dd728017ef8537797ecab
zecc529613a068fbb059915609dd1560fd33c8a11819a64b86851d7dd4fa22b8dfe6acd9affd00c
z19c0e5dcff0e808ca6b65fd4964db814c4e0ec6575d119b086671f4e1ade0d841448d56f948d48
z6d0a7f30c81c5030d2bb6e2b4efa5e68a6d8d9ef6f8e6266582fbc3ff51434361db32dac82e6ce
z83315001377f252838b72d6f0a67f17dca91dc3d9c6fa0ecf19024a5d147bf041ee5c9a3d55677
zd8eee46cd01fd3c2f431bebeb67e4900c78840e06ca9c626fa3a90214f604af2f3cbfe9cbd8205
za566841d1d8e93f81852da5270e06c113b6c1ab718f562882e2a6948fcc835d9897ad689612110
zf149a04406a5ee7a5a4a58a2176a9526d49241a56c2045a2acaa851de5371bcd26298c6ab36e4b
za0470a8d56526416519bf2f60639e9b83d2c8d7a8a15fdc771e8e9e96205d5345cbc65ccd3af3c
z368bcb60d2aace646e3df535f29d6a4d33790590c0566d6c7754597f5de23a5753e951c873aa1b
z695ed222760ae183e25a01d3ecfc6aaf597ae65e3d7c20b49e72e131a8e3ea33dd504db92094e8
z02e5cc749fed49c50ae24a585f66e72ef0fd96ea6821fba76fc20323c92c8e10d7dbb009c613a4
z6c7eeb512aed5978de8e4d465c446a9d45ef4b5c5b2ce1c8ab6748012d5e045369ae2e1c42e33e
z5dee951b83c56df606c60ef423d44c71a51c48cf6e0dc9aac7102dde87091d2bdff541b879453a
z8d6b238d6c50fe82b609b0c6f7e097b46a7f82ab23a152db5937c3c072e8142d8a8f1a708984c1
z767adc4c514c631d32de342e4a39b52074a75acb28e1d7e8ed8bbca6ffa9b52ca9b14df11a203e
zc73ad4ac6a9668d152cd95a66fda78f9b0f37264bf0b99390e8d7429800825fb6b124d1561051a
z84d499719b062cc3ced412ea4cc194e9f6b656acbc6ecaa39425752efcc38bc5e5a5eb887acb76
zf83eb196b725fd09eb8787d6bf893ecd8171385391c245f562b2625644715153468567101e9f68
z186d08bb204dc8425047b9a57469a59c68d830a206e3533785c03b7f1e52a068a35f39b6e1c654
z99be2b3f9a083fbc95565b0416d486db5e925f56b1796951e6a9db6df5cfa82bc8123444b6a08a
z73781ac159fa82582892809833c513bb1af02d820dfe6ccaa26b3851f867aa152228efcedb3b21
z930dbd51f1a24fdf1f9fbb6076d6155f26bf6692521d5b164421bf76202075675adc1823d44dc2
z4f1a6409c1ca5cfc51d186a224ef4dd706bd6c0a3a4de9ef65fea7b61f98e2dfe7f140fb9bf484
z223fe898c8c15fdd33dfd9f1b7f4ea20b72df58ae77addb53f8e07026e7de4f6d55f5346a51caa
z8920302a73669b6b77319d48cb37e30b5c6ecae12170aac91add0d2b77ee85dda69dd85850c71b
z6635ac4c035dcfabea97945e82104c28733612943abd590b20f1aac89e88d2018b4d2d912b0389
za3e6a80170e6da12aefdc036693d1e78a32b6e0984bed8bdf618aa8c92bc4ab8ecf12a6c8ecd3a
zc224173a4b4896c90e10e1a7ea582a2c9c1eafd3c711d22d100b2135af29bb1abc27fe6469ccbc
z9f06188dea97cb5a04c7cf56dd45fb9f53d2bf2dcacf2ca434ef9707b71307e9093043f77e1ab1
z3592fc348b8f7c3ca6e0d03531570b6158dbee45fdcb26aaca106c5bacdf8a48dcb220c75325fd
zbbe982fb0d272a5fa6c0ea5713fdd2f8996df08df29e976d693a0c5937c34c26d5b12f50e5620a
z224781013011bd3747a46f8d438977bfa6058b128f1ff26cd765b0bddcf5496e2c6aa56df148b5
z1417365d89dfb678d3ce4f1a7a35841de422c5e000a1a79dd1a218a48bae21e90d9e67d2542588
z8ea94a63ab96739f69c6756834bca30a27ad7538d40aaec165d1fe6c421e3dbfb263279b8ed619
z251b57c9845db956c68d91ee0d8bce72fdd34df9f7d09167ca531864cf2702a686afe97ae94cc1
za23dac49c2dc33c894f778bc9f3b51d4c2f3ec3de0c042e96545de07cff7d213832d9c18ac3504
z0fda50218c19b20601c64ed06c811b973f1e54ba2f07612cde854cb1b1afbd448df77425bc4cb0
z00b6a0dd7ef4155c9c4604a103ad8577aa206f03614001b412d0d816cd9815198bf968ee85d3c3
z1d08515b765759baffc7cfeae106134f24783e5f972edf62cde9d18a451179bc66746577700c12
zb7907db9c91361e2448670b13009aa722034faa75629627a9b2f1337b4f5724cb483e122be6363
za4a599ae25f3b19c4e6817e7713428aba38bb4e7aaf5b995b7d5ef07fa7fa901dce5968246461b
zb643c73cdd79985b4daa5d4682d0f7f1d38f0d894b4ba4d17675298ac595f3d861303442aee885
zdc7580494fd6391d01630141bb84ab5f7acf0091894f19b1a73b79061158a734fd53b2892225a6
z07be3e4a9dfc256604b405dadf6391e7dae5d4b0e39759e0260118c2d1608a1eaff9577c11a499
z3be3363cf754293c1fead7d9f246a1a3dad94d448ff171f185b9ba2653330641f57eb665ef1d8b
zc49c4fe19fb498f3d09c4ccbc6f49fe158d5b31995fb802a01ec5df6fe792b2d083a9b5e6437e8
z8732362feccf3a4baaebd177b002063c8d3325c3852965cdf5d15c4472ece0aa5a3dc5af0566ea
z71df26c8a5eabd63f536b206dd2063453485e9fad598c2b0dbaeb97b5b61d98eb94d1c60d36ff0
zb2881c5b0da2e65248c61cce02a0dd6953242428daf8520a02b9e19ac1c60cb1a2abf0e4465c73
z2b75838e7cf643831b92c7fcea0cc9f8280b100f4ea662a0b11566667fcc81534c29caa5d9554c
z23f7fb0aaca7597abd582629df69b839dd1a68779cbba87508235ddbb71bb89bece2589535661e
zb95a96e1a5ea32d8e5ad09f3877e6ce87c1e19ead2bcca0a317e96c6edc8c250a24c1bd47c4011
z8baf46ed3768107989c67cf147dac7442faef46f5e74597085beae1cd4da438e4d60dfc0eb3716
zebc4c8bc3543f310610e596f01d2afc8e6a27e1446452013e44fe32490218a4abc92a2e6f54c36
zc9e8e4b3618d502148a098467a3cdf19e8cb97a777d68b555fbb478375f3ba9262d8bc315a3f78
z779bbafc6dd37b4768d68ff7239f6a4bcd2f03a9c6285e2a6bb45329e216f55d40febddd6f94fe
zea1ecc41b89b4910f0bec92d571e66cfee06db9631d15d0e1dc84d4fce0cfb175317948a64160f
z39111de44f2e04a991f324a85bda1bdc6adb07174a9d8339637547e895a8ad50f0f4f2f464b6ac
z7e79b4ef53c9ab4b21a06aee89eeab700552c3412b1c859bf391b09b8f8c999bbce4291d1474fd
z443a49f54c04e6a6c95f102ff340b5af18c91b557fba52c2afe7a7444019b410607608a9f9859c
z96974b2b86fd71fa7eb25e0b1c73df60853286693e1ac0b906820c88bfd3a30fce4b95efdcc8eb
z9de49ab899088e738b9a8893065300c31b53eb23b989c99a4e4bec307fc303021b9129d15dc397
zdda6fb953dce20627fba800e0ba19cacc957c17884a8dbd843267f594203bdb2f050d0f46f2cde
zea31382b55e7ef05e62eaea9632b8b08c24b93bc6932f6d932e94ab810ea5189a75c753e7890f0
z4679681df463d020cfbbcbd208dffa7b8834f421fa308c690207d3fdb0c6299b2c70a18784126c
zb1cd201d9771a317449ab4542bc6a35bc6cef483564bb7f6cee735198e92cd03286bd7238b42a7
za13ce331e2c841467e8ce41e3ee79bc9eb441482be4025cef6148dbe0247524eeb033ef2bdae0c
z1633d02203a894c777d73e5e2edf12d0d6396d182c11ea7c6ad612812a335a36553122a0baf4a3
za267bfd352039f7a575bb016d81e0ed72d9ada53635c50d7aaa0c5b6361a901c341d2256b16d7b
zae7dab7f2ebd32b3ac4f5d71eef319a6d534f530e2e1e9d8395e1543b98f3e0f1d186fe1def26c
z7264316892da8b7fbd7891dd77213ad81f734dbf0f7ff2cf6c82df0dbf46c06b39b23c76681afd
z45f13ba9582e1dbc76882e4fedd02e48aee755ecffb7ed3f832431319e4b3a31a3e18d0e02a520
zbf3a8c908e660290fbd20e3a8d26ed99a9896d84037b120c12148c4d28bf2a15424309d5b9ec76
z5b11e4e878c6a7536f7bb32504babc0cc38aa8200173b0001dff9da86e8828aaed60d6545c3cfe
zdab534f1967a41e7469a0eb6ab970bd6a9bed6efc4ca7b509d6e454d61748af7a866aa523f3add
z3380ca38aef072dc1fe133e3809a7c9b56584c4a148ed8e40be4461b2e3840b8de30eab58aedba
z316e5f4f9c3cae9bbaf2cf751ac6b2f1da43e4be62516a884a1f735da52ef623fe8ea9aeef7eb6
z25b025591ea2f2dee8a23692107a96b07859c5be9857c080bc03cda4c6cc3a4b2767e4dc57c031
z3c04644a56e944d59d75973fbae86616fd50e8e5d58b61b5dcfc41ad5a6448a122f081d8c79ef7
z4287bf6783998844b35e2f430f048062966a1030d2b01e83bc8d00d72b97dbecae0a868f8f3e0f
z4deedbe2fb73302ebe4cbbc84555f35fa9b3f7b973b13a561495eff77aa18efc557415b47b6d6e
z6bc12049aea26cf8e238602ad88c8787696ebe384cabe8f27fdd0f0e65492c5c6b4d6bbba01293
z673104cae50245b3008de59f8436c3652cab527fd2e19b9b4c7e57abfc702318f918599465a831
zf2ebb69d0b4a9584ffb72047213f99bba0b72bfce669a76cd758d08e4a0fce7864586412e677ab
z25f286aa01ad2ea58c8cc8f81ecb1a7aaf3edf860aa932d3d00971efb3fa88756d1dc6e0fe273b
z5876373827476e3b4a089ab94d73045534ba83e3270cb1c35476751b7259fbbb04e06c64dabae0
zafeda603f5c8b5cf7917191b9082f574d4033069add0f8a9ad519c3367b7a9fbcefb0d76c0f6c6
zb8935d54b13235c9d833059897ef5cb16730c337740eb6218c18e4e841563ef2b5f9a9ca538509
zdfb195fa73ebb07edc4193f837507a50531f559797e221bf83f204899bb25e2b17637488ea3f69
za477071bb5d37cf6da7b1df05f540b9b5ac73463b04dad5fa0e072eb0aa4efe5ac87b1d5b3a9fd
z2867fc0a1e1e76a4959005ebd1e11f52e28a514d5a60bc4efaa6b0cf4730b1e7579b06df9a6f5e
zee1901fb774055beb86678c2a21bead516fd973029df3c578730471a94e69747b78ce5dbd39b9f
zc5516ef888ab5781427d80828296c98018c611dd0f75ce3c498a757136ab98911c50da9cd1abcc
z763d25a288e5dc3496f4c04f5e13db9db6a3bb318ffeaee15aefd8045d3e6151620d7f3628a8ee
z1a65a7d1ced91dae06e6a4fcb88b98b3ec662be42b6a6ae457a367798e7fbeb9382606cc37b6f7
zd68887a67a747e76fadca95239896d290e7dff045ff5cff6ea29a3ebee9f7cc3db4b002aa384b7
zbfa2b3d60a66b69d308dcb254af68b95d1f48d5deb1d0b4cb3333530e83726f94cdde37a1cde64
zd38829313a9c67d5f917fab0aecbf65eb0b8fbd114da725bf4e926f7da23379dd10663190101d4
zafc4bb15002673bb43faa8ae13a91fcbdf2fbb2dda595fb7ecbe185ec30956c7c5c847e5c8e75b
z59fd7c7962a18d3f5e3d79c2fa744bf49cbbb8caa6e9e5a00aeae634ef26a3ef48ed327b90306f
zc2307f5416e2c6988ec2ee8e9b6d56052952f1098b86e00524f7e923527d547615d40b8f2b966f
z14d7780569f151716d955aca0e4f78562ac50a03bf183f58d2b167552da28c1bd9f16e7c290546
z894fc99252cb6251d2d61960dd1dbce74e459b1b86877b0e52cee4e3dcd7f060819dd63a8d798a
z9c0df4322e84a2cc4ec6fdc87049ed38b7146345e83686188c97cfece8c3bd7c3da728c38d512b
z186d2de56c0e62b09bcdeaa316a48d9082e92ea0c82d6652d9973e574e27f1fdeb3807e2a083af
z6c27c70a4c05a5ad7254c67d834ea40852ae7dd337af43a34653950033867c4888bda97f45d7c4
z8e9a9dc76f05da7aac650c28e60cb8d7f015dec4fd44f4c677659b3f2387adc7c2df5df7a67a7e
zd4f8bdc24022fab7382ebe676f9b2f532c0b45fb83be2f9dfeeb85d1576d6a26426f5b9e626954
z128630b75935044592daf2fbe163d1abedf6f58f2d9fe988d2ead056157f177d4de33428d0fcbe
z9670896ad3bc8e05596bcf4bd8959d8f1221cd96650a97216b8a9055ac6b7f98a342f65705bf87
z6777b4f95742e7f901aab24aea81f8cffef591d2ce04634ea74dc4ecf4d673cce6c3e48b8f414e
ze139839fbf4790a67da14048588d5e56c96d67ba15da0939a1427286b779f55e7fc7a755090318
z9fe51defaa6876603e2097318ee1705074fd8e30d09be81acb227a26febacb64d2905d1a70974b
z7fd593006e9f332f445e204e2fadf9917ac633263ce09ae2991b20721b82e318c446cbc0e37d1a
z988d32f5e96a5a29e8e845a9afe15a4e0632fe00c52efa81ab69ab8c6158b7700f58cc1b41b4d1
z776e7a1b65610c41e6d4804372abb293fe9aad44719922de29eaae01fe33e40ab9d945f9d30272
zaf3e0d898724c0e99fc3925ee6e198e83002f2bec633fc92be58f4153f9b28c6006aa5d1133695
z3d75fd92887e3604f6da0c77191c59ee910ca83a7d7188002aafa1d4ea32d439b02bac3d36beec
zb795157ada24cf11b50976a893926caaf496b21da012d5feeab56ab375c2511f86a39660385fb0
za155b967e1ae5b786c6c07c426ca217eddf045e361331d4208cdefea05f31b65f34c5d695d4e20
z7ad02d332e2041f932c6d237355e633449e57e04bc58c2f6381851be02ff95804c2a8440d058a6
z1d426cbb3bd839aa2027fbccae1481f25ac9e79caca911d0fbf7dc151f15455f5b82deed6959b9
z84a1c871618e087714619a9dfb82a11c9295a5ef02f8c06ee37cb63b4044cc67e8203257ecc7d1
z117a04238d5bc199063edf0c8375ac30f838b51c6126c4c08c10d621f8f3a1033f7c921acea817
ze836a9d05fbac0f32eb5258419953d2fb947da2c86ec20f4fc7bd806e2761ae6bed1224b0a9587
zd5aa92eef10862cb4da2e8c070539a40c5449eb5c5d7bda8d4d23c3ec6e6bd1d7aee2b17221766
z1d053c2ae3091134cc9fe37890088c51dccac8665dee24e6070e88d5026f209a8b69658d1609bc
zdc4cb5c5c574077727ab1cbff37494ef797aa794765c26655ac2b8e609cba5dfad29838e86d53d
z16ce95599ac5db7e33cebd726dc06257c6c4750a2529ae1583de07d70e0a6452b82f293e3d3fc1
zddddc462500e1a1eba51106209211b3b4034140f0924e82ad32525503d10f2dd93fd769e034b70
z0208ef5d1e288d6e621b071585433902a6e0990402d6b4240639cf5e1d1cc3802a72574c5349af
z933cb8a414f8daec87b3f37af07dbe2ffb7b3bbf72753cbf666a5975f72c3aedf2216f48a90947
z143044cf4a6e9f19dd04fd6ad14d2acc89977e2542bf8fa4bbe3743e96847aed7b22e43d573e03
z6511909d55d3709c89c4fb1c47c9f093abd7407206ace22125ad90ddefb36b7e4acd7f8df406f2
z3735a3403f0f67c631460d02bd2779c26f6875234298f592a38ddd65c26fac9addcf0dc68845e6
z5d85c117a0baddafb99133315ca6b5251a956d7cf7e56c6c2720993e96f0fea52c1a6d70322f45
ze8413382c1fee14b5061c3d0da6afa497d3cc36951815e94a466f7947765686a36934b01187925
z3b855a21cdfe5eb5f852f8da25d4da6f7d1dcb1745c2a2f49cf47432b45a5942bd9a666d25c0bb
za666bb9e97dfdcb1e7d4df474aee2876b7b2797f78d40f8d78931ee102751f86b2b4662b783f83
zead42567dee54112c8c326324d56330ed7f81b3d70b25d0cd240f6ff165c459da503a6ed0144ca
ze168889bb12b34957cf4f2f21ae140ae1d4d9cd8646051d5263351fa2c21950cf87f1851fd4dcf
ze8ed06a5c8435352e765ef2294014e9f54016b7846c3ce49642457fdc80e65fdc656edcf465e00
z71049b6775af8aa6c61e04faf6a8286e01cc778a7203849351ef390abd49ef18765ea48e78b193
zbcfe4e7a7eef7310f1c574f81d885357b6e67500b628f016f6dfc7a550889634e468ec77b96fa2
z47633c76074563b673fd45d1284350a07ca39f49337a327b42c5e8378adedb9fe49b18dc42ec65
z7b94b23abab016484fbc1536a9eb820584a1de94b1469ed55972870d5df02729b584a18fe747a0
ze80aa7e21e26f5209e6ef8988e476a004517b9ec7d8c7033a08444616b3e3a2604267f780915c5
z955575f08ca5be095783d05a7bd834960a344632c5436883008b07d241ef586ba87c26b13e3b30
za6687d525e2c1ab98a986dfd936f2bbc2d25ae9ba403df2595fc4c6b4b69439c76cc2d4ef8f539
z61959b189de9e766629d716e0559487ecd90794483e48675e4068573505cd0943056c4f78dac97
z7df464fdb8d5eb3dc435878e1065b785749bc40be5d171ff024d9129f15c61c14bcf9d076b90a2
zc2ba46f2c83a9832667f00c004e6da3fbeba8e1d42de0365a16960b5ae006dcf60f30222ef35b0
z889a09b54c8acae473c341620d6947812565c7bbfcc4d3dceba72a146ff7c87eadadb4de6b30d0
z60b88422b5e4dc1f53d54bf1ede0371853a3f3d86df50dcaa157f7b2cc6f5f665002821ee89bdc
z30fb5ad2918928ed2ad08ac330f51175aafacfe2eb9a5a259bee0936c800b9a0605b4b36fb2ad3
z6d8235f72fce0d8e0f186c59998635f162e71c74c0d7a9e7a0e17353f6f3a1e0313a0cda670bd5
z05ab0bf343059761d021599c213f410363b0d2c6eb2941810f271eb63b0a7133d883725141254c
z5097036c0f7fd11d159d4a4969374a42b14af2ae2fc6f7f20454ca92cae0230b85ff66d861f554
zfe13d3694319ed79e61d51748ee777c61137043180e942f2a34884c8d40e4247a20a93c6a995f0
za5a85995e6e569b2e4d8152e2abdab31a90880222ee421f597344e220b75f61f28a106c0e6bb40
z70f0ab5738eb7344aff69efb59c659b5e40a38aabb677bb5fc6c6ea51aaad023893decbc434335
z57c35f836f27b0dd5da4d5b4766741d6fbbd4fe7d82e1fcdf6b589b5abbb7cb75fd9ce1da32a68
z59a006c30dd67e3a288e9d8d4cba614001a9b1bc6ba9b5f1b192d1a6c1cb48c8a596506c2fc293
z70dd0beae37528ce21483bf6f92cf33bbed49385b0023094f2fb046db1e3a0c72803479bcda29c
zf8ca434b4e5beb1bb335d825a6ae03adeee4161d19d2e6d3939301b7b083d3afedbcb8dd39f9f2
z13fc75dc82811bdfa84c7a4efc83f9043cc31f37316a003aaa821ccc639dd96656613b1ded8380
z47b88b69edcf809286eddee6044790c4d27f97ee4e889664edb30ed58d280e061281f30c034b29
z017d72f0f109943a04c2976b27bd842cacda2b7a1b8e2b03f1dacbd7bfb5759b06052422005e1b
z3bce874157cd59afcbacb9e19c8fc09e173b1dc2bfcb369d9bb7dae54af0cb6e2d34d1ceb9d69d
z24c6bf9909c30b26411ec471a42f38067c461a144c8f28830a1cdaa0a0f3926a1e3c00e15d0621
zb9dc112101466b3ac494c50ce610f7bd49ffbd3ad86fabe4f3b174a93c29215d4f2d6f1a7176b5
zf4399ad63a5f4b32b273931831bbffb33c9d6dcf156836003c82d07e9615b20ec56881273a7c0c
zc5ae659106c200e51fd05d925c6030ed92032b4c3d97e6ef0afcf09e47b8107854306440a3a283
z1df581594d077f50babbf09c7686ec857096e9ce6b7bfb50647c59dc6507fc7639d82a54016e8c
zb910fb761285ee1be6a58291efc9e20f416778c5161a4c6db3b469a09ea5d764ddf749b6004a43
zbbefce6d94c0c8ca58186a166295f17a9b811a3f0664ff7675d657479913448bdf887c9773c535
z538355664c73525b70617f4263bfe7359984c75aebc61fb3183782f8e4da15c0731d507c37984d
z13bb5418f2e402589f7746701e65b385ace6f86bf848bac28cfcc504778e2a27cc80a1afb7c0a7
zc4d46ca458c4bd4ee95cc4d45d56968dff39dfad2a5f4d7641a34b11f6cb631035b91ef74becfa
z70db6c31424eb22efffb9402a861554b241aad4dd647fc12e748c8d22f1d5b4e44d642397fe630
z8acd80b19dd6b29e328b1b744157446e1904c4c6061d3382bb4a30208862eeed6035563b674c2a
za3573045c30c2e7fbefb3fb84c3967aef378fa7121100a9a0e798105b89e1deb56ae17266186c6
zec3a7c93938d96812290d8c68523aac727449a0da7b243180529a8c77c48b4a00c522db6af5eeb
z9f926528f97523238a28172e12cddb8acc90cbfecba78a0bd5f75b151978c6cd7055da752442b5
zdd3e8641d64ce57309ce484f13def77dd5ed342751a443ac999a3dd0f6cf062dd31f1e7a373239
z4dcc4646168a0c2a6542e1794710b495c9ee165bbb34692acae6491069d35a0f95bf6ccf1ff540
z0ac7579013fa08f0663467f64285fcc26424542c06f2840e8995c99d570e050eae31a0341fd6d6
zae3d7ef0894d6386e12ebe572fd7a821f9592e0d37cdf69c64fafa1fd0e9e25da6caf5753abd54
z1db26af956786c86aa559f0c79e2d1cd76baa5ea6880fba18f8c044cd6f7cd18b4d6ba79c05f4a
zf492a22724584f1d5463f38cb110b4caf52e6753189717ad862bc2efddf7e2f626346ce365d4dd
z524d1637e351561dec4df29cb67538e1fd957aa9d3f7bc995e16973ccdb2c063c3f2c01325eb91
zbae9e735f223511f03daaef95957749d23fa5a65ade7672139c735cde1ca986db1f4ce889b1056
z166dec27630053f423ace7dc27043551c2c947681e54e7a8f9ef2424f9ca360551de4dc8ea92de
ze32e107bd214fcf3a5ee62d9e4d4cedbe0792f3f70dad1de79feba7593ce3f1b93a77b58d21441
z0127b8633170ffa9d4b256463caa62a160796a26f9343098bd906314af42bbf6f3b80c1bf8adfa
z06bdeb16c199059a8a920b76503c3ec5386427f27afebaf5829aaeb8ecffb200fa621c214b4405
z7cc97ae59d60931eb9ea0c0ea7f4211b21b66fc3f28e9c9134c42ce66e573df3c6bb56830df444
zd0ba965cdf58101ab79afc480a4e6adbc2acca3b19873aa519b0f7e64c20f8e83dfacdc9ea5677
z09071208a2904e289d0b96377b9d7a8fa8e4fa2b9418e73f0fb7212b73d4fdc4d4235610c2faef
z90a5187947b9aee29cdc29b02dfdfa0bb3548cc4ae102f32ff39269a770fc49d88cfa2d90a2c84
z669ffbf2d17138743c3d21397a38b4cc7763fca5f0bc02c1a3e042c179708a1045b1cc5ea178f5
z0dc1d53bdece578cd365cb2f2a08c401a78a876336a14769a120a30d5803fa6b18b88fada08a2d
z092317563fbdfee38ccf73914ff4eb6890330075e4266f081253fb32d192d2abb55c666e499691
zc12e4ba4dc7b95d772aed5ad039baf10c7e8de4659984ac0dab1a126151dfe7f7e06d6640ee3d6
z98269f926c3e629e8f2325b93d325335a7f134fa7d65e9be9c5850ea48f40312416d1d98e4ceaa
z18987f867704f959fe7b05c9b937094aee2ad21bf2086c14eb4cfdd1092321ec831ba375aaa554
zbc24cea7884628ef49fe00cff8ce706cf7ebf4380070df6ebe81c0aaffc142bb150573bbfd6db7
zbb9d6c7bbe07b052867e80babb6698a6668f20e2dcf76ed3561c7e0620d8a0d52ba1cdd8f8b7af
z0d053f96c30150de76be8788d7f6f5f08216eb9c2d9ddc2000d8598f1dcd78a112dd0b0d40ea4e
z59d323bc67f8a6a5b6e98a42a2bd249e072813801fd5ad1fba6b78dad7ff5b4945c74729132fc4
z9cc15b832403d02d432126d307b4664a37a99935441d6a597e749c70781914b1e6cfba8b7b8154
z8ff7339fa14e05e04aae4292a4c13fc368b3171a1c7f4c6aea8285ea81ed6e957f25678f83ed40
zafd91e2b8435a59c44770a62ae641f0a2f9dde9165890de8524927017cf3a1bd1f5bb8ff9314a8
za8eb366cf694af7ab618f22159926a79bc24f14a9d084b94204ec5401f025e80d514c217802d13
z421293b503a574ac7820b3270a12180b85104d09b887157a1ff6c1aa982cddabfca9b32de8ec90
z698afc1d7bf8bc9a0166695ab4c271b963b555fd668e82a861fb4229f3ee0d5fb13e9a02fb5e76
zca63d323116349097f64d4582cb811dd61691fd1eb0a1eeecac1d367ecbb503b62da1811e8324e
zd6419709de7e16dee4d2cc40a1055a497b9402f2d53e06b7cb770dcd9ca5912ef68ff07774cab4
zc7bdb30217e6bd57f1a3497455aed0fdacbb67de17903ced195c16140d7f2ea51d3c7f3d405b06
z49ec8455865d7845ac95288a7f08fb530456306bd7ec1588db27e3531f60eb0b6e07043edd6dd7
zc284747576e27d6f246edf3abcf7d71a647a36d2c492208e16ae768c5f032d6bcede6b5bc3cab6
zfd54f08870545e58aaf0a8d55b59d791effca86a02bf54ba05a5054d2429a562da108310a29af2
zea937a00c0aa975397ae8ed40f3137dcfba44ffcae321bc0805bfd199e30a3890ce93f9da9eceb
za53d81a2871c137bcf87a30dfd9ed528ec621366bc705ab723732c015c814ade850b3f98e7e715
z4a5ae420cb0f1e533a53148df7da4b67803ee7bfa61cb17ec2e209a3fbdfbec7764727ede185e3
z8941ac8624c4d2edf9090b186cef7afd913311d8e5ce9a0e1fcc196e7d6e066a077aa09df2ae01
ze2febd4b84c69615f49318a2d37530fd8da1fb7bacafa4b2606513c0a7179177666aabb7e16b86
z7ce601a624f54bbc458756dead9b1c7dd2adfe5543701302987a67902097397213322f4585af58
zd0c92d89ef7a9116ed01f46cedeb738dccfd545b892305613ec1e32c398e1cd78b5858db86d0d6
z22cd6358e675ea707722274a0562a5ff6bca1ef62de426f03aae19455cafd98fb557b1baddff27
z82cde228343fccde4aed5247315679065e94e6fefe63c3417f1b98357a2ba3232c3d3608ba4d98
za4b6099715dff52947801a0e43e294435bd750934799d360965df7eef90b8e6da0174dd4e36df6
z3a452e38898f09a90b1908813a105da45d9e41e028fb688de0e40733c963544b7e6197227ad722
z9f03b86ffcb0f0fb0b78fca309fb4eaada14cce45ed3fb12189e579fc2473a374f44b3d034acf5
zbb4c43a1369e751509d81efd50ae5b38b59576c5c4079e1436c20d23461b242b75e507e23ee2d2
zdcd53b4fb1c1d53b4488e4bf581f230bed2f39572ba8d713b40a0c4f6bb4af70c4c55edbb4364e
zf1efa8050dcc6f24a012f80498d8474350a913c4b2bf52d837473755e86f1efe07f80008855a11
z971b846b1041d6cfb31f14d301f1f36b033166e1a5683ee644eca9b133cc85c5ac246bdd59889e
z569766358ee49e5f74092fc3c72576e5812564aade083c913d61b50eb8138b0e8224076f24074b
z0f7374a53b7a3eabab960c0a82acbadb78bf415c9d548ed18553c7dde61b5b4771c6dd7bdec117
z9e85dbfcf4e07c59b208ae79042a35877a6fbec7450f4eb1c02dee6fbf5ba2e38c76cdbcca0808
z1f8c960c39197d8787abc7d89c53cf0d7a38ed6dd3f4bedf1d8be1950ed49adfe1ce692dc2e1e6
z6cd75de7340727df887bf0aa878b08b42ccdc3eef1c6fba208d3037d48a2575f6495794178a738
z0af0ff5ec08685ccc7655c4df00fadc4d8344e9b2826c7c3ef8145fa0d14868875015dc5f25ff5
z62a1e1bb0440c83dfef3fcc931b7d038226ba0c12a2bfbff42b2c25dba50eaecd4b8ca9e20e2b9
zdeddbf2872f4f396c5cbdb5ab4021e7c38527200024c6d0b1cbd490a38a91ec979af1221976972
z00726b316c8bdf2511cc5a9ca8e4b359e92b3c68f73c7c73357da3c2c51e2adc0e30d88796bca3
z98ebcd2167964b2c78d71bb829bca665833f2c52b9ac42681da4f265e1792ca7cc32d1c9420e9a
ze93dec4958852f5ac64784a4ffe94121db08bd4c64aeb0c0f6106ec31e6181b7ef6181956d4198
z7a6c9252123af12ce7b06dda80846a6b537c8c8936d8139b090451243c2a3a286075aba62e0f10
zd86d93e08bc6eeaaa1cf3406163c25425802f0a118b46762a3a2d75cd1bb283e5fe16a0e278409
zd7d14fffc60f8cfa4aa916c9617210b06bbca22fd5a82fea714f48e45acb51b8e42cf1c3dc037b
z029003927bd58d6aca030508ea7c50eb2e103f774c88536bbee5e8a188da068d6663aa7e35557e
z2d7054a1773c4cce5da7f25c6626f4eb1cce51377594077ade5b9fdf22f2bba850393c8f28a9d7
z96cae019fa0eec69dfeb6e74289309f72043f376d6e444009ef0cbfc300b553311dca6966857ca
z9fc61d0f2e16d2f22e603f10f14b06661a1688bf61fcb63626155e34a4a3edc91f0695933f91f0
zd608dad21b03cbbac7563b9944326793cd1c8b3ab23c829d03ee5eb49856d95d059a4891bb1fbf
z12f51a68a595d0c65e3495b02722c6aab018d2fbc52752a2d92661cd6e43f47a00bbd670740e0f
zd3a225e6c18b81f95dc92f4d2a6df5e56653b284e8d0092e46953358e7e7e1821cae04f702c661
zd7b931e6a37e33b1d61deb5a4fb8de29702051b78af6f57c9209c3f1b6c2a37bb3fafc16da5ac9
z890e337cb2b640462e45fe8e234735188ab694ff38e053220267e7b922cb169ad5b3ab6e2b9099
z314ba6c953bd6879a4136ca0a6012345f84cf843a1d25d5a8e3fb33bf4a7f69d4cf30a6a14cac7
z14e61989d15b235b806df0585a86da878a5957a5d4220b1c484a7f694c51bd72e9109ce99ea28a
z2961e0ae0d9e2984817433cdce7b8e3978d14a18f8df583668a12c2b31c781b2a99c737a1ab6a4
zbfaa1d9b1b28395aac2ebcda414fd9094c75dc829e58261446487e911a9179c8b5551bdbbce888
z5e04e381ed25e1876a3812e456473586c6fefccf0d7e17241ca94d5d48c854f72f83c699d59786
zf7c4b0bb352c0cf772e2c662d59fb69a59786b49410b54f9760de51702ac296cf485f84b00c8b8
z791b7ac3dcc606a124ca852baac1d5a8397568bcded8588c302cc029e89a9add06c6ce497ddd2f
z242aca9f202978c240310575ba4b85e0cc11e9426ae6a3a5461fe6b5f5d648c562a4615b15ec11
z597e4f51f01ff06c143fd8e11d5194efd731403072c16367c0885f347becfdf7db7c3c4e753742
zdec063cc4bcc3be16021e72dd4b63f301666989688e5a1440965ab7205f3434bd2549c097708b9
zcbb2d82f235f760f70de424b8ed94fad3eb1cc9f749a35c21c59f5e69199bef9f112c701badac1
z68732629c765e18c7081e895865c139787130fc0ebc55210121f11361bda535d58b8c152799bf0
z7548b66694dcd33d5ff2ad592800ff4cd3b9429142bb5e201af32a440e778da33d690a92807622
ze566eec746c1fab676f9f7aa44165172d5408800d1b07d8a0ead8cf563203200bfcc0290e6a70b
zc6ce156cba064ee92205d8c2ec779076f7e84db5f52bd79122a607fdef500f95d1a9ef903c673e
zc2ec5684b3bbefe76eeb8a4f26a5449d952c29c6c9c237b973a5aac6b777a4a510082be7f20844
z8f711143496f4213e4c736889f17f39684f012a60b10cff78143534658fb05db8b27db284f0418
zead1fc5524338c62499e821d0b22b1a5dd4f7a1fd832cd8764829fdb154de61178cb3fc5efbe4c
za80a9cf98ed725def55fcd584ce6dbe2723e155078ee0b56d3619ba97772ef61076ba3752f9571
z168f73a2b7c75ad921c3e6839fe010c8ade6fa1a7edb2bffabecc089533c0c21306f0a40a1922f
zd579de6c51406408f61acdb415d9d8398c84262c43e944816d769a03330a11b96cf3c6aac10928
zb9617d2e91cefe2b442ef3dd318cd4897dd08f96709c07f18c22a6412d06e79569fd3ac8c8a29a
z94b628ddb00272b10aff06054cb4e1080c5e67f600ffa0ddfe123080da2df8c5b6d9be4b82ee18
zfb4078fd0f1987d9132218f80f3655aef0144a3ac3c4ce27cdd025623594a1a8585a916ec3c6dc
z2722ab11a181ca68adda61c56a3f0530066a6a08e5a52558396db2fa0d1b68dad271ad72a27116
z245b9a3b0662e0a631b155b7d955af9721819c0846a141cdbe1e45b3d85bb85e5582dce5da188e
zcba375e63f44f08e581ec84b46d7a4edb7df2fcdaad38ce231980a580269bf3fcaf4cb0fa5bdad
z2b2ff8b08b20eedf0d9ab77203cd1ee1166836951d101022cb677711bd843546fbaa6608f53ea2
zaac7d7845c956f5d696a35bc2dc01a278de8860b85ffcfeec60cd7b2c87e23616a09056ee80d85
z18a2d0e94be5ca6f7f809dbd112a5c5973caeae152c45383e513de5608e6383a6cc098c0f05dc4
z47d7ce6f9b1906f3f610e7bfb40d95b573ceb1ead0c7bc5f7fb80e3d69d4e5f97593b883d3be47
z09a23fe7206ca2940e04ac08b142f18f1f53e081c20adfced7fc98b41f48ceec57cc36ccb9b2c1
zf7e4b7b3ecf75ebe5781cb5d60f4ab3e361fb39cb2190686118b7d49774d98001c79d7079f4087
zfc54c98e3c03447c4563f86baecb3f8e7418ae253be44c3d17e50749adc57012b26b2cf6999cf4
z752f41ef10c89710f991bd9867e51073eebe1c8e97915548580857c5a1c4f2a32c2e1ec57fe796
z5a8c9098ad482ff246dcf13a4926fea405e10a5a2961dec6d684215d0f93d6d42b811911f8831d
z7568fe0c975bac7faf117b50fe9dc47badfeb0c296a133cb627c3f517559e94cf2d37f76eaf019
z47a29a100ca95fbcd079a68414b6b10b13235a7cd9030b77ada9561507e73d832bbf589be616a9
z5baa978c175b0aeea4738bbd06b1c51d39bcc82f28d7d00e796adc0b4f10ac0276057e35c0df64
ze5253dbd09a008dd37d3d422a757ce57c7b5dd4d076b9f2acbfa1290ca08c20c65248d0552f222
z26992d2e8af30b65a3089ba67e7b7936ac879c86743a72526303c82323dbe06bbda5e5cc29dd50
z1bdc73bfa9701b3bf836bb77bb49ca4182f1a84d070fc9e7b6e4387de9592d9bcf197ac7f7db93
z5af7f2d23f45b758547e2bf665c84f30764f3aed7de8952d01a230c02e9023ede155a54fb192ec
zea523dcfd95ec1104c9b4496d3d2717e528281a46f5ca7fe39b62200ac9f2341e88927c1bc6cde
z4d975baca35cd8847cfdbee7838912126b8dea2bf9617525164f32118bdabeced779777fac9904
z40dd18489e55da5fc334c5a05499d011aee16e5e25effc69a552c4c6c9387c06c3fd1274e13d48
za03f28ab131aaf8fa060402183e0367db970334f2bfe8ec9046dce0dead96a8783830e9a5af0cb
zd1fccb8fc5b494df2fefedc3f170d56f44ff6ccdc0572ad9d6a484cfb6357183f011b4d3236979
z26827c41dae7e9ed30816ceca01de6728815271673adb913603dc020324d9f8790bc73b5b7dd02
z263fa985cb3b05f821befacd43a4e10fd59b3425d5ba8a118141d887727c3f7191231e1032db6e
z0c0e702fab8cebbe2af30099d8baf6a0edfd16bc15dd9d4be6032029e04deb7fd324a496cbd1e0
za2a9e1cedc2d75765f2cb5ff1bacccf9473068ad176e76a8bd91d53d36487854572f6321870a02
z638e2ed7b67e5fa3521142b9fb038982559f2f3de24f1a23c32d4d84a068d65c49ad83137ee7c5
z59766357a7105a522bd446d3d747dd54b3e7b798f2f6ed5446bb839597cc27b3398c460cd88caf
z1b91344c0031c9966590c4caa62c70d630813d2d9179e043d308bf4837e847ed5fff7682a1568f
z1a865bcfcc9f36e0b65ac202b7bae39919531785d8ff4fd52e4562d4ca90eb1d52276babd55144
z39e6f726598d6950aecefd2c2418661e16c2d198ef4983d2f76d8b4ab82f1381686d332d0b9e0a
zc0a65592e63afe89e2b0cbabd56e66f1ccdf352b0f836e2119e03f70ab05570b3c039523122761
za01bd09c7faae770644f17ec26a3d3069bf734129234deb5f0edd0e51a2bded14d279ecdeade36
zc5a8af256435d94b50f517ffe4be2dc3f7655e018a37517ae83f941b29f729c6a43bdb17fb02c9
zb5a77a3e7fee4eefcffd985a6a2029eab014cd6db6ab27a329b5f2edf494917163755a0ae22e2d
zbcd9aae55718ea8a21982a702f16fc2fccefacff3e7edf31ae37e91af1aa5b65ce2736d4afa824
zaeb5eb5e4e4e7869dfeb1a9b7efbb85c8b2b62fb5b8457a3a11e728f65abaa0f5edd21c424c70d
z6e553ea690d80b455ee3d57e0cd9cdf53dce6a36ce4ac23046742ff58812808ce1fe40679d9286
z9dc14b7719828fc4d827e244ec6477745931725736f2ed4bce023101e87786db6eedc52a284933
zac411ce9af6aa199c158693321de1f599a73d9f3961d90be5b1ecc7efeb4c91ec283b362615f2d
zf05c0b8d253f632c5a995a7951e1aa4974d621e1d77115bd97952a2bf28d7bb35568f2108755d3
z608773147fd63cee42c2f3b3af0fcffe2eefbda1589b3547711e0d68b15c161c1435afd555b211
z116ee16e5343e1df4d4a99b3008760fb9213edf3d216f0aab35860a2843a832c4a3a465f56b7bb
z3897cff9a09adb221a19b0c5ad12144d73d41127e55f20ec70a577a7e55981b027e935c3974d97
zbf95ea19f218b43203cf8c8ca63f24eb0fa17574b2474a597bd58e791401b7621c6188133b5778
z611d88eed00d2f4843d902e0b0fee8e00aff424e65e50d43bd24b9faa482677ed4d4b9fe8750c6
zfa554f1fee055d8b936d328204f84c5b6957d36fd5a3bb8b5a123d5b912639b49658f04aee5e7a
z6830616bd7a7e8f2ee1879c7966878dec7fdfbdf3b756b957e8a26860ef05241c618dce9127168
zd3c1a74e6159545e8f396ae548e50c5d1415a306ec8d7ca7b6ddf754db7acd2a7f4320e51de8df
z174d72a589896f44fa8ac424805a49d94c7921ed563b87909a66c5754e54e291da19a805be01ac
z6e01c1990ffa29023f71d0f84ee8d264b479aabb5121cdc6c88f621eb948bcfaf0898ee73dd584
z30e1a7d282645a65483de379fb44fbc84aa93dc11fbd6cdf314ce383713bd9f713ceaa1ca518e5
z1c5666903c3a7638d3e58c2c286b44738cfdb7cea579aed54e9d0d4141dc8d9571ea2ef55e9c9f
zdbbaedc2ca2dba7c6dc5aed8687e5912675cbdbb7e7c4d0ca7047334ee3315b2bceb38d2f85555
z7ddd250fddda92d4dbedf7a202300d0ce326bd05130a84228e422d980169d3fd5099cfa52c483e
zeef5b6d0d7398dba18fd9231c1f7a71d8b8620348f34cf1fa3ce1a8e340d9dea3ca3495a0f84ca
zcee153a6b8d2a242b69d8815ddaaff6c5b87b1874f6ae4011130fc234fcb87cd64ae45a869683d
z62d134fd732348525380ee442d1afe0eb685d157b0c1dc8ec0246b6f0f483a3b85555a3c71faf8
zc600ff74c58a08027d98aa0d1767de6d2559d0006f867d042dd4fead325708ff9ed3553aca837b
z200f6515bf207b3ac23ef4b255e2b71630364662f66d3a19ebb5cab4fa40ba23eadb4b9eb290bb
z786a3b2eb97d9f84bf5807129d0e909bb1dc4f371143f7e2044e5b8f8b0aae77c564e7bf86adac
ze6c0191349c1a444a23c3e2396b9d0fc0fb227bfb8d0965564d74094323b422c9ebb6d3c5894eb
z65c4b4a8d078d395acfa64ce1826eb874481d4588ae18907a383d9527f88b485a871ba5321369f
zcb1c115e385e5bdee76a22cd26af39f3de664d6a1edc5c3fb21b3506b1d1156f5f7983f74b1b76
z28e4a37311b409b1173493ebcce8a3f0b13b75989ba8d34d9c4ee516e7750cc7b16773542664d1
z56282f3c480b7b4aeb39adc79ab08eb00d8c17452877263cd0c9336c0b10c089c34523c6fd24cb
zbb723d18d9452bf229943105177a8a563f8fb54f72dd78b004b30f532b2402cfac9172b297a669
z6bf357feaff064170de8dcac261cd4c5efcc04e59b646635f5738954959491484d03f40f6cfdd5
ze9c1a185b9e6de3b5270348433b9023c85989c1e0d020be15a8fceefbdf71650f0a522a69c7491
z8dec370d1cceefce9399e21ebd96c04739d29727ddd7987c623ebb9175d3db1c1c5e5f8039a445
z257a8bde354e3f849549a4ae857649eacbd1e5e8870367e653e5846087b156a7116e109215c73a
zeafeedd5b86261760ff24ec25a66483fc9a3eb50e3ca84a5f92a2ca85f9ab3245f04f5d805a6a0
zb648a2748df35806bdb6db5eb0948dbbede52799f9e7d0eed7b2d0a6c642b68b14f337bc58d8cb
z1a5c285087451cd22911760721aca3da706706dc97506524a736f6e9b29b6a04eb6b60c70e3de9
z23a4e26e6f15eb4e893dc2b0524622fb2c1259cc4ecd0b932db8c7789b9ea0cf4944935e489a0e
z53393ba709c1772b621dc53ed6c3df9ec41d6ea5fabc1ad9f7c38a30466b652da509a3350bd0ea
zce224e98f69de8b0e9f0273de978d2e28bfa2f96f10ac8e3c27e6dceccb6c6ec7170c5d08cffb5
za09238d35f29c29f5d9bf2545af32d3c9e1e11e2e96766477359a2eeda392f12dcf023ffe918df
z3360889c7dfaff3c5e0097b0e0a9a582380c351ba43f573e4eb62daac4ef95f8f318f75c3b89ae
z04b0a209b5f9dd340e41e2f3d10225d5a3f5c1a483cd1a91d6107dc7f6b7854eabda2e0b752ff4
z130d2a1f8f990d5cf12cb53710a0cf50a618bbadc684916deecdc36e4f253be973d9b05c9f6680
z2db23809282f99eb364f2163b9f7f07e997dffb1cab076075d968702f86f97196063878bd8432a
zb9e178df7bbc48d693ce94b3009d7cd1eb7c0d232ffce93a9bee32bb43d8e0af17b29e05f7fb0d
za327e5aec54eb1fa3b0fd7baa1cfbd895cfc935f989941e38c065edf71da91704a19cfc7c163f7
z4130170f6b46703a7c95234c6db52797fa831239c34d26b872b7d4777fd813550d522efd8b245d
ze36eb39131566ca28616f2cbac18f765928d1532e695cd982b087636f84392f79381a77b969727
z7219f598641c8249313861c0c07cb5bb14c292dbe603ab345fcd3ce606c4e598806e7008684bcf
z059bf3a91a864cef3ed825165c75cb9ec96ed821ca3f337bbf5c1298bcd9a977431dd871d126d9
ze443d27f31923fb8f53a31dd6e71afa173c8880b1378f6488809e916d09b6d70a93a7f77b384c8
z5a455381d22be99cc163823ebe751ec93721ddb088b760c397d72f73426461760a8955f3f467f1
zf47473ed961c0dbe5d63175af6181065f1a0930aa0fc1313116142e701c7de4d65b5b2960a0f6e
zbd9fc7fb33104711a09bd685a5e47ed55c4eadf487a830c33ab287dd0b55ba87149f4732a3bbe4
z3ff2ce6a9d0f12fd6c6494c755009ff61162f0bde4b6cfebabc416017847fab5bfb813d962540f
z351bf569fd56176bd2d1da69f821ca8d860337fa2543156984f8b9ba7c1c55a8b4e614972da88e
z7117bf0fc5e8d276d25c50fd14d09238445a91dca83aad20d842ef31d1f1b54555700a3b3ef8c8
z227d36e1c9558ff26e4fd193d6f3d2791df8adb020dacabe529983f711db99dbc9a95fd106bc33
z3077a6e59757fdbccbe4e6b500df227707967003a96c6e3b88c5283dd0c6003a8087a73e0d944d
z07d9406045fca4e9a8c19fccb22d7bd1063c66c073a6e685c9e9b1bd98585a73bfbb09ae48bda8
z7f5aea630d7fb7bddcafaec9bdb2fcbe113cc52f9bcf52c5555033455284c35b213d79351c2eda
z80206848346fe1255428515ff2e9ad2c39bd4238f5630469259e4e3fc4c85a4cc3d211bc1b80b4
z9e63d6b335c3f04dcfb3a9b78f07d1a161d81dac0ce7fc4902a7adfcc2907b2bc729137cbfa041
ze5b7ad6c527f0afb3c31da521b2996d094a057bc154e933096f24193f15edb6a9082cf60e11f10
zec9e4c834398bc207d9cfb62766e6adf1378824689f735c4d26dbbfe64413d30dc79fa4cea2143
z3202c5ca31fca83f9f0f68ca2e29347c8af81054cf42ada56bdd9e58632561419fa053ad817457
z9569d231458cf02f1cf1ea34f2c6818df1a9a7733254f0c7efd12c9cf77ab1981470b0a23c3312
za03c89c5030f5a6ba3fd2c81fb1769659d13e8aa9bd5f631123bdef37bc5df142621f03b9db41e
za53cf5b2275e23edb0b8600c3283209d91c5939ae5a5595863ee2c736f0c37d17e0d7912f4231d
z120a4f441d47970ee4acb43a1bcff8e3228fbdb2a9839372ff499e470b0d624db77972cfec1182
zc75c11adce84540a19c58d5e78d962eb6181d57be11e1c2cf6f063878972a72dea747a33a3b0e1
zec756f7b892d1115899ee4e5a4f0613a9a65e716070959ae28acd44c2d30699004ed0a15bf873f
zb0f2867140fe5b1a4b023e79d21b2c560bdd9e41d616549dba225bff6971486874051f523aca4c
zf626266ceb172310564fe36c7f0ffdc7592b12e8f6ac25445cf0b61ee7a3e6e1b7072b81bd6566
z021bae60797000c6c9ade52d0ca2b9caa717ad2c0071240af51fdf67a7a2b71497ae355b542490
z06414502774a4b0a034eed6a031bb62ce5db1d8c0b67fa55d72f8839ed4b46dbc0e304a9061e87
zfa2462602470374c629d5345de143bebad55c81a3a3b9e591e75264eacdde58407b25ed741993d
z2b7aa307d120e922a38cc701dadb3b5bdf83da6c0954285b2e3df4ae1026de9a96f241d9a29cee
zb76182c0648f85cac8bd5be9e123426f4264070380b19e066e7ec9c946ffb21e257e8562d2ede0
zc6a943fdcaae4405cb37213ddeebc67f0c85dfa205c76ce144c57ee3d5bed41a474d2a5d01a62f
zd37ac7231adbb8b6c1ca3fb44493b71bd01db08fa28a03b701edc030703bb1d63a462f4b9aaf20
z2c68c0b9ffc5d93a29e196741289f4032ca3479a4d7c7a571eae756fed85ebe487c571ff3817c9
z20134248c6853388cd04fd86b432e2b05653035212ffa473c44300cb2b556fc05372238c62d180
z9cf80aa71c83d482621f9a984e1bfa29c74970aea905a8320c954722eb680f46559982027487ce
z63e175864e815bddffd88dff66c94015acfdb29de9afa0f0e78912c603b8db6005b3234e347900
z445ee58cd6b7514fd500a43af0eb87bd37cecf357ff9097a0b7a37c79e729299f41cd9adcb81be
z49d457fb04fc4df7b2edcadf61ae0f3fafcb6f0cf0533733ad79490f967494ffcfafdf6f8b469a
z1358d1165e446d5dd73d1e04900548d52d337f96f3453f3ea7f652b1011941b98558723c57b716
z2aa4bfccee35450d775ff1c09ab6c46c9413d3c870ad0cd085876588026d5274ff247d0ccd00a7
zc7cda9a318547f9991ae18751bc506763543d2acdec5193c7d8c68db8831e2f35249ffb262fa6f
z96020bb311aca4fca247fee85f777c358dae7a217a361e870f004fed9ae62388278e4d30f7c25d
z2a4b1c5875ee945354d3f9e791a373bbf3b7391e4967c768c6b7d283ef1ebe54f9c16dbf4eebef
zc8e11fcf170e1bf7cf6ec311c9c9f1ba81ef239cbbe0b2a770d5898c6ec3aa43dfe74f1aed13af
z79fde12515f7604148fe5fc89aa29f1c9655e012e7fc2952c2ef2b51d57317ff08dacc5921a88b
zfd1bca069d798c699a4da4c03eb7461fd410c7dbd473b9be4e508996cab5da4b35b8fbb9e18090
zeac5004bcaa17d37863a5e76c834ddf2ed6103814aec44b40ae316aa9a63d76196f401e6645dd2
zbac5aff574109232052e6102dd2c56bbafa8cc9bedc53c8f69c7c1db939b347a4d2f95ba443b93
z399e75b8aa4058de6842c9bc9c55b6ead75df6232214cc6a96460a53a732bd8e02fd387747a986
z5a37f1c273de904f96e3bde61ed0324d238a7a6c486c19126779423d44a4edf8b5c0925fddf3d6
z5a46b47fe169acb130a875b5c551c841fa48d923c61b52615498843787406fa3c999a6ddfe862d
z5ab43ac1d2cd187a28233e9dccc440e445e9dc7a6104501cc78db38d0ae8a91d23e4f490679682
z3c256825f0c4d6e658996666a298f7ac355ad41443a85829c7b306d40a2639946fc33b632bd3f4
zd2d51082a6f4fb3800aabe764f4bf98efee9afa3abd7c8a0692804629e1571eeb67648002db9fb
zd0d426fa37b12cae103d7b8a269ab135caff7096d86d245d0b86d5cf44f17369c54748775fb3e8
z5f477d19f1c28178b0a4fdc1b8d2b741da76666b049e2cfa6db4516308450a678d9fd4ed38a104
z15cc213b15681ff6ca8f22ebe98854ae796200af43830b2ce54c61c17ddee7b3d6d262b02849bf
z8db48ab4d9dca1b9cdaae2b99e473e018bca73c21cd20d20abc690fc04b6e61df0d9f6a4c14db6
z14e81b79872baf67cb97adbdc93c80b5c78c47653644b9b22b9fbc3fc18cf21205b867d0602289
z05c3b44f6ece118badebdec74b45813e33c1aa4253372b1ce1ae2f736b4706522ae1caf62755bf
z91b63a31b450aae202de3cb74da4fc4338ca805b773750b37e55c5dea9575b6cc0e22dc231f1cb
zf397efcbea0909d7a509d56b78e454015d6c211d967e68f5b112f5f89bd4aa6c6de1109737537c
z885c0eca46723b4afbfc73213b8df758a0592fbd5addbba25dffc1faadeffc154f707030026da9
z120a03f82e596093ebf8b8a0bc10241eb63bdfbfeee6de8921443718fe30ca2212bb899016a0f1
zbdba94acf38f502273547e2275eea757af0248c8a8a89a892295f6e2846b90dda3de6ded0db7c1
z989e6da24de1e67e54cc31518a58caf086c6d3a3c6d5e1c4e6f98ca4aaa77ad33cfd4812e94388
z142b71fbaaf8d7cda231611a9cba95b33cb525d12b5e23394a8ca9bf982ee45c39666a554074cd
zee0b0e1e19b9c51431bf465ed473d2509b9a3cebb70a83e5b028446bc6e074db86264c6433796f
zcb6f4fe18b9537466a08cf4508f04f7bcc829fafe481ad89eabf9997e9f87a3d9b2e3e3a0bca73
z0ae9f2e478ee1438948abaf16c1f2541b14088ff5716c7f60fd3624c5a267ad716377b123f299e
z3258f32e9c65755db1396e3531ad795364eb3b1673afbaa15a1e50c59ae7baeed27bec21fcbe6d
z55589b200ad78044bfa226e6b1c0175fe42493c722330ecd7669d8f2b9b5405b6c0fdb30de25de
z9cca70d49de7f7ee808765fcaa93a8457755c4cd67197bb81b27e724c10b3e9178ac7390a521a0
zb83b936f8948e79241d6aa7115c59bdeb5fa6b1f3170f4651d4a475e0d0a5f2d104736cc03068b
zfdd06f8bc1d9c331414c7be1ade7ef47a9e2d279891770fdc7714aefcf7e99d233d322d6cb8b45
zfd0f7eb5df32e00231ba718ad19e6dece6e07ce9875ccf4e8a211f4759df743a2a5327c258a420
z007e2f2e37a9d60bea851640582def45bfbbaca8d344e11883c7d55b13388dd72ba7d6f3ae106d
ze7cfa941dc49a9bd0b6f87666d0ce92652fe3fafb82921bb5ed11d1d82dc3252b1dd1062a80424
zf340087cc2a8cd458b795f63461fbabd2e8c94f4e62b3e95e510caa4169899d30c32dd7a002e0c
z9d7b35d224cc07165a44507d2f74f5af884505fdc339a4bcf6d6e9f6fe59aac4e68c38de097abe
zad97feec24f86d776e5d93d79f489c85e59a38f4d2884cb978bd73e42198104ff70825e5969714
z5b1ec3a8c2019701a82dfac3f0dc33d467c5a1a1a190ba279b2da10eefd7bd6de0078ff1840dd2
za4f6e405bfd3c830cf0c2b7220ff2832e4fe32d232e1a79315c43454ac854500d98df05ff794ff
z90327197cb87c532477f910857842c58b4afe9d874d7644f46e5dc51a5162749e5ad640a0d8074
zfce5448856c598975bf7afe39f8fdb9cedd0b254ab1a6261f14b78685552313e90cd25fadc8f24
zce82808fa735dc46d15bb19bc1cf47a50729b938370cc8c2da53db7b4e076275099d843d18f013
z25103b29439e0db50ff25733fc743c88ffa0b4713e80bf1f49bc9d563b3cc59118778d50882369
ze7f9171af9b36e94774d476d99dd03e8390efc5fccf2af3620014789a5d15a2ef9ebd1d05b09cf
zdc504067717dc4fd633da7b346b5b0afdba6ac9f98202d0008df156b27f193dac9ead1f065baa2
z83376814e674a30fb236d5da655665de7882e0bd89a579d67d68fbbd7276b3bb51399a746d94a7
z6c36170924891e602f7bc953c6c622b35bf64dd0605e80f049bf7d125708d3bb6963281a52620f
zb6701a3961b168ea84c920ecdf9d0f204b6dadf71e3d693bd918f360f926c7fea1edb0b697fa61
zb8f8c15acceb6e9e690a0ad6078377b463402b903e00794153e61ae59447f3a52d35b5c493d876
zd69ad65973a2973719bbd7a17263a9ceed95e8788cbbd96b2e400899773b68c57c982f9b55c698
zc149aebef309b16f04440217921943145109b5dd64937b395efee480a5f7898dcf65dea24e24fa
zdbc275a486ac9a54cc3f4ab768dea8e0c8848a647bbe873a8d24435496ced4d7d661e6635dde1c
zdb82b8a0c045352c4c19740fd9e15807ac5e0804b0159fe1707fe0d38b15275ed889a344bd99b0
z5bbc132ec1dea2a9ece657192ed8e88051801b9e69722bf2fb42f74c9eae8dac18df072ffec42c
z174b5eea44af7a0dd0bed2ab9d99664fcd9a681cf46eac81312972c19fec45fbf26682fb57a90e
za45a22cc72373c86381225fe551f1c2d9a7e17c0810602279e7abb5c203406faf82976b490b26e
z220e71009ae003c3e07da7ce92e9291e838492381e99f7755e1282275eab92c0973d2be1875515
z50e1f6cdebaa96e58b0a533b5cd26af04af72e71c78cb9c83431be772fdada7635ec5f12946266
zf70ea3f51d5a0c6de7eadc644d19a93ba4ff4da09d71c33fa73471931dc8bb73663d29a2e77799
z0d35abfbecb9305e441dd56ddc115075e0f24433fb3b7016945af41e7ae6c023aaad8d6545a1bb
z8b76265d23fed352df8f7f0251f120fa2144170ec661d696b59b9ce8d9ffa66844c4be1a5c1701
z26b02895c1445869bd61b086df553786cff2169b686513565d6f829cba05d11f652fe3471257e4
z8c5f5d6c4093f9da18b8640a510e6dc58c3fd19bff0ffce582a084abec008e8b924739d8c4c81e
z7f414e07b476fd8b8291a792e6bebd76f581b9bc60780d394926888ecfdbfbdbc3f462a9e8ea0f
z49ec17697d0025516525d2a5fc93d2b7e7f982a70b65b72c84f3cb972d330fa40ac623fd0b3159
z468888d5fce546060c210c09225bde0f7f2580d99fd7390fc4800c123b5c8f135c4dbf4f94d4bb
z7d9abe794ed0d3c7b8bcc28127799efabf1b2f2917a750b50fa7959ca5d20b5993bbf07b9eca04
zfe03631972fc4e23392443fc29836b566e3ce56a6a25044e94a8e84075d944a75951645a55cea7
z14cad45e8d016b19f94e916f5743bd6ecd7794695cab2031c8ab940bb408455cb56ac5093c51c0
z911144ed8235d58412c4baefb603b690af835ef6c02a3372aa36c0635cc85cad3a41064c75356d
zd57120578d720cc3492191cd3b5f24ba5553aabcb6836107551df8098a41c93072af3fc8479081
zd26c0d6e2030d2b5c85b8b80e62235702dc2ca31b212c8b6f5020d941c9531e00f1c0ef65511c0
z61860a10188895f14f0e53473485c4fbdc2a743eddb94c031221cef8ccf4f70397806b2a8ba8b2
zf84f944f986ed5ad92dc59b0c2e73d5c2f64cc2c24e57adf2ace841688dec8376508749997f165
z5a5f53bad3b19caab5b18fb2748ac4d993eee2a265a75cf4af8922bdc7ccef7dac71b84eb1ec49
zde9c771cb8ee424cbfd5a535e3d2b4018466efa9c8953de759470aae6488ba48763b64a7780fa1
z4ad817f1c3151fc5b16855cd08a528ae6aa284328f5eece7719567703e257d41ab9c3b65306e57
zd03ecc7df5118d557a252329e4301aceeccb675b13bf92c721ba7d37d7aee417d4476d7f8f76e2
z9c2a8b27d571cb3a23b28e720ea27a98646ee04d0260f8618bde7312872dfc5d53f1b063828462
z88967aee41e6e817c0acaeee3b00c6f139e9971ae8c6dd3f3de961d61552293337b6d0ead949fb
z768fab4ef38f0f0881c51028daef7ea286c3c8c8755998b789f70c5c9a86c21ee89b5e06717f0c
ze303ee8503ce4aa6280c4af7a0645cdd053311f7178c04c38cb5dcdb519370dcfbfe5b85bbcdc7
z769364e046341424a89a3c58691d5bb547adb74454aa13d21fcd3c065d2a62d0882c02c7449098
zec73b94d3f80fa3aa05a8d57115611b80a3d0f0b606fe0939b626d0e6229b48d44c76ba7ed8c99
zd4342d7d5aa12a9f51f2555bbfd93c28e6c06992bee2d04ddf04a54aedd1b90c3978d765160c0b
zd82352edd38daaa92063aa2011bdd94ed3fd4c7d9ed5833fc86bd6cf080c9c799c08ff2fa3148b
z09a378bfea4a7ba8642a92fbaea1519dfd063d780003fbee8f0d7c1c412c8fc7ec2992db7fa692
z9a72587f26f9ea64cb6a7a871fadfb6e8d13737765763191251ad5fd580845c2c3e6c3e7e0be78
zd7d22b592fbf0d7e5ff52afb281344f8b7555cd2ef5fcaef92b458e3b46f94e36dc9d57b00e379
z4810b38becdb729a35bde1241085a2b3f6195add94147f3457266b63399cc92a43b2d81c90083f
z50a7bb76eb2e12f92e9320edd9f57daca1e1d44f79962de666a69b35af492e3ca9d9b7f0c4f5d5
zf705dfc7dd061acb8a920da8df7f8ef4f088f6579b8a55d0390f0741c572d88f5d9760c7ad1a75
zbf825fcab8e5616aa54084662f1645dc915485c577ee4875eccf4601fa294cf633e115b78b8faf
z167f85be9061ce0fdcd258452bfb026e28d5608435e0da2e7c5f4849115e911a06e21991d7dc37
zfb32c3abd6c3edfc30d635aba191fb908dc953dd8616fa41e829be4f6615841047e54625517373
z26b3048533be482ceb5271453c52762e2c4b1390d3d313ae7536887adb68a03b88c66f7a50492d
zd6f6637d060368828186cc0585d530692d40bebb10d4ceba9adb25db6eda331ca7d68a16b66468
z8da3d6bdf056cb2043437c431c35b710eae39f909f86c38d4b95818c6063a6cbf62571ca7c0cc8
z22a3459307030b106aba53ceff7a5720001493b8f4b4390a2d0a3b7046511a3b6742bc3ef9242c
z1e2b122e6a7227a4a9c80dee1537f87a1e0e2441d6936a22d11eda9e6d12bbaa9389d0b55a0fae
z5ac9b746d4ece4126c8e8a19b0a7f74c166d1bd9fa1a58fce2e81e460abda7ecfb5aeccc0d51f1
zdf0e6b5169ffb0a10b18ed39aacad4588c84627190fb8b982e32095a2f7e22c13a54703751f43d
z39e750cfb26fecdf5be58cbb89cb3b6ef84e175d148d8169ca55e11ce1ce2b54398d1b26218980
z40f5eba0d6b8e0732a70c0541259b183ffa70ac481ee5e8889ff63f676a68363715ef83b508c13
z18e163525b9c3c27f71a40a6e00317634a4ad6b44df5b6b3ee24552c5a482d3c0819090df7b136
z05e2212d96253bdba30f172ea6a2a9b582b8e7b992d064ff4d38e62e1c8fa3c93c8413ccbe5a0b
zbc6b64d894966e7a6c0cdfdc9818a2154f196c79dc42544970e930c249ca0b8f603307c7826ae9
zd849184a4848e96d37290162083d69fd8ff59f8f2f1a9c5942190b38646e9698a3ef0c9894018a
zfcb39a3f7db2a34ef881f66e6ef7c65d60e9fa4d49e04cd783a395111b71aeb611eec3a4156811
z4bdefa31f48df212fbd91e6f39fbcfa6a975e87645934a520ecb0670518afaf5a28342ce23aa98
zec60228161b23cae52545ba672b7edbb305d72743dd62a75d1509b265e484e31177e32faa9fd3a
z2c6ce838690151682d599215851e413a3c09a17e7bcc8649ca80481a59a29fdd91ca97923059c0
ze8202f2e2b7565bc3baae9f22f39f09df63fb83a6496f9fea2b19565de71ca1a09d6ec6d1d24ba
z06de9123b0c97f8a026d69e4b07c396dae7d58952bcfe23648476f39b8c16f625358202d7b244b
zf36697c3cf95d1089700e5dc0aa49d6cff16617b9acbccf7a18cd4c5c9d21952b018bbded812a5
z7c0fd9d51ccc241084fa6cb3fe7fa118d78946f5ae26b8b6b7b0af9880d1ebbd35a5776cf908be
z79e3735b4bc2b244c1e474475c1c3205c7ab9f9160dea7bdb8c10f29555891e237e99b62916f25
z03b36609d29bdf30b50bd8d554503b2324f064969715bb4d38a3288a4ec554c427fa2bf912275e
z0c7b847d9c391478d7120deea3e30c0c7d265997ff6083461d781d3904711f0285f2ca70d72611
z094a1d59eb5a4e6b9d782b8a0a03062946460cd9889d76b8d96a4076c628827a0a01b599f4f4f9
z55af39cd7d453705854391068b062f1fa08f3843f3c4466825f83a1cd357106f97374d9c87cea1
z8437331a57278c337db7a605a6c8e32aad459448941faddd8bd67c4e81ec6c92a41b92c09e0597
z73f38cab8d1c6a49412e712811c49dfaab6028e174f77cc2784f4284c5cd6b3892e589500fe19a
zaf367d738fc2ba5fb94651044e591d3cb26eddf12d19d57aca45106df21d8d9cce464da829e9ec
zdecbfcea9b290bd932acb6f88f620f5d0ea71a34fad88971e45906d0088f21fc94ebe715194e73
ze71cff685cd0e76394a7bc670e7ed812cc079fd55189453bcebc917d7731ebf7010c4e74e7de1f
zc9b946ba22630bedfa6266af6e364828684749bd258653bed51d6eab865adcbb073703e895e888
zc956dbfb466ac9167f5fff9afeba6b57290bd67baa51c299db90b6aa83106900b7f5301228555d
z9a6184b6b56fa42365152c3f965265d032419e5b13f2eb8527fbc2bdc9801e3d82c07d5b9de1e3
ze96a0574bf2106b554f5ad35f04b474a5d8ebcca5ab4d0f2bcca77dd6572150661797b1813f65b
z41517e1aab07da14bea7d7eb556e43c0d976f505131884159d8f6cfa8cb98a972dc3adfffb57a0
z87e1baaa5b8365470d64b710bbb082aeec05ffda71c329ba75155207eeccca0092306e47b406d7
zd497c9db8080dc99bb7559f3c477b51368c2cd8cc4ccf345b9da7715abcfc4cb8cc2f2f1235305
z6253f2ef984eb30ca8e2d799bdba4a67110a1b8be761b99598469084e9747ea9ffc061d7bb01d6
z7ab0978172a417ff9cd6b94a134e772a24f1e976b9f1e06957b6cdefee418fb3e12ffe08a762d2
zd436e0a8e45db2e867bd392d64318f38a5b23711c21fcd3af5dcc30c3ea0d0555fd2fd0dfc8a2c
z4838125f41d6fa668d3487998e4567d75846ac50b14eadadcba67ac9e9a5281cb2975d40efc87e
z0e51587077cd75eb710c54ccd70fdab905e858f56264aeb900293d56d822e801ceeda21b26028b
z140e3d546529e94eb783dd5940c017fffcae9a42a52406331bb082d02819e99da25813e819ee53
z1de4f65d6f04b7d59a563a3db87ed9f92cfa62138ec8226d25629b09a69bcfd9fed2d50295a0c0
z4e6da14692cfcf90a950b4cc68a25af35e5e74646a16e0f747cb6e26cae52415b6b110b5a10a0b
zf4b0d110ca424e6070644cdcc2970c2a71eed6e047f48115412efed296bbced959b6cb2224ff64
z29ac4eec47ba11dd65263b13f11ddde26eaf22c862f3aafd3e2920b60659b76d44e59592549b29
zee9f35aea87b05225d2cc9008683e15d3961892d787c8b3e6baa23708232cd54baaa2af8967e2b
z590c102496a5e028181df8770d84a08615f0e7a823902720ce8c859dbe1fe5e3ff44eb87d47b5c
z7b02145ab44f6d0551536c515d645ffd1308bdd2c75d3884d656b8b3ec0a7e1fee6f86166f02fe
z0cc6647e6b62d8524cb3cc1b35bfbceb66d292b698e5872e94d03bcc0df9a6d53349fcc6e33966
z4e5e71fb646d5d26d3cfc63f6ebca27dc2727b85e8757a83171975873395081cab922fe689b65f
z2ebc05eb58fbaa64ab6156c732378588a53c45fb98b3dc2667c7c835190cdd2372e56255426a48
zeb9eb7478f524f5a22ce3e4a595e69467e5266987f5c6f6ce9fca158ed13548c9ab47113e7fca2
zb658f249a7b2e8f0328a048fb67d53ec18208604f52033ce6af5438cd3887845672c49ca73d481
ze1042f18764b54e7c758da98abcd8977bbf56e81dcc993df0814220576dd25ae0abfd9c1b04f50
z480fb389820297f3406bbdd9b13b33d08bdcc09e08ed05d435fe0ab2dbdd3682e2c9bcbb181950
z0a15235c945916586f54f4abeae6918882c8ec96e472b95c7497f9e87d89abc7d1bb66253ab074
ze1d91ffcc21c23cf8045685a52b315dfb3e59283fbce5b584dfaf4a67a8b16b884c100342c6002
z050a8313c06b77a8c454ca7896b17f9b03ffdeee819413441c0e5104528f98e32d1f792551073a
z30720629689cea75a78b5afc37f56a34c440a068e699bdb4f7323b07afe538b75b5a0513aba870
zeab258ab248e3ed98d9f5b09845970a3275a33a4b3c89a66bf850b7c186602b095dee55195b532
zba3db5cbaa230e3157fcc50af475f4f492d05b1c76c59d76544381475f7edbbeb0b729ff5327b3
z07512779d9537df6b5090fc0881fbb85f5e6211fe899e3ffb4ec6871ccb6dd8b0b5ca540082e05
zfac6213dbe56077e576c4917255ad45380a7937e28e64f4f2ffe8a088a46215e603c9df1d9822e
z76cf3cc9e0a42624b9be5cfca4704eaf4563f334c7e914188a2fddbde524179c7a94fa3caafc04
z6e3e0af43a720dd61e1e14f399e6fa15eee294fec9d7649ff33894b96a70c6e2b41ed39b5e51bd
zb775d6f2ce61c9c27d3293b7bcda518e7f2733a6b90702f0097888e3984eb536e9808043134c40
z0039ca6e00998309e705a9555d146805236e277b5df4536758a46c34ff389ad03ffba231740ea4
zc4728dd73b8ba8227c5e615ad099d3ea60384b9d70717f9d8c8cefb907fb68382253a43338238a
ze781f1f2039dd86f6a367197962023967070d08c3bc8ff20b384eae4cfba9fa8e728116a8070f0
ze1eaad9820d2fda75367b066327a28eed1442bb610dc8147d242a12042ed5d6e03c2ae4393f3aa
zf7a5ef56eda598d1eceb59129ae8613541c2f658252da5070f73032ea7c060959dfb388ceb8f90
zff432354ad6bc8cbc4604b8beee8955e5d967316824bae59960425739f6ce3249971ed549b557e
z2b50601cdfc666c517d6aa05824e3598f93eda3865e9d7aa98bc98765fdb17084cd0f1b43cfbea
z0149fd966caad2a5fe51a0fea1a92bd71d098f8b62fde4664a026d9f1024cf3143bca7bf096b3d
zb2c5f2bad3e62e41919e95213aca68c9ef3313c09eb8f6729fbbd7f96a2f732335c69ff7891f67
zc5621a1b449106820d068233da3e7ba430d328f7eb084f8134c121bfe476ce7d30047e2e328731
z90cc4833485e7b63aff4b97364cc9f31f79c431f6b04e30f2517a941e0ec7a5b79e1d0c3dae0ef
z62f4d54027c52589ade48e7ca7dc76554209a705d5a0bd3f64cbc05ee2a17cb3c3a4a0984041db
z3cd797decadbfef0b813638a6e2068d9c023ef76f1e437a2dbfaf34de7dbdc8965e5a998baf199
z9141c88a39acb98b3ff40011ac179be4100ea610bd728f025e34016a84b2232d5fd5445de84cd0
z23a5d36d99307f9633b356be382a7d0dc3072bee39c153a913f3d7ead6139efb12f468e0591d46
z0569184c0d294a7824db0d3129a300de5583f8a23c1fe86f8270880e17c7f71908434097259415
z2245072d115c6810f7dfe032ade7275327c777bc929b4bccebe87ab5b3e323b9a16e2ab509635b
zed16b2c4973bd3020cccb959f6ecc065e10e5c387ae6aa42489d1702ed6526e98131d53e45e772
z7c1d54215e7f83b130ae2a0a5accc17075507c56ef56ed3da37840ce9ad7582782f0354844323d
z2e2d281f4ab6fe0e7c5f20fce4f56aa6aa05a5922ee3150c7758bf089bf31186be4569ae00e238
ze2b272ecaf03b1655c09927c638f6a567a99f0417d54c4e542c0a4c83cd304049e225a36c12d88
z42d797645c9d03393c86d25e80e382c4731d40437ad2dfade2fcea5e4825e57ba532e9d7230cfb
za809a380741eb9b0f052760cc20d19ccb7fb3616ca77ed0c621f2391df394904e162c5108f9f6e
z5f844866f469cfc23532ec4fa480ec56672945b8ac88f9ee826d87aa98bece47d081901fb55a79
z73a74c942755ba76d157b249f3ab0704d962ab15a4b65b20c8364496026e8105ea9f54b887827a
z5d66c730667a52674794cb65137f73a7d840d3bcbd8ce1c3b39f97b8263d4c31fa7ec00368e8c2
z21557ab4327e50871f9588ade57c8aa421dbfa127a96425f30ff8a021fbe2f2ed96acf2513091d
zc8a8ead3c5ada243debe588e77bcbb9728df8377b2a9aa70d8b7fd87d8cd4caf6706d1d0c578a9
z296a886b28c3479b34f982a2135cc1b57b62b6bf995035de6388fb76e4e93b46ea432385d6c07b
z0d50b5665c3bc3a516c51c746c7d9a79a684ca5ee39bb4b424fae3d96bd5b5562afabc94620410
z10e29eba8ac6f8af0956bc3c8c997bad7179876b2b0aeb5a0ddccefbe543205fb3c1cb6a58430c
z18917854100b4183ed5c233e7a3e2a0591b3ddc046747530a23ed026a8b02af67cfd5e07db1997
z23b531856eb2f8ef04a4618448be625a010dc1d88f41bcf09706bdab0c6bc88948fe629cb877c0
z66e412cca688cb1cba679286be8957865800427cae6b39881c2764a1ff3f9b730bdc71ac6fb0fe
z31a6abc076c6853db2e64cfdc0ba938d08e7f1ebb489ce4fb29228465b7dba02e1c7b67ea9e8f2
z8e45459a642756725bae123edcc316f6abe6b4dce36e7a154fe4942c1969a759940d8a919d383d
z8ae2afa2cad00b7dac022959b3cebf9fac459854dd9f89c58d472f96577646d9cd20e71b1d180a
z1fa349ef79837dec1fb46a9e5a34926474f1d5b2c631cc8b778105a7f9b93ca8aec572ab0c3681
zd964dea1116bbe8caa9415c1119e21c12b86bd6476cd76965f6567a0385823f5aaa547f954bfa8
ze90d985e037f0c5603f974cafb0c7073c9149a041cb027695748acc159a273caf951764a40d9b0
zddcc4501ba254bb590225c597883c5b3d7164cc68d8ecfac782c659f8fe18965f8703ab8ab9d52
z29cab611d8610a6c54cab4d246e5a1837ba87cb3722e8a26d6a3d61b0ed31e7476a9d4a6f4780b
z7b8c9734f8202b05357948fa9a2d86a63600ba3bde059658701f6a51e34bfed6987b6f455a111a
z72da95a471c9688047cc0229765e325ab2ac8bea578ba5b57308bae558ab8f9e4777d172271e3e
z4033e6bdce9cdc0b4c8199d249e2e5a6822dafb23fbd3596b5fd8ba5857f0d29fd601c6cb022b7
z06c5fbb045c0521973e283a14a4b23d1617c4c56a776c9862f004c568254b36dd719c51459f8ca
z7b2e87a822f7d3e5e7b6daa1360f858e77f62193ef625f20675a023bb4f9e62de7ad40c3513d9e
zd1352ed4277f91e47a9780455ddd25a65c503900f863659f7613ca623e4132565d8059468fed6e
z629065b416a1d6fb5256f967b1bc45bb31dcfb650596ff50e34a871e144b1cc83c6edd75eeaaa8
z4d5354da77c903e7295773337e3b69df809861c69e6033c030a59944ca25fc9a293b376c68b933
z9a5537d31ad8dcfd10c6bfd080538a13fa5e22c6eb86e71dee9b6ff4a111466bc83e6e044b13f7
zc7b2113b485b2d209e7140049819d8cb202bdb8c5d72c605b920f2227fc759c3660f659edc90e1
zbf6a47096edd4884fcf498d913e270769b54c505522d03edf4844fa16b06edd7d64d27e55fa008
z44f6318c0fcba3a8973f6cd32dbf8ff8e803eba5a7237f4a752f75402d20513d8b0dbd875cfedb
z6336fe3f4e58e1c07c9467106559bef2c91777f1d001e09f340327e3abe339793be10023fc2ce2
zf8f4c24aff3f9b4ffa9eec09d186203e212b86ec09766346912d49586b419c9ecda236e62cd941
z85f28515f89b2099174fdd5dfe41cc4e83d91231375244458a419d53603c769feb57cc313dacaa
za15328efb4464d26fe6a7922f53f91c421846c84d771c4956ba2d935f51751baf7cd70a5af3ee2
z2e6228230a59a0f8dc6538e1a65f83628b16ff7904b4f999df40c402d176693c09aeede58ed44d
z7961d34619f0c10804146b61b6a771860f7f5c88c8e501ae68464cce153fa94d97b3b5c4c44ed7
z0f2f849ac296972b10f09ee225fb46d018be789e9ced257d9c59b59d8193dd5acf5b214d4d3b62
z84ac401f70d1e4de0de6ee4a9b936dcdca9dc1d9b91ef922843d0c5530979ab5698864356b4c86
z31dcfb386e0a0c410e3290e4c865f07ca7ae2447ff6ddd2d14efa531181872ef65c8e44f74605d
z0c83e0041e135d33c37d6c01e510c03bfed36693128e264a9f5e3c644d8cbc744f2e2fa857050f
zb951968ae75fa48b7a880c1ca5caef355b43527a5de603751991dec74d807697324d43e2b6f639
z83843dbe7b4351b1272f6d8a83a7ba6db10542df6a553ba0642f9fb218ddb64da565939937c111
zb9017717581848e1ad2a440ae48796f96bd07a28b7ee17deb1474fc9fabd56bfb5e613501f5fe6
z7a1a72b3b230d6c2841340c8ee07862c29e2aeaeecfafbf273cfd9fff4a268d5aa5009a9728b13
zb6b8d7191bc0bb135d74c5f741ef4272be1285267b6e11ef764aead26c32bac81a4e83e9e003b8
z2f9730c7f13fd2311f7b07529681fa6657ff2b9f30b903fe743e7d5bb3b231cfdf09aa96f04b9b
z0dca21f32e3a457f54faeb5d1dd894f61134f8d5bba82862583ee4147d650e9ebcfa992465dd46
zff1e7ee0796ef2a16cb3b83e0b44aad2a18379c9fdcf1d28bb942a7b4f4704ff831269f1f7a253
zdfdff11b8fc9840d70ae5c7d631231f92bf261fd59904ddc81a2325bb8aabb2310336fd8b28e8b
z9ced68f176a666ebd8a78860d3faf68ebbbfd184558c880dbc5680971490e844e9fd28b5e1030a
zc65141194c88c480dfd348d6ce411c93e0efa903eef201851eb91e411f02dd7fb798d26a6dbf2e
z268a5b068a11b642ef76691cd23c070f07f0126b36e0d7b6661b8e7f6c532a16fedd38def3a401
z11bb026a40d9e14c6f532ceca1b8092ef07af85e319a33e8f06fa9723d8364e12a990e54fb3700
z83fcc85a648d7c37ab6de888f888847fbede595d34bb2263cfc3475e83b4ca7debd14ffb4f2ab4
za68203e86777febac9cf54ed2730d53f23180daeab54e98c2f0a8a46ae9d82bfb18891535ff6ac
z42f45f04bd2bb64efb1aa3a08da5a90b3f87bdd48a33f2d3f32f25588884b84f402e1cd4be852a
z383df66f01ed01a61c8b2bd4998681cbe6d4c3dc8aa04c580e992c19725d438ddafff0249ce91b
zaff68be77a6f1a444bf5d4cb2e9ac4f94dcc3546d240a6b5c29f809aaea1798d284204c501f086
z63e43ad7bbacb413ab9f336415afe8d34e08e3033bd5f15859c3f770bc24c31700885a49aee57c
z02d8fa345ba4c5f5bd59a0f2ae6e05b5877b5a7d8c39989c243c97a48ed11d9775876e834c629f
z5a5ff39840a1a5ac52dc8596cad24c5b63ecbb019c601e87fb2150574bb8cc7f5c7ed1507d1800
z27c7c7667ca73e282f4388993a30141b13258206e54d302767c4795d11ecbd3e835c0b8cd9633c
z4d0c403ba475c6828fc8dfab631c009287a5fcf04f7de5a0395d6615af14a75599e1dd7568d930
zb4b6ea7b19a10294bc0741222deccc922563a8b8d5ba551480117534a98789786b258c69bf4cad
z889ce692ee59e8b93e552922cbc1fc71b2dd56fe776f07fee97de88a5e1f0249e11348daead352
z1ddac69ca76fdef88ec40fc3560bbda38f1910913ff822dd2ca92c68f5b40b2e9191d6047c0075
z89444d68f2fcb94a0419d950679ea240d52737cd13a3c703cb17de19601e4df369c8bd0d0f9b4e
z8423cf7bf93a684f90d6c5dfcdd492bddb68547688ad2a138e7f30764b5cc971e1a689cc942fc6
z00909194bc5721f74e917d04f135508a4df0b62caf2af5f985df4544eaf20a1023940b3c632054
zbd2cdc9450e355c2d420ba04caa24207992a05dabf114b5a061cf6dafd51476d1778d2afe76359
z168e3c48d2ed8a29d3b8be505828d23351dcaf12d825cca29c964336d07403a39d3662038d4196
zfa42dbb46d81bfd6d366f9b4cacd71a9c208d800b85974f11a667335bb857166ae1ae31f12686a
z29cc5457be93b01ea0499eb5f62c3ea060b645a42579f787e52b798eeccc4d6dcb8a7ab2580a56
z1695affc5b343790c8b01a7d5e8d0f4ab2b1b196e044b06aebe7f3bea217d857ad18641e7ee16f
z184c07d368d625c3b911da75b5b2178a0d69f9b4146ab1467d76a3cd337a7c4b59f7e44e2d5dfe
zf778ed2d0223949f81249cc9b5152c52ec1246d23819bd9ac1ce9d56a8a50c5f96acdbfceadc0b
z3b4b4c0c3ac3c80ef2cadbdfd34a5670e707c7c051ab19edffc01d222179cdc27b37767ce21337
z20f1c65a46dca7b7765af1d6498a5e246d68b3878a36f5028b88ec6a3bcc811fbb761a60397081
z48d79220897a200bd3bfa0b46021600d64c352944b5757a9cc19ca5b7cb0e2e058931be3b304f8
z55dbd095616f8658402b1283166b0ec7f2fb27eaf847eced4d50c27155ccf7d69b8c91c0951cc6
z966c54e1ab0dc6ee7b019b8cce98ef1169318264ac1a4c777ba387d4b15f3ffdf8481a7f548f3a
z3a79e3bf77ab3d89f6193f548ffbc7568d0cea2f4a155380e10dce6c5905a0beb8a0c650063a83
z30262075fcca6230bcb6293fe27f7664b36f29e1b2cc76db71b326bef2e0e76bb1b0d8bcad757f
z7dbf756d05a48c43d1f8264cfe51892bb75cf6c9f2d1e8ae07a3c63c4d38d2a37a9273f96c7cc3
za671bffc99120d8b75fcdd2d40b0b99d0dbc82f67111bca15af98fd3a01b4933ce55b3117e57da
z7737294455174410469caaad6cb876a1b07d65b932e4d543e45a9c5eedadc71766d9a023ee63a5
zf423430a6a8a38147d3fcbccffb565b6f5fc9156a4342ab9a910c79e8d9e525c12ab1fbadf23d0
z07eb7c314832957c61573bc91b806e36bf8fc95e53fa51b0069a3e9cef6584018e9efcc9c2535d
zc97f7419e620359bdea03d61616b682f0cf0e752e88835a54d4bac19c13f5fbfc61b497fec4c1e
zba2ca9e576c054ce255f3d7dc912293c7246e26442307c4a5461b746729bfb0de43ef464777e78
z6b7d831a6306b5ac6c1816cae18c8c52a0ef2a1fc6383a5da68adc777bcaedbde54b2a057c0e3d
zbd768908dfafa1b42dead4e2560f57ab2c31594c1bb376c53a0e7b5f00c983934070dd37adf414
zebac429d1a46d1a3dfabd184a69483710d2f9a29360a37b2cb6ee8bb5e19597bcf1686a00c5fd7
z7987204fc77c8cf19e8499c7aef8b26bd4bb3331092d72256b610ad76d041d42ff855179f7afa5
z48c4f17a8f8b5f6d4c782f8e27b04c68d3f29b8280fb2fe69bbec9f54ef2f79a05322431f5d6f3
zeaea925f6754747a2cd5807c2ad73a9f73fbb2a0267f8b01072ae1933e6d2d353bab04c89cccac
z49899fb12dc88cf7fcc9787625a8c164013797e8e8deca9a2fa47eb95a084fcefa81b74a3089af
z394b4e07788383f56ac01f939d627f50d340734a33e85c656a0244af9818e8829cccf43c584be6
z4c4b483e0d6ce004655f935b96b0ea4dccaf4287b87bb286be11a56dd5a9a11b368919d7e07ccf
z355a0716d3356160bb9a3057346688483db6da0899cbefaf637cbc51a8fe9209abccfc404a47fa
z308cde397a5ad2290d136c20118452879177a6926be9b8fcaacf6464371061138f03132285bace
z8756c120ec0ce96263b9d1bd15e6a394c07b7ce275af14dd0abd4ebe607a2801b262315b6ae811
z349f8a1738138cf63c509c5522438f4d553c68fcdd0628ff1e1a35cdc048e43c748ff2f64f7c47
z1f39bea0b3cce7b55d737b0fb06a219f6e5329737bc37dce66e5d1e09729304760abff792d659d
z77a68a13615dcf04dae1bf5b384aa755cb9fa48e346de3c71cd75bd9b0adb1674891301bf09bf1
ze89431d5cadb630d2fc9e0cb4b97f8ca6828e35271ea47a2edefb541c6b48bf79c5fb7fc65722e
zcb18304fe3cfe3fb437d9acc32d8c3b00acb29cce123c0aea7755b719a94a42b22164fa3644683
zd24a3be13cf0e66590723c10861dc665a9864837f64ee680aa4e1fbcc99fafb68b115d37fec24f
zba47240b8814b10e52bc3a749b57f341107c1aaf5abd52acc8d05512cfc07dd1a186282c2d9499
z1d64c021e4d50decd7df9f1f8ace6e30dccab1f835a44077132d372cd62084f4b2638354bd7e14
z2f13b6a39a9c492944978ac09cd05054120280e28abc9202414dbc68aec7a100e56c1f930afe33
zc73767404facd089540ec89e7946b0fa692f8dd6a1f179373eb29515f34a92f3a09a590ede36c6
zbe6601658e1fc9418023623bd7b2cdfda79b2a4c2b7b97c0e7a764d107aa77ac0eafbf321d66b0
z63a244dc5b27979ba0ed3ab8dbc79f6b99587e34aa576c82b847131fb6ada2c31307dd26b46cb2
z73cfe5b0438bdaf2aae027bc10b93d75249e16d6f94f3850325ce4fc55ba4c1bbf27ef561de665
z57c72cb66ad402451d873f6a09d9a3438484109c5d45353da4741096487e5703a0cf6c1e26cbc5
zd823cd24c0a0c371d1754d1cbe3cf9ad17cd77e375f5a76a136351348343017761ef46ad8594e0
z105481a018c39a7c7d7ed71a898c245261a0ff33eebae94921a9d3210a7c063497bc274c3861dc
z5c51349fb21a2849ecf8c06c58363e422743037cf277247ced92e2562aacd1c88199125c8b119c
zaf6db674dd5acdd4e73e163e89f16d8f62b4c01d592e2b984dfe2459d03bd63c1e4fd9ee9c4720
z100531612620ce7825548b2dcc28643c7daf486e503b893a457db4d83daf7e2f8dcd12199aeae7
zfb9d71bc112210bc2dc8e4c1a59760778671627e4d358deaedac0d0eae251a0999e6c5ecd078df
z3fb29454cc0f6ae09b70ddf61931ccc2b2b51f635375f0587af80d5c29d7c2bd0a8835749aeea7
z096f4cdaea5cce40e62485fd3410b1d302b7f1422372a383743c06a3d0f6b65c625b202e835d2e
za438ef7c9350efdc85deaf7505eaa7948aa0cfe51b63d30b395750815142d586877fdbe9dcd4f2
z3192273acc067821d820930d17686bd7673b4c235f2c8311d41b7ca4217766f80744b9938a87fd
z92c5ee531ab416a54baa7579e4d34cfb01d2aa7267ce84e58565d09bdcc9e8d6fbf7d8f118d2fa
zb920c33023a89143851a9703ecc6f9b91c6f0defc9cd63296fbf8b2eb26923a20d1aa140e0a45e
z20dff08cf6f3273cfffa0a626b63d4409f3f97ffc8235e42086391c562789a4add04dc55848b3c
z26d366d37d1870ba71ececfc29670742b06f78a0aeb0bfabbc7edcaf10f27abd0c758c6a89c841
ze65bbea3dbd586a3f55a717923eb16673fa8914d69d660c6136a9746e764aef298cb1d0ddf633e
zf0e1bc8359ade87465cd1e4f8222d511c3840a865b9a8e78fb621dfa7b9b0d0f7510512362ee05
zfe39a8c4a360fa9d53c671a3171784f61f8ff5eca91c1e4fdf6a5d675fa73cd99059c4b4e2dcf5
z29cac9cab69ec4fee1b87214cfc5741e06f7ae474575e0ed5ec315e5cfc6c0c01c9f0578b47d45
z236276d0afd7c3c4beebd8bc250fe471fcc28f5962c862d2d281368ea3c88fba8b84107bf9b249
z91f4a21a26c59e804fd0c9fded1150113be5a2a7caf51590a52dce66fc310363d98601194e5536
ze03447ce82d9da47b8f5ee0843f5b159118f3f81ba0b5e2324c8d55af48f59c69e9dacdc91e04f
z6247fcb18abd196553bda4bcf07c0b3548215a9965d00a8e4d4e1e4ab01e93c7c195fd54caab93
z16b06e896addd8dd1a4cff7dc181ef92278d793729b0a4f27e86a18e7c1e65b786bae84c7122df
z9a39db6659fcfc4ffb2e039ec77390416e7be985d8d6931516b4d61362cf9b4db4864dec28de77
z9f8e31fd5f17203c06ff43001a1153308ba8a3fcb13fa5700d723866d54e69f32b887c85f48ffa
z3298aded3289eeed85f04f970a60da2d4b5f8a352ee57bd0ed25b66a45cca5cff45c7a6ab88251
z3eb4ef5a9ffc1b132065c76faddacb96c6308187d308d206d8267f0e467b2b91fa36b21c15abb0
z757084a5052d298304bc62f941d8132790f21e369436ca043261912d62aae16f5279ce6205c995
z790dd2c3b384ffb92ff6bcfb3e716cbfda21e9fd923a8003d59747755272ee672cc9a7cf97dafe
z73666aa5e2260050079245bb250d18922d356bbb2d4a11c9e0093b33b3e7aba9ab27b88b6c9e22
z15a76512dc4fd9025345721015fb15ed645bef5f53b044a5526d5c2071a3e0732bf5eb3e4fbff0
z5ebd19f4812390fc721056b377730143bbef50dcdaaaa9dd0a94c1b9ae5b767df1b2e9caba008f
z2f0c8349615c69ba119f6cf6897fbefd5a260923a192b243734d873680b7eeb66d9af3a9ae6d9e
z80480d0f533c9998f8a184e12e8a52e5181a0853127873db0651159de50c6e740171671a2352e1
z429373090ca1c5c3bb2d9610d174dcd3e4f30e29f9d63cd639208d4f55d9a7a8e4a434c2781cf4
z9fbd6b8e73357f6ae1bd34777d56a47ceabe40b3d75d3cbb70a1fca9ed8c96b3223da77e2dd1cc
z85da1fb3e87fe3b328b82298bbbaea249a0c935036c706c852f5e8727772542df32000a6325efd
zd11a29b1f5a52b2dece15628658b86e3615e7ec5e3194f62106e31d6985b9993c3e87678301bbd
z6e3fbe1ece2d4b5d5119d37394c04bef4e82729369d149c3ac14157f2d77cb3558f09e3e48da05
zb32c4efcabd093fdc4742f0a24d8590709f3789c941dca243c84a6706abc76a11a5de7639745e0
z01cc7d57aad9d4bedc02ffc9a32609e7b77348e3806938b9c3602419a38306605bd4c04424c311
z48b83c8d7d3bfcca6ede5d720df7c7f3b128614b1ec56bb603cb8a1831de18a5614a885645fb98
zece2a11a30dcae236c24f511c7f42a18fc3da7e4bd528ba78d57a4a116a4d5cc9a7794ed3af683
ze377345e3f8dba4d93b15d24600fe4bcda051875439eeb8db5b5de1f5efed5ccd1199292c951f5
za289ae01106df76e6faf3de6c1181b2b9710cb2f39ec39e6a10d8d4a319f6c8286c0ce1456ea6d
zeab5edfc78c44183a97ec17c808edcb358096f89eb85233971dbb3ae497836439ed08a30ed6025
z36d26651dd3c974d8cf211a47c05d93ba36dad8c4b21117ebb20da1a00cf4d3767af6685fb1b13
z4b4d446bcc68948cb3e7941b66fde5bbf3c93a9d4ed804d2e8126c8398c1f89f373a382880fce1
za9eba08e0e32a0c1ac5c40da9ccd77fe4d2b5edd6af0b7190305a464770eb9c307b73d40045aa2
z039db0ca0c212f7fceb55267749e36da8dd276acae2fa291f909fc268d59f1fe99c5675270a0dd
z1b6e88047cee365e0b242fe404793fb79476cfef088e1b1c6516d8b258af307f095ad6979b1889
z4f215342f9628da2b8e42bfbf673bb4cffeb14a2572746c87c208bff2e839eaf009367bc46a073
z48a8e28e92e12f6f9c214a6fc8558c559da9a2c8bddbb72f18f1b0c8ec5315dec4a3a9cc411e2b
z89a803fcf1191991c62527d6318231d8b2977491a439b29f6e326c8e15c463a044ff9434ca5b47
za6dace5c8a8fabf04e4f25214552a45dcf24fc233067695cf96835e2d0ed41d74c51d868fa106a
z47083782b8c16b44d7d8b37695ef0b010cba1d8f92b759f1b58c345ce3cdc1d3eaa770fb298d0a
z1907cde4c51fbe400599f4ccda889f962d96e94aa6bf5bbbbb164724e6ec5bfdc715ff756e847e
z8cdc754968883d72e2ea2c926084771b6aae74885b704c71c4ffb61f8439407568e047f9c52b3e
zf40dc50a5a0d99d61816edbf762bf5218bd7a217fdab2d367d93177981297e7c9cf3b85e2b6147
zac340295818621d4a59e0192292862572d6edb6f37d129c6c8c40faa6cf1d4408d6bed002404f0
z242188d0b18a8e0cab355ea7414e05f138e951edf795d3d010aaeb66cb5258bb659caeae9732b1
z1bca6999969caf8860942192dddb774146b9e13e494637fd530d2b15dddaca211e3b301c9a9048
zbedb60328781d6180f84b502547eb2254a8e7f760610b0bbf2219971965cf4f8fc015fd918ce6e
z6756448dcaf6c6c8397e35d1e3529f7a324d7db4856d8e24a5b35e749113c584f34eb02d037e6a
z1442a7b65a38b1ffea696951500561fd796cfb15955517c467a0dd921634ad7e7fe531e9cda396
z28e5c731555a056134eba99a80f011f3ee342196d79596bb368eacc0753a80889ff40a47c447c9
zf8bb26ef09a536948b6c1a1bac2e6999eec199268e54b4867a7de2b64225df86d2f7cbda1dfc6e
z7434c2f93b165f2afbfe4f7e3bc4ad80a1e30febd1632d86aaaa39158a1a9df4d1e428ae18164e
ze0706687eb1312c10aeda6704d29f23134b0515cf8c9dd6e56976d28ead40e0f321d2fd73efeaa
z0bc70b18669356f0a22678f26bd0393be93b11d9fd3fcf230491475add3188c7873bb2091be739
z5b9181146b349c352c5d277f491b7c9ea58d84297c48d7517cb990c7181b6d63270f4baa0495b3
zfe829980c2d32144269c5b48b15ab0a8541ffc56586426eff5c9c3661c4b79225d7986a173df1e
zf5d05dae5241ad4f5a30aedc87fb6a94607d2fa54e24548c4d2dd8443d9493b2c09c5b12fe595b
z94ec0b01e818d975a2c5f2f78b9275b46002ba3059e64622ea18d14e2723f5ca444554737bf228
ze138738aae746e3cdfa8849dc01ce0573a50314423fc197cc03008b08af66d9937e36ee9ab6357
z985c8f821e8ccbf82490af10b73913f718b37cf98a70660884c8fcce827ab506f88d1775735094
zff7d0175e1493e0ca00c5864d46988e80b481568bd19306e7e006d4e5f51ee4b92f00cb254b293
z0c904ff7434e9d081d3dbccf41501571aefedb466b3429380905fc73e0c846d38a3d5b2724c488
zfb081b9648d6c62c724049cc98345a836b5c68116db0a86916dfbd3d9a931c4b4d5aa88424a78c
z6a5b2875e6564c661e8df85b914d9bb5a729c04a4141fa5b0dd4d90103aa14e09f5d00c6b023ab
z2c844898406cf3c78c9ac46c178f703e24d2bfcb97f75a8a63f3ba4710105fb0417cfff777c97c
z6d15d5f59a93b66016a52bb21de70e5519d17abde8d17c8fea9aff3e55fabfadf21a44d21d879b
ze7372c16208e4c7db2201e12421343d8ef63da9d2a0f501df4c3e9f8d64fc540499bcdb903c749
z926ece276523d90f23feb904c7ef5309e3b2c7fcf70c3d919aa2cfcb9ef368e78ab2d1669af5b9
z77e2c3d0fd4883e3d641a75569961b760c0a86a661c5dc6bc2a1deeac706ddee2f792fadf27417
za4595b3f56765b694b18ddc9f818319c7dd8b50915038740e4b17755480d253d57ac3e786822df
z8d774b3daaa6b3802471a7a8af2aa8c8ff78812fb80df6539ac2066d130c107d727e8aa7f9502d
zb6a354d4b47e6d593d03751dc603af45a4b33a51d274ba1db417279f8830c76596a153ee85fc46
zf6f1b5ec7797cbd4c1264d6d48846feb6b1d1c3d078e305355c06b00b11a4dc50730c6f08be117
z7317769587ecaa5b4a0b9edc6226ed30616bf056f9cefeb60f20cf89ca801630e610373e93c28d
zef9ac33c6f3dea9bdd6ab14a8ab14ca41e49655da14867e45cfe4ad259fd32bf67f3679a2c5ce5
z901301cb969e9813247858910df107b7e1b64e12ff5af3abf517476e5bbfbe764e8a5ba04f1278
z60933883d9e4792b145b3224f9da8ebd644660711eb5630364ee7a7c18f27b85b4ace25341ed29
ze545d62601c5c2ca369e143ab2324752e72385da7037dbb09dbc159bd062562d256ca624859e3b
z049002818fcc2840e13affcd505779e92c5133034b5d2fcdcacb17526d42fea1446abc0bb1b0f3
z0fc499a0284453ef247ad709dce045ed5647c541eff2d6510ed258320ea02940f41cfdafd4003a
z658579b4793db26a76687a4806d450475b7eca5c6e81960bf1e21a39e14bafc164ce2719579692
z7614b5c2e9d97d032048dcbb37bb7f4825ac68b479a949fd6e166a1ce323ec9a6876949606331f
zc25e9451e5d69e8a3bbd28d47bfa6e5ef9c254a0bacaa3f7d9d1251abc1f5d7fb1abbf2c367297
zf3b0e3e34905415ab11bbf70f6386f1e7122d09d5b3549169ae52e33239b48976c695a61b7ffb8
zfb01032d38a07fbb56cd7cf55e2615f65fb585732dfa71dad3b60a96126dd2e2db03161eb89bbb
z4d19fdf969056967c47a45596d648a09eca8093e065f5785b6ae0436d61088301d0b0986d47e36
z74fb1c33cda0899cd11611ad357865b076b72093105520db5a7359f41cba4db156f21579b3c174
zb71130e92331580b0b0ade7d46e51dd6641c841d73e18f22ec2ca01b5953fe80544e9cd5bf1956
z7dfef616f7b63df5623b445eee25ccc7fb716763bf10baaed15254cfabef7b6c608b41055e79da
z02545df76eaf03568d947e8f1d0bc8ae99837be5936345bc22b29a2a72192593325d91c7f1cf9a
zedab55fceae6a813f4dcdb2d1d738d782f810b35786d0e7f7d3e0b10677ac80434f94a308183df
z840d7741c6805ab33c18b4584cf610d37327c4dc48c5d2aea605c65b1a775148ce96325a92e73f
z1b004da27c6a53aa22c8436f5035413c00e9122d323fcd79ca3946c22999298d2390bcae663a34
z64899dea88f6ba0fe3e2ff70139f888e833246a7a02b1d10509cd97dfbb8557daa34602e8e0e40
ze411d140cd76cf57637b8605f62d65afc9d7da8eb11c7a1dee4f6ef0c480684318b54d1353a7c5
zcc29d0f005ab9b43d6996208fd60fccd591bd6c5348a212c5a78a31edc8daf30bb56a5689a683f
z1e2d79027cbe51857360090463710ae7a40d53dd0a8a27a6a07f86d4908c3aa97acab18876b589
z3986f90fdaeeea3627088914d753132497486463321c7e3ffe552c04b33be731331805fb18f5c4
z8d44cb78204efaac3ed5d13e4b2d1093432a5fe920b7aee5b5b8dc7676df30d29fbdf7d7f4b95e
z0ccb8da935222be0cae291a194ae0bba2acf1f87b236694fcd101a499273328694c020b7c9707f
z7faf87a5c64b99d4f8a2857d8d8a44fd730715bd049d2827e2a8e473d80d6db77ba70005baff42
zbbbbf5364a9ef3d86f68c6beaf9d5534a2145fe882415e163d96c53cfa6c235ce58f176c280349
z05b3961a682a548dde8dcf1549503d34424bc05e9daeba9d28221260f8b0ba0d77925e0311d6ad
za821c72da3b50bdd131e977acf2ef8025673e3e535b135f6c685b0771ead097928b3cb9c62ad1a
ze184b1affa66b3e1ce41c6463b65497b2df72a198010331a1f87f57cdd6649f2b2a6932c6d3c87
z03e324c927fc67939470edf5215421711087a24d3af51d5f412ca2fc4d4e33b4f5c89821c18493
z608968531bfb98399199e10b6f2726c385e5baa8611a85106c2abbc61c403a7de977401616255c
z8f3bc7612ca91bfed143ad3adebdb1b8f2cee283da5d61567bf17604f5bbd9b82f9783766f0ccc
z20f231b4345e0db0214bf9ecb012a135fa2186dd4cf9378eec9b262f7baedeada7fe697d917a4d
z6d526a7315c20df43ff91f50847bd84e38bea008a30a6b1c9d2b3dbd01576d2c5140aa44d65e98
z1b07b29767e1e17e989bf9d3b245ea8988eb203d9eee5958b9a891d55f6e9ae42780ea62c30b14
z83d178a739f9fabdbf3eaa30bb2ead9579682e5834e2f8520375b69315145856e42dcea709548e
z86823a99ae9e4223efb4ed9a1072da87a89f1ee5447bd0d5792b2001841da0cc8f9940b3e49377
z2ffaacf011ae08cdeb3b892adb10cdb04b8ba294120525aa946a7c4d2213a2823e1d257e8cf442
z259ad2a5ee58102e34ed45a7b19199eaddbf6b5fcc3d525e19f375e6afa775a1da0ba3caa60809
zf8492f9635c4ec201aff12a5d1887b3ca0d9f885e1621e2afe44d70fdba1c5d19d34d8c42ba07e
z8999d154823719670cafddbda0eaa461f971253973c5aea98c8dfd8ad0fac998daffd789207f9b
z1f51c9f17d81e86c328676691b219ff9edd1e94b8d7c9347b76b0643cb98c964049d22ffd363f0
zbaa5a4a9bf1eb59e0860a2fa1ee6d3a5f54437d3bc494294125eea8d5d9b0042ed698f6972058e
z872330a003717b261abeed2a5ee8af993af51f5a44923e70fb35c348e4551de34965cc3d244e93
zd7427aae5625f33569dfb73750f77ef1d6515068839776e550aab39cf5f276b7afd0162bd326ee
z066b0d30014b340db9ea65bdc774cdf5bfe419289f85d8b444b3b9313f2cedfc1ce534fdb010cc
zae7df21540acb3265cd75641fd2decf0e569a44e3793ba7ae6ba66c6c81a5240bedd1dfb06f212
z8a9cb8349d975765586be70b58945bdeec0c3e36d0e760aeaa2ef1f6ad71f127865f5f39413238
z095531eddad5ef89c5f8d840961c4eb389c1f5f4eba19fa2e6b23d3a3e2f6478a9bb5a14b3fbe5
z50bcd0e1d4e017c3ef9b856b9d519c5f3890bf2a4898d2a22656d9bdce9aefe34b1d2829aeb091
z2d27f1a80e35ff4c831c9aa8b55869974d4e46f92229374aeb015fe49e01dac1aa03b4d264deaa
z3af1273d4c8560cc3d68339f8efc626225d362c5ab08fa097e459fe82d3a2e7b8dfd14ab20f5af
z128075ee421927fb53a911d6a5481eb965a03489d64b9486eb4a5db77bb6fd379a368ddfdf85f9
z1a1809f380f16a0816e5f8f60102dbf32936967f67f3ae40025469415e90641d0253c653f5033c
z5bf5a9da3c1fd9c30caf4aae4a4439dc97d2999bb5321f46577232924fff983220174c680218f5
z22febdf1d570bc0e769982e99c78dfb8516269e4ea638da708d5a352d05dfbd5be931d529e633f
z69835b95127ee0c07ba8e53b1f7977e2f56e3ec4a8b0b0abb31de48e8c0c0801d175fc411d3249
z1ce7176d53295c623984995b720306a549e54c0e38a7d583e10e0c568fc4376ab5fcacf5925535
z95418a81b1076e27c352a22858ac85894f375c2cc9d3c061a5b410bce68b5b51d05069f37b79ca
zd89394942f6102ccbbfa57cb3659feea27d3ba38fd5aeaa0775fd773330919c212e4212067780d
z8e062d3741e5fab91b44e5965a9cf2b78b9df0e94b3fb98f5706381f84cdd1a629de6a6b49170b
zde39a720f5223294a32ff861d76c6a83fe40c09210886ae7b2901132528260f06096a51bbd923f
z5e46dacf1dafd30329b02f7704e7c3473d8cacca1724dac9f450447212dec00e404455f68bf78d
z35860e9f2547ef3b29745ac586eb88aa8db45db74f8c3785785302a83cc00da10395a77e9ea7cd
z0ad4c753c3d0dc967ad6b7df3b44525a4b837b824b8d9579ab0b8c26ccfbbb5cd0a088aebbaf4b
z344323830177d7ed700b2c5019581a8fbaa2ff3c38370e3a4bffad854e8c1ad9fb1aab3f2bf19d
z0c68b26705352455625f76b5236777cb319fe9101b7dad9cd5ce42f94ae290c04bdbb5d1584fa2
ze49a434bcca766aa01a0e03f609d51e6d7c26c817096b013182294e2be6688e913a3e7afbc7e94
z3f924d85fcc44ba8f1946d0907fc573ac1a4197dea1523d8be9ea3a9af70bf0da1f258ec586f70
z9171c791147497e58653f63c6f6f6c42a45bf07d33476be6b362f170520ca04be2257fea5eff25
z0232043804f3fc3d0ecb7d61c02b5f3cd7f3f3906ddf258fbf6db944c95892d8b78c52404a2270
z8870ba3a2a558834d06d5774c9f0190c7f372d06df7ca5e44d509f065fef2f25abd6075b425db3
zd2bc5cc9959f3a3847ecfee66d157c95aff1158be10f7c1885af199c648bd8b28a99e01317e400
z252a3240b79327166ee63ce3c94a6b3b527855833eb550607b03e12bf18b9478fea35b8b1b1915
zc761b47f96eacaf5ed62fefdd91eaa86a5ee797c82575322f392e1b57fc50a3fa0d3e861ab494c
zc8557d65fedd974bf3bfdfcbbf5780625931a5fd7e297c2e361c3f3e315c0b0ed626ec4a0427e1
zc20f090b22d89576735ee3b93f108ae2b49b92fc436f84000562a7a4571b6736193306a53ac970
z558e715757c67b7ed544e0bf8ee9e971ea6365978d7dbfcfbc27c5001d94839fb3b126b63e786c
ze7bd69ba6226e9f8c3d2423a69147aa288d49df7f593db11f50c34b5771ab16e0fcf44774b8086
zdfbfd16198d688309ff8141cbe9d36b938711c44542c354cdf62a7aa13df654b2a5f597e6692c9
z9ee775bf01e10949d051977665c3ff86a8404dae44c80ab9e62cfc956145958fd3f413e76d25d0
z15f76c058fec14af0ac603dbfadd973f6ce93383364b3f0f5995e174cc54f7d92649d7ef15dbd9
z648ef5cf89e39eef197b5a769fe4a046b35bcd492b45e2477472e49170572eeb7f01a1be1aecdf
zd1f9996e9adf1bcefb6e6b7d7056036325029507c6f1ddbb65ede9210b03b9a1fd49508ef7d181
ze8fc9587612a7978bd155edaf362cb7241fe78072554df77ea98f88c6d62e30d42e56340654890
zebbd36d7fd2c4c3c5b9742abf8ec1934e3a13982fa6e1b4640ebeb61ab508c55a74e68547d92a6
z00fabe1569eafce817b49e17ed36b0973425c6af04d1b657b1d2b22e0d9fe88888c62c1354e6ce
zc4ec717d2f6fe0d4efba92f0627a513220b0b594fcc285f407444032bbb552c50ad06caf9ffec9
zda44d59028e05f54d1494888d41e6aa114ea0e978f172c0656d4dfeaf28c7ad502ff02a384d588
z4a31a86c91755135246eba2f09c6404e1f60e5110c5b51c8495284d245c171f3982e0af34e977c
z64e1700ba46f8137fa6c326cd90ac6b87442431c7a71924f11b818d10a2327023a4dd860d73804
z5350807b957679550f0fdad4f7b5a83b0fec5a333c4e4d41fd9369ef2c740fbcf305dfefb7b650
z339ad3efadea522d03b8f1e9f878aedfdd976610df8625b4bff90cd4c55224740632e61de2ec07
zeb311185b183561fffc7537719d794319176b3670ea47f3f14360ce07a9d976d784c0be0c16e12
z1d1769c70928175bf488e96658e085012823fda29aa7e04420bdfce86a47185faba3b42091d8a7
zbf0755b3172b54da23d5e2d2791588f6eace1910d465731510b8d5f35f30ebfad9675a3cf87766
zb0516c352e18ea77109501502e5dc8a6f10dc5bf326ddc643540fa6da847aeee2abc22a5f37ad9
zb8e245b77c6dccc895df7e3d40d1e50bc32b77803ec114821624d633d9c4243caced672782229d
z3919022c5583e564f2cdda480a3407d794c303bca793ce3c9620724bf261ea13c89d3a7fa96719
z5eb13a284db9351b4a4652f07fa889fb51604f612a0585038747653e28ca85c00b9d8a8b2b8638
zd9dc36e8ac6689b8bdb903d1ddfdbf4c5de475037feef54901e234b5c6d50a588f2f0b5ab5ed50
z33cc2889189cb1d062e5107ea4bce0a4221afd333909b12a276f56f13a39e7c6d99a7753b6c090
z528fb007d01a084726c41d7d8755ce2a5bf0f28a208cd32a4804c6e0de7a5f5d8071ea243f021f
ze0c431b5ce0c95328a3b99def9789193c204ecfb04d22919b8e668b3b3f95918865eadf2405321
za7db4a4da3540c6bb9662f7dedececc34330a7b99c089b29c03c9cf9dd57180ca87eb96ce1cffa
zef4623062fa4ec5b75560f3f0755eb1968f0538905c082e255941a46552ef4b3ba9661c5d66eb9
z4150c53ae7134884a3a9702107fe2650c0976a3dade56778452e031e578a21ea999ad16da3861d
zb7a4cc4983cab9bb927142b856e32d5b11a30fe833e8a429780620a0ade62bc041ee5caafb4bf3
z29edb33daae6aaa2594acc9140e989e561363f37f3497c1ba9abae6669233b4e22303dbfe85709
z0d360847efa3af608961223125e1a0cc98402a8ae0063734c5c212e64985a6ebb162ba2009f0ce
z69265131d4f206b2ce21793b6cb3957775adc5f3e61dac7d94de47ccd28d7049f43c4b6a0206fa
zb5c761f9d5199df169994c10035bb85d34ac9ff26541f7cb4791610188a794a45499bdb4867cf6
z8959864350fa2d182e6eaf90ad10ebea2e77e8b57d34517e6121069aaae5a6dcad11cb6308c38d
z041b3f7783ab61667a831258e8dc0feaa9dc8fb93fe77a3f62585dc5ab240e5d2b5cd5ce31b25a
zfb9f6bae57a33f2ce0896afecba04d0da9d6d312743dc232f41abeaf8fc281395b96b6bb092690
z1ed706adfd3d97e8fd4f0d5f1d5f74c4e6a54c692b2fcff88ec4f46f396893712318147b26e5ec
z3ef3788dd8113d89060b218088f3bf386e62a905c3a4471dd1ea9bf93da443bd07c069be9a394c
ze07f519bea20094dc0dbf6dab4f65430eeb935e755191f51a6ca11fb9b63a3a7d6ac449d6c0ee1
zf5c55f967f341cd89e233179571544c7a022c48cd4fc5f2934930626a2587f435b7255c42c3734
z342b004e5c0e707701a81c702ebee4418b1c6d28c95bd9ba9992ebc5721048d7608d4078c242ee
z21a5cbdd7c38b570a9a8cae559c9d9f1b98811f3a7b561a00251c4c1f2eee9823aa64f94c9f769
z262642059c0d821977170ad928cf9a188088c6f32d7d14ee133c1672868f8ccbda1de3144cdcb0
z03dbad48e28019cb40823d11a51c00deb8ef16e468bd8f1160e82f69195e9ceb229d467dc1f603
z2e244c299f05baa8da425e49ede163627a028922cc53b747f8a973b834d86e1a7b717d57ab75c0
zcced493c382559576a0dfbd20e4b5403f709a0271a65e1eaeab27beaa605551b85f6f11d8b60ee
z5a1e296559738b5df150d7f05664e56aa846725f0606a7a734b15fc9f3014788e84a53c038c712
z38f0ee1e1420f37f251cc6b5cc8c9ec7c519c9d139f17135082e8e4a958359f1a5cc2fc70f14f5
z315f66ec52b2661655a293b4e8bae847ccba41f7bebc77f8d3240e75cf5f15dd2777a594471640
zb2f1dfc16bc667867f527b5afc8b5b1d14c360b68ec5ee3f129cc30836d7f9945488fc0ed026f2
z6d42c27150dfad424f1335456e2181006f384ce878964e6ff5b27df58dcbfba6e56abb420b0ad1
z1074786ace332f8142e92fc0cb6e77c92e6060499228c8c37f291dc34c37fa78eb513f2a27df80
z9443ff9491da968d62935a126cf556a6cbbecbab220766bc098e2da08c807ce69d390891b321cd
zc126ed6a82d126501583c25c70fdb2fd8acb2c4819a2e92998ab9804e2a29d16e44d4efd483166
zc524bb55b04c05f604e568dd6d9acc0c6931fe1ca9a979676edc410435aa6268db94b9ed8c9e28
z02e03cce12a4d6e6564d46d04b837a6f9164c7be92664e10a23e73549fa68672cdd8ba881f6a93
z3a8b454a998a07df45c627f2bd4254d5ee0dfe3b3bb6c5d465ad3e9288b85d2b3ae5ab7effb7c9
z542a31fcb568c98230582245a03bd84a1eed55173b0fe4173ad4df1a9b924883d10e61a4747ba4
zd48bbe172113696292a8bee7913abfa3413759aa18b65e5efbbc3636aa731fd3f99306503ea6a0
zbace3b0d36a4b23df145fa71b61d13adc25438d6a44cc3336610ca3ba7a7d3a5f94b49177b17aa
zff2bb7f9d1c007f4a99ed963a6b0b7773bcacc200208eaf7f01c880068f90eedaaedd2c9452c98
z3fbc51929a88c006ecb7437e032d7943e6307fbb1558a0c25180472743cf4d49f9e2afce24b080
z8257935e53184edb950db57c8b0833ce86474245a8cf661fa6d8b38cd580f5ce86a0ca56be2143
z8da94bf092b9d650418842fbbce26a21286b433867fe1e9c329fe710d8d89231b2134acb3ac29a
z1b85f2e7f8bb2c171321814de863b855103b20be7ee4f03d4cfaa5e4e2f4d0ed5b6cacc047b609
z38ce4645a49ee9999b00a4d46966843ded49661a131a32846b18e8ceeb94f0ef1cd20eda922246
z3edf684bb225e16db9e2a9e613cf28e54937f9558eeddaf9f4cb1f990b57ed75ad77f9015bf07c
z256b0190ed7b75b49c8755857428e93fd748adbf4bec02fec57421b2b22a2f8fceec0deca97040
z18eb270f23f7c2c25ce0e87b974248a28a71e8e9018ddc11e5fdc89e17effc134f92982aeb7ed2
ze084da6477eb185920e2a7ced55d63eae41ec6028a2739c191ce55b097e89b1702f732d5776b05
zca7cde1141da4e12c418eb72c78ec241cab3894dd2c4024c20714fa857541afe475732293c7f58
z8013957577a92db5313fe9fe125338386f78361f95d93f12a94293f97b6d6c15c485515145fec7
zc91167d5fd0561e52b74971ea9073238120cb3a8b2e01c4ce8ec61df1aa6a7c1a6301583008beb
z42631971fc4b4859b6b79191b9cdd8e769a2278849bfe60c0ff770f89b95427dad650c1ceed844
za449e75ee98e0ec4376b501bedb27b7c5e877a277114052776112d035738ccbbf557708dc72f5b
zab7614921dadb39990869c8e8f0236fc4e701a20a375a9b5c631c42d3f4c20b5fbbc9bd70398d6
ze78ec60fa6a1c535aab68360b598b5b6a80bbb063a8a9b8bc83f733291a4545380b9e4777c39a7
z3a000e533d4b6b65e175f59d4c60bb5b463f3ad619d8f8ad4b754624cd59b0f979f2792432e699
z745efde6fc3ea3ecc5add6154d70db29f6d02fe993fc73d1d64643c65692677bc38822b184d18c
z8892ab0442bc993c7d325615564b7b79ca516acafd27e20043d2aac072d59a6afeee55fd3af370
z1e5b66994c2f15cfb0efdc9f651ec37879f354a5bc3fab3d6ef7a058f8f0a23dc0d6ad8d99ccf0
zdb1a163dcda3f73b3ea090403b03a8b32a0f8819870861d3566986313999c397a1e665f7670ac2
z953f2f104ec8132f00b4bf261d489e9058b2fb686117920e39a7dad24985317d2d29656f228add
z0fd6c08b1faab3a5e58babde6f1169369a656132790de5d7fa37a1a1b33b23831bf2c54ad53dfb
zd2f2073b6202f67472d19befa687ecc6abbe8a3572a9ce02d4293b3917daa898cca48c33928cce
z3fc72421cd9a2d661f4e652998c70d89c2b6dce56d68ab9059eef1873f00f0da1bfd3d5b3b4b64
zc5d87216a824718c50c398c23d526376a710b6672fb82c588d0a8d39ffe3e17fe8604bff3b2eb8
zf65e3ca28b100a094b089359fbcf92fd2510b554ef4b0f2b90810990be9fe8936045a6bb9d8612
zc5dec6611288058ace396fdd899f8b31bf9137b67e16be3ef6b093f4be9be1f955ef4b1c0b1a89
zfecd6689c322153f5a0f7433a684d00f1e9d3f70f16e9db7a3e21e145b8a1614844182256eef49
z0ad09beba53f6176276b06aa7efbb8dd04bc3c2dabb7733fd62b072cebe845dcc38a4217c6d8d0
z99ad9da4d09e566a4cbe63ec6aa86533e75d2c9113441b4c4ff5df1fda7e0f794387f99b86e536
zcfbcaeb3404ef769c79625b84b8992d32628003f36540c77d44bedc266ee8bbb7b0f0854cb892b
z3f3b1eede48aa90bd20948a6cf9abdab8d3d7b0786b089f35ab7799f147a2b99979c0907dc89a7
zc6c34a5a9f6619bcca71f15081871cfdcbce8d4e383445df3fe9e0a780b47a0d8aae0b57c47b8a
z93efc6c47c9fc47bf049baa80a48830e468f22f655260cbb81d78633084b0d5e56cf43eb96f767
z060e4d0754f01a1d402f0ceef96ea1234addd418f3756d7ace8ba2a3505d7b337fa47c8101dbc1
z90aecc9f3cf664f25bbd06471d4f7784b54caf6b0df74dec7e0b7dfe53aaaf0d5942fb41c3a1c1
z855649f26f0491642f55cf4bd38b0850257fa8bb7f190f4e03471a737fef1e705721ec8a969a42
ze9b84db614b31d3979a577e1ccc844059588c3e7f19f9eb8618fbe6e4198048239fb51b09d962f
zbe4a26849189f147522fa2c846f5c07691b24b6f6c7d59ecef4bba429ed293793216d38d14288c
z1a63ed1f7445d7f11a4a14d2f0fb8c319ec1dfcfd4b75a83fe172eac5a6872e53a2aaca5642620
z17dc10b0f221962cbb222618f48eaa897f6ba99c27f035cd276fdc42835a04c17abe45d72088c1
za83921f143634fe1bf9ae735785b910669950f0aa10679e32757b334afc54fec89b2959f124773
z02c3794ee47f6c3c679b293ac3050c202cdcc29405f31400743cdcd7cf83aa0a98d3b51208397f
z4c105bfd6cae19d4c0fb154c4334393d1ad7b82c1cd3db7fe28f4aa35f5bbdeb8ac79f7fa77d50
z837961daeafbc340e28bbc7947e20ec336a0051abedb50d3b85a1b054d5e2ade57daea4b0c9868
z907bf4a95935a9a19fb69448d9a8d9d2dbb7c978d0d3cb2b83017f63feef78d813e01b01644cc7
z89a87019d88c0ff544b1bb66e1716932f6b5004401b5d7be8a1a992c4e4e06c5cb59f9ccfdf981
z4f878854c1347939038fc7f263af55191c462ddfd7d8be76c4adec78cdd1a3d934a97dd54425cb
z72f0b00bbe49818cef81a619aefa64204da00a6ed85f3515ace4f334a62a92746da48ebaf4a692
z4f0332c036398de8573250e5e6ac26992c0508c6ab7be358256f79cbbe3641a83ab5a9515656f2
ze48b415dde7476b4715d62e566a92bf3017c3291d7c68340e1ea49bd0b6e6fd880dfec63ba63bd
z6d80888d0a8e4464de881594f17fff64706063e2f3c4cd23bc912ccfe3d49db143de9488eb6b10
z412d4a8aa48cc70b60a795f6b2f115513206c1e229c7e0c7b10bc5ad079c2d114c6ea75f919959
z3acf5d5a4d0dfd8e210965bf9214ba4e1598e9235bc51065ab1cf3bdc32adbbc50af04483fa431
z6f529ec7a3f22df93f1a5fd2e5eda7743f26601a5b5f22a03a3e30d717a20a46fee61728879b88
zc36ae689c11901f15fd5b9bda6c6d7d200ddc72de9ac838cb6b39bc495450cfa3b55b5afbd4f38
zb3cb12665a9169897da4e8aff8dfaa28f2b483ee476aece30c55a1e87b469b415f6c38e18588da
z8f65a7e30882aa2b7df58dae7fd444dd2a34ce8edb79a1634dc920e7b59a67374337b386d6b4ee
z9bb384fd5553b6e575d26f2c579b9e0503f0656f9905de35c94601227cc9a80d117742452fa91a
z0800fb5789d4c477ec2b40930d239f00a65bb126a394e9d1836208a01b23ddcb487f2f0ae96620
zf5f74909cd0155493cc89f6a6b2f2483d871818a2386ccbac86e0c24bc08696d62e556a8ad150d
z56cae9da57b574496d6764f00fb64be97a34fa6e40a080de00114178eb0530cbd417c1e890e819
z92aa86eb4e55b641ff606ef29a031b3d6a8a2ecb21c2db19989608ff3a00c98296c5928e533459
zc536e34892ea618776b3c8aaf393e498ad7af171eda90c22aa5a20430af3ef33fa6cf302c298dd
z8317f557fa32700af89eb97d47c1d325731949958428a5ec0e5121a229768f129b68b87c141d14
z0bc4398e879a71bb5e5c5ccab917d104b973ccd89ea327fa24ed68452d2af161d348a4308d9ad1
za25f483beadedf7c80259b41d9bf0256df21ab224076a31967ccec2759ac789381fcadf4ffb09d
za7cc4a824cb6b1589a24479ead7389740c62420c7db133d81fa019a4645af6fc4ed8bb89060376
z515c3587ee210cf32051874b8f222420b426e2b81792d331bf466e33515a81296424141dad13bc
zcd7e6176faf6c73cfd40607785c893a52df69691a1e7f3c37ae827d664b1affff34c8e9be3979d
zcae584108d387ce85342506f8d1fdbf0c45e4211161f544e07a5d1b4a7fae6046fbe5d43e9bf75
zc0b5e864e4dfa0c40e5b42e03a7ea637bff29ed9dfa2bd7ec0038b0883d3eac5febd943f04bc8e
z6c2f7722cf37f8a53242261f0e22e814a82bec983b7e5916f49a35fc7284d054919ee27ca8a2df
zc6eb1194bb68e8a7bfbc0b90b93b98e471c9df3fe0339595d1b738b74d46e97189fdb932daa509
zc7996ef9cc63c24026deaabfa6bc9c54ccb674c4745ca3023c9ebf5be7542a8bb795e4f72bfb38
z57402c596e217b48d29905d86933da9b87990aad9f896319c36b5a06c5c65891fab14c387c85fa
z2840f21ae99ed31d290ee521e505bd9fab667884afd3ccb8f13d40e7ff9bf78f47bdcf32eb62fd
z0cb934a6dac1f97268661283a86651d52cdc30d53b176db265b6ec97becf766f1d07fb6738eaba
z7e4e947851cb79530a56d5037a9ad67a6e4fddecc9f678f7d0c28fa168ebc5091bf03e27f4ac26
z05078b72ef10b10adad6cf2377e07766d746b607040a20e8c220afb042bbe382e0962f97a5aded
z3f68539f28445c980c57fba085dbd67f9bc95438cc3f56fd1cf5c1503239988417239866a00e0e
z121632eb8b98081c61485e17b132a7f65b283e8a2f8c80c840665755b3b7d98bf2629205e5cea6
z48dcbea7046764cff7c04682702c95d88611a092cc2d2c7f11652db824593be9c4f9c6931ad36e
z04eec60e52bfddd0fc70855dc60b04c51a235de7b8626d79438c409ec562b35c5f3f88eaef0875
z2101dd778eac81c8048391047e893b2f5a1ccbbeb556cb2b845326f878008d475e9d2b6369aded
z1b5b1ec39737108d8a8c0962930553ba9bb69d3ed97ec2a16d14cf5b066e8bffc6ff230ed287bb
z0edbe31d96c1c83b408ec8fdb3cfb7e28fea85e6d329475809064fcd7ee4c4cc6032acbdd01d62
z28eae47036b1957882920bda532cab8a9e14870bcba1f5d3b03fadefa8bdd0c9287c4c5c9c7a7e
z3c07643a8a4e9493eb9f5ec5f01c34e593d17fc2c00904d422e250f3cc9290c8d36c0e1982c49b
zdebe3d8f375c6e7049172306db85711b122ad7a3c700e65bec7f6c97040477b3bb364786bcb495
z7f6966e54fea22e7d8227bb2dfbb200a79708a6b3a7aabe5558d953651376c224a311b3746a54d
z4c787966c4afffaa5da14c6cd9d75f190d81e31638f23978a5c61daf40bbddef2a9947ee493f35
ze7fa84a77f0468083a9c2de80ac840d4d171baf8feac4319975b15d0b31631c464ba3bcdca9341
z53556aa9720240062afd74285d589adcb833d0441cd015520364a5d00e7057270807df115111a6
z3ffecbbfcc716d340fa5dbdb2a9fea039816e8cf931a152db44380ac366dff8b6b58ec00776794
zb61d562571b36e8dfa059d38764b7b71bb0984b468fbe47e22354651f85b30d81d45b9ca67aa50
z578baae6f213768613f592ebf87594f786313b57003e44c7dfa4fbf4ebec32b9ce502b4aa1a106
z2e5b6f47c0dd31f7c4acd603cedd7d09393ac0d8144ea4073af7b8710e0ddc5d87c1d323c33924
z8d1bf5fa115c4cb77efb48edee6893c86831dbb4de13e887fce975a8afd7d379cab13fadea8802
z0ca55436a85d4ed2d90682fce87fa219b6c58652ab95aee4c2a5b77bba63f4a362297a0093bebc
z8d4298019212e0bdac26612dc7c3e50faeb1e131554f3c188fbb1eefb47fe02e61005d775471d7
z5c4dce5b3266191d3bcbed1f210e5b9cb41769cd6be092c62e3a3df42833aeaea3d9360a3f8bfd
zff8fdb6aa89a44af7db47ce229e55b27428cb44d068690404d36343800e3681a5dde2af10a9ff9
z267d0aac04df992bc044ee3bb636562b5740a26ec9ff40ca13e61c87ae28b393ee4c113660f185
z2c0a3ea206a01aab990b293f4d1d70de1c2832751e1f738224ccfaa447cc2343bedd5ed78ec4bd
za7207e122386eb787d8f924b91bcee2131f7a86bcd5ccff521692fc54425cba38b024ff9362394
z6ace98d193354c97a83c1d3c294ee364ae6152f04b65a73f0f4cb55ed8e3bf16a7d3285a6f7aa4
z5ec432010e30f5e2ea55a18dc12ea72b2012d7071b3472ec1175f5e5606f7abd709091307049cc
zd90ee18da0bb4fe5cc0af10da166f5b0f6d48c1c02574c842fd1ef9f72633a6d5898fe7cfd1bb5
zcd5a738d18c67c20fd973f5e0feb875792131849ab4a8a57ff3571ac1f734d7475697d452e588c
z5a956a0ed0e9cad6f196d1e21dd3782e1dc09e34f48dabaa15744dfba5ca33e6c2a2bbd9faeaad
zd6da90b3accafc32d098af536cd7187c8a5fd4b0d80c2459bf3e6f996b6b3ca30029ef1a0fb969
zb3dfac26e52b2c3e834a0675cefbf0bbcfcf1b32bf84df305cc5193f080f6c2b69755d57a2d80f
zb71d76dd68b89c6d5a0694e35db330de5b66c448e7fe37fbdea40a5a99b902c6a0675fa984a7e5
zed4ede7c1258924f04502d327020287dc97efc0332a089b2eb19158f99e795a943d233cc61932d
z72057e1220062e4eee679a245624e31b7722b0d923c8852778828ec9ac6f8125109b4ea890ae21
z098303807adbb0b87cfc0b0c910d06fda7aa481214f79cb310cdacabe5a0793f602e56455b6da3
z6e67b0e84cc8f9c1e91ad99f719c6cf2a2bfe9bb30fdc4470a791649e33ca8def28fe849c91ca9
z9685cfce6eccb8d2c7f2c941534a1aa555fb2a7c5c1f7cd319ccb832efa45e8d08dc88b3e9e6c7
zf077f989ffd87945dac07d70c3b37327b88328fe4a46019fb419d5d0d8b16fc9b1349d4c517e41
z55cca5e52a786e49d20dc0d6337645cb0d514c06965abd2c3b722fca86acabe2ee4b06e0e6cb40
z60b09615d24b4600b945bf9467aaa9d8ee38bc06d7723566e4540b20d7c546a16b9db34087d316
z8647da4e2e6d209e8d8a4167de6e252f07ee3e1dda998665362f72761d1e40ea0cf5a8240c646f
za09a1509a14fd1f09f6f5ebcdef4659c45b528ed360b1603ef86c7171dcdb99629513c45c372ef
z4467c21780dee2d54c28f4ea8282c8783c79833c7f85b855978a87accbc5c87815a98d124b45f5
z62996f02a7e81155d9360d7feafa8f4312abe313d1f9400b69a17c706123401eca2b850ef514d5
zc76588f1adfb20f7570b81c5a76f046428486f5fcac563fa5c129b5dc3721d9bdabadcf69a1ac9
z16329961f9e450fb410f5c4edd6662be55a8e43aa1dce3f86d225b04ba45b23402b3e7ad0e50ed
z65e8aecb5d6d0fc32bb23ad1eac9aa0789c1b38bb50eec3a925b60a698ee6ff7338816c1859afe
z55b21c12eb96ca6f6f4f6e472ce935030b03b3c2035246f8893d05c8980ea1d7d375eeaf136f2c
z386633a299514f67916d50a95ee64c2c5b155e93b018a4f60e700a0d34ae65a7122af29b3da58a
z6bc248bbdcf22d30eb1258d3efca025d7260ad321659d98adcf6c2190cfefade221f6735d8ff8d
zf602afc2f9c29e61ad7674807d4390333fda9d0d69fd81aa9ff96fbba2eb64a00ee203e5a1526e
z63da17c2bdbe84141a58b09cedf49400e9b6ba971cdce17f46afe3129793debb3d227a411e30d7
z402f692e5f55b7d2530e04fff957b34fcb95f03c74937f81ff4e82d053cd0808363fa417155d0d
zcad2b9e83331a83ad8bae6f80397a85326672774a73216d9b932654f4291d53cf3c3505df20394
zb54f573b62fd75c875449bc28a8aca08f3ce2528ba54959e0319a7b9c3287b66fa028deb88886d
zb44cfb2b94cacb732b6867432e92f9a962dd792400b5b8cf7b9f662c13ceb1098423e790774bba
z2329e3c015ad6d448e3d2c81356f2f6773bd8be86ae0848906511df7a1ffdd85064590aa33b483
zedb759ead1e8d3a58e3fa33383f2206e19c27596c1f7d7b231e90c53c3dca273e2756799eb9d94
zc751936ce6cb5dd7e0e2fcaf9824596cac5e32105a6b855edf9de2f026d948fb3ddad7b6eb00e2
zeaa9efde71a4f6afd69380c7672b6bc8dd17aef0a256d4401e1924d95445b7b4f0069520db7c84
za582eca25885f752fc7bdbc076da93204449f0aa6acdffa82f689c4d5da475828a374d87b74d9c
z6fcf534c6d9b80b88a8013552e63e3986d12d280f140d508a7ab890bb9af6964c0275130230fe1
zeabb07c4aa87d25ded1a84e0512a047cc39fb167b6488a8930235938c215e412e2012ad0469c12
zb5265818affd3bec4d3bb84042de0ffb7f3fb13729e1da8cb9432861a1f57f7c5d6a9fc733391c
z134364eb3464c593cce6a42ed7ad7477ef3ea8863c6d6ce955ddf10ff91af95a200789a746f498
z6f44a94d7d0bab3f4231bf19f4bbcc98fc550ff8bac58ab3e79d6df17b992ce721bbaa52f1cf8f
zedb22a7130d05022e550337e8e99e8b4e465fe5cbfc0eab14705fb4f88d3bbcc5ae8b607882e53
z6d9dcfd15c1a78f8628c0061a4ce89927ab7c053ab93e8b7ada5ac5bc340ac7b306a0f93e9e179
zf22d1f8bf21878eba2c466298c007c75eb9706c977f752dd3a40ca21a8287f2f11e877b4623975
z59891555425f4c202a755667f912e4c25305beea339432dc6669bd5e3aea13a909c6c6f6c4242e
z28aecf4b2c330c66b4b0a50d85905b2795042b3cbcd4f156639dfaa1ab6e37fe47c616d976fe98
z7b5e7725da69b048e86776ce0c0ea1d8367c416814c85bd0bca0ff934c39779fbdde093274c4ce
z6638f9930345b351fe50792e51041c54609f99ad710db638fe906312075477122f0ef196f7e6dc
z3da0b4e2b4d3f31f8a5acbcd71735335f6b3032c60049b6e57b5941b29830fbb89e46c11928f99
z7c02b7fc88c944d07f0164fca5ed652b27cf26b699d39a9e53bdcf99676467946ba81b48a27b32
zbb9403985332e88b93e79aec40f79273ab139fcdcb26c8ec4182dcfa8edf0230638e32968e50f6
za716289bc4a5791c413031c2b6b736b3ddc029d8f9d4253fe61d5a1f2d9bb9ee4f8db539e140b3
zbab8528968b12b034401169ec49b021933160282d212016289229ba7a3b960f4799a13fdc81136
ze8be87df476230e900e5d70e1e64fdf62ab5703e8f8abeb4fee8e98134ab79ddc1e4a3415dbb07
z0aff996db3eb251e357fb7f9881f72cd8552833b1f6e5813ed910ecd1e82c4f29858a180dbb75e
z816ec4f65ee4ed3d94cfd2290d4e23154f98063b358334134255f89cd69ef01d8805612b8df3ee
z3cadea0e3c9eed6c661e7092eeccc2904f851cc35b6807e27f3fe9603fb529588243efd032cd88
z5df36793a53153cfdcac16deff23eef36669a1109375b505fc43c158b06d5a791dc392eb3b413d
ze0762f117e899b593bb3af8127516dc6a12d3b65a1818237bdd5935dfe2056e77c6a30773e0902
z23ac097f3927339386828702014a53187bb62c40bd30bf608a2824896024133f08f18c772a7099
z42de068471253b78d2f7bed8fe47ffade8c72b2219984ce2108c941d184cc5fb96019b009fa28a
z07c6cf47763f60be841828811a02ffb9152f2b7f020228cc9eb8467c414aaf4d1a0687f94c0a4e
z2b3a24b9d4335f4826e63d97672bb6579d629cafe8236669ec396ac723ace6d416107711d5ad2d
z7910fe964f39292149bd7a41dc131dbaac45c20050f82caaf2eec7d132344d568bd8e4641bb678
zc4e7de69e6962d701e36244b63d29e6354c5934a6773443190484f43d259eb981094f33fda1d68
zbb9693661e3bb6bd509edb2b0151076eb4206d1eb480cb436b231eb210d3bfe959b5b5427cc6ba
z2a5b8cecaf23d0a3aacda82654c22db831e500e9a41632a61eb922a0b8f32dec936ff0ef1604ed
zfdef877ce00f422b8c6be97a9c543841f73fb322dc9c5b5a82699565a9e2e1d74ec2ee3c9d2422
z98434eee1355ce2ea85ad284ef781713b3721f44540aad79e5601029612367599d01352c29274b
z311bb1d5398a7b4ab5be61474f2d28e9ca9194eb726966c086e6058155fca485edeb81481db363
zeff82abd9d8796021c766e7980ffa992f5a75c031b918bc46b55fdabb6eed3f48d8f7891babee2
zf11ad5256f8019de4cc130baa6bd318a113c9757da9ac7c3f3bed318e215cc6537e779c72ffa38
z447422c8b7ebabe6385464e95a1ceedb67911fa0edbec07152ebd00a28261e9477bc9b236a1725
z1752f1f9444a00e306c44c7c4cac6d69a7436819372652410ffcce42093f7439b38dfbf064b40c
z3b3f0233d712867141aec93254bcd528410879af900b8c19f236c964c74e383c877c14ddb48fe9
zef2a69f6ca51246ffae0e21d0ba868ef43531f78dfa10e3e02dc01790acf940665646ebc308a58
z34ea136d9782c73e00457d5220da1300f3db7978f2d7a045c26e28557d73594fc137bc10001c01
z5be19fe7e76f6ae71aa5ea3b18a68d87d7a45be1ec6b2f2f579987a5c03b5d3b1137c4004e89a7
z1e4f15c9c66e9d4a930e767e8c341d45c116266681b3e49df2c2d021487eba74286ac74a1a6cae
z417878021473b39d75e68244ceb9cbf3868d5641ab970406d58fca3430bf19eb3b2c126a60a601
z0207cf0b3a78bc5010f824ee3efcb36a601b29e35732c07e48bfd3eddd5ee0fbf718baea353817
z2c98b1cbfcbc11a68a29df6662290bd67197a4a4166957de3a5115369b0ea0bd83c0e7864f00ec
z6ba0ce061f0825d3fbaf39a8adf792413b77b6ca168112470cedd34680e87da3ed07542c2f1ac3
z1e18ea3e6f9f482d1bffb2596e84467e02746c398106b042eb3f5ac7a8651478cc6380527aa89b
zcc69fec8f26412e7614fa688c4607f5312e7bc701ee11c173d9de770afbf535f56e46c2da25907
z26fe8075b2013269ac0b3877319cc6b3c8eccd8606a0ea13a4bc759409c32de986d5121073fbc4
zc6c6467bd8a874902fb8947e009a1a0ed56aa8785ccf6e8eac645dce50e3d872fd381d7ba16a5e
z2772aca410464bbf574cdef266308c5cb7f90a369eeecee735076406d3ea5e98f02a2ec4a17589
z45cb376d1861abfa6e700aece0531300c21d1f06d420f9ccbfcaf2af1a6a9ce7fa8db888ece875
zd1b119dacd6b18cb125e7d4b4dd6411ee2ee58df99f10fddf4e4a4d5f570ac0bd0098b72ebfda5
zc6f2f35f1f5b4eb97a110ff4d7c0ef397195d407aaf32452af12c23f95fb8adf88e7648edae051
z2f4cddf75b440b4e81860cfc9a0e65ea477ea6c50af79c5c292a97e10a2d237452d7d7c61d835f
z316b369fde0dd3a44f1266c0124e60f6026e2f125f1f43916aa13778fbefc9af026fa138e415d5
z1ccd0dcefc28f2266bd582cd99bbecf259373f40ae99b65889fd2cf55642d0f624706afe5730b1
z00103bcf26b6a284fdb3bf094295d8617a976fb1edb022fda0c77195e9f3907e30a50f74486544
z2774cccc017eaf55eec390a251c6437d176c34d116f1c56ce9bdb6efb4c03d9d78483727ab03c4
z27124818306ccf2a7134b8ff938fbce9d48de7fda573cd3aaf70d6b27097333643e75bf71db251
zcbb520965d72c0bbc5c853667f7d29cdb0f5e14d8843584e48a17aae1ad9008788dbb48811acd1
zb8e47e44220b4d539fded834af28ae528c8f07615f152093bf364bf8ff932f77406164b02a5e0f
z741e910d0d7c63f201cf874d25147f22a84b6c6ea218adb797e1bac74d86cdabeff82a2599376e
ze9d702b6de3d97b41aa8c0d02439c62f0c12dfff6c5e32300b195c24f3ac38676e53dbd3933559
z430ddf9e5ecdf534ed71e05d15ad0a043bcd2430dbe33d217b640800de8bde133b70c1dc6b6bf2
zdce6f3a6dc552c6c40e450f1de84d79e5677aa2a7686c152193c2c2f114cfd7aca99c130bf0a56
zcce30f893a3dd0400fd8b0124af4e0590a63f0a12b0474dfa8d7bc772d7a20ef7c7f6e2a8c7125
zd31e031de62d9c8a767f296c924d0f1c947bcc75173efed1de45dd0dd91f09c604e068dded764f
z4c111192fd8bcb7d701c5c9198d856e3bd60c4c029205f3e3d45b5a9876dace6f61c5ef72974f8
zbe1ff7fd6d664d8ccbe596a4107d69c85c6a986ce459bcbc5eeef744adc14b31e6589e680f2ba0
zdc544bc68112c702e3f8e742262218b0fcbeed4df2e8885ef6781bc4fac2af2480c4cda4b96e62
zd6b197a0b00ddeb132ea1566b9e0350a1ec4ef9f7e4143cca0daf876206c06ff801e2f8b549f27
zc51a6f59f3d2c66eba5cceef93c77005694d5ee1af15d96f85836d10ba771088230be1198bc21d
z9ac131b7d5f0cf51ebc87aff5b69b15311e0c4ca26d6d1e467665f81ccdfb6f39660cac3302ab8
ze6477febcbeb99364638becf263eeac3eb274e930e5334dd89445da24605014d07e0461a75ce3b
z1a8385dfa4556bf6d615164d02a91dba2f40c0bbb1af115355cf174343e7348b2087218202652d
z6f240a4157467a256e75124ab42df060b5ac6b83ad1aa8fe5cb8f89022c738b2cb5efe92961533
ze4208a3ee36f424f41c4bdeba255742f49c64aaa58818346b269098729e29c4231fcec9e7fe7bf
z6ff9df7720b3963fc1f010acb35de6821619bba12736e147837a70bc88e2abc80881708330eca2
z6b461999c6410c005734d0020b14349bcf667497f8b2f9d5c6596d9bddb1cb059fad5fe59bbbaf
zd84498b1be803ca6744e961cdbb909cc03ff30aa1ddb5dd400e206b71504e7cba43fb5d16ed866
ze6fcc4a84206fb070eb653f1217b01d8565b0bd1e02d2ec701955f1f13ac72067c2bbea7a6a97a
zb977f90282f881b048f2ba6ce6f73c901a7a49f6eb317058d0bee65d9f90151cb8e6ca1eca4f93
zd391b29f6762d3ba202d3b8d901be2a6cc4c8128050d94e53886ac2063fb2632135803153633a3
z35f4d146d6a3827415e08a60f39d93835272f6fcb0edcc17bcf2480b30f9fc8de4488c8edeecdd
z7d591b12912e97dbccad13e57859dc1f723ff2158a0d7c8eb72e063b721c1cbf5d3c98a0b7bde9
z7e4e3249ec7e7d139b8af6fad8198367b267121724aa1339e6c1eeb4cbcf67aa4d3d780bfbcce4
za02d73312c6d28ad34b027999247a519382a78c162b488950409432e216d2962cff2a918406578
z9eed7449cabc3ed8974822a08751a597478d1700c94c7422c9e11dd455ee8a0707887886ae9d7c
zc3627d064c9331d973e42d1414bf335c750a82401aef83016932dc03f768a52ad376f5d4f716b3
z0593ba9d24e8b3a620f47f422229b45c511e70400f9cabca5da5e34fb6e41bcef4877c7cc31e0d
z16689144c72aac58dd243687e4222a32459b4d18d5ce6fc490865b7e663ce25ee1cc3f0c520804
zc5e4540553c91e2d8df1e9da2d80e87603f3421edc04e1f236cea4bdc1f3d17907d7c23b67a5f9
z178174d7861958d1fa1747f324527880f1e452759019ce52567a708398deb311dd6b42d02c87a2
z9fe979eb5638ecab9a0cad39d5b529fdc5436224108382dd0b04535884c243c599d17a58a1d6fb
z1681837226ed7e2a799903d7a474f2508f8f7018410afffdb0dcb1f1d749afa0c5a886c6e07473
zdc70803dc975d4e2eaeb7853f592aeb77a482878015ccc3adc31bb100ec033211cfd6e7f5db934
ze7ba1178803c67864a2a126eb53a0afd6bb5e3db1972834808e7d68eb81d7863c69d4adf89cd0b
zba28122c757eb82a0f1a5ab2d12cf253b0b7d9d481a68e5c64ef2c6120d14ecb12554dddc074bc
zd428f3d413a7fd1beef2941b8e177136fa453a7f54bc9d3fae4cd25997d7b8cc9e3496c5c0c9fa
z682b7a1218e4c6b22f77d246c758eddcba12b171ec95a502dd365295ab5efc9e1481730e74b58d
zf0b9f3051c36f6a9aef4b2cdd605c4cfb6c5bd3b77059a662368a4f8df240de0d0b122ea4a616e
zf6777be5d87e2d294ed08bedd67d9d789296e88ffd6d3f223ac1e27498541da577d5cbef82a52b
zbbc3d72ca73fc5ad8707f597df86e85ccc346b95c596ec58c24bc5be1d8503d95a0c86f1b6e253
z46e1e9622eff2f2bca2efa7db9a07c8eff3dd5aab9fb14484ce443e5191b70904cdbb446c822bf
zd31748cf7bc54cda98af9f448edbb4abc462db632819c9fa37b7bd3cd0e3cc7285b0ffaea3d0b3
z541890b77fa3fdd0c28acc64607fd4e29f66300a44f5768f6b9c338aa1f17f52b6a5db6d9a635c
zb2ac392ca21e868391d82bb050b84033e891101fc492c7fb78a02c308aed41950f42798bfd49b3
z33e586cc250037f447d46857aa5978decd50009572bf1068810a761ed6fc2214850f985c0389e2
z2b2aca17ca0ca26af207d0141fd7efd6cacf023fe4a36be1df67d060b424eb07bc80df85461703
z86c398d659d4cfd40e43f3a2d85e2ccb034e45f439d81d58eeafe7b2cb58682fdd2f32ee3d372c
z7eca9fa289424d08b5ba2c9633393dee074a7284f02a7166b391d0fea3129982d6214999550bcc
z6db099ca6bef1063acc4371452364515a4d49d57ec16b165981e3365adf70e6606226f0885c9ab
ze01ea7fe33a816b9207baeaecfe005eee145ea901999a6de5d2bd599162214502068f8270f2b4b
ze5bc97d46e4ac96542da022a5e057764afa8a8c8956fc5751155e759205c7c057082cf18c8724a
zdd273cc899826ae860eee6a8a8750315987922cf2c1d6a8c6e7b258389bffff57989c52348901c
zeecf1820b2dd55efb70c0f8b83dde91169a46cf19d06574b6e48870553d5c33ddda776d1da374a
z68354b847d9b82796186b33a253f87f075cffb5e6a8548388f6d1f7811cfcb5247a0d2b34f4ef7
zb28fbbc85929a40ae107d757b78ddfb19918b8db47e3536c890a03c73f2d23eca1324480ad1e5e
z4577c6817fc9baec423e82c463128d17a1fa14437d45c4935620291f66f0a31e385f6203c8db32
z3b31f9a73d1151f75c18d0b689d86a3ddad2b11d3c17c9bce8fc47b10daf384380735363598287
z28c7fb35b5d5bb36566c2fad4de177c2a2b535c5c9db95108161d05125ff1b7d7c3eae2ba96b3e
z1d4bac21e026bca2e236e357666f5c113cc430a6095a9a8d2088c7ea641b14206a5ca44423b9ff
z32dc9d7dc6188f93d280b0a918a8d955782434156f33d9b0360fd59f7df2469506e8b5727de23f
zfd44074e815b1d3104e844fa60eb02cd99631b8258ca99fe2bd169df5fd5061eb3004b5fccfe52
z2738eaee2ddfc9e1be3ef0c0b7e0f53cc56d9b22a0857698c1c8119e310d287ca92031a70d643f
zc1fbd551ae48c62c90e3ec74fe9500f78316ed02b30d7676a9051beefc3a21e4095ee4c4258237
ze14f3151f516853e043fa53be2d5e76f610ae51db6f10b2db9815af99361bb243eee7ffc04bb9d
ze4aa757f68bd4ed1ce7e9a8645736616fbde58dfd6eded0bfc3b412fabfbb3f59488011faba420
z9cd85b345e7aa25981aa6cb50e172f4294f3041001f45f5832978ce7f5828955307fa7cd381a32
z97ec12cb208526ee40c8add04c9fed1de0197aee2f95b1ea938fe1e9d7626761a714d9d2f3a990
z5fdb3c47dfa300790440667be1d4fb0627034d16174bd2a77c2663f2816ec8f3d6e4f4795a863c
zd18231fdd6fe04fb8237c618f94851d3624d75ad7811a9553022dd7448633299988a162305b93e
za823da2941e23d528a57ab94c3ca827c44efcfcdc7c9f47dd01657d33f3d60eb56add4928d2907
z480903135f07e8f43052c41bff7700b05b6d8e0737146f116ff7dea8e4a3388d7385b34b4a103c
zc696bc592d760829f6a5fc5569f8e7299e0e1a5fa51ccb63459fc6bfaf85544c890ad4b88e85ab
z480086b9a04695f9e6f0d1f8f938f20d2ebf2a28d9d09cad45134ae237a0520b90de2ac1560162
z96cffb4127139cce1e2292f0af1b19c9931c594b5ff8dbeb15a26106b9cf299ad6ac8d1a8cc6f9
zcdcff622d8da671c5ec5b50c51138d52ad1019b1cfbe5e84e8c2a2823cf6d3d0349fd2a4ea3ffc
zd7d4f6e34945618ed7f7e56b30ded98866641cfc6b74f62622643729d3925c76ac3715fd2b20a5
zcfbb8a74993e9bc199b25b5eba55ac540c95f9198f36b965de554589a171957b81c7461ae528e1
zb52f5927579d89e3c1b78ce1dc0c9b850132b23d64da685804523040aba9868e21ff661fc0263e
z0b985aab493a59abb848a858c08fb40a170d4fc976f5b447f29740fce0346ed35c304ed91ebd04
z029931709c709c1287693c791f0d0e155b5f9285d15f034127b5d14c7ae362a8d25e36fde8b5f8
z8db3015aab09ab448638763f4741cfeb8f446f21b8db070ae3a90de9d4c5f2192b67e7e8953073
z3838c2fc4fea9aa3265d0685991805964954fe90054c98fa67771dd08823bda5f51c9fca85b361
z90bfcbf5f9fe3e40dcc8f09db5aaabc12b8095cfeff6037ec934d56c9a9b89831849db629902ce
z6aa3ac1eb2ac7c40804c487904673e4bfdcbe404c7efb01ee419fe2a4801100ffd506cc08acb2a
zdae13cb7eff8a4a71fe7366a2d3f4a771789750d3ea4124c3c1d640963b82aa5667494ed03af1c
zc93f47f4d197ab126914314d515b32ec53037c39edcae1deb2196332c91b0110a70459cc59ddc7
zcd4b6c674d6fc3f5583749ad6cb2952341649ab7eee304e0d66aba906966d99de17c330e3f1066
zbbc935b1a5994574a92a5ec7d6b1cf74e62f748601f1f823a4a8ec59ec221125995979257519ef
za75792f9180ec889bc836183509ced3bdf6f1d16e7847ebe114ac3313d3d3db8664412b4424e98
z81646b6fd1eb3177e19b400aebfe4724704e2a980fb5036f37fe641905b10e42a7cc8086b0ddc9
z40cf07362996314363ca9a06ba3fcdf57bb6a17101aa33732a26a539daa25a7af254371c274f93
z32b8e3ceecb6264ba99b2dfbc4eb1aee8fed9c15f6b467f161eabcbded2db5e5fde59480de603f
za25d1a0f2a77fe86846879ccc3e37f7b84150102b3a673d9f03aeeade607236aee9ffa455c2e5e
z0a24dc0fb9e99b1c2e0a574e339a16c96b36089223ee927e0027e962f27985eefab496da2772c5
z2782cad7411522d368134d3c019e3107608a296758dcf999536f1b01aa1b66d1d9dae760fcc218
zd0546de6d4adbe38155d01c0ef695e4c8043b2a24334e54620f36c9a7fcb998621945aae2340f1
zf8f1ca1f3515fc75ffbc413fe0678f96ae42488a9f1eb7f4933477a0ea3f71179212d815ff408d
z1a5b74053d152c5541f459051cc42d8002270818aad3ac8cb2e71a9151dbea8ffaedcf7de4316e
z8bc031fd42a7e412cbf8edc9bf1baafd64675080284d680b6e6c6b229c8659b4b8ac981a5e5dec
za872b9778e1fc144fd99b23f2517df9d525bc028f51f02c8eabf3f1fea43bbe0e4995ecf9634a7
z5258462534468a19927c19bbc1dce07e2e0e2eff80d2daadb8b20f45cbe8ff6491a79f9f3e2263
z5857310c4c480c334a1f9f14ab8220cd50936960d1401a1eb36a98b664758b23fde2c431861bce
z908a0306aa50da155134ae07687cdddec5d93ad18cb29fb81c1bc1cc30923040ecd41d27874d5c
ze60dc4dadad7482ae9125ce1158876038b7d23772775386edfdbae89b25cf364f2f864658a1c3c
za2a08099510c854c0b3079e591cd132f01711532f2661614b978236ac49e58550182c1b196e967
z038e48998fbe88dca611c26e98716769d6e49750dd83fcbf4ff9f8aa4b97745fcd42db65338503
z410da647fba858c7da8d4ec4bcbfed26ddd8dab181bf4a7bf72746e8449d33c49b0c5bc4790224
z3d7e0822ac7afcfccaea914851f731b029e7155c37af1333aebb65aadea57d65971b6052cebf7b
z3fb65ce8a65ac751cdf3b2caff13e8e17dca565c9ff873d155051d03dd104ea934edc9a21b073c
z6ace060e5da1af9c398371e3abe05974ef0612d13404b53edd30b6f09bbe5db04913dabc36d722
zbdf0cc6ba3d90a8a484baac429e88195ed50e4e54ca94ce1580bd69d95a0f81b1c70ccace80602
z26b320f15c0dfa1e8a29fa2d645a8fb4890db9d2f816a0428dc6f7828d002bde999234ace7f871
z2fcc68ae031991c24348387990f7b4ed3998dcc99a8fd4aeecf4c1683bb353e2365462d24fbbff
z34597a9c27a5c4c1139c331627721c333c36a0f92bc6620f8f14cedcbaa5d7a37e38bf06d21588
z0b45fcc8d18f9c95467f22ecd621eec11d09b5d63c4327e11d5c2bf8cee3eaf711e3be02f83102
z37456800ca1281ef969461312d67530abd680289e453975c712b0063e1246dc242ce429ff697a7
z83c1edb49bee9939d6ed2cdab5dc81f0189ac54ee8131fc50fe82b0e0dae7b0ca47279e01cef63
zeace2b9c29e2b277b0cdc2da76d089c37bbc0242cb295c2bc22fb2326e8a85794e40da9a0e6542
z76e4b937f402968c47c9ae5a3784b0a085f2f16d8204412d2b1d77b9249c0fe815cde024fc6540
zeee3854698b9d199f9eb02b4ea3423ffff0c769df8af4f6c227ac3cbe2967fe6f242ae6f5dd951
zc746a8f00bcd7c7290c122788050111f2fd905afaf4b944c3dfd1d16686e8dd838e6c5fb18f81a
zb7070c70b2b91cbd638f5c922aba42c33252118d2ff5d566c05071d2c6c6aed567ac96c35f3b26
z669fcc1ae479c87f993440ff7f6cdcaa8b0cfa7b43b098ce56d275e4094802c4450d051deea3c7
z024fac6c45cd879ccc32b5ad698932af52ad9254f20adbd7f3b7618d1d0ddfbbffde47eb9c385d
ze0b32f0b9ea1710e4c2ebc05e17d7e507fb2bde7b58c7c932c4ba24b4d6a13ce173be2dbe537f9
zc78f3899925f2aa322af0debd86423a6d3de0cf821808e2b1bcf57658e8406a19d254faddcc9fe
z02a90a0fd36f6321ed154a3c356cf9a3e97abef081da41d0ac84ec2a9121b3d05f815c2153e85a
z5402ccab171e45987ce0b2c2e6c3ca6baea1282cdbde28e84a8ac8cb3c228c44bb4968a3e5efa6
zdcff8bc276f911939e79700c4b8aa8054bc88f7c397da696a0468bface202cdcd3f32156b831a1
zb143b6caa6549cb60b726d8472f47277808fc1242927eaad2233daee5d9be258627453cea83a61
z7961f020d7c16f494f61b515701b8abe06bcb4f5a39a34481db1f999ce1bc4e1f6144ef71e0d30
zb2cea6775964f6d24a61fb66c8d2b1cd41c119697a5835f340cd3781754702ef091f2276d3e09f
z0a26bb18613a34781c01b8eca35f2d416e27a5efb894402005667bef11467921a28bfdf21fee62
z8aa2fed7c021fd280677967d2ebbe689afdd72debe075b7031539ae42e2e410590f36dcedb4cef
z65254ef754aec5064450fb33aa6daff56de1b34a156103c2fb363e2b8ea17d6146f69e4803f636
zf88ad43ee91af1eb8dd1b44800849215c24156ad6301d485f8aadafefbdc7a799cada55a728b48
zffdc9e8a786b0da358bd0ca35905018df77473759d467006928230dbe75296d6f7790cf518535a
z412d5d5385b2c5d9253d6053b0fee10cd7f71a8aecebdae446d401fededa0a24b67e8c0d899187
z654721cd5b83484aae0056ee1d3d94669ca6d930b83a5ea4f2c925ddf55b6b973ac870db3019b3
zd1db77c7c614b33afb6c6654f640d36b075b48388eb7bf20353b55f061c146dfa844f05d9c6657
z73151787ef774a1938092de17abd6a1d3a04bc5fae7edeed83a1179aec8e3c2835d9298eea72fd
z24ee823305a591e37162e84a2ffc291cd4910ffb6846425b143f209625a9c8fdf035303bdc9839
z89059e05803ff36f99158e13c1e924e524cdb314ec89283cd367e945a164f2b08811ebc2ceb8cb
z885a75a1d5723d47ba6dcef9b1c17321c42646eabcbd734875931f0b311ff0701fa524951cac42
z28f99fe8e8d5b060d7678b914b45b2c0e5966aa176b6abd27da6b895aa4c0ea2231d1dcdaa2420
zbca4ca4df71d88a32a4dad7c7e2cecb03cf6c1e84a1b8b9ca6c53d42e074bd873d666d697ffc13
z3f1caf8977fe344a55b12e4ddc4964309ccbad79e351c020fbd77f6034ed441b0776419f9acbfe
zbd014bcaa25e8389149f8a4fc44de3698a827d0c1cfb9db850e553ef989c970ae1ad485e3c5787
za2a3048b4d944b01282bbf13a542b53c0795341151bbcd3c5e85c9bcbf2edc769af10cf6c06d4c
zb2fb834e5e523b471e7ef05005663cd6b1f523334e125fa459bc2059bfbf85404a6055d886fbad
z975085b8045f52e38b867a0a07c35240ed4564b20734537fb25748f2087d8312cb7e421c33888a
zd2f41b1337afd731689fff52fe7c5d10acbc7b28bbf904dfcf2e6ca5bb6c7cb6852df1713d7a60
z05688295ecac4387ba04cf0dd3ebeaeeba10b030b6cadd15fd5a3ef1ea6978e6d71b4add517ed5
ze9dcfbf20afde3b99b151847318a590a8422ce06de2d8cff7e02272d76b8288ea8a7eb141c0201
ze295e9bead7935e2289779e1d00e97813a61fb0be3e1bad800d52c73df3806aad2108c99fa264e
z5543edea6a4683b571924109d2f57cefdfd171cf153a785ecbbb1cf6d6b46ef6f51ece7993f21d
z4c0f91991feb0a017e715d4bacb2b6342ab02304237c1ec94eb4df52e228fc7cb41be06c99d249
z340235652c451896fcb3eabecd92ddc930d5120662b111b2b2a5a701abb96cd95644bf7e091227
z57affe4a19bd20994cb088e94f45a3136c7776b068b2361ffe58ccc4e02c854a2bc617cf885fa1
zc2aafe31691b4c6515748c3dc487cb43014424e71598339ff8311513e70d214a41bc389b8a83fc
za0bd5999695b418718a0e6df9b48fc8dbf3f715d31d8abaf506d6eabf2b3c498d41ab6498720c1
zf368d498005b8bde1da44591bebe09d184162d5a2a022d996b18af54cc4c18ed90039f26ca7d0f
z33d8df34ab74d89a837e65ad4ef9b76cdf08927af8a0f7862d83245e6b1de9c5dbf1e0dd9e4222
ze82444514b7a6a1af4196e04fe505fd9e6ed4ef78fe396efe43278c0540873e6e5f7fab033b4d7
z2c43ef9d25e43ebe06d70d0f6f9507c4f806380d6d4d58bd094f95d860355528d7f30733c8926b
za0e6572c6d7b35e3480156adcae84452a7adf77c402ecc7e9356cec06c9605790ad81340d68e37
ze3b30f09eb99d39e8f0447356e6ff06c6e9f50087e63576634d391633b3ed74ba3ef4fe3371ae5
zfe0e6193bf35ec063063fa6e997f69fbff586aade8c9cc2acde228ab9614da88ceb139dbe9a7bc
z31c8c862f38b5bb5a2093e8ff6c82ec9fdd6a877cd386986519acded849a853900d73394e551c2
z5b7bb1c7be173c21e00c9d46bab5f4a011b5e9eca0353cda888b6154db7eb82f5bf67dc426b470
zd56b1897c1e91010d1a8a2a42da79bea25c50ecb969b34c8c37f71d246d3d9ef74c89a54f866d2
zecd4f2df43288ddd3cc44b82cc64d7c4626c95a467645f85719c172658b6b8cd2b6f2bead76f82
z7ab6db6023df175915dadbce92d8627419b04cbe98fc419df4ada81e512c7195b1bbf173e06a5f
zf3d81c3a0134c64f4255c90e0a988ad417d5efa2af22aadaa2bad688033e8c06850f2d05adce66
zf2c9bcba7cdac2c4cba286fba1ed9f65c2bc49c5e3daad0593ace303ca48ed16bbeae2aeafcf2e
zaaa62907fd4f85932b9bae341d8a51d50ee63a2883d29a52b730c71a2e1bdca0001814e041fede
ze606124e7ab8dc6b47e0407b9271e555df3863eff3b745af2276daae99f887bcfa94c11a0def36
z4033ca420d0fe2281c24801d2133dc7b9eb6a05acd68d826b1ff59cd2d00a07f225e770c1b853f
z16bb8a9e5335c1452f2124fb6bf4d6e40fe0d2151830b8d145b5046ef8026a4dba8c53366739d9
z1f342409c442fa14a673effb07d7535566ee0d58d2bbffd64c1621498fd446ceb5079246138d30
zf8f7607e7db4f659ef137abbcaa3ab0c9f358d1d85355437102cf074da6433474f457c1d74d6e0
z20f99255400282f857d6d31a390f07f4471cefcfb4ea16274210d69507637402d3fd539bb90871
z564c81e1dde812c4ff6761f6d51d92169e2da30c3c424d2afb72ca3d561b937508eb9206de4eef
zcca74b5e2b62cc00027f0594292001bc3cb241069ce96fe056d46e68c0c1b91e509ff4b71eb130
z49ff525da1e2a7a76a88341c7401182b5e7f041f2ed0358045f74abc61dbcf34e4c83d0fdf77e3
z1f1125c0a6f24b799bb3a5a583638322b57c7d24df856fda033116bcdeb6f5d92e04d827b43c6c
z2f0fb38392f7a841087e955a5143a64ccfcd0ed753cac5e4ea5430496ef5f09382fe580e05b486
z7040d5e6c1a281c31dab7309e3cfa79fe25086ef6c52aef5c5f7d33b9936825108a9ca05dfb774
z45272d824d5acd22a08e80452ff3a475b5ba46f0a0c798918912a073ac87a401d3557ff9e5c117
z2096a50676b0e27a77917b3ebf10dc7aae12741a168fd044e1739d8c28f038702a4b7218fb0ae2
z50107af15a3c6316db3d6b541795c744ce3bddc133426c6656009cdc5d2a3bb4dfa1751bd7a14a
z405c389979d5b3c83890da968605f837205ac16be62b780415e8b4f9a053618fd3928786ce9c77
zfb29fe27c3f16bf207b05221f4f2d215ca45739769403ba28855da8d686783d67f838239ebbfbf
z0d3e3d1fb8a0874ac02758cd389d2a4e10391e58a4a4bd4ac36626712581b85b33fa456293db9f
zc6719898e4e7ed547a8b4e29a40e384e70f30103dcdd6645f666205dadde9801bbde461ce98264
z1bd70f7b6f058013e246c92513fcfd96499950bf1a0a2693cdcc4964e20ccf92b69a0010b1a297
z1a52c3523c789f24eaed7d68baaf22441d7163db410be6504270b2b3ca7cd7b3887c4dda361273
z92dbe73143742e3ae287f9d56c4a1f688c3398908080fce02255ea33f4ec2fcc5e33181c51fd15
zeb2028893871b4323b5d372f9dd720eb493bbecf0571c242bf444e56885439611332428b728115
z2963ab796fde29b980b94905b023f46069d7c4d470b4b4d012032705d695f41f8342559c255ef1
z081372d986396898b992eedecf601715e27c62c454858f16f77ef447b1a76f1f7573015b1c37ab
ze4adec2adee35b41f6b5c2c0cdff7584ce4f3429c0cc3ecc89fd0e284da7ac2a5c35e972001452
z48c946b07fa95a8f96146c052e73b9596db4d72f0b832ab9489d6655ea0675e750d5dc098169e2
zb02b43c87c57702d8fbcfa9fe3a03fbc349f82d8d3e0f12e29c3d68d104310d32035520b6a5dd5
zcb2b88c41063c2c5c68d7adcbf4f4c17fe8090f75161763a1a78383bb1e752037f527252a95830
zd2f450e05257697ff0c80edfb82f59866e7d4606e374b1f6d5a31867426245a494081105890e6a
z07e9b63ac3a304686f240b678bc97f52e1da7a042618c8a6adf82f107f63067702f1bf467e3009
z92100788855aa14d30b948eeca86978aa70dee1ebc41c1c9c0953e083ded605b784def6cd727d5
z361d8302d6457b766ec7982c19a9ab5b0c96eb8cd6c6b1119618c754ff4d9cf1d7d5952d265c46
z3bdb0c4bbe49a4dabcfb235d39a055275e0cdb51326f9910f55eca88c0a7d28e542c68f842a1b8
zf78efd1a2eaac0d9787df058fc0fc341b7158806d937962d996cc7b62e496f9ed20e607aa1c3b8
z761160bc587bb9798bf05287e61d184ead80a480f9c6bfa04dd9d8e40fbc4b3d1c6e49c2a100f3
zbdfa33e7b7b0377aa3451407ecfa74b8f99d230c1e86db3143fc424aa2cc9782ec1b46ef6658dd
zae4d009ec7c5800502f3bda3e80bae90666088556fee97af527c764535447f07fc6e3c642d367c
zf53f51570212ec4827a205c2ba2a26adc421279b5250ec5cf511f2986f77746ab2990ad64db11a
zd18c6aa2ed43e2e8993f3ddb297f8f7eeacd4169dd1ee0c64939cf14f7126e9a4ef334f5b0f098
zeb69bca8556a117fc9d06dd0988a63a859928696bd376965e0057385710b2627cb349b083c3d95
zd6e80d6016b5028d4a694486d66190efed2d33437ef2d11206c46e488b8a7fde7e872876ca457c
z61519dffc664bd44e94637e2df80299150510e79e9e2e0a7e4526bc8a412b9b582840365207056
za5020fef3f909754fafcb199635d9ce04861805336fecf50077de019052d3058b6d8669cada4e9
z97db411883adc3fdb6f9f5cd77045d2e5b714aa33c7e9f5139300cfa091c815620e3be4c642e78
z94cf5f5329af17bd6883e3da8e783e020c69e785ea9376a15e77e641df46368808ba61b1cce8e3
z86d4c7d588611f16d9df42129abe78262ecea5ee89c9be117edad7ea43d982f63025e15d6feb8f
z7e20ef6ffb49a63c22449077714ef5cf007845cb46994837c3e686961d9bd46ae79f8911495a19
z7cc48003db70c65769ace386a1c28e7dced2743deb46c020e6f73afdc63df10f327587c64567de
z615e13b2b2dd28a5fba5370128a630b3c6b5334f829375c5acdc0f43d047a2470d7444ff32a9ed
zd7d64a7fb6516d24336802ff7f04ca2fa847e04eec9e9f27f4324d1df67aca5f4dff7a151c6b6a
z07cfbcc293d573bf57d229414e9d867f67b7a2c1856bcb6231e903f3fb8a6d78b70613cf3d1ccb
z9f27ec91ffea4b39954c561fa2fabb91aef1b2725d57db0346109e56775a6f17ad32e9f85f7e35
zda4381dca06ea64a1e4d060e603d0c859681146fea3c7ed1410181f840b0fc049d269fe86768fb
z3a118f00d8d34a00d2e08a9dad84d37e4fb4b28345b73a8b0ef6f69a6f747dcb0945b271ce379e
z98219904fd261e6540f5268a6b76d3769f8a3052ea6cbb10e09f2042728362cfbe12ee3804a4d5
z140f256f9f5fece93e80041b1759cb26478511a51b9661d92a412a13ec18117b282962bdb432e7
zbf1b6b55b60b85b6ede9d5a8ec5996bc849bfadb6d94f22a396554046dfef3d3f9a0a448c196c3
z13f04b1d0f97c7f7b12bd27f603d064e696193fba178bdb570941472b371f8add9a7e1a1c93dda
zef71ccd624ac009c90fdacc307a8a13b8a526ecd3c2dbcb753279da1557c8a3c0f23f330f3654e
zdfc79a261d1fd7b77020cff824e435f6b3d328996050a1e96f00314f96da11deda0f1383cbef63
z882e2fa57ae54ed3770ea16b6fd6bf89d441dc3c16752b79c7139f4bc58bfba2ae7aac7e356569
zd258876fa47180f497b82435d0ab48fb4115eef458bce69be68c4632190e88bc7d68b2d36d4b53
zd3a8b6d324f5993e5b1ff4da0caf480494b343d100ea99668cc6d359fed3b965746fa1436642ef
z3bd28ad85b5d866b9d0b7220eef7748b71b11bb938eae7f8557b4778bec722e892b11266ab00e5
z505868a6acfdf1ff81e2d01fea24cff5d8671c56fb63f63b78dd2abf01d1045452fe1cbb728dab
z99e734f2a9aa0f4f4fa94aba3fe34019fef264e9531ddc113bb16545b508f584826283d728c455
z99a5304d447f499866a7fdcaec4050f68da9bd411f39d3295709ad98f289cd6fd13eda0acd016d
z1613f9b505e7f5227cbc2f7ca43e57e005c05bea3e81d6645bb761f3bfe12677d3b1e9c065cb20
zb0af22c91ab41e3076f32aa80115b4029abd2b3d90302da0d6c65631974fe9403c538a6a07282d
z7c1b6fbbae9395efc56de9f2d40651d26cd37b55ea2af784c8d4823e206172f60bb2217916caaf
zd8b241655047c98a1dc7abd98edce301de67721b7bbb2046bac8dc17443b782635f7252805afb7
zaf7656f72669651d4f47137c483d4274bd5fa8fbbd743b905bec047aac4ad066d48db6469f5655
z60cae68192cb08c7046bf45795489be304bda4db7b449fcff21d9c95ef5d2a864679430965d805
zbff1748b836ad1733afb446e5b537924b4e9d36b7809f6397685fb81d54b0f57efffdee0b8c6c4
zac774913b24c9498239b328b99725ab7e3fbf217925c27539ac21f8f0149e34835ea77e6ed588d
z80077f5de64f8f5afc4ea6bbf5eec6a89d5c39028eb117373b644ce2630073e26304c37fa87383
zc0c397af2592dee7fcf884c439a7b1b1404d3a6bb13264a9c633f04c0118f351e13ffa96f92901
z5e506e2bf1bd4b74aae46913179a7f08ede3c58ea381670ae0787fe9655c30de382886c5f22308
z4228dfd68f374485b3c993d3bf15b64f29ec45f1a38df9d24e34f06977e33217d60e55e116bb06
z36edd251860c8cf97b6b762b0b25f6134419dfdc5e1cb9edd414427af98c390e8c9fe96b09fb29
z824995c2b99daee87cd195140eef2fc0a56a887489aa43a3f326f8674767bc647925dcc956bc8e
z5fe7f750204789b692a823d255c27a43be8f53dd5c9ea056ad4f7dc7210e660fd27f17e1a960b7
z3055f357aea37410c87a1910c1a8c3604d7db961bcb5ac25239b840f3c24657fd3e059a5e20104
z6f1db1083f936140b1d809cee81bbeb6172ee65b61c82f9e00b7621f522eceaaa9ec37eff3ce24
zb3389fc3380cfb5bc40c6b9ef2028965cedc8924285330fa17f65fd5c79fbf0c19313419fd0fb0
z658839cec9ca6030fc9811a7178c2db3b0a480e801b5f1caf13d8c7a657c6ec27d92134503ff2f
zeb6162852b0b2f93aeed0cba24e60cce7bfe2997bb370b1e1db7885e2ddb2050ed70b679b8a578
z6702f1d31246999ed2ca41ce7e842b960f95bcf093beaf457102f14f315f67852a00356a38d93c
zfa2723725919697d58460e7232427f1f7a582f5c1dfbd17e70a616f79cf917278e319b86fb2701
zb4055eb9b1052a79120902380b84f7af3fd81284fd49e4fc8cd32d8d0424bf3514ca8ca3076247
z267fc0b6055c438e370d96a5d9fa68920955c8c4257d06afb129f7b9d18be7a3332299ee176479
z344e79412765248d31b70cfdb464b0608c74339efd15aa63191966c00f806d395334d0bd8fa38b
z365721dd2e1d425c0fc53bb43fc4ad2087ff55f95ed82562f97ec7c7d599eb953a785934182bf8
zbf3c11ecdf914232b54373a66483a903170fadce007b8817596b4afd6b08060db9f111cdec688b
z530cab45a5fe8a07ad43d288cf9ac16e5825bba02ff458ceef7e60182e65b6e9a3aa8369c2723e
za02ae27cccaf5ad3225378f05083cf9f5bdf2d456196e462562f388d7f41275a5f1c91a0fb1d3b
z62eb7a2b941ddf30a7a0acdc98cbe05b60434ae0006e5e4c39b13853d5d1801d2983de354aaf42
z74773abdc525e27a4707be248cd16e145bd18587bfea2fac3a8739f4890a6857ba28cc35b2a4c0
zcf38bc6a952f0841a1e2edbd4b28cf2e2f1766d7b4d6f534e4015704d54918146ec828de0b994b
z9ab56ba97852d6fe559da61bc34390a5456e8df6511d26f4513d491eb74127116e4cb1057b6786
z56fea9b227c1e5e6b0626d6a7336e12aaf3d820366f7c6be7bc23c25fab8babdc3d5a3495ae10e
z9780b2196bf0b65884031e727ab2d6fcfe8f64b8c401c771cef64e70e7a62c732086df608ca488
z662dc5dd220eaab7c66283cf2f0c707759f9ba00f0804932d66317186aa798876f0a5713090ecb
z17f31233a9282e7fc08a05dd61f373c31cf30303a92b2511af5da6400df79ed09ddac03051b664
z057b1c2ec6a7bdd21d5df6ab30d3991ce6880dddf0419c586f60e2dbcb2296c6624eb3bcde7280
zac54fecafa44652e38e967dba753304d9620e81301a404df125c9146af79941d688052e42bb94c
zc0c025552b719a0b28148a810b7a1eedadfeec6bcb825b5f7f8c98b504e0eaf43613595ca11b4f
z2e46c39724dd7025245af1c2500db457564005bdbb198da8c26e543d8dc0c74ccb9db06831c992
ze56a0d0c84be19d15517a3f7525d3997c884034af12b5bccf4a7ce51e2f878f296c684c206a84e
z311cdc24f6c77d47589d2b98a316314489d745f6be9161e709d00373233f6d231377039f04c95b
zd161799e7f7b44d3d3bca69a31c58bed9191cbf9a23f67f993a1c394bec5ba8abd6e4dcf0ec644
z85e5ee2ce9c3cec22f1607a86c01aa17f8acd59a2616d76522b37da8c126be299bdda6fab3081f
zff23f02fd775fe3d05c9d249a750b1abd81c9ada486620c58bc46d3a6d53cfe689190514ce73b1
z55240fec6a28dd4d5252167f5b80b39a116677e5881eab9fc1aaead97b350ec3b6aa1980a54ddf
z44a274474cbb6c3d0b75de2f5bffd889181c29f5bb8b365e7684e567e79e3735a78bb02a927159
z630eae8af924c9748b1ec265835c66ece84e4165039d18a7613bd498a1126244c3b595be03c4a6
z5c89cb6598a3cdab1e0bf4f2031f60969a24680b96d968f16f5df79d2c36f8aace7d6199132cc5
z7f838bcdab277e3ca76e197236a1fcfefe1740d58bc74e6e0af9c5a5b48271a59023e25a475f00
zd9917eb75bead79350fd0c38ebf51dcfcd1b3f42fa9051c4000131010b2390606bddf30ce4ed88
z61be446db497ac43ece2bc287ad13d6ee03c14825fac48aee97141e6c3571e89bd3cbc7eafa8c5
z3bd86c3cf036244bd0e10adc36767207966005a6ea60ac2d0f565a1b4d7d4bdfe0fc02aee99fea
zb4a596fca460dc03a0262b215741f1db39dfdff984816f10e4b919fdf9a520b50a4695df4a0401
z724258337cff33765d59de6ef9d6285d235046c5aeacd0c32fd82bc30c658b4f5cb121a0c99738
z6932e890b9b06fdeb834663ede376b6426753aba5c311025c583d743ba941ccf99338497a65e8b
zcf01908dab383a03247a2e0669fbb0bc0651951ad36c0d99b04132c03ba17693a31c335f475748
zaa66e40a701e5b9c309cdb7da98b6c22542de425444c89270df2847b9d1cf4c646f5e154e93b07
zca1a0a08552106130063a54b666ca869b36ddffc7faccd8be281c98b815bc0a6c9abf24d13fba3
ze8d62c814fcce98dffab08fedb32b0e4d5f4c2db33f1824f01adb44ca4cdc0db34a7ac88705d2f
z336831190e5d5dfc113b5123585717f79e90147cf2867671e6ab15aed39b0a5f00848d9757f17b
za0bd146ccb30802a62ff6d6837e39df5f911e5b81d7bb01970b4009b9e5958c1cdfa7e5d87367f
z74ff42c2a732f393bce21d2d3fdd60b2adb2db4790196304cf4ebc71d8ae60a1bf83595e966b11
zca3b4dc37f58ed7d5943aca668e78e74473e883d67bb7691ea410a929bb19d9aef094884c95594
zd2c29cb49f4a670af286ed86c70c8eb7894e3b77afb27e10d6b1a65951486898538f7b341cd88a
zfed1cabe5dc3eaf789ee3e7b369ef1f7fb3b0e51c0c7c94ecf097027c0cbf524e4cc32823a1e3f
zac3307e5d1fcf9071504081ead0ccc933291731461a5937784e5bc83e192500b3db59f3fe1aa46
z18f6a6d4433e8d23d1fc0a0e43b55e1a1ebeaef43d5fce85de51a31bc65f3ac12c705307de2687
za8fffe975ebd1616e12653ab0f14ff7a6d01f491fca32496fb167056cceb40b12d398b48467f85
ze328073c1230e527417a0ec03f11829e919d635f0dcf43d7146f566689e5a390107177f225a09a
z6c554b50fa19561aabb2ace25c93baeaf7b7ba6a03d7f9a87e715285f31b5bc10b83bce1bb8018
z83b15daf84de220764a44f4f4f443a79056ecf928d8daa634955d5ec77ed3c4c84705c8ae775a5
z16db64555c8bc767d079efad9d360e113e1df76009bd96db3353f28f995ab9e24446a16c14f881
z506419408369c0e636552433ff4b12ec2cddb06cb4dd891a98f44ab9e9aedc6fa197376d72fac1
z1c6924ba6263f273be08fa91d77db62a4115c02cfaeb9ceec98bac8d1f89ab47658bd0ce44c03d
z78476d0b28b369e46e690c6f1fa33913aa6cd74bb88bf7af648bcb14ba9fe4c8aa6924cae2689c
z5c96c9dcc5fbc67ab2dbf9d45a83c6c8d93bc2d02660a7b5cf48c32cc18905e1c05386485e9bbb
z10e23f98978dd1a4b614fed2d5dda97b6f2d16019103ae5a14bc8907578e4c17b0575ccd571f35
zb9a8861ddad33749d83bb11b99839213e21e832fd93ed73fbdd95ce132c4aff710e444cdbf799d
zb93bc05c6ab3f8dc2bc68f9148cca0dee00e32d6f2a8e231ca4458cdeaaf813c46e3aece34ac8b
z575d1357211a0499c5fd75488bd7963a7a234e8f38633a0bd4991fa99426eeac67853ca1a5efb9
z0ed56c8dbf21d105dbb22a658665c304f6e17fb2a8397ed70638542b091d01a6323f0a94f19d42
zf5f8088a46aa5fb6337decb796afb83d5d2116d01ba73b028272eaf2ea1d8cd97cfb67a1e81c7f
z855ad3f3b7dca2d6bf83edb87a52e08615b1dfb7de1fb81175f4b68f376d6e3a042665e17d819f
zfeda9ce4657169b01e1c0e388419f0f5d58ec443827bad8c6f3584ca92f57fddad8622433f0894
z270454819b52dfee32c2da5921e1e741a9283bbb4ef6f0ace07a2bb443c6b138ce8fff277f05b3
z84b778a7080778802dcfd810f589dffeb3b12567a95d1b014c5e5c814c24506cfadfc2cb7ed595
zde9969baeb986c42d8cbff21308c46177a7d94004d48e59e8cdc08067c231d996245fb4f23bdd8
zd1abb8a66d2fd5b10802ab32e2a5178a0b492a5b5b8743928dbd56784151f3daaa96ee470ee473
ze761607a1d6160d0fb692b4c461efb7ed970227d71a12e5e87ba75ace6ef81514186f36c614b78
z3b6de0791479fac2937906afd21b85450724381c467838f278e136442048be023bcf6378fbc10b
zf02f8a77419f750dad04ee5fa9e98cdf2f0dc59bea467d2990dbc75d0434200241461ff56e3114
z72fe471410f792529eb91aeb1c0d0847fafbf9d49b7f5d48aa1e8b87eb4bc15c84a48bd0424762
z73979f642aadbde7046ca7f41f95fd4f37c9301e1d9774deba41524239360cb97b86f27d6f815a
zabca030d5756b53d94de4140c12a5e63894698b4cf52b5a5d1027dec33274cf7bd93aaf1cd4c9e
z34c7d6f934abf14a3d6bef89176b82a173fb871f798e2d63f74d798be7e9e99cf173b84dcee566
zed58eb0f6eaecabf6b708d0dd391600866c85f26ec8a6dfb8e291a4e600d6100cd2ec0d91479df
z5afd55b7dcef18779f63cb652a156316202d40637ba09aa617e2fbdf9fbd2a9b8d5d14701eb4db
zbe4c206253445f0e203bd12b9c6bed148f2ff7e3a5b938982ef5de17ba7b2ecc6c61128b056be9
z4370cf362d2c60abe88b25a8622d3ed3aafce24c3ceb70703c8716cf544d0069e9604361de01e9
zaeedde1d9962bd0457400f2f8f3178972f81f2aee0b027710ba2b042aaff6ad8653ab3131ffc36
z4c039cf3d701deae7a8178bf5ede9a71a1fd6abcc009b81f91c38e113bef53d3526e73fd681579
z140bf0e076007679d9048efea0bd80b86ee93647cb695f04518cbd436382f403a9499630a6dfeb
z9591defa8628d955d92aa15b82ed2e9a058efff9e039ba7d419771e6c8fba0082df69a770048f1
z2199d25bcfe5877799dee65799e0cc7098d3fc3b08e0910d5b49aacdd8a32f8c85b07a95687d04
z25fb6ad8e8467dbfd5483696e0d922a6800e608fd912aa102a663667bba23e44442c981d2f93f4
z0208718a7ac22abd1f42f05cc47b784d294a0deea2eac986358ca66143da7d7a6a2173230f1c47
z7b28400ec9f3770704453d436228357dfef764ee21676954e749a82fb1583c3ff8ad254080891e
zb513c09e3c345389f1507d8791e3cc5825cefc7cf22625b8d04c4a65c5eb6258a20cb652c6403a
z8d7a84df4054dd81d8ab6fae8500f9dbe6eb8643aa356dc56c7fb854b4742ebb260a16b92e1383
z01651810a83943fbcc20372d4f7ae7e7a1a5df061dff28fccb9247d7b87b661a61bf4a8140e6e9
z1bf50ccf8a517937326c94f32eb8b0bac19469bdb41c112f67bb05d0096ef17ad1c7c86b585242
z35cdd2a818a713db3954eb3cfca4ce4a959774abedc410e6a853f16de4e1e51185fe8d4afbf24d
z88cd04ffbe1f3d54f403e9c7d60eebb29aa26466f869d8fef5ce40f20a97ba0d14ba88d55987aa
z9b1e47af31e1041cfd1bcd3c1ad22c0d9b633fd7d20e976af28369c63bf9fdaa95136554a2a0d0
z68c8aade9362cfaff2d58f62a3dc92d8c5971b53ab66153a74b81f6b31783e42d88848ce4dd0c0
z8092bf45ce51ef624bd000bc2e6c6d2d9281fca3d42d0ed9e872bc9591e6daf43b958beca0c27b
zb092cd64c2d07f32382a4cb5c1d106e1a0e4a3282ceea5e5f2fa006f62c73f1b9b82ed137f940b
z14fd9a6c78fd1d7c28177b15b326f7fcd59ffaaaae8cafe35f337897b321656b9904a0a81258b6
zf3999cf88965fcecbf88529b83a2decddae0e495a69365c9e7b1ac065d8b76d1812e62bbf12233
zab2975e7089794ee26dd78fce325fb58dd898d4b8f391c3ad7129d1e3fb83655d005461794de04
zbf6070027ffedbed4788ee7829a09e7d35fdfc36d6e82b1510763095aab0b0256718ffb13530e5
zb0bbd86f5f8d128ff8bca9d37560f2800d53b853796546710094ecfa4014ea0c694cec403d440e
z802439f21e8666b329408c8d0680f916705d2a282df163848767ef8e02212f134a489623e7113c
zc9a39929d70fe6e589171ca184aca37a163d9ba902b355870bf4e63d970cb6d99d831382dcb7e6
z6b109720be0d6971bcaeab7ce9efef6c81935d7169f22f7a4df50fca9b49ddf4e2103b53150b0e
zf559bdc89889c4ff215a1228d8bd58f2959f8e6e222bf115a55154298c7292db30ece4e92c6843
za24245c4ff21aef7d0985530d0703e6b208cbbc817fa66ee30a833bfce82def8d8eeb159584839
zfd77e3bc88e2184861b810c060fffbe93e67c2f785e236af5479f810e7557e1d974d5721cdf739
za49a5257c12407ec4ee686b2f7e1fef9eae0f0eb5dc4d02e4bc3eff03f70f0ade8ee56592cf3ba
z8a0208af33ad81c59bbe73fe6a7c1bda97b2a37214cc5ba21062b5de757e8bc64497bd16a3d3d2
zb899c233c0078e4a5563a0abfcb06621eca9ae7fd7dc4faae501132323dd911db55a483855b012
z925aef6599808803fa135ddb1194a4406e642be7fc8417f146cd7b36a875c7e07af916a29087e0
zdba3c0589c9b800c6c2264ce481035d6123478048184818bdb4a68bfa2e79c48c00e5ce579564d
z36e51d7edc20c3b52a6d9d4c50c45978fc1b5e0f9278c42ad4a084049f1aef59632039d6e67000
z62265120aea495523de6ec7befb7a6dca5cfd196a594d47dfb039171410d56b4d78236d2c5d5e4
z5f4169b50ccb8439a32fd1f0cd2f56ef9bca9bf86ed24c870621bd175ec01c1921a4c3ab7c5f17
z0f4b87d6dc3691e6f4deea372081e603e6eb7076c695ceea7721aa5af2967f5f01b5b6e9baf52e
z5257bb9a788c98551461cf4450e07042b1a6171d60c186b3ecedb96d471c494431e57d0a53e5f3
z61a222a0c892759ea83a975d4fc651a9980f1b5be2f6bbb12437cf57ee74de5e8d7f0fb42a07a7
zbb6734c4180a9f3e02a7df9e4e5be086deff38d63490444fecf5d599398294e2f226788b108842
ze5e550926f5c1a2092fa09ce1b4bd80d4507d5b8a80ee3d5ff503bf32b7b7f9b9fed25f80c65f4
z50e021314c06a2df4334747c43656d46edd0bce599a5583a641889ff098af6294a554795cc14b3
z354d2b57011505bec73e76d644dc93f43edabc0f14ee95704397f9de7d2120d063df66da56ce9b
zf888ff88f2af572d08c72c73e63e7878a63491316b630ffc71d3dab6181a45f941e44a9a50f85a
z927e36a87fee0260f4d43ec36d57d28fd2097cecdc90a6152076c0d4d4c5beb512c7f452bc1e0d
z2fccb2f2afe5e9f556cc8244bf89b175e793e9bc2b8484ecefe9a1ce2ad22c60a84f4fea05d9ae
z1b16036b6297499faac791857c1cf8d1562a9fc6bec0eb15a471246a9c9ef1cdc11e020dba2b98
za5c5ec7427ac35dfbc72edc2e0e078a9f268c7aaef7eb30144d3ccc8ed17b36fba3adb8df22526
z6a6626e421dcd7f81fc1e5432a7a21dceefb66bf5863a0b83bb0c383d535b59bc167324121fb05
z5e2303023153aa63d72c96d9342acd7ff5ed66fa2b04f439b1c6c75f53a5980187ae0d2a6bd0a3
z8b3e9475e8f07331c1ab690d88c0af7fb3b50e6ea98f0db54213a27f3a31da9f320ab2c8bda240
z748d41a609c58bdeca0de9b7ccef4fd922d0f88c0f052db0d00470cf9ef63fec1ac7cfd3909ddf
zf5277a7568a6220d1f589f94f8faf0f987ff48022e89ac9d61b8893eb92508fc66d1454cd2af86
z9ecaef1bb93f9fa7278323145abe796a7505df50aa1f6047f44b7d6dfeb346333cc9b43b3420de
ze9dbe2c6da257533cacbd556cca24fa6ea5eb2f4494bf89611c7aa20b6ae1a1075318569e14ec1
z017a54aa117f8fe8c761697eed82bb5e66fc354fffd4289c155a9d0f0cab5274567a8e87ea6c56
z397871c38571e56f7e6b5d9fbc89a88bed6d9fd04840e71d42195c59ade8cc2dfed266b561745a
z903d372e5d1aa860a745dbd432888c77ee886fdae40873c24673a59fdbbc0fad48b92a6058f92a
z9fd89c5b030bef6a093cd305e90b168214ee1841e4234c2f2170c4b04a329de94ebeb8697eb1e8
z8d30a6ea84844e3499acb8a18e7a7de7bba6ce9d4bbb445f7771dcb9b5519251f7626643761e29
z3b9a341ddba5da927f00883d69dc34a88d7d3d227b6f63d288d24eaee63c7ce1e71e7f4a545cbf
z54be5bee40e1abdaa45f097052c7e397610a650b508ec42e22a05f396642cd06350def8c8a4eb2
z6cb5eb29ef6d201732acb3346556f8216ea04e0f84ac3c8395ea87070d8b9de1ce47e0576f49fe
z4554ba974666e5803b1981a740f425028afaac7711b33733ec35bd4d050503911c6249d2f85f61
ze4c08042a6474da172acbbd30cb9aab5fc5de1f19d56d64227910085406ab48a1ff592ae902747
z2349b559a1aae1ccc5593cef6659d8ad4c49e10982f1ec6bac667fbaa5f1303369dfa906181bda
z17925cd411495f9c71d5f1ce87a81f0f5e24673c26db04c80944a11d5c050075767600c17ea540
zcc3dc4eb7ef3176514557eb34e9eb328b2c8576e92f0b0954a80010a3d9a706e075f4e57300787
z8034c301fb60749f66713bfcd79ac63838b32e8e974ef80648c9ab9c1b3b949575aaa49b9623c2
zdcb109cea4857f736c0a178b75c01898c1f33e116120377fa2ede32971692f01dc84edbff15ab6
z4266026f241d3b4f97b25fef451de58a77abaeb68dd83f378b0ea5883a79992f9f181d0cd9df08
zf9ffd2f3ec3a06c13b7ee156b3447d2788b46bce20bf4e971459342095d97719c19eecad3443e5
zbf7d03c2bbb8654cf77ee12ee8325c526e57d9f8d453c49bfa73fc68279d09bf0606448893db8d
zb47f28d4496da0eee260d72f9ec02b66112568956b7c502f72c3d05fc77ffcb2641881217f1c11
z577ac7b5181673257763845775bf04fb45622074d4a2af9fa5af36bd190e19daf453a57b8392cc
z30dc2bd4e6dc56ea4413936e13d93795203b3e55e4b1e397be19c10122747297c19c9d7e0f5a34
z2b361772e7676721f18e98e19dec729641294ff28b1b9fedc08e37131a2cf0b41fc776a39c677f
z00e21ccfe0b08f9914ca451e92e93c5d1a514bd592d067ae5198531af84a0fff6aaa18c5e2a9a1
z17fa137bf747f2cf7fd2f7ce4d97e0743d1ad49d3270ddfd2cd04ebe37838163dd4514f3a0106a
z06e777b040754767118ba1185617027936f7b49b7e729383e80e76a5b6c303a9b29f9693227b2e
z324678637aaa5be547794554078b7ee25fe4b12aee0208cfc6b4a24d9d00f2fb8f91af1f893048
za78a6b6b9a500176906889ecca5dbe3bab2be1f2c169030c78c055d3da2ba567fbc2f8adb2563f
zb92748610484c356f1db1b682ceec345d880aee95795a11ce74bf82c163340837a9f4e430b01ec
z77e866182fc2cfb804859d93e777fdce9a3730bb2954e9e85da5632098b368e085090b6dfea1b1
z77cd019cf22e62a791d5caaea1aeb76cf384be6956c07bf2bad367e67052baedd8412600820c3d
z8595dbe387431737f7041c7bc1bae327b141fdbd4d3d4a39f41f2b0d4be9cbc08a36e47579e3cf
zbaaced896d265a73b1046ed65e3935473217a16ec109d3b39545f242d5c121b1fcd35812c5c5f1
zef70e91c93f7b5ca2adf1d8b5623a9e47e6ecf75efee3cdbbe08369d575e7e8de1da76917b0f01
zaef1588684ac452e059a153f2245c0c1ad127f28dcdf135b9058f7c0e3b9e15f789a925fa4f05d
z306b4e48252febc45bd22bdca642dbc9c5b38b593061c2a2fa640bb9f15232923e7a0f4dca2fb5
z9c594b15c18c3674635605d293b356a1e9db0b68241d42f78c098baa6c625d50d1b4bbb3a29d56
z8aa32a91defcd9a1d5ec6f3bf1b0a9964248c84aa5ef7541dbe723d80b0cef8b73d7d99d224bc3
zb88ae5b60b86c2933aee65ddfacd55b0100d7d5a2045a7ca22512cefed2e247a848ad9b5dcefd3
z207d4270346c5756ca7a705aa77bfa0e0daf2507f4c3c39555f6140aa57a9144103433c389a234
z2a1f1d3ec265f19473e5261b24c3dec2d14d39699a2ac5f31990f183954d127a49d8cf5e25324e
z90d899da6125e6b653de64b5b21272e2f970e2ef0473466f0b90b288532e46361a37a963c919d9
zac92b4e4dc539d1f281a51e8d18f3efc7d465f69f20cdcc9a8077ce128ce6a36b7002a3bcfbe25
z81430870a9b4ef0a6c6f9490d33f38f78d70ea13d3df42d555f7dde00cb92e96f3cb2737c3ffa6
z379e34288b88edd2ff78cf8ca2664a6bae03e0f98dec6103fb28456b7a736ccac98100be5eba8e
z3cad8a62f53ef76504f9d0338ef1cc9d5e7f744668cb694fb5b144c7d4b90d48922ddc143ff8e7
zb9a8d24e2bc197a6561999ce341e09619b0363507e579da2142774d02cab393772848216a5c916
zb5ca0570996e61264abbc52951f492451a27cf755eb67b6b7f86d3eb0ec0b7e480120ddbba7768
z0cf07dda142bcf7f232ca21101d3c32bce2104e90e3434530bb398f5acc16bd7c27654d551b581
za5806d177970f99e793d636adb92c66e857a04eecccdba90d1cbe2b27c3caf13a7fd76e2f720b6
ze6acf7a09cc0748fbc1586fb70e99e620c7ab7382c3647ea207d851d30b0c9bf192db62782137d
zefbbc312eb29ca89218f6e0c8dfa3383d2da083e68a1b8691a36ce5d1e6554024b72a7a0cf965c
z2bb5c1c30ca87ae378ad46751a4e554e3d884ba3f27c384040e244094d6613901ddd06d06d0c90
z1eb7c2602e77b11091314aff4495584ebcf99c19262f042ef833258b8a5e8ba54c57f8bffdeb97
z0cecdedb2c9f005888c131c45b8213357185d040f155d2e9a8d977352b2d8c7002a7ccc1bf50d5
zf60b70037428db60767d1bc5f2e384fd39ad107ccff2bb921d42f148fd5b6ca6a4fefc2d8aff20
z337c09a61e7a23aa9dfe5854fc99d7e6a9e3d5a1c917a73b071ef09d1bbc5241b64f41381bfaa4
zebe134be51f1379e4e8d43ec6dd0cb7abb4276888c1519d989d6276660d889505e1a50e19eeefc
z42c61c2e74c072fefe84fa62e61c0506cf1b4640f0bbf36fe8212cb35b0a53e729545f752af0e1
z7db05b166188fff11b26e31ee539d863d7b45589e3441fe574b4b94247b0700fe9e78132b535a6
z670a176f7167a5dfa35d4d46325161a63d0c4e8bed9264b2e5c37ff6faecd7f4b61f2324c52d53
z3e446575e9768f6b1c8aaa0f6468f58db1ad6821a7c8220398086b6dcd509077ac48cf2a1bffae
z55f9813bb627133e17b988000f012a48a098d302d5712a938315cc011887cbbd963d049ee1a317
zc44c52e8549bb863f83d3073bab56bdf3c53b747c10d845da2e18d999240170a9a23dd97b6c862
z21688ee2d592a4f16f213347bee196653879953c8b170825cb2c0216ea931b39d0a8788db94666
z1035eb3ce1c3bffe70eb604d29d52ad9c3cf43d89a43ac0ce2cf2d81d8bb2e846bb4fce5d177cd
z8075a063293440a5ca7a0ab8bd61d6d6e1ee6368d1f45320720cfb4956922c554ed5825bd071e4
zda6e51b1cac5468288c271813e04ba443878dacabd39c4074ed706d5113c77039f827fe2c3f1e9
z85df695e4c2734870361448d7552d39d1676dd66c072c827d75942097b00240ebbb934d6a930d7
z25a64d0a3c12200632018630967030ee671f901c826d910d576031a1f8669a90fd5499b01d93b4
zff9004af5e50f21c49080a696f4e8a7ffdcaaec20e4f0549605d609c3ccdafb1440987b4026898
z8dc386bb7874f5b0c8c4293dc0e39722e8a0ce9003f9ca74e4b9cd6501231f30415e5d7a6da551
zdd3805e25a9eaae1993d86a64a6ed38b0d5755eb0a2a841ae2dfd7c69e70019b7b9f849a3daafa
ze2c98bea86fc17f8d3111924df1b9e4abffab47fe8d0982885b5de2a0aee40d1c6ab3c03035364
z7944391abd64094b2400ac78bdf1c7f7388de96cf746e9543b1630a27aa7fe9871513f874f23cc
z7673153aa1d5cec1603f2917d057782c16d61f0ecbe9551daaad12cce60128a5d188ea6a2f6724
za3d498cf108940a4c0cd9689a3f5bae0e3e07dcdebe69f67cff35570415aa966d5c5c711978f99
z98074d6ba40f35dc0bfadfe96434947f1d3e9c2b8a412fbdcb88539bf805412ac2086c552da149
zf759e1ebe8ab7ba6b2486727cde82c0216b36cf05ee79012a691a8d4b27bb6322625ff76e59ce9
z61b37da5d49437a953edc51fb2d804c3b91bb15be7f526fd868504b5dac5568e07c5e7e0f61d60
z682c9f09e45335fc39d769b349ef2e256729dfc2c7f2ef4be0ac8b7632417839613c9ab384984c
z3e82f463d41adc00efdf9ced1b5bc934973ecab7a8b5d316234e25741eb316421072cbfdef78de
z482ef31a75af01139c2ae5541968abd756f5815a27027405bfb6a5078f4064a43b4281678481a6
zda4524df7fd913d3fb8b1bd0a99e97c1752299fd4298c64d94a339f154c617b57da3225a257f1c
z0db31723896283281a63674183b30ba2d80998f1447a47a8aae44177d0a70284c8df8d401dd503
z688882093505e4468d28837fe6dc04a26ad5a5fe4e65e7df6a0fcd038f415564ab820908b06961
zfeec75ab7af7946bc0661ac6acaa6c3e49225c5166c50f67bbbea983be2eafa8167610c457964f
z44f640b2a8e022232c0dc107b80104d4e341e59a30686e55e863e43465c02535613fc66651d08e
z76167ad8ee4654a5e71130c8ec681a38ae3a614812975ad31dd5081498cd564ad797a51596ad95
zbc89b9caba8a01650ddc590fe316b0b0b548b30fd3c0a51602f10c8df6e8e7e7ee1188e5cd9637
z2e013a8985b6d956a5079242796495e36259ea6b39a7bfc030e7a63f5e23c230e884085ee52420
zad1fdf15479bab6842e8111967c671d97a69b5611855bb80c4ee1dee08d696c8b9be58ddd628a0
z05bcb4af4a9336214f66affb00aa7c5669e9e4a312555f783b4a790be9531656ee954e08a0cae2
z573f5f6718e0be0f27a052f582552e1d738c9fd914ac052b2ca39456c5bc72e6aba489d559eb3e
z204293c93118f62f743d6d9ec6e46ec539f2150a661b7757915d2a2b2633bf65425080d9edecf7
zbc93633710733e1a5ef646d953273d0cbdfaa42106de39b2370bcd65d8aa5b351ccc21d764b964
zf4c566f01ae70ff3eaa36d7b7ccb680433e49aa20539bd93f52aa6e922aed8ffc06acf5ece7f26
z88bbabfc21b43615ba8de52e1802dd54a5cc0d07e99d08c54860d26526813a83daa5dcb4be0e96
zf374cca3a8b7e08696330430c12fa0e0d528fd130240611bc2524d33fedae5a6b8557e79f319b7
zd591515c7ec77397e7cfbe596dbc8d9d09b3bbf9712b6a0dd702acdfb361d385e890592d8f657a
z7eddbea7cb37c692478ec9dca05d9d893b4bfc67ba99be77378da58008c1b3ec8f5302ae89103d
zdedd1b663821a903c23c31df5434097c5d9595406f2459d8ed7a3e95f8aadecfda23542ba35b97
z5e1dc4114db8d5c3057d564b89ce72931af97bf15878376dea3d842e4e9c086cb9294f37d5e6cc
zb9305876ee366e15f740aa5640e616905639f0beeb9e7e15942b24fd7d3125a83e295ee85b4ea6
z4298f0ae8195bb2f80d86bf32e152f1ba352c9c968dfbfe19f474e89faf8b32a94cbb62e658d84
z6553b54b14c4c6a53cddb65bae199f9e129c7bc9968e788e8519069a47aaec53c745cb3d955f9b
z6a5a6cf32a09be79c6835db3af3aa29feb0456485cb31491814d776cc2773f842caa92ce349355
z7d9284edca74f5d081b9e7693271a003f311b673e6899abfe09355cae5f52d991976e768337bb4
z10de7f2645596ef8d204731b48d8b7ced82893bbfdafa12bce67fd833b6d446afc4a4605c5e034
z554d53dabd143c287ac32349cae11eee939391c5c2bf5b65961016dca8d7c95d4f21bf2169220c
z320f2f2e020d5b407851e290c29f24baef8a097474e1dbd7ced9ccc0b9acc5445d64142e5d0cc5
za2782c16abb6708208e98284b903f5bd2688efaf2f2847ffa6eb80452d714a4210cbdeab91815f
zf98cd262071c95cc0f4aa7c5cb4375236712ce3e60adf6e74bd8f36e25aae90a11809641549438
zb1c668694e6fae14797bece651d8f6b3934bff09888d69fb0229951a0043a01d4e01eedc709111
zb300d0f3027606baae33a231005974d0d760b6084d59f8ac96e9132dc6989b36d6948726e22f08
z69551e8e9177d9d8f043d9c6518f2bd38cd67907cf915877c2b703c242354e851e38f7c85c95b3
zf2bb986c7081dddf004faaead3c3cd61fbe53fd0d45bab1c7f2e680d30513fd2ac7705dac8dd87
z02bf33360e09920dfb65c90c4db107abb16dffa4ba726dd49c3a2c1e9f696f42488efd5f70b7c1
z0f865ec8e7412eefbb3b4690ac3f5b6067064bc7f9238c795cf139c3050af6c06fb33c4fea2c52
z4e3c904dc616744607b94013915b5f699aba61a000dad3328d552bdbe095a433289b7d1217e6af
z22eef5c49e664972cb1983a0aa6b2a665fe8dcd34aa1e0d7a3e5f5b13789d2c2d26981328bbd54
ze130e090280b04a6cddf0c2527e4f41dfdf0f367782a96050442405ef6fc4dcf1c587c0a4f45fe
z17e052a7816f982bb8fc99c9390738f768ee0df68163e3d971842bee79b8d8233073972800f356
z0461dbc83c74183659990b4f85b62ce1127f52d4157f431f19e48b1ac21381a9c869ed6ff49b07
z05ec33c8f3c1e5aacd4ebc7e22d11d183ac4f25d9d1b755b2a093e685080fd431bef95cdc65104
z20a702ec3d9f7bc521ec2e2953da21afb5f779c914d4345588fd2d13e53efbbb1e8e358e45edf4
z56ffad68853dc700909202d788143e24cf640e11f4955fc71e648beadc9b7b149d3e3de57a73a3
za9ea435e051ea39eb9685aa57d665375d82afaeace8a7878d1a8d0144f20af5fd5e8364dc8e35e
z0f467d7fb63783763ad47ac547cdb66dfc17d1dc9e98a4022652236b0ae2cd0b7528559c5c35aa
zd95aacea1efbffa42773bbea30f688de2b15d4a61f70662d04381f0fe2575eecfa41951e21fe31
z3c0bf54fda7bd92f7992f1b41784836b4e9c45725a71d5a7657d1b73212e07a392b40a6e6be97b
zbd75984c5c00be23a23ec67ea58130f469cd7168dc1e3347f11ac1d261db7eca9336d4898fdd88
zf5120d37a80c5ae12d56bbfdfca3da7e99848fffce0ea5c55525bbaeaa935580d7bcd8eb32b87a
z7259d4adc1df289ed0fb3133f4955b92f8ebac78d283fbe484c8eb9f5dfd6306a55b05dc765c38
zcee74dfa5cd68aa33637ed7848681112c0a1c5b693c39d52fe770a9224f8e2b628a41c96453c91
z868826af5b96b73a28e833ec0417a8edc984aed2a49ce6fe214b58e861f2a19d90ac30afa52c6e
za741c9c29d84712c5f6eca454906ef5c44eee662a03ec90766fe962ec88611f9682eaaad66c218
z9c4d4490fcd0626e42a5e51071bc9f8848d37936fac8c1ee14b95b59b3289f359879d05ab52979
z2c73f09b861e3eda88d97b7b58afd08a517456929666d7b4e7839294385c194e52f3fec2140b22
z2cd9778e13778cb5bc4728bc48fcab41c1e0b70a1bcc14379c5ea8a9c6bae7089927030c3cd5b4
z88fe8eacf5403cbcee7ec738bee901ff09cfa588dce6ca7b7847895a5d4ea1c060279dd3a76171
z0933bc0184e1d5dbbf61f0ff534eba52fe0a8590182a12eda6dc42c909176550f7eb3a09e17277
z23ce650233c87f98be0f8b7136b5efbf7ce60de9fb36e2217b5003b196ca304dd58d28d07229ff
z199ca0f76d9f477f285582666a9251139870e409bd5996c28b590b419a3a2a718adeb485297938
zea434bdd4db59767aa42db38ba7278c889ec51568a3cca5dd9993c4605edc16f5d8f1e20106123
zd00b1965b0db41c0ce9851f4f8beadd71b7ef062ac20ab7bbccdc422040759d349b16c1a3c337b
zc08f2f95205089662fb58bd9fdc6396a0a50b01cf0925863824ecea87cd040eb523870905c8f7f
z779e2e648c360fbb84fc9ebba76ac88dded84933af4680f730e2d0a7a5c34da54e2ee4f2285c05
z1a070c0689c1557ff1ba8044b63084ea4a156c4bfeee285f6094293be50eca931db40a1b6d7cbe
z6b333c8731e92e85ad43df4a5ace3efae060c1aefea4c074607c26f11297e63bc19971aef65421
ze6cd8439f126d0536d2f986bc3d90f82f4757a5d0f46205f99c83888f544bfe43c5dbc575ac209
za8dd3581ece48bcef026fa4e992ebebc6c44425a83be02fcc63e8ff666915244b57db5de0246e1
z720c1cd8b5b304df75aaf67091573af18ca54b6e71c19b20b06476237b4cd1e889a3b20791aa85
z7d5f22845f0ca1f4b52d1a0b563578491727131b62102593b342cbdb76c20f84f2de992e553596
zf1932d01b2828bae0ce4f2ea477c0028ed378534f385d00dd5b38d12ee4872512b0a9158182a07
zee894f445a10e5b182c8c35053c2338edfe94db51d51d8f4fc6b31518b4c8ee841867016987a5d
z33d5aee852e5fd822ccbd81d709cdb10a0d04979ef6e70ba637b59ebf9a02fd549a4df0ba2f5cc
z784124ba191ca0e537534e36adb4d34aaace818f33e0606e85bd1b98f5158330de3c951e891248
z68c5df89a2a396e0536bf7271c30d64b25686e203da5e06606a0e5850021c9e9376206f27b47fc
z04569f01e020d9c726a2400af346d654856efac909d5b05fc59ff6fc4b42abc24993e7c0ca31f2
z01a1386e05b854216413c69168e147fd51f86b1fbb71a0786da44f666c01ee03f2ff7d9448241a
z288c2ad3f275e8edcc36440075d33e77c07edefa6fa5e9b15a0bfaee7f78cb650508a06370a95b
z24c47d62df12c026bfb14f964d46a6bb59f59bb9faa658745dcff78deb4edf2784cc6be768372b
z98fe3c1bad3d12f24473ee27928ddb53ca27f58452b6cf31ffb0cf05f3c67b53dffe7cf5b3b0ed
z563a5491b47ed63cc72ec59b55148d9ab23ddbda68497f6ca939028ad377a394683dbcedf80964
z99ca873593e2d9bb7e865b3762d4ce35f2a302f81b43390712239ae20b6daa88e64a6139a52ab7
zf5842e4f734ac5f65c5a7a402a2cd47bfb40690d73f3d84fb272a40e26f9546ac2d80c71bd9e3f
zf4e4f0cd91152ff77a625b7fd69266d2325fe042ed29e45f85fb63d6d15a850e1249a5d0ba70af
za0f32765ff1afc41789651e15c71316a0f5b4f91a5505273c7a14bc2fdbae4dee4c439070a19ce
zdceff9869c857d8dc93579b7f8425457f774076d72407326a39d1332aaca783ccd9225e4c981c9
z3a283e158078ab0d1cbac7c7b5fe51fa43ca65b09be0a8ab3a2868dad14f2d37637f7026ee7d20
zcde727bea3149c6ef5f84a5414c92503a5fdabe04fb18b1bb36fc972ae8b3cd73a8454a118e665
z2a86f1e102ba48f20a1482616e0246f7ac3e24f2dca6f333deef45af2a6541749632c174a9cba0
z6ca7ab1f2eb2ffb2959a9dcfafbf38457dec2a3f7d09dd134a7e211e21d5f2b4380270d60fb2cd
zc9da7f02c4d09ff9353c380757d072cd3fe98cb0e0742251ee0058f25766301bced9fc89f2ec4d
z72cef9e037edc6a0a8b1b8036b5bbbb9d37a60cca0b9a95f72cc74b18fcbff9e662fa2fd50a3b5
zbe11f0d54eae4640181cf19b618fa226dc66f5b99d67f5ab66aa307021a2aff87231080babc782
zc86ec5a4c7abeaaf62c6881b9d30268a7e800889639a7c40b4dc2e3326eaa7fd949300c5718aef
z4cb88e2641ec85f2f6a78a32696177cc8c3b2535aaf71c697dbbe7f55732c01a860df8d5603819
z233ec70a99fa4cc4815229922bb9715c4a21adea4728cc6dadded8fb3abf21638381ca78d74b6c
zb34bb000bc6073e94d475dcac01325799e1510227bec43952174bf4552e0daf5ada00d7bcae2b2
zf0ca88a13224ef8a38df67224d4bb7b3a03ef18d7fb9adcebfe5f814ab57536268c9b0de37530e
z916c0bd0cf11a6f81acb22ffca513bf1d17e3eee7ce4cdc6c468eed0123da4c261fee108ecba14
z8b83f3acff885187e4f8ac92fb8a96906f02c757232398cd19f1842bd265daa8671ead3033959f
z5ec05d7cb4a20d64ce7728b0a58f73184d59f5f9d00f613011a6d0acc2d0d81ff122621e60f4ab
z2d1b12db7e669275b94afd16fc9925097930c505dbf3aba6cdbd913c792eec8f6ba1dcbc989339
z961ec0681334f1d2affe2d80c463c8ec4a568aa08721f44757caa4ee93be06569839decbe538c6
z93e8dc5245914414ddf593c53d00f5a0989b3dfbddf56d2f6ec816a25496a97e34541a237fe0e2
z75ac294693052b57c74ba200f0fc73bcf3be704245b1252a5f23095ca5e1c442018fcdd9c2ba38
z550850a50940244ef4d62460345b6b4dbf63d687a3da85dfbc227d0f12a0a8c2db24b9de89eff3
z0e80d7927b9c8ccc8d357f9b6881719eda02a1438bd9571e6f4cb7a014ae9604180039880abd34
z8e795ee162913ddbbddab2b69afa350591e8de108666015ca9d6ce3ad89650e4103a8a78807ec7
z5e5324f70decfc37b32211e214929a18f630119c5de13cadd264575dc0df17cf150332ae314d00
z107e1047a75c099d12a51368c38fcecc7e262b872c2b4badea618a838b2fb67e16aa6355800d61
za1105d04b57bbaa9de00e948081790197f3f991b069a581de1734424a282182581d034ab02d7a7
z7328bca9f8946583ab78329ad476dd4f2f377c8e9234f6f5cdb83687ada73b442bbbdf08f1be3e
z4a7b24f73b388b0350d374774e9a46bf31adbe0b88bf4b79e3fceffc3ac74bdae54cfdfb9c93f4
z412806d7d94e9420a8feab5d17150ddfe92d4de3bd3888ca406fdab1b28f59065fbddf5f2d3884
zf0b85ed621ba73dfdb2fa6633d235730f7bcb5f7a119753b2ac221f3246de38e67f861cc85cd78
zca9268b264ccd071c33a698c5c6f232d01fcedd86ca6cae5e0820e9c137eeed2dd0938d0e4b9c4
z25ec41131f28e81dfa7dd7c53f7f2a7a193569f67b4b6e73b547f3db96a52d6b71b66d0d507b45
z9dcb02dc480ffae4e38daa990b8e4f91b666b1ea337960d7a425e3b66c57c96cbafe0320bfa02f
zf3fefac84c108e61874b1058e89b1c5174de126644a50d176c4fa30c8f45c3226f9647422da4d8
ze709553f65a0a0a4bc76850f47e3cdfa30ada4e7d2ef4419eae2e1b8b5a316bd02963cd346566d
z2d576bd595b09c650dd42abe0125fd2e984c00bcba79d70b23a7271d409b55fabb7230053ff6a0
z57c5a956a081c74d7fd252ebf58aff6a1e1758caf6069133a2b4900b776d96011473b1b10a13ee
z1ad7859a5f98a04774bfdd0a34fe0289857742d1e2d85671122fb99aa86e169b91d28ff7fa15cc
z151f3b25426ddd9df7bba6313ca564f3798736c8fe949af9b7df40f8c7df42ce08786a0a55a36a
zff4f84af82a1196ac92ac3e1fbfae69ce7e6187b5cc8b5aad7e78bf1f1a816ba3fdff6d93c0183
z83e6bdb644cc3ee4d132e5945b1c03d4b0ac2df0171657d4ba35077b47cbf708c2cb0264557dd3
z33041e6292580de43f65b576ef7aa7ce7383a7ef6597f2bf887a42ac26ee58766f2b5feb668fd0
zb3f03e547a48e9bef62f9684c5b720f474f4d38a8336bd53504e6c594b099d77ff912ca79a8917
za1e72130e038b7a0ddadc3af4cbf3b82c305933cea3edbb8c1eba89f320956a80a591c9c73c63c
z67252b45fddf75b4943e0a8fb55516b01c0ecb8dbbefd618b7a1b26940ff77535d5ff08292f3fb
zbe7d1f2804aced62919b75f43b1e02b8c4eabedc9772974f0ff876f3ed7ad0950b470e4104b261
zbb5665bcef386f861ccab6c8be602f71bf5adf4d6af13788726af78ccb4c4aad2b28a5bbbe2075
z77b38ca4131edfbea39b41bdf581de4b2e46c1124b841ad37bb8a4de906987adfd6892bba039b5
z3cc046d2cd8737d9b6c11265a1c51201d1d91e35608d073513cea2902a1c185f5cbf1532eef4b1
ze7fca156ff17858c7ca92de9e1a72e3d710d766b02078a8e3648575edead7b2155fe324bde1b85
zf2533ea5b95ddde63970996d3719abf315a6ddafb0d37f5262fe98dd483a8a4d4eeae41d13e40b
zb0d452dbec22586eb38dd9b0f2fe06f4def0b0a21490ef17e89f89cf08abf5617d105236dfe043
zb92d3d2137cfc7737b5f2beb992bbff36124255e4b6e4a541563f36bee3f943f27643a1a80b2ad
zf26e47c48d518e1fdad4ec20d5a44fd391dfa082ee07fda2021f274099d641e9a0582800bbe22a
z48ac6387898b8bd0f1aa7d7887bc044fd7e41726823b7b52a8b47cb503ef4543e1a5f9c862b09b
zbd74aa7b2bef3d0aabb6bad2463e7b668e7ce105dea80336d16063d78fb9c96f751c735e2c3b55
z7bcad37891455c78fb4b61a3c5c99233de0767c939125820c51ef1978ffdb0eca6236525af40af
zf2fc9496375252c75ced5995e94f68231d8c71b63dd57f3537c6ce8800d9b8a5749594f79b1897
z48028b690ed40f5f5260d8b50990e95e692e43a4594ece7fc95757641d861ab8c029fe4500760b
z8e0e6496a2937ddae15dbae940cc9567a326f2bf7e08654e333d2609d62a0bdc01fac5e9ca3d83
zafa8da479865111ddf53cb318340f5f11fa4837192ae8d1e9e8e31132ae2bd1142b023eab02313
zd6f842a3e34bc676ce5df4da3c7c51756e69d3c038892521e5b6f26399a87cf02a859e36c3744b
z546f8366b838843502d02bcc096d2fae2ff2cc89b063be226af4ca600f787d836d8cb4ba1269cf
ze0426ba4bedd6240eb830271a009bb92424fdd6cf703981f1e0577c6e4c6a7f3e8463aae0c281d
z749afb513ad9f8367d06d762238492e35cee199f55d983eba2b160ee23a947c011a82c26cf8538
zcc65ee48e79fa06c8a03566f9e60e778e34ec5d3d7533d5cfd4472bed53cd39d4775f73788b3eb
zcb59f47f9f0f5fe407a9be8745de90e1c50e7c939a01bae828339928bcfd01080e26b5d3209475
ze33ed2132aef30da628fc36513f00466b4ecd2829f99933211e836c9f9912fa80707369ba27a5b
zfebe77be136a3506e99598ade8d9048c8ee25ce0e5584c06c5b96818aa86a728a60b7ee2759d96
zf77b6c964e67e81e143c9b763b4cec88d18abd8442ee6e182f0c5bc89b39b74abf877601206f8d
z2a7367e2114ebe7d470160a5a0ad4b421a8d63c170ad65d5443b8fa8f036c4c0d3325bb3a772c8
z648af71b056df3999fe6e2bcf2a9023a5cbe5db9de210b16e3d19e4313ed9db2d95e17d77c64b2
z38282a7825f7c2837ec8ca87ca8962fcc5d91ae879a780a8406db1bda7de21e7cccec3d17c5a97
z268e76e37f0795e72ba0c3ff23ad2677a1fa359b71a45e970675e2894046ea853093a0044d6847
ze2a918a06606a18a0c69f883f12c44c7005da90d054123112e2bd273a0eff441c7d3ad8dca90ad
zb90f2a26e64fa249add9af08c1d81511a581027cc6944ccb5ade89a4c231a54fa667621d86231a
z1dd00208982fb0af89f83d2ce01657b425a82ff58ddff89dffa5924f02c03285f902476f3270ed
z0a5fb07fef5d94e7dac649c7f5d804f4a69a9bd245007e8286913e3fcf6fdb99a9e85194207914
z18e861a75a9983bbd76951248114ae48c4c6dea9face036385e28c5a731ad1a2d91c5f71274d68
z174d1cf8dde9bb21187bf5611722c44e211fd2a16df9c5fc198dc0c8bf7db3c0c71f5d469b73ca
zcef8f46eef947ce8582bea137b7bf29c536f52973faddd652ec2f8931dd68ddb8af37e524af041
zcf5ea62d5f00b56f01365a9eed03a519f8bd76c2083a48e24f9f36a3d363862529c7ff44223c7a
zf78cd4f5a6535041c63c75cfed472755f22c6cc2c3ac73af7d29c344caad76bb56bf1498c27bd3
z3b03cf76f0b78803c97dd88ff672b0f3f35ebc1000b27d6a1a850cf03d6aed86f2df69fa211d80
zf80f8b6fe65c42b93de3703703d6ea32aac4b10f1783dff940b081cdc06f0bf13bd17de11af675
z7d6aa136dd986329134b2acd8d8f3ff96693bd29d607371f7358d6ce104684a9c46820efed3681
zc7dcdb5450aa90103da7172f61717b6aa841c35e1b0425766ff64037929458f679726e62a9aac0
z390f5f2b82a19de1075632c0b8fa2e8334634eac1646f614929506f144630ec44035f60eed1add
z763c39d3f21c21f5c20bf001370cbbcfe28c32af34c146b80fb71d8caa9cf8c53387eb9c4d2dfa
z71543dc942fc69f5b0eb7db512b6e18e53242cd724adb8232f8f4124407f03a5c65a9bb729fc7c
z2208bd50219751f9697338f860e8d978c82dd57f9ded9403cf06f513d0c4648f97ce88bedfa7ec
z9eabab1893814bb0c7412cb874c17cab7d76c856b2031dd9889ae7e13dace37999714825ddb5db
zcde965f0ffec25220a0be39d3e3d7e8676d3217cc667a1b205ae9680a900b7181b86f42bbc2ba5
z1feca7879bca0bcc7bb20e2ab3b09cbb419c45fe40bbc8d690524c07fe415e1ad5b2eb04b4877e
z174e734e57e9005597770383248f29dfc3cf607f64f45b8805a16e4dc4145587d2457a1a8beeba
z45dd8a3055171a290dd398c3b24706e539e4e049db6e14e2ec8ce84cfacb6ead328d9a846558cd
z7d6735e92242ce6b36f45cdf443a83ed011119a0d21f94e18254c94fb69330a8f605d09f117d69
zd4a3ef2f6db26ea18df7e052bf0dd3d0b6c2eefcf905337e5d9a66bbae5a80f4287533b8e3f5a5
zab7e80fc4b1a67d5a1bb128416f5a323501591604dacd92f06655d1da5c62162ec6fb750959d7f
zb4b900212dd7c36040ef12cf15c3fee86f32872b7ff97977d2c311bb9cf4ea7727a4ac206fa2a2
z7f04cd004594656094906721774532944d3e810e3e22ed00c5735395c1faa492bc0cf02d74aaba
zcbfb48f81ffaf3d1616945a5ed04a99a724abd76cd3760cdcb1977d2958f4b3de8826da8f07369
zb00f7222d4e705b87d3f84cb02937ed4f389e1fdeb8453342b4376b9805d1d375faa9ac9aaa5c9
z9513640e3481bbf81a347fc9a828da1265fa6dd031c32f2633c3cb568de91e442039433f5896b8
z91a3074ad9db278833766143406c509a7e1c7b7b74b556e34e89d9cef7351aac45b09e8a12cb7c
z03d7e0289f2adc70fc196900efb60e0157528c41d12224a214a46fd424890490713307b29dbcbe
z917e52e0f8fbd01e55938b483642c12466f42504f9bab4a601da25f3b30aa3ca89caba908f640d
z80db69e25f27ac4dc2a0fa5b26a885856e570f9c82d879e79d410388d3f59bb2543e3c9f792126
zc9574dad8c51b7c25c86a95cae2f9c391ea673f0ecfdacd3e55047f76959db25c6577a64777d5b
zcfd6cf877f06b016fa83ee40dda74b32a05bc20ed0d9f7dd9e8e65b52d3d4e36de87718aa89395
zf422b6f397bfd179ca734549e5e693b6f0f58a4c198a6d6c7070a4a3d67a1613aad7d1a5010fd4
zc12a393769bf78c0b2bed92b8d5ecca9b1fc0f4c2e160d374648d661a0048c537b5257a1255d08
zf956bd2df38e4529fb0611b6e865ef131e44e7dcc212a5e2a120e9208300d19d980fc49e7a8926
z0c952d18e8ad07ab4a198494be1566eea195c534290806d894819f95f8875a80f36cf12934b6b6
z6f87acb0d38ce6187ec7b1cccae3427ce3a2d0c5aacece95c86a5506a763c91c75a24e4967caee
z1522b5dea0a7eea4255c1e4f3027574d01dc29aeea9a29ee78d8188643e45bca45883212aa15f1
zb8798dfc03fe562df54d13776a91668ab27edc32fc3783e77deae89514224fc4a935346ca4c75b
z6585c5f5b4de53e3e5638d74baff1e7ae66affb740be2e39e19eeffb72c7498c9e66c6b2ee9c52
zaa6ab88515331ba5dbfa7ae439025a4dd283761e7b6d856735c5099d2db7f3e3ebe242012b9bd2
zb60cebb020439337c992ffcf9a8d221c9118d95c56618369a565d91b35c7ab593b8f55935c3320
za40bfbf870370f700fb31c32c0d109b08bef36579e3637dbb835d61c3f554e624f58886eb023e5
zc442e9a78df7c234718b59186d79f2235ab83f20dd569741234e3ee3ce5fed6f0608069fd4c4e6
z907a65e500f47a9067b0bc408de94871bfaa21e08ec2dd44af5a729d89998ee12b1b640958ae99
z3e6904f4ebf8493b11701230bc3577de69a7207d4f93c242df952163bbc7313b27944db8ca6220
z5e2f02ab7dac6c35efba3886bbc552d4256156d6b7d3038a1dd2f176ddac5b36de735a41e51502
zada5267dede4e9e8b132ec5892b7c6d057d17d221680ce15dd229f2c4ee7dae3808a85ae044a6f
za39fd627f55bddee69fbbaed9442d92dbd4cac39a1b0b55ba93da6ffc35cfcfb738c17017eb3b4
ze64fc0c42498c4c05ae1345111a8049eb7239f8738faab37d83f8a1beff9494850c2979954c6e9
z1f3ea6e712bae914b3f96ccd4a231c047a06cbc33bfa7b5f120de411d5d981db19c44de3ae2c4a
ze312e35c0ba2fbfa51d95fb216035be9927d40b3f8a346d8399f01d0b8a8efbaf7a1d347449500
z7509561dd4d809c3c924443be422b0bf2f3ffec8f8c584e77691e85fbd29ee5d0005142208d3fc
z0d7008e5935f773e505ab617b83df2997abf91af4b5c2a2c720ad54e1c479afde4400182fb1a69
z1742b5698386722b16510b31a9473e7982e0e615ccfaba2623b1c39809c684938237a98d23c996
za74fb6201fbf026938649ecccd211a6731e1895a263dd28c5a7329fd08a9cc74bd1713e771f7d4
zc12bb5b4df6de978b55293d5ed824dc3a7fdc9cf7ec973aa8677c58601cc1dad458b1ae188ac7d
za68e2ed913177bbd1f4540644a61fbb29eb1fd6dfce14fa1fa7cdd92faae49ba0e00c2fbaf18cb
z9820d755c6fd28e1e8e54bb7034e7a256212a6edaa52306ce3e4f890443d4773a49e778c8ceee5
zc62ea63d5316636287da638b8af0a49007caaf27a9ff5eb83ed36bab5a057b1089a4f0995832ec
z3eb2833b51ee5bab0f08686e22e6c31e8b7e1249c5508937595e5a64ad3e59ebbacc8ae3109162
zb4d1d7c78853d47e40a59eed6d4c697c24c4bbc6a3cb0d307a7bff371e40eece900fe71da5faa4
zbd9662619a3419723105a0ffa90def4e3fab690f862c71c242c23bd41d01649f12c93297ff0858
zbdab12f0db26ab5035989c4e449ad38dc8d3a5f6811e930c7d73ab840294bf878f0867de01cf3a
z646dfdb342e7e0520857672b8ff1d77b2247734a53906cc6f8f5189ca512e8128a810e96e4b107
zbef8194a3df92ad8c53a7dd8b098a6c1bca4bc549cad657cce8ffb5c6d36d1b41ec33ef0817130
z7f185d859422eb68d39a464cbd6a41c6d814d4a5b7f940f394ab346e86d1124e9f3914129e4e41
z61015702f60d8e85e0b468a009427dc8a9df354b3bd1a5d12fe446aacc42a61421ad71900b49ed
z8c87fa5fa70168302771c68feddb5f1d4fdca47cf43de6a9c70877b97134ff997db05617395a96
zf98b398b7d52c39d400a7a46902498e7ba8c1b95a006ff956179d2de2c35d1fdf22ca853d5e3d2
z28a5cc9c444a60fb699494d9cccf179b3fee37c944894650139e40d21b1013078dcf95ce40caa1
z86349765c0c117d8d22436cc0be0c669cbc7af38611d49679978236a842ec2b398fcba3d491327
z6f2fda74cc289cff072a5d6fa4dd96f317a44d4c9f6290f7d65311dfc91658d4fa9e69e595ea9f
zc71fe674ec3d4d7f7e533c19a329bd6af02ca7d7ff963de5e21a58c65666519861b8058cb3d626
z6b5778833b62353b055a87e796d646a6799b8a93dc02cb9482a9e093b72e5fc4f76343f4e25dda
z86ca419b6e33d491c3f88485cdf585282d2c6149accdd0ee5c8fa42e8fe24eb43480c824535d35
z8f24f52b1de20b7bbfcdcb13c20ea19f7b7ab153a207aa5d2819bb6074dc12318872e083711c3c
zd40f931b80b1b9fb03964074ca02c2619e11a56949de272687b4f6e1a7da15860d01705402febc
zab1121918370f4e81c946bc6643449bfb5ce32a096048cc41edb307cdea800e7ef1c1926505bf9
z03d00c698c3c15e8a0cac41d4aef745fd80501290a60d42a4318afa64f52d61021ca935fec189f
z1f061d7dcd9e841b7be5bb8abfd922ab1da2ab70709f94d4662c1634a435b0a382cc6be178923a
zde5f3b8e89fb18b1a7a5f7bc18cb3ddf4fbba36e6c821c29bd549af6359d2d1126687e494e513c
zf478ab2491b8e0f921a7424a7d196474c85769fd88fa297f4713663af6989b83c9c388fc7cd5f7
zb721402ca6f4a60735f9419c163350b96bf216997e56622a89e53f7ce15414afd070fae03e4387
z06b4246aeb859ce9f65218e66968d8aeec30fdda15342511dde8c627d770c6b2a5cb08ecdd0a80
z58a349df23e89989ebb2eede861c6359776ee10df29fd5194572f659e4c43c57d86f6c432ccd8e
z174627e34e4e97aaab0a815802afa51801b60845f3815c700eced7be5a451b81d6660f54efe7dc
za5d4104e3e87e2974a63ff8527a06b2d3850419a53d2bf6674f2c1305a9bbc199a0c1aeda978d3
zc450772381be4b1e43078851b855e40de43137260abbb19099725c625dae64f7b43e7455fa28ee
z600a0afbd0f10c096b72fb2d4ba1f5f7a4c2b3924fdce8bbf6ae7df22f7b019691261091fce1fd
z498920f9c0baf6aa08f7c50da652f2e60ee55ba59fa73202906a6957985f75f72f522678fb3612
z98ee639f024c440ccf9bca1aa9b9ea919bdb7505aae80922970111b7d0780cc89d9555d6c0325a
z584796b14c9c42e82a209724b01f7cd0d7bf3965cfc248bf3a32d0850e183f60bc73d0e3d15bc5
zed515838cf81f611c994cfefe7d636481e995b94d479039dd4863c41778728b2aeaff9df1ab2f0
zc31485c74838c96b96d7c88ca1c5bba37b822fc05c0e920853413284660a0c90ed39ac51d67335
z608a87b51d8ccac7bae9d58ee18e92864488a88472ae2e37c4c8b5aa344d4aa66051cc6e8ef004
z40a46d305bff7b06768621cc43aa70886f1188c2812add9d2221ed46c5d9d5aaeccfbc38777a24
zd7ac1f4a2812eb4bce6b2eb7be18a76cdc2ff269d050285ecf2b00f7c869476cf721a2972f4798
z4a1003b7feef04f2c82059109407b389199859e0f557a3d70551f458ef5a880182f18ff8f74ff8
zf61f15da430e06b578845bf90b907ef3269e860516593e8f60c6bd65faa194ffdd2b08e04117d3
z360403f74c29b14876a213fbfc64fc19fefb1dfcfb9d35f023c64f924298b9fa92eefdac50a09a
z1b7ab357d1fc14f44c3c788c2dab533ec6241f0d3d635b486aa5c9f484b5beb4a097ac9e79b226
zcd862effd7eca853161121f4e806a1479ee6efbf6c59ced9856f99e332705abc3b2eca410576da
z61303e30c2d6c2878b4faad5787b461334b3fff342f65efa96aab936624ee2b3048894a5850588
z9edbb846503f573568a3de53d8d69078071e82d14c3ab3988c8d763343c6002f69328c771169e5
z2f8c04e8647b48050b5d0ccb274f50ec50521cd901fdc7e34541e0d8ec17743ee1e7fe3c9945e3
ze0f719d012eab1b8de7de02e9a6671fac1dfcb70ee99d6bcb431a2d2da5c9554514828ee197b9d
z3721d32657f4a339524afa74b24c31661eb31157c06b2228cc3e27f3c81d48372bd5a708c2c0ec
zd077f93c103f6e5898941c30821d0851034305ba7fc028e5f808d6544dc544857c6cbecec9a416
z93fb5a3638496bc8900a445ab9580f597cc76c1a624fb6b843d09bb4b51df6612495094dc84d64
z58ca4d016d004416ce33957db45403ccd71a128edf67aa558a1c4a7682408ab96adbf87f5092af
z5d6e4cc1d9030d7dc129cc9614c8cf0eef7840678cc2e22d85affd07bf306249bdd381896eaa55
z798ee05761063b2bebe0e6506e987694b4b4da0f40d2afe6ea956519ad1702805b6576e2fd8625
zb6e7f4be4d00cda1b34f360f55437a8a8e0a7374fa0daac2b512b3ff5b5043f369cc1925a152d5
z51219db43f9070c3f14fbcc4637e185bcf4a5f0cc87e1d67b1dd194a58dd7c70802c148c09c091
zdae4d10fbb341a6b05a7add88935ffc6753c6aef9544ed5897ca9dc9668099fb6bb67d5e009b59
z56b54f1ba160429778c4a6aa3db3f2fc090970eaba579447c30dff168e68dcd784246d3cf8289b
z68d0f49174bf92e73e38363a933bc76f962454fa081ee515fc5e18ef8b31614d2f5bffd3e35506
zfaf3708c2eed90a5e65a38f78a6123bcb9b9b92f39f1172e70b3381fb81b05fb095c6df72e4733
z31288ca82940b5e45be3bfd8b4b166698ebd2879e95cbe549866a335b1756b7197d2f93d307a42
z2c5e454374ca25c0224c6faaa1b056ad72f0f99269f806be92967884ed64272de685cef152f2e3
zae859c961d93c093e0823ba4a18020f40f8eeb691e00cb71a1a6e93c11920cdef975667c060029
z10f3b9287e4512fb6bed9a17edc0aca9cab55393685c1524395515e5521c63bcdf25d1130dea7d
zfdd4b129d9095352a14df0bf4ff30882da9f81746508fd5c2155eef028997a4d9706201571e6bb
zc60d475ec2bd6f4198be5549923b9c55d14cf61b22d825733e88f0c41fe0b66850108a727c7c4c
z75f80e33acbdc9c58e6db81e3cf21b027341a054b7173f543a6b55c80a966398989b7b2fb1d3b7
z38cf185fca741049ad42a5f4888fd7466574b17339ceba9ffdcab9f41815a9e69320f9ce0bdeeb
z9ac4b0b88df6dd18c1cb887b794e2890efb37cd8238c7e086bfceb26a4b6df8ffb213332696e33
zb8116ef302f9973cd7f005929d37ed3c01b4407e9c7d7693eb8c467eb92ee0279f1fbb4400592b
z9d9264a01f2adb5eef80224485a1e4ce3ccd6dba6feab67661465f278e7d0abf3e5645bf755e82
z16604ca30f2fcabbf54b9606e955130e5dc6effa7eaaec28838f9d03b17126289b7fb56360b4b4
z91c94fa7cf9713d91b8cf0e8ba1c0d1d693b7b7c1b580f475234f1d79c372db15a8132c50424ca
ze5feee1997e9e290f1d53109b4ee385c9653b0caef68a0e89eb937696aeb54123510c7baf822e2
z56820a4582f50f777f5caad2fd6220f7db711293765182a49912ef6e0d51e70993d16e849cdd6e
za5625a1497bb0ab452815f6792d6c845ed4ab8f7b9f9f935f40f0ce73837084ba960037251c1c6
z18c9958e27e2e08d07a07526f793005ef0acc423cbc3c2eb07cad99daed24ced12e6940a26b357
z2975d11daa86d08728ba119f582f67968ac0b0234f224636608f944429c156de87248d777202c8
z6753951922337722b8088a5476bc630667f37ea1f29157e42ec059670af11ae454ca5032f5257f
zd4924f09fd9b7aca0b60d2dd0fb16e514c535fb34422fdb4921cc5f3c904809f0b3ba1468f3767
zb2b7f50ccc7a2d6674700665dda6d962969b653bbf24a225441ed57b7212ae8dee8f4535b0f8ce
z5f173f49f40e991d68d10ceb724f3a1a77acc31f3b43b7968ac0bf0b951896961357c2b0e38897
z5e7186aa9d1765c03de86abb1cddced28c95929983b97199346adfe53e1ebe1b5927b38d24b3ec
z1544b50bf86b45261c94dcf2112344bf1ac142dc8b7461f426b8f745153c8a2bc54029a80c79be
z93dcaf4a84dfa54ff3b5130525046feb1b73ece8c20e18739bd4008fb3f55cb2ad5a5150cdf090
z126a2baacb1726461b5481b9b0cd6edf387c65ca7bf853c4e97ffb75c55688b538d113c7f3afc8
zdf3f0d6123b5d0122e76bcd6fbb1ea08e74b82264310d44dfcee95bc8dc9eb716ac72ca89f7804
zee91d547413f57bf85f73a5c09fc2e4bfe443c9f2008dc5b134759c72a130e1cc5dfcd5bf83952
zaaf4c099039320fc80c0389a9019ffe8e058f50154c49b714f3e993eadb4eedfe2f9136312048b
z97c014b3c6572b0bee48e3bc45453c5d56417f7a17ad9d763d0a2da5c49358f2d40e7a1616ee5a
z1ad750bb8f4db84418386b73fa95cf18ad99d1a0e71c201b4d6b03601cf83aee91397dd751aeac
zdeb0bf25ee1449854e4ceb52f3cdfabb8dda510c52bbcd7a190f74ff5719116e8a1152b13a762a
z60429e6e12b5a3b6660e4a538afa1cbd65d3f1d48f884a8fab4c211c89d329c2386ea950a56fc7
z0cac6db7cbf57b56f0fee26b5887462ef614a83a872d6bd1913b7215ad68e105a3a945164f719b
z74d4ff492a4c42da05ab1a3f6c8b37f9464d96f7b1c4e1877259c2a0e621293c9d78f563492283
zd76f0c41475e566882a551a457f328879608a2cd1f251c52fc2cf66c196591c0143f66824f9eba
zc983d3c3c84abaab37948e531d9c9a45c2e2dad54bd971ad6d9d39b46c8e9f5a46cdb47623e6b3
z32d1537df0a582dd8686f2f594703cba69e5a19bd0ae4ee5895c0f9a671c387400aac54141e8cb
z96cbbad419e211649c60d085779ff702be609f842fcfb707e0c6f8c1d19a49dd750ed62d05defa
z9363a481100fc44d6ec1ce3e2bdc5d3472b5023fadcd47fd1fc1090ae70730e3a90761f53d07c3
z1f9d516380cf7ddeab8a7b8b8f9f3e9b0e34ba4068a32c1bea2d37e122df4cee3f754d04f90edb
za71b7c5f5147b3625bddcdd67979a5af586db5aead9a9949e9824cdafaff75540de08832b03e06
z6d6315e8ff21a9d996f6558afd4b666cbd956ec9ddc302f97e5c0ddd16f2f941d193b345a45a68
z067eeeef9e866a53d19c7d2aca58df5baad74ea618cd77e2bc66a99a27dad5d853ab2d59cfef12
za633f1d2cf042166392e3ab51f2bb917733e61e4640a3ce87b5d8475438e3b1f3ec29842896695
z4792e0e556f061b9f3d86a6762d293b37bfc240ef7e62cafd7a720109e5f394d1a36585e8123f9
z9d51061e44c0e9bc9ac9e9e1c1d05c4dc96300fd53cddc8311d3300e81fa39626c312b1fe08eee
z9bb8aa19329e1b8b5e7792264eeab2359006a7ab5bad4250ec04cdfc3e62192eeb2bb072e934b3
z3833e9778dd54e78e62988c6ab8d5517f050b4b745ee0c91260bee13cd0df40ade9b15fe42fc62
zf2715331baa14ccb3cd990f1ef04ca3924193d04ad5a52b07567769bd760a0c96c3dd38898b2bb
ze4bec0ec78f128d8898c50407db160aadbd1eb817f7ca241d572c317866cbf05603ac7b73b9c2e
z087c42bd771a82f5bcd1ee1b1ec625bc08a4810e73bbe062263d9a8b7cbea353fd8d3426c761aa
zdac319edfb41ba26e1c5e5b8a147e0541b59c10ad850e095a356a4f356c36e85ae022055d004c9
z3c502c9cbf01645fda77c7aa37336fdeba391fb0758d4e1f2dd283a880b8016abfb08ab230881c
zc3f09a141a15cedc38229b520255cec41a75f638a7747d191ee83e9732366d26b4e31cc3afc564
za36a2024ef7fc4211748794e84611539767af0eec01a718291767278b5bac74d863cce3928df93
z6b69c57ddbeb630371f83b23d07981b892d6d2fc2bd028952b54a8908afa7c8fe049333872c112
zff58904b1749b44f8e9b1bd4f1985d0d2ae08f91b09aee9230cb59357430ed30aa5ac46dc346bf
z1570ba99a59df578900e83e81f4c10067413a59f41e46a4321387d0ee846ce7fc5549f1d5b9197
z4df478ebf76f163e63c3077536d9ba98e84aa37d24038de111390afcacc320c608c5a6f45e73c5
z9ac3ccc23ec0b033c5ffb9670290f8b6b1896bf69f18c39faf2db0288ab04842d654aef2146703
zbe36fd0e0e58ff6e0fe43493cb4dcfbe2860c2f65ee9eaa624a99c9a74de2074fa7e5a62f871d0
za8145643b3c8103a36eda663fd66640fefa854d254ec982d302e6b11c2a05f1b2e23b897ae7efe
z8146310e99b8f00b8cd8814e603327bc9d3dbd37ae76f24a30162e8a9bdf5926c66bbb97005f33
z2c9b7dffb71a6b27eb8025a37db553e95f60bd8770b74d4438e769c72e069ff7b450ba9265374d
zeea04d2987207b8ba9b9899efd9ab1899cc0244596e9d6b8ba29db0b86d8188ffe941e0bfc0d6e
zb0f7ba6085f5f14c154e36b13d7249c7a39e1336045e5c9988e472b78440286175f58fa0ebd379
z5d8813783dbc15aa1e36d66365c10d088f43d2a9dfe4afe10c244e8b4ff7d82bd0b9bc5e908a41
z1695b8a5de65bf8a27ac324a7bf4b478f803aa0326d3e08958aa4a057b1b9972600fc427580d25
z5c5cfc1b749cedffff67aa9693ba115856a0d983fbb9f0a441f37d94327a64aae9f94e6b67760b
z16b76c70cd7745a3f643c1f2eb82933806f694fd59df80a36b7cb07d58385402ddd6d19ba84b8a
zc88561c3adec0c8edcc845966a2b3e59aa18ad07cdfd5f404943d72d8fc448ad1201a77ffc6326
z4e394f47493704e74f24692532332e675271fe96b5296eb4de9d0adc7e333f72534ac2b18b1281
z3147aa3ce7012ba74848d0d250e69a86cf668832d26bd07eda6cc4771c0319b3b8fff475ea5469
za2ca72bcf43d943936fc5e970499759f547cf8e2a79b86ce9cd5b2af31678d508a7536bc6516d5
z68a378e549d42d3a992ebe05fdc84b74b56159bbbdb31f36791e1359a7ac6b856ae683c9992641
za78bf3899e20664565af3e49b8be86a59a5fde6e0d71bff089af5f41b0ab59d0d59af50d93831c
zb2907a346790bbff01642b574ec4b1d94d47c2ca365b63e761d9fdfdaf7de1dc0904dafd4957ff
zdd1e2b859306dd31aea2f346b7f0cd01b81f043823a934431d43855be09bc2b7a48e63de403dfb
z4c041b325794ce62b820c8ce537a6ab6570982a60fba6f32c8c96d9a74d31e7f354d3700cb1d40
zecbe8a092e77d0b0c8ab67ba9c12c48d531d42e29ac908585603acaf438705c6075dc7dd1085ab
z9768f22bf9d37e56c1f0ca69ec040dd7187ef62b546f4822c87c2e4d24bb2560a3f1e77a5e3393
zb23f7a19c5bb47feca840607e90dfe4933d7d1faedc9625422b5c038e6fadc66a629703f817c74
z10ab58aa8ed361c20c9d8d3459e96f53fab74088639d3a6792757a2f71239784722ba3abaf3bf0
zcc3f4f1d1ea7cc78d96a94060f9d7965d5a3dc3738bcb1df203662389b8deeb39358bd728e97ea
z10a38def961ddf8a6fbd07d37f30973b3a629caecce14f1f066454af8f8cc87c13d3666bf5831b
z1f1777a167e77e6356608ac932c55f07f026d5e52f392981e66e6ec37a7d10438bb40de7e36876
zbdc96ffe52b104724b9c7cfb0f3a516cf3c03adf4d747d5bd70c2fa398bdc4ba536ba455783215
zf039a64643c4e213352b45ef9bea4fd61b2fc7306684c75154ff293a2e9141fcdeb4b8bf1c034d
z678e69ebb7e630b8f56784088ce8d559ae56a4fabb96ac58f041dee205d18e9c50d72e29d2198c
zcb45447bb94c8fc70368fa5a64c92abb4b2c27830a4647e4450ddd2f123afadf0958921d64989d
zf30db4fcd8a6e4f1abb3ac61f4825cc0edc40d0af3343b0128834ce4ffb7d7ad3d5e19f5d5a29f
z0cf3cd93e165226403f8765f57faaf6462ada7b70a8e2faa9fb697f68509466d72159c891aa85d
z029f0e0a11aea176ee53ee8235af5f10908987ff6c4a3f0f64ef1c6e53ea20751244ea2ebf7cf4
z54b576e4675b3b960b2fb381536a28e208381e1a404a745f12ef48c292692190106ee12995d96f
za7af8dc8a69411e71a51107a43fbf3fc44b909ade0eb206d7ff131bb6be4ce335f0be022189885
z8c39689b2e3e0ec7d43909103accf2ddfd9386529bcb0b9f7ccd4163f88339f5d37b3e7132b76d
z6dfd6c3a370dce7eada0c3ffd391a62c5e287b9a5610679621e67e3f4a4e094329188031fb4306
zd7064ddc66d6bf2867134fd7841811a9390bf02ee889e178d2c3313e233044c9c92000c9f684c3
z360c7320ec9737053e37c45e3c8457174b391b8860888518e032ac733aa9699152e91103e8a6c5
z40614bf5c40f4dd297954a284dba9e48635e8c375836b8cf227ce3314c819073b9e1d5b2a9f463
zc224f1c7a58c52c24fc4463f54eb5005638c5acc4ada97e3b8342c08bca719a2e60da1b206e356
za6f2d315b7d5ab430c0b2137ef24e0900667f9e8888a286eec31fbc3c85017a9b24894d752e645
zcf376eb41c8f9f85c0f67e133cd74059e4a4aadc2c18815969ca61fc8698c2268c00b3c8e6bd8b
z3ee7133aed78db3188f369c5d2c3b187fdd595ff0cde18b00d9f98e54642101490d0151566dc31
z3d114d144e436876d89052e80b1a7687facce32eba9be779311ea4ded6d2bc413f28d0cca39a54
z38b4827eccef8ee92709649a4cfc263f25ed48b7f3538bffef49dfaed2b7b7a4a3511b0c52abae
z6b3f0bf3c61c5a2e732bcb2ddb6478654408f31ce2895f254849ec59546d3619a0b4e9a28183a2
z4eb44eb7294c8a32f1929ac5be006b4630221f831820af902e90aed64597c48a8f6103c858e50a
z1498525456f4c3e32bccf85b706de39553cea861fac3ac260fc633ac9ed03e4e725089159bbb6c
z792f62691ba7f88947a124999f7954637cc9685ca55bf714f9d798c6fc6df1e2e913c6f466b667
z6ed3caa086f616c89d5de6c6c0e512e58be0703dc91c16de1cc99950a31a352015e7125df5fa55
zc719d3e44749c2ba5498f0c10cf7ac4defae47eb91f02872adadf9f69efdd4cfcb931fd3dcc3f0
zc4515bdf48b7abe1884d88c613d90c646da691d5f4c5fb55645f1f42d283721df22567cb47d09f
zcf2c443b00df31655069a138b8500903df44c37fd1f03bca8b3b187996f79cfca3362e460b006a
z772b5ab8cef9bcedb631e3d535896d82d08c9b2af17962e3838bafaeb96ea0f2030d1fc4515ea7
z24dac643befc379b4d05031cdee8182d82d4d70f1f5589a3483fc2be75a861bb58359fa1666cfd
z9164e8dfb77bfa6b7cf9d3a558d3485c17bbc34adf64692508e02775ecf23285113881208ee5cb
zecf6c6635d5c2af0a4e8b272cf41c74a113dc48814301f05da3b325f3e1ab4ef341492b6e8a70d
z42948b0bfe599a729e4be70efe6b6bf7ae3953ea29fa04563034cf965cbc0380e75d03fc11e761
z5317053b01a1855730e08bf846fbdb9f02e7df16288776597b2fb38b7a09e25cf6b0e91792918a
zdfb59cc0de96999a07eab66461b3a6bf4de91eeefff39d09e909779221c20a1842b503a2e9e678
z0d9a6512ecbbf74c69b42077f78c8572a5e6289f82f1737d722499590d0555091c4d64149e72cf
z62d3f65756c3cc4498fbde947415b5034b80512bacb39db051d1cf68168024cc5d8ae5dde2fc66
z729f8879fda1a845280df04d722d22e4d2fc039594b8ccf42164a90a849ce41398f33603e97969
z9ecb8bafb33ccee17b81e05a2a83fa2ba2cfdb4c52bef561a5aaad5ff90248921a10f77db1fd7d
z965b10f3359bf73db52af4d192fe119625681884afb24086daa497fc15fe3b83ace21c936fa781
z8c046cc2f7a6bc553162aaad06e03a986591b5910b5012797069ac8da82ba3fdb281d97df4db6f
zcfb221bb4492347389eb8316e70a518982c7ba2d75dea5dc8b81881549fbd371938dc7f2097867
z4b79cab152a5fb457b8e481e7333fa44188b4d18824874ff0c8ef1b9e8903ca1c6cce55edec386
z5bd9923099deae09d10aa840ce08511aa55c81202542222683982e4fcbeb45f1fd19236f915db6
zeb5bfc5397741ffef2168312cb995dc65946e984eec455da9003a5a6f277c71767e80549f20fa6
z20573b11f0448e61572ffafb03b5f960071b144eb98de82741d91327af8fa3ce80da392351322a
zde379de98294fd407792d21de9a30e8a4eeed7e6d6407eb3ab6edbe75bad584816b8eb94e363a5
zacad25341072bca723e584b5acc743e19dc91aec05ded389d1a1842ff74c56d4d010a728bb9484
zcd580795ad977b535b6328339aa8b0449a33b939803b6ad245a98e581b5c21b2658d26adfea061
z387a6793fb0aed12fa6a4ccd2a608c137b12760595500ea7cb7adb0ae44b5a066ea7a26f246334
zf6488eb626a5e0f4ca9df84d77827141da211e2d120f330b4785d49c718a029ee994a6cf8bc41e
zcf792683244aece73b6e49996b5c6d2098b05a17814ca8cfb46098d1f7095f308335ac4f68c418
z872741616c5090cf4519ef67167c853932334dd1d1d69da826a5ab1ccb9b7156b2639ce6fc4c02
z9cb57022efe125e62e6f5fcf7a7e741a59d69df8e9619e6989c61b422cbd6a9c32035bdecb9b43
zd836c1b29c23e02bbc8b2a33320ce07e96f7490f770970225e6b7a470d7591d4c41cb39d2a47e2
z31207a94d731d3895346916096289eb270190407c10869682dbaa825fc98866188a2507bfcb5f0
z819c3a9ee0806e9d72ec591bee59432ce729e34244a8daf92ca291ec61ded21bfb0d20af36169b
z430f71ad05e0200911f60bf2d4b9c6b9109270dd2063744b3c0bdc9dcb9655405d8c39fd10a320
z77e7fa2dc84b142eb600d08db17896bb64e8dafadb225fbe1a77ae6a7a0b1944265cbd3860f9ca
z505f382df476aa3e5f35ea493bf2e041684b5d650cb65ddea3edb5e8619e4fce5687b35c70bac9
z56107bf555922b97a660640a5b4dfec79f19926b7ef22a08f2e8b8ca3695a03442504427db8e14
za7a07931478e6c7eb310e99ebac374a99bfbe62b6bb130d22c099fb9f006013707f6e851dd369f
z88a55262ed7ebdce9a65f7223b06788e5c36e1cc31523e7824c18e3402a58591db4d97392e97d7
zc8dc9f56881a3ef1ff3abfcfbfe5b239e68aabff6ba415044257a76f6976034aa443bb66015bd5
z1ddb55acf0ead9046244bf16352ff72c53d52c790723154f539d9c4183c3126497c2b281bb2331
z0ef26c5a6f85c3da3447077bd61bcdc18c7f9f8f05b4c7bb167869748e66b2a479b21c234cb2f0
z09ae4bd6a14a6811fdf8da7261323671465c91084b746eb72298316662476531bef7c88ac1c578
zb7a30274032d337851ed9eddda4ea5ad2d9d549be80db7fcff58b1bdecd0160f87b5042b502dea
z24851e5529dba30c76b8b49ba73bc2123514cb78e32e7c158d352b66cd3ad8e790349b170e2ad1
z76c918e2284d30cf7b99bf8c02625b70cef932082c84682d7cbf960e1c087d1647028316706998
z2f361bdd5ef4133425c70455699da1d110c532f0a2b3b1059a394cd216e51470e306da9f4fcc88
z1d6ac9d59f0d12527d867bf983a70b155aec6a2d96cb6fece157b07164e6b0eb5e4428484ed74c
z67b8462794ea594274e2f4a9fbd8d770d1d94e3dcc137a967f79fe7cc9bffa461b14d4aa475e1d
z8f308c592b44492c930fc0f1b789203c7a6e02ba4ebd1e637b35dbab3a24bf7f70c8e32fe73805
z6d0729e6a11560c9ca9c6e73264f0d16f62cf815966756e934bcf3cb12905899ab95516c2cd218
z955084aaaba9fdb92a5e13d5f97f60356684fb8402b4efa5784b4ca65de072016a0cec8f998922
z11a61f3aebb407b47967562416eae90633646308f46b33e8c54a2068041482f55b187790bc1f61
ze262f39956a58ae6ec08e595319ed7a6304e322eb3e5d8ab4b8bfe62c46565861d6e16aaa1ba2d
za7d42bf5a8576b9f4343a45ff187805684da5a37890a4c56ee6c6723bc21b41d5db2463af32682
z104c6a3692e6d5635b0cd3063db0a9debddfd6867cfbbbfbc4166c499830f9eb06e7ac1c0aa2d7
z2c1e2c04e13738a61f4e37cbed27d3d4ea2a1c31afb5ebb4638c1e3f355a2f24381bf54cf7c04c
z0363f83cf3336b9e90909d49b40facb1f839eb6cfed853fdbd8efe463d9fc838eff9aced7d26aa
z5aac2e6254e005d57649e2b112311acae5efa39951a745bf2f1eec67777cd30286fa8695fe320b
z65daa998efe90c33720584111737a1602cc863efae27d99add0b0068ca48c4f3d27d71c45091de
z379f4dcd11425ad204e4fdbc7ddfd5b1fa51602fe12b8d6237f4cca1ef53b42a4e7800c7db9637
z69520714f198ed06c269a7c6a6be3f18aa3699c16b2a6b9a618b1b3a5bd77d63bb8341400f9934
z253067e0ef9953d908c0374b905c71f30151597e78448590bc7ef99c76eb63eef2e10dd1aa7477
zbf28a9c3cdb5d0552fd245e64bb4006fd90b42fee7cad5eed9f3ca31f08033d859a391b19cdf36
z74077aa3efb4c38f7c97b8ab081de7361c470e1a4067fc5d6fd2f30689ea758fa04cf6662c24fb
zd5df0fd8cf39044efe0e9e035bff0ae251a70c98444adfc7a77ac3d6e611483423db7ac444c6c6
zd40adc791a299bca3a04edb2eb7705c23cab3c2092d858aed70706eee46c7c3516ff9ede38588c
zb5446eb3b6ce1e87d8a0fb106721c4b29050dca81922abff9816c2c32d06aeaa99ad8abef29ab5
z8afe4a1bc0d071ef21f0585332635da409624e209c0d04ff9aa9769a767af8a1001b53d550c110
zfbd4f93f7ec0b74b189b6fa2ad08756e9054a1889cc8230fc9b97196913a4f5009b4de205a5178
ze64fb639e6b25f5086ceee2130ac58cedb2799f9564d09470b90bfeea39c0d4b7eb196a7fa9644
z5cd9de5075698f9c9daabb3b9ebf1bd462b2220e6312821ff5ca07cbc3501aacc908326576c27a
ze333f5a304336c7c0e71c527fa661ea57e94bc6b0791bf4bbb312df67a7627977df5080bf2e30d
z1be2b7be370d538dc3d63d83e7580d0288e44083c39a775b9f738f48be1f1bc065b6a7f3bda390
z43aa576d69ab86fb32e298d441886a477f44fb193cc260cd72848110bdca151f2c07bd25592005
z0557a839d09c9276b0c6a9cd36927392c3b9000830a22eeebbfc6dd263016419bf33407d25f43c
zc66e25bd6ba3e9d510fd645d856fc221f660d9adf94c775388655b9db80c5a08d5b8ce7a11cc45
z95238b71ec1416e826314eede48be54dcaf082743aa2fbab75cba639ef5335e07de8026dd21643
zd7196da4445d5f13442e0f15e2e1bacb843c415809fb1cc12317f3f468dba25f36b6d78fbe5137
zd1418a3fc1186ed41eaef883c5356844d41f506b933d63564ba0db2313ea8fa5082fcdbbd9ca55
zcbe50d27c20bce8a4d2d0c8c312d5907fba2286a6ed710fecee633cf42e0ab88f5822399456ad7
zfbf9b6d0b9265db1361e516a4d3b7c843ff9f509a8be1770ac4d0f7d24cd471d1df1379976c7a7
zda36854246972fdaaefd8a926e6ac86f56173aab60ba0f55464bea756a890ac3efebe215e5b6c1
ze27aa4d439087e9b7e13dc4a042fac01616ab8f5aad5a07bec436de95a5a5bfc01935358a2160f
zc225f363b738b670cb187b08a11fcae00ffada189a51d84ded607d836af59c007298661c77ca17
z42051f19e8647a210e5b37ce029106d7bee73bcba71c802d0272d79a002ba1cc20aee074457246
z60c33599b352be253dfb922a23504eb36d143ac1a79bcf31279646058e94ac401fce70083658e8
z8036132dc74b563925e34b542c1c90a9fd6e2dc9a2d34901df1b034161b183e55d7791f0086478
zdf8812d577a59d68a45cbd223f71be1b433c7f528e4cd9c56a99dcd73d58adb0486550e73675d9
z5713da790c76a33e525765dfc4282f783006c24c6d46d38640eee1ed10b5a79202dd1e9dbf0a79
z99d8ef00201a211d38b474c3c33df13efaef4344a2674b69fb12428a0c3c4e5a189a4e07185b3b
zc1d8df64d20db957238032b5bcce0da519fb4fb8deaeef8b6469069506a9aa07449c5052838052
z54601617a1f89232816fc62e868937b725745acb6b539d94745195faa26d4f2d4cb85e9ee487db
zaace5417cf99a98a210fc847bd7b35f5ef577c3df0eb609be5844a8f144aa01d5eead06c4b3a02
z89adaeecc2219a9d5e94ee98cd317028614145808a218631c172ee422a798368df38f296685aec
zc3c62a3079faca17acebe99a67b871cf21e66ef5b4616387bfaefed026d1e0e1f77a72e8c5732a
z754b8605dde3f891f6a9d9f4633fe062a9e6d963731caebebc5c01cec685e6f8337a7cbcfa0d40
z3ce926d42f6a7641bd21b4c9b3ed810c8bcd082c726f0eaaff896616a6d5ee8efef867a7c0f57c
z2f6d762bc004fd61c0f433be248e1d9c537996c5c8048c86943d871861c297c0fa0b48f82db4db
zd772c3b6d2f75da609717ebc494c87daf790cc289dfc4667b1885dccfab3a61084e2b6baf35b48
z34b34e05da8b09428060407c608312897af874a1f0f10b34ccb1e406a874c512f2150b94cb2ef6
z38c6c24c854fbd699d64d32f6e9841e4c29300cccb645a59b5cb55dfa554bbe10ab2110217316a
z14f4a2caca85c7e0d3485fc60690c407ed2856c349c5cf45a631d61174638d37b61ffa3461a16c
zb47427ba4cec22830e88ddb73d0b0f8a13909b1a817cfc31b0ad65e584122270771e8e19b453b4
ze9689099f1a88fd93715361f1880b3410f625f260651dc58c841280b080cc9fbd03e61b5414a8a
z503ff471ceb5c64f508286b41e46f7fe6047df085378cdb8dd3f65339fbc15715c039757233b47
z7585de2f8783bcfbad7273129b9b7fd02f7e63576a89a12b56dd423dce1f8f10af3b7c44101926
zcc5d4031e0908be426e774b2a13bd89ced9447fd782ba26157ff3ae15ff1baa0cce950e6d85f0d
ze0e6f155e4d56833cc770e4cb412660b09e2194ec0153cef89d1c735363d65a45d22edada6d5e6
z7a2d8adaaa4a0b92fd38d24fdccfa9c9b02425a6a793417f62f2ac3a2fd91ddca71be51a4b7645
zbfee91891a23b52978744f73bcaccd41e1508f000d68b34e92a21466172cd14bc478e30ec3eb17
zd365eceaa42ec6e82836867f9104b605d0c4c4e3ffdc0e524af0961becb8edb3a3a7379f6da52c
zf6b6c7a8b80bdff401ecbffe776425995450d502b7016473d187ed8c42538f918c3f6c692b9092
z90c16e701c220403e4302e3089a17608e3df68f3077f7e6e402c4f5aa62bf4d3e21c1a9df18c63
z88db700eb8bc06e83a158cafc583fe97d79eb3f39023f6cecbbfe5fc78598f3e361ca40640796b
z3cc356e75c62b1675bfaa8c20769046f9d14953a257794fcd2fbde639e64f5271a3155a18045c3
z52d91427dcb8aa0def79af7f33c0435e45ade07d624bbebf990038583ed7073d1247a8b7f2b14d
z245f82637943f691af3b101439ee5da4b9e6fbd411feb464c2aa7d86cd6d9c1c6f80ae8a212530
z1594a679129bedf5dcfa99be2c96f0283543fa156471fc65195ed5dc8d1cd2c60dc1a1141a2f79
zb20d4aac949696506e4d15f4b821f5f8a3f43ead904dc2308b4beab17e1192514f62e6f473abf7
zb564c1872d037b0cfa6f491d97bd70b20a2c52c06d20dca391308e30ee6cb11434ac6f1606d6bf
z38786327610c3ce228a15490b4dbdc61aad43335cba158c9a68564e476e357c6c901094b8e27fe
z0f759c7315bb3630683c72a7a19e6f445e00f70d3fd92f955e98b38cc7b5ac0aa5efef76a15962
z3cd11ab4ec66602554021848fb489eaec862b69ffce7f7e8e3c3297aeedc1e052716128d2862d4
zf7d26c58928392e7cdce1614f32ae22c01100230f647145e73397acc2c3d1db85864d81834eafd
zba1eb2bdab2019618936911e0893909086ec22b767ecb9181639bf4d54f539e5800d4e62f482f9
zd55b5aef4222871243208370d885d6924aa4eac90c27b506493da9d87308a619f71f519cfe9455
zc7c680eca63ac6fed6633ad9a876c140ccd57baea0136741bf55594b9fcea9b09f54b1e96f736b
z0dc3872dfb395007f1305ea895d547c99d220c892edc66481d7ba49e88d904cfcf4491f75b574f
za721beac2c23b0f7ede2f46361af758a13af70e05f66c201837657fc3965af6737e4204bff2852
z5df2cbd654091b187b416346cea4f11867b8444b7c017f5fba358e24bd96c73c0cfa6d444e516a
z6894eba1ac0bb456897735f58d48fde59472ff318aecb8d0874edc5b39d9e1f033fafe8ce56d21
z4f41693e62e72f4bc9036dfd0b45300787d4abf4913421b255b9810d8d06a4dbd672a9140d0043
z915c75e80db1166cfd90805c05bda599105404710da132e93ca11230b43ca8c2a4d1c1051368a1
zb6d4842da2e49f5393fbf732105f92553274acd090be27cce2739b75a1192031ddbd9eab4ca5ab
z5a85d4a4f09f48cac89c52340f879d96bc7509e33b4764b1faddc8e2fdad1e9a259c5abac06ac9
zd9533c774378380f5d34f2a16f0fcf98ebda1aeaf7910786c2a1981274918d700ee9d4cab99dd3
zd01e79839c2607a4aea6cbedd781c8a16d1dd8b052ad0b5831aedc029fb18fe6022929ea3c4d4f
zc4f2e279a4c13e49584385c669966a21b25cc9f0f306649e477b8b5d911b7d57bf36b159e28e0e
z7de8b014846e4010ef7ab350c1c5746d751d75dab11bd986528c35400b8d037988013b166951a5
zf9d67f570ec4170091380e36dceb2ecbc11818464eac8a9f6bc5093921135099bee1e1d406df07
zf43327725d51ee5183cd96bba3354cb439346b9feac32e2b8bc4ddb7045c71dd1ab7cf05be52cd
z493157d69e06bd37e601ee73a0432ed7c78446b582b7c37a21db9bb328cefb18b26e66d683c324
z088b4361cda4f0947e417ae3690decfae7d1a45fa98e674bacc111f19314de3119ac29568de358
z94c18dbb4a7cebf729396660f80327509146891263dfcb15e7468f8cbc6e3714feb020d1fc3442
ze315ca8e94685650c19920d47ceb74c24224776e522363895892b6c896955ca48156139213189e
zc70cc26794f750c6e18d03a9c292a0c8439ae19ca2849598576afb25bfd079fb6876bcd3ce09d0
zfa01c5e5934815b49b78602fd4677ed08b8c36cbe76bae3b093d1e2c12a239ea859f6d9b752e3d
zcfca224073cf5f23630216e35a8fe0a061261a97adba79a3f70f454cd76d0501e020abcfe2f2b1
z58b7a692bc0904c776707b9e649a923211763a5dc9324ae3ee387e6dd5dfc155f9f730bc870111
z56622c2c4e6274a05cf5a473774983b88c4b638681a1b643787b3ea87a1ae64013dcbd849247f9
zbcfb4467bca314cec81d498b9f61f5aec9d33ec7bb72c5ecca93816a251ba26d694f039413dabd
zb9b9d897216879896640a46928540a91381f0e22906ec2a90cd7678f60084b924d3ecf3797b981
zb06c4e14e6448f197ced6e5f2a1e6e498d8adf457e433d1f5d1a8d02b7721e723d165cfb61a4dc
zd0226b72a3dc3d584c30acbc5d8327923c7216d5dd928d79aa319e597f79eb750c0cb52b315ad0
zad4ae8f8b40b154bdba20152299c2c1bc01603e34953c70674c10f163a4001ef7d8599f4052bde
z5927e48b7cd55443a76af3a6802b6a975a697ceeeee72b674f04f86a59bd981a698e80ff4fcaf1
z175c1fa0635c8d81ae7a67a20fd39aea9e400c7754bebe553e77c7cd32f5eb5457a44e6533b935
z79798c256810ca6f2606d4239a0550a5462581738ef60fbf461cf873e052289652f468ceca0166
z74422342f78ecad78f3c9668b05666dff02b631b6b1c737eee3babeb25db5795a003e01d164aec
z3cef34c9666c015eba769be029ac5ed5ebb11ae10d8b73efefcabf36a723e01cb458c30ea84cc6
z9109755dbbec208a126458461102783811a3b3537bd9e07579d082e8eec584480bbd313bffff33
zcc0a3acf047b39295f891c7d8664c0be88cc08fa47211e3409cb28f4552eb8aae4d09e13b94926
zb317963301351047cd64116ea346f5b1ae9b031e672c66f84d98b60e8affef3fe698fece3f7df4
z36f81c79150b0fe6f1533223a4fc0d181db41e5bb077f5a37b9a70123e83459758d4a5d9038301
zfdef2f822e35fa5bad0d6f5d7dca4906d3c28636ca1b10e89d88a1bbb387a8e30bd27da02c030b
zb8fc2c3003261aaa73e6760223e00fd8d6422b4e22e36bad7fdb62e00e1e26f3450bdf5b3fd18f
z6c7edfb4c58e69ad15759fd26230315f5ab1459665e522912dae1efb5985a67440166f5d55d700
z214bfe85f709012158af17ee45678b3c68629f91b7964b1acb382d3d090a3ee40bd80d965b05e0
z3bc8d77fd859ec6be6dd01ba233ac4b26e8830d768361acec5660e92cf4b87bd7e3356835dce89
zfd73e8c12af045976082b23eeac506ca1a1c5669616b95704f88bd50936bab51ff9ffe15600fe9
zbd298e3bbb16bcb44e118115aaf5a24cd5827ee786a672fc322a1a3d4c1a755bb49c189e2b71a2
zcc85ec1793c2f76733c073ab7c9434ee55581e6059c594e21461fdb3bfc733fb9b7515a66a0d94
z6a037687392ff756d3783f61704fae5c5586676c047b9df7d822410e8f1247f2c07ce996fa2123
zd9d190555bbc1109308877c6e4b98fd34db645a4e8d032c01bf94194477d5ec9158d6d1e2833a7
zaef6f952c209883e02f97b9c3da96db181bef73c454a5f6233c6083cdcec1ad84ae1ec56a853e5
z23cf9f1b3d8e16a939025d567a0099d973b57ce3584a8e18cd06d7099ada29ec76cc9ef09a2856
z02f8334f060055be2fefb238e1d4058cb686a4da083c3f62d330f75bad7ca23ae4c1c040b93d76
z4fd3d716befeb8b13685f0181a7fe0175bf314b209d0e9b51701c3d3c07449529ee8248742e7bd
z0c14671788a50eac36f5c1fc318cc3ccc94f834410231ed4a47bd9f3021968f8327cfed7542372
ze7a8565e86a4b6662bcbf2e4422473eb6613113b703bfec1220ed7aa759f4d0f25369ab939c687
z820ad1754f69c46ec692edc0581efb2e1fcbfa0a5e7adad1882fd504dfb3933a8e2ec50e82365f
z3056a53cef4edde9b82fd7cc28b3c5db9963ac777c6bc2e32b85db2663729f9210b3af75bd7941
zb8819c0293fb5a7f6c9cb7df8a6663aa943fea4b149fb230740d1322efb036414c5fd724d6005d
zc39958f76b359abe43daaf2d5649b0ed66eaa5102c5777700e14eeaebc854c8535e1c0981126ec
zd2fad7b3424a5471a96f89c7fe399bd806aae49109f06709bf3f6e3497816feb1bc608645c7af7
za7a69f8abfb4536b616f6a11b4336b811cf641d8efa8b13425484eef9b6329d36d6ccb978c94e4
zca976195a1ca67d211821f82f91d870e2191517eb14f4e1f7445dcd4b729dd60c1e3df7814a956
z0d047b2541b42b2889ac56933d542daafa88da55e622e66fc1d434c0435da6c17734e9d8e39023
z70fc62f2b968698b36d0f71a119167f2916625c03dcff32398f12108356d9d231753ff7b1e0dcd
zfe5a88e2651f179611b378a5ed31b1b68143564282e51084748893881832d675a77b8f5bd9028b
z08c07e00c60252204cf1a8fd0d3a0c772b870325f3d1678a1a636e194e47d57b2417ccb91f5235
z2b7668821da6ebd96b14d825da4e4dfeb0a09fcfa7f36ce24b7eb4f3615945f52efdb1561efa62
z1203062158936ab6e61cfcabef5996ba0322cf90236ec5ce3b66aafa908e530a4b05cf78baa54a
z1984a462a1f156035c9438893588c4f22458fee61440bb81b2c6a589faab85fd35f14f21284679
zba4e4c1928fad53875af33e1e2164be33b00a6f0aa33695b971f267f0004d77d47a4e1adeac39c
zfad904710998572379383353660772606b24d9bd16f8c202d074234b147ef09bebcae7db87422e
zc496b7f178e24b474250d76b993d5cc189d5227ad9a5352f63b9c8eba2aa227e66fdf836a1f9e5
z2b997e386e1ff6be2f41b9b605230b4239e59d598b9c3e39cb6152588f6ac19709674b4c36d30d
z24d9e99d3d39446259a80f02fc802eae65c745a6a4dab06ae203ec18e5560805bcea519fd10979
z3ca6622eb2ffbf74016d057d5105234bd640e2d6b8b9f10cf4daf831278b57c3bea16f77d1ed5d
z849c4f90d73d7450dcc429b347bd72813994e73a8b28ebf0fb871a5fd62f6cb4770e28212727d4
z6d635fbde679cbaa7982b1cb779f54af683b20428f0dc503dd5783cff196aa64f2f6db7c343e44
z70ca5c51dfa4ab42e77c9c109456a07497ab53e550d1a83e5bdbe181784bd43935ebd6bbdd7714
z60c65538b17a672b2f4b57e7d4209c26701b421a877afb147c64914a76b8f10ac387675c5db616
z09b6a18467d3332c988a2daee3628b4768654b6eb4420acdc2b2e0d4ed16d041069e5780975271
zc36415e77cd56800a34af7fd130cf280c36137bb96723514e16c015aa77dec98809d4837fbc493
z8a20afb36f37262b662a57498d773435efc240b2e44858f1f721cbcda45b65f5e87c503d9287f1
z6e29246fbd95608b30717bf0f6b40de166efb77778e6d3ba6ff75c1f57aae90aaa8fab1d96451f
zace03343275db68f340898bc204f43477a44267ed1920015845d19348d78e58fdcddbfc12ca840
z43a649bcad9802d312345099ed5b867a982897e98614398a2b96d76e278f852bdb62b8d0d8b386
ze6ada701e966497f1635aae1922737f6529fe25c6e4b03a6a5fa112a8d046e58da49b72e5264c1
z1b0595e9b8b4eb73fd3fce631879c319fd9f5a6f217b6d48111edd14899979870ca7ea29530da8
z8784baa9387cd20e5cf91817c52a0bfcb52ef50df0fbf4d36fba1d58998d3bdf1b1b3f1f2d8266
zbb73ebaa1293eef6ee4643ca043762c379a716acf327f64a7fe120d4e596c316c736aaf8ae46f5
za50db4dc88e0392d67cb7b9a733c27a1fd58810b4fe275ec8160233785ecb4eeca181d112d2b91
z7afec1c54205baa816e62ed1761998d4b8ee8fd4bc441cf7f6caa35f533814079924d7ed05dd38
z06790064dd8528ca6ec641d22a2973a8930389ae45e03ed7b2e58f83a0f7f76259141efa31e473
zd5b491184944dc70ebd8b1865c8c932f0c3a4b385251d37ef68d09e0bb6198461092fd9d32db1e
z3fe2a90ca38c1f59450b706b27d57aeeaa97dd8a4603ffbc62004362355a97822cc5d87b0de55b
zb483a38eafe3f0785d7264720f35ec390f556377609d0b3d94343cfa96df12e2f4c33ea02c5ebd
ze830c9c598963e2c1a6adbaa5bdf8f9d02b95a7c7123fa12b791cf933d3528a81d7146c0f8c2da
z68889af9d108b98d1872b07e8d61526cfd02316ae9aba64760cff5f9365962ac2b5c4b4cef903d
zef210d9cae3b0ab9be0328d8de5f4ebe3484bfa8bfd89add8a3f050bc0810ae27ab5484d7e2359
zc1006c2f9cc861202dbfbee32eddd6ffeed56ed98ad134fccccd67bed9c70340d70d4a8eb73c24
zed5d04301d562d2189525dd462553150afb3afe6d702fd4cd977b852277643b2962dcc228c9b55
z17120b810bde90743c5e9dd8bee77a5fe5dd6f06b276ba77435c9723422cc6cfe9831c808a80c9
z1518111ae745568573620b566edfa14b90dbbdd05d14cd8491a3d8fe54b89b9d33630687a656e6
z069e057538303349d35a3311cc1040c2e57b9efd67edbbca3d44d7de122b7de64d605338f101c2
zec183d154859b3e5ef52ac42fc01cfd04eeeabc95186c2801684cc7c80db11042dd288fcd863a0
zb55c6a80a3d426c4a94a7aae156941fc5ed1950a36288c8db4eb381d109313597c1646e9bff013
z7316deda907e4d303f151ec11dc83f1cf4b2ba39b390802fd75644d84c5641205df54fe1b2c70c
zbe3fe4d15d65804344e9b2eddd5f30a6aa5e699bc475d39bf8f4f65a2500f6b38e0a32226eb364
z58287210f513cb1e6b3a838110f03d7753ef42cff99919a2aa2d3001ea58825161f0ad311ba253
z8c72a5df40ae88b671ff700d22313f145e9d044103216d1750fc9dcae6c041f7607adc5ad40210
zc567845bc99b6c6518312536f91a2b304b37f91de846d3f9051fe038a12f55b2d41e5bfee26aae
z39d1398a5676caa1c7132330ca8c62179a96e8c93dc7a3fec04c01a7976740b68096054d36c2fc
zd385b6fe9bea9829900e1980445b762e5d9609ddbbada7c72a622369e8fc16225ffa97e793c84b
z27ead4872e9af9b5553ee24a40bb4b18e57449f9a32bd714aa73b632cc06ec8864b4a4dfebf887
z288c3ff60931febe399498cb2345572697caa80042235f13ec4d2b2692488651d4f6cc1f54e30b
z8c8104ec21b4cb808c5648b5f471c1763a7b821367d9095289f8495ccb2a05016c12eb8abe85f8
z7262f2aa39646ddf38eca1ab10471b88ceaf1271745e29c20741ac2cc4164c2431e9ab2695b487
z95a9f48733a28a88cd17588037ee56024d084f35849e4bef7d7a643060fff0dcc945d27f8dc416
z392544823b5f2a83acaad3fe7633aebb959d8a7d018507e461d4eb63622a8c4cdec7d181e9a829
z6402bc9867b79b641528f74daca7f719958fe563461558933c3ea31100d6671527d5bdd8c324c0
zf70744f647af2088c51ecd6f70e5057e35b180920aaa76dc00129e541e23ff3cab5e478c286bf6
z02b4bd1f7cec3ae192dd5002b0fa5744f8cb31e77d07876a881f36db50e7a9e2c5b4fcff1c0f05
z5bc0977c654ba48d40cb889c5a3d92e44415e5a6b456826aff278c63e1e05b0be5648187a9a2be
zf2be449520d2fa7663c4dc1d71410f9fea2df60d23ccafa2f532bba3d64ec78e5797e6b4d66c7c
zecdb8af4fd8bfcb9dba6fc1f4400f770b251189ed8f6b95617de4202226df0d93504d6fa101c64
zc9f67936daf182fbebb344e955cc95d23d8ab54446ac02861fd0dd929ca74f0b5af72a4a16d464
zb84d3edfd5a95e2c047e6d2bab4bee408f05aff02c2ecb3bf3b2b2e1cce2bd3a57f77fc8b849d9
zacf679def8144637c25e3f1a4fc71826b6a9f15e9ba1d6350caa0db1bab01a9b6eedb7dc632cc0
z732ab4df8739a73a81a233182a30c6db38421b5bb6f1bfec27bf42046eb7882f608d9d0e558e9a
z81f9b411b222a6b782af2329cfe7973b1b7f96f37b2006a89eda1207a8aaaa117e0dd0506c9565
za353981828b1ec4067381e31a8d0f5e442ecef996e10c37adff77648d25487b90bc4bcc752363d
z5f1657192aa125f4a9b2d9761928d96806dec3bc8fe5557cf00b848a708d17deec79d5fe62a631
z92f48807138d89669be6b86fc27f6038f786d738bba8b1c30fe609e606002e164dfe000e124f5b
z75bc41c27728c931c5526ad2c204e6ba3680d06b16af7a2b9c4918edd4600c01b659ede43af5bd
ze70dfd8b07e033c6dfd8c20c3f8dabe1aa724bcab303b0cd22bd1299a7c7f8e980a3435afc3d38
z0e3eb474b88f2e4418d37c0b14754aef29c0d4b5f67ab8de86db5fe2340cc1468b8b9062457cf7
z2945a76eb091243698e14b515f1794fde8db3d67a82ed1d0659f8e205d23147d2851b83afd16ad
z2497eb8e31e1d47c6286713ae1468f5ce4eae34b1490dc20ccf3959a66e439b3a77d068dcde037
zf274c549ddd0678dd1ef0f5a7de853eb6edcb29ee65b94137667edf9e27e873134dcca0ad2bbd1
z362574f24b98329f3c3d9ffd41996b87d7569f32cbea0cd2217f4ed68c7af00bf8c2802fc16fc3
z35fe5e016808750975c87c46e6425b43a4bd50f6771fc9bef950cbdc259f9f960f969c75db9958
ze6de2207207938486a0e025b809a6e55fadc1e1839a7e22f8aa3bbdc36b4759fcd47083b62c564
z1c747fa264e3758208a6e504e9791b1d386fef098d6c03bbd6cb35c5d9d2bdc6748d07742ac061
z5e5389856832adee914237ca17c33e9ebfc169ec6269020555c686552482e939a4635595a13685
z2347823f362e245d29183491a9396e4d29c74bd7647b9d46a563ab2fa5aa8db7a6a184372ce576
z627cf4e93b3a9669d8311f6fa3e3715335f3e37a1e9bd2f1f2fb44fbb3ae4d6fe24a31f87d7eae
zbecfccfe5f0030ffb205ce39e423965692c964509bb98eb514ec4973d938dd724e21a000a5dff6
z3b413376fa4a08b20c3d292b26bcab11af78653427fbb3fc0851ca99d6d2e47f2ec920d4ecd50e
z0ebe3ba7549112793fc1cf19e6949168fe5d52d517c932aa3fb97ea298f1a7460ed26874c5e00c
z478812c4ac3d7dcbb334b5630f0215adfdf1d8c80a936f9358da06bfd25c1952948ca873f006f7
z3372ecefb078c0fa8e47cfd9b11fd2d555b30d3ab947ad91b13c5b9152cd161036ed6d7d5d4512
z8ebde5533b13483a7a5d427cc0bbfb5db508b53fa206d8a34a6451cf056c7fc3620a3a6f826788
z0dbbf831b948bf61f0bf09ce11d01e153738f7358e882bedfeeb628316341f001ab6023a178b23
zee290d1c234cb645557a14630f524c3ae4c24822b8f9f4b00aeddb8afad40b383e95eeddabd476
z2ecb2cd5ddef38d1f54464cb3b245603515d20227be49219757ee4fe14175181d6954fe3fce9b5
z6394976a2303513e6d37533237099e1abc4a5a161bcf3c73fb413172b538b7856df7e41c4d7e59
z8cae8c5a030be2cfa0ba62dd60dd1a5238e239b00f839d4785014bbdc67e77bce4ee8e13b3caf1
z773d5f1fbf8975f93d0a351c752bcd4fbf8c2164bb5feef4f57bb88a1f403f21716a99624224ea
z23618ec964372cec7f21ea9ecd39dafb2507d4309b52f5cc6d7aab506057f2dd5ca605c58104c5
zcf6f37a201d12d368fe6050c1c04977b8712bcd36caf6eea554890a0ecaab525b8b13dc70f132e
z0fa943ae8aa1d9f742f189529f68f0aba58cf042ba8775ef383d5414b1a812eb29a6463d2aadbd
z9704de57f9faef0f367be506ea1f4c62501ea40d492a8ec29d3a2d2530dc250de9279e2f773d7b
zc9c98717030ef8b8a5905c345136d9ee32ad7303f928bea11b7b43a2bd82ed9a602327122fe797
zf857c42b845be32402e2493ba81fdd3f46492f5cda17afdbad62a80aff13d0aa4ce0661cf61163
ze8a49f3a829fb75b62d06438134d1802a5ffd0547748abfc63970f54f0f0bfb4dac8a54401c592
ze8934dc3cd2f01793c4ef66d0d97444015a4a5466fe398185998e6360ed7ffcf3e3b60540114be
z72b18d47043ccaa8a37f75c1c2c70a8818187a036080fff14228fef563cdadd80ec706eaf28ab6
zc70f7c810f118f1565c30bee6649fb8a8747bb35b8627e4f192f55bbbe18875cd769377b778ebd
z9b7c998224cc1f98a3a4880c48399f31a60db8b8b9d6fedab3586374a907bea93cf76cfe4ed979
z026f9d8aa1ad5577d2b38401e08c5fd64a7a00a3aefd6d811dfda59aff5753b1f1159d17d6e7a8
z68d2f50cb18726d4545f08a7ae6755d41d08d080a12806a6f4766e54e9e95c5eee9d8fdf08b12f
zbc239f31132f1d39c991ee972b69f8d7529afbf9f209e6550d875cb50c15784e28c3f90f6aa8f4
zb97a804bcdb83d7edcfcd4126f4b7b90639478de03e4fff3bf982310d20db8d2a26c9a9920951b
z42fe62464b02dc05eed37c12b84fca04cd1bf4c224e0554553525f42cc7ec3b3763d4a9c5caeb0
zb6b5c3877c80e13297035e5592f5bfa3e7448b4a81ef6029542cb7d4586863fc173de8d47c7f98
z502ce6be4aef9c31df9593e08ab83e44d2db13b5136b27c38c417a86a1055cc70c7203ac00b051
z6a763662c9dfa49d89ed18db68b71e5222614a3d647c1f8af7302991cd0bb917c058afb3fb3b04
z2c89743eba38e13bfd6bcab3bb62e4f87170052bb7c7817f3506985aa45477c2f648b195c22286
zb0cad865ed56510c44c616508aa10025e42147de9675b183daeb4e4b3771560a23ecfba2edc768
z42041b7a31c506760695230f1d828bea4e5e9cab7d4d69e2362aeb85c1da9b6c581db1d0559afd
z1b54f3f77e454438f0f9713e56003eb2cd3c5c57e8aa99ee8ac4a33e830c6d617c41857db8da5d
z5a1f245a131b5f0be7c2f4cb67ea6f22a4a91f241d05219e37b62385239999f92251705c887750
zc4abe176b7a85bde3f0d488d0862c97cc04104bff99b2912d3d2f2cccfa18795ef66850c9016c4
z46d0f761142817654b26a29a2bfd8415581e3dec4dc886ac90aca5957c726892d885ad2923425b
zd5afa1d36e4e62a62df8f4a6ed109262397ac99d59f76bb3c52573aaccde5d19137eb5631290d9
z7fc9062ff135ffa805754d6de170065ed9e50db80d0ac0bc7233849bf06ac75c273a2fc8c410b0
z14818ff829e4e5a8935e540df624c004e8ac9cd9148b780e07de0d6662a3fedd4041b668f764f5
z683a59d74a26773bc94785de72da8fc236e14a25cdcab0161748a9a1f6845c7714b8d3ffcb02e0
zfee6920ede163aec5e6edee115b0cb8aab196bdc8002c400ddd83b3947fd42d7440e7ef72c20ef
z1007f826c5b3e41e0888cccbdd5596cfa7c9f1c4977cea84ab913d6adf310a3ececd02a3eff816
z33a6ff701fe08a6e2cb690d967d9138a573f76ff67e399af3dcee60a64a24be2f8752ffb67a248
zad2da56ed1f376d44749a75f52820834f4eff9695b1a98b83d3440ba5b7154b7f9a5bca616521d
z176b736d161bc612b4f1703c705ff1b268ed3e4aed79f722f1f95dd38094685745e9a4f69767ad
ze1bfcaee3c7ae16fde2f9891976579f069aa59fdeb682eedd8cfeee2568a943b59a05e29525713
za2deb396b2b90d95bb44ba85f6916410102217991d4352f23a52925a6c1a2b70599a7ccee41017
zf33f670d7096181a7133b1dbacd73899da9e64c7f1f3f1107994537a5b24d48b290928a508b0ad
z273e583f72e01c86a38137c64e38db9555a5db1178c96f75a91d7ffae8eed3730a1c192d18202b
z11fcc7a78e57e9dcf9603409664bb2023d792fd68eda5ec3a098707e7924b9d03502bf8bca5be6
z50e9c27a6f4df6ad6776dd7a33ee368b607cf09a2c9d953a71ade00c8b6f9e65e239547cf247f4
z3145919c6d60855b1a15ab186b6d09556a31c8af9aec5cce4686746ba1c044206251d070cea1d7
z487a55089726b8bd0d1e7c5aaf9568b9e0960c8df8ceddb3b1aa1f92f2691901b09ec06282b2e4
zc9c1cd335892ea3ab2c5ab2b99881f1b739eaa375c2564ba949ceefab145984f0afa2fc9110816
zb0ae92461a4b7fa5de89f49697773350cdcd0b8799b463a209850b0d54fe63065ebba56fb9eb61
zaaf825cd176d800bb5c8de0c8898916f3208b30a6122354347d673bec449e5090e7a69d3a67250
z2aa1e72b823cc3eea9dd3408cd02e231ad9067d9944d99a6605993406fafb1432bb662a17e215c
z8cf3dfc270225761d271fcbaadd2845456026296567fd8ccd72882f387b8571abe7c94e2a5fa6d
z7dbf0836589bbc4cf9b7125cfdc8b9643257831f7c01327a2a1de1a25e1938a646002bbf73f3a0
zcc27accc6c8da937c089c07d6dc52011afbcbdae975b567044edf8fa9cf35fe267c745c82dbb8a
z0bda433f03c0e2e4a977cf1f23c143aa1241a865fe0b71b7edcbc10bd7a7f64b5567c029684f8b
zc9dc3fbe74c6731ba83fa135ad6460e70a25be2ee25f256163e59085abaf45d5040dd4d51f6bee
zc81e1477d56133c61101e61fce81c55eb871297d9e32b0a4dcbd0ed9388175a67355f5db346ac0
z874fa597c23b31d5453d77b5db74d2964db053b62ab9bf058081b280022093eaed7f68c21492b7
z29d3aa88c0fecc52574c5e2c621905f450ffd27471253204888cd0668105e6522168c90fb88342
z5040c4f7158fe4e07b3e89eacd80d7229fcc832f6599a8793dceff896d4c0925817786992ffca0
zccf06c53f9297d94e83a32edea0c4f989f416cb411032aeb6a7df882f9b3e3e29b0574cf3303e7
z1cddf80f6b8dca5569763464926b9c8b1fe9077ed114006564244072627d5443800c367956a319
z1cd30d03bb5deb2d50d8aaeea65409b62f3ce9bb21fda1f667061a40a8c9041b3ecb9e925a3f26
z31f59852e5582962f92b31c03148a5f5e74bf9a500c40e8ee469c4384bc06f5aafb4704b82bda6
zf6ae1e928ded1736b47a2a0af1ee91dcee3fa9a7da8e4fdb7509f49de417b119fb4e20a6531920
z38854bb6e2b8ae657f408aa1da560cb10a7ca63657ffc144743a5d2b4f107fde93e45fa566cd26
z1cc1f89f50294c4c9c5b05ef05aabcdf14f45f3b6a24dad7cf17a434edb98d51d931deb701d4db
z9b088a235713d95d4031735525a56dbf19dda503d4adcbd8919657b95c2e7d9b335f8309f856c0
zb95ddc41e98b5a706740df38622b6709a4b7a0e60ffcceee2989c061832a023a20a1402ab23d5b
zde11cd33ac1dbb4c6932a0fe8cce0edaa407ce66f5154209d7b383b6ce8bb135d5e0038657bb8d
z08930c5207dad8afc49ff0977b15f49838b0c24ec77e31c43b301670579ade0a5a1469fd027a7d
zceaf2f2563b0b4c950e8c963ccee6928b0927475f9c568f911ac7b9aa51de5f7ee706dd887b26f
zd1980a1467ec3bcaa0e61fdf6754a96ed438326b14fa9a75532437c513e35749c7a44b84842e98
z9f929999cfc0d0f075c26b36543dec7ccb78a1c3e393dcd53d0f1c113d08f5e969784f879539c8
z980358a68068df3b99d2952500e32d35cb7cfc3f97f9d9402743f5039a7fe39141765140a900bb
z124339e7a50b20cf1828a871b23835d9b433c87693b7f94ec4435f0d442003daae26cb65225a34
z6e6ceba827b04a979c3cb28ef08453b45b5bcf0ddcdb584d3ea28a34dfbb7c0b7ba37e29cccb3e
z3d57b2708e3bb2009fddedb5fd12e2cc2bf639cf60da8220a247f4d27e0f845b9bb9c18731be22
ze1290e62f2cc650dde43a9c3870fa82d314d085f6790a70aceef83af1c1b3701a1f954f0fec5e0
zde35ef49460cbbf10c77e2bc6ba4a4bd4258b33fd04899357b3fdcde883dbf20619a439768538d
z98758ec626bfb4a6659a8a515e0b569e5523e248892bbf87d82874a57691b27df236feba53e9d1
zd5bddcc5c99ccee594f9c1b5ecc45aeef896eb6a3a25655e1a88bba4aa44b97fbaa898ae1e6b07
z629bf4cdd0b07056de7fc9f3395dffa4f0257312c2ece2dfd434e6dd0537c31ee6cb07bc63419e
z660735cc26a75219227bb88e42659c03fce90ba51ca2ac6cde17ed943d89f437d1d1684416c7cd
zb3dc373b40240f1ecf4733a39345bda25faca0c562c1a372b0b1ee79a6ff9dd2f32f227f668036
z7aef776a877c225f0d0c568ba89f69d07b1dbbe75b068e7f0350ec08d43ee25dead5fa6fed7587
z9123a52948b19ef95c5af08aa96f5a35d2ac2e5a81038454500d82dd2848ddbbfd46ae91239ce9
z08cce3e5b241b18c9c672a86c3d373c4fc2a7f277799d0217cbe5e0ba906aac5a0380a17b67904
zdc87db4e8865d74903850db042a349de5f33c22fbce73d10396a390da56941dcc31d7e56b26015
z73547fdf673e5679a56f59b4350aeb11a2ebfa6688d7d37d5ffea5c16b5d8a5411cc4fecca4421
z754a43bea6a9a5770405f55f17e837ce9b2acf4e12dd9d74306d254d9b2d946308988a877bbd83
ze14f238dd5ca13e67ac437ab52742b903f0048eec9e767eacef7a1f77f7dab88758f1087d3b839
z095e2460dd4df376d803da89c5d33e9f1c90b39b29b05ad9d2740a3515aec721f985e475431a22
zffb4d52b1cd3e71014f3bc783887566338632aaf10f397992884789a7456634e701ea9ebf4807e
z7dbe6b68772ad8e936978d555341652832f2584d475cef886d925a856815991203662b04cddbc9
z92c61bafe3fafe2cb4ca2aab8c34f57c0fbb21c457c1e0966459440ad5a2f34fb9475972e4239d
zd6dd7078e07bb55bdc8cdb22007b062bc4d820dc1d3c28ede39586e534c6df316f51a1f27e2824
za0d1678e3929b7ea3d988637da913bb7852809dd0fd9f9a31a30e32d4bb6795228c673587d50d0
z52e0d29ae84337d08a0712e1859675ddfcbf0d7a1b3aeb7b98c0ca5caa4eebe41db503f953ae67
zac28fd2d89a3fd91b495c37f3f1da7ae6cbb57b9c4507b73c28634cad23683fbac8c5b65b6b3b8
z6dccbfbb438b37d543d85f4c8d4b7010871d4e36c8e8fd522af6519e4ab5d845fccec6570c90a7
z9d0960929b1f95cac693aa9be78993501db651cba3f39bf20b935689310921fed15530f11e8017
zbfab781e10abe53c65d955804a3d4979aa907fc73d3fef7e2beb45f49845228cc864e348134fb2
z96c092c416b7b5db598aad77421c7ce1b0fcc06baa9e104de881e57845cb33c96a297365766277
z13ad2ba3ac1fac68d8640cc7c274804c32605e268269d6ecfe4a59e80d3e290b829707441eba90
zca6ff115d8cb9151541e94868c1e68436682c1c096e56ffafa66e013c9ee5c3e53a410ed3d0ad6
z46165260fa0f1698d4067e68cbd0d04abb115f03e97ce54d340e44ec919f68eefbde284bf3edef
z213ecfd513f64276f981c85c10a0b73b3e2564459839ded65bdea9534ec7cecb34b0c34b4c35a9
zf035dc3ef35f86455a264112c461344d936f967ccac57616a40fd2e778992ca15615aa9b9f33f4
z4a44430f88e1661c02c53e418cd8227619e92af064f3d4ee4da73b8651778103b4170349e50416
z0a5a0f57cd9813a542e69920269de725cd7552c387addb170416abda46f4e61ff2768199e61ff9
zc4b874db8c809d9965f443f5b72be434dcd9d43aeba7d834aee294f78c0c4c9d92073448641ffb
zee88012452230bdbede80cfc73c6d2154fa1525f5e58028ae026eadcf86e5fe8660b7396a376b4
z60ad839b8dd83d784a0d7ed4f3a0607ec8f0fb0a9b5e21e54349767239edb5ae6342966ad30314
zfd5fba966c15df39f25021c05ad6b6b6667805b928e74e292633c5f2f6b7a0099212e3b38859a1
z2f50aa685acf81ecfd81172199422f24a9c61b50f73b4f8df3c98a5a4001b7c92e88a0b34da782
z07834614f7878c1715b67041b966a1e6aee38cc7ad6b7f68975b0eb3df11e4d0a25fe97edd196c
z15dfe20764ca8b24446b49d68ed499e7c2fcf8b8c03a2535c9b9e141f862b1709be9631e9220be
z78c3bd4a409d64a9b800894d1d63938d8e535df808a72c8c9b1a04cbcfaaafca1de11388f4274b
za37fc94f4a20e2345a786c9c15d832bfc1797facdafeaed0270d5372fb74986dbb1457da6a37c5
zf108813b89d32a4e758774d340b6f121f8c82141adeb4e3db97c7b34326d166f03379821f02e9e
z1428d7a1ebed2f6c6ba35bfd1d5682a7b42d4c2e1528484f17b9cc2b0a57eb1512465012aaa9ab
z7a47809dbf9d856a509e84edddf6952725f4ff9790bff86a9bce058538a8626ad9a3b7b5c922a0
z641fbeea562ddfa1bc4dcafc3c229df8b09c9c3134f2d1340c96d1be7a9d48b9fecf9c4c334bf8
z5d79a90f24a6a274c3a9886b2f4f37d259954aa29a92b68d1e43fb7301501d40e5b16018cbbe68
zcbdab5e3ac23638889faace3106133f41e274aee0bfcbd423955b9e4b5e5271349d8d0e0b91ca2
z3d3c8f41893db544af0c58173562010189df0482bd1dcf775323ce199fff78efbda64c8128050b
z1115e95405763488ddfcf39dcc01a2ae647388a9ca61b06eeb4647d78c18ab69cdfe46bd1acb8a
z6af72244c9428b2418011e259dd6385e3e39c8659e908403965525f856104f01c8e17f64004fed
zd45a452a60a0634ed86e83f71c994e21a1bc85b10aa1e642f7eed1f5724ee17a517afeac64735e
z2e148d3c81df44d9a512bc2d91e157907b41d0a8c79baa8fd25aa6bcfe6dc55402cfd89b7064ce
z6ef8a88d1ce48bd6acfe102ffc377dcf5ca7ae9fc85c50eda7359e113beb98d572acad80062593
z0bcbd921aa9a2f6aa36a2d3dbaca2a21fce4a01c0600154cc17720182c811025f5813c717f8ef2
z57b9bd69e9efa0657dd52b8f1c006b920882f05039073e55dd0cd587230a0241abb2c6ca6afdfb
zcee09f41945a49cea60967216bb5bc744a083658c8b0f07ea144c6813ab3f53436753c9d299abf
ze1f0514eb9aea4b24c690ea5ac7f8c090f49d59ea3455ee8e3f8a51ad427790e1af41b6f3c06b3
z41308a16611d021439fd6b889a539b652a2a0f0d2c38b6653f94e9fc0765e7e30a71aaf3c72c4d
ze76c3ca41437922530945bc817c8fbe031419066fb80b29e914484f980e0cbfe5f9bf009f4e9a5
z09c8409d1309cc7112f9b8e0bb38b7e5eaacad9c7f9e2a5834d04d72f2711b8f8ad1910bc4e754
z095249805f7c13eb41e77a211d89aaedb0806a8f3b26e68ba03141602290e90b8002496f1cdfb6
z1363ab5d6d10c3903397cb438d441812cd59ff87afdf8403544574a6c1f0dd3c1d364ba749312e
z1a15fa54ba1db61b9be01e9b4d4209e4688aa683b726cadc6a15b48da37129d9851b758835ba4c
z2b5b974ed9d1981e9eda323fe2b01945c2f61837910e53b6acd55a19ad87f1c6f77359174d5123
z3ef88a46b055736d37ff8c4638dcb7d2d8ebac304ef503275d22579e4c2bf3c1972cd38d046a02
zcee773e29990b08f03d1fc3ea5203fb40b0c799a591a2f15d0f60189449328e9dec835bad2bfba
zd60c1b703ab87e2a8a4dbfe9d0577b7c0c08515c07ce322d0cdd2d63fa78886ac6e5e9be73c1ce
zad5b6cc0e39f0e58d5eeae85fbf1958b13c9ea08692989c4015d09870abf9f0d60d1063d3bd8ee
z6c45a4c1372c2a6584e07f0e8ae3764cfb17194d75c067aecb627f1f2706525b105b0aa489f526
zea358197b9e8ed8574c3b696f0c00214da15c81039e4d71b10316227fa6719d7fc6e1f3320005a
zdc5ea8defbd69a8b7065971d21421e44ba8a80c2b8fd270f99ea5dd8103016229cdd80dfa330d6
z8ca04c05d7ee6d714e555cf7b5ffce672af80815b8d9df113b596e654fd2a5bf8231a060088a2b
z39c607202de38187a7836f6f1479f064b282c140252314e0783f809d6e9475c58ae6c800e62f2f
z4ca550d47117b84f77e51842b780ac897fb3c956baf0a34110e844fc411d5011df747c6f36e1c2
za400715bd123a952786cc859e9492cbf0e806c80266799d71bd58dd287a6fb0b7ba9fbf7604118
z9e51c404e45e13bc0fa5a7d79a346f02ea965507d48e702b1bef87dcbe874c59e27ce2d9545fa8
z0d28c927ee44dfde020e62e784642cb997a4553e3d122f7f735356abafdabc97b243ec23b598b5
z050c1b3b9023a26bfd0641e5c3c6e1af26d95832051e8d39b4a6e232d94b7a4f95ed6837bd7760
z29f61e1260b1853b36dff26a56094a978e8b51fefed5e0fb018612dd559e5a902bb9f8ea5d7922
z0c804d3f38df38b6beb5328dca1c2f5a51ec4f71697c1c2b0b54fdf30344ec4972c62995eafa4e
z13c45f3b1559abb1e71955af55f5e01acb9e3d9d372ddbd8516ffb9a72208be83f365ad22c0040
z6800aa8dc6dd2cb42c31b2714d7e20187eeb0e9b263b310dcb4efe186cb9e16a2256f5a056d42c
z109ac1473c10c82be66680a3a73b58054ad4d6558e3beaf1fe97604435d02a385313b36d154a51
z6873392d1e8df79864f7befbb4a7433fd58b1bd1cc9c9379096386c1ad6d26de9486b741623d59
z8f064edba8b5efe187931f730df99ecbf4d792f93bf673cf0c352d2a33dbb76c1a5a6e39f4d2e6
z0a6c81500f6ca9e4c5c25ec7cfeb5b7ebc92dd99801a13b300062c1e37780b9ec43b1130fe7303
ze0fbcd005f646c2aeac7446377ca59a669f6ac80d8863aa252d4de9cb9e730ba7c5a3b6215a1d7
z22938c54e5d4c69bb26e45a781630108631df6e9e9b23da4167982ac7c70ec0c852c60422c8804
z1c4a304f51200f9ab81b4c1c71e6bb39bb57fe707394dc1dd3e839d6331c2362206ad88b6c58af
z70c22a880c19bc696350e61b2b01a48614bbdbbef10f562692d202e950a256c45a67a6b26278df
z49df54fec7d98ff5049f34313fbe50a23cfc4d27aad7c20c8ac0d086c2604a02d09b997309d30e
z3a1eaa9eb5ceda28f1963c277a985956eb334cb4436388d84f33cccb27a4bbcea22747a51e6906
z77025a7e730c61c54dbd0f8d88ce7046352f2c90cf655aa6065c56e7ffbc229a8c19e59c22a188
zcc07c13224ccbb49d8acfb098fddc9c9694d3674a15adac03607a15acb9ad4f7d6cfae83dad0f3
zb044268e0cf5c70a123099c6a0eb28250fb121583d7d4e94e128a54b5889bb245e38ada27ac5b6
z4a5187a2343f9c42961c8bc2cc6f42ad44c640d6edd50056751898ffc97554499246334290cdac
z907039bbd650a24cb7fab4f7c058ba10070daf3ba85451be3d022e331b57e24e73789c2ec4814e
z9c59d46ace949c1bf827d06aa57c0ff2c2738734993c9f56b326a30b9b2307f67ada7d622b6811
z5ce7493858471558f45fbae389a3a828af99118b8259a846586c60c495b9f5b30cc792887cbf95
z917ae00006760525b575c352a18f5bf665bccf7a8698fd1b3cc4f4807d7d8adf350fcd2db08fe2
z14430411812f73f50ff3531ce9eb9ef3964b1afff31e2ed66137d16b60de2f86da12af9881f9df
z071875520f4155db6761750fb7c1fc453db46656fcc8caca16f07cb48e064682c667513d1630c6
zba205ae143563719983f200beaf7ba1850f6db830b73cab00a1bc499e363ab459ab642e3935983
z420e5116e7906e40256dfaff37b91762ccef461db8c05f5ceb39183e6ac714d5d56762f0125e75
zcb98a36fe31ca0b892126c143fda5c63d39f08cad39af327901b32a97a6de6c8f95689bc3072db
z7077ad29a5302be78c4c08456f398fede4f9ac4d28132e6cae0cca8d24720ef93a60e49b53ed72
z45ae1ee0b897f490682519036e5b0441a1d8e5fdfb14257a83494e276d085f31bda5918f4c4285
z9fc9cf2c42f410c4dd335691703953557fd5f3764991de3b8c04c2c157cfb1f3b8deafc9510215
z144a61de85d1b2a45074eddd7ef00afb6886557f31c9c9d14a104ee91b474d7edf6dc95f5b266b
zd81938f5ca5e18a2cfc6111ea5ed1a4ab080d0ba0768b98bbba425dea6d1aafbb292473dfb73a3
z258d3624befb76073f32f90d094a21df59caf893d0960f1327c97de93ffb54e3b04bf21958e079
z9dffb031ad88bf1dc0b5bb2c835d1d599c17be14b3677206a6764096b476e8a922f44bbe5a5cba
zb5f79b3b5dc942aa48081ccfc1cfdd7a76d70abb78b6779bb52ea3c8c798a88f3ef8c9f0bb34b9
z5bde3c3b85739662b625b7fe50ee5d7d38cd98fece49d5e9704659e62a6fa2b96b08e2f8c56ec3
zf273714cba12a7d53b88a0268db33e6b51fb5ff515cc306c0d74ff47ab31013cb3a1d869f68fce
z9888019d1c58a6d3fb3b161549f398c031872d49eff08640d22bd9f9a60c533f55d72c3f7f3b27
z7b3a64f8100d7c6d2d5af7b435d13f7ff4079753929c8868a3388efb290c780d066a180ec33c97
z0519f3c32a36bb06c913bd8a2c1cd909c278dc8dfa056701d9fb34eec42f4ce74fcbd965c6b203
zad95c96e68fb93f0139193e301bc59758d7ff99c22e663fa48058ddce6e5760b5d4784a6600f3f
z797b6a15b7e5aba7423f061ef031e9da655571106b3d052dbef5913bcc6bb6612369c60a64210b
z28cacd9b5a786d9bf07eb35cdfa19657830300aee38c534c0fb132b227cd5e9e5f3d1009139b09
z0c57eeeccabb08684c370201608de85d5e16cce1fe2016341029dff9c6b0294c13146db711da32
zb03b24f994fe5c1faf23de703c5f0e9b63095b5eb4f9673da2776fb02fd8f481b9485b816a26d5
z13d2b60b1ac8658256db91945ea96a209f24b46f4e23b274aa874e76e859c6850ef3d5a6d59110
za18a018553d64dd61929fedc6ec4d7a2749a571d0b9246d502efa02f96de451ab83c7656e77d63
z2e96bc55647a6d6ad4b682e7115fb9c6db3a2b442d8e332dbfa555fc704a29f666e28ef1526659
z8db751321beeba10fc91d016bc23337f6b41a94e036644a8549866f939bd26c3338bd7244d6919
z0c06ee958034cc20de10f95ae2704396514a98e2a5fb7c8d4a50debcb85efdb7ffd4cb3fe247f0
z7ca980286d257727f3559c88be4562395e075228fb59b0c6ad17cad408a040614f02e55ba23eeb
z764b60902fc31963d2389c0185b819f339d5a047e7188bf564879b58a558a25c921cbbba6f39da
z868a8ef7c41f2a227d669edb347570c5e890d70641ad24e19612715db69dff9d6e0784f3d0a05f
zbfc8cc541163e45fe2621810da0f13876939c3789efcb3e8f79d7e44705a39c8c3456616ca9c40
z6e07557390b55340d0c94c7418dfeb0b1ca90a94b2cea6a54009a1462fc22129894dad18031ba4
z866ac8d28a2c28d44f0f0f0a4b73b855633d51cf7274a3613a8277d3c0d7f009f7eca1b0ee1f6f
z622070506bd7d988d74f6b48ecae195438c56e97483f19e9369513b1883302a956ce61d388a286
z5484c8661434cf1caad8a094ff9f37b2d9188466c2f91b8305989b42d2fa76ec8d7aaad0c186cb
z99c4290bce020f149b8a38ca9532c32a2568ba295a57b68a13addd1e35e53ac3a46faceb875fa1
z8bedcde27cc636a907ec5a57d0f7115d30e3bddebd7dbd66f5611d7b0ad0188c43c173c09f78f9
z886f7cd7a9e5f8be90032d5404f130b260319246f6babffb48571f6186eedd0b8b0323abde608d
z90708d2263af54b2a0468836b9493106731978b0acbcaa4f01e0fd69ba049d90fc0105e9dd01cb
z4d26d0f5c0a8a7a152f4605b9b798abf3bd4045f2ea13854c5e6f283fa8b15f9e84fa97525f577
z64ee01e7cde6974e19a80b5da3ccfd4abf1659baa473597d48b76be4e90cc1e5c229ed9ed55d65
z54183633b404bcb1660dab902e95dde29cf1b17797f0d531dc361a2c5712e6ef6c7606f41f536b
z253c3bfc4ffe09bc54ad96578513abb5e3d3d27913a370e0f86c18aa10be97264c8d759b82b2e6
zda9bf35a102ca0657e2b6d24c6a5dde306a294ed8a5b5bbbdb1303bdd3a4d1f6ed448ba41b8590
zfb211ac30c66ddae9f37b602025f77b1ce8305fc172c2a8c77e3021a8f0d9628534d323b967dd5
za60836d5264a1fbb69de6b387d718e301e03ea5c00e3137e342e723e4a5f4607bef0febffc1bc2
zef52ecc99778be02e5c7b6684cc863702d3ae14e1e1631772899407745cb1dfba0392b62295083
z9cd9313acf4d60577dbbe34da5aedbf52cc8122504239f1ecc89a4d92c3110138a2a4284449af9
zdb4d923b72c50dfa40a8a75a919b4737146406bdbc6946c2b19ee33d6cb5698618fb3fe8579ca9
z93f1cca1b60ea336f61ef276250f325c28567db6ab84de59e949c0b988e39ccce0266a8bc88198
z54b85a3e4200c2e5422fce035406648c1fcbc1f194ba9c40297a8c17c5618b4fa2be4c1e27e516
z0bc3a354289b7a61374e4d3651699807e311ee73dc1e440f3d5124f6731916240c3de6bde0ee3c
z7f9663afd56f5dc97f49d35a1e89f6d0c6a404a7a3ea0484f980e977d38c26d3cf32554f8e6789
z450fea8679e6a981d4e5819da90907b811337389d586b38677ad287a68ea3ea796ac40d815d9ba
z78cd4be68ece1534d3dc4b403e570768f6c30bf8427069eb9dd0dc3f0854648684abb7f370c423
z897ff654fb95e42502f304784d9833362687c49d57a10e2df4a24fd3f9c714cb9c8835027d77cb
z02c627bcb3edaf7d000c7f2deb39c408999e52d74d6b3f7eb61bc81c15ba5e64bce396baa52552
za8aef160e3cb28d55f0a4a02f08971773c001df4c3094a8b05f8a72ad028d4f3f070b9ab9ed4aa
z45896f245b14ba7427cdafdefbc71e1557183146af359c984b13e4fcb92f352ba2dfbc5233b96b
zdcec518a1be6beb87cca0c7a93a2a74a9e4cacc3ba463ab09ea852e164dce7b4884097fdff0f70
zfbf2abddea81910c3e45e185ca616f5233e77450e00bb9ef73cb0de276ffc2ff4934279cfc15c2
ze9c26f1922ead521d73e04e9cdae6d61b0b52a3aef315a19a628d7c6ba2f210418cab4bc055f5d
z9633a30797394e9cc3b58625d808aa00da8de99b13e0b907ccc38952a19ef7737d6d38a72c0d37
z6149b2e2d56dfc00fa4ea76ccb4fbdfa528050eb533e72fdb0966b17e7a99d51393f312c3da217
z10c6de7de982d55dd6bb93bb9e41d9ce46123752880cbbda6c3687b9cd97863f41844dac914b0c
zc82d8e809b03563ad495c495c8568a32f6305e4066fe5a074c751b16db7f7f5b9d4ee0c184b24a
ze7792e2a0feeb86d644522bb2bd3a26872960c3c753d55e10f95f1840c0900bca6ec10c2ec79b7
zfbb83748f499d78a6af4511bb636d402b2fd68daaafaefa0fc34049d35baa5d67c05f686abaa4d
z0f9d0ba93fc4c28301ad39701420b5f42d3506e5ae1a1344d3ac38b2d120289e6011a27b51b1df
z4f0925f86f01ae1f3b7e8cb00deb57f6e42aaf5a01af4d70ac372995bd8d4c0ac1ec6b959e0576
za2b4c3383ea58af38deb8d0798ebed18fb6b5ebfddf8654d0a95d12e26bf47c5c6d76915e3ecd0
ze59cf9fe8836d0f18462ab312347e2b24546d4f1c502784b9848fe7ead8bc3cc7bcc691eaed2fc
zb53a6ca9d992e072e093864072eb9e0e18a4fc0682acc5fabc1613da4934a82b2d0af873eb9cde
z4a45a2cc4639f7e3e2bb4d7c3a1cded0569ee410b0f5e32e55e75727e3de4b464164a956e58566
z2b5054b5a27c8e6faed2cb2d913b2e99ee808f57ac46b75ac00db842ec1a29592b57ae79ea37d7
zcccb00ec7c559422ff256f199d5f6846594b76e115f33a56b548b6f2707d0e60c2cd9f3864a184
z04a1b4be26d9ffa0c51c1b51c98eefd7e9e40d4a22035ed0a40487ea5d3c7b5dcbc6c14b163fb3
zc1f77d6a6fa144098c592fc92dff574c0951935aabaf2e78a9e921290c7fe1dfaf8b6d09fc1897
z10e20b6ce3d832141bf4eb128d69888239b3e3bac930fd40604bb1b8d105d4438a2bc176e7e16e
z200fcd583f7fc39cbb2089af119feea83282fad8194d145464e4705cfe937874e373b9cc664f4b
z792481251b2026b0781d9d7f002e0c28f94b430e42eaa7c8cb885ca2993da5dd0c1b16d7310e36
zbf7b83af78a0d0e86f0c08668273d578897bdbeca32d5708e556c8d8715f97909f970e2cac1063
z510281dd62de4c289448c5b9962a5153425b4532dea272786b6266545a853484d50f291badbdd8
za1c363c820a0685e766ae6b3522e34f165236a26b35e98b2b972433bf6b1259fc86dd2f6143f17
zc8a169a1016a6222e62c03709efbf8ce2ae6bc34d9db2e8f2800cf1f8077f0311dbf475e6d669d
zab835fae6f0b957c5a2f45d5a58282e6c208b25cef4cbf2c5c45ea71734cb45f4781d5c02f94cd
zeb4f5c38d7bcdd8d1d7c044d26b7d76d4269c1b20529d1f5ac58e5689f23c635539c74cd32bc27
za6ed81290c83680f8add21c0105694c4a99ee31c69813a95a3d0fc02390a7e173e4cd1db42bebb
zdf94da1833b5fce93f6d5f9ef809a5bb8168ecc1c3c4892a7deba3f2365e5bce7158b9749ed004
z9382475fde3530fb05a7d8e66f21ec2151c3e7472c293d1ac22e1fb4b3b55fea8d4e741f225078
z8cc440fb4ff8e6a3c5ca8e114dd3b190611c53da44c30b3e5c55092744c4dc3f3f260de008e045
z40d166593c59bd60db7ddad469965ed10013eaf6d5593d248c6274796e90994c37bc34186270dd
zbbed9859170f07f9e3809761e342c1aedefa9eeeec7665f809912a1c8c4931b5dfb903581f9c17
z3a70212a29606d3cea68196bc66f421b6188beb0edd879fd76f7a0f37bddab83f978a411264e7e
zf5b55814be0039d6fcbddbcb99a8dc684ee3c2af98a7a7d76a3913b16d4922c96df4b5660cdf0a
zb09ea77009234d6d8a2781983361eaf9181ea0ee614a5e9344ad1fef610e4c3ab0c147f127637e
zf460748f7cafa01a25f7ec0bf9b03dba24c8ced187409a58a8ba96bb934bf25ae6132130d0cb48
za48034606fc7348fa8cc2d113f13734d672108e58f8d665ea55d714da44fb2f762a13721ec0845
z44d3c3144fc8471dddf2ac1b5c336b6408046f07cdee2390a878f8c626098b943ee1e38cdcddc6
za041befed889729efce4c125e653171a2f36bc436da3f8d10721845ef582537e0306a27e86bd82
zc503a643139b8565b7c110ca6f59ea1c55ee4360313a1e4e23a6fc9e8333e5b9b05f9c762a40e0
z45456772623347b269557e0fec08d4fcc286235247b5624a26b60d33e048b03f91394df2e850e1
z6a382fbf8db3f0022b0475f0281d90610ff7c58d5e2e1cfe360fd00156bcf3c5657b46a0b16d34
za1c4dc9810a5c3eca79879a71e43c0afbb233d31980c171a54d5ff785cdc79432b0d39c8525d69
zb975de80eddf200bb36a00126f8e0291e93541d9684f7aeb698ef20feff3e3f02c7d8186d2fcf3
zd085c052a7989c48101ede63aa15b3c69dff37619251e9186f136121bfd110ee721003e2ac4b05
z778c7bbf8709e8bd1b89c5659d34c02997ffbb71f235bf8dc8f14c0322b6311050a1095fca6851
z37047eb14a25f242aab94929428bbdaa055a8ecc9cb710c3e027d0808840a5513c0a9d552fec64
z8ab6dba667d8236773f5f0df3430b4e5711346d1931a6e222a851f5fd030295b18c256d7b42a0e
zfe49c9137f0ce98693f847921357037a9d01e0de4516e9c7427a867659e418a5bf746e41066ba1
z54e49054b5fea00b4ffbe6b2197acea699f7d80467a30afc6feb42bf0818ed3f31add2b90959ed
z56ed3b84eb72f7e5b20886c14006dbe3be412df4d00d0a5299104c7d550c4bcc862e9ce8fb4fd5
z3e90430583d3b4b95943e4d45e855c5d06f13a2959f0c138f6af66e2d33d54c848af834603fa01
zac17c93c13bdc6e28216393375f271b3e321eb41ed9e67d00454d2dac41eca3fc5c773ea0da513
zdcb1a7747801c1db58f227d2239762f398e22928c85b1f37e8a4fc3c0655a4f33b65ac54381641
ze77e7bae16c46ad951a36fa9c54f77e8f45fbfc88639536591e903d5ada86eb39d9339c4afeacc
z14c4df67ac1a9d200a351bc200beda46385bfb1c2f86019dbe085f2e3829800bed9c8e8dbba595
z448414562d5a7a2b1e6da898aec60cde67649e131f143b7822d21fef42a0d132594addd21c5bc6
z970112ffb327cca964688bec47d045fb58a418ae237a2922fae55ec40909be547d63b04ceb1d4b
z4e7a579c0ed91ea84638e8e72009b067b8109d4205d9e0356f9f3a1edf2bb0694a89bb8e1fb787
z0dd6a210a6031aba09b9c7f1141a0a732e2d69230bce4206f24d5e3330beeaddf7aab4dcc0b7f2
z318505ce51674c266c32a6565a83de5870d52bb8f23ed0bb8f684c3673dc45a5f3c2d84c5d02c2
zd6ff30c1622b1ba7ed812eecbdc37016edbad75e8513cf8a32ef2d233f22c457b08d4617257c0e
zbb46203af9ee114949ff00d5cb77deedbf883697904d7e3deab1024200b90ad9387e3ed633131c
z9d5621831e872fedc80909d1161d3cc0bbd9a0efdc245f0c6e34d479b175f281514a602b574fbd
z500f14f55b57df1154118d8049272c1ab046482f3a425a331b0ed538743af97d2cf3d49a29ad33
zb288bceb408c99ec7fe30c9e4a70a2d00adfc2861d3b9efee44c36760fad552b2b85832940073a
z590f193f75c155da301be350dc2b0ab34ee735d11908ff9487776587ec3fe88eaa546d99f3c30f
zbe53d61545d4a0c6b03495db0b2d9f63876783fa964dc92e4887919a64699f565373101081006f
zc899840b33eb222f1319144e4c7056d87e1e07430a8a662b5fac82533be1a2b5f2cfeac7e5d785
z8e8df1084ba03bf3133b131f558275386f6ddabb4d6856da8abc5029a42939d789940280fbda7a
z36243bfae7dc61b25ea9bed23c860b2aeef48cd365de48eebdbd21fc6631ac0dcc7493d320811e
z336b2976a59e47b78fca8df5417137608c9f0181229c5d15e8e4756e920c07afd9af599cb90525
z6fe9f3731df9cd0a089a8c340360c41d78b0eca185e94036b0cbe32de90dc83b8d5ec6bcdb501f
z3b726a5d72b2c19adbedce9ff3f18ad24dd46aa3685208f2230f8e1ff1663f71018400d71ca7cf
zac78b76099c37a33d1aac89e92c91b39491a8d3e02200b8d1dea5fbc9406dd81a08494b60791cd
zea58f1c0004e6998e2a2dfcbc6ab1ef9f8b402a58c027abba4dff5a3a7ed938d040bbedbe3ec59
zc7e2bee65e51345d3257360403bbef45f99e01799203aa4798603875453daff7c0b9a87980d5a4
zb4455c52ba8a493f070907cce81900becd8d0ee92fe6196c89ecaa9823237588c733972628d1b7
z1ff7efd31173267a09cec9a771ab9cb313e5eebfd505fb018002a8d4c5a2e76c9ce503a55c303e
z4e50b56ef1346e6e780137a22b305b96f8550a1d126ac7a178b68821e75d57cef0e0f32d49633f
z01518e454e0d4887f3652861534b303cf6de3f98968efce5df2d44b409e9e4d390913391621e69
z17552f6b9b470786b94214fd2fd60cb80b865bc70548bc5e1eedfcc0b9950dd7122523912dc208
z8574168ce5d9b5eb018fe3b5fb50c71f000d80e3c037f0c63674e782772cdd0481ec6d0d92b8c0
ze0da5e52bd4f068644aa554d1734b00a54d2c53b6cebe42c53ed4f4d45748c848ab964992ae8e0
z85e3f49c32b4693035dd3e10dea968746014c052eb70ad32d17972f299892621bc831edbfa3a75
z300b535db0083a12beb569a359a9e577f7d6125606e5103da5c8166718b02425bf2c3475c015b5
zc79a1db0e069b2c2f147880c137c105d8b7956677058b4fc351241c09dc02481250fe2c2185ccd
z74f41780e5badfa4e1885c8e12e89befa704cbc4b3a18b4af2f55bf33aff3fba485a75cdc51d89
z0f80a2ef507534178c03bd34f91e2121268fdf381a47aee887a5035ba62054423fdcbd75f210fe
z8b9e25d5433b2ec4dcf95c13eb9a827f2296c1ac121834e9ab701d671d42e958af436e8bb84d71
z505d5f62ee058475d3380997f4a9f12e82ca3d0e0419bc4a0d97a8c0d9e346fc4bc6e1df6850dc
z14c7f7b2db0e2b37cd1a408dab4cc56c8762eb818bf2e094c56ed2b13c2f7e137b54457458913a
ze084ac54eca3dd9c19edc7c2912d60c4ea255da202390b1e522ca80ef027d2ebf0a8f20bba661d
z671bdf4d985ccbfa75daaf4d6829d40021389774d867c953ea391780a72c53ff01dd68d3a5cf7e
zefcf9646d18e2c7800444f586b88a51e6cd5ac2caa9b4d7d1c2a553fd4702ba7f00b9c358a21ed
z0f2443cbeda2f30c5227099002c3710a14855a1d3c54bb961085cb7987b9e40c71287ae9e5cf4c
zdd520c332ca359eb71763b8d8f2f8089b119a79b4a25aa79dee42b4056aee2e517a7365d4aa3c6
z8a165adb52286d3b0076e21c315de48eef329491da59d1adc1a2b6a1bfc35383f95e7e607c7b21
z4948a157b492ff18d69249cbfe54461b7b13587af9b2366ceb6826c663fb9b2c7928acbb9396a2
zce2a0aa329f1a957ceb6cd95f0f7d614e1676767e9c4a757f39a0ee80511f453c98aa46893cd6d
zb459daa0de89a4d234ea0ecc3bfaa4413b0b96cc5bcb5dbe9615fce91c924deb8d91ab18f623c4
z9baf4f9e3112e1646b69b8824f89f917fcc490d883ba95403e7897612f26785e024de9d1eafaf7
z22acd2d2c2062171662d23155dc66720584e0d71b6c4fdcacc50781fb6ca79a6bcd7a9182d901b
zeaf3f09a76eb5dad79af9d7d0be1bdab6cfb505d4c8eedcb948f7d77929c525ec7576ffd149220
z28517ef46c877e0a6d12bbf88058adbaaabe6d7f33e0b5b86c006a2ba5a3c8c3456761ba691291
zc44203389fe735f88a89c9b00ca151548b7ec977f39d7506184cefd727b29230c73158a234abd3
z846c0d8682e1d43cec109bf8b0014d99b12b8191860c268e7f381dd7fe13344d68a4348d0a1d34
zea841c437afbc3a593ac5fe3b8cedb51bebee13c30096bef911e9004bdc998a85fad6f552014bc
z884515983a5182831e4d20408d6c2638d1f7e273a68ae9ce012b8d1a6477218632d72f5476edc5
z362dfdd9a56f03c86fc73780b951e8f124b485fa99ae5a468e76758896063f578d4b8ba7f2e4ad
zd1d47f1d5fc68e607a80f16d4fc7510afa3140b2364c8b498e080841a34a60416248a4799714ac
z8a565976d4d91a5cb90031a51de0ab027ffb9c5c7d4a5a1706d80c7c1478e15aeec31a6c789ee3
z603339331528ee13ad16663a08c0e47fe320959c182886fe63d76364fbaa50412c0faa076535f7
z9388b2c6714b197696bc9017d51f89eed582051e012dedcc44a13c1f085398d2360b7dfb9be274
z1cf669440168a2709cb1f155dfde18bf250a24e7cb0a8282b612bbf5aa91fccb131c488ae45b86
z3cf72245ccb98c846283db223697f72f68f68b2e7dbe21ab69acc920fa3249145be8af953810ec
ze5c3675b26a6e17b71e30e1bdd6aa565a2385faea820282b774e47efefd7e571cc3b5e459d9753
z9471685deeefadf2c8e3039c440324629eb619610eeb8567bdba68a80510abf8fff9a3b8269547
zd7ab986ed328851a8de2d576f7ebfac44bc9882d872da99b373f0827c8dbe7da322eb022fab0a0
z1e4877c55102373bb8744220b4ec7a462518c759451f6cadf35d8493e38472ad657e4c2c8ef2e3
zfb1e5a3c3366c08326c471f492cfd9aaf47a31e471aa36dc2285a4bbd24966fc032b9fdccec49b
z9373a235230d1d141eab29c4a6c84c8eb33aaa4c8ee18257efac9a87aade1cd458c937b0be9967
z0c0bd6a5ed7e550b2bef7f397811617a9e43d081ae18d4daf444ba487490b801ebb6aa95b24a9d
zb76065406baed1f3594fff0879566a421dc082b23569684b1669b41d7008987ad07bf6b5d65b8e
z748f916ad745937547ab30d9746d11d981ff38dec39de14dfd62b07ed7251043d618df997c5967
z20737ea4b5be6d399c36f28ce516eab1a1385612a935a4a16170073f3a5bf45daddfc14dd40599
z2227ba05f002d890611902c566b6ce4023dfb2be7d264c14b15915c30abe03534c38217b8cbfbd
zf3ae70106cbca05aef2234266e4bbff54c365e3760cf1ac4d3e565c4cbb271fab2bc0780e23dd1
z27f6ac2cd1bd54ded93782edb9089ca8cbf192b0448a05741007c21bc7cb8bff704d3ba8c6d3b6
ze0c3bf8a1e2b025b9b3e4de9c23c3d5354a5e377055717ea5c89eb0399c2e2d25cbef990ddedb7
z795ffc47554711309bc2c4182151ffe879608594ab1b6ff2ecfc615c4db4b28bd9bd374abbe29b
z9dee9845c138c6c8f46ec925a4718e9c18a5eee6802a0fc5134073467921e73ff72e468e1c6b8c
z566a892489e43dbd595ee2361673f78e26af8aebef652b71207e31a3846df79d7045abe317be73
z94ac5401350a69f1d43c437609d9767d060baf8a49b2a181b831ad4333cc74cf819dbe14ed9f73
zacbb45def59fcf70c5709d85f89a9ae3ac9201b9d8f96c85a26c19a76f9aeef08a21390b4bc8c0
z641b5354c7efaf605a71edb05ec183a6090b3658b9cfa4f8b8a71d0192a3edc0711bea98efc89b
z109bb5a073f3fce0290d26cb183384aa619f25fc120788e1d73d03c8a9c69358b26139443caa4f
z584372d69eb3faf511993414d8ef3475547719abf7bebf299747f0bfa6db15316776d2fe17984b
zfd3bbec835f50770b6a7c78d4ee896dba244d7d87af292bc0f92f4e8b6c60366ce943d3378c3da
za453e7caf45ce691fea4d1392c8b578ae3f922771600733cf45e1a787b8da52558b5ab74e2f0bb
z3be781bf825b501ca67de56bcaac0a219a6b6d92bf4102f4957d795ebed8a73fa1a4fbc31d65af
z38315612ced89c361014c1e5dd8ed0b4b695e92426149829588d71ad3e9120994bb7e7917f91b1
z9e325797b81fa0a9e917062793933ffe97a9b0557efd89d527092b715ffe0a2200cd7814dcc1df
z575413d1c58f22a8389e0250fff27b5ff93074529549b6f1c8babef47e139e75151836b8b45a4f
zea4c85f7a5da3111e7384beb192ca111fc736cb617fbd08b10d3d5b4a4a1626df934c6c56cb947
z29f33d4e360f8b4c0ec8e14e30615736d94f7b29538822295deece962c2c19800d461312c63b3f
z7e1d07e5b7f01912c10799c645b40997f290fa2c047ba56b35e8008d40495d9f5d8a3a18f99ffd
z91d20e71361ed7d60059ce7944c43d0b91d6d413917b8993acd6cf5709006f666030197787916e
z05c71d9457713f6ae028aee5e955bcbe3462deca07ca4bb17b69e4c0b4ab2f9c689b3d0423707a
z4a9129e0fab7c0aea14c9e728cc31b61bb069a45449dd85c8b5a546764309103f447b5537443dc
z068c80e7cfca282d6ef9ecb891a886427de6ab3770b68d552bad5cb5fc3336fd14c79b4c9651be
z5466fe1dd69354867ec7f6b4a5558aec47997e181ccd85976a792c39177d4c60e8b9c799b4041a
zab11f57190860d7c18d60e83718025c26e0e916770f25d82a66692c6b258190c8f36f5a591e650
zb0361bb429c11abc3a1d7b4071d162bf9dea918360247040432ed4692aa120082145ff36780e6b
z6ffb374ffca639354c9ecf48b5b71791d830cacdbe35fbf5f078c996086b15944deb152faeb7ff
z69e68bf2fd12f54363981c1933b1f414af332db29c2b2beedf219b6253bb087c6eb13b446f446b
z136875e0f10be7abdefd99c216b3985bbd8b7719cb2d98994643c7b6c6cb95f1fbc25a3fbb328d
zf03cce7db909af53d041f93189127d3a883f633924801b977345abc8dc57bc548951be6ea9f5ef
z0dfac5b41ce27df9c340c940416aae11817ed12cb960a71a394272930a3a35a78b81e8be18fb2e
zf3a4a1357622b5f447f362674eece366f3100d1bdfabc9cd5e5f8a5c731493e74a0310c21dead7
zcbe088583c4ae565d383ac4bea013599536728e9e6c1d84040a41e55aa2dabae2f19fc30f58336
zbcd046d67338184d355b2a373ac46e0fcd0d03e39be61c3cdd32ff123fa0ee47a714e0763721ba
z5e75d98a2f6167467ef8c90ea5406a57608370353c08cdb862a4094908439779abd24b2afa6cbf
zc99cc1db3a19ac654d65d9ed5f04e46494d6a40d6504d01782e3686eed6ef1076464aba96b92e7
z390cc8e900aa2b53298e3ecd5f62af5dff9f7858ce1862e1bc1ee94c8d0a0e4cddad9f64acbe16
z9d584bf99e5088df0dab75598a73c55400be77128cb8b4bc11dab75205306ec07615844abe9d3e
za7b12eaec4f0858a1f71208fa59085a4c183b468c3eece163345e9282824707aab3aba5344033e
z77d943ec9b1ed6c952b30b6ccd8da7232add1ce1ccbee9773f92c6a3e0592c63f464f6b974f7c1
zafeaf1050f2185afdefb9fae61e2bb448f45b91215f7511481d040bc5db917c8ddbe370785da77
z95269bc767530c040f2b8e0908ce86d99a802c0d8ad2794ad738661d3fc60617988508ef1458b8
z0d44a08fb145ba6b9766604e8b2a54fa7f859fd01f88bd4007df03cfb5bae2790de17a1c07e642
zf0f790ddea4f6e63197aa648eebebd20fdb4d988d87f6e5ad96b6ab0e863cb6a059d9f7cefa282
z0a40c85efb82254115b31c6f66dd329e9e9779685c61ffaf9c34a3d7fa8670b1d2ecad117a0be4
z213d981ba9788698d02ad3f49086f2ee59088c8729d9a38b31931928cb3fa05fb05590ff498699
zd7a6623d7711194bac6d1931a20edbb7aa883045b155451722f3c6f892fed053d173c7197790f3
z25159720ca0cba3e65b3abab87382327166a04da4f83f9747f971ee94092a28398bda1a34e596f
ze83ec430984e0aacf0159ca3fa83bf894886600b930294b57fbd93ded9ea234ddb05bb4033790b
zccd42e4bb75c5eec79a263c4ca1e0347ef28261612e53858661f823f893d4d0940a65560aa773f
z72868d51fc57f99f14bcb4ed4e6baac6e6d8ad62a5e33d6988d1bc882ba6836ead47034d456b53
z29bd475d03d3e16c940255f4961403c730e434ac0417d077d853200a92be33d47b01512f1ba9a7
zbdbcd20fe21e9e5fa51fd6607df01c02be8c01784f45718166854ae54382dea7a89e70c4eb3983
z9b0a15e498798f74932d1b5e4042510b1c4c2be39d16c7b0729b4c377b417d6d22b7d8424d0b2e
z492c85d1592fdb85fdf4bb9fc4682c68f9398c6d3892cc57bdc831276413d2b0401e731ca2a1ba
zfd15b23abcc9facd89798424c9f6155096169d4118c0567a95eaebdb2ea910cd81e40464b1f40b
z626e85917cb5d44697723214e49e9468f62a75414961702d44bc0c0e1b60b96e6bb60807805ad6
zdca780649f7e377f265f859b9ff60fbebb0705a8ef0f951fc2da4aae65706c7555693c941511c7
z47a40955940e93e34d180441259706f8d48638b08e91f83541923c49e70e9aa9a74e5287e432ed
z88ce5f630a52e0284a962b1b4edc9b77408e30b9249365cb21a0a2d06bb2fc107444c974d96ab4
z5206937410bec0646db201f117a0e09131af4344aed805a11d70f73348b1f3af9394465f05f3b7
z2a21c66adbfcef9d51a821193593c371ef48bfe674bfaeb626e9ff1418e157ac4bc1e61ef42635
ze16b1b976565bbbc05b6477b85f6c3a0bc683a7bd400847deaee7fbc03c0de9f9bf7b980bd16fe
ze09a11d22e7b061ef06ea0a99da917a47c1224737b495d528ab6bd316b51620327f2c5f8b5926b
z9b37b6d0a7025fa3b2825731cec20c35e5e6ae80ac0a237b45ca2c0ff887d1885f70ae72e7eb2c
z76976dee3684946d9a4af1e7bdcea49156d72c1c16c36c45333ae75a446eca94d556b817f88cc4
zca3954eee4ab10e953646894e9d321d4aa22160927bdb756bf59f3a288c825e41017aaf03ea0d2
z052bf1387a702e977d65d6fd3a6a4be2124f1df044c5dca56d8a5e614a8b8c4ba4cb37e89a458e
z7dd4c13bffa74f52b0c0c124f26966ef00d9959da6fcb386a71d17ea083fc1bb488781ebec521f
zc05d4a2fe5c91cdf6e36a51c1c7e7abf8532f8a50a8e70e7803b8f70611d3d4497e211684a859a
z669a953f516c23be2726d1b94ce55d21a404c5684c0f9692ba2fd7cd775a3cb6a50993abd9d9df
z83daf6ce08104e28bd35b440b46184c1ba15709ab98b9e6e140700059b0435a582e40a33093c80
z60ed6771b6b7d123207227fb0863bf86fa4d73a88996460c214df735c6a5fc1f60733117a470a4
z385fc45228ce32550c52461935221088244665646ba0f31dcf6bf4913af1d82af6612c9fe74038
zf14b0bf3a4981b7352856d9d862d4da19c68d8b15e45ae5abe9d8da7163d048a7d6326e37f1f52
zeabc08bb961b510773e88f542b0466d011dbb449f6c43c460fbbb0f294d1938c1bf944ecdea98d
z1f39af0cd35091b35b7f106887cf78a6a3afd4f7f9bd7eeb5d740f7a72074743bfc8df0d8bc395
zb03a324d71442b5650563d4c10a51ffa4551b19c726eb220aeaed085b293868b7ed8283b76c26d
z9624730c1644172989742630d80dbcb368754ad02105560e81cab3dddf4c19f2631ed27943312d
z8debc4cd8bdbe42abd234de2760f11af858325f8a18b3d702706c25fa919460873eae1c48dba0b
zef1b685828b41150d29b9219ac73f2add39f8cbf3cb5e98d498c6f156ef50110b9d6816e32ccee
zeb199a0ad63d681d16fe5c80e6cf05e792215d562f84798d5ace78708c59b59aad94de4419161a
zacc996712b05142bdaf4efcfe79251f952cc59e367fcda72fbcca4fc33d0543c79dc82dd9f6e17
zf43ee67ec0616b2f89a1123584862681551e587a85157600a4496e0398bd8df6e816ffb9f6eee1
ze508cb60c98af7c955401723c1c16fc7923117ac0b418bedaf1436dd9a1d6adf1aca872c36cd09
z3c1ae4f25279f7fe10092feecaf8bd79d830e9c7631dbcb7f864a41c79bd1679f54fa099e6bffa
z5cf367ec81daa9f33e749b9c27b5ed5a94fa79c37fb7701f7c8ade11403b7db973c290b3fbacdb
z968f11926c5c7ca2d277ba68341ce4b5a5d5ad0d767dba6b3163bdfc01fced90e6c8c683e81a65
z9f7704d7407366804488ef10615335a42e65da95b22d8ceee91c257bb6af9187f4a9812ed044a6
zc148d7e84178053ec7a2ea6f2ad6f325ebe346d359c4f260b19bc932f9cf642f7f3f59e09649a8
z139883dbeb6907fdabcec791acd4babca7727bea014f2b71c4356909088c12d2aa45b823b754c2
z842a931074abfb955cc8bae11743e11f44bf4b8df250a3988b51a5cbcebcd1bdabfa5f51ec7fb0
z35711be244244dd1668b63ee0f3fb474536a937b3315db69d0f2cc244fcc7fb75259a1ccbb8503
zf5cb24acf86cb602e3ee161abee3e171ffdd9ba11deaa52bedb7295cb12ba577f79eb65b4a5069
z6deaafb4de79d5d8776414394f81d25c7dfbbd37a9cffcbd1e570706f91bcdaa13f88e124ec9a9
z1718a1432713b79044c9050e7361d2ff298aa4af29b065323faec4c75cfd11d01f224cc6286423
z011e1dd565e70a96f5297e0da992beb915c0f410485c8208c9fc7a57784d654a67a28080da566b
z871d6a84475a4eb3cc45f54c169123dd9966e04f1fb87033eaf3247c5c335aff83f623a3b08ded
ze5deb2d3e307eff6183908c6f4ec500e44624be09037b469eb9ad77b5b93014950f0035295e3f5
zf77138c0c27a6226ea8120ae9bd82642efbbda6a3394020d2ebf75206bbe2a5816ed187136a17f
z5d1aef5771e5c0cc7a80b7833330b617918b1ea1c7a0f88a02f908a5b143b0228e8caaf701c032
z11712f04733a17466030cd7b75b41a2767da1fa4af2fea6f1be7573f1fe1f2bdd39631b8f57e3c
z69e0d90e24f3b617c96ae31232e6079557f0d159c4aa3f7c35d4d18c86823bf2c12cb04f672cd0
z33e64c099a6809aeb063701e7d1daa2cb41078cd0e138d6b540b85aab8c61a4b90e78b3c6ccc57
zee3995227f8a6afe78fccaae37828153c132e499ac94084635d4d8b29d29bfc2537761bdb1d97f
z0b43d156d63364bac76e23ce58d2facc8c8c27946fa1990a3dc259cb4d6abc05921999832aa690
z0257d27e5e00b0a7b9900752622d68a62853b222e5501ce9c7ee8c30e96d525a88e148273292f3
z81218c05f2ca8358bd4e53099628c25496525e2e2123f7803a054bfc61247dea37568ebf38575d
ze6e4ad2982f657e3827915e902f065c4f3e8bdc72389d809d835939c802a9640678aa46a4a23db
z562336d36a487153d6030a352c4925a8f4d8779c5b72c9a6784fd3c55ff7851bc31085f372d86e
z8b528589b07f205e28327723a072c68bb858b1212220a8f51306349e734d6ce736caad7fcc910e
z510c4ba2788835b59e9619567872e0660047ccaf2eb24a1b72b1476a33bb8a98bb32b52035f132
zcfc3e01e40fbd04d65d79ee1b36ccefed0dcb38266aab194ca79c4f935a36924107ec06be1284c
z9b28cad3262bc1d1d8704a2cc0fb20ee85f539c61390c89afea0671bde9f740162c99249b930b2
zb73a70f0c9be895b45fde6a5ca7477e86343595edaa1ca370662432d6fb199bff2d05f57aa51b5
z725280804159dded4efa956d6acb48ac7ee933f18afae3e95b59aea1e941d657bb98d97b690a3a
za8dd0a16c7d588be79b051472c2205ae1ddfaa91e955cdb54995d0aa11f84d9679c19279edc4ed
z287a4cb07ecb1917b85a6badd1868de55fd123f93d3ab803e0b3428997e629666b2c5d2f3714b4
z20ae5bb540188a2b9882056b926cea0b8668c91c655a3f3e9c3f761c4fc926c5b69641c72a2847
zcb8d1746772d197431549ca3d505c50aa6aa04abe02b5fdc74937ce32fa7169b783303956f85da
z296ae4d2c6ef2777041cb9c72cab2cfeb82ee0d078518998066759c40d5d40271d58bdf38132db
zbd882531066015b8e50710337ca261a93e4cc6c3f3b1f069876f8ae830bf1fe48be004d367789d
z445e042a93c5a46f7e6af170edafc928d1a4a5be5de887700eec3d90d3b1561673e8fd836dd9c7
zc5c6172628e7e01c38769087f4f3464e2bdeeb72bd9824a507c56ace94d0f24903cc206ebb2f4e
z3d4b4444db3aaf6abd9ad7e9903dc45c4b98d475a79614e6eca50030e0bac3477cbe5693a8bebb
z2960dcb63e2c5d7c64ab191c9b6775dda35176ce19e72a2c5916950fb5efe1620a7d7a49dd7ae3
z71e546d54f4902bd025bd8a31f8480395b426b7fb42bd6416e5bda0411f60cb6f3fcd678facefb
z7b01241c1b5ccf86d4da021c8f9956d1fc48570487b2563a9b7f5ae5b81de4c48c4e44be48a7bc
zfc99bd0d650cdfbb8bc8eaaa9fa417a64eac69af9cc05dfcdd20b9ae3feaef2f25632f3a261512
z6320ae2319dbc1aa5b2e8ede35e3ad82ea833f67cad882f795cac6902f5ea4ea4767b0504cb199
zee23b04cf8de3edf2cc3c82cecc4506927bc2d72dca7ef3a6c79b8999c30c6d71358533a3e6e34
zd593ff7d7e4e72059e4e0c9a4acba8de9e9ee52ffdc959c07ed8144ab9d2d2cee3121352ec2554
z9e5b95c72df107702d2c90bf963a3b7fe8ca3ffbdc21616e909504c784097fdd95e332e955ac2f
z89892bceb028d272222ac780a35a210dd1d42b0eee0594fefd4d0f4954043acac59db6d14474ee
z05b53bdd774ca45b8f1421aa7cef4ae666674bb42b4618b80d4fa57bf566e3a9ee1e0961b85610
z20b9340cbdd89ba578496dc0f0041201aab2b1a2ca308a560d5e8b03c71d42d533023674ae15dc
zdf9c5970543d5cf476dcd9b94d50140e97345a131fe673ce0b35b3ac0b8c4c33ed59fa848afe65
z58acd1602a6eb55fe95bc224704325e344bd8e4122efa66d3ed57bd9ed7faef1641929872d96c6
za6c6d3534333e5791e1dac9bd64892f6f2fa44478ab2cb579ede290b3e43a529aa949988591cae
z2de0b3c91ae861b9af73eb7a0b77c7760597b6699ae5b71a2ef0a691328cc5c50070071d8939c5
zabf46d41046e21f330217c387d3e01732bd78a899b72a81ffa1ad67170b168e8c6b995ec9fab26
z5cbe736938be1e43b3d4821c81e5a0f02b708033882f0528e3b901dcfaf94bcaeb817fa2e1e1e9
z98d1dd0cef3b9e203bcd9e4115e9c761e258ff9df0db4ed5ffdecfd2e8a0acbe9d33ba1cfda36f
z89826db4dd8f3d5fbac04170f9f1be14edaf539775c32d1c352b8c43a0b4c2afc8c5ecadea3615
z480106bd5981bfee2fc4da84ee41245c7fbcf2eba333ad46b816ea1bd67fa7e4ac12cea6e0df64
zed399c51245c79245ac8f7d707c42ecb768502212b9ae490298d67d3f5386ecb2ae070cc7b158a
z259ec4c029b42a81cf306126abc9122657eb0fb973da2d51aeb4c94841fab98e0005fd39e92e1e
zd764679f59db56ba4cd04dc882a1ad3286edea045f05f24023995531a947cabb2d8f06ab68a94c
zf09664835e67e0433550ad78bd8f164bb223dfb9cf9924efd11a1dee29f4da4fd1bfa91aca943e
z3ffcc04d27f07e829655b01bc783c74a414b6f5d1f79f05e31b1027a257aafb3777f1b6fb03e47
z637893aaa243ba114b13a7665bf52ad470c117ab379cc16321e7a011c2bd4ca9d5b39a5f70be7e
zbd761564d8b5f225e2d1f16297fb2aeca2f6fdc54a022f3f7afdc0ee1bffefbc08cca41c4fb271
z8e05c67a5c45391e8be3116e029cba861a2a4a846425b775353a4eb9b9deab1c170d29623260b3
z3dece0862af20f1b84a0532bc4fde0459bb8fdbcaade8d4e75cd92bfdaaab4035e0fc260bc01e2
z6bf1cbe1db6e57c0d5d24910948b9bee2c52c4f8461dde18be44cc995b11aa3fdddd0ce95c2e04
z999e38841bc367fc96a580696a56625886530d0b759abe660ab43f37d7bf702194b2e7a435afbb
zb6c84c2b18222c3e561cac56da5285e52f8a932045e27b8fadd4c5597e7b9ee6db546b48f916cc
zfa2b69aa24d47ba49b6589596b5096768d780665484d2c3884be026b1648dc63b570620c9556b0
z0994c1f3849103bfe4124930108726f2caf39682fbba172fda9a344ecfcd14d3eea91871ce49f2
z138c23d7988f8dce8ecd6e2efa43b4c5a5e3b4f42b745ce51bd9b884da792cdd863565256f343e
z027496213bb1650f1bb6d188f736dd8f6fa3d54ae412892c7bcd478c891632bca86d9289e8d10f
zcd047f2227781e94fd09b61e4bfca0600927f9669013bb814ef021d432d3b7ae6898a8bd191121
z54b090fa69d1a0fd4aaa17e5b380fa3b1885283d974b5f32309bd25750f5bbf0361cee99e8371a
z3dcc325b222e35c9ea1c9d20b59874bf7ba778aa2e63eb7efb28150a8bd4aff5cc718bbface2ea
zdd17a6590ed8f0bf5900839c4e60e805e1a94d9b9d35606da5a825ec381581d078baa77f2587bf
z09326de36d0d8e2b053115e553cefe5e3e181975dcae3945ab38b711e1bce08fafa74daa8391e6
z13ba62e980c5ef01d536d5bc4a62f4b2ddd6b7ad580057afe0bdfc84832ea74dc437dad3f7afd3
z1df3a2f171242a805e32c82f5fc20d430b49d6dcb55832eabcb890071e1a5949aaaba190b58961
zb56701b5b8d61d738b847226df21f74782fdd4801049d97acef66a958bea50fbb7c9ddb211f1cb
z5b7c34b55cbbce243132586afe5239c21eba900e63e7528f4249d6e3b842a112845f309838902c
z180051a18c23790b000e0ad7745d37ead7e0793182a932a0c36f9dcf350ffd0d9ea430485d1dfb
z6160c250618c49d79ce5b86f2affbf7a0614cf01eebbe1a1689ac148c8301e5096150a25d4b0a0
zb749d97faef8f6bbb09a818918661d9be05e4918fa98e0077df1fed52f185e379b3aaad00940d9
zceb99207e9d847557bba3b8a48198a8a555e62694627d41f808ac50d16a42bc583051497d23469
z6cd5836b4480ff94ab493f56684f1ea098b9a0810579a7b817b2bf6af1537a7e1081b665c60a43
z5454ce83ebab6b2325e97ad38653227c3f6981255321d78f7ecfda8caa9f4f71f6a00d4daf4e1a
zc265dc598b4f42fa1769fa4902ac9a43506a16b5929bac8ab9b08b83a0b394eebdd3db18ad1212
z7db341a343c7136c69ba2cc5bce2e01aae9ed7fd5c3e2b3031c9fc351ac3ff6582bb9c807ed8df
z0a7b508f5ce522d2f749c1f33caf72f73202329fd30fb27353dddc0e86cbcb6134f230996fcf36
zc3e348099a464071d2cfed3ed4d8e224365615d1a9336ac5a7b9c3454fd29eb2f3754443339307
z7845e3c82bfcb5019202135ad696ac79ce89d594f13ab9c47137963d734da07999c252b4072858
z8723b35cbe1c07c07aec105db33b48416219fd3c340a4f65ee756ebf668184a0b1a67af2296876
z17e3b6ecf03046f843e9e1068a2719fef10747f1d1500ed576f98afb076b20d2aa1e62593b0ba3
zab783e7a30c28e6dc361145b8b8036d60ff54eb4877995445eb165cf1f89c6aedbb4a33c72bc09
zf215be74c8df286bbb2addaf542a10eae3602b6d81ce8e417a0e1daa0308818f3c2a49a09899a8
z1f639988b96e9992cdb73bf671447ea6288960cd7b2648a999e98fb7bd10fc4a05aaa83c451e41
ze0bd5e5060ed335072fcc18f00a6a68a36c4b4a32b170fe794245e50062666de8592e3fa47575e
z24e6783a58ce6c2aa9c0b2583d504b82d615e1ba0dd326493324e56aeb62a95ad192e49307ccba
z91a44f19122285b628ed14623a1ea9608451677449ba092c4d2eb4fd44150142d6de823cd7546e
za5515b7d25586f0648f5be7e064ee9f92ab305bbd2298e6526c2225ebe095cc1a7f7a3f6c093ef
z0c789dd6a06585eeda00faaa7476274de316a68314b3487f425425ee1c874778b67fd9579b35d4
z72a498939245abfeb53ac122c300553d0ba73c4831d551579fd1905ea0f7cf39e58ce03e0bd3c4
ze34cfa01ce6366390838c6f5641a9745c79623c195820f8f1507e2923e6d3c662ab4bfdce648d3
z2aea08d328d87137172a1ccd66246e4a29ad679a5eb02e1f5b6555a513ea80f9d078ea0928a768
z1383617a4f7a04dfa1c5af9d00fb27002998f24340aa35aaeef659a615b741bb9719c97d3cf9c7
z9cb6cecdce265e04a1fc135f4a83560515af0bde66d038d0936a3ab8bea3c658e735d8f8683e08
z0ad452d8c8785863dcf4d5a08823faab8dad2e5a092fe23012907510be5e8496048f1c927af43b
z61744f509d06949043ca0953bf7d4458d638c7f409e3108f9d2ecad71bcace7c15a75563420ede
zc14e6fad0a284a78d74b0ef12c31f551fd8a46131ce012efd74d13e14cd41e5accd3be5fdd0b74
zd342fc5912d7dc88814b890557abb16d3df2a319fd1421d0843862c818e5642a83d1f4dd5dfba4
z3b982d166d5cf20e554796293150d27ef18aa9ab6c9432124d50b924b12516a563db97a2ea08c8
z9aeba0ef95ffc2a6a19e832ebb2e7123566c59a038161c6adcc9736d4e1b0126a82069e60f8d9f
z4ab8e35185f75c3db2c9e44410d90f8519d12f3d1556d30338a744c60c805d8790be304ece88a4
z6e84b4d55118186205c78deb75ac64a0f1881f2cc0b8f3f7d31bcfc9b4a74b16fe27b7f9a076d9
z000290cfd6f55f64979557b6c3acc62cb933592e590c53f77944948f44a0087deb39c18d4708de
z897574b7243febfa557f432f063fef9884b20ac7e1e3443a7b112c133e63dfa7bc95af71a5a081
z6c12dbd99330a18ddce7da67fc78b0a00fcf10610235c2c8350b68482cf8386c40a6c9d81ec4bd
z65e5b42aeb0736ff58e0660442cb04d0c62a0db4291f1bc602d3cb5e1e574c88a5b8674b5b4b6b
z99e7d68a1ab5547a7e7698da05f4cebfc6befba0c900a9e60dc18087f8b562843f1e80fbf8c1b3
zba8b42f14d39f7735b7e420dc156ee64d4ddfcda084ebe97cb66e7bcd6e66a1f918477b194ac0b
z95bf8535c7361f54f575ef1670d39046cc856ce06e057b13e676441522e9af4e9a4140322ffe65
zef2cebbc220f1a18836095962fd19a91efc3ed5c4b486f7345c6a27288a7eb6db415b6347e1103
z54c6c154ee154084ffc5e4b3eec831581eec74539fd9efe243d70b6837661a68830a2ce24ac377
ze620672da37406d7d9f0836b081c42b15fbe5b1d5505f07eac9241e84235882a9e5d62c26f2228
z8a364abb104f5ae692a53dc76055b8bfb41d374a84029ab7b89d1c48d440b9a49764d36b905897
z0d523e5d42b19d0fc9bc884f60fc59222525d1df4c918d484f0d685751c08187feca54a5ca1c0c
z22b2f04faa0fb3b4daf9c082dfcda8ea0a1c915f742aeea19208ec443541e45675b1b3611c46e9
z9718d3713a63d0973155ac958ab8990edae8454b19106d3d8ddf1ab206be20d05a38e28045555c
z36dbfa8246bbfa92b8cbc396bf8b7b3eb3fedea946191307276e463999dd4cea67c6c4f88b832b
z40d12d5c2806c9d58d0354dbd4500193a915fbbaf49eaf36e479536fbf2c9ae833969c9e80af48
zfd05505138cf5d9f26c775deec5539401649ff0d4c985dd467382dca9b452b9435912bf34f737e
z3dc3847336a46c33c9b5fd9906dda07078867d56a3737ca3849287ca1b34c254f4cc06233fc96a
zaf4ff5ab84a651605df617945a96d8a2b1aa73a6020ee891ba57df2f42278e5c89a6633b793a60
z8ee64ee69336b97088b9d5a3781e6db373fe7212fcb0cff2d5a2518dc3b8fd2c615c806602938d
zbf7333fb1d95cd37459aaf65f12330aca4b1558bf48bbd1471c29f8150f38eaea904e03e24b2a9
z5e52d7de55f9a9921524a9405eb2c17e770d1f267601a8569f4aec0add5eb1884f20c569176b4f
z5381374023f6a9c0f9e09c188b6d20d662b2de4c658c1d50065c29a696171e8618bb101cafb21b
zfb1e6fbf509ea969fd8ae34b52b1688ab99d3d85e2e41a1480e819609ee31bdb968d6760fcc635
z49df734628d885e7ddf8c22786f681c530dd7d0bd4d1c109d95eb54e8a207bb3014ad0cc6406c4
zce35c860503eaabbb7812f376c6576312e48b96ce7776ee61645a28a99898e194ce7c642f8cc85
z650415d110edaeb7f9cb69e3701885c421197603f5139a0a4098d21b0df0ff44299c8f73f02dad
z801048a864a16ab216dc37b64465c5b88010f55f03dba70f571f99181a3f118ea5b63287e6b76b
z10764520dac0e1971966e3b3491f24abb088e1589e3c2b024a3ebe431908c33a2807b0e465f169
z85694394bc638c5e5970678d5e7f13d5e59be43a7872a45ec0e1e59f32df6b6aec84425f4ac53c
z2273c3fa59972a874f517729f63b5ed98dbc0699f8de185ef07c6f94b1abca3568d56405bfd9bc
zdefd416da38d6460856230e23c237416ba79fdbcb6f4f6369790551068b52ce7ced960571a72db
zcb818e9730bef017a13e862c4c58214cbc8aa7af11ab74b318b9ff8c06bdc14d1ce688f00b8895
zc46870432d333bc16a3d18e46077eab0d1092e0c4cfe79e991ecca814aacf9818dd8bd85b3eae3
z14c0bf0b0988f98fc6e84afd65330815cc3d05f8835aad3f6ffe8ac1dbb7968aab302f270865e2
zcc465fd2c470dccb008e40a9b62a3ed38f612705c6f4e24fded658e8fe5fec361225349551b765
z44cc946781019a457ee1f8e636d67c7a709961d60f025312691d07daf235ca5dda89ac92b020ff
z8d460973dbce4e7c98af8e5c804a97cd4c16543f01a68613a885a0c3f96dc64edb8384ff6985e1
zf7e77b6d7973c24a41340652c79fc1a45907a5cedea112303daf5c0279c1007c8dafe7d1f0633f
z046e45cfa02a59e590405ead7ab78585fd70da68aa2326b331e0861025f4e6cf990d4543cb9def
z497fb2608b1db5cf13651a320d5331d04bb1d748259300f6d8ec1e9444e2bad001368a5119d405
z477af52b3eed19e7cafa424b450b6d4446002929404c3b6d223b9989f6df42ed0917bf3cb47535
zd75df5719fc95d2a479dfe60f0bdd7c58bb6cdb378a7fe919928933de1691e770d066e60e0cafc
z247dce479b55372b88ad50619f0377212d3291edd852f1b35f54e5167afb94b14cc3d290e11175
za31e2fff044821ad32831f024586fa1ff6d281318afa5f0c73bc8437aa522d565c70d296f5d89a
ze406e2e4ce1015577f11119c33d7dbc0c1a0521968aa1783a6e700a69748eae652aa27cb21ca29
zac5a62aabeaa12621753750312d5aa62a5abc7b5f363559cb331107cbd9c19240ed92d3a14a122
z7b14ada38a610f1c613fd918ac1d391e15d665ff1a16c7b767cd196351aa26cd6cf639896d737e
zd734a52e33a0e5016d9619da01ef6fcc8d51a629554730f94354b888255103611db5bd413e4c30
za703205685ce270bb9780aa4e2d38257a66c06c45d6d2d23085aacd11929474b099d7e5952ab02
z82590703b06e85ced0d36fd29cfec19b7040ed5f2221e3fea19a74e9f4f11d5eb78f360df0c247
ze506c251de50e36258b07d77c0b5cd1566537dad5ae4a2a2facaaf80ad79d0213a4755dc6a303a
z03140474b6c9b95c7bbc3921d94a855117a579159a44f7cd34cecf3164fdcf1abc1363ab98fd90
z6e98568367eaa8bfd5102325e43578961c93336b4f2edb4ed1a8bccdd4b30865d1c655d4560e70
zb22c6b3a5f6586707b149b301f29240969f6e0ffa031b2b7cfc695f8367a33489db014c73305a2
zaa58ddafdca849c52951ced399d546f668fa84e5a9ceb6a15c0fecda52f325a64b97f14394b606
zc5d07c0c9e636687fcdb290f82c4aed3088a48bf21fcecaca78884de84ce4a4c14079ef3824db3
z0c799a7de740addc776c58be4c01f4fb7760a5afb4e5d5ee77e23784e67a0f7cbb0bbdf11ee1e3
zf818e6ecf17c8d66fa14875370708d4a4f22fcbe54b474f21fe747777e63aab4209b86d6ff8ad8
z5f6c1fecf67d0ebd8bac4315f7471fcd355128bff657c39a4fadba98c74db13625c31cafd2534f
z845890f38e57ba8996bb7a1980e0a6451900dd2a77c8ae0e405336937f468ddd476ce09cd9cfc8
zb765dcccfbdc561ef2423d450a09aeaa8cbe51e8c5e6337962e493dc25ce0c2f6f9a09fd0a39d3
z5bcdc1cf5b4eb775d4dd386a45306889e5b65c71944d9d2221bfe766cb480690ffc9335b0733fd
z58d333576e24ca637b0de62241c4a4294b8d4af009066227c2f82e3c86f8cbe5956550f29b18a8
z52a67a3d15b2924c6c4aa01c4ef1ce9bfbc276765a5d5551b776992efb369b760c79f89223b53c
zd6c74e883cec65a2e63c5964bd4142e22281ccc6abb4f7889681fe3ff2c54f7b7d1b55e06e0662
zb280d2cefc53c5b30dc767ea29da3f0e1c31250ad50f9aa774c087f0dac013c3fe9c1f6f6c7d8c
z563e2dcc01dca46f3b0c63c6e9af938cba3d5c560191ce196cb5175488ca46e7bfb3be9b2fdf19
z2a9ab1675265ae74518203992d0d90e7ab408977de917dbcb6e01c7027721566c4e979f51a3895
z211f9bc49d44516097575f94ec6e71e601e64d4f2b648d457f277c25ef0f230de389ef6970e0ef
zde9cddf3c3071ba998626da38aeb4f8d7f03edf9c3485e5856c8c23efac9b7cfacc11d88e82790
zd76e46f08af49b59c241cd579ae1f97fcb32295505bc27af04d24188a35ba132f37f26ab5eb075
zf3ab248a103ae216141a2788c81caf035bc2254dae7e817d28bd72ac1d4ca84219aad87b70684c
zbb910d853bac5923f664340c23a5211ad66a3db205fdccdc295db5d9c4886ac0efe48616f3435b
z8515dbd694b64b9394cade4b97553d0ea0d3bc99c9d6e8103df754ce73f28c37d482d202ab5469
z0ae8ce0c8178417c695434d5139e3461f6b4d5f1ce0e340df511181fe53e979078bfaf7d213cf9
zbbf4bdd019fc23e8ff6e02a4355e54c5599874a0184416a9800ce2cbdf9141519a00c3698c4da0
z4b2e9ff0e4a5385673ea53bf28e69511e292019eea481f877e521f3996d08a0069b9cfda18c155
z7e97f8b55f0aecbed5cf2711d29ed18707ef5e54cde3f7b1f996d6f143cb8863972ec0b81a1130
zdcb4e63d45ddfbce369e46c696947eab5fe6923ce1d35b3caf951e4d485b3d81fcc2c5e4fe1772
z39c003bcd5e384808734731f89987eb13ea3a25ae71c77fbb7e6fd6576896cbe4cc60318f53da9
za2a981d9937e372e0866df845e3ae665c80d98d2d798f800e13ba3149ae75770d6f721e822b85f
zba320e9ab23f8517f21b199599380472c3ad35b98033119d33c1ee2b4de1ab48d50d99afcae06a
ze39fb96b269651664adc3d78e080092d1c6b221c59a5ae1e7c9099377d925e50092b6c857d2239
zdbf8d34a67a587b1140794d89577dd062e84acc18a2c68177cdfd9ad1877bf2921f1c0700b5c19
z54d636dfcd0d6c48342b891f99ce2cf242b5abb247a00a664ca7d9dac5850e51caff11ea6bf1d3
z640f5f971bcbd3067d6b81bac4bf099e976816cf6af6e9c9fdad6ab4b631adaaf05b365e676a4d
z04456a53c79f9e651c20f9b2368d8e7c569d2db0efab6b613d48e8996d2a9034a295c641208bac
z445f7ec6c0c2713774680cc31d90fb67071424dd60486245c9bbf6a14ae523605b3016e315b5d6
z2551bcdd7c5d54fdef1a802e4c98dc41d89ff17322bb7a68f355dbd89097492ed74ead719beaea
z306c658e466878f4c0347a9ea5ad76d0fc99006a35692219246b0397b01c73191265c8b4bfc6c5
z4e2a7dad2337ca109d59dfbc756246c40d7ad2c04e9c9fb1bec8d0c887b00a00130aaa9376a07f
z19bd5c0a4483dce72e43d5a69a173e89d6fc84cc5a19d7bbb73d8c96b9fba91d7b5f6c526cedb4
z987415206d3fd795f50a9eae3ae2783415d4bec79fb5a2da255da15c6f51f0340ba688bc26a665
za54c6936136ef2508252dae8f7f3e1c4749f5e2cdbe3c1796645bc647833c41213a0c63c6dd4d2
z624b8148cb4474cd7c61aa9eb775d2a36965a1914017ec1fe5914099e3a19a3d3123305c3fd48c
zdd811396376080c5a5c06bdbcef9b885f33f8cd412027b03cc8cbe7ee6b9b883c9def221f565b5
zaa581a05ba19b02db1718e840e2bb7689185d6cb2efb02647a34b236af525d0da8a9514a34d0ae
ze044f8bae776735bbf16178019ae1240f65eed5edf5e26255ea6906e449d54388ffbab0d54feb2
zd6a4cd0712ccd008c1e198520b61d5283efea1b9331430ee7242e9a16b28a9af205892bab0d887
zc3beda8b09d1eb243b526042c0cc6bce5c8f0c8229572d64f1c79ca12b749cb3b4133fe5e46019
zafb28264dae1410da892fd74d74a16d7a11dbf0ab4ad86a57582eaa1075abb015d343d711b7dff
z1ea1229ec102c95ccc762671bebb0694c2ca87fe4eee8045ad84fb07d0d258e634a22fc9ee6996
z0694684b8ade1ab06c563524c030f476ee105bdbf304afabd5be3daab451bab5d17dd8f659c2ae
z0167e4d0cd1fc26eda91d038a40f69c829af1295f394255ef9698231c33aa1422889cdd64b60ba
z98b4297ed05d2852fa0ac1fdd0f021f890965188726e489c5f49b3836a4ead3f6128df09730e39
zc476b74f35b5949a637545b13f97d44b36d35a34e6c95cd7a9f509340a00fa757fa358eaba2324
zea65701b891b6653acd7f2357a2012298d0f4d6e6d12063ace7b15240d0062fa3998ccd312dee0
z5bf5c2051163cf6a5e078abcbfadb11954376c8cd47c457ff3a443a499cc3c7fe4ec512e6b2758
zf90f143d67c2a09c4a2d449892b3389c9ef6053dee706b3b288a4f040d4ad9ed96a7217f76fa83
zcbd1a007aba0a0ead3d96a22d31dcc2b797c08f421293dfd0a805de1ea1756222582943044713b
z8cd00dac1c0cdfb93f3c38c04ce67fdc6e299e3d7ded51356d95a23d0980ef7c68985264ec805e
z1b7a8d73418805b5c5eb6784326abfea5d47fcea512c0d2f257cb9eec21c65c7c95e4175a93960
z79d7eef7b72e4059d94f4907c98a4014f30910e23fdc0eed79d2dbf612e42de0ced5818f6ea457
z0ad7a2b5179381913bbf5762a1f2946fc75b9e4808cadd14b6936f86c9e091b0d5ad25bf4b312c
zd7c353ab4dbe78707d4ea5bec764a021f7bf1cec657e61a1fcab40f2df1d523d27ca71d33bba0b
z9aad15d2084a633906200bc1dcf55b4d7941762c1d18d296ea1ea2b94bf76598d124ebb7411757
zf8c79365d7f1ea2be63a554249accb68ad23d178e0a546797d34a7375fd1a01ae61e34b22a1e15
z85fa8479d7e3eceb19892fbfb8339df7350b659f89f7dcaefd4eddbf4cc01e4a3ac686fd6aa113
z613edf5d2b08d9876e7e7e2203f1afe7ea5c73405a32bf80d2c3a08df0a91d3eb2ec5ed186e666
z80cdab37dd1d4eee8b075daec85126a4cdf0ea0b601d0085d53d9d39cf51b3efb620ea1c78f523
z6a55955494d06b574e6beaeca580d347c433720c702fe7e0acc12186e8c1065655bf4cec70454c
zcba35f18488a981e5599f4bdd08444c82a6459cbe83b4ce78c76abcf01506f0f36a7b051a68d51
zbf73d83b9bf94951b5866dc25f6f02711fd6071efeddbab9705b895f75fbfe32385f8c210f6c5c
z7ec0b75f20272684cf4f3afb9da01faf5eec72da56ed7d85a270b7bfe6d7addc345bca9df92d3b
z9fe8f09e56ecb906e7a4d188d1c3885b702488fbbabdc57915d1332d21e21b4993b06d340d2ab7
z92861643dbee81e8817625c6d0a854dd00468db17fce13702f2362299d0a6ed3ee9fbc5e5582e2
z0eaf276e8aac95563d3c2664b2edd62ee812ac4b107d7f7a85a960b57baa9c2365945b270815ec
z680d3dee826680b23b379714c2ca327eeba8cf844c47584b89c4aae50019e85eaeed5ee8bdf284
z9c3bac5d574470b396a9b5e02a8df4f90369d632881e0ddb5bc1e68dfed8de4dd0e7790d5dac61
z83ce1ea8b1eebd637a37d990a9a8651ab00aff688632d7138342813be65a355286ec7f61e6a4af
zb5f6651c90e74f7e0084bf354f4573c7d943c9221f28d4fd166d74918cfded1200c97032319aae
z31d1940dd76d95cbc6ab3f82f39508c9f8848f6dcd633272047c2738a68271769c9188dcc86476
z9c7b281e91aae2a6030979f79b968e96a724c9db0b51af98200c292315eff4084b087c5b19234c
zf08fb94f3c847532b54e7bec71d2b6493906b08ba15ac11cab852266c712e586c5111fdf11dbab
z1029983e1004360d437597b68613e5f357fce74149f284b4415076fe4c3caa4e3f788a0cdb7fe3
za67f7f72137911c594ecf4b1891b32c6acb23ed8ea7ca15efb45cfa81a7d8bb18f0d10b527b28c
zd61ec24fde8a389a616cbc11c826fddf97682f1fb530148bc91c469b73685e51a0fede5a07247c
z32f743098d49d616064e9263a9d362c6a1db07d3ffe04026c48d59454f09e182c6a6f4b4f6b651
z59aefc952cbab763f04a6e4ffe556e41a0c7d3e9d0eda37d412feaed1d8bd9e357c2a68c7ac4d5
z29eb9081605478eedf4e78f134d8eefb2e09420cf8626dd645e5a6cc1d0715e6c1e7bc0c896aa2
z054c8ec1e0df88021e200bde4e6539f98ac9185da0040c72ba54799ce90caaa37c7b0dbe5f4180
z307ca26c3c3740d16f51a76941ebf64ff60427d9c19eb7287fe91291411faa8f48d2e80e832bb2
zd4073b6f0217101f21ba786239a724908a4aeb632e39f6ca53d75c3af070320caa815874442e0e
zea0985d5d079bcb5d922830efd6849f372b9a747a731a37fa14d60636d09ef031d776d4b715a75
z0bf3b1c0adce827168240bc2cdc756a919b22b327a4110761732ce2f43925f0fb250aba751b92c
z2b66a3c583b8f4f875fdafaa55e62b7a0174269720b4288443fcebb458a336419dedd46058b999
z0d832fb15f36146738bfd5ba6c739a0c44044e07d1657749d02320405cbb3c345f042966f75696
z54867f87f99b26301ccbc61f07b608bec049c4ffc2cec8153433a56b77e8d504a82079d167036a
zdb3c8027e5d9e107275ec6ef33d07aeb3b7d71a35e3fd8e80ec8d4e0526e5a4b65b053b58ed4e7
z046ef2ee213978edefdfeba406b62b4a3aa96d0e3dab01a9d278ab6a07c6b98fb927b0b107e924
z8a33658cdf5c5d8685593d7d612639f9598746914fda14e09f3e072c73a493b809dbe23bfa21fb
z26f0d830bdfd8fc5c25faaefd448ae2ff42c23338e15c2d7dc3f412c9f46cb6a94489d06207421
zff1a8a9625f046ac937d509fc83ab5392fee373d6cc44d39a711de3d8c890ca662a272da3e8ba0
zd62366b712f1c2ba1a3c10da00be6a73a9f005dcb5d5498bc7fdd107be8981044e52cf694cf28c
ze66c988c76b9080501510aa96730d54e3a82702cafe184680b07d0be6183a7831169be46e61ad8
zbd2e8680e2ecec1b8c6dc71f549e2250e94bf285a77943770b01be3651282ac21e05eac42c6bb0
z4bde889136efd3659b5799d64c3821f40e1a1940858a79c2df36f3b4557220c4aa8dba7065b91c
z23ad020307da5d466ca44c297b2dc320e31ff7c15d19ae70a2d874591a4a51289986fc1d7b528c
zafc12716f77dc06434a58afebe78d66b46853b9c2ee8ceb40adf48202a30a9fde0c009f7d79c02
zc9da60801deeb13f8bd8b95ada1970e58a1903fe52a5dbd13795812f542a5e3b88417a42017eea
zc3c10886eb5f3870014e51310b15b88aba0e2be774e23be584adce00bae67e723f2f780f4dea8d
zb4fa4508a5630f2c9e50c622cf8a7264916c90f1835b2396dc9b72f9f6743b7d7dc61af74dd36d
z5e1bb0d656708928d64a95ba29be4163f6a6a05c900842b08ed6b5e65c25cfba80ebabd2ea92d4
zbc40316c9ff1e89d5b0bac025adfe1e48b00e7cbc8da5c4f958cab9de56ad20cd2b01aae865807
za6700eb5299235a96b5c0ea02b68aafe283668967618315dcd130b6d99eed91f984124e82d4835
z0343b9d4a47180828c8c44ddd7bf3b27f0f26bf4ef55099eb7e9daafb6110163e3404cccc7a5d8
zd14cab95102bb1561a1b1b356c8f667f4474d301ca4df95c9d0afe4792e8a39db3318a2aa88a90
z94fbfd7d05aeb22fab79c8a3876cb6a85f0427b6da3f2282718df1b74b7dc080fafa8e0c69f787
zca07e6f77acccc3ea195f12f22683c62a4e80e7165c0bf3d22e8f11bac50ec3c719511606090e1
z6136a2e55039cbf0b553c68556a78c06d6301ddcaaf71b972ee0095e76870c624fde0c222ede23
z9770c33db38e6d298ee2b8d8c117ee52c0b0057c5424310c337ac477f8f9b2e9107ec656b52858
zf1bc7d98806b2c54318fa6ea6d04742d82c33b0f02089cadc13e002942e7bed32ff88cbdb532a9
z36f9f14434b94ddf2d7b35490f8139390f809ba39448e25f63acc1f6b12e6f4fd98000d1caa352
z0401b3b58f83e6c76770935d0857fe7e0c8a428f2f93e839f9a4f9a280b6c718353bb96878bf91
z5f4e1be5502b0867fcdcd1a3a9fcebeb3ea273842d1c6e57c2ff7d028405b904d687f316c40b26
zfca00dfbae6d2b5b0137bd4ca3e75ac049fe78cf0359aa6040b005675f41081d09a72f82ea3b10
z9eee9a0993930b6b247f66389daa735d9abf59cf593c01b0653698b92f3430dfa87157d94b28cc
zf50aecf4c9c2bf688d1740161c561026dfca24e0dc5182742dcd14a523a68382af33bdea7c676d
ze82b9a44cdbd16436ab47b63944ffa4c51f4fd4c1977655ff6743b9e5c8d663f84d5e9ff077266
z202b6b0b48aee9c6410ea665f1ca122d2deb19232d66aff16a63d82d9f5a291e30
`end_protected_0in
`else
`ifdef MODEL_TECH
`include "qvl_usb_1_1_logic.mti.svp"
`endif // MODEL_TECH
`endif // encrypted_0in
