-- ----------------------------------------------------------------------------
--
--  Copyright (c) Mentor Graphics Corporation, 1982-1996, All Rights Reserved.
--                       UNPUBLISHED, LICENSED SOFTWARE.
--            CONFIDENTIAL AND PROPRIETARY INFORMATION WHICH IS THE
--          PROPERTY OF MENTOR GRAPHICS CORPORATION OR ITS LICENSORS.
--
-- PackageName :  synth_regpak 
-- Comments    : Synthesizable RegPak (Synth_RegPak) contains same
--             : functions and procedures as std_regpak. Only one of these
--             : packages should be referenced at one time.
--             :  
-- Comments    : 
--             :
-- Assumptions : none
-- Limitations : none
-- Known Errors: none
-- ----------------------------------------------------------------------------
-- >>>>>>>>>>>>>>>>>>>>>>> COPYRIGHT NOTICE <<<<<<<<<<<<<<<<<<<<<<<<<<<
-- ----------------------------------------------------------------------------
-- Mentor Graphics Corporation owns the sole copyright to this software.
-- Under International Copyright laws you (1) may not make a copy of this
-- software except for the purposes of maintaining a single archive copy, 
-- (2) may not derive works herefrom, (3) may not distribute this work to
-- others. These rights are provided for information clarification, 
-- other restrictions of rights may apply as well.
--
-- This is an "Unpublished" work.
-- ----------------------------------------------------------------------------
-- >>>>>>>>>>>>>>>>>>>>>>> License   NOTICE <<<<<<<<<<<<<<<<<<<<<<<<<<<
-- ----------------------------------------------------------------------------
-- This software is further protected by specific source code and/or
-- object code licenses provided by Mentor Graphics Corporation. Use of this
-- software other than as provided in the licensing agreement constitues
-- an infringement. No modification or waiver of any right(s) shall be 
-- given other than by the written authorization of an officer of The 
-- Mentor Graphics Corporation.
-- ----------------------------------------------------------------------------
-- >>>>>>>>>>>>>>>>>>>>>>> Proprietary Information <<<<<<<<<<<<<<<<<<<<
-- ----------------------------------------------------------------------------
-- This source code contains proprietary information of Mentor Graphics 
-- Corporation and shall not be disclosed other than as provided in the software
-- licensing agreement.
-- ----------------------------------------------------------------------------
-- >>>>>>>>>>>>>>>>>>>>>>>>>>>>> Warrantee <<<<<<<<<<<<<<<<<<<<<<<<<<<<
-- ----------------------------------------------------------------------------
-- Mentor Graphics Corporation MAKES NO WARRANTY OF ANY KIND WITH REGARD TO 
-- THE USE OF THIS SOFTWARE, EITHER EXPRESSED OR IMPLIED, INCLUDING, BUT NOT
-- LIMITED TO, THE IMPLIED WARRANTIES OF MERCHANTABILITY OR FITNESS
-- FOR A PARTICULAR PURPOSE.
-- ----------------------------------------------------------------------------
-- Modification History :    ( Refer to Testbench for Validation comments )
-- ----------------------------------------------------------------------------
--   Version No: | Author:|  Mod. Date:| Changes Made:                    
--    Beta 2.000 |   mkd  |  07/19/92  | Beta release
--    v1.610     |   wrm  |  04/14/93  | production release
--    v1.700 B   |   wrm  |  05/03/93  | Beta release - no change
--    v1.700     |   wrm  |  05/25/93  | production release - no change
--    v1.800     |   wrm  |  07/28/93  | production release - no change
--    v2.000     |   wrm  |  07/21/94  | production release
--    v2.040     |   niu  |  08/16/94  | Exemplar Synthesis supported - infinite loop
--    v2.045     |   niu  |  08/18/94  | Exemplar Synthesis supported - exit statement
--    v2.050     |   niu  |  08/19/94  | Exemplar Synthesis supported - static POS 
--    v2.060	 |   niu  |  03/20/95  | Fix bug in To_Integer (didn't work with 'L''H',
--		 |	  |	       | Unrecoginze 'X' 'U' in vector)
--    v2.100     |   wrm  |  01/10/95  | Production release
--    v2.2       |   bmc  |  07/25/96  | Updated for Mentor Graphics Release
-- ----------------------------------------------------------------------------
-- synopsys translate_off
LIBRARY ieee;
-- synopsys translate_on
use ieee.std_logic_1164.all;

Package synth_regpak is

    -------------------------------------------------------------------
    -- Provide for mathematical operations in popular formats
    -------------------------------------------------------------------

     TYPE regmode_type IS ( TwosComp, Unsigned );
     CONSTANT IntegerBitLength : INTEGER := 32;  -- Implementation Machine Length of Integers;
     CONSTANT DefaultRegMode   : regmode_type := TwosComp;
-- synopsys synthesis_off
    CONSTANT WarningsOn     : Boolean := true;
    CONSTANT DefaultRegDelay : TIME := 0 ns;  
-- synopsys synthesis_on
     -------------------------------------------------------------------------------
     --     Function Name : Overloaded "+" operator
     -- 1.3.3    
     --     Purpose       : Addition operator for logic vectors.
     --     
     --     Parameters    :     result            left              right
     --                       std_logic_vector    std_logic_vector  std_logic_vector
     --     
     --     NOTE          : Addition is performed in DefaultRegMode  which is set
     --                     to Two's complement. 
     --                     The operands may be of different length. The length of
     --                     the result equals the length of the longer operand.
     --     
     --                     Any overflow condition and carry_out is ignored
     --     Use           : 
     --                      VARIABLE a,b,c : std_logic_vector ( 7 downto 0 );
     --                      c := a + b;
     --                      c := a + B"0101";  -- c = a + 5;
     --                      c := a + B"101";   -- c = a + (-3)
     --
     --     See Also      : RegAdd, RegSub, RegInc, RegDec, RegNegate
     -------------------------------------------------------------------------------
     FUNCTION  "+" ( CONSTANT addend       : IN std_logic_vector;
		     CONSTANT augend       : IN std_logic_vector
		   ) RETURN std_logic_vector;
     -------------------------------------------------------------------------------
     --     Function Name : Overloaded "+" operator
     -- 1.3.4
     --     Purpose       : Addition operator for logic vectors.
     --
     --     Parameters    :     result         left                   right
     --                       std_logic_vector    std_logic_vector  Integer
     --
     --     NOTE          : The addition operation is performed assuming all
     --                     operands and results are in DefaultRegMode which
     --                     is set to Two's complement.
     --
     --                     The augend is converted to Std_logic_vector of length
     --                     equal to the addend. The length of 
     --                     the result equals the length of the addend.
     --
     --                     Any overflow condition is reported.
     --     Use           :
     --                      VARIABLE a,c : std_logic_vector ( 7 downto 0 );
     --                      VARIABLE b: Integer; 
     --                      c := a + b;
     --                      c := a + 5;
     --
     --     See Also      : RegAdd, RegSub, RegInc, RegDec, RegNegate
     -------------------------------------------------------------------------------
     FUNCTION  "+" ( CONSTANT addend       : IN std_logic_vector;
		     CONSTANT augend       : IN Integer
		   ) RETURN std_logic_vector;
     -------------------------------------------------------------------------------
     --     Function Name : Overloaded "+" operator
     --  1.3.5
     --     Purpose       : Addition operator for logic vectors.
     --
     --     Parameters    :     result         left       right
     --                       std_logic_vector   Integer   std_logic_vector
     --
     --     NOTE          : The addition operation is performed assuming all
     --                     operands and results are 
     --                        
     --                     The addend is converted to Std_logic_vector of length
     --                     equal to the augend. The length of 
     --                     the result equals the length of the augend
     --
     --                     Any overflow condition is ignored.
     --     Use           :
     --                      VARIABLE a: Integer; 
     --                      VARIABLE b,c : std_logic_vector ( 7 downto 0 );
     --                      c := a + b;
     --                      c := 5 + b;
     --
     --     See Also      : RegAdd, RegSub, RegInc, RegDec, RegNegate
     -------------------------------------------------------------------------------
     FUNCTION  "+" ( CONSTANT addend       : IN Integer;
		     CONSTANT augend       : IN std_logic_vector
		   ) RETURN std_logic_vector;
     -------------------------------------------------------------------------------
     --     Function Name : Overloaded "+" operator
     -- 1.3.3    
     --     Purpose       : Addition operator for std_ulogic_vectors.
     --     
     --     Parameters    :     result            left              right
     --                     std_ulogic_vector  std_ulogic_vector  std_ulogic_vector
     --     
     --     NOTE          : Addition is performed in DefaultRegMode  which is set
     --                     to Two's complement. 
     --                     The operands may be of different length. The length of
     --                     the result equals the length of the longer operand.
     --     
     --                     Any overflow condition and carry_out is ignored
     --     Use           : 
     --                      VARIABLE a,b,c : std_ulogic_vector ( 7 downto 0 );
     --                      c := a + b;
     --                      c := a + B"0101";  -- c = a + 5;
     --                      c := a + B"101";   -- c = a + (-3)
     --
     --     See Also      : RegAdd, RegSub, RegInc, RegDec, RegNegate
     -------------------------------------------------------------------------------
     FUNCTION  "+" ( CONSTANT addend       : IN std_ulogic_vector;
		     CONSTANT augend       : IN std_ulogic_vector
		   ) RETURN std_ulogic_vector;
     -------------------------------------------------------------------------------
     --     Function Name : Overloaded "+" operator
     -- 1.3.4
     --     Purpose       : Addition operator for std_ulogic vectors.
     --
     --     Parameters    :     result         left                   right
     --                    std_ulogic_vector  std_ulogic_vector    Integer
     --
     --     NOTE          : The addition operation is performed assuming all
     --                     operands and results are signed Two's complement integers.
     --
     --                     The augend is converted to Std_ulogic_vector of length
     --                     equal to the addend. The length of 
     --                     the result equals the length of the addend.
     --
     --                     Any overflow condition is reported.
     --     Use           :
     --                      VARIABLE a,c : std_ulogic_vector ( 7 downto 0 );
     --                      VARIABLE b: Integer; 
     --                      c := a + b;
     --                      c := a + 5;
     --
     --     See Also      : RegAdd, RegSub, RegInc, RegDec, RegNegate
     -------------------------------------------------------------------------------
     FUNCTION  "+" ( CONSTANT addend       : IN std_ulogic_vector;
		     CONSTANT augend       : IN Integer
		   ) RETURN std_ulogic_vector;
     -------------------------------------------------------------------------------
     --     Function Name : Overloaded "+" operator
     --  
     --     Purpose       : Addition operator for std_ulogic vectors.
     --
     --     Parameters    :     result         left       right
     --                    std_ulogic_vector   Integer   std_ulogic_vector
     --
     --     NOTE          : The addition operation is performed assuming all
     --                     operands and results are signed Two's complement integers.
     --
     --                     The addend is converted to Std_ulogic_vector of length
     --                     equal to the augend. The length of 
     --                     the result equals the length of the augend
     --
     --                     Any overflow condition is ignored.
     --     Use           :
     --                      VARIABLE a: Integer; 
     --                      VARIABLE b,c : std_ulogic_vector ( 7 downto 0 );
     --                      c := a + b;
     --                      c := 5 + b;
     --
     --     See Also      : RegAdd, RegSub, RegInc, RegDec, RegNegate
     -------------------------------------------------------------------------------
     FUNCTION  "+" ( CONSTANT addend       : IN Integer;
		     CONSTANT augend       : IN std_ulogic_vector
		   ) RETURN std_ulogic_vector;
     ---------------------------------------------------------------------------------
     --     Function Name : Overloaded "+" operator
     -- 1.3.6 
     --     Purpose       : Addition operator for bit vectors.
     --
     --     Parameters    :     result         left       right
     --                        bit_vector    bit_vector   bit_vector 
     --
     --     NOTE          : The addition operation is performed assuming all
     --                     operands and results are signed Two's complement integers.
     --
     --                     The operands may be of different length. The length of
     --                     the result equals the length of the longer operand.
     --
     --                     Any overflow condition is ignored.
     --     Use           :
     --                      VARIABLE a,b,c : bit_vector ( 7 downto 0 );
     --                      c := a + b;
     --                      c := a + B"0101";  -- c = a + 5;
     --                      c := a + B"101";   -- c = a + (-3)
     --
     --     See Also      : RegAdd, RegSub, RegInc, RegDec, RegNegate
    -------------------------------------------------------------------------------
     FUNCTION  "+" ( CONSTANT addend       : IN bit_vector;
		     CONSTANT augend       : IN bit_vector
		   ) RETURN bit_vector;
     ---------------------------------------------------------------------------------
     --     Function Name : Overloaded "+" operator
     -- 1.3.7
     --     Purpose       : Addition operator for bit vectors.
     --
     --     Parameters    :     result         left       right
     --                        bit_vector    bit_vector   Integer 
     --
     --     NOTE          : The addition operation is performed assuming all
     --                     operands and results are signed Two's complement integers.
     --
     --                     The augend is converted to bit_vector of length
     --                     equal to the addend. The length of 
     --                     the result equals the length of the addend.
     --
     --                     Any overflow condition is ignored.
     --     Use           :
     --                      VARIABLE a,c : bit_vector ( 7 downto 0 );
     --                      VARIABLE b: Integer; 
     --                      c := a + b;
     --                      c := a + 5;
     --
     --     See Also      : RegAdd, RegSub, RegInc, RegDec, RegNegate
    -------------------------------------------------------------------------------
     FUNCTION  "+" ( CONSTANT addend       : IN bit_vector;
		     CONSTANT augend       : IN Integer
		   ) RETURN bit_vector;
     ---------------------------------------------------------------------------------
     --     Function Name : Overloaded "+" operator
     -- 1.3.8
     --     Purpose       : Addition operator for bit vectors.
     --
     --     Parameters    :     result         left       right
     --                        bit_vector    Integer   bit_vector 
     --
     --     NOTE          : The addition operation is performed assuming all
     --                     operands and results are signed Two's complement integers.
     --
     --                     The addend is converted to bit_vector of length
     --                     equal to the augend. The length of 
     --                     the result equals the length of the augend
     --
     --                     Any overflow condition is ignored.
     --     Use           :
     --                      VARIABLE a: Integer; 
     --                      VARIABLE b,c : bit_vector ( 7 downto 0 );
     --                      c := a + b;
     --                      c := 5 + b; 
     --
     --     See Also      : RegAdd, RegSub, RegInc, RegDec, RegNegate
    -------------------------------------------------------------------------------
     FUNCTION  "+" ( CONSTANT addend       : IN Integer;
		     CONSTANT augend       : IN bit_vector
		   ) RETURN bit_vector;

     -------------------------------------------------------------------------------
     --     Function Name : Overloaded "-" operator
     -- 1.3.11    
     --     Purpose       : Subtraction operator for logic vectors.
     --     
     --     Parameters    :     result         left       right
     --                       std_logic_vector    std_logic_vector  std_logic_vector
     --     
     --     NOTE          : The subtraction operation is performed assuming all
     --                     operands and results are signed Two's complement integers.
     --
     --                     The operands may be of different length. The length of
     --                     the result equals the length of the longer operand.
     --     
     --                     Any underflow condition is ignored.
     --     Use           : 
     --                      VARIABLE a,b,c : std_logic_vector ( 7 downto 0 );
     --                      c := a - b;
     --                      c := a - "0101";  -- c = a - 5;
     --                      c := a - "101";   -- c = a - (-3)
     --     
     --     See Also      : RegAdd, RegSub, RegInc, RegDec, RegNegate
     -------------------------------------------------------------------------------
     FUNCTION  "-" ( CONSTANT minuend      : IN std_logic_vector;
		     CONSTANT subtrahend   : IN std_logic_vector
		   ) RETURN std_logic_vector;
     -------------------------------------------------------------------------------
     --     Function Name : Overloaded "-" operator
     -- 1.3.12
     --     Purpose       : Subtraction operator for logic vectors.
     --
     --     Parameters    :     result         left       right
     --                       std_logic_vector    INTEGER  std_logic_vector
     --
     --     NOTE          : The subtraction operation is performed assuming all
     --                     operands and results are signed Two's complement integers.
     --
     --                     The minuend is converted to std_logic_vector of length
     --                     equal to the subtrahend. The length of the result
     --                     equals the length of the subtrahend.
     --
     --                     Any overflow condition is ignored.
     --     Use           :
     --                      VARIABLE a: Integer;
     --                      VARIABLE b,c : std_logic_vector ( 7 downto 0 );
     --                      c := a - b;
     --                      c := 5 - b;
     --
     --     See Also      : RegAdd, RegSub, RegInc, RegDec, RegNegate
     -------------------------------------------------------------------------------
     FUNCTION  "-" ( CONSTANT minuend      : IN Integer;
		     CONSTANT subtrahend   : IN std_logic_vector
		   ) RETURN std_logic_vector;
     -------------------------------------------------------------------------------
     --     Function Name : Overloaded "-" operator
     -- 1.3.13
     --     Purpose       : Subtraction operator for logic vectors.
     --
     --     Parameters    :     result         left       right
     --                       std_logic_vector    std_logic_vector  Integer
     --
     --     NOTE          : The subtraction operation is performed assuming all
     --                     operands and results are signed Two's complement integers.
     --
     --                     The subtrahend is converted to std_logic_vector of length
     --                     equal to the minuend. The length of the result
     --                     equals the length of the minuend.
     --
     --                     Any overflow condition is ignored.
     --     Use           :
     --                      VARIABLE a,c : std_logic_vector ( 7 downto 0 );
     --                      VARIABLE b: Integer;
     --                      c := a - b;
     --                      c := a - 5;
     --
     --     See Also      : RegAdd, RegSub, RegInc, RegDec, RegNegate
     -------------------------------------------------------------------------------
     FUNCTION  "-" ( CONSTANT minuend      : IN std_logic_vector;
		     CONSTANT subtrahend   : IN Integer
		   ) RETURN std_logic_vector;
     -------------------------------------------------------------------------------
     --     Function Name : Overloaded "-" operator
     --     
     --     Purpose       : Subtraction operator for ulogic vectors.
     --     
     --     Parameters    :     result         left                right
     --                    std_ulogic_vector  std_ulogic_vector  std_ulogic_vector
     --     
     --     NOTE          : The subtraction operation is performed assuming all
     --                     operands and results are signed Two's complement integers.
     --
     --                     The operands may be of different length. The length of
     --                     the result equals the length of the longer operand.
     --     
     --                     Any underflow condition is ignored.
     --     Use           : 
     --                      VARIABLE a,b,c : std_ulogic_vector ( 7 downto 0 );
     --                      c := a - b;
     --                      c := a - "0101";  -- c = a - 5;
     --                      c := a - "101";   -- c = a - (-3)
     --     
     --     See Also      : RegAdd, RegSub, RegInc, RegDec, RegNegate
     -------------------------------------------------------------------------------
     FUNCTION  "-" ( CONSTANT minuend      : IN std_ulogic_vector;
		     CONSTANT subtrahend   : IN std_ulogic_vector
		   ) RETURN std_ulogic_vector;
     -------------------------------------------------------------------------------
     --     Function Name : Overloaded "-" operator
     -- 1.3.12
     --     Purpose       : Subtraction operator for ulogic vectors.
     --
     --     Parameters    :     result         left       right
     --                    std_ulogic_vector  INTEGER  std_ulogic_vector
     --
     --     NOTE          : The subtraction operation is performed assuming all
     --                     operands and results are signed Two's complement integers.
     --
     --                     The minuend is converted to std_ulogic_vector of length
     --                     equal to the subtrahend. The length of the result
     --                     equals the length of the subtrahend.
     --
     --                     Any overflow condition is ignored.
     --     Use           :
     --                      VARIABLE a: Integer;
     --                      VARIABLE b,c : std_logic_vector ( 7 downto 0 );
     --                      c := a - b;
     --                      c := 5 - b;
     --
     --     See Also      : RegAdd, RegSub, RegInc, RegDec, RegNegate
     -------------------------------------------------------------------------------
     FUNCTION  "-" ( CONSTANT minuend      : IN Integer;
		     CONSTANT subtrahend   : IN std_ulogic_vector
		   ) RETURN std_ulogic_vector;
     -------------------------------------------------------------------------------
     --     Function Name : Overloaded "-" operator
     -- 1.3.13
     --     Purpose       : Subtraction operator for ulogic vectors.
     --
     --     Parameters    :     result         left              right
     --                     std_ulogic_vector std_ulogic_vector  Integer
     --
     --     NOTE          : The subtraction operation is performed assuming all
     --                     operands and results are signed Two's complement integers.
     --
     --                     The subtrahend is converted to std_ulogic_vector of length
     --                     equal to the minuend. The length of the result
     --                     equals the length of the minuend.
     --
     --                     Any overflow condition is ignored.
     --     Use           :
     --                      VARIABLE a,c : std_ulogic_vector ( 7 downto 0 );
     --                      VARIABLE b: Integer;
     --                      c := a - b;
     --                      c := a - 5;
     --
     --     See Also      : RegAdd, RegSub, RegInc, RegDec, RegNegate
     -------------------------------------------------------------------------------
     FUNCTION  "-" ( CONSTANT minuend      : IN std_ulogic_vector;
		     CONSTANT subtrahend   : IN Integer
		   ) RETURN std_ulogic_vector;
     -------------------------------------------------------------------------------
     --     Function Name : Overloaded "-" operator
     -- 1.3.14 
     --     Purpose       : Subtraction operator for bit vectors.
     --
     --     Parameters    :     result         left       right
     --                       bit_vector    bit_vector  bit_vector
     --
     --     NOTE          : The subtraction operation is performed assuming all
     --                     operands and results are signed Two's complement integers.
     --
     --                     The operands may be of different length. The length of
     --                     the result equals the length of the longer operand.
     --
     --                     Any underflow condition is ignored.
     --     Use           :
     --                      VARIABLE a,b,c : bit_vector ( 7 downto 0 );
     --                      c := a - b;
     --                      c := a - B"0101";  -- c = a - 5;
     --                      c := a - B"101";   -- c = a - (-3)
     --
     --     See Also      : RegAdd, RegSub, RegInc, RegDec, RegNegate
     -------------------------------------------------------------------------------
     FUNCTION  "-" ( CONSTANT minuend      : IN bit_vector;
		     CONSTANT subtrahend   : IN bit_vector
		   ) RETURN bit_vector;
     -------------------------------------------------------------------------------
     --     Function Name : Overloaded "-" operator
     -- 1.3.15
     --     Purpose       : Subtraction operator for logic vectors.
     --
     --     Parameters    :     result         left       right
     --                       bit_vector    bit_vector  Integer
     --
     --     NOTE          : The subtraction operation is performed assuming all
     --                     operands and results are signed Two's complement integers.
     --
     --                     The subtrahend is converted to bit_vector of length
     --                     equal to the minuend. The length of the result
     --                     equals the length of the minuend.
     --
     --                     Any overflow condition is ignored.
     --     Use           :
     --                      VARIABLE a,c : bit_vector ( 7 downto 0 );
     --                      VARIABLE b: Integer;
     --                      c := a - b;
     --                      c := a - 5;
     --
     --     See Also      : RegAdd, RegSub, RegInc, RegDec, RegNegate
     -------------------------------------------------------------------------------
     FUNCTION  "-" ( CONSTANT minuend      : IN bit_vector;
		     CONSTANT subtrahend   : IN Integer
		   ) RETURN bit_vector;
     -------------------------------------------------------------------------------
     --     Function Name : Overloaded "-" operator
     -- 1.3.16
     --     Purpose       : Subtraction operator for bit vectors.
     --
     --     Parameters    :     result         left       right
     --                       bit_vector    INTEGER  bit_vector
     --
     --     NOTE          : The subtraction operation is performed assuming all
     --                     operands and results are signed Two's complement integers.
     --
     --                     The minuend is converted to bit_vector of length
     --                     equal to the subtrahend. The length of the result
     --                     equals the length of the subtrahend.
     --
     --                     Any overflow condition is ignored.
     --     Use           :
     --                      VARIABLE a: Integer;
     --                      VARIABLE b,c : bit_vector ( 7 downto 0 );
     --                      c := a - b;
     --                      c := 5 - b;
     --
     --     See Also      : RegAdd, RegSub, RegInc, RegDec, RegNegate
     -------------------------------------------------------------------------------
     FUNCTION  "-" ( CONSTANT minuend      : IN Integer;
		     CONSTANT subtrahend   : IN bit_vector
		   ) RETURN bit_vector;
     -------------------------------------------------------------------------------
     --     Function Name : Overloaded "-" operator
     -- 1.4.5
     --     Purpose       : Unary minus operator for bit vectors.
     --
     --     Parameters    :     result         v 
     --                       bit_vector    bit_vector 
     --
     --     NOTE          : The  minus  operation is performed assuming 
     --                     operand and result are signed Two's complement integers.
     --     Use           :
     --                      VARIABLE a,c : bit_vector ( 7 downto 0 );
     --                      c :=  - a;
     --
     --     See Also      :  RegNegate
     -------------------------------------------------------------------------------
     FUNCTION "-"  (CONSTANT subtrahend   : IN bit_vector
		   ) RETURN bit_vector;
     -------------------------------------------------------------------------------
     --     Function Name : Overloaded "-" operator
     -- 1.4.6
     --     Purpose       : Unary minus operator for logic vectors.
     --
     --     Parameters    :     result              operand 
     --                       std_logic_vector    std_logic_vector 
     --
     --     NOTE          : The  minus  operation is performed assuming 
     --                     operand and result are in signed Two's complement notation.
     --
     --     Use           :
     --                      VARIABLE a,c : std_logic_vector ( 7 downto 0 );
     --                      c :=  - a;
     --
     --     See Also      :  RegNegate
     -------------------------------------------------------------------------------
     FUNCTION "-"  (CONSTANT subtrahend   : IN std_logic_vector
		   ) RETURN std_logic_vector;
     -------------------------------------------------------------------------------
     --     Function Name : Overloaded "-" operator
     --
     --     Purpose       : Unary minus operator for ulogic vectors.
     --
     --     Parameters    :     result              operand 
     --                       std_ulogic_vector    std_ulogic_vector 
     --
     --     NOTE          : The  minus  operation is performed assuming 
     --                     operand and result are in signed Two's complement notation.
     --
     --     Use           :
     --                      VARIABLE a,c : std_ulogic_vector ( 7 downto 0 );
     --                      c :=  - a;
     --
     --     See Also      :  RegNegate
     -------------------------------------------------------------------------------
     FUNCTION "-"  (CONSTANT subtrahend   : IN std_ulogic_vector
		   ) RETURN std_ulogic_vector;
     -------------------------------------------------------------------------------
     --     Function Name : Overloaded "*" operator
     --    
     --     Purpose       : Multiplication operator for logic vectors.
     --     
     --     Parameters    :     result         left       right
     --                       std_logic_vector    std_logic_vector  std_logic_vector
     --     
     --     NOTE          : The multiplication operation is performed assuming all
     --                     operands and results are signed Two's complement integers.
     --
     --                     The operands may be of different length. The length of
     --                     the result equals the length of the longer operand.
     --     
     --                     A temporary result is computed of sufficient length
     --                     to avoid overflow. The high order bits of this temporary
     --                     vector are truncated to form the required length result.
     --                     No indication is given if the magnitude of the computed
     --                     result exceeds the size of the returned result vector.
     --     Use           : 
     --                      VARIABLE a,b,c : std_logic_vector ( 7 downto 0 );
     --                      c := a * b;
     --                      c := a * B"1101";  -- c = a * (-3)
     --     
     --     See Also      : RegMult, RegDiv
     -------------------------------------------------------------------------------
     FUNCTION  "*" ( CONSTANT multiplicand : IN std_logic_vector;
		     CONSTANT multiplier   : IN std_logic_vector
		   ) RETURN std_logic_vector;
     -------------------------------------------------------------------------------
     --     Function Name : Overloaded "*" operator
     -- 1.5.4
     --     Purpose       : Multiplication operator for logic vectors.
     --
     --     Parameters    :     result           left                right
     --                       std_logic_vector    std_logic_vector  Integer
     --
     --     NOTE          : The multiplication operation is performed assuming all
     --                     operands and results are signed Two's complement integers.
     --
     --                     The multiplier is converted to std_logic_vector of length
     --                     equal to the multiplicand. The length of the result
     --                     equals the length of the multiplicand.
     --
     --                     A temporary result is computed of sufficient length
     --                     to avoid overflow. The high order bits of this temporary
     --                     vector are truncated to form the required length result.
     --                     No indication is given if the magnitude of the computed
     --                     result exceeds the size of the returned result vector.
     --     Use           :
     --                      VARIABLE a,c : std_logic_vector ( 7 downto 0 );
     --                      VARIABLE b: Integer;
     --                      c := a * b;
     --                      c := a * 5; 
     --
     --     See Also      : RegMult, RegDiv
   -------------------------------------------------------------------------------
     FUNCTION  "*" ( CONSTANT multiplicand : IN std_logic_vector;
		     CONSTANT multiplier   : IN Integer
		   ) RETURN std_logic_vector;
     -------------------------------------------------------------------------------
     --     Function Name : Overloaded "*" operator
     -- 1.5.5
     --     Purpose       : Multiplication operator for logic vectors.
     --
     --     Parameters    :     result           left                right
     --                       std_logic_vector    Integer     std_logic_vector
     --
     --     NOTE          : The multiplication operation is performed assuming all
     --                     operands and results are signed Two's complement integers.
     --
     --                     The multiplicand is converted to std_logic_vector of length
     --                     equal to the multiplier. The length of the result
     --                     equals the length of the multiplier.
     --
     --                     A temporary result is computed of sufficient length
     --                     to avoid overflow. The high order bits of this temporary
     --                     vector are truncated to form the required length result.
     --                     No indication is given if the magnitude of the computed
     --                     result exceeds the size of the returned result vector.
     --     Use           :
     --                      VARIABLE a,c : std_logic_vector ( 7 downto 0 );
     --                      VARIABLE b: Integer;
     --                      c := a * b;
     --                      c := a * 5; 
     --
     --     See Also      : RegMult, RegDiv
     -------------------------------------------------------------------------------
     FUNCTION  "*" ( CONSTANT multiplicand : IN Integer;
		     CONSTANT multiplier   : IN std_logic_vector
		   ) RETURN std_logic_vector;
     -------------------------------------------------------------------------------
     --     Function Name : Overloaded "*" operator
     --    
     --     Purpose       : Multiplication operator for ulogic vectors.
     --     
     --     Parameters    :     result         left       right
     --                    std_ulogic_vector    std_ulogic_vector  std_ulogic_vector
     --     
     --     NOTE          : The multiplication operation is performed assuming all
     --                     operands and results are signed Two's complement integers.
     --
     --                     The operands may be of different length. The length of
     --                     the result equals the length of the longer operand.
     --     
     --                     A temporary result is computed of sufficient length
     --                     to avoid overflow. The high order bits of this temporary
     --                     vector are truncated to form the required length result.
     --                     No indication is given if the magnitude of the computed
     --                     result exceeds the size of the returned result vector.
     --     Use           : 
     --                      VARIABLE a,b,c : std_ulogic_vector ( 7 downto 0 );
     --                      c := a * b;
     --                      c := a * B"1101";  -- c = a * (-3)
     --     
     --     See Also      : RegMult, RegDiv
     -------------------------------------------------------------------------------
     FUNCTION  "*" ( CONSTANT multiplicand : IN std_ulogic_vector;
		     CONSTANT multiplier   : IN std_ulogic_vector
		   ) RETURN std_ulogic_vector;
     -------------------------------------------------------------------------------
     --     Function Name : Overloaded "*" operator
     -- 1.5.4
     --     Purpose       : Multiplication operator for logic vectors.
     --
     --     Parameters    :     result           left                right
     --                     std_ulogic_vector    std_ulogic_vector  Integer
     --
     --     NOTE          : The multiplication operation is performed assuming all
     --                     operands and results are signed Two's complement integers.
     --
     --                     The multiplier is converted to std_ulogic_vector of length
     --                     equal to the multiplicand. The length of the result
     --                     equals the length of the multiplicand.
     --
     --                     A temporary result is computed of sufficient length
     --                     to avoid overflow. The high order bits of this temporary
     --                     vector are truncated to form the required length result.
     --                     No indication is given if the magnitude of the computed
     --                     result exceeds the size of the returned result vector.
     --     Use           :
     --                      VARIABLE a,c : std_ulogic_vector ( 7 downto 0 );
     --                      VARIABLE b: Integer;
     --                      c := a * b;
     --                      c := a * 5; 
     --
     --     See Also      : RegMult, RegDiv
   -------------------------------------------------------------------------------
     FUNCTION  "*" ( CONSTANT multiplicand : IN std_ulogic_vector;
		     CONSTANT multiplier   : IN Integer
		   ) RETURN std_ulogic_vector;
     -------------------------------------------------------------------------------
     --     Function Name : Overloaded "*" operator
     -- 1.5.5
     --     Purpose       : Multiplication operator for logic vectors.
     --
     --     Parameters    :     result           left                right
     --                       std_ulogic_vector    Integer     std_ulogic_vector
     --
     --     NOTE          : The multiplication operation is performed assuming all
     --                     operands and results are signed Two's complement integers.
     --
     --                     The multiplicand is converted to std_ulogic_vector of 
     --                     length equal to the multiplier. The length of the 
     --                     result equals the length of the multiplier.
     --
     --                     A temporary result is computed of sufficient length
     --                     to avoid overflow. The high order bits of this temporary
     --                     vector are truncated to form the required length result.
     --                     No indication is given if the magnitude of the computed
     --                     result exceeds the size of the returned result vector.
     --     Use           :
     --                      VARIABLE a,c : std_ulogic_vector ( 7 downto 0 );
     --                      VARIABLE b: Integer;
     --                      c := a * b;
     --                      c := a * 5; 
     --
     --     See Also      : RegMult, RegDiv
     -------------------------------------------------------------------------------
     FUNCTION  "*" ( CONSTANT multiplicand : IN Integer;
		     CONSTANT multiplier   : IN std_ulogic_vector
		   ) RETURN std_ulogic_vector;
 --+-----------------------------------------------------------------------------
 --|     Function Name : Overloaded "*" operator
 --|
 --|     Purpose       : Multiplication operator for bit vectors.
 --|
 --|     Parameters    :     result         left       right
 --|                       BIT_VECTOR    BIT_VECTOR  BIT_VECTOR
 --|
 --|     NOTE          : The multiplication operation is performed assuming all
 --|                     operands and results are signed Two's complement integers.
 --|
 --|                     The operands may be of different length. The length of
 --|                     the result equals the length of the longer operand.
 --|
 --|                     A temporary result is computed of sufficient length
 --|                     to avoid overflow. The high order bits of this temporary
 --|                     vector are truncated to form the required length result.
 --|                     No indication is given if the magnitude of the computed
 --|                     result exceeds the size of the returned result vector.
 --|     Use           :
 --|                      VARIABLE a,b,c : bit_vector ( 7 downto 0 );
 --|                      c := a * b;
 --|                      c := a * B"1101";  -- c = a * (-3)
 --|
 --|     See Also      : RegMult, RegDiv
 --|-----------------------------------------------------------------------------
     FUNCTION  "*" ( CONSTANT multiplicand : IN BIT_VECTOR;
		     CONSTANT multiplier   : IN BIT_VECTOR
		   ) RETURN BIT_VECTOR;
 --+-----------------------------------------------------------------------------
 --|     Function Name : Overloaded "*" operator
 --| 1.5.7
 --|     Purpose       : Multiplication operator for bit vectors.
 --|
 --|     Parameters    :     result         left       right
 --|                       BIT_VECTOR    BIT_VECTOR  INTEGER
 --|
 --|     NOTE          : The multiplication operation is performed assuming all
 --|                     operands and results are signed Two's complement integers.
 --|
 --|                     The multiplier is converted to bit_vector of length
 --|                     equal to the multiplicand. The length of the result
 --|                     equals the length of the multiplicand.
 --|
 --|                     A temporary result is computed of sufficient length
 --|                     to avoid overflow. The high order bits of this temporary
 --|                     vector are truncated to form the required length result.
 --|                     No indication is given if the magnitude of the computed
 --|                     result exceeds the size of the returned result vector.
 --|     Use           :
 --|                      VARIABLE a,c : BIT_VECTOR ( 7 downto 0 );
 --|                      VARIABLE b: INTEGER;
 --|                      c := a * b;
 --|                      c := a * 5; 
 --|
 --|     See Also      : RegMult, RegDiv
 --|-----------------------------------------------------------------------------
     FUNCTION  "*" ( CONSTANT multiplicand : IN BIT_VECTOR;
		     CONSTANT multiplier   : IN INTEGER
		   ) RETURN BIT_VECTOR;
 --+-----------------------------------------------------------------------------
 --|     Function Name : Overloaded "*" operator
 --| 1.5.8
 --|     Purpose       : Multiplication operator for bit vectors.
 --|
 --|     Parameters    :     result         left       right
 --|                       BIT_VECTOR    INTEGER  BIT_VECTOR
 --|
 --|     NOTE          : The multiplication operation is performed assuming all
 --|                     operands and results are signed Two's complement integers.
 --|
 --|                     The multiplicand is converted to BIT_VECTOR of length
 --|                     equal to the multiplier. The length of the result
 --|                     equals the length of the multiplier.
 --|
 --|                     A temporary result is computed of sufficient length
 --|                     to avoid overflow. The high order bits of this temporary
 --|                     vector are truncated to form the required length result.
 --|                     No indication is given if the magnitude of the computed
 --|                     result exceeds the size of the returned result vector.
 --|     Use           :
 --|                      VARIABLE a : INTEGER;
 --|                      VARIABLE b,c : BIT_VECTOR ( 7 downto 0 );
 --|                      c := a * b;
 --|                      c := 5 * b; 
 --|
 --|     See Also      : RegMult, RegDiv
 --|-----------------------------------------------------------------------------
    FUNCTION  "*" ( CONSTANT multiplicand : IN INTEGER; 
		    CONSTANT multiplier   : IN BIT_VECTOR
		   ) RETURN BIT_VECTOR;

     -------------------------------------------------------------------------------
     --     Function Name : Overloaded "/" operator
     --    
     --     Purpose       : Division operator for logic vectors.
     --     
     --     Parameters    :     result         left       right
     --                       std_logic_vector    std_logic_vector  std_logic_vector
     --     
     --     NOTE          : The division operation is performed assuming all
     --                     operands and results are signed Two's complement integers.
     --
     --                     The operands may be of different length. The length of
     --                     the result equals the length of dividend.
     --     
     --                     Any remainder is ignored - no rounding is applied.
     --
     --                     An ASSERTION message of severity ERROR is issued
     --                     if division by 0 is attempted. In this case the
     --                     return value is 0 (all 0's).
     --     Use           : 
     --                      VARIABLE a,b,c : std_logic_vector ( 7 downto 0 );
     --                      c := a / b;
     --                      c := a / B"1101";  -- c = a / (-3)
     --     Se Also       : RegMult, RegDiv
     ----------------------------------------------------------------------------------
     FUNCTION  "/" ( CONSTANT dividend     : IN std_logic_vector;
		     CONSTANT divisor      : IN std_logic_vector
		   ) RETURN std_logic_vector;
     -------------------------------------------------------------------------------
     --     Function Name : Overloaded "/" operator
     -- 1.5.12
     --     Purpose       : Division operator for logic vectors.
     --
     --     Parameters    :     result         left       right
     --                       std_logic_vector    std_logic_vector  INTEGER
     --
     --     NOTE          : The division operation is performed assuming all
     --                     operands and results are signed Two's complement integers.
     --
     --                     The divisor is converted to std_logic_vector of length
     --                     equal to the dividend. The length of the result
     --                     equals the length of the dividend.
     --
     --                     Any remainder is ignored - no rounding is applied.
     --
     --                     An ASSERTION message of severity ERROR is issued
     --                     if division by 0 is attempted. In this case the
     --                     return value is 0 (all 0's).
     --     Use           :
     --                      VARIABLE a,c : std_logic_vector ( 7 downto 0 );
     --                      VARIABLE b : INTEGER;
     --                      c := a / b;
     --                      c := a / 5; 
     --     Se Also       : RegMult, RegDiv
     --------------------------------------------------------------------------------
     FUNCTION  "/" ( CONSTANT dividend     : IN std_logic_vector;
		     CONSTANT divisor      : IN INTEGER
		   ) RETURN std_logic_vector;
     -------------------------------------------------------------------------------
     --     Function Name : Overloaded "/" operator
     -- 1.5.13
     --     Purpose       : Division operator for logic vectors.
     --
     --     Parameters    :     result         left       right
     --                       std_logic_vector    INTEGER  std_logic_vector
     --
     --     NOTE          : The division operation is performed assuming all
     --                     operands and results are signed Two's complement integers.
     --
     --                     The dividend is converted to std_logic_vector of length
     --                     equal to the divisor. The length of the result
     --                     equals the length of the divisor.
     --
     --                     Any remainder is ignored - no rounding is applied.
     --
     --                     An ASSERTION message of severity ERROR is issued
     --                     if division by 0 is attempted. In this case the
     --                     return value is 0 (all 0's).
     --     Use           :
     --                      VARIABLE a : INTEGER;
     --                      VARIABLE b,c : std_logic_vector ( 7 downto 0 );
     --                      c := a / b;
     --                      c := 5 / b;
     --     Se Also       : RegMult, RegDiv
     --------------------------------------------------------------------------------
     FUNCTION  "/" ( CONSTANT dividend     : IN INTEGER;
		     CONSTANT divisor      : IN std_logic_vector
		   ) RETURN std_logic_vector;
     -------------------------------------------------------------------------------
     --     Function Name : Overloaded "/" operator
     --    
     --     Purpose       : Division operator for ulogic vectors.
     --     
     --     Parameters    :     result         left       right
     --                       std_ulogic_vector    std_ulogic_vector  std_ulogic_vector
     --     
     --     NOTE          : The division operation is performed assuming all
     --                     operands and results are signed Two's complement integers.
     --
     --                     The operands may be of different length. The length of
     --                     the result equals the length of the dividend.
     --     
     --                     Any remainder is ignored - no rounding is applied.
     --
     --                     An ASSERTION message of severity ERROR is issued
     --                     if division by 0 is attempted. In this case the
     --                     return value is 0 (all 0's).
     --     Use           : 
     --                      VARIABLE a,b,c : std_ulogic_vector ( 7 downto 0 );
     --                      c := a / b;
     --                      c := a / B"1101";  -- c = a / (-3)
     --     Se Also       : RegMult, RegDiv
     ---------------------------------------------------------------------------------
     FUNCTION  "/" ( CONSTANT dividend     : IN std_ulogic_vector;
		     CONSTANT divisor      : IN std_ulogic_vector
		   ) RETURN std_ulogic_vector;
     -------------------------------------------------------------------------------
     --     Function Name : Overloaded "/" operator
     -- 1.5.12
     --     Purpose       : Division operator for logic vectors.
     --
     --     Parameters    :     result         left       right
     --                       std_ulogic_vector    std_ulogic_vector  INTEGER
     --
     --     NOTE          : The division operation is performed assuming all
     --                     operands and results are signed Two's complement integers.
     --
     --                     The divisor is converted to std_ulogic_vector of length
     --                     equal to the dividend. The length of the result
     --                     equals the length of the dividend.
     --
     --                     Any remainder is ignored - no rounding is applied.
     --
     --                     An ASSERTION message of severity ERROR is issued
     --                     if division by 0 is attempted. In this case the
     --                     return value is 0 (all 0's).
     --     Use           :
     --                      VARIABLE a,c : std_ulogic_vector ( 7 downto 0 );
     --                      VARIABLE b : INTEGER;
     --                      c := a / b;
     --                      c := a / 5; 
     --     Se Also       : RegMult, RegDiv
   --------------------------------------------------------------------------------
     FUNCTION  "/" ( CONSTANT dividend     : IN std_ulogic_vector;
		     CONSTANT divisor      : IN INTEGER
		   ) RETURN std_ulogic_vector;
     -------------------------------------------------------------------------------
     --     Function Name : Overloaded "/" operator
     -- 1.5.13
     --     Purpose       : Division operator for logic vectors.
     --
     --     Parameters    :     result         left       right
     --                       std_ulogic_vector    INTEGER  std_ulogic_vector
     --
     --     NOTE          : The division operation is performed assuming all
     --                     operands and results are signed Two's complement integers.
     --
     --                     The dividend is converted to std_ulogic_vector of length
     --                     equal to the divisor. The length of the result
     --                     equals the length of the divisor.
     --
     --                     Any remainder is ignored - no rounding is applied.
     --
     --                     An ASSERTION message of severity ERROR is issued
     --                     if division by 0 is attempted. In this case the
     --                     return value is 0 (all 0's).
     --     Use           :
     --                      VARIABLE a : INTEGER;
     --                      VARIABLE b,c : std_ulogic_vector ( 7 downto 0 );
     --                      c := a / b;
     --                      c := 5 / b;
     --     Se Also       : RegMult, RegDiv
     --------------------------------------------------------------------------------
     FUNCTION  "/" ( CONSTANT dividend     : IN INTEGER;
		     CONSTANT divisor      : IN std_ulogic_vector
		   ) RETURN std_ulogic_vector;
 --+-----------------------------------------------------------------------------
 --|     Function Name : Overloaded "/" operator
 --| 1.5.14
 --|     Purpose       : Division operator for bit vectors.  
 --|     Parameters    :     result         left       right
 --|                       BIT_VECTOR    BIT_VECTOR  BIT_VECTOR
 --|
 --|     NOTE          : The division operation is performed assuming all
 --|                     operands and results are signed Two's complement integers.
 --|
 --|                     The operands may be of different length. The length of
 --|                     the result equals the length of the dividend.
 --|
 --|                     Any remainder is ignored - no rounding is applied.
 --|
 --|                     An ASSERTION message of severity ERROR is issued
 --|                     if division by 0 is attempted. In this case the
 --|                     return value is 0 (all 0's).
 --|     Use           :
 --|                      VARIABLE a,b,c : bit_vector ( 7 downto 0 );
 --|                      c := a / b;
 --|                      c := a / B"1101";  -- c = a / (-3)
 --|
 --|     See Also      : RegMult, RegDiv
 --|-----------------------------------------------------------------------------
     FUNCTION  "/" ( CONSTANT dividend     : IN BIT_VECTOR;
		     CONSTANT divisor      : IN BIT_VECTOR
		   ) RETURN BIT_VECTOR;
 --+-----------------------------------------------------------------------------
 --|     Function Name : Overloaded "/" operator
 --| 1.5.15
 --|     Purpose       : Division operator for bit vectors.
 --|     Parameters    :     result         left       right
 --|                       BIT_VECTOR    BIT_VECTOR  INTEGER
 --|
 --|     NOTE          : The division operation is performed assuming all
 --|                     operands and results are signed Two's complement integers.
 --|
 --|                     The divisor is converted to bit_vector of length
 --|                     equal to the dividend. The length of the result
 --|                     equals the length of the dividend.
 --|
 --|                     Any remainder is ignored - no rounding is applied.
 --|
 --|                     An ASSERTION message of severity ERROR is issued
 --|                     if division by 0 is attempted. In this case the
 --|                     return value is 0 (all 0's).
 --|     Use           :
 --|                      VARIABLE a,c : BIT_VECTOR ( 7 downto 0 );
 --|                      VARIABLE b : INTEGER;
 --|                      c := a / b;
 --|                      c := a / 5;
 --| 
 --|     See Also      : RegMult, RegDiv
 --|-----------------------------------------------------------------------------
     FUNCTION  "/" ( CONSTANT dividend     : IN BIT_VECTOR;
		     CONSTANT divisor      : IN INTEGER
		   ) RETURN BIT_VECTOR;
 --+-----------------------------------------------------------------------------
 --|     Function Name : Overloaded "/" operator
 --| 1.5.16
 --|     Purpose       : Division operator for bit vectors.
 --|     Parameters    :     result         left       right
 --|                       BIT_VECTOR    INTEGER  BIT_VECTOR
 --|
 --|     NOTE          : The division operation is performed assuming all
 --|                     operands and results are signed Two's complement integers.
 --|
 --|                     The dividend is converted to bit_vector of length
 --|                     equal to the divisor. The length of the result
 --|                     equals the length of the divisor.
 --|
 --|                     Any remainder is ignored - no rounding is applied.
 --|
 --|                     An ASSERTION message of severity ERROR is issued
 --|                     if division by 0 is attempted. In this case the
 --|                     return value is 0 (all 0's).
 --|     Use           :
 --|                      VARIABLE a : INTEGER;
 --|                      VARIABLE b,c : BIT_VECTOR ( 7 downto 0 );
 --|                      c := a / b;
 --|                      c := 5 / b;
 --|
 --|     See Also      : RegMult, RegDiv
 --|-----------------------------------------------------------------------------
     FUNCTION  "/" ( CONSTANT dividend     : IN INTEGER;
		     CONSTANT divisor      : IN BIT_VECTOR
		   ) RETURN BIT_VECTOR;
     -------------------------------------------------------------------------------
     --     Function Name : Overloaded "mod" operator
     -- 1.5.19
     --     Purpose       : Modulus operator for logic vectors.
     --
     --     Parameters    :     result         left       right
     --                       std_logic_vector    std_logic_vector  std_logic_vector
     --
     --     NOTE          : The modulus operation is performed assuming all
     --                     operands and results are signed Two's complement integers.
     --
     --                     The operands may be of different length. The length of
     --                     the result equals the length of the modulus.
     --
     --                     An ASSERTION message of severity ERROR is issued
     --                     if division by 0 is attempted. In this case the
     --                     return value is 0 (all 0's).
     --     Use           :
     --                      VARIABLE a,b,c : std_logic_vector ( 7 downto 0 );
     --                      c := a mod b;
     --                      c := a mod B"1101";  -- c = a / (-3)
     --     Se Also       : RegRem, RegDiv
     -------------------------------------------------------------------------------
     FUNCTION  "mod" ( CONSTANT dividend     : IN std_logic_vector;
		       CONSTANT modulus      : IN std_logic_vector
		     ) RETURN std_logic_vector;
   -------------------------------------------------------------------------------
     --     Function Name : Overloaded "mod" operator
     -- 1.5.20
     --     Purpose       : Modulus operator for logic vectors.
     --
     --     Parameters    :     result         left       right
     --                       std_logic_vector    std_logic_vector  INTEGER
     --
     --     NOTE          : The modulus operation is performed assuming all
     --                     operands and results are signed Two's complement integers.
     --
     --                     The modulus is converted to std_logic_vector of length
     --                     equal to the dividend. The length of the result
     --                     equals the length of the dividend.
     --
     --                     An ASSERTION message of severity ERROR is issued
     --                     if division by 0 is attempted. In this case the
     --                     return value is 0 (all 0's).
     --     Use           :
     --                      VARIABLE a,c : std_logic_vector ( 7 downto 0 );
     --                      VARIABLE b : INTEGER;
     --                      c := a mod b;
     --                      c := a mod 5;
     --     Se Also       : RegRem, RegDiv
     -------------------------------------------------------------------------------
     FUNCTION  "mod" ( CONSTANT dividend     : IN std_logic_vector;
		       CONSTANT modulus      : IN INTEGER
		     ) RETURN std_logic_vector;
     -------------------------------------------------------------------------------
     --     Function Name : Overloaded "mod" operator
     -- 1.5.21
     --     Purpose       : Modulus operator for logic vectors.
     --
     --     Parameters    :     result         left       right
     --                       std_logic_vector    INTEGER  std_logic_vector
     --
     --     NOTE          : The modulus operation is performed assuming all
     --                     operands and results are signed Two's complement integers.
     --
     --                     The dividend is converted to std_logic_vector of length
     --                     equal to the modulus. The length of the result
     --                     equals the length of the modulus.
     --
     --                     An ASSERTION message of severity ERROR is issued
     --                     if division by 0 is attempted. In this case the
     --                     return value is 0 (all 0's).
     --     Use           :
     --                      VARIABLE a : INTEGER;
     --                      VARIABLE b,c : std_logic_vector ( 7 downto 0 );
     --                      c := a mod b;
     --                      c := 5 mod b;
     --     Se Also       : RegRem, RegDiv
     --------------------------------------------------------------------------------
     FUNCTION  "mod" ( CONSTANT dividend     : IN INTEGER;
		       CONSTANT modulus      : IN std_logic_vector
		     ) RETURN std_logic_vector;
     -------------------------------------------------------------------------------
     --     Function Name : Overloaded "mod" operator
     -- 
     --     Purpose       : Modulus operator for ulogic vectors.
     --
     --     Parameters    :     result         left       right
     --                       std_ulogic_vector    std_ulogic_vector  std_ulogic_vector
     --
     --     NOTE          : The modulus operation is performed assuming all
     --                     operands and results are signed Two's complement integers.
     --
     --                     The operands may be of different length. The length of
     --                     the result equals the length of the modulus.
     --
     --                     An ASSERTION message of severity ERROR is issued
     --                     if division by 0 is attempted. In this case the
     --                     return value is 0 (all 0's).
     --     Use           :
     --                      VARIABLE a,b,c : std_ulogic_vector ( 7 downto 0 );
     --                      c := a mod b;
     --                      c := a mod B"1101";  -- c = a / (-3)
     --     Se Also       : RegRem, RegDiv
     --------------------------------------------------------------------------------
     FUNCTION  "mod" ( CONSTANT dividend     : IN std_ulogic_vector;
		       CONSTANT modulus      : IN std_ulogic_vector
		     ) RETURN std_ulogic_vector;
     -------------------------------------------------------------------------------
     --     Function Name : Overloaded "mod" operator
     -- 
     --     Purpose       : Modulus operator for ulogic vectors.
     --
     --     Parameters    :     result         left       right
     --                       std_ulogic_vector    std_ulogic_vector  INTEGER
     --
     --     NOTE          : The modulus operation is performed assuming all
     --                     operands and results are signed Two's complement integers.
     --
     --                     The modulus is converted to std_ulogic_vector of length
     --                     equal to the dividend. The length of the result
     --                     equals the length of the dividend.
     --
     --                     An ASSERTION message of severity ERROR is issued
     --                     if division by 0 is attempted. In this case the
     --                     return value is 0 (all 0's).
     --     Use           :
     --                      VARIABLE a,c : std_ulogic_vector ( 7 downto 0 );
     --                      VARIABLE b : INTEGER;
     --                      c := a mod b;
     --                      c := a mod 5;
     --     Se Also       : RegRem, RegDiv
     --------------------------------------------------------------------------------
     FUNCTION  "mod" ( CONSTANT dividend     : IN std_ulogic_vector;
		       CONSTANT modulus      : IN INTEGER
		     ) RETURN std_ulogic_vector;
     -------------------------------------------------------------------------------
     --     Function Name : Overloaded "mod" operator
     -- 1.5.21
     --     Purpose       : Modulus operator for ulogic vectors.
     --
     --     Parameters    :     result         left       right
     --                       std_ulogic_vector    INTEGER  std_ulogic_vector
     --
     --     NOTE          : The modulus operation is performed assuming all
     --                     operands and results are signed Two's complement integers.
     --
     --                     The dividend is converted to std_ulogic_vector of length
     --                     equal to the modulus. The length of the result
     --                     equals the length of the modulus.
     --
     --                     An ASSERTION message of severity ERROR is issued
     --                     if division by 0 is attempted. In this case the
     --                     return value is 0 (all 0's).
     --     Use           :
     --                      VARIABLE a : INTEGER;
     --                      VARIABLE b,c : std_ulogic_vector ( 7 downto 0 );
     --                      c := a mod b;
     --                      c := 5 mod b;
     --     Se Also       : RegRem, RegDiv
     --------------------------------------------------------------------------------
     FUNCTION  "mod" ( CONSTANT dividend     : IN INTEGER;
		       CONSTANT modulus      : IN std_ulogic_vector
		     ) RETURN std_ulogic_vector;
     -------------------------------------------------------------------------------
     --     Function Name : Overloaded "mod" operator
     -- 1.5.22
     --     Purpose       : Modulus operator for bit vectors.
     --
     --     Parameters    :     result         left       right
     --                       bit_vector    bit_vector  bit_vector
     --
     --     NOTE          : The modulus operation is performed assuming all
     --                     operands and results are signed Two's complement integers.
     --
     --                     The operands may be of different length. The length of
     --                     the result equals the length of the modulus.
     --
     --                     An ASSERTION message of severity ERROR is issued
     --                     if division by 0 is attempted. In this case the
     --                     return value is 0 (all 0's).
     --     Use           :
     --                      VARIABLE a,b,c : bit_vector ( 7 downto 0 );
     --                      c := a mod b;
     --                      c := a mod B"1101";  -- c = a / (-3)
     --     Se Also       : RegRem, RegDiv
     ---------------------------------------------------------------------------------
     FUNCTION  "mod" ( CONSTANT dividend     : IN bit_vector;
		       CONSTANT modulus      : IN bit_vector
		     ) RETURN bit_vector;
     -------------------------------------------------------------------------------
     --     Function Name : Overloaded "mod" operator
     -- 1.5.23
     --     Purpose       : Modulus operator for bit vectors.
     --
     --     Parameters    :     result         left       right
     --                       bit_vector     bit_vector  INTEGER
     --
     --     NOTE          : The modulus operation is performed assuming all
     --                     operands and results are signed Two's complement integers.
     --
     --                     The modulus is converted to bit_vector of length
     --                     equal to the dividend. The length of the result
     --                     equals the length of the dividend.
     --
     --                     An ASSERTION message of severity ERROR is issued
     --                     if division by 0 is attempted. In this case the
     --                     return value is 0 (all 0's).
     --     Use           :
     --                      VARIABLE a,c : bit_vector ( 7 downto 0 );
     --                      VARIABLE b : INTEGER;
     --                      c := a mod b;
     --                      c := a mod 5;
     --     Se Also       : RegRem, RegDiv
     --------------------------------------------------------------------------------
     FUNCTION  "mod" ( CONSTANT dividend     : IN bit_vector;
		       CONSTANT modulus      : IN INTEGER
		     ) RETURN bit_vector;
     -------------------------------------------------------------------------------
     --     Function Name : Overloaded "mod" operator
     -- 1.5.24
     --     Purpose       : Modulus operator for bit vectors.
     --
     --     Parameters    :     result         left       right
     --                       bit_vector    INTEGER  bit_vector
     --
     --     NOTE          : The modulus operation is performed assuming all
     --                     operands and results are signed Two's complement integers.
     --
     --                     The dividend is converted to bit_vector of length
     --                     equal to the modulus. The length of the result
     --                     equals the length of the modulus.
     --
     --                     An ASSERTION message of severity ERROR is issued
     --                     if division by 0 is attempted. In this case the
     --                     return value is 0 (all 0's).
     --     Use           :
     --                      VARIABLE a : INTEGER;
     --                      VARIABLE b,c : bit_vector ( 7 downto 0 );
     --                      c := a mod b;
     --                      c := 5 mod b;
     --     Se Also       : RegRem, RegDiv
     --------------------------------------------------------------------------------
     FUNCTION  "mod" ( CONSTANT dividend     : IN INTEGER;
		       CONSTANT modulus      : IN bit_vector
		     ) RETURN bit_vector;
     --------------------------------------------------------------------------------
     --     Function Name : Overloaded "rem" operator
     -- 1.5.27
     --     Purpose       : Remainder operator for logic vectors.
     --
     --     Parameters    :     result         left             right
     --                     std_logic_vector  std_logic_vector  std_logic_vector
     --
     --     NOTE          : The division operation is performed assuming all
     --                     operands and results are signed Two's complement integers.
     --
     --                     The operands may be of different length. The length of
     --                     the result equals the length of the dividend.
     --
     --                     An ASSERTION message of severity ERROR is issued
     --                     if division by 0 is attempted. In this case the
     --                     return value is 0 (all 0's).
     --     Use           :
     --                      VARIABLE a,b,c : std_logic_vector ( 7 downto 0 );
     --                      c := a rem b;
     --                      c := a rem B"1101";  -- c = a rem (-3)
     ---------------------------------------------------------------------------------
     FUNCTION  "rem" ( CONSTANT dividend     : IN std_logic_vector;
		       CONSTANT divisor      : IN std_logic_vector
		     ) RETURN std_logic_vector;
     ---------------------------------------------------------------------------------
     --     Function Name : Overloaded "rem" operator
     -- 1.5.28
     --     Purpose       : Remainder operator for logic vectors.
     --
     --     Parameters    :     result         left       right
     --                       std_logic_vector    std_logic_vector  INTEGER
     --
     --     NOTE          : The division operation is performed assuming all
     --                     operands and results are signed Two's complement integers.
     --
     --                     The divisor is converted to std_logic_vector of length
     --                     equal to the dividend. The length of the result
     --                     equals the length of the dividend.
     --
     --                     An ASSERTION message of severity ERROR is issued
     --                     if division by 0 is attempted. In this case the
     --                     return value is 0 (all 0's).
     --     Use           :
     --                      VARIABLE a,c : std_logic_vector ( 7 downto 0 );
     --                      VARIABLE b : INTEGER;
     --                      c := a rem b;
     --                      c := a rem 5;
     --     Se Also       : RegMod, RegDiv
     --------------------------------------------------------------------------------
     FUNCTION  "rem" ( CONSTANT dividend     : IN std_logic_vector;
		       CONSTANT divisor      : IN INTEGER
		     ) RETURN std_logic_vector;
     -------------------------------------------------------------------------------
     --     Function Name : Overloaded "rem" operator
     -- 1.5.29
     --     Purpose       : Remainder operator for logic vectors.
     --
     --     Parameters    :     result         left       right
     --                       std_logic_vector    INTEGER  std_logic_vector
     --
     --     NOTE          : The division operation is performed assuming all
     --                     operands and results are signed Two's complement integers.
     --
     --                     The dividend is converted to std_logic_vector of length
     --                     equal to the divisor. The length of the result
     --                     equals the length of the divisor.
     --
     --                     An ASSERTION message of severity ERROR is issued
     --                     if division by 0 is attempted. In this case the
     --                     return value is 0 (all 0's).
     --     Use           :
     --                      VARIABLE a : INTEGER;
     --                      VARIABLE b,c : std_logic_vector ( 7 downto 0 );
     --                      c := a rem b;
     --                      c := 5 rem b;
     --     Se Also       : RegMod, RegDiv
     ------------------------------------------------------------------------------
     FUNCTION  "rem" ( CONSTANT dividend     : IN INTEGER;
		       CONSTANT divisor      : IN std_logic_vector
		     ) RETURN std_logic_vector;
     -------------------------------------------------------------------------------
     --     Function Name : Overloaded "rem" operator
     -- 
     --     Purpose       : Remainder operator for ulogic vectors.
     --
     --     Parameters    :     result         left             right
     --                     std_ulogic_vector  std_ulogic_vector  std_ulogic_vector
     --
     --     NOTE          : The division operation is performed assuming all
     --                     operands and results are signed Two's complement integers.
     --
     --                     The operands may be of different length. The length of
     --                     the result equals the length of the dividend.
     --
     --                     An ASSERTION message of severity ERROR is issued
     --                     if division by 0 is attempted. In this case the
     --                     return value is 0 (all 0's).
     --     Use           :
     --                      VARIABLE a,b,c : std_ulogic_vector ( 7 downto 0 );
     --                      c := a rem b;
     --                      c := a rem B"1101";  -- c = a rem (-3)
     ---------------------------------------------------------------------------------
     FUNCTION  "rem" ( CONSTANT dividend     : IN std_ulogic_vector;
		       CONSTANT divisor      : IN std_ulogic_vector
		     ) RETURN std_ulogic_vector;
     -------------------------------------------------------------------------------
     --     Function Name : Overloaded "rem" operator
     -- 
     --     Purpose       : Remainder operator for ulogic vectors.
     --
     --     Parameters    :     result         left       right
     --                       std_ulogic_vector    std_ulogic_vector  INTEGER
     --
     --     NOTE          : The division operation is performed assuming all
     --                     operands and results are signed Two's complement integers.
     --
     --                     The divisor is converted to std_ulogic_vector of length
     --                     equal to the dividend. The length of the result
     --                     equals the length of the dividend.
     --
     --                     An ASSERTION message of severity ERROR is issued
     --                     if division by 0 is attempted. In this case the
     --                     return value is 0 (all 0's).
     --     Use           :
     --                      VARIABLE a,c : std_ulogic_vector ( 7 downto 0 );
     --                      VARIABLE b : INTEGER;
     --                      c := a rem b;
     --                      c := a rem 5;
     --     Se Also       : RegMod, RegDiv
     -------------------------------------------------------------------------------
     FUNCTION  "rem" ( CONSTANT dividend     : IN std_ulogic_vector;
		       CONSTANT divisor      : IN INTEGER
		     ) RETURN std_ulogic_vector;
     -------------------------------------------------------------------------------
     --     Function Name : Overloaded "rem" operator
     -- 1.5.29
     --     Purpose       : Remainder operator for ulogic vectors.
     --
     --     Parameters    :     result         left       right
     --                       std_ulogic_vector    INTEGER  std_ulogic_vector
     --
     --     NOTE          : The division operation is performed assuming all
     --                     operands and results are signed Two's complement integers.
     --
     --                     The dividend is converted to std_ulogic_vector of length
     --                     equal to the divisor. The length of the result
     --                     equals the length of the divisor.
     --
     --                     An ASSERTION message of severity ERROR is issued
     --                     if division by 0 is attempted. In this case the
     --                     return value is 0 (all 0's).
     --     Use           :
     --                      VARIABLE a : INTEGER;
     --                      VARIABLE b,c : std_ulogic_vector ( 7 downto 0 );
     --                      c := a rem b;
     --                      c := 5 rem b;
     --     Se Also       : RegMod, RegDiv
     --------------------------------------------------------------------------------
     FUNCTION  "rem" ( CONSTANT dividend     : IN INTEGER;
		       CONSTANT divisor      : IN std_ulogic_vector
		     ) RETURN std_ulogic_vector;
 --+--------------------------------------------------------------------------------
 --|     Function Name : Overloaded "rem" operator
 --| 1.5.30
 --|     Purpose       : Remainder operator for bit vectors.
 --|     Parameters    :     result         left       right
 --|                       BIT_VECTOR    BIT_VECTOR  BIT_VECTOR
 --|
 --|     NOTE          : The division operation is performed assuming all
 --|                     operands and results are signed Two's complement integers.
 --|
 --|                     The operands may be of different length. The length of
 --|                     the result equals the length of the longer operand.
 --|
 --|                     An ASSERTION message of severity ERROR is issued
 --|                     if division by 0 is attempted. In this case the
 --|                     return value is 0 (all 0's).
 --|     Use           :
 --|                      VARIABLE a,b,c : bit_vector ( 7 downto 0 );
 --|                      c := a rem b;
 --|                      c := a rem B"1101";  -- c = a rem (-3)
 --|
 --|     See Also      : RegMod, RegDiv
 --|-----------------------------------------------------------------------------
     FUNCTION  "rem" ( CONSTANT dividend     : IN BIT_VECTOR;
		       CONSTANT divisor      : IN BIT_VECTOR
		     ) RETURN BIT_VECTOR;
 --+-----------------------------------------------------------------------------
 --|     Function Name : Overloaded "rem" operator
 --| 1.5.31
 --|     Purpose       : Remainder operator for bit vectors.
 --|     Parameters    :     result         left       right
 --|                       BIT_VECTOR    BIT_VECTOR  INTEGER
 --|
 --|     NOTE          : The division operation is performed assuming all
 --|                     operands and results are signed Two's complement integers.
 --|
 --|                     The divisor is converted to bit_vector of length
 --|                     equal to the dividend. The length of the result
 --|                     equals the length of the dividend.
 --|
 --|                     An ASSERTION message of severity ERROR is issued
 --|                     if division by 0 is attempted. In this case the
 --|                     return value is 0 (all 0's).
 --|     Use           :
 --|                      VARIABLE a,c : BIT_VECTOR ( 7 downto 0 );
 --|                      VARIABLE b : INTEGER;
 --|                      c := a rem b;
 --|                      c := a rem 5;
 --|
 --|     See Also      : RegMod, RegDiv
 --|-----------------------------------------------------------------------------
     FUNCTION  "rem" ( CONSTANT dividend     : IN BIT_VECTOR;
		       CONSTANT divisor      : IN INTEGER
		     ) RETURN BIT_VECTOR;
 --+-----------------------------------------------------------------------------
 --|     Function Name : Overloaded "rem" operator
 --| 1.5.32
 --|     Purpose       : Remainder operator for bit vectors.
 --|     Parameters    :     result         left       right
 --|                       BIT_VECTOR    INTEGER  BIT_VECTOR
 --|
 --|     NOTE          : The division operation is performed assuming all
 --|                     operands and results are signed Two's complement integers.
 --|
 --|                     The dividend is converted to bit_vector of length
 --|                     equal to the divisor. The length of the result
 --|                     equals the length of the divisor.
 --|
 --|                     An ASSERTION message of severity ERROR is issued
 --|                     if division by 0 is attempted. In this case the
 --|                     return value is 0 (all 0's).
 --|     Use           :
 --|                      VARIABLE a : INTEGER;
 --|                      VARIABLE b,c : BIT_VECTOR ( 7 downto 0 );
 --|                      c := a rem b;
 --|                      c := 5 rem b;
 --|
 --|     See Also      : RegMod, RegDiv
 --|-----------------------------------------------------------------------------
     FUNCTION  "rem" ( CONSTANT dividend     : IN INTEGER;
		       CONSTANT divisor      : IN BIT_VECTOR
		     ) RETURN BIT_VECTOR;
     -------------------------------------------------------------------------------
     --     Function Name : Overloaded "ABS" operator
     -- 1.6.11
     --     Purpose       : Absolute value operator for logic vectors.
     --
     --     Parameters    :     result             operand       
     --                       std_logic_vector    std_logic_vector
     --
     --     Use           :
     --                      VARIABLE a,c : std_logic_vector ( 7 downto 0 );
     --                      c := ABS(a);
     --
     --     See Also      : RegAbs
     -------------------------------------------------------------------------------
     FUNCTION  "ABS" ( CONSTANT operand : IN std_logic_vector
		     ) RETURN std_logic_vector;
     -------------------------------------------------------------------------------
     --     Function Name : Overloaded "ABS" operator
     -- 
     --     Purpose       : Absolute value operator for ulogic vectors.
     --
     --     Parameters    :     result             operand       
     --                       std_ulogic_vector    std_ulogic_vector
     --
     --     Use           :
     --                      VARIABLE a,c : std_ulogic_vector ( 7 downto 0 );
     --                      c := ABS(a);
     --
     --     See Also      : RegAbs
     -------------------------------------------------------------------------------
     FUNCTION  "ABS" ( CONSTANT operand : IN std_ulogic_vector
		     ) RETURN std_ulogic_vector;
     -------------------------------------------------------------------------------
     --     Function Name : Overloaded "ABS" operator
     -- 1.6.12
     --     Purpose       : Absolute value operator for bit vectors.
     --
     --     Parameters    :     result        operand       
     --                       bit_vector    bit_vector
     --
     --     Use           :
     --                      VARIABLE a,c : bit_vector ( 7 downto 0 );
     --                      c := ABS(a);
     --
     --     See Also      : RegAbs
     -------------------------------------------------------------------------------
     FUNCTION  "ABS" ( CONSTANT operand : IN bit_vector
		     ) RETURN bit_vector;

     -------------------------------------------------------------------------------
     --     Function Name : Overloaded "=" operator
     --   1.2.1 and 1.2.3  
     --     Purpose       : Equality relational operator for std_logic_vector : integer.
     --     
     --     Parameters    :     result         left              right
     --                        std_ulogic  std_logic_vector   std_logic_vector
     --                        BOOLEAN     INTEGER            std_logic_vector
     --                        BOOLEAN     std_logic_vector   INTEGER
     --                        std_ulogic  INTEGER            std_logic_vector
     --                        std_ulogic  std_logic_vector   INTEGER
     --                                     
     --     NOTE          : The std_logic_vector operands are assumed to be  
     --                     in  DefaultRegMode. If not they will be converted
     --                     to DefaultRegMode in the compare procedure. 
     --                     These vectors may be of any length.
     --     Use           : 
     --                      VARIABLE a : std_logic_vector ( 7 DOWNTO 0 ) := X"FF";
     --                      VARIABLE b : INTEGER;
     --                      IF ( a = b )  THEN 
     --     
     --     See Also      : RegEqual, RegNotEqual,
     -------------------------------------------------------------------------------
     FUNCTION  "=" ( CONSTANT l  : std_logic_vector;
		     CONSTANT r  : std_logic_vector
		   ) RETURN std_ulogic;
     -------------------------------------------------------------------------------
     FUNCTION  "=" ( CONSTANT l  : std_logic_vector;
		     CONSTANT r  : INTEGER
		   ) RETURN BOOLEAN;
     -- -----------------------------------------------------------------------------
     FUNCTION  "=" ( CONSTANT l  : INTEGER   ;
		     CONSTANT r  : std_logic_vector 
		   ) RETURN BOOLEAN;
     -------------------------------------------------------------------------------
     FUNCTION  "=" ( CONSTANT l  : std_logic_vector;
		     CONSTANT r  : INTEGER
		   ) RETURN std_ulogic;

     -- -----------------------------------------------------------------------------
     FUNCTION  "=" ( CONSTANT l  : INTEGER   ;
		     CONSTANT r  : std_logic_vector 
		   ) RETURN std_ulogic;
     -------------------------------------------------------------------------------
     --     Function Name : Overloaded "=" operator
     --   1.2.1 and 1.2.3  
     --     Purpose       : Equality relational operator for std_ulogic_vector : integer.
     --     
     --     Parameters    :     result         left              right
     --                        std_ulogic  std_ulogic_vector   std_ulogic_vector
     --                        BOOLEAN     INTEGER            std_ulogic_vector
     --                        BOOLEAN     std_ulogic_vector   INTEGER
     --                        std_ulogic  INTEGER            std_ulogic_vector
     --                        std_ulogic  std_ulogic_vector   INTEGER
     --                                     
     --     NOTE          : The std_ulogic_vector operands are assumed to be  
     --                     in  DefaultRegMode. If not they will be converted
     --                     to DefaultRegMode in the compare procedure. 
     --                     These vectors may be of any length.
     --     Use           : 
     --                      VARIABLE a : std_ulogic_vector ( 7 DOWNTO 0 ) := X"FF";
     --                      VARIABLE b : INTEGER;
     --                      IF ( a = b )  THEN 
     --     
     --     See Also      : RegEqual, RegNotEqual,
     -------------------------------------------------------------------------------
     FUNCTION  "=" ( CONSTANT l  : std_ulogic_vector;
		     CONSTANT r  : std_ulogic_vector
		   ) RETURN std_ulogic;
     -------------------------------------------------------------------------------
     FUNCTION  "=" ( CONSTANT l  : std_ulogic_vector;
		     CONSTANT r  : INTEGER
		   ) RETURN BOOLEAN;
     -- -----------------------------------------------------------------------------
     FUNCTION  "=" ( CONSTANT l  : INTEGER   ;
		     CONSTANT r  : std_ulogic_vector 
		   ) RETURN BOOLEAN;
     -------------------------------------------------------------------------------
     FUNCTION  "=" ( CONSTANT l  : std_ulogic_vector;
		     CONSTANT r  : INTEGER
		   ) RETURN std_ulogic;

     -- -----------------------------------------------------------------------------
     FUNCTION  "=" ( CONSTANT l  : INTEGER   ;
		     CONSTANT r  : std_ulogic_vector 
		   ) RETURN std_ulogic;
     -------------------------------------------------------------------------------
     --     Function Name : Overloaded "=" operator
     -- 1.2.2 and 1.2.4
     --     Purpose       : Equality relational operator for bit_vector : integer.
     --
     --     Parameters    :     result         left       right
     --                        BOOLEAN       INTEGER   bit_vector 
     --                        BOOLEAN      bit_vector   INTEGER
     --
     --     NOTE          : The bit_vector operands are assumed to be 
     --                     in  DefaultRegMode. If not they will be converted
     --                     to DefaultRegMode in the compare procedure. 
     --                     These vectors may be of any length.
     --     Use           :
     --                      VARIABLE a : bit_vector ( 7 DOWNTO 0 ) := X"FF";
     --                      VARIABLE b : INTEGER;
     --                      IF ( a = b )  THEN
     --
     --     See Also      : compare, RegLessThan, RegGreaterThan,
     -------------------------------------------------------------------------------
     FUNCTION  "=" ( CONSTANT l  : bit_vector;
		     CONSTANT r  : bit_vector
		   ) RETURN bit;
     -------------------------------------------------------------------------------
     FUNCTION  "=" ( CONSTANT l  : bit_vector;
		     CONSTANT r  : INTEGER
		   ) RETURN BOOLEAN;
     -- -----------------------------------------------------------------------------
     FUNCTION  "=" ( CONSTANT l  : INTEGER   ;
		     CONSTANT r  : bit_vector 
		   ) RETURN BOOLEAN;
     -------------------------------------------------------------------------------
     FUNCTION  "=" ( CONSTANT l  : bit_vector;
		     CONSTANT r  : INTEGER
		   ) RETURN bit;
     -- -----------------------------------------------------------------------------
     FUNCTION  "=" ( CONSTANT l  : INTEGER   ;
		     CONSTANT r  : bit_vector 
		   ) RETURN bit;

     -------------------------------------------------------------------------------
     --     Function Name : Overloaded "/=" operator
     --   1.2.1 and 1.2.3  
     --     Purpose       : Un-equality relational operator for std_logic_vector : integer.
     --     
     --     Parameters    :     result         left              right
     --                        std_ulogic  std_logic_vector   std_logic_vector
     --                        BOOLEAN     INTEGER            std_logic_vector
     --                        BOOLEAN     std_logic_vector   INTEGER
     --                        std_ulogic  INTEGER            std_logic_vector
     --                        std_ulogic  std_logic_vector   INTEGER
     --                                     
     --     NOTE          : The std_logic_vector operands are assumed to be  
     --                     in  DefaultRegMode. If not they will be converted
     --                     to DefaultRegMode in the compare procedure. 
     --                     These vectors may be of any length.
     --     Use           : 
     --                      VARIABLE a : std_logic_vector ( 7 DOWNTO 0 ) := X"FF";
     --                      VARIABLE b : INTEGER;
     --                      IF ( a /= b )  THEN 
     --     
     --     See Also      : RegEqual, RegNotEqual,
     -------------------------------------------------------------------------------
     FUNCTION  "/=" ( CONSTANT l  : std_logic_vector;
		     CONSTANT r  : std_logic_vector
		   ) RETURN std_ulogic;
     -------------------------------------------------------------------------------
     FUNCTION  "/=" ( CONSTANT l  : std_logic_vector;
		     CONSTANT r  : INTEGER
		   ) RETURN BOOLEAN;
     -- -----------------------------------------------------------------------------
     FUNCTION  "/=" ( CONSTANT l  : INTEGER   ;
		     CONSTANT r  : std_logic_vector 
		   ) RETURN BOOLEAN;
     -------------------------------------------------------------------------------
     FUNCTION  "/=" ( CONSTANT l  : std_logic_vector;
		     CONSTANT r  : INTEGER
		   ) RETURN std_ulogic;

     -- -----------------------------------------------------------------------------
     FUNCTION  "/=" ( CONSTANT l  : INTEGER   ;
		     CONSTANT r  : std_logic_vector 
		   ) RETURN std_ulogic;
     -------------------------------------------------------------------------------
     --     Function Name : Overloaded "/=" operator
     --   1.2.1 and 1.2.3  
     --     Purpose       : Un-equality relational operator for std_ulogic_vector : integer.
     --     
     --     Parameters    :     result         left              right
     --                        std_ulogic  std_ulogic_vector   std_ulogic_vector
     --                        BOOLEAN     INTEGER            std_ulogic_vector
     --                        BOOLEAN     std_ulogic_vector   INTEGER
     --                        std_ulogic  INTEGER            std_ulogic_vector
     --                        std_ulogic  std_ulogic_vector   INTEGER
     --                                     
     --     NOTE          : The std_ulogic_vector operands are assumed to be  
     --                     in  DefaultRegMode. If not they will be converted
     --                     to DefaultRegMode in the compare procedure. 
     --                     These vectors may be of any length.
     --     Use           : 
     --                      VARIABLE a : std_ulogic_vector ( 7 DOWNTO 0 ) := X"FF";
     --                      VARIABLE b : INTEGER;
     --                      IF ( a /= b )  THEN 
     --     
     --     See Also      : RegEqual, RegNotEqual,
     -------------------------------------------------------------------------------
     FUNCTION  "/=" ( CONSTANT l  : std_ulogic_vector;
		     CONSTANT r  : std_ulogic_vector
		   ) RETURN std_ulogic;
     -------------------------------------------------------------------------------
     FUNCTION  "/=" ( CONSTANT l  : std_ulogic_vector;
		     CONSTANT r  : INTEGER
		   ) RETURN BOOLEAN;
     -- -----------------------------------------------------------------------------
     FUNCTION  "/=" ( CONSTANT l  : INTEGER   ;
		     CONSTANT r  : std_ulogic_vector 
		   ) RETURN BOOLEAN;
     -------------------------------------------------------------------------------
     FUNCTION  "/=" ( CONSTANT l  : std_ulogic_vector;
		     CONSTANT r  : INTEGER
		   ) RETURN std_ulogic;

     -- -----------------------------------------------------------------------------
     FUNCTION  "/=" ( CONSTANT l  : INTEGER   ;
		     CONSTANT r  : std_ulogic_vector 
		   ) RETURN std_ulogic;
     -------------------------------------------------------------------------------
     --     Function Name : Overloaded "/=" operator
     -- 1.2.2 and 1.2.4
     --     Purpose       : Un-equality relational operator for bit_vector : integer.
     --
     --     Parameters    :     result         left       right
     --                        BOOLEAN       INTEGER   bit_vector 
     --                        BOOLEAN      bit_vector   INTEGER
     --
     --     NOTE          : The bit_vector operands are assumed to be 
     --                     in  DefaultRegMode. If not they will be converted
     --                     to DefaultRegMode in the compare procedure. 
     --                     These vectors may be of any length.
     --     Use           :
     --                      VARIABLE a : bit_vector ( 7 DOWNTO 0 ) := X"FF";
     --                      VARIABLE b : INTEGER;
     --                      IF ( a /= b )  THEN
     --
     --     See Also      : compare, RegLessThan, RegGreaterThan,
     -------------------------------------------------------------------------------
     FUNCTION  "/=" ( CONSTANT l  : bit_vector;
		     CONSTANT r  : bit_vector
		   ) RETURN bit;
     -------------------------------------------------------------------------------
     FUNCTION  "/=" ( CONSTANT l  : bit_vector;
		     CONSTANT r  : INTEGER
		   ) RETURN BOOLEAN;
     -- -----------------------------------------------------------------------------
     FUNCTION  "/=" ( CONSTANT l  : INTEGER   ;
		     CONSTANT r  : bit_vector 
		   ) RETURN BOOLEAN;
     -------------------------------------------------------------------------------
     FUNCTION  "/=" ( CONSTANT l  : bit_vector;
		     CONSTANT r  : INTEGER
		   ) RETURN bit;
     -- -----------------------------------------------------------------------------
     FUNCTION  "/=" ( CONSTANT l  : INTEGER   ;
		     CONSTANT r  : bit_vector 
		   ) RETURN bit;
     -------------------------------------------------------------------------------
     --     Function Name : Overloaded "<" operator
     -- 1.2.18 and 1.2.20     
     --     Purpose       : Less-than relational operator for bit_vectors.
     --     
     --     Parameters    :     result         left       right
     --                        BOOLEAN       INTEGER    bit_vector
     --                        BOOLEAN      bit_vector   INTEGER
     --     
     --     NOTE          : The bit_vector operands are assumed to be 
     --                     in  DefaultRegMode. If not they will be converted
     --                     to DefaultRegMode in the compare procedure. 
     --                     These vectors may be of any length.
     --     Use           :
     --                      VARIABLE a : bit_vector ( 7 DOWNTO 0 ) := X"FF";
     --                      VARIABLE b : INTEGER;
     --                      IF ( a < b )  THEN 
     --     
     --     See Also      : compare, RegLessThan, RegGreaterThan,
     -------------------------------------------------------------------------------
     FUNCTION  "<" ( CONSTANT l  : bit_vector;
		     CONSTANT r  : bit_vector
		   ) RETURN bit;
     -------------------------------------------------------------------------------
     FUNCTION  "<" ( CONSTANT l  : bit_vector;
		     CONSTANT r  : INTEGER
		   ) RETURN BOOLEAN;
     -- -----------------------------------------------------------------------------
     FUNCTION  "<" ( CONSTANT l  : INTEGER   ;
		     CONSTANT r  : bit_vector 
		   ) RETURN BOOLEAN;
     -------------------------------------------------------------------------------
     FUNCTION  "<" ( CONSTANT l  : bit_vector;
		     CONSTANT r  : INTEGER
		   ) RETURN bit;
     -- -----------------------------------------------------------------------------
     FUNCTION  "<" ( CONSTANT l  : INTEGER   ;
		     CONSTANT r  : bit_vector 
		   ) RETURN bit;
     -------------------------------------------------------------------------------
     --     Function Name : Overloaded "<" operator
     --
     --     Purpose       : Less-than relational operator for std_logic_vectors.
     --
     --     Parameters    :     result         left       right
     --                        std_ulogic  std_logic_vector   std_logic_vector
     --                        BOOLEAN     INTEGER            std_logic_vector
     --                        BOOLEAN     std_logic_vector   INTEGER
     --                        std_ulogic  INTEGER            std_logic_vector
     --                        std_ulogic  std_logic_vector   INTEGER
     --
     --     NOTE          : The std_logic_vector operands are assumed to be 
     --                     in  DefaultRegMode. If not they will be converted
     --                     to DefaultRegMode in the compare procedure. 
     --                     These vectors may be of any length.
     --     Use           :
     --                      VARIABLE a : std_logic_vector ( 7 DOWNTO 0 ) := X"FF";
     --                      VARIABLE b : INTEGER;
     --                      IF ( a < b )  THEN
     --
     --     See Also      : compare, RegLessThan, RegGreaterThan,
     -------------------------------------------------------------------------------
     FUNCTION  "<" ( CONSTANT l  : std_logic_vector;
		     CONSTANT r  : std_logic_vector
		   ) RETURN std_ulogic;
     -------------------------------------------------------------------------------
     FUNCTION  "<" ( CONSTANT l  : std_logic_vector;
		     CONSTANT r  : INTEGER
		   ) RETURN BOOLEAN;
     -- -----------------------------------------------------------------------------
     FUNCTION  "<" ( CONSTANT l  : INTEGER   ;
		     CONSTANT r  : std_logic_vector 
		   ) RETURN BOOLEAN;
     -------------------------------------------------------------------------------
     FUNCTION  "<" ( CONSTANT l  : std_logic_vector;
		     CONSTANT r  : INTEGER
		   ) RETURN std_ulogic;
     -- -----------------------------------------------------------------------------
     FUNCTION  "<" ( CONSTANT l  : INTEGER   ;
		     CONSTANT r  : std_logic_vector 
		   ) RETURN std_ulogic;
     -------------------------------------------------------------------------------
     --     Function Name : Overloaded "<" operator
     --
     --     Purpose       : Less-than relational operator for std_logic_vectors.
     --
     --     Parameters    :     result         left       right
     --                        std_ulogic  std_ulogic_vector   std_ulogic_vector
     --                        BOOLEAN     INTEGER            std_ulogic_vector
     --                        BOOLEAN     std_ulogic_vector   INTEGER
     --                        std_ulogic  INTEGER            std_ulogic_vector
     --                        std_ulogic  std_ulogic_vector   INTEGER  
     --
     --     NOTE          : The std_ulogic_vector operands are assumed to be 
     --                     in  DefaultRegMode. If not they will be converted
     --                     to DefaultRegMode in the compare procedure. 
     --                     These vectors may be of any length.
     --     Use           :
     --                      VARIABLE a : std_ulogic_vector ( 7 DOWNTO 0 ) := X"FF";
     --                      VARIABLE b : INTEGER;
     --                      IF ( a < b )  THEN
     --
     --     See Also      : compare, RegLessThan, RegGreaterThan,
     -------------------------------------------------------------------------------
     FUNCTION  "<" ( CONSTANT l  : std_ulogic_vector;
		     CONSTANT r  : std_ulogic_vector
		   ) RETURN std_ulogic;
     -------------------------------------------------------------------------------
     FUNCTION  "<" ( CONSTANT l  : std_ulogic_vector;
		     CONSTANT r  : INTEGER
		   ) RETURN BOOLEAN;
     -- -----------------------------------------------------------------------------
     FUNCTION  "<" ( CONSTANT l  : INTEGER   ;
		     CONSTANT r  : std_ulogic_vector 
		   ) RETURN BOOLEAN;
     -------------------------------------------------------------------------------
     FUNCTION  "<" ( CONSTANT l  : std_ulogic_vector;
		     CONSTANT r  : INTEGER
		   ) RETURN std_ulogic;
     -- -----------------------------------------------------------------------------
     FUNCTION  "<" ( CONSTANT l  : INTEGER   ;
		     CONSTANT r  : std_ulogic_vector 
		   ) RETURN std_ulogic;
     -------------------------------------------------------------------------------
     --     Function Name : Overloaded "<=" operator
     -- 1.2.26 and 1.2.28     
     --     Purpose       : Less-than-or-equal relational operator for bit_vectors.
     --     
     --     Parameters    :     result         left       right
     --                        BOOLEAN       INTEGER    bit_vector
     --                        BOOLEAN      bit_vector   INTEGER
     --     
     --     NOTE          : The bit_vector operands are assumed to be 
     --                     in  DefaultRegMode. If not they will be converted
     --                     to DefaultRegMode in the compare procedure. 
     --                     These vectors may be of any length.
     --     Use           :
     --                      VARIABLE a : bit_vector ( 7 DOWNTO 0 ) := X"FF";
     --                      VARIABLE b : INTEGER;
     --                      IF ( a <= b )  THEN 
     --     
     --     See Also      : compare, RegLessThan, RegGreaterThan,
     -------------------------------------------------------------------------------
     FUNCTION  "<=" ( CONSTANT l  : bit_vector;
		     CONSTANT r  : bit_vector
		   ) RETURN bit;
     -------------------------------------------------------------------------------
     FUNCTION  "<=" ( CONSTANT l  : bit_vector;
		      CONSTANT r  : INTEGER
		    ) RETURN BOOLEAN;
     -- -----------------------------------------------------------------------------
     FUNCTION  "<=" ( CONSTANT l  : INTEGER   ;
		      CONSTANT r  : bit_vector 
		    ) RETURN BOOLEAN;
     -------------------------------------------------------------------------------
     FUNCTION  "<=" ( CONSTANT l  : bit_vector;
		      CONSTANT r  : INTEGER
		    ) RETURN bit;
     -- -----------------------------------------------------------------------------
     FUNCTION  "<=" ( CONSTANT l  : INTEGER   ;
		      CONSTANT r  : bit_vector 
		    ) RETURN bit;
     -------------------------------------------------------------------------------
     --     Function Name : Overloaded "<=" operator
     --    
     --     Purpose       : Less-than-or-equal relational operator for 
     --                     std_logic_vectors.
     --     
     --     Parameters    :     result         left       right
     --                        std_ulogic  std_logic_vector   std_logic_vector
     --                        BOOLEAN     INTEGER            std_logic_vector
     --                        BOOLEAN     std_logic_vector   INTEGER
     --                        std_ulogic  INTEGER            std_logic_vector
     --                        std_ulogic  std_logic_vector   INTEGER 
     --     
     --     NOTE          : The std_logic_vector operands are assumed to be 
     --                     in  DefaultRegMode. If not they will be converted
     --                     to DefaultRegMode in the compare procedure. 
     --                     These vectors may be of any length.
     --     Use           : 
     --                      VARIABLE a : std_logic_vector ( 7 DOWNTO 0 ) := X"FF";
     --                      VARIABLE b : INTEGER;
     --                      IF ( a <= b )  THEN 
     --     
     --     See Also      : compare, RegLessThan, RegGreaterThan,
     -------------------------------------------------------------------------------
     FUNCTION  "<=" ( CONSTANT l  : std_logic_vector;
		      CONSTANT r  : std_logic_vector
		    ) RETURN std_ulogic;
     -------------------------------------------------------------------------------
     FUNCTION  "<=" ( CONSTANT l  : std_logic_vector;
		      CONSTANT r  : INTEGER
		    ) RETURN BOOLEAN;
     -- -----------------------------------------------------------------------------
     FUNCTION  "<=" ( CONSTANT l  : INTEGER   ;
		      CONSTANT r  : std_logic_vector 
		    ) RETURN BOOLEAN;
     -------------------------------------------------------------------------------
     FUNCTION  "<=" ( CONSTANT l  : std_logic_vector;
		      CONSTANT r  : INTEGER
		    ) RETURN std_ulogic;
     -- -----------------------------------------------------------------------------
     FUNCTION  "<=" ( CONSTANT l  : INTEGER   ;
		      CONSTANT r  : std_logic_vector 
		    ) RETURN std_ulogic;
     -------------------------------------------------------------------------------
     --     Function Name : Overloaded "<=" operator
     --    
     --     Purpose       : Less-than-or-equal relational operator for 
     --                     std_ulogic_vectors.
     --     
     --     Parameters    :     result         left       right
     --                        std_ulogic  std_ulogic_vector   std_ulogic_vector
     --                        BOOLEAN     INTEGER            std_ulogic_vector
     --                        BOOLEAN     std_ulogic_vector   INTEGER
     --                        std_ulogic  INTEGER            std_ulogic_vector
     --                        std_ulogic  std_ulogic_vector   INTEGER 
     --     
     --     NOTE          : The std_ulogic_vector operands are assumed to be 
     --                     in  DefaultRegMode. If not they will be converted
     --                     to DefaultRegMode in the compare procedure. 
     --                     These vectors may be of any length.
     --     Use           : 
     --                      VARIABLE a : std_ulogic_vector ( 7 DOWNTO 0 ) := X"FF";
     --                      VARIABLE b : INTEGER;
     --                      IF ( a <= b )  THEN 
     --     
     --     See Also      : compare, RegLessThan, RegGreaterThan,
     -------------------------------------------------------------------------------
     FUNCTION  "<=" ( CONSTANT l  : std_ulogic_vector;
		      CONSTANT r  : std_ulogic_vector
		    ) RETURN std_ulogic;
     -------------------------------------------------------------------------------
     FUNCTION  "<=" ( CONSTANT l  : std_ulogic_vector;
		      CONSTANT r  : INTEGER
		    ) RETURN BOOLEAN;
     -- -----------------------------------------------------------------------------
     FUNCTION  "<=" ( CONSTANT l  : INTEGER   ;
		      CONSTANT r  : std_ulogic_vector 
		    ) RETURN BOOLEAN;
     -------------------------------------------------------------------------------
     FUNCTION  "<=" ( CONSTANT l  : std_ulogic_vector;
		      CONSTANT r  : INTEGER
		    ) RETURN std_ulogic;
     -- -----------------------------------------------------------------------------
     FUNCTION  "<=" ( CONSTANT l  : INTEGER   ;
		      CONSTANT r  : std_ulogic_vector 
		    ) RETURN std_ulogic;

     -------------------------------------------------------------------------------
     --     Function Name : Overloaded ">" operator
     -- 1.2.18 and 1.2.20     
     --     Purpose       : Greater-than relational operator for bit_vectors.
     --     
     --     Parameters    :     result         left       right
     --                        BOOLEAN       INTEGER    bit_vector
     --                        BOOLEAN      bit_vector   INTEGER
     --     
     --     NOTE          : The bit_vector operands are assumed to be 
     --                     in  DefaultRegMode. If not they will be converted
     --                     to DefaultRegMode in the compare procedure. 
     --                     These vectors may be of any length.
     --     Use           :
     --                      VARIABLE a : bit_vector ( 7 DOWNTO 0 ) := X"FF";
     --                      VARIABLE b : INTEGER;
     --                      IF ( a > b )  THEN 
     --     
     --     See Also      : compare, RegLessThan, RegGreaterThan,
     -------------------------------------------------------------------------------
     FUNCTION  ">" ( CONSTANT l  : bit_vector;
		     CONSTANT r  : bit_vector
		   ) RETURN bit;
     -------------------------------------------------------------------------------
     FUNCTION  ">" ( CONSTANT l  : bit_vector;
		     CONSTANT r  : INTEGER
		   ) RETURN BOOLEAN;
     -- -----------------------------------------------------------------------------
     FUNCTION  ">" ( CONSTANT l  : INTEGER   ;
		     CONSTANT r  : bit_vector 
		   ) RETURN BOOLEAN;
     -------------------------------------------------------------------------------
     FUNCTION  ">" ( CONSTANT l  : bit_vector;
		     CONSTANT r  : INTEGER
		   ) RETURN bit;
     -- -----------------------------------------------------------------------------
     FUNCTION  ">" ( CONSTANT l  : INTEGER   ;
		     CONSTANT r  : bit_vector 
		   ) RETURN bit;
     -------------------------------------------------------------------------------
     --     Function Name : Overloaded ">" operator
     --
     --     Purpose       : Greater-than relational operator for std_logic_vectors.
     --
     --     Parameters    :     result         left       right
     --                        std_ulogic  std_logic_vector   std_logic_vector
     --                        BOOLEAN     INTEGER            std_logic_vector
     --                        BOOLEAN     std_logic_vector   INTEGER
     --                        std_ulogic  INTEGER            std_logic_vector
     --                        std_ulogic  std_logic_vector   INTEGER
     --
     --     NOTE          : The std_logic_vector operands are assumed to be 
     --                     in  DefaultRegMode. If not they will be converted
     --                     to DefaultRegMode in the compare procedure. 
     --                     These vectors may be of any length.
     --     Use           :
     --                      VARIABLE a : std_logic_vector ( 7 DOWNTO 0 ) := X"FF";
     --                      VARIABLE b : INTEGER;
     --                      IF ( a > b )  THEN
     --
     --     See Also      : compare, RegLessThan, RegGreaterThan,
     -------------------------------------------------------------------------------
     FUNCTION  ">" ( CONSTANT l  : std_logic_vector;
		     CONSTANT r  : std_logic_vector
		   ) RETURN std_ulogic;
     -------------------------------------------------------------------------------
     FUNCTION  ">" ( CONSTANT l  : std_logic_vector;
		     CONSTANT r  : INTEGER
		   ) RETURN BOOLEAN;
     -- -----------------------------------------------------------------------------
     FUNCTION  ">" ( CONSTANT l  : INTEGER   ;
		     CONSTANT r  : std_logic_vector 
		   ) RETURN BOOLEAN;
     -------------------------------------------------------------------------------
     FUNCTION  ">" ( CONSTANT l  : std_logic_vector;
		     CONSTANT r  : INTEGER
		   ) RETURN std_ulogic;
     -- -----------------------------------------------------------------------------
     FUNCTION  ">" ( CONSTANT l  : INTEGER   ;
		     CONSTANT r  : std_logic_vector 
		   ) RETURN std_ulogic;
     -------------------------------------------------------------------------------
     --     Function Name : Overloaded ">" operator
     --
     --     Purpose       : Greater-than relational operator for std_logic_vectors.
     --
     --     Parameters    :     result         left       right
     --                        std_ulogic  std_ulogic_vector   std_ulogic_vector
     --                        BOOLEAN     INTEGER            std_ulogic_vector
     --                        BOOLEAN     std_ulogic_vector   INTEGER
     --                        std_ulogic  INTEGER            std_ulogic_vector
     --                        std_ulogic  std_ulogic_vector   INTEGER  
     --
     --     NOTE          : The std_ulogic_vector operands are assumed to be 
     --                     in  DefaultRegMode. If not they will be converted
     --                     to DefaultRegMode in the compare procedure. 
     --                     These vectors may be of any length.
     --     Use           :
     --                      VARIABLE a : std_ulogic_vector ( 7 DOWNTO 0 ) := X"FF";
     --                      VARIABLE b : INTEGER;
     --                      IF ( a > b )  THEN
     --
     --     See Also      : compare, RegLessThan, RegGreaterThan,
     -------------------------------------------------------------------------------
     FUNCTION  ">" ( CONSTANT l  : std_ulogic_vector;
		     CONSTANT r  : std_ulogic_vector
		   ) RETURN std_ulogic;
     -------------------------------------------------------------------------------
     FUNCTION  ">" ( CONSTANT l  : std_ulogic_vector;
		     CONSTANT r  : INTEGER
		   ) RETURN BOOLEAN;
     -- -----------------------------------------------------------------------------
     FUNCTION  ">" ( CONSTANT l  : INTEGER   ;
		     CONSTANT r  : std_ulogic_vector 
		   ) RETURN BOOLEAN;
     -------------------------------------------------------------------------------
     FUNCTION  ">" ( CONSTANT l  : std_ulogic_vector;
		     CONSTANT r  : INTEGER
		   ) RETURN std_ulogic;
     -- -----------------------------------------------------------------------------
     FUNCTION  ">" ( CONSTANT l  : INTEGER   ;
		     CONSTANT r  : std_ulogic_vector 
		   ) RETURN std_ulogic;
     -------------------------------------------------------------------------------
     --     Function Name : Overloaded ">=" operator
     -- 1.2.26 and 1.2.28     
     --     Purpose       : Greater-than-or-equal relational operator for bit_vectors.
     --     
     --     Parameters    :     result         left       right
     --                        BOOLEAN       INTEGER    bit_vector
     --                        BOOLEAN      bit_vector   INTEGER
     --     
     --     NOTE          : The bit_vector operands are assumed to be 
     --                     in  DefaultRegMode. If not they will be converted
     --                     to DefaultRegMode in the compare procedure. 
     --                     These vectors may be of any length.
     --     Use           :
     --                      VARIABLE a : bit_vector ( 7 DOWNTO 0 ) := X"FF";
     --                      VARIABLE b : INTEGER;
     --                      IF ( a >= b )  THEN 
     --     
     --     See Also      : compare, RegLessThan, RegGreaterThan,
     -------------------------------------------------------------------------------
     FUNCTION  ">=" ( CONSTANT l  : bit_vector;
		     CONSTANT r  : bit_vector
		   ) RETURN bit;
     -------------------------------------------------------------------------------
     FUNCTION  ">=" ( CONSTANT l  : bit_vector;
		      CONSTANT r  : INTEGER
		    ) RETURN BOOLEAN;
     -- -----------------------------------------------------------------------------
     FUNCTION  ">=" ( CONSTANT l  : INTEGER   ;
		      CONSTANT r  : bit_vector 
		    ) RETURN BOOLEAN;
     -------------------------------------------------------------------------------
     FUNCTION  ">=" ( CONSTANT l  : bit_vector;
		      CONSTANT r  : INTEGER
		    ) RETURN bit;
     -- -----------------------------------------------------------------------------
     FUNCTION  ">=" ( CONSTANT l  : INTEGER   ;
		      CONSTANT r  : bit_vector 
		    ) RETURN bit;
     -------------------------------------------------------------------------------
     --     Function Name : Overloaded ">=" operator
     --    
     --     Purpose       : Greater-than-or-equal relational operator for 
     --                     std_logic_vectors.
     --     
     --     Parameters    :     result         left       right
     --                        std_ulogic  std_logic_vector   std_logic_vector
     --                        BOOLEAN     INTEGER            std_logic_vector
     --                        BOOLEAN     std_logic_vector   INTEGER
     --                        std_ulogic  INTEGER            std_logic_vector
     --                        std_ulogic  std_logic_vector   INTEGER 
     --     
     --     NOTE          : The std_logic_vector operands are assumed to be 
     --                     in  DefaultRegMode. If not they will be converted
     --                     to DefaultRegMode in the compare procedure. 
     --                     These vectors may be of any length.
     --     Use           : 
     --                      VARIABLE a : std_logic_vector ( 7 DOWNTO 0 ) := X"FF";
     --                      VARIABLE b : INTEGER;
     --                      IF ( a >= b )  THEN 
     --     
     --     See Also      : compare, RegLessThan, RegGreaterThan,
     -------------------------------------------------------------------------------
     FUNCTION  ">=" ( CONSTANT l  : std_logic_vector;
		      CONSTANT r  : std_logic_vector
		    ) RETURN std_ulogic;
     -------------------------------------------------------------------------------
     FUNCTION  ">=" ( CONSTANT l  : std_logic_vector;
		      CONSTANT r  : INTEGER
		    ) RETURN BOOLEAN;
     -- -----------------------------------------------------------------------------
     FUNCTION  ">=" ( CONSTANT l  : INTEGER   ;
		      CONSTANT r  : std_logic_vector 
		    ) RETURN BOOLEAN;
     -------------------------------------------------------------------------------
     FUNCTION  ">=" ( CONSTANT l  : std_logic_vector;
		      CONSTANT r  : INTEGER
		    ) RETURN std_ulogic;
     -- -----------------------------------------------------------------------------
     FUNCTION  ">=" ( CONSTANT l  : INTEGER   ;
		      CONSTANT r  : std_logic_vector 
		    ) RETURN std_ulogic;
     -------------------------------------------------------------------------------
     --     Function Name : Overloaded ">=" operator
     --    
     --     Purpose       : Greater-than-or-equal relational operator for 
     --                     std_ulogic_vectors.
     --     
     --     Parameters    :     result         left       right
     --                        std_ulogic  std_ulogic_vector   std_ulogic_vector
     --                        BOOLEAN     INTEGER            std_ulogic_vector
     --                        BOOLEAN     std_ulogic_vector   INTEGER
     --                        std_ulogic  INTEGER            std_ulogic_vector
     --                        std_ulogic  std_ulogic_vector   INTEGER 
     --     
     --     NOTE          : The std_ulogic_vector operands are assumed to be 
     --                     in  DefaultRegMode. If not they will be converted
     --                     to DefaultRegMode in the compare procedure. 
     --                     These vectors may be of any length.
     --     Use           : 
     --                      VARIABLE a : std_ulogic_vector ( 7 DOWNTO 0 ) := X"FF";
     --                      VARIABLE b : INTEGER;
     --                      IF ( a >= b )  THEN 
     --     
     --     See Also      : compare, RegLessThan, RegGreaterThan,
     -------------------------------------------------------------------------------
     FUNCTION  ">=" ( CONSTANT l  : std_ulogic_vector;
		      CONSTANT r  : std_ulogic_vector
		    ) RETURN std_ulogic;
     -------------------------------------------------------------------------------
     FUNCTION  ">=" ( CONSTANT l  : std_ulogic_vector;
		      CONSTANT r  : INTEGER
		    ) RETURN BOOLEAN;
     -- -----------------------------------------------------------------------------
     FUNCTION  ">=" ( CONSTANT l  : INTEGER   ;
		      CONSTANT r  : std_ulogic_vector 
		    ) RETURN BOOLEAN;
     -------------------------------------------------------------------------------
     FUNCTION  ">=" ( CONSTANT l  : std_ulogic_vector;
		      CONSTANT r  : INTEGER
		    ) RETURN std_ulogic;
     -- -----------------------------------------------------------------------------
     FUNCTION  ">=" ( CONSTANT l  : INTEGER   ;
		      CONSTANT r  : std_ulogic_vector 
		    ) RETURN std_ulogic;
--+-----------------------------------------------------------------------------
--|     Function Name  : To_TwosComp
--| 1.8.7
--|     Overloading    : None
--|  
--|     Purpose        : Convert a BIT_VECTOR to Two's Compliment Notation.
--|  
--|     Parameters     :
--|                      SrcReg     - input  BIT_VECTOR, the vector to be read.
--|                      SrcRegMode - input  regmode_type, indicating the format of
--|                                the input BIT_VECTOR.   Default is TwosComp.
--|
--|     Result         : BIT_VECTOR, the vector in Two's complement notation.
--|
--|     Use            :
--|                      VARIABLE vect : BIT_VECTOR ( 15 DOWNTO 0 );
--|                      vect := To_TwosComp ( B"101",  UnSigned ); -- set to +5
--|
--|     See Also       : To_BitVector, To_Integer, To_TwosComp
--|-----------------------------------------------------------------------------
    FUNCTION To_TwosComp  ( CONSTANT SrcReg      : IN BIT_VECTOR;
                            CONSTANT SrcRegMode  : IN regmode_type 
                     -- synopsys synthesis_off
						      := DefaultRegMode
                     -- synopsys synthesis_on

                          ) RETURN BIT_VECTOR;
    -------------------------------------------------------------------------------
    --     Function Name  : To_TwosComp
    -- 1.8.8
    --     Overloading    : None
    --    
    --     Purpose        : Convert an std_logic_vector to Two's Compliment Notation.
    --     
    --     Parameters     : 
    --                      SrcReg    - input  std_logic_vector, the vector to be read.
    --                      SrcRegMode - input  regmode_type, indicating the format of
    --                              the input std_logic_vector.   Default is TwosComp.
    --     
    --     Result         : std_logic_vector, the vector in Two's complement notation.
    --
    --     Use            : 
    --                      VARIABLE vect : std_logic_vector ( 15 DOWNTO 0 );
    --                      vect := To_TwosComp ( B"101", UnSigned ); -- set to +5
    --     
    --     See Also       : To_StdLogicVector, To_Integer, To_TwosComp, From_TwosComp
    -------------------------------------------------------------------------------
    FUNCTION To_TwosComp  ( CONSTANT SrcReg      : IN std_logic_vector;
                            CONSTANT SrcRegMode  : IN regmode_type  
                     -- synopsys synthesis_off
						      := DefaultRegMode 
                     -- synopsys synthesis_on
                          ) RETURN std_logic_vector;
    -------------------------------------------------------------------------------
    --     Function Name  : To_TwosComp
    -- 1.8.8
    --     Overloading    : None
    --    
    --     Purpose        : Convert an std_ulogic_vector to Two's Compliment Notation.
    --     
    --     Parameters     : 
    --                      SrcReg   - input  std_ulogic_vector, the vector to be read.
    --                      SrcRegMode - input  regmode_type, indicating the format of
    --                             the input std_ulogic_vector.   Default is TwosComp.
    --     
    --     Result         : std_ulogic_vector, the vector in Two's complement notation.
    --
    --     Use            : 
    --                      VARIABLE vect : std_ulogic_vector ( 15 DOWNTO 0 );
    --                      vect := To_TwosComp ( B"101", UnSigned ); -- set to +5
    --     
    --     See Also       : To_StdLogicVector, To_Integer, To_TwosComp, From_TwosComp
    -------------------------------------------------------------------------------
    FUNCTION To_TwosComp  ( CONSTANT SrcReg      : IN std_ulogic_vector;
                            CONSTANT SrcRegMode  : IN regmode_type  
                     -- synopsys synthesis_off
						      := DefaultRegMode 
                     -- synopsys synthesis_on
                          ) RETURN std_ulogic_vector;
--+-----------------------------------------------------------------------------
--|     Function Name  : To_Unsign
--| 1.8.11
--|     Overloading    : None
--| 
--|     Purpose        : Convert a BIT_VECTOR to Unsigned Notation.
--| 
--|     Parameters     :
--|                      SrcReg     - input  BIT_VECTOR, the vector to be read.
--|                      SrcRegMode - input  regmode_type, indicating the format of
--|                                the input BIT_VECTOR.   Default is TwosComp.
--|
--|     Result         : BIT_VECTOR, the vector in unsigned notation. 
--|
--|
--|     Use            :
--|                      VARIABLE vect : BIT_VECTOR ( 15 DOWNTO 0 );
--|                      vect := To_Unsign ( B"0101", SignMagnitude ); -- set to +5
--|
--|     See Also       : to_BitVector, to_Integer, To_TwosComp, From_TwosComp
--|-----------------------------------------------------------------------------
    FUNCTION To_Unsign    ( CONSTANT SrcReg      : IN BIT_VECTOR;
                            CONSTANT SrcRegMode  : IN regmode_type  
                     -- synopsys synthesis_off
						      := DefaultRegMode 
                     -- synopsys synthesis_on
                          ) RETURN BIT_VECTOR;
    -------------------------------------------------------------------------------
    --     Function Name  : To_Unsign
    --
    --     Overloading    : None
    --
    --     Purpose        : Convert a std_logic_vector to Unsigned Notation.
    --
    --     Parameters     :
    --                      SrcReg     - input  std_logic_vector, the vector to be read.
    --                      SrcRegMode - input  regmode_type, indicating the format of
    --                              the input std_logic_vector.   Default is TwosComp.
    --
    --     Result         : std_logic_vector, the vector in unsigned notation.
    --
    --     Use            :
    --                      VARIABLE vect : std_logic_vector ( 15 DOWNTO 0 );
    --                      vect := To_Unsign ( B"0l01",SignMagnitude ); -- set to +5
    --
    --     See Also       : To_StdLogicVector, To_Integer, To_TwosComp, From_TwosComp
  -------------------------------------------------------------------------------
    FUNCTION To_Unsign    ( CONSTANT SrcReg      : IN std_logic_vector;
                            CONSTANT SrcRegMode  : IN regmode_type  
                     -- synopsys synthesis_off
						      := DefaultRegMode 
                     -- synopsys synthesis_on
                          ) RETURN std_logic_vector;
   -------------------------------------------------------------------------------
    --     Function Name  : To_Unsign
    --
    --     Overloading    : None
    --
    --     Purpose        : Convert an std_ulogic_vector to Unsigned Notation.
    --
    --     Parameters     :
    --                      SrcReg     - input  std_ulogic_vector, the vector to be read.
    --                      SrcRegMode - input  regmode_type, indicating the format of
    --                              the input std_ulogic_vector.   Default is TwosComp.
    --
    --     Result         : std_ulogic_vector, the vector in unsigned notation.
    --
    --     Use            :
    --                      VARIABLE vect : std_ulogic_vector ( 15 DOWNTO 0 );
    --                      vect := To_Unsign ( "0l01",SignMagnitude ); -- set to +5
    --
    --     See Also       : To_StdLogicVector, To_Integer, To_TwosComp, From_TwosComp
    ---------------------------------------------------------------------------------
    FUNCTION To_Unsign    ( CONSTANT SrcReg      : IN std_ulogic_vector;
                            CONSTANT SrcRegMode  : IN regmode_type  
                     -- synopsys synthesis_off
						      := DefaultRegMode 
                     -- synopsys synthesis_on
                          ) RETURN std_ulogic_vector;
    -------------------------------------------------------------------------------
    --     Function Name  : To_StdLogicVector
    --
    --     Overloading    : Procedure and Function.
    --
    --     Purpose        : Translate an INTEGER into a std_logic_vector.
    --
    --     Parameters     : intg    - input  INTEGER, the value to be translated.
    --                      width   - input  INTEGER, length of the return vector.
    --                                Default is IntegerBitLength  (Machine Integer
    --                                length).
    --                      SrcRegMode - input  regmode_type, indicating the format
    --                                   of the output std_logic_vector.   Default 
    --                                   is TwosComp.
    --
    --     Result        : std_logic_vector, the binary representation of the integer.
    --
    --     NOTE          : An ASSERTION message of severity ERROR if the conversion
    --                      fails:
    --                       * 'intg' is negative and UnSigned format is specified.
    --                         The absolute value of 'intg' is used.
    --                       * The length of 'SrcReg' is insufficient to hold the
    --                         binary value. The low order bits are returned.
    --
    --                      A runtime system error should occur if the value of
    --                      'width'  does not equal the expected return vector
    --                      length (from the context of the function usage).
     --     Use            :
    --                      VARIABLE vect : std_logic_vector ( 15 DOWNTO 0 );
    --
    --                      vect := To_StdLogicVector ( -294, 16, TwosComp );
    --
    --     See Also       : To_StdLogicVector, To_Integer, To_TwosComp
    -------------------------------------------------------------------------------
    FUNCTION To_StdLogicVector ( CONSTANT intg       : IN INTEGER;
                                 CONSTANT width      : IN NATURAL;
                                 CONSTANT SrcRegMode : IN regmode_type  
                     -- synopsys synthesis_off
						      := DefaultRegMode 
                     -- synopsys synthesis_on
                               ) RETURN std_logic_vector;
    -------------------------------------------------------------------------------
    --     Function Name  : To_StdULogicVector
    --
    --     Overloading    : Procedure and Function.
    --
    --     Purpose        : Translate an INTEGER into a std_ulogic_vector.
    --
    --     Parameters     : intg    - input  INTEGER, the value to be translated.
    --                      width   - input  INTEGER, length of the return vector.
    --                                Default is IntegerBitLength  (Machine Integer
    --                                length).
    --                      SrcRegMode - input  regmode_type, indicating the format
    --                                   of the output std_logic_vector.   Default 
    --                                   is TwosComp.
    --
    --     Result        : std_ulogic_vector
    --
    --     NOTE          : An ASSERTION message of severity ERROR if the conversion
    --                      fails:
    --                       * 'intg' is negative and UnSigned format is specified.
    --                         The absolute value of 'intg' is used.
    --                       * The length of 'SrcReg' is insufficient to hold the
    --                         binary value. The low order bits are returned.
    --
    --                      A runtime system error should occur if the value of
    --                      'width'  does not equal the expected return vector
    --                      length (from the context of the function usage).
    --     Use            :
    --                      VARIABLE vect : std_logic_vector ( 15 DOWNTO 0 );
    --
    --                      vect := To_StdLogicVector ( -294, 16, TwosComp );
    --
    --     See Also       : To_StdLogicVector, To_Integer, To_TwosComp
    -------------------------------------------------------------------------------
    FUNCTION To_StdULogicVector ( CONSTANT intg       : IN INTEGER;
                                  CONSTANT width      : IN NATURAL;
                                  CONSTANT SrcRegMode : IN regmode_type  
                     -- synopsys synthesis_off
						      := DefaultRegMode 
                     -- synopsys synthesis_on
                                ) RETURN std_ulogic_vector;
--+-----------------------------------------------------------------------------
--|     Function Name  : To_BitVector
--|
--|     Overloading    : 
--|
--|     Purpose        : Translate an INTEGER into a BIT_VECTOR.
--|
--|     Parameters     : intg    - input  INTEGER, the value to be translated.
--|                      width   - input  NATURAL, length of the return vector.
--|                            Default is IntegerBitLength (Machine integer length).
--|                      SrcRegMode - input  regmode_type, indicating the format of
--|                                the output BIT_VECTOR.   Default is TwosComp.
--|
--|     Result        : BIT_VECTOR, the binary representation of the integer.
--|
--|     NOTE           : An ASSERTION message of severity ERROR if the conversion
--|                      fails:
--|                       * 'intg' is negative and UnSigned format is specified.
--|                         The absolute value of 'intg' is used.
--|                       * The length of 'SrcReg' is insufficient to hold the
--|                         binary value. The low order bits are returned.
--|
--|                      A runtime system error should occur if the value of
--|                      'width' is does not equal the expected return vector
--|                      length (from the context of the function usage).
--|     Use            :
--|                      VARIABLE vect : BIT_VECTOR ( 15 DOWNTO 0 );
--|
--|                      vect := To_BitVector ( -294, 16, TwosComp );
--|
--|     See Also       : To_BitVector, To_Integer, To_TwosComp
--|-----------------------------------------------------------------------------
    FUNCTION To_BitVector ( CONSTANT intg       : IN INTEGER;
                            CONSTANT width      : IN Natural;
                            CONSTANT SrcRegMode : IN regmode_type  
                     -- synopsys synthesis_off
						      := DefaultRegMode 
                     -- synopsys synthesis_on
                          ) RETURN BIT_VECTOR;
--+-----------------------------------------------------------------------------
--|     Procedure Name : To_Integer
--|
--|     Overloading    : 
--|
--|     Purpose        : Interpret BIT_VECTOR as an INTEGER.
--|
--|     Parameters     :
--|                      SrcReg     - input  BIT_VECTOR, the vector to be read.
--|                      SrcRegMode - input  regmode_type, indicating the format of
--|                                the input BIT_VECTOR.   Default is TwosComp.
--|     NOTE           : 
--|                       * Magnitude of the computed integer is to large. The
--|                         input value is considered to large if after removing
--|                         leading 0's (1's for negative numbers) the length
--|                         of the remaining vector is > IntegerBitLength - 1.
--|                         (ie the machine integer length).
--|                      The error return value is INTEGER'LEFT.
--|     Use            :
--|                      VARIABLE vect : BIT_VECTOR ( 15 DOWNTO 0 );
--|
--|                      To_Integer ( vect, TwosComp );
--|
--|     See Also       : To_BitVector, To_Integer, To_TwosComp 
--|---------------------------------------------------------------------------------
     FUNCTION To_Integer  ( CONSTANT SrcReg     : IN BIT_VECTOR;
                            CONSTANT SrcRegMode : IN regmode_type  
                     -- synopsys synthesis_off
						      := DefaultRegMode 
                     -- synopsys synthesis_on
                          ) return INTEGER;
    -------------------------------------------------------------------------------
    --     Procedure Name : To_Integer
    --
    --     Overloading    : Procedure and Function.
    --    
    --     Purpose        : Interpret std_logic_vector as an INTEGER.
    --     
    --     Parameters     : 
    --                      SrcReg     - input  std_logic_vector, the vector to be 
    --                                          converted.
    --                      SrcRegMode - input  regmode_type, indicating the format 
    --                                    of the input std_logic_vector.   
    --                                    Default is DefaultRegMode.
    --     NOTE           : 
    --                      * Magnitude of the computed integer is to large. The 
    --                        input value is considered to large if after removing
    --                        leading 0's (1's for negative numbers)  the length
    --                        of the remaining vector is > IntegerBitLength-1.
    --                        (ie the machine integer length).
    --                        The error return value is INTEGER'LEFT.
    --     Use            : 
    --                      VARIABLE vect : std_logic_vector ( 15 DOWNTO 0 );
    --
    --                      To_Integer ( vect, TwosComp );
    --     
    --     See Also       :  To_Integer, To_TwosComp, To_OnesComp
    -------------------------------------------------------------------------------
    FUNCTION To_Integer   ( CONSTANT SrcReg     : IN std_logic_vector;
                            CONSTANT SrcRegMode : IN regmode_type  
                     -- synopsys synthesis_off
						      := DefaultRegMode 
                     -- synopsys synthesis_on
                          ) RETURN INTEGER;
    -------------------------------------------------------------------------------
    --     Procedure Name : To_Integer
    --
    --     Overloading    : Procedure and Function.
    --    
    --     Purpose        : Interpret std_ulogic_vector as an INTEGER.
    --     
    --     Parameters     : 
    --                      SrcReg     - input  std_ulogic_vector, the vector to be 
    --                                          converted.
    --                      SrcRegMode - input  regmode_type, indicating the format 
    --                                    of the input std_ulogic_vector.   
    --                                    Default is DefaultRegMode.
    --     NOTE           : 
    --                      * Magnitude of the computed integer is to large. The 
    --                        input value is considered to large if after removing
    --                        leading 0's (1's for negative numbers)  the length
    --                        of the remaining vector is > IntegerBitLength-1.
    --                        (ie the machine integer length).
    --                      The error return value is INTEGER'LEFT.
    --     Use            : 
    --                      VARIABLE vect : std_ulogic_vector ( 15 DOWNTO 0 );
    --
    --                      To_Integer ( vect, TwosComp );
    --     
    --     See Also       : To_StdLogicVector, To_Integer, To_TwosComp, To_OnesComp
    -------------------------------------------------------------------------------
    FUNCTION To_Integer   ( CONSTANT SrcReg     : IN std_ulogic_vector;
                            CONSTANT SrcRegMode : IN regmode_type  
                     -- synopsys synthesis_off
						      := DefaultRegMode 
                     -- synopsys synthesis_on
                          )  RETURN INTEGER;
    -------------------------------------------------------------------------------
    --     Procedure Name : RegAbs
    -- 1.6.9
    --     Overloading    : 
    --
    --     Purpose        : converts  std_logic_vector into an absolute value.
    --
    --     Parameters     :
    --                      result     - input-output  std_logic_vector, 
    --                      SrcReg     - input  std_logic_vector, the vector to be read.
    --                      SrcRegMode - input  regmode_type, indicating the format of
    --                              the input std_logic_vector.   Default is TwosComp.
    --
    --     Use            :
    --                      VARIABLE reslt, vect : std_logic_vector ( 15 DOWNTO 0 );
    --
    --                       RegAbs ( reslt,  vect, TwosComp );
    -------------------------------------------------------------------------------
    PROCEDURE RegAbs  ( VARIABLE result     : INOUT std_logic_vector;
                        CONSTANT SrcReg     : IN std_logic_vector;
                        CONSTANT SrcRegMode : IN regmode_type 
                     -- synopsys synthesis_off
						      := DefaultRegMode 
                     -- synopsys synthesis_on
                      );
    -------------------------------------------------------------------------------
    PROCEDURE RegAbs  ( VARIABLE result     : INOUT std_ulogic_vector;
                        CONSTANT SrcReg     : IN std_ulogic_vector;
                        CONSTANT SrcRegMode : IN regmode_type 
                     -- synopsys synthesis_off
						      := DefaultRegMode 
                     -- synopsys synthesis_on
                      );
    -------------------------------------------------------------------------------
    PROCEDURE RegAbs  ( VARIABLE result     : INOUT bit_vector;
                        CONSTANT SrcReg     : IN bit_vector;
                        CONSTANT SrcRegMode : IN regmode_type
                     -- synopsys synthesis_off
						      := DefaultRegMode 
                     -- synopsys synthesis_on
                      ) ;
--+-----------------------------------------------------------------------------
--|     Function Name  : RegAdd
--|
--|     Overloading    : None
--|
--|     Purpose        : Addition of logic vectors.
--|
--|     Parameters     :
--|                      result     - input/output  std_logic_vector,
--|                      carry_out  - OUT    std_ulogic,
--|                      overflow   - OUT    std_ulogic,
--|                      addend     - input  std_logic_vector,
--|                      augend     - input  std_logic_vector,
--|                      carry_in   - input  std_ulogic,
--|                      SrcRegMode - input  regmode_type, indicating the format of
--|                              the input std_logic_vector.   Default is TwosComp.
--|     NOTE           :
--|                      The inputs may be of any length and may be of differing
--|                      lengths.
--|  
--|                    For Synthesis:
--|                      Result is computed with length N (where
--|                      N is the greater of the input vector lengths).
--|                      It is assumed that user will provide result length equal
--|                      to the length of the greater of addend and augend. 
--|                      No error checking has been performed.
--|     Use            :
--|                      VARIABLE x, y, sum : std_logic_vector ( 15 DOWNTO 0);
--|                      VARIABLE carry_in, carry_out , ovf: std_ulogic;
--| 
--|                      RegAdd ( sum, carry_out, ovf,x, y, carry_in, TwosComp );
--| 
--|     See Also       : RegAdd, RegSub, RegMult, RegDiv, RegInc, RegDec, RegNegate
--|-----------------------------------------------------------------------------
    PROCEDURE RegAdd  ( VARIABLE result     : INOUT  std_logic_vector;
                        VARIABLE carry_out  : OUT std_ulogic;
                        VARIABLE overflow   : OUT std_ulogic;
                        CONSTANT addend     : IN std_logic_vector;
                        CONSTANT augend     : IN std_logic_vector;
                        CONSTANT carry_in   : IN std_ulogic;
                        CONSTANT SrcRegMode : IN regmode_type 
                     -- synopsys synthesis_off
						      := DefaultRegMode 
                     -- synopsys synthesis_on
                      ) ;
-------------------------------------------------------------------------------
    PROCEDURE RegAdd  ( VARIABLE result     : INOUT  std_ulogic_vector;
                        VARIABLE carry_out  : OUT std_ulogic;
                        VARIABLE overflow   : OUT std_ulogic;
                        CONSTANT addend     : IN std_ulogic_vector;
                        CONSTANT augend     : IN std_ulogic_vector;
                        CONSTANT carry_in   : IN std_ulogic;
                        CONSTANT SrcRegMode : IN regmode_type 
                     -- synopsys synthesis_off
						      := DefaultRegMode 
                     -- synopsys synthesis_on
                      ) ;
--------------------------------------------------------------------------------
    PROCEDURE RegAdd   (VARIABLE  result     : INOUT  BIT_VECTOR;
                        VARIABLE carry_out  : OUT BIT;
                        VARIABLE overflow   : OUT BIT;
                        CONSTANT addend     : IN BIT_VECTOR;
                        CONSTANT augend     : IN BIT_VECTOR;
                        CONSTANT carry_in   : IN BIT;
                        CONSTANT SrcRegMode : IN regmode_type 
                     -- synopsys synthesis_off
			                         := DefaultRegMode 
                     -- synopsys synthesis_on
                      );
--+-----------------------------------------------------------------------------
--|     Function Name  : RegSub
--|    
--|     Overloading    : None
--|
--|     Purpose        : Subtraction of BIT_VECTORS.
--|                       ( result = minuend - subtrahend )
--|
--|     Parameters     :
--|                      result     - input-output BIT_VECTOR, the computed sum
--|                      borrow_out - output BIT,
--|                      overflow   - output BIT, overflow condition
--|                      minuend - input  BIT_VECTOR,
--|                      subtrahend - input  BIT_VECTOR,
--|                      borrow_in  - input  BIT, borrow from the LSB
--|                      SrcRegMode - input  regmode_type, indicating the format of
--|                                the input BIT_VECTOR.   Default is TwosComp.
--|     NOTE           :
--|                      The inputs may be of any length and may be of differing
--|                      lengths.
--|
--|                      A temporary result is computed with length N (where
--|                      N is the greater of the input vector lengths).
--|     Use            :
--|                      VARIABLE x, y, diff : BIT_VECTOR ( 15 DOWNTO 0);
--|                      VARIABLE n_borrow, borrow_in : BIT;
--|
--|                      RegSub ( diff, n_borrow, x, y, borrow_in, UnSigned );
--|
--|     See Also       : RegAdd, RegSub, RegMult, RegDiv, RegInc, RegDec, RegNegate
--|-----------------------------------------------------------------------------
    PROCEDURE RegSub  ( VARIABLE result     : INOUT BIT_VECTOR;
                        VARIABLE borrow_out : OUT BIT;
                        VARIABLE overflow   : OUT BIT;
                        CONSTANT minuend    :  IN BIT_VECTOR;
                        CONSTANT subtrahend :  IN BIT_VECTOR;
                        CONSTANT borrow_in  :  IN BIT 
                     -- synopsys synthesis_off
                                                    := '0'
                     -- synopsys synthesis_on
                                                            ;
                        CONSTANT SrcRegMode :  IN regmode_type 
                     -- synopsys synthesis_off
						      := DefaultRegMode 
                     -- synopsys synthesis_on
                      );
--------------------------------------------------------------------------------
    PROCEDURE RegSub  ( VARIABLE result     : INOUT std_logic_vector;
                        VARIABLE borrow_out : OUT std_ulogic;
                        VARIABLE overflow   : OUT std_ulogic;
                        CONSTANT minuend    :  IN std_logic_vector;
                        CONSTANT subtrahend :  IN std_logic_vector;
                        CONSTANT borrow_in  :  IN std_ulogic  
                     -- synopsys synthesis_off
                                                    := '0'
                     -- synopsys synthesis_on
                                                            ;
                        CONSTANT SrcRegMode :  IN regmode_type 
                     -- synopsys synthesis_off
						      := DefaultRegMode 
                     -- synopsys synthesis_on
                      );
--------------------------------------------------------------------------------
    PROCEDURE RegSub  ( VARIABLE result     : INOUT std_ulogic_vector;
                        VARIABLE borrow_out : OUT std_ulogic;
                        VARIABLE overflow   : OUT std_ulogic;
                        CONSTANT minuend    :  IN std_ulogic_vector;
                        CONSTANT subtrahend :  IN std_ulogic_vector;
                        CONSTANT borrow_in  :  IN std_ulogic  
                     -- synopsys synthesis_off
                                                    := '0'
                     -- synopsys synthesis_on
                                                            ;
                        CONSTANT SrcRegMode :  IN regmode_type 
                     -- synopsys synthesis_off
						      := DefaultRegMode 
                     -- synopsys synthesis_on
                      );
--+-----------------------------------------------------------------------------
--|     Function Name  : RegMult
--|
--|     Overloading    : None
--|
--|     Purpose        : Multiplication of BIT_VECTORS.
--|
--|     Parameters     :
--|                      result       - output BIT_VECTOR, the computed product
--|                      overflow     - output BIT, overflow condition
--|                      multiplicand - input BIT_VECTOR,
--|                      multiplier   -  input BIT_VECTOR,
--|                      SrcRegMode   - input  regmode_type, indicating the format 
--|                                     of the input BIT_VECTOR.   Default is 
--|                                     DefaultRegMode which is set to TwosComp.
--|     NOTE           :
--|                      The inputs may be of any length and may be of differing
--|                      lengths.
--|
--|    Algorithm       : The multiplication is carried out as follows:
--|
--|                      1) Determine sign of result based on sign of 
--|                         multiploicand and sign  of multiplier.
--|
--|                      2) Convert the multiplicand amd multiplier to Unsigned 
--|                         representation.
--|                      
--|                      3) Perform multiplication based on add and shift algorithm.
--|
--|                      4) Convert the result to the SrcRegMode with appropropriate sign
--|     Result         :
--|                     A  temporary result is computed with length N+M (where
--|                      N,M are the lengths of the multiplicand and multiplier)
--|                      by calling local function Mult_TwosComp or Mult_Unsigned
--|                       
--|                      This computed value is extended or truncated to match
--|                      the width of 'result'. If truncated, the low order bits
--|                      are returned.
--|
--|                      The parameter 'overflow' is set to '1' if the product of the
--|                      two inputs is too large to fit in the parameter result.
--|     Use            :
--|                      VARIABLE x, y, prod : BIT_VECTOR ( 15 DOWNTO 0);
--|                      VARIABLE ovfl : BIT;
--|
--|                      RegMult ( prod, ovfl, x, y, TwosComp );
--|
--|     See Also       : RegAdd, RegSub, RegMult, RegDiv, RegInc, RegDec, RegNegate
--|-----------------------------------------------------------------------------
    PROCEDURE RegMult ( VARIABLE result       : OUT BIT_VECTOR;
                        VARIABLE overflow     : OUT BIT;
                        CONSTANT multiplicand : IN BIT_VECTOR;
                        CONSTANT multiplier   : IN BIT_VECTOR;
                        CONSTANT SrcRegMode   : IN regmode_type
                     -- synopsys synthesis_off
						      := DefaultRegMode 
                     -- synopsys synthesis_on
                      );
--------------------------------------------------------------------------------
    PROCEDURE RegMult ( VARIABLE result       : OUT STD_LOGIC_VECTOR;
                        VARIABLE overflow     : OUT STD_ULOGIC;
                        CONSTANT multiplicand : IN STD_LOGIC_VECTOR;
                        CONSTANT multiplier   : IN STD_LOGIC_VECTOR;
                        CONSTANT SrcRegMode   : IN regmode_type 
                     -- synopsys synthesis_off
						      := DefaultRegMode 
                     -- synopsys synthesis_on
                      );
--------------------------------------------------------------------------------
    PROCEDURE RegMult ( VARIABLE result       : OUT STD_ULOGIC_VECTOR;
                        VARIABLE overflow     : OUT STD_ULOGIC;
                        CONSTANT multiplicand : IN STD_ULOGIC_VECTOR;
                        CONSTANT multiplier   : IN STD_ULOGIC_VECTOR;
                        CONSTANT SrcRegMode   : IN regmode_type
                     -- synopsys synthesis_off
						      := DefaultRegMode 
                     -- synopsys synthesis_on
                      );
--+-----------------------------------------------------------------------------
--|     Function Name  : RegDiv
--|
--|     Overloading    : None
--|
--|     Purpose        : Division of BIT_VECTORS. (Result = dividend / divisor)
--|
--|     Parameters     :
--|                      result     - output BIT_VECTOR,
--|                      remainder  - output BIT_VECTOR,
--|                      ZeroDivide - output BIT,
--|                                   set to '1'  when divide by zero occurred
--|                                          '0'  divide by zero did not occur
--|                      dividend   - input  BIT_VECTOR,
--|                      divisor    - input  BIT_VECTOR,
--|                      SrcRegMode - input  regmode_type, indicating the format of
--|                                the input BIT_VECTOR.   Default is TwosComp.
--|     NOTE           :
--|                      The inputs may be of any length and may be of differing
--|                      lengths.
--|
--|                      For synthesis purposes result and remainder values are 
--|                      computed with  same length as the dividend. 
--|
--|                      The remainder has the same sign as the dividend.
--|     Use            :
--|                      VARIABLE x, y, res, rem : BIT_VECTOR ( 15 DOWNTO 0);
--|                      VARIABLE zflag     : BIT;
--|
--|                      RegDiv ( res, rem,zflag, x, y, TwosComp );
--|
--|     See Also       : RegAdd, RegSub, RegMult, RegDiv, RegInc, RegDec, RegNegate
--|-----------------------------------------------------------------------------
    PROCEDURE RegDiv  ( VARIABLE result     : OUT BIT_VECTOR;
                        VARIABLE remainder  : OUT BIT_VECTOR;
                        VARIABLE ZeroDivide : OUT BIT;
                        CONSTANT dividend   :  IN BIT_VECTOR;
                        CONSTANT divisor    :  IN BIT_VECTOR;
                        CONSTANT SrcRegMode    :  IN regmode_type
                     -- synopsys synthesis_off
						      := DefaultRegMode 
                     -- synopsys synthesis_on
                      ) ;
--------------------------------------------------------------------------------
    PROCEDURE RegDiv  ( VARIABLE result     : OUT STD_LOGIC_VECTOR;
                        VARIABLE remainder  : OUT STD_LOGIC_VECTOR;
                        VARIABLE ZeroDivide : OUT STD_ULOGIC;
                        CONSTANT dividend   :  IN STD_LOGIC_VECTOR;
                        CONSTANT divisor    :  IN STD_LOGIC_VECTOR;
                        CONSTANT SrcRegMode    :  IN regmode_type
                     -- synopsys synthesis_off
						      := DefaultRegMode 
                     -- synopsys synthesis_on
                      );
-------------------------------------------------------------------------------
    PROCEDURE RegDiv  ( VARIABLE result     : OUT STD_ULOGIC_VECTOR;
                        VARIABLE remainder  : OUT STD_ULOGIC_VECTOR;
                        VARIABLE ZeroDivide : OUT STD_ULOGIC;
                        CONSTANT dividend   :  IN STD_ULOGIC_VECTOR;
                        CONSTANT divisor    :  IN STD_ULOGIC_VECTOR;
                        CONSTANT SrcRegMode    :  IN regmode_type
                     -- synopsys synthesis_off
						      := DefaultRegMode 
                     -- synopsys synthesis_on
                      );
--+-----------------------------------------------------------------------------
--|     Function Name  : RegRem
--| 1.5.25
--|     Overloading    : None
--|
--|     Purpose        : Remainder operation of  BIT_VECTORS.
--|
--|     Parameters     :
--|                      result     - output BIT_VECTOR,
--|                      ZeroDivide - output BIT,
--|                                   set to '1'  when divide by zero occurred
--|                                          '0'  divide by zero did not occur
--|                      dividend   - input  BIT_VECTOR,
--|                      divisor    - input  BIT_VECTOR,
--|                      SrcRegMode - input  regmode_type, indicating the format of
--|                                the input BIT_VECTOR.   Default is TwosComp.
--|     NOTE           :
--|                      The inputs may be of any length and may be of differing
--|                      lengths.
--|
--|                      For synthesis purposes quotient and remainder values are 
--|                      computed with  same length as the dividend. 
--|
--|                      The remainder has the same sign as the dividend.
--|     Use            :
--|                      VARIABLE x, y, res : BIT_VECTOR ( 15 DOWNTO 0);
--|                      VARIABLE zflag     : BIT;
--|
--|                      RegRem ( res, zflag, x, y, TwosComp );
--|
--|     See Also       : RegAdd, RegSub, RegMult, RegDiv, RegInc, RegDec, RegNegate
--|-----------------------------------------------------------------------------
    PROCEDURE RegRem  ( VARIABLE result     : OUT BIT_VECTOR;
                        VARIABLE ZeroDivide : OUT BIT;
                        CONSTANT dividend   :  IN BIT_VECTOR;
                        CONSTANT divisor    :  IN BIT_VECTOR;
                        CONSTANT SrcRegMode :  IN regmode_type 
                     -- synopsys synthesis_off
						      := DefaultRegMode 
                     -- synopsys synthesis_on
                      );
--------------------------------------------------------------------------------
    PROCEDURE RegRem  ( VARIABLE result     : OUT STD_LOGIC_VECTOR;
                        VARIABLE ZeroDivide : OUT STD_ULOGIC;
                        CONSTANT dividend   :  IN STD_LOGIC_VECTOR;
                        CONSTANT divisor    :  IN STD_LOGIC_VECTOR;
                        CONSTANT SrcRegMode :  IN regmode_type
                     -- synopsys synthesis_off
						      := DefaultRegMode 
                     -- synopsys synthesis_on
                      );
--------------------------------------------------------------------------------
    PROCEDURE RegRem  ( VARIABLE result     : OUT STD_ULOGIC_VECTOR;
                        VARIABLE ZeroDivide : OUT STD_ULOGIC;
                        CONSTANT dividend   :  IN STD_ULOGIC_VECTOR;
                        CONSTANT divisor    :  IN STD_ULOGIC_VECTOR;
                        CONSTANT SrcRegMode :  IN regmode_type
                     -- synopsys synthesis_off
						      := DefaultRegMode 
                     -- synopsys synthesis_on
                      );
--+-----------------------------------------------------------------------------
--|     Function Name  : RegMod
--| 1.5.17  
--|     Overloading    : None
--| 
--|     Purpose        : Modulus operation of  STD_LOGIC_VECTORS.
--| 
--|     Parameters     :
--|                      result     - output STD_LOGIC_VECTOR,
--|                      ZeroDivide - output STD_ULOGIC,
--|                                   set to '1'  when divide by zero occurred
--|                                          '0'  divide by zero did not occur
--|                      dividend   - input  STD_LOGIC_VECTOR,
--|                      modulus    - input  STD_LOGIC_VECTOR,
--|                      SrcRegMode - input  regmode_type, indicating the format of
--|                                the input STD_LOGIC_VECTOR.   Default is TwosComp.
--|     NOTE           :
--|                      The inputs may be of any length and may be of differing
--|                      lengths.
--|
--|                      For synthesis purposes quotient and modulus values are 
--|                      computed with  same length as the dividend. 
--|
--|                      The mod has the same sign as the modulus operator.
--|     Use            :
--|                      VARIABLE x, y, res : STD_LOGIC_VECTOR ( 15 DOWNTO 0);
--|                      VARIABLE zflag     : STD_ULOGIC;
--|
--|                      RegMod ( res,zflag, x, y, TwosComp );
--|
--|     See Also       : RegAdd, RegSub, RegMult, RegDiv, RegInc, RegDec, RegNegate
--|-----------------------------------------------------------------------------
    PROCEDURE RegMod  ( VARIABLE result     : OUT STD_LOGIC_VECTOR;
                        VARIABLE ZeroDivide : OUT STD_ULOGIC;
                        CONSTANT dividend   : IN STD_LOGIC_VECTOR;
                        CONSTANT modulus    : IN STD_LOGIC_VECTOR;
                        CONSTANT SrcRegMode : IN regmode_type
                     -- synopsys synthesis_off
						      := DefaultRegMode 
                     -- synopsys synthesis_on
                      );
--------------------------------------------------------------------------------
    PROCEDURE RegMod  ( VARIABLE result     : OUT STD_ULOGIC_VECTOR;
                        VARIABLE ZeroDivide : OUT STD_ULOGIC;
                        CONSTANT dividend   : IN STD_ULOGIC_VECTOR;
                        CONSTANT modulus    : IN STD_ULOGIC_VECTOR;
                        CONSTANT SrcRegMode : IN regmode_type
                     -- synopsys synthesis_off
						      := DefaultRegMode 
                     -- synopsys synthesis_on
                      );
--------------------------------------------------------------------------------
    PROCEDURE RegMod  ( VARIABLE result     : OUT BIT_VECTOR;
                        VARIABLE ZeroDivide : OUT BIT;
                        CONSTANT dividend   : IN BIT_VECTOR;
                        CONSTANT modulus    : IN BIT_VECTOR;
                        CONSTANT SrcRegMode : IN regmode_type
                     -- synopsys synthesis_off
						      := DefaultRegMode 
                     -- synopsys synthesis_on
                      );
--+-----------------------------------------------------------------------------
--|     Function Name  : RegShift
--| 
--|     Overloading    : None
--|
--|     Purpose        : Bidirectional logical shift operator for   BIT_VECTORS.
--|
--|     Parameters     :
--|                      SrcReg      - input  BIT_VECTOR, vector to be shifted
--|                      DstReg      - Input_ouput, BIT_VECTOR, shifted result
--|                      ShiftO      - output, BIT, holds the last bit shifted out 
--|                                          of register
--|                      direction   - input, BIT
--|                                     '0'  means right shift
--|                                     '1'  means left shift, default is left shift
--|                      FillVal     - input, BIT, value to fill register with. 
--|                                          default is '0'.
--|                      Nbits       - input , NATURAL, number of positions to shift
--|                                          default is 1.
--|     NOTE           :
--|                      Default values are not allowed for synthesis.
--|
--|     Result         : Shifted bit_vector
--|
--|     Use            :
--|                      VARIABLE acc   : BIT_VECTOR ( 15 DOWNTO 0);
--|                      VARIABLE carry : BIT;
--|
--|                      RegShift ( acc, acc, carry, '1', '0',3 );
--|-----------------------------------------------------------------------------
   PROCEDURE RegShift  ( CONSTANT SrcReg    : IN BIT_VECTOR;
                         VARIABLE DstReg    : INOUT BIT_VECTOR;
                         VARIABLE ShiftO    : OUT BIT; 
                         CONSTANT direction : IN BIT     
                     -- synopsys synthesis_off
						      := '1'
                     -- synopsys synthesis_on
                                                            ;
                         CONSTANT FillVal   : IN BIT  
                     -- synopsys synthesis_off
						      := '0'
                     -- synopsys synthesis_on
                                                            ;
                         CONSTANT Nbits     : IN Natural
                     -- synopsys synthesis_off
						       := 1 
                     -- synopsys synthesis_on
                      ) ;
-------------------------------------------------------------------------------
   PROCEDURE RegShift  ( CONSTANT SrcReg    : IN std_logic_vector;
                         VARIABLE DstReg    : INOUT std_logic_vector;
                         VARIABLE ShiftO    : OUT std_ulogic; 
                         CONSTANT direction : IN std_ulogic
                     -- synopsys synthesis_off
						      := '1'
                     -- synopsys synthesis_on
                                                            ;
                         CONSTANT FillVal   : IN std_ulogic  
                     -- synopsys synthesis_off
						      := '0'
                     -- synopsys synthesis_on
                                                            ;
                         CONSTANT Nbits     : IN Natural
                     -- synopsys synthesis_off
						       := 1 
                     -- synopsys synthesis_on
                      );
-------------------------------------------------------------------------------
   PROCEDURE RegShift  ( CONSTANT SrcReg    : IN std_ulogic_vector;
                         VARIABLE DstReg    : INOUT std_ulogic_vector;
                         VARIABLE ShiftO    : OUT std_ulogic; 
                         CONSTANT direction : IN std_ulogic
                     -- synopsys synthesis_off
						      := '1'
                     -- synopsys synthesis_on
                                                            ;
                         CONSTANT FillVal   : IN std_ulogic  
                     -- synopsys synthesis_off
						      := '0'
                     -- synopsys synthesis_on
                                                            ;
                         CONSTANT Nbits     : IN Natural
                     -- synopsys synthesis_off
						       := 1 
                     -- synopsys synthesis_on
                      );
--+-----------------------------------------------------------------------------
--|     Function Name  : RegInc
--| 
--|     Overloading    : None
--|  
--|     Purpose        : Increment a BIT_VECTOR by 1.
--|  
--|     Parameters     :
--|                      SrcReg     - input  BIT_VECTOR
--|                      SrcRegMode - input  regmode_type, indicating the format of
--|                                the input BIT_VECTOR.   Default is TwosComp.
--|  
--|     Result         : BIT_VECTOR ( SrcReg + 1 )
--| 
--|     NOTE           : The length of the return vector is the same as the
--|                      the input vector.
--|  
--|                      Overflow conditions are ignored. UnSigned numbers wrap
--|                      to 0, signed numbers wrap to the largest negative value.
--|     Use            :
--|                      VARIABLE vect : BIT_VECTOR ( 3 DOWNTO 0 );
--|                      vect := RegInc ( vect, UnSigned )
--| 
--|     See Also       : RegAdd, RegSub, RegMult, RegDiv, RegInc, RegDec, RegNegate
--|-----------------------------------------------------------------------------
    FUNCTION RegInc  ( CONSTANT SrcReg        :  IN BIT_VECTOR;
                       CONSTANT SrcRegMode    :  IN regmode_type
                     -- synopsys synthesis_off
						      := DefaultRegMode 
                     -- synopsys synthesis_on
                     ) RETURN BIT_VECTOR;
    -------------------------------------------------------------------------------
    FUNCTION  RegInc  ( CONSTANT SrcReg        :  IN std_logic_vector;
                        CONSTANT SrcRegMode    :  IN regmode_type
                     -- synopsys synthesis_off
						      := DefaultRegMode 
                     -- synopsys synthesis_on
                      ) RETURN std_logic_vector;
    -------------------------------------------------------------------------------
    FUNCTION  RegInc  ( CONSTANT SrcReg        :  IN std_ulogic_vector;
                        CONSTANT SrcRegMode    :  IN regmode_type 
                     -- synopsys synthesis_off
						      := DefaultRegMode 
                     -- synopsys synthesis_on
                      ) RETURN std_ulogic_vector;
--+-----------------------------------------------------------------------------
--|     Function Name  : RegDec
--|
--|     Overloading    : None
--| 
--|     Purpose        : Decrement a BIT_VECTOR by 1.
--| 
--|     Parameters     :
--|                      SrcReg     - input  BIT_VECTOR
--|                      SrcRegMode - input  regmode_type, indicating the format of
--|                                the input BIT_VECTOR.   Default is TwosComp.
--| 
--|     Result         : BIT_VECTOR ( SrcReg - 1 )
--|
--|     NOTE           : The length of the return vector is the same as the
--|                      the input vector.
--|     Use            :
--|                      VARIABLE vect : BIT_VECTOR ( 3 DOWNTO 0 );
--|                      vect := RegDec ( vect, UnSigned )
--| 
--|     See Also       : RegAdd, RegSub, RegMult, RegDiv, RegInc, RegDec, RegNegate
--|-----------------------------------------------------------------------------
    FUNCTION RegDec  ( CONSTANT SrcReg        :  IN BIT_VECTOR;
                       CONSTANT SrcRegMode    :  IN regmode_type 
                     -- synopsys synthesis_off
						      := DefaultRegMode 
                     -- synopsys synthesis_on
                     ) RETURN BIT_VECTOR;
    -------------------------------------------------------------------------------
    FUNCTION  RegDec  ( CONSTANT SrcReg        :  IN std_logic_vector;
                        CONSTANT SrcRegMode    :  IN regmode_type 
                     -- synopsys synthesis_off
						      := DefaultRegMode 
                     -- synopsys synthesis_on
                      ) RETURN std_logic_vector;
    -------------------------------------------------------------------------------
    FUNCTION  RegDec  ( CONSTANT SrcReg        :  IN std_ulogic_vector;
                        CONSTANT SrcRegMode    :  IN regmode_type 
                     -- synopsys synthesis_off
						      := DefaultRegMode 
                     -- synopsys synthesis_on
                      ) RETURN std_ulogic_vector;
--+-----------------------------------------------------------------------------
--|     Function Name  : RegNegate
--|
--|     Overloading    : None
--|
--|     Purpose        : Negate a BIT_VECTOR ( v := 0 - v )
--|
--|     Parameters     :
--|                      SrcReg     - input  BIT_VECTOR
--|                      SrcRegMode - input  regmode_type, indicating the format of
--|                                the input BIT_VECTOR.   Default is TwosComp.
--|
--|     Result         : BIT_VECTOR ( 0 - SrcReg )
--|
--|     NOTE           : The length of the return vector is the same as the
--|                      the input vector.
--|
--|                      If 'SrcRegMode' is UnSigned the bitwise NOT of 'SrcReg'
--|                      is returned.
--|
--|                      An overflow can occur when 'SrcRegMode' is TwosComp and
--|                      'SrcReg' is the largest negative value (ie "100...00").
--|                      In this case NO error is indicated and the returned
--|                      value is the same as the input.
--|     Use            :
--|                      VARIABLE vect : BIT_VECTOR (15 DOWNTO 0 );
--|                      vect := RegNegate ( vect, TwosComp );
--|
--|     See Also       : RegAdd, RegSub, RegMult, RegDiv, RegInc, RegDec, RegNegate
--|-----------------------------------------------------------------------------
    FUNCTION RegNegate  ( CONSTANT SrcReg      :  IN BIT_VECTOR;
                          CONSTANT SrcRegMode  :  IN regmode_type 
                 -- synopsys synthesis_off
                                                     := DefaultRegMode
                 -- synopsys synthesis_on
                        ) RETURN BIT_VECTOR;
    -------------------------------------------------------------------------------
    FUNCTION  RegNegate  ( CONSTANT SrcReg     :  IN std_logic_vector;
                           CONSTANT SrcRegMode :  IN regmode_type
                 -- synopsys synthesis_off
                                                     := DefaultRegMode
                 -- synopsys synthesis_on
                         ) RETURN std_logic_vector;
    -------------------------------------------------------------------------------
    FUNCTION  RegNegate  ( CONSTANT SrcReg     :  IN std_ulogic_vector;
                           CONSTANT SrcRegMode :  IN regmode_type
                 -- synopsys synthesis_off
                                                     := DefaultRegMode
                 -- synopsys synthesis_on
                         ) RETURN std_ulogic_vector;
    -------------------------------------------------------------------------------
    --     Function Name  : RegFill
    -- 1.7.4
    --     Overloading    : None
    --
    --     Purpose        : Fill an std_logic_vector with a given value
    --
    --     Parameters     :
    --                      SrcReg     - input  std_logic_vector, the  logic vector to be read.
    --                      DstLength  - input  NATURAL, length of the return logic vector.
    --                      FillVal    - input  std_ulogic, default is '0'
    --
    --     Result         : std_logic_vector of length DstLength
    --
    --     NOTE           : The length of the return logic vector  is specified by the
    --                      parameter 'DstLength'. The input logic vector will
    --                      be  filled with the FillVal
    --
    --     Use            :
    --                      VARIABLE vect : std_logic_vector ( 15 DOWNTO 0 );
    --                      vect := RegFill ( "00000101", 16, 'U');
    --
    --     See Also       : SignExtend
   -------------------------------------------------------------------------------
    FUNCTION RegFill   ( CONSTANT SrcReg      : IN std_logic_vector;
                         CONSTANT DstLength   : IN NATURAL;
                         CONSTANT FillVal     : IN std_ulogic
        	-- synopsys synthesis_off
					         := '0'
	        -- synopsys synthesis_on
                       ) RETURN std_logic_vector;
   -------------------------------------------------------------------------------
    FUNCTION RegFill   ( CONSTANT SrcReg      : IN std_ulogic_vector;
                         CONSTANT DstLength   : IN NATURAL;
                         CONSTANT FillVal     : IN std_ulogic
        	-- synopsys synthesis_off
					         := '0'
	        -- synopsys synthesis_on
                       ) RETURN std_ulogic_vector;
   -------------------------------------------------------------------------------
    FUNCTION RegFill   ( CONSTANT SrcReg      : IN bit_vector;
                         CONSTANT DstLength   : IN NATURAL;
                         CONSTANT FillVal     : IN bit  
        	-- synopsys synthesis_off
					         := '0'
	        -- synopsys synthesis_on

                       ) RETURN bit_vector;
    -------------------------------------------------------------------------------
    --     Function Name  : SignExtend
    -- 1.7.1
    --     Overloading    : None
    --    
    --     Purpose        : Sign Extend a logic vector
    --     
    --     Parameters     : 
    --                      SrcReg     - input  std_logic_vector, the vector to be read.
    --                      DstLength  - input  NATURAL, length of the return vector.
    --                      SignBitPos - input  NATURAL, the position of the sign bit.
    --                                    for synthesis purpose it is the MSB (SrcReg'LEFT)

    --                      SrcRegMode  - input regmode_type, indicating the format of
    --                                 the input std_logic_vector.Default is TwosComp.
    --     
    --     Result         : std_logic_vector
    --
    --     NOTE           : The length of the return std_logic_vector is specified by 
    --                      the parameter 'DstLength'. The input std_logic_vector 
    --                      will be sign extended. 
    --
    --                     For synthesis purpose SignBitPos argument is ignored and the  
    --                     the MSB (ie. SrcReg'Left) is considered as a sign bit position.
    --     Use            :
    --                      VARIABLE vect : std_logic_vector ( 15 DOWNTO 0 );
    --                      vect := SignExtend ( "11111101", 16, 7, TwosComp ); -- set to -4
    --
    --     See Also       : RegFill
    -------------------------------------------------------------------------------
    FUNCTION SignExtend   ( CONSTANT SrcReg      : IN std_logic_vector;
                            CONSTANT DstLength   : IN NATURAL;
                            CONSTANT SignBitPos  : IN NATURAL;
                            CONSTANT SrcRegMode  : IN regmode_type 
                     -- synopsys synthesis_off
						      := DefaultRegMode 
                     -- synopsys synthesis_on
                          ) RETURN std_logic_vector;
    -------------------------------------------------------------------------------
    FUNCTION SignExtend   ( CONSTANT SrcReg      : IN std_ulogic_vector;
                            CONSTANT DstLength   : IN NATURAL;
                            CONSTANT SignBitPos  : IN NATURAL;
                            CONSTANT SrcRegMode  : IN regmode_type 
                     -- synopsys synthesis_off
						      := DefaultRegMode 
                     -- synopsys synthesis_on
                          ) RETURN std_ulogic_vector;
    -------------------------------------------------------------------------------
    FUNCTION SignExtend   ( CONSTANT SrcReg      : IN bit_vector;
                            CONSTANT DstLength   : IN NATURAL;
                            CONSTANT SignBitPos  : IN NATURAL;
                            CONSTANT SrcRegMode  : IN regmode_type 
                     -- synopsys synthesis_off
						      := DefaultRegMode 
                     -- synopsys synthesis_on
                          ) RETURN bit_vector;
    -------------------------------------------------------------------------------
    --     Procedure Name : SregAbs
    -- 1.6.9
    --     Overloading    : Procedure .
    --
    --     Purpose        : converts  std_logic_vector into an absolute value.
    --
    --     Parameters     :
    --                      result     - input-output  std_logic_vector, 
    --                      SrcReg     - input  std_logic_vector, the vector to be read.
    --                      SrcRegMode - input  regmode_type, indicating the format of
    --                             the input std_logic_vector.   Default is TwosComp.
    --
    --     Use            :
    --                      SIGNAL reslt, vect : std_logic_vector ( 15 DOWNTO 0 );
    --
    --                       SregAbs ( reslt,  vect, TwosComp );
    -------------------------------------------------------------------------------
    PROCEDURE SregAbs  ( SIGNAL result     : INOUT std_logic_vector;
                        CONSTANT SrcReg     : IN std_logic_vector;
                        CONSTANT SrcRegMode : IN regmode_type 
                     -- synopsys synthesis_off
						      := DefaultRegMode 
                     -- synopsys synthesis_on
                      );
    -------------------------------------------------------------------------------
    PROCEDURE SregAbs  ( SIGNAL result     : INOUT std_ulogic_vector;
                        CONSTANT SrcReg     : IN std_ulogic_vector;
                        CONSTANT SrcRegMode : IN regmode_type 
                     -- synopsys synthesis_off
						      := DefaultRegMode 
                     -- synopsys synthesis_on
                      );
    -------------------------------------------------------------------------------
    PROCEDURE SregAbs  ( SIGNAL result     : INOUT bit_vector;
                        CONSTANT SrcReg     : IN bit_vector;
                        CONSTANT SrcRegMode : IN regmode_type 
                     -- synopsys synthesis_off
						      := DefaultRegMode 
                     -- synopsys synthesis_on
                      );
--+-----------------------------------------------------------------------------
--|     Function Name  : SregAdd
--|
--|     Overloading    : None
--|
--|     Purpose        : Addition of STD_LOGIC_VECTORS.
--|
--|     Parameters     :
--|                      result     - input-output STD_LOGIC_VECTOR, the computed sum
--|                      carry_out  - output STD_ULOGIC,
--|                      overflow   - output STD_ULOGIC, overflow condition
--|                      addend     - input  STD_LOGIC_VECTOR,
--|                      augend     - input  STD_LOGIC_VECTOR,
--|                      carry_in   - input  STD_ULOGIC,  
--|                      SrcRegMode - input  regmode_type, indicating the format of
--|                                the input STD_LOGIC_VECTOR.   Default is TwosComp.
--|
--|     NOTE           :
--|                      The inputs may be of any length and may be of differing
--|                      lengths.
--|                    
--|                    For Synthesis:
--|                      Result is computed with length N (where
--|                      N is the greater of the input vector lengths).
--|                      It is assumed that user will provide result length equal
--|                      to the length of the greater of addend and augend. 
--|                      No error checking has been performed.
--|     Use            :
--|                      SIGNAL x, y, sum : STD_LOGIC_VECTOR ( 15 DOWNTO 0);
--|                      SIGNAL carry_in, carry_out , ovf: STD_ULOGIC;
--| 
--|                      SregAdd ( sum, carry_out, ovf,x, y, carry_in, UnSigned );
--| 
--|     See Also       : SregSub, SregMult, SregDiv
--|-----------------------------------------------------------------------------
    PROCEDURE SregAdd  (SIGNAL result       : INOUT STD_LOGIC_VECTOR;
                        SIGNAL carry_out    : OUT STD_ULOGIC;
                        SIGNAL overflow     : OUT STD_ULOGIC;
                        CONSTANT addend     : IN STD_LOGIC_VECTOR;
                        CONSTANT augend     : IN STD_LOGIC_VECTOR;
                        CONSTANT carry_in   : IN STD_ULOGIC;
                        CONSTANT SrcRegMode : IN regmode_type 
                  -- synopsys synthesis_off
                                                       := DefaultRegMode 
                   -- synopsys synthesis_on
                      );
--------------------------------------------------------------------------------
    PROCEDURE SregAdd  (SIGNAL result       : INOUT STD_ULOGIC_VECTOR;
                        SIGNAL carry_out    : OUT STD_ULOGIC;
                        SIGNAL overflow     : OUT STD_ULOGIC;
                        CONSTANT addend     : IN STD_ULOGIC_VECTOR;
                        CONSTANT augend     : IN STD_ULOGIC_VECTOR;
                        CONSTANT carry_in   : IN STD_ULOGIC;
                        CONSTANT SrcRegMode : IN regmode_type
                  -- synopsys synthesis_off
                                                       := DefaultRegMode 
                   -- synopsys synthesis_on
                      ) ;
--------------------------------------------------------------------------------
    PROCEDURE SregAdd  (SIGNAL result       : INOUT BIT_VECTOR;
                        SIGNAL carry_out    : OUT BIT;
                        SIGNAL overflow     : OUT BIT;
                        CONSTANT addend     : IN BIT_VECTOR;
                        CONSTANT augend     : IN BIT_VECTOR;
                        CONSTANT carry_in   : IN BIT;
                        CONSTANT SrcRegMode : IN regmode_type 
                  -- synopsys synthesis_off
                                                       := DefaultRegMode 
                   -- synopsys synthesis_on
                      );
--+-----------------------------------------------------------------------------
--|     Function Name  : SregSub
--|    
--|     Overloading    : None
--|
--|     Purpose        : Subtraction of STD_LOGIC_VECTORS.
--|                       ( result = minuend - subtrahend )
--|
--|     Parameters     :
--|                      result     - input-output STD_LOGIC_VECTOR, the computed sum
--|                      borrow_out - output STD_ULOGIC,
--|                      overflow   - output STD_ULOGIC, overflow condition
--|                      minuend - input  STD_LOGIC_VECTOR,
--|                      subtrahend - input  STD_LOGIC_VECTOR,
--|                      borrow_in  - input  STD_LOGIC, borrow from the LSB
--|                      SrcRegMode - input  regmode_type, indicating the format of
--|                                the input STD_LOGIC_VECTOR.   Default is TwosComp.
--|     NOTE           :
--|                      The inputs may be of any length and may be of differing
--|                      lengths.
--|
--|                      A  result is computed with length N (where
--|                      N is the greater of the input vector lengths).
--|     Use            :
--|                      SIGNAL x, y, diff : STD_LOGIC_VECTOR ( 15 DOWNTO 0);
--|                      SIGNAL n_borrow, borrow_in : STD_ULOGIC;
--|
--|                      SregSub ( diff, n_borrow, x, y, borrow_in, UnSigned );
--|
--|     See Also       : SregAdd,  SregMult, SregDiv
--|-----------------------------------------------------------------------------
    PROCEDURE SregSub  (SIGNAL result       : INOUT STD_LOGIC_VECTOR;
                        SIGNAL borrow_out   : OUT STD_ULOGIC;
                        SIGNAL overflow     : OUT STD_ULOGIC;
                        CONSTANT minuend    :  IN STD_LOGIC_VECTOR;
                        CONSTANT subtrahend :  IN STD_LOGIC_VECTOR;
                        CONSTANT borrow_in  :  IN STD_ULOGIC  
                  -- synopsys synthesis_off
                                                       := '0'
                  -- synopsys synthesis_on
                                                               ;
                        CONSTANT SrcRegMode :  IN regmode_type
                  -- synopsys synthesis_off
                                                       := DefaultRegMode 
                   -- synopsys synthesis_on
                      );
--------------------------------------------------------------------------------
    PROCEDURE SregSub  (SIGNAL result       : INOUT STD_ULOGIC_VECTOR;
                        SIGNAL borrow_out   : OUT STD_ULOGIC;
                        SIGNAL overflow     : OUT STD_ULOGIC;
                        CONSTANT minuend    :  IN STD_ULOGIC_VECTOR;
                        CONSTANT subtrahend :  IN STD_ULOGIC_VECTOR;
                        CONSTANT borrow_in  :  IN STD_ULOGIC  
                  -- synopsys synthesis_off
                                                       := '0'
                  -- synopsys synthesis_on
                                                               ;
                        CONSTANT SrcRegMode :  IN regmode_type
                  -- synopsys synthesis_off
                                                       := DefaultRegMode 
                   -- synopsys synthesis_on
                      );
--------------------------------------------------------------------------------
    PROCEDURE SregSub  (SIGNAL result       : INOUT BIT_VECTOR;
                        SIGNAL borrow_out   : OUT BIT;
                        SIGNAL overflow     : OUT BIT;
                        CONSTANT minuend    :  IN BIT_VECTOR;
                        CONSTANT subtrahend :  IN BIT_VECTOR;
                        CONSTANT borrow_in  :  IN BIT  
                  -- synopsys synthesis_off
                                                       := '0'
                  -- synopsys synthesis_on
                                                               ;
                        CONSTANT SrcRegMode :  IN regmode_type
                   -- synopsys synthesis_off
                                                       := DefaultRegMode 
                   -- synopsys synthesis_on
                        );
--+-----------------------------------------------------------------------------
--|     Function Name  : SregMult
--|
--|     Overloading    : None
--|
--|     Purpose        : Multiplication of STD_LOGIC_VECTORS.
--|
--|     Parameters     :
--|                      result       - output STD_LOGIC_VECTOR, the computed product
--|                      overflow     - output STD_ULOGIC, overflow condition
--|                      multiplicand - input STD_LOGIC_VECTOR,
--|                      multiplier   -  input STD_LOGIC_VECTOR,
--|                      SrcRegMode   - input  regmode_type, indicating the format 
--|                                     of the input STD_LOGIC_VECTOR.   Default is 
--|                                     DefaultRegMode which is set to TwosComp.
--|     NOTE           :
--|                      The inputs may be of any length and may be of differing
--|                      lengths.
--|
--|    Algorithm       : The multiplication is carried out as follows:
--|
--|                      1) Determine sign of result based on sign of 
--|                         multiploicand and sign  of multiplier.
--|
--|                      2) Convert the multiplicand amd multiplier to Unsigned 
--|                         representation.
--|                      
--|                      3) Perform multiplication based on add and shift algorithm.
--|
--|                      4) Convert the result to the SrcRegMode with appropropriate sign
--|
--|     Result         :
--|                     A  temporary result is computed with length N+M (where
--|                      N,M are the lengths of the multiplicand and multiplier).
--|                      This computed value is extended or truncated to match
--|                      the width of 'result'. If truncated, the low order std_ulogics
--|                      are returned.
--|
--|                      The parameter 'overflow' is set to '1' if the product of the
--|                      of the two inputs too large to fit in the parameter result.
--|     Use            :
--|                      SIGNAL x, y, prod : STD_LOGIC_VECTOR ( 15 DOWNTO 0);
--|                      SIGNAL ovfl : STD_ULOGIC;
--|
--|                      SregMult ( prod, ovfl, x, y, TwosComp );
--|
--|     See Also       : RegAdd, SregSub, SregMult, RegDiv, RegInc, RegDec, RegNegate
--|-----------------------------------------------------------------------------
    PROCEDURE SregMult (SIGNAL result         : OUT STD_LOGIC_VECTOR;
                        SIGNAL overflow       : OUT STD_ULOGIC;
                        CONSTANT multiplicand : IN STD_LOGIC_VECTOR;
                        CONSTANT multiplier   : IN STD_LOGIC_VECTOR;
                        CONSTANT SrcRegMode   : IN regmode_type 
                  -- synopsys synthesis_off
                                                       := DefaultRegMode 
                   -- synopsys synthesis_on
                      );
--------------------------------------------------------------------------------
    PROCEDURE SregMult (SIGNAL result         : OUT STD_ULOGIC_VECTOR;
                        SIGNAL overflow       : OUT STD_ULOGIC;
                        CONSTANT multiplicand : IN STD_ULOGIC_VECTOR;
                        CONSTANT multiplier   : IN STD_ULOGIC_VECTOR;
                        CONSTANT SrcRegMode   : IN regmode_type 
                  -- synopsys synthesis_off
                                                       := DefaultRegMode 
                   -- synopsys synthesis_on
                      );
--------------------------------------------------------------------------------
    PROCEDURE SregMult (SIGNAL result         : OUT BIT_VECTOR;
                        SIGNAL overflow       : OUT BIT;
                        CONSTANT multiplicand : IN BIT_VECTOR;
                        CONSTANT multiplier   : IN BIT_VECTOR;
                        CONSTANT SrcRegMode   : IN regmode_type 
                  -- synopsys synthesis_off
                                                       := DefaultRegMode 
                   -- synopsys synthesis_on
                      );
    -------------------------------------------------------------------------------
    --     Function Name  : SregDiv
    --
    --     Overloading    : None
    --    
    --     Purpose        : Division of std_logic_vectors.(Result = dividend/divisor)
    --     
    --     Parameters     : 
    --                      result     - output std_logic_vector, 
    --                      remainder  - output std_logic_vector,
    --                      ZeroDivide - output std_ulogic,
    --                                   set to '1' when  divide by zero occurred
    --                                          '0'  divide by zero did not occur  
    --                      dividend   - input  std_logic_vector, 
    --                      divisor    - input  std_logic_vector, 
    --                      SrcRegMode - input  regmode_type, indicating the format 
    --                                   of  the input std_logic_vector.   
    --                                   Default is TwosComp.
    --     NOTE           : 
    --                      The inputs may be of any length and may be of differing 
    --                      lengths. 
    --
    --                      For synthesis purposes result and remainder values are 
    --                      computed with  same length as the dividend. 
    --                      The remainder has the same sign as the dividend.
    --     Use            : 
    --                      SIGNAL x, y, res, rem : std_logic_vector ( 15 DOWNTO 0);
    --                      SIGNAL Zflag : std_ulogic;
    --
    --                      SregDiv ( res, rem, Zflag, x, y, TwosComp );
    --     
    --     See Also       : SregAdd, SregSub, SregMult, SregMod, SregRem
    -------------------------------------------------------------------------------
    PROCEDURE SregDiv ( SIGNAL result       : OUT std_logic_vector;
                        SIGNAL remainder    : OUT std_logic_vector;
                        SIGNAL ZeroDivide   : OUT std_ulogic;  
                        CONSTANT dividend   :  IN std_logic_vector;
                        CONSTANT divisor    :  IN std_logic_vector;
                        CONSTANT SrcRegMode :  IN regmode_type
                  -- synopsys synthesis_off
                                                       := DefaultRegMode 
                  -- synopsys synthesis_on
                      );
    -------------------------------------------------------------------------------
    PROCEDURE SregDiv ( SIGNAL result       : OUT std_ulogic_vector;
                        SIGNAL remainder    : OUT std_ulogic_vector;
                        SIGNAL ZeroDivide   : OUT std_ulogic;  
                        CONSTANT dividend   :  IN std_ulogic_vector;
                        CONSTANT divisor    :  IN std_ulogic_vector;
                        CONSTANT SrcRegMode :  IN regmode_type
                  -- synopsys synthesis_off
                                                       := DefaultRegMode 
                  -- synopsys synthesis_on
                      );
    -----------------------------------------------------------------------------
    PROCEDURE SregDiv ( SIGNAL result       : OUT BIT_VECTOR;
                        SIGNAL remainder    : OUT BIT_VECTOR;
                        SIGNAL ZeroDivide   : OUT BIT;
                        CONSTANT dividend   :  IN BIT_VECTOR;
                        CONSTANT divisor    :  IN BIT_VECTOR;
                        CONSTANT SrcRegMode :  IN regmode_type 
                  -- synopsys synthesis_off
                                                       := DefaultRegMode 
                   -- synopsys synthesis_on
                      );
--+-----------------------------------------------------------------------------
--|     Function Name  : SregMod
--| 1.5.17  
--|     Overloading    : None
--| 
--|     Purpose        : Modulus operation of  STD_LOGIC_VECTORS.
--| 
--|     Parameters     :
--|                      result     - output STD_LOGIC_VECTOR,
--|                      ZeroDivide - output STD_ULOGIC,
--|                                   set to '1'  when divide by zero occurred
--|                                          '0'  divide by zero did not occur
--|                      dividend   - input  STD_LOGIC_VECTOR,
--|                      modulus    - input  STD_LOGIC_VECTOR,
--|                      SrcRegMode - input  regmode_type, indicating the format of
--|                                the input STD_LOGIC_VECTOR.   Default is TwosComp.
--|     NOTE           :
--|                      The inputs may be of any length and may be of differing
--|                      lengths.
--|
--|                      For synthesis purposes quotient and modulus values are 
--|                      computed with  same length as the dividend. 
--|
--|                      The mod has the same sign as the modulus operator.
--|     Use            :
--|                      SIGNAL x, y, res : STD_LOGIC_VECTOR ( 15 DOWNTO 0);
--|                      SIGNAL zflag     : STD_ULOGIC;
--|
--|                      SregMod ( res,zflag, x, y, TwosComp );
--|-----------------------------------------------------------------------------
    PROCEDURE SregMod  ( SIGNAL result     : OUT STD_LOGIC_VECTOR;
                        SIGNAL ZeroDivide : OUT STD_ULOGIC;
                        CONSTANT dividend   : IN STD_LOGIC_VECTOR;
                        CONSTANT modulus    : IN STD_LOGIC_VECTOR;
                        CONSTANT SrcRegMode : IN regmode_type
                     -- synopsys synthesis_off
						      := DefaultRegMode 
                     -- synopsys synthesis_on
                      );
-------------------------------------------------------------------------------
    PROCEDURE SregMod  ( SIGNAL result     : OUT STD_ULOGIC_VECTOR;
                         SIGNAL ZeroDivide : OUT STD_ULOGIC;
                         CONSTANT dividend   : IN STD_ULOGIC_VECTOR;
                         CONSTANT modulus    : IN STD_ULOGIC_VECTOR;
                         CONSTANT SrcRegMode : IN regmode_type
                     -- synopsys synthesis_off
						      := DefaultRegMode 
                     -- synopsys synthesis_on
                      );
--- -----------------------------------------------------------------------------
    PROCEDURE SregMod  ( SIGNAL result     : OUT BIT_VECTOR;
                        SIGNAL ZeroDivide : OUT BIT;
                        CONSTANT dividend   : IN BIT_VECTOR;
                        CONSTANT modulus    : IN BIT_VECTOR;
                        CONSTANT SrcRegMode : IN regmode_type
                     -- synopsys synthesis_off
						      := DefaultRegMode 
                     -- synopsys synthesis_on
                      ) ;
--+-----------------------------------------------------------------------------
--|     Function Name  : SregRem
--| 1.5.25
--|     Overloading    : None
--|
--|     Purpose        : Remainder operation of  STD_LOGIC_VECTORS.
--|
--|     Parameters     :
--|                      result     - output STD_LOGIC_VECTOR,
--|                      ZeroDivide - output STD_ULOGIC,
--|                                   set to '1'  when divide by zero occurred
--|                                          '0'  divide by zero did not occur
--|                      dividend   - input  STD_LOGIC_VECTOR,
--|                      divisor    - input  STD_LOGIC_VECTOR,
--|                      SrcRegMode - input  regmode_type, indicating the format of
--|                                the input STD_LOGIC_VECTOR.   Default is TwosComp.
--|     NOTE           :
--|                      The inputs may be of any length and may be of differing
--|                      lengths.
--|
--|                      For synthesis purposes quotient and remainder values are 
--|                      computed with  same length as the dividend. 
--|
--|                      The remainder has the same sign as the dividend.
--|     Use            :
--|                      SIGNAL x, y, res : STD_LOGIC_VECTOR ( 15 DOWNTO 0);
--|                      SIGNAL zflag     : STD_ULOGIC;
--|
--|                      SregRem ( res, zflag, x, y, TwosComp );
--|
--|     See Also       : SeegAdd, SregSub, SregMult, SregDiv
--|-----------------------------------------------------------------------------
    PROCEDURE SregRem ( SIGNAL result       : OUT STD_LOGIC_VECTOR;
                        SIGNAL ZeroDivide   : OUT STD_ULOGIC;
                        CONSTANT dividend   :  IN STD_LOGIC_VECTOR;
                        CONSTANT divisor    :  IN STD_LOGIC_VECTOR;
                        CONSTANT SrcRegMode :  IN regmode_type
                     -- synopsys synthesis_off
						      := DefaultRegMode 
                     -- synopsys synthesis_on
                      );
--------------------------------------------------------------------------------
    PROCEDURE SregRem ( SIGNAL result       : OUT STD_ULOGIC_VECTOR;
                        SIGNAL ZeroDivide   : OUT STD_ULOGIC;
                        CONSTANT dividend   :  IN STD_ULOGIC_VECTOR;
                        CONSTANT divisor    :  IN STD_ULOGIC_VECTOR;
                        CONSTANT SrcRegMode :  IN regmode_type
                     -- synopsys synthesis_off
						      := DefaultRegMode 
                     -- synopsys synthesis_on
                      );
--------------------------------------------------------------------------------
    PROCEDURE SregRem ( SIGNAL result       : OUT BIT_VECTOR;
                        SIGNAL ZeroDivide   : OUT BIT;
                        CONSTANT dividend   :  IN BIT_VECTOR;
                        CONSTANT divisor    :  IN BIT_VECTOR;
                        CONSTANT SrcRegMode :  IN regmode_type
                     -- synopsys synthesis_off
						      := DefaultRegMode 
                     -- synopsys synthesis_on
                      );
--+-----------------------------------------------------------------------------
--|     Function Name  : SregShift
--| 
--|     Overloading    : None
--|
--|     Purpose        : Bidirectional logical shift operator for logic vector.
--|
--|     Parameters     :
--|                      SrcReg      - input  std_logic_vector, vector to be shifted
--|                      DstReg      - ouput, std_logic_vector, shifted result
--|                      ShiftO      - output, std_ulogic, holds the 
--|                                            last bit shifted out 
--|                                          of register
--|                      direction   - input, Std_ulogic
--|                                         '0'  means right shift
--|                                         '1' | 'X'  means left shift, 
--|                                          default is left shift
--|                      FillVal     - input, Std_ulogic, value to fill register with. 
--|                                          default is '0'
--|                      Nbits       - input , NATURAL, number of positions to shift
--|                                          default is 1.
--|
--|     Result         : Shifted std_logic_vector
--|
--|     NOTE           : Defaults not allowed for synthesis.
--|
--|     Use            :
--|                      SIGNAL acc   : std_logic_vector ( 15 DOWNTO 0);
--|                      SIGNAL carry : std_ulogic;
--|
--|                      SregShift ( acc, acc, carry, '1', '0',3 );
--|-----------------------------------------------------------------------------
   PROCEDURE SregShift ( CONSTANT SrcReg    : IN std_logic_vector;
                         SIGNAL DstReg    : INOUT std_logic_vector;
                         SIGNAL ShiftO    : OUT std_ulogic; 
                         CONSTANT direction : IN std_ulogic
                     -- synopsys synthesis_off
						      := '1'
                     -- synopsys synthesis_on
                                                            ;
                         CONSTANT FillVal   : IN std_ulogic  
                     -- synopsys synthesis_off
						      := '0'
                     -- synopsys synthesis_on
                                                            ;
                         CONSTANT Nbits     : IN Natural
                     -- synopsys synthesis_off
						       := 1 
                     -- synopsys synthesis_on
                      ) ;
--------------------------------------------------------------------------------
   PROCEDURE SregShift ( CONSTANT SrcReg    : IN std_ulogic_vector;
                         SIGNAL DstReg    : INOUT std_ulogic_vector;
                         SIGNAL ShiftO    : OUT std_ulogic; 
                         CONSTANT direction : IN std_ulogic
                     -- synopsys synthesis_off
						      := '1'
                     -- synopsys synthesis_on
                                                            ;
                         CONSTANT FillVal   : IN std_ulogic  
                     -- synopsys synthesis_off
						      := '0'
                     -- synopsys synthesis_on
                                                            ;
                         CONSTANT Nbits     : IN Natural
                     -- synopsys synthesis_off
						       := 1 
                     -- synopsys synthesis_on
                      ) ;
--------------------------------------------------------------------------------
   PROCEDURE SregShift ( CONSTANT SrcReg    : IN bit_vector;
                         SIGNAL DstReg    : INOUT bit_vector;
                         SIGNAL ShiftO    : OUT bit; 
                         CONSTANT direction : IN bit
                     -- synopsys synthesis_off
						      := '1'
                     -- synopsys synthesis_on
                                                            ;
                         CONSTANT FillVal   : IN bit  
                     -- synopsys synthesis_off
						      := '0'
                     -- synopsys synthesis_on
                                                            ;
                         CONSTANT Nbits     : IN Natural
                     -- synopsys synthesis_off
						       := 1 
                     -- synopsys synthesis_on
                      );
     -------------------------------------------------------------------------------
     --     Function Name : RegEqual
     -- 1.2.49
     --     Overloading   : Input parameter TYPEs.
     --
     --     Purpose       : Compute equality relation for bit_vector
     --
     --     Parameters    : l       - input bit_vector | INTEGER
     --                     r       - input bit_vector | INTEGER
     --                     SrcRegMode - input regmode_type, indicating the format of
     --                               the bit_vector operands (l,r).
     --                               Default is TwosComp.
     --
     --     Result        : BOOLEAN | bit. 
     --
     --     NOTE          : The operands may be of any length, and may be different
     --                     lengths.
     --
     --                     Overloading not defined for both inputs of INTEGER type.
     --     Use           :
     --                      VARIABLE a, b : bit_vector ( 7 DOWNTO 0 );
     --                      IF ( RegEqual ( a, b, TwosComp)   )  THEN
     --
     --     See Also      : RegLessThanOrEqual, RegGreaterThan, RegGreaterThanOrEqual.
     -------------------------------------------------------------------------------
     FUNCTION RegEqual     ( CONSTANT l          : IN bit_vector;
			     CONSTANT r          : IN bit_vector;
			     CONSTANT SrcRegMode : IN regmode_type
                     -- synopsys synthesis_off
							      := DefaultRegMode 
                     -- synopsys synthesis_on
			   ) RETURN bit;
     -----------------------------------------------------------------------------
     FUNCTION RegEqual    (  CONSTANT l        : IN bit_vector;
			     CONSTANT r        : IN bit_vector;
			     CONSTANT SrcRegMode : IN regmode_type
                     -- synopsys synthesis_off
							      := DefaultRegMode 
                     -- synopsys synthesis_on
			   ) RETURN BOOLEAN;
     -- -----------------------------------------------------------------------------
     FUNCTION RegEqual     ( CONSTANT l          : IN bit_vector;
			     CONSTANT r          : IN INTEGER;
			     CONSTANT SrcRegMode : IN regmode_type
                     -- synopsys synthesis_off
					         	      := DefaultRegMode 
                     -- synopsys synthesis_on
			   ) RETURN BOOLEAN;
     -------------------------------------------------------------------------------
     FUNCTION RegEqual    (  CONSTANT l          : IN INTEGER;
			     CONSTANT r          : IN bit_vector;
			     CONSTANT SrcRegMode : IN regmode_type
                     -- synopsys synthesis_off
					         	      := DefaultRegMode 
                     -- synopsys synthesis_on
			   ) RETURN BOOLEAN;
     -------------------------------------------------------------------------------
     FUNCTION RegEqual     ( CONSTANT l          : IN bit_vector;
			     CONSTANT r          : IN INTEGER;
			     CONSTANT SrcRegMode : IN regmode_type 
                     -- synopsys synthesis_off
					         	      := DefaultRegMode 
                     -- synopsys synthesis_on
			   ) RETURN bit;
     -------------------------------------------------------------------------------
     FUNCTION RegEqual    (  CONSTANT l          : IN INTEGER;
			     CONSTANT r          : IN bit_vector;
			     CONSTANT SrcRegMode : IN regmode_type 
                     -- synopsys synthesis_off
					         	      := DefaultRegMode 
                     -- synopsys synthesis_on
			   ) RETURN bit;
     -------------------------------------------------------------------------------
     --     Function Name : RegEqual
     --
     --     Overloading   : Input parameter TYPEs.
     --    
     --     Purpose       : Compute equality relation for std_logic_vectors
     --     
     --     Parameters    : l       - input std_logic_vector | INTEGER
     --                     r       - input std_logic_vector | INTEGER
     --                     SrcRegMode - input regmode_type, indicating the format of
     --                               the std_logic_vector operands (l,r).
     --                               Default is TwosComp.
     --   					  
     --     Result        : BOOLEAN relation. A TRUE value is returned if: l = r
     --
     --     NOTE          : The operands may be of any length, and may be different
     --                     lengths. 
     --
     --                     Overloading not defined for both inputs of INTEGER type.
     --
     --                    Any time the comparison reaches an index that has an 'X'  
     --                    as an array element, the comparison is deemed indeterminate
     --                    and will return false in case of boolean and '0' incase of
     --                    std_ulogic for synthesis purposes.
     --     Use           : 
     --                      VARIABLE a, b : std_logic_vector ( 7 DOWNTO 0 );
     --                      IF ( RegEqual ( a, b, TwosComp)   )  THEN 
     --     
     --     See Also      :  RegLessThan, RegLessThanOrEqual, RegGreaterThan, 
     --                     RegGreaterThanOrEqual.
     -------------------------------------------------------------------------------
     FUNCTION RegEqual     ( CONSTANT l          : IN std_logic_vector;
			     CONSTANT r          : IN std_logic_vector;
			     CONSTANT SrcRegMode : IN regmode_type
                     -- synopsys synthesis_off
							      := DefaultRegMode 
                     -- synopsys synthesis_on
			   ) RETURN std_ulogic;
     -----------------------------------------------------------------------------
     FUNCTION RegEqual    (  CONSTANT l        : IN std_logic_vector;
			     CONSTANT r        : IN std_logic_vector;
			     CONSTANT SrcRegMode : IN regmode_type
                     -- synopsys synthesis_off
							      := DefaultRegMode 
                     -- synopsys synthesis_on
			   ) RETURN BOOLEAN;
     -- -----------------------------------------------------------------------------
     FUNCTION RegEqual     ( CONSTANT l          : IN std_logic_vector;
			     CONSTANT r          : IN INTEGER;
			     CONSTANT SrcRegMode : IN regmode_type
                     -- synopsys synthesis_off
					         	      := DefaultRegMode 
                     -- synopsys synthesis_on
			   ) RETURN BOOLEAN;
     -------------------------------------------------------------------------------
     FUNCTION RegEqual    (  CONSTANT l          : IN INTEGER;
			     CONSTANT r          : IN std_logic_vector;
			     CONSTANT SrcRegMode : IN regmode_type
                     -- synopsys synthesis_off
					         	      := DefaultRegMode 
                     -- synopsys synthesis_on
			   ) RETURN BOOLEAN;
     -------------------------------------------------------------------------------
     FUNCTION RegEqual     ( CONSTANT l          : IN std_logic_vector;
			     CONSTANT r          : IN INTEGER;
			     CONSTANT SrcRegMode : IN regmode_type 
                     -- synopsys synthesis_off
					         	      := DefaultRegMode 
                     -- synopsys synthesis_on
			   ) RETURN std_ulogic;
     -------------------------------------------------------------------------------
     FUNCTION RegEqual    (  CONSTANT l          : IN INTEGER;
			     CONSTANT r          : IN std_logic_vector;
			     CONSTANT SrcRegMode : IN regmode_type 
                     -- synopsys synthesis_off
					         	      := DefaultRegMode 
                     -- synopsys synthesis_on
			   ) RETURN std_ulogic;
     -------------------------------------------------------------------------------
     --     Function Name : RegEqual
     --
     --     Overloading   : Input parameter TYPEs.
     --    
     --     Purpose       : Compute equality relation for std_ulogic_vectors
     --     
     --     Parameters    : l       - input std_ulogic_vector | INTEGER
     --                     r       - input std_ulogic_vector | INTEGER
     --                     SrcRegMode - input regmode_type, indicating the format of
     --                               the std_ulogic_vector operands (l,r).
     --                               Default is TwosComp.
     --     
     --     Result        : BOOLEAN relation. A TRUE value is returned if: l =  r
     --
     --     NOTE          : The operands may be of any length, and may be different
     --                     lengths. 
     --
     --                     Overloading not defined for both inputs of INTEGER type.
     --
     --
     --                     Any time the comparison reaches an index that has an 'X' as an
     --                     array element, the comparison is deemed indeterminate and will 
     --                     return false in case of boolean and '0' incase of std_ulogic for
     --                     synthesis purposes.
     --     Use           : 
     --                      VARIABLE a, b : std_ulogic_vector ( 7 DOWNTO 0 );
     --                      IF ( RegEqual ( a, b, TwosComp)   )  THEN 
     --     
     --     See Also      :  RegLessThan, RegLessThanOrEqual, RegGreaterThan, 
     --                     RegGreaterThanOrEqual.
     -------------------------------------------------------------------------------
     FUNCTION RegEqual     ( CONSTANT l          : IN std_ulogic_vector;
			     CONSTANT r          : IN std_ulogic_vector;
			     CONSTANT SrcRegMode : IN regmode_type
                     -- synopsys synthesis_off
							      := DefaultRegMode 
                     -- synopsys synthesis_on
			   ) RETURN std_ulogic;
     -----------------------------------------------------------------------------
     FUNCTION RegEqual    (  CONSTANT l        : IN std_ulogic_vector;
			     CONSTANT r        : IN std_ulogic_vector;
			     CONSTANT SrcRegMode : IN regmode_type
                     -- synopsys synthesis_off
							      := DefaultRegMode 
                     -- synopsys synthesis_on
			   ) RETURN BOOLEAN;
     -- -----------------------------------------------------------------------------
     FUNCTION RegEqual     ( CONSTANT l          : IN std_ulogic_vector;
			     CONSTANT r          : IN INTEGER;
			     CONSTANT SrcRegMode : IN regmode_type
                     -- synopsys synthesis_off
					         	      := DefaultRegMode 
                     -- synopsys synthesis_on
			   ) RETURN BOOLEAN;
     -------------------------------------------------------------------------------
     FUNCTION RegEqual    (  CONSTANT l          : IN INTEGER;
			     CONSTANT r          : IN std_ulogic_vector;
			     CONSTANT SrcRegMode : IN regmode_type
                     -- synopsys synthesis_off
					         	      := DefaultRegMode 
                     -- synopsys synthesis_on
			   ) RETURN BOOLEAN;
     -------------------------------------------------------------------------------
     FUNCTION RegEqual     ( CONSTANT l          : IN std_ulogic_vector;
			     CONSTANT r          : IN INTEGER;
			     CONSTANT SrcRegMode : IN regmode_type 
                     -- synopsys synthesis_off
					         	      := DefaultRegMode 
                     -- synopsys synthesis_on
			   ) RETURN std_ulogic;
     -------------------------------------------------------------------------------
     FUNCTION RegEqual    (  CONSTANT l          : IN INTEGER;
			     CONSTANT r          : IN std_ulogic_vector;
			     CONSTANT SrcRegMode : IN regmode_type 
                     -- synopsys synthesis_off
					         	      := DefaultRegMode 
                     -- synopsys synthesis_on
			   ) RETURN std_ulogic;
     -------------------------------------------------------------------------------
     --     Function Name : RegNotEqual
     -- 1.2.49
     --     Overloading   : Input parameter TYPEs.
     --
     --     Purpose       : Compute un-equality relation for bit_vector
     --
     --     Parameters    : l       - input bit_vector | INTEGER
     --                     r       - input bit_vector | INTEGER
     --                     SrcRegMode - input regmode_type, indicating the format of
     --                               the bit_vector operands (l,r).
     --                               Default is TwosComp.
     --
     --     Result        : BOOLEAN | bit. 
     --
     --     NOTE          : The operands may be of any length, and may be different
     --                     lengths.
     --
     --                     Overloading not defined for both inputs of INTEGER type.
     --     Use           :
     --                      VARIABLE a, b : bit_vector ( 7 DOWNTO 0 );
     --                      IF ( RegNotEqual ( a, b, TwosComp)   )  THEN
     --
     --     See Also      : RegLessThanOrEqual, RegGreaterThan, RegGreaterThanOrEqual.
     -------------------------------------------------------------------------------
     FUNCTION RegNotEqual     ( CONSTANT l          : IN bit_vector;
			     CONSTANT r          : IN bit_vector;
			     CONSTANT SrcRegMode : IN regmode_type
                     -- synopsys synthesis_off
							      := DefaultRegMode 
                     -- synopsys synthesis_on
			   ) RETURN bit;
     -----------------------------------------------------------------------------
     FUNCTION RegNotEqual    (  CONSTANT l        : IN bit_vector;
			     CONSTANT r        : IN bit_vector;
			     CONSTANT SrcRegMode : IN regmode_type
                     -- synopsys synthesis_off
							      := DefaultRegMode 
                     -- synopsys synthesis_on
			   ) RETURN BOOLEAN;
     -- -----------------------------------------------------------------------------
     FUNCTION RegNotEqual     ( CONSTANT l          : IN bit_vector;
			     CONSTANT r          : IN INTEGER;
			     CONSTANT SrcRegMode : IN regmode_type
                     -- synopsys synthesis_off
					         	      := DefaultRegMode 
                     -- synopsys synthesis_on
			   ) RETURN BOOLEAN;
     -------------------------------------------------------------------------------
     FUNCTION RegNotEqual    (  CONSTANT l          : IN INTEGER;
			     CONSTANT r          : IN bit_vector;
			     CONSTANT SrcRegMode : IN regmode_type
                     -- synopsys synthesis_off
					         	      := DefaultRegMode 
                     -- synopsys synthesis_on
			   ) RETURN BOOLEAN;
     -------------------------------------------------------------------------------
     FUNCTION RegNotEqual     ( CONSTANT l          : IN bit_vector;
			     CONSTANT r          : IN INTEGER;
			     CONSTANT SrcRegMode : IN regmode_type 
                     -- synopsys synthesis_off
					         	      := DefaultRegMode 
                     -- synopsys synthesis_on
			   ) RETURN bit;
     -------------------------------------------------------------------------------
     FUNCTION RegNotEqual    (  CONSTANT l          : IN INTEGER;
			     CONSTANT r          : IN bit_vector;
			     CONSTANT SrcRegMode : IN regmode_type 
                     -- synopsys synthesis_off
					         	      := DefaultRegMode 
                     -- synopsys synthesis_on
			   ) RETURN bit;
     -------------------------------------------------------------------------------
     --     Function Name : RegNotEqual
     --
     --     Overloading   : Input parameter TYPEs.
     --    
     --     Purpose       : Compute un-equality relation for std_logic_vectors
     --     
     --     Parameters    : l       - input std_logic_vector | INTEGER
     --                     r       - input std_logic_vector | INTEGER
     --                     SrcRegMode - input regmode_type, indicating the format of
     --                               the std_logic_vector operands (l,r).
     --                               Default is TwosComp.
     --   					  
     --     Result        : BOOLEAN relation. A TRUE value is returned if: l = r
     --
     --     NOTE          : The operands may be of any length, and may be different
     --                     lengths. 
     --
     --                     Overloading not defined for both inputs of INTEGER type.
     --
     --                     Any time the comparison reaches an index that has an 'X'
     --                     as an array element, the comparison is deemed indeterminate
     --                     and will return false in case of boolean and '0' incase of
     --                     std_ulogic for synthesis purposes.
     --     Use           : 
     --                      VARIABLE a, b : std_logic_vector ( 7 DOWNTO 0 );
     --                      IF ( RegNotEqual ( a, b, TwosComp)   )  THEN 
     --     
     --     See Also      :  RegLessThan, RegLessThanOrEqual, RegGreaterThan, 
     --                     RegGreaterThanOrEqual.
     -------------------------------------------------------------------------------
     FUNCTION RegNotEqual     ( CONSTANT l          : IN std_logic_vector;
			     CONSTANT r          : IN std_logic_vector;
			     CONSTANT SrcRegMode : IN regmode_type
                     -- synopsys synthesis_off
							      := DefaultRegMode 
                     -- synopsys synthesis_on
			   ) RETURN std_ulogic;
     -----------------------------------------------------------------------------
     FUNCTION RegNotEqual    (  CONSTANT l        : IN std_logic_vector;
			     CONSTANT r        : IN std_logic_vector;
			     CONSTANT SrcRegMode : IN regmode_type
                     -- synopsys synthesis_off
							      := DefaultRegMode 
                     -- synopsys synthesis_on
			   ) RETURN BOOLEAN;

     -- -----------------------------------------------------------------------------
     FUNCTION RegNotEqual     ( CONSTANT l          : IN std_logic_vector;
			     CONSTANT r          : IN INTEGER;
			     CONSTANT SrcRegMode : IN regmode_type
                     -- synopsys synthesis_off
					         	      := DefaultRegMode 
                     -- synopsys synthesis_on
			   ) RETURN BOOLEAN;
     -------------------------------------------------------------------------------
     FUNCTION RegNotEqual    (  CONSTANT l          : IN INTEGER;
			     CONSTANT r          : IN std_logic_vector;
			     CONSTANT SrcRegMode : IN regmode_type
                     -- synopsys synthesis_off
					         	      := DefaultRegMode 
                     -- synopsys synthesis_on
			   ) RETURN BOOLEAN;
     -------------------------------------------------------------------------------
     FUNCTION RegNotEqual     ( CONSTANT l          : IN std_logic_vector;
			     CONSTANT r          : IN INTEGER;
			     CONSTANT SrcRegMode : IN regmode_type 
                     -- synopsys synthesis_off
					         	      := DefaultRegMode 
                     -- synopsys synthesis_on
			   ) RETURN std_ulogic;
     -------------------------------------------------------------------------------
     FUNCTION RegNotEqual    (  CONSTANT l          : IN INTEGER;
			     CONSTANT r          : IN std_logic_vector;
			     CONSTANT SrcRegMode : IN regmode_type 
                     -- synopsys synthesis_off
					         	      := DefaultRegMode 
                     -- synopsys synthesis_on
			   ) RETURN std_ulogic;
     -------------------------------------------------------------------------------
     --     Function Name : RegNotEqual
     --
     --     Overloading   : Input parameter TYPEs.
     --    
     --     Purpose       : Compute un-equality relation for std_ulogic_vectors
     --     
     --     Parameters    : l       - input std_ulogic_vector | INTEGER
     --                     r       - input std_ulogic_vector | INTEGER
     --                     SrcRegMode - input regmode_type, indicating the format of
     --                               the std_ulogic_vector operands (l,r).
     --                               Default is TwosComp.
     --     
     --     Result        : BOOLEAN relation. A TRUE value is returned if: l =  r
     --
     --     NOTE          : The operands may be of any length, and may be different
     --                     lengths. 
     --
     --                     Overloading not defined for both inputs of INTEGER type.
     --
     --                     Any time the comparison reaches an index that has an 'X' as
     --                     an array element, the comparison is deemed indeterminate  
     --                     and will return false in case of boolean and '0' incase of
     --                     std_ulogic for synthesis purposes.
     --     Use           : 
     --                      VARIABLE a, b : std_ulogic_vector ( 7 DOWNTO 0 );
     --                      IF ( RegNotEqual ( a, b, TwosComp)   )  THEN 
     --     
     --     See Also      : RegLessThan, RegLessThanOrEqual, RegGreaterThan, 
     --                     RegGreaterThanOrEqual.
     -------------------------------------------------------------------------------
     FUNCTION RegNotEqual     ( CONSTANT l          : IN std_ulogic_vector;
			     CONSTANT r          : IN std_ulogic_vector;
			     CONSTANT SrcRegMode : IN regmode_type
                     -- synopsys synthesis_off
							      := DefaultRegMode 
                     -- synopsys synthesis_on
			   ) RETURN std_ulogic;
     -----------------------------------------------------------------------------
     FUNCTION RegNotEqual    (  CONSTANT l        : IN std_ulogic_vector;
			     CONSTANT r        : IN std_ulogic_vector;
			     CONSTANT SrcRegMode : IN regmode_type
                     -- synopsys synthesis_off
							      := DefaultRegMode 
                     -- synopsys synthesis_on
			   ) RETURN BOOLEAN;

     -- -----------------------------------------------------------------------------
     FUNCTION RegNotEqual     ( CONSTANT l          : IN std_ulogic_vector;
			     CONSTANT r          : IN INTEGER;
			     CONSTANT SrcRegMode : IN regmode_type
                     -- synopsys synthesis_off
					         	      := DefaultRegMode 
                     -- synopsys synthesis_on
			   ) RETURN BOOLEAN;
     -------------------------------------------------------------------------------
     FUNCTION RegNotEqual    (  CONSTANT l          : IN INTEGER;
			     CONSTANT r          : IN std_ulogic_vector;
			     CONSTANT SrcRegMode : IN regmode_type
                     -- synopsys synthesis_off
					         	      := DefaultRegMode 
                     -- synopsys synthesis_on
			   ) RETURN BOOLEAN;
     -------------------------------------------------------------------------------
     FUNCTION RegNotEqual     ( CONSTANT l          : IN std_ulogic_vector;
			     CONSTANT r          : IN INTEGER;
			     CONSTANT SrcRegMode : IN regmode_type 
                     -- synopsys synthesis_off
					         	      := DefaultRegMode 
                     -- synopsys synthesis_on
			   ) RETURN std_ulogic;
     -------------------------------------------------------------------------------
     FUNCTION RegNotEqual    (  CONSTANT l          : IN INTEGER;
			     CONSTANT r          : IN std_ulogic_vector;
			     CONSTANT SrcRegMode : IN regmode_type 
                     -- synopsys synthesis_off
					         	      := DefaultRegMode 
                     -- synopsys synthesis_on
			   ) RETURN std_ulogic;
     -------------------------------------------------------------------------------
     --     Function Name : RegLessThan
     -- 1.2.49
     --     Overloading   : Input parameter TYPEs.
     --
     --     Purpose       : Compute a less than relation for bit_vector
     --
     --     Parameters    : l       - input bit_vector | INTEGER
     --                     r       - input bit_vector | INTEGER
     --                     SrcRegMode - input regmode_type, indicating the format of
     --                               the bit_vector operands (l,r).
     --                               Default is TwosComp.
     --
     --     Result        : BOOLEAN | bit. 
     --
     --     NOTE          : The operands may be of any length, and may be different
     --                     lengths.
     --
     --                     Overloading not defined for both inputs of INTEGER type.
     --     Use           :
     --                      VARIABLE a, b : bit_vector ( 7 DOWNTO 0 );
     --                      IF ( RegLessThan ( a, b, TwosComp)   )  THEN
     --
     --     See Also      : RegLessThanOrEqual, RegGreaterThan, RegGreaterThanOrEqual.
     -------------------------------------------------------------------------------
     FUNCTION RegLessThan  ( CONSTANT l          : IN bit_vector;
			     CONSTANT r          : IN bit_vector;
			     CONSTANT SrcRegMode : IN regmode_type
                     -- synopsys synthesis_off
						      := DefaultRegMode 
                     -- synopsys synthesis_on
			   ) RETURN bit;
     -------------------------------------------------------------------------------
     FUNCTION RegLessThan  ( CONSTANT l          : IN bit_vector;
			     CONSTANT r          : IN bit_vector;
			     CONSTANT SrcRegMode : IN regmode_type
                     -- synopsys synthesis_off
						      := DefaultRegMode 
                     -- synopsys synthesis_on
			   ) RETURN BOOLEAN;
     -- -----------------------------------------------------------------------------
     FUNCTION RegLessThan  ( CONSTANT l          : IN bit_vector;
			     CONSTANT r          : IN INTEGER;
			     CONSTANT SrcRegMode : IN regmode_type
                     -- synopsys synthesis_off
						      := DefaultRegMode 
                     -- synopsys synthesis_on
			   ) RETURN BOOLEAN;
     -------------------------------------------------------------------------------
     FUNCTION RegLessThan (  CONSTANT l          : IN INTEGER;
			     CONSTANT r          : IN bit_vector;
			     CONSTANT SrcRegMode : IN regmode_type
                     -- synopsys synthesis_off
						      := DefaultRegMode 
                     -- synopsys synthesis_on
			   ) RETURN BOOLEAN;
     -------------------------------------------------------------------------------
     FUNCTION RegLessThan  ( CONSTANT l          : IN bit_vector;
			     CONSTANT r          : IN INTEGER;
			     CONSTANT SrcRegMode : IN regmode_type
                     -- synopsys synthesis_off
						      := DefaultRegMode 
                     -- synopsys synthesis_on
			   ) RETURN bit;
     -------------------------------------------------------------------------------
     FUNCTION RegLessThan (  CONSTANT l          : IN INTEGER;
			     CONSTANT r          : IN bit_vector;
			     CONSTANT SrcRegMode : IN regmode_type
                     -- synopsys synthesis_off
						      := DefaultRegMode 
                     -- synopsys synthesis_on
			   ) RETURN bit;
     -------------------------------------------------------------------------------
     --     Function Name : RegLessThan
     --
     --     Overloading   : Input parameter TYPEs.
     --    
     --     Purpose       : Compute a less than relation for std_logic_vectors
     --     
     --     Parameters    : l       - input std_logic_vector | INTEGER
     --                     r       - input std_logic_vector | INTEGER
     --                     SrcRegMode - input regmode_type, indicating the format of
     --                               the std_logic_vector operands (l,r).
     --                               Default is TwosComp.
     --     
     --     Result        : BOOLEAN | std_ulogic
     --
     --     NOTE          : The operands may be of any length, and may be different
     --                     lengths. 
     --
     --                     Overloading not defined for both inputs of INTEGER type.
     --
     --                     Any time the comparison reaches an index that has an 'X' as an
     --                     array element, the comparison is deemed indeterminate and will 
     --                     return false in case of boolean and '0' incase of
     --                     std_ulogic for synthesis purposes.
     --     Use           : 
     --                      VARIABLE a, b : std_logic_vector ( 7 DOWNTO 0 );
     --                      IF ( RegLessThan ( a, b, TwosComp)   )  THEN 
     --     
     --     See Also      : RegLessThanOrEqual, RegGreaterThan, RegGreaterThanOrEqual.
     -------------------------------------------------------------------------------
     FUNCTION RegLessThan  ( CONSTANT l          : IN std_logic_vector;
			     CONSTANT r          : IN std_logic_vector;
			     CONSTANT SrcRegMode : IN regmode_type
                     -- synopsys synthesis_off
						      := DefaultRegMode 
                     -- synopsys synthesis_on
			   ) RETURN std_ulogic;
     -----------------------------------------------------------------------------
     FUNCTION RegLessThan (  CONSTANT l          : IN std_logic_vector;
			     CONSTANT r          : IN std_logic_vector;
			     CONSTANT SrcRegMode : IN regmode_type
                     -- synopsys synthesis_off
						      := DefaultRegMode 
                     -- synopsys synthesis_on
			   ) RETURN BOOLEAN;
     -- -----------------------------------------------------------------------------
     FUNCTION RegLessThan  ( CONSTANT l          : IN std_logic_vector;
			     CONSTANT r          : IN INTEGER;
			     CONSTANT SrcRegMode : IN regmode_type
                     -- synopsys synthesis_off
						      := DefaultRegMode 
                     -- synopsys synthesis_on
			   ) RETURN BOOLEAN;
     -------------------------------------------------------------------------------
     FUNCTION RegLessThan (  CONSTANT l          : IN INTEGER;
			     CONSTANT r          : IN std_logic_vector;
			     CONSTANT SrcRegMode : IN regmode_type
                     -- synopsys synthesis_off
						      := DefaultRegMode 
                     -- synopsys synthesis_on

			   ) RETURN BOOLEAN;
     -------------------------------------------------------------------------------
     FUNCTION RegLessThan  ( CONSTANT l          : IN std_logic_vector;
			     CONSTANT r          : IN INTEGER;
			     CONSTANT SrcRegMode : IN regmode_type
                     -- synopsys synthesis_off
						      := DefaultRegMode 
                     -- synopsys synthesis_on

			   ) RETURN std_ulogic;
     -------------------------------------------------------------------------------
     FUNCTION RegLessThan (  CONSTANT l          : IN INTEGER;
			     CONSTANT r          : IN std_logic_vector;
			     CONSTANT SrcRegMode : IN regmode_type
                     -- synopsys synthesis_off
						      := DefaultRegMode 
                     -- synopsys synthesis_on

			   ) RETURN std_ulogic;
     -------------------------------------------------------------------------------
     --     Function Name : RegLessThan
     --
     --     Overloading   : Input parameter TYPEs.
     --    
     --     Purpose       : Compute a less than relation for std_ulogic_vectors
     --     
     --     Parameters    : l       - input std_ulogic_vector | INTEGER
     --                     r       - input std_ulogic_vector | INTEGER
     --                     SrcRegMode - input regmode_type, indicating the format of
     --                               the std_ulogic_vector operands (l,r).
     --                               Default is TwosComp.
     --     
     --     Result        : BOOLEAN | std_ulogic
     --
     --     NOTE          : The operands may be of any length, and may be different
     --                     lengths. 
     --
     --                     Overloading not defined for both inputs of INTEGER type.
     --
     --                     Any time the comparison reaches an index that has an 'X' as an
     --                     array element, the comparison is deemed indeterminate and will 
     --                     return false in case of boolean and '0' incase of 
     --                     std_ulogic for synthesis purposes.
     --     Use           : 
     --                      VARIABLE a, b : std_ulogic_vector ( 7 DOWNTO 0 );
     --                      IF ( RegLessThan ( a, b, TwosComp)   )  THEN 
     --     
     --     See Also      : RegLessThanOrEqual,RegGreaterThan,RegGreaterThanOrEqual.
     -------------------------------------------------------------------------------
     FUNCTION RegLessThan  ( CONSTANT l          : IN std_ulogic_vector;
			     CONSTANT r          : IN std_ulogic_vector;
			     CONSTANT SrcRegMode : IN regmode_type
                     -- synopsys synthesis_off
						      := DefaultRegMode 
                     -- synopsys synthesis_on

			   ) RETURN std_ulogic;
     -----------------------------------------------------------------------------
     FUNCTION RegLessThan (  CONSTANT l          : IN std_ulogic_vector;
			     CONSTANT r          : IN std_ulogic_vector;
			     CONSTANT SrcRegMode : IN regmode_type
                     -- synopsys synthesis_off
						      := DefaultRegMode 
                     -- synopsys synthesis_on

			   ) RETURN BOOLEAN;
     -- -----------------------------------------------------------------------------
     FUNCTION RegLessThan  ( CONSTANT l          : IN std_ulogic_vector;
			     CONSTANT r          : IN INTEGER;
			     CONSTANT SrcRegMode : IN regmode_type
                     -- synopsys synthesis_off
						      := DefaultRegMode 
                     -- synopsys synthesis_on

			   ) RETURN BOOLEAN;
     -------------------------------------------------------------------------------
     FUNCTION RegLessThan (  CONSTANT l          : IN INTEGER;
			     CONSTANT r          : IN std_ulogic_vector;
			     CONSTANT SrcRegMode : IN regmode_type
                     -- synopsys synthesis_off
						      := DefaultRegMode 
                     -- synopsys synthesis_on
			   ) RETURN BOOLEAN;
     -------------------------------------------------------------------------------
     FUNCTION RegLessThan  ( CONSTANT l          : IN std_ulogic_vector;
			     CONSTANT r          : IN INTEGER;
			     CONSTANT SrcRegMode : IN regmode_type
                     -- synopsys synthesis_off
						      := DefaultRegMode 
                     -- synopsys synthesis_on
			   ) RETURN std_ulogic;
     -------------------------------------------------------------------------------
     FUNCTION RegLessThan (  CONSTANT l          : IN INTEGER;
			     CONSTANT r          : IN std_ulogic_vector;
			     CONSTANT SrcRegMode : IN regmode_type
                     -- synopsys synthesis_off
						      := DefaultRegMode 
                     -- synopsys synthesis_on
			   ) RETURN std_ulogic;
     -------------------------------------------------------------------------------
     --     Function Name : RegLessThanOrEqual
     -- 1.2.51
     --     Overloading   : Input parameter TYPEs.
     --
     --     Purpose       : Compute a less than or equal relation for bit_vectors
     --
     --     Parameters    : l       - input bit_vector | INTEGER
     --                     r       - input bit_vector | INTEGER
     --                     SrcRegMode - input regmode_type, indicating the format of
     --                               the bit_vector operands (l,r).
     --                               Default is TwosComp.
     --
     --     Result        : BOOLEAN | bit
     --
     --     NOTE          : The operands may be of any length, and may be different
     --                     lengths.
     --
     --                     Overloading not defined for both inputs of INTEGER type.
     --     Use           :
     --                      VARIABLE a, b : bit_vector ( 7 DOWNTO 0 );
     --                      IF ( RegLessThanOrEqual ( a, b, TwosComp)   )  THEN
     --
     --     See Also      : RegLessThan,RegGreaterThan,  RegGreaterThanOrEqual.
     -------------------------------------------------------------------------------
     FUNCTION RegLessThanOrEqual ( CONSTANT l          : IN bit_vector;
				   CONSTANT r          : IN bit_vector;
				   CONSTANT SrcRegMode : IN regmode_type
                     -- synopsys synthesis_off
							      := DefaultRegMode 
                     -- synopsys synthesis_on
				 ) RETURN bit;
     -----------------------------------------------------------------------------
     FUNCTION RegLessThanOrEqual ( CONSTANT l          : IN bit_vector;
				   CONSTANT r          : IN bit_vector;
 			           CONSTANT SrcRegMode : IN regmode_type
                     -- synopsys synthesis_off
							      := DefaultRegMode 
                     -- synopsys synthesis_on
				 ) RETURN BOOLEAN;
     -- -----------------------------------------------------------------------------
     FUNCTION RegLessThanOrEqual ( CONSTANT l          : IN bit_vector;
				   CONSTANT r          : IN INTEGER;
			     CONSTANT SrcRegMode : IN regmode_type
                     -- synopsys synthesis_off
						      := DefaultRegMode 
                     -- synopsys synthesis_on
				 ) RETURN BOOLEAN;
     -------------------------------------------------------------------------------
     FUNCTION RegLessThanOrEqual ( CONSTANT l          : IN INTEGER;
				   CONSTANT r          : IN bit_vector;
  			           CONSTANT SrcRegMode : IN regmode_type
                     -- synopsys synthesis_off
					         	      := DefaultRegMode 
                     -- synopsys synthesis_on
				 ) RETURN BOOLEAN;
     -------------------------------------------------------------------------------
     FUNCTION RegLessThanOrEqual ( CONSTANT l          : IN bit_vector;
				   CONSTANT r          : IN INTEGER;
  			           CONSTANT SrcRegMode : IN regmode_type
                     -- synopsys synthesis_off
					         	      := DefaultRegMode 
                     -- synopsys synthesis_on
				 ) RETURN bit;
     -------------------------------------------------------------------------------
     FUNCTION RegLessThanOrEqual ( CONSTANT l          : IN INTEGER;
				   CONSTANT r          : IN bit_vector;
  			           CONSTANT SrcRegMode : IN regmode_type
                     -- synopsys synthesis_off
					         	      := DefaultRegMode 
                     -- synopsys synthesis_on
				 ) RETURN bit;
     -- ----------------------------------------------------------------------------
     --     Function Name : RegLessThanOrEqual
     --    
     --     Purpose       : Compute a less than or equal relation for std_logic_vectors
     --     
     --     Parameters    : l       - input std_logic_vector | INTEGER
     --                     r       - input std_logic_vector | INTEGER
     --                     SrcRegMode - input regmode_type, indicating the format of
     --                               the std_logic_vector operands (l,r).
     --                               Default is TwosComp.
     --     
     --     Result        : BOOLEAN | std_ulogic
     --
     --     NOTE          : The operands may be of any length, and may be different
     --                     lengths. 
     --
     --                     Overloading not defined for both inputs of INTEGER type.
     --                     Any time the comparison reaches an index that has an 'X' as an
     --                     array element, the comparison is deemed indeterminate and will 
     --                     return false in case of boolean and '0' incase of 
     --                     std_ulogic for synthesis purposes.
     --     Use           : 
     --                      VARIABLE a, b : std_logic_vector ( 7 DOWNTO 0 );
     --                      IF ( RegLessThanOrEqual ( a, b, TwosComp)   )  THEN 
     --     
     --     See Also      : RegLessThan, RegGreaterThan, RegGreaterThanOrEqual.
     -------------------------------------------------------------------------------
     FUNCTION RegLessThanOrEqual ( CONSTANT l          : IN std_logic_vector;
				   CONSTANT r          : IN std_logic_vector;
  			           CONSTANT SrcRegMode : IN regmode_type
                     -- synopsys synthesis_off
					         	      := DefaultRegMode 
                     -- synopsys synthesis_on
				 ) RETURN std_ulogic;
     -----------------------------------------------------------------------------
     FUNCTION RegLessThanOrEqual ( CONSTANT l          : IN std_logic_vector;
				   CONSTANT r          : IN std_logic_vector;
  			           CONSTANT SrcRegMode : IN regmode_type
                     -- synopsys synthesis_off
					         	      := DefaultRegMode 
                     -- synopsys synthesis_on
				 ) RETURN BOOLEAN;
     -- -----------------------------------------------------------------------------
     FUNCTION RegLessThanOrEqual ( CONSTANT l          : IN std_logic_vector;
				   CONSTANT r          : IN INTEGER;
  			           CONSTANT SrcRegMode : IN regmode_type
                     -- synopsys synthesis_off
					         	      := DefaultRegMode 
                     -- synopsys synthesis_on
				 ) RETURN BOOLEAN;
     -------------------------------------------------------------------------------
     FUNCTION RegLessThanOrEqual ( CONSTANT l          : IN INTEGER;
				   CONSTANT r          : IN std_logic_vector;
  			           CONSTANT SrcRegMode : IN regmode_type
                     -- synopsys synthesis_off
					         	      := DefaultRegMode 
                     -- synopsys synthesis_on
				 ) RETURN BOOLEAN;
     -------------------------------------------------------------------------------
     FUNCTION RegLessThanOrEqual ( CONSTANT l          : IN std_logic_vector;
				   CONSTANT r          : IN INTEGER;
  			           CONSTANT SrcRegMode : IN regmode_type
                     -- synopsys synthesis_off
					         	      := DefaultRegMode 
                     -- synopsys synthesis_on
				 ) RETURN std_ulogic;
     -------------------------------------------------------------------------------
     FUNCTION RegLessThanOrEqual ( CONSTANT l          : IN INTEGER;
				   CONSTANT r          : IN std_logic_vector;
  			           CONSTANT SrcRegMode : IN regmode_type
                     -- synopsys synthesis_off
					         	      := DefaultRegMode 
                     -- synopsys synthesis_on
				 ) RETURN std_ulogic;
     -- ----------------------------------------------------------------------------
     --     Function Name : RegLessThanOrEqual
     --    
     --     Purpose       : Compute a less than or equal relation for std_ulogic_vectors
     --     
     --     Parameters    : l       - input std_ulogic_vector | INTEGER
     --                     r       - input std_ulogic_vector | INTEGER
     --                     SrcRegMode - input regmode_type, indicating the format of
     --                               the std_ulogic_vector operands (l,r).
     --                               Default is TwosComp.
     --     
     --     Result        : BOOLEAN | std_ulogic
     --
     --     NOTE          : The operands may be of any length, and may be different
     --                     lengths. 
     --
     --                     Overloading not defined for both inputs of INTEGER type.
     --
     --                     Any time the comparison reaches an index that has an 'X' as an
     --                     array element, the comparison is deemed indeterminate and will 
     --                     return false in case of boolean and '0' incase of 
     --                     std_ulogic for synthesis purposes.
     --     Use           : 
     --                      VARIABLE a, b : std_ulogic_vector ( 7 DOWNTO 0 );
     --                      IF ( RegLessThanOrEqual ( a, b, TwosComp)   )  THEN 
     --     
     --     See Also      : RegLessThan, RegGreaterThan,   RegGreaterThanOrEqual.
     -------------------------------------------------------------------------------
     FUNCTION RegLessThanOrEqual ( CONSTANT l          : IN std_ulogic_vector;
				   CONSTANT r          : IN std_ulogic_vector;
  			           CONSTANT SrcRegMode : IN regmode_type
                     -- synopsys synthesis_off
					         	      := DefaultRegMode 
                     -- synopsys synthesis_on
				 ) RETURN std_ulogic;
     -----------------------------------------------------------------------------
     FUNCTION RegLessThanOrEqual ( CONSTANT l          : IN std_ulogic_vector;
				   CONSTANT r          : IN std_ulogic_vector;
  			           CONSTANT SrcRegMode : IN regmode_type
                     -- synopsys synthesis_off
					         	      := DefaultRegMode 
                     -- synopsys synthesis_on
				 ) RETURN BOOLEAN;
     -- -----------------------------------------------------------------------------
     FUNCTION RegLessThanOrEqual ( CONSTANT l          : IN std_ulogic_vector;
				   CONSTANT r          : IN INTEGER;
  			           CONSTANT SrcRegMode : IN regmode_type
                     -- synopsys synthesis_off
					         	      := DefaultRegMode 
                     -- synopsys synthesis_on
				 ) RETURN BOOLEAN;
     -------------------------------------------------------------------------------
     FUNCTION RegLessThanOrEqual ( CONSTANT l          : IN INTEGER;
				   CONSTANT r          : IN std_ulogic_vector;
  			           CONSTANT SrcRegMode : IN regmode_type
                     -- synopsys synthesis_off
					         	      := DefaultRegMode 
                     -- synopsys synthesis_on
				 ) RETURN BOOLEAN;
     -------------------------------------------------------------------------------
     FUNCTION RegLessThanOrEqual ( CONSTANT l          : IN std_ulogic_vector;
				   CONSTANT r          : IN INTEGER;
  			           CONSTANT SrcRegMode : IN regmode_type
                     -- synopsys synthesis_off
					         	      := DefaultRegMode 
                     -- synopsys synthesis_on
				 ) RETURN std_ulogic;
     -------------------------------------------------------------------------------
     FUNCTION RegLessThanOrEqual ( CONSTANT l          : IN INTEGER;
				   CONSTANT r          : IN std_ulogic_vector;
  			           CONSTANT SrcRegMode : IN regmode_type
                     -- synopsys synthesis_off
					         	      := DefaultRegMode 
                     -- synopsys synthesis_on
				 ) RETURN std_ulogic;

     -------------------------------------------------------------------------------
     --     Function Name : RegGreaterThan
     -- 1.2.53
     --     Overloading   : Input parameter TYPEs.
     --
     --     Purpose       : Compute a greater than relation for bit_vectors
     --
     --     Parameters    : l       - input bit_vector | INTEGER
     --                     r       - input bit_vector | INTEGER
     --                     SrcRegMode - input regmode_type, indicating the format of
     --                               the bit_vector operands (l,r).
     --                               Default is TwosComp.
     --
     --     Result        : BOOLEAN | bit
     --
     --     NOTE          : The operands may be of any length, and may be different
     --                     lengths.
     --
     --                     Overloading not defined for both inputs of INTEGER type.
     --     Use           :
     --                      VARIABLE a, b : bit_vector ( 7 DOWNTO 0 );
     --                      IF ( RegGreaterThan ( a, b, TwosComp)   )  THEN
     --
     --     See Also      : RegLessThan, RegLessThanOrEqual, RegGreaterThanOrEqual.
     -------------------------------------------------------------------------------
     FUNCTION RegGreaterThan ( CONSTANT l          : IN bit_vector;
			       CONSTANT r          : IN bit_vector;
		               CONSTANT SrcRegMode : IN regmode_type
                     -- synopsys synthesis_off
							      := DefaultRegMode 
                     -- synopsys synthesis_on
				 ) RETURN bit;
     -----------------------------------------------------------------------------
     FUNCTION RegGreaterThan    ( CONSTANT l          : IN bit_vector;
				   CONSTANT r          : IN bit_vector;
 			           CONSTANT SrcRegMode : IN regmode_type
                     -- synopsys synthesis_off
							      := DefaultRegMode 
                     -- synopsys synthesis_on
				 ) RETURN BOOLEAN;
     -- -----------------------------------------------------------------------------
     FUNCTION RegGreaterThan ( CONSTANT l          : IN bit_vector;
			       CONSTANT r          : IN INTEGER;
			       CONSTANT SrcRegMode : IN regmode_type
                     -- synopsys synthesis_off
						      := DefaultRegMode 
                     -- synopsys synthesis_on
				 ) RETURN BOOLEAN;
     -------------------------------------------------------------------------------
     FUNCTION RegGreaterThan ( CONSTANT l          : IN INTEGER;
				   CONSTANT r          : IN bit_vector;
  			           CONSTANT SrcRegMode : IN regmode_type
                     -- synopsys synthesis_off
					         	      := DefaultRegMode 
                     -- synopsys synthesis_on
				 ) RETURN BOOLEAN;
     -------------------------------------------------------------------------------
     FUNCTION RegGreaterThan ( CONSTANT l          : IN bit_vector;
			       CONSTANT r          : IN INTEGER;
  			       CONSTANT SrcRegMode : IN regmode_type
                     -- synopsys synthesis_off
					         	      := DefaultRegMode 
                     -- synopsys synthesis_on
				 ) RETURN bit;
     -------------------------------------------------------------------------------
     FUNCTION RegGreaterThan ( CONSTANT l          : IN INTEGER;
			       CONSTANT r          : IN bit_vector;
  			       CONSTANT SrcRegMode : IN regmode_type
                     -- synopsys synthesis_off
					         	      := DefaultRegMode 
                     -- synopsys synthesis_on
				 ) RETURN bit;
     -- ----------------------------------------------------------------------------
     --     Function Name : RegGreaterThan
     --
     --     Overloading   : Input parameter TYPEs.
     --    
     --     Purpose       : Compute a greater than relation for std_logic_vectors
     --     
     --     Parameters    : l       - input std_logic_vector | INTEGER
     --                     r       - input std_logic_vector | INTEGER
     --                     SrcRegMode - input regmode_type, indicating the format of
     --                               the std_logic_vector operands (l,r).
     --                               Default is TwosComp.
     --     
     --     Result        : BOOLEAN | std_ulogic
     --
     --     NOTE          : The operands may be of any length, and may be different
     --                     lengths. 
     --
     --                     Overloading not defined for both inputs of INTEGER type.
     --
     --                     Any time the comparison reaches an index that has an 'X' as an
     --                     array element, the comparison is deemed indeterminate and will 
     --                     return false in case of boolean and '0' incase of 
     --                     std_ulogic for synthesis purposes.
     --     Use           : 
     --                      VARIABLE a, b : std_logic_vector ( 7 DOWNTO 0 );
     --                      IF ( RegGreaterThan ( a, b, TwosComp)   )  THEN 
     --     
     --     See Also      : RegLessThan, RegLessThanOrEqual,RegGreaterThanOrEqual.
     -------------------------------------------------------------------------------
     FUNCTION RegGreaterThan  ( CONSTANT l          : IN std_logic_vector;
				CONSTANT r          : IN std_logic_vector;
				CONSTANT SrcRegMode : IN regmode_type 
                     -- synopsys synthesis_off
							      := DefaultRegMode 
                     -- synopsys synthesis_on
				 ) RETURN std_ulogic;
     -----------------------------------------------------------------------------
     FUNCTION RegGreaterThan    ( CONSTANT l          : IN std_logic_vector;
				   CONSTANT r          : IN std_logic_vector;
 			           CONSTANT SrcRegMode : IN regmode_type
                     -- synopsys synthesis_off
							      := DefaultRegMode 
                     -- synopsys synthesis_on
				 ) RETURN BOOLEAN;
     -- -----------------------------------------------------------------------------
     FUNCTION RegGreaterThan ( CONSTANT l          : IN std_logic_vector;
				   CONSTANT r          : IN INTEGER;
			     CONSTANT SrcRegMode : IN regmode_type
                     -- synopsys synthesis_off
						      := DefaultRegMode 
                     -- synopsys synthesis_on
				 ) RETURN BOOLEAN;
     -------------------------------------------------------------------------------
     FUNCTION RegGreaterThan ( CONSTANT l          : IN INTEGER;
				   CONSTANT r          : IN std_logic_vector;
  			           CONSTANT SrcRegMode : IN regmode_type
                     -- synopsys synthesis_off
					         	      := DefaultRegMode 
                     -- synopsys synthesis_on
				 ) RETURN BOOLEAN;
     -------------------------------------------------------------------------------
     FUNCTION RegGreaterThan ( CONSTANT l          : IN std_logic_vector;
				   CONSTANT r          : IN INTEGER;
  			           CONSTANT SrcRegMode : IN regmode_type
                     -- synopsys synthesis_off
					         	      := DefaultRegMode 
                     -- synopsys synthesis_on
				 ) RETURN std_ulogic;
     -------------------------------------------------------------------------------
     FUNCTION RegGreaterThan ( CONSTANT l          : IN INTEGER;
				   CONSTANT r          : IN std_logic_vector;
  			           CONSTANT SrcRegMode : IN regmode_type
                     -- synopsys synthesis_off
					         	      := DefaultRegMode 
                     -- synopsys synthesis_on
				 ) RETURN std_ulogic;
     -- ----------------------------------------------------------------------------
     --     Function Name : RegGreaterThan
     --
     --     Overloading   : Input parameter TYPEs.
     --    
     --     Purpose       : Compute a greater than relation for std_logic_vectors
     --     
     --     Parameters    : l       - input std_ulogic_vector | INTEGER
     --                     r       - input std_ulogic_vector | INTEGER
     --                     SrcRegMode - input regmode_type, indicating the format of
     --                               the std_ulogic_vector operands (l,r).
     --                               Default is TwosComp.
     --     
     --     Result        : BOOLEAN | std_ulogic
     --
     --     NOTE          : The operands may be of any length, and may be different
     --                     lengths. 
     --
     --                     Overloading not defined for both inputs of INTEGER type.
     --
     --                     Any time the comparison reaches an index that has an 'X' as an
     --                     array element, the comparison is deemed indeterminate and will 
     --                     return false in case of boolean and '0' incase of 
     --                     std_ulogic for synthesis purposes.
     --     Use           : 
     --                      VARIABLE a, b : std_ulogic_vector ( 7 DOWNTO 0 );
     --                      IF ( RegGreaterThan ( a, b, TwosComp)   )  THEN 
     --     
     --     See Also      : RegLessThan, RegLessThanOrEqual, RegGreaterThanOrEqual.
     -------------------------------------------------------------------------------
     FUNCTION RegGreaterThan  ( CONSTANT l          : IN std_ulogic_vector;
				CONSTANT r          : IN std_ulogic_vector;
				CONSTANT SrcRegMode : IN regmode_type 
                     -- synopsys synthesis_off
							      := DefaultRegMode 
                     -- synopsys synthesis_on
				 ) RETURN std_ulogic;
     -----------------------------------------------------------------------------
     FUNCTION RegGreaterThan    ( CONSTANT l          : IN std_ulogic_vector;
				   CONSTANT r          : IN std_ulogic_vector;
 			           CONSTANT SrcRegMode : IN regmode_type
                     -- synopsys synthesis_off
							      := DefaultRegMode 
                     -- synopsys synthesis_on
				 ) RETURN BOOLEAN;
     -- -----------------------------------------------------------------------------
     FUNCTION RegGreaterThan ( CONSTANT l          : IN std_ulogic_vector;
				   CONSTANT r          : IN INTEGER;
			     CONSTANT SrcRegMode : IN regmode_type
                     -- synopsys synthesis_off
						      := DefaultRegMode 
                     -- synopsys synthesis_on
				 ) RETURN BOOLEAN;
     -------------------------------------------------------------------------------
     FUNCTION RegGreaterThan ( CONSTANT l          : IN INTEGER;
				   CONSTANT r          : IN std_ulogic_vector;
  			           CONSTANT SrcRegMode : IN regmode_type
                     -- synopsys synthesis_off
					         	      := DefaultRegMode 
                     -- synopsys synthesis_on
				 ) RETURN BOOLEAN;
     -------------------------------------------------------------------------------
     FUNCTION RegGreaterThan ( CONSTANT l          : IN std_ulogic_vector;
				   CONSTANT r          : IN INTEGER;
  			           CONSTANT SrcRegMode : IN regmode_type
                     -- synopsys synthesis_off
					         	      := DefaultRegMode 
                     -- synopsys synthesis_on
				 ) RETURN std_ulogic;
     -------------------------------------------------------------------------------
     FUNCTION RegGreaterThan ( CONSTANT l          : IN INTEGER;
			       CONSTANT r          : IN std_ulogic_vector;
  			       CONSTANT SrcRegMode : IN regmode_type
                     -- synopsys synthesis_off
					         	      := DefaultRegMode 
                     -- synopsys synthesis_on
				 ) RETURN std_ulogic;
     -------------------------------------------------------------------------------
     --     Function Name : RegGreaterThanOrEqual
     -- 1.2.53
     --     Overloading   : Input parameter TYPEs.
     --
     --     Purpose       : Compute a greater-than-or-equal relation for bit_vectors
     --
     --     Parameters    : l       - input bit_vector | INTEGER
     --                     r       - input bit_vector | INTEGER
     --                     SrcRegMode - input regmode_type, indicating the format of
     --                               the bit_vector operands (l,r).
     --                               Default is TwosComp.
     --
     --     Result        : BOOLEAN | bit
     --
     --     NOTE          : The operands may be of any length, and may be different
     --                     lengths.
     --
     --                     Overloading not defined for both inputs of INTEGER type.
     --     Use           :
     --                      VARIABLE a, b : bit_vector ( 7 DOWNTO 0 );
     --                      IF ( RegGreaterThanOrEqual ( a, b, TwosComp)   )  THEN
     --
     --     See Also      : RegLessThan, RegLessThanOrEqual, RegGreaterThan,
     -------------------------------------------------------------------------------
     FUNCTION RegGreaterThanOrEqual ( CONSTANT l          : IN bit_vector;
			       CONSTANT r          : IN bit_vector;
		               CONSTANT SrcRegMode : IN regmode_type
                     -- synopsys synthesis_off
							      := DefaultRegMode 
                     -- synopsys synthesis_on
				 ) RETURN bit;
     -----------------------------------------------------------------------------
     FUNCTION RegGreaterThanOrEqual    ( CONSTANT l          : IN bit_vector;
				   CONSTANT r          : IN bit_vector;
 			           CONSTANT SrcRegMode : IN regmode_type
                     -- synopsys synthesis_off
							      := DefaultRegMode 
                     -- synopsys synthesis_on
				 ) RETURN BOOLEAN;
     -- -----------------------------------------------------------------------------
     FUNCTION RegGreaterThanOrEqual ( CONSTANT l          : IN bit_vector;
				   CONSTANT r          : IN INTEGER;
			     CONSTANT SrcRegMode : IN regmode_type
                     -- synopsys synthesis_off
						      := DefaultRegMode 
                     -- synopsys synthesis_on
				 ) RETURN BOOLEAN;
     -------------------------------------------------------------------------------
     FUNCTION RegGreaterThanOrEqual ( CONSTANT l          : IN INTEGER;
				   CONSTANT r          : IN bit_vector;
  			           CONSTANT SrcRegMode : IN regmode_type
                     -- synopsys synthesis_off
					         	      := DefaultRegMode 
                     -- synopsys synthesis_on
				 ) RETURN BOOLEAN;
     -------------------------------------------------------------------------------
     FUNCTION RegGreaterThanOrEqual ( CONSTANT l          : IN bit_vector;
				   CONSTANT r          : IN INTEGER;
  			           CONSTANT SrcRegMode : IN regmode_type
                     -- synopsys synthesis_off
							      := DefaultRegMode 
                     -- synopsys synthesis_on
				 ) RETURN bit;
     -------------------------------------------------------------------------------
     FUNCTION RegGreaterThanOrEqual ( CONSTANT l          : IN INTEGER;
 				   CONSTANT r          : IN bit_vector;
  			           CONSTANT SrcRegMode : IN regmode_type
                     -- synopsys synthesis_off
					         	      := DefaultRegMode 
                     -- synopsys synthesis_on
				 ) RETURN bit;
     -- ----------------------------------------------------------------------------
     --     Function Name : RegGreaterThanOrEqual
     --
     --     Overloading   : Input parameter TYPEs.
     --    
     --     Purpose       : Compute a greater-than-or-equal relation for std_logic_vectors
     --     
     --     Parameters    : l       - input std_logic_vector | INTEGER
     --                     r       - input std_logic_vector | INTEGER
     --                     SrcRegMode - input regmode_type, indicating the format of
     --                               the std_logic_vector operands (l,r).
     --                               Default is TwosComp.
     --     
     --     Result        : BOOLEAN | std_ulogic
     --
     --     NOTE          : The operands may be of any length, and may be different
     --                     lengths. 
     --
     --                     Overloading not defined for both inputs of INTEGER type.
     --
     --                     Any time the comparison reaches an index that has an 'X' as an
     --                     array element, the comparison is deemed indeterminate and will 
     --                     return false in case of boolean and '0' incase of 
     --                     std_ulogic for synthesis purposes.
     --     Use           : 
     --                      VARIABLE a, b : std_logic_vector ( 7 DOWNTO 0 );
     --                      IF ( RegGreaterThanOrEqual ( a, b, TwosComp)   )  THEN 
     --     
     --     See Also      : RegLessThan, RegLessThanOrEqual, RegGreaterThan, 
     -------------------------------------------------------------------------------
     FUNCTION RegGreaterThanOrEqual  ( CONSTANT l          : IN std_logic_vector;
				CONSTANT r          : IN std_logic_vector;
				CONSTANT SrcRegMode : IN regmode_type 

                     -- synopsys synthesis_off
							      := DefaultRegMode 
                     -- synopsys synthesis_on
				 ) RETURN std_ulogic;
     -----------------------------------------------------------------------------
     FUNCTION RegGreaterThanOrEqual    ( CONSTANT l          : IN std_logic_vector;
   				         CONSTANT r          : IN std_logic_vector;
 			                 CONSTANT SrcRegMode : IN regmode_type
                     -- synopsys synthesis_off
							      := DefaultRegMode 
                     -- synopsys synthesis_on
				       ) RETURN BOOLEAN;
     -- -----------------------------------------------------------------------------
     FUNCTION RegGreaterThanOrEqual ( CONSTANT l          : IN std_logic_vector;
				      CONSTANT r          : IN INTEGER;
			              CONSTANT SrcRegMode : IN regmode_type
                     -- synopsys synthesis_off
						      := DefaultRegMode 
                     -- synopsys synthesis_on
				    ) RETURN BOOLEAN;
     -------------------------------------------------------------------------------
     FUNCTION RegGreaterThanOrEqual ( CONSTANT l          : IN INTEGER;
				      CONSTANT r          : IN std_logic_vector;
  			              CONSTANT SrcRegMode : IN regmode_type
                     -- synopsys synthesis_off
					         	      := DefaultRegMode 
                     -- synopsys synthesis_on
				    ) RETURN BOOLEAN;
     -------------------------------------------------------------------------------
     FUNCTION RegGreaterThanOrEqual ( CONSTANT l          : IN std_logic_vector;
				      CONSTANT r          : IN INTEGER;
  			              CONSTANT SrcRegMode : IN regmode_type
                     -- synopsys synthesis_off
					         	      := DefaultRegMode 
                     -- synopsys synthesis_on
				    ) RETURN std_ulogic;
     -------------------------------------------------------------------------------
     FUNCTION RegGreaterThanOrEqual ( CONSTANT l          : IN INTEGER;
				      CONSTANT r          : IN std_logic_vector;
  			              CONSTANT SrcRegMode : IN regmode_type
                     -- synopsys synthesis_off
					         	      := DefaultRegMode 
                     -- synopsys synthesis_on
				    ) RETURN std_ulogic;
     -- ----------------------------------------------------------------------------
     --     Function Name : RegGreaterThanOrEqual
     --
     --     Overloading   : Input parameter TYPEs.
     --    
     --     Purpose       : Compute a greater-than-or-equal relation for std_ulogic_vectors
     --     
     --     Parameters    : l       - input std_ulogic_vector | INTEGER
     --                     r       - input std_ulogic_vector | INTEGER
     --                     SrcRegMode - input regmode_type, indicating the format of
     --                               the std_ulogic_vector operands (l,r).
     --                               Default is TwosComp.
     --     
     --     Result        : BOOLEAN | std_ulogic
     --
     --     NOTE          : The operands may be of any length, and may be different
     --                     lengths. 
     --
     --                     Overloading not defined for both inputs of INTEGER type.
     --
     --                     Any time the comparison reaches an index that has an 'X' as an
     --                     array element, the comparison is deemed indeterminate and will 
     --                     return false in case of boolean and '0' incase of 
     --                     std_ulogic for synthesis purposes.
     --     Use           : 
     --                      VARIABLE a, b : std_ulogic_vector ( 7 DOWNTO 0 );
     --                      IF ( RegGreaterThanOrEqual ( a, b, TwosComp)   )  THEN 
     --     
     --     See Also      : RegLessThan, RegLessThanOrEqual, RegGreaterThan, 
     -------------------------------------------------------------------------------
     FUNCTION RegGreaterThanOrEqual  ( CONSTANT l          : IN std_ulogic_vector;
				       CONSTANT r          : IN std_ulogic_vector;
				       CONSTANT SrcRegMode : IN regmode_type 
                     -- synopsys synthesis_off
							      := DefaultRegMode 
                     -- synopsys synthesis_on
             			     ) RETURN std_ulogic;
     -----------------------------------------------------------------------------
     FUNCTION RegGreaterThanOrEqual  ( CONSTANT l          : IN std_ulogic_vector;
				       CONSTANT r          : IN std_ulogic_vector;
 			               CONSTANT SrcRegMode : IN regmode_type
                     -- synopsys synthesis_off
							      := DefaultRegMode 
                     -- synopsys synthesis_on
				     ) RETURN BOOLEAN;
     -- -----------------------------------------------------------------------------
     FUNCTION RegGreaterThanOrEqual ( CONSTANT l          : IN std_ulogic_vector;
				   CONSTANT r          : IN INTEGER;
			     CONSTANT SrcRegMode : IN regmode_type
                     -- synopsys synthesis_off
						      := DefaultRegMode 
                     -- synopsys synthesis_on
				 ) RETURN BOOLEAN;
     -------------------------------------------------------------------------------
     FUNCTION RegGreaterThanOrEqual ( CONSTANT l          : IN INTEGER;
				      CONSTANT r          : IN std_ulogic_vector;
  			              CONSTANT SrcRegMode : IN regmode_type
                     -- synopsys synthesis_off
					         	      := DefaultRegMode 
                     -- synopsys synthesis_on
				    ) RETURN BOOLEAN;
     -------------------------------------------------------------------------------
     FUNCTION RegGreaterThanOrEqual ( CONSTANT l          : IN std_ulogic_vector;
				      CONSTANT r          : IN INTEGER;
  			              CONSTANT SrcRegMode : IN regmode_type
                     -- synopsys synthesis_off
					         	      := DefaultRegMode 
                     -- synopsys synthesis_on
				    ) RETURN std_ulogic;
     -------------------------------------------------------------------------------
     FUNCTION RegGreaterThanOrEqual ( CONSTANT l          : IN INTEGER;
				      CONSTANT r          : IN std_ulogic_vector;
  			              CONSTANT SrcRegMode : IN regmode_type
                     -- synopsys synthesis_off
					         	      := DefaultRegMode 
                     -- synopsys synthesis_on
				   ) RETURN std_ulogic;

end synth_regpak;
--
--
--
Package body synth_regpak is
-- synopsys synthesis_off
     CONSTANT max_string_len : INTEGER := 256;  -- for To_String

     TYPE map01   IS ARRAY(BIT, BIT) OF BIT;
     TYPE X01map2  IS ARRAY(std_ulogic, std_ulogic ) OF X01;

     CONSTANT tbl_lt : X01map2 := (
    --      ---------------------------------------------------------
    --      |  U    X    0    1    Z    W    L    H    -        |   |  
    --      ---------------------------------------------------------
            ( 'X', 'X', 'X', 'X', 'X', 'X', 'X', 'X', 'X' ), -- | U |
            ( 'X', 'X', 'X', 'X', 'X', 'X', 'X', 'X', 'X' ), -- | X |
            ( 'X', 'X', '0', '1', 'X', 'X', '0', '1', 'X' ), -- | 0 |
            ( 'X', 'X', '0', '0', 'X', 'X', '0', '0', 'X' ), -- | 1 |
            ( 'X', 'X', 'X', 'X', 'X', 'X', 'X', 'X', 'X' ), -- | Z |
            ( 'X', 'X', 'X', 'X', 'X', 'X', 'X', 'X', 'X' ), -- | W |
            ( 'X', 'X', '0', '1', 'X', 'X', '0', '1', 'X' ), -- | L |
            ( 'X', 'X', '0', '0', 'X', 'X', '0', '0', 'X' ), -- | H |
            ( 'X', 'X', 'X', 'X', 'X', 'X', 'X', 'X', 'X' )  -- | - |
        );

     CONSTANT tbl_eq : X01map2 := (
    --      ---------------------------------------------------------
    --      |  U    X    0    1    Z    W    L    H    -        |   |  
    --      ---------------------------------------------------------
            ( 'X', 'X', 'X', 'X', 'X', 'X', 'X', 'X', 'X' ), -- | U |
            ( 'X', 'X', 'X', 'X', 'X', 'X', 'X', 'X', 'X' ), -- | X |
            ( 'X', 'X', '1', '0', 'X', 'X', '1', '0', 'X' ), -- | 0 |
            ( 'X', 'X', '0', '1', 'X', 'X', '0', '1', 'X' ), -- | 1 |
            ( 'X', 'X', 'X', 'X', 'X', 'X', 'X', 'X', 'X' ), -- | Z |
            ( 'X', 'X', 'X', 'X', 'X', 'X', 'X', 'X', 'X' ), -- | W |
            ( 'X', 'X', '1', '0', 'X', 'X', '1', '0', 'X' ), -- | L |
            ( 'X', 'X', '0', '1', 'X', 'X', '0', '1', 'X' ), -- | H |
            ( 'X', 'X', 'X', 'X', 'X', 'X', 'X', 'X', 'X' )  -- | - |
        );

     CONSTANT tbl_lt_bit : map01 := (  '0' => ( '0' => '0', '1' => '1'),
      		         	     '1' => ( '0' => '0', '1' => '0') );

     CONSTANT tbl_eq_bit : map01 := ( '0' => ( '0' => '1', '1' => '0'),
				    '1' => ( '0' => '0', '1' => '1'));

-- synopsys synthesis_on
-- -----------------------------------------------------------------------------------
-- ----------------------------------------------------------------------------------
--        L O C A L   F U N C T I O N S   AND   P R O C E D U R E S
-- ----------------------------------------------------------------------------------
-- ----------------------------------------------------------------------------------
--    
     ---------------------------------------------------------------------------------
     --     Function Name  : MAXIMUM
     -- hidden
     --     Overloading    :
     --
     --     Purpose        : To determine the max of two inetgers
     --
     --     Parameters     : i1    - input  integer
     --                      i2    - input integer
     --
     --     Result        : Integer, max of i1 , i2
     --
     -- ------------------------------------------------------------------------------
     FUNCTION MAXIMUM  ( CONSTANT i1 : IN INTEGER;
			 CONSTANT i2 : IN INTEGER
		       ) RETURN INTEGER IS
     BEGIN
	IF i1 < i2 THEN 
	   RETURN i2; 
        ELSE 
           RETURN i1;
	END IF;
     END MAXIMUM;
     ---------------------------------------------------------------------------------
     --     Function Name  : MINIMUM
     -- hidden
     --     Overloading    :
     --
     --     Purpose        : To determine the min of two inetgers
     --
     --     Parameters     : i1    - input  integer
     --                      i2    - input integer
     --
     --     Result        : Integer, min of i1 , i2
     --
     -- ------------------------------------------------------------------------------
     FUNCTION MINIMUM  ( CONSTANT i1 : IN INTEGER;
			 CONSTANT i2 : IN INTEGER
		       ) RETURN INTEGER IS
     BEGIN
	IF i1 > i2 THEN 
	    RETURN i2; 
        ELSE
            RETURN i1;
	END IF;
     END MINIMUM;

     -- ------------------------------------------------------------------------------
     FUNCTION All_Zero   ( CONSTANT bv : IN bit_vector
                 	 ) RETURN boolean IS
	VARIABLE bv_copy : BIT_VECTOR(bv'LENGTH -1 DOWNTO 0);
	VARIABLE result  : BOOLEAN;
     BEGIN
	bv_copy := bv;
        result  := TRUE;
	convt_loop: FOR I in bv'LENGTH - 1 DOWNTO 0 LOOP
		IF (bv_copy(i) /= '0') THEN
			result := FALSE;
--			EXIT convt_loop;
			return result;
		END IF;
 	end LOOP convt_loop;
	return result;
     END All_Zero;
     -- ------------------------------------------------------------------------------
     FUNCTION All_Zero   ( CONSTANT sv : IN std_logic_vector
                 	 ) RETURN boolean IS
	VARIABLE sv_copy : std_logic_vector(sv'LENGTH -1 DOWNTO 0);
	VARIABLE result  : BOOLEAN;
     BEGIN
	sv_copy := sv;
        result  := TRUE;
	convt_loop: FOR I in sv'LENGTH - 1 DOWNTO 0 LOOP
		IF (sv_copy(i) /= '0') THEN
			result := FALSE;
--			EXIT convt_loop;
			return result;
		END IF;
 	end LOOP convt_loop;
	return result;
     END All_Zero;
     -- ------------------------------------------------------------------------------
     FUNCTION All_Zero   ( CONSTANT sv : IN std_ulogic_vector
                 	 ) RETURN boolean IS
	VARIABLE sv_copy : std_ulogic_vector(sv'LENGTH -1 DOWNTO 0);
	VARIABLE result  : BOOLEAN;
     BEGIN
	sv_copy := sv;
        result  := TRUE;
	convt_loop: FOR I in sv'LENGTH - 1 DOWNTO 0 LOOP
		IF (sv_copy(i) /= '0') THEN
			result := FALSE;
--			EXIT convt_loop;
			return result;
		END IF;
 	end LOOP convt_loop;
	return result;
     END All_Zero;
     -- ------------------------------------------------------------------------------
     -- return true if no one ecnountered 
     -- false otherwise
     FUNCTION No_One   ( CONSTANT bv : IN bit_vector
                 	 ) RETURN boolean IS
	VARIABLE bv_copy : bit_vector(bv'LENGTH -1 DOWNTO 0);
	VARIABLE result  : BOOLEAN;
     BEGIN
        bv_copy := bv;
        result := TRUE;
	convt_loop: FOR I in bv'LENGTH - 1 DOWNTO 0 LOOP
		IF (bv_copy(i) = '1') THEN
			result := FALSE;
--			EXIT convt_loop;
			return result;
		END IF;
 	end LOOP convt_loop;
	return result;
     END No_One;
     -- ------------------------------------------------------------------------------
     -- return true if no one ecnountered 
     -- false otherwise
     FUNCTION No_One   ( CONSTANT sv : IN std_logic_vector
                 	 ) RETURN boolean IS
	VARIABLE sv_copy : std_logic_vector(sv'LENGTH -1 DOWNTO 0);
	VARIABLE result  : BOOLEAN;
     BEGIN
        sv_copy := sv;
        result := TRUE;
	convt_loop: FOR I in sv'LENGTH - 1 DOWNTO 0 LOOP
		IF (sv_copy(i) = '1') THEN
			result := FALSE;
--			EXIT convt_loop;
			return result;	
		END IF;
 	end LOOP convt_loop;
	return result;
     END No_One;
     -- ------------------------------------------------------------------------------
     -- return true if no one ecnountered 
     -- false otherwise
     FUNCTION No_One   ( CONSTANT sv : IN std_ulogic_vector
                 	 ) RETURN boolean IS
	VARIABLE sv_copy : std_ulogic_vector(sv'LENGTH -1 DOWNTO 0);
	VARIABLE result  : BOOLEAN;
     BEGIN
        sv_copy := sv;
        result := TRUE;
	convt_loop: FOR I in sv'LENGTH - 1 DOWNTO 0 LOOP
		IF (sv_copy(i) = '1') THEN
			result := FALSE;
--			EXIT convt_loop;
			return result;
		END IF;
 	end LOOP convt_loop;
	return result;
     END No_One;
     -------------------------------------------------------------------------------
     --     Function Name  : To_Bit_loc
     -- hidden
     --     Overloading    : 
     --
     --     Purpose        : Translate  a  boolean into a bit .
     --
     --     Parameters     :  b    - input  boolean value to be translated.
     --
     --     Result        : bit,
     --
     --     Use            :
     --                      VARIABLE  lt : bit ;
     --                      VARIABLE  ok : boolean := true;
     --
     --                        lt := To_Bit_loc(ok);
     -- ------------------------------------------------------------------------------
     FUNCTION To_Bit_loc ( b:boolean
		      ) RETURN bit IS
     BEGIN
	if (b = true) then
		return('1');
        else 
		return ('0');
        end if;

     END To_Bit_loc;
     -------------------------------------------------------------------------------
     --     Function Name  : To_StdUlogic_loc
     -- hidden
     --     Overloading    : 
     --
     --     Purpose        : Translate  a  boolean into an std_ulogic .
     --
     --     Parameters     :  b    - input  boolean value to be translated.
     --
     --     Result        : std_ulogic,
     --
     --     Use            :
     --                      VARIABLE  lt : std_ulogic ;
     --                      VARIABLE  ok : boolean := true;
     --
     --                        lt := To_StdULogic_loc(ok);
     -- ------------------------------------------------------------------------------
     FUNCTION To_StdUlogic_loc ( b:boolean
             		       ) RETURN std_ulogic IS
     BEGIN
	if (b = true) then
		return('1');
        else 
		return ('0');
        end if;

     END To_StdUlogic_loc;
 --+-----------------------------------------------------------------------------
 --|     Procedure Name : Return_Boolean_TwosComp
 --|  hidden
 --|     Overloading    :
 --|     Purpose        :boolean type propagation function.
 --|
 --|     Parameters     :
 --|                      A          - input  BIT_VECTOR 
 --|                      B          - input  BIT_VECTOR 
 --|
 --|     Result         : Boolean
 --|-----------------------------------------------------------------------------
     FUNCTION Return_Boolean_TwosComp   ( CONSTANT A       : IN  BIT_VECTOR;
			                  CONSTANT B       : IN  BIT_VECTOR
			               )  return BOOLEAN IS
	variable Z:Boolean;       
	-- pragma return_port_name Z     
     BEGIN
	return(Z);
     END Return_Boolean_TwosComp;		        
 --+-----------------------------------------------------------------------------
 --|     Procedure Name : Return_Boolean_TwosComp
 --|  hidden
 --|     Overloading    :
 --|     Purpose        :boolean type propagation function.
 --|
 --|     Parameters     :
 --|                      A          - input  STD_LOGIC_VECTOR 
 --|                      B          - input  STD_LOGIC_VECTOR 
 --|
 --|     Result         : Boolean
 --|-----------------------------------------------------------------------------
     FUNCTION Return_Boolean_TwosComp   ( CONSTANT A     : IN  STD_LOGIC_VECTOR;
			                  CONSTANT B     : IN  STD_LOGIC_VECTOR
			                ) return BOOLEAN IS
	variable Z:Boolean;       
	-- pragma return_port_name Z     
     BEGIN
	return(Z);
     END Return_Boolean_TwosComp;		        
 --+-----------------------------------------------------------------------------
 --|     Procedure Name : Return_Boolean_TwosComp
 --|  hidden
 --|     Overloading    :
 --|     Purpose        :boolean type propagation function.
 --|
 --|     Parameters     :
 --|                      A          - input  STD_ULOGIC_VECTOR 
 --|                      B          - input  STD_ULOGIC_VECTOR 
 --|
 --|     Result         : Boolean
 --|-----------------------------------------------------------------------------
     FUNCTION Return_Boolean_TwosComp    ( CONSTANT A     : IN  STD_ULOGIC_VECTOR;
			                   CONSTANT B     : IN  STD_ULOGIC_VECTOR
			                 ) return BOOLEAN IS
	variable Z:Boolean;       
	-- pragma return_port_name Z     
     BEGIN
	return(Z);
     END Return_Boolean_TwosComp;		        
 --+-----------------------------------------------------------------------------
 --|     Procedure Name : Return_Boolean_Unsigned
 --|  hidden
 --|     Overloading    :
 --|     Purpose        :boolean type propagation function.
 --|
 --|     Parameters     :
 --|                      A          - input  BIT_VECTOR 
 --|                      B          - input  BIT_VECTOR 
 --|
 --|     Result         : Boolean
 --|-----------------------------------------------------------------------------
     FUNCTION Return_Boolean_Unsigned    ( CONSTANT A      : IN  BIT_VECTOR;
			                   CONSTANT B      : IN  BIT_VECTOR
			                 ) return BOOLEAN IS
	variable Z:Boolean;       
	-- pragma return_port_name Z     
     BEGIN
	return(Z);
     END Return_Boolean_Unsigned;		        
 --+-----------------------------------------------------------------------------
 --|     Procedure Name : Return_Boolean_Unsigned
 --|  hidden
 --|     Overloading    :
 --|     Purpose        :boolean type propagation function.
 --|
 --|     Parameters     :
 --|                      A          - input  STD_LOGIC_VECTOR 
 --|                      B          - input  STD_LOGIC_VECTOR 
 --|
 --|     Result         : Boolean
 --|-----------------------------------------------------------------------------
     FUNCTION Return_Boolean_Unsigned   ( CONSTANT A     : IN  STD_LOGIC_VECTOR;
			                  CONSTANT B     : IN  STD_LOGIC_VECTOR
			                ) return BOOLEAN IS
	variable Z:Boolean;       
	-- pragma return_port_name Z     
     BEGIN
	return(Z);
     END Return_Boolean_Unsigned;		        
 --+-----------------------------------------------------------------------------
 --|     Procedure Name : Return_Boolean_Unsigned
 --|  hidden
 --|     Overloading    :
 --|     Purpose        :boolean type propagation function.
 --|
 --|     Parameters     :
 --|                      A          - input  STD_ULOGIC_VECTOR 
 --|                      B          - input  STD_ULOGIC_VECTOR 
 --|
 --|     Result         : Boolean
 --|-----------------------------------------------------------------------------
     FUNCTION Return_Boolean_Unsigned    ( CONSTANT A    : IN  STD_ULOGIC_VECTOR;
			                   CONSTANT B    : IN  STD_ULOGIC_VECTOR
			                 ) return BOOLEAN IS
	variable Z:Boolean;       
	-- pragma return_port_name Z     
     BEGIN
	return(Z);
     END Return_Boolean_Unsigned;		        
 --+-----------------------------------------------------------------------------
 --|     Procedure Name : LessThan_TwosComp
 --|  hidden
 --|     Overloading    :
 --|
 --|     Purpose        : Compute the relation less than  for BIT_VECTORS.
 --|
 --|     Parameters     :
 --|                      A          - input  BIT_VECTOR 
 --|                      B          - input  BIT_VECTOR 
 --|
 --|     NOTE           : The operands must be of same Aength with mode TwosComp.
 --|
 --|     Assumptions    : Both inputs must have range (msb downto 0)
 --|
 --|     Result         : Boolean
 --|
 --|     Use            :
 --|                      VARIABLE a, b : BIT_VECTOR ( 7 DOWNTO 0 );
 --|                      VARIABLE lt : boolean;
 --|                      lt := LessThan_TwosComp (l, r );
 --|
 --|-----------------------------------------------------------------------------
     FUNCTION LessThan_TwosComp    ( CONSTANT A        : IN  BIT_VECTOR;
			             CONSTANT B        : IN  BIT_VECTOR
			          )  return BOOLEAN IS
       VARIABLE vl       : bit_vector (A'length - 1 downto 0);
       VARIABLE vr       : bit_vector (B'length - 1 downto 0);
       VARIABLE indx     : INTEGER;       
	-- pragma map_to_operator LT_TC_OP
	-- pragma type_function Return_Boolean_TwosComp         
	-- pragma return_port_name Z
     BEGIN
	-- synopsys synthesis_off
        vl := A;
        vr := B;
       -- complement the sign bit
	vl(A'length - 1) := NOT vl(A'length - 1);
	vr(B'length - 1) := NOT vr(B'length - 1);
       -- perform comparison in a short circuit fashion
       -- Find the most significant differing bit : If equal use LSB
	 FOR i IN A'length - 1 DOWNTO 0 LOOP
	   indx := i;
--	   EXIT WHEN  vl(i) /= vr(i) ; 
		if (vl(i) /= vr(i)) then
			return ( tbl_lt_bit ( vl(indx), vr(indx) ) = '1');
		end if;
	 END LOOP;
     -- Compute the relationships based on the value of the differing bit
--	 return ( tbl_lt_bit ( vl(indx), vr(indx) ) = '1');
		return FALSE;
	-- synopsys synthesis_on
     END LessThan_TwosComp;
 --+-----------------------------------------------------------------------------
 --|     Procedure Name : LessThan_TwosComp
 --|  hidden
 --|     Overloading    :
 --|
 --|     Purpose        : Compute the relation less than  for STD_LOGIC_VECTORS.
 --|
 --|     Parameters     :
 --|                      A          - input  STD_LOGIC_VECTOR 
 --|                      B          - input  STD_LOGIC_VECTOR 
 --|
 --|     NOTE           : The operands must be of same Aength with mode TwosComp.
 --|                     
 --|                      Any time the comparison reaches an index that has an 'X' as an
 --|                      array element, the comparison is deemed indeterminate and  
 --|                      will return boolean false.
 --|
 --|     Assumptions    : Both inputs must have range (msb downto 0)
 --|
 --|     Result         : Boolean
 --|
 --|     Use            : VARIABLE a, b : STD_LOGIC_VECTOR ( 7 DOWNTO 0 );
 --|                      VARIABLE lt : boolean;
 --|                      lt := LessThan_TwosComp (l, r );
 --|-----------------------------------------------------------------------------
     FUNCTION LessThan_TwosComp      ( CONSTANT A       : IN  STD_LOGIC_VECTOR;
			               CONSTANT B       : IN  STD_LOGIC_VECTOR
			             ) return BOOLEAN IS
       VARIABLE vl       : std_logic_vector (A'length - 1 downto 0);
       VARIABLE vr       : std_logic_vector (B'length - 1 downto 0);
       VARIABLE indx     : INTEGER;       
	-- pragma map_to_operator LT_TC_OP
	-- pragma type_function Return_Boolean_TwosComp         
	-- pragma return_port_name Z
     BEGIN
	-- synopsys synthesis_off
        vl := A;
        vr := B;
       -- complement the sign bit
	vl(A'length - 1) := NOT vl(A'length - 1);
	vr(B'length - 1) := NOT vr(B'length - 1);
       -- perform comparison in a short circuit fashion
       -- Find the most significant differing bit : If equal use LSB
	 FOR i IN A'length - 1 DOWNTO 0 LOOP
	   indx := i;
--	   EXIT WHEN ( vl(i) /= vr(i) OR vl(i) = 'X' OR vr(i) = 'X');
		if( vl(i) /= vr(i) OR vl(i) = 'X' OR vr(i) = 'X')then
			if (vl(indx) = 'X' OR vr(indx) = 'X') Then
				ASSERT NOT WarningsOn
					REPORT "  --- Comparison is indeterminate will return " &
						" false in case of boolean and '0' in case of std_ulogic "
					SEVERITY WARNING;
			END IF;
			-- Compute the relationships based on the value of the differing bit
			return ( tbl_lt ( vl(indx), vr(indx) ) = '1');
		end if;
	 END LOOP;
--	if (vl(indx) = 'X' OR vr(indx) = 'X') Then
--	    ASSERT NOT WarningsOn
--	    REPORT "  --- Comparison is indeterminate will return " &
--		   " false in case of boolean and '0' in case of std_ulogic "
--	    SEVERITY WARNING;
--	 END IF;
       -- Compute the relationships based on the value of the differing bit
--	 return ( tbl_lt ( vl(indx), vr(indx) ) = '1');
		return FALSE;
       -- synopsys synthesis_on
     END LessThan_TwosComp;
 --+-----------------------------------------------------------------------------
 --|     Procedure Name : LessThan_TwosComp
 --|  hidden
 --|     Overloading    :
 --|
 --|     Purpose        : Compute the relation less than  for STD_ULOGIC_VECTORS.
 --|
 --|     Parameters     :
 --|                      A          - input  STD_ULOGIC_VECTOR 
 --|                      B          - input  STD_ULOGIC_VECTOR 
 --|
 --|     NOTE           : The operands must be of same Aength with mode TwosComp.
 --|                     
 --|                      Any time the comparison reaches an index that has an 'X' as an
 --|                      array element, the comparison is deemed indeterminate and will 
 --|                      return boolean false.
 --|
 --|     Assumptions    : Both inputs must have range (msb downto 0)
 --|
 --|     Result         : Boolean
 --|
 --|     Use            : VARIABLE a, b : STD_ULOGIC_VECTOR ( 7 DOWNTO 0 );
 --|                      VARIABLE lt : boolean;
 --|                      lt := LessThan_TwosComp (l, r );
 --|-----------------------------------------------------------------------------
     FUNCTION LessThan_TwosComp    ( CONSTANT A         : IN  STD_ULOGIC_VECTOR;
			             CONSTANT B         : IN  STD_ULOGIC_VECTOR
			           ) return BOOLEAN IS
       VARIABLE vl       : std_ulogic_vector (A'length - 1 downto 0);
       VARIABLE vr       : std_ulogic_vector (B'length - 1 downto 0);
       VARIABLE indx     : INTEGER;       
	-- pragma map_to_operator LT_TC_OP
	-- pragma type_function Return_Boolean_TwosComp         
	-- pragma return_port_name Z
     BEGIN
	-- synopsys synthesis_off
        vl := A;
        vr := B;
       -- complement the sign bit
	vl(A'length - 1) := NOT vl(A'length - 1);
	vr(B'length - 1) := NOT vr(B'length - 1);
       -- perform comparison in a short circuit fashion
       -- Find the most significant differing bit : If equal use LSB
	 FOR i IN A'length - 1 DOWNTO 0 LOOP
	   indx := i;
--	   EXIT WHEN ( vl(i) /= vr(i) OR vl(i) = 'X' OR vr(i) = 'X');
		if( vl(i) /= vr(i) OR vl(i) = 'X' OR vr(i) = 'X')then
			if (vl(indx) = 'X' OR vr(indx) = 'X') Then
				ASSERT NOT WarningsOn
					REPORT "  --- Comparison is indeterminate will return " &
						" false in case of boolean and '0' in case of std_ulogic "
					SEVERITY WARNING;
			END IF;
			-- Compute the relationships based on the value of the differing bit
				return ( tbl_lt ( vl(indx), vr(indx) ) = '1');
		end if;
	 END LOOP;
--	if (vl(indx) = 'X' OR vr(indx) = 'X') Then
--	    ASSERT NOT WarningsOn
--	    REPORT "  --- Comparison is indeterminate will return " &
--		   " false in case of boolean and '0' in case of std_ulogic "
--	    SEVERITY WARNING;
--	 END IF;
     -- Compute the relationships based on the value of the differing bit
--	 return ( tbl_lt ( vl(indx), vr(indx) ) = '1');
		return FALSE;
	-- synopsys synthesis_on
     END LessThan_TwosComp;
 --+-----------------------------------------------------------------------------
 --|     Function Name : LessThan_Unsigned
 --|  hidden
 --|     Overloading    :
 --|
 --|     Purpose        : Compute the less than relation for BIT_VECTORS.
 --|
 --|     Parameters     :
 --|                      A          - input  BIT_VECTOR 
 --|                      B          - input  BIT_VECTOR 
 --|
 --|     NOTE           : The operands must be of same length with mode Unsigned.
 --|
 --|     Assumptions    : Both inputs must have range (msb downto 0)
 --|
 --|     Result         : Boolean
 --|
 --|     Use            : VARIABLE a, b : BIT_VECTOR ( 7 DOWNTO 0 );
 --|                      VARIABLE lt : boolean;
 --|                      lt := LessThan_Unsigned (l, r );
 --|-----------------------------------------------------------------------------
     FUNCTION LessThan_Unsigned       ( CONSTANT A          : IN  BIT_VECTOR;
			                CONSTANT B          : IN  BIT_VECTOR
			              ) return BOOLEAN IS
 	VARIABLE indx     : INTEGER;
	-- pragma map_to_operator LT_UNS_OP
	-- pragma type_function Return_Boolean_Unsigned         
	-- pragma return_port_name Z
     BEGIN
	-- synopsys synthesis_off
       -- perform comparison in a short circuit fashion
       -- Find the most significant differing bit : If equal use LSB
	 FOR i IN A'length - 1 DOWNTO 0 LOOP
	   indx := i;
--	   EXIT WHEN  A(i) /= B(i) ; 
		if (A(i) /= B(i)) then
			return( tbl_lt_bit ( A(indx), B(indx) ) = '1');
		end if;
	 END LOOP;

     -- Compute the relationships based on the value of the differing bit
--	 return( tbl_lt_bit ( A(indx), B(indx) ) = '1');
		return FALSE;
	-- synopsys synthesis_on
     END LessThan_Unsigned;
 --+-----------------------------------------------------------------------------
 --|     Function Name : LessThan_Unsigned
 --|  hidden
 --|     Overloading    :
 --|
 --|     Purpose        : Compute the less than relation for STD_LOGIC_VECTORS.
 --|
 --|     Parameters     :
 --|                      A          - input  STD_LOGIC_VECTOR 
 --|                      B          - input  STD_LOGIC_VECTOR 
 --|
 --|     NOTE           : The operands must be of same length with mode Unsigned.
 --|                      Any time the comparison reaches an index that has an 'X' as an
 --|                      array element, the comparison is deemed indeterminate and will 
 --|                      return boolean false.
 --|
 --|     Assumptions    : Both inputs must have range (msb downto 0)
 --|
 --|     Result         : Boolean
 --|
 --|     Use            : VARIABLE a, b : STD_LOGIC_VECTOR ( 7 DOWNTO 0 );
 --|                      VARIABLE lt : boolean;
 --|                      lt := LessThan_Unsigned (l, r );
 --|-----------------------------------------------------------------------------
     FUNCTION LessThan_Unsigned     ( CONSTANT A          : IN  STD_LOGIC_VECTOR;
			              CONSTANT B          : IN  STD_LOGIC_VECTOR
			            ) return BOOLEAN IS
 	VARIABLE indx     : INTEGER;
	-- pragma map_to_operator LT_UNS_OP
	-- pragma type_function Return_Boolean_Unsigned         
	-- pragma return_port_name Z
     BEGIN
	-- synopsys synthesis_off
       -- perform comparison in a short circuit fashion
       -- Find the most significant differing bit : If equal use LSB
	 FOR i IN A'length - 1 DOWNTO 0 LOOP
	   indx := i;
--	   EXIT WHEN ( A(i) /= B(i) OR A(i) = 'X' OR B(i) = 'X');
		if( A(i) /= B(i) OR A(i) = 'X' OR B(i) = 'X')then
			if (A(indx) = 'X' OR B(indx) = 'X') Then
				ASSERT NOT WarningsOn
					REPORT "   --- Comparison is indeterminate will return " &
						" false in case of boolean and '0' in case of std_ulogic "
					SEVERITY WARNING;
			END IF;
			-- Compute the relationships based on the value of the differing bit
			return( tbl_lt ( A(indx), B(indx) ) = '1');
		end if;
	 END LOOP;
--	if (A(indx) = 'X' OR B(indx) = 'X') Then
--	    ASSERT NOT WarningsOn
--	    REPORT "   --- Comparison is indeterminate will return " &
--		   " false in case of boolean and '0' in case of std_ulogic "
--	    SEVERITY WARNING;
--	 END IF;
     -- Compute the relationships based on the value of the differing bit
--	 return( tbl_lt ( A(indx), B(indx) ) = '1');
		return FALSE;
	-- synopsys synthesis_on
     END LessThan_Unsigned;
 --+-----------------------------------------------------------------------------
 --|     Function Name : LessThan_Unsigned
 --|  hidden
 --|     Overloading    :
 --|
 --|     Purpose        : Compute the less than relation for STD_ULOGIC_VECTORS.
 --|
 --|     Parameters     :
 --|                      A          - input  STD_ULOGIC_VECTOR 
 --|                      B          - input  STD_ULOGIC_VECTOR 
 --|
 --|     NOTE           : The operands must be of same length with mode Unsigned.
 --|
 --|                      Any time the comparison reaches an index that has an 'X' as an
 --|                      array element, the comparison is deemed indeterminate and will 
 --|                      return boolean false.
 --|
 --|     Assumptions    : Both inputs must have range (msb downto 0)
 --|
 --|     Result         : Boolean
 --|
 --|     Use            : VARIABLE a, b : STD_ULOGIC_VECTOR ( 7 DOWNTO 0 );
 --|                      VARIABLE lt : boolean;
 --|                      lt := LessThan_Unsigned (l, r );
 --|-----------------------------------------------------------------------------
     FUNCTION LessThan_Unsigned    ( CONSTANT A          : IN  STD_ULOGIC_VECTOR;
			             CONSTANT B          : IN  STD_ULOGIC_VECTOR
			           ) return BOOLEAN IS
 	VARIABLE indx     : INTEGER;
	-- pragma map_to_operator LT_UNS_OP
	-- pragma type_function Return_Boolean_Unsigned         
	-- pragma return_port_name Z
     BEGIN
       -- synopsys synthesis_off
       -- perform comparison in a short circuit fashion
       -- Find the most significant differing bit : If equal use LSB
	 FOR i IN A'length - 1 DOWNTO 0 LOOP
	   indx := i;
--	   EXIT WHEN ( A(i) /= B(i) OR A(i) = 'X' OR B(i) = 'X');
		if( A(i) /= B(i) OR A(i) = 'X' OR B(i) = 'X')then
			if (A(indx) = 'X' OR B(indx) = 'X') Then
				ASSERT NOT WarningsOn
					REPORT "  --- Comparison is indeterminate will return " &
						" false in case of boolean and '0' in case of std_ulogic "
					SEVERITY WARNING;
			END IF;
			-- Compute the relationships based on the value of the differing bit
			return( tbl_lt ( A(indx), B(indx) ) = '1');
		end if;
	 END LOOP;
--	if (A(indx) = 'X' OR B(indx) = 'X') Then
--	    ASSERT NOT WarningsOn
--	    REPORT "  --- Comparison is indeterminate will return " &
--		   " false in case of boolean and '0' in case of std_ulogic "
--	    SEVERITY WARNING;
--	 END IF;
     -- Compute the relationships based on the value of the differing bit
--	 return( tbl_lt ( A(indx), B(indx) ) = '1');
		return FALSE;
	-- synopsys synthesis_on
     END LessThan_Unsigned;
 --+-----------------------------------------------------------------------------
 --|     Function Name : LessThanOrEqual_TwosComp
 --|  hidden
 --|     Overloading    :
 --|
 --|     Purpose        : Compute the  less than or equal  relation 
 --|                      for BIT_VECTORS.
 --|
 --|     Parameters     :
 --|                      A          - input  BIT_VECTOR 
 --|                      B          - input  BIT_VECTOR 
 --|
 --|     NOTE           : The operands must be of same length with mode TwosComp.
 --|
 --|     Assumptions    : Both inputs must have range (msb downto 0)
 --|
 --|     Result         : Boolean
 --|
 --|     Use            : VARIABLE a, b : BIT_VECTOR ( 7 DOWNTO 0 );
 --|                      VARIABLE lte : boolean;
 --|                      lte := LessThanOrEqual_TwosComp (l, r );
 --|-----------------------------------------------------------------------------
     FUNCTION LessThanOrEqual_TwosComp   ( CONSTANT A      : IN  BIT_VECTOR;
			                   CONSTANT B      : IN  BIT_VECTOR
     			                 )  return BOOLEAN IS
       VARIABLE vl       : bit_vector (A'length - 1 downto 0);
       VARIABLE vr       : bit_vector (B'length - 1 downto 0);
       VARIABLE indx     : INTEGER;
       VARIABLE lt, eq   : Boolean;
	-- pragma map_to_operator LEQ_TC_OP
	-- pragma type_function Return_Boolean_TwosComp
	-- pragma return_port_name Z
     BEGIN
	-- synopsys synthesis_off
        vl := A;
        vr := B;
       -- complement the sign bit
	vl(A'length - 1) := NOT vl(B'length - 1);
	vr(B'length - 1) := NOT vr(B'length - 1);
       -- perform comparison in a short circuit fashion
       -- Find the most significant differing bit : If equal use LSB
	 FOR i IN A'length - 1 DOWNTO 0 LOOP
	   indx := i;
--	   EXIT WHEN  vl(i) /= vr(i) ; 
		if (vl(i) /= vr(i) )then 
			-- Compute the relationships based on the value of the differing bit
			lt := (tbl_lt_bit (vl(indx), vr(indx)) = '1');
			eq := (tbl_eq_bit (vl(indx), vr(indx)) = '1');
			return ( lt OR eq);
		end if;
	 END LOOP;
       -- Compute the relationships based on the value of the differing bit
--         lt := (tbl_lt_bit (vl(indx), vr(indx)) = '1');
--         eq := (tbl_eq_bit (vl(indx), vr(indx)) = '1');
--         return ( lt OR eq);
		return TRUE;
	-- synopsys synthesis_on
     END LessThanOrEqual_TwosComp;
 --+-----------------------------------------------------------------------------
 --|     Function Name : LessThanOrEqual_TwosComp
 --|  hidden
 --|     Overloading    :
 --|
 --|     Purpose        : Compute the  less than or equal  relation 
 --|                      for STD_LOGIC_VECTORS.
 --|
 --|     Parameters     :
 --|                      A          - input  STD_LOGIC_VECTOR 
 --|                      B          - input  STD_LOGIC_VECTOR 
 --|
 --|     NOTE           : The operands must be of same length with mode TwosComp.
 --|
 --|                      Any time the comparison reaches an index that has an 'X' as an
 --|                      array element, the comparison is deemed indeterminate and will 
 --|                      return boolean false.
 --|
 --|     Assumptions    : Both inputs must have range (msb downto 0)
 --|
 --|     Result         : Boolean
 --|
 --|     Use            : VARIABLE a, b : STD_LOGIC_VECTOR ( 7 DOWNTO 0 );
 --|                      VARIABLE lte : boolean;
 --|                      lte := LessThanOrEqual_TwosComp (l, r );
 --|-----------------------------------------------------------------------------
     FUNCTION LessThanOrEqual_TwosComp   ( CONSTANT A     : IN  STD_LOGIC_VECTOR;
			                   CONSTANT B     : IN  STD_LOGIC_VECTOR
     			                 ) return BOOLEAN IS
       VARIABLE vl       : std_logic_vector (A'length - 1 downto 0);
       VARIABLE vr       : std_logic_vector (B'length - 1 downto 0);
       VARIABLE indx     : INTEGER;
       VARIABLE lt, eq   : Boolean;
	-- pragma map_to_operator LEQ_TC_OP
	-- pragma type_function Return_Boolean_TwosComp
	-- pragma return_port_name Z
     BEGIN
	-- synopsys synthesis_off
        vl := A;
        vr := B;
       -- complement the sign bit
	vl(A'length - 1) := NOT vl(B'length - 1);
	vr(B'length - 1) := NOT vr(B'length - 1);
       -- perform comparison in a short circuit fashion
       -- Find the most significant differing bit : If equal use LSB
	 FOR i IN A'length - 1 DOWNTO 0 LOOP
	   indx := i;
--	   EXIT WHEN ( vl(i) /= vr(i) OR vl(i) = 'X' OR vr(i) = 'X');
		if ( vl(i) /= vr(i) OR vl(i) = 'X' OR vr(i) = 'X') then
			if (vl(indx) = 'X' OR vr(indx) = 'X') Then
				ASSERT NOT WarningsOn
					REPORT "  --- Comparison is indeterminate will return " &
						" false in case of boolean and '0' in case of std_ulogic "
					SEVERITY WARNING;
			END IF;
			-- Compute the relationships based on the value of the differing bit
			lt := (tbl_lt (vl(indx), vr(indx)) = '1');
			eq := (tbl_eq (vl(indx), vr(indx)) = '1');
			return ( lt OR eq);
		end if;
	 END LOOP;
--	if (vl(indx) = 'X' OR vr(indx) = 'X') Then
--	    ASSERT NOT WarningsOn
--	    REPORT "  --- Comparison is indeterminate will return " &
--		   " false in case of boolean and '0' in case of std_ulogic "
--	    SEVERITY WARNING;
--	 END IF;
       -- Compute the relationships based on the value of the differing bit
--         lt := (tbl_lt (vl(indx), vr(indx)) = '1');
--         eq := (tbl_eq (vl(indx), vr(indx)) = '1');
--         return ( lt OR eq);
		return TRUE;
	-- synopsys synthesis_on
     END LessThanOrEqual_TwosComp;
 --+-----------------------------------------------------------------------------
 --|     Function Name : LessThanOrEqual_TwosComp
 --|  hidden
 --|     Overloading    :
 --|
 --|     Purpose        : Compute the  less than or equal  relation 
 --|                      for STD_ULOGIC_VECTORS.
 --|
 --|     Parameters     :
 --|                      A          - input  STD_ULOGIC_VECTOR 
 --|                      B          - input  STD_ULOGIC_VECTOR 
 --|
 --|     NOTE           : The operands must be of same length with mode TwosComp.
 --|
 --|                      Any time the comparison reaches an index that has an 'X' as an
 --|                      array element, the comparison is deemed indeterminate and will 
 --|                      return boolean false.
 --|
 --|     Assumptions    : Both inputs must have range (msb downto 0)
 --|
 --|     Result         : Boolean
 --|
 --|     Use            : VARIABLE a, b : STD_ULOGIC_VECTOR ( 7 DOWNTO 0 );
 --|                      VARIABLE lte : boolean;
 --|                      lte := LessThanOrEqual_TwosComp (l, r );
 --|-----------------------------------------------------------------------------
     FUNCTION LessThanOrEqual_TwosComp   ( CONSTANT A    : IN  STD_ULOGIC_VECTOR;
			                   CONSTANT B    : IN  STD_ULOGIC_VECTOR
     			                 ) return BOOLEAN IS
       VARIABLE vl       : std_ulogic_vector (A'length - 1 downto 0);
       VARIABLE vr       : std_ulogic_vector (B'length - 1 downto 0);
       VARIABLE indx     : INTEGER;
       VARIABLE lt, eq   : Boolean;
	-- pragma map_to_operator LEQ_TC_OP
	-- pragma type_function Return_Boolean_TwosComp
	-- pragma return_port_name Z
     BEGIN
	-- synopsys synthesis_off
        vl := A;
        vr := B;
       -- complement the sign bit
	vl(A'length - 1) := NOT vl(B'length - 1);
	vr(B'length - 1) := NOT vr(B'length - 1);
       -- perform comparison in a short circuit fashion
       -- Find the most significant differing bit : If equal use LSB
	 FOR i IN A'length - 1 DOWNTO 0 LOOP
	   indx := i;
--	   EXIT WHEN ( vl(i) /= vr(i) OR vl(i) = 'X' OR vr(i) = 'X');
		if( vl(i) /= vr(i) OR vl(i) = 'X' OR vr(i) = 'X')then
			if (vl(indx) = 'X' OR vr(indx) = 'X') Then
				ASSERT NOT WarningsOn
					REPORT "   --- Comparison is indeterminate will return " &
						" false in case of boolean and '0' in case of std_ulogic "
					SEVERITY WARNING;
			END IF;
			-- Compute the relationships based on the value of the differing bit
			lt := (tbl_lt (vl(indx), vr(indx)) = '1');
			eq := (tbl_eq (vl(indx), vr(indx)) = '1');
			return ( lt OR eq);
		end if;
	 END LOOP;
--	if (vl(indx) = 'X' OR vr(indx) = 'X') Then
--	    ASSERT NOT WarningsOn
--	    REPORT "   --- Comparison is indeterminate will return " &
--		   " false in case of boolean and '0' in case of std_ulogic "
--	    SEVERITY WARNING;
--	 END IF;

       -- Compute the relationships based on the value of the differing bit
--         lt := (tbl_lt (vl(indx), vr(indx)) = '1');
--         eq := (tbl_eq (vl(indx), vr(indx)) = '1');
--         return ( lt OR eq);
		return TRUE;
	-- synopsys synthesis_on
     END LessThanOrEqual_TwosComp;
 --+-----------------------------------------------------------------------------
 --|     Function Name : LessThanOrEqual_Unsigned
 --|  hidden
 --|     Overloading    :
 --|
 --|     Purpose        : Compute the less than  or equal relation for BIT_VECTORS.
 --|
 --|     Parameters     :
 --|                      A          - input  BIT_VECTOR 
 --|                      B          - input  BIT_VECTOR 
 --|
 --|     NOTE           : The operands must be of same length with mode Unsigned.
 --|
 --|     Assumptions    : Both inputs must have range (msb downto 0)
 --|
 --|     Result         : Boolean
 --|
 --|     Use            : VARIABLE a, b : BIT_VECTOR ( 7 DOWNTO 0 );
 --|                      VARIABLE lt : boolean;
 --|                      lt := LessThanOrEqual_Unsigned (l, r );
 --|-----------------------------------------------------------------------------
     FUNCTION LessThanOrEqual_Unsigned   ( CONSTANT A          : IN  BIT_VECTOR;
			                    CONSTANT B          : IN  BIT_VECTOR
           		                 )  return BOOLEAN IS
        VARIABLE indx     : INTEGER;
 	VARIABLE lt, eq    : Boolean;	
	-- pragma map_to_operator LEQ_UNS_OP
	-- pragma type_function Return_Boolean_Unsigned
	-- pragma return_port_name Z
     BEGIN
	-- synopsys synthesis_off
       -- perform comparison in a short circuit fashion
       -- Find the most significant differing bit : If equal use LSB
	 FOR i IN A'length - 1 DOWNTO 0 LOOP
	   indx := i;
--	   EXIT WHEN  A(i) /= B(i) ; 
		if (A(i) /= B(i)) then
			-- Compute the relationships based on the value of the differing bit
			lt := (tbl_lt_bit (A(indx), B(indx)) = '1');
			eq := (tbl_eq_bit (A(indx), B(indx)) = '1');
			return ( lt OR eq);
		end if;
	 END LOOP;
     -- Compute the relationships based on the value of the differing bit
--         lt := (tbl_lt_bit (A(indx), B(indx)) = '1');
--         eq := (tbl_eq_bit (A(indx), B(indx)) = '1');
--         return ( lt OR eq);
		return TRUE;
	-- synopsys synthesis_on
     END LessThanOrEqual_Unsigned;
 --+-----------------------------------------------------------------------------
 --|     Function Name : LessThanOrEqual_Unsigned
 --|  hidden
 --|     Overloading    :
 --|
 --|     Purpose        : Compute the less than  or equal relation for STD_LOGIC_VECTORS.
 --|
 --|     Parameters     :
 --|                      A          - input  STD_LOGIC_VECTOR 
 --|                      B          - input  STD_LOGIC_VECTOR 
 --|
 --|     NOTE           : The operands must be of same length with mode Unsigned.
 --|
 --|                      Any time the comparison reaches an index that has an 'X' as an
 --|                      array element, the comparison is deemed indeterminate and will 
 --|                      return boolean false.
 --|
 --|     Assumptions    : Both inputs must have range (msb downto 0)
 --|
 --|     Result         : Boolean
 --|
 --|     Use            : VARIABLE a, b : STD_LOGIC_VECTOR ( 7 DOWNTO 0 );
 --|                      VARIABLE lt : boolean;
 --|                      lt := LessThanOrEqual_Unsigned (l, r );
 --|-----------------------------------------------------------------------------
     FUNCTION LessThanOrEqual_Unsigned   ( CONSTANT A    : IN  STD_LOGIC_VECTOR;
			                   CONSTANT B    : IN  STD_LOGIC_VECTOR
           		                 ) return BOOLEAN IS
        VARIABLE indx     : INTEGER;
 	VARIABLE lt, eq    : Boolean;	
	-- pragma map_to_operator LEQ_UNS_OP
	-- pragma type_function Return_Boolean_Unsigned
	-- pragma return_port_name Z
     BEGIN
	-- synopsys synthesis_off
       -- perform comparison in a short circuit fashion
       -- Find the most significant differing bit : If equal use LSB
	 FOR i IN A'length - 1 DOWNTO 0 LOOP
	   indx := i;
--	   EXIT WHEN ( A(i) /= B(i) OR A(i) = 'X' OR B(i) = 'X');
		if ( A(i) /= B(i) OR A(i) = 'X' OR B(i) = 'X') then
			if (A(indx) = 'X' OR B(indx) = 'X') Then
				ASSERT NOT WarningsOn
					REPORT "  --- Comparison is indeterminate will return " &
						" false in case of boolean and '0' in case of std_ulogic "
					SEVERITY WARNING;
			END IF;
			-- Compute the relationships based on the value of the differing bit
			lt := (tbl_lt (A(indx), B(indx)) = '1');
			eq := (tbl_eq (A(indx), B(indx)) = '1');
			return ( lt OR eq);
		end if;
	 END LOOP;
--	if (A(indx) = 'X' OR B(indx) = 'X') Then
--	    ASSERT NOT WarningsOn
--	    REPORT "  --- Comparison is indeterminate will return " &
--		   " false in case of boolean and '0' in case of std_ulogic "
--	    SEVERITY WARNING;
--	 END IF;
     -- Compute the relationships based on the value of the differing bit
--         lt := (tbl_lt (A(indx), B(indx)) = '1');
--         eq := (tbl_eq (A(indx), B(indx)) = '1');
--         return ( lt OR eq);
		return TRUE;
	-- synopsys synthesis_on
     END LessThanOrEqual_Unsigned;
 --+-----------------------------------------------------------------------------
 --|     Function Name : LessThanOrEqual_Unsigned
 --|  hidden
 --|     Overloading    :
 --|
 --|     Purpose        : Compute the less than  or equal relation for STD_ULOGIC_VECTORS.
 --|
 --|     Parameters     :
 --|                      A          - input  STD_ULOGIC_VECTOR 
 --|                      B          - input  STD_ULOGIC_VECTOR 
 --|
 --|     NOTE           : The operands must be of same length with mode Unsigned.
 --|
 --|                      Any time the comparison reaches an index that has an 'X' as an
 --|                      array element, the comparison is deemed indeterminate and will 
 --|                      return boolean false.
 --|
 --|     Assumptions    : Both inputs must have range (msb downto 0)
 --|
 --|     Result         : Boolean
 --|
 --|     Use            : VARIABLE a, b : STD_ULOGIC_VECTOR ( 7 DOWNTO 0 );
 --|                      VARIABLE lt : boolean;
 --|                      lt := LessThanOrEqual_Unsigned (l, r );
 --|-----------------------------------------------------------------------------
     FUNCTION LessThanOrEqual_Unsigned   ( CONSTANT A     : IN  STD_ULOGIC_VECTOR;
			                   CONSTANT B     : IN  STD_ULOGIC_VECTOR
           		                 )  return BOOLEAN IS
        VARIABLE indx     : INTEGER;
 	VARIABLE lt, eq    : Boolean;	
	-- pragma map_to_operator LEQ_UNS_OP
	-- pragma type_function Return_Boolean_Unsigned
	-- pragma return_port_name Z
     BEGIN
	-- synopsys synthesis_off
       -- perform comparison in a short circuit fashion
       -- Find the most significant differing bit : If equal use LSB
	 FOR i IN A'length - 1 DOWNTO 0 LOOP
	   indx := i;
--	   EXIT WHEN ( A(i) /= B(i) OR A(i) = 'X' OR B(i) = 'X');
		if( A(i) /= B(i) OR A(i) = 'X' OR B(i) = 'X')then
			if (A(indx) = 'X' OR B(indx) = 'X') Then
				ASSERT NOT WarningsOn
					REPORT "  --- Comparison is indeterminate will return " &
						" false in case of boolean and '0' in case of std_ulogic "
					SEVERITY WARNING;
			END IF;
			-- Compute the relationships based on the value of the differing bit
			lt := (tbl_lt (A(indx), B(indx)) = '1');
			eq := (tbl_eq (A(indx), B(indx)) = '1');
			return ( lt OR eq);
		end if;
	 END LOOP;
--	if (A(indx) = 'X' OR B(indx) = 'X') Then
--	    ASSERT NOT WarningsOn
--	    REPORT "  --- Comparison is indeterminate will return " &
--		   " false in case of boolean and '0' in case of std_ulogic "
--	    SEVERITY WARNING;
--	 END IF;
     -- Compute the relationships based on the value of the differing bit
--         lt := (tbl_lt (A(indx), B(indx)) = '1');
--         eq := (tbl_eq (A(indx), B(indx)) = '1');
--         return ( lt OR eq);
		return TRUE;
	-- synopsys synthesis_on
     END LessThanOrEqual_Unsigned;
 --+-----------------------------------------------------------------------------
 --|     Function Name : Equal
 --|  hidden
 --|     Overloading    :
 --|
 --|     Purpose        : Compute the relation Equal for BIT_VECTORS.
 --|
 --|     Parameters     : L          - input  BIT_VECTOR 
 --|                      R          - input  BIT_VECTOR 
 --|
 --|     NOTE           : The operands must be of same length with mode TwosComp.
 --|
 --|     Assumptions    : Both inputs must have range (msb downto 0)
 --|
 --|     Result         : Boolean
 --|
 --|     Use            : VARIABLE a, b : BIT_VECTOR ( 7 DOWNTO 0 );
 --|                      VARIABLE eq : boolean;
 --|                      eq := Equal (l, r );
 --|-----------------------------------------------------------------------------
     FUNCTION Equal   ( CONSTANT L          : IN  BIT_VECTOR;
	       		CONSTANT R          : IN  BIT_VECTOR
 		     )  return BOOLEAN IS
       VARIABLE indx     : INTEGER;
	-- pragma built_in  SYN_EQL
     BEGIN
	-- synopsys synthesis_off
       -- perform comparison in a short circuit fashion
       -- Find the most significant differing bit : If equal use LSB
	 FOR i IN L'length - 1 DOWNTO 0 LOOP
	   indx := i;
--	   EXIT WHEN  L(i) /= R(i) ; 
		if (L(i) /= R(i)) then
			-- Compute the relationships based on the value of the differing bit
			return( tbl_eq_bit (L(indx), R(indx) ) = '1');
		end if;
	 END LOOP;
     -- Compute the relationships based on the value of the differing bit
--	 return( tbl_eq_bit (L(indx), R(indx) ) = '1');
		return TRUE;
	-- synopsys synthesis_on
     END Equal;
 --+-----------------------------------------------------------------------------
 --|     Function Name : Equal
 --|  hidden
 --|     Overloading    :
 --|
 --|     Purpose        : Compute the relation Equal for STD_LOGIC_VECTORS.
 --|
 --|     Parameters     : L          - input  STD_LOGIC_VECTOR 
 --|                      R          - input  STD_LOGIC_VECTOR 
 --|
 --|     NOTE           : The operands must be of same length with mode TwosComp.
 --|
 --|                      Any time the comparison reaches an index that has an 'X' as an
 --|                      array element, the comparison is deemed indeterminate and will 
 --|                      return boolean false.
 --|
 --|     Assumptions    : Both inputs must have range (msb downto 0)
 --|
 --|     Result         : Boolean
 --|
 --|     Use            : VARIABLE a, b : STD_LOGIC_VECTOR ( 7 DOWNTO 0 );
 --|                      VARIABLE eq : boolean;
 --|                      eq := Equal (l, r );
 --|-----------------------------------------------------------------------------
     FUNCTION Equal   ( CONSTANT L          : IN  STD_LOGIC_VECTOR;
	       		CONSTANT R          : IN  STD_LOGIC_VECTOR
 		     )  return BOOLEAN IS
       VARIABLE indx     : INTEGER;
	-- pragma built_in  SYN_EQL
     BEGIN
	-- synopsys synthesis_off
       -- perform comparison in a short circuit fashion
       -- Find the most significant differing bit : If equal use LSB
	 FOR i IN L'length - 1 DOWNTO 0 LOOP
	   indx := i;
--	   EXIT WHEN ( L(i) /= R(i) OR L(i) = 'X' OR R(i) = 'X');
		if( L(i) /= R(i) OR L(i) = 'X' OR R(i) = 'X')then
			if (L(indx) = 'X' OR R(indx) = 'X') Then
				ASSERT NOT WarningsOn
					REPORT " Equal  --- Comparison is indeterminate will return " &
						" false in case of boolean and '0' in case of std_ulogic "
				SEVERITY WARNING;
			END IF;
			-- Compute the relationships based on the value of the differing bit
			return( tbl_eq (L(indx), R(indx) ) = '1');
		end if;
	 END LOOP;
--	if (L(indx) = 'X' OR R(indx) = 'X') Then
--	    ASSERT NOT WarningsOn
--	    REPORT " Equal  --- Comparison is indeterminate will return " &
--		   " false in case of boolean and '0' in case of std_ulogic "
--	    SEVERITY WARNING;
--	 END IF;
     -- Compute the relationships based on the value of the differing bit
--	 return( tbl_eq (L(indx), R(indx) ) = '1');
		return TRUE;
	-- synopsys synthesis_on
     END Equal;
 --+-----------------------------------------------------------------------------
 --|     Function Name : Equal
 --|  hidden
 --|     Overloading    :
 --|
 --|     Purpose        : Compute the relation Equal for STD_ULOGIC_VECTORS.
 --|
 --|     Parameters     : L          - input  STD_ULOGIC_VECTOR 
 --|                      R          - input  STD_ULOGIC_VECTOR 
 --|
 --|     NOTE           : The operands must be of same length with mode TwosComp.
 --|
 --|                      Any time the comparison reaches an index that has an 'X' as an
 --|                      array element, the comparison is deemed indeterminate and will 
 --|                      return boolean false.
 --|
 --|     Assumptions    : Both inputs must have range (msb downto 0)
 --|
 --|     Result         : Boolean
 --|
 --|     Use            : VARIABLE a, b : STD_ULOGIC_VECTOR ( 7 DOWNTO 0 );
 --|                      VARIABLE eq : boolean;
 --|                      eq := Equal (l, r );
 --|-----------------------------------------------------------------------------
     FUNCTION Equal   ( CONSTANT L          : IN  STD_ULOGIC_VECTOR;
	       		CONSTANT R          : IN  STD_ULOGIC_VECTOR
 		     )  return BOOLEAN IS
       VARIABLE indx     : INTEGER;
	-- pragma built_in  SYN_EQL
     BEGIN
	-- synopsys synthesis_off
       -- perform comparison in a short circuit fashion
       -- Find the most significant differing bit : If equal use LSB
	 FOR i IN L'length - 1 DOWNTO 0 LOOP
	   indx := i;
--	   EXIT WHEN ( L(i) /= R(i) OR L(i) = 'X' OR R(i) = 'X');
		if( L(i) /= R(i) OR L(i) = 'X' OR R(i) = 'X')then
			if (L(indx) = 'X' OR R(indx) = 'X') Then
				ASSERT NOT WarningsOn
					REPORT " Equal  --- Comparison is indeterminate will return " &
						" false in case of boolean and '0' in case of std_ulogic "
					SEVERITY WARNING;
			END IF;
			-- Compute the relationships based on the value of the differing bit
			return( tbl_eq (L(indx), R(indx) ) = '1');
		end if;
	 END LOOP;
--	if (L(indx) = 'X' OR R(indx) = 'X') Then
--	    ASSERT NOT WarningsOn
--	    REPORT " Equal  --- Comparison is indeterminate will return " &
--		   " false in case of boolean and '0' in case of std_ulogic "
--	    SEVERITY WARNING;
--	 END IF;
     -- Compute the relationships based on the value of the differing bit
--	 return( tbl_eq (L(indx), R(indx) ) = '1');
		return TRUE;
	-- synopsys synthesis_on
     END Equal;
 --+-----------------------------------------------------------------------------
 --|     Function Name : NotEqual
 --|  hidden
 --|     Overloading    :
 --|
 --|     Purpose        : Compute the not Equal relation for BIT_VECTORS.
 --|
 --|     Parameters     : L          - input  BIT_VECTOR 
 --|                      R          - input  BIT_VECTOR 
 --|
 --|     NOTE           : The operands must be of same length with mode Unsigned.
 --|
 --|     Assumptions    : Both inputs must have range (msb downto 0)
 --|
 --|     Result         : Boolean
 --|
 --|     Use            : VARIABLE a, b : BIT_VECTOR ( 7 DOWNTO 0 );
 --|                      VARIABLE neq : boolean;
 --|                      neq := NotEqual (l, r );
 --|-----------------------------------------------------------------------------
     FUNCTION NotEqual          ( CONSTANT L          : IN  BIT_VECTOR;
			          CONSTANT R          : IN  BIT_VECTOR
			        )  return BOOLEAN IS
       VARIABLE indx     : INTEGER;
	-- pragma built_in  SYN_NEQ
     BEGIN
	-- synopsys synthesis_off
       -- perform comparison in a short circuit fashion
       -- Find the most significant differing bit : If equal use LSB
	 FOR i IN L'length - 1 DOWNTO 0 LOOP
	   indx := i;
--	   EXIT WHEN  L(i) /= R(i) ; 
		if (L(i) /= R(i)) then
			-- Compute the relationships based on the value of the differing bit
			return ( NOT ( tbl_eq_bit ( L(indx), R(indx) ) = '1'));
		end if;
	 END LOOP;
     -- Compute the relationships based on the value of the differing bit
--	 return ( NOT ( tbl_eq_bit ( L(indx), R(indx) ) = '1'));
		return FALSE;
	-- synopsys synthesis_on
     END NotEqual;
 --+-----------------------------------------------------------------------------
 --|     Function Name : NotEqual
 --|  hidden
 --|     Overloading    :
 --|
 --|     Purpose        : Compute the not Equal relation for STD_LOGIC_VECTORS.
 --|
 --|     Parameters     : L          - input  STD_LOGIC_VECTOR 
 --|                      R          - input  STD_LOGIC_VECTOR 
 --|
 --|     NOTE           : The operands must be of same length with mode Unsigned.
 --|
 --|                      Any time the comparison reaches an index that has an 'X' as an
 --|                      array element, the comparison is deemed indeterminate and will 
 --|                      return boolean false.
 --|
 --|     Assumptions    : Both inputs must have range (msb downto 0)
 --|
 --|     Result         : Boolean
 --|
 --|     Use            : VARIABLE a, b : STD_LOGIC_VECTOR ( 7 DOWNTO 0 );
 --|                      VARIABLE neq : boolean;
 --|                      neq := NotEqual (l, r );
 --|-----------------------------------------------------------------------------
     FUNCTION NotEqual          ( CONSTANT L          : IN  STD_LOGIC_VECTOR;
			          CONSTANT R          : IN  STD_LOGIC_VECTOR
			        )  return BOOLEAN IS
       VARIABLE indx     : INTEGER;
	-- pragma built_in  SYN_NEQ
     BEGIN
	-- synopsys synthesis_off
       -- perform comparison in a short circuit fashion
       -- Find the most significant differing bit : If equal use LSB
	 FOR i IN L'length - 1 DOWNTO 0 LOOP
	   indx := i;
--	   EXIT WHEN ( L(i) /= R(i) OR L(i) = 'X' OR R(i) = 'X');
		if( L(i) /= R(i) OR L(i) = 'X' OR R(i) = 'X')then
			if (L(indx) = 'X' OR R(indx) = 'X') Then
				ASSERT NOT WarningsOn
					REPORT " NotEqual  --- Comparison is indeterminate will return " &
						" false in case of boolean and '0' in case of std_ulogic "
					SEVERITY WARNING;
				return false;
			else
				-- Compute the relationships based on the value of the differing bit
				return ( NOT ( tbl_eq ( L(indx), R(indx) ) = '1'));
			end if;
		end if;
	 END LOOP;
--	if (L(indx) = 'X' OR R(indx) = 'X') Then
--	      ASSERT NOT WarningsOn
--	      REPORT " NotEqual  --- Comparison is indeterminate will return " &
--		   " false in case of boolean and '0' in case of std_ulogic "
--	      SEVERITY WARNING;
--              return false;
--         else
        -- Compute the relationships based on the value of the differing bit
--	      return ( NOT ( tbl_eq ( L(indx), R(indx) ) = '1'));
--         end if;
		return FALSE;
	-- synopsys synthesis_on
     END NotEqual;
 --+-----------------------------------------------------------------------------
 --|     Function Name : NotEqual
 --|  hidden
 --|     Overloading    :
 --|
 --|     Purpose        : Compute the not Equal relation for STD_ULOGIC_VECTORS.
 --|
 --|     Parameters     : L          - input  STD_ULOGIC_VECTOR 
 --|                      R          - input  STD_ULOGIC_VECTOR 
 --|
 --|     NOTE           : The operands must be of same length with mode Unsigned.
 --|
 --|                      Any time the comparison reaches an index that has an 'X' as an
 --|                      array element, the comparison is deemed indeterminate and will 
 --|                      return boolean false.
 --|
 --|     Assumptions    : Both inputs must have range (msb downto 0)
 --|
 --|     Result         : Boolean
 --|
 --|     Use            : VARIABLE a, b : STD_ULOGIC_VECTOR ( 7 DOWNTO 0 );
 --|                      VARIABLE neq : boolean;
 --|                      neq := NotEqual (l, r );
 --|-----------------------------------------------------------------------------
     FUNCTION NotEqual          ( CONSTANT L          : IN  STD_ULOGIC_VECTOR;
			          CONSTANT R          : IN  STD_ULOGIC_VECTOR
			        )  return BOOLEAN IS
       VARIABLE indx     : INTEGER;
	-- pragma built_in  SYN_NEQ
     BEGIN
	-- synopsys synthesis_off
       -- perform comparison in a short circuit fashion
       -- Find the most significant differing bit : If equal use LSB
	 FOR i IN L'length - 1 DOWNTO 0 LOOP
	   indx := i;
--	   EXIT WHEN ( L(i) /= R(i) OR L(i) = 'X' OR R(i) = 'X');
		if( L(i) /= R(i) OR L(i) = 'X' OR R(i) = 'X')then
			if (L(indx) = 'X' OR R(indx) = 'X') Then
				ASSERT NOT WarningsOn
					REPORT " NotEqual  --- Comparison is indeterminate will return " &
						" false in case of boolean and '0' in case of std_ulogic "
					SEVERITY WARNING;
				return false;
			else
				-- Compute the relationships based on the value of the differing bit
				return ( NOT ( tbl_eq ( L(indx), R(indx) ) = '1'));
			end if;
		end if;
	 END LOOP;
--	if (L(indx) = 'X' OR R(indx) = 'X') Then
--  	      ASSERT NOT WarningsOn
--	      REPORT " NotEqual  --- Comparison is indeterminate will return " &
--		   " false in case of boolean and '0' in case of std_ulogic "
--	      SEVERITY WARNING;
--              return false;
--        else
        -- Compute the relationships based on the value of the differing bit
--	      return ( NOT ( tbl_eq ( L(indx), R(indx) ) = '1'));
--        end if;
		return FALSE;	
	-- synopsys synthesis_on
     END NotEqual;
    -------------------------------------------------------------------------------
    --     Function Name  : RegFill_Zero
    -- 1.7.3
    --     Overloading    : None
    --
    --     Purpose        : Fill the most significant bits of a register with a '0'
    --
    --     Parameters     :
    --                      ARG     - input  std_logic_vector, the vector to be read.
    --                      SIZE  - input  INTEGER, length of the return vector.
    --
    --     Result         : std_logic_vector
    --
    --     NOTE           : The length of the return bit vector  is specified by the
    --                      parameter 'SIZE'. The input logic vector will
    --                      be  filled with the '0'.
    --     Use            :
    --                      VARIABLE vect : std_logic_vector ( 15 DOWNTO 0 );
    --                      vect := RegFill_Zero ( "00000101", 16);
    -------------------------------------------------------------------------------
    FUNCTION RegFill_Zero   ( CONSTANT ARG    : IN std_logic_vector;
                              CONSTANT SIZE   : IN INTEGER
                            ) RETURN std_logic_vector IS
      VARIABLE result : std_logic_vector (SIZE - 1 DOWNTO 0);
      VARIABLE  reg   : std_logic_vector (ARG'LENGTH - 1 DOWNTO 0);
      -- synopsys built_in SYN_ZERO_EXTEND
    BEGIN
      -- synopsys synthesis_off
      --  null range check
      reg := ARG;
      IF (ARG'LENGTH = 0) THEN
         IF (SIZE = 0) THEN
            ASSERT FALSE
            REPORT " RegFill_Zero --- input  has null range and" &
                " Destination also has null range. "
            SEVERITY ERROR;
            RETURN result ;
         ELSE
            ASSERT FALSE
            REPORT " RegFill_Zero --- input  has null range"
            SEVERITY ERROR;
            result := (OTHERS => '0');
            RETURN result ;
         END IF;
 
      ELSIF (SIZE = 0) THEN
          ASSERT false
          REPORT "RegFill_Zero --- Destination has null range "
          SEVERITY ERROR;
          RETURN result;
 
      ELSIF (SIZE <= ARG'LENGTH) THEN
                        -- no need to sign extend
         ASSERT (SIZE = ARG'LENGTH)
         REPORT " RegFill_Zero ---  Destination length is less than source"
         SEVERITY ERROR;
         RETURN reg;        -- return the input data without any change

       ELSE
           result(ARG'LENGTH - 1 DOWNTO 0) := reg;
        -- Fill the MSB's of result with the given fill value.
          For i IN SIZE - 1 DOWNTO ARG'LENGTH  Loop
             result(i) := '0';
          END LOOP;
       END IF;
       RETURN  To_X01(result);
      -- synopsys synthesis_on
    END RegFill_Zero;
    -------------------------------------------------------------------------------
    --     Function Name  : SignExtend_TwosComp
    -- 1.7.2
    --     Overloading    : None
    --
    --     Purpose        : Sign Extend an std_logic_vector
    --
    --     Parameters     :
    --                      ARG     - input  std_logic_vector, the vector to be read.
    --                      SIZE  - input  INTEGER, length of the return vector.
    --
    --     Result         : std_logic_vector, the extened std_logic_vector
    --
    --     NOTE           : The length of the return logic vector  is specified by the
    --                      parameter 'SIZE'. The input logic vector will 
    --                      be sign extended. 
    --                
    --                      Sign-position is the Most Significant Bit (MSB)
     --     Use            :
    --                      VARIABLE vect : std_logic_vector ( 15 DOWNTO 0 );
    --                      vect := SignExtend_TwosComp ( "11111101", 16); -- set to -4
     -------------------------------------------------------------------------------
    FUNCTION SignExtend_TwosComp   ( CONSTANT ARG    : IN std_logic_vector;
                                     CONSTANT SIZE   : IN INTEGER
                                   ) RETURN std_logic_vector IS
      VARIABLE result   : std_logic_vector (SIZE - 1 DOWNTO 0); 
      VARIABLE reg      : std_logic_vector (ARG'LENGTH - 1 DOWNTO 0);
      VARIABLE sign     : std_ulogic;
      VARIABLE sign_pos : INTEGER;
      -- synopsys built_in SYN_SIGN_EXTEND
    --
    BEGIN
    -- synopsys synthesis_off
       result     := (OTHERS => '0');
       reg        := ARG;
       -- Internally ARG is copied  to reg which  is defined ARG'LENGTH - 1 downto 0
       -- There sign bit position is now ARG'LENGTH - 1. This will take care of ascending
       -- as well as descending range input ARG.
      sign_pos := ARG'LENGTH - 1;
     --  null range check
      IF (ARG'LENGTH = 0) THEN
         IF (SIZE = 0) THEN
            ASSERT FALSE
            REPORT " SignExtend_TwosComp --- input register has null range" &
                " Destination has also null range "
            SEVERITY ERROR;
            RETURN result ;
         ELSE 
            ASSERT FALSE
            REPORT " SignExtend_TwosComp --- input register has null range" 
            SEVERITY ERROR;
            RETURN result ;
         END IF;

      ELSIF (SIZE = 0) THEN
          ASSERT false
          REPORT "SignExtend_TwosComp --- Destination length of zero was passed "
          SEVERITY ERROR;
          RETURN result;

      ELSIF (SIZE <= ARG'LENGTH) THEN
                        -- no need to sign extend
         ASSERT (SIZE = ARG'LENGTH)
         REPORT " SignExtend_TwosComp ---  Destination length is not greater than source"
         SEVERITY ERROR;
         RETURN reg;        -- return the input data without any change
 
      ELSE
          --  save the sign bit
          sign := reg(sign_pos);
         -- Copy the source register to variable result up to the sign position - 1.
            For i IN sign_pos - 1 DOWNTO 0 LOOP
               result(i) := reg(i);
            END LOOP;
      
         -- Extend the sign depending on the regmode. TwosComp
            For i IN SIZE - 1 DOWNTO sign_pos Loop
                   result(i) := sign;
            END LOOP;
      END IF;
      RETURN ( To_X01(result));
    -- synopsys synthesis_on	
    END SignExtend_TwosComp;
--+-----------------------------------------------------------------------------
--|     Function Name  : Add_TwosComp
--|  hidden function
--|     Overloading    : None
--|
--|     Purpose        : Two's Complement Addition of STD_LOGIC_VECTORS.
--|
--|     Parameters     :
--|                      A     - input  STD_LOGIC_VECTOR,
--|                      B     - input  STD_LOGIC_VECTOR,
--|     NOTE           : 
--|                      This function is implemented based on hardware design of a
--|                      Two's complement adder.
--|                      The inputs may be of any length  but both A and B
--|                      must have same lengths.
--|                    
--|                    
--|     Assumptions    : Both inputs must have range (msb downto 0)
--|
--|     Result         : returns bit_vector of the same length as A and B.
--|
--|     Use            : VARIABLE x, y, sum : STD_LOGIC_VECTOR ( 15 DOWNTO 0);
--|                      sum:=Add_TwosComp (x, y);
--|-----------------------------------------------------------------------------
     FUNCTION  Add_TwosComp  ( CONSTANT A     :  IN Std_Logic_Vector;
                               CONSTANT B     :  IN Std_Logic_Vector
                             )  RETURN Std_Logic_Vector IS 
      VARIABLE r        : Std_Logic_Vector ( A'LENGTH - 1  DOWNTO 0 );
      VARIABLE p        : STD_ULOGIC;
      VARIABLE g        : STD_ULOGIC;
      VARIABLE carry    : STD_ULOGIC;
      -- pragma map_to_operator ADD_TC_OP
      -- pragma return_port_name Z      
    BEGIN
	-- initialization
	p     := '1';
	g     := '0';
	carry := '0';  -- for twoscomp add set carry in '0'
	-- perform addition
      FOR n IN 0 TO A'LENGTH - 1 LOOP
             p := p AND (A(n) OR B(n));                        -- Cpropagate
             g := (A(n) AND B(n)) OR ( g AND (A(n) OR B(n)));  -- Cgenerate
          r(n) :=  A(n) XOR B(n) XOR carry;                    -- individual bit sums
         carry :=  g OR (p AND carry);                         -- carry
      END LOOP;
      RETURN r;
    END Add_TwosComp;
--+-----------------------------------------------------------------------------
--|     Function Name  : Add_Unsigned
--|  hidden procedure 
--|     Overloading    : None
--|
--|     Purpose        : Addition of unsigned STD_LOGIC_VECTORS.
--|
--|     Parameters     :
--|                      A     - input  STD_LOGIC_VECTOR,
--|                      B     - input  STD_LOGIC_VECTOR,
--|     NOTE           : 
--|                      This function is implemented based on hardware design of a
--|                      Two's complement adder.
--|                      The inputs may be of any length  but both A and B
--|                      must have same lengths.
--|                    
--|     Assumptions    : Both inputs must have range (msb downto 0)
--|
--|     Result         : returns bit_vector of the same length as A and B.
--|
--|     Use            : VARIABLE x, y, sum : STD_LOGIC_VECTOR ( 15 DOWNTO 0);
--|                      sum:=Add_Unsigned (x, y);
--|-----------------------------------------------------------------------------
     FUNCTION  Add_Unsigned  ( CONSTANT A     :  IN Std_Logic_Vector;
                               CONSTANT B     :  IN Std_Logic_Vector
                             )  RETURN Std_Logic_Vector IS 
      VARIABLE r        : Std_Logic_Vector ( A'LENGTH - 1  DOWNTO 0 );
      VARIABLE p        : STD_ULOGIC;
      VARIABLE g        : STD_ULOGIC;
      VARIABLE carry    : STD_ULOGIC;
      -- pragma map_to_operator ADD_UNS_OP
      -- pragma return_port_name Z      
    BEGIN
	-- initialization
	p     := '1';
	g     := '0';
	carry := '0';  -- for Unsigned add set carry in '0'
	-- perform addition
      FOR n IN 0 TO A'LENGTH - 1 LOOP
             p := p AND (A(n) OR B(n));                        -- Cpropagate
             g := (A(n) AND B(n)) OR ( g AND (A(n) OR B(n)));  -- Cgenerate
          r(n) :=  A(n) XOR B(n) XOR carry;                    -- individual bit sums
         carry :=  g OR (p AND carry);                         -- carry
      END LOOP;
      RETURN r;
    END Add_Unsigned;
--+-----------------------------------------------------------------------------
--|     Function Name  : Add_TwosComp_VHDL_TECH
--|  hidden procedure
--|     Overloading    : None
--|
--|     Purpose        : Two's Complement Addition of LOGIC VECTORS.
--|
--|     Parameters     :
--|                      result     - output std_logic_vector, the computed sum
--|                      carry_out  - output std_logic, 
--|                      overflow   - output std_logic, overflow condition
--|                      addend     - input  std_logic_vector,
--|                      augend     - input  std_logic,
--|                      carry_in   - input std_logic,
--|     NOTE           :
--|                      This procedure is implemented based on hardware design of a
--|                      Two's complement adder. 
--|                      The inputs may be of any length  but both addend and augend
--|                      must have same lengths.
--|
--|     Use            : VARIABLE x, y, sum : std_logic_vector ( 15 DOWNTO 0);
--|                      VARIABLE carry, ovf : std_ulogic;
--|
--|                      Add_TwosComp_VHDL_TECH ( sum, carry, ovf, x, y, '0' );
--|-----------------------------------------------------------------------------
    PROCEDURE Add_TwosComp_VHDL_TECH  ( VARIABLE result     : OUT std_logic_vector;
                              VARIABLE carry_out  : OUT std_ulogic;
                              VARIABLE overflow   : OUT std_ulogic;
                              CONSTANT addend     :  IN std_logic_vector;
                              CONSTANT augend     :  IN std_logic_vector;
                              CONSTANT carry_in   :  IN std_ulogic
                             ) IS
      CONSTANT reglen   : INTEGER := addend'LENGTH;
      VARIABLE a        : std_logic_vector ( reglen - 1  DOWNTO 0 );
      VARIABLE b        : std_logic_vector ( augend'LENGTH - 1  DOWNTO 0 );
      VARIABLE r        : std_logic_vector ( reglen - 1  DOWNTO 0 );
      VARIABLE p        : std_ulogic;
      VARIABLE g        : std_ulogic;
      VARIABLE c_iminus : std_ulogic;
      VARIABLE carry    : std_ulogic;
    BEGIN
	-- initialization
        a     := addend;
        b     := augend;
	p     := '1';
	g     := '0';
	carry := carry_in;
	-- perform addition
    -- check the length of addend and augend
    -- synopsys translate_off
      ASSERT   (addend'LENGTH = augend'LENGTH)
      REPORT " Add_TwosComp_VHDL_TECH --- operand lenght not same "
      SEVERITY ERROR;
    -- synopsys translate_on
    -- perform the add using a simple ripple carry bit wise add.
      FOR n IN 0 TO reglen - 1 LOOP
           c_iminus := carry;
             p := p AND (a(n) OR b(n));                        -- Cpropagate
             g := (a(n) AND b(n)) OR ( g AND (a(n) OR b(n)));  -- Cgenerate
          r(n) :=  a(n) XOR b(n) XOR carry;                    -- individual bit sums
         carry :=  g OR (p AND carry);                         -- carry
      END LOOP;
      carry_out := To_X01(carry);
    -- set overflow if carry_in and carry_out of sign bit are different.
         overflow := To_X01(c_iminus XOR carry);
         result   := To_X01( r);
        RETURN;
    END Add_TwosComp_VHDL_TECH;
--+-----------------------------------------------------------------------------
--|     Function Name  : Add_Unsigned_VHDL_TECH
--|  hidden procedure
--|     Overloading    : None
--|
--|     Purpose        : Addition of LOGIC VECTORS in unsigned mode.
--|
--|     Parameters     :
--|                      result     - output std_logic_vector, the computed sum
--|                      carry_out  - output std_ulogic,
--|                      overflow   - output std_logic, overflow condition
--|                      addend     - input  std_logic_vector,
--|                      augend     - input  std_logic_vector,
--|                      carry_in   - input std_ulogic,
--|     NOTE           :
--|                      The inputs may be of any length  but both addend and augend
--|                      must have same lengths.
--|
--|     Use            : VARIABLE x, y, sum : std_logic_vector ( 15 DOWNTO 0);
--|                      VARIABLE carry, ovf : std_ulogic;
--|
--|                      Add_Unsigned ( sum, carry, ovf, x, y, '0' );
--|-----------------------------------------------------------------------------
    PROCEDURE Add_Unsigned_VHDL_TECH  ( VARIABLE result     : OUT std_logic_vector;
                              VARIABLE carry_out  : OUT std_ulogic;
                              VARIABLE overflow   : OUT std_ulogic;
                              CONSTANT addend     :  IN std_logic_vector;
                              CONSTANT augend     :  IN std_logic_vector;
                              CONSTANT carry_in   :  IN std_ulogic
                -- synopsys synthesis_off
                                                       := '0'
                 -- synopsys synthesis_on
                             ) IS
 
      CONSTANT reglen : INTEGER := addend'LENGTH;
      VARIABLE a      : std_logic_vector ( reglen - 1  DOWNTO 0 );
      VARIABLE b      : std_logic_vector ( augend'LENGTH - 1  DOWNTO 0 );
      VARIABLE r      : std_logic_vector ( reglen - 1  DOWNTO 0 );
      VARIABLE p      : std_ulogic;
      VARIABLE g      : std_ulogic;
      VARIABLE carry  : std_ulogic;
    BEGIN
	-- initialization
        a     := addend;
        b     := augend;
	p     := '1';
	g     := '0';
	carry := carry_in;
	-- perform addition
    -- check the length of addend and augend
    -- synopsys translate_off
      ASSERT   (addend'LENGTH = augend'LENGTH)
      REPORT " Add_Unsigned --- operand lenght not same "
      SEVERITY ERROR;
     -- synopsys translate_on
    -- perform the add using a simple ripple carry bit wise add.
      FOR n IN 0 TO reglen - 1 LOOP
             p := p AND (a(n) OR b(n));                        -- Cpropagate
             g := (a(n) AND b(n)) OR ( g AND (a(n) OR b(n)));  -- Cgenerate
          r(n) :=  a(n) XOR b(n) XOR carry;                    -- individual bit sums
         carry :=  g OR (p AND carry);                         -- carry
      END LOOP;
      carry_out := To_X01(carry);
    -- set overflow if carry_in and carry_out of last bit postition are different.
         overflow := To_X01(carry);
         result := To_X01(r);
        RETURN;
    END Add_Unsigned_VHDL_TECH;
--+-----------------------------------------------------------------------------
--|     Function Name  : Sub_TwosComp
--|  hidden procedure
--|     Overloading    : None
--|
--|     Purpose        : Two's Complement subtraction of STD_LOGIC_VECTORS.
--|
--|     Parameters     :
--|                      A     - input  STD_LOGIC_VECTOR,
--|                      B     - input  STD_LOGIC_VECTOR,
--|     NOTE           : 
--|                      This function is implemented based on hardware design of a
--|                      Two's complement adder/subtractor
--|
--|                      The inputs may be of any length  but both A and B
--|                      must have same lengths.
--|                      
--|     Assumptions    : Both inputs must have range (msb downto 0)
--|
--|     Result         : returns STD_LOGIC_vector of the same length as A and B.
--|
--|     Use            : VARIABLE x, y, sum : STD_LOGIC_VECTOR ( 15 DOWNTO 0);
--|                       sum:= Sub_TwosComp (x, y);
--|-----------------------------------------------------------------------------
     FUNCTION  Sub_TwosComp  ( CONSTANT A     :  IN STD_LOGIC_VECTOR;
                               CONSTANT B     :  IN STD_LOGIC_VECTOR
                             )  RETURN STD_LOGIC_VECTOR IS 
      VARIABLE r        : STD_LOGIC_VECTOR ( A'LENGTH - 1  DOWNTO 0 );
      VARIABLE bb        : STD_LOGIC_VECTOR (B 'LENGTH - 1  DOWNTO 0 );
      VARIABLE p        : STD_ULOGIC;
      VARIABLE g        : STD_ULOGIC;
      VARIABLE carry    : STD_ULOGIC;
    -- pragma map_to_operator SUB_TC_OP
    -- pragma return_port_name Z
    BEGIN
        -- The operation of (a - b - borrow_in) when a,b are Two's complement
        -- numbers can be computed
        --  as   a + (NOT b + 1) - borrow_in
        --  or   a + (NOT b) + (1-borrow_in)
        --  or   a + (NOT b) + (NOT borrow_in)
    	-- initialization
        bb    := B;
	p     := '1';
	g     := '0';
	carry := '1'; -- for twoscomp sub set carry in '1'  := NOT Borrow_in 
	-- perform operation
       FOR n IN 0 TO A'LENGTH - 1 LOOP
          bb(n) := NOT bb(n);
             p := p AND (A(n) OR bb(n));                        -- Cpropagate
             g := (A(n) AND bb(n)) OR ( g AND (A(n) OR bb(n)));  -- Cgenerate
          r(n) :=  A(n) XOR bb(n) XOR carry;                    -- individual bit sums
         carry :=  g OR (p AND carry);                         -- carry
       END LOOP;
       RETURN r;
    END Sub_TwosComp;
--+-----------------------------------------------------------------------------
--|     Function Name  : Sub_Unsigned
--|  hidden procedure
--|     Overloading    : None
--|
--|     Purpose        : Subtraction of STD_LOGIC_VECTORS.
--|
--|     Parameters     :
--|                      A     - input  STD_LOGIC_VECTOR,
--|                      B     - input  STD_LOGIC_VECTOR,
--|     NOTE           : 
--|                      The inputs may be of any length  but both A  and B
--|                      must have same lengths.
--|                      
--|     Assumptions    : Both inputs must have range (msb downto 0)
--|
--|     Result         : returns STD_LOGIC_VECTOR of the same length as A and B.
--|
--|     Use            : VARIABLE x, y, sum : STD_LOGIC_VECTOR ( 15 DOWNTO 0);
--|                      sum := Sub_Unsigned ( x, y);
--|-----------------------------------------------------------------------------
     FUNCTION  Sub_Unsigned  ( CONSTANT A     :  IN STD_LOGIC_VECTOR;
                               CONSTANT B     :  IN STD_LOGIC_VECTOR
                             )  RETURN STD_LOGIC_VECTOR IS 
      VARIABLE r        : STD_LOGIC_VECTOR ( A'LENGTH - 1  DOWNTO 0 );
      VARIABLE bb        : STD_LOGIC_VECTOR (B 'LENGTH - 1  DOWNTO 0 );
      VARIABLE p        : STD_ULOGIC;
      VARIABLE g        : STD_ULOGIC;
      VARIABLE carry    : STD_ULOGIC;
    -- pragma map_to_operator SUB_UNS_OP
    -- pragma return_port_name Z

    BEGIN
    -- In unsigned mode number is positive, two's comp of positive
    -- is same as unsigned number 
    -- The operation of (a - b - borrow_in) when a,b are Two's complement
    -- numbers can be computed
    --  as   a + (NOT b + 1) - borrow_in
    --  or   a + (NOT b) + (1-borrow_in)
    --  or   a + (NOT b) + (NOT borrow_in)
    -- Initilizations
	p   := '1';
        g   := '0';
        bb  := B;
    -- perform the subtract
      carry :=  '1' ;          -- carry := NOT borrow_in;
      FOR n IN 0 TO A'LENGTH - 1 LOOP
          bb(n) := NOT bb(n);
             p := p AND (A(n) OR bb(n));                         -- Cpropagate
             g := (A(n) AND bb(n)) OR ( g AND (A(n) OR bb(n)));   -- Cgenerate
          r(n) :=  A(n) XOR bb(n) XOR carry;                     -- individual bit sums
         carry :=  g OR (p AND carry);                         -- carry
      END LOOP;
       RETURN r;
    END Sub_Unsigned; 
--+-----------------------------------------------------------------------------
--|     Function Name  : Sub_TwosComp_VHDL_TECH
--|  hidden procedure
--|     Overloading    : None
--|
--|     Purpose        : Two's Complement subtraction of logic vectors.
--|
--|     Parameters     :
--|                      result     - output std_logic_vector, the computed sum
--|                      borrow_out   - output std_logic,
--|                      underflow   - output std_logic, overflow condition
--|                      addend     - input  std_logic_vector,
--|                      augend     - input  std_logic_vector,
--|                      borrow_in   - input std_logic,
--|     NOTE           :
--|                      This procedure is implemented based on hardware design of a
--|                      Two's complement subtractor.
--|                      The inputs may be of any length  but both addend and augend
--|                      must have same lengths.
--|
--|     Use            : VARIABLE x, y, sum : std_logic_vector ( 15 DOWNTO 0);
--|                      VARIABLE borrow, ovf : std_ulogic;
--|
--|                      Sub_TwosComp ( sum, borrow, ovf, x, y, '0' );
--|-----------------------------------------------------------------------------
    PROCEDURE Sub_TwosComp_VHDL_TECH  ( VARIABLE result     : OUT std_logic_vector;
                                        VARIABLE borrow_out : OUT std_ulogic;
                                        VARIABLE underflow  : OUT std_ulogic;
                                        CONSTANT minuend    :  IN std_logic_vector;
                                        CONSTANT subtrahend :  IN std_logic_vector;
                                        CONSTANT borrow_in  :  IN std_ulogic  
                 -- synopsys synthesis_off
                                                        := '0'
                 -- synopsys synthesis_on
                                     ) IS
      CONSTANT reglen   : INTEGER :=  minuend'LENGTH;
      VARIABLE a        : std_logic_vector ( reglen - 1  DOWNTO 0 );
      VARIABLE b        : std_logic_vector ( subtrahend'LENGTH - 1  DOWNTO 0 );
      VARIABLE r        : std_logic_vector ( reglen - 1  DOWNTO 0 );
      VARIABLE p        : std_ulogic;
      VARIABLE g        : std_ulogic;
      VARIABLE c_iminus : std_ulogic;
      VARIABLE carry    : std_ulogic;
    BEGIN
	-- Initializations     
	a   := minuend;
        b   := subtrahend;
        p   := '1';
        g   := '0';
       -- synopsys translate_off
      -- check the length of minuend and subtrahend
      ASSERT   (minuend'LENGTH = subtrahend'LENGTH)
      REPORT " Sub_TwosComp_VHDL_TECH --- operand length not same "
      SEVERITY ERROR;
        -- synopsys translate_on
 
    -- The operation of (a - b - borrow_in) when a,b are Two's complement
    -- numbers can be computed
    --  as   a + (NOT b + 1) - borrow_in
    --  or   a + (NOT b) + (1-borrow_in)
    --  or   a + (NOT b) + (NOT borrow_in)
 
    -- perform the subtract
      carry := NOT borrow_in;
      FOR n IN 0 TO reglen - 1 LOOP
          c_iminus := carry;
          b(n) := NOT b(n);
             p := p AND (a(n) OR b(n));                         -- Cpropagate
             g := (a(n) AND b(n)) OR ( g AND (a(n) OR b(n)));   -- Cgenerate
          r(n) :=  a(n) XOR b(n) XOR carry;                     -- individual bit sums
         carry :=  g OR (p AND carry);                         -- carry
      END LOOP;
      borrow_out := To_X01(NOT carry);
      -- set overflow if carry_in and carry_out of sign bit are different.
         underflow := To_X01( c_iminus XOR carry);
         result := To_X01(r);
       RETURN;
    END Sub_TwosComp_VHDL_TECH;
--+-----------------------------------------------------------------------------
--|     Function Name  : Sub_Unsigned_VHDL_TECH
--|  hidden procedure
--|     Overloading    : None
--|
--|     Purpose        :Subtraction of logic vectors.
--|
--|     Parameters     :
--|                      result     - output std_logic_vector, the computed sum
--|                      borrow_out   - output std_ulogic,
--|                      underflow   - output std_ulogic, overflow condition
--|                      addend     - input  std_logic_vector,
--|                      augend     - input  std_logic_vector,
--|                      borrow_in   - input std_ulogic,
--|     NOTE           :
--|                      The inputs may be of any length  but both addend and augend
--|                      must have same lengths.
--|
--|     Use            : VARIABLE x, y, sum : std_logic_vector ( 15 DOWNTO 0);
--|                      VARIABLE borrow, ovf : std_ulogic;
--|
--|                      Sub_Unsigned_VHDL_TECH ( sum, borrow, ovf, x, y, '0' );
--|-----------------------------------------------------------------------------
    PROCEDURE Sub_Unsigned_VHDL_TECH  ( VARIABLE result     : OUT std_logic_vector;
                              VARIABLE borrow_out : OUT std_ulogic;
                              VARIABLE underflow  : OUT std_ulogic;
                              CONSTANT minuend    :  IN std_logic_vector;
                              CONSTANT subtrahend :  IN std_logic_vector;
                              CONSTANT borrow_in  :  IN std_ulogic 
                 -- synopsys synthesis_off
                                                        := '0'
                 -- synopsys synthesis_on
                            ) IS
      CONSTANT reglen : INTEGER :=  minuend'LENGTH;
      VARIABLE a      : std_logic_vector ( reglen - 1  DOWNTO 0 );
      VARIABLE b      : std_logic_vector ( subtrahend'LENGTH - 1  DOWNTO 0 );
      VARIABLE r      : std_logic_vector ( reglen - 1  DOWNTO 0 );
      VARIABLE p      : std_ulogic;
      VARIABLE g      : std_ulogic;
      VARIABLE carry  : std_ulogic;
    BEGIN
	-- Initializations     
	a   := minuend;
        b   := subtrahend;
        p   := '1';
        g   := '0';
       -- synopsys translate_off
       -- check the length of minuend and subtrahend
      ASSERT   (minuend'LENGTH = subtrahend'LENGTH)
      REPORT " Sub_TwosComp --- operand length not same "
      SEVERITY ERROR;
      -- synopsys translate_on
 
    -- The operation of (a - b - borrow_in) when a,b are Two's complement
    -- numbers can be computed
    --  as   a + (NOT b + 1) - borrow_in
    --  or   a + (NOT b) + (1-borrow_in)
    --  or   a + (NOT b) + (NOT borrow_in)
 
    -- perform the subtract
      carry := NOT borrow_in;
      FOR n IN 0 TO reglen - 1 LOOP
          b(n) := NOT b(n);
             p := p AND (a(n) OR b(n));                         -- Cpropagate
             g := (a(n) AND b(n)) OR ( g AND (a(n) OR b(n)));   -- Cgenerate
          r(n) :=  a(n) XOR b(n) XOR carry;                     -- individual bit sums
         carry :=  g OR (p AND carry);                         -- carry
      END LOOP;
      borrow_out := To_X01(NOT carry);
         underflow := To_X01(NOT carry);
         result := To_X01(r);
        RETURN;
    END Sub_Unsigned_VHDL_TECH;
--+-----------------------------------------------------------------------------
--|     Function Name  : RegAdd_Syn
--|
--|     Overloading    : None
--|
--|     Purpose        : Addition of logic vectors.
--|
--|     Parameters     :
--|                      result     - output std_logic_vector, the computed sum
--|                      addend     - input  std_logic_vector,
--|                      augend     - input  std_logic_vector,
--|                      SrcRegMode - input  regmode_type, indicating the format of
--|                                the input std_logic_vector.   Default is TwosComp.
--|
--|     NOTE           :
--|                      The inputs may be of any length and may be of differing
--|                      lengths.
--|  
--|                    For Synthesis:
--|                      Result is computed with length N (where
--|                      N is the greater of the input vector lengths).
--|                      It is assumed that user will provide result length equal
--|                      to the length of the greater of addend and augend. 
--|                      No error checking has been performed.
--|     Use            :
--|                      VARIABLE x, y, sum : std_logic_vector ( 15 DOWNTO 0);
--| 
--|                      RegAdd_Syn ( sum, x, y, TwosComp );
--|-----------------------------------------------------------------------------
    PROCEDURE RegAdd_Syn  ( VARIABLE result     : INOUT std_logic_vector;
                            CONSTANT addend     : IN std_logic_vector;
                            CONSTANT augend     : IN std_logic_vector;
                            CONSTANT SrcRegMode : IN regmode_type
                 -- synopsys synthesis_off
					           := DefaultRegMode 
                 -- synopsys synthesis_on
                      ) IS

	CONSTANT reslen       : INTEGER := MAXIMUM ( addend'LENGTH, augend'LENGTH );
	VARIABLE a, b, r      : STD_LOGIC_VECTOR ( reslen - 1 DOWNTO 0 );
	VARIABLE  result_copy : STD_LOGIC_VECTOR ( result'Length - 1 DOWNTO 0 );
     BEGIN 
      -- synopsys translate_off
      --   Null range check
      --   if result vector is a null range
        IF ( result'LENGTH = 0) THEN
             ASSERT false
             REPORT " RegAdd_Syn ---  Destination has null range. "
             SEVERITY ERROR;
             RETURN;
      --   if addend or augned or both have null range no need to add
        ELSIF (addend'LENGTH = 0) AND (augend'LENGTH = 0) THEN
             ASSERT false
             REPORT " RegAdd_Syn --- both addend  and augend has null range "
             SEVERITY ERROR;
             result_copy :=  (OTHERS => '0');
             result := result_copy; 
             RETURN;      
        END IF;
      -- synopsys translate_on
      -- if one of the addend or augend is null 
        IF (addend'LENGTH = 0) THEN
      -- synopsys translate_off
             ASSERT false
             REPORT " RegAdd_Syn --- addend has null range "
             SEVERITY ERROR;
      -- synopsys translate_on
             a :=  ( OTHERS => '0');     -- treat it as	zero's            
             b := augend;

        ELSIF (augend'LENGTH = 0) THEN 
      -- synopsys translate_off
             ASSERT false
             REPORT " RegAdd_Syn ---  augend has null range "
             SEVERITY ERROR;
      -- synopsys translate_on
             b :=  (OTHERS => '0');                 
             a := addend;
                 -- inputs are  not null so sign extend them to the same length.  
        ELSE
             a := SignExtend(addend , reslen, addend'LEFT, SrcRegMode);
             b := SignExtend(augend , reslen, augend'LEFT, SrcRegMode);

        END IF;	
       -- Compute the add operation
	if (SrcRegMode = TwosComp) Then
		r := Add_TwosComp (a, b); 
        else
		r := Add_Unsigned (a, b);
        end if;
        result_copy := r(result'length - 1 downto 0);
        result := To_X01(result_copy);
        return;
     END RegAdd_Syn;
--+-----------------------------------------------------------------------------
--|     Function Name  : RegAdd_Syn
--|
--|     Overloading    : None
--|
--|     Purpose        : Addition of logic vectors.
--|
--|     Parameters     :
--|                      result     - output std_ulogic_vector, the computed sum
--|                      addend     - input  std_ulogic_vector,
--|                      augend     - input  std_ulogic_vector,
--|                      SrcRegMode - input  regmode_type, indicating the format of
--|                                the input std_ulogic_vector.   Default is TwosComp.
--|
--|     NOTE           : The inputs may be of any length and may be of differing
--|                      lengths.
--|  
--|                    For Synthesis:
--|                      Result is computed with length N (where
--|                      N is the greater of the input vector lengths).
--|                      It is assumed that user will provide result length equal
--|                      to the length of the greater of addend and augend. 
--|                      No error checking has been performed.
--|     Use            :
--|                      VARIABLE x, y, sum : std_ulogic_vector ( 15 DOWNTO 0);
--| 
--|                      RegAdd_Syn ( sum, x, y, TwosComp );
--|-----------------------------------------------------------------------------
    PROCEDURE RegAdd_Syn  ( VARIABLE result     : INOUT std_ulogic_vector;
                            CONSTANT addend     : IN std_ulogic_vector;
                            CONSTANT augend     : IN std_ulogic_vector;
                            CONSTANT SrcRegMode : IN regmode_type
                 -- synopsys synthesis_off
					           := DefaultRegMode 
                 -- synopsys synthesis_on
                      ) IS
	VARIABLE  reslt : STD_LOGIC_VECTOR ( result'Length - 1 DOWNTO 0 );
	VARIABLE  a_copy : std_logic_vector ( addend'Length - 1 DOWNTO 0 );
	VARIABLE  b_copy : std_logic_vector ( augend'Length - 1 DOWNTO 0 );
   BEGIN 
	a_copy := To_StdLogicVector(addend);
        b_copy := To_StdLogicVector(augend);
        RegAdd_Syn (reslt, a_copy, b_copy, SrcRegMode);
        result := To_StdULogicVector(reslt);
        return;
   END RegAdd_Syn;
--+-----------------------------------------------------------------------------
--|     Function Name  : RegAdd_Syn
--|
--|     Overloading    : None
--|
--|     Purpose        : Addition of BIT_VECTORS.
--|
--|     Parameters     :
--|                      result     - input-output BIT_VECTOR, the computed sum
--|                      addend     - input  BIT_VECTOR,
--|                      augend     - input  BIT_VECTOR,
--|                      SrcRegMode - input  regmode_type, indicating the format of
--|                                the input BIT_VECTOR.   Default is TwosComp.
--|
--|     NOTE           : The inputs may be of any length and may be of differing
--|                      lengths.
--|                    
--|                    For Synthesis:
--|                      Result is computed with length N (where
--|                      N is the greater of the input vector lengths).
--|                      It is assumed that user will provide result length equal
--|                      to the length of the greater of addend and augend. 
--|                      No error checking has been performed.
--|     Use            :
--|                      VARIABLE x, y, sum : BIT_VECTOR ( 15 DOWNTO 0);
--|                      VARIABLE carry_out , ovf: BIT;
--| 
--|                      RegAdd_Syn ( sum, carry_out, ovf,x, y, UnSigned );
--|-----------------------------------------------------------------------------
   PROCEDURE RegAdd_Syn  ( VARIABLE result     : INOUT BIT_VECTOR;
                           CONSTANT addend     : IN BIT_VECTOR;
                           CONSTANT augend     : IN BIT_VECTOR;
                           CONSTANT SrcRegMode : IN regmode_type 
                 -- synopsys synthesis_off
                                                        := DefaultRegMode 
                 -- synopsys synthesis_on
                      ) IS
	VARIABLE  reslt : std_logic_vector ( result'Length - 1 DOWNTO 0 );
	VARIABLE  a_copy : std_logic_vector ( addend'Length - 1 DOWNTO 0 );
	VARIABLE  b_copy : std_logic_vector ( augend'Length - 1 DOWNTO 0 );
   BEGIN 
	a_copy := To_StdLogicVector(addend);
        b_copy := To_StdLogicVector(augend);
        RegAdd_Syn (reslt, a_copy, b_copy, SrcRegMode);
        result := To_BitVector(reslt);
        return;
   END RegAdd_Syn;
--+-----------------------------------------------------------------------------
--|     Function Name  : RegSub_Syn
--|    
--|     Overloading    : None
--|
--|     Purpose        : Subtraction of logic vectors.
--|                       ( result = minuend - subtrahend )
--|
--|     Parameters     :
--|                      result     - input_output std_logic_vector, the computed diff
--|                      minuend    - input  std_logic_vector,
--|                      subtrahend - input  std_logic_vector,
--|                      SrcRegMode - input  regmode_type, indicating the format of
--|                                   the input std_logic_vector.   Default is TwosComp.
--|
--|     NOTE           : The inputs may be of any length and may be of differing
--|                      lengths.
--|
--|                      A temporary result is computed with length N (where
--|                      N is the greater of the input vector lengths).
--|     Use            :
--|                      VARIABLE x, y, diff : std_logic_vector ( 15 DOWNTO 0);
--|                      RegSub_Syn ( diff,  x, y, UnSigned );
--|-----------------------------------------------------------------------------
    PROCEDURE RegSub_Syn  ( VARIABLE result     : INOUT std_logic_vector;
                            CONSTANT minuend    :  IN std_logic_vector;
                            CONSTANT subtrahend :  IN std_logic_vector;
                            CONSTANT SrcRegMode :  IN regmode_type
                 -- synopsys synthesis_off
                                                      := DefaultRegMode 
                 -- synopsys synthesis_on
                      ) IS
      CONSTANT reslen       : INTEGER := MAXIMUM (minuend'LENGTH, subtrahend'LENGTH);
      VARIABLE a, b, r      : STD_LOGIC_VECTOR ( reslen - 1 DOWNTO 0 );
      VARIABLE reslt_copy   : STD_LOGIC_VECTOR ( result'length-1 downto 0);
    BEGIN
    -- synopsys translate_off
     --   Null range check
     --   if result vector is a null range
       IF ( result'LENGTH = 0) THEN
             ASSERT false
             REPORT " RegSub_Syn ---  Destination has null range. " &
                    " cannot save result. "
             SEVERITY ERROR;
             RETURN;

     --   if both minuend and subtrahend  have null range no need to subtract
       ELSIF  (minuend'LENGTH = 0) AND (subtrahend'LENGTH = 0) THEN
             ASSERT false
             REPORT " RegSub_Syn --- both minuend and subtrahend has null range "
             SEVERITY ERROR;
             reslt_copy :=  (OTHERS => '0');
             result := reslt_copy;
             RETURN;
       END IF;
     -- synopsys translate_on
     -- if one of the minuend or subtrahend is null
       IF (minuend'LENGTH = 0) THEN
    -- synopsys translate_off
             ASSERT false
             REPORT " RegSub_Syn --- minuend has null range "
             SEVERITY ERROR;
    -- synopsys translate_on
             a :=  ( OTHERS => '0');     -- treat it as zero's
             b :=  subtrahend ;
 
       ELSIF (subtrahend'LENGTH = 0) THEN
    -- synopsys translate_off
             ASSERT false
             REPORT " RegSub_Syn ---  subtrahend has null range "
             SEVERITY ERROR;
    -- synopsys translate_on
             b :=  (OTHERS => '0');
             a := minuend ;
  
                 -- inputs are  not null so sign extend them to the same length.
       ELSE
             a := SignExtend(minuend , reslen, minuend'LEFT, SrcRegMode);
             b := SignExtend(subtrahend , reslen, subtrahend'LEFT, SrcRegMode);
 
       END IF;
       -- compute the subtraction
	if (SrcRegMode = TwosComp) Then
		r:= Sub_TwosComp (a, b); 
        else
		r:= Sub_Unsigned (a, b);
        end if;
        reslt_copy := r(result'length -1 downto 0);
        result := To_X01(reslt_copy);
        return;
     END RegSub_Syn;
--+-----------------------------------------------------------------------------
--|     Function Name  : RegSub_Syn
--|    
--|     Overloading    : None
--|
--|     Purpose        : Subtraction of ulogic vectors.
--|                       ( result = minuend - subtrahend )
--|
--|     Parameters     :
--|                      result     - input_output std_ulogic_vector, the computed diff
--|                      minuend    - input  std_ulogic_vector,
--|                      subtrahend - input  std_ulogic_vector,
--|                      SrcRegMode - input  regmode_type, indicating the format of
--|                                   the input std_ulogic_vector.   Default is TwosComp.
--|
--|     NOTE           : The inputs may be of any length and may be of differing
--|                      lengths.
--|
--|                      A temporary result is computed with length N (where
--|                      N is the greater of the input vector lengths).
--|     Use            :
--|                      VARIABLE x, y, diff : std_ulogic_vector ( 15 DOWNTO 0);
--|
--|                      RegSub_Syn ( diff, x, y,  UnSigned );
--|-----------------------------------------------------------------------------
    PROCEDURE RegSub_Syn  ( VARIABLE result     : INOUT std_ulogic_vector;
                            CONSTANT minuend    :  IN std_ulogic_vector;
                            CONSTANT subtrahend :  IN std_ulogic_vector;
                            CONSTANT SrcRegMode :  IN regmode_type
                 -- synopsys synthesis_off
                                                      := DefaultRegMode 
                 -- synopsys synthesis_on
                      ) IS
        VARIABLE reslt  : std_logic_vector ( result'length-1 downto 0);
	VARIABLE  a_copy : std_logic_vector ( minuend'Length - 1 DOWNTO 0 );
	VARIABLE  b_copy : std_logic_vector ( subtrahend'Length - 1 DOWNTO 0 );
   BEGIN 
	a_copy := To_StdLogicVector(minuend);
        b_copy := To_StdLogicVector(subtrahend);
        RegSub_Syn (reslt, a_copy, b_copy, SrcRegMode);
        result := To_StdULogicVector(reslt);
        return;
   END RegSub_Syn;
--+-----------------------------------------------------------------------------
--|     Function Name  : RegSub_Syn
--|    
--|     Overloading    : None
--|
--|     Purpose        : Subtraction of BIT_VECTORS.
--|                       ( result = minuend - subtrahend )
--|
--|     Parameters     :
--|                      result     - input-output BIT_VECTOR, the computed sum
--|                      minuend - input  BIT_VECTOR,
--|                      subtrahend - input  BIT_VECTOR,
--|                      SrcRegMode - input  regmode_type, indicating the format of
--|                                the input BIT_VECTOR.   Default is TwosComp.
--|
--|     NOTE           :
--|                      The inputs may be of any length and may be of differing
--|                      lengths.
--|
--|                      A temporary result is computed with length N (where
--|                      N is the greater of the input vector lengths).
--|     Use            :
--|                      VARIABLE x, y, diff : BIT_VECTOR ( 15 DOWNTO 0);
--|
--|                      RegSub_Syn ( diff, x, y, UnSigned );
--|-----------------------------------------------------------------------------
    PROCEDURE RegSub_Syn  ( VARIABLE result     : INOUT BIT_VECTOR;
                            CONSTANT minuend    :  IN BIT_VECTOR;
                            CONSTANT subtrahend :  IN BIT_VECTOR;
                            CONSTANT SrcRegMode :  IN regmode_type
                 -- synopsys synthesis_off
                                                      := DefaultRegMode 
                 -- synopsys synthesis_on
                      ) IS
        VARIABLE reslt  : std_logic_vector ( result'length-1 downto 0);
	VARIABLE  a_copy : std_logic_vector ( minuend'Length - 1 DOWNTO 0 );
	VARIABLE  b_copy : std_logic_vector ( subtrahend'Length - 1 DOWNTO 0 );
   BEGIN 
	a_copy := To_StdLogicVector(minuend);
        b_copy := To_StdLogicVector(subtrahend);
        RegSub_Syn (reslt, a_copy, b_copy, SrcRegMode);
        result     := To_BitVector(reslt);
        return;
    END RegSub_Syn;
--+-----------------------------------------------------------------------------
--|     Function Name  : Mult_TwosComp_ARG
--| hidden function
--|     Overloading    : None
--|
--|     Purpose        : Type propagation function
--|
--|     Parameters     : A - input STD_LOGIC_VECTOR,
--|                      B   -  input STD_LOGIC_VECTOR,
--|-----------------------------------------------------------------------------
    FUNCTION Mult_TwosComp_ARG (  CONSTANT A : IN STD_LOGIC_VECTOR;
                                  CONSTANT B : IN STD_LOGIC_VECTOR
                               ) return STD_LOGIC_VECTOR IS
      VARIABLE Z      : STD_LOGIC_VECTOR( (A'LENGTH + B'LENGTH - 1) downto 0);
	-- pragma return_port_name Z     
     BEGIN 
	return (Z);
     END Mult_TwosComp_ARG;
--+-----------------------------------------------------------------------------
--|     Function Name  : Mult_TwosComp
--| hidden function
--|     Overloading    : None
--|
--|     Purpose        : Multiplication of STD_LOGIC_VECTORS.
--|
--|     Parameters     :
--|                      A - input STD_LOGIC_VECTOR,
--|                      B   -  input STD_LOGIC_VECTOR,
--|     NOTE           :
--|                      The inputs may be of any length and may be of differing
--|                      lengths.
--|
--|     Assumptions    : Both inputs must have range (msb downto 0)
--|
--|    Algorithm       : The multiplication is carried out as follows:
--|
--|                      1) Determine sign of result based on sign of 
--|                         multiploicand and sign  of B.
--|
--|                      2) Convert the A amd B to Unsigned 
--|                         representation.
--|                      
--|                      3) Perform multiplication based on add and shift algorithm.
--|
--|     Result         :
--|                     A  result is computed with length N+M (where
--|                      N,M are the lengths of the A and B).
--|     Use            :
--|                      VARIABLE x, y, prod : STD_LOGIC_VECTOR ( 15 DOWNTO 0);
--|
--|                       prod := Mult_TwosComp (x, y);
--|-----------------------------------------------------------------------------
    FUNCTION Mult_TwosComp (  CONSTANT A : IN STD_LOGIC_VECTOR;
                              CONSTANT B : IN STD_LOGIC_VECTOR
                           ) return STD_LOGIC_VECTOR IS

      CONSTANT reslen      : INTEGER := A'LENGTH + B'LENGTH;
      VARIABLE r           : STD_LOGIC_VECTOR ( reslen - 1  DOWNTO 0 );
      VARIABLE rega        : STD_LOGIC_VECTOR ( A'LENGTH - 1 DOWNTO 0 );
      VARIABLE regb        : STD_LOGIC_VECTOR ( B'LENGTH -1  DOWNTO 0 );
      VARIABLE carry       : STD_ULOGIC;
      VARIABLE nxt_c       : STD_ULOGIC;
      VARIABLE sign_bit    : STD_ULOGIC;
      VARIABLE i           : INTEGER;
	-- pragma map_to_operator MULT_TC_OP
	-- pragma type_function Mult_TwosComp_ARG
	-- pragma return_port_name Z     

     BEGIN 
	-- initialization       
        r    := (OTHERS => '0');
        rega := A;
        regb := B;
	-- inputs are  not null so determine the sign and convert 
	-- the inputs to unsigned  representation.
	sign_bit := rega(rega'LEFT) XOR regb(regb'LEFT);    
	IF (rega(rega'LEFT) /= '0') THEN
		rega := To_Unsign (rega, TwosComp);     
	END IF;

	IF ( regb(regb'LEFT)  /= '0' ) THEN
        	regb := To_Unsign (regb, TwosComp);      
	END IF;
        -- perform the multiply using shift and add.
        -- for each bit of the regb
        FOR k IN 0 TO B'LENGTH - 1 LOOP
        -- if the regb bit is '1' then add the shifted rega
           IF (regb(k) = '1') THEN
               i := k;       -- 'i' is LSB position in result for this add
               carry := '0';
               FOR n IN 0 TO rega'LENGTH - 1 LOOP
                  nxt_c := (rega(n) AND r(i)) OR ( carry AND (rega(n) OR r(i))); -- carry compute
                  r(i) :=  rega(n) XOR r(i) XOR carry;                       -- bit sum
                  carry := nxt_c;
                  i := i + 1;
               END LOOP;
               r(i) := carry;            -- carry out is added to result
           END IF;
        END LOOP;
        -- if the result should be negative, then negate
         IF (sign_bit /='0')  THEN
         	return ( RegNegate (r, TwosComp) );         
         ELSE
		return r;
         END IF;
     END Mult_TwosComp;
--+-----------------------------------------------------------------------------
--|     Function Name  : RegMult_TwosComp
--| hidden procedure
--|     Overloading    : None
--|
--|     Purpose        : Multiplication of STD_LOGIC_VECTORS.
--|
--|     Parameters     :
--|                      result       - output STD_LOGIC_VECTOR, the computed product
--|                      overflow     - output STD_ULOGIC, overflow condition
--|                      multiplicand - input STD_LOGIC_VECTOR,
--|                      multiplier   -  input STD_LOGIC_VECTOR,
--|
--|     NOTE           :
--|                      The inputs may be of any length and may be of differing
--|                      lengths.
--|
--|    Algorithm       : The multiplication is carried out as follows:
--|
--|                      1) Determine sign of result based on sign of 
--|                         multiploicand and sign  of multiplier.
--|
--|                      2) Convert the multiplicand amd multiplier to Unsigned 
--|                         representation.
--|                      
--|                      3) Perform multiplication based on add and shift algorithm.
--|
--|     Result         :
--|                     A  temporary result is computed with length N+M (where
--|                      N,M are the lengths of the multiplicand and multiplier)
--|                      by calling local function Mult_TwosComp or Mult_Unsigned
--|                       
--|                      This computed value is extended or truncated to match
--|                      the width of 'result'. If truncated, the low order bits
--|                      are returned.
--|
--|                      The parameter 'overflow' is set to '1' if the product of the
--|                      two inputs is too large to fit in the parameter result.
--|
--|     Use            :
--|                      VARIABLE x, y, prod : STD_LOGIC_VECTOR ( 15 DOWNTO 0);
--|                      VARIABLE ovfl : STD_ULOGIC;
--|
--|                      RegMult_TwosComp ( prod, ovfl, x, y);
--|-----------------------------------------------------------------------------
    PROCEDURE RegMult_TwosComp ( VARIABLE result       : OUT STD_LOGIC_VECTOR;
                                 VARIABLE overflow     : OUT STD_ULOGIC;
                                 CONSTANT multiplicand : IN STD_LOGIC_VECTOR;
                                 CONSTANT multiplier   : IN STD_LOGIC_VECTOR
                              ) IS
      CONSTANT reslen      : INTEGER := multiplicand'LENGTH + multiplier'LENGTH;
      VARIABLE r           : STD_LOGIC_VECTOR ( reslen - 1  DOWNTO 0 );
      VARIABLE rega        : STD_LOGIC_VECTOR ( multiplicand'LENGTH - 1 DOWNTO 0 );
      VARIABLE regb        : STD_LOGIC_VECTOR ( multiplier'LENGTH -1  DOWNTO 0 );
      VARIABLE carry       : STD_ULOGIC;
      VARIABLE nxt_c       : STD_ULOGIC;
      VARIABLE sign_bit    : STD_ULOGIC;
      VARIABLE overflo     : STD_ULOGIC;  
      VARIABLE i           : INTEGER;
      VARIABLE reslt_copy : STD_LOGIC_VECTOR ( result'length - 1 downto 0 );
     BEGIN 
     --  Initializations
        r        := (OTHERS => '0');
        rega     := multiplicand;
        regb     := multiplier;
        overflo  := '0';
     -- synopsys translate_off
     --   Null range check
     --   if result vector is a null range
       IF ( result'LENGTH = 0) THEN
             ASSERT false
             REPORT " RegMult ---  Destination  to hold the product has null range. "
             SEVERITY ERROR;
             overflow := overflo;
             RETURN;
     --   if both multiplicand  and multiplier  have null range no need to multiply
       ELSIF (multiplicand'LENGTH = 0) AND (multiplier'LENGTH = 0) THEN
             ASSERT false
             REPORT " RegMult --- both multiplicand  and multiplier has null range "
             SEVERITY ERROR;
             reslt_copy :=  (OTHERS => '0');
             result := reslt_copy;                   -- result is filled with zeros
             overflow := overflo;       
             RETURN;      

     -- if one of the multiplicand  or multiplier is null 
       ELSIF (multiplicand'LENGTH = 0) THEN
             ASSERT false
             REPORT " RegMult --- multiplicand  has null range "
             SEVERITY ERROR;
                                 -- treat multiplicand as zero so result is zero 
             reslt_copy := (OTHERS => '0');
             result := reslt_copy;
             overflow := overflo;
             RETURN;
       ELSIF (multiplier'LENGTH = 0) THEN
             ASSERT false
             REPORT " RegMult --- multiplier  has null range "
             SEVERITY ERROR;
                                 -- treat multiplier as zero so result is zero 
             reslt_copy := (OTHERS => '0');
             result := reslt_copy;
             overflow := overflo;
             RETURN;
       END IF;
           
	-- synopsys translate_on
	sign_bit := rega(rega'LEFT) XOR regb(regb'LEFT);    
	-- call function mult_twoscomp 
	r := Mult_TwosComp(rega, regb);
	-- Determine the length of the result to be returned
	--
	IF (result'LENGTH < reslen)   THEN
	                reslt_copy := r(result'LENGTH - 1 DOWNTO 0); 
        	        IF (sign_bit = '0') THEN     -- positive result
                	      FOR j IN result'LENGTH  - 1 TO reslen - 2 LOOP
                        	 if (r(j) = '1') THEN
	                           overflo := '1';
        	                 END IF;
--                	         EXIT WHEN (r(j) = '1');
				if(r(j) = '1')then
					result := reslt_copy;
					overflow := overflo;
					RETURN;
				end if;
	                      END LOOP;
                                              
        	        ELSE                          -- negative result  -128 is valid
                	       FOR j IN result'LENGTH  TO reslen - 2 LOOP
                        	  if (r(j) = '0') THEN
	                             overflo := '1';
        	                  END IF;
--                	         EXIT WHEN (r(j) = '0');
				if (r(j) = '0') then
					result := reslt_copy;
					overflow := overflo;
					RETURN;
				end if;
	                       END LOOP;
        	        END IF;
                                         
	ELSIF (result'LENGTH > reslen) THEN                -- sign extend the product
		reslt_copy := SignExtend(r, result'LENGTH, r'Left, TwosComp);
        ELSE
		reslt_copy := r;                              -- equal length
	END IF;
        result := reslt_copy;
        overflow := overflo;
        RETURN;
    END RegMult_TwosComp;
--+-----------------------------------------------------------------------------
--|     Function Name  : Mult_Unsigned
--| hidden function
--|     Overloading    : None
--|
--|     Purpose        : Multiplication of STD_LOGIC_VECTORS.
--|
--|     Parameters     :
--|                      A - input STD_LOGIC_VECTOR,
--|                      B   -  input STD_LOGIC_VECTOR,
--|     NOTE           :
--|                      The inputs may be of any length and may be of differing
--|                      lengths.
--|
--|     Assumptions    : Both inputs must have range (msb downto 0)
--|
--|                      Perform multiplication based on add and shift algorithm.
--|
--|     Result         :
--|                     A  result is computed with length N+M (where
--|                      N,M are the lengths of the A and B).
--|     Use            :
--|                      VARIABLE x, y, prod : STD_LOGIC_VECTOR ( 15 DOWNTO 0);
--|
--|                       prod := Mult_Unsigned (x, y);
--|-----------------------------------------------------------------------------
    FUNCTION Mult_Unsigned (  CONSTANT A : IN STD_LOGIC_VECTOR;
                              CONSTANT B : IN STD_LOGIC_VECTOR
                           ) return STD_LOGIC_VECTOR IS
      CONSTANT reslen      : INTEGER := A'LENGTH + B'LENGTH;
      VARIABLE r           : STD_LOGIC_VECTOR ( reslen - 1  DOWNTO 0 );
      VARIABLE carry       : STD_ULOGIC;
      VARIABLE nxt_c       : STD_ULOGIC;
      VARIABLE sign_bit    : STD_ULOGIC;
      VARIABLE i           : INTEGER;
	-- pragma map_to_operator MULT_UNS_OP
	-- pragma return_port_name Z     
     BEGIN 
	-- initialization       
        r    := (OTHERS => '0');
        FOR k IN 0 TO B'LENGTH - 1 LOOP
        -- if the B bit is '1' then add the shifted A
           IF (B(k) = '1') THEN
               i := k;       -- 'i' is LSB position in result for this add
               carry := '0';
               FOR n IN 0 TO A'LENGTH - 1 LOOP
                  nxt_c := (A(n) AND r(i)) OR ( carry AND (A(n) OR r(i))); -- carry compute
                  r(i) :=  A(n) XOR r(i) XOR carry;                       -- bit sum
                  carry := nxt_c;
                  i := i + 1;
               END LOOP;
               r(i) := carry;            -- carry out is added to result
           END IF;
        END LOOP;
	return r;
     END Mult_Unsigned;
--+-----------------------------------------------------------------------------
--|     Function Name  : RegMult_Unsigned
--|
--|     Overloading    : None
--|
--|     Purpose        : Multiplication of STD_LOGIC_VECTORS.
--|
--|     Parameters     :
--|                      result       - output STD_LOGIC_VECTOR, the computed product
--|                      overflow     - output STD_ULOGIC, overflow condition
--|                      multiplicand - input STD_LOGIC_VECTOR,
--|                      multiplier   -  input STD_LOGIC_VECTOR,
--|
--|     NOTE           :
--|                      The inputs may be of any length and may be of differing
--|                      lengths.
--|
--|    Algorithm       : The multiplication is carried out as follows:
--|
--|                      1) Determine sign of result based on sign of 
--|                         multiploicand and sign  of multiplier.
--|
--|                      2) Convert the multiplicand amd multiplier to Unsigned 
--|                         representation.
--|                      
--|                      3) Perform multiplication based on add and shift algorithm.
--|
--|     Result         :
--|                     A  temporary result is computed with length N+M (where
--|                      N,M are the lengths of the multiplicand and multiplier)
--|                      by calling local function Mult_TwosComp or Mult_Unsigned
--|                       
--|                      This computed value is extended or truncated to match
--|                      the width of 'result'. If truncated, the low order bits
--|                      are returned.
--|
--|                      The parameter 'overflow' is set to '1' if the product of the
--|                      two inputs is too large to fit in the parameter result.
--|
--|     Use            :
--|                      VARIABLE x, y, prod : STD_LOGIC_VECTOR ( 15 DOWNTO 0);
--|                      VARIABLE ovfl : STD_ULOGIC;
--|
--|                      RegMult_Unsigned( prod, ovfl, x, y);
--|-----------------------------------------------------------------------------
    PROCEDURE RegMult_Unsigned ( VARIABLE result       : OUT STD_LOGIC_VECTOR;
                                 VARIABLE overflow     : OUT STD_ULOGIC;
                                 CONSTANT multiplicand : IN STD_LOGIC_VECTOR;
                                 CONSTANT multiplier   : IN STD_LOGIC_VECTOR
                               ) IS
      CONSTANT reslen      : INTEGER := multiplicand'LENGTH + multiplier'LENGTH;
      VARIABLE r           : STD_LOGIC_VECTOR ( reslen - 1  DOWNTO 0 );
      VARIABLE rega        : STD_LOGIC_VECTOR ( multiplicand'LENGTH - 1 DOWNTO 0 );
      VARIABLE regb        : STD_LOGIC_VECTOR ( multiplier'LENGTH -1  DOWNTO 0 );
      VARIABLE carry       : STD_ULOGIC;
      VARIABLE nxt_c       : STD_ULOGIC;
      VARIABLE sign_bit    : STD_ULOGIC;
      VARIABLE overflo     : STD_ULOGIC;  
      VARIABLE i           : INTEGER;
      VARIABLE reslt_copy : STD_LOGIC_VECTOR ( result'length - 1 downto 0 );
     BEGIN 
     --  Initializations
        r        := (OTHERS => '0');
        rega     := multiplicand;
        regb     := multiplier;
        overflo  := '0';
     -- synopsys translate_off
     --   Null range check
     --   if result vector is a null range
       IF ( result'LENGTH = 0) THEN
             ASSERT false
             REPORT " RegMult ---  Destination  to hold the product has null range. "
             SEVERITY ERROR;
             overflow := overflo;
             RETURN;
     --   if both multiplicand  and multiplier  have null range no need to multiply
       ELSIF (multiplicand'LENGTH = 0) AND (multiplier'LENGTH = 0) THEN
             ASSERT false
             REPORT " RegMult --- both multiplicand  and multiplier has null range "
             SEVERITY ERROR;
             reslt_copy :=  (OTHERS => '0');
             result := reslt_copy;                   -- result is filled with zeros
             overflow := overflo;       
             RETURN;      

     -- if one of the multiplicand  or multiplier is null 
       ELSIF (multiplicand'LENGTH = 0) THEN
             ASSERT false
             REPORT " RegMult --- multiplicand  has null range "
             SEVERITY ERROR;
                                 -- treat multiplicand as zero so result is zero 
             reslt_copy := (OTHERS => '0');
             result := reslt_copy;
             overflow := overflo;
             RETURN;
       ELSIF (multiplier'LENGTH = 0) THEN
             ASSERT false
             REPORT " RegMult --- multiplier  has null range "
             SEVERITY ERROR;
                                 -- treat multiplier as zero so result is zero 
             reslt_copy := (OTHERS => '0');
             result := reslt_copy;
             overflow := overflo;
             RETURN;
       END IF;
           
	-- synopsys translate_on
	-- call function  mult_unsigned 
	r := Mult_Unsigned(rega, regb);
	-- Determine the length of the result to be returned
	--
	IF (result'LENGTH < reslen)   THEN
               reslt_copy := r(result'LENGTH - 1 DOWNTO 0); 
               FOR j IN result'LENGTH TO reslen - 1 LOOP
                   if (r(j) /= '0') THEN
                        overflo := '1';
                   END IF;
--                   EXIT WHEN (r(j) /= '0');
			if(r(j) /= '0')then
				result := reslt_copy;
				overflow := overflo;
				RETURN;
			end if;
               END LOOP;
	ELSIF (result'LENGTH > reslen) THEN                -- zero extend the product
		reslt_copy := RegFill_Zero(r, result'LENGTH);
        ELSE
		reslt_copy := r;                              -- equal length
	END IF;
        result := reslt_copy;
        overflow := overflo;
        RETURN;
    END RegMult_Unsigned;
--+-----------------------------------------------------------------------------
--|     Function Name  : RegShift_Left
--| 
--|     Overloading    : None
--|
--|     Purpose        : Logical shift left operator for   BIT_VECTORS.
--|
--|     Parameters     :
--|                      SrcReg      - input  BIT_VECTOR, vector to be shifted
--|                      DstReg      - Input_ouput, BIT_VECTOR, shifted result
--|                      ShiftO      - output, BIT, holds the last bit shifted out 
--|                                          of register
--|                      FillVal    -- input BIT, value to be shifted in
--|                      Nbits       - input , NATURAL, number of positions to shift
--|                                          default is 1.
--|
--|     Result         : Shifted bit_vector
--|
--|     Use            : VARIABLE acc   : BIT_VECTOR ( 15 DOWNTO 0);
--|                      VARIABLE carry : BIT;
--|
--|                      RegShift_Left ( acc, acc, carry,'0', 3 );
--|-----------------------------------------------------------------------------
   PROCEDURE RegShift_Left  ( CONSTANT SrcReg    : IN BIT_VECTOR;
                              VARIABLE DstReg    : INOUT BIT_VECTOR;
                              VARIABLE ShiftO    : OUT BIT; 
                              CONSTANT FillVal   : IN BIT;
                              CONSTANT Nbits     : IN Natural 
		-- synopsys synthesis_off
                                                          := 1
		-- synopsys synthesis_on
                      ) IS 
      VARIABLE r         : BIT_VECTOR (SrcReg'Length - 1 DOWNTO 0);
      VARIABLE src_copy  : BIT_VECTOR (SrcReg'Length - 1 DOWNTO 0 );
   BEGIN
    -- initialization
      src_copy := SrcReg;
     -- None of the registers is null, perform shift operation
	for i IN Nbits - 1 downto 0 Loop
		r(i) := FillVal;
        end loop;
	for i IN SrcReg'Length - 1 downto Nbits Loop
		r(i) := src_copy(i - Nbits);
        end loop;
        ShiftO := src_copy(SrcReg'Length - Nbits);
        DstReg := r;
        RETURN;
   END RegShift_Left;
--+-----------------------------------------------------------------------------
--|     Function Name  : RegShift_Left
--| 
--|     Overloading    : None
--|
--|     Purpose        : Logical shift left operator for   STD_LOGIC_VECTORS.
--|
--|     Parameters     :
--|                      SrcReg      - input  STD_LOGIC_VECTOR, vector to be shifted
--|                      DstReg      - Input_ouput, STD_LOGIC_VECTOR, shifted result
--|                      ShiftO      - output, std_ulogic, holds the last bit shifted out 
--|                                          of register
--|                      FillVal    -- input std_ulogic, value to be shifted in
--|                      Nbits       - input , NATURAL, number of positions to shift
--|                                          default is 1.
--|
--|     Result         : Shifted std_logic_vector
--|
--|     Use            : VARIABLE acc   : STD_LOGIC_VECTOR ( 15 DOWNTO 0);
--|                      VARIABLE carry : std_ulogic;
--|
--|                      RegShift_Left ( acc, acc, carry, '0', 3 );
--|-----------------------------------------------------------------------------
   PROCEDURE RegShift_Left  ( CONSTANT SrcReg    : IN STD_LOGIC_VECTOR;
                              VARIABLE DstReg    : INOUT STD_LOGIC_VECTOR;
                              VARIABLE ShiftO    : OUT STD_ULOGIC; 
                              CONSTANT FillVal   : IN STD_ULOGIC;
                              CONSTANT Nbits     : IN Natural 
		-- synopsys synthesis_off
                                                          := 1
		-- synopsys synthesis_on
                      ) IS 
      VARIABLE r         : STD_LOGIC_VECTOR (SrcReg'Length - 1 DOWNTO 0);
      VARIABLE src_copy  : STD_LOGIC_VECTOR (SrcReg'Length - 1 DOWNTO 0 );

   BEGIN
    -- initialization
      src_copy := SrcReg;
     -- None of the registers is null, perform shift operation
	for i IN Nbits - 1 downto 0 Loop
		r(i) := FillVal;
        end loop;
	for i IN SrcReg'Length - 1 downto Nbits Loop
		r(i) := src_copy(i - Nbits);
        end loop;
        ShiftO := src_copy(SrcReg'Length - Nbits);
        DstReg := r;
        RETURN;
   END RegShift_Left;
--+-----------------------------------------------------------------------------
--|     Function Name  : RegShift_Left
--| 
--|     Overloading    : None
--|
--|     Purpose        : Logical shift left operator for   STD_ULOGIC_VECTORS.
--|
--|     Parameters     :
--|                      SrcReg      - input  STD_ULOGIC_VECTOR, vector to be shifted
--|                      DstReg      - Input_ouput, STD_ULOGIC_VECTOR, shifted result
--|                      ShiftO      - output, std_ulogic, holds the last bit shifted out 
--|                                          of register
--|                      FillVal    -- input std_ulogic, value to be shifted in
--|                      Nbits       - input , NATURAL, number of positions to shift
--|                                          default is 1.
--|
--|     Result         : Shifted std_ulogic_vector
--|
--|     Use            : VARIABLE acc   : STD_ULOGIC_VECTOR ( 15 DOWNTO 0);
--|                      VARIABLE carry : std_ulogic;
--|
--|                      RegShift_Left ( acc, acc, carry, '0', 3 );
--|-----------------------------------------------------------------------------
   PROCEDURE RegShift_Left  ( CONSTANT SrcReg    : IN STD_ULOGIC_VECTOR;
                              VARIABLE DstReg    : INOUT STD_ULOGIC_VECTOR;
                              VARIABLE ShiftO    : OUT STD_ULOGIC; 
                              CONSTANT FillVal   : IN STD_ULOGIC;
                              CONSTANT Nbits     : IN Natural 
		-- synopsys synthesis_off
                                                          := 1
		-- synopsys synthesis_on
                      ) IS 
      VARIABLE r         : STD_ULOGIC_VECTOR (SrcReg'Length - 1 DOWNTO 0);
      VARIABLE src_copy  : STD_ULOGIC_VECTOR (SrcReg'Length - 1 DOWNTO 0 );

   BEGIN
    -- initialization
      src_copy := SrcReg;
     -- None of the registers is null, perform shift operation
	for i IN Nbits - 1 downto 0 Loop
		r(i) := FillVal;
        end loop;
	for i IN SrcReg'Length - 1 downto Nbits Loop
		r(i) := src_copy(i - Nbits);
        end loop;
        ShiftO := src_copy(SrcReg'Length - Nbits);
        DstReg := r;
        RETURN;
   END RegShift_Left;
--+-----------------------------------------------------------------------------
--|     Function Name  : RegShift_right
--| 
--|     Overloading    : None
--|
--|     Purpose        : Logical shift right operator for   BIT_VECTORS.
--|
--|     Parameters     :
--|                      SrcReg      - input  BIT_VECTOR, vector to be shifted
--|                      DstReg      - Input_ouput, BIT_VECTOR, shifted result
--|                      ShiftO      - output, BIT, holds the last bit shifted out 
--|                                          of register
--|                      FillVal    -- input BIT, value to be shifted in
--|                      Nbits       - input , NATURAL, number of positions to shift
--|                                          default is 1.
--|
--|     Result         : Shifted bit_vector
--|
--|     Use            : VARIABLE acc   : BIT_VECTOR ( 15 DOWNTO 0);
--|                      VARIABLE carry : BIT;
--|
--|                      RegShift_right ( acc, acc, carry, '0', 1);
--|-----------------------------------------------------------------------------
   PROCEDURE RegShift_right  ( CONSTANT SrcReg    : IN BIT_VECTOR;
                               VARIABLE DstReg    : INOUT BIT_VECTOR;
                               VARIABLE ShiftO    : OUT BIT; 
                               CONSTANT FillVal   : IN BIT;
                               CONSTANT Nbits     : IN Natural 
		-- synopsys synthesis_off
                                                          := 1
		-- synopsys synthesis_on
                      ) IS 
      VARIABLE r         : BIT_VECTOR (SrcReg'Length - 1 DOWNTO 0);
      VARIABLE src_copy  : BIT_VECTOR (SrcReg'Length - 1 DOWNTO 0 );
    BEGIN
    -- initialization
      src_copy := SrcReg;
    -- shift right
       For i In SrcReg'LENGTH - 1 downto SrcReg'Length - Nbits Loop
		r(i) := FillVal;
       end loop;
       For i IN SrcReg'LENGTH - Nbits - 1 downto 0  Loop
		r(i) := src_copy(i+ Nbits);
       end Loop;
       ShiftO := src_copy(Nbits - 1);
       DstReg := r;
       RETURN;
    END RegShift_Right;
--+-----------------------------------------------------------------------------
--|     Function Name  : RegShift_right
--| 
--|     Overloading    : None
--|
--|     Purpose        : Logical shift right operator for   STD_LOGIC_VECTORS.
--|
--|     Parameters     :
--|                      SrcReg      - input  STD_LOGIC_VECTOR, vector to be shifted
--|                      DstReg      - Input_ouput, STD_LOGIC_VECTOR, shifted result
--|                      ShiftO      - output, std_ulogic, holds the last bit shifted out 
--|                                          of register
--|                      FillVal    -- input std_ulogic, value to be shifted in
--|                      Nbits       - input , NATURAL, number of positions to shift
--|                                          default is 1.
--|
--|     Result         : Shifted std_logic_vector
--|
--|     Use            : VARIABLE acc   : STD_LOGIC_VECTOR ( 15 DOWNTO 0);
--|                      VARIABLE carry : std_ulogic;
--|
--|                      RegShift_right ( acc, acc, carry, '0', 1);
--|-----------------------------------------------------------------------------
   PROCEDURE RegShift_right  ( CONSTANT SrcReg    : IN STD_LOGIC_VECTOR;
                               VARIABLE DstReg    : INOUT STD_LOGIC_VECTOR;
                               VARIABLE ShiftO    : OUT std_ulogic; 
                               CONSTANT FillVal   : IN std_ulogic;
                               CONSTANT Nbits     : IN Natural 
		-- synopsys synthesis_off
                                                          := 1
		-- synopsys synthesis_on
                      ) IS 
      VARIABLE r         : STD_LOGIC_VECTOR (SrcReg'Length - 1 DOWNTO 0);
      VARIABLE src_copy  : STD_LOGIC_VECTOR (SrcReg'Length - 1 DOWNTO 0 );
    BEGIN
    -- initialization
      src_copy := SrcReg;
    -- shift right
       For i In SrcReg'LENGTH - 1 downto SrcReg'Length - Nbits Loop
		r(i) := FillVal;
       end loop;
       For i IN SrcReg'LENGTH - Nbits - 1 downto 0  Loop
		r(i) := src_copy(i+ Nbits);
       end Loop;
       ShiftO := src_copy(Nbits - 1);
       DstReg := r;
       RETURN;
    END RegShift_Right;
--+-----------------------------------------------------------------------------
--|     Function Name  : RegShift_right
--| 
--|     Overloading    : None
--|
--|     Purpose        : Logical shift right operator for   STD_ULOGIC_VECTORS.
--|
--|     Parameters     :
--|                      SrcReg      - input  STD_ULOGIC_VECTOR, vector to be shifted
--|                      DstReg      - Input_ouput, STD_ULOGIC_VECTOR, shifted result
--|                      ShiftO      - output, std_ulogic, holds the last bit shifted out 
--|                                          of register
--|                      FillVal    -- input std_ulogic, value to be shifted in
--|                      Nbits       - input , NATURAL, number of positions to shift
--|                                          default is 1.
--|
--|     Result         : Shifted std_ulogic_vector
--|
--|     Use            : VARIABLE acc   : STD_ULOGIC_VECTOR ( 15 DOWNTO 0);
--|                      VARIABLE carry : std_ulogic;
--|
--|                      RegShift_right ( acc, acc, carry, '0', 1);
--|-----------------------------------------------------------------------------
   PROCEDURE RegShift_right  ( CONSTANT SrcReg    : IN STD_ULOGIC_VECTOR;
                               VARIABLE DstReg    : INOUT STD_ULOGIC_VECTOR;
                               VARIABLE ShiftO    : OUT std_ulogic; 
                               CONSTANT FillVal   : IN std_ulogic;
                               CONSTANT Nbits     : IN Natural 
		-- synopsys synthesis_off
                                                          := 1
		-- synopsys synthesis_on
                      ) IS 
      VARIABLE r         : STD_ULOGIC_VECTOR (SrcReg'Length - 1 DOWNTO 0);
      VARIABLE src_copy  : STD_ULOGIC_VECTOR (SrcReg'Length - 1 DOWNTO 0 );
    BEGIN
    -- initialization
      src_copy := SrcReg;
    -- shift right
       For i In SrcReg'LENGTH - 1 downto SrcReg'Length - Nbits Loop
		r(i) := FillVal;
       end loop;
       For i IN SrcReg'LENGTH - Nbits - 1 downto 0  Loop
		r(i) := src_copy(i+ Nbits);
       end Loop;
       ShiftO := src_copy(Nbits - 1);
       DstReg := r;
       RETURN;
    END RegShift_Right;
     -------------------------------------------------------------------------------
     --     Function Name : Overloaded "+" operator
     -- 1.3.3    
     --     Purpose       : Addition operator for logic vectors.
     --     
     --     Parameters    :     result            left              right
     --                       std_logic_vector    std_logic_vector  std_logic_vector
     --     
     --     NOTE          : Addition is performed in DefaultRegMode  which is set
     --                     to Two's complement. 
     --                     The operands may be of different length. The length of
     --                     the result equals the length of the longer operand.
     --     
     --                     Any overflow condition and carry_out is ignored
     --     
     --     Use           : 
     --                      VARIABLE a,b,c : std_logic_vector ( 7 downto 0 );
     --                      c := a + b;
     --                      c := a + B"0101";  -- c = a + 5;
     --                      c := a + B"101";   -- c = a + (-3)
     --
     --     See Also      : RegAdd, RegSub, RegInc, RegDec, RegNegate
     -------------------------------------------------------------------------------
     FUNCTION  "+" ( CONSTANT addend       : IN std_logic_vector;
		     CONSTANT augend       : IN std_logic_vector
		   ) RETURN std_logic_vector IS
       CONSTANT reslen    : INTEGER := MAXIMUM (addend'LENGTH, augend'LENGTH);
       VARIABLE result    : std_logic_vector (reslen - 1 DOWNTO 0); 
     BEGIN
     --
     -- Use the RegAdd_Syn procedure notation
	 RegAdd_Syn ( result, addend, augend, DefaultRegMode);
	 RETURN result;
     END;
     -------------------------------------------------------------------------------
     --     Function Name : Overloaded "+" operator
     -- 1.3.4
     --     Purpose       : Addition operator for logic vectors.
     --
     --     Parameters    :     result         left                   right
     --                       std_logic_vector    std_logic_vector  Integer
     --
     --     NOTE          : The addition operation is performed assuming all
     --                     operands and results are in DefaultRegMode which
     --                     is set to Two's complement.
     --
     --                     The augend is converted to Std_logic_vector of length
     --                     equal to the addend. The length of 
     --                     the result equals the length of the addend.
     --
     --                     Any overflow condition is reported.
     --
     --     Use           :
     --                      VARIABLE a,c : std_logic_vector ( 7 downto 0 );
     --                      VARIABLE b: Integer; 
     --                      c := a + b;
     --                      c := a + 5;
     --
     --     See Also      : RegAdd, RegSub, RegInc, RegDec, RegNegate
     -------------------------------------------------------------------------------
     FUNCTION  "+" ( CONSTANT addend       : IN std_logic_vector;
		     CONSTANT augend       : IN Integer
		   ) RETURN std_logic_vector IS
       VARIABLE result    : std_logic_vector (addend'LENGTH - 1 DOWNTO 0); 
       VARIABLE aug_copy  : std_logic_vector (addend'LENGTH - 1 DOWNTO 0); 
     BEGIN
       -- Convert augend from Integer to std_logic_vector
	aug_copy := To_StdLogicVector(augend, addend'LENGTH, DefaultRegMode);	     		
       -- Use the RegAdd_Syn procedure with DefaultRegMode mode
	RegAdd_Syn (result, addend, aug_copy,  DefaultRegMode);
	RETURN result;
     END;
     -------------------------------------------------------------------------------
     --     Function Name : Overloaded "+" operator
     --  1.3.5
     --     Purpose       : Addition operator for logic vectors.
     --
     --     Parameters    :     result         left       right
     --                       std_logic_vector   Integer   std_logic_vector
     --
     --     NOTE          : The addition operation is performed assuming all
     --                     operands and results are 
     --                        
     --
     --                     The addend is converted to Std_logic_vector of length
     --                     equal to the augend. The length of 
     --                     the result equals the length of the augend
     --
     --                     Any overflow condition is ignored.
     --
     --     Use           :
     --                      VARIABLE a: Integer; 
     --                      VARIABLE b,c : std_logic_vector ( 7 downto 0 );
     --                      c := a + b;
     --                      c := 5 + b;
     --
     --     See Also      : RegAdd, RegSub, RegInc, RegDec, RegNegate
     -------------------------------------------------------------------------------
     FUNCTION  "+" ( CONSTANT addend       : IN Integer;
		     CONSTANT augend       : IN std_logic_vector
		   ) RETURN std_logic_vector IS
       VARIABLE result 	 : std_logic_vector (augend'LENGTH - 1 DOWNTO 0); 
       VARIABLE a_copy 	 : std_logic_vector (augend'LENGTH - 1 DOWNTO 0); 
     BEGIN
     -- Convert addend from Integer to std_logic_vector
	a_copy := To_StdLogicVector(addend, augend'LENGTH, DefaultRegMode);
     -- Use the RegAdd_Syn procedure with  DefaultRegMode mode
	RegAdd_Syn (result, a_copy, augend, DefaultRegMode);
	RETURN result;
     END;
     -------------------------------------------------------------------------------
     --     Function Name : Overloaded "+" operator
     -- 1.3.3    
     --     Purpose       : Addition operator for std_ulogic_vectors.
     --     
     --     Parameters    :     result            left              right
     --                     std_ulogic_vector  std_ulogic_vector  std_ulogic_vector
     --     
     --     NOTE          : Addition is performed in DefaultRegMode  which is set
     --                     to Two's complement. 
     --                     The operands may be of different length. The length of
     --                     the result equals the length of the longer operand.
     --     
     --                     Any overflow condition and carry_out is ignored
     --     
     --     Use           : 
     --                      VARIABLE a,b,c : std_ulogic_vector ( 7 downto 0 );
     --                      c := a + b;
     --                      c := a + B"0101";  -- c = a + 5;
     --                      c := a + B"101";   -- c = a + (-3)
     --
     --     See Also      : RegAdd, RegSub, RegInc, RegDec, RegNegate
     -------------------------------------------------------------------------------
     FUNCTION  "+" ( CONSTANT addend       : IN std_ulogic_vector;
		     CONSTANT augend       : IN std_ulogic_vector
		   ) RETURN std_ulogic_vector IS
       CONSTANT reslen    : INTEGER := MAXIMUM (addend'LENGTH, augend'LENGTH);
       VARIABLE result    : std_ulogic_vector (reslen - 1 DOWNTO 0); 
     BEGIN
     -- Use the RegAdd_Syn procedure with  DefaultRegMode notation
	RegAdd_Syn (result, addend, augend, DefaultRegMode);
	RETURN result;
     END;
     -------------------------------------------------------------------------------
     --     Function Name : Overloaded "+" operator
     -- 1.3.4
     --     Purpose       : Addition operator for std_ulogic vectors.
     --
     --     Parameters    :     result         left                   right
     --                    std_ulogic_vector  std_ulogic_vector    Integer
     --
     --     NOTE          : The addition operation is performed assuming all
     --                     operands and results are signed Two's complement integers.
     --
     --                     The augend is converted to Std_ulogic_vector of length
     --                     equal to the addend. The length of 
     --                     the result equals the length of the addend.
     --
     --                     Any overflow condition is reported.
     --
     --     Use           :
     --                      VARIABLE a,c : std_ulogic_vector ( 7 downto 0 );
     --                      VARIABLE b: Integer; 
     --                      c := a + b;
     --                      c := a + 5;
     --
     --     See Also      : RegAdd, RegSub, RegInc, RegDec, RegNegate
     -------------------------------------------------------------------------------
     FUNCTION  "+" ( CONSTANT addend       : IN std_ulogic_vector;
		     CONSTANT augend       : IN Integer
		   ) RETURN std_ulogic_vector IS
       VARIABLE result    : std_ulogic_vector (addend'LENGTH - 1 DOWNTO 0); 
       VARIABLE aug_copy  : std_ulogic_vector (addend'LENGTH - 1 DOWNTO 0); 
     BEGIN
     -- Convert augend from Integer to std_ulogic_vector
	aug_copy := To_StdULogicVector(augend,addend'LENGTH,DefaultRegMode);
     -- Use the RegAdd_Syn procedure with DefaultRegMode 
	RegAdd_Syn (result, addend, aug_copy, DefaultRegMode);
	RETURN result;
     END;
     -------------------------------------------------------------------------------
     --     Function Name : Overloaded "+" operator
     --  
     --     Purpose       : Addition operator for std_ulogic vectors.
     --
     --     Parameters    :     result         left       right
     --                    std_ulogic_vector   Integer   std_ulogic_vector
     --
     --     NOTE          : The addition operation is performed assuming all
     --                     operands and results are signed Two's complement integers.
     --
     --                     The addend is converted to Std_ulogic_vector of length
     --                     equal to the augend. The length of 
     --                     the result equals the length of the augend
     --
     --                     Any overflow condition is ignored.
     --
     --     Use           :
     --                      VARIABLE a: Integer; 
     --                      VARIABLE b,c : std_ulogic_vector ( 7 downto 0 );
     --                      c := a + b;
     --                      c := 5 + b;
     --
     --     See Also      : RegAdd, RegSub, RegInc, RegDec, RegNegate
     -------------------------------------------------------------------------------
     FUNCTION  "+" ( CONSTANT addend       : IN Integer;
		     CONSTANT augend       : IN std_ulogic_vector
		   ) RETURN std_ulogic_vector IS
       VARIABLE result 	 : std_ulogic_vector (augend'LENGTH - 1 DOWNTO 0); 
       VARIABLE a 	 : std_ulogic_vector (augend'LENGTH - 1 DOWNTO 0); 
     BEGIN
     -- Convert addend from Integer to std_ulogic_vector
	a := To_StdULogicVector(addend, augend'LENGTH, DefaultRegMode);
     -- Use the RegAdd_Syn procedure with   DefaultRegMode
	RegAdd_Syn (result, a, augend, DefaultRegMode);
	RETURN result;
     END;
     ---------------------------------------------------------------------------------
     --     Function Name : Overloaded "+" operator
     -- 1.3.6 
     --     Purpose       : Addition operator for bit vectors.
     --
     --     Parameters    :     result         left       right
     --                        bit_vector    bit_vector   bit_vector 
     --
     --     NOTE          : The addition operation is performed assuming all
     --                     operands and results are signed Two's complement integers.
     --
     --                     The operands may be of different length. The length of
     --                     the result equals the length of the longer operand.
     --
     --                     Any overflow condition is ignored.
     --
     --     Use           :
     --                      VARIABLE a,b,c : bit_vector ( 7 downto 0 );
     --                      c := a + b;
     --                      c := a + B"0101";  -- c = a + 5;
     --                      c := a + B"101";   -- c = a + (-3)
     --
     --     See Also      : RegAdd, RegSub, RegInc, RegDec, RegNegate
    -------------------------------------------------------------------------------
     FUNCTION  "+" ( CONSTANT addend       : IN bit_vector;
		     CONSTANT augend       : IN bit_vector
		   ) RETURN bit_vector IS
       CONSTANT reslen : INTEGER := MAXIMUM (addend'LENGTH, augend'LENGTH);
       VARIABLE result : bit_vector (reslen - 1  DOWNTO 0);
     BEGIN
     -- Use the RegAdd_Syn with   DefaultRegMode 
	RegAdd_Syn (result, addend, augend, DefaultRegMode);
	return result;
     END;
     ---------------------------------------------------------------------------------
     --     Function Name : Overloaded "+" operator
     -- 1.3.7
     --     Purpose       : Addition operator for bit vectors.
     --
     --     Parameters    :     result         left       right
     --                        bit_vector    bit_vector   Integer 
     --
     --     NOTE          : The addition operation is performed assuming all
     --                     operands and results are signed Two's complement integers.
     --
     --                     The augend is converted to bit_vector of length
     --                     equal to the addend. The length of 
     --                     the result equals the length of the addend.
     --
     --                     Any overflow condition is ignored.
     --
     --     Use           :
     --                      VARIABLE a,c : bit_vector ( 7 downto 0 );
     --                      VARIABLE b: Integer; 
     --                      c := a + b;
     --                      c := a + 5;
     --
     --     See Also      : RegAdd, RegSub, RegInc, RegDec, RegNegate
    -------------------------------------------------------------------------------
     FUNCTION  "+" ( CONSTANT addend       : IN bit_vector;
		     CONSTANT augend       : IN Integer
		   ) RETURN bit_vector IS
       VARIABLE result    : bit_vector (addend'LENGTH - 1  DOWNTO 0);
       VARIABLE aug_cpy   : bit_vector (addend'LENGTH - 1  DOWNTO 0);
     BEGIN
     -- Convert augend from Integer to bit_vector
	aug_cpy := To_BitVector(augend, addend'LENGTH, DefaultRegMode);
     -- Use the RegAdd_Syn procedure with  DefaultRegMode 
	RegAdd_Syn (result, addend, aug_cpy, DefaultRegMode);
	RETURN result;
     END;
     ---------------------------------------------------------------------------------
     --     Function Name : Overloaded "+" operator
     -- 1.3.8
     --     Purpose       : Addition operator for bit vectors.
     --
     --     Parameters    :     result         left       right
     --                        bit_vector    Integer   bit_vector 
     --
     --     NOTE          : The addition operation is performed assuming all
     --                     operands and results are signed Two's complement integers.
     --
     --                     The addend is converted to bit_vector of length
     --                     equal to the augend. The length of 
     --                     the result equals the length of the augend
     --
     --                     Any overflow condition is ignored.
     --
     --     Use           :
     --                      VARIABLE a: Integer; 
     --                      VARIABLE b,c : bit_vector ( 7 downto 0 );
     --                      c := a + b;
     --                      c := 5 + b; 
     --
     --     See Also      : RegAdd, RegSub, RegInc, RegDec, RegNegate
    -------------------------------------------------------------------------------
     FUNCTION  "+" ( CONSTANT addend       : IN Integer;
		     CONSTANT augend       : IN bit_vector
		   ) RETURN bit_vector IS
       VARIABLE result : bit_vector (augend'LENGTH - 1  DOWNTO 0);
       VARIABLE a_copy : bit_vector (augend'LENGTH - 1  DOWNTO 0);
     BEGIN
     -- Convert addend from Integer to bit_vector
	a_copy := To_BitVector(addend, augend'LENGTH, DefaultRegMode);
     -- Use the RegAdd_Syn procedure with  DefaultRegMode 
	RegAdd_Syn (result, a_copy, augend, DefaultRegMode );
	RETURN result;
     END;
     -------------------------------------------------------------------------------
     --     Function Name : Overloaded "-" operator
     -- 1.3.11    
     --     Purpose       : Subtraction operator for logic vectors.
     --     
     --     Parameters    :     result         left       right
     --                       std_logic_vector    std_logic_vector  std_logic_vector
     --     
     --     NOTE          : The subtraction operation is performed assuming all
     --                     operands and results are signed Two's complement integers.
     --
     --                     The operands may be of different length. The length of
     --                     the result equals the length of the longer operand.
     --     
     --                     Any underflow condition is ignored.
     --     
     --     Use           : 
     --                      VARIABLE a,b,c : std_logic_vector ( 7 downto 0 );
     --                      c := a - b;
     --                      c := a - B"0101";  -- c = a - 5;
     --                      c := a - B"101";   -- c = a - (-3)
     --     
     --     See Also      : RegAdd, RegSub, RegInc, RegDec, RegNegate
     -------------------------------------------------------------------------------
     FUNCTION  "-" ( CONSTANT minuend      : IN std_logic_vector;
		     CONSTANT subtrahend   : IN std_logic_vector
		   ) RETURN std_logic_vector IS
       CONSTANT reslen     : INTEGER := MAXIMUM (minuend'LENGTH, subtrahend'LENGTH);
       VARIABLE result     : std_logic_vector (reslen - 1 DOWNTO 0); 
     BEGIN
     -- Use the RegSub_Syn procedure with  DefaultRegMode 
	RegSub_Syn ( result, minuend, subtrahend, DefaultRegMode );
	RETURN result;
     END;
     -------------------------------------------------------------------------------
     --     Function Name : Overloaded "-" operator
     -- 1.3.12
     --     Purpose       : Subtraction operator for logic vectors.
     --
     --     Parameters    :     result         left       right
     --                       std_logic_vector    INTEGER  std_logic_vector
     --
     --     NOTE          : The subtraction operation is performed assuming all
     --                     operands and results are signed Two's complement integers.
     --
     --                     The minuend is converted to std_logic_vector of length
     --                     equal to the subtrahend. The length of the result
     --                     equals the length of the subtrahend.
     --
     --                     Any overflow condition is ignored.
     --
     --     Use           :
     --                      VARIABLE a: Integer;
     --                      VARIABLE b,c : std_logic_vector ( 7 downto 0 );
     --                      c := a - b;
     --                      c := 5 - b;
     --
     --     See Also      : RegAdd, RegSub, RegInc, RegDec, RegNegate
     -------------------------------------------------------------------------------
     FUNCTION  "-" ( CONSTANT minuend      : IN Integer;
		     CONSTANT subtrahend   : IN std_logic_vector
		   ) RETURN std_logic_vector IS
       VARIABLE result     : std_logic_vector (subtrahend'LENGTH - 1 DOWNTO 0); 
       VARIABLE a_copy     : std_logic_vector (subtrahend'LENGTH - 1 DOWNTO 0); 
     BEGIN
     -- Convert minuend from Integer to std_logic_vector
	a_copy := To_StdLogicVector(minuend, subtrahend'LENGTH, DefaultRegMode);
     -- Use the RegSub_Syn procedure with DefaultRegMode 
       RegSub_Syn (result, a_copy, subtrahend, DefaultRegMode);
       RETURN result;
     END;
     -------------------------------------------------------------------------------
     --     Function Name : Overloaded "-" operator
     -- 1.3.13
     --     Purpose       : Subtraction operator for logic vectors.
     --
     --     Parameters    :     result         left       right
     --                       std_logic_vector    std_logic_vector  Integer
     --
     --     NOTE          : The subtraction operation is performed assuming all
     --                     operands and results are signed Two's complement integers.
     --
     --                     The subtrahend is converted to std_logic_vector of length
     --                     equal to the minuend. The length of the result
     --                     equals the length of the minuend.
     --
     --                     Any overflow condition is ignored.
     --
     --     Use           :
     --                      VARIABLE a,c : std_logic_vector ( 7 downto 0 );
     --                      VARIABLE b: Integer;
     --                      c := a - b;
     --                      c := a - 5;
     --
     --     See Also      : RegAdd, RegSub_Syn, RegInc, RegDec, RegNegate
     -------------------------------------------------------------------------------
     FUNCTION  "-" ( CONSTANT minuend      : IN std_logic_vector;
		     CONSTANT subtrahend   : IN Integer
		   ) RETURN std_logic_vector IS
       VARIABLE result        : std_logic_vector (minuend'LENGTH - 1 DOWNTO 0); 
       VARIABLE b_copy        : std_logic_vector (minuend'LENGTH - 1 DOWNTO 0); 
     BEGIN
     -- Convert subtrahend from Integer to std_logic_vector
	b_copy := To_StdLogicVector(subtrahend, minuend'LENGTH, DefaultRegMode);
     -- Use the RegSub_Syn procedure with DefaultRegMode 
       RegSub_Syn (result, minuend, b_copy,  DefaultRegMode);
       RETURN result;
     END;
     -------------------------------------------------------------------------------
     --     Function Name : Overloaded "-" operator
     --     
     --     Purpose       : Subtraction operator for ulogic vectors.
     --     
     --     Parameters    :     result         left                right
     --                    std_ulogic_vector  std_ulogic_vector  std_ulogic_vector
     --     
     --     NOTE          : The subtraction operation is performed assuming all
     --                     operands and results are signed Two's complement integers.
     --
     --                     The operands may be of different length. The length of
     --                     the result equals the length of the longer operand.
     --     
     --                     Any underflow condition is ignored.
     --     
     --     Use           : 
     --                      VARIABLE a,b,c : std_ulogic_vector ( 7 downto 0 );
     --                      c := a - b;
     --                      c := a - B"0101";  -- c = a - 5;
     --                      c := a - B"101";   -- c = a - (-3)
     --     
     --     See Also      : RegAdd, RegSub, RegInc, RegDec, RegNegate
     -------------------------------------------------------------------------------
     FUNCTION  "-" ( CONSTANT minuend      : IN std_ulogic_vector;
		     CONSTANT subtrahend   : IN std_ulogic_vector
		   ) RETURN std_ulogic_vector IS
       CONSTANT reslen     : INTEGER := MAXIMUM (minuend'LENGTH, subtrahend'LENGTH);
       VARIABLE result     : std_ulogic_vector (reslen - 1 DOWNTO 0); 
     BEGIN
     -- Use the RegSub_Syn procedure with  DefaultRegMode 
	RegSub_Syn ( result, minuend, subtrahend, DefaultRegMode );
	RETURN result;
     END;
     -------------------------------------------------------------------------------
     --     Function Name : Overloaded "-" operator
     -- 1.3.12
     --     Purpose       : Subtraction operator for ulogic vectors.
     --
     --     Parameters    :     result         left       right
     --                    std_ulogic_vector  INTEGER  std_ulogic_vector
     --
     --     NOTE          : The subtraction operation is performed assuming all
     --                     operands and results are signed Two's complement integers.
     --
     --                     The minuend is converted to std_ulogic_vector of length
     --                     equal to the subtrahend. The length of the result
     --                     equals the length of the subtrahend.
     --
     --                     Any overflow condition is ignored.
     --
     --     Use           :
     --                      VARIABLE a: Integer;
     --                      VARIABLE b,c : std_logic_vector ( 7 downto 0 );
     --                      c := a - b;
     --                      c := 5 - b;
     --
     --     See Also      : RegAdd, RegSub, RegInc, RegDec, RegNegate
     -------------------------------------------------------------------------------
     FUNCTION  "-" ( CONSTANT minuend      : IN Integer;
		     CONSTANT subtrahend   : IN std_ulogic_vector
		   ) RETURN std_ulogic_vector IS
       VARIABLE result      : std_ulogic_vector (subtrahend'LENGTH - 1 DOWNTO 0); 
       VARIABLE a_cpy       : std_ulogic_vector (subtrahend'LENGTH - 1 DOWNTO 0); 
     BEGIN
     -- Convert minuend from Integer to std_ulogic_vector
	a_cpy := To_StdULogicVector(minuend, subtrahend'LENGTH, DefaultRegMode);
     -- Use the RegSub_Syn procedure with DefaultRegMode 
	RegSub_Syn (result, a_cpy, subtrahend, DefaultRegMode);
	RETURN result;
     END;
     -------------------------------------------------------------------------------
     --     Function Name : Overloaded "-" operator
     -- 1.3.13
     --     Purpose       : Subtraction operator for ulogic vectors.
     --
     --     Parameters    :     result         left              right
     --                     std_ulogic_vector std_ulogic_vector  Integer
     --
     --     NOTE          : The subtraction operation is performed assuming all
     --                     operands and results are signed Two's complement integers.
     --
     --                     The subtrahend is converted to std_ulogic_vector of length
     --                     equal to the minuend. The length of the result
     --                     equals the length of the minuend.
     --
     --                     Any overflow condition is ignored.
     --
     --     Use           :
     --                      VARIABLE a,c : std_ulogic_vector ( 7 downto 0 );
     --                      VARIABLE b: Integer;
     --                      c := a - b;
     --                      c := a - 5;
     --
     --     See Also      : RegAdd, RegSub, RegInc, RegDec, RegNegate
     -------------------------------------------------------------------------------
     FUNCTION  "-" ( CONSTANT minuend      : IN std_ulogic_vector;
		     CONSTANT subtrahend   : IN Integer
		   ) RETURN std_ulogic_vector IS
       VARIABLE result        : std_ulogic_vector (minuend'LENGTH - 1 DOWNTO 0); 
       VARIABLE b_cpy        : std_ulogic_vector (minuend'LENGTH - 1 DOWNTO 0); 
     BEGIN
     -- Convert subtrahend from Integer to std_logic_vector
	b_cpy := To_StdULogicVector(subtrahend, minuend'LENGTH, DefaultRegMode);
     -- Use the RegSub_Syn procedure with DefaultRegMode 
       RegSub_Syn (result, minuend, b_cpy, DefaultRegMode);
	 RETURN result;
     END;
     -------------------------------------------------------------------------------
     --     Function Name : Overloaded "-" operator
     -- 1.3.14 
     --     Purpose       : Subtraction operator for bit vectors.
     --
     --     Parameters    :     result         left       right
     --                       bit_vector    bit_vector  bit_vector
     --
     --     NOTE          : The subtraction operation is performed assuming all
     --                     operands and results are signed Two's complement integers.
     --
     --                     The operands may be of different length. The length of
     --                     the result equals the length of the longer operand.
     --
     --                     Any underflow condition is ignored.
     --
     --     Use           :
     --                      VARIABLE a,b,c : bit_vector ( 7 downto 0 );
     --                      c := a - b;
     --                      c := a - B"0101";  -- c = a - 5;
     --                      c := a - B"101";   -- c = a - (-3)
     --
     --     See Also      : RegAdd, RegSub, RegInc, RegDec, RegNegate
     -------------------------------------------------------------------------------
     FUNCTION  "-" ( CONSTANT minuend      : IN bit_vector;
		     CONSTANT subtrahend   : IN bit_vector
		   ) RETURN bit_vector IS
       CONSTANT reslen     : INTEGER := MAXIMUM (minuend'LENGTH, subtrahend'LENGTH);
       VARIABLE result     : bit_vector (reslen - 1  DOWNTO 0);
     BEGIN
     -- Use the RegSub_Syn procedure with DefaultRegMode
	 RegSub_Syn (result, minuend, subtrahend, DefaultRegMode);
	 RETURN result;
     END;
     -------------------------------------------------------------------------------
     --     Function Name : Overloaded "-" operator
     -- 1.3.15
     --     Purpose       : Subtraction operator for logic vectors.
     --
     --     Parameters    :     result         left       right
     --                       bit_vector    bit_vector  Integer
     --
     --     NOTE          : The subtraction operation is performed assuming all
     --                     operands and results are signed Two's complement integers.
     --
     --                     The subtrahend is converted to bit_vector of length
     --                     equal to the minuend. The length of the result
     --                     equals the length of the minuend.
     --
     --                     Any overflow condition is ignored.
     --
     --     Use           :
     --                      VARIABLE a,c : bit_vector ( 7 downto 0 );
     --                      VARIABLE b: Integer;
     --                      c := a - b;
     --                      c := a - 5;
     --
     --     See Also      : RegAdd, RegSub, RegInc, RegDec, RegNegate
     -------------------------------------------------------------------------------
     FUNCTION  "-" ( CONSTANT minuend      : IN bit_vector;
		     CONSTANT subtrahend   : IN Integer
		   ) RETURN bit_vector IS
       VARIABLE result       : bit_vector (minuend'LENGTH - 1  DOWNTO 0);
       VARIABLE b_cpy        : bit_vector (minuend'LENGTH - 1  DOWNTO 0);	
     BEGIN
     -- Convert subtrahend from Integer to bit_vector
	b_cpy := To_BitVector(subtrahend, minuend'LENGTH, DefaultRegMode);
     -- Use the RegSub_Syn procedure with DefaultRegMode
	RegSub_Syn (result, minuend, b_cpy, DefaultRegMode);
	RETURN result;
     END;
     -------------------------------------------------------------------------------
     --     Function Name : Overloaded "-" operator
     -- 1.3.16
     --     Purpose       : Subtraction operator for bit vectors.
     --
     --     Parameters    :     result         left       right
     --                       bit_vector    INTEGER  bit_vector
     --
     --     NOTE          : The subtraction operation is performed assuming all
     --                     operands and results are signed Two's complement integers.
     --
     --                     The minuend is converted to bit_vector of length
     --                     equal to the subtrahend. The length of the result
     --                     equals the length of the subtrahend.
     --
     --                     Any overflow condition is ignored.
     --
     --     Use           :
     --                      VARIABLE a: Integer;
     --                      VARIABLE b,c : bit_vector ( 7 downto 0 );
     --                      c := a - b;
     --                      c := 5 - b;
     --
     --     See Also      : RegAdd, RegSub, RegInc, RegDec, RegNegate
     -------------------------------------------------------------------------------
     FUNCTION  "-" ( CONSTANT minuend      : IN Integer;
		     CONSTANT subtrahend   : IN bit_vector
		   ) RETURN bit_vector IS
       VARIABLE result     : bit_vector (subtrahend'LENGTH - 1  DOWNTO 0);
       VARIABLE a_cpy      : bit_vector (subtrahend'LENGTH - 1  DOWNTO 0);
     BEGIN
     -- Convert minuend from Integer to bit_vector
	a_cpy := To_BitVector(minuend, subtrahend'LENGTH, DefaultRegMode);
     -- Use the RegSub_Syn procedure with  DefaultRegMode notation
	RegSub_Syn (result, a_cpy, subtrahend, DefaultRegMode);
	 RETURN result;
     END;
     -------------------------------------------------------------------------------
     --     Function Name : Overloaded "-" operator
     -- 1.4.5
     --     Purpose       : Unary minus operator for bit vectors.
     --
     --     Parameters    :     result         v 
     --                       bit_vector    bit_vector 
     --
     --     NOTE          : The  minus  operation is performed assuming 
     --                     operand and result are signed Two's complement integers.
     --
     --     Use           :
     --                      VARIABLE a,c : bit_vector ( 7 downto 0 );
     --                      c :=  - a;
     --
     --     See Also      :  RegNegate
     -------------------------------------------------------------------------------
     FUNCTION "-"  (CONSTANT subtrahend   : IN bit_vector
		   ) RETURN bit_vector IS
       VARIABLE reg    : bit_vector (subtrahend'LENGTH - 1  DOWNTO 0);
     BEGIN
        reg := subtrahend;
        IF ((reg(subtrahend'LENGTH - 1) /= '0') AND
                 (No_One(reg(subtrahend'LENGTH - 2 downto 0)))) THEN
            -- synopsys translate_off                 
                  ASSERT false
                  REPORT "Unary '-'   ---  2's comp bit_vector  cannot be converted."
                     & " Returning the same vector."
                  SEVERITY Error;   
           -- synopsys translate_on
                return (reg);
        ELSE
           -- Use the RegNegate procedure with default  DefaultRegMode notation
      	       return( RegNegate (subtrahend,  DefaultRegMode));
        END IF;
     END;
     -------------------------------------------------------------------------------
     --     Function Name : Overloaded "-" operator
     -- 1.4.6
     --     Purpose       : Unary minus operator for logic vectors.
     --
     --     Parameters    :     result              operand 
     --                       std_logic_vector    std_logic_vector 
     --
     --     NOTE          : The  minus  operation is performed assuming 
     --                     operand and result are in signed Two's complement notation.
     --
     --     Use           :
     --                      VARIABLE a,c : std_logic_vector ( 7 downto 0 );
     --                      c :=  - a;
     --
     --     See Also      :  RegNegate
     -------------------------------------------------------------------------------
     FUNCTION "-"  (CONSTANT subtrahend   : IN std_logic_vector
		   ) RETURN std_logic_vector IS
       VARIABLE reg    : std_logic_vector (subtrahend'LENGTH - 1  DOWNTO 0);
     BEGIN
        reg := subtrahend;
        IF ((reg(subtrahend'LENGTH - 1) /= '0') AND
                 (No_One(reg(subtrahend'LENGTH - 2 downto 0)))) THEN
            -- synopsys translate_off                 
                  ASSERT false
                  REPORT "Unary '-'   ---  2's comp bit_vector  cannot be converted."
                     & " Returning the same vector."
                  SEVERITY Error;   
           -- synopsys translate_on
                return (reg);
        ELSE
           -- Use the RegNegate procedure with default  DefaultRegMode notation
      	       return( RegNegate (subtrahend,  DefaultRegMode));
        END IF;
     END;
     -------------------------------------------------------------------------------
     --     Function Name : Overloaded "-" operator
     --
     --     Purpose       : Unary minus operator for ulogic vectors.
     --
     --     Parameters    :     result              operand 
     --                       std_ulogic_vector    std_ulogic_vector 
     --
     --     NOTE          : The  minus  operation is performed assuming 
     --                     operand and result are in signed Two's complement notation.
     --
     --     Use           :
     --                      VARIABLE a,c : std_ulogic_vector ( 7 downto 0 );
     --                      c :=  - a;
     --
     --     See Also      :  RegNegate
     -------------------------------------------------------------------------------
     FUNCTION "-"  (CONSTANT subtrahend   : IN std_ulogic_vector
		   ) RETURN std_ulogic_vector IS
       VARIABLE reg    : std_ulogic_vector (subtrahend'LENGTH - 1  DOWNTO 0);
     BEGIN
        reg := subtrahend;
        IF ((reg(subtrahend'LENGTH - 1) /= '0') AND
                 (No_One(reg(subtrahend'LENGTH - 2 downto 0)))) THEN
            -- synopsys translate_off                 
                  ASSERT false
                  REPORT "Unary '-'   ---  2's comp bit_vector  cannot be converted."
                     & " Returning the same vector."
                  SEVERITY Error;   
           -- synopsys translate_on
                return (reg);
        ELSE
           -- Use the RegNegate procedure with default  DefaultRegMode notation
      	       return( RegNegate (subtrahend,  DefaultRegMode));
        END IF;
     END;
     -------------------------------------------------------------------------------
     --     Function Name : Overloaded "*" operator
     --    
     --     Purpose       : Multiplication operator for logic vectors.
     --     
     --     Parameters    :     result         left       right
     --                       std_logic_vector    std_logic_vector  std_logic_vector
     --     
     --     NOTE          : The multiplication operation is performed assuming all
     --                     operands and results are signed Two's complement integers.
     --
     --                     The operands may be of different length. The length of
     --                     the result equals the length of the longer operand.
     --     
     --                     A temporary result is computed of sufficient length
     --                     to avoid overflow. The high order bits of this temporary
     --                     vector are truncated to form the required length result.
     --                     No indication is given if the magnitude of the computed
     --                     result exceeds the size of the returned result vector.
     --     
     --     Use           : 
     --                      VARIABLE a,b,c : std_logic_vector ( 7 downto 0 );
     --                      c := a * b;
     --                      c := a * B"1101";  -- c = a * (-3)
     --     
     --     See Also      : RegMult, RegDiv
     -------------------------------------------------------------------------------
     FUNCTION  "*" ( CONSTANT multiplicand : IN std_logic_vector;
		     CONSTANT multiplier   : IN std_logic_vector
		   ) RETURN std_logic_vector IS
       CONSTANT reslen   : INTEGER := MAXIMUM (multiplicand'LENGTH, multiplier'LENGTH);
       VARIABLE result   : std_logic_vector ( reslen - 1 DOWNTO 0 );
       VARIABLE overflow : std_ulogic;
     BEGIN
     -- Use the general multiplication procedure
	 RegMult ( result, overflow, multiplicand, multiplier, DefaultRegMode);
	 RETURN result;
     END;
     -------------------------------------------------------------------------------
     --     Function Name : Overloaded "*" operator
     -- 1.5.4
     --     Purpose       : Multiplication operator for logic vectors.
     --
     --     Parameters    :     result           left                right
     --                       std_logic_vector    std_logic_vector  Integer
     --
     --     NOTE          : The multiplication operation is performed assuming all
     --                     operands and results are signed Two's complement integers.
     --
     --                     The multiplier is converted to std_logic_vector of length
     --                     equal to the multiplicand. The length of the result
     --                     equals the length of the multiplicand.

     --
     --                     A temporary result is computed of sufficient length
     --                     to avoid overflow. The high order bits of this temporary
     --                     vector are truncated to form the required length result.
     --                     No indication is given if the magnitude of the computed
     --                     result exceeds the size of the returned result vector.
     --
     --     Use           :
     --                      VARIABLE a,c : std_logic_vector ( 7 downto 0 );
     --                      VARIABLE b: Integer;
     --                      c := a * b;
     --                      c := a * 5; 
     --
     --     See Also      : RegMult, RegDiv
   -------------------------------------------------------------------------------
     FUNCTION  "*" ( CONSTANT multiplicand : IN std_logic_vector;
		     CONSTANT multiplier   : IN Integer
		   ) RETURN std_logic_vector IS
       VARIABLE result        : std_logic_vector ( multiplicand'LENGTH - 1 DOWNTO 0 );
       VARIABLE b_copy        : std_logic_vector ( multiplicand'LENGTH - 1 DOWNTO 0 );
       VARIABLE overflow      : std_ulogic;
     BEGIN
     -- Convert multiplier from Integer to std_logic_vector
	b_copy := To_StdLogicVector(multiplier, multiplicand'LENGTH, DefaultRegMode);
     -- Use the general multiplication procedure
	 RegMult ( result, overflow, multiplicand, b_copy, DefaultRegMode);
	 RETURN result;
     END;
     -------------------------------------------------------------------------------
     --     Function Name : Overloaded "*" operator
     -- 1.5.5
     --     Purpose       : Multiplication operator for logic vectors.
     --
     --     Parameters    :     result           left                right
     --                       std_logic_vector    Integer     std_logic_vector
     --
     --     NOTE          : The multiplication operation is performed assuming all
     --                     operands and results are signed Two's complement integers.
     --
     --                     The multiplicand is converted to std_logic_vector of length
     --                     equal to the multiplier. The length of the result
     --                     equals the length of the multiplier.

     --
     --                     A temporary result is computed of sufficient length
     --                     to avoid overflow. The high order bits of this temporary
     --                     vector are truncated to form the required length result.
     --                     No indication is given if the magnitude of the computed
     --                     result exceeds the size of the returned result vector.
     --
     --     Use           :
     --                      VARIABLE a,c : std_logic_vector ( 7 downto 0 );
     --                      VARIABLE b: Integer;
     --                      c := a * b;
     --                      c := a * 5; 
     --
     --     See Also      : RegMult, RegDiv
     -------------------------------------------------------------------------------
     FUNCTION  "*" ( CONSTANT multiplicand : IN Integer;
		     CONSTANT multiplier   : IN std_logic_vector
		   ) RETURN std_logic_vector IS
       VARIABLE result          : std_logic_vector ( multiplier'LENGTH - 1 DOWNTO 0 );
       VARIABLE a_copy          : std_logic_vector ( multiplier'LENGTH - 1 DOWNTO 0 );
       VARIABLE overflow        : std_ulogic;
     BEGIN
     -- Convert multiplicand from Integer to std_logic_vector
	a_copy := To_StdLogicVector(multiplicand, multiplier'LENGTH, DefaultRegMode);
     -- Use the general multiplication procedure
	RegMult ( result, overflow, a_copy, multiplier, DefaultRegMode);
	RETURN result;
     END;
     -------------------------------------------------------------------------------
     --     Function Name : Overloaded "*" operator
     --    
     --     Purpose       : Multiplication operator for ulogic vectors.
     --     
     --     Parameters    :     result         left       right
     --                    std_ulogic_vector    std_ulogic_vector  std_ulogic_vector
     --     
     --     NOTE          : The multiplication operation is performed assuming all
     --                     operands and results are signed Two's complement integers.
     --
     --                     The operands may be of different length. The length of
     --                     the result equals the length of the longer operand.
     --     
     --                     A temporary result is computed of sufficient length
     --                     to avoid overflow. The high order bits of this temporary
     --                     vector are truncated to form the required length result.
     --                     No indication is given if the magnitude of the computed
     --                     result exceeds the size of the returned result vector.
     --     
     --     Use           : 
     --                      VARIABLE a,b,c : std_ulogic_vector ( 7 downto 0 );
     --                      c := a * b;
     --                      c := a * B"1101";  -- c = a * (-3)
     --     
     --     See Also      : RegMult, RegDiv
     -------------------------------------------------------------------------------
     FUNCTION  "*" ( CONSTANT multiplicand : IN std_ulogic_vector;
		     CONSTANT multiplier   : IN std_ulogic_vector
		   ) RETURN std_ulogic_vector IS
       CONSTANT reslen   : INTEGER := MAXIMUM (multiplicand'LENGTH, multiplier'LENGTH);
       VARIABLE result   : std_ulogic_vector ( reslen - 1 DOWNTO 0 );
       VARIABLE overflow : std_ulogic;
     BEGIN
     -- Use the general multiplication procedure
	 RegMult ( result, overflow, multiplicand, multiplier, DefaultRegMode );
	 RETURN result;
     END;
     -------------------------------------------------------------------------------
     --     Function Name : Overloaded "*" operator
     -- 1.5.4
     --     Purpose       : Multiplication operator for logic vectors.
     --
     --     Parameters    :     result           left                right
     --                     std_ulogic_vector    std_ulogic_vector  Integer
     --
     --     NOTE          : The multiplication operation is performed assuming all
     --                     operands and results are signed Two's complement integers.
     --
     --                     The multiplier is converted to std_ulogic_vector of length
     --                     equal to the multiplicand. The length of the result
     --                     equals the length of the multiplicand.

     --
     --                     A temporary result is computed of sufficient length
     --                     to avoid overflow. The high order bits of this temporary
     --                     vector are truncated to form the required length result.
     --                     No indication is given if the magnitude of the computed
     --                     result exceeds the size of the returned result vector.
     --
     --     Use           :
     --                      VARIABLE a,c : std_ulogic_vector ( 7 downto 0 );
     --                      VARIABLE b: Integer;
     --                      c := a * b;
     --                      c := a * 5; 
     --
     --     See Also      : RegMult, RegDiv
   -------------------------------------------------------------------------------
     FUNCTION  "*" ( CONSTANT multiplicand : IN std_ulogic_vector;
		     CONSTANT multiplier   : IN Integer
		   ) RETURN std_ulogic_vector IS
       VARIABLE result        : std_ulogic_vector ( multiplicand'LENGTH - 1 DOWNTO 0 );
       VARIABLE b_cpy         : std_ulogic_vector ( multiplicand'LENGTH - 1 DOWNTO 0 );
       VARIABLE overflow      : std_ulogic;
     BEGIN
     -- Convert multiplier from Integer to std_ulogic_vector
	b_cpy := To_StdULogicVector(multiplier, multiplicand'LENGTH, DefaultRegMode);
     -- Use the general multiplication procedure
	 RegMult ( result, overflow, multiplicand, b_cpy , DefaultRegMode);
	 RETURN result;
     END;
     -------------------------------------------------------------------------------
     --     Function Name : Overloaded "*" operator
     -- 1.5.5
     --     Purpose       : Multiplication operator for logic vectors.
     --
     --     Parameters    :     result           left                right
     --                       std_ulogic_vector    Integer     std_ulogic_vector
     --
     --     NOTE          : The multiplication operation is performed assuming all
     --                     operands and results are signed Two's complement integers.
     --
     --                     The multiplicand is converted to std_ulogic_vector of length
     --                     equal to the multiplier. The length of the result
     --                     equals the length of the multiplier.

     --
     --                     A temporary result is computed of sufficient length
     --                     to avoid overflow. The high order bits of this temporary
     --                     vector are truncated to form the required length result.
     --                     No indication is given if the magnitude of the computed
     --                     result exceeds the size of the returned result vector.
     --
     --     Use           :
     --                      VARIABLE a,c : std_ulogic_vector ( 7 downto 0 );
     --                      VARIABLE b: Integer;
     --                      c := a * b;
     --                      c := a * 5; 
     --
     --     See Also      : RegMult, RegDiv
     -------------------------------------------------------------------------------
     FUNCTION  "*" ( CONSTANT multiplicand : IN Integer;
		     CONSTANT multiplier   : IN std_ulogic_vector
		   ) RETURN std_ulogic_vector IS
       VARIABLE result          : std_ulogic_vector ( multiplier'LENGTH - 1 DOWNTO 0 );
       VARIABLE a_cpy          : std_ulogic_vector ( multiplier'LENGTH - 1 DOWNTO 0 );
       VARIABLE overflow        : std_ulogic;
     BEGIN
     -- Convert multiplicand from Integer to std_ulogic_vector
	a_cpy := To_StdULogicVector(multiplicand, multiplier'LENGTH, DefaultRegMode);
     -- Use the general multiplication procedure
	 RegMult ( result, overflow, a_cpy, multiplier, DefaultRegMode);
	 RETURN result;
     END;
 --+-----------------------------------------------------------------------------
 --|     Function Name : Overloaded "*" operator
 --|
 --|     Purpose       : Multiplication operator for bit vectors.
 --|
 --|     Parameters    :     result         left       right
 --|                       BIT_VECTOR    BIT_VECTOR  BIT_VECTOR
 --|
 --|     NOTE          : The multiplication operation is performed assuming all
 --|                     operands and results are signed Two's complement integers.
 --|
 --|                     The operands may be of different length. The length of
 --|                     the result equals the length of the longer operand.
 --|
 --|                     A temporary result is computed of sufficient length
 --|                     to avoid overflow. The high order bits of this temporary
 --|                     vector are truncated to form the required length result.
 --|                     No indication is given if the magnitude of the computed
 --|                     result exceeds the size of the returned result vector.
 --|
 --|     Use           :
 --|                      VARIABLE a,b,c : bit_vector ( 7 downto 0 );
 --|                      c := a * b;
 --|                      c := a * B"1101";  -- c = a * (-3)
 --|
 --|     See Also      : RegMult, RegDiv
 --|-----------------------------------------------------------------------------
     FUNCTION  "*" ( CONSTANT multiplicand : IN BIT_VECTOR;
		     CONSTANT multiplier   : IN BIT_VECTOR
		   ) RETURN BIT_VECTOR IS
       CONSTANT reslen   : INTEGER := MAXIMUM (multiplicand'LENGTH, multiplier'LENGTH);
       VARIABLE result   : BIT_VECTOR ( reslen - 1 DOWNTO 0 );
       VARIABLE overflow : BIT;
     BEGIN
     -- Use the general multiplication procedure
	 RegMult ( result, overflow, multiplicand, multiplier, DefaultRegMode);
	 RETURN result;
     END;
 --+-----------------------------------------------------------------------------
 --|     Function Name : Overloaded "*" operator
 --| 1.5.7
 --|     Purpose       : Multiplication operator for bit vectors.
 --|
 --|     Parameters    :     result         left       right
 --|                       BIT_VECTOR    BIT_VECTOR  INTEGER
 --|
 --|     NOTE          : The multiplication operation is performed assuming all
 --|                     operands and results are signed Two's complement integers.
 --|
 --|                     The multiplier is converted to bit_vector of length
 --|                     equal to the multiplicand. The length of the result
 --|                     equals the length of the multiplicand.
 --|
 --|                     A temporary result is computed of sufficient length
 --|                     to avoid overflow. The high order bits of this temporary
 --|                     vector are truncated to form the required length result.
 --|                     No indication is given if the magnitude of the computed
 --|                     result exceeds the size of the returned result vector.
 --|
 --|     Use           :
 --|                      VARIABLE a,c : BIT_VECTOR ( 7 downto 0 );
 --|                      VARIABLE b: INTEGER;
 --|                      c := a * b;
 --|                      c := a * 5; 
 --|
 --|     See Also      : RegMult, RegDiv
 --|-----------------------------------------------------------------------------
     FUNCTION  "*" ( CONSTANT multiplicand : IN BIT_VECTOR;
		     CONSTANT multiplier   : IN INTEGER
		   ) RETURN BIT_VECTOR IS
       VARIABLE result       : BIT_VECTOR ( multiplicand'LENGTH - 1 DOWNTO 0 );
       VARIABLE b_copy       : BIT_VECTOR ( multiplicand'LENGTH - 1 DOWNTO 0 );
       VARIABLE overflow     : BIT;
     BEGIN
     -- Convert multiplier from Integer to BIT_VECTOR and
	b_copy := To_BitVector(multiplier, multiplicand'LENGTH, DefaultRegMode);
     --  Use the general multiplication procedure
	 RegMult ( result, overflow, multiplicand, b_copy, DefaultRegMode );
	 RETURN result;
     END;
 --+-----------------------------------------------------------------------------
 --|     Function Name : Overloaded "*" operator
 --| 1.5.8
 --|     Purpose       : Multiplication operator for bit vectors.
 --|
 --|     Parameters    :     result         left       right
 --|                       BIT_VECTOR    INTEGER  BIT_VECTOR
 --|
 --|     NOTE          : The multiplication operation is performed assuming all
 --|                     operands and results are signed Two's complement integers.
 --|
 --|                     The multiplicand is converted to BIT_VECTOR of length
 --|                     equal to the multiplier. The length of the result
 --|                     equals the length of the multiplier.
 --|
 --|                     A temporary result is computed of sufficient length
 --|                     to avoid overflow. The high order bits of this temporary
 --|                     vector are truncated to form the required length result.
 --|                     No indication is given if the magnitude of the computed
 --|                     result exceeds the size of the returned result vector.
 --|
 --|     Use           :
 --|                      VARIABLE a : INTEGER;
 --|                      VARIABLE b,c : BIT_VECTOR ( 7 downto 0 );
 --|                      c := a * b;
 --|                      c := 5 * b; 
 --|
 --|     See Also      : RegMult, RegDiv
 --|-----------------------------------------------------------------------------
    FUNCTION  "*" ( CONSTANT multiplicand : IN INTEGER; 
		    CONSTANT multiplier   : IN BIT_VECTOR
		   ) RETURN BIT_VECTOR IS
       VARIABLE result         : BIT_VECTOR ( multiplier'LENGTH - 1 DOWNTO 0 );
       VARIABLE a_copy         : BIT_VECTOR ( multiplier'LENGTH - 1 DOWNTO 0 );
       VARIABLE overflow       : BIT;
     BEGIN
     -- Convert multiplicand from Integer to BIT_VECTOR
	a_copy := To_BitVector(multiplicand, multiplier'LENGTH, DefaultRegMode);
     -- Use the general multiplication procedure
	 RegMult ( result, overflow, a_copy, multiplier, DefaultRegMode );
	 RETURN result;
     END;
     -------------------------------------------------------------------------------
     --     Function Name : Overloaded "/" operator
     --    
     --     Purpose       : Division operator for logic vectors.
     --     
     --     Parameters    :     result         left       right
     --                       std_logic_vector    std_logic_vector  std_logic_vector
     --     
     --     NOTE          : The division operation is performed assuming all
     --                     operands and results are signed Two's complement integers.
     --
     --                     The operands may be of different length. The length of
     --                     the result equals the length of dividend.
     --     
     --                     Any remainder is ignored - no rounding is applied.
     --
     --                     An ASSERTION message of severity ERROR is issued
     --                     if division by 0 is attempted. In this case the
     --                     return value is 0 (all 0's).
     --     
     --     Use           : 
     --                      VARIABLE a,b,c : std_logic_vector ( 7 downto 0 );
     --                      c := a / b;
     --                      c := a / B"1101";  -- c = a / (-3)
     --     Se Also       : RegMult, RegDiv
     ----------------------------------------------------------------------------------
     FUNCTION  "/" ( CONSTANT dividend     : IN std_logic_vector;
		     CONSTANT divisor      : IN std_logic_vector
		   ) RETURN std_logic_vector IS
       VARIABLE result    : std_logic_vector ( dividend'LENGTH - 1 DOWNTO 0 );
       VARIABLE remainder : std_logic_vector(dividend'LENGTH - 1 DOWNTO 0);
       VARIABLE zflag     : std_ulogic;
     BEGIN
     -- Use the general division procedure 
	 RegDiv ( result, remainder, zflag, dividend, divisor, DefaultRegMode); 
	 RETURN result; 
     END;
     -------------------------------------------------------------------------------
     --     Function Name : Overloaded "/" operator
     -- 1.5.12
     --     Purpose       : Division operator for logic vectors.
     --
     --     Parameters    :     result         left       right
     --                       std_logic_vector    std_logic_vector  INTEGER
     --
     --     NOTE          : The division operation is performed assuming all
     --                     operands and results are signed Two's complement integers.
     --
     --                     The divisor is converted to std_logic_vector of length
     --                     equal to the dividend. The length of the result
     --                     equals the length of the dividend.
     --
     --                     Any remainder is ignored - no rounding is applied.
     --
     --                     An ASSERTION message of severity ERROR is issued
     --                     if division by 0 is attempted. In this case the
     --                     return value is 0 (all 0's).
     --
     --     Use           :
     --                      VARIABLE a,c : std_logic_vector ( 7 downto 0 );
     --                      VARIABLE b : INTEGER;
     --                      c := a / b;
     --                      c := a / 5; 
     --     Se Also       : RegMult, RegDiv
     --------------------------------------------------------------------------------
     FUNCTION  "/" ( CONSTANT dividend     : IN std_logic_vector;
		     CONSTANT divisor      : IN INTEGER
		   ) RETURN std_logic_vector IS
       VARIABLE result     : std_logic_vector ( dividend'LENGTH - 1 DOWNTO 0 );
       VARIABLE remainder  : std_logic_vector (dividend'LENGTH - 1 DOWNTO 0);
       VARIABLE bv         : std_logic_vector (dividend'LENGTH - 1 DOWNTO 0);
       VARIABLE zflag      : std_ulogic;
     BEGIN
     -- Convert divisor from Integer to std_logic_vector
	bv := To_StdLogicVector(divisor, dividend'LENGTH, DefaultRegMode);
     -- Use the general division procedure
	 RegDiv ( result, remainder, zflag, dividend, bv,  DefaultRegMode );
	 RETURN result;
     END;
     -------------------------------------------------------------------------------
     --     Function Name : Overloaded "/" operator
     -- 1.5.13
     --     Purpose       : Division operator for logic vectors.
     --
     --     Parameters    :     result         left       right
     --                       std_logic_vector    INTEGER  std_logic_vector
     --
     --     NOTE          : The division operation is performed assuming all
     --                     operands and results are signed Two's complement integers.
     --
     --                     The dividend is converted to std_logic_vector of length
     --                     equal to the divisor. The length of the result
     --                     equals the length of the divisor.
     --
     --                     Any remainder is ignored - no rounding is applied.
     --
     --                     An ASSERTION message of severity ERROR is issued
     --                     if division by 0 is attempted. In this case the
     --                     return value is 0 (all 0's).
     --
     --     Use           :
     --                      VARIABLE a : INTEGER;
     --                      VARIABLE b,c : std_logic_vector ( 7 downto 0 );
     --                      c := a / b;
     --                      c := 5 / b;
     --     Se Also       : RegMult, RegDiv
     --------------------------------------------------------------------------------
     FUNCTION  "/" ( CONSTANT dividend     : IN INTEGER;
		     CONSTANT divisor      : IN std_logic_vector
		   ) RETURN std_logic_vector IS
       VARIABLE result      : std_logic_vector ( divisor'LENGTH - 1 DOWNTO 0 );
       VARIABLE remainder   : std_logic_vector (divisor'LENGTH - 1 DOWNTO 0);
       VARIABLE av          : std_logic_vector (divisor'LENGTH - 1 DOWNTO 0);
       VARIABLE zflag       : std_ulogic;
     BEGIN
     -- Convert dividend from Integer to std_logic_vector
      av := To_StdLogicVector(dividend, divisor'LENGTH, DefaultRegMode);
     -- Use the general division procedure
	 RegDiv ( result, remainder,zflag, av, divisor, DefaultRegMode );
	 RETURN result;
     END;
     -------------------------------------------------------------------------------
     --     Function Name : Overloaded "/" operator
     --    
     --     Purpose       : Division operator for ulogic vectors.
     --     
     --     Parameters    :     result         left       right
     --                       std_ulogic_vector    std_ulogic_vector  std_ulogic_vector
     --     
     --     NOTE          : The division operation is performed assuming all
     --                     operands and results are signed Two's complement integers.
     --
     --                     The operands may be of different length. The length of
     --                     the result equals the length of the dividend.
     --     
     --                     Any remainder is ignored - no rounding is applied.
     --
     --                     An ASSERTION message of severity ERROR is issued
     --                     if division by 0 is attempted. In this case the
     --                     return value is 0 (all 0's).
     --     
     --     Use           : 
     --                      VARIABLE a,b,c : std_ulogic_vector ( 7 downto 0 );
     --                      c := a / b;
     --                      c := a / B"1101";  -- c = a / (-3)
     --     Se Also       : RegMult, RegDiv
     ---------------------------------------------------------------------------------
     FUNCTION  "/" ( CONSTANT dividend     : IN std_ulogic_vector;
		     CONSTANT divisor      : IN std_ulogic_vector
		   ) RETURN std_ulogic_vector IS
       VARIABLE result    : std_ulogic_vector ( dividend'length - 1 DOWNTO 0 );
       VARIABLE remainder : std_ulogic_vector(dividend'length - 1 DOWNTO 0);
       VARIABLE zflag     : std_ulogic;
     BEGIN
     -- Use the general division procedure 
	 RegDiv ( result, remainder, zflag, dividend, divisor, DefaultRegMode); 
	 RETURN result; 
     END;
     -------------------------------------------------------------------------------
     --     Function Name : Overloaded "/" operator
     -- 1.5.12
     --     Purpose       : Division operator for logic vectors.
     --
     --     Parameters    :     result         left       right
     --                       std_ulogic_vector    std_ulogic_vector  INTEGER
     --
     --     NOTE          : The division operation is performed assuming all
     --                     operands and results are signed Two's complement integers.
     --
     --                     The divisor is converted to std_ulogic_vector of length
     --                     equal to the dividend. The length of the result
     --                     equals the length of the dividend.
     --
     --                     Any remainder is ignored - no rounding is applied.
     --
     --                     An ASSERTION message of severity ERROR is issued
     --                     if division by 0 is attempted. In this case the
     --                     return value is 0 (all 0's).
     --
     --     Use           :
     --                      VARIABLE a,c : std_ulogic_vector ( 7 downto 0 );
     --                      VARIABLE b : INTEGER;
     --                      c := a / b;
     --                      c := a / 5; 
     --     Se Also       : RegMult, RegDiv
   --------------------------------------------------------------------------------
     FUNCTION  "/" ( CONSTANT dividend     : IN std_ulogic_vector;
		     CONSTANT divisor      : IN INTEGER
		   ) RETURN std_ulogic_vector IS
       VARIABLE result     : std_ulogic_vector ( dividend'LENGTH - 1 DOWNTO 0 );
       VARIABLE remainder  : std_ulogic_vector (dividend'LENGTH - 1 DOWNTO 0);
       VARIABLE bv         : std_ulogic_vector (dividend'LENGTH - 1 DOWNTO 0);
       VARIABLE zflag      : std_ulogic;
     BEGIN
     -- Convert divisor from Integer to std_ulogic_vector
	bv := To_StdULogicVector(divisor, dividend'LENGTH, DefaultRegMode);
     -- Use the general division procedure
	 RegDiv ( result, remainder, zflag,dividend, bv, DefaultRegMode );
	 RETURN result;
     END;
     -------------------------------------------------------------------------------
     --     Function Name : Overloaded "/" operator
     -- 1.5.13
     --     Purpose       : Division operator for logic vectors.
     --
     --     Parameters    :     result         left       right
     --                       std_ulogic_vector    INTEGER  std_ulogic_vector
     --
     --     NOTE          : The division operation is performed assuming all
     --                     operands and results are signed Two's complement integers.
     --
     --                     The dividend is converted to std_ulogic_vector of length
     --                     equal to the divisor. The length of the result
     --                     equals the length of the divisor.
     --
     --                     Any remainder is ignored - no rounding is applied.
     --
     --                     An ASSERTION message of severity ERROR is issued
     --                     if division by 0 is attempted. In this case the
     --                     return value is 0 (all 0's).
     --
     --     Use           :
     --                      VARIABLE a : INTEGER;
     --                      VARIABLE b,c : std_ulogic_vector ( 7 downto 0 );
     --                      c := a / b;
     --                      c := 5 / b;
     --     Se Also       : RegMult, RegDiv
     --------------------------------------------------------------------------------
     FUNCTION  "/" ( CONSTANT dividend     : IN INTEGER;
		     CONSTANT divisor      : IN std_ulogic_vector
		   ) RETURN std_ulogic_vector IS
       VARIABLE result      : std_ulogic_vector ( divisor'LENGTH - 1 DOWNTO 0 );
       VARIABLE remainder   : std_ulogic_vector(divisor'LENGTH - 1 DOWNTO 0);
       VARIABLE av          : std_ulogic_vector(divisor'LENGTH - 1 DOWNTO 0);
       VARIABLE zflag       : std_ulogic;
     BEGIN
     -- Convert dividend from Integer to std_ulogic_vector
	av := To_StdULogicVector(dividend, divisor'LENGTH, DefaultRegMode);
     -- Use the general division procedure
	 RegDiv ( result, remainder, zflag, av, divisor, DefaultRegMode );
	 RETURN result;
     END;
 --+-----------------------------------------------------------------------------
 --|     Function Name : Overloaded "/" operator
 --| 1.5.14
 --|     Purpose       : Division operator for bit vectors.  
 --|     Parameters    :     result         left       right
 --|                       BIT_VECTOR    BIT_VECTOR  BIT_VECTOR
 --|
 --|     NOTE          : The division operation is performed assuming all
 --|                     operands and results are signed Two's complement integers.
 --|
 --|                     The operands may be of different length. The length of
 --|                     the result equals the length of the dividend.
 --|
 --|                     Any remainder is ignored - no rounding is applied.
 --|
 --|                     An ASSERTION message of severity ERROR is issued
 --|                     if division by 0 is attempted. In this case the
 --|                     return value is 0 (all 0's).
 --|
 --|     Use           :
 --|                      VARIABLE a,b,c : bit_vector ( 7 downto 0 );
 --|                      c := a / b;
 --|                      c := a / B"1101";  -- c = a / (-3)
 --|
 --|     See Also      : RegMult, RegDiv
 --|-----------------------------------------------------------------------------
     FUNCTION  "/" ( CONSTANT dividend     : IN BIT_VECTOR;
		     CONSTANT divisor      : IN BIT_VECTOR
		   ) RETURN BIT_VECTOR IS
       VARIABLE result    : BIT_VECTOR ( dividend'LENGTH - 1 DOWNTO 0 );
       VARIABLE remainder : BIT_VECTOR(dividend'LENGTH - 1 DOWNTO 0);
       VARIABLE zflag     : BIT;
     BEGIN
     -- Use the general division procedure
	 RegDiv ( result, remainder, zflag, dividend, divisor, DefaultRegMode );
	 RETURN result;
     END;
 --+-----------------------------------------------------------------------------
 --|     Function Name : Overloaded "/" operator
 --| 1.5.15
 --|     Purpose       : Division operator for bit vectors.
 --|     Parameters    :     result         left       right
 --|                       BIT_VECTOR    BIT_VECTOR  INTEGER
 --|
 --|     NOTE          : The division operation is performed assuming all
 --|                     operands and results are signed Two's complement integers.
 --|
 --|                     The divisor is converted to bit_vector of length
 --|                     equal to the dividend. The length of the result
 --|                     equals the length of the dividend.
 --|
 --|                     Any remainder is ignored - no rounding is applied.
 --|
 --|                     An ASSERTION message of severity ERROR is issued
 --|                     if division by 0 is attempted. In this case the
 --|                     return value is 0 (all 0's).
 --|
 --|     Use           :
 --|                      VARIABLE a,c : BIT_VECTOR ( 7 downto 0 );
 --|                      VARIABLE b : INTEGER;
 --|                      c := a / b;
 --|                      c := a / 5;
 --| 
 --|     See Also      : RegMult, RegDiv
 --|-----------------------------------------------------------------------------
     FUNCTION  "/" ( CONSTANT dividend     : IN BIT_VECTOR;
		     CONSTANT divisor      : IN INTEGER
		   ) RETURN BIT_VECTOR IS
       VARIABLE result    : BIT_VECTOR ( dividend'LENGTH - 1 DOWNTO 0 );
       VARIABLE remainder : BIT_VECTOR (dividend'LENGTH - 1 DOWNTO 0);
       VARIABLE bv        : BIT_VECTOR (dividend'LENGTH - 1 DOWNTO 0);
       VARIABLE zflag     : BIT;
     BEGIN
     -- Convert divisor from Integer to bit_vector
	bv := To_BitVector(divisor, dividend'LENGTH, DefaultRegMode);
     -- Use the general division procedure
	 RegDiv ( result, remainder, zflag,dividend, bv, DefaultRegMode );
	 RETURN result;
     END;
 --+-----------------------------------------------------------------------------
 --|     Function Name : Overloaded "/" operator
 --| 1.5.16
 --|     Purpose       : Division operator for bit vectors.
 --|     Parameters    :     result         left       right
 --|                       BIT_VECTOR    INTEGER  BIT_VECTOR
 --|
 --|     NOTE          : The division operation is performed assuming all
 --|                     operands and results are signed Two's complement integers.
 --|
 --|                     The dividend is converted to bit_vector of length
 --|                     equal to the divisor. The length of the result
 --|                     equals the length of the divisor.
 --|
 --|                     Any remainder is ignored - no rounding is applied.
 --|
 --|                     An ASSERTION message of severity ERROR is issued
 --|                     if division by 0 is attempted. In this case the
 --|                     return value is 0 (all 0's).
 --|
 --|
 --|     Use           :
 --|                      VARIABLE a : INTEGER;
 --|                      VARIABLE b,c : BIT_VECTOR ( 7 downto 0 );
 --|                      c := a / b;
 --|                      c := 5 / b;
 --|
 --|     See Also      : RegMult, RegDiv
 --|-----------------------------------------------------------------------------
     FUNCTION  "/" ( CONSTANT dividend     : IN INTEGER;
		     CONSTANT divisor      : IN BIT_VECTOR
		   ) RETURN BIT_VECTOR IS
       VARIABLE result     : BIT_VECTOR(divisor'LENGTH - 1 DOWNTO 0);
       VARIABLE remainder  : BIT_VECTOR(divisor'LENGTH - 1 DOWNTO 0);
       VARIABLE av         : BIT_VECTOR(divisor'LENGTH - 1 DOWNTO 0);
       VARIABLE zflag      : BIT;
     BEGIN
     -- Convert dividend from Integer to bit_vector
	av := To_BitVector(dividend, divisor'LENGTH, DefaultRegMode);
     -- Use the general divison procedure
	 RegDiv ( result, remainder, zflag, av, divisor, DefaultRegMode );
	 RETURN result;
     END;
     -------------------------------------------------------------------------------
     --     Function Name : Overloaded "mod" operator
     -- 1.5.19
     --     Purpose       : Modulus operator for logic vectors.
     --
     --     Parameters    :     result         left       right
     --                       std_logic_vector    std_logic_vector  std_logic_vector
     --
     --     NOTE          : The modulus operation is performed assuming all
     --                     operands and results are signed Two's complement integers.
     --
     --                     The operands may be of different length. The length of
     --                     the result equals the length of the modulus.
     --
     --                     An ASSERTION message of severity ERROR is issued
     --                     if division by 0 is attempted. In this case the
     --                     return value is 0 (all 0's).
     --
     --     Use           :
     --                      VARIABLE a,b,c : std_logic_vector ( 7 downto 0 );
     --                      c := a mod b;
     --                      c := a mod B"1101";  -- c = a / (-3)
     --     Se Also       : RegRem, RegDiv
     -------------------------------------------------------------------------------
     FUNCTION  "mod" ( CONSTANT dividend     : IN std_logic_vector;
		       CONSTANT modulus      : IN std_logic_vector
		     ) RETURN std_logic_vector IS
       VARIABLE result   : std_logic_vector ( modulus'LENGTH - 1 DOWNTO 0 );
       VARIABLE zflag    : std_ulogic;
     BEGIN
     -- Use the general modulus procedure
	 RegMod ( result, zflag, dividend, modulus, DefaultRegMode);
	 RETURN result;
     END;
   -------------------------------------------------------------------------------
     --     Function Name : Overloaded "mod" operator
     -- 1.5.20
     --     Purpose       : Modulus operator for logic vectors.
     --
     --     Parameters    :     result         left       right
     --                       std_logic_vector    std_logic_vector  INTEGER
     --
     --     NOTE          : The modulus operation is performed assuming all
     --                     operands and results are signed Two's complement integers.
     --
     --                     The modulus is converted to std_logic_vector of length
     --                     equal to the dividend. The length of the result
     --                     equals the length of the dividend.
     --
     --                     An ASSERTION message of severity ERROR is issued
     --                     if division by 0 is attempted. In this case the
     --                     return value is 0 (all 0's).
     --
     --     Use           :
     --                      VARIABLE a,c : std_logic_vector ( 7 downto 0 );
     --                      VARIABLE b : INTEGER;
     --                      c := a mod b;
     --                      c := a mod 5;
     --     Se Also       : RegRem, RegDiv
   --------------------------------------------------------------------------------
     FUNCTION  "mod" ( CONSTANT dividend     : IN std_logic_vector;
		       CONSTANT modulus      : IN INTEGER
		     ) RETURN std_logic_vector IS
       VARIABLE result     : std_logic_vector ( dividend'LENGTH - 1 DOWNTO 0 );
       VARIABLE bv     : std_logic_vector ( dividend'LENGTH - 1 DOWNTO 0 );
       VARIABLE zflag      : std_ulogic;
     BEGIN
     -- Convert modulus from Integer to std_logic_vector
	bv := To_StdLogicVector(modulus, dividend'LENGTH, DefaultRegMode);
     -- Use the general modulus procedure
	 RegMod ( result, zflag, dividend, bv, DefaultRegMode );
	 RETURN result;
     END;
     -------------------------------------------------------------------------------
     --     Function Name : Overloaded "mod" operator
     -- 1.5.21
     --     Purpose       : Modulus operator for logic vectors.
     --
     --     Parameters    :     result         left       right
     --                       std_logic_vector    INTEGER  std_logic_vector
     --
     --     NOTE          : The modulus operation is performed assuming all
     --                     operands and results are signed Two's complement integers.
     --
     --                     The dividend is converted to std_logic_vector of length
     --                     equal to the modulus. The length of the result
     --                     equals the length of the modulus.
     --
     --                     An ASSERTION message of severity ERROR is issued
     --                     if division by 0 is attempted. In this case the
     --                     return value is 0 (all 0's).
     --
     --     Use           :
     --                      VARIABLE a : INTEGER;
     --                      VARIABLE b,c : std_logic_vector ( 7 downto 0 );
     --                      c := a mod b;
     --                      c := 5 mod b;
     --     Se Also       : RegRem, RegDiv
     --------------------------------------------------------------------------------
     FUNCTION  "mod" ( CONSTANT dividend     : IN INTEGER;
		       CONSTANT modulus      : IN std_logic_vector
		     ) RETURN std_logic_vector IS
       VARIABLE result      : std_logic_vector ( modulus'LENGTH - 1 DOWNTO 0 );
       VARIABLE av          : std_logic_vector ( modulus'LENGTH - 1 DOWNTO 0 );
       VARIABLE zflag       : std_ulogic;
     BEGIN
     -- Convert dividend from Integer to std_logic_vector
	av := To_StdLogicVector(dividend, modulus'LENGTH, DefaultRegMode);
     -- Use the general modulus procedure
	 RegMod ( result, zflag, av, modulus, DefaultRegMode );
	 RETURN result;
     END;
     -------------------------------------------------------------------------------
     --     Function Name : Overloaded "mod" operator
     -- 
     --     Purpose       : Modulus operator for ulogic vectors.
     --
     --     Parameters    :     result         left       right
     --                       std_ulogic_vector    std_ulogic_vector  std_ulogic_vector
     --
     --     NOTE          : The modulus operation is performed assuming all
     --                     operands and results are signed Two's complement integers.
     --
     --                     The operands may be of different length. The length of
     --                     the result equals the length of the modulus.
     --
     --                     An ASSERTION message of severity ERROR is issued
     --                     if division by 0 is attempted. In this case the
     --                     return value is 0 (all 0's).
     --
     --     Use           :
     --                      VARIABLE a,b,c : std_ulogic_vector ( 7 downto 0 );
     --                      c := a mod b;
     --                      c := a mod B"1101";  -- c = a / (-3)
     --     Se Also       : RegRem, RegDiv
     --------------------------------------------------------------------------------
     FUNCTION  "mod" ( CONSTANT dividend     : IN std_ulogic_vector;
		       CONSTANT modulus      : IN std_ulogic_vector
		     ) RETURN std_ulogic_vector IS
       VARIABLE result   : std_ulogic_vector ( modulus'LENGTH - 1 DOWNTO 0 );
       VARIABLE zflag    : std_ulogic;
     BEGIN
     -- Use the general modulus procedure
	 RegMod ( result, zflag, dividend, modulus, DefaultRegMode );
	 RETURN result;
     END;
   -------------------------------------------------------------------------------
     --     Function Name : Overloaded "mod" operator
     -- 
     --     Purpose       : Modulus operator for ulogic vectors.
     --
     --     Parameters    :     result         left       right
     --                       std_ulogic_vector    std_ulogic_vector  INTEGER
     --
     --     NOTE          : The modulus operation is performed assuming all
     --                     operands and results are signed Two's complement integers.
     --
     --                     The modulus is converted to std_ulogic_vector of length
     --                     equal to the dividend. The length of the result
     --                     equals the length of the dividend.
     --
     --                     An ASSERTION message of severity ERROR is issued
     --                     if division by 0 is attempted. In this case the
     --                     return value is 0 (all 0's).
     --
     --     Use           :
     --                      VARIABLE a,c : std_ulogic_vector ( 7 downto 0 );
     --                      VARIABLE b : INTEGER;
     --                      c := a mod b;
     --                      c := a mod 5;
     --     Se Also       : RegRem, RegDiv
   --------------------------------------------------------------------------------
     FUNCTION  "mod" ( CONSTANT dividend     : IN std_ulogic_vector;
		       CONSTANT modulus      : IN INTEGER
		     ) RETURN std_ulogic_vector IS
       VARIABLE result     : std_ulogic_vector ( dividend'LENGTH - 1 DOWNTO 0 );
       VARIABLE bu         : std_ulogic_vector ( dividend'LENGTH - 1 DOWNTO 0 );
       VARIABLE zflag      : std_ulogic;
     BEGIN
     -- Convert modulus from Integer to std_ulogic_vector
	bu := To_StdULogicVector(modulus, dividend'LENGTH, DefaultRegMode);
     -- Use the general modulus procedure
	 RegMod ( result, zflag, dividend, bu, DefaultRegMode );
	 RETURN result;
     END;
     -------------------------------------------------------------------------------
     --     Function Name : Overloaded "mod" operator
     -- 1.5.21
     --     Purpose       : Modulus operator for ulogic vectors.
     --
     --     Parameters    :     result         left       right
     --                       std_ulogic_vector    INTEGER  std_ulogic_vector
     --
     --     NOTE          : The modulus operation is performed assuming all
     --                     operands and results are signed Two's complement integers.
     --
     --                     The dividend is converted to std_ulogic_vector of length
     --                     equal to the modulus. The length of the result
     --                     equals the length of the modulus.
     --
     --                     An ASSERTION message of severity ERROR is issued
     --                     if division by 0 is attempted. In this case the
     --                     return value is 0 (all 0's).
     --
     --     Use           :
     --                      VARIABLE a : INTEGER;
     --                      VARIABLE b,c : std_ulogic_vector ( 7 downto 0 );
     --                      c := a mod b;
     --                      c := 5 mod b;
     --     Se Also       : RegRem, RegDiv
     --------------------------------------------------------------------------------
     FUNCTION  "mod" ( CONSTANT dividend     : IN INTEGER;
		       CONSTANT modulus      : IN std_ulogic_vector
		     ) RETURN std_ulogic_vector IS
       VARIABLE result      : std_ulogic_vector ( modulus'LENGTH - 1 DOWNTO 0 );
       VARIABLE au          : std_ulogic_vector ( modulus'LENGTH - 1 DOWNTO 0 );
       VARIABLE zflag       : std_ulogic;
     BEGIN
     -- Convert dividend from Integer to std_ulogic_vector
	au := To_StdULogicVector(dividend, modulus'LENGTH, DefaultRegMode);
     -- Use the general modulus procedure
	 RegMod ( result, zflag,au, modulus, DefaultRegMode );
	 RETURN result;
     END;
     -------------------------------------------------------------------------------
     --     Function Name : Overloaded "mod" operator
     -- 1.5.22
     --     Purpose       : Modulus operator for bit vectors.
     --
     --     Parameters    :     result         left       right
     --                       bit_vector    bit_vector  bit_vector
     --
     --     NOTE          : The modulus operation is performed assuming all
     --                     operands and results are signed Two's complement integers.
     --
     --                     The operands may be of different length. The length of
     --                     the result equals the length of the dividend
     --
     --                     An ASSERTION message of severity ERROR is issued
     --                     if division by 0 is attempted. In this case the
     --                     return value is 0 (all 0's).
     --
     --     Use           :
     --                      VARIABLE a,b,c : bit_vector ( 7 downto 0 );
     --                      c := a mod b;
     --                      c := a mod B"1101";  -- c = a / (-3)
     --     Se Also       : RegRem, RegDiv
     ---------------------------------------------------------------------------------
     FUNCTION  "mod" ( CONSTANT dividend     : IN bit_vector;
		       CONSTANT modulus      : IN bit_vector
		     ) RETURN bit_vector IS
       VARIABLE result   : bit_vector ( dividend'LENGTH - 1 DOWNTO 0 );
       VARIABLE zflag    : BIT;
     BEGIN
     -- Use the general modulus procedure
	 RegMod ( result, zflag, dividend, modulus, DefaultRegMode );
	 RETURN result;
     END;
     -------------------------------------------------------------------------------
     --     Function Name : Overloaded "mod" operator
     -- 1.5.23
     --     Purpose       : Modulus operator for bit vectors.
     --
     --     Parameters    :     result         left       right
     --                       bit_vector     bit_vector  INTEGER
     --
     --     NOTE          : The modulus operation is performed assuming all
     --                     operands and results are signed Two's complement integers.
     --
     --                     The modulus is converted to bit_vector of length
     --                     equal to the dividend. The length of the result
     --                     equals the length of the dividend.
     --
     --                     An ASSERTION message of severity ERROR is issued
     --                     if division by 0 is attempted. In this case the
     --                     return value is 0 (all 0's).
     --
     --     Use           :
     --                      VARIABLE a,c : bit_vector ( 7 downto 0 );
     --                      VARIABLE b : INTEGER;
     --                      c := a mod b;
     --                      c := a mod 5;
     --     Se Also       : RegRem, RegDiv
     --------------------------------------------------------------------------------
     FUNCTION  "mod" ( CONSTANT dividend     : IN bit_vector;
		       CONSTANT modulus      : IN INTEGER
		     ) RETURN bit_vector IS
       VARIABLE result     : bit_vector ( dividend'LENGTH - 1 DOWNTO 0 );
       VARIABLE bv         : bit_vector ( dividend'LENGTH - 1 DOWNTO 0 );
       VARIABLE zflag      : bit;
     BEGIN
     -- Convert modulus from Integer to bit_vector
	bv := To_BitVector(modulus, dividend'LENGTH, DefaultRegMode);
     -- Use the general modulus procedure
	 RegMod ( result, zflag, dividend, bv,  DefaultRegMode );
	 RETURN result;
     END;
     -------------------------------------------------------------------------------
     --     Function Name : Overloaded "mod" operator
     -- 1.5.24
     --     Purpose       : Modulus operator for bit vectors.
     --
     --     Parameters    :     result         left       right
     --                       bit_vector    INTEGER  bit_vector
     --
     --     NOTE          : The modulus operation is performed assuming all
     --                     operands and results are signed Two's complement integers.
     --
     --                     The dividend is converted to bit_vector of length
     --                     equal to the modulus. The length of the result
     --                     equals the length of the modulus.
     --
     --                     An ASSERTION message of severity ERROR is issued
     --                     if division by 0 is attempted. In this case the
     --                     return value is 0 (all 0's).
     --
     --     Use           :
     --                      VARIABLE a : INTEGER;
     --                      VARIABLE b,c : bit_vector ( 7 downto 0 );
     --                      c := a mod b;
     --                      c := 5 mod b;
     --     Se Also       : RegRem, RegDiv
     --------------------------------------------------------------------------------
     FUNCTION  "mod" ( CONSTANT dividend     : IN INTEGER;
		       CONSTANT modulus      : IN bit_vector
		     ) RETURN bit_vector IS
       VARIABLE result     : bit_vector ( modulus'LENGTH - 1 DOWNTO 0 );
       VARIABLE av         : bit_vector ( modulus'LENGTH - 1 DOWNTO 0 );
       VARIABLE zflag      : BIT;
     BEGIN
     -- Convert dividend from Integer to bit_vector
	av := To_BitVector(dividend, modulus'LENGTH, DefaultRegMode);
     -- Use the general division procedure
	RegMod ( result, zflag, av, modulus, DefaultRegMode);
	RETURN result;
     END;
     -------------------------------------------------------------------------------
     --     Function Name : Overloaded "rem" operator
     -- 1.5.27
     --     Purpose       : Remainder operator for logic vectors.
     --
     --     Parameters    :     result         left             right
     --                     std_logic_vector  std_logic_vector  std_logic_vector
     --
     --     NOTE          : The division operation is performed assuming all
     --                     operands and results are signed Two's complement integers.
     --
     --                     The operands may be of different length. The length of
     --                     the result equals the length of the dividend.
     --
     --                     An ASSERTION message of severity ERROR is issued
     --                     if division by 0 is attempted. In this case the
     --                     return value is 0 (all 0's).
     --
     --     Use           :
     --                      VARIABLE a,b,c : std_logic_vector ( 7 downto 0 );
     --                      c := a rem b;
     --                      c := a rem B"1101";  -- c = a rem (-3)
     -----------------------------------------------------------------------------------
     FUNCTION  "rem" ( CONSTANT dividend     : IN std_logic_vector;
		       CONSTANT divisor      : IN std_logic_vector
		     ) RETURN std_logic_vector IS
       VARIABLE result   : std_logic_vector ( dividend'LENGTH - 1 DOWNTO 0 );
       VARIABLE zflag    : std_ulogic;
     BEGIN
     -- Use the general remainder procedure
	 RegRem ( result,zflag,  dividend, divisor, DefaultRegMode );
	 RETURN result;
     END;
     ---------------------------------------------------------------------------------
     --     Function Name : Overloaded "rem" operator
     -- 1.5.28
     --     Purpose       : Remainder operator for logic vectors.
     --
     --     Parameters    :     result         left       right
     --                       std_logic_vector    std_logic_vector  INTEGER
     --
     --     NOTE          : The division operation is performed assuming all
     --                     operands and results are signed Two's complement integers.
     --
     --                     The divisor is converted to std_logic_vector of length
     --                     equal to the dividend. The length of the result
     --                     equals the length of the dividend.
     --
     --                     An ASSERTION message of severity ERROR is issued
     --                     if division by 0 is attempted. In this case the
     --                     return value is 0 (all 0's).
     --
     --     Use           :
     --                      VARIABLE a,c : std_logic_vector ( 7 downto 0 );
     --                      VARIABLE b : INTEGER;
     --                      c := a rem b;
     --                      c := a rem 5;
     --     Se Also       : RegMod, RegDiv
     --------------------------------------------------------------------------------
     FUNCTION  "rem" ( CONSTANT dividend     : IN std_logic_vector;
		       CONSTANT divisor      : IN INTEGER
		     ) RETURN std_logic_vector IS
       VARIABLE result     : std_logic_vector ( dividend'LENGTH - 1 DOWNTO 0 );
       VARIABLE bv         : std_logic_vector ( dividend'LENGTH - 1 DOWNTO 0 );
       VARIABLE zflag      : std_ulogic;
     BEGIN
     -- Convert divisor from Integer to std_logic_vector
	bv := To_StdLogicVector(divisor, dividend'LENGTH, DefaultRegMode);
     -- Use the general remainder procedure
	 RegRem ( result, zflag, dividend, bv, DefaultRegMode );
	 RETURN result;
     END;
     -------------------------------------------------------------------------------
     --     Function Name : Overloaded "rem" operator
     -- 1.5.29
     --     Purpose       : Remainder operator for logic vectors.
     --
     --     Parameters    :     result         left       right
     --                       std_logic_vector    INTEGER  std_logic_vector
     --
     --     NOTE          : The division operation is performed assuming all
     --                     operands and results are signed Two's complement integers.
     --
     --                     The dividend is converted to std_logic_vector of length
     --                     equal to the divisor. The length of the result
     --                     equals the length of the divisor.
     --
     --                     An ASSERTION message of severity ERROR is issued
     --                     if division by 0 is attempted. In this case the
     --                     return value is 0 (all 0's).
     --
     --     Use           :
     --                      VARIABLE a : INTEGER;
     --                      VARIABLE b,c : std_logic_vector ( 7 downto 0 );
     --                      c := a rem b;
     --                      c := 5 rem b;
     --     Se Also       : RegMod, RegDiv
     ------------------------------------------------------------------------------
     FUNCTION  "rem" ( CONSTANT dividend     : IN INTEGER;
		       CONSTANT divisor      : IN std_logic_vector
		     ) RETURN std_logic_vector IS
       VARIABLE result      : std_logic_vector ( divisor'LENGTH - 1 DOWNTO 0 );
       VARIABLE av          : std_logic_vector ( divisor'LENGTH - 1 DOWNTO 0 );
       VARIABLE zflag       : std_ulogic;
     BEGIN
     -- Convert dividend from Integer to std_logic_vector
	av := To_StdLogicVector(dividend, divisor'LENGTH, DefaultRegMode);
     -- Use the general remainder procedure
	RegRem ( result, zflag, av, divisor, DefaultRegMode );
	RETURN result;
     END;
     -------------------------------------------------------------------------------
     --     Function Name : Overloaded "rem" operator
     -- 
     --     Purpose       : Remainder operator for ulogic vectors.
     --
     --     Parameters    :     result         left             right
     --                     std_ulogic_vector  std_ulogic_vector  std_ulogic_vector
     --
     --     NOTE          : The division operation is performed assuming all
     --                     operands and results are signed Two's complement integers.
     --
     --                     The operands may be of different length. The length of
     --                     the result equals the length of the dividend.
     --
     --                     An ASSERTION message of severity ERROR is issued
     --                     if division by 0 is attempted. In this case the
     --                     return value is 0 (all 0's).
     --
     --     Use           :
     --                      VARIABLE a,b,c : std_ulogic_vector ( 7 downto 0 );
     --                      c := a rem b;
     --                      c := a rem B"1101";  -- c = a rem (-3)
     ---------------------------------------------------------------------------------
     FUNCTION  "rem" ( CONSTANT dividend     : IN std_ulogic_vector;
		       CONSTANT divisor      : IN std_ulogic_vector
		     ) RETURN std_ulogic_vector IS
       VARIABLE result   : std_ulogic_vector ( dividend'LENGTH - 1 DOWNTO 0 );
       VARIABLE zflag    : std_ulogic;
     BEGIN
     -- Use the general remainder procedure
	 RegRem ( result, zflag, dividend, divisor, DefaultRegMode );
	 RETURN result;
     END;
     -------------------------------------------------------------------------------
     --     Function Name : Overloaded "rem" operator
     -- 
     --     Purpose       : Remainder operator for ulogic vectors.
     --
     --     Parameters    :     result         left       right
     --                       std_ulogic_vector    std_ulogic_vector  INTEGER
     --
     --     NOTE          : The division operation is performed assuming all
     --                     operands and results are signed Two's complement integers.
     --
     --                     The divisor is converted to std_ulogic_vector of length
     --                     equal to the dividend. The length of the result
     --                     equals the length of the dividend.
     --
     --                     An ASSERTION message of severity ERROR is issued
     --                     if division by 0 is attempted. In this case the
     --                     return value is 0 (all 0's).
     --
     --     Use           :
     --                      VARIABLE a,c : std_ulogic_vector ( 7 downto 0 );
     --                      VARIABLE b : INTEGER;
     --                      c := a rem b;
     --                      c := a rem 5;
     --     Se Also       : RegMod, RegDiv
     -------------------------------------------------------------------------------
     FUNCTION  "rem" ( CONSTANT dividend     : IN std_ulogic_vector;
		       CONSTANT divisor      : IN INTEGER
		     ) RETURN std_ulogic_vector IS
       VARIABLE result     : std_ulogic_vector ( dividend'LENGTH - 1 DOWNTO 0 );
       VARIABLE bu         : std_ulogic_vector ( dividend'LENGTH - 1 DOWNTO 0 );
       VARIABLE zflag      : std_ulogic;
     BEGIN
     -- Convert divisor from Integer to std_ulogic_vector
	bu := To_StdULogicVector(divisor, dividend'LENGTH, DefaultRegMode);
     -- Use the general remainder procedure
	 RegRem ( result, zflag,  dividend, bu, DefaultRegMode );
	 RETURN result;
     END;
     -------------------------------------------------------------------------------
     --     Function Name : Overloaded "rem" operator
     -- 1.5.29
     --     Purpose       : Remainder operator for ulogic vectors.
     --
     --     Parameters    :     result         left       right
     --                       std_ulogic_vector    INTEGER  std_ulogic_vector
     --
     --     NOTE          : The division operation is performed assuming all
     --                     operands and results are signed Two's complement integers.
     --
     --                     The dividend is converted to std_ulogic_vector of length
     --                     equal to the divisor. The length of the result
     --                     equals the length of the divisor.
     --
     --                     An ASSERTION message of severity ERROR is issued
     --                     if division by 0 is attempted. In this case the
     --                     return value is 0 (all 0's).
     --
     --     Use           :
     --                      VARIABLE a : INTEGER;
     --                      VARIABLE b,c : std_ulogic_vector ( 7 downto 0 );
     --                      c := a rem b;
     --                      c := 5 rem b;
     --     Se Also       : RegMod, RegDiv
     --------------------------------------------------------------------------------
     FUNCTION  "rem" ( CONSTANT dividend     : IN INTEGER;
		       CONSTANT divisor      : IN std_ulogic_vector
		     ) RETURN std_ulogic_vector IS
       VARIABLE result      : std_ulogic_vector ( divisor'LENGTH - 1 DOWNTO 0 );
       VARIABLE au          : std_ulogic_vector ( divisor'LENGTH - 1 DOWNTO 0 );
       VARIABLE zflag       : std_ulogic;
     BEGIN
     -- Convert dividend from Integer to std_ulogic_vector
	au := To_StdULogicVector(dividend, divisor'LENGTH, DefaultRegMode);
     -- Use the general remainder procedure
	 RegRem ( result, zflag, au, divisor, DefaultRegMode );
	 RETURN result;
     END;
 --+-----------------------------------------------------------------------------
 --|     Function Name : Overloaded "rem" operator
 --| 1.5.30
 --|     Purpose       : Remainder operator for bit vectors.
 --|     Parameters    :     result         left       right
 --|                       BIT_VECTOR    BIT_VECTOR  BIT_VECTOR
 --|
 --|     NOTE          : The division operation is performed assuming all
 --|                     operands and results are signed Two's complement integers.
 --|
 --|                     The operands may be of different length. The length of
 --|                     the result equals the length of the longer operand.
 --|
 --|                     An ASSERTION message of severity ERROR is issued
 --|                     if division by 0 is attempted. In this case the
 --|                     return value is 0 (all 0's).
 --|
 --|     Use           :
 --|                      VARIABLE a,b,c : bit_vector ( 7 downto 0 );
 --|                      c := a rem b;
 --|                      c := a rem B"1101";  -- c = a rem (-3)
 --|
 --|     See Also      : RegMod, RegDiv
 --|-----------------------------------------------------------------------------
     FUNCTION  "rem" ( CONSTANT dividend     : IN BIT_VECTOR;
		       CONSTANT divisor      : IN BIT_VECTOR
		     ) RETURN BIT_VECTOR IS
       VARIABLE result   : BIT_VECTOR ( dividend'LENGTH - 1 DOWNTO 0 );
       VARIABLE zflag    : BIT;
     BEGIN
     -- Use the general remainder procedure
	 RegRem ( result, zflag, dividend, divisor, DefaultRegMode );
	 RETURN result;
     END;
 --+-----------------------------------------------------------------------------
 --|     Function Name : Overloaded "rem" operator
 --| 1.5.31
 --|     Purpose       : Remainder operator for bit vectors.
 --|     Parameters    :     result         left       right
 --|                       BIT_VECTOR    BIT_VECTOR  INTEGER
 --|
 --|     NOTE          : The division operation is performed assuming all
 --|                     operands and results are signed Two's complement integers.
 --|
 --|                     The divisor is converted to bit_vector of length
 --|                     equal to the dividend. The length of the result
 --|                     equals the length of the dividend.
 --|
 --|                     An ASSERTION message of severity ERROR is issued
 --|                     if division by 0 is attempted. In this case the
 --|                     return value is 0 (all 0's).
 --|
 --|
 --|     Use           :
 --|                      VARIABLE a,c : BIT_VECTOR ( 7 downto 0 );
 --|                      VARIABLE b : INTEGER;
 --|                      c := a rem b;
 --|                      c := a rem 5;
 --|
 --|     See Also      : RegMod, RegDiv
 --|-----------------------------------------------------------------------------
     FUNCTION  "rem" ( CONSTANT dividend     : IN BIT_VECTOR;
		       CONSTANT divisor      : IN INTEGER
		     ) RETURN BIT_VECTOR IS
       VARIABLE result    : BIT_VECTOR ( dividend'LENGTH - 1 DOWNTO 0 );
       VARIABLE bv        : BIT_VECTOR ( dividend'LENGTH - 1 DOWNTO 0 );
       VARIABLE zflag     : BIT;
     BEGIN
     -- Convert divisor from Integer to bit_vector
	bv := To_BitVector(divisor, dividend'LENGTH, DefaultRegMode);
     -- Use the general remainder procedure
	 RegRem ( result, zflag, dividend, bv, DefaultRegMode );
	 RETURN result;
     END;
 --+-----------------------------------------------------------------------------
 --|     Function Name : Overloaded "rem" operator
 --| 1.5.32
 --|     Purpose       : Remainder operator for bit vectors.
 --|     Parameters    :     result         left       right
 --|                       BIT_VECTOR    INTEGER  BIT_VECTOR
 --|
 --|     NOTE          : The division operation is performed assuming all
 --|                     operands and results are signed Two's complement integers.
 --|
 --|                     The dividend is converted to bit_vector of length
 --|                     equal to the divisor. The length of the result
 --|                     equals the length of the divisor.
 --|
 --|                     An ASSERTION message of severity ERROR is issued
 --|                     if division by 0 is attempted. In this case the
 --|                     return value is 0 (all 0's).
 --|
 --|
 --|     Use           :
 --|                      VARIABLE a : INTEGER;
 --|                      VARIABLE b,c : BIT_VECTOR ( 7 downto 0 );
 --|                      c := a rem b;
 --|                      c := 5 rem b;
 --|
 --|     See Also      : RegMod, RegDiv
 --|-----------------------------------------------------------------------------
     FUNCTION  "rem" ( CONSTANT dividend     : IN INTEGER;
		       CONSTANT divisor      : IN BIT_VECTOR
		     ) RETURN BIT_VECTOR IS
       VARIABLE result     : BIT_VECTOR(divisor'LENGTH - 1 DOWNTO 0);
       VARIABLE av         : BIT_VECTOR(divisor'LENGTH - 1 DOWNTO 0);
       VARIABLE zflag      : BIT;
     BEGIN
     -- Convert dividend from Integer to bit_vector
	av := To_BitVector(dividend, divisor'LENGTH, DefaultRegMode);
     -- Use the general remainder procedure
	 RegRem ( result, zflag, av, divisor, DefaultRegMode );
	 RETURN result;
     END;
     -------------------------------------------------------------------------------
     --     Function Name : Overloaded "ABS" operator
     -- 1.6.11
     --     Purpose       : Absolute value operator for logic vectors.
     --
     --     Parameters    :     result             operand       
     --                       std_logic_vector    std_logic_vector
     --
     --
     --     Use           :
     --                      VARIABLE a,c : std_logic_vector ( 7 downto 0 );
     --                      c := ABS(a);
     --
     --     See Also      : RegAbs
     -------------------------------------------------------------------------------
     FUNCTION  "ABS" ( CONSTANT operand : IN std_logic_vector
		     ) RETURN std_logic_vector IS
       VARIABLE result   : std_logic_vector ( operand'LENGTH - 1 DOWNTO 0 );
     BEGIN
     --
     -- Use the general absolute value  procedure with DefaultRegMode mode
	 RegAbs ( result, operand, DefaultRegMode);
	 RETURN result;
     END;
     -------------------------------------------------------------------------------
     --     Function Name : Overloaded "ABS" operator
     -- 
     --     Purpose       : Absolute value operator for ulogic vectors.
     --
     --     Parameters    :     result             operand       
     --                       std_ulogic_vector    std_ulogic_vector
     --
     --
     --     Use           :
     --                      VARIABLE a,c : std_ulogic_vector ( 7 downto 0 );
     --                      c := ABS(a);
     --
     --     See Also      : RegAbs
     -------------------------------------------------------------------------------
     FUNCTION  "ABS" ( CONSTANT operand : IN std_ulogic_vector
		     ) RETURN std_ulogic_vector IS
       VARIABLE result   : std_ulogic_vector ( operand'LENGTH - 1 DOWNTO 0 );
     BEGIN
     --
     -- Use the general absolute value  procedure with DefaultRegMode mode
	 RegAbs ( result, operand, DefaultRegMode);
	 RETURN result;
     END;
     -------------------------------------------------------------------------------
     --     Function Name : Overloaded "ABS" operator
     -- 1.6.12
     --     Purpose       : Absolute value operator for bit vectors.
     --
     --     Parameters    :     result        operand       
     --                       bit_vector    bit_vector
     --
     --
     --     Use           :
     --                      VARIABLE a,c : bit_vector ( 7 downto 0 );
     --                      c := ABS(a);
     --
     --     See Also      : RegAbs
     -------------------------------------------------------------------------------
     FUNCTION  "ABS" ( CONSTANT operand : IN bit_vector
		     ) RETURN bit_vector IS
       VARIABLE result   : bit_vector ( operand'LENGTH - 1 DOWNTO 0 );
     BEGIN
     -- Use the general absolute value  procedure with DefaultRegMode Mode
	 RegAbs ( result, operand, DefaultRegMode);
	 RETURN result;
     END;
     -------------------------------------------------------------------------------
     --     Function Name : Overloaded "=" operator
     --   1.2.1 and 1.2.3  
     --     Purpose       : Equality relational operator for std_logic_vector : integer.
     --     
     --     Parameters    :     result         left              right
     --                        std_ulogic  std_logic_vector   std_logic_vector
     --                        BOOLEAN     INTEGER            std_logic_vector
     --                        BOOLEAN     std_logic_vector   INTEGER
     --                        std_ulogic  INTEGER            std_logic_vector
     --                        std_ulogic  std_logic_vector   INTEGER
     --                                     
     --     NOTE          : The std_logic_vector operands are assumed to be  
     --                     in  DefaultRegMode. If not they will be converted
     --                     to DefaultRegMode in the compare procedure. 
     --                     These vectors may be of any length.
     --
     --     Use           : 
     --                      VARIABLE a : std_logic_vector ( 7 DOWNTO 0 ) := X"FF";
     --                      VARIABLE b : INTEGER;
     --                      IF ( a = b )  THEN 
     --     
     --     See Also      : RegEqual, RegNotEqual,
     -------------------------------------------------------------------------------
     FUNCTION  "=" ( CONSTANT l  : std_logic_vector;
		     CONSTANT r  : std_logic_vector
		   ) RETURN std_ulogic IS
       VARIABLE eq : std_ulogic;
     BEGIN
	-- Use RegEqual with DefaultRegMode mode
	eq := RegEqual (l,r, DefaultRegMode);
	return eq;
     END;
     -------------------------------------------------------------------------------
     FUNCTION  "=" ( CONSTANT l  : std_logic_vector;
		     CONSTANT r  : INTEGER
		   ) RETURN BOOLEAN IS
	VARIABLE eq  : boolean;
	VARIABLE rv  : std_logic_vector (IntegerBitLength - 1 downto 0);
     BEGIN
        -- Convert to std_logic_vector for comparison to allow any length input vector.
	rv := To_StdLogicVector (r, IntegerBitLength, DefaultRegMode);
	-- Use RegEqual with DefaultRegMode mode
	eq := RegEqual (l, rv, DefaultRegMode);
	RETURN eq;
     END;
     -- -----------------------------------------------------------------------------
     FUNCTION  "=" ( CONSTANT l  : INTEGER   ;
		     CONSTANT r  : std_logic_vector 
		   ) RETURN BOOLEAN IS
        VARIABLE eq  : boolean;
	VARIABLE lv  : std_logic_vector (IntegerBitLength - 1 downto 0);
     BEGIN
        -- Convert to std_logic_vectors for comparison to allow any length input vector.
	lv := To_StdLogicVector (l, IntegerBitLength, DefaultRegMode);
	-- Use RegEqual with DefaultRegMode mode
	eq := RegEqual (lv, r, DefaultRegMode);
	RETURN eq;
     END;
     -------------------------------------------------------------------------------
     FUNCTION  "=" ( CONSTANT l  : std_logic_vector;
		     CONSTANT r  : INTEGER
		   ) RETURN std_ulogic IS
	VARIABLE eq   : std_ulogic;
	VARIABLE rv  : std_logic_vector (IntegerBitLength - 1 downto 0);
     BEGIN
        -- Convert to std_logic_vector for comparison to allow any length input vector.
	rv := To_StdLogicVector (r, IntegerBitLength, DefaultRegMode);
	-- Use RegEqual with DefaultRegMode mode
	eq := RegEqual (l, rv,  DefaultRegMode);
	RETURN eq;
     END;
     -- -----------------------------------------------------------------------------
     FUNCTION  "=" ( CONSTANT l  : INTEGER   ;
		     CONSTANT r  : std_logic_vector 
		   ) RETURN std_ulogic IS
	VARIABLE eq  : std_ulogic;
	VARIABLE lv  : std_logic_vector (IntegerBitLength - 1 downto 0);
     BEGIN
        -- Convert to std_logic_vector for comparison to allow any length input vector.
	lv := To_StdLogicVector (l, IntegerBitLength, DefaultRegMode);
	-- Use RegEqual with DefaultRegMode mode
	eq := RegEqual (lv,  r, DefaultRegMode);
	RETURN eq;
     END;
     -------------------------------------------------------------------------------
     --     Function Name : Overloaded "=" operator
     --   1.2.1 and 1.2.3  
     --     Purpose       : Equality relational operator for std_ulogic_vector : integer.
     --     
     --     Parameters    :     result         left              right
     --                        std_ulogic  std_ulogic_vector   std_ulogic_vector
     --                        BOOLEAN     INTEGER            std_ulogic_vector
     --                        BOOLEAN     std_ulogic_vector   INTEGER
     --                        std_ulogic  INTEGER            std_ulogic_vector
     --                        std_ulogic  std_ulogic_vector   INTEGER
     --                                     
     --     NOTE          : The std_ulogic_vector operands are assumed to be  
     --                     in  DefaultRegMode. If not they will be converted
     --                     to DefaultRegMode in the compare procedure. 
     --                     These vectors may be of any length.
     --
     --     Use           : 
     --                      VARIABLE a : std_ulogic_vector ( 7 DOWNTO 0 ) := X"FF";
     --                      VARIABLE b : INTEGER;
     --                      IF ( a = b )  THEN 
     --     
     --     See Also      : RegEqual, RegNotEqual,
     -------------------------------------------------------------------------------
     FUNCTION  "=" ( CONSTANT l  : std_ulogic_vector;
		     CONSTANT r  : std_ulogic_vector
		   ) RETURN std_ulogic IS
       VARIABLE eq : std_ulogic;
     BEGIN
	-- Use RegEqual with DefaultRegMode mode
	eq := RegEqual (l,r, DefaultRegMode);
	return eq;
     END;
     -------------------------------------------------------------------------------
     FUNCTION  "=" ( CONSTANT l  : std_ulogic_vector;
		     CONSTANT r  : INTEGER
		   ) RETURN BOOLEAN IS
	VARIABLE eq  : boolean;
	VARIABLE rv  : std_ulogic_vector (IntegerBitLength - 1 downto 0);
     BEGIN
        -- Convert to std_ulogic_vectors for comparison to allow any length input vector.
	rv := To_StdULogicVector (r, IntegerBitLength, DefaultRegMode);
	-- Use RegEqual with DefaultRegMode mode
	eq := RegEqual (l, rv, DefaultRegMode);
	RETURN eq;
     END;
     -- -----------------------------------------------------------------------------
     FUNCTION  "=" ( CONSTANT l  : INTEGER   ;
		     CONSTANT r  : std_ulogic_vector 
		   ) RETURN BOOLEAN IS
        VARIABLE eq  : boolean;
	VARIABLE lv  : std_ulogic_vector (IntegerBitLength - 1 downto 0);
     BEGIN
        -- Convert to std_ulogic_vectors for comparison to allow any length input vector.
	lv := To_StdULogicVector (l, IntegerBitLength, DefaultRegMode);
	-- Use RegEqual with DefaultRegMode mode
	eq := RegEqual (lv, r, DefaultRegMode);
	RETURN eq;
     END;
     -------------------------------------------------------------------------------
     FUNCTION  "=" ( CONSTANT l  : std_ulogic_vector;
		     CONSTANT r  : INTEGER
		   ) RETURN std_ulogic IS
        VARIABLE eq   : std_ulogic;
	VARIABLE rv  : std_ulogic_vector (IntegerBitLength - 1 downto 0);
     BEGIN
        -- Convert to std_ulogic_vectors for comparison to allow any length input vector.
	rv := To_StdULogicVector (r, IntegerBitLength, DefaultRegMode);
 	-- Use RegEqual with DefaultRegMode mode
	eq := RegEqual (l, rv, DefaultRegMode);
	RETURN eq;
     END;
     -- -----------------------------------------------------------------------------
     FUNCTION  "=" ( CONSTANT l  : INTEGER   ;
		     CONSTANT r  : std_ulogic_vector 
		   ) RETURN std_ulogic IS
        VARIABLE eq : std_ulogic;
	VARIABLE lv  : std_ulogic_vector (IntegerBitLength - 1 downto 0);
     BEGIN
        -- Convert to std_ulogic_vectors for comparison to allow any length input vector.
	lv := To_StdULogicVector (l, IntegerBitLength, DefaultRegMode);
	-- Use RegEqual with DefaultRegMode mode
	eq := RegEqual (lv, r, DefaultRegMode);
	RETURN eq;
     END;
     -------------------------------------------------------------------------------
     --     Function Name : Overloaded "=" operator
     -- 1.2.2 and 1.2.4
     --     Purpose       : Equality relational operator for bit_vector : integer.
     --
     --     Parameters    :     result         left       right
     --                        BOOLEAN       INTEGER   bit_vector 
     --                        BOOLEAN      bit_vector   INTEGER
     --
     --     NOTE          : The bit_vector operands are assumed to be 
     --                     in  DefaultRegMode. If not they will be converted
     --                     to DefaultRegMode in the compare procedure. 
     --                     These vectors may be of any length.
     --
     --     Use           :
     --                      VARIABLE a : bit_vector ( 7 DOWNTO 0 ) := X"FF";
     --                      VARIABLE b : INTEGER;
     --                      IF ( a = b )  THEN
     --
     --     See Also      :  RegLessThan, RegGreaterThan,
     -------------------------------------------------------------------------------
     FUNCTION  "=" ( CONSTANT l  : bit_vector;
		     CONSTANT r  : bit_vector
		   ) RETURN bit IS
	VARIABLE eq : BIT;    
     BEGIN
	-- Use RegEqual with DefaultRegMode mode
	eq := RegEqual (l,r, DefaultRegMode);
	return eq;
     END;
     -------------------------------------------------------------------------------
     FUNCTION  "=" ( CONSTANT l  : bit_vector;
		     CONSTANT r  : INTEGER
		   ) RETURN BOOLEAN IS
	VARIABLE eq  : Boolean;
	VARIABLE rv  : bit_vector (IntegerBitLength - 1 downto 0);
     BEGIN
        -- Convert to bit_vector for comparison to allow any length input vector.
	rv := To_BitVector (r, IntegerBitLength, DefaultRegMode);
	-- Use RegEqual with DefaultRegMode mode
	eq := RegEqual (l, rv, DefaultRegMode);
	return eq;
     END;
     -- -----------------------------------------------------------------------------
     FUNCTION  "=" ( CONSTANT l  : INTEGER   ;
		     CONSTANT r  : bit_vector 
		   ) RETURN BOOLEAN IS
        VARIABLE eq  : boolean;
	VARIABLE lv  : bit_vector (IntegerBitLength - 1 downto 0);
     BEGIN
        -- Convert to bit_vector for comparison to allow any length input vector.
	lv := To_BitVector (l, IntegerBitLength, DefaultRegMode);
	-- Use RegEqual with DefaultRegMode mode
	eq := RegEqual (lv, r, DefaultRegMode);
	return eq;
     END;
     -------------------------------------------------------------------------------
     FUNCTION  "=" ( CONSTANT l  : bit_vector;
		     CONSTANT r  : INTEGER
		   ) RETURN bit IS
        VARIABLE eq : bit;
	VARIABLE rv  : bit_vector (IntegerBitLength - 1 downto 0);
     BEGIN
        -- Convert to bit_vector for comparison to allow any length input vector.
	rv := To_BitVector (r, IntegerBitLength, DefaultRegMode);
 	-- Use RegEqual with DefaultRegMode mode
	eq := RegEqual (l, rv, DefaultRegMode);
	return eq;
     END;
     -- -----------------------------------------------------------------------------
     FUNCTION  "=" ( CONSTANT l  : INTEGER   ;
		     CONSTANT r  : bit_vector 
		   ) RETURN bit IS
          VARIABLE eq    :bit;
	VARIABLE lv  : bit_vector (IntegerBitLength - 1 downto 0);
     BEGIN
        -- Convert to bit_vector for comparison to allow any length input vector.
	lv := To_BitVector (l, IntegerBitLength, DefaultRegMode);
	-- Use RegEqual with DefaultRegMode mode
	eq := RegEqual (lv,  r, DefaultRegMode);
	return eq;
     END;
     -------------------------------------------------------------------------------
     --     Function Name : Overloaded "/=" operator
     --   1.2.1 and 1.2.3  
     --     Purpose       : Un-equality relational operator for std_logic_vector : integer.
     --     
     --     Parameters    :     result         left              right
     --                        std_ulogic  std_logic_vector   std_logic_vector
     --                        BOOLEAN     INTEGER            std_logic_vector
     --                        BOOLEAN     std_logic_vector   INTEGER
     --                        std_ulogic  INTEGER            std_logic_vector
     --                        std_ulogic  std_logic_vector   INTEGER
     --                                     
     --     NOTE          : The std_logic_vector operands are assumed to be  
     --                     in  DefaultRegMode. If not they will be converted
     --                     to DefaultRegMode.
     --                     These vectors may be of any length.
     --
     --     Use           : 
     --                      VARIABLE a : std_logic_vector ( 7 DOWNTO 0 ) := X"FF";
     --                      VARIABLE b : INTEGER;
     --                      IF ( a /= b )  THEN 
     --     
     --     See Also      : RegEqual, RegNotEqual,
     -------------------------------------------------------------------------------
     FUNCTION  "/=" ( CONSTANT l  : std_logic_vector;
		     CONSTANT r  : std_logic_vector
		   ) RETURN std_ulogic IS
       VARIABLE neq : std_ulogic;
     BEGIN
	-- Use RegNotEqual with DefaultRegMode mode
	neq := RegNotEqual (l,r, DefaultRegMode);
	return neq;
     END;
     -------------------------------------------------------------------------------
     FUNCTION  "/=" ( CONSTANT l  : std_logic_vector;
		     CONSTANT r  : INTEGER
		   ) RETURN BOOLEAN IS
	VARIABLE neq  : boolean;
	VARIABLE rv  : std_logic_vector (IntegerBitLength - 1 downto 0);
     BEGIN
        -- Convert to std_logic_vector for comparison to allow any length input vector.
	rv := To_StdLogicVector (r, IntegerBitLength, DefaultRegMode);
	-- Use RegNotEqual with DefaultRegMode mode
	neq := RegNotEqual (l, rv, DefaultRegMode);
	RETURN neq;
     END;
     -- -----------------------------------------------------------------------------
     FUNCTION  "/=" ( CONSTANT l  : INTEGER   ;
		     CONSTANT r  : std_logic_vector 
		   ) RETURN BOOLEAN IS
        VARIABLE neq  : boolean;
	VARIABLE lv  : std_logic_vector (IntegerBitLength - 1 downto 0);
     BEGIN
        -- Convert to std_logic_vector for comparison to allow any length input vector.
	lv := To_StdLogicVector (l, IntegerBitLength, DefaultRegMode);
	-- Use RegNotEqual with DefaultRegMode mode
	neq := RegNotEqual (lv, r, DefaultRegMode);
	RETURN neq;
     END;
     -------------------------------------------------------------------------------
     FUNCTION  "/=" ( CONSTANT l  : std_logic_vector;
		     CONSTANT r  : INTEGER
		   ) RETURN std_ulogic IS
	VARIABLE neq   : std_ulogic;
	VARIABLE rv  : std_logic_vector (IntegerBitLength - 1 downto 0);
     BEGIN
        -- Convert to std_logic_vector for comparison to allow any length input vector.
	rv := To_StdLogicVector (r, IntegerBitLength, DefaultRegMode);
	-- Use RegNotEqual with DefaultRegMode mode
	neq := RegNotEqual (l, rv,  DefaultRegMode);
	RETURN neq;
     END;
     -- -----------------------------------------------------------------------------
     FUNCTION  "/=" ( CONSTANT l  : INTEGER   ;
		     CONSTANT r  : std_logic_vector 
		   ) RETURN std_ulogic IS
	VARIABLE neq  : std_ulogic;
	VARIABLE lv  : std_logic_vector (IntegerBitLength - 1 downto 0);
     BEGIN
        -- Convert to std_logic_vector for comparison to allow any length input vector.
	lv := To_StdLogicVector (l, IntegerBitLength, DefaultRegMode);
	-- Use RegNotEqual with DefaultRegMode mode
	neq := RegNotEqual (lv,  r, DefaultRegMode);
	RETURN neq;
     END;
     -------------------------------------------------------------------------------
     --     Function Name : Overloaded "/=" operator
     --   1.2.1 and 1.2.3  
     --     Purpose       : Un-Equality relational operator for std_ulogic_vector : integer.
     --     
     --     Parameters    :     result         left              right
     --                        std_ulogic  std_ulogic_vector   std_ulogic_vector
     --                        BOOLEAN     INTEGER            std_ulogic_vector
     --                        BOOLEAN     std_ulogic_vector   INTEGER
     --                        std_ulogic  INTEGER            std_ulogic_vector
     --                        std_ulogic  std_ulogic_vector   INTEGER
     --                                     
     --     NOTE          : The std_ulogic_vector operands are assumed to be  
     --                     in  DefaultRegMode. If not they will be converted
     --                     to DefaultRegMode.
     --                     These vectors may be of any length.
     --
     --     Use           : 
     --                      VARIABLE a : std_ulogic_vector ( 7 DOWNTO 0 ) := X"FF";
     --                      VARIABLE b : INTEGER;
     --                      IF ( a /= b )  THEN 
     --     
     --     See Also      : RegEqual, RegNotEqual,
     -------------------------------------------------------------------------------
     FUNCTION  "/=" ( CONSTANT l  : std_ulogic_vector;
		     CONSTANT r  : std_ulogic_vector
		   ) RETURN std_ulogic IS
       VARIABLE neq : std_ulogic;
     BEGIN
	-- Use RegNotEqual with DefaultRegMode mode
	neq := RegNotEqual (l,r, DefaultRegMode);
	return neq;
     END;
     -------------------------------------------------------------------------------
     FUNCTION  "/=" ( CONSTANT l  : std_ulogic_vector;
		     CONSTANT r  : INTEGER
		   ) RETURN BOOLEAN IS
	VARIABLE neq  : boolean;
	VARIABLE rv  : std_ulogic_vector (IntegerBitLength - 1 downto 0);
     BEGIN
        -- Convert to std_ulogic_vectors for comparison to allow any length input vector.
	rv := To_StdULogicVector (r, IntegerBitLength, DefaultRegMode);
	-- Use RegNotEqual with DefaultRegMode mode
	neq := RegNotEqual (l, rv, DefaultRegMode);
	RETURN neq;
     END;
     -- -----------------------------------------------------------------------------
     FUNCTION  "/=" ( CONSTANT l  : INTEGER   ;
		     CONSTANT r  : std_ulogic_vector 
		   ) RETURN BOOLEAN IS
        VARIABLE neq  : boolean;
	VARIABLE lv  : std_ulogic_vector (IntegerBitLength - 1 downto 0);
     BEGIN
        -- Convert to std_ulogic_vectors for comparison to allow any length input vector.
	lv := To_StdULogicVector (l, IntegerBitLength, DefaultRegMode);
	-- Use RegNotEqual with DefaultRegMode mode
	neq := RegNotEqual (lv, r, DefaultRegMode);
	RETURN neq;
     END;
     -------------------------------------------------------------------------------
     FUNCTION  "/=" ( CONSTANT l  : std_ulogic_vector;
		     CONSTANT r  : INTEGER
		   ) RETURN std_ulogic IS
        VARIABLE neq   : std_ulogic;
	VARIABLE rv  : std_ulogic_vector (IntegerBitLength - 1 downto 0);
     BEGIN
        -- Convert to std_ulogic_vectors for comparison to allow any length input vector.
	rv := To_StdULogicVector (r, IntegerBitLength, DefaultRegMode);
 	-- Use RegNotEqual with DefaultRegMode mode
	neq := RegNotEqual (l, rv, DefaultRegMode);
	RETURN neq;
     END;
     -- -----------------------------------------------------------------------------
     FUNCTION  "/=" ( CONSTANT l  : INTEGER   ;
		     CONSTANT r  : std_ulogic_vector 
		   ) RETURN std_ulogic IS
        VARIABLE neq : std_ulogic;
	VARIABLE lv  : std_ulogic_vector (IntegerBitLength - 1 downto 0);
     BEGIN
        -- Convert to std_ulogic_vectors for comparison to allow any length input vector.
	lv := To_StdULogicVector (l, IntegerBitLength, DefaultRegMode);
	-- Use RegNotEqual with DefaultRegMode mode
	neq := RegNotEqual (lv, r, DefaultRegMode);
	RETURN neq;
     END;
     -------------------------------------------------------------------------------
     --     Function Name : Overloaded "/=" operator
     -- 1.2.2 and 1.2.4
     --     Purpose       : Un-Equality relational operator for bit_vector : integer.
     --
     --     Parameters    :     result         left       right
     --                        BOOLEAN       INTEGER   bit_vector 
     --                        BOOLEAN      bit_vector   INTEGER
     --
     --     NOTE          : The bit_vector operands are assumed to be 
     --                     in  DefaultRegMode. If not they will be converted
     --                     to DefaultRegMode .
     --                     These vectors may be of any length.
     --
     --     Use           :
     --                      VARIABLE a : bit_vector ( 7 DOWNTO 0 ) := X"FF";
     --                      VARIABLE b : INTEGER;
     --                      IF ( a /= b )  THEN
     --
     --     See Also      :  RegLessThan, RegGreaterThan,
     -------------------------------------------------------------------------------
     FUNCTION  "/=" ( CONSTANT l  : bit_vector;
		     CONSTANT r  : bit_vector
		   ) RETURN bit IS
	VARIABLE neq : BIT;    
     BEGIN
	-- Use RegNotEqual with DefaultRegMode mode
	neq := RegNotEqual (l,r, DefaultRegMode);
	return neq;
     END;
     -------------------------------------------------------------------------------
     FUNCTION  "/=" ( CONSTANT l  : bit_vector;
		     CONSTANT r  : INTEGER
		   ) RETURN BOOLEAN IS
	VARIABLE neq  : Boolean;
	VARIABLE rv  : bit_vector (IntegerBitLength - 1 downto 0);
     BEGIN
        -- Convert to bit_vector for comparison to allow any length input vector.
	rv := To_BitVector (r, IntegerBitLength, DefaultRegMode);
	-- Use RegNotEqual with DefaultRegMode mode
	neq := RegNotEqual (l, rv, DefaultRegMode);
	return neq;
     END;
     -- -----------------------------------------------------------------------------
     FUNCTION  "/=" ( CONSTANT l  : INTEGER   ;
		     CONSTANT r  : bit_vector 
		   ) RETURN BOOLEAN IS
        VARIABLE neq  : boolean;
	VARIABLE lv  : bit_vector (IntegerBitLength - 1 downto 0);
     BEGIN
        -- Convert to bit_vector for comparison to allow any length input vector.
	lv := To_BitVector (l, IntegerBitLength, DefaultRegMode);
	-- Use RegNotEqual with DefaultRegMode mode
	neq := RegNotEqual (lv, r, DefaultRegMode);
	return neq;
     END;
     -------------------------------------------------------------------------------
     FUNCTION  "/=" ( CONSTANT l  : bit_vector;
		     CONSTANT r  : INTEGER
		   ) RETURN bit IS
        VARIABLE neq : bit;
	VARIABLE rv  : bit_vector (IntegerBitLength - 1 downto 0);
     BEGIN
        -- Convert to bit_vector for comparison to allow any length input vector.
	rv := To_BitVector (r, IntegerBitLength, DefaultRegMode);
 	-- Use RegNotEqual with DefaultRegMode mode
	neq := RegNotEqual (l, rv, DefaultRegMode);
	return neq;
     END;
     -- -----------------------------------------------------------------------------
     FUNCTION  "/=" ( CONSTANT l  : INTEGER   ;
		     CONSTANT r  : bit_vector 
		   ) RETURN bit IS
          VARIABLE neq    :bit;
	VARIABLE lv  : bit_vector (IntegerBitLength - 1 downto 0);
     BEGIN
        -- Convert to bit_vector for comparison to allow any length input vector.
	lv := To_BitVector (l, IntegerBitLength, DefaultRegMode);
	-- Use RegNotEqual with DefaultRegMode mode
	neq := RegNotEqual (lv,  r, DefaultRegMode);
	return neq;
     END;
     --------------------------------------------------------------------------------
     --     Function Name : Overloaded "<" operator
     -- 1.2.18 and 1.2.20     
     --     Purpose       : Less-than relational operator for bit_vectors.
     --     
     --     Parameters    :     result         left       right
     --                        BOOLEAN       INTEGER    bit_vector
     --                        BOOLEAN      bit_vector   INTEGER
     --     
     --     NOTE          : The bit_vector operands are assumed to be 
     --                     in  DefaultRegMode. If not they will be converted
     --                     to DefaultRegMode.
     --                     These vectors may be of any length.
     --
     --     Use           :
     --                      VARIABLE a : bit_vector ( 7 DOWNTO 0 ) := X"FF";
     --                      VARIABLE b : INTEGER;
     --                      IF ( a < b )  THEN 
     --     
     --     See Also      :   RegLessThan, RegGreaterThan,
     -------------------------------------------------------------------------------
     FUNCTION  "<" ( CONSTANT l  : bit_vector;
		     CONSTANT r  : bit_vector
		   ) RETURN bit IS
	VARIABLE lt : BIT;    
     BEGIN
	-- Use RegLessThan with DefaultRegMode mode
	lt := RegLessThan (l,r, DefaultRegMode);
	return lt;
     END;
     -------------------------------------------------------------------------------
     FUNCTION  "<" ( CONSTANT l  : bit_vector;
		     CONSTANT r  : INTEGER
		   ) RETURN BOOLEAN IS
        VARIABLE lt  : Boolean;
	VARIABLE rv  : bit_vector (IntegerBitLength - 1 downto 0);
     BEGIN
        -- Convert to bit_vector for comparison to allow any length input vector.
	rv := To_BitVector (r, IntegerBitLength, DefaultRegMode);
	-- Use RegLessThan with DefaultRegMode mode
	lt := RegLessThan (l, rv , DefaultRegMode);
	return lt;
     END;
     -- -----------------------------------------------------------------------------
     FUNCTION  "<" ( CONSTANT l  : INTEGER   ;
		     CONSTANT r  : bit_vector 
		   ) RETURN BOOLEAN IS
        VARIABLE lt    : boolean;
	VARIABLE lv  : bit_vector (IntegerBitLength - 1 downto 0);
     BEGIN
        -- Convert to bit_vector for comparison to allow any length input vector.
	lv := To_BitVector (l, IntegerBitLength, DefaultRegMode);
	-- Use RegLessThan with DefaultRegMode mode
	lt := RegLessThan (lv, r, DefaultRegMode);
	return lt;
     END;
     -------------------------------------------------------------------------------
     FUNCTION  "<" ( CONSTANT l  : bit_vector;
		     CONSTANT r  : INTEGER
		   ) RETURN bit IS
       VARIABLE lt : bit;
	VARIABLE rv  : bit_vector (IntegerBitLength - 1 downto 0);
     BEGIN
        -- Convert to bit_vector for comparison to allow any length input vector.
	rv := To_BitVector (r, IntegerBitLength, DefaultRegMode);
	-- Use RegLessThan with DefaultRegMode mode
	lt := RegLessThan (l, rv, DefaultRegMode);
	return lt;
     END;
     -- -----------------------------------------------------------------------------
     FUNCTION  "<" ( CONSTANT l  : INTEGER   ;
		     CONSTANT r  : bit_vector 
		   ) RETURN bit IS
        VARIABLE lt  : bit;
	VARIABLE lv  : bit_vector (IntegerBitLength - 1 downto 0);
     BEGIN
        -- Convert to bit_vector for comparison to allow any length input vector.
	lv := To_BitVector (l, IntegerBitLength, DefaultRegMode);
	-- Use RegLessThan with DefaultRegMode mode
	lt := RegLessThan (lv, r, DefaultRegMode);
	return lt;
     END;
     -------------------------------------------------------------------------------
     --     Function Name : Overloaded "<" operator
     --
     --     Purpose       : Less-than relational operator for std_logic_vectors.
     --
     --     Parameters    :     result         left       right
     --                        std_ulogic  std_logic_vector   std_logic_vector
     --                        BOOLEAN     INTEGER            std_logic_vector
     --                        BOOLEAN     std_logic_vector   INTEGER
     --                        std_ulogic  INTEGER            std_logic_vector
     --                        std_ulogic  std_logic_vector   INTEGER
     --
     --     NOTE          : The std_logic_vector operands are assumed to be 
     --                     in  DefaultRegMode. If not they will be converted
     --                     to DefaultRegMode.
     --                     These vectors may be of any length.
     --
     --     Use           :
     --                      VARIABLE a : std_logic_vector ( 7 DOWNTO 0 ) := X"FF";
     --                      VARIABLE b : INTEGER;
     --                      IF ( a < b )  THEN
     --
     --     See Also      :   RegLessThan, RegGreaterThan,
     -------------------------------------------------------------------------------
     FUNCTION  "<" ( CONSTANT l  : std_logic_vector;
		     CONSTANT r  : std_logic_vector
		   ) RETURN std_ulogic IS
       VARIABLE lt : std_ulogic;
     BEGIN
	-- Use RegLessThan with DefaultRegMode mode
	lt := RegLessThan (l,r, DefaultRegMode);
	return lt;
     END;
     -------------------------------------------------------------------------------
     FUNCTION  "<" ( CONSTANT l  : std_logic_vector;
		     CONSTANT r  : INTEGER
		   ) RETURN BOOLEAN IS
        VARIABLE lt  : boolean;
	VARIABLE rv  : std_logic_vector (IntegerBitLength - 1 downto 0);
     BEGIN
        -- Convert to bit_vector for comparison to allow any length input vector.
	rv := To_StdLogicVector (r, IntegerBitLength, DefaultRegMode);
	-- Use RegLessThan with DefaultRegMode mode
	lt := RegLessThan (l, rv, DefaultRegMode);
	RETURN lt;
     END;
     -- -----------------------------------------------------------------------------
     FUNCTION  "<" ( CONSTANT l  : INTEGER   ;
		     CONSTANT r  : std_logic_vector 
		   ) RETURN BOOLEAN IS
        VARIABLE lt  : boolean;
	VARIABLE lv  : std_logic_vector (IntegerBitLength - 1 downto 0);
     BEGIN
        -- Convert to bit_vector for comparison to allow any length input vector.
	lv := To_StdLogicVector (l, IntegerBitLength, DefaultRegMode);
	-- Use RegLessThan with DefaultRegMode mode
	lt := RegLessThan (lv, r, DefaultRegMode);
	RETURN lt;
     END;
     -------------------------------------------------------------------------------
     FUNCTION  "<" ( CONSTANT l  : std_logic_vector;
		     CONSTANT r  : INTEGER
		   ) RETURN std_ulogic IS
        VARIABLE lt   : std_ulogic;
	VARIABLE rv  : std_logic_vector (IntegerBitLength - 1 downto 0);
     BEGIN
        -- Convert to bit_vector for comparison to allow any length input vector.
	rv := To_StdLogicVector (r, IntegerBitLength, DefaultRegMode);
	-- Use RegLessThan with DefaultRegMode mode
	lt := RegLessThan (l, rv, DefaultRegMode);
	RETURN lt;
     END;
     -- -----------------------------------------------------------------------------
     FUNCTION  "<" ( CONSTANT l  : INTEGER   ;
		     CONSTANT r  : std_logic_vector 
		   ) RETURN std_ulogic IS
        VARIABLE lt : std_ulogic;
	VARIABLE lv  : std_logic_vector (IntegerBitLength - 1 downto 0);
     BEGIN
        -- Convert to bit_vector for comparison to allow any length input vector.
	lv := To_StdLogicVector (l, IntegerBitLength, DefaultRegMode);
	-- Use RegLessThan with DefaultRegMode mode
	lt := RegLessThan (lv, r, DefaultRegMode);
	RETURN lt;
     END;
     -------------------------------------------------------------------------------
     --     Function Name : Overloaded "<" operator
     --
     --     Purpose       : Less-than relational operator for std_logic_vectors.
     --
     --     Parameters    :     result         left       right
     --                        std_ulogic  std_ulogic_vector   std_ulogic_vector
     --                        BOOLEAN     INTEGER            std_ulogic_vector
     --                        BOOLEAN     std_ulogic_vector   INTEGER
     --                        std_ulogic  INTEGER            std_ulogic_vector
     --                        std_ulogic  std_ulogic_vector   INTEGER  
     --
     --     NOTE          : The std_ulogic_vector operands are assumed to be 
     --                     in  DefaultRegMode. If not they will be converted
     --                     to DefaultRegMode.
     --                     These vectors may be of any length.
     --
     --     Use           :
     --                      VARIABLE a : std_ulogic_vector ( 7 DOWNTO 0 ) := X"FF";
     --                      VARIABLE b : INTEGER;
     --                      IF ( a < b )  THEN
     --
     --     See Also      :   RegLessThan, RegGreaterThan,
     -------------------------------------------------------------------------------
     FUNCTION  "<" ( CONSTANT l  : std_ulogic_vector;
		     CONSTANT r  : std_ulogic_vector
		   ) RETURN std_ulogic IS
       VARIABLE lt : std_ulogic;
     BEGIN
	-- Use RegLessThan with DefaultRegMode mode
	lt := RegLessThan (l,r, DefaultRegMode);
	return lt;
     END;
     -------------------------------------------------------------------------------
     FUNCTION  "<" ( CONSTANT l  : std_ulogic_vector;
		     CONSTANT r  : INTEGER
		   ) RETURN BOOLEAN IS
        VARIABLE lt  : boolean;
	VARIABLE rv  : std_ulogic_vector (IntegerBitLength - 1 downto 0);
     BEGIN
        -- Convert to bit_vector for comparison to allow any length input vector.
	rv := To_StdULogicVector (r, IntegerBitLength, DefaultRegMode);
	-- Use RegLessThan with DefaultRegMode mode
	lt := RegLessThan (l, rv, DefaultRegMode);
	RETURN lt;
     END;
     -- -----------------------------------------------------------------------------
     FUNCTION  "<" ( CONSTANT l  : INTEGER   ;
		     CONSTANT r  : std_ulogic_vector 
		   ) RETURN BOOLEAN IS
        VARIABLE lt  : boolean;
	VARIABLE lv  : std_ulogic_vector (IntegerBitLength - 1 downto 0);
     BEGIN
        -- Convert to bit_vector for comparison to allow any length input vector.
	lv := To_StdULogicVector (l, IntegerBitLength, DefaultRegMode);
	-- Use RegLessThan with DefaultRegMode mode
	lt := RegLessThan (lv, r, DefaultRegMode);
	RETURN lt;
     END;
     -------------------------------------------------------------------------------
     FUNCTION  "<" ( CONSTANT l  : std_ulogic_vector;
		     CONSTANT r  : INTEGER
		   ) RETURN std_ulogic IS
       VARIABLE lt   : std_ulogic;
	VARIABLE rv  : std_ulogic_vector (IntegerBitLength - 1 downto 0);
     BEGIN
        -- Convert to bit_vector for comparison to allow any length input vector.
	rv := To_StdULogicVector (r, IntegerBitLength, DefaultRegMode);
	-- Use RegLessThan with DefaultRegMode mode
	lt := RegLessThan (l, rv, DefaultRegMode);
	RETURN lt;
     END;
     -- -----------------------------------------------------------------------------
     FUNCTION  "<" ( CONSTANT l  : INTEGER   ;
		     CONSTANT r  : std_ulogic_vector 
		   ) RETURN std_ulogic IS
        VARIABLE lt : std_ulogic;
	VARIABLE lv  : std_ulogic_vector (IntegerBitLength - 1 downto 0);
     BEGIN
        -- Convert to bit_vector for comparison to allow any length input vector.
	lv := To_StdULogicVector (l, IntegerBitLength, DefaultRegMode);
	-- Use RegLessThan with DefaultRegMode mode
	lt := RegLessThan (lv, r, DefaultRegMode);
	RETURN lt;
     END;
     -------------------------------------------------------------------------------
     --     Function Name : Overloaded "<=" operator
     -- 1.2.26 and 1.2.28     
     --     Purpose       : Less-than-or-equal relational operator for bit_vectors.
     --     
     --     Parameters    :     result         left       right
     --                        BOOLEAN       INTEGER    bit_vector
     --                        BOOLEAN      bit_vector   INTEGER
     --     
     --     NOTE          : The bit_vector operands are assumed to be 
     --                     in  DefaultRegMode. If not they will be converted
     --                     to DefaultRegMode.
     --                     These vectors may be of any length.
     --
     --     Use           :
     --                      VARIABLE a : bit_vector ( 7 DOWNTO 0 ) := X"FF";
     --                      VARIABLE b : INTEGER;
     --                      IF ( a <= b )  THEN 
     --     
     --     See Also      :   RegLessThan, RegGreaterThan,
     -------------------------------------------------------------------------------
     FUNCTION  "<=" ( CONSTANT l  : bit_vector;
		     CONSTANT r  : bit_vector
		   ) RETURN bit IS
       VARIABLE leq : bit;
     BEGIN
	-- Use RegLessThanOrEqual with DefaultRegMode mode
	leq := RegLessThanOrEqual (l,r, DefaultRegMode);
	return leq;
     END;
     -------------------------------------------------------------------------------
     FUNCTION  "<=" ( CONSTANT l  : bit_vector;
		     CONSTANT r  : INTEGER
		   ) RETURN BOOLEAN IS
        VARIABLE leq  : Boolean;
	VARIABLE rv  : bit_vector (IntegerBitLength - 1 downto 0);
     BEGIN
        -- Convert to bit_vector for comparison to allow any length input vector.
	rv := To_BitVector (r, IntegerBitLength, DefaultRegMode);
	-- Use RegLessThanOrEqual with DefaultRegMode mode
	leq := RegLessThanOrEqual (l, rv , DefaultRegMode);
	return leq;
     END;
     -- -----------------------------------------------------------------------------
     FUNCTION  "<=" ( CONSTANT l  : INTEGER   ;
		     CONSTANT r  : bit_vector 
		   ) RETURN BOOLEAN IS
        VARIABLE leq    : boolean;
	VARIABLE lv  : bit_vector (IntegerBitLength - 1 downto 0);
     BEGIN
        -- Convert to bit_vector for comparison to allow any length input vector.
	lv := To_BitVector (l, IntegerBitLength, DefaultRegMode);
	-- Use RegLessThanOrEqual with DefaultRegMode mode
	leq := RegLessThanOrEqual (lv, r, DefaultRegMode);
	return leq;
     END;
     -------------------------------------------------------------------------------
     FUNCTION  "<=" ( CONSTANT l  : bit_vector;
		     CONSTANT r  : INTEGER
		   ) RETURN bit IS
       VARIABLE leq : bit;
	VARIABLE rv  : bit_vector (IntegerBitLength - 1 downto 0);
     BEGIN
        -- Convert to bit_vector for comparison to allow any length input vector.
	rv := To_BitVector (r, IntegerBitLength, DefaultRegMode);
	-- Use RegLessThanOrEqual with DefaultRegMode mode
	leq := RegLessThanOrEqual (l, rv, DefaultRegMode);
	return leq;
     END;
     -- -----------------------------------------------------------------------------
     FUNCTION  "<=" ( CONSTANT l  : INTEGER   ;
		     CONSTANT r  : bit_vector 
		   ) RETURN bit IS
        VARIABLE leq  : bit;
	VARIABLE lv  : bit_vector (IntegerBitLength - 1 downto 0);
     BEGIN
        -- Convert to bit_vector for comparison to allow any length input vector.
	lv := To_BitVector (l, IntegerBitLength, DefaultRegMode);
	-- Use RegLessThanOrEqual with DefaultRegMode mode
	leq := RegLessThanOrEqual (lv, r, DefaultRegMode);
	return leq;
     END;
     -------------------------------------------------------------------------------
     --     Function Name : Overloaded "<=" operator
     --
     --     Purpose       : Less-than-or-equal relational operator for std_logic_vectors.
     --
     --     Parameters    :     result         left       right
     --                        std_ulogic  std_logic_vector   std_logic_vector
     --                        BOOLEAN     INTEGER            std_logic_vector
     --                        BOOLEAN     std_logic_vector   INTEGER
     --                        std_ulogic  INTEGER            std_logic_vector
     --                        std_ulogic  std_logic_vector   INTEGER
     --
     --     NOTE          : The std_logic_vector operands are assumed to be 
     --                     in  DefaultRegMode. If not they will be converted
     --                     to DefaultRegMode.
     --                     These vectors may be of any length.
     --
     --     Use           :
     --                      VARIABLE a : std_logic_vector ( 7 DOWNTO 0 ) := X"FF";
     --                      VARIABLE b : INTEGER;
     --                      IF ( a <= b )  THEN
     --
     --     See Also      :   RegLessThanOrEqual, RegGreaterThan,
     -------------------------------------------------------------------------------
     FUNCTION  "<=" ( CONSTANT l  : std_logic_vector;
		     CONSTANT r  : std_logic_vector
		   ) RETURN std_ulogic IS
       VARIABLE leq : std_ulogic;
     BEGIN
	-- Use RegLessThanOrEqual with DefaultRegMode mode
	leq := RegLessThanOrEqual (l,r, DefaultRegMode);
	return leq;
     END;
     -------------------------------------------------------------------------------
     FUNCTION  "<=" ( CONSTANT l  : std_logic_vector;
		     CONSTANT r  : INTEGER
		   ) RETURN BOOLEAN IS
        VARIABLE leq  : boolean;
	VARIABLE rv  : std_logic_vector (IntegerBitLength - 1 downto 0);
     BEGIN
        -- Convert to bit_vector for comparison to allow any length input vector.
	rv := To_StdLogicVector (r, IntegerBitLength, DefaultRegMode);
	-- Use RegLessThanOrEqual with DefaultRegMode mode
	leq := RegLessThanOrEqual (l, rv, DefaultRegMode);
	RETURN leq;
     END;
     -- -----------------------------------------------------------------------------
     FUNCTION  "<=" ( CONSTANT l  : INTEGER   ;
		     CONSTANT r  : std_logic_vector 
		   ) RETURN BOOLEAN IS
        VARIABLE leq  : boolean;
	VARIABLE lv  : std_logic_vector (IntegerBitLength - 1 downto 0);
     BEGIN
        -- Convert to bit_vector for comparison to allow any length input vector.
	lv := To_StdLogicVector (l, IntegerBitLength, DefaultRegMode);
	-- Use RegLessThanOrEqual with DefaultRegMode mode
	leq := RegLessThanOrEqual (lv, r, DefaultRegMode);
	RETURN leq;
     END;
     -------------------------------------------------------------------------------
     FUNCTION  "<=" ( CONSTANT l  : std_logic_vector;
		     CONSTANT r  : INTEGER
		   ) RETURN std_ulogic IS
        VARIABLE leq   : std_ulogic;
	VARIABLE rv  : std_logic_vector (IntegerBitLength - 1 downto 0);
     BEGIN
        -- Convert to bit_vector for comparison to allow any length input vector.
	rv := To_StdLogicVector (r, IntegerBitLength, DefaultRegMode);
	-- Use RegLessThanOrEqual with DefaultRegMode mode
	leq := RegLessThanOrEqual (l, rv, DefaultRegMode);
	RETURN leq;
     END;
     -- -----------------------------------------------------------------------------
     FUNCTION  "<=" ( CONSTANT l  : INTEGER   ;
		     CONSTANT r  : std_logic_vector 
		   ) RETURN std_ulogic IS
        VARIABLE leq : std_ulogic;
	VARIABLE lv  : std_logic_vector (IntegerBitLength - 1 downto 0);
     BEGIN
        -- Convert to bit_vector for comparison to allow any length input vector.
	lv := To_StdLogicVector (l, IntegerBitLength, DefaultRegMode);
	-- Use RegLessThanOrEqual with DefaultRegMode mode
	leq := RegLessThanOrEqual (lv, r, DefaultRegMode);
	RETURN leq;
     END;
     -------------------------------------------------------------------------------
     --     Function Name : Overloaded "<=" operator
     --
     --     Purpose       : Less-than-or-equal relational operator for std_logic_vectors.
     --
     --     Parameters    :     result         left       right
     --                        std_ulogic  std_ulogic_vector   std_ulogic_vector
     --                        BOOLEAN     INTEGER            std_ulogic_vector
     --                        BOOLEAN     std_ulogic_vector   INTEGER
     --                        std_ulogic  INTEGER            std_ulogic_vector
     --                        std_ulogic  std_ulogic_vector   INTEGER  
     --
     --     NOTE          : The std_ulogic_vector operands are assumed to be 
     --                     in  DefaultRegMode. If not they will be converted
     --                     to DefaultRegMode.
     --                     These vectors may be of any length.
     --
     --     Use           :
     --                      VARIABLE a : std_ulogic_vector ( 7 DOWNTO 0 ) := X"FF";
     --                      VARIABLE b : INTEGER;
     --                      IF ( a <= b )  THEN
     --
     --     See Also      :   RegLessThanOrEqual, RegGreaterThan,
     -------------------------------------------------------------------------------
     FUNCTION  "<=" ( CONSTANT l  : std_ulogic_vector;
		     CONSTANT r  : std_ulogic_vector
		   ) RETURN std_ulogic IS
       VARIABLE leq : std_ulogic;
     BEGIN
	-- Use RegLessThanOrEqual with DefaultRegMode mode
	leq := RegLessThanOrEqual (l,r, DefaultRegMode);
	return leq;
     END;
     -------------------------------------------------------------------------------
     FUNCTION  "<=" ( CONSTANT l  : std_ulogic_vector;
		     CONSTANT r  : INTEGER
		   ) RETURN BOOLEAN IS
        VARIABLE leq  : boolean;
	VARIABLE rv  : std_ulogic_vector (IntegerBitLength - 1 downto 0);
     BEGIN
        -- Convert to bit_vector for comparison to allow any length input vector.
	rv := To_StdULogicVector (r, IntegerBitLength, DefaultRegMode);
	-- Use RegLessThanOrEqual with DefaultRegMode mode
	leq := RegLessThanOrEqual (l, rv, DefaultRegMode);
	RETURN leq;
     END;
     -- -----------------------------------------------------------------------------
     FUNCTION  "<=" ( CONSTANT l  : INTEGER   ;
		     CONSTANT r  : std_ulogic_vector 
		   ) RETURN BOOLEAN IS
        VARIABLE leq  : boolean;
	VARIABLE lv  : std_ulogic_vector (IntegerBitLength - 1 downto 0);
     BEGIN
        -- Convert to bit_vector for comparison to allow any length input vector.
	lv := To_StdULogicVector (l, IntegerBitLength, DefaultRegMode);
	-- Use RegLessThanOrEqual with DefaultRegMode mode
	leq := RegLessThanOrEqual (lv, r, DefaultRegMode);
	RETURN leq;
     END;
     -------------------------------------------------------------------------------
     FUNCTION  "<=" ( CONSTANT l  : std_ulogic_vector;
		     CONSTANT r  : INTEGER
		   ) RETURN std_ulogic IS
       VARIABLE leq   : std_ulogic;
	VARIABLE rv  : std_ulogic_vector (IntegerBitLength - 1 downto 0);
     BEGIN
        -- Convert to bit_vector for comparison to allow any length input vector.
	rv := To_StdULogicVector (r, IntegerBitLength, DefaultRegMode);
	-- Use RegLessThanOrEqual with DefaultRegMode mode
	leq := RegLessThanOrEqual (l, rv, DefaultRegMode);
	RETURN leq;
     END;
     -- -----------------------------------------------------------------------------
     FUNCTION  "<=" ( CONSTANT l  : INTEGER   ;
		     CONSTANT r  : std_ulogic_vector 
		   ) RETURN std_ulogic IS
        VARIABLE leq : std_ulogic;
	VARIABLE lv  : std_ulogic_vector (IntegerBitLength - 1 downto 0);
     BEGIN
        -- Convert to bit_vector for comparison to allow any length input vector.
	lv := To_StdULogicVector (l, IntegerBitLength, DefaultRegMode);
	-- Use RegLessThanOrEqual with DefaultRegMode mode
	leq := RegLessThanOrEqual (lv, r, DefaultRegMode);
	RETURN leq;
     END;

     --------------------------------------------------------------------------------
     --     Function Name : Overloaded ">" operator
     -- 1.2.18 and 1.2.20     
     --     Purpose       : Greater-than relational operator for bit_vectors.
     --     
     --     Parameters    :     result         left       right
     --                        BOOLEAN       INTEGER    bit_vector
     --                        BOOLEAN      bit_vector   INTEGER
     --     
     --     NOTE          : The bit_vector operands are assumed to be 
     --                     in  DefaultRegMode. If not they will be converted
     --                     to DefaultRegMode.
     --                     These vectors may be of any length.
     --
     --     Use           :
     --                      VARIABLE a : bit_vector ( 7 DOWNTO 0 ) := X"FF";
     --                      VARIABLE b : INTEGER;
     --                      IF ( a > b )  THEN 
     --     
     --     See Also      :   RegGreaterThan, RegGreaterThan,
     -------------------------------------------------------------------------------
     FUNCTION  ">" ( CONSTANT l  : bit_vector;
		     CONSTANT r  : bit_vector
		   ) RETURN bit IS
	VARIABLE gt : BIT;    
     BEGIN
	-- Use RegGreaterThan with DefaultRegMode mode
	gt := RegGreaterThan (l,r, DefaultRegMode);
	return gt;
     END;
     -------------------------------------------------------------------------------
     FUNCTION  ">" ( CONSTANT l  : bit_vector;
		     CONSTANT r  : INTEGER
		   ) RETURN BOOLEAN IS
        VARIABLE gt  : Boolean;
	VARIABLE rv  : bit_vector (IntegerBitLength - 1 downto 0);
     BEGIN
        -- Convert to bit_vector for comparison to allow any length input vector.
	rv := To_BitVector (r, IntegerBitLength, DefaultRegMode);
	-- Use RegGreaterThan with DefaultRegMode mode
	gt := RegGreaterThan (l, rv , DefaultRegMode);
	return gt;
     END;
     -- -----------------------------------------------------------------------------
     FUNCTION  ">" ( CONSTANT l  : INTEGER   ;
		     CONSTANT r  : bit_vector 
		   ) RETURN BOOLEAN IS
        VARIABLE gt    : boolean;
	VARIABLE lv  : bit_vector (IntegerBitLength - 1 downto 0);
     BEGIN
        -- Convert to bit_vector for comparison to allow any length input vector.
	lv := To_BitVector (l, IntegerBitLength, DefaultRegMode);
	-- Use RegGreaterThan with DefaultRegMode mode
	gt := RegGreaterThan (lv, r, DefaultRegMode);
	return gt;
     END;
     -------------------------------------------------------------------------------
     FUNCTION  ">" ( CONSTANT l  : bit_vector;
		     CONSTANT r  : INTEGER
		   ) RETURN bit IS
       VARIABLE gt : bit;
	VARIABLE rv  : bit_vector (IntegerBitLength - 1 downto 0);
     BEGIN
        -- Convert to bit_vector for comparison to allow any length input vector.
	rv := To_BitVector (r, IntegerBitLength, DefaultRegMode);
	-- Use RegGreaterThan with DefaultRegMode mode
	gt := RegGreaterThan (l, rv, DefaultRegMode);
	return gt;
     END;
     -- -----------------------------------------------------------------------------
     FUNCTION  ">" ( CONSTANT l  : INTEGER   ;
		     CONSTANT r  : bit_vector 
		   ) RETURN bit IS
        VARIABLE gt  : bit;
	VARIABLE lv  : bit_vector (IntegerBitLength - 1 downto 0);
     BEGIN
        -- Convert to bit_vector for comparison to allow any length input vector.
	lv := To_BitVector (l, IntegerBitLength, DefaultRegMode);
	-- Use RegGreaterThan with DefaultRegMode mode
	gt := RegGreaterThan (lv, r, DefaultRegMode);
	return gt;
     END;
     -------------------------------------------------------------------------------
     --     Function Name : Overloaded ">" operator
     --
     --     Purpose       : Greater-than relational operator for std_logic_vectors.
     --
     --     Parameters    :     result         left       right
     --                        std_ulogic  std_logic_vector   std_logic_vector
     --                        BOOLEAN     INTEGER            std_logic_vector
     --                        BOOLEAN     std_logic_vector   INTEGER
     --                        std_ulogic  INTEGER            std_logic_vector
     --                        std_ulogic  std_logic_vector   INTEGER
     --
     --     NOTE          : The std_logic_vector operands are assumed to be 
     --                     in  DefaultRegMode. If not they will be converted
     --                     to DefaultRegMode.
     --                     These vectors may be of any length.
     --
     --     Use           :
     --                      VARIABLE a : std_logic_vector ( 7 DOWNTO 0 ) := X"FF";
     --                      VARIABLE b : INTEGER;
     --                      IF ( a > b )  THEN
     --
     --     See Also      :   RegLessThan, RegGreaterThan,
     -------------------------------------------------------------------------------
     FUNCTION  ">" ( CONSTANT l  : std_logic_vector;
		     CONSTANT r  : std_logic_vector
		   ) RETURN std_ulogic IS
       VARIABLE gt : std_ulogic;
     BEGIN
	-- Use RegGreaterThan with DefaugtRegMode mode
	gt := RegGreaterThan (l,r, DefaultRegMode);
	return gt;
     END;
     -------------------------------------------------------------------------------
     FUNCTION  ">" ( CONSTANT l  : std_logic_vector;
		     CONSTANT r  : INTEGER
		   ) RETURN BOOLEAN IS
        VARIABLE gt  : boolean;
	VARIABLE rv  : std_logic_vector (IntegerBitLength - 1 downto 0);
     BEGIN
        -- Convert to bit_vector for comparison to allow any length input vector.
	rv := To_StdLogicVector (r, IntegerBitLength, DefaultRegMode);
	-- Use RegGreaterThan with DefaultRegMode mode
	gt := RegGreaterThan (l, rv, DefaultRegMode);
	RETURN gt;
     END;
     -- -----------------------------------------------------------------------------
     FUNCTION  ">" ( CONSTANT l  : INTEGER   ;
		     CONSTANT r  : std_logic_vector 
		   ) RETURN BOOLEAN IS
        VARIABLE gt  : boolean;
	VARIABLE lv  : std_logic_vector (IntegerBitLength - 1 downto 0);
     BEGIN
        -- Convert to bit_vector for comparison to allow any length input vector.
	lv := To_StdLogicVector (l, IntegerBitLength, DefaultRegMode);
	-- Use RegGreaterThan with DefaultRegMode mode
	gt := RegGreaterThan (lv, r, DefaultRegMode);
	RETURN gt;
     END;
     -------------------------------------------------------------------------------
     FUNCTION  ">" ( CONSTANT l  : std_logic_vector;
		     CONSTANT r  : INTEGER
		   ) RETURN std_ulogic IS
        VARIABLE gt   : std_ulogic;
	VARIABLE rv  : std_logic_vector (IntegerBitLength - 1 downto 0);
     BEGIN
        -- Convert to bit_vector for comparison to allow any length input vector.
	rv := To_StdLogicVector (r, IntegerBitLength, DefaultRegMode);
	-- Use RegGreaterThan with DefaultRegMode mode
	gt := RegGreaterThan (l, rv, DefaultRegMode);
	RETURN gt;
     END;
     -- -----------------------------------------------------------------------------
     FUNCTION  ">" ( CONSTANT l  : INTEGER   ;
		     CONSTANT r  : std_logic_vector 
		   ) RETURN std_ulogic IS
        VARIABLE gt : std_ulogic;
	VARIABLE lv  : std_logic_vector (IntegerBitLength - 1 downto 0);
     BEGIN
        -- Convert to bit_vector for comparison to allow any length input vector.
	lv := To_StdLogicVector (l, IntegerBitLength, DefaultRegMode);
	-- Use RegGreaterThan with DefaultRegMode mode
	gt := RegGreaterThan (lv, r, DefaultRegMode);
	RETURN gt;
     END;
     -------------------------------------------------------------------------------
     --     Function Name : Overloaded ">" operator
     --
     --     Purpose       : Greater-than relational operator for std_logic_vectors.
     --
     --     Parameters    :     result         left       right
     --                        std_ulogic  std_ulogic_vector   std_ulogic_vector
     --                        BOOLEAN     INTEGER            std_ulogic_vector
     --                        BOOLEAN     std_ulogic_vector   INTEGER
     --                        std_ulogic  INTEGER            std_ulogic_vector
     --                        std_ulogic  std_ulogic_vector   INTEGER  
     --
     --     NOTE          : The std_ulogic_vector operands are assumed to be 
     --                     in  DefaultRegMode. If not they will be converted
     --                     to DefaultRegMode.
     --                     These vectors may be of any length.
     --
     --     Use           :
     --                      VARIABLE a : std_ulogic_vector ( 7 DOWNTO 0 ) := X"FF";
     --                      VARIABLE b : INTEGER;
     --                      IF ( a > b )  THEN
     --
     --     See Also      :   RegLessThan, RegGreaterThan,
     -------------------------------------------------------------------------------
     FUNCTION  ">" ( CONSTANT l  : std_ulogic_vector;
		     CONSTANT r  : std_ulogic_vector
		   ) RETURN std_ulogic IS
       VARIABLE gt : std_ulogic;
     BEGIN
	-- Use RegGreaterThan with DefaultRegMode mode
	gt := RegGreaterThan (l,r, DefaultRegMode);
	return gt;
     END;
     -------------------------------------------------------------------------------
     FUNCTION  ">" ( CONSTANT l  : std_ulogic_vector;
		     CONSTANT r  : INTEGER
		   ) RETURN BOOLEAN IS
        VARIABLE gt  : boolean;
	VARIABLE rv  : std_ulogic_vector (IntegerBitLength - 1 downto 0);
     BEGIN
        -- Convert to bit_vector for comparison to allow any length input vector.
	rv := To_StdULogicVector (r, IntegerBitLength, DefaultRegMode);
	-- Use RegGreaterThan with DefaultRegMode mode
	gt := RegGreaterThan (l, rv, DefaultRegMode);
	RETURN gt;
     END;
     -- -----------------------------------------------------------------------------
     FUNCTION  ">" ( CONSTANT l  : INTEGER   ;
		     CONSTANT r  : std_ulogic_vector 
		   ) RETURN BOOLEAN IS
        VARIABLE gt  : boolean;
	VARIABLE lv  : std_ulogic_vector (IntegerBitLength - 1 downto 0);
     BEGIN
        -- Convert to bit_vector for comparison to allow any length input vector.
	lv := To_StdULogicVector (l, IntegerBitLength, DefaultRegMode);
	-- Use RegGreaterThan with DefaultRegMode mode
	gt := RegGreaterThan (lv, r, DefaultRegMode);
	RETURN gt;
     END;
     -------------------------------------------------------------------------------
     FUNCTION  ">" ( CONSTANT l  : std_ulogic_vector;
		     CONSTANT r  : INTEGER
		   ) RETURN std_ulogic IS
       VARIABLE gt   : std_ulogic;
	VARIABLE rv  : std_ulogic_vector (IntegerBitLength - 1 downto 0);
     BEGIN
        -- Convert to bit_vector for comparison to allow any length input vector.
	rv := To_StdULogicVector (r, IntegerBitLength, DefaultRegMode);
	-- Use RegGreaterThan with DefaultRegMode mode
	gt := RegGreaterThan (l, rv, DefaultRegMode);
	RETURN gt;
     END;
     -- -----------------------------------------------------------------------------
     FUNCTION  ">" ( CONSTANT l  : INTEGER   ;
		     CONSTANT r  : std_ulogic_vector 
		   ) RETURN std_ulogic IS
        VARIABLE gt : std_ulogic;
	VARIABLE lv  : std_ulogic_vector (IntegerBitLength - 1 downto 0);
     BEGIN
        -- Convert to bit_vector for comparison to allow any length input vector.
	lv := To_StdULogicVector (l, IntegerBitLength, DefaultRegMode);
	-- Use RegGreaterThan with DefaultRegMode mode
	gt := RegGreaterThan (lv, r, DefaultRegMode);
	RETURN gt;
     END;
     -------------------------------------------------------------------------------
     --     Function Name : Overloaded ">=" operator
     -- 1.2.26 and 1.2.28     
     --     Purpose       : Greater-than-or-equal relational operator for bit_vectors.
     --     
     --     Parameters    :     result         left       right
     --                        BOOLEAN       INTEGER    bit_vector
     --                        BOOLEAN      bit_vector   INTEGER
     --     
     --     NOTE          : The bit_vector operands are assumed to be 
     --                     in  DefaultRegMode. If not they will be converted
     --                     to DefaultRegMode.
     --                     These vectors may be of any length.
     --
     --     Use           :
     --                      VARIABLE a : bit_vector ( 7 DOWNTO 0 ) := X"FF";
     --                      VARIABLE b : INTEGER;
     --                      IF ( a >= b )  THEN 
     --     
     --     See Also      :   RegLessThan, RegGreaterThan,
     -------------------------------------------------------------------------------
     FUNCTION  ">=" ( CONSTANT l  : bit_vector;
		     CONSTANT r  : bit_vector
		   ) RETURN bit IS
       VARIABLE geq : bit;
     BEGIN
	-- Use RegGreaterThanOrEqual with DefaultRegMode mode
	geq := RegGreaterThanOrEqual (l,r, DefaultRegMode);
	return geq;
     END;
     -------------------------------------------------------------------------------
     FUNCTION  ">=" ( CONSTANT l  : bit_vector;
		     CONSTANT r  : INTEGER
		   ) RETURN BOOLEAN IS
        VARIABLE geq  : Boolean;
	VARIABLE rv  : bit_vector (IntegerBitLength - 1 downto 0);
     BEGIN
        -- Convert to bit_vector for comparison to allow any length input vector.
	rv := To_BitVector (r, IntegerBitLength, DefaultRegMode);
	-- Use RegGreaterThanOrEqual with DefaultRegMode mode
	geq := RegGreaterThanOrEqual (l, rv , DefaultRegMode);
	return geq;
     END;
     -- -----------------------------------------------------------------------------
     FUNCTION  ">=" ( CONSTANT l  : INTEGER   ;
		     CONSTANT r  : bit_vector 
		   ) RETURN BOOLEAN IS
        VARIABLE geq    : boolean;
	VARIABLE lv  : bit_vector (IntegerBitLength - 1 downto 0);
     BEGIN
        -- Convert to bit_vector for comparison to allow any length input vector.
	lv := To_BitVector (l, IntegerBitLength, DefaultRegMode);
	-- Use RegGreaterThanOrEqual with DefaultRegMode mode
	geq := RegGreaterThanOrEqual (lv, r, DefaultRegMode);
	return geq;
     END;
     -------------------------------------------------------------------------------
     FUNCTION  ">=" ( CONSTANT l  : bit_vector;
		     CONSTANT r  : INTEGER
		   ) RETURN bit IS
       VARIABLE geq : bit;
	VARIABLE rv  : bit_vector (IntegerBitLength - 1 downto 0);
     BEGIN
        -- Convert to bit_vector for comparison to allow any length input vector.
	rv := To_BitVector (r, IntegerBitLength, DefaultRegMode);
	-- Use RegGreaterThanOrEqual with DefaultRegMode mode
	geq := RegGreaterThanOrEqual (l, rv, DefaultRegMode);
	return geq;
     END;
     -- -----------------------------------------------------------------------------
     FUNCTION  ">=" ( CONSTANT l  : INTEGER   ;
		     CONSTANT r  : bit_vector 
		   ) RETURN bit IS
        VARIABLE geq  : bit;
	VARIABLE lv  : bit_vector (IntegerBitLength - 1 downto 0);
     BEGIN
        -- Convert to bit_vector for comparison to allow any length input vector.
	lv := To_BitVector (l, IntegerBitLength, DefaultRegMode);
	-- Use RegGreaterThanOrEqual with DefaultRegMode mode
	geq := RegGreaterThanOrEqual (lv, r, DefaultRegMode);
	return geq;
     END;
     -------------------------------------------------------------------------------
     --     Function Name : Overloaded ">=" operator
     --
     --     Purpose       : Greater-than-or-equal relational operator for std_logic_vectors.
     --
     --     Parameters    :     result         left       right
     --                        std_ulogic  std_logic_vector   std_logic_vector
     --                        BOOLEAN     INTEGER            std_logic_vector
     --                        BOOLEAN     std_logic_vector   INTEGER
     --                        std_ulogic  INTEGER            std_logic_vector
     --                        std_ulogic  std_logic_vector   INTEGER
     --
     --     NOTE          : The std_logic_vector operands are assumed to be 
     --                     in  DefaultRegMode. If not they will be converted
     --                     to DefaultRegMode.
     --                     These vectors may be of any length.
     --
     --     Use           :
     --                      VARIABLE a : std_logic_vector ( 7 DOWNTO 0 ) := X"FF";
     --                      VARIABLE b : INTEGER;
     --                      IF ( a >= b )  THEN
     --
     --     See Also      :   RegLessThanOrEqual, RegGreaterThan,
     -------------------------------------------------------------------------------
     FUNCTION  ">=" ( CONSTANT l  : std_logic_vector;
		     CONSTANT r  : std_logic_vector
		   ) RETURN std_ulogic IS
       VARIABLE geq : std_ulogic;
     BEGIN
	-- Use RegGreaterThanOrEqual with DefaultRegMode mode
	geq := RegGreaterThanOrEqual (l,r, DefaultRegMode);
	return geq;
     END;
     -------------------------------------------------------------------------------
     FUNCTION  ">=" ( CONSTANT l  : std_logic_vector;
		     CONSTANT r  : INTEGER
		   ) RETURN BOOLEAN IS
        VARIABLE geq  : boolean;
	VARIABLE rv  : std_logic_vector (IntegerBitLength - 1 downto 0);
     BEGIN
        -- Convert to bit_vector for comparison to allow any length input vector.
	rv := To_StdLogicVector (r, IntegerBitLength, DefaultRegMode);
	-- Use RegGreaterThanOrEqual with DefaultRegMode mode
	geq := RegGreaterThanOrEqual (l, rv, DefaultRegMode);
	RETURN geq;
     END;
     -- -----------------------------------------------------------------------------
     FUNCTION  ">=" ( CONSTANT l  : INTEGER   ;
		     CONSTANT r  : std_logic_vector 
		   ) RETURN BOOLEAN IS
        VARIABLE geq  : boolean;
	VARIABLE lv  : std_logic_vector (IntegerBitLength - 1 downto 0);
     BEGIN
        -- Convert to bit_vector for comparison to allow any length input vector.
	lv := To_StdLogicVector (l, IntegerBitLength, DefaultRegMode);
	-- Use RegGreaterThanOrEqual with DefaultRegMode mode
	geq := RegGreaterThanOrEqual (lv, r, DefaultRegMode);
	RETURN geq;
     END;
     -------------------------------------------------------------------------------
     FUNCTION  ">=" ( CONSTANT l  : std_logic_vector;
		     CONSTANT r  : INTEGER
		   ) RETURN std_ulogic IS
        VARIABLE geq   : std_ulogic;
	VARIABLE rv  : std_logic_vector (IntegerBitLength - 1 downto 0);
     BEGIN
        -- Convert to bit_vector for comparison to allow any length input vector.
	rv := To_StdLogicVector (r, IntegerBitLength, DefaultRegMode);
	-- Use RegGreaterThanOrEqual with DefaultRegMode mode
	geq := RegGreaterThanOrEqual (l, rv, DefaultRegMode);
	RETURN geq;
     END;
     -- -----------------------------------------------------------------------------
     FUNCTION  ">=" ( CONSTANT l  : INTEGER   ;
		     CONSTANT r  : std_logic_vector 
		   ) RETURN std_ulogic IS
        VARIABLE geq : std_ulogic;
	VARIABLE lv  : std_logic_vector (IntegerBitLength - 1 downto 0);
     BEGIN
        -- Convert to bit_vector for comparison to allow any length input vector.
	lv := To_StdLogicVector (l, IntegerBitLength, DefaultRegMode);
	-- Use RegGreaterThanOrEqual with DefaultRegMode mode
	geq := RegGreaterThanOrEqual (lv, r, DefaultRegMode);
	RETURN geq;
     END;
     -------------------------------------------------------------------------------
     --     Function Name : Overloaded ">=" operator
     --
     --     Purpose       : Greater-than-or-equal relational operator for std_logic_vectors.
     --
     --     Parameters    :     result         left       right
     --                        std_ulogic  std_ulogic_vector   std_ulogic_vector
     --                        BOOLEAN     INTEGER            std_ulogic_vector
     --                        BOOLEAN     std_ulogic_vector   INTEGER
     --                        std_ulogic  INTEGER            std_ulogic_vector
     --                        std_ulogic  std_ulogic_vector   INTEGER  
     --
     --     NOTE          : The std_ulogic_vector operands are assumed to be 
     --                     in  DefaultRegMode. If not they will be converted
     --                     to DefaultRegMode.
     --                     These vectors may be of any length.
     --
     --     Use           :
     --                      VARIABLE a : std_ulogic_vector ( 7 DOWNTO 0 ) := X"FF";
     --                      VARIABLE b : INTEGER;
     --                      IF ( a >= b )  THEN
     --
     --     See Also      :   RegLessThanOrEqual, RegGreaterThan,
     -------------------------------------------------------------------------------
     FUNCTION  ">=" ( CONSTANT l  : std_ulogic_vector;
		     CONSTANT r  : std_ulogic_vector
		   ) RETURN std_ulogic IS
       VARIABLE geq : std_ulogic;
     BEGIN
	-- Use RegGreaterThanOrEqual with DefaultRegMode mode
	geq := RegGreaterThanOrEqual (l,r, DefaultRegMode);
	return geq;
     END;
     -------------------------------------------------------------------------------
     FUNCTION  ">=" ( CONSTANT l  : std_ulogic_vector;
		     CONSTANT r  : INTEGER
		   ) RETURN BOOLEAN IS
        VARIABLE geq  : boolean;
	VARIABLE rv  : std_ulogic_vector (IntegerBitLength - 1 downto 0);
     BEGIN
        -- Convert to bit_vector for comparison to allow any length input vector.
	rv := To_StdULogicVector (r, IntegerBitLength, DefaultRegMode);
	-- Use RegGreaterThanOrEqual with DefaultRegMode mode
	geq := RegGreaterThanOrEqual (l, rv, DefaultRegMode);
	RETURN geq;
     END;
     -- -----------------------------------------------------------------------------
     FUNCTION  ">=" ( CONSTANT l  : INTEGER   ;
		     CONSTANT r  : std_ulogic_vector 
		   ) RETURN BOOLEAN IS
        VARIABLE geq  : boolean;
	VARIABLE lv  : std_ulogic_vector (IntegerBitLength - 1 downto 0);
     BEGIN
        -- Convert to bit_vector for comparison to allow any length input vector.
	lv := To_StdULogicVector (l, IntegerBitLength, DefaultRegMode);
	-- Use RegGreaterThanOrEqual with DefaultRegMode mode
	geq := RegGreaterThanOrEqual (lv, r, DefaultRegMode);
	RETURN geq;
     END;
     -------------------------------------------------------------------------------
     FUNCTION  ">=" ( CONSTANT l  : std_ulogic_vector;
		     CONSTANT r  : INTEGER
		   ) RETURN std_ulogic IS
       VARIABLE geq   : std_ulogic;
	VARIABLE rv  : std_ulogic_vector (IntegerBitLength - 1 downto 0);
     BEGIN
        -- Convert to bit_vector for comparison to allow any length input vector.
	rv := To_StdULogicVector (r, IntegerBitLength, DefaultRegMode);
	-- Use RegGreaterThanOrEqual with DefaultRegMode mode
	geq := RegGreaterThanOrEqual (l, rv, DefaultRegMode);
	RETURN geq;
     END;
     -- -----------------------------------------------------------------------------
     FUNCTION  ">=" ( CONSTANT l  : INTEGER   ;
		     CONSTANT r  : std_ulogic_vector 
		   ) RETURN std_ulogic IS
        VARIABLE geq : std_ulogic;
	VARIABLE lv  : std_ulogic_vector (IntegerBitLength - 1 downto 0);
     BEGIN
        -- Convert to bit_vector for comparison to allow any length input vector.
	lv := To_StdULogicVector (l, IntegerBitLength, DefaultRegMode);
	-- Use RegGreaterThanOrEqual with DefaultRegMode mode
	geq := RegGreaterThanOrEqual (lv, r, DefaultRegMode);
	RETURN geq;
     END;
--+-----------------------------------------------------------------------------
--|     Function Name  : To_TwosComp_FromUnsign
--| 1.8.7
--|     Overloading    : None
--|  
--|     Purpose        : Convert a STD_ULOGIC_VECTOR to Two's Compliment Notation.
--|  
--|     Parameters     :
--|                      ARG     - input  STD_LOGIC_VECTOR, the vector to be read.
--|                      SIZE    - input INTEGER
--|
--|     Result         : STD_LOGIC_VECTOR, the vector in Two's complement notation.
--|
--|
--|     Use            :
--|                      VARIABLE vect : STD_LOGIC_VECTOR ( 15 DOWNTO 0 );
--|                      vect := To_TwosComp_FromUnsign ( "0101", 4); -- set to +5
--|
--|     See Also       : To_BitVector, To_Integer, To_TwosComp
--|-----------------------------------------------------------------------------
    FUNCTION To_TwosComp_FromUnsig  ( CONSTANT ARG      : IN STD_LOGIC_VECTOR;
                                      CONSTANT SIZE     : IN INTEGER
                                    ) RETURN STD_LOGIC_VECTOR IS

	VARIABLE reg_copy  : STD_LOGIC_VECTOR (ARG'LENGTH - 1 DOWNTO 0);
	VARIABLE result    : STD_LOGIC_VECTOR (ARG'LENGTH - 1 DOWNTO 0);
	-- synopsys built_in SYN_ZERO_EXTEND
    BEGIN
	-- synopsys synthesis_off        
       --  Check for null input
        reg_copy := ARG;
        IF (ARG'LENGTH = 0) THEN
            ASSERT false
            REPORT " To_TwosComp --- input register has zero length,  "
	     & " Returning vector with zero length "
            SEVERITY ERROR;
            RETURN reg_copy;

        ELSE
          result := reg_copy;
         -- if MSB is '1' or 'X' then the number is larger than what
         -- could be accommodated in the  register.
           IF (reg_copy(ARG'LENGTH -1) /= '0') THEN
                ASSERT false
                REPORT "To_TwosComp - MSB of unsigned std_logic_vector "
                   & " is not '0'. it cannot be converted "
               SEVERITY Error; 
          END IF;
        END IF;
        RETURN result;
 	-- synopsys synthesis_on
    END To_TwosComp_FromUnsig;

--+-----------------------------------------------------------------------------
--|     Function Name  : To_TwosComp
--| 1.8.7
--|     Overloading    : None
--|  
--|     Purpose        : Convert a STD_LOGIC_VECTOR to Two's Compliment Notation.
--|  
--|     Parameters     :
--|                      SrcReg     - input  STD_LOGIC_VECTOR, the vector to be read.
--|                      SrcRegMode - input  regmode_type, indicating the format of
--|                                the input STD_LOGIC_VECTOR.   Default is TwosComp.
--|
--|     Result         : STD_LOGIC_VECTOR, the vector in Two's complement notation.
--|
--|
--|     Use            :
--|                      VARIABLE vect : STD_LOGIC_VECTOR ( 15 DOWNTO 0 );
--|                      vect := To_TwosComp ( "0101",  UnSigned ); -- set to +5
--|
--|     See Also       : To_BitVector, To_Integer, To_TwosComp
--|-----------------------------------------------------------------------------
    FUNCTION To_TwosComp  ( CONSTANT SrcReg      : IN STD_LOGIC_VECTOR;
                            CONSTANT SrcRegMode  : IN regmode_type
                     -- synopsys synthesis_off
						      := DefaultRegMode 
                     -- synopsys synthesis_on
                          ) RETURN STD_LOGIC_VECTOR IS

    BEGIN
	if (SrcRegMode = Unsigned) THEN
		return (To_TwosComp_FromUnsig(SrcReg, SrcReg'LENGTH));
	else
		return(SrcReg);
	end if;
    END To_TwosComp;
--+-----------------------------------------------------------------------------
--|     Function Name  : To_TwosComp
--| 1.8.7
--|     Overloading    : None
--|  
--|     Purpose        : Convert a STD_ULOGIC_VECTOR to Two's Compliment Notation.
--|  
--|     Parameters     :
--|                      SrcReg     - input  STD_ULOGIC_VECTOR, the vector to be read.
--|                      SrcRegMode - input  regmode_type, indicating the format of
--|                                the input STD_ULOGIC_VECTOR.   Default is TwosComp.
--|
--|     Result         : STD_ULOGIC_VECTOR, the vector in Two's complement notation.
--|
--|
--|     Use            :
--|                      VARIABLE vect : STD_ULOGIC_VECTOR ( 15 DOWNTO 0 );
--|                      vect := To_TwosComp ( "0101",  UnSigned ); -- set to +5
--|
--|     See Also       : To_BitVector, To_Integer, To_TwosComp
--|-----------------------------------------------------------------------------
    FUNCTION To_TwosComp  ( CONSTANT SrcReg      : IN STD_ULOGIC_VECTOR;
                            CONSTANT SrcRegMode  : IN regmode_type
                     -- synopsys synthesis_off
						      := DefaultRegMode 
                     -- synopsys synthesis_on
                          ) RETURN STD_ULOGIC_VECTOR IS
	VARIABLE reslt : std_logic_vector(SrcReg'length - 1 downto 0);
    BEGIN
	reslt := To_TwosComp( To_StdLogicVector(SrcReg), SrcRegMode);
	return  To_StdULogicVector(reslt);
    END To_TwosComp;
--+-----------------------------------------------------------------------------
--|     Function Name  : To_TwosComp
--| 1.8.7
--|     Overloading    : None
--|  
--|     Purpose        : Convert a BIT_VECTOR to Two's Compliment Notation.
--|  
--|     Parameters     :
--|                      SrcReg     - input  BIT_VECTOR, the vector to be read.
--|                      SrcRegMode - input  regmode_type, indicating the format of
--|                                the input BIT_VECTOR.   Default is TwosComp.
--|
--|     Result         : BIT_VECTOR, the vector in Two's complement notation.
--|
--|
--|     Use            :
--|                      VARIABLE vect : BIT_VECTOR ( 15 DOWNTO 0 );
--|                      vect := To_TwosComp ( B"0101",  UnSigned ); -- set to +5
--|
--|     See Also       : To_BitVector, To_Integer, To_TwosComp
--|-----------------------------------------------------------------------------
    FUNCTION To_TwosComp  ( CONSTANT SrcReg      : IN BIT_VECTOR;
                            CONSTANT SrcRegMode  : IN regmode_type
                     -- synopsys synthesis_off
						      := DefaultRegMode 
                     -- synopsys synthesis_on
                          ) RETURN BIT_VECTOR IS

	VARIABLE reslt : std_logic_vector(SrcReg'length - 1 downto 0);
    BEGIN
	reslt := To_TwosComp( To_StdLogicVector(SrcReg), SrcRegMode);
	return  To_BitVector(reslt);
    END To_TwosComp;
--+-----------------------------------------------------------------------------
--|     Function Name  : To_Unsign_FromTwosComp
--| 1.8.11
--|     Overloading    : None
--| 
--|     Purpose        : Convert a STD_LOGIC_VECTOR to Unsigned Notation.
--| 
--|     Parameters     :
--|                      ARG     - input  STD_LOGIC_VECTOR, the vector to be read.
--|                      SIZE    - input  Integer
--|
--|     Result         : STD_LOGIC_VECTOR, the vector in unsigned notation. 
--|
--|
--|     Use            :
--|                      VARIABLE vect : STD_LOGIC_VECTOR ( 15 DOWNTO 0 );
--|                      vect := To_Unsign_FromTwosComp ( "0101", 4); -- set to +5
--|
--|     See Also       : to_BitVector, to_Integer, To_TwosComp, From_TwosComp
--|-----------------------------------------------------------------------------
    FUNCTION To_Unsign_FromTwosComp  ( CONSTANT ARG      : IN STD_LOGIC_VECTOR;
                                       CONSTANT SIZE     : IN INTEGER
                                     ) RETURN STD_LOGIC_VECTOR IS
      VARIABLE reg_copy : STD_LOGIC_VECTOR (ARG'LENGTH - 1 DOWNTO 0);
      VARIABLE result    : STD_LOGIC_VECTOR (ARG'LENGTH - 1 DOWNTO 0);
    BEGIN
	reg_copy := ARG;  		 
	-- synopsys translate_off  
      --  Check for null input
      IF (ARG'LENGTH = 0) THEN

          ASSERT false
          REPORT " To_Unsign --- input register has null range "
          SEVERITY ERROR;
          RETURN reg_copy;

      ELSE
	-- synopsys translate_on      
        result := reg_copy;
          -- convert to unsigned representation.
          -- if a negative value, take two's comp it
          -- will become unsigned
            IF (reg_copy(ARG'LENGTH - 1) /= '0') THEN
              -- if largest negative number then no conversion required
    	          IF ( NOT All_Zero(reg_copy(ARG'LENGTH-2 DOWNTO 0))) THEN
                     result := RegNegate ( reg_copy, TwosComp);
                  END IF;   
            END IF;
       -- synopsys translate_off
       END IF;
       -- synopsys translate_on
       RETURN result;
    END To_Unsign_FromTwosComp;
    -------------------------------------------------------------------------------
    --     Function Name  : To_Unsign
    --
    --     Overloading    : None
    --
    --     Purpose        : Convert a std_logic_vector to Unsigned Notation.
    --
    --     Parameters     :
    --                      SrcReg     - input  std_logic_vector, the vector to be read.
    --                      SrcRegMode - input  regmode_type, indicating the format of
    --                                the input std_logic_vector.   Default is TwosComp.
    --
    --     Result         : std_logic_vector, the vector in unsigned notation.
    --
    --
    --     Use            :
    --                      VARIABLE vect : std_logic_vector ( 15 DOWNTO 0 );
    --                      vect := To_Unsign ( "0l01", TwosComp ); -- set to +5
    --
    --     See Also       : To_StdLogicVector, To_Integer, To_TwosComp, From_TwosComp
  -------------------------------------------------------------------------------
    FUNCTION To_Unsign    ( CONSTANT SrcReg      : IN std_logic_vector;
                            CONSTANT SrcRegMode  : IN regmode_type  
                     -- synopsys synthesis_off
						      := DefaultRegMode 
                     -- synopsys synthesis_on
                          ) RETURN std_logic_vector IS
      VARIABLE reg_copy : std_logic_vector (SrcReg'LENGTH - 1 DOWNTO 0);
    BEGIN
	reg_copy := SrcReg;
	if (SrcRegMode = TwosComp) then
		return(To_Unsign_FromTwosComp(reg_copy, SrcReg'LENGTH));
	else 
		return(reg_copy);
        end if;
    END To_Unsign;
   -------------------------------------------------------------------------------
    --     Function Name  : To_Unsign
    --
    --     Overloading    : None
    --
    --     Purpose        : Convert an std_ulogic_vector to Unsigned Notation.
    --
    --     Parameters     :
    --                      SrcReg     - input  std_ulogic_vector, the vector to be read.
    --                      SrcRegMode - input  regmode_type, indicating the format of
    --                                the input std_ulogic_vector.   Default is TwosComp.
    --
    --     Result         : std_ulogic_vector, the vector in unsigned notation.
    --
    --
    --     Use            :
    --                      VARIABLE vect : std_ulogic_vector ( 15 DOWNTO 0 );
    --                      vect := To_Unsign ( "0l01",TwosComp ); -- set to +5
    --
    --     See Also       : To_StdLogicVector, To_Integer, To_TwosComp, From_TwosComp
  -------------------------------------------------------------------------------
    FUNCTION To_Unsign    ( CONSTANT SrcReg      : IN std_ulogic_vector;
                            CONSTANT SrcRegMode  : IN regmode_type  
                     -- synopsys synthesis_off
						      := DefaultRegMode 
                     -- synopsys synthesis_on
                          ) RETURN std_ulogic_vector IS
	VARIABLE reslt_copy : std_logic_vector (SrcReg'LENGTH - 1 DOWNTO 0);
    BEGIN
	reslt_copy := To_Unsign( To_StdLogicVector(SrcReg), SrcRegMode);
        return To_StdULogicVector(reslt_copy);
    END To_Unsign;
--+-----------------------------------------------------------------------------
--|     Function Name  : To_Unsign
--| 1.8.11
--|     Overloading    : None
--| 
--|     Purpose        : Convert a BIT_VECTOR to Unsigned Notation.
--| 
--|     Parameters     :
--|                      SrcReg     - input  BIT_VECTOR, the vector to be read.
--|                      SrcRegMode - input  regmode_type, indicating the format of
--|                                the input BIT_VECTOR.   Default is TwosComp.
--|
--|     Result         : BIT_VECTOR, the vector in unsigned notation. 
--|
--|
--|     Use            :
--|                      VARIABLE vect : BIT_VECTOR ( 15 DOWNTO 0 );
--|                      vect := To_Unsign ( B"0101", SignMagnitude ); -- set to +5
--|
--|     See Also       : to_BitVector, to_Integer, To_TwosComp, From_TwosComp
--|-----------------------------------------------------------------------------
    FUNCTION To_Unsign    ( CONSTANT SrcReg      : IN BIT_VECTOR;
                            CONSTANT SrcRegMode  : IN regmode_type  
                     -- synopsys synthesis_off
						      := DefaultRegMode 
                     -- synopsys synthesis_on
                          ) RETURN BIT_VECTOR IS

	VARIABLE reslt_copy : std_logic_vector (SrcReg'LENGTH - 1 DOWNTO 0);
    BEGIN
	reslt_copy := To_Unsign( To_StdLogicVector(SrcReg), SrcRegMode);
        return To_BitVector(reslt_copy);
    END To_Unsign;
    -------------------------------------------------------------------------------
    --     Function Name  : To_StdLogicVector_TwosComp
    --
    --     Overloading    : Procedure and Function.
    --
    --     Purpose        : Translate an INTEGER into a std_logic_vector.
    --
    --     Parameters     : ARG    - input  INTEGER, the value to be translated.
    --                      SIZE   - input  INTEGER, length of the return vector.
    --                                Default is IntegerBitLength  (Machine Integer
    --                                length).
    --
    --     Result        : std_logic_vector, the binary representation of the integer.
    --
    --     NOTE          : An ASSERTION message of severity ERROR if the conversion
    --                      fails:
    --                       * 'ARG' is negative and UnSigned format is specified.
    --                         The absolute value of 'ARG' is used.
    --                       * The length of 'SrcReg' is insufficient to hold the
    --                         binary value. The low order bits are returned.
    --
    --                      A runtime system error should occur if the value of
    --                      'SIZE'  does not equal the expected return vector
    --                      length (from the context of the function usage).
    --
   --     Use            :
    --                      VARIABLE vect : std_logic_vector ( 15 DOWNTO 0 );
    --
    --                      vect := To_StdLogicVector_TwosComp ( -294, 16);
    --
    --     See Also       : To_StdLogicVector, To_Integer, To_TwosComp
    -------------------------------------------------------------------------------
    FUNCTION To_StdLogicVector_TwosComp ( CONSTANT ARG       : IN INTEGER;
                                          CONSTANT SIZE      : IN INTEGER
                                        ) RETURN std_logic_vector IS
      CONSTANT bmap         : std_logic_vector(0 TO 1) := "01";
      VARIABLE result       : std_logic_vector (SIZE-1 DOWNTO 0);
      VARIABLE value        : INTEGER;
      VARIABLE maglen, temp : INTEGER;
      VARIABLE negative     : BOOLEAN;
      VARIABLE good         : BOOLEAN;
      -- synopsys built_in SYN_INTEGER_TO_SIGNED

    BEGIN
    -- synopsys synthesis_off
        -- Initializations
	 result   := (OTHERS=>'0');
         value    := ARG;
         negative := FALSE;
         good     := TRUE;
    -- if formatting the logic vector as an unsigned number, the full vector
    -- can be used for the magnitude of the value. Otherwise reduce the size
    -- of the magnitude by 1 to allow for the sign bit.
        maglen := SIZE - 1;

    -- if the input integer value is negative, set the NEGATIVE flag true
    -- and use the absolute value of the integer. Furthermore, if the logic vector
    -- is to be formatted as an unsigned value, set the GOOD status to FALSE.  

       IF (value < 0) Then
          negative := TRUE;                -- set negative flag
          value    := - value;             -- make value positive
       END IF;

       -- Convert the positive integer value to an unsigned logic vector
    -- NOTE: for positive numbers, all formats are the same
    -- if the integer is to big for the return register set GOOD to FALSE.

--      FOR i IN 0 TO IntegerBitLength - 1 LOOP
      FOR i IN 0 TO SIZE - 1 LOOP
--         EXIT WHEN value <= 0;
	if (value <= 0) then
		IF negative THEN
			result := RegNegate(result, TwosComp);
		END IF;
		RETURN result;
	end if;
         temp := value / 2;
         result(i) := bmap(value - (temp*2));
         value := temp;
         IF (i > maglen) THEN 
              good := FALSE; 
         END IF;
      END LOOP;
      ASSERT value=0 
      REPORT "To_StdLogicVector_TwosComp ---  IntegerBitLength too small to hold " &
             " the std_logic  value of the input integer "
      SEVERITY FAILURE;

      IF negative THEN
          result := RegNegate(result, TwosComp);
      END IF;

      RETURN result;
    -- synopsys synthesis_on
    END To_StdLogicVector_TwosComp;

    -------------------------------------------------------------------------------
    --     Function Name  : To_StdLogicVector_Unsigned
    --
    --     Overloading    : Procedure and Function.
    --
    --     Purpose        : Translate an INTEGER into a std_logic_vector.
    --
    --     Parameters     : ARG    - input  INTEGER, the value to be translated.
    --                      SIZE   - input  INTEGER, length of the return vector.
    --                                Default is IntegerBitLength  (Machine Integer
    --                                length).
    --
    --     Result        : std_logic_vector, the binary representation of the integer.
    --
    --     NOTE          : An ASSERTION message of severity ERROR if the conversion
    --                      fails:
    --                       * 'ARG' is negative and UnSigned format is specified.
    --                         The absolute value of 'ARG' is used.
    --                       * The length of 'SrcReg' is insufficient to hold the
    --                         binary value. The low order bits are returned.
    --
    --                      A runtime system error should occur if the value of
    --                      'SIZE'  does not equal the expected return vector
    --                      length (from the context of the function usage).
    --
   --     Use            :
    --                      VARIABLE vect : std_logic_vector ( 15 DOWNTO 0 );
    --
    --                      vect := To_StdLogicVector_Unsigned ( -294, 16);
    --
    --     See Also       : To_StdLogicVector, To_Integer, To_TwosComp
    -------------------------------------------------------------------------------
    FUNCTION To_StdLogicVector_Unsigned ( CONSTANT ARG       : IN INTEGER;
                                          CONSTANT SIZE      : IN INTEGER
                                        ) RETURN std_logic_vector IS
      CONSTANT bmap         : std_logic_vector(0 TO 1) := "01";
      VARIABLE result       : std_logic_vector (SIZE-1 DOWNTO 0);
      VARIABLE value        : INTEGER;
      VARIABLE maglen, temp : INTEGER;
      VARIABLE negative     : BOOLEAN;
      VARIABLE good         : BOOLEAN;
      -- synopsys built_in SYN_INTEGER_TO_UNSIGNED

    BEGIN
    -- synopsys synthesis_off
        -- Initializations
	 result   := (OTHERS=>'0');
         value    := ARG;
         negative := FALSE;
         good     := TRUE;
    -- if formatting the logic vector as an unsigned number, the full vector
    -- can be used for the magnitude of the value. Otherwise reduce the size
    -- of the magnitude by 1 to allow for the sign bit.
        maglen := SIZE;
 
    -- if the input integer value is negative, set the NEGATIVE flag true
    -- and use the absolute value of the integer. Furthermore, if the logic vector
    -- is to be formatted as an unsigned value, set the GOOD status to FALSE.  

      IF (value < 0) Then
          negative := TRUE;                -- set negative flag
          value    := - value;             -- make value positive
          ASSERT not WarningsOn 
          REPORT " To_StdLogicVector --- negative integer with unsigned mode "
          SEVERITY WARNING;
       END IF;

       -- Convert the positive integer value to an unsigned logic vector
    -- NOTE: for positive numbers, all formats are the same
    -- if the integer is to big for the return register set GOOD to FALSE.

      FOR i IN 0 TO IntegerBitLength - 1 LOOP
--         EXIT WHEN value <= 0;
		if (value <= 0) then
			IF negative THEN
				result := RegNegate(result, Unsigned);
			END IF;
			RETURN result;
		end if;
         temp := value / 2;
         result(i) := bmap(value - (temp*2));
         value := temp;
         IF (i > maglen - 1) THEN
              good := FALSE;
         END IF;
      END LOOP;
      ASSERT value=0 
      REPORT "To_StdLogicVector ---  IntegerBitLength too small to hold " &
             " the std_logic  value of the input integer "
      SEVERITY FAILURE;

      IF negative THEN
          result := RegNegate(result, Unsigned);
      END IF;
      RETURN result;
    -- synopsys synthesis_on
    END To_StdLogicVector_Unsigned;

    -------------------------------------------------------------------------------
    --     Function Name  : To_StdLogicVector
    --
    --     Overloading    : Procedure and Function.
    --
    --     Purpose        : Translate an INTEGER into a std_logic_vector.
    --
    --     Parameters     : intg    - input  INTEGER, the value to be translated.
    --                      width   - input  INTEGER, length of the return vector.
    --                                Default is IntegerBitLength  (Machine Integer
    --                                length).
    --                      SrcRegMode - input  regmode_type, indicating the format
    --                                   of the output std_logic_vector.   Default 
    --                                   is TwosComp.
    --
    --     Result        : std_logic_vector, the binary representation of the integer.
    --
    --     NOTE          : An ASSERTION message of severity ERROR if the conversion
    --                      fails:
    --                       * 'intg' is negative and UnSigned format is specified.
    --                         The absolute value of 'intg' is used.
    --                       * The length of 'SrcReg' is insufficient to hold the
    --                         binary value. The low order bits are returned.
    --
    --                      A runtime system error should occur if the value of
    --                      'width'  does not equal the expected return vector
    --                      length (from the context of the function usage).
    --
   --     Use            :
    --                      VARIABLE vect : std_logic_vector ( 15 DOWNTO 0 );
    --
    --                      vect := To_StdLogicVector ( -294, 16, TwosComp );
    --
    --     See Also       : To_StdLogicVector, To_Integer, To_TwosComp
    -------------------------------------------------------------------------------
    FUNCTION To_StdLogicVector ( CONSTANT intg       : IN INTEGER;
                                 CONSTANT width      : IN NATURAL;
                                 CONSTANT SrcRegMode : IN regmode_type  
                     -- synopsys synthesis_off
						      := DefaultRegMode 
                     -- synopsys synthesis_on
                               ) RETURN std_logic_vector IS

    BEGIN
    --
	if (SrcRegMode = Unsigned) Then 
		return (To_StdLogicVector_Unsigned(intg, width));
        else
		return (To_StdLogicVector_TwosComp(intg, width));
        end if;

    END To_StdLogicVector;
    -------------------------------------------------------------------------------
    --     Function Name  : To_StdULogicVector_TwosComp
    --
    --     Overloading    : Procedure and Function.
    --
    --     Purpose        : Translate an INTEGER into a std_logic_vector.
    --
    --     Parameters     : ARG    - input  INTEGER, the value to be translated.
    --                      SIZE   - input  INTEGER, length of the return vector.
    --                                Default is IntegerBitLength  (Machine Integer
    --                                length).
    --
    --     Result        : std_logic_vector, the binary representation of the integer.
    --
    --     NOTE          : An ASSERTION message of severity ERROR if the conversion
    --                      fails:
    --                       * 'ARG' is negative and UnSigned format is specified.
    --                         The absolute value of 'ARG' is used.
    --                       * The length of 'SrcReg' is insufficient to hold the
    --                         binary value. The low order bits are returned.
    --
    --                      A runtime system error should occur if the value of
    --                      'SIZE'  does not equal the expected return vector
    --                      length (from the context of the function usage).
    --
   --     Use            :
    --                      VARIABLE vect : std_logic_vector ( 15 DOWNTO 0 );
    --
    --                      vect := To_StdULogicVector_TwosComp ( -294, 16);
    --
    --     See Also       : To_StdULogicVector, To_Integer, To_TwosComp
    -------------------------------------------------------------------------------
    FUNCTION To_StdULogicVector_TwosComp ( CONSTANT ARG       : IN INTEGER;
                                          CONSTANT SIZE      : IN INTEGER
                                        ) RETURN std_ulogic_vector IS
      CONSTANT bmap         : std_ulogic_vector(0 TO 1) := "01";
      VARIABLE result       : std_ulogic_vector (SIZE-1 DOWNTO 0);
      VARIABLE value        : INTEGER;
      VARIABLE maglen, temp : INTEGER;
      VARIABLE negative     : BOOLEAN;
      VARIABLE good         : BOOLEAN;
      -- synopsys built_in SYN_INTEGER_TO_SIGNED

    BEGIN
    -- synopsys synthesis_off
        -- Initializations
	 result   := (OTHERS=>'0');
         value    := ARG;
         negative := FALSE;
         good     := TRUE;
    -- if formatting the logic vector as an unsigned number, the full vector
    -- can be used for the magnitude of the value. Otherwise reduce the size
    -- of the magnitude by 1 to allow for the sign bit.
        maglen := SIZE - 1;

    -- if the input integer value is negative, set the NEGATIVE flag true
    -- and use the absolute value of the integer. Furthermore, if the logic vector
    -- is to be formatted as an unsigned value, set the GOOD status to FALSE.  

       IF (value < 0) Then
          negative := TRUE;                -- set negative flag
          value    := - value;             -- make value positive
       END IF;

       -- Convert the positive integer value to an unsigned logic vector
    -- NOTE: for positive numbers, all formats are the same
    -- if the integer is to big for the return register set GOOD to FALSE.

--      FOR i IN 0 TO IntegerBitLength - 1 LOOP
      FOR i IN 0 TO SIZE - 1 LOOP
--         EXIT WHEN value <= 0;
		if (value <= 0) then
			IF negative THEN
				result := RegNegate(result, TwosComp);
			END IF;
			RETURN result;
		end if;
         temp := value / 2;
         result(i) := bmap(value - (temp*2));
         value := temp;
         IF (i > maglen) THEN 
              good := FALSE; 
         END IF;
      END LOOP;
      ASSERT value=0 
      REPORT "To_StdULogicVector_TwosComp ---  IntegerBitLength too small to hold " &
             " the std_logic  value of the input integer "
      SEVERITY FAILURE;

      IF negative THEN
          result := RegNegate(result, TwosComp);
      END IF;

      RETURN result;
    -- synopsys synthesis_on
    END To_StdULogicVector_TwosComp;

    -------------------------------------------------------------------------------
    --     Function Name  : To_StdULogicVector_Unsigned
    --
    --     Overloading    : Procedure and Function.
    --
    --     Purpose        : Translate an INTEGER into a std_ulogic_vector.
    --
    --     Parameters     : ARG    - input  INTEGER, the value to be translated.
    --                      SIZE   - input  INTEGER, length of the return vector.
    --                                Default is IntegerBitLength  (Machine Integer
    --                                length).
    --
    --     Result        : std_ulogic_vector, the binary representation of the integer.
    --
    --     NOTE          : An ASSERTION message of severity ERROR if the conversion
    --                      fails:
    --                       * 'ARG' is negative and UnSigned format is specified.
    --                         The absolute value of 'ARG' is used.
    --                       * The length of 'SrcReg' is insufficient to hold the
    --                         binary value. The low order bits are returned.
    --
    --                      A runtime system error should occur if the value of
    --                      'SIZE'  does not equal the expected return vector
    --                      length (from the context of the function usage).
    --
   --     Use            :
    --                      VARIABLE vect : std_ulogic_vector ( 15 DOWNTO 0 );
    --
    --                      vect := To_StdULogicVector_Unsigned ( -294, 16);
    --
    --     See Also       : To_StdULogicVector, To_Integer, To_TwosComp
    -------------------------------------------------------------------------------
    FUNCTION To_StdULogicVector_Unsigned ( CONSTANT ARG       : IN INTEGER;
                                          CONSTANT SIZE      : IN INTEGER
                                        ) RETURN std_ulogic_vector IS
      CONSTANT bmap         : std_ulogic_vector(0 TO 1) := "01";
      VARIABLE result       : std_ulogic_vector (SIZE-1 DOWNTO 0);
      VARIABLE value        : INTEGER;
      VARIABLE maglen, temp : INTEGER;
      VARIABLE negative     : BOOLEAN;
      VARIABLE good         : BOOLEAN;
	-- synopsys built_in SYN_INTEGER_TO_UNSIGNED
    BEGIN
    -- synopsys synthesis_off
        -- Initializations
	 result   := (OTHERS=>'0');
         value    := ARG;
         negative := FALSE;
         good     := TRUE;
    -- if formatting the logic vector as an unsigned number, the full vector
    -- can be used for the magnitude of the value. Otherwise reduce the size
    -- of the magnitude by 1 to allow for the sign bit.
        maglen := SIZE;
 
    -- if the input integer value is negative, set the NEGATIVE flag true
    -- and use the absolute value of the integer. Furthermore, if the logic vector
    -- is to be formatted as an unsigned value, set the GOOD status to FALSE.  

      IF (value < 0) Then
          negative := TRUE;                -- set negative flag
          value    := - value;             -- make value positive
          ASSERT not WarningsOn 
          REPORT " To_StdULogicVector --- negative integer with unsigned mode "
          SEVERITY WARNING;
       END IF;

       -- Convert the positive integer value to an unsigned logic vector
    -- NOTE: for positive numbers, all formats are the same
    -- if the integer is to big for the return register set GOOD to FALSE.

      FOR i IN 0 TO IntegerBitLength - 1 LOOP
--         EXIT WHEN value <= 0;
		if (value <= 0) then
			IF negative THEN
				result := RegNegate(result, Unsigned);
			END IF;
			RETURN result;
		end if;
         temp := value / 2;
         result(i) := bmap(value - (temp*2));
         value := temp;
         IF (i > maglen - 1) THEN
              good := FALSE;
         END IF;
      END LOOP;
      ASSERT value=0 
      REPORT "To_StdULogicVector ---  IntegerBitLength too small to hold " &
             " the std_logic  value of the input integer "
      SEVERITY FAILURE;

      IF negative THEN
          result := RegNegate(result, Unsigned);
      END IF;
      RETURN result;
    -- synopsys synthesis_on
    END To_StdULogicVector_Unsigned;


    -------------------------------------------------------------------------------
    --     Function Name  : To_StdULogicVector
    --
    --     Overloading    : Procedure and Function.
    --
    --     Purpose        : Translate an INTEGER into a std_ulogic_vector.
    --
    --     Parameters     : intg    - input  INTEGER, the value to be translated.
    --                      width   - input  INTEGER, length of the return vector.
    --                                Default is IntegerBitLength  (Machine Integer
    --                                length).
    --                      SrcRegMode - input  regmode_type, indicating the format
    --                                   of the output std_ulogic_vector.   Default 
    --                                   is TwosComp.
    --
    --     Result        : std_ulogic_vector
    --
    --     NOTE          : An ASSERTION message of severity ERROR if the conversion
    --                      fails:
    --                       * 'intg' is negative and UnSigned format is specified.
    --                         The absolute value of 'intg' is used.
    --                       * The length of 'SrcReg' is insufficient to hold the
    --                         binary value. The low order bits are returned.
    --
    --                      A runtime system error should occur if the value of
    --                      'width'  does not equal the expected return vector
    --                      length (from the context of the function usage).
    --
   --     Use            :
    --                      VARIABLE vect : std_logic_vector ( 15 DOWNTO 0 );
    --
    --                      vect := To_StdULogicVector ( -294, 16, TwosComp );
    --
    --     See Also       : To_StdLogicVector, To_Integer, To_TwosComp
    -------------------------------------------------------------------------------
    FUNCTION To_StdULogicVector ( CONSTANT intg       : IN INTEGER;
                                  CONSTANT width      : IN NATURAL ;
                                  CONSTANT SrcRegMode : IN regmode_type  
                     -- synopsys synthesis_off
						      := DefaultRegMode 
                     -- synopsys synthesis_on
                                ) RETURN std_ulogic_vector IS
    BEGIN
    --
	if (SrcRegMode = Unsigned) Then 
		return (To_StdULogicVector_Unsigned(intg, width));
        else
		return (To_StdULogicVector_TwosComp(intg, width));
        end if;

    END To_StdULogicVector;

--+-----------------------------------------------------------------------------
--|     Function Name  : To_BitVector_TwosComp
--|
--|     Overloading    : 
--|
--|     Purpose        : Translate an INTEGER into a BIT_VECTOR in TwosComp Mode
--|
--|     Parameters     : ARG    - input  INTEGER, the value to be translated.
--|                      SIZE   - input  INTEGER, length of the return vector.
--|
--|     Result        : BIT_VECTOR, the binary representation of the integer.
--|
--|     NOTE           : An ASSERTION message of severity ERROR if the conversion
--|                      fails:
--|                       * 'ARG' is negative and UnSigned format is specified.
--|                         The absolute value of 'ARG' is used.
--|                       * The length of 'SrcReg' is insufficient to hold the
--|                         binary value. The low order bits are returned.
--|
--|                      A runtime system error should occur if the value of
--|                      'SIZE' is does not equal the expected return vector
--|                      length (from the context of the function usage).
--|
--|     Use            :
--|                      VARIABLE vect : BIT_VECTOR ( 15 DOWNTO 0 );
--|
--|                      vect := To_BitVector_TwosComp ( -294, 16);
--|
--|     See Also       : To_BitVector, To_Integer, To_TwosComp
--|-----------------------------------------------------------------------------
    FUNCTION To_BitVector_TwosComp ( CONSTANT ARG       : IN INTEGER;
                            CONSTANT SIZE      : IN INTEGER
                          ) RETURN BIT_VECTOR IS
      VARIABLE result   : BIT_VECTOR (SIZE-1 DOWNTO 0);
      VARIABLE value    : INTEGER;
      VARIABLE maglen   : Integer;     -- magnitude length
      VARIABLE temp     : Integer;
      VARIABLE negative : Boolean;
      VARIABLE good     : Boolean;
      -- synopsys built_in SYN_INTEGER_TO_SIGNED

    BEGIN
	-- synopsys synthesis_off
        -- Initializations
	result   := (OTHERS=>'0');
        value    := ARG;
        negative := FALSE;
        good     := TRUE;
        maglen := SIZE - 1;
	IF (value < 0) Then
          negative := TRUE;                -- set negative flag
          value    := - value;             -- make value positive
        END IF;

       -- Convert the positive integer value to an unsigned bit vector
       -- NOTE: for positive numbers, all formats are the same
       -- if the integer is to big for the return register set GOOD to FALSE.

--        FOR i IN 0 TO IntegerBitLength - 1 LOOP
        FOR i IN 0 TO SIZE - 1 LOOP
--		EXIT WHEN value <= 0;
		if (value <= 0) then
			IF negative THEN
				result := RegNegate(result, TwosComp);
			END IF;
			RETURN result;
		end if;
           temp := value / 2;
--           result(i) := BIT'VAL(value - (temp*2));
		if ((value-(temp*2)) = 0) then
			result(i) := '0';
		else
			result(i) := '1';
		end if;
           value := temp;
           IF (i > maglen) THEN 
              good := FALSE; 
           END IF;
        END LOOP;
        ASSERT value=0 
        REPORT "To_BitVector ---  IntegerBitLength too small to hold " &
             " the binary value of the input integer "
        SEVERITY FAILURE;

       IF negative THEN
          result := RegNegate(result, TwosComp);
       END IF;
       RETURN result;
       -- synopsys synthesis_on
    END To_BitVector_TwosComp;
--+-----------------------------------------------------------------------------
--|     Function Name  : To_BitVector_Unsigned
--|
--|     Overloading    : 
--|
--|     Purpose        : Translate an INTEGER into a BIT_VECTOR in Unsigned Mode
--|
--|     Parameters     : ARG    - input  INTEGER, the value to be translated.
--|                      SIZE   - input  INTEGER, length of the return vector.

--|
--|     Result        : BIT_VECTOR, the binary representation of the integer.
--|
--|     NOTE           : An ASSERTION message of severity ERROR if the conversion
--|                      fails:
--|                       * 'ARG' is negative and UnSigned format is specified.
--|                         The absolute value of 'ARG' is used.
--|                       * The length of 'SrcReg' is insufficient to hold the
--|                         binary value. The low order bits are returned.
--|
--|                      A runtime system error should occur if the value of
--|                      'SIZE' is does not equal the expected return vector
--|                      length (from the context of the function usage).
--|
--|     Use            :
--|                      VARIABLE vect : BIT_VECTOR ( 15 DOWNTO 0 );
--|
--|                      vect := To_BitVector_Unsigned ( -294, 16);
--|
--|     See Also       : To_BitVector, To_Integer, To_Unsigned
--|-----------------------------------------------------------------------------
    FUNCTION To_BitVector_Unsigned ( CONSTANT ARG       : IN INTEGER;
                            CONSTANT SIZE      : IN INTEGER
                          ) RETURN BIT_VECTOR IS
      VARIABLE result   : BIT_VECTOR (SIZE-1 DOWNTO 0);
      VARIABLE value    : INTEGER;
      VARIABLE maglen   : Integer;     -- magnitude length
      VARIABLE temp     : Integer;
      VARIABLE negative : Boolean;
      VARIABLE good     : Boolean;
      -- synopsys built_in SYN_INTEGER_TO_UNSIGNED

    BEGIN
	-- synopsys synthesis_off
        -- Initializations
	result   := (OTHERS=>'0');
        value    := ARG;
        negative := FALSE;
        good     := TRUE;
        maglen := SIZE;
	IF (value < 0) Then
          negative := TRUE;                -- set negative flag
          value    := - value;             -- make value positive
           ASSERT not WarningsOn 
           REPORT " To_BitVector --- negative integer with unsigned mode "
           SEVERITY WARNING;
        END IF;

       -- Convert the positive integer value to an unsigned bit vector
    -- NOTE: for positive numbers, all formats are the same
    -- if the integer is to big for the return register set GOOD to FALSE.

      FOR i IN 0 TO IntegerBitLength - 1 LOOP
--         EXIT WHEN value <= 0;
		if (value <= 0) then
			IF negative THEN
				result := RegNegate(result, Unsigned);
			END IF;
			RETURN result;
		end if;
         temp := value / 2;
         result(i) := BIT'VAL(value - (temp*2));
         value := temp;
         IF (i > maglen - 1) THEN
              good := FALSE;
         END IF;
      END LOOP;
      ASSERT value=0 
      REPORT "To_BitVector ---  IntegerBitLength too small to hold " &
             " the binary value of the input integer "
      SEVERITY FAILURE;

      IF negative THEN
          result := RegNegate(result, Unsigned);
      END IF;

      RETURN result;
       -- synopsys synthesis_on
    END To_BitVector_Unsigned;
--+-----------------------------------------------------------------------------
--|     Function Name  : To_BitVector
--|
--|     Overloading    : 
--|
--|     Purpose        : Translate an INTEGER into a BIT_VECTOR.
--|
--|     Parameters     : intg    - input  INTEGER, the value to be translated.
--|                      width   - input  NATURAL, length of the return vector.
--|                            Default is IntegerBitLength (Machine integer length).
--|                      SrcRegMode - input  regmode_type, indicating the format of
--|                                the output BIT_VECTOR.   Default is TwosComp.
--|
--|     Result        : BIT_VECTOR, the binary representation of the integer.
--|
--|     NOTE           : An ASSERTION message of severity ERROR if the conversion
--|                      fails:
--|                       * 'intg' is negative and UnSigned format is specified.
--|                         The absolute value of 'intg' is used.
--|                       * The length of 'SrcReg' is insufficient to hold the
--|                         binary value. The low order bits are returned.
--|
--|                      A runtime system error should occur if the value of
--|                      'width' is does not equal the expected return vector
--|                      length (from the context of the function usage).
--|
--|     Use            :
--|                      VARIABLE vect : BIT_VECTOR ( 15 DOWNTO 0 );
--|
--|                      vect := To_BitVector ( -294, 16, TwosComp );
--|
--|     See Also       : To_BitVector, To_Integer, To_TwosComp
--|-----------------------------------------------------------------------------
    FUNCTION To_BitVector ( CONSTANT intg       : IN INTEGER;
                            CONSTANT width      : IN Natural;
                            CONSTANT SrcRegMode : IN regmode_type  
                     -- synopsys synthesis_off
						      := DefaultRegMode 
                     -- synopsys synthesis_on
                          ) RETURN BIT_VECTOR IS
    BEGIN
    --
	if (SrcRegMode = Unsigned) Then 
		return (To_BitVector_Unsigned(intg, width));
        else
		return (To_BitVector_TwosComp(intg, width));
        end if;
    END To_BitVector;
--+-----------------------------------------------------------------------------
--|     Procedure Name : To_Integer_FromTwosComp
--|
--|     Overloading    : 
--|
--|     Purpose        : Interpret BIT_VECTOR as an INTEGER.
--|
--|     Parameters     :
--|                      ARG     - input  BIT_VECTOR, the vector to be read.
--|
--|     NOTE           : 
--|                       * Magnitude of the computed integer is to large. The
--|                         input value is considered to large if after removing
--|                         leading 0's (1's for negative numbers) the length
--|                         of the remaining vector is > IntegerBitLength - 1.
--|                         (ie the machine integer length).
--|                      The error return value is INTEGER'LEFT.
--|
--|     Use            :
--|                      VARIABLE vect : BIT_VECTOR ( 15 DOWNTO 0 );
--|
--|                      To_Integer ( vect, 16);
--|
--|     See Also       : To_BitVector, To_Integer, To_TwosComp 
--|-----------------------------------------------------------------------------
     FUNCTION To_Integer_FromTwosComp  ( CONSTANT ARG    : IN BIT_VECTOR
                                       ) return INTEGER IS
 
	VARIABLE reg_copy   	: BIT_VECTOR(ARG'LENGTH - 1 DOWNTO 0);
	VARIABLE result 	: INTEGER;
	-- synopsys built_in SYN_SIGNED_TO_INTEGER
    BEGIN
	-- synopsys synthesis_off
	-- initializations  
	reg_copy := ARG;
	result   := 0;
     --  Check for null input
	IF (ARG'LENGTH = 0) THEN
          ASSERT false
          REPORT " To_Integer (Bit_Vector case) --- input register has null range, " 
                 & "  returning zero  result  "
          SEVERITY ERROR;
          RETURN 0;
        END IF;

        -- now convert the magnitude part of the bit vector to a positive integer.
        -- if the magnitude part is positive convert with this loop
        IF (reg_copy(ARG'LENGTH - 1)='0') THEN
        -- Convert Unsigned
           FOR i IN ARG'LENGTH-2 DOWNTO 0 LOOP
              IF ((i>=IntegerBitLength - 1) AND (reg_copy(i)='1'))   THEN -- number too big
       	         assert false
	         report " To_Integer (BitVector case) -- attempt to convert a vector "
		       & "larger than or 32 bit  "
	         severity error;
		return 0;
	      END IF;		
--              result := result + result + BIT'POS(reg_copy(i));  -- shift and add
		if (reg_copy(i)='0') then
			result := result + result + 0;  -- shift and add
		elsif (reg_copy(i)='1') then
			result := result + result + 1;  -- shift and add
		end if;
           END LOOP;
  
        -- if the magnitude part is negative convert with this loop
        -- (the bits of the input vector are complemented)
        ELSE  -- Convert Negative number
            FOR i IN ARG'LENGTH-2 DOWNTO 0 LOOP
               IF ((i>=IntegerBitLength - 1) AND (reg_copy(i)='0')) THEN  -- number too big
       	         assert false
	         report " To_Integer (BitVector case) -- attempt to convert a vector "
		       & "larger than 32 bit.  "
	         severity error;
		return 0;
	       END IF;		
--               result := result + result - BIT'POS(reg_copy(i)) + 1; -- shift and add complemented bit
		if (reg_copy(i)='0') then
			result := result + result - 0 + 1; -- shift and add complemented bit
		elsif (reg_copy(i)='1') then
			result := result + result - 1 + 1; -- shift and add complemented bit
		end if;
            END LOOP;
           -- adjust (add 1) for 2's comp numbers
               IF (result = INTEGER'HIGH) THEN              -- number to big
       	         assert false
	         report " To_Integer (BitVector case) -- attempt to convert a vector "
		       & "larger than or 32 bit  "
	         severity error;
		return 0;
	      END IF;		
              result := result + 1;
            -- since this is a negative number, make it so.
            result := - result;
        END IF;
		return result;
	-- synopsys synthesis_on    
    END To_Integer_FromTwosComp;

--+-----------------------------------------------------------------------------
--|     Procedure Name : To_Integer_FromUnsign
--|
--|     Overloading    : 
--|
--|     Purpose        : Interpret BIT_VECTOR as an INTEGER.
--|
--|     Parameters     :
--|                      ARG     - input  BIT_VECTOR, the vector to be read.
--|
--|     NOTE           : 
--|                       * Magnitude of the computed integer is to large. The
--|                         input value is considered to large if after removing
--|                         leading 0's (1's for negative numbers) the length
--|                         of the remaining vector is > IntegerBitLength - 1.
--|                         (ie the machine integer length).
--|                      The error return value is INTEGER'LEFT.
--|
--|     Use            :
--|                      VARIABLE vect : BIT_VECTOR ( 15 DOWNTO 0 );
--|
--|                      To_Integer ( vect);
--|
--|     See Also       : To_BitVector, To_Integer, To_TwosComp 
--|-----------------------------------------------------------------------------
     FUNCTION To_Integer_FromUnsign   ( CONSTANT ARG    : IN BIT_VECTOR
                                       ) return INTEGER IS
 
	VARIABLE reg_copy   	: BIT_VECTOR(ARG'LENGTH - 1 DOWNTO 0);
	VARIABLE result 	: INTEGER;
	-- synopsys built_in SYN_UNSIGNED_TO_INTEGER
    BEGIN
	-- synopsys synthesis_off
	-- initializations  
	reg_copy := ARG;
	result   := 0;
     	--  Check for null input
	IF (ARG'LENGTH = 0) THEN
          ASSERT false
          REPORT " To_Integer (Bit_Vector case) --- input register has null range, " 
                 & "  returning zero  result  "
          SEVERITY ERROR;
          RETURN result;
        END IF;

        -- if the input vector is unsigned, the leading bit is data. 
        -- Now convert the magnitude part of the bit vector to a positive integer.
        -- Convert Unsigned
           FOR i IN ARG'LENGTH DOWNTO 1 LOOP
              IF ((i>=IntegerBitLength) AND (reg_copy(i-1)='1'))   THEN -- number too big
       	         assert false
	         report " To_Integer (BitVector case) -- attempt to convert a vector "
		       & "larger than or 32 bit  "
	         severity error;
		return 0;
	      END IF;		
--              result := result + result + BIT'POS(reg_copy(i-1));  -- shift and add
		if (reg_copy(i-1)='0') then
			result := result + result + 0;  -- shift and add
		elsif (reg_copy(i-1)='1') then
			result := result + result + 1;  -- shift and add
		end if;
           END LOOP;
		return result;
	-- synopsys synthesis_on    
    END To_Integer_FromUnsign;


--+-----------------------------------------------------------------------------
--|     Procedure Name : To_Integer
--|
--|     Overloading    : 
--|
--|     Purpose        : Interpret BIT_VECTOR as an INTEGER.
--|
--|     Parameters     :
--|                      SrcReg     - input  BIT_VECTOR, the vector to be read.
--|                      SrcRegMode - input  regmode_type, indicating the format of
--|                                the input BIT_VECTOR.   Default is TwosComp.
--|
--|     NOTE           : 
--|                       * Magnitude of the computed integer is to large. The
--|                         input value is considered to large if after removing
--|                         leading 0's (1's for negative numbers) the length
--|                         of the remaining vector is > IntegerBitLength - 1.
--|                         (ie the machine integer length).
--|                      The error return value is INTEGER'LEFT.
--|
--|     Use            :
--|                      VARIABLE vect : BIT_VECTOR ( 15 DOWNTO 0 );
--|
--|                      To_Integer ( vect, TwosComp );
--|
--|     See Also       : To_BitVector, To_Integer, To_TwosComp 
--|-----------------------------------------------------------------------------
     FUNCTION To_Integer  ( CONSTANT SrcReg     : IN BIT_VECTOR;
                            CONSTANT SrcRegMode : IN regmode_type
                     -- synopsys synthesis_off
						      := DefaultRegMode 
                     -- synopsys synthesis_on
                          ) return INTEGER IS
 
     BEGIN
	if (SrcRegMode = TwosComp) then
		return(To_Integer_FromTwosComp(SrcReg));
	else 
		return(To_Integer_FromUnsign(SrcReg));
	end if;
    END To_Integer;

--+-----------------------------------------------------------------------------
--|     Procedure Name : To_Integer_FromTwosComp
--|
--|     Overloading    : 
--|
--|     Purpose        : Interpret STD_LOGIC_VECTOR as an INTEGER.
--|
--|     Parameters     :
--|                      ARG     - input  STD_LOGIC_VECTOR, the vector to be read.
--|
--|     NOTE           : 
--|                       * Magnitude of the computed integer is to large. The
--|                         input value is considered to large if after removing
--|                         leading 0's (1's for negative numbers) the length
--|                         of the remaining vector is > IntegerBitLength - 1.
--|                         (ie the machine integer length).
--|                      The error return value is INTEGER'LEFT.
--|
--|     Use            :
--|                      VARIABLE vect : STD_LOGIC_VECTOR ( 15 DOWNTO 0 );
--|
--|                      To_Integer ( vect, 16);
--|
--|     See Also       : To_BitVector, To_Integer, To_TwosComp 
--|-----------------------------------------------------------------------------
     FUNCTION To_Integer_FromTwosComp  ( CONSTANT ARG    : IN STD_LOGIC_VECTOR
                                       ) return INTEGER IS
 
	VARIABLE reg_copy   : STD_LOGIC_VECTOR(ARG'LENGTH - 1 DOWNTO 0);
	VARIABLE result : INTEGER;
	-- synopsys built_in SYN_SIGNED_TO_INTEGER
    BEGIN
	-- synopsys synthesis_off
	-- initializations  
	reg_copy := ARG;
	result   := 0;
     --  Check for null input
	IF (ARG'LENGTH = 0) THEN
          ASSERT false
          REPORT " To_Integer (Std_Logic_Vector case) --- input register has null range, " 
                 & "  returning zero  result  "
          SEVERITY ERROR;
          RETURN 0;
        END IF;

          -- now convert the magnitude part of the logic vector to a positive integer.
          -- if the magnitude part is positive convert with this loop
            IF (reg_copy(ARG'LENGTH - 1)='0') THEN
              -- Convert Unsigned
                FOR i IN ARG'LENGTH - 2 DOWNTO 0 LOOP
                                            -- number too big
                  IF ((i>=IntegerBitLength - 1) AND (reg_copy(i)='1'))   THEN 
         	       assert false
	               report " To_Integer (Std_logic_vector case) -- attempt to convert a vector "
		         & "larger than or 32 bit  "
	               severity error;
			return 0;
                  END IF;		
--                  result := result + result + std_logic'POS(reg_copy(i)) - 2;  -- shift and add
			if ((reg_copy(i)='0') or (reg_copy(i)='L')) then
				result := result + result + 2 - 2;  -- shift and add
			elsif ((reg_copy(i)='1') or (reg_copy(i)='H')) then
				result := result + result + 3 - 2;  -- shift and add
			else
--				result := result + result + 4 - 2;  -- shift and add
				ASSERT false
				REPORT " To_Integer (Std_Logic_Vector case) -- input vector has element "
					& "other than 0, 1, L, H "
				SEVERITY ERROR;
				result := 0;
				return result;
			end if;
               END LOOP;
                  -- if the magnitude part is negative convert with this loop 
                  -- (the bits of the input vector are complemented)
            ELSE  -- Convert Negative number
                FOR i IN ARG'LENGTH - 2 DOWNTO 0 LOOP
                    IF ((i>=IntegerBitLength - 1) AND (reg_copy(i)='0'))   THEN 
         	       assert false
	               report " To_Integer (Std_logic_vector case) -- attempt to convert a vector "
		         & "larger than or 32 bit  "
	               severity error;
			return 0;
                    END IF;		
                   -- shift and add complemented bit
--                    result := result + result - std_logic'POS(reg_copy(i)) + 3; 
			if ((reg_copy(i)='0') or (reg_copy(i)='L'))then
				result := result + result - 2 + 3; 
			elsif ((reg_copy(i)='1') or (reg_copy(i)='H'))then
				result := result + result - 3 + 3; 
			else
--				result := result + result - 4 + 3; 
				ASSERT false
				REPORT " To_Integer (Std_Logic_Vector case) -- input vector has element "
					& "other than 0, 1, L, H "
				SEVERITY ERROR;
				result := 0;
				return result;
			end if;
               END LOOP;
               -- adjust (add 1) for 2's comp numbers
               IF (result = INTEGER'HIGH) THEN              -- number to big
         	       assert false
	               report " To_Integer (Std_logic_vector case) -- attempt to convert a vector "
		         & "larger than or 32 bit  "
	               severity error;
			return 0;
                END IF;		
                result := result + 1;
               -- since this is a negative number, make it so.
                result := - result;
            END IF;
		return result;
	-- synopsys synthesis_on    
    END To_Integer_FromTwosComp;

--+-----------------------------------------------------------------------------
--|     Procedure Name : To_Integer_FromUnsign
--|
--|     Overloading    : 
--|
--|     Purpose        : Interpret STD_LOGIC_VECTOR as an INTEGER.
--|
--|     Parameters     :
--|                      ARG     - input  STD_LOGIC_VECTOR, the vector to be read.
--|
--|     NOTE           : 
--|                       * Magnitude of the computed integer is to large. The
--|                         input value is considered to large if after removing
--|                         leading 0's (1's for negative numbers) the length
--|                         of the remaining vector is > IntegerBitLength - 1.
--|                         (ie the machine integer length).
--|                      The error return value is INTEGER'LEFT.
--|
--|     Use            :
--|                      VARIABLE vect : STD_LOGIC_VECTOR ( 15 DOWNTO 0 );
--|
--|                      To_Integer ( vect);
--|
--|     See Also       : To_BitVector, To_Integer, To_TwosComp 
--|-----------------------------------------------------------------------------
     FUNCTION To_Integer_FromUnsign   ( CONSTANT ARG    : IN STD_LOGIC_VECTOR
                                       ) return INTEGER IS
 
	VARIABLE reg_copy   	: STD_LOGIC_VECTOR(ARG'LENGTH - 1 DOWNTO 0);
	VARIABLE result 	: INTEGER;
	-- synopsys built_in SYN_UNSIGNED_TO_INTEGER
    BEGIN
	-- synopsys synthesis_off
	-- initializations  
	reg_copy := ARG;
	result   := 0;
     	--  Check for null input
	IF (ARG'LENGTH = 0) THEN
          ASSERT false
          REPORT " To_Integer (Std_Logic_Vector case) --- input register has null range, " 
                 & "  returning zero  result  "
          SEVERITY ERROR;
          RETURN result;
        END IF;

	-- if the input vector is unsigned, the leading bit is data.
	-- now convert the magnitude part of the logic vector to a positive integer.
	-- if the magnitude part is positive convert with this loop
            FOR i IN ARG'LENGTH DOWNTO 1 LOOP
                  IF ((i>=IntegerBitLength) AND (reg_copy(i-1)='1'))   THEN 
                                            -- number too big
         	       assert false
	               report " To_Integer (Std_logic_vector case) -- attempt to convert a vector "
		         & "larger than or 32 bit  "
	               severity error;
			return 0;
                  END IF;		
--                  result := result + result + std_logic'POS(reg_copy(i-1)) - 2;  -- shift and add
			if ((reg_copy(i-1)='0') or (reg_copy(i-1)='L')) then
				result := result + result + 2 - 2;  -- shift and add
			elsif ((reg_copy(i-1)='1') or (reg_copy(i-1)='H')) then
				result := result + result + 3 - 2;  -- shift and add
			else
--				result := result + result + 4 - 2;  -- shift and add
				ASSERT false
				REPORT " To_Integer (Std_Logic_Vector case) -- input vector has element "
					& "other than 0, 1, L, H "
				SEVERITY ERROR;
				result := 0;
				return result;
			end if;
            END LOOP;
		return result;
	-- synopsys synthesis_on    
    END To_Integer_FromUnsign;

    -------------------------------------------------------------------------------
    --     Procedure Name : To_Integer
    --
    --     Overloading    : Procedure and Function.
    --    
    --     Purpose        : Interpret std_logic_vector as an INTEGER.
    --     
    --     Parameters     : 
    --                      SrcReg     - input  std_logic_vector, the vector to be 
    --                                          converted.
    --                      SrcRegMode - input  regmode_type, indicating the format 
    --                                    of the input std_logic_vector.   
    --                                    Default is DefaultRegMode.
    --     
    --     NOTE           : 
    --                      * Magnitude of the computed integer is to large. The 
    --                        input value is considered to large if after removing
    --                        leading 0's (1's for negative numbers)  the length
    --                        of the remaining vector is > IntegerBitLength-1.
    --                        (ie the machine integer length).
    --                      The error return value is INTEGER'LEFT.
    --
    --     Use            : 
    --                      VARIABLE vect : std_logic_vector ( 15 DOWNTO 0 );
    --
    --                      To_Integer ( vect, TwosComp );
    --     
    --     See Also       :  To_Integer, To_TwosComp, To_OnesComp
    -------------------------------------------------------------------------------
    FUNCTION To_Integer   ( CONSTANT SrcReg     : IN std_logic_vector;
                            CONSTANT SrcRegMode : IN regmode_type 
                     -- synopsys synthesis_off
						      := DefaultRegMode 
                     -- synopsys synthesis_on
                          ) RETURN INTEGER IS
                             
     BEGIN
	if (SrcRegMode = TwosComp) then
		return(To_Integer_FromTwosComp(SrcReg));
	else 
		return(To_Integer_FromUnsign(SrcReg));
	end if;
    END To_Integer;
--+-----------------------------------------------------------------------------
--|     Procedure Name : To_Integer_FromTwosComp
--|
--|     Overloading    : 
--|
--|     Purpose        : Interpret STD_ULOGIC_VECTOR as an INTEGER.
--|
--|     Parameters     :
--|                      ARG     - input  STD_ULOGIC_VECTOR, the vector to be read.
--|
--|     NOTE           : 
--|                       * Magnitude of the computed integer is to large. The
--|                         input value is considered to large if after removing
--|                         leading 0's (1's for negative numbers) the length
--|                         of the remaining vector is > IntegerBitLength - 1.
--|                         (ie the machine integer length).
--|                      The error return value is INTEGER'LEFT.
--|
--|     Use            :
--|                      VARIABLE vect : STD_ULOGIC_VECTOR ( 15 DOWNTO 0 );
--|
--|                      To_Integer ( vect, 16);
--|
--|     See Also       : To_BitVector, To_Integer, To_TwosComp 
--|-----------------------------------------------------------------------------
     FUNCTION To_Integer_FromTwosComp  ( CONSTANT ARG    : IN STD_ULOGIC_VECTOR
                                       ) return INTEGER IS
 
	VARIABLE reg_copy   : STD_ULOGIC_VECTOR(ARG'LENGTH - 1 DOWNTO 0);
	VARIABLE result : INTEGER;
	-- synopsys built_in SYN_SIGNED_TO_INTEGER
    BEGIN
	-- synopsys synthesis_off
	-- initializations  
	reg_copy := ARG;
	result   := 0;
     --  Check for null input
	IF (ARG'LENGTH = 0) THEN
          ASSERT false
          REPORT " To_Integer (Std_Ulogic_Vector case) --- input register has null range, " 
                 & "  returning zero  result  "
          SEVERITY ERROR;
          RETURN 0;
        END IF;

          -- now convert the magnitude part of the logic vector to a positive integer.
          -- if the magnitude part is positive convert with this loop
            IF (reg_copy(ARG'LENGTH - 1)='0') THEN
              -- Convert Unsigned
                FOR i IN ARG'LENGTH-2 DOWNTO 0 LOOP
                                            -- number too big
                  IF ((i>=IntegerBitLength - 1) AND (reg_copy(i)='1'))   THEN 
         	       assert false
	               report " To_Integer (std_ulogic_vector case) -- attempt to convert a vector "
		         & "larger than or 32 bit  "
	               severity error;
			return 0;
                  END IF;		
--                  result := result + result + std_ulogic'POS(reg_copy(i)) - 2;  -- shift and add
			if ((reg_copy(i)='0') or (reg_copy(i)='L')) then
				result := result + result + 2 - 2;  -- shift and add
			elsif ((reg_copy(i)='1') or (reg_copy(i)='H'))then
				result := result + result + 3 - 2;  -- shift and add
			else
--				result := result + result + 4 - 2;  -- shift and add
				ASSERT false
				REPORT " To_Integer (Std_Ulogic_Vector case) -- input vector has element "
					& "other than 0, 1, L, H "
				SEVERITY ERROR;
				result := 0;
				return result;
			end if;
               END LOOP;
                  -- if the magnitude part is negative convert with this loop 
                  -- (the bits of the input vector are complemented)
            ELSE  -- Convert Negative number
                FOR i IN ARG'LENGTH - 2 DOWNTO 0 LOOP
                    IF ((i>=IntegerBitLength - 1) AND (reg_copy(i)='0'))   THEN 
         	       assert false
	               report " To_Integer (std_ulogic_vector case) -- attempt to convert a vector "
		         & "larger than or 32 bit  "
	               severity error;
			return 0;
                    END IF;		
                   -- shift and add complemented bit
--                    result := result + result - std_ulogic'POS(reg_copy(i)) + 3; 
			if ((reg_copy(i)='0') or (reg_copy(i)='L')) then
				result := result + result - 2 + 3;  -- shift and add
			elsif ((reg_copy(i)='1') or (reg_copy(i)='H'))then
				result := result + result - 3 + 3;  -- shift and add
			else
--				result := result + result - 4 + 3;  -- shift and add
				ASSERT false
				REPORT " To_Integer (Std_Ulogic_Vector case) -- input vector has element "
					& "other than 0, 1, L, H "
				SEVERITY ERROR;
				result := 0;
				return result;
			end if;
               END LOOP;
               -- adjust (add 1) for 2's comp numbers
               IF (result = INTEGER'HIGH) THEN              -- number to big
         	       assert false
	               report " To_Integer (std_ulogic_vector case) -- attempt to convert a vector "
		         & "larger than or 32 bit  "
	               severity error;
			return 0;
                END IF;		
                result := result + 1;
               -- since this is a negative number, make it so.
                result := - result;
            END IF;
		return result;
	-- synopsys synthesis_on    
    END To_Integer_FromTwosComp;
--+-----------------------------------------------------------------------------
--|     Procedure Name : To_Integer_FromUnsign
--|
--|     Overloading    : 
--|
--|     Purpose        : Interpret STD_ULOGIC_VECTOR as an INTEGER.
--|
--|     Parameters     :
--|                      ARG     - input  STD_ULOGIC_VECTOR, the vector to be read.
--|
--|     NOTE           : 
--|                       * Magnitude of the computed integer is to large. The
--|                         input value is considered to large if after removing
--|                         leading 0's (1's for negative numbers) the length
--|                         of the remaining vector is > IntegerBitLength - 1.
--|                         (ie the machine integer length).
--|                      The error return value is INTEGER'LEFT.
--|
--|     Use            :
--|                      VARIABLE vect : STD_ULOGIC_VECTOR ( 15 DOWNTO 0 );
--|
--|                      To_Integer ( vect);
--|
--|     See Also       : To_BitVector, To_Integer, To_TwosComp 
--|-----------------------------------------------------------------------------
     FUNCTION To_Integer_FromUnsign   ( CONSTANT ARG    : IN STD_ULOGIC_VECTOR
                                       ) return INTEGER IS
 
	VARIABLE reg_copy   	: STD_ULOGIC_VECTOR(ARG'LENGTH - 1 DOWNTO 0);
	VARIABLE result 	: INTEGER;
	-- synopsys built_in SYN_UNSIGNED_TO_INTEGER
    BEGIN
	-- synopsys synthesis_off
	-- initializations
	reg_copy := ARG;
	result   := 0;
	--  Check for null input
	IF (ARG'LENGTH = 0) THEN
          ASSERT false
          REPORT " To_Integer (Std_Ulogic_Vector case) --- input register has null range, " 
                 & "  returning zero  result  "
          SEVERITY ERROR;
          RETURN result;
        END IF;

	-- if the input vector is unsigned, the leading bit is data. 
	-- now convert the magnitude part of the logic vector to a positive integer.
	-- if the magnitude part is positive convert with this loop
            FOR i IN ARG'LENGTH DOWNTO 1 LOOP
                  IF ((i>=IntegerBitLength) AND (reg_copy(i-1)='1'))   THEN 
                                            -- number too big
         	       assert false
	               report " To_Integer (std_ulogic_vector case) -- attempt to convert a vector "
		         & "larger than or 32 bit  "
	               severity error;
			return 0;
                  END IF;		
--                  result := result + result + std_ulogic'POS(reg_copy(i-1)) - 2;  -- shift and add
			if ((reg_copy(i-1) = '0') or (reg_copy(i-1)='L'))then
				result := result + result + 2 - 2;  -- shift and add
			elsif ((reg_copy(i-1) = '1') or (reg_copy(i-1)='H'))then
				result := result + result + 3 - 2;  -- shift and add
			else
--				result := result + result + 4 - 2;  -- shift and add
				ASSERT false
				REPORT " To_Integer (Std_Ulogic_Vector case) -- input vector has element "
					& "other than 0, 1, L, H "
				SEVERITY ERROR;
				result := 0;
				return result;
			end if;
            END LOOP;
           return result;
	-- synopsys synthesis_on    
    END To_Integer_FromUnsign;

    -------------------------------------------------------------------------------
    --     Procedure Name : To_Integer
    --
    --     Overloading    : Procedure and Function.
    --    
    --     Purpose        : Interpret std_ulogic_vector as an INTEGER.
    --     
    --     Parameters     : 
    --                      SrcReg     - input  std_ulogic_vector, the vector to be 
    --                                          converted.
    --                      SrcRegMode - input  regmode_type, indicating the format 
    --                                    of the input std_ulogic_vector.   
    --                                    Default is DefaultRegMode.
    --     
    --     NOTE           : 
    --                      * Magnitude of the computed integer is to large. The 
    --                        input value is considered to large if after removing
    --                        leading 0's (1's for negative numbers)  the length
    --                        of the remaining vector is > IntegerBitLength-1.
    --                        (ie the machine integer length).
    --                      The error return value is INTEGER'LEFT.
    --
    --     Use            : 
    --                      VARIABLE vect : std_ulogic_vector ( 15 DOWNTO 0 );
    --
    --                      To_Integer ( vect, TwosComp );
    --     
    --     See Also       : To_StdLogicVector, To_Integer, To_TwosComp, To_OnesComp
    -------------------------------------------------------------------------------
    FUNCTION To_Integer   ( CONSTANT SrcReg     : IN std_ulogic_vector;
                            CONSTANT SrcRegMode : IN regmode_type 
                     -- synopsys synthesis_off
						      := DefaultRegMode 
                     -- synopsys synthesis_on
                          )  RETURN INTEGER IS
     BEGIN
	if (SrcRegMode = TwosComp) then
		return(To_Integer_FromTwosComp(SrcReg));
	else 
		return(To_Integer_FromUnsign(SrcReg));
	end if;
    END To_Integer;
    -------------------------------------------------------------------------------
    --     Function Name  : RegFill
    -- 1.7.4
    --     Overloading    : None
    --
    --     Purpose        : Fill an std_logic_vector with a given value
    --
    --     Parameters     :
    --                      SrcReg     - input  std_logic_vector, the  logic vector to be read.
    --                      DstLength  - input  NATURAL, length of the return logic vector.
    --                      FillVal    - input  std_ulogic, default is '0'
    --
    --     Result         : std_logic_vector of length DstLength
    --
    --     NOTE           : The length of the return logic vector  is specified by the
    --                      parameter 'DstLength'. The input logic vector will
    --                      be  filled with the FillVal
    --
    --     Use            :
    --                      VARIABLE vect : std_logic_vector ( 15 DOWNTO 0 );
    --                      vect := RegFill ( "00000101", 16, 'U');
    --
    --     See Also       : SignExtend
   -------------------------------------------------------------------------------
    FUNCTION RegFill   ( CONSTANT SrcReg      : IN std_logic_vector;
                         CONSTANT DstLength   : IN NATURAL;
                         CONSTANT FillVal     : IN std_ulogic  
        	-- synopsys synthesis_off
					         := '0'
	        -- synopsys synthesis_on
                       ) RETURN std_logic_vector IS
      VARIABLE result : std_logic_vector (DstLength - 1 DOWNTO 0);
      VARIABLE reg    : std_logic_vector (SrcReg'LENGTH - 1 DOWNTO 0);
      VARIABLE len    : integer;
    BEGIN
  	len := DstLength;
	if (FillVal = '0') Then
		result := RegFill_Zero(SrcReg, len);
                return result;
         else
		-- initializations
       	         result := (OTHERS => '0');
	         reg    := SrcReg;
        	-- synopsys translate_off
		--  null range check
	        IF (SrcReg'LENGTH = 0) THEN
			IF (DstLength = 0) THEN
        		        ASSERT FALSE
                		REPORT " RegFill --- input  has null range and" &
		                 " Destination also has null range. "
        		        SEVERITY ERROR;
                		RETURN result ;
		        ELSE
        		        ASSERT FALSE
                		REPORT " RegFill --- input  has null range"
	                	SEVERITY ERROR;
	        	        result := (OTHERS => FillVal);
			       	RETURN result ;
		        END IF;
 
       		ELSIF (DstLength = 0) THEN
	        	    ASSERT false
	        	    REPORT "RegFill --- Destination has null range "
		            SEVERITY ERROR;
        		    RETURN result;
 
	        ELSIF (DstLength <= SrcReg'LENGTH) THEN
                        -- no need to sign extend
        		   ASSERT (DstLength = SrcReg'LENGTH)
	        	   REPORT " RegFill ---  Destination length is less than source"
	        	   SEVERITY ERROR;
		           RETURN reg;        -- return the input data without any change

	       	ELSE
		      -- synopsys translate_on
	        	   result(SrcReg'LENGTH - 1 DOWNTO 0) := reg;
		        -- Fill the MSB's of result with the given fill value.
        		  For i IN DstLength - 1 DOWNTO SrcReg'LENGTH  Loop
	        	     result(i) := FillVal;
	        	  END LOOP;
	      -- synopsys translate_off
        	END IF;
	      -- synopsys translate_on
	      -- convert to X01
	        RETURN (To_X01(result));
 	end if;
    END RegFill;
    -------------------------------------------------------------------------------
    --     Function Name  : RegFill
    -- 
    --     Overloading    : None
    --
    --     Purpose        : Fill an std_ulogic_vector with a given value
    --
    --     Parameters     :
    --                      SrcReg     - input  std_ulogic_vector, the  logic vector to be read.
    --                      DstLength  - input  NATURAL, length of the return logic vector.
    --                      FillVal    - input  std_ulogic,  default is '0'
    --
    --     Result         : std_ulogic_vector of length DstLength
    --
    --     NOTE           : The length of the return logic vector  is specified by the
    --                      parameter 'DstLength'. The input logic vector will
    --                      be  filled with the FillVal
    --
    --     Use            :
    --                      VARIABLE vect : std_ulogic_vector ( 15 DOWNTO 0 );
    --                      vect := RegFill ( "00000101", 16, 'U');
    --
    --     See Also       : SignExtend
   -------------------------------------------------------------------------------
    FUNCTION RegFill   ( CONSTANT SrcReg      : IN std_ulogic_vector;
                         CONSTANT DstLength   : IN NATURAL;
                         CONSTANT FillVal     : IN std_ulogic
        	-- synopsys synthesis_off
					         := '0'
	        -- synopsys synthesis_on
                       ) RETURN std_ulogic_vector IS
	VARIABLE reslt  : std_logic_vector (DstLength - 1 DOWNTO 0);
	VARIABLE reg    : std_logic_vector (SrcReg'Length - 1 DOWNTO 0);
    BEGIN
	reg := To_StdLogicVector(SrcReg);
	reslt := RegFill (reg, DstLength, FillVal);
        return To_StdULogicVector(reslt);       
    END RegFill;
    -------------------------------------------------------------------------------
    --     Function Name  : RegFill
    -- 1.7.3
    --     Overloading    : None
    --
    --     Purpose        : Fill the most significant bits of a register with a given value
    --
    --     Parameters     :
    --                      SrcReg     - input  bit_vector, the vector to be read.
    --                      DstLength  - input  NATURAL, length of the return vector.
    --                      FillVal    - input  bit,  default is '0'
    --
    --     Result         : bit_vector
    --
    --     NOTE           : The length of the return bit vector  is specified by the
    --                      parameter 'DstLength'. The input bit vector will
    --                      be  filled with the FillVal
    --
    --     Use            :
    --                      VARIABLE vect : bit_vector ( 15 DOWNTO 0 );
    --                      vect := RegFill ( B"00000101", 16, '0');
    --                    or 
    --                      vect := RegFill ( B"00000101", 16);
    --
    --     See Also       : SignExtend
   -------------------------------------------------------------------------------
    FUNCTION RegFill   ( CONSTANT SrcReg      : IN bit_vector;
                         CONSTANT DstLength   : IN NATURAL;
                         CONSTANT FillVal     : IN bit  
        	-- synopsys synthesis_off
					         := '0'
	        -- synopsys synthesis_on
                       ) RETURN bit_vector IS
	VARIABLE reslt  : std_logic_vector (DstLength - 1 DOWNTO 0);
	VARIABLE reg    : std_logic_vector (SrcReg'Length - 1 DOWNTO 0);
	VARIABLE FVal   : std_ulogic;
    BEGIN
	reg := To_StdLogicVector(SrcReg);
        FVal := To_StdULogic(FillVal);
	reslt := RegFill (reg, DstLength, FVal);
        return To_BitVector(reslt);       
    END RegFill;
    -------------------------------------------------------------------------------
    --     Function Name  : SignExtend
    -- 1.7.1
    --     Overloading    : None
    --    
    --     Purpose        : Sign Extend a logic vector
    --     
    --     Parameters     : 
    --                      SrcReg     - input  std_logic_vector, the vector to be read.
    --                      DstLength  - input  NATURAL, length of the return vector.
    --                      SignBitPos - input  NATURAL, the position of the sign bit.
    --                                    for synthesis purpose it is the MSB (SrcReg'LEFT)
    --                      SrcRegMode    - input  regmode_type, indicating the format of
    --                                   the input std_logic_vector.   Default is TwosComp.
    --     
    --     Result         : std_logic_vector
    --
    --     NOTE           : The length of the return std_logic_vector  is specified by the
    --                      parameter 'DstLength'. The input std_logic_vector will 
    --                      be sign extended. 
    --
    --                      For synthesis purpose SignBitPos argument is ignored and the MSB 
    --                      ( ie. SrcReg'Left) is considered as a sign bit position.
    --
    --     Use            :
    --                      VARIABLE vect : std_logic_vector ( 15 DOWNTO 0 );
    --                      vect := SignExtend ( "11111101", 16,TwosComp ); -- set to -4
    --     
    --     See Also       : RegFill
    -------------------------------------------------------------------------------
    FUNCTION SignExtend   ( CONSTANT SrcReg      : IN std_logic_vector;
                            CONSTANT DstLength   : IN NATURAL;
                            CONSTANT SignBitPos  : IN NATURAL;
                            CONSTANT SrcRegMode  : IN regmode_type
                     -- synopsys synthesis_off
						      := DefaultRegMode 
                     -- synopsys synthesis_on
                          ) RETURN std_logic_vector IS
	variable len : integer;
    Begin
	len := DstLength;

	if (SrcRegMode = TwosComp) THEN     
		return ( SignExtend_TwosComp(SrcReg, len));
	else
		return ( RegFill_Zero(SrcReg, len));
	end if;
   
    END SignExtend;
    -------------------------------------------------------------------------------
    --     Function Name  : SignExtend
    -- 1.7.1
    --     Overloading    : None
    --    
    --     Purpose        : Sign Extend a logic vector
    --     
    --     Parameters     : 
    --                      SrcReg     - input  std_ulogic_vector, the vector to be read.
    --                      DstLength  - input  NATURAL, length of the return vector.
    --                      SignBitPos - input  NATURAL, the position of the sign bit.
    --                                    for synthesis purpose it is the MSB (SrcReg'LEFT)
    --                      SrcRegMode    - input  regmode_type, indicating the format of
    --                                   the input std_ulogic_vector.   Default is TwosComp.
    --     
    --     Result         : std_ulogic_vector
    --
    --     NOTE           : The length of the return std_ulogic_vector  is specified by the
    --                      parameter 'DstLength'. The input std_ulogic_vector will 
    --                      be sign extended. 
    --
    --                      For synthesis purpose SignBitPos argument is ignored and the MSB 
    --                      ( ie. SrcReg'Left) is considered as a sign bit position.
    --
    --     Use            :
    --                      VARIABLE vect : std_ulogic_vector ( 15 DOWNTO 0 );
    --                      vect := SignExtend ( "11111101", 16,7,TwosComp ); -- set to -4
    --     
    --     See Also       : RegFill
    -------------------------------------------------------------------------------
    FUNCTION SignExtend   ( CONSTANT SrcReg      : IN std_ulogic_vector;
                            CONSTANT DstLength   : IN NATURAL;
                            CONSTANT SignBitPos  : IN NATURAL;
                            CONSTANT SrcRegMode  : IN regmode_type
                     -- synopsys synthesis_off
						      := DefaultRegMode 
                     -- synopsys synthesis_on
                          ) RETURN std_ulogic_vector IS
	VARIABLE reslt_copy : std_logic_vector (DstLength - 1 downto 0);     
	VARIABLE reg    : std_logic_vector (SrcReg'Length - 1 DOWNTO 0);
    BEGIN
	reg := To_StdLogicVector(SrcReg);
	reslt_copy := SignExtend( reg, DstLength, SignBitPos, SrcRegMode);
        return To_StdULogicVector(reslt_copy);         
    END SignExtend;
    -------------------------------------------------------------------------------
    --     Function Name  : SignExtend
    -- 1.7.1
    --     Overloading    : None
    --    
    --     Purpose        : Sign Extend a bit vector
    --     
    --     Parameters     : 
    --                      SrcReg     - input  bit_vector, the vector to be read.
    --                      DstLength  - input  NATURAL, length of the return vector.
    --                      SignBitPos - input  NATURAL, the position of the sign bit.
    --                                    for synthesis purpose it is the MSB (SrcReg'LEFT)
    --                      SrcRegMode    - input  regmode_type, indicating the format of
    --                                   the input bit_vector.   Default is TwosComp.
    --     
    --     Result         : bit_vector, the extened bit vector
    --
    --     NOTE           : The length of the return bit vector  is specified by the
    --                      parameter 'DstLength'. The input bit vector will 
    --                      be sign extended. 
    --
    --                      For synthesis purpose SignBitPos argument is ignored and the MSB 
    --                      ( ie. SrcReg'Left) is considered as a sign bit position.
    --     Use            :
    --                      VARIABLE vect : bit_vector ( 15 DOWNTO 0 );
    --                      vect := SignExtend ( B"11111101", 16, 7,TwosComp ); -- set to -4
    --     
    -------------------------------------------------------------------------------
    FUNCTION SignExtend   ( CONSTANT SrcReg      : IN bit_vector;
                            CONSTANT DstLength   : IN NATURAL;
                            CONSTANT SignBitPos  : IN NATURAL;
                            CONSTANT SrcRegMode  : IN regmode_type
                     -- synopsys synthesis_off
						      := DefaultRegMode 
                     -- synopsys synthesis_on
                          ) RETURN bit_vector IS
	VARIABLE reslt_copy : std_logic_vector (DstLength - 1 downto 0);     
	VARIABLE reg    : std_logic_vector (SrcReg'Length - 1 DOWNTO 0);
    BEGIN
	reg := To_StdLogicVector(SrcReg);
	reslt_copy := SignExtend( reg, DstLength, SignBitPos, SrcRegMode);
        return To_BitVector(reslt_copy);         
    END SignExtend;
    -------------------------------------------------------------------------------
    --     Procedure Name : RegAbs
    -- 1.6.9
    --     Overloading    : Procedure .
    --
    --     Purpose        : converts  std_logic_vector into an absolute value.
    --
    --     Parameters     :
    --                      result     - input-output  std_logic_vector, 
    --                      SrcReg     - input  std_logic_vector, the vector to be read.
    --                      SrcRegMode - input  regmode_type, indicating the format of
    --                                the input std_logic_vector.   Default is TwosComp.
    --
    --
    --     Use            :
    --                      VARIABLE reslt, vect : std_logic_vector ( 15 DOWNTO 0 );
    --
    --                       RegAbs ( reslt,  vect, TwosComp );
    --
    -------------------------------------------------------------------------------
    PROCEDURE RegAbs  ( VARIABLE result     : INOUT std_logic_vector;
                        CONSTANT SrcReg     : IN std_logic_vector;
                        CONSTANT SrcRegMode : IN regmode_type 
                     -- synopsys synthesis_off
						      := DefaultRegMode 
                     -- synopsys synthesis_on
                      ) IS
       VARIABLE result_copy : std_logic_vector (result'LENGTH - 1 DOWNTO 0);
       VARIABLE reg          : std_logic_vector (SrcReg'LENGTH - 1 DOWNTO 0);
    --
    BEGIN
    --
    	result_copy := result;  
        reg         := SrcReg;
  -- synopsys translate_off
    --   Null range check
    --   if result vector is a null range
       IF ( result'LENGTH = 0) THEN
             ASSERT false
             REPORT " RegAbs ---  Destination has null range. "
             SEVERITY ERROR;
             RETURN;
     -- if the input is of null range 
       ELSIF (SrcReg'LENGTH = 0) THEN
             ASSERT false
             REPORT " RegAbs --- input has null range "
             SEVERITY ERROR;
             result_copy := (OTHERS => '0');
             result := result_copy;
             RETURN;
        END IF;
  -- synopsys translate_on
        IF (SrcRegMode = TwosComp) THEN  
              -- if a negative value, take two's comp it
              -- will become absolute
               IF (reg(SrcReg'LENGTH - 1) /= '0') THEN
                   -- if not largest negative number
                     IF ( No_One(reg(SrcReg'LENGTH - 2 downto 0))) THEN
                        -- synopsys translate_off
                            ASSERT false
                            REPORT "RegAbs  --  2's comp vector  cannot be converted. "
                            SEVERITY Error;   
                        -- synopsys translate_on
                       ELSE
                             reg := RegNegate ( reg, TwosComp);
                       END IF;
                END IF;
          
          ELSE  -- Unsigned  
              null;
          END IF;
          result_copy(SrcReg'LENGTH - 1 downto 0) := reg;
          result := result_copy;
         RETURN;
    END RegAbs;
    -------------------------------------------------------------------------------
    --     Procedure Name : RegAbs
    -- 
    --     Overloading    : Procedure .
    --
    --     Purpose        : converts  std_ulogic_vector into an absolute value.
    --
    --     Parameters     :
    --                      result     - input- output  std_ulogic_vector, 
    --                      SrcReg     - input  std_ulogic_vector, the vector to be read.
    --                      SrcRegMode - input  regmode_type, indicating the format of
    --                                the input std_ulogic_vector.   Default is TwosComp.
    --
    --
    --     Use            :
    --                      VARIABLE reslt, vect : std_ulogic_vector ( 15 DOWNTO 0 );
    --
    --                       RegAbs ( reslt,  vect, TwosComp );
    --
    -------------------------------------------------------------------------------
    PROCEDURE RegAbs  ( VARIABLE result     : INOUT std_ulogic_vector;
                        CONSTANT SrcReg     : IN std_ulogic_vector;
                        CONSTANT SrcRegMode : IN regmode_type 
                     -- synopsys synthesis_off
						      := DefaultRegMode 
                     -- synopsys synthesis_on
                      ) IS
       VARIABLE reslt_copy  : std_logic_vector (result'LENGTH - 1 DOWNTO 0);
       VARIABLE reg_copy    : std_logic_vector (SrcReg'LENGTH - 1 DOWNTO 0);
    BEGIN
        reg_copy := To_StdLogicVector(SrcReg);
	RegAbs(reslt_copy, reg_copy, SrcRegMode);
        result := To_StdULogicVector(reslt_copy);         
        return;
    END RegAbs;
    -------------------------------------------------------------------------------
    --     Function Name  : RegAbs
    --
    --     Procedure Name : RegAbs
    -- 1.6.10
    --     Overloading    : Procedure .
    --
    --     Purpose        : converts  bit_vectors into an absolute value.
    --
    --     Parameters     :
    --                      result     - input-output  bit_vector, 
    --                      SrcReg     - input  bit_vector, the vector to be read.
    --                      SrcRegMode - input  regmode_type, indicating the format of
    --                                the input bit_vector.   Default is TwosComp.
    --
    --
    --     Use            :
    --                      VARIABLE reslt, vect : bit_vector ( 15 DOWNTO 0 );
    --
    --                       RegAbs ( reslt,  vect, TwosComp );
    --
    -------------------------------------------------------------------------------
    PROCEDURE RegAbs  ( VARIABLE result     : INOUT bit_vector;
                        CONSTANT SrcReg     : IN bit_vector;
                        CONSTANT SrcRegMode : IN regmode_type
                     -- synopsys synthesis_off
						      := DefaultRegMode 
                     -- synopsys synthesis_on
                      ) IS
       VARIABLE reslt_copy  : std_logic_vector (result'LENGTH - 1 DOWNTO 0);
       VARIABLE reg_copy    : std_logic_vector (SrcReg'LENGTH - 1 DOWNTO 0);
    BEGIN
        reg_copy := To_StdLogicVector(SrcReg);
	RegAbs(reslt_copy, reg_copy, SrcRegMode);
        result := To_BitVector(reslt_copy);         
        return;
    END RegAbs;
--+-----------------------------------------------------------------------------
--|     Function Name  : RegAdd
--|
--|     Overloading    : None
--|
--|     Purpose        : Addition of logic vectors.
--|
--|     Parameters     :
--|                      result     - output std_logic_vector, the computed sum
--|                      carry_out  - output std_logic,
--|                      overflow   - output std_logic,
--|                      addend     - input  std_logic_vector,
--|                      augend     - input  std_logic_vector,
--|                      carry_in   - input  std_logic, carry into the LSB.
--|                      SrcRegMode - input  regmode_type, indicating the format of
--|                              the input std_logic_vector.   Default is TwosComp.
--|     NOTE           :
--|                      The inputs may be of any length and may be of differing
--|                      lengths.
--|  
--|                    For Synthesis:
--|                      Result is computed with length N (where
--|                      N is the greater of the input vector lengths).
--|                      It is assumed that user will provide result length equal
--|                      to the length of the greater of addend and augend. 
--|                      No error checking has been performed.
--|     Use            :
--|                      VARIABLE x, y, sum : std_logic_vector ( 15 DOWNTO 0);
--|                      VARIABLE carry_in, carry_out , ovf: std_ulogic;
--| 
--|                      RegAdd ( sum, carry_out, ovf,x, y, carry_in, TwosComp );
--| 
--|     See Also       : RegAdd, RegSub, RegMult, RegDiv, RegInc, RegDec, RegNegate
--|-----------------------------------------------------------------------------
    PROCEDURE RegAdd  ( VARIABLE result     : INOUT std_logic_vector;
                        VARIABLE carry_out  : OUT std_ulogic;
                        VARIABLE overflow   : OUT std_ulogic;
                        CONSTANT addend     : IN std_logic_vector;
                        CONSTANT augend     : IN std_logic_vector;
                        CONSTANT carry_in   : IN std_ulogic;
                        CONSTANT SrcRegMode : IN regmode_type
                 -- synopsys synthesis_off
					           := DefaultRegMode 
                 -- synopsys synthesis_on
                      ) IS

	CONSTANT reslen       : INTEGER := MAXIMUM ( addend'LENGTH, augend'LENGTH );
	VARIABLE a, b, r      : STD_LOGIC_VECTOR ( reslen - 1 DOWNTO 0 );
	VARIABLE  result_copy : STD_LOGIC_VECTOR ( result'Length - 1 DOWNTO 0 );
     BEGIN 
      -- synopsys translate_off
      --   Null range check
      --   if result vector is a null range
        IF ( result'LENGTH = 0) THEN
             ASSERT false
             REPORT " RegAdd ---  Destination has null range. "
             SEVERITY ERROR;
             RETURN;
      --   if addend or augned or both have null range no need to add
        ELSIF (addend'LENGTH = 0) AND (augend'LENGTH = 0) THEN
             ASSERT false
             REPORT " RegAdd --- both addend  and augend has null range "
             SEVERITY ERROR;
             result_copy :=  (OTHERS => '0');
             IF (carry_in = '1') THEN
                 IF (SrcRegMode = TwosComp OR SrcRegMode = Unsigned) THEN
                        result_copy(0) := '1';
                 END IF;
             END IF;
             result := result_copy; 
             carry_out := '0';
             overflow := '0';       
             RETURN;      
        END IF;
      -- synopsys translate_on
      -- if one of the addend or augend is null 
        IF (addend'LENGTH = 0) THEN
      -- synopsys translate_off
             ASSERT false
             REPORT " RegAdd --- addend has null range "
             SEVERITY ERROR;
      -- synopsys translate_on
             a :=  ( OTHERS => '0');     -- treat it as	zero's            
             b := augend;

        ELSIF (augend'LENGTH = 0) THEN 
      -- synopsys translate_off
             ASSERT false
             REPORT " RegAdd ---  augend has null range "
             SEVERITY ERROR;
      -- synopsys translate_on
             b :=  (OTHERS => '0');                 
             a := addend;
                 -- inputs are  not null so sign extend them to the same length.  
        ELSE
             a := SignExtend(addend , reslen, addend'LEFT, SrcRegMode);
             b := SignExtend(augend , reslen, augend'LEFT, SrcRegMode);

        END IF;	
       -- Compute the add operation
	if (SrcRegMode = TwosComp) Then
		Add_TwosComp_VHDL_TECH (result,carry_out, overflow, a, b, carry_in); 
        else
		Add_Unsigned_VHDL_TECH (result,carry_out, overflow, a, b, carry_in);
        end if;
        RETURN;
     END RegAdd;
--+-----------------------------------------------------------------------------
--|     Function Name  : RegAdd
--|
--|     Overloading    : None
--|
--|     Purpose        : Addition of logic vectors.
--|
--|     Parameters     :
--|                      result     - output std_ulogic_vector, the computed sum
--|                      carry_out  - output std_logic,
--|                      overflow   - output std_logic,
--|                      addend     - input  std_ulogic_vector,
--|                      augend     - input  std_ulogic_vector,
--|                      carry_in   - input  std_logic, carry into the LSB.
--|                      SrcRegMode - input  regmode_type, indicating the format of
--|                             the input std_ulogic_vector.   Default is TwosComp.
--|     NOTE           :
--|                      The inputs may be of any length and may be of differing
--|                      lengths.
--|  
--|                    For Synthesis:
--|                      Result is computed with length N (where
--|                      N is the greater of the input vector lengths).
--|                      It is assumed that user will provide result length equal
--|                      to the length of the greater of addend and augend. 
--|                      No error checking has been performed.
--|     Use            :
--|                      VARIABLE x, y, sum : std_ulogic_vector ( 15 DOWNTO 0);
--|                      VARIABLE carry_in, carry_out , ovf: std_ulogic;
--| 
--|                      RegAdd ( sum, carry_out, ovf,x, y, carry_in, TwosComp );
--| 
--|     See Also       : RegAdd, RegSub, RegMult, RegDiv, RegInc, RegDec, RegNegate
--|-----------------------------------------------------------------------------
    PROCEDURE RegAdd  ( VARIABLE result     : INOUT std_ulogic_vector;
                        VARIABLE carry_out  : OUT std_ulogic;
                        VARIABLE overflow   : OUT std_ulogic;
                        CONSTANT addend     : IN std_ulogic_vector;
                        CONSTANT augend     : IN std_ulogic_vector;
                        CONSTANT carry_in   : IN std_ulogic;
                        CONSTANT SrcRegMode : IN regmode_type
                 -- synopsys synthesis_off
					           := DefaultRegMode 
                 -- synopsys synthesis_on
                      ) IS
	VARIABLE  reslt_copy : STD_LOGIC_VECTOR ( result'Length - 1 DOWNTO 0 );
	VARIABLE  a          : STD_LOGIC_VECTOR ( addend'Length - 1 DOWNTO 0 );
	VARIABLE  b          : STD_LOGIC_VECTOR ( augend'Length - 1 DOWNTO 0 );
     BEGIN 
	a := To_StdLogicVector(addend);
        b := To_StdLogicVector(augend);
        RegAdd(reslt_copy, carry_out, overflow, a, b, carry_in, SrcRegMode); 
        result := To_StdULogicVector(reslt_copy);
        return;
     END RegAdd;
--+-----------------------------------------------------------------------------
--|     Function Name  : RegAdd
--|
--|     Overloading    : None
--|
--|     Purpose        : Addition of BIT_VECTORS.
--|
--|     Parameters     :
--|                      result     - input-output BIT_VECTOR, the computed sum
--|                      carry_out  - output BIT,
--|                      overflow   - output BIT, overflow condition
--|                      addend     - input  BIT_VECTOR,
--|                      augend     - input  BIT_VECTOR,
--|                      carry_in   - input  BIT,  
--|                      SrcRegMode - input  regmode_type, indicating the format of
--|                                the input BIT_VECTOR.   Default is TwosComp.
--|     NOTE           :
--|                      The inputs may be of any length and may be of differing
--|                      lengths.
--|
--|                    For Synthesis:
--|                      Result is computed with length N (where
--|                      N is the greater of the input vector lengths).
--|                      It is assumed that user will provide result length equal
--|                      to the length of the greater of addend and augend. 
--|                      No error checking has been performed.
--|     Use            :
--|                      VARIABLE x, y, sum : BIT_VECTOR ( 15 DOWNTO 0);
--|                      VARIABLE carry_in, carry_out , ovf: BIT;
--| 
--|                      RegAdd ( sum, carry_out, ovf,x, y, carry_in, UnSigned );
--| 
--|     See Also       : RegAdd, RegSub, RegMult, RegDiv, RegInc, RegDec, RegNegate
--|-----------------------------------------------------------------------------
    PROCEDURE RegAdd  ( VARIABLE result     : INOUT BIT_VECTOR;
                        VARIABLE carry_out  : OUT BIT;
                        VARIABLE overflow   : OUT BIT;
                        CONSTANT addend     : IN BIT_VECTOR;
                        CONSTANT augend     : IN BIT_VECTOR;
                        CONSTANT carry_in   : IN BIT;
                        CONSTANT SrcRegMode : IN regmode_type 
                 -- synopsys synthesis_off
                                                        := DefaultRegMode 
                 -- synopsys synthesis_on
                      ) IS
	VARIABLE  reslt_copy   : std_logic_vector ( result'Length - 1 DOWNTO 0 );
        VARIABLE  c_out, ovflo : Std_ulogic;
        VARIABLE  c_in         : Std_ulogic;
	VARIABLE  a            : STD_LOGIC_VECTOR ( addend'Length - 1 DOWNTO 0 );
	VARIABLE  b            : STD_LOGIC_VECTOR ( augend'Length - 1 DOWNTO 0 );
     BEGIN 
	a := To_StdLogicVector(addend);
        b := To_StdLogicVector(augend);
        c_in := To_StdULogic(carry_in);
        RegAdd(reslt_copy, c_out, ovflo, a, b, c_in, SrcRegMode); 
        result    := To_BitVector(reslt_copy);
        carry_out := To_Bit(c_out);
        overflow  := To_Bit(ovflo);
        return;
    END RegAdd;
--+-----------------------------------------------------------------------------
--|     Function Name  : RegSub
--|    
--|     Overloading    : None
--|
--|     Purpose        : Subtraction of logic vectors.
--|                       ( result = minuend - subtrahend )
--|
--|     Parameters     :
--|                      result     - input_output std_logic_vector, the computed diff
--|                      borrow_out - output std_logic,
--|                      overflow   - output std_logic, overflow condition
--|                      minuend    - input  std_logic_vector,
--|                      subtrahend - input  std_logic_vector,
--|                      borrow_in  - input  std_logic, borrow from the LSB
--|                      SrcRegMode - input  regmode_type, indicating the format of
--|                               the input std_logic_vector.   Default is TwosComp.
--|     NOTE           :
--|                      The inputs may be of any length and may be of differing
--|                      lengths.
--|
--|                      A temporary result is computed with length N (where
--|                      N is the greater of the input vector lengths).
--|     Use            :
--|                      VARIABLE x, y, diff : std_logic_vector ( 15 DOWNTO 0);
--|                      VARIABLE n_borrow, borrow_in : std_ulogic;
--|
--|                      RegSub ( diff, n_borrow, x, y, borrow_in, UnSigned );
--|
--|     See Also       : RegAdd, RegSub, RegMult, RegDiv, RegInc, RegDec, RegNegate
--|-----------------------------------------------------------------------------
    PROCEDURE RegSub  ( VARIABLE result     : INOUT std_logic_vector;
                        VARIABLE borrow_out : OUT std_ulogic;
                        VARIABLE overflow   : OUT std_ulogic;
                        CONSTANT minuend    :  IN std_logic_vector;
                        CONSTANT subtrahend :  IN std_logic_vector;
                        CONSTANT borrow_in  :  IN std_ulogic
                 -- synopsys synthesis_off
                                                       := '0'
                 -- synopsys synthesis_on
                                                               ;
                        CONSTANT SrcRegMode :  IN regmode_type
                 -- synopsys synthesis_off
                                                      := DefaultRegMode 
                 -- synopsys synthesis_on
                      ) IS
      CONSTANT reslen       : INTEGER := MAXIMUM (minuend'LENGTH, subtrahend'LENGTH);
      VARIABLE a, b, r      : STD_LOGIC_VECTOR ( reslen - 1 DOWNTO 0 );
      VARIABLE reslt_copy   : STD_LOGIC_VECTOR ( result'length-1 downto 0);
    BEGIN
    -- synopsys translate_off
     --   Null range check
     --   if result vector is a null range
       IF ( result'LENGTH = 0) THEN
             ASSERT false
             REPORT " RegSub ---  Destination has null range. " &
                    " cannot save result. "
             SEVERITY ERROR;
             RETURN;

     --   if both minuend and subtrahend  have null range no need to subtract
       ELSIF  (minuend'LENGTH = 0) AND (subtrahend'LENGTH = 0) THEN
             ASSERT false
             REPORT " RegSub --- both minuend and subtrahend has null range "
             SEVERITY ERROR;
             reslt_copy :=  (OTHERS => '0');
             borrow_out := '0';
             IF (borrow_in /= '0') THEN
                 IF (SrcRegMode = TwosComp OR SrcRegMode = Unsigned) THEN
                        reslt_copy := (OTHERS =>'1');
                        borrow_out := '1';
                 END IF;
             END IF;
             result := reslt_copy;
             overflow := '0';
             RETURN;
       END IF;
     -- synopsys translate_on
     -- if one of the minuend or subtrahend is null
       IF (minuend'LENGTH = 0) THEN
    -- synopsys translate_off
             ASSERT false
             REPORT " RegSub --- minuend has null range "
             SEVERITY ERROR;
    -- synopsys translate_on
             a :=  ( OTHERS => '0');     -- treat it as zero's
             b :=  subtrahend ;
 
       ELSIF (subtrahend'LENGTH = 0) THEN
    -- synopsys translate_off
             ASSERT false
             REPORT " RegSub ---  subtrahend has null range "
             SEVERITY ERROR;
    -- synopsys translate_on
             b :=  (OTHERS => '0');
             a := minuend ;
  
                 -- inputs are  not null so sign extend them to the same length.
       ELSE
             a := SignExtend(minuend , reslen, minuend'LEFT, SrcRegMode);
             b := SignExtend(subtrahend , reslen, subtrahend'LEFT, SrcRegMode);
 
       END IF;
       -- compute the subtraction
	if (SrcRegMode = TwosComp) Then
		Sub_TwosComp_VHDL_TECH (result,borrow_out, overflow, a, b, borrow_in); 
        else
		Sub_Unsigned_VHDL_TECH (result,borrow_out, overflow, a, b, borrow_in);
        end if;
	return;
     END RegSub;
--+-----------------------------------------------------------------------------
--|     Function Name  : RegSub
--|    
--|     Overloading    : None
--|
--|     Purpose        : Subtraction of ulogic vectors.
--|                       ( result = minuend - subtrahend )
--|
--|     Parameters     :
--|                      result     - input_output std_ulogic_vector, the computed diff
--|                      borrow_out - output std_logic,
--|                      overflow   - output std_logic, overflow condition
--|                      minuend    - input  std_ulogic_vector,
--|                      subtrahend - input  std_ulogic_vector,
--|                      borrow_in  - input  std_logic, borrow from the LSB
--|                      SrcRegMode - input  regmode_type, indicating the format of
--|                              the input std_ulogic_vector.   Default is TwosComp.
--|     NOTE           :
--|                      The inputs may be of any length and may be of differing
--|                      lengths.
--|
--|                      A temporary result is computed with length N (where
--|                      N is the greater of the input vector lengths).
--|     Use            :
--|                      VARIABLE x, y, diff : std_ulogic_vector ( 15 DOWNTO 0);
--|                      VARIABLE n_borrow, borrow_in : std_ulogic;
--|
--|                      RegSub ( diff, n_borrow, x, y, borrow_in, UnSigned );
--|
--|     See Also       : RegAdd, RegSub, RegMult, RegDiv, RegInc, RegDec, RegNegate
--|-----------------------------------------------------------------------------
    PROCEDURE RegSub  ( VARIABLE result     : INOUT std_ulogic_vector;
                        VARIABLE borrow_out : OUT std_ulogic;
                        VARIABLE overflow   : OUT std_ulogic;
                        CONSTANT minuend    :  IN std_ulogic_vector;
                        CONSTANT subtrahend :  IN std_ulogic_vector;
                        CONSTANT borrow_in  :  IN std_ulogic 
                 -- synopsys synthesis_off
                                                       := '0'
                 -- synopsys synthesis_on
                                                               ;
                        CONSTANT SrcRegMode :  IN regmode_type
                 -- synopsys synthesis_off
                                                      := DefaultRegMode 
                 -- synopsys synthesis_on
                      ) IS
        VARIABLE reslt_copy    : STD_LOGIC_VECTOR ( result'length-1 downto 0);
	VARIABLE  a            : STD_LOGIC_VECTOR ( minuend'Length - 1 DOWNTO 0 );
	VARIABLE  b            : STD_LOGIC_VECTOR (subtrahend'Length - 1 DOWNTO 0 );
     BEGIN 
	a := To_StdLogicVector(minuend);
        b := To_StdLogicVector(subtrahend);
	RegSub(reslt_copy, borrow_out, overflow, a, b, borrow_in, SrcRegMode); 
	result := To_StdULogicVector(reslt_copy);
	return;
    END RegSub;
--+-----------------------------------------------------------------------------
--|     Function Name  : RegSub
--|    
--|     Overloading    : None
--|
--|     Purpose        : Subtraction of BIT_VECTORS.
--|                       ( result = minuend - subtrahend )
--|
--|     Parameters     :
--|                      result     - input-output BIT_VECTOR, the computed sum
--|                      borrow_out - output BIT,
--|                      overflow   - output BIT, overflow condition
--|                      minuend - input  BIT_VECTOR,
--|                      subtrahend - input  BIT_VECTOR,
--|                      borrow_in  - input  BIT, borrow from the LSB
--|                      SrcRegMode - input  regmode_type, indicating the format of
--|                                the input BIT_VECTOR.   Default is TwosComp.
--|     NOTE           :
--|                      The inputs may be of any length and may be of differing
--|                      lengths.
--|
--|                      A temporary result is computed with length N (where
--|                      N is the greater of the input vector lengths).
--|     Use            :
--|                      VARIABLE x, y, diff : BIT_VECTOR ( 15 DOWNTO 0);
--|                      VARIABLE n_borrow, borrow_in : BIT;
--|
--|                      RegSub ( diff, n_borrow, x, y, borrow_in, UnSigned );
--|
--|     See Also       : RegAdd, RegSub, RegMult, RegDiv, RegInc, RegDec, RegNegate
--|-----------------------------------------------------------------------------
    PROCEDURE RegSub  ( VARIABLE result     : INOUT BIT_VECTOR;
                        VARIABLE borrow_out : OUT BIT;
                        VARIABLE overflow   : OUT BIT;
                        CONSTANT minuend    :  IN BIT_VECTOR;
                        CONSTANT subtrahend :  IN BIT_VECTOR;
                        CONSTANT borrow_in  :  IN BIT 
                 -- synopsys synthesis_off
                                                       := '0'
                 -- synopsys synthesis_on
                                                               ;
                        CONSTANT SrcRegMode :  IN regmode_type
                 -- synopsys synthesis_off

                                                      := DefaultRegMode 
                 -- synopsys synthesis_on
                      ) IS
        VARIABLE reslt_copy    : std_logic_vector( result'length-1 downto 0);
        VARIABLE b_out, undflo, b_in : std_ulogic;
	VARIABLE  a            : STD_LOGIC_VECTOR ( minuend'Length - 1 DOWNTO 0 );
	VARIABLE  b            : STD_LOGIC_VECTOR (subtrahend'Length - 1 DOWNTO 0 );
     BEGIN 
	a    := To_StdLogicVector(minuend);
        b    := To_StdLogicVector(subtrahend);
        b_in := To_StdUlogic(borrow_in);
	RegSub(reslt_copy, b_out, undflo, a, b, b_in, SrcRegMode); 

	result := To_BitVector(reslt_copy);
	borrow_out := To_Bit(b_out);
	overflow  := To_Bit(undflo);
	return;
    END RegSub;
--+-----------------------------------------------------------------------------
--|     Function Name  : RegMult
--|
--|     Overloading    : None
--|
--|     Purpose        : Multiplication of STD_LOGIC_VECTORS.
--|
--|     Parameters     :
--|                      result       - output STD_LOGIC_VECTOR, the computed product
--|                      overflow     - output STD_ULOGIC, overflow condition
--|                      multiplicand - input STD_LOGIC_VECTOR,
--|                      multiplier   -  input STD_LOGIC_VECTOR,
--|                      SrcRegMode   - input  regmode_type, indicating the format 
--|                                     of the input STD_LOGIC_VECTOR.   Default is 
--|                                     DefaultRegMode which is set to TwosComp.
--|     NOTE           :
--|                      The inputs may be of any length and may be of differing
--|                      lengths.
--|
--|    Algorithm       : The multiplication is carried out as follows:
--|
--|                      1) Determine sign of result based on sign of 
--|                         multiploicand and sign  of multiplier.
--|
--|                      2) Convert the multiplicand amd multiplier to Unsigned 
--|                         representation.
--|                      
--|                      3) Perform multiplication based on add and shift algorithm.
--|
--|                      4) Convert the result to the SrcRegMode with appropropriate sign
--|
--|     Result         :
--|                     A  temporary result is computed with length N+M (where
--|                      N,M are the lengths of the multiplicand and multiplier)
--|                      by calling local function Mult_TwosComp or Mult_Unsigned
--|                       
--|                      This computed value is extended or truncated to match
--|                      the width of 'result'. If truncated, the low order bits
--|                      are returned.
--|
--|                      The parameter 'overflow' is set to '1' if the product of the
--|                      two inputs is too large to fit in the parameter result.
--|     Use            :
--|                      VARIABLE x, y, prod : STD_LOGIC_VECTOR ( 15 DOWNTO 0);
--|                      VARIABLE ovfl : STD_ULOGIC;
--|
--|                      RegMult ( prod, ovfl, x, y, TwosComp );
--|
--|     See Also       : RegAdd, RegSub, RegMult, RegDiv, RegInc, RegDec, RegNegate
--|-----------------------------------------------------------------------------
    PROCEDURE RegMult ( VARIABLE result       : OUT STD_LOGIC_VECTOR;
                        VARIABLE overflow     : OUT STD_ULOGIC;
                        CONSTANT multiplicand : IN STD_LOGIC_VECTOR;
                        CONSTANT multiplier   : IN STD_LOGIC_VECTOR;
                        CONSTANT SrcRegMode   : IN regmode_type
                 -- synopsys synthesis_off
                                                      := DefaultRegMode 
                 -- synopsys synthesis_on
                      ) IS
     Begin
	if (SrcRegMode = TwosComp) THEN
		RegMult_TwosComp(result, overflow, multiplicand, multiplier);
	else 
		RegMult_Unsigned(result, overflow, multiplicand, multiplier);
	end if;
        RETURN;
    END RegMult;
--+-----------------------------------------------------------------------------
--|     Function Name  : RegMult
--|
--|     Overloading    : None
--|
--|     Purpose        : Multiplication of STD_ULOGIC_VECTORS.
--|
--|     Parameters     :
--|                      result       - output STD_ULOGIC_VECTOR, the computed product
--|                      overflow     - output STD_ULOGIC, overflow condition
--|                      multiplicand - input STD_ULOGIC_VECTOR,
--|                      multiplier   -  input STD_ULOGIC_VECTOR,
--|                      SrcRegMode   - input  regmode_type, indicating the format 
--|                                     of the input STD_ULOGIC_VECTOR.   Default is 
--|                                     DefaultRegMode which is set to TwosComp.
--|     NOTE           :
--|                      The inputs may be of any length and may be of differing
--|                      lengths.
--|
--|    Algorithm       : The multiplication is carried out as follows:
--|
--|                      1) Determine sign of result based on sign of 
--|                         multiploicand and sign  of multiplier.
--|
--|                      2) Convert the multiplicand amd multiplier to Unsigned 
--|                         representation.
--|                      
--|                      3) Perform multiplication based on add and shift algorithm.
--|
--|                      4) Convert the result to the SrcRegMode with appropropriate sign
--|
--|     Result         :
--|                     A  temporary result is computed with length N+M (where
--|                      N,M are the lengths of the multiplicand and multiplier)
--|                      by calling local function Mult_TwosComp or Mult_Unsigned
--|                       
--|                      This computed value is extended or truncated to match
--|                      the width of 'result'. If truncated, the low order bits
--|                      are returned.
--|
--|                      The parameter 'overflow' is set to '1' if the product of the
--|                      two inputs is too large to fit in the parameter result.
--|     Use            :
--|                      VARIABLE x, y, prod : STD_ULOGIC_VECTOR ( 15 DOWNTO 0);
--|                      VARIABLE ovfl : STD_ULOGIC;
--|
--|                      RegMult ( prod, ovfl, x, y, TwosComp );
--|
--|     See Also       : RegAdd, RegSub, RegMult, RegDiv, RegInc, RegDec, RegNegate
--|-----------------------------------------------------------------------------
    PROCEDURE RegMult ( VARIABLE result       : OUT STD_ULOGIC_VECTOR;
                        VARIABLE overflow     : OUT STD_ULOGIC;
                        CONSTANT multiplicand : IN STD_ULOGIC_VECTOR;
                        CONSTANT multiplier   : IN STD_ULOGIC_VECTOR;
                        CONSTANT SrcRegMode   : IN regmode_type
                 -- synopsys synthesis_off
                                                      := DefaultRegMode 
                 -- synopsys synthesis_on
                      ) IS

	VARIABLE reslt : STD_LOGIC_VECTOR (result'length - 1 downto 0);
	VARIABLE  a    : STD_LOGIC_VECTOR ( multiplicand'Length - 1 DOWNTO 0 );
	VARIABLE  b    : STD_LOGIC_VECTOR (multiplier'Length - 1 DOWNTO 0 );
     BEGIN 
	a    := To_StdLogicVector(multiplicand);
        b    := To_StdLogicVector(multiplier);
	RegMult(reslt, overflow, a, b, SrcRegMode);
        result := To_StdULogicVector(reslt);
        RETURN;
    END RegMult;
--+-----------------------------------------------------------------------------
--|     Function Name  : RegMult
--|
--|     Overloading    : None
--|
--|     Purpose        : Multiplication of BIT_VECTORS.
--|
--|     Parameters     :
--|                      result       - output BIT_VECTOR, the computed product
--|                      overflow     - output BIT, overflow condition
--|                      multiplicand - input BIT_VECTOR,
--|                      multiplier   -  input BIT_VECTOR,
--|                      SrcRegMode   - input  regmode_type, indicating the format 
--|                                     of the input BIT_VECTOR.   Default is 
--|                                     DefaultRegMode which is set to TwosComp.
--|     NOTE           :
--|                      The inputs may be of any length and may be of differing
--|                      lengths.
--|
--|    Algorithm       : The multiplication is carried out as follows:
--|
--|                      1) Determine sign of result based on sign of 
--|                         multiploicand and sign  of multiplier.
--|
--|                      2) Convert the multiplicand amd multiplier to Unsigned 
--|                         representation.
--|                      
--|                      3) Perform multiplication based on add and shift algorithm.
--|
--|                      4) Convert the result to the SrcRegMode with appropropriate sign
--|
--|     Result         :
--|                     A  temporary result is computed with length N+M (where
--|                      N,M are the lengths of the multiplicand and multiplier)
--|                      by calling local function Mult_TwosComp or Mult_Unsigned
--|                       
--|                      This computed value is extended or truncated to match
--|                      the width of 'result'. If truncated, the low order bits
--|                      are returned.
--|
--|                      The parameter 'overflow' is set to '1' if the product of the
--|                      two inputs is too large to fit in the parameter result.
--|     Use            :
--|                      VARIABLE x, y, prod : BIT_VECTOR ( 15 DOWNTO 0);
--|                      VARIABLE ovfl : BIT;
--|
--|                      RegMult ( prod, ovfl, x, y, TwosComp );
--|
--|     See Also       : RegAdd, RegSub, RegMult, RegDiv, RegInc, RegDec, RegNegate
--|-----------------------------------------------------------------------------
    PROCEDURE RegMult ( VARIABLE result       : OUT BIT_VECTOR;
                        VARIABLE overflow     : OUT BIT;
                        CONSTANT multiplicand : IN BIT_VECTOR;
                        CONSTANT multiplier   : IN BIT_VECTOR;
                        CONSTANT SrcRegMode   : IN regmode_type
                 -- synopsys synthesis_off
                                                      := DefaultRegMode 
                 -- synopsys synthesis_on

                      ) IS
	VARIABLE reslt : STD_LOGIC_VECTOR (result'length - 1 downto 0);
	VARIABLE ovflo : STD_ULOGIC;
	VARIABLE  a    : STD_LOGIC_VECTOR ( multiplicand'Length - 1 DOWNTO 0 );
	VARIABLE  b    : STD_LOGIC_VECTOR (multiplier'Length - 1 DOWNTO 0 );
     BEGIN 
	a    := To_StdLogicVector(multiplicand);
        b    := To_StdLogicVector(multiplier);
	RegMult(reslt, ovflo, a, b, SrcRegMode);
        result   := To_BitVector(reslt);
        overflow := To_Bit(ovflo);
        RETURN;
    END RegMult;
--+-----------------------------------------------------------------------------
--|     Function Name  : RegDiv
--|
--|     Overloading    : None
--|
--|     Purpose        : Division of STD_LOGIC_VECTORS. (Result = dividend / divisor)
--|
--|     Parameters     :
--|                      result     - output STD_LOGIC_VECTOR,
--|                      remainder  - output STD_LOGIC_VECTOR,
--|                      ZeroDivide - output STD_ULOGIC,
--|                                   set to '1'  when divide by zero occurred
--|                                          '0'  divide by zero did not occur
--|                      dividend   - input  STD_LOGIC_VECTOR,
--|                      divisor    - input  STD_LOGIC_VECTOR,
--|                      SrcRegMode - input  regmode_type, indicating the format of
--|                                the input STD_LOGIC_VECTOR.   Default is TwosComp.
--|     NOTE           :
--|                      The inputs may be of any length and may be of differing
--|                      lengths.
--|
--|                      For synthesis purposes result and remainder values are 
--|                      computed with  same length as the dividend. 
--|
--|                      The remainder has the same sign as the dividend.
--|     Use            :
--|                      VARIABLE x, y, res, rem : STD_LOGIC_VECTOR ( 15 DOWNTO 0);
--|                      VARIABLE zflag     : STD_ULOGIC;
--|
--|                      RegDiv ( res, rem,zflag, x, y, TwosComp );
--|
--|     See Also       : RegAdd, RegSub, RegMult, RegDiv, RegInc, RegDec, RegNegate
--|-----------------------------------------------------------------------------
    PROCEDURE RegDiv  ( VARIABLE result     : OUT STD_LOGIC_VECTOR;
                        VARIABLE remainder  : OUT STD_LOGIC_VECTOR;
                        VARIABLE ZeroDivide : OUT STD_ULOGIC;
                        CONSTANT dividend   :  IN STD_LOGIC_VECTOR;
                        CONSTANT divisor    :  IN STD_LOGIC_VECTOR;
                        CONSTANT SrcRegMode    :  IN regmode_type
                     -- synopsys synthesis_off
						      := DefaultRegMode 
                     -- synopsys synthesis_on
                      ) IS
      CONSTANT len           : INTEGER := 2 * dividend'LENGTH;
      VARIABLE res_copy      : STD_LOGIC_VECTOR(result'LENGTH - 1 DOWNTO 0);
      VARIABLE rem_copy      : STD_LOGIC_VECTOR(remainder'LENGTH - 1 DOWNTO 0);
      VARIABLE dividend_copy : STD_LOGIC_VECTOR(dividend'LENGTH - 1 DOWNTO 0);
      VARIABLE divisor_copy  : STD_LOGIC_VECTOR(divisor'LENGTH - 1 DOWNTO 0);
      VARIABLE regr          : STD_LOGIC_VECTOR(len  DOWNTO 0);
      VARIABLE rega          : STD_LOGIC_VECTOR(len  DOWNTO 0);
      VARIABLE regd          : STD_LOGIC_VECTOR(len  DOWNTO 0);
      VARIABLE regb          : STD_LOGIC_VECTOR(dividend'LENGTH - 1  DOWNTO 0);   -- quotient
      VARIABLE sign_res      : std_ulogic;                        -- sign of result
      VARIABLE sign_rem      : std_ulogic;                        -- sign of remainder
      VARIABLE shiftout      : STD_ULOGIC;
     BEGIN 
    -- Initializations
       dividend_copy   := dividend;
       divisor_copy    := divisor;
       regr            := (OTHERS => '0');
       rega            := (OTHERS => '0');
       regd            := (OTHERS => '0');
      
     -- synopsys translate_off
     --   Null range check
     --   if result vector or remainder vector has a null range
       IF (( result'LENGTH = 0) OR (remainder'LENGTH = 0)) THEN
             ASSERT false
             REPORT " RegDiv  ---  Destination   has null range. "
             SEVERITY ERROR;
             RETURN;
     --   if both dividend  divisor  have null range no need to divide
       ELSIF (dividend'LENGTH = 0) AND (divisor'LENGTH = 0) THEN
             ASSERT false
             REPORT " RegDiv --- both dividend  and divisor has null range "
             SEVERITY ERROR;
             res_copy :=  (OTHERS => '0');
             result := res_copy;                   -- result is filled with zeros
             rem_copy :=  (OTHERS => '0');
             remainder := rem_copy;                -- remainder is filled with zeros
             RETURN;      

     -- if one of the dividend  or divisor is null 
       ELSIF (dividend'LENGTH = 0) THEN
             ASSERT false
             REPORT " RegDiv ---  dividend  has null range "
             SEVERITY ERROR;
                                 -- treat dividend as zero so result is zero 
             res_copy := (OTHERS => '0');
             result := res_copy;
             rem_copy :=  (OTHERS => '0');
             remainder := rem_copy;                -- remainder is filled with zeros
             RETURN;
       ELSIF (divisor'LENGTH = 0) THEN
             ASSERT false
             REPORT " RegDiv --- divisor  has null range "
             SEVERITY ERROR;
                                 -- treat result as zero 
             res_copy := (OTHERS => '0');
             result := res_copy;
             rem_copy :=  (OTHERS => '0');
             remainder := rem_copy;                -- remainder is filled with zeros
             RETURN;
       END IF;
    -- synopsys translate_on
    -- check for divide by zero
      IF (All_Zero(divisor_copy))  THEN
    -- synopsys translate_off              
           ASSERT false
           REPORT " RegDiv  ---  divide by zero  "
           SEVERITY ERROR;
    -- synopsys translate_on           
           res_copy := (OTHERS => '0');
           result := res_copy;
           rem_copy :=  (OTHERS => '0');
           remainder := rem_copy;                -- remainder is filled with zeros
	   ZeroDivide := '1';	
      ELSE

          -- inputs are  not null so determine the sign and convert 
          -- the inputs to unsigned  representation.
            sign_res := dividend(dividend'LEFT) XOR divisor(divisor'LEFT);
            sign_rem := dividend(dividend'LEFT);
            dividend_copy := To_Unsign(dividend_copy, SrcRegMode);
            divisor_copy := To_Unsign(divisor_copy, SrcRegMode);  
      
           -- put dividend to rega  and divisor to regd
             for i IN dividend'Length - 1 downto 0 Loop
		  rega(i) := dividend_copy(i);
             end Loop;
             for i IN divisor'Length - 1 downto 0 Loop
		  regd(i) := divisor_copy(i);
             end Loop;

            -- Perform division by binary restoring algorithm
            --    initialize 
            -- load rega to regr, 
            -- regd  gets regd shifted left by nd bits
            -- regb  gets all zerso
             regr := rega;                
            -- left shift regd by dividend'LENGTH ( length of divisor) bits, fill with zero's
             RegShift_Left(regd, regd, shiftout, '0', dividend'LENGTH);
             regb := (OTHERS =>'0');

             For i IN 0 TO dividend'LENGTH - 1 LOOP
                                                -- regr := 2*regr - regd
                 RegShift_Left(regr, regr, shiftout,  '0', 1);
                 RegSub_Syn (regr,  regr,  regd, TwosComp);                 
                 IF (regr(regr'LEFT) /= '0')   THEN
                                               -- regr := regr + regd
                     RegAdd_Syn(regr, regr, regd, TwosComp);
                     RegShift_Left(regb, regb, shiftout, '0', 1);
                 ELSE
                                                   -- regb := 2*regb + 1;
                      RegShift_Left(regb, regb, shiftout, '0', 1);
                      regb := RegInc(regb, Unsigned);
                 END IF;
             END LOOP;
             -- if the result and remainder should be negative
	     -- modyfying for synthesis	
             IF (( sign_res /= '0' ) AND (SrcRegMode /= Unsigned)) THEN
                  regb := RegNegate(regb, SrcRegMode);
                  res_copy := regb;
             ELSE 
                  res_copy := regb;
             END IF;

            IF ((sign_rem /= '0') AND (SrcRegMode /= Unsigned)) THEN
                 regr := RegNegate(regr, SrcRegMode);
            END IF;
                -- remainder is in most significant N bits, shift right N bits 
            RegShift_Right(regr, regr, shiftout,  regr(len), dividend'LENGTH);
           -- remainder length
            rem_copy := regr(dividend'LENGTH - 1 downto 0);
            result := To_X01(res_copy);
            remainder := To_X01( rem_copy);
            ZeroDivide := '0';	
        END IF;
       -- That's all
        RETURN;
   END RegDiv;         
--+-----------------------------------------------------------------------------
--|     Function Name  : RegDiv
--|
--|     Overloading    : None
--|
--|     Purpose        : Division of STD_ULOGIC_VECTORS. (Result = dividend / divisor)
--|
--|     Parameters     :
--|                      result     - output STD_ULOGIC_VECTOR,
--|                      remainder  - output STD_ULOGIC_VECTOR,
--|                      ZeroDivide - output STD_ULOGIC,
--|                                   set to '1'  when divide by zero occurred
--|                                          '0'  divide by zero did not occur
--|                      dividend   - input  STD_ULOGIC_VECTOR,
--|                      divisor    - input  STD_ULOGIC_VECTOR,
--|                      SrcRegMode - input  regmode_type, indicating the format of
--|                                the input STD_ULOGIC_VECTOR.   Default is TwosComp.
--|     NOTE           :
--|                      The inputs may be of any length and may be of differing
--|                      lengths.
--|
--|                      For synthesis purposes result and remainder values are 
--|                      computed with  same length as the dividend. 
--|
--|                      The remainder has the same sign as the dividend.
--|     Use            :
--|                      VARIABLE x, y, res, rem : STD_ULOGIC_VECTOR ( 15 DOWNTO 0);
--|                      VARIABLE zflag     : STD_ULOGIC;
--|
--|                      RegDiv ( res, rem,zflag, x, y, TwosComp );
--|
--|     See Also       : RegAdd, RegSub, RegMult, RegDiv, RegInc, RegDec, RegNegate
--|-----------------------------------------------------------------------------
    PROCEDURE RegDiv  ( VARIABLE result     : OUT STD_ULOGIC_VECTOR;
                        VARIABLE remainder  : OUT STD_ULOGIC_VECTOR;
                        VARIABLE ZeroDivide : OUT STD_ULOGIC;
                        CONSTANT dividend   :  IN STD_ULOGIC_VECTOR;
                        CONSTANT divisor    :  IN STD_ULOGIC_VECTOR;
                        CONSTANT SrcRegMode    :  IN regmode_type
                     -- synopsys synthesis_off
						      := DefaultRegMode 
                     -- synopsys synthesis_on
                      ) IS
        VARIABLE reslt    : STD_LOGIC_VECTOR(result'LENGTH - 1 DOWNTO 0);
        VARIABLE remaind  : STD_LOGIC_VECTOR(remainder'LENGTH - 1 DOWNTO 0);
        VARIABLE  a_copy  : STD_LOGIC_VECTOR (dividend'Length - 1 DOWNTO 0 );
	VARIABLE  b_copy  : STD_LOGIC_VECTOR (divisor'Length - 1 DOWNTO 0 );
     BEGIN 
	a_copy    := To_StdLogicVector(dividend);
        b_copy    := To_StdLogicVector(divisor);
        RegDiv(reslt, remaind, ZeroDivide, a_copy, b_copy, SrcRegMode);
	result := To_StdULogicVector(reslt);
        remainder := To_StdUlogicVector(remaind);        
        RETURN;
   END RegDiv;         
--+-----------------------------------------------------------------------------
--|     Function Name  : RegDiv
--|
--|     Overloading    : None
--|
--|     Purpose        : Division of BIT_VECTORS. (Result = dividend / divisor)
--|
--|     Parameters     :
--|                      result     - output BIT_VECTOR,
--|                      remainder  - output BIT_VECTOR,
--|                      ZeroDivide - output BIT,
--|                                   set to '1'  when divide by zero occurred
--|                                          '0'  divide by zero did not occur
--|                      dividend   - input  BIT_VECTOR,
--|                      divisor    - input  BIT_VECTOR,
--|                      SrcRegMode - input  regmode_type, indicating the format of
--|                                the input BIT_VECTOR.   Default is TwosComp.
--|     NOTE           :
--|                      The inputs may be of any length and may be of differing
--|                      lengths.
--|
--|                      For synthesis purposes result and remainder values are 
--|                      computed with  same length as the dividend. 
--|
--|                      The remainder has the same sign as the dividend.
--|     Use            :
--|                      VARIABLE x, y, res, rem : BIT_VECTOR ( 15 DOWNTO 0);
--|                      VARIABLE zflag     : BIT;
--|
--|                      RegDiv ( res, rem,zflag, x, y, TwosComp );
--|
--|     See Also       : RegAdd, RegSub, RegMult, RegDiv, RegInc, RegDec, RegNegate
--|-----------------------------------------------------------------------------
    PROCEDURE RegDiv  ( VARIABLE result     : OUT BIT_VECTOR;
                        VARIABLE remainder  : OUT BIT_VECTOR;
                        VARIABLE ZeroDivide : OUT BIT;
                        CONSTANT dividend   :  IN BIT_VECTOR;
                        CONSTANT divisor    :  IN BIT_VECTOR;
                        CONSTANT SrcRegMode    :  IN regmode_type
                     -- synopsys synthesis_off
						      := DefaultRegMode 
                     -- synopsys synthesis_on
                      ) IS

        VARIABLE reslt    : STD_LOGIC_VECTOR(result'LENGTH - 1 DOWNTO 0);
        VARIABLE remaind  : STD_LOGIC_VECTOR(remainder'LENGTH - 1 DOWNTO 0);
        VARIABLE Zdiv     : STD_ULOGIC;
        VARIABLE  a_copy  : STD_LOGIC_VECTOR (dividend'Length - 1 DOWNTO 0 );
	VARIABLE  b_copy  : STD_LOGIC_VECTOR (divisor'Length - 1 DOWNTO 0 );
     BEGIN 
	a_copy    := To_StdLogicVector(dividend);
        b_copy    := To_StdLogicVector(divisor);
        RegDiv(reslt, remaind, Zdiv, a_copy, b_copy, SrcRegMode);
	result := To_BitVector(reslt);
        remainder := To_BitVector(remaind);        
        ZeroDivide := To_Bit(Zdiv);
        RETURN;
   END RegDiv;
--+-----------------------------------------------------------------------------
--|     Function Name  : RegRem
--| 1.5.25
--|     Overloading    : None
--|
--|     Purpose        : Remainder operation of  STD_LOGIC_VECTORS.
--|
--|     Parameters     :
--|                      result     - output STD_LOGIC_VECTOR,
--|                      ZeroDivide - output STD_ULOGIC,
--|                                   set to '1'  when divide by zero occurred
--|                                          '0'  divide by zero did not occur
--|                      dividend   - input  STD_LOGIC_VECTOR,
--|                      divisor    - input  STD_LOGIC_VECTOR,
--|                      SrcRegMode - input  regmode_type, indicating the format of
--|                                the input STD_LOGIC_VECTOR.   Default is TwosComp.
--|     NOTE           :
--|                      The inputs may be of any length and may be of differing
--|                      lengths.
--|
--|                      For synthesis purposes quotient and remainder values are 
--|                      computed with  same length as the dividend. 
--|
--|                      The remainder has the same sign as the dividend.
--|     Use            :
--|                      VARIABLE x, y, res : STD_LOGIC_VECTOR ( 15 DOWNTO 0);
--|                      VARIABLE zflag     : STD_ULOGIC;
--|
--|                      RegRem ( res, zflag, x, y, TwosComp );
--|
--|     See Also       : RegAdd, RegSub, RegMult, RegDiv, RegInc, RegDec, RegNegate
--|-----------------------------------------------------------------------------
    PROCEDURE RegRem  ( VARIABLE result     : OUT STD_LOGIC_VECTOR;
                        VARIABLE ZeroDivide : OUT STD_ULOGIC;
                        CONSTANT dividend   :  IN STD_LOGIC_VECTOR;
                        CONSTANT divisor    :  IN STD_LOGIC_VECTOR;
                        CONSTANT SrcRegMode :  IN regmode_type
                     -- synopsys synthesis_off
						      := DefaultRegMode 
                     -- synopsys synthesis_on
                      ) IS
      CONSTANT len       : INTEGER := 2 * dividend'LENGTH;
      VARIABLE res_copy : STD_LOGIC_VECTOR(result'LENGTH - 1 DOWNTO 0);
      VARIABLE dividend_copy : STD_LOGIC_VECTOR(dividend'LENGTH - 1 DOWNTO 0);
      VARIABLE divisor_copy  : STD_LOGIC_VECTOR(divisor'LENGTH - 1 DOWNTO 0);
      VARIABLE regr      : STD_LOGIC_VECTOR(len  DOWNTO 0);
      VARIABLE rega      : STD_LOGIC_VECTOR(len  DOWNTO 0);
      VARIABLE regd      : STD_LOGIC_VECTOR(len  DOWNTO 0);
      VARIABLE regb      : STD_LOGIC_VECTOR(dividend'LENGTH - 1 DOWNTO 0);   -- quotient
      VARIABLE sign_res  : STD_ULOGIC;              -- sign of result
      VARIABLE shiftout  : STD_ULOGIC;
     BEGIN 
    -- Initializations
       dividend_copy   := dividend;
       divisor_copy    := divisor;
       regr            := (OTHERS => '0');
       rega            := (OTHERS => '0');
       regd            := (OTHERS => '0');
     -- synopsys translate_off
     --   Null range check
     --   if result vector null range
       IF ( result'LENGTH = 0)  THEN
             ASSERT false
             REPORT " RegRem  ---  Destination   has null range. "
             SEVERITY ERROR;
             RETURN;
     --   if both dividend   and divisor   have null range no need to divide
       ELSIF (dividend'LENGTH = 0) AND (divisor'LENGTH = 0) THEN
             ASSERT false
             REPORT " RegRem --- both dividend  and divisor has null range "
             SEVERITY ERROR;
             res_copy :=  (OTHERS => '0');
             result := res_copy;                   -- result is filled with zeros
             RETURN;      
     -- if one of the dividend  or divisor is null 
       ELSIF (dividend'LENGTH = 0) THEN
             ASSERT false
             REPORT " RegRem ---  dividend  has null range "
             SEVERITY ERROR;
                                 -- treat dividend as zero so result is zero 
             res_copy := (OTHERS => '0');
             result := res_copy;
             RETURN;
       ELSIF (divisor'LENGTH = 0) THEN
             ASSERT false
             REPORT " RegRem --- divisor  has null range "
             SEVERITY ERROR;
                                 -- treat result as zero 
             res_copy := (OTHERS => '0');
             result := res_copy;
             RETURN;
       END IF;
     -- synopsys translate_on           
    -- check for divide by zero
      IF (All_Zero(divisor_copy))  THEN
     -- synopsys translate_off
          ASSERT false
          REPORT " RegRem  ---  divide by zero  "
          SEVERITY ERROR;
     -- synopsys translate_on
          res_copy := (OTHERS => '0');
          result := res_copy;
          ZeroDivide := '1';	
      ELSE
        -- inputs are  not null so determine the sign and convert 
        -- the inputs to unsigned  representation.
          sign_res := dividend(dividend'LEFT); -- sign of dividend is sign of result
          dividend_copy := To_Unsign (dividend_copy, SrcRegMode);     
          divisor_copy := To_Unsign(divisor_copy, SrcRegMode);  
          -- put dividend to rega  and divisor to regd
            for i IN dividend'Length - 1 downto 0 Loop
		rega(i) := dividend_copy(i);
            end Loop;
            for i IN divisor'Length - 1 downto 0 Loop
	        regd(i) := divisor_copy(i);
            end Loop;
           -- Perform division by binary restoring algorithm
           --    initialize 
           -- load rega to regr, 
           -- regd  gets regd shifted left by dividend'length bits
           -- regb  gets all zerso
            regr := rega;                
              -- left shift regd by dividend'LENGTH  bits, fill with zero's
            RegShift_Left(regd, regd, shiftout, '0', dividend'LENGTH);
            regb := (OTHERS =>'0');
            For i IN 0 TO dividend'LENGTH - 1 LOOP
                                                -- regr := 2*regr - regd
                RegShift_Left(regr, regr, shiftout,  '0', 1);
                RegSub_Syn (regr,  regr,  regd, TwosComp);                 
                IF (regr(regr'LEFT) /= '0')   THEN
                                               -- regr := regr + regd
                    RegAdd_Syn(regr, regr, regd,  TwosComp);
                    RegShift_Left(regb, regb, shiftout, '0', 1);
                ELSE
                                                 -- regb := 2*regb + 1;
                    RegShift_Left(regb, regb, shiftout, '0', 1);
                    regb := RegInc(regb, Unsigned);
                END IF;
             END LOOP;
           -- if the result  should be negative 
             IF (( sign_res /= '0') AND (SrcRegMode /= Unsigned)) THEN
                 regr := RegNegate(regr, SrcRegMode);
                 -- most significant of regr holds result
                 RegShift_Right(regr, regr, shiftout, regr(len), dividend'LENGTH);
             ELSE           
                 -- most significant of regr holds result
                 RegShift_Right(regr, regr, shiftout, regr(len), dividend'LENGTH);
             END IF;
             res_copy := regr(dividend'LENGTH - 1 downto 0);                
             result := To_X01(res_copy);
             ZeroDivide := '0';	
         END IF;
         RETURN;
    END RegRem;
--+-----------------------------------------------------------------------------
--|     Function Name  : RegRem
--| 1.5.25
--|     Overloading    : None
--|
--|     Purpose        : Remainder operation of  STD_ULOGIC_VECTORS.
--|
--|     Parameters     :
--|                      result     - output STD_ULOGIC_VECTOR,
--|                      ZeroDivide - output STD_ULOGIC,
--|                                   set to '1'  when divide by zero occurred
--|                                          '0'  divide by zero did not occur
--|                      dividend   - input  STD_ULOGIC_VECTOR,
--|                      divisor    - input  STD_ULOGIC_VECTOR,
--|                      SrcRegMode - input  regmode_type, indicating the format of
--|                                the input STD_ULOGIC_VECTOR.   Default is TwosComp.
--|     NOTE           :
--|                      The inputs may be of any length and may be of differing
--|                      lengths.
--|
--|                      For synthesis purposes result is 
--|                      computed with  same length as the dividend. 
--|
--|                      The remainder has the same sign as the dividend.
--|     Use            :
--|                      VARIABLE x, y, res : STD_ULOGIC_VECTOR ( 15 DOWNTO 0);
--|                      VARIABLE zflag     : STD_ULOGIC;
--|
--|                      RegRem ( res, zflag, x, y, TwosComp );
--|
--|     See Also       : RegAdd, RegSub, RegMult, RegDiv, RegInc, RegDec, RegNegate
--|-----------------------------------------------------------------------------
    PROCEDURE RegRem  ( VARIABLE result     : OUT STD_ULOGIC_VECTOR;
                        VARIABLE ZeroDivide : OUT STD_ULOGIC;
                        CONSTANT dividend   :  IN STD_ULOGIC_VECTOR;
                        CONSTANT divisor    :  IN STD_ULOGIC_VECTOR;
                        CONSTANT SrcRegMode :  IN regmode_type
                     -- synopsys synthesis_off
						      := DefaultRegMode 
                     -- synopsys synthesis_on
                      ) IS
        VARIABLE reslt : STD_LOGIC_VECTOR(result'LENGTH - 1 DOWNTO 0);
        VARIABLE  a_copy  : STD_LOGIC_VECTOR (dividend'Length - 1 DOWNTO 0 );
	VARIABLE  b_copy  : STD_LOGIC_VECTOR (divisor'Length - 1 DOWNTO 0 );
     BEGIN 
	a_copy    := To_StdLogicVector(dividend);
        b_copy    := To_StdLogicVector(divisor);
	RegRem(reslt, ZeroDivide, a_copy, b_copy, SrcRegMode);
        result := To_StdULogicVector(reslt);
        RETURN;
    END RegRem;
--+-----------------------------------------------------------------------------
--|     Function Name  : RegRem
--| 1.5.25
--|     Overloading    : None
--|
--|     Purpose        : Remainder operation of  BIT_VECTORS.
--|
--|     Parameters     :
--|                      result     - output BIT_VECTOR,
--|                      ZeroDivide - output BIT,
--|                                   set to '1'  when divide by zero occurred
--|                                          '0'  divide by zero did not occur
--|                      dividend   - input  BIT_VECTOR,
--|                      divisor    - input  BIT_VECTOR,
--|                      SrcRegMode - input  regmode_type, indicating the format of
--|                                the input BIT_VECTOR.   Default is TwosComp.
--|     NOTE           :
--|                      The inputs may be of any length and may be of differing
--|                      lengths.
--|
--|                      For synthesis purposes result is 
--|                      computed with  same length as the dividend. 
--|
--|                      The remainder has the same sign as the dividend.
--|     Use            :
--|                      VARIABLE x, y, res : BIT_VECTOR ( 15 DOWNTO 0);
--|                      VARIABLE zflag     : BIT;
--|
--|                      RegRem ( res, zflag, x, y, TwosComp );
--|
--|     See Also       : RegAdd, RegSub, RegMult, RegDiv, RegInc, RegDec, RegNegate
--|-----------------------------------------------------------------------------
    PROCEDURE RegRem  ( VARIABLE result     : OUT BIT_VECTOR;
                        VARIABLE ZeroDivide : OUT BIT;
                        CONSTANT dividend   :  IN BIT_VECTOR;
                        CONSTANT divisor    :  IN BIT_VECTOR;
                        CONSTANT SrcRegMode :  IN regmode_type 
                     -- synopsys synthesis_off
						      := DefaultRegMode 
                     -- synopsys synthesis_on
                      ) IS
        VARIABLE reslt    : STD_LOGIC_VECTOR(result'LENGTH - 1 DOWNTO 0);
        VARIABLE Zdiv     : STD_ULOGIC;
        VARIABLE  a_copy  : STD_LOGIC_VECTOR (dividend'Length - 1 DOWNTO 0 );
	VARIABLE  b_copy  : STD_LOGIC_VECTOR (divisor'Length - 1 DOWNTO 0 );
     BEGIN 
	a_copy    := To_StdLogicVector(dividend);
        b_copy    := To_StdLogicVector(divisor);
        RegRem(reslt, Zdiv, a_copy, b_copy, SrcRegMode);
	result := To_BitVector(reslt);
        ZeroDivide := To_Bit(Zdiv);
        return;
    END RegRem;
--+-----------------------------------------------------------------------------
--|     Function Name  : RegMod
--| 1.5.17  
--|     Overloading    : None
--| 
--|     Purpose        : Modulus operation of  STD_LOGIC_VECTORS.
--| 
--|     Parameters     :
--|                      result     - output STD_LOGIC_VECTOR,
--|                      ZeroDivide - output STD_ULOGIC,
--|                                   set to '1'  when divide by zero occurred
--|                                          '0'  divide by zero did not occur
--|                      dividend   - input  STD_LOGIC_VECTOR,
--|                      modulus    - input  STD_LOGIC_VECTOR,
--|                      SrcRegMode - input  regmode_type, indicating the format of
--|                                the input STD_LOGIC_VECTOR.   Default is TwosComp.
--|     NOTE           :
--|                      The inputs may be of any length and may be of differing
--|                      lengths.
--|
--|                      For synthesis purposes quotient and modulus values are 
--|                      computed with  same length as the dividend. 
--|
--|                      The mod has the same sign as the modulus operator.
--|     Use            :
--|                      VARIABLE x, y, res : STD_LOGIC_VECTOR ( 15 DOWNTO 0);
--|                      VARIABLE zflag     : STD_ULOGIC;
--|
--|                      RegMod ( res,zflag, x, y, TwosComp );
--|
--|     See Also       : RegAdd, RegSub, RegMult, RegDiv, RegInc, RegDec, RegNegate
--|-----------------------------------------------------------------------------
    PROCEDURE RegMod  ( VARIABLE result     : OUT STD_LOGIC_VECTOR;
                        VARIABLE ZeroDivide : OUT STD_ULOGIC;
                        CONSTANT dividend   : IN STD_LOGIC_VECTOR;
                        CONSTANT modulus    : IN STD_LOGIC_VECTOR;
                        CONSTANT SrcRegMode : IN regmode_type
                     -- synopsys synthesis_off
						      := DefaultRegMode 
                     -- synopsys synthesis_on
                      ) IS

      VARIABLE res_copy      : STD_LOGIC_VECTOR(result'LENGTH - 1 DOWNTO 0);
      VARIABLE res           : STD_LOGIC_VECTOR(result'LENGTH - 1 DOWNTO 0);
      VARIABLE remainderb     : STD_LOGIC_VECTOR(result'LENGTH - 1 DOWNTO 0);
      VARIABLE divid_copy : STD_LOGIC_VECTOR(dividend'LENGTH - 1 DOWNTO 0);
      VARIABLE modulus_copy  : STD_LOGIC_VECTOR(modulus'LENGTH - 1 DOWNTO 0);
      VARIABLE zeroflag      : STD_ULOGIC;
      VARIABLE c_out         : STD_ULOGIC;
      VARIABLE uvflo         : STD_ULOGIC;
     BEGIN 
	-- Initializations
        divid_copy    := dividend;
        modulus_copy  := modulus;
     -- synopsys translate_off	
     --   Null range check
     --   if result vector or remainderb vector has a null range
       IF ( result'LENGTH = 0) THEN
             ASSERT false
             REPORT " RegMod  ---  Destination   has null range. "
             SEVERITY ERROR;
             RETURN;
     --   if both dividend   and modulus   have null range no need to divide
       ELSIF (dividend'LENGTH = 0) AND (modulus'LENGTH = 0) THEN
             ASSERT false
             REPORT " RegMod --- both dividend  and modulus has null range "
             SEVERITY ERROR;
             res_copy :=  (OTHERS => '0');
             result := res_copy;            -- result is filled with zeros
             RETURN;      

     -- if one of the dividend  or divisor is null 
       ELSIF (dividend'LENGTH = 0) THEN
             ASSERT false
             REPORT " RegMod ---  dividend  has null range "
             SEVERITY ERROR;
                              -- treat dividend as zero so result is zero 
             res_copy := (OTHERS => '0');
             result := res_copy;
             RETURN;
       ELSIF (modulus'LENGTH = 0) THEN
             ASSERT false
             REPORT " RegMod --- modulus  has null range "
             SEVERITY ERROR;
                                 -- treat result as zero 
             res_copy := (OTHERS => '0');
             result := res_copy;
             RETURN;
       END IF;
      -- synopsys translate_on           
    -- check for divide by zero
      IF (All_Zero(modulus_copy))  THEN 
      -- synopsys translate_off
           ASSERT false
           REPORT " RegMod  ---  divide by zero  "
           SEVERITY ERROR;
      -- synopsys translate_on
           res_copy := (OTHERS => '0');
           result := res_copy;
           ZeroDivide := '1';	
       ELSE
        -- Use procedure RegDiv to calculate the remainderb
        -- Then mod is calculated
          RegDiv(res, remainderb, zeroflag, divid_copy, modulus_copy, SrcRegMode);
          res_copy := remainderb;
          IF ( (SrcRegMode /= Unsigned) AND ( dividend(dividend'LEFT) = '0')) THEN 
                                                                  -- dividend positive
              IF (ALL_Zero(remainderb)) THEN
                  null;
              ELSIF (modulus(modulus'LEFT) /= '0') THEN   -- negative modulus
                   RegAdd(res_copy, c_out, uvflo, modulus_copy, remainderb, '0', SrcRegMode); 
              END IF;
           ELSIF ((SrcRegMode /= Unsigned) AND (dividend(dividend'LEFT) /= '0')) THEN
                                      -- negative dividend
              IF (All_Zero(remainderb)) THEN
                  null;
               ELSIF (modulus_copy(modulus_copy'LEFT ) = '0') THEN      -- positive modulus
                   RegAdd(res_copy, c_out, uvflo, modulus_copy, remainderb, '0', SrcRegMode);
               END IF;
           END IF;
           result := res_copy;    -- copy internal res_copy to result
           ZeroDivide := '0';	
       END IF;
       RETURN;
    END RegMod;
--+-----------------------------------------------------------------------------
--|     Function Name  : RegMod
--| 1.5.17  
--|     Overloading    : None
--| 
--|     Purpose        : Modulus operation of  STD_ULOGIC_VECTORS.
--| 
--|     Parameters     :
--|                      result     - output STD_ULOGIC_VECTOR,
--|                      ZeroDivide - output STD_ULOGIC,
--|                                   set to '1'  when divide by zero occurred
--|                                          '0'  divide by zero did not occur
--|                      dividend   - input  STD_ULOGIC_VECTOR,
--|                      modulus    - input  STD_ULOGIC_VECTOR,
--|                      SrcRegMode - input  regmode_type, indicating the format of
--|                                the input STD_ULOGIC_VECTOR.   Default is TwosComp.
--|     NOTE           :
--|                      The inputs may be of any length and may be of differing
--|                      lengths.
--|
--|                      For synthesis purposes quotient and modulus values are 
--|                      computed with  same length as the dividend. 
--|
--|                      The mod has the same sign as the modulus operator.
--|     Use            :
--|                      VARIABLE x, y, res : STD_ULOGIC_VECTOR ( 15 DOWNTO 0);
--|                      VARIABLE zflag     : STD_ULOGIC;
--|
--|                      RegMod ( res,zflag, x, y, TwosComp );
--|
--|     See Also       : RegAdd, RegSub, RegMult, RegDiv, RegInc, RegDec, RegNegate
--|-----------------------------------------------------------------------------
    PROCEDURE RegMod  ( VARIABLE result     : OUT STD_ULOGIC_VECTOR;
                        VARIABLE ZeroDivide : OUT STD_ULOGIC;
                        CONSTANT dividend   : IN STD_ULOGIC_VECTOR;
                        CONSTANT modulus    : IN STD_ULOGIC_VECTOR;
                        CONSTANT SrcRegMode : IN regmode_type
                     -- synopsys synthesis_off
						      := DefaultRegMode 
                     -- synopsys synthesis_on
                      ) IS
        VARIABLE reslt    : STD_LOGIC_VECTOR(result'LENGTH - 1 DOWNTO 0);
        VARIABLE  d_copy  : STD_LOGIC_VECTOR (dividend'Length - 1 DOWNTO 0 );
	VARIABLE  m_copy  : STD_LOGIC_VECTOR (modulus'Length - 1 DOWNTO 0 );
     BEGIN 
	d_copy    := To_StdLogicVector(dividend);
        m_copy    := To_StdLogicVector(modulus);
 	RegMod(reslt, ZeroDivide, d_copy, m_copy, SrcRegMode);
        result := To_StdULogicVector(reslt);
        RETURN;
    END RegMod;
--+-----------------------------------------------------------------------------
--|     Function Name  : RegMod
--| 1.5.17  
--|     Overloading    : None
--| 
--|     Purpose        : Modulus operation of  BIT_VECTORS.
--| 
--|     Parameters     :
--|                      result     - output BIT_VECTOR,
--|                      ZeroDivide - output BIT,
--|                                   set to '1'  when divide by zero occurred
--|                                          '0'  divide by zero did not occur
--|                      dividend   - input  BIT_VECTOR,
--|                      modulus    - input  BIT_VECTOR,
--|                      SrcRegMode - input  regmode_type, indicating the format of
--|                                the input BIT_VECTOR.   Default is TwosComp.
--|     NOTE           :
--|                      The inputs may be of any length and may be of differing
--|                      lengths.
--|
--|                      For synthesis purposes quotient and modulus values are 
--|                      computed with  same length as the dividend. 
--|
--|                      The mod has the same sign as the modulus operator.
--|     Use            :
--|                      VARIABLE x, y, res : BIT_VECTOR ( 15 DOWNTO 0);
--|                      VARIABLE zflag     : BIT;
--|
--|                      RegMod ( res,zflag, x, y, TwosComp );
--|
--|     See Also       : RegAdd, RegSub, RegMult, RegDiv, RegInc, RegDec, RegNegate
--|-----------------------------------------------------------------------------
    PROCEDURE RegMod  ( VARIABLE result     : OUT BIT_VECTOR;
                        VARIABLE ZeroDivide : OUT BIT;
                        CONSTANT dividend   : IN BIT_VECTOR;
                        CONSTANT modulus    : IN BIT_VECTOR;
                        CONSTANT SrcRegMode : IN regmode_type
                     -- synopsys synthesis_off
						      := DefaultRegMode 
                     -- synopsys synthesis_on
                      ) IS

        VARIABLE reslt    : STD_LOGIC_VECTOR(result'LENGTH - 1 DOWNTO 0);
        VARIABLE Zdiv     : STD_ULOGIC;
        VARIABLE  d_copy  : STD_LOGIC_VECTOR (dividend'Length - 1 DOWNTO 0 );
	VARIABLE  m_copy  : STD_LOGIC_VECTOR (modulus'Length - 1 DOWNTO 0 );
     BEGIN 
	d_copy    := To_StdLogicVector(dividend);
        m_copy    := To_StdLogicVector(modulus);
        RegMod(reslt, Zdiv, d_copy, m_copy, SrcRegMode);
	result := To_BitVector(reslt);
        ZeroDivide := To_Bit(Zdiv);
        RETURN;
    END RegMod;
--+-----------------------------------------------------------------------------
--|     Function Name  : RegShift
--| 
--|     Overloading    : None
--|
--|     Purpose        : Bidirectional logical shift operator for   BIT_VECTORS.
--|
--|     Parameters     :
--|                      SrcReg      - input  BIT_VECTOR, vector to be shifted
--|                      DstReg      - Input_ouput, BIT_VECTOR, shifted result
--|                      ShiftO      - output, BIT, holds the last bit shifted out 
--|                                          of register
--|                      direction   - input, BIT
--|                                     '0'  means right shift
--|                                     '1'  means left shift, default is left shift
--|                      FillVal     - input, BIT, value to fill register with. 
--|                                          default is '0'
--|                      Nbits       - input , NATURAL, number of positions to shift
--|                                          default is 1.
--|     NOTE           : 
--|                      Defaults not allowed for synthesis.
--|
--|     Result         : Shifted bit_vector
--|
--|     Use            : VARIABLE acc   : BIT_VECTOR ( 15 DOWNTO 0);
--|                      VARIABLE carry : BIT;
--|
--|                      RegShift ( acc, acc, carry, '1', '0',3 );
--|-----------------------------------------------------------------------------
   PROCEDURE RegShift  ( CONSTANT SrcReg    : IN BIT_VECTOR;
                         VARIABLE DstReg    : INOUT BIT_VECTOR;
                         VARIABLE ShiftO    : OUT BIT; 
                         CONSTANT direction : IN BIT     
                     -- synopsys synthesis_off
						      := '1'
                     -- synopsys synthesis_on
                                                            ;
                         CONSTANT FillVal   : IN BIT  
                     -- synopsys synthesis_off
						      := '0'
                     -- synopsys synthesis_on
                                                            ;
                         CONSTANT Nbits     : IN Natural
                     -- synopsys synthesis_off
						       := 1 
                     -- synopsys synthesis_on
                      ) IS 
      VARIABLE r         : BIT_VECTOR (SrcReg'LENGTH - 1 DOWNTO 0);
      VARIABLE src_copy  : BIT_VECTOR (SrcReg'LENGTH - 1 DOWNTO 0 );
      VARIABLE dst_copy  : BIT_VECTOR (DstReg'LENGTH - 1 DOWNTO 0 );
   BEGIN
       src_copy   := SrcReg;
       dst_copy   := DstReg;
 -- synopsys translate_off    
    --  Null range Check
    --  if input vector is of zero length
       IF ( SrcReg'LENGTH = 0) THEN
           ASSERT false
           REPORT " RegShift --- input bit_vector   is null  "
           SEVERITY ERROR;
           dst_copy := (OTHERS => FillVal);
           DstReg    := dst_copy;
           ShiftO := '0';
           Return;
       ELSIF (DstReg'LENGTH = 0) THEN
           ASSERT false
           REPORT " RegShift --- output vector is  null  "
           SEVERITY ERROR;
         -- set shift out bit at least
           IF ( direction /= '0') THEN
               ShiftO := src_copy(SrcReg'LENGTH - Nbits);
           ELSE 
               ShiftO := src_copy(Nbits - 1);
           END IF;
           RETURN;
      END IF;
-- synopsys translate_on
    -- None of the registers is null, perform shift operation
      IF (direction /= '0') THEN                                 --  left shift
           RegShift_Left(src_copy, r, ShiftO, FillVal, Nbits);
      ELSE                                                       -- right shift
           RegShift_Right(src_copy, r, ShiftO, FillVal, Nbits);
      END IF;
      -- determine length of the result
      IF (DstReg'LENGTH <= SrcReg'LENGTH) THEN
		for i IN DstReg'Length - 1 downto 0 Loop
			dst_copy(i) := r(i);
                end loop;
      ELSE
		for i IN SrcReg'LENGTH - 1 downto 0 Loop
			dst_copy(i) := r(i);
                end loop;
      END IF;
      DstReg := dst_copy;
      RETURN;
   END RegShift;
--+-----------------------------------------------------------------------------
--|     Function Name  : RegShift
--| 
--|     Overloading    : None
--|
--|     Purpose        : Bidirectional logical shift operator for logic vector.
--|
--|     Parameters     :
--|                      SrcReg      - input  std_logic_vector, vector to be shifted
--|                      DstReg      - ouput, std_logic_vector, shifted result
--|                      ShiftO      - output, std_ulogic, holds the 
--|                                            last bit shifted out 
--|                                          of register
--|                      direction   - input, Std_ulogic
--|                                         '0'  means right shift
--|                                         '1' | 'X'  means left shift, 
--|                                          default is left shift
--|                      FillVal     - input, Std_ulogic, value to fill register with. 
--|                                          default is '0'
--|                      Nbits       - input , NATURAL, number of positions to shift
--|                                          default is 1.
--|
--|     Result         : Shifted std_logic_vector
--|
--|     NOTE           : Defaults not allowed for synthesis.
--|
--|     Use            : VARIABLE acc   : std_logic_vector ( 15 DOWNTO 0);
--|                      VARIABLE carry : std_ulogic;
--|
--|                      RegShift ( acc, acc, carry, '1', '0',3 );
--|-----------------------------------------------------------------------------
   PROCEDURE RegShift  ( CONSTANT SrcReg    : IN std_logic_vector;
                         VARIABLE DstReg    : INOUT std_logic_vector;
                         VARIABLE ShiftO    : OUT std_ulogic; 
                         CONSTANT direction : IN std_ulogic
                     -- synopsys synthesis_off
						      := '1'
                     -- synopsys synthesis_on
                                                            ;
                         CONSTANT FillVal   : IN std_ulogic  
                     -- synopsys synthesis_off
						      := '0'
                     -- synopsys synthesis_on
                                                            ;
                         CONSTANT Nbits     : IN Natural
                     -- synopsys synthesis_off
						       := 1 
                     -- synopsys synthesis_on
                      ) IS 
      VARIABLE r         : STD_LOGIC_VECTOR (SrcReg'LENGTH - 1 DOWNTO 0);
      VARIABLE src_copy  : STD_LOGIC_VECTOR (SrcReg'LENGTH - 1 DOWNTO 0 );
      VARIABLE dst_copy  : STD_LOGIC_VECTOR (DstReg'LENGTH - 1 DOWNTO 0 );
   BEGIN
       src_copy   := SrcReg;
       dst_copy   := DstReg;
 -- synopsys translate_off    
    --  Null range Check
    --  if input vector is of zero length
       IF ( SrcReg'LENGTH = 0) THEN
           ASSERT false
           REPORT " RegShift --- input bit_vector   is null  "
           SEVERITY ERROR;
           dst_copy := (OTHERS => FillVal);
           DstReg    := dst_copy;
           ShiftO := '0';
           Return;
       ELSIF (DstReg'LENGTH = 0) THEN
           ASSERT false
           REPORT " RegShift --- output vector is  null  "
           SEVERITY ERROR;
         -- set shift out bit at least
           IF ( direction /= '0') THEN
               ShiftO := src_copy(SrcReg'LENGTH - Nbits);
           ELSE 
               ShiftO := src_copy(Nbits - 1);
           END IF;
           RETURN;
      END IF;
-- synopsys translate_on
    -- None of the registers is null, perform shift operation
      IF (direction /= '0') THEN                                 --  left shift
           RegShift_Left(src_copy, r, ShiftO, FillVal, Nbits);
      ELSE                                                       -- right shift
           RegShift_Right(src_copy, r, ShiftO, FillVal, Nbits);
      END IF;
      -- determine length of the result
      IF (DstReg'LENGTH <= SrcReg'LENGTH) THEN
		for i IN DstReg'Length - 1 downto 0 Loop
			dst_copy(i) := r(i);
                end loop;
      ELSE
		for i IN SrcReg'LENGTH - 1 downto 0 Loop
			dst_copy(i) := r(i);
                end loop;
      END IF;
      DstReg := dst_copy;
      RETURN;
   END RegShift;
--+-----------------------------------------------------------------------------
--|     Function Name  : RegShift
--| 
--|     Overloading    : None
--|
--|     Purpose        : Bidirectional logical shift operator for logic vector.
--|
--|     Parameters     :
--|                      SrcReg      - input  std_ulogic_vector, vector to be shifted
--|                      DstReg      - ouput, std_ulogic_vector, shifted result
--|                      ShiftO      - output, std_ulogic, holds the 
--|                                            last bit shifted out 
--|                                          of register
--|                      direction   - input, Std_ulogic
--|                                         '0'  means right shift
--|                                         '1' | 'X'  means left shift, 
--|                                          default is left shift
--|                      FillVal     - input, Std_ulogic, value to fill register with. 
--|                                          default is '0'
--|                      Nbits       - input , NATURAL, number of positions to shift
--|                                          default is 1.
--|
--|     Result         : Shifted std_ulogic_vector
--|
--|     NOTE           : Defaults not allowed for synthesis.
--|
--|     Use            : VARIABLE acc   : std_ulogic_vector ( 15 DOWNTO 0);
--|                      VARIABLE carry : std_ulogic;
--|
--|                      RegShift ( acc, acc, carry, '1', '0',3 );
--|-----------------------------------------------------------------------------
   PROCEDURE RegShift  ( CONSTANT SrcReg    : IN std_ulogic_vector;
                         VARIABLE DstReg    : INOUT std_ulogic_vector;
                         VARIABLE ShiftO    : OUT std_ulogic; 
                         CONSTANT direction : IN std_ulogic
                     -- synopsys synthesis_off
						      := '1'
                     -- synopsys synthesis_on
                                                            ;
                         CONSTANT FillVal   : IN std_ulogic  
                     -- synopsys synthesis_off
						      := '0'
                     -- synopsys synthesis_on
                                                            ;
                         CONSTANT Nbits     : IN Natural
                     -- synopsys synthesis_off
						       := 1 
                     -- synopsys synthesis_on
                      ) IS 
      VARIABLE r         : STD_ULOGIC_VECTOR (SrcReg'LENGTH - 1 DOWNTO 0);
      VARIABLE src_copy  : STD_ULOGIC_VECTOR (SrcReg'LENGTH - 1 DOWNTO 0 );
      VARIABLE dst_copy  : STD_ULOGIC_VECTOR (DstReg'LENGTH - 1 DOWNTO 0 );
   BEGIN
       src_copy   := SrcReg;
       dst_copy   := DstReg;
 -- synopsys translate_off    
    --  Null range Check
    --  if input vector is of zero length
       IF ( SrcReg'LENGTH = 0) THEN
           ASSERT false
           REPORT " RegShift --- input bit_vector   is null  "
           SEVERITY ERROR;
           dst_copy := (OTHERS => FillVal);
           DstReg    := dst_copy;
           ShiftO := '0';
           Return;
       ELSIF (DstReg'LENGTH = 0) THEN
           ASSERT false
           REPORT " RegShift --- output vector is  null  "
           SEVERITY ERROR;
         -- set shift out bit at least
           IF ( direction /= '0') THEN
               ShiftO := src_copy(SrcReg'LENGTH - Nbits);
           ELSE 
               ShiftO := src_copy(Nbits - 1);
           END IF;
           RETURN;
      END IF;
-- synopsys translate_on
    -- None of the registers is null, perform shift operation
      IF (direction /= '0') THEN                                 --  left shift
           RegShift_Left(src_copy, r, ShiftO, FillVal, Nbits);
      ELSE                                                       -- right shift
           RegShift_Right(src_copy, r, ShiftO, FillVal, Nbits);
      END IF;
      -- determine length of the result
      IF (DstReg'LENGTH <= SrcReg'LENGTH) THEN
		for i IN DstReg'Length - 1 downto 0 Loop
			dst_copy(i) := r(i);
                end loop;
      ELSE
		for i IN SrcReg'LENGTH - 1 downto 0 Loop
			dst_copy(i) := r(i);
                end loop;
      END IF;
      DstReg := dst_copy;
      RETURN;
   END RegShift;
    -------------------------------------------------------------------------------
    --     Function Name  : RegInc
    --
    --     Overloading    : None
    --    
    --     Purpose        : Increment a std_logic_vector by 1.
    --     
    --     Parameters     : 
    --                      SrcReg     - input  std_logic_vector
    --                      SrcRegMode - input  regmode_type, indicating the format of
    --                             the input std_logic_vector.   Default is TwosComp.
    --     
    --     Result         : std_logic_vector ( SrcReg + 1 )
    --
    --     NOTE           : The length of the return vector is the same as the
    --                      the input vector.
    --                      
    --                      Overflow conditions are ignored. UnSigned numbers wrap
    --                      to 0, signed numbers wrap to the largest negative value.
    --     Use            : 
    --                      VARIABLE vect : std_logic_vector ( 3 DOWNTO 0 );
    --                      vect := RegInc ( vect, UnSigned )
    --     
    --     See Also       : RegAdd, RegSub, RegMult, RegDiv, RegInc, RegDec, RegNegate
    -------------------------------------------------------------------------------
    FUNCTION  RegInc  ( CONSTANT SrcReg        :  IN std_logic_vector;
                        CONSTANT SrcRegMode    :  IN regmode_type 
                 -- synopsys synthesis_off
                                                      := DefaultRegMode 
                 -- synopsys synthesis_on
                      ) RETURN std_logic_vector IS
      VARIABLE result  : std_logic_vector(SrcReg'Length - 1 DOWNTO 0);
      VARIABLE reg     : std_logic_vector(SrcReg'Length - 1 DOWNTO 0);
      VARIABLE incby   : std_logic_vector(SrcReg'Length - 1 DOWNTO 0);
      VARIABLE overflo : std_ulogic;
      VARIABLE carry   : std_ulogic;

    BEGIN
      -- synopsys translate_off
      --  if input source register has null range then 
       IF (SrcReg'LENGTH = 0) THEN
           result := SrcReg;
           ASSERT FALSE
           REPORT " RegInc --- Source register has null range "
           SEVERITY ERROR;
           return result;
       END IF;
	-- synopsys translate_on
	--  increment by 1
        reg      := SrcReg;
        incby    := (OTHERS => '0');
        incby(0) := '1';
        RegAdd_Syn(result, reg, incby, SrcRegMode);
	RETURN  To_X01(result);
    END RegInc;
    -------------------------------------------------------------------------------
    --     Function Name  : RegInc
    --
    --     Overloading    : None
    --    
    --     Purpose        : Increment a std_ulogic_vector by 1.
    --     
    --     Parameters     : 
    --                      SrcReg     - input  std_ulogic_vector
    --                      SrcRegMode - input  regmode_type, indicating the format of
    --                             the input std_ulogic_vector.   Default is TwosComp.
    --     
    --     Result         : std_ulogic_vector ( SrcReg + 1 )
    --
    --     NOTE           : The length of the return vector is the same as the
    --                      the input vector.
    --                      
    --                      Overflow conditions are ignored. UnSigned numbers wrap
    --                      to 0, signed numbers wrap to the largest negative value.
    --     Use            : 
    --                      VARIABLE vect : std_ulogic_vector ( 3 DOWNTO 0 );
    --                      vect := RegInc ( vect, UnSigned )
    --     
    --     See Also       : RegAdd, RegSub, RegDec, RegNegate
    -------------------------------------------------------------------------------
    FUNCTION  RegInc  ( CONSTANT SrcReg        :  IN std_ulogic_vector;
                        CONSTANT SrcRegMode    :  IN regmode_type
                 -- synopsys synthesis_off
                                                      := DefaultRegMode 
                 -- synopsys synthesis_on
                      ) RETURN std_ulogic_vector IS
	VARIABLE result  : std_logic_vector(SrcReg'Length - 1 DOWNTO 0);
	VARIABLE reg     : std_logic_vector(SrcReg'Length - 1 DOWNTO 0);
    BEGIN
	reg := To_StdLogicVector(SrcReg);
        result:= RegInc(reg , SrcRegMode);
        return (To_StdULogicVector(result));
    END RegInc;
--+-----------------------------------------------------------------------------
--|     Function Name  : RegInc
--| 
--|     Overloading    : None
--|  
--|     Purpose        : Increment a BIT_VECTOR by 1.
--|  
--|     Parameters     :
--|                      SrcReg     - input  BIT_VECTOR
--|                      SrcRegMode - input  regmode_type, indicating the format of
--|                                the input BIT_VECTOR.   Default is TwosComp.
--|  
--|     Result         : BIT_VECTOR ( SrcReg + 1 )
--| 
--|     NOTE           : The length of the return vector is the same as the
--|                      the input vector.
--|  
--|                      Overflow conditions are ignored. UnSigned numbers wrap
--|                      to 0, signed numbers wrap to the largest negative value.
--|     Use            :
--|                      VARIABLE vect : BIT_VECTOR ( 3 DOWNTO 0 );
--|                      vect := RegInc ( vect, UnSigned )
--| 
--|     See Also       : RegAdd, RegSub, RegMult, RegDiv, RegInc, RegDec, RegNegate
--|-----------------------------------------------------------------------------
    FUNCTION RegInc  ( CONSTANT SrcReg        :  IN BIT_VECTOR;
                       CONSTANT SrcRegMode    :  IN regmode_type
                 -- synopsys synthesis_off
                                                      := DefaultRegMode 
                 -- synopsys synthesis_on
                     ) RETURN BIT_VECTOR IS
	VARIABLE result  : std_logic_vector(SrcReg'Length - 1 DOWNTO 0);
	VARIABLE reg     : std_logic_vector(SrcReg'Length - 1 DOWNTO 0);
    BEGIN
	reg := To_StdLogicVector(SrcReg);
        result := RegInc( reg, SrcRegMode);
	RETURN  To_BitVector(result);
    END RegInc;
    -------------------------------------------------------------------------------
    --     Function Name  : RegDec
    --
    --     Overloading    : None
    --    
    --     Purpose        : Decrement a std_logic_vector by 1.
    --     
    --     Parameters     : 
    --                      SrcReg     - input  std_logic_vector
    --                      SrcRegMode - input  regmode_type, indicating the format of
    --                              the input std_logic_vector.   Default is TwosComp.
    --     
    --     Result         : std_logic_vector ( SrcReg - 1 )
    --
    --     NOTE           : The length of the return vector is the same as the
    --                      the input vector.
    --     Use            : 
    --                      VARIABLE vect : std_logic_vector ( 3 DOWNTO 0 );
    --                      vect := RegDec ( vect, UnSigned )
    --
    --     See Also       : RegAdd, RegSub, RegMult, RegDiv, RegInc, RegDec, RegNegate
    -------------------------------------------------------------------------------
    FUNCTION  RegDec  ( CONSTANT SrcReg        :  IN std_logic_vector;
                        CONSTANT SrcRegMode    :  IN regmode_type
                 -- synopsys synthesis_off
                                                      := DefaultRegMode 
                 -- synopsys synthesis_on
                      ) RETURN std_logic_vector IS
      VARIABLE result    : std_logic_vector(SrcReg'Length - 1 DOWNTO 0);
      VARIABLE  reg      : std_logic_vector(SrcReg'Length - 1 DOWNTO 0);
      VARIABLE decby     : std_logic_vector(SrcReg'Length - 1 DOWNTO 0);
      VARIABLE underflow : std_ulogic;
      VARIABLE borrow    : std_ulogic;
    
    BEGIN
      -- synopsys translate_off
	--  if input source register has null range then 
        IF (SrcReg'LENGTH = 0) THEN
             ASSERT FALSE
             REPORT " RegDec --- Source register has null range "
             SEVERITY ERROR;
             result := SrcReg;
             return result;
	END IF;
      -- synopsys translate_on
	--  decrement by 1
        reg      := SrcReg;
        decby   := (OTHERS => '0');
        decby(0) := '1';        
       	RegSub_Syn(result, reg, decby, SrcRegMode);
	RETURN  To_X01(result);
    END RegDec;
    -------------------------------------------------------------------------------
    --     Function Name  : RegDec
    --
    --     Overloading    : None
    --    
    --     Purpose        : Decrement a std_ulogic_vector by 1.
    --     
    --     Parameters     : 
    --                      SrcReg     - input  std_ulogic_vector
    --                      SrcRegMode - input  regmode_type, indicating the format of
    --                            the input std_ulogic_vector.   Default is TwosComp.
    --     
    --     Result         : std_ulogic_vector ( SrcReg - 1 )
    --
    --     NOTE           : The length of the return vector is the same as the
    --                      the input vector.
    --     Use            : 
    --                      VARIABLE vect : std_ulogic_vector ( 3 DOWNTO 0 );
    --                      vect := RegDec ( vect, UnSigned )
    --     
    --     See Also       : RegAdd, RegSub, RegMult, RegDiv, RegInc, RegDec, RegNegate
    -------------------------------------------------------------------------------
    FUNCTION  RegDec  ( CONSTANT SrcReg        :  IN std_ulogic_vector;
                        CONSTANT SrcRegMode    :  IN regmode_type
                 -- synopsys synthesis_off
                                                      := DefaultRegMode 
                 -- synopsys synthesis_on
                      ) RETURN std_ulogic_vector IS
	VARIABLE result  : std_logic_vector(SrcReg'Length - 1 DOWNTO 0);
	VARIABLE reg     : std_logic_vector(SrcReg'Length - 1 DOWNTO 0);
    BEGIN
	reg := To_StdLogicVector(SrcReg);
        result:= RegDec(reg , SrcRegMode);
        return (To_StdULogicVector(result));
    END RegDec;
--+-----------------------------------------------------------------------------
--|     Function Name  : RegDec
--|
--|     Overloading    : None
--| 
--|     Purpose        : Decrement a BIT_VECTOR by 1.
--| 
--|     Parameters     :
--|                      SrcReg     - input  BIT_VECTOR
--|                      SrcRegMode - input  regmode_type, indicating the format of
--|                                the input BIT_VECTOR.   Default is TwosComp.
--| 
--|     Result         : BIT_VECTOR ( SrcReg - 1 )
--|
--|     NOTE           : The length of the return vector is the same as the
--|                      the input vector.
--|     Use            :
--|                      VARIABLE vect : BIT_VECTOR ( 3 DOWNTO 0 );
--|                      vect := RegDec ( vect, UnSigned )
--| 
--|     See Also       : RegAdd, RegSub, RegMult, RegDiv, RegInc, RegDec, RegNegate
--|-----------------------------------------------------------------------------
    FUNCTION RegDec  ( CONSTANT SrcReg        :  IN BIT_VECTOR;
                       CONSTANT SrcRegMode    :  IN regmode_type
                 -- synopsys synthesis_off
                                                      := DefaultRegMode 
                 -- synopsys synthesis_on
                     ) RETURN BIT_VECTOR IS

	VARIABLE result  : std_logic_vector(SrcReg'Length - 1 DOWNTO 0);
	VARIABLE reg     : std_logic_vector(SrcReg'Length - 1 DOWNTO 0);
    BEGIN
	reg := To_StdLogicVector(SrcReg);
        result:= RegDec(reg , SrcRegMode);
        return (To_BitVector(result));
   END RegDec;
    -------------------------------------------------------------------------------
    --     Function Name  : RegNegate
    --
    --     Overloading    : None
    --    
    --     Purpose        : Negate a std_logic_vector ( v := 0 - v )
    --     
    --     Parameters     : 
    --                      SrcReg     - input  std_logic_vector
    --                      SrcRegMode - input  regmode_type, indicating the format of
    --                                the input std_logic_vector.   Default is TwosComp.
    --     
    --     Result         : std_logic_vector ( 0 - SrcReg )
    --
    --     NOTE           : The length of the return vector is the same as the
    --                      the input vector.
    --                      
    --                      If 'SrcRegMode' is UnSigned the bitwise NOT of 'SrcReg'
    --                      is returned.
    --
    --                      An overflow can occur when 'SrcRegMode' is TwosComp and
    --                      'SrcReg' is the largest negative value (ie "100...00").
    --                      In this case NO error is indicated and the returned
    --                      value is the same as the input.
    --     Use            : 
    --                      VARIABLE vect : std_logic_vector (15 DOWNTO 0 );
    --                      vect := RegNegate ( vect, TwosComp );
    --                      vect := RegNegate ( vect );
    --     
    --     See Also       : RegAdd, RegSub, RegMult, RegDiv, RegInc, RegDec, RegNegate
    -------------------------------------------------------------------------------
    FUNCTION  RegNegate  ( CONSTANT SrcReg     :  IN std_logic_vector;
                           CONSTANT SrcRegMode :  IN regmode_type := DefaultRegMode
                         ) RETURN std_logic_vector IS
      VARIABLE result : std_logic_vector(SrcReg'Length - 1 DOWNTO 0);
      VARIABLE by_one : std_logic_vector(SrcReg'Length - 1 DOWNTO 0);
    BEGIN
    -- check for null range of SrcReg 
      IF (SrcReg'LENGTH = 0) THEN
	-- synopsys translate_off
         ASSERT false
          REPORT " RegNegate --- source register has null range "
          SEVERITY ERROR; 
        -- synopsys translate_on
          result := SrcReg;
          return (result);
      END IF;

      result := NOT SrcReg;
      IF (SrcRegMode = TwosComp) THEN
	 by_one := (OTHERS => '0');
         by_one(0) := '1';
         return (Add_TwosComp(result, by_one)); 
      ELSE   
         return(result);
      END IF;
    END RegNegate;
    -------------------------------------------------------------------------------
    --     Function Name  : RegNegate
    --
    --     Overloading    : None
    --    
    --     Purpose        : Negate a std_ulogic_vector ( v := 0 - v )
    --     
    --     Parameters     : 
    --                      SrcReg     - input  std_ulogic_vector
    --                      SrcRegMode - input  regmode_type, indicating the format of
    --                                the input std_ulogic_vector.   Default is TwosComp.
    --     
    --     Result         : std_ulogic_vector ( 0 - SrcReg )
    --
    --     NOTE           : The length of the return vector is the same as the
    --                      the input vector.
    --                      
    --                      If 'SrcRegMode' is UnSigned the bitwise NOT of 'SrcReg'
    --                      is returned.
    --
    --                      An overflow can occur when 'SrcRegMode' is TwosComp and
    --                      'SrcReg' is the largest negative value (ie "100...00").
    --                      In this case NO error is indicated and the returned
    --                      value is the same as the input.
    --     Use            : 
    --                      VARIABLE vect : std_ulogic_vector (15 DOWNTO 0 );
    --                      vect := RegNegate ( vect, TwosComp );
    --                      vect := RegNegate ( vect );
    --     
    --     See Also       : RegAdd, RegSub, RegMult, RegDiv, RegInc, RegDec, RegNegate
    -------------------------------------------------------------------------------
    FUNCTION  RegNegate  ( CONSTANT SrcReg     :  IN std_ulogic_vector;
                           CONSTANT SrcRegMode :  IN regmode_type := DefaultRegMode
                         ) RETURN std_ulogic_vector IS
        VARIABLE reslt   : std_logic_vector(SrcReg'Length - 1 DOWNTO 0);
	VARIABLE reg     : std_logic_vector(SrcReg'Length - 1 DOWNTO 0);
    BEGIN
	reg := To_StdLogicVector(SrcReg);
	reslt := RegNegate(reg, SrcRegMode);
        return To_StdULogicVector(reslt);
    END RegNegate;
--+-----------------------------------------------------------------------------
--|     Function Name  : RegNegate
--|
--|     Overloading    : None
--|
--|     Purpose        : Negate a BIT_VECTOR ( v := 0 - v )
--|
--|     Parameters     :
--|                      SrcReg     - input  BIT_VECTOR
--|                      SrcRegMode - input  regmode_type, indicating the format of
--|                                the input BIT_VECTOR.   Default is TwosComp.
--|
--|     Result         : BIT_VECTOR ( 0 - SrcReg )
--|
--|     NOTE           : The length of the return vector is the same as the
--|                      the input vector.
--|
--|                      If 'SrcRegMode' is UnSigned the bitwise NOT of 'SrcReg'
--|                      is returned.
--|
--|                      An overflow can occur when 'SrcRegMode' is TwosComp and
--|                      'SrcReg' is the largest negative value (ie "100...00").
--|                      In this case NO error is indicated and the returned
--|                      value is the same as the input.
--|     Use            :
--|                      VARIABLE vect : BIT_VECTOR (15 DOWNTO 0 );
--|                      vect := RegNegate ( vect, TwosComp );
--|
--|     See Also       : RegAdd, RegSub, RegMult, RegDiv, RegInc, RegDec, RegNegate
--|-----------------------------------------------------------------------------
    FUNCTION RegNegate  ( CONSTANT SrcReg      :  IN BIT_VECTOR;
                          CONSTANT SrcRegMode  :  IN regmode_type 
                 -- synopsys synthesis_off
                                                     := DefaultRegMode
                 -- synopsys synthesis_on
                        ) RETURN BIT_VECTOR IS
        VARIABLE reslt : STD_LOGIC_VECTOR(SrcReg'Length - 1 DOWNTO 0);
	VARIABLE reg     : std_logic_vector(SrcReg'Length - 1 DOWNTO 0);
    BEGIN
	reg := To_StdLogicVector(SrcReg);
        reslt := RegNegate(reg, SrcRegMode);
        return (To_BitVector(reslt));
    END RegNegate;

    -- ----------------------------------------------------------------------------
    -- ----------------------------------------------------------------------------
    --    Adding procedure to handle signals
    -- ----------------------------------------------------------------------------
    -------------------------------------------------------------------------------
    --     Procedure Name : SregAbs
    -- 1.6.9
    --     Overloading    : Procedure .
    --
    --     Purpose        : converts  std_logic_vector into an absolute value.
    --
    --     Parameters     :
    --                      result     - input-output  std_logic_vector, 
    --                      SrcReg     - input  std_logic_vector, the vector to be read.
    --                      SrcRegMode - input  regmode_type, indicating the format of
    --                                the input std_logic_vector.   Default is TwosComp.
    --
    --     Use            :
    --                      SIGNAL reslt, vect : std_logic_vector ( 15 DOWNTO 0 );
    --
    --                       SregAbs ( reslt,  vect, TwosComp );
    -------------------------------------------------------------------------------
    PROCEDURE SregAbs  ( SIGNAL result     : INOUT std_logic_vector;
                        CONSTANT SrcReg     : IN std_logic_vector;
                        CONSTANT SrcRegMode : IN regmode_type 
                     -- synopsys synthesis_off
						      := DefaultRegMode 
                     -- synopsys synthesis_on
                      ) IS
       VARIABLE reslt_copy : std_logic_vector (result'LENGTH - 1 DOWNTO 0);
    BEGIN
	RegAbs(reslt_copy, SrcReg, SrcRegMode);
        result    <= reslt_copy 
                     -- synopsys synthesis_off
				after DefaultRegDelay
                     -- synopsys synthesis_on
                                                    ;
        return;
    END SregAbs;
    -------------------------------------------------------------------------------
    --     Procedure Name : SregAbs
    -- 1.6.9
    --     Overloading    : Procedure .
    --
    --     Purpose        : converts  std_ulogic_vector into an absolute value.
    --
    --     Parameters     :
    --                      result     - input-output  std_ulogic_vector, 
    --                      SrcReg     - input  std_ulogic_vector, the vector to be read.
    --                      SrcRegMode - input  regmode_type, indicating the format of
    --                                the input std_ulogic_vector.   Default is TwosComp.
    --
    --     Use            :
    --                      SIGNAL reslt, vect : std_ulogic_vector ( 15 DOWNTO 0 );
    --
    --                       SregAbs ( reslt,  vect, TwosComp );
    -------------------------------------------------------------------------------
    PROCEDURE SregAbs  ( SIGNAL result     : INOUT std_ulogic_vector;
                        CONSTANT SrcReg     : IN std_ulogic_vector;
                        CONSTANT SrcRegMode : IN regmode_type 
                     -- synopsys synthesis_off
						      := DefaultRegMode 
                     -- synopsys synthesis_on
                      ) IS
       VARIABLE reslt_copy : std_logic_vector (result'LENGTH - 1 DOWNTO 0);
    BEGIN
	RegAbs(reslt_copy, To_StdLogicVector(SrcReg), SrcRegMode);
        result    <= To_StdULogicVector(reslt_copy)
                     -- synopsys synthesis_off
						after DefaultRegDelay
                     -- synopsys synthesis_on
                        		                            ;
        return;
    END SregAbs;
    -------------------------------------------------------------------------------
    --     Procedure Name : SregAbs
    -- 1.6.9
    --     Overloading    : Procedure .
    --
    --     Purpose        : converts  bit_vector into an absolute value.
    --
    --     Parameters     :
    --                      result     - input-output  bit_vector, 
    --                      SrcReg     - input  bit_vector, the vector to be read.
    --                      SrcRegMode - input  regmode_type, indicating the format of
    --                                the input bit_vector.   Default is TwosComp.
    --
    --     Use            :
    --                      SIGNAL reslt, vect : bit_vector ( 15 DOWNTO 0 );
    --
    --                       SregAbs ( reslt,  vect, TwosComp );
    -------------------------------------------------------------------------------
    PROCEDURE SregAbs  ( SIGNAL result     : INOUT bit_vector;
                        CONSTANT SrcReg     : IN bit_vector;
                        CONSTANT SrcRegMode : IN regmode_type 
                     -- synopsys synthesis_off
						      := DefaultRegMode 
                     -- synopsys synthesis_on
                      ) IS

       VARIABLE reslt_copy : std_logic_vector (result'LENGTH - 1 DOWNTO 0);
    BEGIN
	RegAbs(reslt_copy, To_StdLogicVector(SrcReg), SrcRegMode);
        result    <= To_BitVector(reslt_copy)
                     -- synopsys synthesis_off
             				after DefaultRegDelay
                     -- synopsys synthesis_on
                                                             ;
        return;
    END SregAbs;
--+-----------------------------------------------------------------------------
--|     Function Name  : SregAdd
--|
--|     Overloading    : None
--|
--|     Purpose        : Addition of STD_LOGIC_VECTORS.
--|
--|     Parameters     :
--|                      result     - input-output STD_LOGIC_VECTOR, the computed sum
--|                      carry_out  - output STD_ULOGIC,
--|                      overflow   - output STD_ULOGIC, overflow condition
--|                      addend     - input  STD_LOGIC_VECTOR,
--|                      augend     - input  STD_LOGIC_VECTOR,
--|                      carry_in   - input  STD_ULOGIC,  
--|                      SrcRegMode - input  regmode_type, indicating the format of
--|                                the input STD_LOGIC_VECTOR.   Default is TwosComp.
--|     NOTE           :
--|                      The inputs may be of any length and may be of differing
--|                      lengths.
--| 
--|                    For Synthesis:
--|                      Result is computed with length N (where
--|                      N is the greater of the input vector lengths).
--|                      It is assumed that user will provide result length equal
--|                      to the length of the greater of addend and augend. 
--|                      No error checking has been performed.
--|     Use            :
--|                      SIGNAL x, y, sum : STD_LOGIC_VECTOR ( 15 DOWNTO 0);
--|                      SIGNAL carry_in, carry_out , ovf: STD_ULOGIC;
--| 
--|                      SregAdd ( sum, carry_out, ovf,x, y, carry_in, UnSigned );
--| 
--|     See Also       : SregSub, SregMult, SregDiv
--|-----------------------------------------------------------------------------
    PROCEDURE SregAdd  (SIGNAL result       : INOUT STD_LOGIC_VECTOR;
                        SIGNAL carry_out    : OUT STD_ULOGIC;
                        SIGNAL overflow     : OUT STD_ULOGIC;
                        CONSTANT addend     : IN STD_LOGIC_VECTOR;
                        CONSTANT augend     : IN STD_LOGIC_VECTOR;
                        CONSTANT carry_in   : IN STD_ULOGIC;
                        CONSTANT SrcRegMode : IN regmode_type
                  -- synopsys synthesis_off
                                                       := DefaultRegMode 
                   -- synopsys synthesis_on
                      ) IS

       VARIABLE reslt_copy  : STD_LOGIC_VECTOR ( result'length-1 downto 0 );
       VARIABLE a_copy      : STD_LOGIC_VECTOR ( addend'length-1 downto 0 );
       VARIABLE b_copy      : STD_LOGIC_VECTOR ( augend'length-1 downto 0 );
       VARIABLE carry_loc    : std_ulogic; 
       VARIABLE overflow_loc : std_ulogic;
     BEGIN 
	RegAdd(reslt_copy, carry_loc, overflow_loc, addend, augend, carry_in, SrcRegMode);

        result    <=  reslt_copy
                     -- synopsys synthesis_off
             				after DefaultRegDelay
                     -- synopsys synthesis_on
                                                             ;
        carry_out <= carry_loc 
                     -- synopsys synthesis_off
             				after DefaultRegDelay
                     -- synopsys synthesis_on
                                                             ;
        overflow <= overflow_loc
                     -- synopsys synthesis_off
             				after DefaultRegDelay
                     -- synopsys synthesis_on
                                                             ;
        return;
     END SregAdd;
--+-----------------------------------------------------------------------------
--|     Function Name  : SregAdd
--|
--|     Overloading    : None
--|
--|     Purpose        : Addition of STD_ULOGIC_VECTORS.
--|
--|     Parameters     :
--|                      result     - input-output STD_ULOGIC_VECTOR, the computed sum
--|                      carry_out  - output STD_ULOGIC,
--|                      overflow   - output STD_ULOGIC, overflow condition
--|                      addend     - input  STD_ULOGIC_VECTOR,
--|                      augend     - input  STD_ULOGIC_VECTOR,
--|                      carry_in   - input  STD_ULOGIC,  
--|                      SrcRegMode - input  regmode_type, indicating the format of
--|                                the input STD_ULOGIC_VECTOR.   Default is TwosComp.
--|     NOTE           :
--|                      The inputs may be of any length and may be of differing
--|                      lengths.
--| 
--|                    For Synthesis:
--|                      Result is computed with length N (where
--|                      N is the greater of the input vector lengths).
--|                      It is assumed that user will provide result length equal
--|                      to the length of the greater of addend and augend. 
--|                      No error checking has been performed.
--|     Use            :
--|                      SIGNAL x, y, sum : STD_ULOGIC_VECTOR ( 15 DOWNTO 0);
--|                      SIGNAL carry_in, carry_out , ovf: STD_ULOGIC;
--| 
--|                      SregAdd ( sum, carry_out, ovf,x, y, carry_in, UnSigned );
--| 
--|     See Also       : SregSub, SregMult, SregDiv
--|-----------------------------------------------------------------------------
    PROCEDURE SregAdd  (SIGNAL result       : INOUT STD_ULOGIC_VECTOR;
                        SIGNAL carry_out    : OUT STD_ULOGIC;
                        SIGNAL overflow     : OUT STD_ULOGIC;
                        CONSTANT addend     : IN STD_ULOGIC_VECTOR;
                        CONSTANT augend     : IN STD_ULOGIC_VECTOR;
                        CONSTANT carry_in   : IN STD_ULOGIC;
                        CONSTANT SrcRegMode : IN regmode_type
                  -- synopsys synthesis_off
                                                       := DefaultRegMode 
                   -- synopsys synthesis_on
                      ) IS
       VARIABLE reslt_copy  : STD_LOGIC_VECTOR ( result'length-1 downto 0 );
       VARIABLE a_copy      : STD_LOGIC_VECTOR ( addend'length-1 downto 0 );
       VARIABLE b_copy      : STD_LOGIC_VECTOR ( augend'length-1 downto 0 );
       VARIABLE carry_loc    : std_ulogic; 
       VARIABLE overflow_loc : std_ulogic;

     BEGIN 
	a_copy := To_StdLogicVector(addend);
	b_copy := To_StdLogicVector(augend);

	RegAdd(reslt_copy, carry_loc, overflow_loc, a_copy, b_copy, carry_in, SrcRegMode);

        result    <= To_StdULogicVector(reslt_copy) 
                     -- synopsys synthesis_off
             				after DefaultRegDelay
                     -- synopsys synthesis_on
                                                             ;
        carry_out <= carry_loc 
                     -- synopsys synthesis_off
             				after DefaultRegDelay
                     -- synopsys synthesis_on
                                                             ;
        overflow <= overflow_loc
                     -- synopsys synthesis_off
             				after DefaultRegDelay
                     -- synopsys synthesis_on
                                                             ;
        return;
     END SregAdd;
--+-----------------------------------------------------------------------------
--|     Function Name  : SregAdd
--|
--|     Overloading    : None
--|
--|     Purpose        : Addition of BIT_VECTORS.
--|
--|     Parameters     :
--|                      result     - input-output BIT_VECTOR, the computed sum
--|                      carry_out  - output BIT,
--|                      overflow   - output BIT, overflow condition
--|                      addend     - input  BIT_VECTOR,
--|                      augend     - input  BIT_VECTOR,
--|                      carry_in   - input  BIT,  
--|                      SrcRegMode - input  regmode_type, indicating the format of
--|                                the input BIT_VECTOR.   Default is TwosComp.
--|     NOTE           :
--|                      The inputs may be of any length and may be of differing
--|                      lengths.
--|
--|                    For Synthesis:
--|                      Result is computed with length N (where
--|                      N is the greater of the input vector lengths).
--|                      It is assumed that user will provide result length equal
--|                      to the length of the greater of addend and augend. 
--|                      No error checking has been performed.
--|     Use            :
--|                      SIGNAL x, y, sum : BIT_VECTOR ( 15 DOWNTO 0);
--|                      SIGNAL carry_in, carry_out , ovf: BIT;
--| 
--|                      SregAdd ( sum, carry_out, ovf,x, y, carry_in, UnSigned );
--| 
--|     See Also       : SregSub, SregMult, SregDiv
--|-----------------------------------------------------------------------------
    PROCEDURE SregAdd  (SIGNAL result       : INOUT BIT_VECTOR;
                        SIGNAL carry_out    : OUT BIT;
                        SIGNAL overflow     : OUT BIT;
                        CONSTANT addend     : IN BIT_VECTOR;
                        CONSTANT augend     : IN BIT_VECTOR;
                        CONSTANT carry_in   : IN BIT;
                        CONSTANT SrcRegMode : IN regmode_type
                  -- synopsys synthesis_off
                                                       := DefaultRegMode 
                   -- synopsys synthesis_on
                      ) IS
       VARIABLE reslt_copy  : std_logic_vector ( result'length-1 downto 0 );
       VARIABLE carry_loc    : std_ulogic; 
       VARIABLE overflow_loc : std_ulogic;
       VARIABLE a_copy      : STD_LOGIC_VECTOR ( addend'length-1 downto 0 );
       VARIABLE b_copy      : STD_LOGIC_VECTOR ( augend'length-1 downto 0 );
       VARIABLE c_in        : std_ulogic; 
     BEGIN 
	a_copy := To_StdLogicVector(addend);
	b_copy := To_StdLogicVector(augend);
        c_in   := To_StdULogic(carry_in);

	RegAdd(reslt_copy, carry_loc, overflow_loc, a_copy, b_copy, c_in, SrcRegMode);
        result    <= To_BitVector(reslt_copy)
                     -- synopsys synthesis_off
             				after DefaultRegDelay
                     -- synopsys synthesis_on
                                                             ;
        carry_out <= To_Bit(carry_loc)
                     -- synopsys synthesis_off
             				after DefaultRegDelay
                     -- synopsys synthesis_on
                                                             ;
        overflow  <= To_Bit(overflow_loc)
                     -- synopsys synthesis_off
             				after DefaultRegDelay
                     -- synopsys synthesis_on
                                                             ;
        return;
     END SregAdd;
--+-----------------------------------------------------------------------------
--|     Function Name  : SregSub
--|    
--|     Overloading    : None
--|
--|     Purpose        : Subtraction of STD_LOGIC_VECTORS.
--|                       ( result = minuend - subtrahend )
--|
--|     Parameters     :
--|                      result     - input-output STD_LOGIC_VECTOR, the computed sum
--|                      borrow_out - output STD_ULOGIC,
--|                      overflow   - output STD_ULOGIC, overflow condition
--|                      minuend - input  STD_LOGIC_VECTOR,
--|                      subtrahend - input  STD_LOGIC_VECTOR,
--|                      borrow_in  - input  STD_LOGIC, borrow from the LSB
--|                      SrcRegMode - input  regmode_type, indicating the format of
--|                                the input STD_LOGIC_VECTOR.   Default is TwosComp.
--|     NOTE           :
--|                      The inputs may be of any length and may be of differing
--|                      lengths.
--|
--|                      A  result is computed with length N (where
--|                      N is the greater of the input vector lengths).
--|     Use            :
--|                      SIGNAL x, y, diff : STD_LOGIC_VECTOR ( 15 DOWNTO 0);
--|                      SIGNAL n_borrow, borrow_in : STD_ULOGIC;
--|
--|                      SregSub ( diff, n_borrow, x, y, borrow_in, UnSigned );
--|
--|     See Also       : SregAdd,  SregMult, SregDiv
--|-----------------------------------------------------------------------------
    PROCEDURE SregSub  (SIGNAL result       : INOUT STD_LOGIC_VECTOR;
                        SIGNAL borrow_out   : OUT STD_ULOGIC;
                        SIGNAL overflow     : OUT STD_ULOGIC;
                        CONSTANT minuend    :  IN STD_LOGIC_VECTOR;
                        CONSTANT subtrahend :  IN STD_LOGIC_VECTOR;
                        CONSTANT borrow_in  :  IN STD_ULOGIC  
                  -- synopsys synthesis_off
                                                       := '0'
                  -- synopsys synthesis_on
                                                               ;
                        CONSTANT SrcRegMode :  IN regmode_type
                  -- synopsys synthesis_off
                                                       := DefaultRegMode 
                   -- synopsys synthesis_on
                      ) IS
	VARIABLE reslt_copy   : STD_LOGIC_VECTOR ( result'length-1 downto 0 ); 
	VARIABLE borrow_loc   : std_ulogic;
	VARIABLE overflow_loc : std_ulogic;
     BEGIN 

	RegSub(reslt_copy, borrow_loc, overflow_loc, minuend, subtrahend, borrow_in, SrcRegMode);

        result     <= reslt_copy 
                     -- synopsys synthesis_off
             				after DefaultRegDelay
                     -- synopsys synthesis_on
                                                             ;
        borrow_out <= borrow_loc
                     -- synopsys synthesis_off
             				after DefaultRegDelay
                     -- synopsys synthesis_on
                                                             ;
        overflow   <= overflow_loc
                     -- synopsys synthesis_off
             				after DefaultRegDelay
                     -- synopsys synthesis_on
                                                             ;
        RETURN;
    END SregSub;
--+-----------------------------------------------------------------------------
--|     Function Name  : SregSub
--|    
--|     Overloading    : None
--|
--|     Purpose        : Subtraction of STD_ULOGIC_VECTORS.
--|                       ( result = minuend - subtrahend )
--|
--|     Parameters     :
--|                      result     - input-output STD_ULOGIC_VECTOR, the computed sum
--|                      borrow_out - output STD_ULOGIC,
--|                      overflow   - output STD_ULOGIC, overflow condition
--|                      minuend - input  STD_ULOGIC_VECTOR,
--|                      subtrahend - input  STD_ULOGIC_VECTOR,
--|                      borrow_in  - input  STD_ULOGIC, borrow from the LSB
--|                      SrcRegMode - input  regmode_type, indicating the format of
--|                                the input STD_ULOGIC_VECTOR.   Default is TwosComp.
--|
--|     NOTE           :
--|                      The inputs may be of any length and may be of differing
--|                      lengths.
--|
--|                      A  result is computed with length N (where
--|                      N is the greater of the input vector lengths).
--|     Use            :
--|                      SIGNAL x, y, diff : STD_ULOGIC_VECTOR ( 15 DOWNTO 0);
--|                      SIGNAL n_borrow, borrow_in : STD_ULOGIC;
--|
--|                      SregSub ( diff, n_borrow, x, y, borrow_in, UnSigned );
--|
--|     See Also       : SregAdd,  SregMult, SregDiv
--|-----------------------------------------------------------------------------
    PROCEDURE SregSub  (SIGNAL result       : INOUT STD_ULOGIC_VECTOR;
                        SIGNAL borrow_out   : OUT STD_ULOGIC;
                        SIGNAL overflow     : OUT STD_ULOGIC;
                        CONSTANT minuend    :  IN STD_ULOGIC_VECTOR;
                        CONSTANT subtrahend :  IN STD_ULOGIC_VECTOR;
                        CONSTANT borrow_in  :  IN STD_ULOGIC  
                  -- synopsys synthesis_off
                                                       := '0'
                  -- synopsys synthesis_on
                                                               ;
                        CONSTANT SrcRegMode :  IN regmode_type
                  -- synopsys synthesis_off
                                                       := DefaultRegMode 
                   -- synopsys synthesis_on
                      ) IS
	VARIABLE reslt_copy   : STD_LOGIC_VECTOR ( result'length-1 downto 0 ); 
	VARIABLE borrow_loc   : std_ulogic;
	VARIABLE overflow_loc : std_ulogic;
	VARIABLE a_copy      : STD_LOGIC_VECTOR ( minuend'length-1 downto 0 );
	VARIABLE b_copy      : STD_LOGIC_VECTOR ( subtrahend'length-1 downto 0 );
     BEGIN 
	a_copy := To_StdLogicVector(minuend);
	b_copy := To_StdLogicVector(subtrahend);

	RegSub(reslt_copy, borrow_loc, overflow_loc, a_copy, b_copy, borrow_in, SrcRegMode);

        result     <= To_StdULogicVector(reslt_copy)
                     -- synopsys synthesis_off
             				after DefaultRegDelay
                     -- synopsys synthesis_on
                                                             ;
        borrow_out <= borrow_loc
                     -- synopsys synthesis_off
             				after DefaultRegDelay
                     -- synopsys synthesis_on
                                                             ;
        overflow   <= overflow_loc 
                     -- synopsys synthesis_off
             				after DefaultRegDelay
                     -- synopsys synthesis_on
                                                             ;
        RETURN;
    END SregSub;
--+-----------------------------------------------------------------------------
--|     Function Name  : SregSub
--|    
--|     Overloading    : None
--|
--|     Purpose        : Subtraction of BIT_VECTORS.
--|                       ( result = minuend - subtrahend )
--|
--|     Parameters     :
--|                      result     - input-output BIT_VECTOR, the computed sum
--|                      borrow_out - output BIT,
--|                      overflow   - output BIT, overflow condition
--|                      minuend - input  BIT_VECTOR,
--|                      subtrahend - input  BIT_VECTOR,
--|                      borrow_in  - input  BIT, borrow from the LSB
--|                      SrcRegMode - input  regmode_type, indicating the format of
--|                                the input BIT_VECTOR.   Default is TwosComp.
--|     NOTE           :
--|                      The inputs may be of any length and may be of differing
--|                      lengths.
--|
--|                      Result is computed with length N (where
--|                      N is the greater of the input vector lengths).
--|     Use            :
--|                      SIGNAL x, y, diff : BIT_VECTOR ( 15 DOWNTO 0);
--|                      SIGNAL n_borrow, borrow_in : BIT;
--|
--|                      SregSub ( diff, n_borrow, x, y, borrow_in, UnSigned );
--|
--|     See Also       : SregAdd,  SregMult, SregDiv
--|-----------------------------------------------------------------------------
    PROCEDURE SregSub  (SIGNAL result       : INOUT BIT_VECTOR;
                        SIGNAL borrow_out   : OUT BIT;
                        SIGNAL overflow     : OUT BIT;
                        CONSTANT minuend    :  IN BIT_VECTOR;
                        CONSTANT subtrahend :  IN BIT_VECTOR;
                        CONSTANT borrow_in  :  IN BIT  
                  -- synopsys synthesis_off
                                                       := '0'
                  -- synopsys synthesis_on
                                                               ;
                        CONSTANT SrcRegMode :  IN regmode_type
                  -- synopsys synthesis_off
                                                       := DefaultRegMode 
                   -- synopsys synthesis_on
                        ) IS
        VARIABLE reslt_copy   : std_logic_vector ( result'length-1 downto 0 ); 
        VARIABLE borrow_loc   : std_ulogic;
        VARIABLE overflow_loc : std_ulogic;
	VARIABLE b_in        : std_ulogic;
	VARIABLE a_copy      : STD_LOGIC_VECTOR ( minuend'length-1 downto 0 );
	VARIABLE b_copy      : STD_LOGIC_VECTOR ( subtrahend'length-1 downto 0 );
     BEGIN 
	a_copy := To_StdLogicVector(minuend);
	b_copy := To_StdLogicVector(subtrahend);
        b_in   := To_StdULogic(borrow_in);

	RegSub(reslt_copy, borrow_loc, overflow_loc, a_copy, b_copy, b_in, SrcRegMode);

        result    <= To_BitVector(reslt_copy)
                     -- synopsys synthesis_off
             				after DefaultRegDelay
                     -- synopsys synthesis_on
                                                             ;
        borrow_out <= To_Bit(borrow_loc) 
                     -- synopsys synthesis_off
             				after DefaultRegDelay
                     -- synopsys synthesis_on
                                                             ;
        overflow  <= To_Bit(overflow_loc)
                     -- synopsys synthesis_off
             				after DefaultRegDelay
                     -- synopsys synthesis_on
                                                             ;
        return;
    END SregSub;
--+-----------------------------------------------------------------------------
--|     Function Name  : SregMult
--|
--|     Overloading    : None
--|
--|     Purpose        : Multiplication of STD_LOGIC_VECTORS.
--|
--|     Parameters     :
--|                      result       - output STD_LOGIC_VECTOR, the computed product
--|                      overflow     - output STD_ULOGIC, overflow condition
--|                      multiplicand - input STD_LOGIC_VECTOR,
--|                      multiplier   -  input STD_LOGIC_VECTOR,
--|                      SrcRegMode   - input  regmode_type, indicating the format 
--|                                     of the input STD_LOGIC_VECTOR.   Default is 
--|                                     DefaultRegMode which is set to TwosComp.
--|     NOTE           :
--|                      The inputs may be of any length and may be of differing
--|                      lengths.
--|
--|    Algorithm       : The multiplication is carried out as follows:
--|
--|                      1) Determine sign of result based on sign of 
--|                         multiploicand and sign  of multiplier.
--|
--|                      2) Convert the multiplicand amd multiplier to Unsigned 
--|                         representation.
--|                      
--|                      3) Perform multiplication based on add and shift algorithm.
--|
--|                      4) Convert the result to the SrcRegMode with appropropriate sign
--|
--|     Result         :
--|                     A  temporary result is computed with length N+M (where
--|                      N,M are the lengths of the multiplicand and multiplier).
--|                      This computed value is extended or truncated to match
--|                      the width of 'result'. If truncated, the low order std_ulogics
--|                      are returned.
--|
--|                      The parameter 'overflow' is set to '1' if the product of the
--|                      of the two inputs too large to fit in the parameter result.
--|     Use            :
--|                      SIGNAL x, y, prod : STD_LOGIC_VECTOR ( 15 DOWNTO 0);
--|                      SIGNAL ovfl : STD_ULOGIC;
--|
--|                      SregMult ( prod, ovfl, x, y, TwosComp );
--|
--|     See Also       : RegAdd, SregSub, SregMult, RegDiv, RegInc, RegDec, RegNegate
--|-----------------------------------------------------------------------------
    PROCEDURE SregMult (SIGNAL result         : OUT STD_LOGIC_VECTOR;
                        SIGNAL overflow       : OUT STD_ULOGIC;
                        CONSTANT multiplicand : IN STD_LOGIC_VECTOR;
                        CONSTANT multiplier   : IN STD_LOGIC_VECTOR;
                        CONSTANT SrcRegMode   : IN regmode_type 
                  -- synopsys synthesis_off
                                                       := DefaultRegMode 
                   -- synopsys synthesis_on
                      ) IS
      VARIABLE reslt_copy  : STD_LOGIC_VECTOR ( result'length  - 1  DOWNTO 0 );
      VARIABLE overflo     : STD_ULOGIC;
     BEGIN 
	RegMult(reslt_copy, overflo, multiplicand, multiplier, SrcRegMode);

        result <= reslt_copy 
                     -- synopsys synthesis_off
             				after DefaultRegDelay
                     -- synopsys synthesis_on
                                                             ;
        overflow <= overflo 
                     -- synopsys synthesis_off
             				after DefaultRegDelay
                     -- synopsys synthesis_on
                                                             ;
        RETURN;
    END SregMult;
--+-----------------------------------------------------------------------------
--|     Function Name  : SregMult
--|
--|     Overloading    : None
--|
--|     Purpose        : Multiplication of STD_ULOGIC_VECTORS.
--|
--|     Parameters     :
--|                      result       - output STD_ULOGIC_VECTOR, the computed product
--|                      overflow     - output STD_ULOGIC, overflow condition
--|                      multiplicand - input STD_ULOGIC_VECTOR,
--|                      multiplier   -  input STD_ULOGIC_VECTOR,
--|                      SrcRegMode   - input  regmode_type, indicating the format 
--|                                     of the input STD_ULOGIC_VECTOR.   Default is 
--|                                     DefaultRegMode which is set to TwosComp.
--|     NOTE           :
--|                      The inputs may be of any length and may be of differing
--|                      lengths.
--|
--|    Algorithm       : The multiplication is carried out as follows:
--|
--|                      1) Determine sign of result based on sign of 
--|                         multiploicand and sign  of multiplier.
--|
--|                      2) Convert the multiplicand amd multiplier to Unsigned 
--|                         representation.
--|                      
--|                      3) Perform multiplication based on add and shift algorithm.
--|
--|                      4) Convert the result to the SrcRegMode with appropropriate sign
--|
--|     Result         :
--|                     A  temporary result is computed with length N+M (where
--|                      N,M are the lengths of the multiplicand and multiplier).
--|                      This computed value is extended or truncated to match
--|                      the width of 'result'. If truncated, the low order std_ulogics
--|                      are returned.
--|
--|                      The parameter 'overflow' is set to '1' if the product of the
--|                      of the two inputs too large to fit in the parameter result.
--|     Use            :
--|                      SIGNAL x, y, prod : STD_ULOGIC_VECTOR ( 15 DOWNTO 0);
--|                      SIGNAL ovfl : STD_ULOGIC;
--|
--|                      SregMult ( prod, ovfl, x, y, TwosComp );
--|
--|     See Also       : RegAdd, SregSub, SregMult, RegDiv, RegInc, RegDec, RegNegate
--|-----------------------------------------------------------------------------
    PROCEDURE SregMult (SIGNAL result         : OUT STD_ULOGIC_VECTOR;
                        SIGNAL overflow       : OUT STD_ULOGIC;
                        CONSTANT multiplicand : IN STD_ULOGIC_VECTOR;
                        CONSTANT multiplier   : IN STD_ULOGIC_VECTOR;
                        CONSTANT SrcRegMode   : IN regmode_type 
                  -- synopsys synthesis_off
                                                       := DefaultRegMode 
                   -- synopsys synthesis_on
                      ) IS
        VARIABLE reslt       : STD_LOGIC_VECTOR ( result'length  - 1  DOWNTO 0 );
        VARIABLE overflo     : STD_ULOGIC;
	VARIABLE a_copy      : STD_LOGIC_VECTOR (multiplicand'length-1 downto 0 );
	VARIABLE b_copy      : STD_LOGIC_VECTOR (multiplier'length-1 downto 0 );
     BEGIN 
	a_copy := To_StdLogicVector(multiplicand);
	b_copy := To_StdLogicVector(multiplier);

	RegMult(reslt, overflo, a_copy, b_copy, SrcRegMode);

        result   <= To_StdULogicVector(reslt)
                     -- synopsys synthesis_off
             				after DefaultRegDelay
                     -- synopsys synthesis_on
                                                             ;
        overflow <= overflo
                     -- synopsys synthesis_off
             				after DefaultRegDelay
                     -- synopsys synthesis_on
                                                             ;
        RETURN;
    END SregMult;
--+-----------------------------------------------------------------------------
--|     Function Name  : SregMult
--|
--|     Overloading    : None
--|
--|     Purpose        : Multiplication of BIT_VECTORS.
--|
--|     Parameters     :
--|                      result       - output BIT_VECTOR, the computed product
--|                      overflow     - output BIT, overflow condition
--|                      multiplicand - input BIT_VECTOR,
--|                      multiplier   -  input BIT_VECTOR,
--|                      SrcRegMode   - input  regmode_type, indicating the format 
--|                                     of the input BIT_VECTOR.   Default is 
--|                                     DefaultRegMode which is set to TwosComp.
--|     NOTE           :
--|                      The inputs may be of any length and may be of differing
--|                      lengths.
--|
--|    Algorithm       : The multiplication is carried out as follows:
--|
--|                      1) Determine sign of result based on sign of 
--|                         multiploicand and sign  of multiplier.
--|
--|                      2) Convert the multiplicand amd multiplier to Unsigned 
--|                         representation.
--|                      
--|                      3) Perform multiplication based on add and shift algorithm.
--|
--|                      4) Convert the result to the SrcRegMode with appropropriate sign
--|
--|     Result         :
--|                     A  temporary result is computed with length N+M (where
--|                      N,M are the lengths of the multiplicand and multiplier).
--|                      This computed value is extended or truncated to match
--|                      the width of 'result'. If truncated, the low order bits
--|                      are returned.
--|
--|                      The parameter 'overflow' is set to '1' if the product of the
--|                      of the two inputs too large to fit in the parameter result.
--|     Use            :
--|                      SIGNAL x, y, prod : BIT_VECTOR ( 15 DOWNTO 0);
--|                      SIGNAL ovfl : BIT;
--|
--|                      SregMult ( prod, ovfl, x, y, TwosComp );
--|
--|     See Also       : RegAdd, SregSub, SregMult, RegDiv, RegInc, RegDec, RegNegate
--|-----------------------------------------------------------------------------
    PROCEDURE SregMult (SIGNAL result         : OUT BIT_VECTOR;
                        SIGNAL overflow       : OUT BIT;
                        CONSTANT multiplicand : IN BIT_VECTOR;
                        CONSTANT multiplier   : IN BIT_VECTOR;
                        CONSTANT SrcRegMode   : IN regmode_type 
                  -- synopsys synthesis_off
                                                       := DefaultRegMode 
                   -- synopsys synthesis_on
                      ) IS

        VARIABLE reslt       : STD_LOGIC_VECTOR ( result'length  - 1  DOWNTO 0 );
        VARIABLE overflo     : STD_ULOGIC;
	VARIABLE a_copy      : STD_LOGIC_VECTOR (multiplicand'length-1 downto 0 );
	VARIABLE b_copy      : STD_LOGIC_VECTOR (multiplier'length-1 downto 0 );
     BEGIN 
	a_copy := To_StdLogicVector(multiplicand);
	b_copy := To_StdLogicVector(multiplier);

        RegMult(reslt, overflo, a_copy, b_copy, SrcRegMode);
     
        result   <= To_BitVector(reslt) 
                     -- synopsys synthesis_off
             				after DefaultRegDelay
                     -- synopsys synthesis_on
                                                             ;
        overflow <= To_Bit(overflo) 
                     -- synopsys synthesis_off
             				after DefaultRegDelay
                     -- synopsys synthesis_on
                                                             ;
        RETURN;
    END SregMult;
--+-----------------------------------------------------------------------------
--|     Function Name  : SregDiv
--|
--|     Overloading    : None
--|
--|     Purpose        : Division of BIT_VECTORS. (Result = dividend / divisor)
--|
--|     Parameters     :
--|                      result     - output BIT_VECTOR,
--|                      remainder  - output BIT_VECTOR,
--|                      ZeroDivide - output BIT,
--|                                   set to '1'  when divide by zero occurred
--|                                          '0'  divide by zero did not occur
--|                      dividend   - input  BIT_VECTOR,
--|                      divisor    - input  BIT_VECTOR,
--|                      SrcRegMode - input  regmode_type, indicating the format of
--|                                the input BIT_VECTOR.   Default is TwosComp.
--|     NOTE           :
--|                      The inputs may be of any length and may be of differing
--|                      lengths.
--|
--|                      For synthesis purposes result and remainder values are 
--|                      computed with  same length as the dividend. 
--|
--|                      The remainder has the same sign as the dividend.
--|     Use            :
--|                      SIGNAL x, y, res, rem : BIT_VECTOR ( 15 DOWNTO 0);
--|                      SIGNAL Zflag : BIT;
--|
--|                      SregDiv ( res, rem,Zflag, x, y, TwosComp );
--|
--|     See Also       : SregAdd, SregSub, SregMult, SregMod, SregRem
--|-----------------------------------------------------------------------------
    PROCEDURE SregDiv ( SIGNAL result       : OUT BIT_VECTOR;
                        SIGNAL remainder    : OUT BIT_VECTOR;
                        SIGNAL ZeroDivide   : OUT BIT;
                        CONSTANT dividend   :  IN BIT_VECTOR;
                        CONSTANT divisor    :  IN BIT_VECTOR;
                        CONSTANT SrcRegMode    :  IN regmode_type 
                  -- synopsys synthesis_off
                                                       := DefaultRegMode 
                   -- synopsys synthesis_on
                      ) IS
        VARIABLE remaind : STD_LOGIC_VECTOR(remainder'LENGTH - 1 DOWNTO 0);
        VARIABLE reslt   : STD_LOGIC_VECTOR(result'LENGTH - 1 DOWNTO 0);
        VARIABLE Zdiv    : STD_ULOGIC;
	VARIABLE a_copy  : STD_LOGIC_VECTOR (dividend'length-1 downto 0 );
	VARIABLE b_copy  : STD_LOGIC_VECTOR (divisor'length-1 downto 0 );
     BEGIN 
	a_copy := To_StdLogicVector(dividend);
	b_copy := To_StdLogicVector(divisor);

	RegDiv(reslt, remaind, Zdiv, a_copy, b_copy, SrcRegMode);

        result     <= To_BitVector(reslt) 
                     -- synopsys synthesis_off
             				after DefaultRegDelay
                     -- synopsys synthesis_on
                                                             ;
        remainder  <= To_BitVector(remaind)
                     -- synopsys synthesis_off
             				after DefaultRegDelay
                     -- synopsys synthesis_on
                                                             ;
        ZeroDivide <= To_Bit(Zdiv) 
                     -- synopsys synthesis_off
             				after DefaultRegDelay
                     -- synopsys synthesis_on
                                                             ;
        RETURN;
    END SRegDiv;
    -------------------------------------------------------------------------------
    --     Function Name  : SregDiv
    --
    --     Overloading    : None
    --    
    --     Purpose        : Division of std_logic_vectors.(Result = dividend/divisor)
    --     
    --     Parameters     : 
    --                      result     - output std_logic_vector, 
    --                      remainder  - output std_logic_vector,
    --                      ZeroDivide - output std_ulogic,
    --                                   set to '1' when  divide by zero occurred
    --                                          '0'  divide by zero did not occur  
    --                      dividend   - input  std_logic_vector, 
    --                      divisor    - input  std_logic_vector, 
    --                      SrcRegMode - input  regmode_type, indicating the format 
    --                                   of  the input std_logic_vector.   
    --                                   Default is TwosComp.
    --     NOTE           : 
    --                      The inputs may be of any length and may be of differing 
    --                      lengths. 
    --
    --                      For synthesis purposes result and remainder values are 
    --                      computed with  same length as the dividend. 
    --                      The remainder has the same sign as the dividend.
    --     Use            : 
    --                      SIGNAL x, y, res, rem : std_logic_vector ( 15 DOWNTO 0);
    --                      SIGNAL Zflag : std_ulogic;
    --
    --                      SregDiv ( res, rem, Zflag, x, y, TwosComp );
    --     
    --     See Also       : SregAdd, SregSub, SregMult, SregMod, SregRem
    -------------------------------------------------------------------------------
    PROCEDURE SregDiv ( SIGNAL result       : OUT std_logic_vector;
                        SIGNAL remainder    : OUT std_logic_vector;
                        SIGNAL ZeroDivide   : OUT std_ulogic;  
                        CONSTANT dividend   :  IN std_logic_vector;
                        CONSTANT divisor    :  IN std_logic_vector;
                        CONSTANT SrcRegMode :  IN regmode_type
                  -- synopsys synthesis_off
                                                       := DefaultRegMode 
                  -- synopsys synthesis_on
                      ) IS

      VARIABLE remaind : STD_LOGIC_VECTOR(remainder'LENGTH - 1 DOWNTO 0);
      VARIABLE reslt   : STD_LOGIC_VECTOR(result'LENGTH - 1 DOWNTO 0);
      VARIABLE Zdiv    : STD_ULOGIC;

     BEGIN 
	RegDiv(reslt, remaind, Zdiv, dividend, divisor, SrcRegMode);

        result     <= reslt
                     -- synopsys synthesis_off
             				after DefaultRegDelay
                     -- synopsys synthesis_on
                                                             ;
        remainder  <= remaind 
                     -- synopsys synthesis_off
             				after DefaultRegDelay
                     -- synopsys synthesis_on
                                                             ;
        ZeroDivide <= Zdiv 
                     -- synopsys synthesis_off
             				after DefaultRegDelay
                     -- synopsys synthesis_on
                                                             ;
        RETURN;
   END SRegDiv;
    -------------------------------------------------------------------------------
    --     Function Name  : SregDiv
    --
    --     Overloading    : None
    --    
    --     Purpose        : Division of std_ulogic_vectors.(Result = dividend/divisor)
    --     
    --     Parameters     : 
    --                      result     - output std_ulogic_vector, 
    --                      remainder  - output std_ulogic_vector,
    --                      ZeroDivide - output std_ulogic,
    --                                   set to '1' when  divide by zero occurred
    --                                          '0'  divide by zero did not occur  
    --                      dividend   - input  std_ulogic_vector, 
    --                      divisor    - input  std_ulogic_vector, 
    --                      SrcRegMode - input  regmode_type, indicating the format 
    --                                   of  the input std_ulogic_vector.   
    --                                   Default is TwosComp.
    --     NOTE           : 
    --                      The inputs may be of any length and may be of differing 
    --                      lengths. 
    --
    --                      For synthesis purposes result and remainder values are 
    --                      computed with  same length as the dividend. 
    --                      The remainder has the same sign as the dividend.
    --     Use            : 
    --                      SIGNAL x, y, res, rem : std_ulogic_vector ( 15 DOWNTO 0);
    --                      SIGNAL Zflag : std_ulogic;
    --
    --                      SregDiv ( res, rem, Zflag, x, y, TwosComp );
    --     
    --     See Also       : SregAdd, SregSub, SregMult, SregMod, SregRem
    -------------------------------------------------------------------------------
    PROCEDURE SregDiv ( SIGNAL result       : OUT std_ulogic_vector;
                        SIGNAL remainder    : OUT std_ulogic_vector;
                        SIGNAL ZeroDivide   : OUT std_ulogic;  
                        CONSTANT dividend   :  IN std_ulogic_vector;
                        CONSTANT divisor    :  IN std_ulogic_vector;
                        CONSTANT SrcRegMode :  IN regmode_type
                  -- synopsys synthesis_off
                                                       := DefaultRegMode 
                  -- synopsys synthesis_on
                      ) IS
	VARIABLE remaind : STD_LOGIC_VECTOR(remainder'LENGTH - 1 DOWNTO 0);
	VARIABLE reslt   : STD_LOGIC_VECTOR(result'LENGTH - 1 DOWNTO 0);
	VARIABLE Zdiv    : STD_ULOGIC;
	VARIABLE a_copy  : STD_LOGIC_VECTOR (dividend'length-1 downto 0 );
	VARIABLE b_copy  : STD_LOGIC_VECTOR (divisor'length-1 downto 0 );
     BEGIN 
	a_copy := To_StdLogicVector(dividend);
	b_copy := To_StdLogicVector(divisor);

	RegDiv(reslt, remaind, Zdiv, a_copy, b_copy, SrcRegMode);

        result     <= To_StdULogicVector(reslt) 
                     -- synopsys synthesis_off
             				after DefaultRegDelay
                     -- synopsys synthesis_on
                                                             ;
        remainder  <= To_StdULogicVector(remaind)
                     -- synopsys synthesis_off
             				after DefaultRegDelay
                     -- synopsys synthesis_on
                                                             ;
        ZeroDivide <= Zdiv 
                     -- synopsys synthesis_off
             				after DefaultRegDelay
                     -- synopsys synthesis_on
                                                             ;
        RETURN;
   END SRegDiv;
--+-----------------------------------------------------------------------------
--|     Function Name  : SregMod
--| 1.5.17  
--|     Overloading    : None
--| 
--|     Purpose        : Modulus operation of  BIT_VECTORS.
--| 
--|     Parameters     :
--|                      result     - output BIT_VECTOR,
--|                      ZeroDivide - output BIT,
--|                                   set to '1'  when divide by zero occurred
--|                                          '0'  divide by zero did not occur
--|                      dividend   - input  BIT_VECTOR,
--|                      modulus    - input  BIT_VECTOR,
--|                      SrcRegMode - input  regmode_type, indicating the format of
--|                                the input BIT_VECTOR.   Default is TwosComp.
--|     NOTE           :
--|                      The inputs may be of any length and may be of differing
--|                      lengths.
--|
--|                      For synthesis purposes quotient and modulus values are 
--|                      computed with  same length as the dividend. 
--|
--|                      The mod has the same sign as the modulus operator.
--|     Use            :
--|                      SIGNAL x, y, res : BIT_VECTOR ( 15 DOWNTO 0);
--|                      SIGNAL zflag     : BIT;
--|
--|                      SregMod ( res,zflag, x, y, TwosComp );
--|
--|     See Also       : SregAdd, SregSub, SregMult, SregDiv
--|-----------------------------------------------------------------------------
    PROCEDURE SregMod  ( SIGNAL result     : OUT BIT_VECTOR;
                        SIGNAL ZeroDivide : OUT BIT;
                        CONSTANT dividend   : IN BIT_VECTOR;
                        CONSTANT modulus    : IN BIT_VECTOR;
                        CONSTANT SrcRegMode : IN regmode_type
                     -- synopsys synthesis_off
						      := DefaultRegMode 
                     -- synopsys synthesis_on
                      ) IS
	VARIABLE reslt   : STD_LOGIC_VECTOR(result'LENGTH - 1 DOWNTO 0);
	VARIABLE Zdiv    : STD_ULOGIC;
	VARIABLE d_copy  : STD_LOGIC_VECTOR (dividend'length-1 downto 0 );
	VARIABLE m_copy  : STD_LOGIC_VECTOR (modulus'length-1 downto 0 );
     BEGIN 
	d_copy := To_StdLogicVector(dividend);
	m_copy := To_StdLogicVector(modulus);

	RegMod(reslt, Zdiv, d_copy, m_copy, SrcRegMode);

        result     <= To_BitVector(reslt)
	-- synopsys synthesis_off        
                                               after DefaultRegDelay
	-- synopsys synthesis_on        
                                                         ;	
        ZeroDivide <= To_Bit(Zdiv)
	-- synopsys synthesis_off        
                                               after DefaultRegDelay
	-- synopsys synthesis_on        
                                                         ;	
        RETURN;
    END SregMod;
--+-----------------------------------------------------------------------------
--|     Function Name  : SregMod
--| 1.5.17  
--|     Overloading    : None
--| 
--|     Purpose        : Modulus operation of  STD_LOGIC_VECTORS.
--| 
--|     Parameters     :
--|                      result     - output STD_LOGIC_VECTOR,
--|                      ZeroDivide - output STD_ULOGIC,
--|                                   set to '1'  when divide by zero occurred
--|                                          '0'  divide by zero did not occur
--|                      dividend   - input  STD_LOGIC_VECTOR,
--|                      modulus    - input  STD_LOGIC_VECTOR,
--|                      SrcRegMode - input  regmode_type, indicating the format of
--|                                the input STD_LOGIC_VECTOR.   Default is TwosComp.
--|     NOTE           :
--|                      The inputs may be of any length and may be of differing
--|                      lengths.
--|
--|                      For synthesis purposes quotient and modulus values are 
--|                      computed with  same length as the dividend. 
--|
--|                      The mod has the same sign as the modulus operator.
--|     Use            :
--|                      SIGNAL x, y, res : STD_LOGIC_VECTOR ( 15 DOWNTO 0);
--|                      SIGNAL zflag     : STD_ULOGIC;
--|
--|                      SregMod ( res,zflag, x, y, TwosComp );
--|
--|     See Also       : SregAdd, SregSub, SregMult, SregDiv
--|-----------------------------------------------------------------------------
    PROCEDURE SregMod  ( SIGNAL result     : OUT STD_LOGIC_VECTOR;
                        SIGNAL ZeroDivide : OUT STD_ULOGIC;
                        CONSTANT dividend   : IN STD_LOGIC_VECTOR;
                        CONSTANT modulus    : IN STD_LOGIC_VECTOR;
                        CONSTANT SrcRegMode : IN regmode_type
                     -- synopsys synthesis_off
						      := DefaultRegMode 
                     -- synopsys synthesis_on
                      ) IS
	VARIABLE reslt   : STD_LOGIC_VECTOR(result'LENGTH - 1 DOWNTO 0);
	VARIABLE Zdiv    : STD_ULOGIC;
     BEGIN 
	RegMod(reslt, Zdiv, dividend, modulus, SrcRegMode);

        result     <= reslt
	-- synopsys synthesis_off        
                                               after DefaultRegDelay
	-- synopsys synthesis_on        
                                                         ;	
        ZeroDivide <= Zdiv 
	-- synopsys synthesis_off        
                                               after DefaultRegDelay
	-- synopsys synthesis_on        
                                                         ;	
        RETURN;
    END SregMod;
--+-----------------------------------------------------------------------------
--|     Function Name  : SregMod
--| 1.5.17  
--|     Overloading    : None
--| 
--|     Purpose        : Modulus operation of  STD_ULOGIC_VECTORS.
--| 
--|     Parameters     :
--|                      result     - output STD_ULOGIC_VECTOR,
--|                      ZeroDivide - output STD_ULOGIC,
--|                                   set to '1'  when divide by zero occurred
--|                                          '0'  divide by zero did not occur
--|                      dividend   - input  STD_ULOGIC_VECTOR,
--|                      modulus    - input  STD_ULOGIC_VECTOR,
--|                      SrcRegMode - input  regmode_type, indicating the format of
--|                                the input STD_ULOGIC_VECTOR.   Default is TwosComp.
--|     NOTE           :
--|                      The inputs may be of any length and may be of differing
--|                      lengths.
--|
--|                      For synthesis purposes quotient and modulus values are 
--|                      computed with  same length as the dividend. 
--|
--|                      The mod has the same sign as the modulus operator.
--|     Use            :
--|                      SIGNAL x, y, res : STD_ULOGIC_VECTOR ( 15 DOWNTO 0);
--|                      SIGNAL zflag     : STD_ULOGIC;
--|
--|                      SregMod ( res,zflag, x, y, TwosComp );
--|
--|     See Also       : SregAdd, SregSub, SregMult, SregDiv 
--|-----------------------------------------------------------------------------
    PROCEDURE SregMod  ( SIGNAL result     : OUT STD_ULOGIC_VECTOR;
                        SIGNAL ZeroDivide : OUT STD_ULOGIC;
                        CONSTANT dividend   : IN STD_ULOGIC_VECTOR;
                        CONSTANT modulus    : IN STD_ULOGIC_VECTOR;
                        CONSTANT SrcRegMode : IN regmode_type
                     -- synopsys synthesis_off
						      := DefaultRegMode 
                     -- synopsys synthesis_on
                      ) IS
	VARIABLE reslt   : STD_LOGIC_VECTOR(result'LENGTH - 1 DOWNTO 0);
	VARIABLE Zdiv    : STD_ULOGIC;
	VARIABLE d_copy  : STD_LOGIC_VECTOR (dividend'length-1 downto 0 );
	VARIABLE m_copy  : STD_LOGIC_VECTOR (modulus'length-1 downto 0 );
     BEGIN 
	d_copy := To_StdLogicVector(dividend);
	m_copy := To_StdLogicVector(modulus);

	RegMod(reslt, Zdiv, d_copy, m_copy, SrcRegMode);

        result     <= To_StdULogicVector(reslt) 
	-- synopsys synthesis_off        
                                               after DefaultRegDelay
	-- synopsys synthesis_on        
                                                         ;	
        ZeroDivide <= Zdiv 
	-- synopsys synthesis_off        
                                               after DefaultRegDelay
	-- synopsys synthesis_on        
                                                         ;	
        RETURN;
    END SregMod;
--+-----------------------------------------------------------------------------
--|     Function Name  : SregRem
--| 1.5.25
--|     Overloading    : None
--|
--|     Purpose        : Remainder operation of  BIT_VECTORS.
--|
--|     Parameters     :
--|                      result     - output BIT_VECTOR,
--|                      ZeroDivide - output BIT,
--|                                   set to '1'  when divide by zero occurred
--|                                          '0'  divide by zero did not occur
--|                      dividend   - input  BIT_VECTOR,
--|                      divisor    - input  BIT_VECTOR,
--|                      SrcRegMode - input  regmode_type, indicating the format of
--|                                the input BIT_VECTOR.   Default is TwosComp.
--|     NOTE           :
--|                      The inputs may be of any length and may be of differing
--|                      lengths.
--|
--|                      For synthesis purposes quotient and remainder values are 
--|                      computed with  same length as the dividend. 
--|
--|                      The remainder has the same sign as the dividend.
--|     Use            :
--|                      VARIABLE x, y, res : BIT_VECTOR ( 15 DOWNTO 0);
--|                      VARIABLE zflag     : BIT;
--|
--|                      SregRem ( res, zflag, x, y, TwosComp );
--|
--|     See Also       : SeegAdd, SregSub, SregMult, SregDiv
--|-----------------------------------------------------------------------------
    PROCEDURE SregRem ( SIGNAL result       : OUT BIT_VECTOR;
                        SIGNAL ZeroDivide   : OUT BIT;
                        CONSTANT dividend   :  IN BIT_VECTOR;
                        CONSTANT divisor    :  IN BIT_VECTOR;
                        CONSTANT SrcRegMode :  IN regmode_type
                     -- synopsys synthesis_off
						      := DefaultRegMode 
                     -- synopsys synthesis_on
                      ) IS

        VARIABLE reslt   : STD_LOGIC_VECTOR(result'LENGTH - 1 DOWNTO 0);
        VARIABLE Zdiv    : STD_ULOGIC;
	VARIABLE a_copy  : STD_LOGIC_VECTOR (dividend'length-1 downto 0 );
	VARIABLE b_copy  : STD_LOGIC_VECTOR (divisor'length-1 downto 0 );
     BEGIN 
	a_copy := To_StdLogicVector(dividend);
	b_copy := To_StdLogicVector(divisor);

	RegRem(reslt, Zdiv, a_copy, b_copy, SrcRegMode);

        result     <= To_BitVector(reslt)
	-- synopsys synthesis_off        
                                               after DefaultRegDelay
	-- synopsys synthesis_on        
                                                         ;	
        ZeroDivide <= To_Bit(Zdiv)
	-- synopsys synthesis_off        
                                               after DefaultRegDelay
	-- synopsys synthesis_on        
                                                         ;	
        RETURN;
    END SregRem;
--+-----------------------------------------------------------------------------
--|     Function Name  : SregRem
--| 1.5.25
--|     Overloading    : None
--|
--|     Purpose        : Remainder operation of  STD_LOGIC_VECTORS.
--|
--|     Parameters     :
--|                      result     - output STD_LOGIC_VECTOR,
--|                      ZeroDivide - output STD_ULOGIC,
--|                                   set to '1'  when divide by zero occurred
--|                                          '0'  divide by zero did not occur
--|                      dividend   - input  STD_LOGIC_VECTOR,
--|                      divisor    - input  STD_LOGIC_VECTOR,
--|                      SrcRegMode - input  regmode_type, indicating the format of
--|                                the input STD_LOGIC_VECTOR.   Default is TwosComp.
--|     NOTE           :
--|                      The inputs may be of any length and may be of differing
--|                      lengths.
--|
--|                      For synthesis purposes quotient and remainder values are 
--|                      computed with  same length as the dividend. 
--|
--|                      The remainder has the same sign as the dividend.
--|     Use            :
--|                      VARIABLE x, y, res : STD_LOGIC_VECTOR ( 15 DOWNTO 0);
--|                      VARIABLE zflag     : STD_ULOGIC;
--|
--|                      SregRem ( res, zflag, x, y, TwosComp );
--|
--|     See Also       : SeegAdd, SregSub, SregMult, SregDiv
--|-----------------------------------------------------------------------------
    PROCEDURE SregRem ( SIGNAL result       : OUT STD_LOGIC_VECTOR;
                        SIGNAL ZeroDivide   : OUT STD_ULOGIC;
                        CONSTANT dividend   :  IN STD_LOGIC_VECTOR;
                        CONSTANT divisor    :  IN STD_LOGIC_VECTOR;
                        CONSTANT SrcRegMode :  IN regmode_type
                     -- synopsys synthesis_off
						      := DefaultRegMode 
                     -- synopsys synthesis_on
                      ) IS
      VARIABLE reslt   : STD_LOGIC_VECTOR(result'LENGTH - 1 DOWNTO 0);
      VARIABLE Zdiv    : STD_ULOGIC;

     BEGIN 
	RegRem(reslt,  Zdiv, dividend, divisor, SrcRegMode);

        result     <= reslt
	-- synopsys synthesis_off        
                                               after DefaultRegDelay
	-- synopsys synthesis_on        
                                                         ;	
        ZeroDivide <= Zdiv 
	-- synopsys synthesis_off        
                                               after DefaultRegDelay
	-- synopsys synthesis_on        
                                                         ;	
        RETURN;
    END SregRem;
--+-----------------------------------------------------------------------------
--|     Function Name  : SregRem
--| 1.5.25
--|     Overloading    : None
--|
--|     Purpose        : Remainder operation of  STD_ULOGIC_VECTORS.
--|
--|     Parameters     :
--|                      result     - output STD_ULOGIC_VECTOR,
--|                      ZeroDivide - output STD_ULOGIC,
--|                                   set to '1'  when divide by zero occurred
--|                                          '0'  divide by zero did not occur
--|                      dividend   - input  STD_ULOGIC_VECTOR,
--|                      divisor    - input  STD_ULOGIC_VECTOR,
--|                      SrcRegMode - input  regmode_type, indicating the format of
--|                                the input STD_ULOGIC_VECTOR.   Default is TwosComp.
--|     NOTE           :
--|                      The inputs may be of any length and may be of differing
--|                      lengths.
--|
--|                      For synthesis purposes quotient and remainder values are 
--|                      computed with  same length as the dividend. 
--|
--|                      The remainder has the same sign as the dividend.
--|     Use            :
--|                      VARIABLE x, y, res : STD_ULOGIC_VECTOR ( 15 DOWNTO 0);
--|                      VARIABLE zflag     : STD_ULOGIC;
--|
--|                      SregRem ( res, zflag, x, y, TwosComp );
--|
--|     See Also       : SeegAdd, SregSub, SregMult, SregDiv
--|-----------------------------------------------------------------------------
    PROCEDURE SregRem ( SIGNAL result       : OUT STD_ULOGIC_VECTOR;
                        SIGNAL ZeroDivide   : OUT STD_ULOGIC;
                        CONSTANT dividend   :  IN STD_ULOGIC_VECTOR;
                        CONSTANT divisor    :  IN STD_ULOGIC_VECTOR;
                        CONSTANT SrcRegMode :  IN regmode_type
                     -- synopsys synthesis_off
						      := DefaultRegMode 
                     -- synopsys synthesis_on
                      ) IS
        VARIABLE reslt   : STD_LOGIC_VECTOR(result'LENGTH - 1 DOWNTO 0);
        VARIABLE Zdiv    : STD_ULOGIC;
	VARIABLE a_copy  : STD_LOGIC_VECTOR (dividend'length-1 downto 0 );
	VARIABLE b_copy  : STD_LOGIC_VECTOR (divisor'length-1 downto 0 );
     BEGIN 
	a_copy := To_StdLogicVector(dividend);
	b_copy := To_StdLogicVector(divisor);

	RegRem(reslt, Zdiv, a_copy, b_copy, SrcRegMode);

        result     <= To_StdULogicVector(reslt) 
	-- synopsys synthesis_off        
                                               after DefaultRegDelay
	-- synopsys synthesis_on        
                                                         ;	
        ZeroDivide <= Zdiv  
	-- synopsys synthesis_off        
                              after DefaultRegDelay
	-- synopsys synthesis_on        
                                        ;	
        RETURN;
    END SregRem;
--+-----------------------------------------------------------------------------
--|     Function Name  : SregShift
--| 
--|     Overloading    : None
--|
--|     Purpose        : Bidirectional logical shift operator for logic vector.
--|
--|     Parameters     :
--|                      SrcReg      - input  bit_vector, vector to be shifted
--|                      DstReg      - ouput, bit_vector, shifted result
--|                      ShiftO      - output, bit, holds the 
--|                                            last bit shifted out 
--|                                          of register
--|                      direction   - input, bit
--|                                         '0'  means right shift
--|                                         '1' | 'X'  means left shift, 
--|                                          default is left shift
--|                      FillVal     - input, bit, value to fill register with. 
--|                                          default is '0'
--|                      Nbits       - input , NATURAL, number of positions to shift
--|                                          default is 1.
--|
--|     Result         : Shifted bit_vector
--|
--|     NOTE           : Defaults not allowed for synthesis.
--|
--|     Use            :
--|                      SIGNAL acc   : bit_vector ( 15 DOWNTO 0);
--|                      SIGNAL carry : bit;
--|
--|                      SregShift ( acc, acc, carry, '1', '0',3 );
--|-----------------------------------------------------------------------------
   PROCEDURE SregShift ( CONSTANT SrcReg    : IN bit_vector;
                         SIGNAL DstReg    : INOUT bit_vector;
                         SIGNAL ShiftO    : OUT bit; 
                         CONSTANT direction : IN bit
                     -- synopsys synthesis_off
						      := '1'
                     -- synopsys synthesis_on
                                                            ;
                         CONSTANT FillVal   : IN bit  
                     -- synopsys synthesis_off
						      := '0'
                     -- synopsys synthesis_on
                                                            ;
                         CONSTANT Nbits     : IN Natural
                     -- synopsys synthesis_off
						       := 1 
                     -- synopsys synthesis_on
                      ) IS 
	CONSTANT dlen      : INTEGER := DstReg'LENGTH;
        VARIABLE r         : BIT_VECTOR (SrcReg'LENGTH - 1 DOWNTO 0);
        VARIABLE src_copy  : BIT_VECTOR (SrcReg'LENGTH - 1 DOWNTO 0 );
        VARIABLE dst_copy  : BIT_VECTOR (DstReg'LENGTH - 1 DOWNTO 0 );
        VARIABLE Shiftout  : BIT;
   BEGIN
       src_copy   := SrcReg;
       dst_copy   := DstReg;
 -- synopsys translate_off    
    --  Null range Check
    --  if input vector is of zero length
       IF ( SrcReg'LENGTH = 0) THEN
           ASSERT false
           REPORT " SregShift --- input bit_vector   is null  "
           SEVERITY ERROR;
           dst_copy := (OTHERS => FillVal);
           DstReg    <= dst_copy after DefaultRegDelay;
           ShiftO <= '0' after DefaultRegDelay;
           Return;
       ELSIF (DstReg'LENGTH = 0) THEN
           ASSERT false
           REPORT " SregShift --- output vector is  null  "
           SEVERITY ERROR;
         -- set shift out bit at least
           IF ( direction /= '0') THEN
               ShiftO <= src_copy(SrcReg'LENGTH - Nbits) after DefaultRegDelay;
           ELSE 
               ShiftO <= src_copy(Nbits - 1) after DefaultRegDelay;
           END IF;
           RETURN;
      END IF;
-- synopsys translate_on
    -- None of the registers is null, perform shift operation
      IF (direction /= '0') THEN                                 --  left shift
           RegShift_Left(src_copy, r, Shiftout, FillVal, Nbits);
      ELSE                                                       -- right shift
           RegShift_Right(src_copy, r, Shiftout, FillVal, Nbits);
      END IF;
      -- determine length of the result
      IF (dlen <= SrcReg'LENGTH) THEN
		for i IN dlen - 1 downto 0 Loop
			dst_copy(i) := r(i);
                end loop;
      ELSE
		for i IN SrcReg'LENGTH - 1 downto 0 Loop
			dst_copy(i) := r(i);
                end loop;
      END IF;
      DstReg <= dst_copy 
-- synopsys translate_off     
			after DefaultRegDelay
-- synopsys translate_on
       						;
      ShiftO <= Shiftout
-- synopsys translate_off     
			after DefaultRegDelay
-- synopsys translate_on
       						;
      RETURN;
   END SregShift;
--+-----------------------------------------------------------------------------
--|     Function Name  : SregShift
--| 
--|     Overloading    : None
--|
--|     Purpose        : Bidirectional logical shift operator for logic vector.
--|
--|     Parameters     :
--|                      SrcReg      - input  std_logic_vector, vector to be shifted
--|                      DstReg      - ouput, std_logic_vector, shifted result
--|                      ShiftO      - output, std_ulogic, holds the 
--|                                            last bit shifted out 
--|                                          of register
--|                      direction   - input, Std_ulogic
--|                                         '0'  means right shift
--|                                         '1' | 'X'  means left shift, 
--|                                          default is left shift
--|                      FillVal     - input, Std_ulogic, value to fill register with. 
--|                                          default is '0'
--|                      Nbits       - input , NATURAL, number of positions to shift
--|                                          default is 1.
--|
--|     Result         : Shifted std_logic_vector
--|
--|     NOTE           : Defaults not allowed for synthesis.
--|
--|     Use            :
--|                      SIGNAL acc   : std_logic_vector ( 15 DOWNTO 0);
--|                      SIGNAL carry : std_ulogic;
--|
--|                      SregShift ( acc, acc, carry, '1', '0',3 );
--|-----------------------------------------------------------------------------
   PROCEDURE SregShift ( CONSTANT SrcReg    : IN std_logic_vector;
                         SIGNAL DstReg    : INOUT std_logic_vector;
                         SIGNAL ShiftO    : OUT std_ulogic; 
                         CONSTANT direction : IN std_ulogic
                     -- synopsys synthesis_off
						      := '1'
                     -- synopsys synthesis_on
                                                            ;
                         CONSTANT FillVal   : IN std_ulogic  
                     -- synopsys synthesis_off
						      := '0'
                     -- synopsys synthesis_on
                                                            ;
                         CONSTANT Nbits     : IN Natural
                     -- synopsys synthesis_off
						       := 1 
                     -- synopsys synthesis_on
                      ) IS 
	CONSTANT dlen      : INTEGER := DstReg'LENGTH;
        VARIABLE r         : STD_LOGIC_VECTOR (SrcReg'LENGTH - 1 DOWNTO 0);
        VARIABLE src_copy  : STD_LOGIC_VECTOR (SrcReg'LENGTH - 1 DOWNTO 0 );
        VARIABLE dst_copy  : STD_LOGIC_VECTOR (DstReg'LENGTH - 1 DOWNTO 0 );
        VARIABLE Shiftout  : STD_ULOGIC;
   BEGIN
       src_copy   := SrcReg;
       dst_copy   := DstReg;
 -- synopsys translate_off    
    --  Null range Check
    --  if input vector is of zero length
       IF ( SrcReg'LENGTH = 0) THEN
           ASSERT false
           REPORT " SregShift --- input bit_vector   is null  "
           SEVERITY ERROR;
           dst_copy := (OTHERS => FillVal);
           DstReg    <= dst_copy after DefaultRegDelay;
           ShiftO <= '0' after DefaultRegDelay;
           Return;
       ELSIF (DstReg'LENGTH = 0) THEN
           ASSERT false
           REPORT " SregShift --- output vector is  null  "
           SEVERITY ERROR;
         -- set shift out bit at least
           IF ( direction /= '0') THEN
               ShiftO <= src_copy(SrcReg'LENGTH - Nbits) after DefaultRegDelay;
           ELSE 
               ShiftO <= src_copy(Nbits - 1) after DefaultRegDelay;
           END IF;
           RETURN;
      END IF;
-- synopsys translate_on
    -- None of the registers is null, perform shift operation
      IF (direction /= '0') THEN                                 --  left shift
           RegShift_Left(src_copy, r, Shiftout, FillVal, Nbits);
      ELSE                                                       -- right shift
           RegShift_Right(src_copy, r, Shiftout, FillVal, Nbits);
      END IF;
      -- determine length of the result
      IF (dlen <= SrcReg'LENGTH) THEN
		for i IN dlen - 1 downto 0 Loop
			dst_copy(i) := r(i);
                end loop;
      ELSE
		for i IN SrcReg'LENGTH - 1 downto 0 Loop
			dst_copy(i) := r(i);
                end loop;
      END IF;
      DstReg <= dst_copy 
		-- synopsys translate_off     
			after DefaultRegDelay
		-- synopsys translate_on
       						;
      ShiftO <= Shiftout
		-- synopsys translate_off     
			after DefaultRegDelay
		-- synopsys translate_on
       						;
      RETURN;
   END SregShift;
--+-----------------------------------------------------------------------------
--|     Function Name  : SregShift
--| 
--|     Overloading    : None
--|
--|     Purpose        : Bidirectional logical shift operator for logic vector.
--|
--|     Parameters     :
--|                      SrcReg      - input  std_ulogic_vector, vector to be shifted
--|                      DstReg      - ouput, std_ulogic_vector, shifted result
--|                      ShiftO      - output, std_ulogic, holds the 
--|                                            last bit shifted out 
--|                                          of register
--|                      direction   - input, Std_ulogic
--|                                         '0'  means right shift
--|                                         '1' | 'X'  means left shift, 
--|                                          default is left shift
--|                      FillVal     - input, Std_ulogic, value to fill register with. 
--|                                          default is '0'
--|                      Nbits       - input , NATURAL, number of positions to shift
--|                                          default is 1.
--|
--|     Result         : Shifted std_ulogic_vector
--|
--|     NOTE           : Defaults not allowed for synthesis.
--|
--|     Use            :
--|                      SIGNAL acc   : std_ulogic_vector ( 15 DOWNTO 0);
--|                      SIGNAL carry : std_ulogic;
--|
--|                      SregShift ( acc, acc, carry, '1', '0',3 );
--|-----------------------------------------------------------------------------
   PROCEDURE SregShift ( CONSTANT SrcReg    : IN std_ulogic_vector;
                         SIGNAL DstReg    : INOUT std_ulogic_vector;
                         SIGNAL ShiftO    : OUT std_ulogic; 
                         CONSTANT direction : IN std_ulogic
                     -- synopsys synthesis_off
						      := '1'
                     -- synopsys synthesis_on
                                                            ;
                         CONSTANT FillVal   : IN std_ulogic  
                     -- synopsys synthesis_off
						      := '0'
                     -- synopsys synthesis_on
                                                            ;
                         CONSTANT Nbits     : IN Natural
                     -- synopsys synthesis_off
						       := 1 
                     -- synopsys synthesis_on
                      ) IS 
	CONSTANT dlen      : INTEGER := DstReg'LENGTH;
        VARIABLE r         : STD_ULOGIC_VECTOR (SrcReg'LENGTH - 1 DOWNTO 0);
        VARIABLE src_copy  : STD_ULOGIC_VECTOR (SrcReg'LENGTH - 1 DOWNTO 0 );
        VARIABLE dst_copy  : STD_ULOGIC_VECTOR (DstReg'LENGTH - 1 DOWNTO 0 );
        VARIABLE Shiftout  : STD_ULOGIC;
   BEGIN
       src_copy   := SrcReg;
       dst_copy   := DstReg;
 -- synopsys translate_off    
    --  Null range Check
    --  if input vector is of zero length
       IF ( SrcReg'LENGTH = 0) THEN
           ASSERT false
           REPORT " SregShift --- input bit_vector   is null  "
           SEVERITY ERROR;
           dst_copy := (OTHERS => FillVal);
           DstReg    <= dst_copy after DefaultRegDelay;
           ShiftO <= '0' after DefaultRegDelay;
           Return;
       ELSIF (DstReg'LENGTH = 0) THEN
           ASSERT false
           REPORT " SregShift --- output vector is  null  "
           SEVERITY ERROR;
         -- set shift out bit at least
           IF ( direction /= '0') THEN
               ShiftO <= src_copy(SrcReg'LENGTH - Nbits) after DefaultRegDelay;
           ELSE 
               ShiftO <= src_copy(Nbits - 1) after DefaultRegDelay;
           END IF;
           RETURN;
      END IF;
-- synopsys translate_on
    -- None of the registers is null, perform shift operation
      IF (direction /= '0') THEN                                 --  left shift
           RegShift_Left(src_copy, r, Shiftout, FillVal, Nbits);
      ELSE                                                       -- right shift
           RegShift_Right(src_copy, r, Shiftout, FillVal, Nbits);
      END IF;
      -- determine length of the result
      IF (dlen <= SrcReg'LENGTH) THEN
		for i IN dlen - 1 downto 0 Loop
			dst_copy(i) := r(i);
                end loop;
      ELSE
		for i IN SrcReg'LENGTH - 1 downto 0 Loop
			dst_copy(i) := r(i);
                end loop;
      END IF;
      DstReg <= dst_copy 
		-- synopsys translate_off     
			after DefaultRegDelay
		-- synopsys translate_on
       						;
      ShiftO <= Shiftout 
		-- synopsys translate_off     
			after DefaultRegDelay
		-- synopsys translate_on
       						;
      RETURN;
   END SregShift;
     -------------------------------------------------------------------------------
     --     Function Name : RegEqual
     -- 1.2.49
     --     Overloading   : Input parameter TYPEs.
     --
     --     Purpose       : Compute equality relation for bit_vector
     --
     --     Parameters    : l       - input bit_vector | INTEGER
     --                     r       - input bit_vector | INTEGER
     --                     SrcRegMode - input regmode_type, indicating the format of
     --                               the bit_vector operands (l,r).
     --                               Default is TwosComp.
     --
     --     Result        : BOOLEAN | bit. 
     --
     --     NOTE          : The operands may be of any length, and may be different
     --                     lengths.
     --
     --                     Overloading not defined for both inputs of INTEGER type.
     --     Use           :
     --                      VARIABLE a, b : bit_vector ( 7 DOWNTO 0 );
     --                      IF ( RegEqual ( a, b, TwosComp)   )  THEN
     --
     --     See Also      : RegLessThanOrEqual, RegGreaterThan, RegGreaterThanOrEqual.
     -------------------------------------------------------------------------------
     FUNCTION RegEqual     ( CONSTANT l          : IN bit_vector;
			     CONSTANT r          : IN bit_vector;
			     CONSTANT SrcRegMode : IN regmode_type
                     -- synopsys synthesis_off
							      := DefaultRegMode 
                     -- synopsys synthesis_on
			   ) RETURN bit IS
       CONSTANT resltlen : INTEGER := MAXIMUM (l'LENGTH, r'LENGTH);
       VARIABLE vl, vr   : BIT_VECTOR (resltlen - 1 DOWNTO 0);
     BEGIN
        -- synopsys translate_off
	-- Null range check
	IF ( (l'LENGTH = 0) AND (r'LENGTH = 0) ) THEN   
	      ASSERT false 
	      REPORT "  --- Both left and right vectors have null range "
	      SEVERITY ERROR;
              return( '0');
         ELSIF( l'LENGTH = 0) THEN        -- left input is of null range
    	      ASSERT false
	      REPORT " --- left input has null range "
	      SEVERITY ERROR;
              return('0');

         ELSIF( r'LENGTH = 0) THEN        -- right  input is of null range
	      ASSERT false
	      REPORT " --- right input has null range "
	      SEVERITY ERROR;
              RETURN ('0');
         END IF;
	-- synopsys translate_on        
 	-- input are not null so sign extend them to the same length
	vl := SignExtend(l, resltlen, l'LEFT, SrcRegMode);
	vr := SignExtend(r, resltlen, r'LEFT, SrcRegMode);
       	return( To_Bit_loc( Equal(vl, vr)));
     END RegEqual; 
     -----------------------------------------------------------------------------
     FUNCTION RegEqual    (  CONSTANT l        : IN bit_vector;
			     CONSTANT r        : IN bit_vector;
			     CONSTANT SrcRegMode : IN regmode_type
                     -- synopsys synthesis_off
							      := DefaultRegMode 
                     -- synopsys synthesis_on
			   ) RETURN BOOLEAN IS
       CONSTANT resltlen : INTEGER := MAXIMUM (l'LENGTH, r'LENGTH);
       VARIABLE vl, vr   : BIT_VECTOR (resltlen - 1 DOWNTO 0);
     BEGIN
        -- synopsys translate_off
	-- Null range check
	IF ( (l'LENGTH = 0) AND (r'LENGTH = 0) ) THEN   
	      ASSERT false 
	      REPORT "  --- Both left and right vectors have null range "
	      SEVERITY ERROR;
              return( false);
         ELSIF( l'LENGTH = 0) THEN        -- left input is of null range
    	      ASSERT false
	      REPORT " --- left input has null range "
	      SEVERITY ERROR;
              return(false);

         ELSIF( r'LENGTH = 0) THEN        -- right  input is of null range
	      ASSERT false
	      REPORT " --- right input has null range "
	      SEVERITY ERROR;
              RETURN (false);
         END IF;
	-- synopsys translate_on        
 	-- input are not null so sign extend them to the same length
	vl := SignExtend(l, resltlen, l'LEFT, SrcRegMode);
	vr := SignExtend(r, resltlen, r'LEFT, SrcRegMode);
	return ( Equal(vl, vr));
     END RegEqual; 
     -- -----------------------------------------------------------------------------
     FUNCTION RegEqual     ( CONSTANT l          : IN bit_vector;
			     CONSTANT r          : IN INTEGER;
			     CONSTANT SrcRegMode : IN regmode_type
                     -- synopsys synthesis_off
					         	      := DefaultRegMode 
                     -- synopsys synthesis_on
			   ) RETURN BOOLEAN IS
	VARIABLE vl, vr    : bit_vector(IntegerBitLength - 1 DOWNTO 0);
     BEGIN
	-- synopsys translate_off
	-- Null range check
	 IF( l'LENGTH = 0) THEN        -- left input is of null range
    	      ASSERT false
	      REPORT " --- left input has null range "
	      SEVERITY ERROR;
              return(false);
         END IF;
	-- synopsys translate_on        
	-- input are not null so sign extend them to the same length
        -- Convert to bit_vector for comparison to allow any length input vector.
        vr := To_BitVector ( r, IntegerBitLength, SrcRegMode );
 	vl := SignExtend(l, IntegerBitLength, l'LEFT, SrcRegMode);
       	return (Equal(vl, vr));
     END RegEqual; 
     -------------------------------------------------------------------------------
     FUNCTION RegEqual    (  CONSTANT l          : IN INTEGER;
			     CONSTANT r          : IN bit_vector;
			     CONSTANT SrcRegMode : IN regmode_type
                     -- synopsys synthesis_off
					         	      := DefaultRegMode 
                     -- synopsys synthesis_on
			   ) RETURN BOOLEAN IS
       VARIABLE vl, vr    : bit_vector(IntegerBitLength - 1 DOWNTO 0);
     BEGIN
	-- synopsys translate_off
	-- Null range check
	 IF( r'LENGTH = 0) THEN        -- right input is of null range
    	      ASSERT false
	      REPORT " --- left input has null range "
	      SEVERITY ERROR;
              return(false);
         END IF;
	-- synopsys translate_on        
	-- input are not null so sign extend them to the same length
        -- Convert to bit_vector for comparison to allow any length input vector.
        vl := To_BitVector ( l, IntegerBitLength, SrcRegMode );
 	vr := SignExtend(r, IntegerBitLength, r'LEFT, SrcRegMode);
	return (Equal(vl, vr));
     END RegEqual; 
     -------------------------------------------------------------------------------
     FUNCTION RegEqual     ( CONSTANT l          : IN bit_vector;
			     CONSTANT r          : IN INTEGER;
			     CONSTANT SrcRegMode : IN regmode_type 
                     -- synopsys synthesis_off
					         	      := DefaultRegMode 
                     -- synopsys synthesis_on
			   ) RETURN bit IS
	VARIABLE vl, vr    : bit_vector(IntegerBitLength - 1 DOWNTO 0);
     BEGIN
	-- synopsys translate_off
	-- Null range check
	 IF( l'LENGTH = 0) THEN        -- left input is of null range
    	      ASSERT false
	      REPORT " --- left input has null range "
	      SEVERITY ERROR;
              return('0');
         END IF;
	-- synopsys translate_on        
	-- input are not null so sign extend them to the same length
        -- Convert to bit_vector for comparison to allow any length input vector.
        vr := To_BitVector ( r, IntegerBitLength, SrcRegMode );
 	vl := SignExtend(l, IntegerBitLength, l'LEFT, SrcRegMode);
       	return ( To_Bit_loc(Equal(vl, vr)));
     END RegEqual; 
     -------------------------------------------------------------------------------
     FUNCTION RegEqual    (  CONSTANT l          : IN INTEGER;
			     CONSTANT r          : IN bit_vector;
			     CONSTANT SrcRegMode : IN regmode_type 
                     -- synopsys synthesis_off
					         	      := DefaultRegMode 
                     -- synopsys synthesis_on
			   ) RETURN bit IS
       VARIABLE vl, vr    : bit_vector(IntegerBitLength - 1 DOWNTO 0);
     BEGIN
	-- synopsys translate_off
	-- Null range check
	 IF( r'LENGTH = 0) THEN        -- right input is of null range
    	      ASSERT false
	      REPORT " --- left input has null range "
	      SEVERITY ERROR;
              return('0');
         END IF;
	-- synopsys translate_on        
	-- input are not null so sign extend them to the same length
        -- Convert to bit_vector for comparison to allow any length input vector.
        vl := To_BitVector ( l, IntegerBitLength, SrcRegMode );
 	vr := SignExtend(r, IntegerBitLength, r'LEFT, SrcRegMode);
	return (To_Bit_loc(Equal(vl, vr)));
     END RegEqual; 
     -------------------------------------------------------------------------------
     --     Function Name : RegEqual
     --
     --     Overloading   : Input parameter TYPEs.
     --    
     --     Purpose       : Compute equality relation for std_logic_vectors
     --     
     --     Parameters    : l       - input std_logic_vector | INTEGER
     --                     r       - input std_logic_vector | INTEGER
     --                     SrcRegMode - input regmode_type, indicating the format of
     --                               the std_logic_vector operands (l,r).
     --                               Default is TwosComp.
     --     
     --     Result        : BOOLEAN relation. A TRUE value is returned if: l = r
     --
     --     NOTE          : The operands may be of any length, and may be different
     --                     lengths. 
     --
     --                     Overloading not defined for both inputs of INTEGER type.
     --
     --                     Any time the comparison reaches an index that has an 'X' as an
     --                     array element, the comparison is deemed indeterminate and will 
     --                     return false in case of boolean and '0' incase of 
     --                     std_ulogic for synthesis purposes.
     --     Use           : 
     --                      VARIABLE a, b : std_logic_vector ( 7 DOWNTO 0 );
     --                      IF ( RegEqual ( a, b, TwosComp)   )  THEN 
     --     
     --     See Also      :  RegLessThan, RegLessThanOrEqual, RegGreaterThan, 
     --                     RegGreaterThanOrEqual.
     -------------------------------------------------------------------------------
     FUNCTION RegEqual     ( CONSTANT l          : IN std_logic_vector;
			     CONSTANT r          : IN std_logic_vector;
			     CONSTANT SrcRegMode : IN regmode_type
                     -- synopsys synthesis_off
							      := DefaultRegMode 
                     -- synopsys synthesis_on
			   ) RETURN std_ulogic IS
       CONSTANT resltlen : INTEGER := MAXIMUM (l'LENGTH, r'LENGTH);
       VARIABLE vl, vr   : std_logic_vector (resltlen - 1 DOWNTO 0);
     BEGIN
        -- synopsys translate_off
	-- Null range check
	IF ( (l'LENGTH = 0) AND (r'LENGTH = 0) ) THEN   
	      ASSERT false 
	      REPORT "  --- Both left and right vectors have null range "
	      SEVERITY ERROR;
              return( '0');
         ELSIF( l'LENGTH = 0) THEN        -- left input is of null range
    	      ASSERT false
	      REPORT " --- left input has null range "
	      SEVERITY ERROR;
              return('0');

         ELSIF( r'LENGTH = 0) THEN        -- right  input is of null range
	      ASSERT false
	      REPORT " --- right input has null range "
	      SEVERITY ERROR;
              RETURN ('0');
         END IF;
	-- synopsys translate_on        
 	-- input are not null so sign extend them to the same length
	vl := SignExtend(l, resltlen, l'LEFT, SrcRegMode);
	vr := SignExtend(r, resltlen, r'LEFT, SrcRegMode);
       	return( To_StdULogic_loc( Equal(vl, vr)));
     END RegEqual; 
     -----------------------------------------------------------------------------
     FUNCTION RegEqual    (  CONSTANT l        : IN std_logic_vector;
			     CONSTANT r        : IN std_logic_vector;
			     CONSTANT SrcRegMode : IN regmode_type
                     -- synopsys synthesis_off
							      := DefaultRegMode 
                     -- synopsys synthesis_on
			   ) RETURN BOOLEAN IS
       CONSTANT resltlen : INTEGER := MAXIMUM (l'LENGTH, r'LENGTH);
       VARIABLE vl, vr   : STD_LOGIC_VECTOR (resltlen - 1 DOWNTO 0);
     BEGIN
        -- synopsys translate_off
	-- Null range check
	IF ( (l'LENGTH = 0) AND (r'LENGTH = 0) ) THEN   
	      ASSERT false 
	      REPORT "  --- Both left and right vectors have null range "
	      SEVERITY ERROR;
              return( false);
         ELSIF( l'LENGTH = 0) THEN        -- left input is of null range
    	      ASSERT false
	      REPORT " --- left input has null range "
	      SEVERITY ERROR;
              return(false);

         ELSIF( r'LENGTH = 0) THEN        -- right  input is of null range
	      ASSERT false
	      REPORT " --- right input has null range "
	      SEVERITY ERROR;
              RETURN (false);
         END IF;
	-- synopsys translate_on        
 	-- input are not null so sign extend them to the same length
	vl := SignExtend(l, resltlen, l'LEFT, SrcRegMode);
	vr := SignExtend(r, resltlen, r'LEFT, SrcRegMode);
	return ( Equal(vl, vr));
     END RegEqual; 
     -- -----------------------------------------------------------------------------
     FUNCTION RegEqual     ( CONSTANT l          : IN std_logic_vector;
			     CONSTANT r          : IN INTEGER;
			     CONSTANT SrcRegMode : IN regmode_type
                     -- synopsys synthesis_off
					         	      := DefaultRegMode 
                     -- synopsys synthesis_on
			   ) RETURN BOOLEAN IS
	VARIABLE vl, vr    : std_logic_vector(IntegerBitLength - 1 DOWNTO 0);
     BEGIN
	-- synopsys translate_off
	-- Null range check
	 IF( l'LENGTH = 0) THEN        -- left input is of null range
    	      ASSERT false
	      REPORT " --- left input has null range "
	      SEVERITY ERROR;
              return(false);
         END IF;
	-- synopsys translate_on        
	-- input are not null so sign extend them to the same length
        -- Convert to std_logic_vector for comparison to allow any length input vector.
        vr := To_StdLogicVector ( r, IntegerBitLength, SrcRegMode );
 	vl := SignExtend(l, IntegerBitLength, l'LEFT, SrcRegMode);
       	return (Equal(vl, vr));
     END RegEqual; 
     -------------------------------------------------------------------------------
     FUNCTION RegEqual    (  CONSTANT l          : IN INTEGER;
			     CONSTANT r          : IN std_logic_vector;
			     CONSTANT SrcRegMode : IN regmode_type
                     -- synopsys synthesis_off
					         	      := DefaultRegMode 
                     -- synopsys synthesis_on
			   ) RETURN BOOLEAN IS
       VARIABLE vl, vr    : std_logic_vector(IntegerBitLength - 1 DOWNTO 0);
     BEGIN
	-- synopsys translate_off
	-- Null range check
	 IF( r'LENGTH = 0) THEN        -- right input is of null range
    	      ASSERT false
	      REPORT " --- left input has null range "
	      SEVERITY ERROR;
              return(false);
         END IF;
	-- synopsys translate_on        
	-- input are not null so sign extend them to the same length
        -- Convert to std_logic_vector for comparison to allow any length input vector.
        vl := To_StdLogicVector ( l, IntegerBitLength, SrcRegMode );
 	vr := SignExtend(r, IntegerBitLength, r'LEFT, SrcRegMode);
	return (Equal(vl, vr));
     END RegEqual; 
     -------------------------------------------------------------------------------
     FUNCTION RegEqual     ( CONSTANT l          : IN std_logic_vector;
			     CONSTANT r          : IN INTEGER;
			     CONSTANT SrcRegMode : IN regmode_type 
                     -- synopsys synthesis_off
					         	      := DefaultRegMode 
                     -- synopsys synthesis_on
			   ) RETURN std_ulogic IS
	VARIABLE vl, vr    : std_logic_vector(IntegerBitLength - 1 DOWNTO 0);
     BEGIN
	-- synopsys translate_off
	-- Null range check
	 IF( l'LENGTH = 0) THEN        -- left input is of null range
    	      ASSERT false
	      REPORT " --- left input has null range "
	      SEVERITY ERROR;
              return('0');
         END IF;
	-- synopsys translate_on        
	-- input are not null so sign extend them to the same length
        -- Convert to std_logic_vector for comparison to allow any length input vector.
        vr := To_StdLogicVector ( r, IntegerBitLength, SrcRegMode );
 	vl := SignExtend(l, IntegerBitLength, l'LEFT, SrcRegMode);
       	return ( To_StdULogic_loc(Equal(vl, vr)));
     END RegEqual; 
     -------------------------------------------------------------------------------
     FUNCTION RegEqual    (  CONSTANT l          : IN INTEGER;
			     CONSTANT r          : IN std_logic_vector;
			     CONSTANT SrcRegMode : IN regmode_type 
                     -- synopsys synthesis_off
					         	      := DefaultRegMode 
                     -- synopsys synthesis_on
			   ) RETURN std_ulogic IS
       VARIABLE vl, vr    : std_logic_vector(IntegerBitLength - 1 DOWNTO 0);
     BEGIN
	-- synopsys translate_off
	-- Null range check
	 IF( r'LENGTH = 0) THEN        -- right input is of null range
    	      ASSERT false
	      REPORT " --- left input has null range "
	      SEVERITY ERROR;
              return('0');
         END IF;
	-- synopsys translate_on        
	-- input are not null so sign extend them to the same length
        -- Convert to std_logic_vector for comparison to allow any length input vector.
        vl := To_StdLogicVector ( l, IntegerBitLength, SrcRegMode );
 	vr := SignExtend(r, IntegerBitLength, r'LEFT, SrcRegMode);
	return (To_StdULogic_loc(Equal(vl, vr)));
     END RegEqual; 
     -------------------------------------------------------------------------------
     --     Function Name : RegEqual
     --
     --     Overloading   : Input parameter TYPEs.
     --    
     --     Purpose       : Compute equality relation for std_ulogic_vectors
     --     
     --     Parameters    : l       - input std_ulogic_vector | INTEGER
     --                     r       - input std_ulogic_vector | INTEGER
     --                     SrcRegMode - input regmode_type, indicating the format of
     --                               the std_ulogic_vector operands (l,r).
     --                               Default is TwosComp.
     --     
     --     Result        : BOOLEAN relation. A TRUE value is returned if: l = r
     --
     --     NOTE          : The operands may be of any length, and may be different
     --                     lengths. 
     --
     --                     Overloading not defined for both inputs of INTEGER type.
     --
     --                     Any time the comparison reaches an index that has an 'X' as an
     --                     array element, the comparison is deemed indeterminate and will 
     --                     return false in case of boolean and '0' incase of 
     --                     std_ulogic for  synthesis purposes.
     --     Use           : 
     --                      VARIABLE a, b : std_ulogic_vector ( 7 DOWNTO 0 );
     --                      IF ( RegEqual ( a, b, TwosComp)   )  THEN 
     --     
     --     See Also      :  RegLessThan, RegLessThanOrEqual, RegGreaterThan, 
     --                     RegGreaterThanOrEqual.
     -------------------------------------------------------------------------------
     FUNCTION RegEqual     ( CONSTANT l          : IN std_ulogic_vector;
			     CONSTANT r          : IN std_ulogic_vector;
			     CONSTANT SrcRegMode : IN regmode_type
                     -- synopsys synthesis_off
							      := DefaultRegMode 
                     -- synopsys synthesis_on
			   ) RETURN std_ulogic IS
       CONSTANT resltlen : INTEGER := MAXIMUM (l'LENGTH, r'LENGTH);
       VARIABLE vl, vr   : std_ulogic_vector (resltlen - 1 DOWNTO 0);
     BEGIN
        -- synopsys translate_off
	-- Null range check
	IF ( (l'LENGTH = 0) AND (r'LENGTH = 0) ) THEN   
	      ASSERT false 
	      REPORT "  --- Both left and right vectors have null range "
	      SEVERITY ERROR;
              return( '0');
         ELSIF( l'LENGTH = 0) THEN        -- left input is of null range
    	      ASSERT false
	      REPORT " --- left input has null range "
	      SEVERITY ERROR;
              return('0');

         ELSIF( r'LENGTH = 0) THEN        -- right  input is of null range
	      ASSERT false
	      REPORT " --- right input has null range "
	      SEVERITY ERROR;
              RETURN ('0');
         END IF;
	-- synopsys translate_on        
 	-- input are not null so sign extend them to the same length
	vl := SignExtend(l, resltlen, l'LEFT, SrcRegMode);
	vr := SignExtend(r, resltlen, r'LEFT, SrcRegMode);
       	return( To_StdULogic_loc( Equal(vl, vr)));
     END RegEqual; 
     -----------------------------------------------------------------------------
     FUNCTION RegEqual    (  CONSTANT l        : IN std_ulogic_vector;
			     CONSTANT r        : IN std_ulogic_vector;
			     CONSTANT SrcRegMode : IN regmode_type
                     -- synopsys synthesis_off
							      := DefaultRegMode 
                     -- synopsys synthesis_on
			   ) RETURN BOOLEAN IS
       CONSTANT resltlen : INTEGER := MAXIMUM (l'LENGTH, r'LENGTH);
       VARIABLE vl, vr   : STD_ULOGIC_VECTOR (resltlen - 1 DOWNTO 0);
     BEGIN
        -- synopsys translate_off
	-- Null range check
	IF ( (l'LENGTH = 0) AND (r'LENGTH = 0) ) THEN   
	      ASSERT false 
	      REPORT "  --- Both left and right vectors have null range "
	      SEVERITY ERROR;
              return( false);
         ELSIF( l'LENGTH = 0) THEN        -- left input is of null range
    	      ASSERT false
	      REPORT " --- left input has null range "
	      SEVERITY ERROR;
              return(false);

         ELSIF( r'LENGTH = 0) THEN        -- right  input is of null range
	      ASSERT false
	      REPORT " --- right input has null range "
	      SEVERITY ERROR;
              RETURN (false);
         END IF;
	-- synopsys translate_on        
 	-- input are not null so sign extend them to the same length
	vl := SignExtend(l, resltlen, l'LEFT, SrcRegMode);
	vr := SignExtend(r, resltlen, r'LEFT, SrcRegMode);
	return ( Equal(vl, vr));
     END RegEqual; 
     -- -----------------------------------------------------------------------------
     FUNCTION RegEqual     ( CONSTANT l          : IN std_ulogic_vector;
			     CONSTANT r          : IN INTEGER;
			     CONSTANT SrcRegMode : IN regmode_type
                     -- synopsys synthesis_off
					         	      := DefaultRegMode 
                     -- synopsys synthesis_on
			   ) RETURN BOOLEAN IS
	VARIABLE vl, vr    : std_ulogic_vector(IntegerBitLength - 1 DOWNTO 0);
     BEGIN
	-- synopsys translate_off
	-- Null range check
	 IF( l'LENGTH = 0) THEN        -- left input is of null range
    	      ASSERT false
	      REPORT " --- left input has null range "
	      SEVERITY ERROR;
              return(false);
         END IF;
	-- synopsys translate_on        
	-- input are not null so sign extend them to the same length
        -- Convert to std_ulogic_vector for comparison to allow any length input vector.
        vr := To_StdULogicVector ( r, IntegerBitLength, SrcRegMode );
 	vl := SignExtend(l, IntegerBitLength, l'LEFT, SrcRegMode);
       	return (Equal(vl, vr));
     END RegEqual; 
     -------------------------------------------------------------------------------
     FUNCTION RegEqual    (  CONSTANT l          : IN INTEGER;
			     CONSTANT r          : IN std_ulogic_vector;
			     CONSTANT SrcRegMode : IN regmode_type
                     -- synopsys synthesis_off
					         	      := DefaultRegMode 
                     -- synopsys synthesis_on
			   ) RETURN BOOLEAN IS
       VARIABLE vl, vr    : std_ulogic_vector(IntegerBitLength - 1 DOWNTO 0);
     BEGIN
	-- synopsys translate_off
	-- Null range check
	 IF( r'LENGTH = 0) THEN        -- right input is of null range
    	      ASSERT false
	      REPORT " --- left input has null range "
	      SEVERITY ERROR;
              return(false);
         END IF;
	-- synopsys translate_on        
	-- input are not null so sign extend them to the same length
        -- Convert to std_ulogic_vector for comparison to allow any length input vector.
        vl := To_StdULogicVector ( l, IntegerBitLength, SrcRegMode );
 	vr := SignExtend(r, IntegerBitLength, r'LEFT, SrcRegMode);
	return (Equal(vl, vr));
     END RegEqual; 
     -------------------------------------------------------------------------------
     FUNCTION RegEqual     ( CONSTANT l          : IN std_ulogic_vector;
			     CONSTANT r          : IN INTEGER;
			     CONSTANT SrcRegMode : IN regmode_type 
                     -- synopsys synthesis_off
					         	      := DefaultRegMode 
                     -- synopsys synthesis_on
			   ) RETURN std_ulogic IS
	VARIABLE vl, vr    : std_ulogic_vector(IntegerBitLength - 1 DOWNTO 0);
     BEGIN
	-- synopsys translate_off
	-- Null range check
	 IF( l'LENGTH = 0) THEN        -- left input is of null range
    	      ASSERT false
	      REPORT " --- left input has null range "
	      SEVERITY ERROR;
              return('0');
         END IF;
	-- synopsys translate_on        
	-- input are not null so sign extend them to the same length
        -- Convert to std_ulogic_vector for comparison to allow any length input vector.
        vr := To_StdULogicVector ( r, IntegerBitLength, SrcRegMode );
 	vl := SignExtend(l, IntegerBitLength, l'LEFT, SrcRegMode);
       	return ( To_StdULogic_loc(Equal(vl, vr)));
     END RegEqual; 
     -------------------------------------------------------------------------------
     FUNCTION RegEqual    (  CONSTANT l          : IN INTEGER;
			     CONSTANT r          : IN std_ulogic_vector;
			     CONSTANT SrcRegMode : IN regmode_type 
                     -- synopsys synthesis_off
					         	      := DefaultRegMode 
                     -- synopsys synthesis_on
			   ) RETURN std_ulogic IS
       VARIABLE vl, vr    : std_ulogic_vector(IntegerBitLength - 1 DOWNTO 0);
     BEGIN
	-- synopsys translate_off
	-- Null range check
	 IF( r'LENGTH = 0) THEN        -- right input is of null range
    	      ASSERT false
	      REPORT " --- left input has null range "
	      SEVERITY ERROR;
              return('0');
         END IF;
	-- synopsys translate_on        
	-- input are not null so sign extend them to the same length
        -- Convert to std_ulogic_vector for comparison to allow any length input vector.
        vl := To_StdULogicVector ( l, IntegerBitLength, SrcRegMode );
 	vr := SignExtend(r, IntegerBitLength, r'LEFT, SrcRegMode);
	return (To_StdULogic_loc(Equal(vl, vr)));
     END RegEqual; 
     -------------------------------------------------------------------------------
     --     Function Name : RegNotEqual
     -- 1.2.49
     --     Overloading   : Input parameter TYPEs.
     --
     --     Purpose       : Compute un-equality relation for bit_vector
     --
     --     Parameters    : l       - input bit_vector | INTEGER
     --                     r       - input bit_vector | INTEGER
     --                     SrcRegMode - input regmode_type, indicating the format of
     --                               the bit_vector operands (l,r).
     --                               Default is TwosComp.
     --
     --     Result        : BOOLEAN | bit. 
     --
     --     NOTE          : The operands may be of any length, and may be different
     --                     lengths.
     --
     --                     Overloading not defined for both inputs of INTEGER type.
     --
     --     Use           :
     --                      VARIABLE a, b : bit_vector ( 7 DOWNTO 0 );
     --                      IF ( RegNotEqual ( a, b, TwosComp)   )  THEN
     --
     --     See Also      : RegLessThanOrEqual, RegGreaterThan, RegGreaterThanOrEqual.
     -------------------------------------------------------------------------------
     FUNCTION RegNotEqual     ( CONSTANT l          : IN bit_vector;
			     CONSTANT r          : IN bit_vector;
			     CONSTANT SrcRegMode : IN regmode_type
                     -- synopsys synthesis_off
							      := DefaultRegMode 
                     -- synopsys synthesis_on
			   ) RETURN bit IS
       CONSTANT resltlen : INTEGER := MAXIMUM (l'LENGTH, r'LENGTH);
       VARIABLE vl, vr   : BIT_VECTOR (resltlen - 1 DOWNTO 0);
     BEGIN
        -- synopsys translate_off
	-- Null range check
	IF ( (l'LENGTH = 0) AND (r'LENGTH = 0) ) THEN   
	      ASSERT false 
	      REPORT "  --- Both left and right vectors have null range "
	      SEVERITY ERROR;
              return( '0');
         ELSIF( l'LENGTH = 0) THEN        -- left input is of null range
    	      ASSERT false
	      REPORT " --- left input has null range "
	      SEVERITY ERROR;
              return('0');

         ELSIF( r'LENGTH = 0) THEN        -- right  input is of null range
	      ASSERT false
	      REPORT " --- right input has null range "
	      SEVERITY ERROR;
              RETURN ('0');
         END IF;
	-- synopsys translate_on        
 	-- input are not null so sign extend them to the same length
	vl := SignExtend(l, resltlen, l'LEFT, SrcRegMode);
	vr := SignExtend(r, resltlen, r'LEFT, SrcRegMode);
       	return( To_Bit_loc( NotEqual(vl, vr)));
     END RegNotEqual; 
     -----------------------------------------------------------------------------
     FUNCTION RegNotEqual    (  CONSTANT l        : IN bit_vector;
			     CONSTANT r        : IN bit_vector;
			     CONSTANT SrcRegMode : IN regmode_type
                     -- synopsys synthesis_off
							      := DefaultRegMode 
                     -- synopsys synthesis_on
			   ) RETURN BOOLEAN IS
       CONSTANT resltlen : INTEGER := MAXIMUM (l'LENGTH, r'LENGTH);
       VARIABLE vl, vr   : BIT_VECTOR (resltlen - 1 DOWNTO 0);
     BEGIN
        -- synopsys translate_off
	-- Null range check
	IF ( (l'LENGTH = 0) AND (r'LENGTH = 0) ) THEN   
	      ASSERT false 
	      REPORT "  --- Both left and right vectors have null range "
	      SEVERITY ERROR;
              return( false);
         ELSIF( l'LENGTH = 0) THEN        -- left input is of null range
    	      ASSERT false
	      REPORT " --- left input has null range "
	      SEVERITY ERROR;
              return(false);

         ELSIF( r'LENGTH = 0) THEN        -- right  input is of null range
	      ASSERT false
	      REPORT " --- right input has null range "
	      SEVERITY ERROR;
              RETURN (false);
         END IF;
	-- synopsys translate_on        
 	-- input are not null so sign extend them to the same length
	vl := SignExtend(l, resltlen, l'LEFT, SrcRegMode);
	vr := SignExtend(r, resltlen, r'LEFT, SrcRegMode);
	return ( NotEqual(vl, vr));
     END RegNotEqual; 
     -- -----------------------------------------------------------------------------
     FUNCTION RegNotEqual     ( CONSTANT l          : IN bit_vector;
			     CONSTANT r          : IN INTEGER;
			     CONSTANT SrcRegMode : IN regmode_type
                     -- synopsys synthesis_off
					         	      := DefaultRegMode 
                     -- synopsys synthesis_on
			   ) RETURN BOOLEAN IS
	VARIABLE vl, vr    : bit_vector(IntegerBitLength - 1 DOWNTO 0);
     BEGIN
	-- synopsys translate_off
	-- Null range check
	 IF( l'LENGTH = 0) THEN        -- left input is of null range
    	      ASSERT false
	      REPORT " --- left input has null range "
	      SEVERITY ERROR;
              return(false);
         END IF;
	-- synopsys translate_on        
	-- input are not null so sign extend them to the same length
        -- Convert to bit_vector for comparison to allow any length input vector.
        vr := To_BitVector ( r, IntegerBitLength, SrcRegMode );
 	vl := SignExtend(l, IntegerBitLength, l'LEFT, SrcRegMode);
       	return (NotEqual(vl, vr));
     END RegNotEqual; 
     -------------------------------------------------------------------------------
     FUNCTION RegNotEqual    (  CONSTANT l          : IN INTEGER;
			     CONSTANT r          : IN bit_vector;
			     CONSTANT SrcRegMode : IN regmode_type
                     -- synopsys synthesis_off
					         	      := DefaultRegMode 
                     -- synopsys synthesis_on
			   ) RETURN BOOLEAN IS
       VARIABLE vl, vr    : bit_vector(IntegerBitLength - 1 DOWNTO 0);
     BEGIN
	-- synopsys translate_off
	-- Null range check
	 IF( r'LENGTH = 0) THEN        -- right input is of null range
    	      ASSERT false
	      REPORT " --- left input has null range "
	      SEVERITY ERROR;
              return(false);
         END IF;
	-- synopsys translate_on        
	-- input are not null so sign extend them to the same length
        -- Convert to bit_vector for comparison to allow any length input vector.
        vl := To_BitVector ( l, IntegerBitLength, SrcRegMode );
 	vr := SignExtend(r, IntegerBitLength, r'LEFT, SrcRegMode);
	return (NotEqual(vl, vr));
     END RegNotEqual; 
     -------------------------------------------------------------------------------
     FUNCTION RegNotEqual     ( CONSTANT l          : IN bit_vector;
			     CONSTANT r          : IN INTEGER;
			     CONSTANT SrcRegMode : IN regmode_type 
                     -- synopsys synthesis_off
					         	      := DefaultRegMode 
                     -- synopsys synthesis_on
			   ) RETURN bit IS
	VARIABLE vl, vr    : bit_vector(IntegerBitLength - 1 DOWNTO 0);
     BEGIN
	-- synopsys translate_off
	-- Null range check
	 IF( l'LENGTH = 0) THEN        -- left input is of null range
    	      ASSERT false
	      REPORT " --- left input has null range "
	      SEVERITY ERROR;
              return('0');
         END IF;
	-- synopsys translate_on        
	-- input are not null so sign extend them to the same length
        -- Convert to bit_vector for comparison to allow any length input vector.
        vr := To_BitVector ( r, IntegerBitLength, SrcRegMode );
 	vl := SignExtend(l, IntegerBitLength, l'LEFT, SrcRegMode);
       	return ( To_Bit_loc(NotEqual(vl, vr)));
     END RegNotEqual; 
     -------------------------------------------------------------------------------
     FUNCTION RegNotEqual    (  CONSTANT l          : IN INTEGER;
			     CONSTANT r          : IN bit_vector;
			     CONSTANT SrcRegMode : IN regmode_type 
                     -- synopsys synthesis_off
					         	      := DefaultRegMode 
                     -- synopsys synthesis_on
			   ) RETURN bit IS
       VARIABLE vl, vr    : bit_vector(IntegerBitLength - 1 DOWNTO 0);
     BEGIN
	-- synopsys translate_off
	-- Null range check
	 IF( r'LENGTH = 0) THEN        -- right input is of null range
    	      ASSERT false
	      REPORT " --- left input has null range "
	      SEVERITY ERROR;
              return('0');
         END IF;
	-- synopsys translate_on        
	-- input are not null so sign extend them to the same length
        -- Convert to bit_vector for comparison to allow any length input vector.
        vl := To_BitVector ( l, IntegerBitLength, SrcRegMode );
 	vr := SignExtend(r, IntegerBitLength, r'LEFT, SrcRegMode);
	return (To_Bit_loc(NotEqual(vl, vr)));
     END RegNotEqual; 
     -------------------------------------------------------------------------------
     --     Function Name : RegNotEqual
     --
     --     Overloading   : Input parameter TYPEs.
     --    
     --     Purpose       : Compute un-equality relation for std_logic_vectors
     --     
     --     Parameters    : l       - input std_logic_vector | INTEGER
     --                     r       - input std_logic_vector | INTEGER
     --                     SrcRegMode - input regmode_type, indicating the format of
     --                               the std_logic_vector operands (l,r).
     --                               Default is TwosComp.
     --     
     --     Result        : BOOLEAN relation. A TRUE value is returned if: l = r
     --
     --     NOTE          : The operands may be of any length, and may be different
     --                     lengths. 
     --
     --                     Overloading not defined for both inputs of INTEGER type.
     --
     --                     Any time the comparison reaches an index that has an 'X' as an
     --                     array element, the comparison is deemed indeterminate and will 
     --                     return false in case of boolean and '0' incase of 
     --                     std_ulogic for   synthesis purposes.
     --     Use           : 
     --                      VARIABLE a, b : std_logic_vector ( 7 DOWNTO 0 );
     --                      IF ( RegNotEqual ( a, b, TwosComp)   )  THEN 
     --     
     --     See Also      :  RegLessThan, RegLessThanOrEqual, RegGreaterThan, 
     --                     RegGreaterThanOrEqual.
     -------------------------------------------------------------------------------
     FUNCTION RegNotEqual     ( CONSTANT l          : IN std_logic_vector;
			     CONSTANT r          : IN std_logic_vector;
			     CONSTANT SrcRegMode : IN regmode_type
                     -- synopsys synthesis_off
							      := DefaultRegMode 
                     -- synopsys synthesis_on
			   ) RETURN std_ulogic IS
       CONSTANT resltlen : INTEGER := MAXIMUM (l'LENGTH, r'LENGTH);
       VARIABLE vl, vr   : std_logic_vector (resltlen - 1 DOWNTO 0);
     BEGIN
        -- synopsys translate_off
	-- Null range check
	IF ( (l'LENGTH = 0) AND (r'LENGTH = 0) ) THEN   
	      ASSERT false 
	      REPORT "  --- Both left and right vectors have null range "
	      SEVERITY ERROR;
              return( '0');
         ELSIF( l'LENGTH = 0) THEN        -- left input is of null range
    	      ASSERT false
	      REPORT " --- left input has null range "
	      SEVERITY ERROR;
              return('0');

         ELSIF( r'LENGTH = 0) THEN        -- right  input is of null range
	      ASSERT false
	      REPORT " --- right input has null range "
	      SEVERITY ERROR;
              RETURN ('0');
         END IF;
	-- synopsys translate_on        
 	-- input are not null so sign extend them to the same length
	vl := SignExtend(l, resltlen, l'LEFT, SrcRegMode);
	vr := SignExtend(r, resltlen, r'LEFT, SrcRegMode);
       	return( To_StdULogic_loc( NotEqual(vl, vr)));
     END RegNotEqual; 
     -----------------------------------------------------------------------------
     FUNCTION RegNotEqual    (  CONSTANT l        : IN std_logic_vector;
			     CONSTANT r        : IN std_logic_vector;
			     CONSTANT SrcRegMode : IN regmode_type
                     -- synopsys synthesis_off
							      := DefaultRegMode 
                     -- synopsys synthesis_on
			   ) RETURN BOOLEAN IS
       CONSTANT resltlen : INTEGER := MAXIMUM (l'LENGTH, r'LENGTH);
       VARIABLE vl, vr   : STD_LOGIC_VECTOR (resltlen - 1 DOWNTO 0);
     BEGIN
        -- synopsys translate_off
	-- Null range check
	IF ( (l'LENGTH = 0) AND (r'LENGTH = 0) ) THEN   
	      ASSERT false 
	      REPORT "  --- Both left and right vectors have null range "
	      SEVERITY ERROR;
              return( false);
         ELSIF( l'LENGTH = 0) THEN        -- left input is of null range
    	      ASSERT false
	      REPORT " --- left input has null range "
	      SEVERITY ERROR;
              return(false);

         ELSIF( r'LENGTH = 0) THEN        -- right  input is of null range
	      ASSERT false
	      REPORT " --- right input has null range "
	      SEVERITY ERROR;
              RETURN (false);
         END IF;
	-- synopsys translate_on        
 	-- input are not null so sign extend them to the same length
	vl := SignExtend(l, resltlen, l'LEFT, SrcRegMode);
	vr := SignExtend(r, resltlen, r'LEFT, SrcRegMode);
	return ( NotEqual(vl, vr));
     END RegNotEqual; 
     -- -----------------------------------------------------------------------------
     FUNCTION RegNotEqual     ( CONSTANT l          : IN std_logic_vector;
			     CONSTANT r          : IN INTEGER;
			     CONSTANT SrcRegMode : IN regmode_type
                     -- synopsys synthesis_off
					         	      := DefaultRegMode 
                     -- synopsys synthesis_on
			   ) RETURN BOOLEAN IS
	VARIABLE vl, vr    : std_logic_vector(IntegerBitLength - 1 DOWNTO 0);
     BEGIN
	-- synopsys translate_off
	-- Null range check
	 IF( l'LENGTH = 0) THEN        -- left input is of null range
    	      ASSERT false
	      REPORT " --- left input has null range "
	      SEVERITY ERROR;
              return(false);
         END IF;
	-- synopsys translate_on        
	-- input are not null so sign extend them to the same length
        -- Convert to std_logic_vector for comparison to allow any length input vector.
        vr := To_StdLogicVector ( r, IntegerBitLength, SrcRegMode );
 	vl := SignExtend(l, IntegerBitLength, l'LEFT, SrcRegMode);
       	return (NotEqual(vl, vr));
     END RegNotEqual; 
     -------------------------------------------------------------------------------
     FUNCTION RegNotEqual    (  CONSTANT l          : IN INTEGER;
			     CONSTANT r          : IN std_logic_vector;
			     CONSTANT SrcRegMode : IN regmode_type
                     -- synopsys synthesis_off
					         	      := DefaultRegMode 
                     -- synopsys synthesis_on
			   ) RETURN BOOLEAN IS
       VARIABLE vl, vr    : std_logic_vector(IntegerBitLength - 1 DOWNTO 0);
     BEGIN
	-- synopsys translate_off
	-- Null range check
	 IF( r'LENGTH = 0) THEN        -- right input is of null range
    	      ASSERT false
	      REPORT " --- left input has null range "
	      SEVERITY ERROR;
              return(false);
         END IF;
	-- synopsys translate_on        
	-- input are not null so sign extend them to the same length
        -- Convert to std_logic_vector for comparison to allow any length input vector.
        vl := To_StdLogicVector ( l, IntegerBitLength, SrcRegMode );
 	vr := SignExtend(r, IntegerBitLength, r'LEFT, SrcRegMode);
	return (NotEqual(vl, vr));
     END RegNotEqual; 
     -------------------------------------------------------------------------------
     FUNCTION RegNotEqual     ( CONSTANT l          : IN std_logic_vector;
			     CONSTANT r          : IN INTEGER;
			     CONSTANT SrcRegMode : IN regmode_type 
                     -- synopsys synthesis_off
					         	      := DefaultRegMode 
                     -- synopsys synthesis_on
			   ) RETURN std_ulogic IS
	VARIABLE vl, vr    : std_logic_vector(IntegerBitLength - 1 DOWNTO 0);
     BEGIN
	-- synopsys translate_off
	-- Null range check
	 IF( l'LENGTH = 0) THEN        -- left input is of null range
    	      ASSERT false
	      REPORT " --- left input has null range "
	      SEVERITY ERROR;
              return('0');
         END IF;
	-- synopsys translate_on        
	-- input are not null so sign extend them to the same length
        -- Convert to std_logic_vector for comparison to allow any length input vector.
        vr := To_StdLogicVector ( r, IntegerBitLength, SrcRegMode );
 	vl := SignExtend(l, IntegerBitLength, l'LEFT, SrcRegMode);
       	return ( To_StdULogic_loc(NotEqual(vl, vr)));
     END RegNotEqual; 
     -------------------------------------------------------------------------------
     FUNCTION RegNotEqual    (  CONSTANT l          : IN INTEGER;
			     CONSTANT r          : IN std_logic_vector;
			     CONSTANT SrcRegMode : IN regmode_type 
                     -- synopsys synthesis_off
					         	      := DefaultRegMode 
                     -- synopsys synthesis_on
			   ) RETURN std_ulogic IS
       VARIABLE vl, vr    : std_logic_vector(IntegerBitLength - 1 DOWNTO 0);
     BEGIN
	-- synopsys translate_off
	-- Null range check
	 IF( r'LENGTH = 0) THEN        -- right input is of null range
    	      ASSERT false
	      REPORT " --- left input has null range "
	      SEVERITY ERROR;
              return('0');
         END IF;
	-- synopsys translate_on        
	-- input are not null so sign extend them to the same length
        -- Convert to std_logic_vector for comparison to allow any length input vector.
        vl := To_StdLogicVector ( l, IntegerBitLength, SrcRegMode );
 	vr := SignExtend(r, IntegerBitLength, r'LEFT, SrcRegMode);
	return (To_StdULogic_loc(NotEqual(vl, vr)));
     END RegNotEqual; 
     -------------------------------------------------------------------------------
     --     Function Name : RegNotEqual
     --
     --     Overloading   : Input parameter TYPEs.
     --    
     --     Purpose       : Compute un-equality relation for std_ulogic_vectors
     --     
     --     Parameters    : l       - input std_ulogic_vector | INTEGER
     --                     r       - input std_ulogic_vector | INTEGER
     --                     SrcRegMode - input regmode_type, indicating the format of
     --                               the std_ulogic_vector operands (l,r).
     --                               Default is TwosComp.
     --     
     --     Result        : BOOLEAN relation. A TRUE value is returned if: l = r
     --
     --     NOTE          : The operands may be of any length, and may be different
     --                     lengths. 
     --
     --                     Overloading not defined for both inputs of INTEGER type.
     --
     --                     Any time the comparison reaches an index that has an 'X' as an
     --                     array element, the comparison is deemed indeterminate and will 
     --                     return false in case of boolean and '0' incase of 
     --                     std_ulogic for synthesis purposes.
     --
     --     Use           : 
     --                      VARIABLE a, b : std_ulogic_vector ( 7 DOWNTO 0 );
     --                      IF ( RegNotEqual ( a, b, TwosComp)   )  THEN 
     --     
     --     See Also      :  RegLessThan, RegLessThanOrEqual, RegGreaterThan, 
     --                     RegGreaterThanOrEqual.
     -------------------------------------------------------------------------------
     FUNCTION RegNotEqual     ( CONSTANT l          : IN std_ulogic_vector;
			     CONSTANT r          : IN std_ulogic_vector;
			     CONSTANT SrcRegMode : IN regmode_type
                     -- synopsys synthesis_off
							      := DefaultRegMode 
                     -- synopsys synthesis_on
			   ) RETURN std_ulogic IS
       CONSTANT resltlen : INTEGER := MAXIMUM (l'LENGTH, r'LENGTH);
       VARIABLE vl, vr   : std_ulogic_vector (resltlen - 1 DOWNTO 0);
     BEGIN
        -- synopsys translate_off
	-- Null range check
	IF ( (l'LENGTH = 0) AND (r'LENGTH = 0) ) THEN   
	      ASSERT false 
	      REPORT "  --- Both left and right vectors have null range "
	      SEVERITY ERROR;
              return( '0');
         ELSIF( l'LENGTH = 0) THEN        -- left input is of null range
    	      ASSERT false
	      REPORT " --- left input has null range "
	      SEVERITY ERROR;
              return('0');

         ELSIF( r'LENGTH = 0) THEN        -- right  input is of null range
	      ASSERT false
	      REPORT " --- right input has null range "
	      SEVERITY ERROR;
              RETURN ('0');
         END IF;
	-- synopsys translate_on        
 	-- input are not null so sign extend them to the same length
	vl := SignExtend(l, resltlen, l'LEFT, SrcRegMode);
	vr := SignExtend(r, resltlen, r'LEFT, SrcRegMode);
       	return( To_StdULogic_loc( NotEqual(vl, vr)));
     END RegNotEqual; 
     -----------------------------------------------------------------------------
     FUNCTION RegNotEqual    (  CONSTANT l        : IN std_ulogic_vector;
			     CONSTANT r        : IN std_ulogic_vector;
			     CONSTANT SrcRegMode : IN regmode_type
                     -- synopsys synthesis_off
							      := DefaultRegMode 
                     -- synopsys synthesis_on
			   ) RETURN BOOLEAN IS
       CONSTANT resltlen : INTEGER := MAXIMUM (l'LENGTH, r'LENGTH);
       VARIABLE vl, vr   : STD_ULOGIC_VECTOR (resltlen - 1 DOWNTO 0);
     BEGIN
        -- synopsys translate_off
	-- Null range check
	IF ( (l'LENGTH = 0) AND (r'LENGTH = 0) ) THEN   
	      ASSERT false 
	      REPORT "  --- Both left and right vectors have null range "
	      SEVERITY ERROR;
              return( false);
         ELSIF( l'LENGTH = 0) THEN        -- left input is of null range
    	      ASSERT false
	      REPORT " --- left input has null range "
	      SEVERITY ERROR;
              return(false);

         ELSIF( r'LENGTH = 0) THEN        -- right  input is of null range
	      ASSERT false
	      REPORT " --- right input has null range "
	      SEVERITY ERROR;
              RETURN (false);
         END IF;
	-- synopsys translate_on        
 	-- input are not null so sign extend them to the same length
	vl := SignExtend(l, resltlen, l'LEFT, SrcRegMode);
	vr := SignExtend(r, resltlen, r'LEFT, SrcRegMode);
	return ( NotEqual(vl, vr));
     END RegNotEqual; 
     -- -----------------------------------------------------------------------------
     FUNCTION RegNotEqual     ( CONSTANT l          : IN std_ulogic_vector;
			     CONSTANT r          : IN INTEGER;
			     CONSTANT SrcRegMode : IN regmode_type
                     -- synopsys synthesis_off
					         	      := DefaultRegMode 
                     -- synopsys synthesis_on
			   ) RETURN BOOLEAN IS
	VARIABLE vl, vr    : std_ulogic_vector(IntegerBitLength - 1 DOWNTO 0);
     BEGIN
	-- synopsys translate_off
	-- Null range check
	 IF( l'LENGTH = 0) THEN        -- left input is of null range
    	      ASSERT false
	      REPORT " --- left input has null range "
	      SEVERITY ERROR;
              return(false);
         END IF;
	-- synopsys translate_on        
	-- input are not null so sign extend them to the same length
        -- Convert to std_ulogic_vector for comparison to allow any length input vector.
        vr := To_StdULogicVector ( r, IntegerBitLength, SrcRegMode );
 	vl := SignExtend(l, IntegerBitLength, l'LEFT, SrcRegMode);
       	return (NotEqual(vl, vr));
     END RegNotEqual; 
     -------------------------------------------------------------------------------
     FUNCTION RegNotEqual    (  CONSTANT l          : IN INTEGER;
			     CONSTANT r          : IN std_ulogic_vector;
			     CONSTANT SrcRegMode : IN regmode_type
                     -- synopsys synthesis_off
					         	      := DefaultRegMode 
                     -- synopsys synthesis_on
			   ) RETURN BOOLEAN IS
       VARIABLE vl, vr    : std_ulogic_vector(IntegerBitLength - 1 DOWNTO 0);
     BEGIN
	-- synopsys translate_off
	-- Null range check
	 IF( r'LENGTH = 0) THEN        -- right input is of null range
    	      ASSERT false
	      REPORT " --- left input has null range "
	      SEVERITY ERROR;
              return(false);
         END IF;
	-- synopsys translate_on        
	-- input are not null so sign extend them to the same length
        -- Convert to std_ulogic_vector for comparison to allow any length input vector.
        vl := To_StdULogicVector ( l, IntegerBitLength, SrcRegMode );
 	vr := SignExtend(r, IntegerBitLength, r'LEFT, SrcRegMode);
	return (NotEqual(vl, vr));
     END RegNotEqual; 
     -------------------------------------------------------------------------------
     FUNCTION RegNotEqual     ( CONSTANT l          : IN std_ulogic_vector;
			     CONSTANT r          : IN INTEGER;
			     CONSTANT SrcRegMode : IN regmode_type 
                     -- synopsys synthesis_off
					         	      := DefaultRegMode 
                     -- synopsys synthesis_on
			   ) RETURN std_ulogic IS
	VARIABLE vl, vr    : std_ulogic_vector(IntegerBitLength - 1 DOWNTO 0);
     BEGIN
	-- synopsys translate_off
	-- Null range check
	 IF( l'LENGTH = 0) THEN        -- left input is of null range
    	      ASSERT false
	      REPORT " --- left input has null range "
	      SEVERITY ERROR;
              return('0');
         END IF;
	-- synopsys translate_on        
	-- input are not null so sign extend them to the same length
        -- Convert to std_ulogic_vector for comparison to allow any length input vector.
        vr := To_StdULogicVector ( r, IntegerBitLength, SrcRegMode );
 	vl := SignExtend(l, IntegerBitLength, l'LEFT, SrcRegMode);
       	return ( To_StdULogic_loc(NotEqual(vl, vr)));
     END RegNotEqual; 
     -------------------------------------------------------------------------------
     FUNCTION RegNotEqual    (  CONSTANT l          : IN INTEGER;
			     CONSTANT r          : IN std_ulogic_vector;
			     CONSTANT SrcRegMode : IN regmode_type 
                     -- synopsys synthesis_off
					         	      := DefaultRegMode 
                     -- synopsys synthesis_on
			   ) RETURN std_ulogic IS
       VARIABLE vl, vr    : std_ulogic_vector(IntegerBitLength - 1 DOWNTO 0);
     BEGIN
	-- synopsys translate_off
	-- Null range check
	 IF( r'LENGTH = 0) THEN        -- right input is of null range
    	      ASSERT false
	      REPORT " --- left input has null range "
	      SEVERITY ERROR;
              return('0');
         END IF;
	-- synopsys translate_on        
	-- input are not null so sign extend them to the same length
        -- Convert to std_ulogic_vector for comparison to allow any length input vector.
        vl := To_StdULogicVector ( l, IntegerBitLength, SrcRegMode );
 	vr := SignExtend(r, IntegerBitLength, r'LEFT, SrcRegMode);
	return (To_StdULogic_loc(NotEqual(vl, vr)));
     END RegNotEqual; 
     -------------------------------------------------------------------------------
     --     Function Name : RegLessThan
     -- 1.2.49
     --     Overloading   : Input parameter TYPEs.
     --
     --     Purpose       : Compute a less than relation for bit_vector
     --
     --     Parameters    : l       - input bit_vector | INTEGER
     --                     r       - input bit_vector | INTEGER
     --                     SrcRegMode - input regmode_type, indicating the format of
     --                               the bit_vector operands (l,r).
     --                               Default is TwosComp.
     --
     --     Result        : BOOLEAN | bit. 
     --
     --     NOTE          : The operands may be of any length, and may be different
     --                     lengths.
     --
     --                     Overloading not defined for both inputs of INTEGER type.
     --     Use           :
     --                      VARIABLE a, b : bit_vector ( 7 DOWNTO 0 );
     --                      IF ( RegLessThan ( a, b, TwosComp)   )  THEN
     --
     --     See Also      : RegLessThanOrEqual, RegGreaterThan, RegGreaterThanOrEqual.
     -------------------------------------------------------------------------------
     FUNCTION RegLessThan  ( CONSTANT l          : IN bit_vector;
			     CONSTANT r          : IN bit_vector;
			     CONSTANT SrcRegMode : IN regmode_type
                     -- synopsys synthesis_off
						      := DefaultRegMode 
                     -- synopsys synthesis_on
			   ) RETURN bit IS
       CONSTANT resltlen : INTEGER := MAXIMUM (l'LENGTH, r'LENGTH);
       VARIABLE vl, vr   : BIT_VECTOR (resltlen - 1 DOWNTO 0);
     BEGIN
        -- synopsys translate_off
	-- Null range check
	IF ( (l'LENGTH = 0) AND (r'LENGTH = 0) ) THEN   
	      ASSERT false 
	      REPORT "  --- Both left and right vectors have null range "
	      SEVERITY ERROR;
              return( '0');
         ELSIF( l'LENGTH = 0) THEN        -- left input is of null range
    	      ASSERT false
	      REPORT " --- left input has null range "
	      SEVERITY ERROR;
              return('1');

         ELSIF( r'LENGTH = 0) THEN        -- right  input is of null range
	      ASSERT false
	      REPORT " --- right input has null range "
	      SEVERITY ERROR;
              RETURN ('0');
         END IF;
	-- synopsys translate_on        
 	-- input are not null so sign extend them to the same length
	vl := SignExtend(l, resltlen, l'LEFT, SrcRegMode);
	vr := SignExtend(r, resltlen, r'LEFT, SrcRegMode);

	IF (SrcRegMode = TwosComp) THEN
        	return( To_Bit_loc( LessThan_TwosComp(vl, vr)));
        ELSE
		return( To_Bit_loc (LessThan_Unsigned(vl, vr)));
	END IF;
     END RegLessThan; 
     -----------------------------------------------------------------------------
     FUNCTION RegLessThan (  CONSTANT l        : IN bit_vector;
			     CONSTANT r        : IN bit_vector;
			     CONSTANT SrcRegMode : IN regmode_type
                     -- synopsys synthesis_off
						      := DefaultRegMode 
                     -- synopsys synthesis_on
			   ) RETURN BOOLEAN IS

       CONSTANT resltlen : INTEGER := MAXIMUM (l'LENGTH, r'LENGTH);
       VARIABLE vl, vr   : BIT_VECTOR (resltlen - 1 DOWNTO 0);
     BEGIN
        -- synopsys translate_off
	-- Null range check
	IF ( (l'LENGTH = 0) AND (r'LENGTH = 0) ) THEN   
	      ASSERT false 
	      REPORT "  --- Both left and right vectors have null range "
	      SEVERITY ERROR;
              return( false);
         ELSIF( l'LENGTH = 0) THEN        -- left input is of null range
    	      ASSERT false
	      REPORT " --- left input has null range "
	      SEVERITY ERROR;
              return(true);

         ELSIF( r'LENGTH = 0) THEN        -- right  input is of null range
	      ASSERT false
	      REPORT " --- right input has null range "
	      SEVERITY ERROR;
              RETURN (false);
         END IF;
	-- synopsys translate_on        
 	-- input are not null so sign extend them to the same length
	vl := SignExtend(l, resltlen, l'LEFT, SrcRegMode);
	vr := SignExtend(r, resltlen, r'LEFT, SrcRegMode);

	IF (SrcRegMode = TwosComp) THEN
        	return(LessThan_TwosComp(vl, vr));
        ELSE
		return (LessThan_Unsigned(vl, vr));
	END IF;
     END RegLessThan; 
     -- -----------------------------------------------------------------------------
     FUNCTION RegLessThan  ( CONSTANT l          : IN bit_vector;
			     CONSTANT r          : IN INTEGER;
			     CONSTANT SrcRegMode : IN regmode_type
                     -- synopsys synthesis_off
						      := DefaultRegMode 
                     -- synopsys synthesis_on
			   ) RETURN BOOLEAN IS
       VARIABLE vl, vr    : bit_vector(IntegerBitLength - 1 DOWNTO 0);
     BEGIN
	-- synopsys translate_off
	-- Null range check
	 IF( l'LENGTH = 0) THEN        -- left input is of null range
    	      ASSERT false
	      REPORT " --- left input has null range "
	      SEVERITY ERROR;
              return(true);
         END IF;
	-- synopsys translate_on        
	-- input are not null so sign extend them to the same length
        -- Convert to bit_vector for comparison to allow any length input vector.
        vr := To_BitVector ( r, IntegerBitLength, SrcRegMode );
 	vl := SignExtend(l, IntegerBitLength, l'LEFT, SrcRegMode);
	IF (SrcRegMode = TwosComp) THEN
        	return(LessThan_TwosComp(vl, vr));
        ELSE
		return (LessThan_Unsigned(vl, vr));
	END IF;
     END RegLessThan; 
     -------------------------------------------------------------------------------
     FUNCTION RegLessThan (  CONSTANT l          : IN INTEGER;
			     CONSTANT r          : IN bit_vector;
			     CONSTANT SrcRegMode : IN regmode_type
                     -- synopsys synthesis_off
						      := DefaultRegMode 
                     -- synopsys synthesis_on
			   ) RETURN BOOLEAN IS
       VARIABLE vl, vr    : bit_vector(IntegerBitLength - 1 DOWNTO 0);
     BEGIN
	-- synopsys translate_off
	-- Null range check
	 IF( r'LENGTH = 0) THEN        -- right input is of null range
    	      ASSERT false
	      REPORT " --- left input has null range "
	      SEVERITY ERROR;
              return(false);
         END IF;
	-- synopsys translate_on        
	-- input are not null so sign extend them to the same length
        -- Convert to bit_vector for comparison to allow any length input vector.
        vl := To_BitVector ( l, IntegerBitLength, SrcRegMode );
 	vr := SignExtend(r, IntegerBitLength, r'LEFT, SrcRegMode);
	IF (SrcRegMode = TwosComp) THEN
        	return(LessThan_TwosComp(vl, vr));
        ELSE
		return (LessThan_Unsigned(vl, vr));
	END IF;
     END RegLessThan; 
     -------------------------------------------------------------------------------
     FUNCTION RegLessThan  ( CONSTANT l          : IN bit_vector;
			     CONSTANT r          : IN INTEGER;
			     CONSTANT SrcRegMode : IN regmode_type
                     -- synopsys synthesis_off
						      := DefaultRegMode 
                     -- synopsys synthesis_on
			   ) RETURN bit IS
       VARIABLE vl, vr    : bit_vector(IntegerBitLength - 1 DOWNTO 0);
     BEGIN
        -- synopsys translate_off
	-- Null range check
         IF( l'LENGTH = 0) THEN        -- left input is of null range
    	      ASSERT false
	      REPORT " --- left input has null range "
	      SEVERITY ERROR;
              return('1');
         END IF;
	-- synopsys translate_on        
	-- input are not null so sign extend them to the same length
        -- Convert to bit_vector for comparison to allow any length input vector.
 	vl := SignExtend(l, IntegerBitLength, l'LEFT, SrcRegMode);
        vr := To_BitVector ( r, IntegerBitLength, SrcRegMode );

	IF (SrcRegMode = TwosComp) THEN
        	return( To_Bit_loc( LessThan_TwosComp(vl, vr)));
        ELSE
		return( To_Bit_loc (LessThan_Unsigned(vl, vr)));
	END IF;
    END RegLessThan; 
     -------------------------------------------------------------------------------
     FUNCTION RegLessThan (  CONSTANT l          : IN INTEGER;
			     CONSTANT r          : IN bit_vector;
			     CONSTANT SrcRegMode : IN regmode_type
                     -- synopsys synthesis_off
						      := DefaultRegMode 
                     -- synopsys synthesis_on
			   ) RETURN bit IS
       VARIABLE vl, vr    : bit_vector(IntegerBitLength - 1 DOWNTO 0);
     BEGIN
        -- synopsys translate_off
	-- Null range check
         IF( r'LENGTH = 0) THEN        -- left input is of null range
    	      ASSERT false
	      REPORT " --- left input has null range "
	      SEVERITY ERROR;
              return('0');
         END IF;
	-- synopsys translate_on        
	-- input are not null so sign extend them to the same length
        -- Convert to bit_vector for comparison to allow any length input vector.
        vl := To_BitVector ( l, IntegerBitLength, SrcRegMode );
 	vr := SignExtend(r, IntegerBitLength, r'LEFT, SrcRegMode);

	IF (SrcRegMode = TwosComp) THEN
        	return( To_Bit_loc( LessThan_TwosComp(vl, vr)));
        ELSE
		return( To_Bit_loc (LessThan_Unsigned(vl, vr)));
	END IF;
    END RegLessThan; 
     -------------------------------------------------------------------------------
     --     Function Name : RegLessThan
     --
     --     Overloading   : Input parameter TYPEs.
     --    
     --     Purpose       : Compute a less than relation for std_logic_vectors
     --     
     --     Parameters    : l       - input std_logic_vector | INTEGER
     --                     r       - input std_logic_vector | INTEGER
     --                     SrcRegMode - input regmode_type, indicating the format of
     --                               the std_logic_vector operands (l,r).
     --                               Default is TwosComp.
     --     
     --     Result        : BOOLEAN | std_ulogic
     --
     --     NOTE          : The operands may be of any length, and may be different
     --                     lengths. 
     --
     --                     Overloading not defined for both inputs of INTEGER type.
     --
     --                     Any time the comparison reaches an index that has an 'X' as an
     --                     array element, the comparison is deemed indeterminate and will 
     --                     return false in case of boolean and '0' incase of 
     --                     std_ulogic for synthesis purposes.
     --
     --     Use           : 
     --                      VARIABLE a, b : std_logic_vector ( 7 DOWNTO 0 );
     --                      IF ( RegLessThan ( a, b, TwosComp)   )  THEN 
     --     
     --     See Also      : RegLessThanOrEqual,RegGreaterThan,RegGreaterThanOrEqual.
     -------------------------------------------------------------------------------
     FUNCTION RegLessThan  ( CONSTANT l          : IN std_logic_vector;
			     CONSTANT r          : IN std_logic_vector;
			     CONSTANT SrcRegMode : IN regmode_type
                     -- synopsys synthesis_off
						      := DefaultRegMode 
                     -- synopsys synthesis_on
			   ) RETURN std_ulogic IS
       CONSTANT resltlen : INTEGER := MAXIMUM (l'LENGTH, r'LENGTH);
       VARIABLE vl, vr   : STD_LOGIC_VECTOR (resltlen - 1 DOWNTO 0);
     BEGIN
        -- synopsys translate_off
	-- Null range check
	IF ( (l'LENGTH = 0) AND (r'LENGTH = 0) ) THEN   
	      ASSERT false 
	      REPORT "  --- Both left and right vectors have null range "
	      SEVERITY ERROR;
              return( '0');
         ELSIF( l'LENGTH = 0) THEN        -- left input is of null range
    	      ASSERT false
	      REPORT " --- left input has null range "
	      SEVERITY ERROR;
              return('1');

         ELSIF( r'LENGTH = 0) THEN        -- right  input is of null range
	      ASSERT false
	      REPORT " --- right input has null range "
	      SEVERITY ERROR;
              RETURN ('0');
         END IF;
	-- synopsys translate_on        
 	-- input are not null so sign extend them to the same length
	vl := SignExtend(l, resltlen, l'LEFT, SrcRegMode);
	vr := SignExtend(r, resltlen, r'LEFT, SrcRegMode);

	IF (SrcRegMode = TwosComp) THEN
        	return( To_StdULogic_loc( LessThan_TwosComp(vl, vr)));
        ELSE
		return( To_StdULogic_loc(LessThan_Unsigned(vl, vr)));
	END IF;
     END RegLessThan; 
     -----------------------------------------------------------------------------
     FUNCTION RegLessThan (  CONSTANT l        : IN std_logic_vector;
			     CONSTANT r        : IN std_logic_vector;
			     CONSTANT SrcRegMode : IN regmode_type
                     -- synopsys synthesis_off
						      := DefaultRegMode 
                     -- synopsys synthesis_on
			   ) RETURN BOOLEAN IS

       CONSTANT resltlen : INTEGER := MAXIMUM (l'LENGTH, r'LENGTH);
       VARIABLE vl, vr   : STD_LOGIC_VECTOR (resltlen - 1 DOWNTO 0);
     BEGIN
        -- synopsys translate_off
	-- Null range check
	IF ( (l'LENGTH = 0) AND (r'LENGTH = 0) ) THEN   
	      ASSERT false 
	      REPORT "  --- Both left and right vectors have null range "
	      SEVERITY ERROR;
              return( false);
         ELSIF( l'LENGTH = 0) THEN        -- left input is of null range
    	      ASSERT false
	      REPORT " --- left input has null range "
	      SEVERITY ERROR;
              return(true);

         ELSIF( r'LENGTH = 0) THEN        -- right  input is of null range
	      ASSERT false
	      REPORT " --- right input has null range "
	      SEVERITY ERROR;
              RETURN (false);
         END IF;
	-- synopsys translate_on        
 	-- input are not null so sign extend them to the same length
	vl := SignExtend(l, resltlen, l'LEFT, SrcRegMode);
	vr := SignExtend(r, resltlen, r'LEFT, SrcRegMode);

	IF (SrcRegMode = TwosComp) THEN
        	return(LessThan_TwosComp(vl, vr));
        ELSE
		return (LessThan_Unsigned(vl, vr));
	END IF;
     END RegLessThan; 
     -- -----------------------------------------------------------------------------
     FUNCTION RegLessThan  ( CONSTANT l          : IN std_logic_vector;
			     CONSTANT r          : IN INTEGER;
			     CONSTANT SrcRegMode : IN regmode_type
                     -- synopsys synthesis_off
						      := DefaultRegMode 
                     -- synopsys synthesis_on
			   ) RETURN BOOLEAN IS
       VARIABLE vl, vr    : std_logic_vector(IntegerBitLength - 1 DOWNTO 0);
     BEGIN
	-- synopsys translate_off
	-- Null range check
	 IF( l'LENGTH = 0) THEN        -- left input is of null range
    	      ASSERT false
	      REPORT " --- left input has null range "
	      SEVERITY ERROR;
              return(true);
         END IF;
	-- synopsys translate_on        
	-- input are not null so sign extend them to the same length
        -- Convert to std_logic_vector for comparison to allow any length input vector.
        vr := To_StdLogicVector ( r, IntegerBitLength, SrcRegMode );
 	vl := SignExtend(l, IntegerBitLength, l'LEFT, SrcRegMode);
	IF (SrcRegMode = TwosComp) THEN
        	return(LessThan_TwosComp(vl, vr));
        ELSE
		return (LessThan_Unsigned(vl, vr));
	END IF;
     END RegLessThan; 
     -------------------------------------------------------------------------------
     FUNCTION RegLessThan (  CONSTANT l          : IN INTEGER;
			     CONSTANT r          : IN std_logic_vector;
			     CONSTANT SrcRegMode : IN regmode_type
                     -- synopsys synthesis_off
						      := DefaultRegMode 
                     -- synopsys synthesis_on
			   ) RETURN BOOLEAN IS
       VARIABLE vl, vr    : std_logic_vector(IntegerBitLength - 1 DOWNTO 0);
     BEGIN
	-- synopsys translate_off
	-- Null range check
	 IF( r'LENGTH = 0) THEN        -- right input is of null range
    	      ASSERT false
	      REPORT " --- left input has null range "
	      SEVERITY ERROR;
              return(false);
         END IF;
	-- synopsys translate_on        
	-- input are not null so sign extend them to the same length
        -- Convert to std_logic_vector for comparison to allow any length input vector.
        vl := To_StdLogicVector ( l, IntegerBitLength, SrcRegMode );
 	vr := SignExtend(r, IntegerBitLength, r'LEFT, SrcRegMode);
	IF (SrcRegMode = TwosComp) THEN
        	return(LessThan_TwosComp(vl, vr));
        ELSE
		return (LessThan_Unsigned(vl, vr));
	END IF;
     END RegLessThan; 
     -------------------------------------------------------------------------------
     FUNCTION RegLessThan  ( CONSTANT l          : IN std_logic_vector;
			     CONSTANT r          : IN INTEGER;
			     CONSTANT SrcRegMode : IN regmode_type
                     -- synopsys synthesis_off
						      := DefaultRegMode 
                     -- synopsys synthesis_on
			   ) RETURN std_ulogic IS
       VARIABLE vl, vr    : std_logic_vector(IntegerBitLength - 1 DOWNTO 0);
     BEGIN
        -- synopsys translate_off
	-- Null range check
         IF( l'LENGTH = 0) THEN        -- left input is of null range
    	      ASSERT false
	      REPORT " --- left input has null range "
	      SEVERITY ERROR;
              return('1');
         END IF;
	-- synopsys translate_on        
	-- input are not null so sign extend them to the same length
        -- Convert to std_logic_vector for comparison to allow any length input vector.
 	vl := SignExtend(l, IntegerBitLength, l'LEFT, SrcRegMode);
        vr := To_StdLogicVector ( r, IntegerBitLength, SrcRegMode );

	IF (SrcRegMode = TwosComp) THEN
        	return( To_StdULogic_loc( LessThan_TwosComp(vl, vr)));
        ELSE
		return( To_StdULogic_loc (LessThan_Unsigned(vl, vr)));
	END IF;
     END RegLessThan; 
     -------------------------------------------------------------------------------
     FUNCTION RegLessThan (  CONSTANT l          : IN INTEGER;
			     CONSTANT r          : IN std_logic_vector;
			     CONSTANT SrcRegMode : IN regmode_type
                     -- synopsys synthesis_off
						      := DefaultRegMode 
                     -- synopsys synthesis_on
			   ) RETURN std_ulogic IS
       VARIABLE vl, vr    : std_logic_vector(IntegerBitLength - 1 DOWNTO 0);
     BEGIN
        -- synopsys translate_off
	-- Null range check
         IF( r'LENGTH = 0) THEN        -- left input is of null range
    	      ASSERT false
	      REPORT " --- left input has null range "
	      SEVERITY ERROR;
              return('0');
         END IF;
	-- synopsys translate_on        
	-- input are not null so sign extend them to the same length
        -- Convert to std_logic_vector for comparison to allow any length input vector.
        vl := To_StdLogicVector ( l, IntegerBitLength, SrcRegMode );
 	vr := SignExtend(r, IntegerBitLength, r'LEFT, SrcRegMode);

	IF (SrcRegMode = TwosComp) THEN
        	return( To_StdULogic_loc( LessThan_TwosComp(vl, vr)));
        ELSE
		return( To_StdULogic_loc (LessThan_Unsigned(vl, vr)));
	END IF;
     END RegLessThan; 
     -------------------------------------------------------------------------------
     --     Function Name : RegLessThan
     --
     --     Overloading   : Input parameter TYPEs.
     --    
     --     Purpose       : Compute a less than relation for std_ulogic_vectors
     --     
     --     Parameters    : l       - input std_ulogic_vector | INTEGER
     --                     r       - input std_ulogic_vector | INTEGER
     --                     SrcRegMode - input regmode_type, indicating the format of
     --                               the std_ulogic_vector operands (l,r).
     --                               Default is TwosComp.
     --     
     --     Result        : BOOLEAN | std_ulogic
     --
     --     NOTE          : The operands may be of any length, and may be different
     --                     lengths. 
     --
     --                     Overloading not defined for both inputs of INTEGER type.
     --
     --                     Any time the comparison reaches an index that has an 'X' as an
     --                     array element, the comparison is deemed indeterminate and will 
     --                     return false in case of boolean and '0' incase of 
     --                     std_ulogic for synthesis purposes.
     --     Use           : 
     --                      VARIABLE a, b : std_ulogic_vector ( 7 DOWNTO 0 );
     --                      IF ( RegLessThan ( a, b, TwosComp)   )  THEN 
     --     
     --     See Also      : RegLessThanOrEqual, RegGreaterThan, RegGreaterThanOrEqual.
     -------------------------------------------------------------------------------
     FUNCTION RegLessThan  ( CONSTANT l          : IN std_ulogic_vector;
			     CONSTANT r          : IN std_ulogic_vector;
			     CONSTANT SrcRegMode : IN regmode_type
                     -- synopsys synthesis_off
						      := DefaultRegMode 
                     -- synopsys synthesis_on
			   ) RETURN std_ulogic IS
       CONSTANT resltlen : INTEGER := MAXIMUM (l'LENGTH, r'LENGTH);
       VARIABLE vl, vr   : STD_ULOGIC_VECTOR (resltlen - 1 DOWNTO 0);
     BEGIN
        -- synopsys translate_off
	-- Null range check
	IF ( (l'LENGTH = 0) AND (r'LENGTH = 0) ) THEN   
	      ASSERT false 
	      REPORT "  --- Both left and right vectors have null range "
	      SEVERITY ERROR;
              return( '0');
         ELSIF( l'LENGTH = 0) THEN        -- left input is of null range
    	      ASSERT false
	      REPORT " --- left input has null range "
	      SEVERITY ERROR;
              return('1');

         ELSIF( r'LENGTH = 0) THEN        -- right  input is of null range
	      ASSERT false
	      REPORT " --- right input has null range "
	      SEVERITY ERROR;
              RETURN ('0');
         END IF;
	-- synopsys translate_on        
 	-- input are not null so sign extend them to the same length
	vl := SignExtend(l, resltlen, l'LEFT, SrcRegMode);
	vr := SignExtend(r, resltlen, r'LEFT, SrcRegMode);

	IF (SrcRegMode = TwosComp) THEN
        	return( To_StdULogic_loc( LessThan_TwosComp(vl, vr)));
        ELSE
		return( To_StdULogic_loc(LessThan_Unsigned(vl, vr)));
	END IF;
      END RegLessThan; 
     -----------------------------------------------------------------------------
     FUNCTION RegLessThan (  CONSTANT l        : IN std_ulogic_vector;
			     CONSTANT r        : IN std_ulogic_vector;
			     CONSTANT SrcRegMode : IN regmode_type
                     -- synopsys synthesis_off
						      := DefaultRegMode 
                     -- synopsys synthesis_on
			   ) RETURN BOOLEAN IS
       CONSTANT resltlen : INTEGER := MAXIMUM (l'LENGTH, r'LENGTH);
       VARIABLE vl, vr   : STD_ULOGIC_VECTOR (resltlen - 1 DOWNTO 0);
     BEGIN
        -- synopsys translate_off
	-- Null range check
	IF ( (l'LENGTH = 0) AND (r'LENGTH = 0) ) THEN   
	      ASSERT false 
	      REPORT "  --- Both left and right vectors have null range "
	      SEVERITY ERROR;
              return( false);
         ELSIF( l'LENGTH = 0) THEN        -- left input is of null range
    	      ASSERT false
	      REPORT " --- left input has null range "
	      SEVERITY ERROR;
              return(true);

         ELSIF( r'LENGTH = 0) THEN        -- right  input is of null range
	      ASSERT false
	      REPORT " --- right input has null range "
	      SEVERITY ERROR;
              RETURN (false);
         END IF;
	-- synopsys translate_on        
 	-- input are not null so sign extend them to the same length
	vl := SignExtend(l, resltlen, l'LEFT, SrcRegMode);
	vr := SignExtend(r, resltlen, r'LEFT, SrcRegMode);

	IF (SrcRegMode = TwosComp) THEN
        	return(LessThan_TwosComp(vl, vr));
        ELSE
		return (LessThan_Unsigned(vl, vr));
	END IF;
    END RegLessThan; 
     -- -----------------------------------------------------------------------------
     FUNCTION RegLessThan  ( CONSTANT l          : IN std_ulogic_vector;
			     CONSTANT r          : IN INTEGER;
			     CONSTANT SrcRegMode : IN regmode_type
                     -- synopsys synthesis_off
						      := DefaultRegMode 
                     -- synopsys synthesis_on
			   ) RETURN BOOLEAN IS
       VARIABLE vl, vr    : std_ulogic_vector(IntegerBitLength - 1 DOWNTO 0);
     BEGIN
	-- synopsys translate_off
	-- Null range check
	 IF( l'LENGTH = 0) THEN        -- left input is of null range
    	      ASSERT false
	      REPORT " --- left input has null range "
	      SEVERITY ERROR;
              return(true);
         END IF;
	-- synopsys translate_on        
	-- input are not null so sign extend them to the same length
        -- Convert to std_ulogic_vector for comparison to allow any length input vector.
        vr := To_StdULogicVector ( r, IntegerBitLength, SrcRegMode );
 	vl := SignExtend(l, IntegerBitLength, l'LEFT, SrcRegMode);
	IF (SrcRegMode = TwosComp) THEN
        	return(LessThan_TwosComp(vl, vr));
        ELSE
		return (LessThan_Unsigned(vl, vr));
	END IF;
     END RegLessThan; 
     -------------------------------------------------------------------------------
     FUNCTION RegLessThan (  CONSTANT l          : IN INTEGER;
			     CONSTANT r          : IN std_ulogic_vector;
			     CONSTANT SrcRegMode : IN regmode_type
                     -- synopsys synthesis_off
						      := DefaultRegMode 
                     -- synopsys synthesis_on
			   ) RETURN BOOLEAN IS
       VARIABLE vl, vr    : std_ulogic_vector(IntegerBitLength - 1 DOWNTO 0);
     BEGIN
	-- synopsys translate_off
	-- Null range check
	 IF( r'LENGTH = 0) THEN        -- right input is of null range
    	      ASSERT false
	      REPORT " --- left input has null range "
	      SEVERITY ERROR;
              return(false);
         END IF;
	-- synopsys translate_on        
	-- input are not null so sign extend them to the same length
        -- Convert to std_ulogic_vector for comparison to allow any length input vector.
        vl := To_StdULogicVector ( l, IntegerBitLength, SrcRegMode );
 	vr := SignExtend(r, IntegerBitLength, r'LEFT, SrcRegMode);
	IF (SrcRegMode = TwosComp) THEN
        	return(LessThan_TwosComp(vl, vr));
        ELSE
		return (LessThan_Unsigned(vl, vr));
	END IF;
     END RegLessThan; 
     -------------------------------------------------------------------------------
     FUNCTION RegLessThan  ( CONSTANT l          : IN std_ulogic_vector;
			     CONSTANT r          : IN INTEGER;
			     CONSTANT SrcRegMode : IN regmode_type
                     -- synopsys synthesis_off
						      := DefaultRegMode 
                     -- synopsys synthesis_on
			   ) RETURN std_ulogic IS
       VARIABLE vl, vr    : std_ulogic_vector(IntegerBitLength - 1 DOWNTO 0);
     BEGIN
        -- synopsys translate_off
	-- Null range check
         IF( l'LENGTH = 0) THEN        -- left input is of null range
    	      ASSERT false
	      REPORT " --- left input has null range "
	      SEVERITY ERROR;
              return('1');
         END IF;
	-- synopsys translate_on        
	-- input are not null so sign extend them to the same length
        -- Convert to std_ulogic_vector for comparison to allow any length input vector.
 	vl := SignExtend(l, IntegerBitLength, l'LEFT, SrcRegMode);
        vr := To_StdULogicVector ( r, IntegerBitLength, SrcRegMode );

	IF (SrcRegMode = TwosComp) THEN
        	return( To_StdULogic_loc( LessThan_TwosComp(vl, vr)));
        ELSE
		return( To_StdULogic_loc (LessThan_Unsigned(vl, vr)));
	END IF;
     END RegLessThan; 
     -------------------------------------------------------------------------------
     FUNCTION RegLessThan (  CONSTANT l          : IN INTEGER;
			     CONSTANT r          : IN std_ulogic_vector;
			     CONSTANT SrcRegMode : IN regmode_type
                     -- synopsys synthesis_off
						      := DefaultRegMode 
                     -- synopsys synthesis_on
			   ) RETURN std_ulogic IS
       VARIABLE vl, vr    : std_ulogic_vector(IntegerBitLength - 1 DOWNTO 0);
     BEGIN
        -- synopsys translate_off
	-- Null range check
         IF( r'LENGTH = 0) THEN        -- left input is of null range
    	      ASSERT false
	      REPORT " --- left input has null range "
	      SEVERITY ERROR;
              return('0');
         END IF;
	-- synopsys translate_on        
	-- input are not null so sign extend them to the same length
        -- Convert to std_ulogic_vector for comparison to allow any length input vector.
        vl := To_StdULogicVector (l, IntegerBitLength, SrcRegMode );
 	vr := SignExtend(r, IntegerBitLength, r'LEFT, SrcRegMode);

	IF (SrcRegMode = TwosComp) THEN
        	return( To_StdULogic_loc( LessThan_TwosComp(vl, vr)));
        ELSE
		return( To_StdULogic_loc (LessThan_Unsigned(vl, vr)));
	END IF;
     END RegLessThan; 
     -------------------------------------------------------------------------------
     --     Function Name : RegLessThanOrEqual
     -- 1.2.51
     --     Overloading   : Input parameter TYPEs.
     --
     --     Purpose       : Compute a less than or equal relation for bit_vectors
     --
     --     Parameters    : l       - input bit_vector | INTEGER
     --                     r       - input bit_vector | INTEGER
     --                     SrcRegMode - input regmode_type, indicating the format of
     --                               the bit_vector operands (l,r).
     --                               Default is TwosComp.
     --
     --     Result        : BOOLEAN | bit
     --
     --     NOTE          : The operands may be of any length, and may be different
     --                     lengths.
     --
     --                     Overloading not defined for both inputs of INTEGER type.
     --     Use           :
     --                      VARIABLE a, b : bit_vector ( 7 DOWNTO 0 );
     --                      IF ( RegLessThanOrEqual ( a, b, TwosComp)   )  THEN
     --
     --     See Also      : RegLessThan, RegGreaterThan, RegGreaterThanOrEqual.
     -------------------------------------------------------------------------------
     FUNCTION RegLessThanOrEqual ( CONSTANT l          : IN bit_vector;
				   CONSTANT r          : IN bit_vector;
				   CONSTANT SrcRegMode : IN regmode_type
                     -- synopsys synthesis_off
							      := DefaultRegMode 
                     -- synopsys synthesis_on
				 ) RETURN bit IS
       CONSTANT resltlen : INTEGER := MAXIMUM (l'LENGTH, r'LENGTH);
       VARIABLE vl, vr   : BIT_VECTOR (resltlen - 1 DOWNTO 0);
     BEGIN
        -- synopsys translate_off
	-- Null range check
	IF ( (l'LENGTH = 0) AND (r'LENGTH = 0) ) THEN   
	      ASSERT false 
	      REPORT "  --- Both left and right vectors have null range "
	      SEVERITY ERROR;
              return( '0');
         ELSIF( l'LENGTH = 0) THEN        -- left input is of null range
    	      ASSERT false
	      REPORT " --- left input has null range "
	      SEVERITY ERROR;
              return('1');

         ELSIF( r'LENGTH = 0) THEN        -- right  input is of null range
	      ASSERT false
	      REPORT " --- right input has null range "
	      SEVERITY ERROR;
              RETURN ('0');
         END IF;
	-- synopsys translate_on        
 	-- input are not null so sign extend them to the same length
	vl := SignExtend(l, resltlen, l'LEFT, SrcRegMode);
	vr := SignExtend(r, resltlen, r'LEFT, SrcRegMode);

	IF (SrcRegMode = TwosComp) THEN
        	return( To_Bit_loc( LessThanOrEqual_TwosComp(vl, vr)));
        ELSE
		return( To_Bit_loc (LessThanOrEqual_Unsigned(vl, vr)));
	END IF;
     END RegLessThanOrEqual; 
     -----------------------------------------------------------------------------
     FUNCTION RegLessThanOrEqual ( CONSTANT l          : IN bit_vector;
				   CONSTANT r          : IN bit_vector;
 			           CONSTANT SrcRegMode : IN regmode_type
                     -- synopsys synthesis_off
							      := DefaultRegMode 
                     -- synopsys synthesis_on
				 ) RETURN BOOLEAN IS
       CONSTANT resltlen : INTEGER := MAXIMUM (l'LENGTH, r'LENGTH);
       VARIABLE vl, vr   : BIT_VECTOR (resltlen - 1 DOWNTO 0);
     BEGIN
        -- synopsys translate_off
	-- Null range check
	IF ( (l'LENGTH = 0) AND (r'LENGTH = 0) ) THEN   
	      ASSERT false 
	      REPORT "  --- Both left and right vectors have null range "
	      SEVERITY ERROR;
              return( false);
         ELSIF( l'LENGTH = 0) THEN        -- left input is of null range
    	      ASSERT false
	      REPORT " --- left input has null range "
	      SEVERITY ERROR;
              return(true);

         ELSIF( r'LENGTH = 0) THEN        -- right  input is of null range
	      ASSERT false
	      REPORT " --- right input has null range "
	      SEVERITY ERROR;
              RETURN (false);
         END IF;
	-- synopsys translate_on        
 	-- input are not null so sign extend them to the same length
	vl := SignExtend(l, resltlen, l'LEFT, SrcRegMode);
	vr := SignExtend(r, resltlen, r'LEFT, SrcRegMode);

	IF (SrcRegMode = TwosComp) THEN
        	return ( LessThanOrEqual_TwosComp(vl, vr));
        ELSE
		return ( LessThanOrEqual_Unsigned(vl, vr));
	END IF;
     END RegLessThanOrEqual; 
     -- -----------------------------------------------------------------------------
     FUNCTION RegLessThanOrEqual ( CONSTANT l          : IN bit_vector;
				   CONSTANT r          : IN INTEGER;
			     CONSTANT SrcRegMode : IN regmode_type
                     -- synopsys synthesis_off
						      := DefaultRegMode 
                     -- synopsys synthesis_on
				 ) RETURN BOOLEAN IS
	VARIABLE vl, vr    : bit_vector(IntegerBitLength - 1 DOWNTO 0);
     BEGIN
	-- synopsys translate_off
	-- Null range check
	 IF( l'LENGTH = 0) THEN        -- left input is of null range
    	      ASSERT false
	      REPORT " --- left input has null range "
	      SEVERITY ERROR;
              return(true);
         END IF;
	-- synopsys translate_on        
	-- input are not null so sign extend them to the same length
        -- Convert to bit_vector for comparison to allow any length input vector.
        vr := To_BitVector ( r, IntegerBitLength, SrcRegMode );
 	vl := SignExtend(l, IntegerBitLength, l'LEFT, SrcRegMode);
	IF (SrcRegMode = TwosComp) THEN
        	return(LessThanOrEqual_TwosComp(vl, vr));
        ELSE
		return (LessThanOrEqual_Unsigned(vl, vr));
	END IF;
     END RegLessThanOrEqual; 
     -------------------------------------------------------------------------------
     FUNCTION RegLessThanOrEqual ( CONSTANT l          : IN INTEGER;
				   CONSTANT r          : IN bit_vector;
  			           CONSTANT SrcRegMode : IN regmode_type
                     -- synopsys synthesis_off
					         	      := DefaultRegMode 
                     -- synopsys synthesis_on
				 ) RETURN BOOLEAN IS
       VARIABLE vl, vr    : bit_vector(IntegerBitLength - 1 DOWNTO 0);
     BEGIN
	-- synopsys translate_off
	-- Null range check
	 IF( r'LENGTH = 0) THEN        -- right input is of null range
    	      ASSERT false
	      REPORT " --- left input has null range "
	      SEVERITY ERROR;
              return(false);
         END IF;
	-- synopsys translate_on        
	-- input are not null so sign extend them to the same length
        -- Convert to bit_vector for comparison to allow any length input vector.
        vl := To_BitVector ( l, IntegerBitLength, SrcRegMode );
 	vr := SignExtend(r, IntegerBitLength, r'LEFT, SrcRegMode);
	IF (SrcRegMode = TwosComp) THEN
        	return(LessThanOrEqual_TwosComp(vl, vr));
        ELSE
		return (LessThanOrEqual_Unsigned(vl, vr));
	END IF;
     END RegLessThanOrEqual; 
     -------------------------------------------------------------------------------
     FUNCTION RegLessThanOrEqual ( CONSTANT l          : IN bit_vector;
				   CONSTANT r          : IN INTEGER;
  			           CONSTANT SrcRegMode : IN regmode_type
                     -- synopsys synthesis_off
					         	      := DefaultRegMode 
                     -- synopsys synthesis_on
				 ) RETURN bit IS
       VARIABLE vl, vr    : bit_vector(IntegerBitLength - 1 DOWNTO 0);
     BEGIN
        -- synopsys translate_off
	-- Null range check
         IF( l'LENGTH = 0) THEN        -- left input is of null range
    	      ASSERT false
	      REPORT " --- left input has null range "
	      SEVERITY ERROR;
              return('1');
         END IF;
	-- synopsys translate_on        
	-- input are not null so sign extend them to the same length
        -- Convert to bit_vector for comparison to allow any length input vector.
 	vl := SignExtend(l, IntegerBitLength, l'LEFT, SrcRegMode);
        vr := To_BitVector ( r, IntegerBitLength, SrcRegMode );

	IF (SrcRegMode = TwosComp) THEN
        	return( To_Bit_loc( LessThanOrEqual_TwosComp(vl, vr)));
        ELSE
		return( To_Bit_loc (LessThanOrEqual_Unsigned(vl, vr)));
	END IF;
     END RegLessThanOrEqual; 
     -------------------------------------------------------------------------------
     FUNCTION RegLessThanOrEqual ( CONSTANT l          : IN INTEGER;
				   CONSTANT r          : IN bit_vector;
  			           CONSTANT SrcRegMode : IN regmode_type
                     -- synopsys synthesis_off
					         	      := DefaultRegMode 
                     -- synopsys synthesis_on
				 ) RETURN bit IS
       VARIABLE vl, vr    : bit_vector(IntegerBitLength - 1 DOWNTO 0);
     BEGIN
        -- synopsys translate_off
	-- Null range check
         IF( r'LENGTH = 0) THEN        -- left input is of null range
    	      ASSERT false
	      REPORT " --- left input has null range "
	      SEVERITY ERROR;
              return('0');
         END IF;
	-- synopsys translate_on        
	-- input are not null so sign extend them to the same length
        -- Convert to bit_vector for comparison to allow any length input vector.
        vl := To_BitVector ( l, IntegerBitLength, SrcRegMode );
 	vr := SignExtend(r, IntegerBitLength, r'LEFT, SrcRegMode);

	IF (SrcRegMode = TwosComp) THEN
        	return( To_Bit_loc( LessThanOrEqual_TwosComp(vl, vr)));
        ELSE
		return( To_Bit_loc (LessThanOrEqual_Unsigned(vl, vr)));
	END IF;
     END RegLessThanOrEqual; 
     -- ----------------------------------------------------------------------------
     --     Function Name : RegLessThanOrEqual
     --    
     --     Purpose       : Compute a less than or equal relation for std_logic_vectors
     --     
     --     Parameters    : l       - input std_logic_vector | INTEGER
     --                     r       - input std_logic_vector | INTEGER
     --                     SrcRegMode - input regmode_type, indicating the format of
     --                               the std_logic_vector operands (l,r).
     --                               Default is TwosComp.
     --     
     --     Result        : BOOLEAN | std_ulogic
     --
     --     NOTE          : The operands may be of any length, and may be different
     --                     lengths. 
     --
     --                     Overloading not defined for both inputs of INTEGER type.
     --
     --                     Any time the comparison reaches an index that has an 'X' as an
     --                     array element, the comparison is deemed indeterminate and will 
     --                     return false in case of boolean and '0' incase of 
     --                     std_ulogic for synthesis purposes.
     --     Use           : 
     --                      VARIABLE a, b : std_logic_vector ( 7 DOWNTO 0 );
     --                      IF ( RegLessThanOrEqual ( a, b, TwosComp)   )  THEN 
     --     
     --     See Also      : RegLessThan, RegGreaterThan, RegGreaterThanOrEqual.
     -------------------------------------------------------------------------------
     FUNCTION RegLessThanOrEqual ( CONSTANT l          : IN std_logic_vector;
				   CONSTANT r          : IN std_logic_vector;
  			           CONSTANT SrcRegMode : IN regmode_type
                     -- synopsys synthesis_off
					         	      := DefaultRegMode 
                     -- synopsys synthesis_on
				 ) RETURN std_ulogic IS
       CONSTANT resltlen : INTEGER := MAXIMUM (l'LENGTH, r'LENGTH);
       VARIABLE vl, vr   : STD_LOGIC_VECTOR (resltlen - 1 DOWNTO 0);
     BEGIN
        -- synopsys translate_off
	-- Null range check
	IF ( (l'LENGTH = 0) AND (r'LENGTH = 0) ) THEN   
	      ASSERT false 
	      REPORT "  --- Both left and right vectors have null range "
	      SEVERITY ERROR;
              return( '0');
         ELSIF( l'LENGTH = 0) THEN        -- left input is of null range
    	      ASSERT false
	      REPORT " --- left input has null range "
	      SEVERITY ERROR;
              return('1');

         ELSIF( r'LENGTH = 0) THEN        -- right  input is of null range
	      ASSERT false
	      REPORT " --- right input has null range "
	      SEVERITY ERROR;
              RETURN ('0');
         END IF;
	-- synopsys translate_on        
 	-- input are not null so sign extend them to the same length
	vl := SignExtend(l, resltlen, l'LEFT, SrcRegMode);
	vr := SignExtend(r, resltlen, r'LEFT, SrcRegMode);

	IF (SrcRegMode = TwosComp) THEN
        	return( To_StdULogic_loc( LessThanOrEqual_TwosComp(vl, vr)));
        ELSE
		return( To_StdULogic_loc(LessThanOrEqual_Unsigned(vl, vr)));
	END IF;
     END RegLessThanOrEqual; 
     -----------------------------------------------------------------------------
     FUNCTION RegLessThanOrEqual ( CONSTANT l          : IN std_logic_vector;
				   CONSTANT r          : IN std_logic_vector;
 			           CONSTANT SrcRegMode : IN regmode_type
                     -- synopsys synthesis_off
							      := DefaultRegMode 
                     -- synopsys synthesis_on
				 ) RETURN BOOLEAN IS
       CONSTANT resltlen : INTEGER := MAXIMUM (l'LENGTH, r'LENGTH);
       VARIABLE vl, vr   : STD_LOGIC_VECTOR (resltlen - 1 DOWNTO 0);
     BEGIN
        -- synopsys translate_off
	-- Null range check
	IF ( (l'LENGTH = 0) AND (r'LENGTH = 0) ) THEN   
	      ASSERT false 
	      REPORT "  --- Both left and right vectors have null range "
	      SEVERITY ERROR;
              return(false);
         ELSIF( l'LENGTH = 0) THEN        -- left input is of null range
    	      ASSERT false
	      REPORT " --- left input has null range "
	      SEVERITY ERROR;
              return(true);

         ELSIF( r'LENGTH = 0) THEN        -- right  input is of null range
	      ASSERT false
	      REPORT " --- right input has null range "
	      SEVERITY ERROR;
              RETURN (false);
         END IF;
	-- synopsys translate_on        
 	-- input are not null so sign extend them to the same length
	vl := SignExtend(l, resltlen, l'LEFT, SrcRegMode);
	vr := SignExtend(r, resltlen, r'LEFT, SrcRegMode);

	IF (SrcRegMode = TwosComp) THEN
        	return ( LessThanOrEqual_TwosComp(vl, vr));
        ELSE
		return ( LessThanOrEqual_Unsigned(vl, vr));
	END IF;
     END RegLessThanOrEqual; 
     -- -----------------------------------------------------------------------------
     FUNCTION RegLessThanOrEqual ( CONSTANT l          : IN std_logic_vector;
				   CONSTANT r          : IN INTEGER;
  			           CONSTANT SrcRegMode : IN regmode_type
                     -- synopsys synthesis_off
					         	      := DefaultRegMode 
                     -- synopsys synthesis_on
				 ) RETURN BOOLEAN IS
       VARIABLE vl, vr    : std_logic_vector(IntegerBitLength - 1 DOWNTO 0);
     BEGIN
	-- synopsys translate_off
	-- Null range check
	 IF( l'LENGTH = 0) THEN        -- left input is of null range
    	      ASSERT false
	      REPORT " --- left input has null range "
	      SEVERITY ERROR;
              return(true);
         END IF;
	-- synopsys translate_on        
	-- input are not null so sign extend them to the same length
        -- Convert to std_logic_vector for comparison to allow any length input vector.
        vr := To_StdLogicVector ( r, IntegerBitLength, SrcRegMode );
 	vl := SignExtend(l, IntegerBitLength, l'LEFT, SrcRegMode);
	IF (SrcRegMode = TwosComp) THEN
        	return(LessThanOrEqual_TwosComp(vl, vr));
        ELSE
		return (LessThanOrEqual_Unsigned(vl, vr));
	END IF;
     END RegLessThanOrEqual; 
     -------------------------------------------------------------------------------
     FUNCTION RegLessThanOrEqual ( CONSTANT l          : IN INTEGER;
				   CONSTANT r          : IN std_logic_vector;
  			           CONSTANT SrcRegMode : IN regmode_type
                     -- synopsys synthesis_off
					         	      := DefaultRegMode 
                     -- synopsys synthesis_on
				 ) RETURN BOOLEAN IS
       VARIABLE vl, vr    : std_logic_vector(IntegerBitLength - 1 DOWNTO 0);
     BEGIN
	-- synopsys translate_off
	-- Null range check
	 IF( r'LENGTH = 0) THEN        -- right input is of null range
    	      ASSERT false
	      REPORT " --- left input has null range "
	      SEVERITY ERROR;
              return(false);
         END IF;
	-- synopsys translate_on        
	-- input are not null so sign extend them to the same length
        -- Convert to std_logic_vector for comparison to allow any length input vector.
        vl := To_StdLogicVector ( l, IntegerBitLength, SrcRegMode );
 	vr := SignExtend(r, IntegerBitLength, r'LEFT, SrcRegMode);
	IF (SrcRegMode = TwosComp) THEN
        	return(LessThanOrEqual_TwosComp(vl, vr));
        ELSE
		return (LessThanOrEqual_Unsigned(vl, vr));
	END IF;
     END RegLessThanOrEqual; 
     -------------------------------------------------------------------------------
     FUNCTION RegLessThanOrEqual ( CONSTANT l          : IN std_logic_vector;
				   CONSTANT r          : IN INTEGER;
  			           CONSTANT SrcRegMode : IN regmode_type
                     -- synopsys synthesis_off
					         	      := DefaultRegMode 
                     -- synopsys synthesis_on
				 ) RETURN std_ulogic IS
       VARIABLE vl, vr    : std_logic_vector(IntegerBitLength - 1 DOWNTO 0);
     BEGIN
        -- synopsys translate_off
	-- Null range check
         IF( l'LENGTH = 0) THEN        -- left input is of null range
    	      ASSERT false
	      REPORT " --- left input has null range "
	      SEVERITY ERROR;
              return('1');
         END IF;
	-- synopsys translate_on        
	-- input are not null so sign extend them to the same length
        -- Convert to std_logic_vector for comparison to allow any length input vector.
 	vl := SignExtend(l, IntegerBitLength, l'LEFT, SrcRegMode);
        vr := To_StdLogicVector ( r, IntegerBitLength, SrcRegMode );

	IF (SrcRegMode = TwosComp) THEN
        	return( To_StdULogic_loc( LessThanOrEqual_TwosComp(vl, vr)));
        ELSE
		return( To_StdULogic_loc (LessThanOrEqual_Unsigned(vl, vr)));
	END IF;
     END RegLessThanOrEqual; 
     -------------------------------------------------------------------------------
     FUNCTION RegLessThanOrEqual (  CONSTANT l          : IN INTEGER;
     				     CONSTANT r          : IN std_logic_vector;
				     CONSTANT SrcRegMode : IN regmode_type
                     -- synopsys synthesis_off
							      := DefaultRegMode 
                     -- synopsys synthesis_on
				   ) RETURN std_ulogic IS
       VARIABLE vl, vr    : std_logic_vector(IntegerBitLength - 1 DOWNTO 0);
     BEGIN
        -- synopsys translate_off
	-- Null range check
         IF( r'LENGTH = 0) THEN        -- left input is of null range
    	      ASSERT false
	      REPORT " --- left input has null range "
	      SEVERITY ERROR;
              return('0');
         END IF;
	-- synopsys translate_on        
	-- input are not null so sign extend them to the same length
        -- Convert to std_logic_vector for comparison to allow any length input vector.
        vl := To_StdLogicVector ( l, IntegerBitLength, SrcRegMode );
 	vr := SignExtend(r, IntegerBitLength, r'LEFT, SrcRegMode);

	IF (SrcRegMode = TwosComp) THEN
        	return( To_StdULogic_loc( LessThanOrEqual_TwosComp(vl, vr)));
        ELSE
		return( To_StdULogic_loc (LessThanOrEqual_Unsigned(vl, vr)));
	END IF;
     END RegLessThanOrEqual; 
     -- ----------------------------------------------------------------------------
     --     Function Name : RegLessThanOrEqual
     --    
     --     Purpose       : Compute a less than or equal relation for std_ulogic_vectors
     --     
     --     Parameters    : l       - input std_ulogic_vector | INTEGER
     --                     r       - input std_ulogic_vector | INTEGER
     --                     SrcRegMode - input regmode_type, indicating the format of
     --                               the std_ulogic_vector operands (l,r).
     --                               Default is TwosComp.
     --     
     --     Result        : BOOLEAN | std_ulogic
     --
     --     NOTE          : The operands may be of any length, and may be different
     --                     lengths. 
     --
     --                     Overloading not defined for both inputs of INTEGER type.
     --
     --                     Any time the comparison reaches an index that has an 'X' as an
     --                     array element, the comparison is deemed indeterminate and will 
     --                     return false in case of boolean and '0' incase of 
     --                     std_ulogic for synthesis purposes.
     --     Use           : 
     --                      VARIABLE a, b : std_ulogic_vector ( 7 DOWNTO 0 );
     --                      IF ( RegLessThanOrEqual ( a, b, TwosComp)   )  THEN 
     --     
     --     See Also      : RegLessThan, RegGreaterThan,   RegGreaterThanOrEqual.
     -------------------------------------------------------------------------------
     FUNCTION RegLessThanOrEqual ( CONSTANT l          : IN std_ulogic_vector;
				   CONSTANT r          : IN std_ulogic_vector;
  			           CONSTANT SrcRegMode : IN regmode_type
                     -- synopsys synthesis_off
					         	      := DefaultRegMode 
                     -- synopsys synthesis_on
				 ) RETURN std_ulogic IS
       CONSTANT resltlen : INTEGER := MAXIMUM (l'LENGTH, r'LENGTH);
       VARIABLE vl, vr   : STD_ULOGIC_VECTOR (resltlen - 1 DOWNTO 0);
     BEGIN
        -- synopsys translate_off
	-- Null range check
	IF ( (l'LENGTH = 0) AND (r'LENGTH = 0) ) THEN   
	      ASSERT false 
	      REPORT "  --- Both left and right vectors have null range "
	      SEVERITY ERROR;
              return( '0');
         ELSIF( l'LENGTH = 0) THEN        -- left input is of null range
    	      ASSERT false
	      REPORT " --- left input has null range "
	      SEVERITY ERROR;
              return('1');

         ELSIF( r'LENGTH = 0) THEN        -- right  input is of null range
	      ASSERT false
	      REPORT " --- right input has null range "
	      SEVERITY ERROR;
              RETURN ('0');
         END IF;
	-- synopsys translate_on        
 	-- input are not null so sign extend them to the same length
	vl := SignExtend(l, resltlen, l'LEFT, SrcRegMode);
	vr := SignExtend(r, resltlen, r'LEFT, SrcRegMode);

	IF (SrcRegMode = TwosComp) THEN
        	return( To_StdULogic_loc( LessThanOrEqual_TwosComp(vl, vr)));
        ELSE
		return( To_StdULogic_loc (LessThanOrEqual_Unsigned(vl, vr)));
	END IF;
     END RegLessThanOrEqual; 
     -----------------------------------------------------------------------------
     FUNCTION RegLessThanOrEqual ( CONSTANT l          : IN std_ulogic_vector;
				   CONSTANT r          : IN std_ulogic_vector;
 			           CONSTANT SrcRegMode : IN regmode_type
                     -- synopsys synthesis_off
							      := DefaultRegMode 
                     -- synopsys synthesis_on
				 ) RETURN BOOLEAN IS
       CONSTANT resltlen : INTEGER := MAXIMUM (l'LENGTH, r'LENGTH);
       VARIABLE vl, vr   : STD_ULOGIC_VECTOR (resltlen - 1 DOWNTO 0);
     BEGIN
        -- synopsys translate_off
	-- Null range check
	IF ( (l'LENGTH = 0) AND (r'LENGTH = 0) ) THEN   
	      ASSERT false 
	      REPORT "  --- Both left and right vectors have null range "
	      SEVERITY ERROR;
              return(false);
         ELSIF( l'LENGTH = 0) THEN        -- left input is of null range
    	      ASSERT false
	      REPORT " --- left input has null range "
	      SEVERITY ERROR;
              return(true);

         ELSIF( r'LENGTH = 0) THEN        -- right  input is of null range
	      ASSERT false
	      REPORT " --- right input has null range "
	      SEVERITY ERROR;
              RETURN (false);
         END IF;
	-- synopsys translate_on        
 	-- input are not null so sign extend them to the same length
	vl := SignExtend(l, resltlen, l'LEFT, SrcRegMode);
	vr := SignExtend(r, resltlen, r'LEFT, SrcRegMode);

	IF (SrcRegMode = TwosComp) THEN
        	return ( LessThanOrEqual_TwosComp(vl, vr));
        ELSE
		return ( LessThanOrEqual_Unsigned(vl, vr));
	END IF;
     END RegLessThanOrEqual; 
     -- -----------------------------------------------------------------------------
     FUNCTION RegLessThanOrEqual ( CONSTANT l          : IN std_ulogic_vector;
				   CONSTANT r          : IN INTEGER;
  			           CONSTANT SrcRegMode : IN regmode_type
                     -- synopsys synthesis_off
					         	      := DefaultRegMode 
                     -- synopsys synthesis_on
				 ) RETURN BOOLEAN IS
       VARIABLE vl, vr    : std_ulogic_vector(IntegerBitLength - 1 DOWNTO 0);
     BEGIN
	-- synopsys translate_off
	-- Null range check
	 IF( l'LENGTH = 0) THEN        -- left input is of null range
    	      ASSERT false
	      REPORT " --- left input has null range "
	      SEVERITY ERROR;
              return(true);
         END IF;
	-- synopsys translate_on        
	-- input are not null so sign extend them to the same length
        -- Convert to std_ulogic_vector for comparison to allow any length input vector.
        vr := To_StdULogicVector ( r, IntegerBitLength, SrcRegMode );
 	vl := SignExtend(l, IntegerBitLength, l'LEFT, SrcRegMode);
	IF (SrcRegMode = TwosComp) THEN
        	return(LessThanOrEqual_TwosComp(vl, vr));
        ELSE
		return (LessThanOrEqual_Unsigned(vl, vr));
	END IF;
     END RegLessThanOrEqual; 
     -------------------------------------------------------------------------------
     FUNCTION RegLessThanOrEqual ( CONSTANT l          : IN INTEGER;
				   CONSTANT r          : IN std_ulogic_vector;
  			           CONSTANT SrcRegMode : IN regmode_type
                     -- synopsys synthesis_off
					         	      := DefaultRegMode 
                     -- synopsys synthesis_on
				 ) RETURN BOOLEAN IS
       VARIABLE vl, vr    : std_ulogic_vector(IntegerBitLength - 1 DOWNTO 0);
     BEGIN
	-- synopsys translate_off
	-- Null range check
	 IF( r'LENGTH = 0) THEN        -- right input is of null range
    	      ASSERT false
	      REPORT " --- left input has null range "
	      SEVERITY ERROR;
              return(false);
         END IF;
	-- synopsys translate_on        
	-- input are not null so sign extend them to the same length
        -- Convert to std_ulogic_vector for comparison to allow any length input vector.
        vl := To_StdULogicVector ( l, IntegerBitLength, SrcRegMode );
 	vr := SignExtend(r, IntegerBitLength, r'LEFT, SrcRegMode);
	IF (SrcRegMode = TwosComp) THEN
        	return(LessThanOrEqual_TwosComp(vl, vr));
        ELSE
		return (LessThanOrEqual_Unsigned(vl, vr));
	END IF;
     END RegLessThanOrEqual; 
     -------------------------------------------------------------------------------
     FUNCTION RegLessThanOrEqual ( CONSTANT l          : IN std_ulogic_vector;
				   CONSTANT r          : IN INTEGER;
  			           CONSTANT SrcRegMode : IN regmode_type
                     -- synopsys synthesis_off
					         	      := DefaultRegMode 
                     -- synopsys synthesis_on
				 ) RETURN std_ulogic IS
       VARIABLE vl, vr    : std_ulogic_vector(IntegerBitLength - 1 DOWNTO 0);
     BEGIN
        -- synopsys translate_off
	-- Null range check
         IF( l'LENGTH = 0) THEN        -- left input is of null range
    	      ASSERT false
	      REPORT " --- left input has null range "
	      SEVERITY ERROR;
              return('1');
         END IF;
	-- synopsys translate_on        
	-- input are not null so sign extend them to the same length
        -- Convert to std_ulogic_vector for comparison to allow any length input vector.
 	vl := SignExtend(l, IntegerBitLength, l'LEFT, SrcRegMode);
        vr := To_StdULogicVector ( r, IntegerBitLength, SrcRegMode );

	IF (SrcRegMode = TwosComp) THEN
        	return( To_StdULogic_loc( LessThanOrEqual_TwosComp(vl, vr)));
        ELSE
		return( To_StdULogic_loc (LessThanOrEqual_Unsigned(vl, vr)));
	END IF;
     END RegLessThanOrEqual; 
     -------------------------------------------------------------------------------
     FUNCTION RegLessThanOrEqual  (  CONSTANT l          : IN INTEGER;
     				     CONSTANT r          : IN std_ulogic_vector;
				     CONSTANT SrcRegMode : IN regmode_type
                     -- synopsys synthesis_off
							      := DefaultRegMode 
                     -- synopsys synthesis_on
				   ) RETURN std_ulogic IS
       VARIABLE vl, vr    : std_ulogic_vector(IntegerBitLength - 1 DOWNTO 0);
     BEGIN
        -- synopsys translate_off
	-- Null range check
         IF( r'LENGTH = 0) THEN        -- left input is of null range
    	      ASSERT false
	      REPORT " --- left input has null range "
	      SEVERITY ERROR;
              return('0');
         END IF;
	-- synopsys translate_on        
	-- input are not null so sign extend them to the same length
        -- Convert to std_ulogic_vector for comparison to allow any length input vector.
        vl := To_StdULogicVector ( l, IntegerBitLength, SrcRegMode );
 	vr := SignExtend(r, IntegerBitLength, r'LEFT, SrcRegMode);

	IF (SrcRegMode = TwosComp) THEN
        	return( To_StdULogic_loc( LessThanOrEqual_TwosComp(vl, vr)));
        ELSE
		return( To_StdULogic_loc (LessThanOrEqual_Unsigned(vl, vr)));
	END IF;
     END RegLessThanOrEqual; 
     -------------------------------------------------------------------------------
     --     Function Name : RegGreaterThan
     -- 1.2.53
     --     Overloading   : Input parameter TYPEs.
     --
     --     Purpose       : Compute a greater than relation for bit_vectors
     --
     --     Parameters    : l       - input bit_vector | INTEGER
     --                     r       - input bit_vector | INTEGER
     --                     SrcRegMode - input regmode_type, indicating the format of
     --                               the bit_vector operands (l,r).
     --                               Default is TwosComp.
     --
     --     Result        : BOOLEAN | bit
     --
     --     NOTE          : The operands may be of any length, and may be different
     --                     lengths.
     --
     --                     Overloading not defined for both inputs of INTEGER type.
     --
     --     Use           :
     --                      VARIABLE a, b : bit_vector ( 7 DOWNTO 0 );
     --                      IF ( RegGreaterThan ( a, b, TwosComp)   )  THEN
     --
     --     See Also      :  RegLessThan, RegLessThanOrEqual, RegGreaterThanOrEqual.
     -------------------------------------------------------------------------------
     FUNCTION RegGreaterThan ( CONSTANT l          : IN bit_vector;
			       CONSTANT r          : IN bit_vector;
		               CONSTANT SrcRegMode : IN regmode_type
                     -- synopsys synthesis_off
							      := DefaultRegMode 
                     -- synopsys synthesis_on
				 ) RETURN bit IS
       CONSTANT resltlen : INTEGER := MAXIMUM (l'LENGTH, r'LENGTH);
       VARIABLE vl, vr   : BIT_VECTOR (resltlen - 1 DOWNTO 0);
     BEGIN
        -- synopsys translate_off
	-- Null range check
	IF ( (l'LENGTH = 0) AND (r'LENGTH = 0) ) THEN   
	      ASSERT false 
	      REPORT "  --- Both left and right vectors have null range "
	      SEVERITY ERROR;
              return( '0');
         ELSIF( l'LENGTH = 0) THEN        -- left input is of null range
    	      ASSERT false
	      REPORT " --- left input has null range "
	      SEVERITY ERROR;
              return('0');

         ELSIF( r'LENGTH = 0) THEN        -- right  input is of null range
	      ASSERT false
	      REPORT " --- right input has null range "
	      SEVERITY ERROR;
              RETURN ('1');
         END IF;
	-- synopsys translate_on        
 	-- input are not null so sign extend them to the same length
	vl := SignExtend(l, resltlen, l'LEFT, SrcRegMode);
	vr := SignExtend(r, resltlen, r'LEFT, SrcRegMode);

	IF (SrcRegMode = TwosComp) THEN
        	return (To_Bit_loc(NOT (LessThanOrEqual_TwosComp(vl, vr))));
        ELSE
		return (To_Bit_loc(NOT (LessThanOrEqual_Unsigned(vl, vr))));
	END IF;
     END RegGreaterThan; 
     -----------------------------------------------------------------------------
     FUNCTION RegGreaterThan    ( CONSTANT l          : IN bit_vector;
				   CONSTANT r          : IN bit_vector;
 			           CONSTANT SrcRegMode : IN regmode_type
                     -- synopsys synthesis_off
							      := DefaultRegMode 
                     -- synopsys synthesis_on
				 ) RETURN BOOLEAN IS
       CONSTANT resltlen : INTEGER := MAXIMUM (l'LENGTH, r'LENGTH);
       VARIABLE vl, vr   : BIT_VECTOR (resltlen - 1 DOWNTO 0);
     BEGIN
        -- synopsys translate_off
	-- Null range check
	IF ( (l'LENGTH = 0) AND (r'LENGTH = 0) ) THEN   
	      ASSERT false 
	      REPORT "  --- Both left and right vectors have null range "
	      SEVERITY ERROR;
              return( false);
         ELSIF( l'LENGTH = 0) THEN        -- left input is of null range
    	      ASSERT false
	      REPORT " --- left input has null range "
	      SEVERITY ERROR;
              return(false);

         ELSIF( r'LENGTH = 0) THEN        -- right  input is of null range
	      ASSERT false
	      REPORT " --- right input has null range "
	      SEVERITY ERROR;
              RETURN (true);
         END IF;
	-- synopsys translate_on        
 	-- input are not null so sign extend them to the same length
	vl := SignExtend(l, resltlen, l'LEFT, SrcRegMode);
	vr := SignExtend(r, resltlen, r'LEFT, SrcRegMode);

	IF (SrcRegMode = TwosComp) THEN
        	return (NOT (LessThanOrEqual_TwosComp(vl, vr)));
        ELSE
		return (NOT (LessThanOrEqual_Unsigned(vl, vr)));
	END IF;
     END RegGreaterThan; 
     -- -----------------------------------------------------------------------------
     FUNCTION RegGreaterThan ( CONSTANT l          : IN bit_vector;
				   CONSTANT r          : IN INTEGER;
			     CONSTANT SrcRegMode : IN regmode_type
                     -- synopsys synthesis_off
						      := DefaultRegMode 
                     -- synopsys synthesis_on
				 ) RETURN BOOLEAN IS
	VARIABLE vl, vr    : bit_vector(IntegerBitLength - 1 DOWNTO 0);
     BEGIN
	-- synopsys translate_off
	-- Null range check
	 IF( l'LENGTH = 0) THEN        -- left input is of null range
    	      ASSERT false
	      REPORT " --- left input has null range "
	      SEVERITY ERROR;
              return(false);
         END IF;
	-- synopsys translate_on        
	-- input are not null so sign extend them to the same length
        -- Convert to bit_vector for comparison to allow any length input vector.
        vr := To_BitVector ( r, IntegerBitLength, SrcRegMode );
 	vl := SignExtend(l, IntegerBitLength, l'LEFT, SrcRegMode);

	IF (SrcRegMode = TwosComp) THEN
        	return (NOT (LessThanOrEqual_TwosComp(vl, vr)));
        ELSE
		return (NOT (LessThanOrEqual_Unsigned(vl, vr)));
	END IF;
     END RegGreaterThan; 
     -------------------------------------------------------------------------------
     FUNCTION RegGreaterThan ( CONSTANT l          : IN INTEGER;
				   CONSTANT r          : IN bit_vector;
  			           CONSTANT SrcRegMode : IN regmode_type
                     -- synopsys synthesis_off
					         	      := DefaultRegMode 
                     -- synopsys synthesis_on
				 ) RETURN BOOLEAN IS
       VARIABLE vl, vr    : bit_vector(IntegerBitLength - 1 DOWNTO 0);
     BEGIN
	-- synopsys translate_off
	-- Null range check
	 IF( r'LENGTH = 0) THEN        -- right input is of null range
    	      ASSERT false
	      REPORT " --- left input has null range "
	      SEVERITY ERROR;
              return(true);
         END IF;
	-- synopsys translate_on        
	-- input are not null so sign extend them to the same length
        -- Convert to bit_vector for comparison to allow any length input vector.
        vl := To_BitVector ( l, IntegerBitLength, SrcRegMode );
 	vr := SignExtend(r, IntegerBitLength, r'LEFT, SrcRegMode);
	IF (SrcRegMode = TwosComp) THEN
        	return (NOT (LessThanOrEqual_TwosComp(vl, vr)));
        ELSE
		return (NOT (LessThanOrEqual_Unsigned(vl, vr)));
	END IF;
     END RegGreaterThan; 
     -------------------------------------------------------------------------------
     FUNCTION RegGreaterThan ( CONSTANT l          : IN bit_vector;
				   CONSTANT r          : IN INTEGER;
  			           CONSTANT SrcRegMode : IN regmode_type
                     -- synopsys synthesis_off
					         	      := DefaultRegMode 
                     -- synopsys synthesis_on
				 ) RETURN bit IS
       VARIABLE vl, vr    : bit_vector(IntegerBitLength - 1 DOWNTO 0);
     BEGIN
        -- synopsys translate_off
	-- Null range check
         IF( l'LENGTH = 0) THEN        -- left input is of null range
    	      ASSERT false
	      REPORT " --- left input has null range "
	      SEVERITY ERROR;
              return('0');
         END IF;
	-- synopsys translate_on        
	-- input are not null so sign extend them to the same length
        -- Convert to bit_vector for comparison to allow any length input vector.
 	vl := SignExtend(l, IntegerBitLength, l'LEFT, SrcRegMode);
        vr := To_BitVector ( r, IntegerBitLength, SrcRegMode );

	IF (SrcRegMode = TwosComp) THEN
        	return( To_Bit_loc (NOT ( LessThanOrEqual_TwosComp(vl, vr))));
        ELSE
		return( To_Bit_loc (NOT (LessThanOrEqual_Unsigned(vl, vr))));
	END IF;
     END RegGreaterThan; 
     -------------------------------------------------------------------------------
     FUNCTION RegGreaterThan ( CONSTANT l          : IN INTEGER;
				   CONSTANT r          : IN bit_vector;
  			           CONSTANT SrcRegMode : IN regmode_type
                     -- synopsys synthesis_off
					         	      := DefaultRegMode 
                     -- synopsys synthesis_on
				 ) RETURN bit IS
       VARIABLE vl, vr    : bit_vector(IntegerBitLength - 1 DOWNTO 0);
     BEGIN
        -- synopsys translate_off
	-- Null range check
         IF( r'LENGTH = 0) THEN        -- left input is of null range
    	      ASSERT false
	      REPORT " --- left input has null range "
	      SEVERITY ERROR;
              return('1');
         END IF;
	-- synopsys translate_on        
	-- input are not null so sign extend them to the same length
        -- Convert to bit_vector for comparison to allow any length input vector.
        vl := To_BitVector ( l, IntegerBitLength, SrcRegMode );
 	vr := SignExtend(r, IntegerBitLength, r'LEFT, SrcRegMode);

	IF (SrcRegMode = TwosComp) THEN
        	return( To_Bit_loc( NOT(  LessThanOrEqual_TwosComp(vl, vr))));
        ELSE
		return( To_Bit_loc( NOT (LessThanOrEqual_Unsigned(vl, vr))));
	END IF;
     END RegGreaterThan; 
     -- ----------------------------------------------------------------------------
     --     Function Name : RegGreaterThan
     --
     --     Overloading   : Input parameter TYPEs.
     --    
     --     Purpose       : Compute a greater than relation for std_logic_vectors
     --     
     --     Parameters    : l       - input std_logic_vector | INTEGER
     --                     r       - input std_logic_vector | INTEGER
     --                     SrcRegMode - input regmode_type, indicating the format of
     --                               the std_logic_vector operands (l,r).
     --                               Default is TwosComp.
     --     
     --     Result        : BOOLEAN | std_ulogic
     --
     --     NOTE          : The operands may be of any length, and may be different
     --                     lengths. 
     --
     --                     Overloading not defined for both inputs of INTEGER type.
     --
     --                     Any time the comparison reaches an index that has an 'X' as
     --                     an array element, the comparison is deemed indeterminate  
     --                     and will return false in case of boolean and '0' incase of 
     --                     std_ulogic for synthesis purposes.
     --     Use           : 
     --                      VARIABLE a, b : std_logic_vector ( 7 DOWNTO 0 );
     --                      IF ( RegGreaterThan ( a, b, TwosComp)   )  THEN 
     --     
     --     See Also      : RegLessThan, RegLessThanOrEqual, RegGreaterThan, 
     --                     RegGreaterThanOrEqual.
     -------------------------------------------------------------------------------
     FUNCTION RegGreaterThan  ( CONSTANT l          : IN std_logic_vector;
				CONSTANT r          : IN std_logic_vector;
				CONSTANT SrcRegMode : IN regmode_type 

                     -- synopsys synthesis_off
							      := DefaultRegMode 
                     -- synopsys synthesis_on
				 ) RETURN std_ulogic IS
       CONSTANT resltlen : INTEGER := MAXIMUM (l'LENGTH, r'LENGTH);
       VARIABLE vl, vr   : STD_LOGIC_VECTOR (resltlen - 1 DOWNTO 0);
     BEGIN
        -- synopsys translate_off
	-- Null range check
	IF ( (l'LENGTH = 0) AND (r'LENGTH = 0) ) THEN   
	      ASSERT false 
	      REPORT "  --- Both left and right vectors have null range "
	      SEVERITY ERROR;
              return( '0');
         ELSIF( l'LENGTH = 0) THEN        -- left input is of null range
    	      ASSERT false
	      REPORT " --- left input has null range "
	      SEVERITY ERROR;
              return('0');

         ELSIF( r'LENGTH = 0) THEN        -- right  input is of null range
	      ASSERT false
	      REPORT " --- right input has null range "
	      SEVERITY ERROR;
              RETURN ('1');
         END IF;
	-- synopsys translate_on        
 	-- input are not null so sign extend them to the same length
	vl := SignExtend(l, resltlen, l'LEFT, SrcRegMode);
	vr := SignExtend(r, resltlen, r'LEFT, SrcRegMode);

	IF (SrcRegMode = TwosComp) THEN
        	return( To_StdULogic_loc (LessThan_TwosComp(vr, vl)));
        ELSE
		return( To_StdULogic_loc (LessThan_Unsigned(vr, vl)));
	END IF;
     END RegGreaterThan; 
     -----------------------------------------------------------------------------
     FUNCTION RegGreaterThan    ( CONSTANT l          : IN std_logic_vector;
				   CONSTANT r          : IN std_logic_vector;
 			           CONSTANT SrcRegMode : IN regmode_type
                     -- synopsys synthesis_off
							      := DefaultRegMode 
                     -- synopsys synthesis_on
				 ) RETURN BOOLEAN IS
       CONSTANT resltlen : INTEGER := MAXIMUM (l'LENGTH, r'LENGTH);
       VARIABLE vl, vr   : STD_LOGIC_VECTOR (resltlen - 1 DOWNTO 0);
     BEGIN
        -- synopsys translate_off
	-- Null range check
	IF ( (l'LENGTH = 0) AND (r'LENGTH = 0) ) THEN   
	      ASSERT false 
	      REPORT "  --- Both left and right vectors have null range "
	      SEVERITY ERROR;
              return( false);
         ELSIF( l'LENGTH = 0) THEN        -- left input is of null range
    	      ASSERT false
	      REPORT " --- left input has null range "
	      SEVERITY ERROR;
              return(false);

         ELSIF( r'LENGTH = 0) THEN        -- right  input is of null range
	      ASSERT false
	      REPORT " --- right input has null range "
	      SEVERITY ERROR;
              RETURN (true);
         END IF;
	-- synopsys translate_on        
 	-- input are not null so sign extend them to the same length
	vl := SignExtend(l, resltlen, l'LEFT, SrcRegMode);
	vr := SignExtend(r, resltlen, r'LEFT, SrcRegMode);

	IF (SrcRegMode = TwosComp) THEN
        	return(LessThan_TwosComp(vr, vl));
        ELSE
		return( LessThan_Unsigned(vr, vl));
	END IF;
     END RegGreaterThan; 
     -- -----------------------------------------------------------------------------
     FUNCTION RegGreaterThan ( CONSTANT l          : IN std_logic_vector;
				   CONSTANT r          : IN INTEGER;
			     CONSTANT SrcRegMode : IN regmode_type
                     -- synopsys synthesis_off
						      := DefaultRegMode 
                     -- synopsys synthesis_on
				 ) RETURN BOOLEAN IS
	VARIABLE vl, vr    : std_logic_vector(IntegerBitLength - 1 DOWNTO 0);
     BEGIN
	-- synopsys translate_off
	-- Null range check
	 IF( l'LENGTH = 0) THEN        -- left input is of null range
    	      ASSERT false
	      REPORT " --- left input has null range "
	      SEVERITY ERROR;
              return(false);
         END IF;
	-- synopsys translate_on        
	-- input are not null so sign extend them to the same length
        -- Convert to std_logic_vector for comparison to allow any length input vector.
        vr := To_StdLogicVector ( r, IntegerBitLength, SrcRegMode );
 	vl := SignExtend(l, IntegerBitLength, l'LEFT, SrcRegMode);

	IF (SrcRegMode = TwosComp) THEN
        	return( LessThan_TwosComp(vr, vl));
        ELSE
		return( LessThan_Unsigned(vr, vl));
	END IF;

     END RegGreaterThan; 
     -------------------------------------------------------------------------------
     FUNCTION RegGreaterThan ( CONSTANT l          : IN INTEGER;
				   CONSTANT r          : IN std_logic_vector;
  			           CONSTANT SrcRegMode : IN regmode_type
                     -- synopsys synthesis_off
					         	      := DefaultRegMode 
                     -- synopsys synthesis_on
				 ) RETURN BOOLEAN IS
       VARIABLE vl, vr    : std_logic_vector(IntegerBitLength - 1 DOWNTO 0);
     BEGIN
	-- synopsys translate_off
	-- Null range check
	 IF( r'LENGTH = 0) THEN        -- right input is of null range
    	      ASSERT false
	      REPORT " --- left input has null range "
	      SEVERITY ERROR;
              return(true);
         END IF;
	-- synopsys translate_on        
	-- input are not null so sign extend them to the same length
        -- Convert to std_logic_vector for comparison to allow any length input vector.
        vl := To_StdLogicVector ( l, IntegerBitLength, SrcRegMode );
 	vr := SignExtend(r, IntegerBitLength, r'LEFT, SrcRegMode);

	IF (SrcRegMode = TwosComp) THEN
        	return( LessThan_TwosComp(vr, vl));
        ELSE
		return( LessThan_Unsigned(vr, vl));
	END IF;
     END RegGreaterThan; 
     -------------------------------------------------------------------------------
     FUNCTION RegGreaterThan ( CONSTANT l          : IN std_logic_vector;
				   CONSTANT r          : IN INTEGER;
  			           CONSTANT SrcRegMode : IN regmode_type
                     -- synopsys synthesis_off
					         	      := DefaultRegMode 
                     -- synopsys synthesis_on
				 ) RETURN std_ulogic IS
       VARIABLE vl, vr    : std_logic_vector(IntegerBitLength - 1 DOWNTO 0);
     BEGIN
        -- synopsys translate_off
	-- Null range check
         IF( l'LENGTH = 0) THEN        -- left input is of null range
    	      ASSERT false
	      REPORT " --- left input has null range "
	      SEVERITY ERROR;
              return('0');
         END IF;
	-- synopsys translate_on        
	-- input are not null so sign extend them to the same length
        -- Convert to std_logic_vector for comparison to allow any length input vector.
 	vl := SignExtend(l, IntegerBitLength, l'LEFT, SrcRegMode);
        vr := To_StdLogicVector ( r, IntegerBitLength, SrcRegMode );

	IF (SrcRegMode = TwosComp) THEN
        	return( To_StdULogic_loc (LessThan_TwosComp(vr, vl)));
        ELSE
		return( To_StdULogic_loc (LessThan_Unsigned(vr, vl)));
	END IF;
    END RegGreaterThan; 
     -------------------------------------------------------------------------------
     FUNCTION RegGreaterThan ( CONSTANT l          : IN INTEGER;
				   CONSTANT r          : IN std_logic_vector;
  			           CONSTANT SrcRegMode : IN regmode_type
                     -- synopsys synthesis_off
					         	      := DefaultRegMode 
                     -- synopsys synthesis_on
				 ) RETURN std_ulogic IS
       VARIABLE vl, vr    : std_logic_vector(IntegerBitLength - 1 DOWNTO 0);
     BEGIN
        -- synopsys translate_off
	-- Null range check
         IF( r'LENGTH = 0) THEN        -- left input is of null range
    	      ASSERT false
	      REPORT " --- left input has null range "
	      SEVERITY ERROR;
              return('1');
         END IF;
	-- synopsys translate_on        
	-- input are not null so sign extend them to the same length
        -- Convert to std_logic_vector for comparison to allow any length input vector.
        vl := To_StdLogicVector ( l, IntegerBitLength, SrcRegMode );
 	vr := SignExtend(r, IntegerBitLength, r'LEFT, SrcRegMode);


	IF (SrcRegMode = TwosComp) THEN
        	return( To_StdULogic_loc (LessThan_TwosComp(vr, vl)));
        ELSE
		return( To_StdULogic_loc (LessThan_Unsigned(vr, vl)));
	END IF;
    END RegGreaterThan; 
     -- ----------------------------------------------------------------------------
     --     Function Name : RegGreaterThan
     --
     --     Overloading   : Input parameter TYPEs.
     --    
     --     Purpose       : Compute a greater than relation for std_logic_vectors
     --     
     --     Parameters    : l       - input std_ulogic_vector | INTEGER
     --                     r       - input std_ulogic_vector | INTEGER
     --                     SrcRegMode - input regmode_type, indicating the format of
     --                               the std_ulogic_vector operands (l,r).
     --                               Default is TwosComp.
     --     
     --     Result        : BOOLEAN | std_ulogic
     --
     --     NOTE          : The operands may be of any length, and may be different
     --                     lengths. 
     --
     --                     Overloading not defined for both inputs of INTEGER type.
     --
     --                     Any time the comparison reaches an index that has an 'X' as
     --                     an array element, the comparison is deemed indeterminate  
     --                     and will return false in case of boolean and '0' incase of
     --                     std_ulogic for synthesis purposes.
     --     Use           : 
     --                      VARIABLE a, b : std_ulogic_vector ( 7 DOWNTO 0 );
     --                      IF ( RegGreaterThan ( a, b, TwosComp)   )  THEN 
     --     
     --     See Also      : RegLessThan, RegLessThanOrEqual, RegGreaterThanOrEqual.
     -------------------------------------------------------------------------------
     FUNCTION RegGreaterThan  ( CONSTANT l          : IN std_ulogic_vector;
				CONSTANT r          : IN std_ulogic_vector;
				CONSTANT SrcRegMode : IN regmode_type 
                     -- synopsys synthesis_off
							      := DefaultRegMode 
                     -- synopsys synthesis_on
				 ) RETURN std_ulogic IS
       CONSTANT resltlen : INTEGER := MAXIMUM (l'LENGTH, r'LENGTH);
       VARIABLE vl, vr   : STD_ULOGIC_VECTOR (resltlen - 1 DOWNTO 0);
     BEGIN
        -- synopsys translate_off
	-- Null range check
	IF ( (l'LENGTH = 0) AND (r'LENGTH = 0) ) THEN   
	      ASSERT false 
	      REPORT "  --- Both left and right vectors have null range "
	      SEVERITY ERROR;
              return( '0');
         ELSIF( l'LENGTH = 0) THEN        -- left input is of null range
    	      ASSERT false
	      REPORT " --- left input has null range "
	      SEVERITY ERROR;
              return('0');

         ELSIF( r'LENGTH = 0) THEN        -- right  input is of null range
	      ASSERT false
	      REPORT " --- right input has null range "
	      SEVERITY ERROR;
              RETURN ('1');
         END IF;
	-- synopsys translate_on        
 	-- input are not null so sign extend them to the same length
	vl := SignExtend(l, resltlen, l'LEFT, SrcRegMode);
	vr := SignExtend(r, resltlen, r'LEFT, SrcRegMode);

	IF (SrcRegMode = TwosComp) THEN
        	return( To_StdULogic_loc (LessThan_TwosComp(vr, vl)));
        ELSE
		return( To_StdULogic_loc (LessThan_Unsigned(vr, vl)));
	END IF;
    END RegGreaterThan; 
     -----------------------------------------------------------------------------
     FUNCTION RegGreaterThan    ( CONSTANT l          : IN std_ulogic_vector;
				   CONSTANT r          : IN std_ulogic_vector;
 			           CONSTANT SrcRegMode : IN regmode_type
                     -- synopsys synthesis_off
							      := DefaultRegMode 
                     -- synopsys synthesis_on
				 ) RETURN BOOLEAN IS
       CONSTANT resltlen : INTEGER := MAXIMUM (l'LENGTH, r'LENGTH);
       VARIABLE vl, vr   : STD_ULOGIC_VECTOR (resltlen - 1 DOWNTO 0);
     BEGIN
        -- synopsys translate_off
	-- Null range check
	IF ( (l'LENGTH = 0) AND (r'LENGTH = 0) ) THEN   
	      ASSERT false 
	      REPORT "  --- Both left and right vectors have null range "
	      SEVERITY ERROR;
              return( false);
         ELSIF( l'LENGTH = 0) THEN        -- left input is of null range
    	      ASSERT false
	      REPORT " --- left input has null range "
	      SEVERITY ERROR;
              return(false);

         ELSIF( r'LENGTH = 0) THEN        -- right  input is of null range
	      ASSERT false
	      REPORT " --- right input has null range "
	      SEVERITY ERROR;
              RETURN (true);
         END IF;
	-- synopsys translate_on        
 	-- input are not null so sign extend them to the same length
	vl := SignExtend(l, resltlen, l'LEFT, SrcRegMode);
	vr := SignExtend(r, resltlen, r'LEFT, SrcRegMode);

	IF (SrcRegMode = TwosComp) THEN
        	return( LessThan_TwosComp(vr, vl));
        ELSE
		return( LessThan_Unsigned(vr, vl));
	END IF;

    END RegGreaterThan; 
     -- -----------------------------------------------------------------------------
     FUNCTION RegGreaterThan ( CONSTANT l          : IN std_ulogic_vector;
				   CONSTANT r          : IN INTEGER;
			     CONSTANT SrcRegMode : IN regmode_type
                     -- synopsys synthesis_off
						      := DefaultRegMode 
                     -- synopsys synthesis_on
				 ) RETURN BOOLEAN IS
	VARIABLE vl, vr    : std_ulogic_vector(IntegerBitLength - 1 DOWNTO 0);
     BEGIN
	-- synopsys translate_off
	-- Null range check
	 IF( l'LENGTH = 0) THEN        -- left input is of null range
    	      ASSERT false
	      REPORT " --- left input has null range "
	      SEVERITY ERROR;
              return(false);
         END IF;
	-- synopsys translate_on        
	-- input are not null so sign extend them to the same length
        -- Convert to std_ulogic_vector for comparison to allow any length input vector.
        vr := To_StdULogicVector ( r, IntegerBitLength, SrcRegMode );
 	vl := SignExtend(l, IntegerBitLength, l'LEFT, SrcRegMode);

	IF (SrcRegMode = TwosComp) THEN
        	return( LessThan_TwosComp(vr, vl));
        ELSE
		return( LessThan_Unsigned(vr, vl));
	END IF;
     END RegGreaterThan; 
     -------------------------------------------------------------------------------
     FUNCTION RegGreaterThan ( CONSTANT l          : IN INTEGER;
				   CONSTANT r          : IN std_ulogic_vector;
  			           CONSTANT SrcRegMode : IN regmode_type
                     -- synopsys synthesis_off
					         	      := DefaultRegMode 
                     -- synopsys synthesis_on
				 ) RETURN BOOLEAN IS
       VARIABLE vl, vr    : std_ulogic_vector(IntegerBitLength - 1 DOWNTO 0);
     BEGIN
	-- synopsys translate_off
	-- Null range check
	 IF( r'LENGTH = 0) THEN        -- right input is of null range
    	      ASSERT false
	      REPORT " --- left input has null range "
	      SEVERITY ERROR;
              return(true);
         END IF;
	-- synopsys translate_on        
	-- input are not null so sign extend them to the same length
        -- Convert to std_ulogic_vector for comparison to allow any length input vector.
        vl := To_StdULogicVector ( l, IntegerBitLength, SrcRegMode );
 	vr := SignExtend(r, IntegerBitLength, r'LEFT, SrcRegMode);

	IF (SrcRegMode = TwosComp) THEN
        	return( LessThan_TwosComp(vr, vl));
        ELSE
		return( LessThan_Unsigned(vr, vl));
	END IF;
     END RegGreaterThan; 
     -------------------------------------------------------------------------------
     FUNCTION RegGreaterThan ( CONSTANT l          : IN std_ulogic_vector;
				   CONSTANT r          : IN INTEGER;
  			           CONSTANT SrcRegMode : IN regmode_type
                     -- synopsys synthesis_off
					         	      := DefaultRegMode 
                     -- synopsys synthesis_on
				 ) RETURN std_ulogic IS
       VARIABLE vl, vr    : std_ulogic_vector(IntegerBitLength - 1 DOWNTO 0);
     BEGIN
        -- synopsys translate_off
	-- Null range check
         IF( l'LENGTH = 0) THEN        -- left input is of null range
    	      ASSERT false
	      REPORT " --- left input has null range "
	      SEVERITY ERROR;
              return('0');
         END IF;
	-- synopsys translate_on        
	-- input are not null so sign extend them to the same length
        -- Convert to std_ulogic_vector for comparison to allow any length input vector.
 	vl := SignExtend(l, IntegerBitLength, l'LEFT, SrcRegMode);
        vr := To_StdULogicVector ( r, IntegerBitLength, SrcRegMode );

	IF (SrcRegMode = TwosComp) THEN
        	return( To_StdULogic_loc (LessThan_TwosComp(vr, vl)));
        ELSE
		return( To_StdULogic_loc (LessThan_Unsigned(vr, vl)));
	END IF;
    END RegGreaterThan; 
     -------------------------------------------------------------------------------
     FUNCTION RegGreaterThan ( CONSTANT l          : IN INTEGER;
				   CONSTANT r          : IN std_ulogic_vector;
  			           CONSTANT SrcRegMode : IN regmode_type
                     -- synopsys synthesis_off
					         	      := DefaultRegMode 
                     -- synopsys synthesis_on
				 ) RETURN std_ulogic IS
       VARIABLE vl, vr    : std_ulogic_vector(IntegerBitLength - 1 DOWNTO 0);
     BEGIN
        -- synopsys translate_off
	-- Null range check
         IF( r'LENGTH = 0) THEN        -- left input is of null range
    	      ASSERT false
	      REPORT " --- left input has null range "
	      SEVERITY ERROR;
              return('1');
         END IF;
	-- synopsys translate_on        
	-- input are not null so sign extend them to the same length
        -- Convert to std_ulogic_vector for comparison to allow any length input vector.
        vl := To_StdULogicVector ( l, IntegerBitLength, SrcRegMode );
 	vr := SignExtend(r, IntegerBitLength, r'LEFT, SrcRegMode);

	IF (SrcRegMode = TwosComp) THEN
        	return( To_StdULogic_loc (LessThan_TwosComp(vr, vl)));
        ELSE
		return( To_StdULogic_loc (LessThan_Unsigned(vr, vl)));
	END IF;

    END RegGreaterThan; 
     -------------------------------------------------------------------------------
     --     Function Name : RegGreaterThanOrEqual
     -- 1.2.53
     --     Overloading   : Input parameter TYPEs.
     --
     --     Purpose       : Compute a greater-than-or-equal relation for bit_vectors
     --
     --     Parameters    : l       - input bit_vector | INTEGER
     --                     r       - input bit_vector | INTEGER
     --                     SrcRegMode - input regmode_type, indicating the format of
     --                               the bit_vector operands (l,r).
     --                               Default is TwosComp.
     --
     --     Result        : BOOLEAN | bit
     --
     --     NOTE          : The operands may be of any length, and may be different
     --                     lengths.
     --
     --                     Overloading not defined for both inputs of INTEGER type.
     --
     --     Use           :
     --                      VARIABLE a, b : bit_vector ( 7 DOWNTO 0 );
     --                      IF ( RegGreaterThanOrEqual ( a, b, TwosComp)   )  THEN
     --
     --     See Also      :  RegLessThan, RegLessThanOrEqual, RegGreaterThan,
     -------------------------------------------------------------------------------
     FUNCTION RegGreaterThanOrEqual ( CONSTANT l          : IN bit_vector;
			       CONSTANT r          : IN bit_vector;
		               CONSTANT SrcRegMode : IN regmode_type
                     -- synopsys synthesis_off
							      := DefaultRegMode 
                     -- synopsys synthesis_on
				 ) RETURN bit IS
       CONSTANT resltlen : INTEGER := MAXIMUM (l'LENGTH, r'LENGTH);
       VARIABLE vl, vr   : BIT_VECTOR (resltlen - 1 DOWNTO 0);
     BEGIN
        -- synopsys translate_off
	-- Null range check
	IF ( (l'LENGTH = 0) AND (r'LENGTH = 0) ) THEN   
	      ASSERT false 
	      REPORT "  --- Both left and right vectors have null range "
	      SEVERITY ERROR;
              return( '0');
         ELSIF( l'LENGTH = 0) THEN        -- left input is of null range
    	      ASSERT false
	      REPORT " --- left input has null range "
	      SEVERITY ERROR;
              return('0');

         ELSIF( r'LENGTH = 0) THEN        -- right  input is of null range
	      ASSERT false
	      REPORT " --- right input has null range "
	      SEVERITY ERROR;
              RETURN ('1');
         END IF;
	-- synopsys translate_on        
 	-- input are not null so sign extend them to the same length
	vl := SignExtend(l, resltlen, l'LEFT, SrcRegMode);
	vr := SignExtend(r, resltlen, r'LEFT, SrcRegMode);

	IF (SrcRegMode = TwosComp) THEN
        	return( To_Bit_loc (NOT (LessThan_TwosComp(vl, vr))));
        ELSE
		return( To_Bit_loc ( NOT(LessThan_Unsigned(vl, vr))));
	END IF;
    END RegGreaterThanOrEqual; 
     -----------------------------------------------------------------------------
     FUNCTION RegGreaterThanOrEqual    ( CONSTANT l          : IN bit_vector;
				   CONSTANT r          : IN bit_vector;
 			           CONSTANT SrcRegMode : IN regmode_type
                     -- synopsys synthesis_off
							      := DefaultRegMode 
                     -- synopsys synthesis_on
				 ) RETURN BOOLEAN IS
       CONSTANT resltlen : INTEGER := MAXIMUM (l'LENGTH, r'LENGTH);
       VARIABLE vl, vr   : BIT_VECTOR (resltlen - 1 DOWNTO 0);
     BEGIN
        -- synopsys translate_off
	-- Null range check
	IF ( (l'LENGTH = 0) AND (r'LENGTH = 0) ) THEN   
	      ASSERT false 
	      REPORT "  --- Both left and right vectors have null range "
	      SEVERITY ERROR;
              return( false);
         ELSIF( l'LENGTH = 0) THEN        -- left input is of null range
    	      ASSERT false
	      REPORT " --- left input has null range "
	      SEVERITY ERROR;
              return(false);

         ELSIF( r'LENGTH = 0) THEN        -- right  input is of null range
	      ASSERT false
	      REPORT " --- right input has null range "
	      SEVERITY ERROR;
              RETURN (true);
         END IF;
	-- synopsys translate_on        
 	-- input are not null so sign extend them to the same length
	vl := SignExtend(l, resltlen, l'LEFT, SrcRegMode);
	vr := SignExtend(r, resltlen, r'LEFT, SrcRegMode);

	IF (SrcRegMode = TwosComp) THEN
        	return (NOT ( LessThan_TwosComp(vl, vr)));
        ELSE
		return ( NOT ( LessThan_Unsigned(vl, vr)));
	END IF;
    END RegGreaterThanOrEqual; 
     -- -----------------------------------------------------------------------------
     FUNCTION RegGreaterThanOrEqual ( CONSTANT l          : IN bit_vector;
				   CONSTANT r          : IN INTEGER;
			     CONSTANT SrcRegMode : IN regmode_type
                     -- synopsys synthesis_off
						      := DefaultRegMode 
                     -- synopsys synthesis_on
				 ) RETURN BOOLEAN IS
	VARIABLE vl, vr    : bit_vector(IntegerBitLength - 1 DOWNTO 0);
     BEGIN
	-- synopsys translate_off
	-- Null range check
	 IF( l'LENGTH = 0) THEN        -- left input is of null range
    	      ASSERT false
	      REPORT " --- left input has null range "
	      SEVERITY ERROR;
              return(false);
         END IF;
	-- synopsys translate_on        
	-- input are not null so sign extend them to the same length
        -- Convert to bit_vector for comparison to allow any length input vector.
        vr := To_BitVector ( r, IntegerBitLength, SrcRegMode );
 	vl := SignExtend(l, IntegerBitLength, l'LEFT, SrcRegMode);
	IF (SrcRegMode = TwosComp) THEN
        	return ( NOT (LessThan_TwosComp(vl, vr)));
        ELSE
		return ( NOT (LessThan_Unsigned(vl, vr)));
	END IF;
     END RegGreaterThanOrEqual; 
     -------------------------------------------------------------------------------
     FUNCTION RegGreaterThanOrEqual ( CONSTANT l          : IN INTEGER;
				   CONSTANT r          : IN bit_vector;
  			           CONSTANT SrcRegMode : IN regmode_type
                     -- synopsys synthesis_off
					         	      := DefaultRegMode 
                     -- synopsys synthesis_on
				 ) RETURN BOOLEAN IS
       VARIABLE vl, vr    : bit_vector(IntegerBitLength - 1 DOWNTO 0);
     BEGIN
	-- synopsys translate_off
	-- Null range check
	 IF( r'LENGTH = 0) THEN        -- right input is of null range
    	      ASSERT false
	      REPORT " --- left input has null range "
	      SEVERITY ERROR;
              return(true);
         END IF;
	-- synopsys translate_on        
	-- input are not null so sign extend them to the same length
        -- Convert to bit_vector for comparison to allow any length input vector.
        vl := To_BitVector ( l, IntegerBitLength, SrcRegMode );
 	vr := SignExtend(r, IntegerBitLength, r'LEFT, SrcRegMode);
	IF (SrcRegMode = TwosComp) THEN
        	return (NOT (LessThan_TwosComp(vl, vr)));
        ELSE
		return (NOT (LessThan_Unsigned(vl, vr)));
	END IF;
     END RegGreaterThanOrEqual; 
     -------------------------------------------------------------------------------
     FUNCTION RegGreaterThanOrEqual ( CONSTANT l          : IN bit_vector;
				   CONSTANT r          : IN INTEGER;
  			           CONSTANT SrcRegMode : IN regmode_type
                     -- synopsys synthesis_off
					         	      := DefaultRegMode 
                     -- synopsys synthesis_on
				 ) RETURN bit IS
       VARIABLE vl, vr    : bit_vector(IntegerBitLength - 1 DOWNTO 0);
     BEGIN
        -- synopsys translate_off
	-- Null range check
         IF( l'LENGTH = 0) THEN        -- left input is of null range
    	      ASSERT false
	      REPORT " --- left input has null range "
	      SEVERITY ERROR;
              return('0');
         END IF;
	-- synopsys translate_on        
	-- input are not null so sign extend them to the same length
        -- Convert to bit_vector for comparison to allow any length input vector.
 	vl := SignExtend(l, IntegerBitLength, l'LEFT, SrcRegMode);
        vr := To_BitVector ( r, IntegerBitLength, SrcRegMode );

	IF (SrcRegMode = TwosComp) THEN
        	return( To_Bit_loc (NOT ( LessThan_TwosComp(vl, vr))));
        ELSE
		return( To_Bit_loc (NOT (LessThan_Unsigned(vl, vr))));
	END IF;
    END RegGreaterThanOrEqual; 
     -------------------------------------------------------------------------------
     FUNCTION RegGreaterThanOrEqual ( CONSTANT l          : IN INTEGER;
				   CONSTANT r          : IN bit_vector;
  			           CONSTANT SrcRegMode : IN regmode_type
                     -- synopsys synthesis_off
					         	      := DefaultRegMode 
                     -- synopsys synthesis_on
				 ) RETURN bit IS
       VARIABLE vl, vr    : bit_vector(IntegerBitLength - 1 DOWNTO 0);
     BEGIN
        -- synopsys translate_off
	-- Null range check
         IF( r'LENGTH = 0) THEN        -- left input is of null range
    	      ASSERT false
	      REPORT " --- left input has null range "
	      SEVERITY ERROR;
              return('1');
         END IF;
	-- synopsys translate_on        
	-- input are not null so sign extend them to the same length
        -- Convert to bit_vector for comparison to allow any length input vector.
        vl := To_BitVector ( l, IntegerBitLength, SrcRegMode );
 	vr := SignExtend(r, IntegerBitLength, r'LEFT, SrcRegMode);

	IF (SrcRegMode = TwosComp) THEN
        	return( To_Bit_loc( NOT(  LessThan_TwosComp(vl, vr))));
        ELSE
		return( To_Bit_loc( NOT (LessThan_Unsigned(vl, vr))));
	END IF;
    END RegGreaterThanOrEqual; 
     -- ----------------------------------------------------------------------------
     --     Function Name : RegGreaterThanOrEqual
     --
     --     Overloading   : Input parameter TYPEs.
     --    
     --     Purpose       : Compute a greater-than-or-equal relation for std_logic_vectors
     --     
     --     Parameters    : l       - input std_logic_vector | INTEGER
     --                     r       - input std_logic_vector | INTEGER
     --                     SrcRegMode - input regmode_type, indicating the format of
     --                               the std_logic_vector operands (l,r).
     --                               Default is TwosComp.
     --     
     --     Result        : BOOLEAN | std_ulogic
     --
     --     NOTE          : The operands may be of any length, and may be different
     --                     lengths. 
     --
     --                     Overloading not defined for both inputs of INTEGER type.
     --
     --                     Any time the comparison reaches an index that has an 'X' as an
     --                     array element, the comparison is deemed indeterminate and will 
     --                     return false in case of boolean and '0' incase of std_ulogic for
     --                     synthesis purposes.
     --
     --     Use           : 
     --                      VARIABLE a, b : std_logic_vector ( 7 DOWNTO 0 );
     --                      IF ( RegGreaterThanOrEqual ( a, b, TwosComp)   )  THEN 
     --     
     --     See Also      : RegLessThan, RegLessThanOrEqual, RegGreaterThan, 
     --                     RegGreaterThanOrEqual.
     -------------------------------------------------------------------------------
     FUNCTION RegGreaterThanOrEqual  ( CONSTANT l          : IN std_logic_vector;
				CONSTANT r          : IN std_logic_vector;
				CONSTANT SrcRegMode : IN regmode_type 

                     -- synopsys synthesis_off
							      := DefaultRegMode 
                     -- synopsys synthesis_on
				 ) RETURN std_ulogic IS
       CONSTANT resltlen : INTEGER := MAXIMUM (l'LENGTH, r'LENGTH);
       VARIABLE vl, vr   : STD_LOGIC_VECTOR (resltlen - 1 DOWNTO 0);
     BEGIN
        -- synopsys translate_off
	-- Null range check
	IF ( (l'LENGTH = 0) AND (r'LENGTH = 0) ) THEN   
	      ASSERT false 
	      REPORT "  --- Both left and right vectors have null range "
	      SEVERITY ERROR;
              return( '0');
         ELSIF( l'LENGTH = 0) THEN        -- left input is of null range
    	      ASSERT false
	      REPORT " --- left input has null range "
	      SEVERITY ERROR;
              return('0');

         ELSIF( r'LENGTH = 0) THEN        -- right  input is of null range
	      ASSERT false
	      REPORT " --- right input has null range "
	      SEVERITY ERROR;
              RETURN ('1');
         END IF;
	-- synopsys translate_on        
 	-- input are not null so sign extend them to the same length
	vl := SignExtend(l, resltlen, l'LEFT, SrcRegMode);
	vr := SignExtend(r, resltlen, r'LEFT, SrcRegMode);

	IF (SrcRegMode = TwosComp) THEN
        	return( To_StdULogic_loc (LessThanOrEqual_TwosComp(vr, vl)));
        ELSE
		return( To_StdULogic_loc (LessThanOrEqual_Unsigned(vr, vl)));
	END IF;
    END RegGreaterThanOrEqual; 
     -----------------------------------------------------------------------------
     FUNCTION RegGreaterThanOrEqual    ( CONSTANT l          : IN std_logic_vector;
				   CONSTANT r          : IN std_logic_vector;
 			           CONSTANT SrcRegMode : IN regmode_type
                     -- synopsys synthesis_off
							      := DefaultRegMode 
                     -- synopsys synthesis_on
				 ) RETURN BOOLEAN IS
       CONSTANT resltlen : INTEGER := MAXIMUM (l'LENGTH, r'LENGTH);
       VARIABLE vl, vr   : STD_LOGIC_VECTOR (resltlen - 1 DOWNTO 0);
     BEGIN
        -- synopsys translate_off
	-- Null range check
	IF ( (l'LENGTH = 0) AND (r'LENGTH = 0) ) THEN   
	      ASSERT false 
	      REPORT "  --- Both left and right vectors have null range "
	      SEVERITY ERROR;
              return( false);
         ELSIF( l'LENGTH = 0) THEN        -- left input is of null range
    	      ASSERT false
	      REPORT " --- left input has null range "
	      SEVERITY ERROR;
              return(false);

         ELSIF( r'LENGTH = 0) THEN        -- right  input is of null range
	      ASSERT false
	      REPORT " --- right input has null range "
	      SEVERITY ERROR;
              RETURN (true);
         END IF;
	-- synopsys translate_on        
 	-- input are not null so sign extend them to the same length
	vl := SignExtend(l, resltlen, l'LEFT, SrcRegMode);
	vr := SignExtend(r, resltlen, r'LEFT, SrcRegMode);

	IF (SrcRegMode = TwosComp) THEN
        	return( LessThanOrEqual_TwosComp(vr, vl));
        ELSE
		return( LessThanOrEqual_Unsigned(vr, vl));
	END IF;
    END RegGreaterThanOrEqual; 
     -- -----------------------------------------------------------------------------
     FUNCTION RegGreaterThanOrEqual ( CONSTANT l          : IN std_logic_vector;
				   CONSTANT r          : IN INTEGER;
			     CONSTANT SrcRegMode : IN regmode_type
                     -- synopsys synthesis_off
						      := DefaultRegMode 
                     -- synopsys synthesis_on
				 ) RETURN BOOLEAN IS
	VARIABLE vl, vr    : std_logic_vector(IntegerBitLength - 1 DOWNTO 0);
     BEGIN
	-- synopsys translate_off
	-- Null range check
	 IF( l'LENGTH = 0) THEN        -- left input is of null range
    	      ASSERT false
	      REPORT " --- left input has null range "
	      SEVERITY ERROR;
              return(false);
         END IF;
	-- synopsys translate_on        
	-- input are not null so sign extend them to the same length
        -- Convert to std_logic_vector for comparison to allow any length input vector.
        vr := To_StdLogicVector ( r, IntegerBitLength, SrcRegMode );
 	vl := SignExtend(l, IntegerBitLength, l'LEFT, SrcRegMode);

	IF (SrcRegMode = TwosComp) THEN
        	return( LessThanOrEqual_TwosComp(vr, vl));
        ELSE
		return( LessThanOrEqual_Unsigned(vr, vl));
	END IF;
    END RegGreaterThanOrEqual; 
     -------------------------------------------------------------------------------
     FUNCTION RegGreaterThanOrEqual ( CONSTANT l          : IN INTEGER;
				   CONSTANT r          : IN std_logic_vector;
  			           CONSTANT SrcRegMode : IN regmode_type
                     -- synopsys synthesis_off
					         	      := DefaultRegMode 
                     -- synopsys synthesis_on
				 ) RETURN BOOLEAN IS
       VARIABLE vl, vr    : std_logic_vector(IntegerBitLength - 1 DOWNTO 0);
     BEGIN
	-- synopsys translate_off
	-- Null range check
	 IF( r'LENGTH = 0) THEN        -- right input is of null range
    	      ASSERT false
	      REPORT " --- left input has null range "
	      SEVERITY ERROR;
              return(true);
         END IF;
	-- synopsys translate_on        
	-- input are not null so sign extend them to the same length
        -- Convert to std_logic_vector for comparison to allow any length input vector.
        vl := To_StdLogicVector ( l, IntegerBitLength, SrcRegMode );
 	vr := SignExtend(r, IntegerBitLength, r'LEFT, SrcRegMode);

	IF (SrcRegMode = TwosComp) THEN
        	return( LessThanOrEqual_TwosComp(vr, vl));
        ELSE
		return( LessThanOrEqual_Unsigned(vr, vl));
	END IF;
    END RegGreaterThanOrEqual; 
     -------------------------------------------------------------------------------
     FUNCTION RegGreaterThanOrEqual ( CONSTANT l          : IN std_logic_vector;
				   CONSTANT r          : IN INTEGER;
  			           CONSTANT SrcRegMode : IN regmode_type
                     -- synopsys synthesis_off
					         	      := DefaultRegMode 
                     -- synopsys synthesis_on
				 ) RETURN std_ulogic IS
       VARIABLE vl, vr    : std_logic_vector(IntegerBitLength - 1 DOWNTO 0);
     BEGIN
        -- synopsys translate_off
	-- Null range check
         IF( l'LENGTH = 0) THEN        -- left input is of null range
    	      ASSERT false
	      REPORT " --- left input has null range "
	      SEVERITY ERROR;
              return('0');
         END IF;
	-- synopsys translate_on        
	-- input are not null so sign extend them to the same length
        -- Convert to std_logic_vector for comparison to allow any length input vector.
 	vl := SignExtend(l, IntegerBitLength, l'LEFT, SrcRegMode);
        vr := To_StdLogicVector ( r, IntegerBitLength, SrcRegMode );

	IF (SrcRegMode = TwosComp) THEN
        	return( To_StdULogic_loc (LessThanOrEqual_TwosComp(vr, vl)));
        ELSE
		return( To_StdULogic_loc (LessThanOrEqual_Unsigned(vr, vl)));
	END IF;
    END RegGreaterThanOrEqual; 
     -------------------------------------------------------------------------------
     FUNCTION RegGreaterThanOrEqual ( CONSTANT l          : IN INTEGER;
				   CONSTANT r          : IN std_logic_vector;
  			           CONSTANT SrcRegMode : IN regmode_type
                     -- synopsys synthesis_off
					         	      := DefaultRegMode 
                     -- synopsys synthesis_on
				 ) RETURN std_ulogic IS
       VARIABLE vl, vr    : std_logic_vector(IntegerBitLength - 1 DOWNTO 0);
     BEGIN
        -- synopsys translate_off
	-- Null range check
         IF( r'LENGTH = 0) THEN        -- left input is of null range
    	      ASSERT false
	      REPORT " --- left input has null range "
	      SEVERITY ERROR;
              return('1');
         END IF;
	-- synopsys translate_on        
	-- input are not null so sign extend them to the same length
        -- Convert to std_logic_vector for comparison to allow any length input vector.
        vl := To_StdLogicVector ( l, IntegerBitLength, SrcRegMode );
 	vr := SignExtend(r, IntegerBitLength, r'LEFT, SrcRegMode);

	IF (SrcRegMode = TwosComp) THEN
        	return( To_StdULogic_loc (LessThanOrEqual_TwosComp(vr, vl)));
        ELSE
		return( To_StdULogic_loc (LessThanOrEqual_Unsigned(vr, vl)));
	END IF;
    END RegGreaterThanOrEqual; 
     -- ----------------------------------------------------------------------------
     --     Function Name : RegGreaterThanOrEqual
     --
     --     Overloading   : Input parameter TYPEs.
     --    
     --     Purpose       : Compute a greater-than-or-equal relation for std_ulogic_vectors
     --     
     --     Parameters    : l       - input std_ulogic_vector | INTEGER
     --                     r       - input std_ulogic_vector | INTEGER
     --                     SrcRegMode - input regmode_type, indicating the format of
     --                               the std_ulogic_vector operands (l,r).
     --                               Default is TwosComp.
     --     
     --     Result        : BOOLEAN | std_ulogic
     --
     --     NOTE          : The operands may be of any length, and may be different
     --                     lengths. 
     --
     --                     Overloading not defined for both inputs of INTEGER type.
     --
     --                     Any time the comparison reaches an index that has an 'X' as an
     --                     array element, the comparison is deemed indeterminate and will 
     --                     return false in case of boolean and '0' incase of std_ulogic for
     --                     synthesis purposes.
     --
     --     Use           : 
     --                      VARIABLE a, b : std_ulogic_vector ( 7 DOWNTO 0 );
     --                      IF ( RegGreaterThanOrEqual ( a, b, TwosComp)   )  THEN 
     --     
     --     See Also      : RegLessThan, RegLessThanOrEqual, RegGreaterThan, 
     --                     RegGreaterThanOrEqual.
     -------------------------------------------------------------------------------
     FUNCTION RegGreaterThanOrEqual  ( CONSTANT l          : IN std_ulogic_vector;
				CONSTANT r          : IN std_ulogic_vector;
				CONSTANT SrcRegMode : IN regmode_type 

                     -- synopsys synthesis_off
							      := DefaultRegMode 
                     -- synopsys synthesis_on
				 ) RETURN std_ulogic IS
       CONSTANT resltlen : INTEGER := MAXIMUM (l'LENGTH, r'LENGTH);
       VARIABLE vl, vr   : STD_ULOGIC_VECTOR (resltlen - 1 DOWNTO 0);
     BEGIN
        -- synopsys translate_off
	-- Null range check
	IF ( (l'LENGTH = 0) AND (r'LENGTH = 0) ) THEN   
	      ASSERT false 
	      REPORT "  --- Both left and right vectors have null range "
	      SEVERITY ERROR;
              return( '0');
         ELSIF( l'LENGTH = 0) THEN        -- left input is of null range
    	      ASSERT false
	      REPORT " --- left input has null range "
	      SEVERITY ERROR;
              return('0');

         ELSIF( r'LENGTH = 0) THEN        -- right  input is of null range
	      ASSERT false
	      REPORT " --- right input has null range "
	      SEVERITY ERROR;
              RETURN ('1');
         END IF;
	-- synopsys translate_on        
 	-- input are not null so sign extend them to the same length
	vl := SignExtend(l, resltlen, l'LEFT, SrcRegMode);
	vr := SignExtend(r, resltlen, r'LEFT, SrcRegMode);

	IF (SrcRegMode = TwosComp) THEN
        	return( To_StdULogic_loc (LessThanOrEqual_TwosComp(vr, vl)));
        ELSE
		return( To_StdULogic_loc (LessThanOrEqual_Unsigned(vr, vl)));
	END IF;
    END RegGreaterThanOrEqual; 
     -----------------------------------------------------------------------------
     FUNCTION RegGreaterThanOrEqual    ( CONSTANT l          : IN std_ulogic_vector;
				   CONSTANT r          : IN std_ulogic_vector;
 			           CONSTANT SrcRegMode : IN regmode_type
                     -- synopsys synthesis_off
							      := DefaultRegMode 
                     -- synopsys synthesis_on
				 ) RETURN BOOLEAN IS
       CONSTANT resltlen : INTEGER := MAXIMUM (l'LENGTH, r'LENGTH);
       VARIABLE vl, vr   : STD_ULOGIC_VECTOR (resltlen - 1 DOWNTO 0);
     BEGIN
        -- synopsys translate_off
	-- Null range check
	IF ( (l'LENGTH = 0) AND (r'LENGTH = 0) ) THEN   
	      ASSERT false 
	      REPORT "  --- Both left and right vectors have null range "
	      SEVERITY ERROR;
              return( false);
         ELSIF( l'LENGTH = 0) THEN        -- left input is of null range
    	      ASSERT false
	      REPORT " --- left input has null range "
	      SEVERITY ERROR;
              return(false);

         ELSIF( r'LENGTH = 0) THEN        -- right  input is of null range
	      ASSERT false
	      REPORT " --- right input has null range "
	      SEVERITY ERROR;
              RETURN (true);
         END IF;
	-- synopsys translate_on        
 	-- input are not null so sign extend them to the same length
	vl := SignExtend(l, resltlen, l'LEFT, SrcRegMode);
	vr := SignExtend(r, resltlen, r'LEFT, SrcRegMode);

	IF (SrcRegMode = TwosComp) THEN
        	return( LessThanOrEqual_TwosComp(vr, vl));
        ELSE
		return( LessThanOrEqual_Unsigned(vr, vl));
	END IF;
    END RegGreaterThanOrEqual; 
     -- -----------------------------------------------------------------------------
     FUNCTION RegGreaterThanOrEqual ( CONSTANT l          : IN std_ulogic_vector;
				      CONSTANT r          : IN INTEGER;
 				      CONSTANT SrcRegMode : IN regmode_type
                     -- synopsys synthesis_off
						      := DefaultRegMode 
                     -- synopsys synthesis_on
				 ) RETURN BOOLEAN IS
	VARIABLE vl, vr    : std_ulogic_vector(IntegerBitLength - 1 DOWNTO 0);
     BEGIN
	-- synopsys translate_off
	-- Null range check
	 IF( l'LENGTH = 0) THEN        -- left input is of null range
    	      ASSERT false
	      REPORT " --- left input has null range "
	      SEVERITY ERROR;
              return(false);
         END IF;
	-- synopsys translate_on        
	-- input are not null so sign extend them to the same length
        -- Convert to std_ulogic_vector for comparison to allow any length input vector.
        vr := To_StdULogicVector ( r, IntegerBitLength, SrcRegMode );
 	vl := SignExtend(l, IntegerBitLength, l'LEFT, SrcRegMode);

	IF (SrcRegMode = TwosComp) THEN
        	return( LessThanOrEqual_TwosComp(vr, vl));
        ELSE
		return( LessThanOrEqual_Unsigned(vr, vl));
	END IF;
    END RegGreaterThanOrEqual; 
    -------------------------------------------------------------------------------
    FUNCTION RegGreaterThanOrEqual (CONSTANT l          : IN INTEGER;
				    CONSTANT r          : IN std_ulogic_vector;
  			            CONSTANT SrcRegMode : IN regmode_type
                     -- synopsys synthesis_off
						      := DefaultRegMode 
                     -- synopsys synthesis_on
 				  ) RETURN BOOLEAN IS
       VARIABLE vl, vr    : std_ulogic_vector(IntegerBitLength - 1 DOWNTO 0);
     BEGIN
	-- synopsys translate_off
	-- Null range check
	 IF( r'LENGTH = 0) THEN        -- right input is of null range
    	      ASSERT false
	      REPORT " --- left input has null range "
	      SEVERITY ERROR;
              return(true);
         END IF;
	-- synopsys translate_on        
	-- input are not null so sign extend them to the same length
        -- Convert to std_ulogic_vector for comparison to allow any length input vector.
        vl := To_StdULogicVector ( l, IntegerBitLength, SrcRegMode );
 	vr := SignExtend(r, IntegerBitLength, r'LEFT, SrcRegMode);

	IF (SrcRegMode = TwosComp) THEN
        	return( LessThanOrEqual_TwosComp(vr, vl));
        ELSE
		return( LessThanOrEqual_Unsigned(vr, vl));
	END IF;
    END RegGreaterThanOrEqual; 
    -------------------------------------------------------------------------------
    FUNCTION RegGreaterThanOrEqual (CONSTANT l          : IN std_ulogic_vector;
 				    CONSTANT r          : IN INTEGER;
  			            CONSTANT SrcRegMode : IN regmode_type
                     -- synopsys synthesis_off
						      := DefaultRegMode 
                     -- synopsys synthesis_on
				  ) RETURN std_ulogic IS
       VARIABLE vl, vr    : std_ulogic_vector(IntegerBitLength - 1 DOWNTO 0);
     BEGIN
        -- synopsys translate_off
	-- Null range check
         IF( l'LENGTH = 0) THEN        -- left input is of null range
    	      ASSERT false
	      REPORT " --- left input has null range "
	      SEVERITY ERROR;
              return('0');
         END IF;
	-- synopsys translate_on        
	-- input are not null so sign extend them to the same length
        -- Convert to std_ulogic_vector for comparison to allow any length input vector.
 	vl := SignExtend(l, IntegerBitLength, l'LEFT, SrcRegMode);
        vr := To_StdULogicVector ( r, IntegerBitLength, SrcRegMode );

	IF (SrcRegMode = TwosComp) THEN
        	return( To_StdULogic_loc (LessThanOrEqual_TwosComp(vr, vl)));
        ELSE
		return( To_StdULogic_loc (LessThanOrEqual_Unsigned(vr, vl)));
	END IF;
    END RegGreaterThanOrEqual; 
    -----------------------------------------------------------------------------
    FUNCTION RegGreaterThanOrEqual (CONSTANT l          : IN INTEGER;
				    CONSTANT r          : IN std_ulogic_vector;
  			            CONSTANT SrcRegMode : IN regmode_type
                     -- synopsys synthesis_off
						      := DefaultRegMode 
                     -- synopsys synthesis_on
 				  ) RETURN std_ulogic IS
       VARIABLE vl, vr    : std_ulogic_vector(IntegerBitLength - 1 DOWNTO 0);
     BEGIN
        -- synopsys translate_off
	-- Null range check
         IF( r'LENGTH = 0) THEN        -- left input is of null range
    	      ASSERT false
	      REPORT " --- left input has null range "
	      SEVERITY ERROR;
              return('1');
         END IF;
	-- synopsys translate_on        
	-- input are not null so sign extend them to the same length
        -- Convert to std_ulogic_vector for comparison to allow any length input vector.
        vl := To_StdULogicVector ( l, IntegerBitLength, SrcRegMode );
 	vr := SignExtend(r, IntegerBitLength, r'LEFT, SrcRegMode);

	IF (SrcRegMode = TwosComp) THEN
        	return( To_StdULogic_loc (LessThanOrEqual_TwosComp(vr, vl)));
        ELSE
		return( To_StdULogic_loc (LessThanOrEqual_Unsigned(vr, vl)));
	END IF;
    END RegGreaterThanOrEqual; 


end synth_regpak;



