`ifdef encrypted_0in
`protected_0in
ze74c34e226135848fe16db9ffd31815111b6d7fb642c521a3f628cf6da949865580b22efd062a7
ze90adae0e65e66a2c36a587d0a790699161455169ed55a01f2084f11770a774ec4c588039b380f
z6de9c5084882a40b79a175f5c2114b2b6d78b070cb806e1c0aa9258297f4687ab308bc470f0040
zb0b1de382961eeeaf2e279e1462520fc31c119af8f2b214846f56c2b3cd2eadbe4099496abff18
z15cec83ec4a77b868344aa20ba7360908f5c0de2a79abf8b3534b883bb12180f68b5d4beb444cf
z3fba8f13afb0abfe8fcc4294810f75afe452434d2d0f1166236c82f76edf1e12979f04bc35693e
z32ae028996dd85737a8f5adc1ebb94f39c940246e887647b64782cd7ab429b0544c173176cede7
z01dfb26b1f73408344a52b7e1f117f12bb9c8077b34876c2e6fdc085981637012dc9754765e1a9
zc512ce062e0b8fb16a214591f5c81e1353b900a611fe1f4886b57940b41b7f2ce99a7b84b04b90
z916f717e73bd10589c81e207ed77ec660a8cbed5b487fa50acde1b055c8870bd8676023f21ddcf
z9c98cc47cfa2d654ff1365d1f45035a045a66c5dfa82790502623b57a3af03bf0f0c0d35b51558
zb8b5f2d29acf03737a9ca2a053b7a8f06800d50b465c41b30eb585f62f3d0c2c5a43bc54b3c9b8
z81acf2d405b3b2356c7277371175910889302fc7dc38870232426d1efea28b5d258bcaa0f177b1
zc52cddceff94a138a0a137b7dc25b3fe1989f30341fc446d2211451d70bd3bbf5bbfee546509c5
z26e02b5a0f51127073ec2b77ced81a0703594af64f3c2f07171b2c88744c0bc7fe92c155aad2a5
z17dbc975e4de99a315ee01a21f50971e97a55338d08788a1b97a2d3c49a8e6368101e4ec68939c
z98eddf0754a166ed5935f229a7da295f3e081c23877f04b7197c10b9aee8daefd578029c77b9ff
z66fcd8e9c95d80e7c8bf3e2b15322c022ced66b45e03e2f48439bf7dfbbad809f516a56d486e38
z2a783289af1c628a034ec9d251f3b978eea89bda0f8e76acc0018aeb461ec7af18217e03b2dedd
z2da170ce8de08622b3ce1ba248f1a812c10b073f128ec24d126154db3a3c9bb4bd4a6c69e7b4eb
zed63929264f8a4d11a0fe17beca835dc987761137b995ab9ff5242a30c57c18f2e2a4375ab931f
za922db31bf9a08e656b9c816eaec8c24e19379e9e1a24ef382fa0c7df565038e7ab71be007777d
zc029cd9d32b05de4d45d4896fdfa9c41283ea5d0af898b1b5f7dc636be558d37709c2233b0f80e
ze9e7ee2c3784a4e69afa2df23f89ac8f27a326552b5d6325e93b16763e3974c22f008337092ade
z7313e1dfa705d54fff276030f16af20e602c7d7b0a3f714b0cbce8a1f6c5e9f1cfefb236bc78c5
zcd3c43cb50c4d83321e10ce4693d8b3a2f936bd6512281969a317a914544cefe1c95ab1ceb2fa6
zc0809b96e39a2f8a4750e6afadf07f058fe25ca48accc8bf0f00d57988d0f114377c1731d413c7
z40b89b4890ade91d37ae8b990c2ddbfb0160cef122fde3ade96cf013319979da1f8d8a792f26a5
z459841097fd3d3ae02461bb2446944dfdaa8f3b2446e5282a28d21d467622e2513fbc3cbaf56c4
z1e71542c01a97cd29653910c027d62ac374b523f81acaaadff9b9a670a7983149293d98ce63ede
z8a14ff1c8b7849908e04938ca3063aa861f38604423c3407f2d6917a33187bd6d0c97482e43d8e
z34f454d0cbbdb3d987fa47e936280d345e06b0e0ac2d1034717e7c766625ee013cedc00c67e3d7
z867dc2baff74709512921e85b62bc23623c9a39dcb4e9b8ad6fbccbf18506ab33c69fcddd18300
zd77acf123e8a556aa91ca51c29df69f86c3af24a6d0cbc43016eb9cedd4b0bfb030ed345f92a70
zecf93969bc4ad89c39c52f139193ee82af4f64eed6fea89fd370b8053bfe7a9a617fd415a93c77
zbac82123b0816b5034e4b89c34431a60750f4128d7d3a2178861029fdf9bff19f490c163c69e2a
z92b3abefe1133837c90583b47a64490241dcc2dd6a23cb90144ecc3cf3ce81ab10030b53732f0d
z4b4161d9ffe44af47115ab2cf11f7da2cd1d59a930c2347b0a38404fef502be9ce6901476709a2
z8a932370feee928e054851e1253d221846ce1a38658b9ed025d48b90ece1f0b96d6d5639d74f92
zc76bb4908eed366a606c073db81768b7638932c9a41c02124ac32f5248353cd2dfc7b9e836f132
z2aae8d69222f18f2c87ca29ae19da65f666c77a9d95810445eab809eeca27167bcb34e7d372df4
zbd3352ea0fd06c1e2306f1f762cab79dc0ccbfbdb67dba424f4d605f67fe66e656bc9773655dff
z7fb3bb8eaaefd000580befacff1bd994776a507fa3b847ab472d7f3eaf42db71465d214668024b
z71beebb21b08d0767b514e2c06e575140c8f7c80b655c664eb5074a3c6fa60490ba9edf1465d25
z232bd79f331830272ed83a70ec640fa8695c208883321d34aef561b00649d5122b1eeffe88ede6
za03b3332ebac60a26d68888f653445e8f205c9aaa599584e9b61b1bd838c9910a168f256b7b91e
z306c7eb7db78b499b0b8e61bd73776124da763352d2a6964d8a0ae33e9ba8757b2c058e71b2507
zc73c00c08a370f16ff04abfc306b588b9a388f6d858a25d8bff1d45f1a3643bef09e7cbd904a14
z45941297bdd27a3e6400383c5afb8e32f7a3057b80a197fe0550fdc0b77e8cbc453632af4ee215
z874638a8e85fca5da6964e87fde90d85844149757508433bbf0a16b9676d8a7f8ac7c0906ad288
z22e6e64232f4fa17954bce68a2ce22ff771053b5c4be9d6b0e317df6a91e0bbb2db8d0c9360732
zccd65e465be967c491a28faa30e88c432bff2214380111ad07af31c9554166d46641a862e5277d
zd4ff0b1a44e8eea52715027928aa0dd92d009d64e147e8c3f020860401a7818bc3784df78ead6d
z4314833559ae09c714367edb4c187711940597451deb5478222bf652b2a12ad9e069f4a17caa6b
ze7b6868d2c96010f71a0677a99534c283f3318922fe73844166e3924385dcb49d117620cbcc2f0
z1b124350da7586ce906414e2d07341edf2f4c96d8061bd79de89a8ee0d49767b278337caf1f925
z7061e96a1dee2c792c1914c4cd425a7c0c9b4bad9bd4f7ed9518e7ad698dcd80dfbc92d55355b5
z11f597762fecb5be2bd12a2e3d427698559fe71c49e92be088ac39d1d9ce9b55c96164c04fa456
z50cd9ed9ed1765c5edb34542c8b39b5d42e199205b67cdc1d93f1431ae107e0bb2bcd13fc20ad1
z5b4e5578c46ac41e590918cb797cb66546dec842406ad73de12f1d3034ff3f13b0601d6e204a6a
zbd2f4699598fa0a07f8508f9b9a3702ae5cd2e895cc698f99808233c803ab60d7fa41c99933643
z73a8e2fb156f2ae42fc238e543a11cfaf82b34938bf4a22e5347c420baf37204abac00ba569611
z24e44c1260f8cc1d549367a1332d6c3e058b555f94df24308682879af51545fd87729d4826e0a2
zca012158550c659d570a883ddb1f4c4888321acb282844e850d30c38df126df99f455fc261271c
zad59e3927a5d8501964ee17737defbfae60d8bd7e0da659e19d556d83af1b944fa7a47ee7ad765
zfbe06a1766fde8017896357a4f8c67372a93cc55f8e81a9ea7a1da844278852eed9bc65ff8472a
zae2e9a615f901678f309b36d6bd4ba976ebfca2ffb85565185d1c960698955a463b034f4f78827
z6f204169c5401967ce3c7b98d7820c9506b5ad2e9f34d2ed673153d279997db1e87a763acf731a
z3d260d8267fc2f4a2b84e515cb9a358a3be8dc64e603602a812b42004b4b5f2660cbf90b282a93
z2f500b865cca864687c112458f91ed427e4f47c8983092545b747dd66671b039499ac7ef5735df
z8b9cc597a3bc8ef41cbeebf99c298e460a75f677f60446e09e4fc60ca7267f3491c4a76d1788ae
z3d4da7979dfea1b24abf107beabd0145f006ff96e03c75b9c389b0095382879a9aadd74e15eb59
z3dd875bc7b6e3410b00528e2a6f49878d6aa09573513f978c1cdfdacce2a01af2f37e61f85bab4
z6f543bdcb2f080a4b5015bb4becb660afca13b5700978294f5a896c481042974ab3f3facc7a733
zcf357b9bfa2084c7e6d7b1c2c3d20d4b0bae688552ea5e787eb6fd80895fe8940952706fb109f7
ze2e08fcc2a55b81c0d5158204b9573d19626fed7b1192d85de2fbbdc5c6e40328a902d99a49be6
z91ec22108ceb5611331497fb20c1165a92b065d7817fa660d27bf229bd5d4151d46dfeca11caba
z1b220584bc703fe84df14321eb769c6264b84516f134ae239292e89758c3693e2db50169f51c65
z8589e077194ad925b91d7c400aef4fbd9095bdd806535eac21d2524b2fb3287e6c478e8bab8df3
zf999797e1846f3036a41d4f3c31a27df58219e800cb07c9fe7c3f9b733ce9c6c40a1d404c416d1
zd5c62235ed776a4e118e198264a76d526f50384b62db64342f3bc1842594a1327cf53f5aa6cfe7
z1316471a4d5264fd2b2fbda523b989030508e27299c2f5e55ba1c8f790249d5fdc9659cb005c29
zed2eae0dfa296f401d689f241bfdc3627a7c934ccf1f6c5a8947f1265dccaebd54d47ea9c289f7
z2e896ccc42b22f385ca8b75cb543aed8ca168c790759ab0717fe068c24682daa7c9c8c8f75f5b5
z0bb5980391b77105dd4060af99ef9e73156c3d38959860fe24c7873b76f651f0a4262068b33934
z778f892315d1b4651fb6e1bed0a66f9c0c3ea1706c891bfc371eecc2117acb668ab44bf45fa856
z7fc038a76bbf3cf268b7dcecf99d78d541ee44a69b1761caae376c6803ca2bdaefe80c937c1f6c
zce37098cdef53f052512e2cce300b3146ba5453bd224fa150e4751f62f61bc1630f74808887f50
zef3fcc9220fcffe432720d48ec9d1884a10b4128accfb5ed42ea49d572819cb52a894486f4584d
z535264995fb06f9c408c557c1f825af683d5e698e939c6ef4cdffdc403ee547edb2bfb05e01909
z6a82763da8be206919bd118c1a497b04e3437821ef98a569bbff4a19c55dc9f32e30591ad06200
z96e4d563ca7fa0399f9188c1eba94ea7ad2ef48bd86ab52989ee850478c5374efb2eba24fc6a50
zc87396d8f551c3a1e4eb4e066c8a16f2b31d5fbba1c82ea318aae5b0e3494e22dfa56372dc32d8
z4082b2bfa3d53d55034631ce8cfb9f927666d9177cc30b1fd02d8a5d1e656166abde09e9bd563a
z19617debaa104458ab3ae426a6b2c94b069ec2e7dc412a5b48886d61caee0d9ab48cf9fdf24001
za700b2596097352b2b017ea1623a67833a3425ac3e4f2960e1f6006bc6d0f4e93dbc644b0baf63
zd55684703e0f701d11b39c57620cfe9fe1015eb660f5f4831518c8c7899baab7a917ac260b9c47
z5ed11dbb711fb10b0ef139ee8a153f48dd1ae0364be0746ca1bcda569e35efac270c16407c5a30
z6df2f3b0fc2012aaef62e324d0a94bcf0354851a6dda9daf3d5a4af4bc04f423877046290b1baf
z42e1afcf5a67657f7b348f2b0d3c830ccc62644aaf58494b1aac5127c9f56d1d52010c65bd9f24
zb07c366a3daeac4c5a824545cb3e1ca3c832ab7d3d421033a635b2bdc4c5c3b64fcb5621009a86
z2aff039b3c7f7aecf3fc424548a8b28b7ce485f1fb7caf6cbe00362f1003f907f7c05ab01c64e2
z248d5a210b0d563561c3901d10ae696ed082a05faae98aee7f2f2f2c2e3c9ed35f574ccd65c53e
z917b37622c0525cf1a0cd661e699cc11370373e6404b3ef3fdc52eb202f4bed12b03d90243b0f3
zbdab4b64f97536e79a5e171bd7c2d4f25139fd36d64bee46d0a75e28dc147d36ea927a4cb81eeb
zb87fa6a4c60904952e2f8a0355569962b5004f4b78bbbecc6d856e5761fe4bf79d52f364e767eb
ze71ab21046fc5eb526c767b0358a9d1523d7d4bde898015c105198efbd89bf800e621e0e591bee
z57b47adba15d49859060823f6d38b9296fe5680528623b34806c651ec5448b18799636e4364b3b
zbcf09ef837fae97f2a2c4a730cde93f16622ef9f4301fde3468468f624e2338c45d58c434db1d8
zd640ca35aa130a7eecc0d5a667bed5fe462c06ff8c24cd83db27d6c26fd49dcd14f633555a90be
zf4568ac01a98f37d90e98d945cc086d11fe83762604ec8cb71159725e6dd4a4713f4d9c2e342e9
zf98fdc69d5a15e974354c6f47497efc7851beb805467c1b69e00489a454bf4d0850db14799242a
z04ef72625d158d8807904e41a311a29c89890214dfe7cb0693fbe012b4872ba084225ed86d36e9
zbbb77004be6b8e6a992b0e8fda0a331bb52412fd26ca0e9e3eb04a57f13ef4fb4d0fe1820595b2
z738d40426753ef78b19f940a52c99af2b1fc22f18dfcee2fcc0081b0feda341d341dc4c5fe91bd
z76e800ecbde346d65de89dea8876f8e982768d024014bee913d25785a0b8a33cd53b599dcd6430
z232e6c11b4a31cde9b51802fc9dadd057ea11b41dc8b6f014ab5bd4d2bf4668b39ad59c89f5306
z793d3bf9e9d739fd868ae58475ecc341d577ef2093f34757469de8fa5006ffeff86b746e387103
zb6ff3685cc346e25bbf1d1844d08ee76fc692a22604e8f688ce794d54cf4e69f3102f561b158b6
z3a88c94ca4b91626333b9cf55487942cebf3c8fb498b62213f66c0a202b96d8a565614b8780f00
zb2f6512d3e9bd1c560853b9ae11750179ea591f6acbcb9830ff2d66004372fac7f3a40e1e3e1c8
z130a6a261e3c7f644bce8646d056a3d7d0bd249ee2437ba9d0785383d9b806c4d776c78b2e9399
z1b0ea8e789102c93174f6d138872e7a15d632b592c9ec77795f18f1a2e46fb89fb297928a36ea7
z4758fa36339ec5127e8b2152a440ae330f2087d244dcc58974d6003f1631f04a2802d42572a751
ze5fc69a06548ed52605359e881706ee947a4bfbc0d1e0147c53d8db4bea638fa57abf000ec31ab
zf576f48d45ad8fca8facf728ea6f30d99e5071e2c57c4e52af3a1969ab1e58bcdd6894ec455c45
z196e9eb722557ee04040cbd65337115ecae6e606b2de692e10544e8684a476c12718884d483b98
z9007e9be0b094ca6dcab3ea3b094b385ad9af6b9a69e63a9e2b5fb8b55d6dfb0d5dfc3b1fdeebe
zca29bfb6e2be4f9ce8ff654b1b858c48d21c15501d131f9e0794baebc31732403fdecedfa2e2ba
z6ab2b914c275c5e82839170f6f6bdc3e5f4dd7daa6b789e6efb31baf75e38b60871746282d8b9a
z8181ab0d386f759d141dfa9d848048ae87a78b5d6b59a5bf47ecafd266c729003919ad15f8dd60
z513e1b35d1e229a4dadf2336547c1f90a88bb8fed056c31a1585f9f3a9f8a76b40ed0d515ba68a
zbf17bacafdd2e9e00166f9c55265d6f073602f3a2fe5884592b80ae45bc2dcb90e905b9da63f11
zb625dec1945172109dd5c325dac4812c8e42471deaa72daaad330b3ba5a0b7e4bebb337839fb25
z96bc3188d36592bfe4c6fdcea62802c757ff51edf7babceb648f85423973aa399bdec6e54826ca
zc914c51647d258e2f4305c0940d30352d3749013e430cae3ef7dd720403951816c481be5d9bc9a
zf15fd5797b9645ac4802d93257e90faff3003b874437248979ad5206960e6fa867d38996dde9b3
z74ae6b14f6478e66e8c834f2a96e6bf7e022890a8feb6c9bb2e885b883d23507ba9b4fab1e884d
zb8bdf8fd8ab3561a5e1c526dc8bc53e3b1bd673ea5c0d794967a9f9c7f527888a3019e932387bd
z79418447c2dea2d8376a83bec878cb7f5ae5263ee38b0eb452c67ad08e833c1b99529e264ae883
zc40dedf98ca4c15e8232dedde3b41533be15ff6a0546aafc24b8a52843128ae2851dbd5e231987
zf2fb1fae204ce2896d9528463be95492b8e7260b8f92bb67fc8ed6e2321321de1c137e64494736
z7ab63808213abea42f0db41f08929eaa8225b211d6c9d53927ec95e9216b818ec134c288dc079b
z1ba922d4b00a39cdcc8339d042daaf70f5fb99f7f77d00cbb17a7cb2cd3d81f290a34f2c5575d2
zf549751b05b987947753193d699fd4b790c578da45f7eb02001f73b15939d081becf84646eff98
z67f89951f416b2bfaac646766e76030124809b0af519e171cd88190351915ed59ab2b45c6c2f4f
z88bef4d4714585319f5d820adf8cd388a0b5bb5b6aecdf905d5a3b739d6578e0ef5ab7382256f6
z57c23cc9a95535e38f16b3601a65be76223b9f98215ad13adb90ed26950592f4725f813372406e
z90d27b32baaf0d437a1b0f8904afe4d7f8598d5a317d8b8fe3952293214466fe71a39e5ecda0ca
z0da47efa7a0e2b440d03ca3189ca2d20aeacfbe101811c106a125c706270acb333ffa75a88bfc0
zc4f096fafa727d4051a6e31454c30cbdd398ba27ecdfe1e5b39ebcdef428b862da635bea0fb451
z4176fc0e2a899f5c8a6f31495978a66aabafb57c022b2478d2736cacdae309fb0da71d8e4a627a
zcb93c692854fde0ab5c09bfbcddc8c6da1dec7789b3d5d6e2f5404690544140ad710ccf4098ba7
zc473ddd1852cc142ddc683f249612f3db931864b8bdb2c7a5aaa58089055e2e4f58df68b259906
z8fec396faecd8d0cec5fc60849f43645b6000ed9bf406a2680ee20a513fe94717efb781b961040
z09d223b7df6d64a736eee0c87801bf4cfc558fe0405a5ed87e2a33f1e3a4f7c285d1b157243f7b
za6fff62be4b23a191fc21b3a659f359c18228a7a5efb7b22a713b5b5a50f2650ca02ed8d3db80e
zdb7dce1a5f0838e0c06778fcf2a20895a8a22915d97ad4ae3b8f1166a67f44fb2d214ff48bec48
ze06d24220ec9daa2ad63d18aafa2602c158ef62be969ec69c0b54b49b24dd69e25deff5a081759
zf1c83db94391749598fa2e252fab5504709d2135b4db633a12332e4a24ce4de77816ad9ea6183f
zef7527bff615600d10c0abc7babb0a35c638eed296a4cf18bd663a604befaaadf76ca1dfac35f8
z65ad20e7fc7e959a757f7c4f7994b971ddc605dd6aefd750f5aa3f09f72cf5f92e1877155fcdf2
zb992517a306be482e62a1629d82e6b8ec98c1d5906244f43375ab254fd8ff178bed277b2a3c9ef
zff01ad0756b4cc410358ef2e4088f4cc88b4d4a51fd62a2cc4c12c0830dd87d2864b8e8d4868ec
ze53ff7483c2828b8935b1c15424453c1d051abef3c9b344d51f6e457e9a4ab46b2e40362d426fb
z09360911bcb46540b6ac6ff2097634d66c61341eed928fbb2936571e038eff9dd5b622c1b4fe1f
z6c2062a7f3bef7e8e9070fce57b8ccea31089315bb13b3fb7fb59dbbc77f552b7076326d405b5e
zab651b2901050f854eb1f5d4200a3ca304a9e357ebaaea8a1ef36894f84c1f545ac661e9feba4c
zf2a43fd32d322e07052d32774d2f16c019613f7b95d39d7643d1bcfd2a4a108788adf89cef557f
zffa616e7d6f9318397b87be8155944db1cd506ea6977c14c487e52f0309ac54a930bb77d551cae
zf85a5c58e1a48f2e0234388deb54acc7f66a1f34953f272ff4bf6b875b78a2a75ace7a3be63e07
zad0b99962d8bd3b3dd40b32eb32ffbc0859b19e61bef83fc3b14b26047dd522c60ce70470c255b
z07e85e8acc9666bc48ba7683c4d3f3136e1b0b7e682bc23e26b1180b849a8978fcbb9e52aa7915
z24d17190df7baffd144bf23280c2d0b49c137f838ca78f2925e48b657113658bedc70bf0a66e34
z91f98417d7e900e5fb2968269d84d7ae5db786523b7d0a3f02e2c85c8fe2058a6b8380408206c5
z21e23ee69fbb6183f29ae4d5cd01b2d96bfe99df6612e340c1a20e7c7a368d83a421e4de6054d5
z232bbc1e638512d1a2d82945dae2f3a0dc0e140ac0924f4cddf370294e61ddd4b22a8cc16c3acf
z38c4a339b90764730eaf343a467ef1ab50e028f016446d20ce7c2907c0ee109b80838950257767
z2024418267dd50f6db4d17abcc6bb453771274eb3a60ed6e6a1ea009426f0d710a196723d2cf13
z0d720d0a111a52aa08d391ce486c9ee8f0912904c3ad3bc50bd24eb8dc51cf0e3a5cf95281a350
z3c0b329e7bcba2ebe60e0603c01f8f1dc0e677a391daff0a9e5a5a6e377fdcef52d7e8b4c1f496
zad9790a2b1aa267b97950e9bf4ca15150adcb1062f435defa26dd96cb71474d9199ec8771a62dc
z15ae838c05cc03a8a254ead8174eb6ad7ac8763ad68582adc6070875386dcf4b9e209c9c023a86
zf30018d75242436d1540bb3ad3c04b6e19a8355f8d312fa41fc591a6716f4d105df3467bd8f9f4
zb118d40975da15239c459af20e9f87481b0fb2e6840778927755e78eac460dc0998c2186a2e9ac
z0d25b2ef1757998baad7cfc370c15263396528b48d4d4ad05230bc9e93745c7239f969f06fe7e3
z49a18d74894baea469413e864e04e5bf290c0d88966f45e11e74658b0abdf3bc5b584ace518236
z35b2729834386533d8fd4245aa1986643b51beda72ccd39d03bb1e485e544efb3526a3433d0a01
ze002cabcd0c7683b50fadc069c26b1b180df7c24b7628200a0b703eccf57c8465f950b0b6b92e4
zc028d8d3511092dddc27ea695e753ac41cc830e58afc3e75fff7cc1bb45cec5fc8f2614ed6dda7
zd5a4a8ef42669c63be0c4f82e1a5c83edb964aaee99594a18d2cf32e6976cc450201340a8daf23
z95372bf448ac388306f68ff2ef78afb40431ae7dc6d2fd0dfc71f858d85d9f5bf9340aeb824eb5
zbebe5ed36d4fdc51a591a1ae22d330441ba87c7d960027169a5619583f2c5780d35aae75243863
zcc18c6e0c275b97022c9cfd5dd21edc4a3a7b0ba824aff152a618975335fcda1539495365b1cfb
za9f4ac1231c5d2ab2de003183343e4d959ba84f4347dcfb535b7900b96105795a7b2ad42063258
z93e6e8d2523bf87ff3821d6526dd876068e8b593c2c470c018e52dd7eb0ac82dbb719ce3de9a86
zdf69cf2cd3f8ab793f28685cca310ce92eeadd3897abd66c07ac3f23ab47a96becf34793fca0c1
zd283189db0cd361ce979f95ade9bc1cc0ccbf6e7c7adbcb6a172d4747f98c9e1c0a008fa1a400c
z0a04c26d80bebd6bfd11ec2258a6fb5453decf44a07b666c44d963b719cece429554585594ab6e
z2665cd1a9dbd0ca9765416e8032375266f0f6815c46f536487e5cbfa09facad6542df395dd9fe9
z99b5ce6e8b0a4b8d323da9a03a67eaa34afd6b0a16508a089a266bd7da81be34bb2859ee5f3c63
zf18b5db4afbb3c43f55e593107f9534e341d30ef18c8b16085fc6d8fa7999ad2a970b75adad9bd
z5b29263f63154f3b5d1c3ca3140507e7ce4218dfe522262c463772ab5056e5c25858b76eb6c5b5
zb54ba11d66549e305be05ae602dde8e20a011f496f3b8ca7bc8a544af5d71f2af07b5fceda5baa
zed66f7c77af51d507bd11f89d67d6f094aeecbeaf20872d3a1c3dbfa9d664d8396337bf7c31302
zca8921c0ce08ab815a27b7e0f54fe6180fe7fa65dbde044523957d8c66e19b631b90cbf5848d1c
z51187a8464ff590f187c91be7d6c3e896c76f116d383b89eb607a6279b077402eb574be025db62
za7142a987e2bb1ee68d2d4648b4e8b4312c66029ed64bce712ef775752effedef7a182a1c9e850
z4ed002236fbecb4a845ff5212e4c387259d7e8658b04b813d86ea4c8eb3e2efb36c6bcbcacbbc0
zf25f98850ea7ff9d80cca95d4c22cbf4995fb3a69a5ca36349ed3dd1fed9ab5432f786d81b6e02
z861312ff6cf347f33864c8eb92e3fee488b04d9ee158a7635d10fb91f6720f4a24a29d8ebedd90
z9ebf971360762d991589e510014b01675bc0c09341741ea1ad75fc518bb4b78a774371e4f6d595
zc6d8c5a9ee7e8f9839877ae31d818ceea0184a3d6fe8a14ca642843b496aab20830fe301acda82
z048b232f338b6ce3cc5a8006ae5c7a8c759f18ec5cd13d5721c8aae672863827cccea8eafcf816
z83ffafd9bc79adfd9505e2b754a45cffdce15c11c16a13b9d228f00c824ec4df1cbd1791136d99
zabcfddc35d1bfc575467e55ecafd746ef831d09e027f059d9d068e1bae2a9827cd1ced5a9016b0
z6a8d9a030742101409d71b6a774b863065ed39e00306788e5d12dacbd03b8aa1957a53acbeb4b4
zad742898cc00fd0755a316922398c614cce54944fcf0a86dbf9fd1154c965a47bba97294adeba1
z294a07ac82b433b068bdd16f30657e4fcbad1ae66e364919c10cf88fd85ba8a94cc602aa7af47d
z4f0b8135524cce236e3d4698e1df8db98c5ccdd9e102e04dc6b16af48c3ab2933deb89da22c6b5
z1fc93faaa98edc1652a47f2eef91480ef3dcea124fb28acf607af9419af0ee2d2e9381cd2ee264
z23a7c51577d8f7c8511c7e3758569b6dd5220e7766631468e44def0275ba479a986a9ca2843836
zeb73809dc877a3366009c1ea7e1188c8dd46d95a3ddc0901c3ed635a64ad899bcc18587edcad06
z4b363fb75ffa92b08ce861f68eb12e8cd740814b615ef93b37f5abfabbebf9fa662442794a618c
z48046a38577e0aaf7c31b3986b4c928a6a7007e3643ccb56f6c852eb9fb661925fd4981af872e6
zfc4d9f5f408fb61283ee68258827d66fd62081f4354975543c327d61aec9de1a4d265ea0617bec
z0712456803b0191a8af8f64a800bcc96eac09c91df4f14a6a512f780319c218292052201c2f90e
z260f59dd5a935df7b06d45e8f81df3b028a91b212c85194b4a567b90e4883599345af09a19e8e9
z21816027befc5d8182fcacba28c1950614edab8bfc9d1ac69a5f5c594df581bd04cb5c199fe1ca
z6eca6aa0982e45f71a56f87dd8baa9b1f8a209cbb87320739f88199ed43c5bde92cf565b7e669d
za678f3ea2ddceae881678b3822e4288a1a0cdd1f9a822dbe900958a006b3c3a2c03e4b53f85a44
z275675c8cb6d2f547d93d75adafbcb160bbb0bfb90c1c7c757ba9c45760f84f71589c3996ee0ab
z3a3d3732ae5aebf467c289d62f1411233c65735d0f023b6e5d18109d43aa4603b652c14461c24c
z909cbc58ddd3b293858e7510b2d9c6e45d5aa00476287906279e6e826379d10846a5f1b8abe0d9
zcb9ab16282f2da5ce09ab439e5e4456ece9c0dc218d0f1237747605f0330602ff33df7c6ef1875
z7ae837d97310cbfaa694e0c0808113af889086d7ea568d49fa6fb21073193d8f61fc865ed73c39
z519472aa82263157f49632445e14250f023d090f69cd3af60085ef5f267ee7f39093c6271448ca
z5ac715510d22e3de8256cc4052243719670c83a99442567d33f7383b87ade3051bfbb535666b33
zde4bcc169e8bf1088354affa08c387b77951c2e56342696ec5f9dda60b555c95be30b7d5315f03
zcf291ffe47d993c0679813ff8ef9834f0db0d8a442755bac4728bf890848a6e5076cb199ee2646
zc789267981c51151898763192ad695ae712f19da7085e9554ed862749ae74709f7fa856bee5067
z1e13b18d0305b5487c8bb32940387c07ab80eeb9f750fccc002b36e3c17fabfd42220041d9b581
z67719513fa9628c7ffb04b0e6dfe696b26626e309fffef583765c23c87f4bd99e5801840f62be8
zbdf9f477b75bffbe6b045d913599e4e64c613aa3ffc55049fc56e805fc1b7283ab0c226a6225ba
zac931e6904e9e31c1f1df388308baea35640a2fcdec14b343b2dc0b9d28052bf3842b39654fc75
z1976f366893866470f83090a44007075f9bfe561df34680e8d23ef9514ab9a12682da4d7beba59
z66cdba3590d46376ee7d6c66a23c9cc38449e03584683a5cdbd18f6ba5c979f25ca015e681bb1b
zac2f7c5aa7f805d6a119211f0ed8b0118a23b4179a08d85b9b54d415dee58b5536b0af9ea3089a
z2b987b903367ac1d01cbaff6ac7558eba4777aa84fdc4afed5d77d90fc2a88fb07e5a430a47e4d
z78690243a8ce2b26ddcf560776d398645890bf1cb55b6e74b142d4aea95782285ee64263a70863
z868dc704f813fa454dbba529dff1eb0146e5e8c918e66298700d47f33abfe08a96cc2a92c9b9bf
zd6739d939d834adba66c2bbcb5d042eb1c5d90a04aa97d410b7a4ea71f2b690aa765b702592fbb
zb6b1245c421d94f05cd9cb0b29253a74eaaff76b9048769bae529c6b608b67422a59aef20d5a49
z4ab413bbbe8173b6f78140d21d9f4473e0e29bed3ac5f01b90f3dc4b1b79b9e5cf5117890b0a50
z406d01d864439b17f7853f62df5d214ba750090391d07de87ca833256d774820f0137be460ce96
z41cf68836e6732d53fa5c4dd77739f9c9017f0ed9475ce63fe0161df38b00b029e96526ace4b9b
z90012e73361c4adf60f0689a4bde8d256859c9d10671f5e6c0e58d33937e6b197c2d449dd53dec
zc7631884fdae7848fc9fc8759023aca3c8e9cac0d7476caf8e5d573c2b6396f84d2debcb20e030
z8b57be6eb1603182a011d95d6266e8bede875103d4be4fc7b0b479062b6b7c5017eeb3dc201b87
ze98e9d7f12b5d2c214ce04d39fd6a07b3acfe4334b530cd747cb0a3cf0fe83445ccc0c4c49cf22
z39d81d856d12461aa79a5e02a493364d07fe49df958968feee5e522e5d70d132f3df6fc38ae9d4
z57686b6b5674789f7577dddaf9f428ca1c1c278eef7a06bd6a61bc661c8cbe19bb220261d04791
z98097333f1e39e6a38481cd662d57a8798c5fe8d238e28bf941e97f880de8d7399412a3abafff0
ze2e57eb5d16a97da6dac2b1f05dd815cb733931531f61d4ba2107aefe7fd66cf81b738ece6b7ab
z1116217065c885c4085598163c1009b601f2f36a402928b3f6c15d6edb5c5cdfc67323e254a50c
zd95cebc8cf7a583fdd2959d9f19a7142666857153aee52d58e187ca0c9c2cf477a1eba86dad321
z1aee62e0afd4b74603f1ceb6e4b8bfc946a98aea40ed270cb54b2ddeb8f5e909261e1213a832bb
zfb1e83b93b308dd8d3afe91d2cf8ef8a8c3a7556961f85248dbccb2b21a0ee195b90ea11da965e
za168ad28ca898d85c187a7b27440bab5b5ad2b1da05f17c45b03ad769116c09fdfbbfd1c7dec21
z65df5c784acec2b645248648e9150cf6aaf66b0300f80010c1b01101ec7bb247b47e8726f03d43
z7cc0722aaf3718d82fa44ae4e379ddc280fc8ebf7bc7d658eba5f4d6c32359f2f685205c9a3c08
z6280fad1a570b4e43ce39fc1aaea888b77bdb3edae5442833742b53c93a489497d4f598a4a682c
zb1a8432dbb2156b909d2bb02c95e3b36f27229ebb9076bd9a8226df6b094dfe263b3b1477a5cca
z22556ce135d15db6b8d7e9691a0aba0b61d39b3a600e5ebda48421c7164c287e0462d11f5811f4
zbc78babaa2c7b0853e3ec129830a252a6f71c0d87bb06aa831f1ae077b2bcb32248017028e45aa
zbb93f9bb3bb0f32b77cc8d372944e8338ba47c522a9ad8dd07cf941541001ad53a79e2b323b12f
zcc29603e665d70b66937cae80b49196bf2366ca498ee62a72b2ba4449ad90d621c271606300a2d
z1591e8b9f965522b36c2f7833854a1bcd52d141d268b6a84b699ec37ea5a7a076059b81cce5f5f
z9f83be80cb4c5ec897718d4117fea968e01aaadcdf05564687c158267b2af105b0ce7e370e3d2f
za19bd042131f9e67a02bcbaf43f5ebc3ca24557f5b8fca3f6fbd8a85f84b90463d4c6d857e705e
z0c46443981c25b7f7f404405b0dc5d52ec129c06c3c0d3aedaba227f75a37f04584c111e343018
zbdd8af0d2c93190fa0bd053940e5123d98080e56afe3714e3466712ba7d88b1e0e7c26e399eeef
zc71861137da963ff71aa2a98a5cb9c6daed200848c377fd99ed66bbce902248907a6e3dc8707fb
z7c6be6b3dd53ea5aec2f585bde5f7fc7011126f5a7d7cace7c72c4cd3f62160991844ca06d16e5
z22dfbef85c00233f99c0bc4c85b8a9f93f36505c07253c6642bc8a2ebfc8bc1bdf5a654b93ee6c
z8a37485cf42ee6c47eb1db255e450fa518e053aefa643bed51fd1adfc61c41bb522b2f3a47c623
z5ec95695ce15f0fee6ae30d0f7d3e8396b4effc39d76eda0c66cfa7b9a5cbe8c3737b895764b04
z6a155b20f2585f9296938847019531ab845f4567af6f1e705a56761af771fb5a299d16a38c0200
z1e6498e685e133ed464b8c1aab859887f86e674d6433e9d55e7efe1cdd643ca7d826ea9af814e9
z09b1ca7b2fec0a0723c6ea755ed5fd0edc294f03c973dc156b57d4f314cab9d808689af2f42112
zb1df5f406d567ad18c93e22f97d6f3e973f55be5bde97ceea7425985e80b4b2db9fa494f396d8a
zf31f84f66a8db0a8a34452aa60924d346589d8016715854c32abf3633706c2013e9c450bf20e7b
z1ecd448a84db3c294dca469310c3f2047322d1e94747929d7cf09c5dc608c81b8d3630d36428c0
zde2c369ccacbf628d7c408dc0a7078f380db853e063769be0fa95b7e94ca251f20358f89c53b90
zc435bf74eb43a7939930211c47ae79b4168f5422ba91d16eb5bff98240076600717079aae9d0b7
z4b90fab543e6de74be13a959bf2f94ebfbaf6ada4c7abe9534a5690b37c0686947b1a32ba5d993
z5e90015754ce3dfb2f2a7d89bcdfb39ac90f93eeb70219e74d87c28986863bc4ee985fd6b69c34
zff6d7626b11521df2fdbb937559f226e190173178cfee6062d46a409cff565c787d9e1a0d07d5d
z269559c1acc7f517801f74f0e36785c5d630ad2dfd34f6f6453e80543beeb022d19918646febee
za470e8a1ce6c6eef92cdc8a57330924ee518a75fc403496397af2f1966938d3d44ab24b1aac777
z25a69ca444fc685e2ed2f86b156f5787e7a958ccb5a0339a813dbe14a0fe6f1aec06be268c7f58
z16412e24374570248e19bf430c413968d44924c91a33942f661af65b2011158a9424910846216f
z280dfd123bf3302280e89e8437e228662f0d2aa8895588ed9a1dd11a97b65b7ca401f2c5b7b35f
zf06f303c744d6ce4364a517f837d717a3fb87eef493e7cf5ad00901f9910cde52fc49117c03486
zcb5c03c2b19592443c48213783d2a0733e252357658560943e2ec25d2c65b9a61568e60067823f
z6afc54788c65a9045c6b58785f04ef8fcbc8a34864e91cb38e6d8d42cbdcbd5d9c54fb93879a33
z3312586f314a015886e3f833ce07983c222eade3d6177878327ecc130daf79d2d217e01456b422
za9cb4586bd8a8e7ed15363d5ad7e11ebee18654a879a2c6f6e060d2d015372dc5b93522c76388f
z0ad287a9a43d7c8246b28844c00a8da5bfded0d402247c2792d9e76c5665411403d136f39d4080
z8f4e74c654d917a4641fa75b5c67f135d71b803f77f833f65fe3f2d51f7454f005ab2a3c18136a
z9b78f4d735d1d298d2b62c27c35803ca035f981547be0454e3bae7730a1cbf933d163bc4169024
za8828b2633b00dd49281501e0b9dd129a2b6b24f7ab019c7fb5a5b785f5ca12980ebf391158202
z77c80e0c665a6c092291daaed4f4aee30eb76bb5e69ff2c8d2a6a7ba00bc9121ff138591fcd8e0
zdbb18d7f9e7bba8d4c648f66d8f3bfc1bb3fa90e664c79a976d808b3d536613386b489cd00766a
z10acd4daeedb7eb04c672dddc1b268f524b42c3b476ac45334a29b84cba49933c302f0ac3ebe24
zf1e790a4aea1b115b297aea5c1f5638e87c93d8f42335650fd271bbc75a59d217fe1964c122389
z555fbb3ba0505f1881c6b03898fd6fe843968e971cd586ea33fb72bdf41231faa501e130a33ad9
ze94a52e9a2b7eb54f109bb0df7b52074af63ff15966622c1199fbc298ddb6514a92345a7a4ff01
z11bfc5eb2956d34ec2385e88e711e9dc98f5479f02fb61d0a81dd4b6fe51b34ba820c7f43f1241
zba1d0ff887ce5e792bb2a48d866f30e615f84123e0a6a8f9f93327db25163dffb9ccf12e103e2e
z9744f843614443baf37f585886fe61ff72bfa777b8fe3305ce0a36637e079362ebdc8ac94f204d
z6ec03ea294646f573e045a4d4674c80ffd123f94e3c79cff49b37338f83781490211b47eea2e17
z2854363c6b5bc35f7f89f960fee4705ac1842779a7e9031a6527bc29f635b8d557574ae888319d
z312020828201874c88290f8d18a530ef9d7ec359bfbe3fca32d93e8ab63b97ffebc25b5676c9f3
z31b0454ab1cf4f98e647648d5d3a2de398be684596aef0a0a2136a47b6953b73dc7de84098e42c
z69773c46e73dca3a774e7e58e66472c0b8e51a6727e8d34c6ee6da7b7f8b26876cc1851f7dd426
z8b613c3ee4e7904b43ebf8f2221eb7499fc87f0e5270e99f0eac30f65b530cd0a6dc9adc90d8c5
z92cd97aa7c9aa4e4065447061c0da1c4bf9650fb1623c0c045cb8c0ec52033dcb3d27fdbd62e98
zd542ade4fd7189026546c1850d96a22f1959260cf77e031718162f4da85ad5cd9c1733fcd2abaa
z47faee3b7a87908378f3bf4ca3643ca08443c3c609ac9c49e70a30a3cebe888cb7c796790751af
z37e6b6296c815476147d02995ea4fc7fb27bd920df5d591b115ad4a0dd67e02a8cb20c7117c3d4
z938195baa52529c2c13c701100f7de2a8576a7548a5218abb9f038a43c6692fcee765fde3e52b6
z9876121f5802236adb2d740ee9c460ce9e992daf6fd2a9b384ee106802d744b5aa377dd3e3bd5c
z33f69232bfc58aa32994f1ff0c8d1fd129b485c4ff53b301562f6754e17bc128012b1179a29412
z915d1a75e6aac0aac2fdc754cc0761b1470cf52d886a27f975029d4ab4ad81f551d1d137ab0cba
z0041f2e6c9763d7944e61d5ba0e58846d3a1ddeb0374876e4c97cee032308ca42d9baea1ee3add
zb19506c49ec808e94b8876e6a96a4cd2af45e145a5b8a91f188469ff36dcba03b336416625ac70
z0b5d8c6609477af67d5924b0afdd7587e351365edd964a23995b8a063173918470ec11f6a30b15
z3f6e686eb6a06b302e657f56b4b095db5c0a26da0cb7d37234fa072920b4a80e2fdc379a343ddc
z3146371f7f3a67e54307fa7fae1218ac7239825a8b4a48a030fb76acc1addbca2186a37c9ea24f
z5542ec12d5d0fc8aacd12ab9eda4ac10e6c53a464c28aaf7a806941d45216441ae5843d4ddb52a
zfac95628be58a09c35d2855a82800153d755bde08fee2ccbe0721d86b6b3143a6b82c7bf10cb22
z290fd2cf282baf55a8ada12fbd0e775f3b39dbec952cda43223ecf65522c91a83d3cf677b1376f
z852b4257dd66a3f84c9c15ddea58e290d70bf9dac3c089c2e08366bb2b9685279015a47b4e9424
z467d821eb64c4f4da7c30304596a532eef5fc261ba1667562565f22c34d85b887693d17c4f2ee8
z668d3a895e65d7afe721468bf2072b28ff3b799d1cf86d1ab5e2a63f68568b4ca4e4909e83e6b5
zc82be7402097f9e134bdcdb44a092eecf81ce719b8f30040e4b9431a6ea4ad1f521dfcc4c1e06c
z3094315d458c45ac0463c1f60e0d5255ff72d4765294070c70ed8cc3d4584cca51019e33c4b397
z3541821643d64cf3d97c93396e688684f044d6d3acac14439238c7975104d81984912a7c39f9db
z93fc77013aa92a1abab0361b5ceaa016b6890af8455ba09284a8faba0abe6456f0bc407c3b5887
zdc694b52ad9fba138dde70ff76709058710029a623dd3acc22fbe38256824ca90bb2f095bb7c83
z6e9293f9be4a34c85f190436616919e468f43300efce76f6ed6fa0c38c7dba5a696c5507f210f3
z52c11a16a46e172346b4e454d9cda6c2fdcc338fd630f75ac24087d32bce31f7761bbc13aff916
z7078fce8dca2675e862696fe2571098a917b25305fdd759c049be4b1cc20dc6b05ec84cf86294b
zf7bf894c60d79b40e6d404e048fc8af091e843d02b49182db9f751f826ab3c1458077e4ec953a1
zfa64e4d1d8fc990add15c1f9e6f16d48d7201f69033350d0bae76e6b655e5112b6b769f308ebb3
z64e49ba9fa15a6f6b82afda8691ebde5dac1ed191e00377b7dab0cf19b64533332ad97b4d0b912
zb255c5c3351cdbd77a986613d6d6aae97d96da82d23a889f971e6b1bf479f2eccecaa7197cea20
zee349068189b854aee64947042634897f6263180f1f7c9bd3dff6b94a2b0335acbb2547b3c8afe
z38186c6e52ab02766f330abe70b12037de9f10ef5b3a33fcb0b4bf4a3c0273554b852da28e0d48
zbd887145199a2f45c5a52d527880a328740c8007e2c8e1250c326dc23f661dca5f1035871ac43b
z1b74cb655ebdf81eea9721b2795decec0c9ad811baabd400e16925bd6b06b7d36f8f3fa0430ba6
z8a5a8f89a7a7bb38616473b65c392411f007f08e3cc16638792e45f2b22af918cfce8ad71840cf
z6eea70aebf33103c29d86261bafe67b0ec6da951d1cd353c7d25bbbcdc534bafcf096a44116a63
z04e32a0e57060b22a8993c13b6653576d97849a3c4cdf3b910058205ba9afb6175127f1fd44008
z79804da0477d1abbba379f61b1ad1e3afe569e3c5df0c98d05b5ff1d8aeb1b0b7730232d362efa
z69be65afa62df7d152ecbcb48b2b8538a90f83c015f79872da4d691db325177287322de4982fc6
z2f3e445a717f17e5ce10b8383d9722623bf0dd4d5c1bfcaea519af4f74e601b5fd4de144abb94e
zd9b214860412c77518ae3aded08596a516e65760af09a2a678b3806fc3f4299f3360e6ee2694b6
z9695abbf4e6cefb8601a9036f7510213f49d2d0daeec537bf766f930a77651148a36b578919fde
zfdd02586c1efd14fa11ea555c6cb4ac24847ce09ed278eb580d06e04be33b57ef10a03fbfc01dd
z018bdc7131bf1b123803b0b7b13233b1c432c06be8512c7f75e7d8d240ea1fb7a0648cae888108
z64084a1f124039459fa769f59f6c5faecad78ebae1198da11b30bc08765706f3cba873c5d6c562
z2989d386e718ef5338d583e9898611ee64607f93550e79793aedf4abf5998cc71edc9422459be5
z02adc78557fa7c1845441226559ccf6d9c0ae41e84eba51fbda1ef5f88443cfcfe3c0a752b9d35
zd1fdba0e0b8d8521186658e6bf95b97dc358e3ab330db2596d13af3f727e3c06509c4ef8c8e80a
zd4d115ca5a66078860323a76c3bef271ea53fc95cc048af3bb5be8f0fc7c3b6d39ca389650d208
zd75af70d4f08bec149a69adadf4a5988aa0f823cd43ad50593b37a6513cbbbf3535471d494580f
z01e714c1a55dc1e79d77087a6573fcaacb144d093bc6ef5fc82fff4258cf4e573afecbd3f9bcff
z1396fed1f0311a0828ea0b235106aaa478894a5a257c696abf53a4cc5629bc704b0fd4cd42fa97
z747db81bf36e3456a690195f80fda0344a86cd0c5962ae6f302bff62feae095a6a7a697be2bf92
zd6349c2c77117c45bc698a60b4b0f1bf390ee93d94157e459e22efc3ba114c46ce0238caa79ade
ze48ae57f2d2e4321759283c0d775060829e6b238ff24a991f4220109698bc574fab77713d3f36d
zc9d9e0ddc7ba3506bab245cfd78a57c5e85ea183c8d0838803c684c1e39974db2fe06b796bf773
z79cc60e2e3b52112cfafb0d90ab3f16513afbdd8cfa7b250953bbea19bc5c8a99a668d8b65a13f
zfb04922fcd300380c4cf6694962c51bb618c0fb7ebb0df2b71f6f3b1bcb438f12429c76c08da1d
zaf442b34e3b98f6af764abf009309a6d83b0f5cb13757a0050045929b6c333a1a87d09b3be6798
z5821cfcf51c0582589cdaa588a2227de653f0dd8a80f7d659471eb8a7e50dc9a23fcd9bd9b2432
z6a4ab857efb34d45e262d61b35d9c3307f366bb0c9fb4bbb4a9df0b592ae88097902dcd3ed9fa0
za831a6178e0487fe03b7589799ad374439c012187b93e1423a3b1de7f1c2e3e74231a1f9a7f3b3
zd93118e67f56b228c35c1628883c
`end_protected_0in
`else
`ifdef MODEL_TECH
`include "qvl_value_coverage_assertions.mti.svp"
`endif // MODEL_TECH
`endif // encrypted_0in
