`ifdef encrypted_0in
`protected_0in
ze74c34e226135848fe16db9ffd31815111b6d7fb642c521a3f628cf6da949865580b22efd062a7
ze90adae0e65e66a2c36a587d0a790699161455169ed55a01f2084f11770a774ec4c588039b380f
z6de9c5084882a40b79a175f5c2114b2b6d78b070cb806e1c0aa9258297f4687ab308bc470f0040
zb0b1de382961eeeaf2e279e1462520fc31c119af8f2b214846f56c2b3cd2eadbe4099496abff18
z15cec83ec4a77b868344aa20ba7360908f5c0de2a79abf8b3534b883bb12180f68b5d4beb444cf
z3fba8f13afb0abfe8fcc4294810f75afe452434d2d0f1166236c82f76edf1e12979f04bc35693e
z32ae028996dd85737a8f5adc1ebb94f39c940246e887647b64782cd7ab429b0544c173176cede7
z01dfb26b1f73408344a52b7e1f117f12bb9c8077b34876c2e6fdc085981637012dc9754765e1a9
zc512ce062e0b8fb16a214591f5c81e1353b900a611fe1f4886b57940b41b7f2ce99a7b84b04b90
z916f717e73bd10589c81e207ed77ec660a8cbed5b487fa50acde1b055c8870bd8676023f21ddcf
z9c98cc47cfa2d654ff1365d1f45035a045a66c5dfa827905026270f0d55cdcaeacff2a9a621a2e
zad9d2af0fed53751e72de9a2364fe801bf0b44da25a3b2f4f57d013517bfaf4c7605f9b0ab9231
z0b9979d09bcb015ac8013f244488a1dfb590fe968c58bdeb22af8120f5a9d0291d4ad035086848
z6c022ce211cf658a88681cba3311865be47d9efdecae6661e8bf3bc5576623c6d01fa96f50668a
zae09f7f558532ce2c2021afae137c85146e2f306b4ceb08af0c708ee556d3dbf8425d5505d27ca
z4ef16bbe413b61333567858139c345ec6b136fa073b088f7b8579d5a741f15e0848a22f728ecad
z14e192bc11078c0aa71349121bf5425fd35eb6c6cba925cac4a7e409a57ea39cbd5def6a5d3d1a
zc01cf854ed8451b946722092a157dc7ca3d4f345bdc3cb18aac72b5256a257ff22a935526e5c89
z561ad23dc1ef0574bea112e186e5dc961848ad1564376ebff5de88812bc0a3e2c055498a2b3065
z23f2f18c058bbf0ff6aa19642d76a305810f541dbe6beaca18b6eb43a87a741e66c3cfb5567fd8
z31b759f7541b879604303dc4ff485deb7ceedcf81887a8ed5eccbc33817fe451b9b4ba684b9d95
z77ce3b5377ea30c158c4eb296b7b235260f77fefab4d1c0884bcc8b4d7c7895c616cdfa5f14141
zae96606c256f00e8b7f89fb4d39d6de1d893261359fc60bb8a68b6ceb531ee682fcc3fe1522ed8
zebb28b50e04a4034b01b937a929c3263bd753e6c2a1c8e04edb11dd00c6154c4d64a054f2db2b0
za856c16dc9953172247b4b66cdb7b26a3f1d53930ad3e64898347ddfdaa7a94f668742345f7d09
z7cba6f80ea80f36ae4024aae574756fe0eccafc330fa1b6abc9bdeeb4066b2eec6bbbcbf35015e
z2e8f5234e9048e2c0533c3c5cd91405b9e03140460d1d6c025dd04bed2175c6153846c333cb493
z07a31ad763dd977a227dc9c10bd4453234226864c286b40b8b5ba047f4c0bdb8ee2360038d9b7b
z237c4e2fea1217ec758ae0b7e699ba0a9d3f614680bdf7f7a4ea0f6b9fb55bfa3c9a13a1ecd6cb
za030859fa393a5503c251fcca10daa89b52149a0e9d3d780a9b6e6d1889018daa7d97d64780521
zc0d7561bfe56481cc7b7d7f3c7357ce748f67da20aefb9cedd42e694f101d68bae97d64da92c72
zc32ca4cc8b6b043b648d1eedaa519586107334d7ab432770a8660deb30ba0917b1845a8b4fdeb0
z05a1f21c69b9227398b2edbf0595956e32c59e1fe64369d30f88805a84c706ef57c72bf4ba15a8
zbcf1624e104ddabce99495e03de940b6a8a2394857b4a955ef4854b4d4d09cfaae4c2666f75875
z4e71af7c0edb595ff478608280302c4baf9f8703db91391b18e2ad0fbe3cddcaacc6826e5c889b
z2a830b05f101255ca285cbea62233b3717697477a251e1cdefa256003126e9950a6f3f1973681b
zd72d4c949c37e9d0ff239939a2a53b89c004d33478bc38103a71ad0808062ef09d3715e0a396cd
z8160e8475bd12023ab83ce2fb2a323e41ac33474cca3d27de5772144a39efc1089030ed3f4234b
z88e2b755a485cd2dba5719ba58b74a2a1dbc49181da0a0bf914e0a2d3c987092f3869d0b2217aa
zbf67a69438c9f73a51095ee660eaed14e98c10b8bab3ba6e1cf1c12918028fa3ce9f4ab048884b
z9355265e84580942dcc5f82144eacc6f4adc758bbd1ab9f9cdaaedccdce7b179938489910ecb01
z048cc0e9a1e4c89852591514d289094df5b7d72df65fc0412eccb91dfe6e9a4a0802035c0b5226
ze4430939f7e1e68055af909c47d61f940ad536aefe4ed5997330e1410d412c951265a3dcaa8006
z2bd409a7ce71f4fa6c7edda13da8b3414f415297c2673483006b5dcefb885a5da1f603991ec503
z1064bc539859b37f61edcfa02174a4bbdb77fc42e5a050b8de1d9c198c3bc56d8548b00f6be6ea
z984204dd78dc1c9d6658152dbfda11aa3766a77dfc37b08174ae73d41b5aeb9cdf631e7d58c2a9
zcb484e12c87b8764ec4550d9249559fc7f98f85a6fc82b652122bf98cc8f2bb3d4eed0e7212689
z6a1a86247fd9e0678576c0ca22c903f9b2b81f3a9da7866b48f61c4cc5b97fe1f2aadda0485c57
z7e93a1f599fdd9c35a527db2d43e319e48462946d92365ce80cc47f6b8e5845c70c11c1cebc531
z62e6dd06e1eb2804432c609e62be35fec8d1688636f9c64faccf85709c17fbe12098dfed0ef4ff
z40473d7c8c81a6a9c64e25285a9145b2784f6f4e7425b9bf0a4071b4074c60a16e7fe0ef391708
za8099446700debc529cc3749acdf0502b01ae57232d33b54f6d74a819f45138e7a09ab84c415b5
zc7d5fa631dd4645ac5eb11e4015e7194a3b4c2d6eecfd141697ee5e3a3c0c81a915413624f4717
z62ac2df6974855bb46d130443fac5ccc40c91ecc4738307e049a135de3d1a031b9dcf3eea246c4
z71419f827e0bda3be7148421e68ec0735d4e2f23f2123e398014d8c0a13a0b63e9b57e87d4e50c
z46fe36056c227833422d3e7fb6b7a7c2f21d5f1a343bffbd75debaad6a460b5eb0e90b6dab3484
z1905903b0a8e33550a0afffac0ab6cbe963d5945bf779c025128a48d3028a288d193be6ebb3310
z9bebbf2a006c360f6ec79fc2dfadca2048dc4135c36e91b04ab17215f6f0f21097937c3dd9e746
z92031436788d1d501293762d4af4ca25d2f64355ca593d39cf9c3270f31e5b769e4eb962c49031
zfb1e9e038bf5d7a502ce8b4332aad84064268d1e9b415d18c1f43a9947c5344b90f14467dd2538
zcb3eca4e8d0fefb07b99e6e366613755eaf33166d1ddad93d7037a6165fc9d8d9419e5f3adb7f6
z3abcb3765d2a94f99bf214d3dfc02c01cbea8b7242ebd823e810ce6fc7d58f8b4625aaf22c479a
z0c4c7d39b7a121ca7f81250aee510974ccbf4adde53bdca360ad4d47de56590fce66b25acce106
z27de8b2f175a3f0595fb0b4d6a7f2ba445ef390ede820d10c28e89c5f1cd55290226aac5602456
z82a8ac6b1ba4ed7f182f4ed9bbf0e1652b42f727738a9d84b7781b09203fdcb513ac9b915d8ffb
zbd2deff1e2827fce497288694b7f05fa346dac2b39ff6fd11ee02d2cf5ed312035bfee55bdcca2
za5e1f9aa68ec3d88d45e95dda338a6729d399ac464d7c81df38f6705eb58c9ee5f5f2ed751b48b
zaa78395d6c60a148b2dcead3c1ac4b38aff8dbe8f04f9bb47f4ced1bdf7fb8fa440b7a1beda06e
z2dbaf7144e899c23a09053e2eed2047606cc42d436ebf700978a4ce35d857fca5560c708f45a07
z2205b2806cbb0d9e7246f8f6b7fd5aa5083cfc480d1fd87b4804055ebadf5b0c4a7788bb9367e7
z29cb61d579269a4e0813c095d79271cf6d530934d4cb415a9f7a0edf551ca1752572f1d392287e
zf1489e61f761045ebd08cfdd9b5786042fb81b7866ccdec245626eb600ce8aa6db8d8a1f253aac
z46a79b5c023452adaee5ee520fa92dedfa03beae3e2b55d9c88143e6f2080570c477e58b0fd0ca
z3f7cdf5df862ef32beedba0f85cc043c743e26011f7e98274a794dccae49ae91c3879bbc3bad1f
ze062d77d5672f3df1bb1604938a8be6e3a5e84582db1d4e7a371eaf9f6b119c4eb7966d66ec6a6
z0b90078b1c74c4429cf922061f9e451701230389a4403e43164a24a33489da85e2584834f0b795
z3459f87eb6666672f187b95935913808629427e43cc630631ed444f06097ae900a5dba1e4448ea
z97fa629d8ef985afb618e21f11b123e9e77ce6eaf1e9bb5dee3675944a06e68cd8bb40baa674ed
z8a02de4e31a82aa3dba98f84ba88cc2687e3a07a19453dbf3f98f892a18eec5449a1d6371a6ff8
z16c7bbba9fccc3a66586f50465d139e2bc0b66b513a4162e172a5fa69d367a26188c8fc7994a33
zb2657f4bccae33a3cb2f61e227831fe3f69f56a266b337ad55a5c485a80ef4a7c3ab2f06a55245
z8cea69dfba8723dc0a703aafff04ca04cee561ec9b13b5770416ecaf9c77e3a6eb5da3292bcf99
za3a275ebb52b52da5df9f2560690cfdee96ac1a3802687b1aaf28a7c58bc1c4fd570dd53cfd9d1
zf31787d7b93581a50da0c14c3f79317021ce4c0fab9df8c8c2bb7355c58f2774e8931b001d3415
z4e0a6c8c071f53ea6a7865d9600254db20c31c3be9cc429c65ff0158eb477b42a461133a38befb
zdeba4ae59c9e79e28e661c485e40829876d5bb2b30d2076a8f6c94d2feb6138f4830cd864bce51
z081fddc4caf0f95c34cb5d3528002d2340d07d111533beebad4b6a36dc1d1d64120254c3df4311
zd5332be672a337aba09e8151d0d169e38710ed9d9fde58c0fb658b74d68068a894693e1cc9809f
zb7dedc29a3c911c3c908071596ee132785c17f298f771b08a870ea4834f146a79607aef6ff2357
zd50001d83b00f3bbaf46a40347c4203716fb41e0d67f50085d18438f4e10a73d48a8c4d1cbd308
z78254861c76b6da40c94d8640824df950fb11f156e6cffc8ec70d8d543f6fe91f441930094a9bf
zadea9ab0b7656b7ecaaf29a14ffe33aee78844277e316a584c8a9746d0fd27d223cf6632033308
zf675d2fcd2b909e8b2d1b87c1e0ee938211018dadb46ad2887cfb448224b6f8fd35b2f640cba4b
z6c357c125c686730d4a1af49e0c997e3fc5a49d205498d237e85e213897431947b9fc18adb3e6f
z00883e5b4695231baaaabdf3ec397c6086194a77733fd39fa1e3155bcfb1674e786b6812ba6385
z89d2838bed5a8aaee9de4487c9ecbe9222349c716d6edb23444e406fe1966a217dcd93c1851056
z628cea7a3c5b4351c58a674dae225e19bddfbd1bd875f1d46cca197b49640ce55634346ca3a9d8
z0c15986d1581451b17bc1ce53c95064a7f031090b3735d86cb2c3fddde6f94f1fc6c2c39d68cd2
z94dc7101acee30ca37c0f35e13cba608d49c832223870973339985c81c7efc0533288118fdbf61
z11a1837e760520815b0755652b9391b1dc59c9b55423653fc1ba76db586f5fa56e2101211a4b31
zce9b88caf1bc514748f21bc2f93c5fb899e57ca5e2f291afe2d3565a3bdf6d03c96b87f25d728c
z34404de076144e16f08030b4ef49e60f85a1081814f4599ff61073e513da0189076de6a93e9216
zabfbf169ba6faf73d4356c2c7352e780572c271b09317df2c7f8d6ea7ecb83f118db121699974b
zd570d8772f0935007fcf297e45f295fee91a299c9fe5cf705aa2a3642f24095d7a8c82e792b5cb
za9495cddf582daffd447820f3c665430faf7f7a0b430f533354aa851fd39758418801913f7d9ff
z3fb1ca4b8a3b5f6c220537f57d655e79019f5d7dbf403571d3a207c6a2d5db41d282783ccc5069
z0656b287a1c82cc4fd287ae2d275310947f2dad6e7330264bcc9d290c941134b8c9053d4936c17
z0691b9f65324d9e9e68f09b8cdc870776e5355bd42e04853012036e533d81e0d030c2c24995b94
zef5291dbe4d67ba5ce58da830dd5527c01236acb84148ca17fd442fbfeb93469c4b0ff5842ca9a
z3b86189cd5813f38c9b673f333223b22a6f5fe7d1663e11a7ab87379bdaeb3e0a89e76e93e1abe
z6352145abf9dfe76a3707bc18d559222af785fe93acd88112fe7835ebc456f8feb0a19a5531f72
zcafe1f09061200fbb7d4e087c7b7dcbbd9b61f0dd55c2e9eba44f83ba1f8558edc0c91d90e5c6a
z99c84f1d7f0828277aba30584a732ede2ddc8bd5f0d916b703852dfbe49e125005f0bb04957f1e
zc23f52c68e3a45f54acc37e36d069f17abc83fa639bff79eaf2490e9ed06f3b9593bcb5b98e104
z8dd2015e91b0c3f32510d3749c2e90f47d5cbda6936249a26a2ed8db22a366016eadd7cd21d8a8
zd9fe8e5b421ba8edd593dd987eaa7bf058e10ebee38991fc23f93afecff876220312292bbf7f8a
z5a85bfbb9461e2d8bf1b9ff7fb77f980952f8ad0c4e59ff621efc84c2cc88232d1eb0a336a5831
z0547beafda766b21aa655f6ccac02103baa921fd18257a0a62a266e4b3223e91dc89f37790019a
zbffec611c5c002fbbf35a39fb31e99a33db84abd246dd03ecfa808047794832d0ddf7d78bf50c4
zea7e6c13673ad50718a8989aa0cd406877f3200df96e5894e3d98ed44eb53c8bbf28f8c872aaf7
zb6bee10bfde534bd32e96bb22cf6270b56846a2b29fac66fef4623d5e03d74bf8e1d2960f9df3f
z25d471c9bc650e741d3c3471acc48e3c7a812991afaa29f0e12e876723e22a2952c7d702a4ea94
z530358dfafb4a8787cbb14003963b33c0098fa133213a9ddc44cf48f1bfbcc62c336f504e8eece
za55e2d927d396ffa0fd359fd47c3973e5814b30cc6498e179d35ac4d74c0d7e53cdb0150a53a65
za26fff25b8bc72140ab0215b785097f7269b6c5b3fc3d9ce2cbe0ff3840d67267e373b20e60e46
zcca105fa7593318ba119c19cddeadb45f4e55de2c7f55faef30265e465c82d5c15962fce345a3b
z11a9bb0dd034ab2df048a6546c0a3b3c6763750630afdebc949c62e91742b7603251c4588c05d4
z6d353bd55065ad200d3dbf228f096cf793ec920215b11a967b6418995eb6c19e4741bb1b843ebf
zd4f76e056c79681f51a69a89c31a43e9fe0a1478591ea3de3108b86aa985b68ea8522297d4449e
za52bf1a4b8187d4436435940b57d37f1ef7df36212030afed921c86ed0e0d8b7317c9fec54e38a
zbe7a932165742eda5cbca619585b2d7d556f2dd29bec5b22b9131d4d215a79ecd1e9520b6adbe4
z2c182a340713206dd53270e901213fcb2d21fe1c84649c0c8b04d041980b0c4a986b8b4112a592
z02a687487e4f47915542ffb72e9ccd8d96bfc3f6d1784ad34164f3ae2ab247087d947698da5162
z1efae4128535c07b1115001a14d84863e1a0925dd80057e95338009289f2ee6c054ce53cda8a7f
zcf158f2ad4bfeb0b799105ca2cab4c28aeb29d76de672bf8844c62a8de030c235ae3e2d27dffd4
z00a971ea6a6fde7dd85c3e5cc6fe6f4d7d99a659c230397468e8a8bcdb62066201249fe2ca798f
zbf6e6e0d65a49956da60f896b41df63e08950e07947d40e2fcf91992bacfdd1d52ad7b324429e3
z0eb9448a709a683cf410934e9cbb4a7aa015856885a52e3cca14cff24bcfd4bae5e08536f39e60
z3aff203fa760779bdc5a6c746e3d088795e494db9889462a225a301eb5f2c70c87666e51d70adb
z76b9eab7d1e91603a1b326e3cdea8dbb451a6eca3e62411944603c3047a43645b305d7fda3f94a
z46af784aba2ca70feb504e7f98081a0eb07f117cab9f2d51d79d2d6638289799aebbd9042b98dd
z0ddb52da4d7a2c646a50d05a089a7c1a0540e3299b0e90d07de92a1a79a3efe6d9ef119c9c73b6
z0cd1a3c5425a8468f06bf786471946ca0f8f4ac4df1da5b766fd371058b89b1a3fa057b9cb02cf
zebc81dcbddeb27afd22fada557bbf73068f9de151c34a2d1a5ee5372727a9c232b34a7f101ba02
zbc69c0842e681ade337e45ed0a8c9c51864009f755e0b8f9ffd93f8ba9cca77af181dea71c02f1
z25e40ce812b79e01def1fc5474d205f0395f6dc3c9a51d06c2115c38d3f94d79c0550a03b73fed
z996401768cb04be0fb93212f7835ed7bf113071f34ac8697e06d95faca4bff2f78f03b86008645
z22bc85936860cd1343b46e0f2c90e7ce9f0496d16acb07c38fed29e3e9a222a55908c3310d34a0
zdaf4d3541e270e6467b48d3bb4eee45800c74776e77f5c076cc5d5fa34703e89138df3ff30e269
z6c17a0dbe6966df1fbd1b4deb06d8e70a8542bdde2f4709fc32529416c18ddb180c0cbf24026b8
zb182caaab8774a8718928ee09f7b3fd0ec9497de26c0b29d31e493901f3b2b28dc00cd9deb04c6
z71e7068d4f1239edc74a3b93d5517630cb393cf685f4fdf30984270379d01b684a1c8a4a110a70
zf2a8514ecb4a9e18a358d0f6319f0849fbbe668e2ad9fbef75e46c9d4581ea634711cfb99cd0f5
z47c38939ba2869e6e2d78a57bd86422f1c1770422e3b55d89de1de80a56bb69ab4e23da95112dd
zd7ae938830c05658e4670e4ae126a60b51e7d3c9d5aedabd3ab4c92651196b580e923ca2b0be2b
zfe944925012cc26e869ae706af25ec23e04637f8cbf8c1df45bad7cda2997e3a347c22d01db833
z09af4cfe569b6adb5e954dd328d0542a79d34bb2f318d63384adc7dff2249e376e009833fd7b28
z181ff60b7abee65429b50be4391a5619cd67cf87098935020352b39e7f0edff7a2831d45c37392
z4c3bd3fd75b2cdcbb6a2373d66561759d152ca570a7035f5374d97050d15192bcde8c8c7a86710
zc1bd53a182bdcf3b31f8a7d9a8f18510449582ff007b541c05c375e1d56eecfe3f72d1caa76266
z7265ff61e70c2d5c145acbd2b98c221f82f71c3cde47404af4e967c915b7b0ee8abba4a1b6a6dc
za3a1ed3b5cb81c03542732927a4d152cf5d22399e29db849ff12b4158086104536935690f53489
z4bafe5e93860bb07942d31417fb667db6f74f3c1acd157692d2c6071f4de18ca87042a460d86ee
z983c63a85bc054d77693fcbd3c70ee7dc1c773cde9dcddd46ff06b3e95367195799e7673d874a3
z8ebcc9869242b1240d95debf8e5405e28a99a9e099afd9c02ff5166574535f58b456eb9ad8d4ba
z0a59a09c8af1f1f701a018a7397fd4b7afd2cd95de4f207eb94c035be61f35e52ec0644883aee3
z734f9e33451cb67f988305ddd04881802318dd827ca8d8dec3b31bc9d3d03eea83ce2f6440917b
zac371b4e2e347e959473ae0c2f22eb88eca0fda3c36f29440464ea07bf27440da2885ed51241a1
z2cb9797b550f53ffce5b6ebf4b870d6834c5da7fd245ffdf83a95ed7663ddbdae1eb472bf140e4
zc4409c1db69289ffce4719ee122fe4388010cb9810b4458fc5dc519a3ef99ed89bd8616ba83221
z333192e97d7466b64000513716812c8704ecddff2c2c22c2ce97febd709d5968a7a48092becf09
z3798bce9a9fa8f70a627e89941a05149a2b7936bc7173504025795a087e4cc88779b1ec402c178
zf69bcd57cb77e404b9e7634ad027308318d121b0226c44903cd42345473e0ca37ecd8a462b40f0
za473a91f68b4cfb6675d1979325d791176b0ee4595aaf88487aad8b2e4c61697207b0a30ccba27
z677d0a1254d8571fb0dcaf0afca34ead1c7fbf78940342960c49e1858cbe3607e7170f3bcf5291
z2ed3b5a82285dcffe80425d9f89485965a213449335c4c1c73cd74cd0900e3a9d1548e6a4e420a
ze6e992344f216c06b04d40baa81a715402f080bfd5977e9eefb5346f10e665c85b529eb4a0e6a9
z1f4bc65f82ca4a8d24d54e4abb5c2175d1016d6ccba7eb5d4c9991c9826668bdb7c4d81a6990a4
z2cda9ff02cde9c6ae2c07c5fd689b15ec378f3aef6134aba0cac3e738eb0fc7b98d06d4ebb470f
z4270bb1e29c06e5b08298186c25cfb4baa7b1c7c7ddc63acf84954def683f552bbd8ffffabbb37
z683747053bd6844891a9a85c304609d1a94ac468d14c1aa10280171cb9b9b894295735c5759f05
z74b383d26d56dea298bfc717a2c8fb79c4a84da8c386e057acd9a5984f482e8a3d0303bcb5b396
z4cbda775540ea3d89ac77a7c04897875541a920d7d2aa5ff6c62448fa42acf3839ac29e137c297
zd0dca880c9926a6c8b76a4d4da86335685ddb435e7983aebc1fbbf8c166ffcd99ecc23d50d1234
z2dabd665945aa5d0062c36994d94f52ce444d2ca7080b3a96e311b64770f4f59f4dc230dd46dbf
z436947ead74eb1bc7f9d2c77323c5fd4ee5adff8c05816be537029b05fba2d43a2921f1ef14376
zf2709929ee34e77f7b66a01b3b0a30a5719823410577958a85907e7e134947c397b8ad8fd7a927
ze1f29cb89841a8997412bac8dce8f547ee20d453a06ab3d21b032289999b18b7912b455334eebb
z80dd8b020b1c94885c7c216f8a88f7059c57f0164e297f110e68540d14111ddd68cafbe1822a07
z58dc0b5a58b02802db5f37a28241cf8a695e668b5d1096c2402d3f94f39cc8ebf711fd44fbbd42
z1dbf71628a931721d41002ca72fb0ee997a8d15b410d54d1a0e50494acc8ccadf63230a5247d19
z0af7ccaa84e64bbbd51ed19fd8919dfc6b27e9af92b72a7828ed630cc86cdd52ce37da42da3d8b
zd6eb6996ab4afbbeadebfc7014bd93ca8493581149bc3b45ea1e1b0f7d599a6156b39b9f7ab279
z586acd628ccf96857c791fe8b54b354466bbf2008adfbabd3756d67aa7582ff7638c61258dbe1c
z86eef5643b57469824dc01439f24a64c9e2016c0593dafa21f299f13ec107ff1205fd21cad3977
zc908289944c690227113b3cfc20cd7a3476ea17f38352c528f3f6ef6191a53babcb85cd387bbe1
z7107866a69c2305b98cb524679e3fdb702760a4056fb6ad46f2bbf70ae7fbafb130810c8b3fd4b
z0adee8382b18aeeef9475a83033127f9342be0a4d98f5a51b99991e1d19bfb2955631e587768df
za136fdb2e005ed9e875a755011dde774f9de3161a9cd0272a8f6140aef8e44fdcd2aeac445c12f
z6675661f9efaa2941460489b7a34da24961eb861304610a417faa888d7ef6dfe0cf9664dbcafb7
z86201ca36863e46271fdcbd35b8d2b2d95f35b90e412ee904bc130a0c0ac3330dfb8794392304c
z556d134ffc87a8e7e0d72a78ac6ed2fdf47e86bae1e734ef07ee06a6db899d92c660634b51c101
z84c277ad0ee40d716c971f7ca198a5834e95ef3de5dfe035de9a16d0443924d18de16affefac1f
z399fe755eb7292a8d3578dbc5b9642c4bbe217e706d1e9099deb39387da2aabb02bde1c7b08bf0
zc3d1f9ad9cedaa6d1a197ab07f36b66789736d4a132d700eeb8511412145b8fd440910861dabce
z2a06c0d963697280f9906b79360cbe4ec991569837ecb16b65148c52fd56ee9cbe76cf09731daf
za50683475bcb1d0e4652d84592cf015e640b0fc4c30c99c86df002d587302b0173d0c635f8b1d1
z0845fdabdbc1321b9f24b7be30f2b665668692408636b74b0f418945cb41e7bc5f6fb1eb152d7b
zbe784ea9edb9376c363b2c506d3d093e7b430125eddbbaf0965ad59455ef0cc01482be13ea0439
z9035178fab01fd1b104efb57ebea9624c348cee9055cab938aa08d0a1169aa4bc189b365aa85d4
z18ac86c648887355f0154a69d1aa03e6399f7bcb4b63812d047dbfd8156a4de26a0f5573be18cb
z2166dc57ad64c13abc39310d6d7b9d569f407551fddac856c308002bee8ffc2ba6021e6ce7776b
z5be9e27a3eb26d4e5a71b671464fe7977a3cb742cae397e0c5cb7a644787a3c833101a5997b4be
z1c8414366438bb90d0481973b15f7ccb3741723fd125a67ac00d387e4ba2413688f04ed33783df
z10760e27ca753dcf9eabd10fba502c0aa1210eddff7c9b23040de6933d9c3940b5ab67b2207878
z369e6538ee024ce05fb947f5f9a6036367513cedd5dbbd7c963cb250c8638ca1caeac3122f05bd
z3a6b7178d93aab97ee9b266fa56842de661c3afed01e0cdb5d96551985e1cb2b28ffaf837a343a
z671f7bb8edf681ed83a2012ea2a7b525b7cabce0a483a76408ec3b382af1d5c9ee27a72d4b1c15
z00794697804c805a399f0434deef02bcc50c0b9f5f1935b2dd70382601ca8551d04362d7dfa1b8
zb8bb1b9543426a3cfdac8ae17ad5e57e98a3f3e7b567bf13898821567369880599d05624c67836
z6b25d173908a7c229b7d501dc1c42ccf33d556eb1b45f0223adf9762452850ec30619ad3c1dd47
z914b29e28a62d0b39735376f41a4a3f01b698cb07d9cf8c3a51b3f465bcb06c8f689c27e99736a
z9ec34f7a0ae52644e49c36729a05071d33068c006209f87420fe293366204535e87f36ad33f1dc
zdb5b1433c8a5e8fe80e5ffb01987d02d9d43bc2c650d8552636415c74f3740a50d80d34fa43c42
z169062bccaf962bc755f5c2875e9b4cb8ecd9435c1431bc1418f8c3e927fd9e62499e0070e8702
z85da277884221041dcae1b76ef97e514ec89261a923f699757e1e1a8d0f7f96ad8b1616e992904
z3b154ed432cb8bb8d393b550ed70fcc9643f0cc5852a3403b0a3137801b517e6cade13b0d6745d
z7dff10f167da8292415703ca4025651775005b8736030394920cc0b8a09b49d6547148ae0f6e23
z5fcb261463fa1af9d8961d4476eb8a49257b251b6ea7a2344be5f59ba6e628bdb4d1daa2069550
zf27d763fa4d2a11be7eff36fe33e132dcbb1bdf0fa84918a8ffe56ca0790aa8b4bac54e095de3c
z15ff563090003e04daa5a404f5ff3bbadc037777cf9ae49a44ddd2ff2c27dfb3b1169b221738b8
z1ef15cf66ac52a13f63cbf94139803133069782b792d7b9b9c93f5577e87b4577292f79fce5b62
z38eaf928fd214241d2f0aa3b3acfc283cb692fe2b5d857ddcc88e618abc4010fca563627b1e026
z6035e0eee20cf2be49875413217dc8e3dad8b604cd42904c13f3cb7449fe0127facfe891f7609d
z2b4318d98546a5242f0f809fc83d820edb7c3696b877da2dbbc46c5676e4673d83ede6fe671baa
zbe78a01cce2b1ba225d4737d1c999859bd3b9eed850a3781da87f151616cc2bf6c0ceb5b2f616b
zcd56787287acf6298fd0505d7c4cc12118b2a8f55cb004ecd2084e6663c8f636e4ed102fb5e6a0
z0b138baa34915c3e6d5550c73132434f0f8c8cb5cf95736e8a34b3f0043094248ce48ccf719d31
z2672c3e7d8a0ae34b7948b3c18cfbd7d6b6a9e3835ddf8925114222c0d6025687387687038add3
z99de316e9d68687994fa7b8dd5cfa83151f5836c0cf6d7624d37563688d1ff57d48fd8c1c648e1
zc03beb0202dc36adcbb60b7303c449aeb487588f4e382cc6084fa7bf05d5b65a9cd4d266bde698
zac2dbde12977d59dacf13bb998d62648e4671e5974967ecadadf8a574687f7818ab052c1189940
z85f3820cc72bc5a92adaa4b51ce55caede72ce7bccbf2bcbf38f2557f76905edd3cb15b34b640b
z417cbfe99fe087fc014e8196d495bbf174195c4e6ec3c47b7e5e455ac9fd9076a556e173d2984a
z1f45920ffd305a441c4464a8f76b7d87e53c04ac37a79ce16adaa45e203eefe434ebb3be1db07d
zf4422943c21007f08441a9b185d36b2180d95b8606f3fe4219ff48776052c2337ed50b1ebd3d7d
z934ba2ab644df3e1cf635e291285b6e3db62d6bf5d5927a4993f2b36896b77c1a6fbfdd38482cc
z0457a58c815fa4441b78181c1a067f8c56cae4300aea01c3542a4e8124bb30e44ee788f148f83c
z3e399d33377128b88fed318e2624a9d2eb01fa0095b08c107cd93f3f3a85c84db22f334d73d1fd
z210e0b0560848025833b831732cee5d733198af239272f0aa1eec2f6f778ddb3a440a158374d52
z1d0ef09321fda19eacc070d3f389746ed1e988787c092b2a29ce820222a83875f4a24756945087
z54bba893a2a4f71d98694656a838008a396c8da9e5fd3aff171e9e984db9c352042c6af78903a5
z0f384a01330a9a86165101f623a6f701009e4cb684012267033c1d2368cae1989fb34aeaac1484
ze5146fcc2139e76491253942819db8b03d8dcc878c588625b66b2e3a4e3990345db7e7b8d5f834
z06eb4b293f7bcc9655e081a470f81ecffbaf037245c081d4d3c3554e54586b0ad8ad2fbb410ac5
za48e65c32141df255abdd258101a3d1c4681d5eaeeb8b154758a8f3ef8650fa0155d657bd558e2
z3bf0c5722964cc4fde3c19b40933aec20699a94fd997a904e4bdf18e7d342e909e62d01a276e09
zef3dd0af3f765f1e2700156f2533009a3dbd819e809a474ca1230130bb6ccb3c67a19658a962a6
z860dad803ed59736820dd047df6e8f9edc6104ee18b1f860fd64764237bbf5345e4249426206e5
zf1da253cae18b6f296380c6f87bdbeb767dcf99d2da720b021d60bd6ffb30a23bebbfdb05110e3
z64b1378a74686abfaf20c1139e1accfa4c645aa26f62825f59d8bf9c193b4b161072f6a828f3c6
z9d56ede446bcbe1a3b9cac6a80a1defcf676092d5b6ee3911a58c23ea1b47779e23e76b0ce8dcd
z6ad762a7d160a8e83d09de7717c768f9fb9308eea5656f0aac17237ad30b63f673877e0a11a740
z60cfe76b007c1573f862f45b51e2029d249401b5eac2818985b25b98548b6f61606dec84347c32
z117f4fdc594aa67d45674ff2c0542ab0ade7641c921e5f5edd0228de01070637689e79e4c23eca
z5848d491c5244ae4a725d3ea39cfdeb66172587661194703052621b110bfec95b2827535ae7ec9
z6939b929db1b5feaf843ee8e31b591403935585a5ba01e961f0297779f62e016e95b7381361e92
z8f19bc79fe43d5397cab26b1a66687b0ef54d9375cdcbfde29c81e974bb3cf864ab613009ff6c4
z2b7d5105fa0348f1281a147280745db078780ceed9eebad9ef991d06aef64754bf6605111c098d
z096c29f862486eddb23db2445fcc5ec14655df631b5d38f395bded0401ba940db8ebd630614b24
ze5ae8b0a2f4933684e5cbae6294c1b933599e5a82dcbde5bac93dd574e24ed934d267332512246
zea9cfcbb4c487b2ec014e03630a7ab55657314e5d67ea82cfe75bf23cbcdd015a564c08fe20869
zbfecf17ee0e12fa3ce77fa2863f6237e99fd9507126d8207383bd9c03a4cf916a171cc6f3c60c0
zd237f8fbb2b9e4605ff730bc3a9750f50595a18dfa35a7ef2861ec7200a4301ef6adfcede7fec4
zde2fd9cc3266445e8775899d205af3ed7ae64d8b859c9a7ece7f4004c6cbd5a56c05274a19dc46
zdd7516a8a233e0a8d24c42a5a912da74a8641f5715751f75250510b97940d1f05ec43db41e470e
zb55886c906f1a98107e30f082cfd9a1cee7b55644a88f6f49764e884b949c8a357777b216b2d5f
z7f5a07d1309ab7559d503a48fa6ea7c463dd5895a2c74a282b8c19f6dec270bef3021428157477
zbef4f3da2519afc8eedbf0acd6b7d1094eb8d174c78fc8c7c2032715fcd8bf404b2e8a13e820ad
z69bbf53d5b45ea6167f4877ae8103debace70483099f4950ed9c8dbb1962833885c11adf97bb44
zb0af52c20143c1d1be21fd9f3c6b5afcf6615fdb2843f16a1338a2b322b7fb22a71cb8f9943d06
zdaee4cb3144dbb787a7459a458d52197eeefaeea585a22317637b305edc7a6747213e90eed7eea
ze612c8bf2388e367ff1357d0586b0403bee96ba9386da799273a252c51e764a53a1df9de7dd0ff
z14db10e3c8440f1a4298becead981ec3d61266650be4e9828335f3612caa43a34a6ec1de9cfcdd
z8ac088525727089f38c72143693ed69999bbd5d13cb9d6cd21a2cd999e926e84a7c5bff5ce09ce
z0c82bcc8289bf2a919b50901993bcde5cc42eeda347e65e88d1394474315fcee64d9e2e58ab034
z272498d7ab422f651def6b05318892d9801794373253241c58a5fa482dc2e9c1399693d4069839
zb05b71fb92f3f7ee601d2747f6757d2fb4410c7fa0bb02d415ef8a9f5afcaa8e3fb8ae9a17614f
zafb00e36f3855f474dee99d741bb4eb486bb8f37b2975c1e0a73170fa417aba5e225c119e3cde0
z53b3f762762377e3d553dac55f637d68fcf73a4b59ec89909f2f65b4d4de21b69a097800d1232d
zcd63004c8abb90b4f9d4d2cae4d71e0792a7a26fb53b04a7845e19b2929f00e54fdb90a2e815d4
z313bbaec4f4b7105a2a965115828ba6647f56ae812c51ae493b2b7fcd3cb13f26c33fc9584e1e4
z2f2c9840ed09e50c3d1e52e11e7a11191a73d3b569768388e9bc0a2fe4adba84360d5335cf4374
ze00430c36c6cf2f1ba3601a152b18da0c6136b3b2f2637f8ff64eab07802a450d63d5d62a2cf87
zb85af4771b60977bcff116215377a978ceca15a6b7a8c21293b1e38733657750421b6d6ce08396
zdb1a29cc16b4262baf30879b373fc2047ec8850c51469255aec6f56e2f91425e310b0138563384
zfa7819b88d4dd013bdfcba356363c8c9b085f7fae05f15886cfe37afb3837bc61bc987ac864b57
zf7590d2104a057d8692ce2d83713f4ca1e936d520b5b8475eb25595773a55385b1c0518b0329d5
z4fb722aa87f03d5594481839dbf447498b901a5cba82350245871b2f2a4bdb0f520bedce17b123
zdf85742fa33829076e0e4558c221768f4682c54ea662852f9b24b4ee7c59d8bd6fc57546e986e8
z8f71224a1c33c655ea617fa54713da8dc24e82940dc07b2a9d57b40fef7069da986622f02ea808
zedfc5e6d8b8d35e2c282cfb8c7b8d39bbd03630ca5393352009cb5f656812c45583778283420a4
z94b57ad4b6731faa8cb648f6edaf9b9f09c17277f47e38d25c85a06899cd4306b65ec848ab5a80
z0628b175d6092a9cbfd96e0954a83b85f5cc111a57d2b5b263e4811f357c98fbf40920648e0d5b
z15dedee8eecc72ac3a722a0d1d1f60b814d7a26a75b3338b63804e577fe4735a655c4e112b3b22
zb783ec0faabf631982550ed091a60da96d49619b954eebdbcd928fd0cc9326380789f1b0e37a44
z365d5b068ac01f57e6e57f5865808b14640950e133539656ea18fc5760b624c2d2ece486ba25f2
z0ebe4acc24a646133f7033601d4917e848bcd07a2a56aebd7669f7fc68ee8cbe79cdc2e9711ca5
z26911a46f30d7bc611cbc57c36b755863f9d07e8049089d7ea3431f9b34a0fd3f568a8fb3826c8
z69dea627c81b54ab93d7a9ab3fd5e7dab262313097819afa1962f81a1d95539be06faf46fbcea0
z5530ca800fb152e3ad27ab6cfd88c3a13b68755735f9a2fa07ee5a0ff76f27a2aaecb8472b5c3d
z8c8691abec4cf055267151fd9f515c4870f13d6ee9ccec15d50886e022aeebdf0a3cbe5a33ab94
zed1043b45c6110b368824e706abeb7f0f507d4cdd3f6a89c5cf892a0c4d72b75e4db3a85761126
zc70d9cc39cfc61a7cfd213b2e7c1f6a024ed2b9b3e7dd7a9b5b476920d371111493d3aa4637169
z81038dbbae66cde5eb91bc83935fc042cc4270ec10346de7ef4152c92467e4fcb70ceb7cfefb22
z742540faeefc39e0a0e9d70ffac716c36d54a59c2f9d1969e12a0c8d032e42d1d57a4d0568cd91
z59b6ecdaad330682982026229160202235872ff3bcc5251a894b020e3df15e90c56650ece538da
z98b336c718d383596e9026dc4995220131ae2b230101b742a4d6dde49797a54f3d99f9e00f1b10
z5934e5b08c9aea73baffedce950c62aeaee36f55ca8f8cf316b45b70c76f52e44e4576251eb5c9
z2296f84dbf09be79cf3387dc3dcb8ac5fbd624d1aea630d1828b40772ebfe10c7e1f8fb7604a98
z393929c236f574b7311d9ecd4783075d662c53edd4f6e3d2c8919a193652c4fa82d5723b034b98
z0defabc7d23c1018c2b952fe62975e8b3f9d44e1becd0ee2b5b95b9d2572a8543c292b7f7b3b98
z481da99e17ea58660b97a4030fa1a7ee56b87b93a908763352a019a732d3534f27b2c3da4ddb55
z9267b69ae5434fba956c81776dee4265400570cfc6d22e42a00c0833cbc618c0587c9be5438343
z90a45146a7db62fa5fd05e3f67752380aff61589012fe1d07bdb475de02bc815af9801464fe519
z334842dca8410dd0e48c35e5f3964f6ff9b6d51d01c795cb23e2f8e26d366b56503e3d9464b4af
zd81f76af145e5237b84de4fb7119115c8bf20523e158c7bd97880057c267dce5d901a1c1494a80
z87285d0445ca60623445d5c56f1aaa9abdc8abf33e087ed18ac6344691afd4fdc0d7ca218373ba
z52d081a2d13012c59fb862e5e5fe8ab4da2f2a5d77901b1e9dd21679f4419c936115965aaed4d6
z11e7b7b434e968d6565eb8b48856fbe3b3bf7d7263cd53c95c270ef8dd7710aea494daa9f11590
zd0e622938a9012f6c9a7833b0b6717dc3e5b05204f60a76603748cc1f33dd18850ffa0f4ec5c16
zca9e0ad0694c07275236fa60a1801d60adb84816bb3489b60324b5f8d0c032f5b444977d611527
z59a28c69e8959819574607de45a493f9c7e9e183e598a02a7ef8ca6e2be9d87c8c8c061e50ed13
z45e4fe46b6f24794d94e90b39482f70eea858c209d66cfc6e48dfb0303ddca54edacbaabc0ed3c
z438caa7ee26f7dbd9ce01b52fe0d31cdcbd583f3bbdb0da34f45f3f6debf606dc7437edda029c2
z194097bd3468733575815c689b7c995200a52d016314203178825e209fd9efb071b9ae3087d3c3
z38d6a24a2c37eb79c8c5050e6e321d614ce1afdd120cdabcabfef2bd3c3040fb87284faa617313
ze328bed8add0ee44cddad310ae3bd555f9c73ecb6f3f5dee8d23a75e0991c2854d2510558c1e9a
zcbf9f6bc99ba60835bc6aa3c724e37f1ab8e75e5bf20731f9bc12051da5f06b21406d2bff6cfa2
z786f9cb2b90dd607e39fd146749b204a98acec327b69d3d4471d3bdd5a2b11803fc64db50db5ac
z2540f7552d6d88c1ba4278501835152e231d78528823f75eaf0e04f86b0b7a04c080ec97268102
zeb3e990c6cd258c9dd5b7ef7d0ff71bedc6a1652980e77c70b61aa85c3afd491ada865583ee018
z9050ffee41f2f8d64778c0493d10f5e5444f2eb539f2f14dec0d76ea9eb8855bc2bb24f50435c3
z3561ae082f5adfeb068c2b2e6a3610bc1385cc1bc234aab191e4fa02ce5c58fdcaa504d51a1260
z1258bd6945702ed627b19e06d8ccfc6e9a9ff4a9795e86425d5de70563eeb1bcd8917344b889a7
z4ea1ad7720d73adb3b0c904c87028f58893172e195ca18fc48291cc7d682f196103637bb0709b6
z08a480e9c8cf804ee6a45c1cfa8a4033400ae359439132a7b1de51d9c46f39c76ec847f1d11ae9
z495dbc43d32f624ae0aa280f3c4c4b5697df3d175e097a40bd79a78ee11f50073c182ce6a59daf
zf20ef8af46d207d7c3f11c6e55e3ebdab539265ac432f0a84a14d5234e0b8d8551f8b9cbae4a27
zfbe9b580f39d4eff3929fa0f501e22c9b31f70dfd76458aa1a6afb5f4c6b2a9916cbccd2827fb2
z58ef32d3b63cc6c3ee27d37d6ed481983e4f1d1826bfdfac1e8256a1e17089d06887447eb4af19
z7bb5cb6a190431b76181caaa921c05b44271e800a8db2c6ebe50da76028a300e6e8459a4c791ed
z69f9984080996521006f05c5186d92361073133df310d206646614b8c4bad1fa49624f0ef29652
z32d62648258e617d822ef47302bfe4cf214888ce0a0b3e7c5736994f7bd4ae4daf3ad6300aae79
z75a0ad5a09feb934ac75e2445b8011da5b86a1708c7857814fd0a229c8d87aabcf5e030301b03d
zae600ff1272d29a0e87cafce306fed0e83652a380d9370a84930d4d03224774d54d2fb49c1e397
zc8acaaaa9d6d67212e90600beeec617ae12e59030bcc1fc729c12329f6229c8251ed90685f1ac8
zbef9693db5af22a4238dd65ce26eb6fbbc08459cb29eb8a337d2047a39ecfb6f90b36cc0a1fbfd
zb5dfc354a02862b7df8a303a0f2da996d3e47478646853ceb26b74cd44e93064cd65894923134c
zccbe6f833a867dda02b90d2aa165c4cefe7c6edd0a5444d46dd613976476cdebc80edbd953720e
z33a745d30dceacec3006ea4d5aadb406e400ca7a63c1f9d0c70b52dc4dfd615150c4d08d9551e6
zc8bf9d0985fc2d761d5c7b0e2addf8fffaff85531df736213c193c75bf1e4bc25b9a9c9569a571
z3c4afecfbfa352f287c9a7b1bf2a402ddcc15b40b577a9c2eac45459d200ab5f0a5e718137c627
z18f3f777bdcdf58638224a5453625244ce7005d6a4c6e453f6526e490336ee5f42d24a1eda0544
zded133f5ec28ffa4e2f3f041e0f505f8382a14adb0f2a135a299e9a5fb21a12d2ce49ba132c114
z8ebfd40b7fc2bc4d3a49b692362b98d208b0695943710608a2a6fc22a8a7bc5c25b0b8188f4181
zee640bcf9ed383523e9ffb361e8a4deff08741ee6b54e44d2e847ce5389b4394f975dc958959a8
z5f823873f2b489de885fb405aa7afa41e964787dda8833b11f795b20af77c4939f7799cc33825d
z66bc7a844c9db45eb687cf75f87dc5f61c1e24376012bc9504bdc7053d20c00bb95fd3df537fc1
z064f629b331b7eb5d89ea47a4d529d6a19a7f8d22883b70bb21b5e112216dcf3d2b8ea98729ee1
z4fc472a8361ce76caab3a96dedb6d97a09289db07d3c80b6259f30bcce2f648c1b7c55cd047660
z0f3caec6963684090dbec24b7a4ba8fa0d6448d89e597ec510a0c7dc77a0db507ba39db19b654a
z5889ae86e17ff7bbf7e3c82dbdffa1d04f660b10bfc3f2d623534cd91f4bbc9cbbf912c920ae9a
z4c470167e45619b035996fa534495dfea30ac3bb66db9bc1946fe55997dbba2c50c771316c3e79
z086721397263f84c5fff7dbdb9ee71485a6dcf95dd83b07cdac9e1dc2efad899a38c9a248ee189
z00895371dfb9f5cbdd013cbf5622d2ea254991d671cd321195979d02e3fb9b3d80901581d0f7bb
zb47fa9a9f16f9ed5413f2437d7672600287f53e99f2dcdb95bd14c0468e1410c8cdc599f128db7
z88af3de559acaa2dc8840e6a8cd3cfaf453210187c71009f8c8d2659b4de75a16fcd7e9fab1184
zfa68978c2b05f2e3b4e92173a67dfbdf7df1ac91eec83f032a80b544640e84130a099e874aa655
zac53b7cf99737f066d1099e3fe1d643048f85377646d629f11cedcbeab4c95037eca56fe84b103
z5beeb5a2a96ef40ce6ceda51ae3791f0fcb482dd5b7a0f7bb50c28921102a64a88468a54c2a5ec
z982afe74d2f55fe11d0d4deaacc2f5de94586a4c8f38ed28786358fde8be9236c9fbda2b3afa16
z8291c2859320e17f2bcea9dccac81ef0949c53dd6346cfeb5d6cafefa810f970a69b23c6d9a4b1
za34b07260ed7738cd1ff36c2bbb8d6a546b6194d39da45d7e83d70a98d280b2896ab589e957952
zafa45907992fec12f04bb98e0e87870dd5afaf1ef91153c334a96c83fae9212f0c2e1bdc74e79b
z9c4eeb9716db2804ef1972be170310e70cad2cfa0a93a2be372c501b3bb5e48503e23b69cca733
zd255af39486e1e6f848aca911b861bd2d5222e474891e47223979aa6da460274c01c9afd728131
zf933b952d69fac8b3d82172d4f2988d72333d058b6fe41290f0a44d769114d732850ef48b5c92d
z2160e6163465c10296a873aca93a20da71d0ec4decd9c05450bb5acba7e75185a25b749c1632d6
z02cf82b18ab85b9f9871474b15444616a5e7ba5816058bc0030c9e657dd8dca39e2cefd31afcbb
zf4d1ef28733d4294b5106f8760484ab1fac70556d90d4cb607d0f2cf2756cda8703ac9b01937b0
z02413bf50768c3ce076c1507cecd8a48cf023ab791af64863330e843b26311ab742b93b4b17003
zd81e5e4d8ab584aceecfcac1c6a41974dfe4ad44be05e1df56925668bff8514cf4255e648b02ad
za35c6ea09538e72e0c507e1d0e3405c55f26bb0cf3736d3affd638f4cbc1cca0ed37ac5a1e5724
zce285d13fd959fb107693fc4a3c24c5b7cfc44fd34ff137d0a7f6bbd46736454649493ec007c18
z225f13d00f4a42adf151ff49fe715a8eafe0a00bffcaecf95a28b2354c66561e78a0a1f1003261
ze3678b512151f4f542a85703c1261b992644fc70947c6a866b58b9993ef0b05e686a680bd74804
zddcd4d97ec8c2e14d75620fbd8a95034e3866f836d217ca3eed591acfa2c692a7abcde4e44556c
zec5aaeec92f091f271b2af21ec91007052475d44e6cfdb70086e16b1dd94a8596143b3e4e10adc
zfbcbbf8a89d29ffb3e13091f19816888644bdc9f37bf58646d2686cee5c55e6a216042c44c1aed
z8cd570c56f388ba8dcc73ddb040d2f97011be18e1b9bf787db49e93325444bac71228242af4ea0
z63112681a630fb3978c379d56228c0cc931ae0a15276f4d7da9574427dbd712c4ce04a7df801b3
z948dc3f00614db71b67a774fdc89f4bc50673566c2d0e421eea04707c53c39f06d672f640cfa7f
z8e6c38e14acd67b1d0da8c4680a957878b815f5747fe986f7bc8571999aea41edb58c576f8fcca
ze517f165322dc5349ffc92cb70cb109e3c98401920fe9e12993ff3f88df281f1b8b61143561a40
z86a6f8578a6583c06ee1ba0444be886b3f1bb9070e227fb59ba0eb579ba06f5b42d0691d164998
z5872c7958b6a0b525ee5f01426de65ef6cdbbb4ee5e38c91fe9166bd90267e7ca5fc555d8a9192
z1f9a98f24fcaab1e0a27d001ee3093a8f309d6e3ee978447efda75781c9071aa9b3b81f59ade95
zb3a27a2caa662419fb49636b9022bdda0960100e56e07ece36468caa2949047b20aab7d2eb4bbd
z56d9d94b5b7cf666f9b2d310f45c3aaf5ce47403644a1d82834d1bc6afa0d530b916bf29f292ba
z28de53b865ccdaa6693b1b6a28334762f67c2712a1de3ea421701af888a1ab7dd474c450dd2247
zf169d93985e3aa06a062d09c362dd32a6c8e64d46db6957e5f61d54de3ce99c56f1feded020f5b
z5abbe9018db8db0f11c5a2627e89455e638dd483087cba452927b8102bcac19976908173f4f3a0
z7d9d5939c3ed385882248ac11e6e816a468b40c816ac8984e7d21faddb90847a5db41362607fe4
z3f8ef299e3d7a7758d84ce4ad0520a5ff91ce515a42284d2f14641d0ce9b70cdb92559afcfa5a9
zf5607271bcceb8129df7e9419ac85203fafbe146949c6e000c7dde179a5aa23bfc2831f307e3b6
zd3e70b915bc2184f8b4adab868837cb74a6a28f33ee1f87ceccd98cf93267c2bdfa9ebcfd47232
zb26718004d50503a0c03e7799febdc1cbe8d398e83d37e1ed11dce6cc32c252ac2b32c2b1737a5
zad2216aa64244681a9d666ce36adc9b3d9b71beeac906129ab830ea8f08893b722ee86874be764
z8ae1443b0c93d4f652c97cdd242962770aa8099089df139ab92d996ee4853d9ca129f67b85bc74
z93f7de2e233ec579f669129f054ddeba99c546f7d1e326ccecebc459d06237ef053ab40a988785
z218b79996c9eacb21b480da2b79859858d564256f542c99454e18a7b0b6cb6e2331c5bac02e149
z4d716195819a1e3e2d8bf4e4a1c0fafb6b5ae0555e753597e17ebdd4bd22f9579953a3d29539e6
ze98731926ee4d16db0ce3fd5c078ae247dd7aca3e020246f460c1b99bd7ba869b52bf8dcd8a271
z5bff5ab1b086b6ddbdd0c80d3d62c3b9a200f5b9cc2f65aab4ac25268e3eda3f820cb5d46f88ca
z0658cfc5839045aefdc39af09d55495e40e2be4e9599ae3d72ff64da5c8c2712611703baafbeb1
z3c6e00b6ef4c73fdcc68ddada3ba43e8b559560b669cc6b88f96e7e465700e11aa82ffd7ff1fa4
z85b199cf36330a1795e90b38ea6dafe178bb845e59cc2462ba2fdb3849fa03fed76b07e066218f
z569392d497d9269378529933beb8ea4ab679bc5857c6d7ed91dd92d8509322bc65baae8318a09c
z4ef2c8d4b513721d5ef828c61d28dac88a6b85be29696f3ea2046a544ce1ee7edaa4528297ef9f
z2dd670e7c9846a407dd3119fa97c9262e8c2945706ff60feceac77a404c17dc9adce9ae30bfed8
z24565513642ce341a55e59a3dd00cd71b715cfcfb1610e972d553ae1c7e6f878f8ebc229b6b911
z77d1a7a53986743497869e39a3c381c0d4d5f623687df3931d725f20da74f2b50c1873fdaa9cdb
z3085e6680095e75e7b6ebcbec98e384f81ed6c324c517f574c98d6b076e790c30376a0de5a175a
zc9c6bd210f006d39d75f0e2fae51384e2abfdeccb257faf014605966723f9b605f7119505d9096
z82d8f3dad542e1993792768555fbdf50655aa2a19a99b9fb64743e49c6a735f2f375f3079d9db6
zb1d939cece61e141477f6ae25b4502fe327fb5b80236907585d5a939a51e3737696a63e5471fd8
zced99a445c2a23638dbe0d80b9837492ce44412be9
`end_protected_0in
`else
`ifdef MODEL_TECH
`include "qvl_bits_on_assertions.mti.svp"
`endif // MODEL_TECH
`endif // encrypted_0in
