`ifdef encrypted_0in
`protected_0in
ze74c34e226135848fe16db9ffd31815111b6d7fb642c521a3f628cf6da949865580b22efd062a7
ze90adae0e65e66a2c36a587d0a790699161455169ed55a01f2084f11770a774ec4c588039b380f
z6de9c5084882a40b79a175f5c2114b2b6d78b070cb806e1c0aa9258297f4687ab308bc470f0040
zb0b1de382961eeeaf2e279e1462520fc31c119af8f2b214846f56c2b3cd2eadbe4099496abff18
z15cec83ec4a77b868344aa20ba7360908f5c0de2a79abf8b3534b883bb12180f68b5d4beb444cf
z3fba8f13afb0abfe8fcc4294810f75afe452434d2d0f1166236c82f76edf1e12979f04bc35693e
z32ae028996dd85737a8f5adc1ebb94f39c940246e887647b64782cd7ab429b0544c173176cede7
z01dfb26b1f73408344a52b7e1f117f12bb9c8077b34876c2e6fdc085981637012dc9754765e1a9
zc512ce062e0b8fb16a214591f5c81e1353b900a611fe1f4886b57940b41b7f2ce99a7b84b04b90
z916f717e73bd10589c81e207ed77ec660a8cbed5b487fa50acde1b055c8870bd8676023f21ddcf
z9c98cc47cfa2d654ff1365d1f45035a045a66c5dfa82790502623b57a3af03bf0f0c0d35b51558
zb8b5f2d29acf03737a9ca2a053b7a8f06800d50b465c41b30eb585f62f3d0c2c5a43bc0dd4407e
z8b71c8dcc082c778e934db418ba934a51b6940c3128e6ca3bed99b5c448e33301cce43bbb16527
zb33aff8e41f054be58098e5324afa737ab3ab85c9e5a105cbc657982b652e62ae1ab29aab7d567
z61be0315875d31cc8d6b8d45bc02c93e7e8d3af266449e91343265d087f5ae05b2ff56c0d36be7
zf1afd86e789e18d86421fcaeca542198fd1cfc7200137c3b5fd73f72c9455538dc60672ee0f775
za18bcfdc993490c24876deeb25a52dd808c493c446e4c2c4b2442331524ef7ac93fd23014a2b27
z4548f52a14da4f9dacc4dd8db336a85e4f796d9ce3bf28d44d807b9401a78f01344f9e8e7e51c9
z914735ea9fa20a7d52dd5b463b5b2fe1c4737139ada619ecf451cfd7357f951bc1bd73d42e5c33
z142a1362f224b1f13a44290c540f894851b90de482f52cf5c30d0a765810b3e5cca1f13c2a2146
z5d706aeebc387fe826084a31a38855e17f8bc1f1e23721542d7006fd2225e57bd8a0d91c4d2588
z0fe2c1100cb41235036d7d3e9fc252f61e32c91ac5495de3fddcb0786f021f4ed6444babdd8cea
z254e7a30da9ec3a5714243e5679ac54314e9ffdb5ac54773456e73c85442d06d885846be6436e8
z83a09b88e2e7847123dc977d3060706fb15c432e2c5f2e5fe60538c22e5285b75928633749a5a7
zeb2a2220d57c5b15d0cd05ff0e26a69f3c43ccaca0708aafe75def249338638723329b0b67df63
z92390bc799e8a28b5f88edfdcb55a84ebefda154d443a8ada19c0679088706308f5be25cfa7551
z31c38da6458df208ad2a01f2f77e158df360ce5853e99def2a82c204fde9dd72a99a265308f54d
z386e28447da03c30ece259dbc8becb9a712f5a02768fbe58cdf7162f252d323c183b35e265da4a
z5e658c64951fbb64624e67f1d4677c4dfb6d5f5560ef47d99c8e12c4600c2fb596a65851c6f3b7
z747ed444e1dbd31630a9b5f3059d5d31116f8481b2e177c5747f6778731954eed28b9848b6b402
z3112f32265f2837710b9f810a91de95784e3a6ea3a6e4b198a616cdb80522e2a86249ffd34ebca
z2a19e00cfe292ca282736916871a564ba747cb9899cf4af21cbf0ed3d37bedc3fb12051e31e0c0
ze611239ed9d3b593f31bdfeb1164cbfd4cd3ba6a81d3b39555076ff21fa17a0acb8146849e1946
z48ae46f9d8c97864ffe99e12aba455c5134eb05ce3123b824be952866311090a1bfdade267b949
ze78eaf320333b64ff38382e06ba4260c286e19856783f566eff472a605b5d620e250b144ca9641
zde2049cc2769de03ca57d13f8c83bcf73ecf7337cd36b1a731b0fb5d3233c353e09727b24880b5
za5c32345691b8e2c02c14689f567c467d79bd72a0655255ca8a18e8c1756f0a196b9415e2d6f7b
z866e4ba1cfc9bc987e624278654aa3d06d49e88e54eac8013e2b10bcc8ee964127404790b0788a
zde0ecdd16a7e926fb51b1f9669087ff8d9bfc1777a9fe530baabc4d8cc4a82389cd340736c12a6
zc1bbf8df28875f26ddb7e530498805106f54a5249d59ecb98cf5afee142faacec2e3a70973b78b
z9a76e19949e7c7e0ebf38f5106246ec8ffba57435e228a6c793b3a90a9663d0e7be18eae1bfae2
z0a101776cdc2d5f3a555d51083bdc56ae6817f55199dca1f6212a8876784769d8b583214725e00
z6bd3bf93b8a3fb6caeae45c5e1ad54146e5569dee9abd9be6263241e17773c9e6ce27cc2f80e48
zb0909d5339c112ee1ac7550c2cca68c3e1b856a81094d788db9c269c07f4b66c17e6698849214a
za8704a6b1b1a6cc3aa01a42599cf4a4df83dadd0bf9d4c78821ee8cc9283f4ec3318b33e9ae9b0
z54f555577daddeccd27d3828b9c2cc6a51d2c4bd30c98848cf05097fbc98428db92f565daa27f2
za9829519ee4ba43083dec26874bc65ed23cd75a0030467440472329516687e69fe543f2a8b2374
zf369d8946e626ba9fe4489b3f57bb767d2770463fa031c168d76a7e855c39996cb111ea6f448fa
z55d6018dc1808082be33e5a88645f404bb23c521b4233bfa813125dad47e537f74ba574a8b665d
z9654c38e67975693771c29fc0992573f76f7e633993be1090924dbaa5495e781989d9dfc141223
z16d1f414efe7c8a54f38d998e1920d8692788749666b09e0c0f599d65e16f581b989d4f9442f26
z4329bdc7557cd9a79f0d6a9263e099bf298107be114c05546d085f26125e8132cf4ae884369bdd
zcf1a3a2ec05a97e816c2c8e7eca8894d8c2f9d89da569ba1f2dc5897a89bd261f664e634125596
z39d2e4e1fed08559aeb4396f988b3db867d4b129e4013d997efe9074aae10f8435ee462908601c
zd69a7e89939829111c9933e1cf341b1db58c0c6d8e90066ffe3493dc7044077a3ef09dab5c1ee4
ze026149ae8b170ac48999b5a2d7f4a55373de29698d7355047b063f3a78e9d4715d0a96e715e45
z73e3ac929217a44d650c4e1a9f05235d37bcd0333f2a35d42cdf930b97365c8ae922bb12f6a792
z94456d32be037007bf512ef2d95c015f77133af357bd949f7125d137d72b4023274461f278c540
z4e3db98d9e17e4ee10a7b448a0dab32097f6e9e202d13e5a305f5d1314deed3c2afc269ac1bd14
z3923b74003e8179e63f754bcc0c912d489838937d964a25272ae96797ae7848fb962d42f82e708
z3910a10ec305b3ba63e2246b665fab942d8d99e79dc7e1269c8a32dadf0042c0588c7a2001d98a
zf1ebc34bf52370fc980f43dd8d40f96aad63578f779cc4226b30fa7b073f41e7fb9e4e79c22652
zaaf6119cd12e0fae0f85fb24de9057844e9ae9891b70a51d6b336994c454843a0dbca9786b22da
z97826c1ed47137ac34874b5b3433cb86351f7719d3c65afe430b86391530df243f00c2df541464
z82c7ceaa81217be9a223225149bd661c5ea199ca9b982cfa3b507c1204b363eb96624a03622ccc
z1932d85637e43dcc2fff6e842341bc973b28dc674e75b430227a0c65d1205b5e92345041935157
z621e7ecd1ffc1e7fecf8fb2d5955af05e4717c47e3aca84511a368b99dce9fe5a029efb7cb2bd9
z87e0749ec91bb065cd006041da164d4f51a478846febf7ae52508495462674d5d37b299f158584
zb3d84d3d0b0d849a1fe62f9898fcba8b731ff61d5ad3fa52bc364b469525cb83b78fd319877de9
zb579d665cddcc716255754f636f052881d3cb141861a167cfee32883148ec4720aa595dda6cf78
z5ea1a8ec9e37a117dc0e01a26f92e9a8cee166acd4458935bd63a0dea5138af31658075f1b8fca
z84b712b54bd48bdd1462c38f222e924ff441ba987cab80a0c0de7b2b3805076c6e3fe9ea80e8b4
z4d7b3e43f8471fbfb60029c8ac18bd46fb9dd986b8351b0fbaf1939b8e8a8748253f3d6e5b10c4
zbe67757d242638ebf5cd7a8e2294578c137b5a9a018a465f9e01b9a711072bd4ea2d8426af2df9
z85a12976db30dc654fb9fb72239772d1e2ebea6b046fbf2ed97aba0d078149cd087038420f2d9e
z6ae9413e75eda5eb23c949c33b28504404764e042a9eca948eaf2518643e7a84c56920bc7c6688
ze1da7ef6bb6ed4e3f87feaa190f0125b9ad12e371abc58c4f75680360a1db8e97dab2c490d6fe9
zb0cc749c6d4e7d2b761987db964eefe0b8f19d46ab2cef4dd2a945c95a6be1a76762762b2e17e9
z97765036c3c3d35f447dadf2a87c83ba049d7cc897f99bb74b232a719e77ef9e8f4d7cc5135e8b
z3107583b8e321ac3d7ba647ffda0465e2290c83a1bc93673ed1d75075f1e1a619e7f436fa6a375
zbf6dc32e826b5c2d9ce45e673f33857f8490c7563e6e679433edc890ff1ba7da2a2be343e85708
zc64f631c25569d18d47a9b3a848913433e1195730561eb8875441a06e2b97749650ed27b32f786
z3c53c5adf0bbb50b265c48f56f73c8739d5fb9c1565ea11a48817f66f935f0aa93f79b2c131d9a
zdc3613c25efe9f3a58b6b624b0ba5a98da0ffdd1006b615b21ffde0e9bb760beeeef0928a1ca9e
z8f3e9ee8c484dafebd5fe9b202d57775e94fe45c3c90816c0dda057d91434aa69abb5d425b22b6
z3adbf3224adc88746688af5196b42b6dead3267127acc07ddd5b2c11fc6fc7d1cf1ec50df08c9c
z5e366b25ecbb16716093fe86e4294bed79752f2d1f50b4e06bb194d4f754bd584598d3ef304911
z8f16034df03d961393f5ce3dcfde675cf195cdf5c2aea45e9937cd75b2fe5c3ffe4a10dbd4c62a
z5581ed34132e27be99c8c9afedee6977abdf1ce6d2be0e883156c6fc65e56c6d70cc30f4357678
z32ed95c8b371b689e12a3f03e425264bd5297a247112f831a1d477adb61ea40e899f0640519deb
zd7df526a65ed9ff1eb2de0b5343b14c0ade2391f8a2deb16a333fd43ed380310a591b3e85658dc
z9320ae63239ff8d1b785cae238d519a577cb53dc984162d74833c77e429b7988c290ca3af32f64
z85704291f3e38dbb939cb2fd3e57e53c97a39dd807f010842e4f06572be689e6ff2730a63826e6
z9ae192fcc1f834cef009bacdca2b1b48b239fb2968e20bd5446f0aa37685667bed91473e449789
zcb58db42ccb3291105fd8957a727e63f157a977ef44b89e2ead0b866d3ec5bf546f82665057bf9
z3cf152d5e580efe9d115c2f0207dde9c11a126521a67997176f347273aadecc0cb4ed730167eab
zb87a3f1557f044f52a39761874062d39da32f1c1f6977588e9365cd8522e8f199b8e9c33b42295
z860bb2c368597b709688f86b299f8540a6bb0d45e99304b87b2c6784ed8cb4408bdf67878a0f8a
zc668a7e329894ce0ec4d00bd9b0e68ddff913f070e7f6e5cb5c8ed285e2b20df2494a641eaf521
zccd96e9d7e5f566d8c92f538878767634b8cea9f6880f1abd61a95a2ca80ccedb0cc02544edfa2
za32b4c616694a672cd20d79ad5784ef3e62ca879fa245a24776412a2bd4226841b5cb261c58fff
z5c2c4d3c610a2402563d37f59476f9186758ae4b30bbece16ee159246d8057d1361debe7690cb2
z995e286bebc47e8d17a3492a59cbaf3bdab3eb0314355e715a96f6e531a56b1e6d428d26f7045d
z39c642109839efb273e949bd2d8c1e1d62298c8a3ea6107bed13fc503e74098bd66860f02621a8
z642a7ff8dbae9b35e3f41636e7a8950aeab77fc6f26c5ebb4222c1a5a0479e4ec2ca951589c432
z563da2fb9fe8c864b6d3e5cfb6c32e7471ca42f3c04cdb8de3ea52a666ed197bfe81375eedf5ec
z026a2b263a772d8d4a305b40bec0ea007a585329e8d191acdb08dea37cc06ef23b0c78621dd828
z839d2b22f6754aad1eeb177c5de237a49b511a4b09dc54ad0d9abdb1a43fa8c6cd467694dee80a
z1618960878010923208e18b10f99234fa704844ca9e9faa8ea52da91a5b86ece9ecdfce40110d3
z2f326a601c2c126b24c6e02b529bd6f4069b74c57db3df346331c1d1d3a74f5531766dd723f5bd
z548da4ef119bd9895d8200e27b3a110bd3de0cfe9a69ed4eec478a8585d1dd14b7ddc52701cd70
z9b0537bd855bab73d0c900eb62d701927325ab8b90837b252edf3b8d4fcb34493acfc873e4742b
z28f89af190986ad18afe034bf8dd9be5cc6da148219b9e0394aff8942d210de4bde7ee054e6d36
zb7c996b787a22bd8585cd1c6ce3980eeb9b56ed6c75cebf08e64cd00aadaea29fdc0ba3309ee6b
z8874d136867e83dfc9d73631103a6a803c5bc2e4eecc55ae5f232c24bbb910b55ce6cab5e1c874
z936abf1e6e4de392df62bdf0dfcf6a495d4435f76bb32398911ea18c7a51378fe3547f2c5e23f0
z9553d16ac566633643e016c905abcd7ca4d6e5eefec276a0aea9d6a4ff22c0ebbe73a328c24257
zc34c20b7889228802ab3b6d4138c543ce36020ff64fda1d13c789a94f18f727aaddf7fdf3e0542
zda705eefe8787e3b72f7f4a6b6c1cdf319cabaa7a3e36b4669483157ab28175194b4e1f378150f
zbb7efb3f273e4d83534d17f991303fd0e3e103a385f3ad383644560841e9fc949c52389f1dd82c
z245652df05fa0d12f6a806afc359e39e88b73369b106783dea0414d62afa5ab1495f808f67ccc4
zf0f84a8b8c39795b9de78a594a79221d90b2cf7e4dc30ccd8888c9a2a3372afcdf4d6d9b79af0e
z27030302060b8d3980a220ab7d11ffa7bad92abc0148be8d17c2dd40855f35be17ce1afbe4e50d
z3fcae23ddbe72d3d34d1583652c762a01d2b395fba6abc1155b476971cd8885d64988f4a9550aa
z76195653a018ab5a05401371ef669d35154fe449d23520bfccbbfe2b7f6c1d1289da8dbb9452e2
z404f70e7f2d7f36cd49491aa5043920a0242c133af4385388ce16d62246941492643ccaaf6298e
z4ab22f68a532492a8d9d69eb19147c61e0f29c9046aab70a870aa1fcb2497e0b2cd5be29df3930
z7b51f7dc94824c7f5576e5ed6b8f8f1940bc1512aef4bfcd0b9510fdfd8928de981b71b6dd621b
zb10c69ef97961c84807ec39e9f910bb0eed0d24f54e99ff4d01888cfaa72afb0ff213a62eabb83
z71fb129c4e8875fa90e52f271f8436ce0ae4bb00da57e539a5765cad58059e546f03bc8c013d13
z13b2f1ad876f0f05ae91b843d7f12a455d3ccdd199f645c7160def2c85becb071f64aab07d1f18
z424c00356ca8cce4582902acd8ec5bb1867f9df785472e392e43062fdac08274d1d486cc9e129d
zc254d45416f7570820e72577f22cf27b496ec9b76a71313ffde60aa55913f3a21d2650ef91c44c
zf2bc6814249a34fee0466471a6ebe7a2048d0ccbdbf6f3ec33ec09d5839614de5953143359682d
z67c86cda1130fa918d8710157d2e5805a67afb652e827abc038eae29ce08050bf3a3f328aa0ed4
zd96b0928733b553d7b9f1fd6eb03ebbad4d7b6b3bd8dacfd200d949b7e6fe3741a6690c03fdfbb
z303b083f85bfafa39527b05e23ac64a30c10f784ae2927aeb462302002934d273be72cab855ea7
z5f1af9e7e6e9ba9cc72002081892a21c6b896d5edc3f2107e11ae9f3ecde044b7d1b1960c100a5
zd35092000122c83d46d02d8c5e2cc315fbf49cdb889c45d318945a70eded8b7604696d85fdfef5
z8e22ef91ff4ff0179b83248e1f5854f6630f2a37450bf4328f946991f146c7f962fd5c52da9d5d
z6189e2a2adf616ec444bf03cf7a665e4afd51da8bdd12ae6c0ef62bf2b417296a9cc0f48d0743b
z12ee370647e013275a86368581b1da0b37b53de32f7430b5ee9ebebd4d0a65aa8f169da64d0f85
z7d9dc56019af09c999ab595720381526c3780291c639d89222ca6f6eb1f4eba97771a6413b59a6
z70879958a0719cb36560cc84b3ae1bfee0a847a3092c9dc75cb54bb5a839af552f8777920241fd
z7af3329f883dcd7c9fe90c1c0e4b0b647aae46298d85914b3fd990a817c7a1990d9e4d1294fb4b
z130dc0532cf4661b91070f9ee0c7ddcea38dedd1cf454d539adff6de2cc93442e66d695443bd33
zafe456eba77c5b0d59535ce707d792b6d2e9b19b095ba1973dc0ac2a4cec346118329513705d08
z6b913e70c61a6a71f7aefc35d9f984898c4dfae8eb04aaa374007a21fd30a1ca258eef1c423085
zef26484c99113295494851403fd86ab9a05272541aad3eb491a955f05cefa91183e09223b6af99
z277b60559014deee74fc76637eb9ea68f0f8c3da9fd44e144ad4726005c59b161233294f3d67f6
zfb58aecf4098c2b24671e4850c6ae1195407b0ca089a97c6fc318e4602675618035d48c8f3bf9e
zd2c19663608098fc22347c604d503a4ad527625f590cf6c42bf97bce0e06140b3e7da8fe5628b1
zf7ddfed56f7f8f887bf3d6356f8cfea980094d2cb14e6d196a1a42dc1ebd895d7e1f57003ec5f8
z03e9bacd5bbb5b557dd75998bd16369344b4f92bbb486b4090e128af601de8c53605c7410bfeaa
z2edd2f75bc3cf94cc4c187713f3a4ad76982410a76ea432160742242280783a200f40588987fd7
z75ebe6d82f3254263700465703fbc3ad6fcd3d9950006d0636e36fb8119ca41e13664f6cfc7495
zea2c65912757e18bc3b1ea7726493c22a1e7a8430fe72fd6af899e8d235162e31e37ebea6e8be9
z895c73384f3e5d1ed0eac25e0c0daa1adfce764c69d96112ce5a4f0993e7ef71da24826348a331
zc4be9ce998af797aee19549417964b9d194fbeafee7167f9b9e1fc939bb0b51216c69a5cc1d3c7
z4e246187d547bbce251b94fe4a305863a71c558cd0abc5e0c2b7239cfaf6bcd983423a3e6e0793
zc27851d3bf9641803a420acfbcc09255927630152c80ddf357d975e31502dcb6f77727eb727190
z92a6c26c88fc66e6f12157ccc5fba6e6ae69450beb8979b8035b53cfe9187b0b9ace053c0ae3b3
z2e75e4b1f5cd97dfa6280f16a78ae281ad42f33b161733d320df06250da56a325a0c2f9fae4901
z448dd378c8a7c315ce8ca1eeb8420a7d71bb7f2a6af0e76ba51460428c4abd90fb8fb6f6a421b4
za7a9058e9f329479ca9fba3b186ed467a3a48d5648e97e3d72f54fb6fd8eeb2ee59acf341341f3
z0ae80f8a5531a39498af741b0b74687a118fb834af7bbcbab3cfd608bfb9bb44fe87fc456dcfab
z7b5feed726f45795253379b7d5909fcab0fb068534d035a82808fdc294154a5be8b3aa8e1e8f0b
zd4faae7f9dfd193d47ec4a8e25e01dbcbd3a61b16627c4648bbd19c2cef077c0859d8273c85933
z6548aadc2cbaf0701568c6dae9058f5fa3c2432038dc01c2463a25336d12d29de94f7029c06211
z569d0f0135c4fc54dcf043758247d597507fb88902ea07dcf5c7883f86dfb572184e6633c34e3e
zab32a49d858ceffce7896e8be11e77137c13dd238b328cf235cd0577ff3daf865ca591a1c3dc4d
zf371defcbb28a1e45b388a6ebed888d05889a4c471acc72bbc01840dcd8106c7ce7e6c06dbe5e1
z606693779153a843bcbf0cf4dc7c36a62cb8b583e88eae3789052e6d4be5020cdba7336ea2f34b
z6a5926657422a3105dddac3c4802822c45b2177dceba7521deedba3c1e59bd39ea592a7af4c60f
z47eb8ecaa43d2e10b4951f5e2db6
`end_protected_0in
`else
`ifdef MODEL_TECH
`include "qvl_coverage_assertions.mti.svp"
`endif // MODEL_TECH
`endif // encrypted_0in
