module tb_divider;
// TODO: Implement divider testbench
endmodule