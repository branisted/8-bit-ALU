`ifdef encrypted_0in
`protected_0in
ze74c34e226135848fe16db9ffd31815111b6d7fb642c521a3f628cf6da949865580b22efd062a7
ze90adae0e65e66a2c36a587d0a790699161455169ed55a01f2084f11770a774ec4c588039b380f
z6de9c5084882a40b79a175f5c2114b2b6d78b070cb806e1c0aa9258297f4687ab308bc470f0040
zb0b1de382961eeeaf2e279e1462520fc31c119af8f2b214846f56c2b3cd2eadbe4099496abff18
z15cec83ec4a77b868344aa20ba7360908f5c0de2a79abf8b3534b883bb12180f68b5d4beb444cf
z3fba8f13afb0abfe8fcc4294810f75afe452434d2d0f1166236c82f76edf1e12979f04bc35693e
z32ae028996dd85737a8f5adc1ebb94f39c940246e887647b64782cd7ab429b0544c173176cede7
z01dfb26b1f73408344a52b7e1f117f12bb9c8077b34876c2e6fdc085981637012dc9754765e1a9
zc512ce062e0b8fb16a214591f5c81e1353b900a611fe1f4886b57940b41b7f2ce99a7b84b04b90
z916f717e73bd10589c81e207ed77ec660a8cbed5b487fa50acde1b055c8870bd8676023f21ddcf
z9c98cc47cfa2d654ff1365d1f45035a045a66c5dfa82790502623b57a3af03bf0f0c0d35b51558
zb8b5f2d29acf03737a9ca2a053b7a8f06800d50b465c41b30eb585f62f3d0c2c5a43bc70d6577a
zc250106fe61d6067e7f6fd2d8c98bd222c93c90eafcd7364b8672ce12246ba12b85bce60d0ce82
z8fca6c8c1afe03b9a6190aadc08b4a295ed8596493a06ac8335d43af360db9101e1b8e9bc17434
z4ca519a2228068041ae415a981cd6214aad8ae2156c8f72f1cf4da47653bfe3d91bc19705088dd
z10869b6e3900abbfa1bf2d0b0fe2e68604d52b2b0bc79e7a1941b7ce45a42e4092434b6ec03ce3
z52230d9426f19dd2d6bae87349535abe873c8f30898cb8ef9a4278b209a2336adfb6876cc2d2ad
z91949406a968b8e3a82609ae69818f310a2c71b2ca992fc6b41ed1dc8bed5a30c85c4cdad74d02
z35dcb6fb21e1aae00d583ffe2cdb07eb79374890d6c81bf7945a65273c76724ee254d20efce509
z4eb1996120383171717a1fcc3501bee2d94259c68c6f242f023932a339d8799a0ffedc069fa88c
z2849e77046814316b4d96c95c83d7f58ebf299a7d51edbd3c77be6752021ceec9968be2376bc19
zdcd0518242456bf82dfd37835b151128189952788261dddf68b00c599ab4c3df50d1e07af20877
z91ab3753043f121fbe26c99c0d9fb88bf6f1faa44f0d742353aebc2201473a5f8e4ea493551d31
z061f8839dfa36f37be636ff790db5ebc9054ed7053404005e9575c71713735b0c445fec8bf1df3
zf5621d82ac1efcf0526f19a7220dfa6c03e501bd0a125bea848b992a12a4c0ac1e63b86f0a4ac7
zafc2512a17c5cb8ed211ada24a10bd540ff389331bced17a5e7574f8fe1cb7e0ea9adb5ccaf11f
zeb0ba8a09e370c71c0398e4471b0a9ef7194eb499593591708854003856a5bb69f37390ad64afd
z43e59e807410c27fac58c5061fca1d9fcc9418d60b458032565ae0ad72e14391fc711ae97cfeb7
z7f97f53610772141836288e9e2a9740e7be2695eee0722fb660bb6998b910739343db66ad08ddb
z2328beb8023e6159232d570f0103bde7d442c567ec58c903729868707171f76a11ef286967e578
z3a4c316ebfc6ed9ce057830dc566d42fdc73342a7c57afa84da414b0d0e16ab2682b91466b107c
zd00f53ae547bbeef9a8c2626c218ea69c438ede07b9416571e49f129919627c454b4563f042704
z714bf763d276b08af0e55ec5ac11665c944b21b0d8263bb19ce621491af3496042eb40b20fa6dd
zcc34234f1d700ac123c2718586cce280df19b7e55ca6458881e289a943a87fbcf4cf10ae59d68d
z808f5a2cbd7f65ebbb125ad06d0cc122c5735d1b5c38633a375ba878e9cc6ce007c07c55c0b58e
zd1830d5367f2710ad06aa7ebc85e1de5f3b99f87d2946e4fad539ce4d4ac4f67ba0ea05acb281a
z7aaf66c28de45d72fbac03eab14fe2b766e14023ecb9c53e35687201045a6d5567972360bbad79
z468083e3994753a2def2275806db83d48a389e64ee4617969341081a8fa1974da21080553fdf75
zf066c6fa322f915b34fc9fafa28c1a73acec695e17ac474a41a1207c670e1571b432f72e97c7e1
z4fcc51d3a64759f8cdd7d255e92a4e96eb38f42979458476f3734eea07bbc2ef48c90ba3218a24
zdcc36f6b3d02129e00cd97f9af336d9478660f1400a2b0cfe4ce8aa4de25422b2555654f5e359d
ze746394a496eefebb41b5938e53f76696e674c25aaa13f8f8b4fb83c92065ee9da24dd919c9156
z44412a6cfa7bd435ca04f238aee6b3054ac66eca82aba633959bfc38bb4a5d27c9ce62a5e53c2c
zeab9328ac4e752846280f81f407967229e54b851b1bf9d745200b16ed7d00526f89e20bb4939d3
z4ffc98b4c74adb69811db134ef7d2e861e686b33e7f5e9f62923c0f9c7dc7fa923ba961fc355a8
zec3114a6832ba1f0d188faea90431237dd73a2181af49bc44db1ffc63a4522042874ac0e8fb2c0
z809da3303eee970e7cd88c1cc5c93dae05f4797f2b6a567e77c2c3dfb8d6771c8985b92654cc52
zc583d53bd09426d93f09745d7c9c69e866efa95df2615b6ce3a80f20427a2f387bf2f75ec6132f
zab582fec2981c5246287d274b8f12f30f69846293c934bd37eeda09dc78adffa33c7f854a59615
z710ffe600626da12a1091d73e95f07a4a06cc61649e6c012609fc750fb70c635c36545c0c227d8
z24214b40e1671566571971b0f753e34b078e0704c82d715d7a2f097328de3555701ac78d9e5625
ze7453d80d5347868ed14da045184246d5a4e1957041c05668b2f8a785363f3b5aec41722c6cdc8
z121e38ba60ee6ea6f025b2c4e0c397167ecb1192a222377fb7ad2d6183adf09a209cb7f21803c9
z6507390bcf43a1bae4c109fc89b3410c0a36d6400ab577c65220ac80707267fa58f88606ed8ab9
z07f015e36dcdd168521f81cb080f5f4bebcc9303946e80ccee3173e4661138a5f15f54dec5a136
zc2a08b62a5e537f0fbc8249109c40ea8ea09c27c9fb13fec17c2ffe5ce1281bad9f3ff50e7f151
z412a1188e8718e9c2f8920277c975240b6ae46de119e9700ada249c3c3ea7c1cb36c8f05599a9b
z29527b683b1fc7127b81f25dd5ae3c058b91bb4e045ad7f7770016752a11b6912353a0a77350e2
z03e0fa166e960cc61c7b0c2ab8b9736077829b61eb5d4d98adeda3b859ad96cd8ef8341eb6811d
z8d73b368506aa1a32c79bef6492d11f897a18529d21b1bf55e5a56b0ec1bf95fa114fbff9cc817
z60b644f4faabbad87abf3ff29f8beb35eb10cbfce16412ffbb0d4f68dba5ae012940c5ccf00ed2
za0a2ccb7ed3a5a684d035ac4527f47adc2f945c9a39f7f37cad3b45da95d6942218877aae718ed
z4e4a2881e13cc7285b9a4fb1b1418818c1b81d26393f9459a46b5280e8d544fdc9308a06b0394d
zd95723500fb8c9138f76ade1477055bb17dafbe39292ec0d3de49b4bd048c601c78d1c8ab586db
z1e265a975f39773cbad38813325d613b916c7f6449535076008f7b62f6ac66cff68864fb94929b
zc3410cf43430f80d1a9e8a3478c127818113e03bedcf656a753446cb216b74158bb65720cc984d
zd5936859272006ccc1f0cf646a07118f23bdd3a9fef2867d42c5ffb006d6abc53d84dbdc0d9cb5
z5ea798d841027ed89f7d4a4ccedb9a6fce9f6f6317111d97891f3b21a7d4109c33a6394aa29cd3
z606a9ff7163daec2adc3ada133561c7de91dd1620e619b8373e5dc19558be688b2c28b70a1f50f
z4f67c4649e092a11db9bdf0b6cb5412c46887eba1b32a2c4634472f2a072d77b98bc1bd4dd98c4
zf45615cb8e8133bc36b2405dac95b3cc130d39ffd783ae9856f3028b55cad13f5a4f0c5f15799f
z595f2171d73166d69dd7213738b8fddd34dadfdc21e43b92ec39bc0d99c313607c424a572ee883
z6a264407fa1945148c2f5130b0858c74f275f9e94127df68f57875809bc258dcb57eae605842d4
zc8047b4ba57c03667deb8579b881f6ec2e1f5082820f1ad8c1de8d01b824cd3cd360cc58ba4ddf
zea973eba788273d9e88234a45f0e5c776d9d87ccd3a511cb56887e3c8436a18136385a13f8c35f
zd203917749f3137a9c7a166ec9ac0811dfa2821bd6327eb67126fb34633a11a7f3ac1181e1083b
z282080082d4da4cf27ec004530ee97687ea76931462b4fd873670cf14a4d82de00521c6205a32f
ze05296a8a153100fe708d1f02918c01caa83eaf7b50086e171fbff529baf13154537bf968c4dc9
z652a6dde96c616849f61c5635d6a075d01088dd0024273a16587162703057a3f4d90e397396aa8
z8442e57f1fce464170242d072faa1e36e747c510d50c6021ecd78c29ccd5135251e33d45175841
zc07a51041924756077a44a303a4820aa4108fdb558a3b52607aa809880b6165e5889fe3748983e
zf4fda4ed162cdf870a2952924237f5637e927847177fe780ee6a69035788b105b18910bc715032
z879a8112544b8b706738a6fce7564eaa54e0b26ffbbe441ce6f8bef640894428afad92475266bc
z76b3ab98bb106b24f7e9ff48023869991e0f41c7dfa47d6f7adab1d4d2cb53ee4b424c5b085cfe
zcf4b017816d745eee55368e4dce8b95a0a6e4c0df71f354c5f47fbc8e54b565560bfde6ea9e1ae
z5417394c2dba468776454366346b2e7b5c5d9b677004ef09effdec9a8117f55a846c2ff81f2d78
zd9e1fb785cd191979e6ff161c87bea7b4bfb6b1df61cc2616b953690f7f15fa06ec4d33e0b4e16
ze191c850fe35157beb979c99416c1cd9062d67c9955eb8c5dfffa860ddb57cfb7739b19e176597
z39506d3deb885e5b6a400976ec03b2dfb605ccce43ee7103c7f66c93b27771a51ca96f2b3e572d
z71956eddcaa0c19a626f77636fe460ac8f113504a144c0b80c26bc6589c32d4c7ce6af5cc0f0c7
z04f90112161cde88c8df51ef8d8a2f4cee594dbc3e160e003a9f7766e870a12d78aabf09e8f854
z50d6d13acc69d3bb4f6cf5332a455387cde4ef21a88e3757288c0c38cdc07ca033be4ca2def529
zbb41de1f6314bad3cb4ff21de0bae633176bd143570e53258178a2a825aede9e620703a379757a
zeb5e4d36847b087a0592a0dc6fc317af27b961953c185de9e49fdec64a3258be60acf077928e6f
zbc2d859857e29ba2064c529ce8043ab359a11601715c4aa770cf0960426b5874e302d172f78e0e
zbe7f8e1def12f80ea2eaab0bd7ed74a9a33f70eaa6d08a84f306054a044af3742fce2eee071369
ze0c23b93ac1b69424762a4939f151753983902fa74c4abe0d2599fff11d7b12eed728550751fa5
ze769d88b18a4dd89dafe0595c63fc83e04ae17d4ab23a5ad5db7dfd626ae6684391b976d405434
zf12fa3eebf4cd9a4d801772fe05d37dfa6f83d682a5d6e650dba31bdb84c3e0fe173a1aa65c8fc
z34ab0f5c07b311ba6d33141c712986e2b598d6a28ad3f1d0cf0fe314ed15160ba98523e4393ff4
z724a19564d06166cb309ad377872ed4973855301878811ff0dbe16b03d67d83f310f121aab5d83
z41ca58c5289ffc0bc9c1282f150bc1fb86bb6a6f1089bb5a82094ddfbd96490806c522da223492
za82eaeea5f65632d01053151a63f3438e5ac3ceaa3900f45a59ab3cb56715ec7465461b4718420
z053c7e3bd61b42a521b7b2118c32f4fd53525fc909c79623a357a7ad69b5f48e3fdc5b3e6ec4cd
z08fc5e44671d6778acbdd143519a4a417f20a3521a05acacc170cc01b04095f17d6a692f98674d
z646d72f0fc10fcb828d74b693044f50ea0a079e54e3bd4218640b18bbbd7cde2301b9e6868a13d
z67fc3db2ba7a5a7865003269ab24da1684a15765f9f8ab839ad8a3daf9b0568cda40e712ac5e68
zf0bfe589220bd19e6e20f8f65a641b4bb1180e31ee15a237c2d1ecf7b8237ed50383765a8ac5d5
z6b43d08a73e51e62cfac72c05c4d09ed7512102750d2d91aace250a75d16c92478bc77c4b6dc9c
z42070d1e9bb840042d09b949df188ee9377ce51f714efb4b83b322a51e275407db717d96c6e8f5
zc14ffe382f11ff706cba9545d5f1b1ca1706fb9561734645f47272a55c9fda9e432b36f5bc19f3
zaafd7ce1deaa3b8b6a61ac968b8ac729fa68911f8333e218e7dfc102124b0bbc54f29ac9440fcd
z2027af58072c137d9edfddec24a261fc61d9dd210970b2f8f6173aca51a119f819dd42d9d1a2dd
zf471a9efb64db18aabc723678d63e0f3ee92d45b373782ffcfd637302349098ae186e12b8ab56f
z2a475834f9ba4f718d7dbf610c3577b61a9be7e1f5a8908f0d20b5bb4d2365f48605fea0028ddd
z5e6b20f5439de97e686ef039d1f5d0934da6eb27591bea73a1596192d3e1e448e7833029ef4acb
zdd0faf3da73a6604e37192cca8c322fc028ff3b1caad2a1d48391b131829f239f87a85793f3a3e
z3150a064505b119cdb2c64113337eece11812835aeee66ab8a06f27a8045efcd8a3fa7a80b35b9
z6d86fda4e7795f24a20b5a10b092a2ec652018562b64ec16409f6d1eb4aaf6debb982918f1dfc9
z37739711f01c9a6b8ca836472dec2e8849896c3d7bf317b4d1ad50e4bfed20834603f86565a49c
z0495ca8cb006aac3f335a2421f0905b4948d53d3434ebdda7f8c0a63844c5e024679d551d8dec5
z3d35825ae0094b71f073c052d9d60dce302de1633ea8117f7394f52f6ba74059cda38023ab8334
zc562277ab087c1a115682f7c829e1e6f7004dd383b07051c9a48500e3588a671d089a00dcfed8a
zdf4763116bfbe320cf759d4f0605cf2f11c4dd577fe20a31b79971cfcf27015be63d7d1b0eced6
z02fc8f8d543614684e84f2ea490ec9b55d990ea567afb373d84be1fa38e200d002efdacf999fc2
za502838d940d328c51a92b63f2f2253e514e1e6a62355c5ff6415307c6179b26cd5bffb2dd3ba4
z1f51d6369799c62f77985f4980a6a888b287a76720b3d79a4fae822817935b48f4e4e5183a8124
z0b41f363ea07722237d793637642b51f94c27ad801ae9842e51d7b9351ce39885df7e0adad658f
zed81563bd2b94ba0322dfbfd73c41d5d33f93770b8822a33c6219c4212f08c908bc1bdb2e8a2b6
z4d030992f13e53bfde51dedc1732cc955eb0678980faf0b3c9b7772590c52681a7af9d37722725
zf4ace8249c19e40d810401f8f40d3a42f4f8a2a137e73da3d59cd983c409a9ca0a6a200cbc59e8
zda9383e9dc9ae247f271d338cf0a5456c6d6639e4373ffe2c20e0f7fb3f27fcf34bc47e06a991d
z2f61d2d2daff1d53e19ec68a93e29f746491f7b3bd39b39e6c5dcb5311c52ee10bca601a820dc2
z33bc2323caaf413f0e88e1b17d44c4ce2b1e0e382748fb79070728163cb9e495f3866348001f19
z61a6cdfb3678cb79795b9ecdb12331a812ff6352780b558297d624c23a795baa8ba4bf37f21bab
z432400ed3eb9300db5f9f30b982a2a4049afa1957810841ea21161fad1439f6a2992b0ccac6183
ze70e41a73c577d63686c49e89561ad4a7f2e604f2b4fa948e65567300e95bbd94b34601ff157f3
z171130145b079c100f530b591a004c20428fddef64fca89efd68b1afab89b1d6221178c755d471
z7a403b0370b388c7b3cfdf1b80561db3e841f7ae24fcc2ea00db3a1552a660dc98b160f4b1a364
z5aabba32f55f2ab1916fe709dd53cafe4b2a16844f65a20c7335ebc135a4677bfcfc1df1caaa8d
zab3dcb00a0b3a62e1b32307b4ffff8d0d2a81acd3c9b2f1f17516266211ed472c9e8e3ecff93f7
z971b52afa6fe6022bbe9e5d66719e56f5715fc995266eb6fb0ed7c73a5d936e0d33a8af992b122
zbc2a2a8fb075ba7427203984f7932e38c4a6d9f124cc72f6f46268f1aab835db372269e49fab6e
z118f75b1def70daae85cdf9de361a3f8d814f6a6bee8eff3c57a9c2a3940e373e05cbedf813419
z436ff5dc677f8e53f447ec779e8fbfdbd6aa96b5b0e57da9fc61de1e2b5c54e35278d3c4d1d97f
z5539e7c333b7e65f45c78fcd1fcb1ad2f47052a4f4bb20897746c4727270ec21e3f5a5cec413f0
z821ef32d548532568ad81bdf2c0407b1b1f7660eae964dfff8ced3522d18165a142a48cabbc29a
zea142e646926709164727e95771d2e7e696b3405ac30da841b0a559a610bae34c4b9c8148d542e
z1ff403dfa54bde8391cd9ff987618ce2aa3ed73fa59b1c5505dd0f90bc4fd31f0859f2a183ada8
z24cd562fcab452de59ee2a4b42bcbe3aad7fc2a24ace9883439d5b981e8f9c66154894b5029332
z97dd5512440df91df71c8d837d722e2cbf36cd7257ef8e94858ee18f6ef7f5902e10701f3ab3a9
z53e3c3ccc45b4084cfe93ec547268aa53a5e371c4392e736cc15887fef77a358420cbaa3a2742b
z3d5d099e8a371d9912604ca27582a0da910266d18ef3f19b59e58653a3c62b4b0c859c4a110959
z7d467346982da5080ed095247768290a4686f9e3b196f1ecc7c93bec4aec79963c122b38168509
z566a0acd128164093986335784476aa8932502fd6554abf55f9297e1798129e5bce6397f157405
z9f2ca39a8a469ae68ab38d3aa05647b926cd31d339dfbb63f3d8be5e0d58e91522a457720ee670
ze9862b500b63493ff9fa43589d4d2742bc97f758216acfb9153101f38a8f417600bec244f3c51a
zdb2841018863014defeaeb740ea7bc11ece7c6ad8adbb6b099819823a41ef32529c9ad61a63a03
z7321087c01fa84e7400d2cb6f65dbb45f4f13ce589095c8c597da5ed6b7495b8c483b857d429c2
zcd76a74a4b30a1fddd31ad41a1352b48d0be938231333279e12c122df08bbfeb4123331b370840
z386a758066ccdd98f70528938ba4c681e205fa65e5cea50dfd1a70f70bd4b7f63d9a75cab7faf3
z348c31c30915d9fed07d6850f6fa8f7ec03c930a3d5d2757e9e88a2629c6fcfc391cf9846f4943
zebb64543fbc05e472401835ef608e8cf8e13ed40aab536eab1caf0b2a16e412b00d3ce36baff35
zcb7aa1e7fef2b0922969aef42f83322faf8aac6a6ce7cf1a399c75a464de583c0ab3936c864299
z388600e2ab215d9a6adb92093f1e8a200976270324ed58bd9cea5146801bf25b794c1bcf58d6fd
z8901f1728c3a11d20a0e8c8002400ebb453d4e9098b5db6a4367d572043a5adb6284fb371712cb
z5b16d116bf63ff0b962e6839710d253d8181cf2afcf85c8d6651f21ccde93cfebb4c9478b5fe6c
ze95f0ff89b9508b6378e6567d9a531df5128097b1ef482cd93869531070df4fbfe2fd36c43fb77
zdae1c493b6076e3df5020a8fef8771e01b4edcd4631393051603fab765a9640f73cd26c7b701f6
z73e58af44c46fc7dc239472cdd852e179524f7e6f57acdfa3d18e06b53636e5dd6b99c80e86864
zef3976ac0bb67e27ea73fc228e6f7de4c06039c664d6686be1f6b200727f8531e4eed7d92c6624
zcdc3576399a46563211d189337b59f77cf5fbd9974cf587d27430704475c0732470dc2005cc2e2
z6312913b509915156a4c9fab03dca812eccfe2ce6e24d2044a24e71972aae1212b592e4eaa469a
z02f63af10f570afcd50913cf9b1136f159dc4b18ea6d8808dba0e231c1f633b96463bed082f054
z5d8deb9f59d6ea4cd86b8215dbef384791875d2a9b7fe017a3c4805bed89dcccf38192bb58a8df
za3efd46686450638b45b63eba41d343b86f8b2c81dd3ecb2bf1223ceb87edf9b4be6379d271b2b
z73d10a68cd6cb31ddf582224709322dcef6394ea91107f2e649943d62faedd7ad78b36e3a49fbd
za83cf79a25ebadb735e26031fc03726d8bb39277047554cba032c3d3c4cbbac82606c5851fc907
zd71a3fe255f1a0774bd1a112a6b32c4aba5c871649da93b554948192cc4475a473090c0ca6576a
z31eac67d8754738e6e8a033ec74099ab0aa96833c1cb891ed0277d4e4ba0992ef7f2c00a001fd1
zcf1ffdf86224da97fd5a72c279481f3985cb70c089ec2fe0fb5e93dac6d2cfdbb8140f690b6806
z6d8542fe603256d1964034766bc544e6a81972ffc35f899d2683f0b06540ed18ef6fa7aec407e1
z154d55b313c158d3eae6eaedcaf9d62ca0e6dbf1d5c73691c35bc5bb2e038d5d01863420dafdc0
zc5c1992fdf74a64d20a1bab4e75c0f849aa5a0e5b8a7248deaffcc7c845aefae7983c88924ab7b
z928135f8303940846089a0db5c335800dc71e3667ceb0ceee42bfd0f3692d068f51c56c6cec53c
zf429d06f4029ab99ef540228376dda82bd74237378bc6e2ab8345c820b0c171c76281bef7062c0
zc4c05b4e48f68cef66f0258701c78ccf5579a31eee5008ae414be61b3458893a2f99d1dd5a7c3a
z30d28cca66576f28981ca5b0e8abdff40a7b0f3dcb7bf518db85f9cdc4373c121221c5172cbdd8
z38986c323d5a99fc7efbdc82c3be93ffbacf551a4eef5a151bbe165ec18c1b677d777377e0f729
z61cb95e7d2f35ba7e6b8b67ee3c937e697a60853cd4f2740ff3127eb4f9095705d02493975c20c
z64ac0ef3deae8f50c76efb915b7e6974f35047a71db3b0dc98304f70913fa348e960338dc3040a
zbef447ec77b4d99ad2f80f50ee00a84371b9a68565df61077398735c3083806fe63730465403cf
z237661c210fde8135635a13a224fc010ee19291f3fda67e0ca5447b2437ca554cd39d798876b02
z34b4e0394f65996ebddb2f64de2f3c25e6e449546ced233e6d2f9909dbbbafd652a566184d291f
za28ecbf656d25f2b7bbc937d78c28fe476c9e7aec68b42991d2f1d944d781632bc331aa6a85732
z8b78c08727f419cd970b3f25be0b9b2b68488e2c540a0c8e1d4f3fcb640f8c3943ba37b579ee15
zf5fee38b478a98b8840f37eefb5b67b9a69d93e47d5e9aefccd54f587b2bb062cd668735fda41b
za48be3be4bdc103a046ec6ba25a3ad15036e085c484edc243a0cf11216c8086fa85be10edfd09b
zc71b740322557d668d89b469db390ecfc2c0973dbbabfa664307ae8f85a4808dc1e5bf5c6c9554
z47756c792f74e3b4b45eba67b600c1bf479e7dff53fdc82720c30b46d0909c5e00e753bf61fefb
za751ada08533d9aad0fd6c4ca9637fa244a5de1d9d2afa01aceff8e783f102dcd887d191a5ea7a
z041e825cd5ee7452053fdd2ff18b1608799874047e7e08610fcb4321cfa5729065d4b1913df304
z2f916fa6db0a01d7b172bd89753f2a86543dbe9c61a42f44fffe7bb8adab35caffa3c93d82694f
z908f9aaa80beaf9601ec44cf4941f03bcc508c2dd0ad41d99f4654812f9c9d6e4192bd800eeab7
za9acb9b2e2c15298979572b3217ac3cdb7799baae492ca6a2638fbb86184c5cb494305a6929f2d
za2d17af53c91437a4a3e2ea9e6d7ab6adee9692937aa1d59a3abbaca9ed9e0aba9f90f65ff9c42
zefab4456412195b6c2e5d878a9afda84eece5f076e9d7f8696e2c4cea09a5a5a016ffa329bcb01
z9a38bf16ed656e321c8b82267833f81af5e39442b19120f3b5025945b50475c5baf79f4bd46f03
z64680416df32cfd63a43aa4870585cc70743144ef8653ffcade9a82f93e51b3bdf337b18f3a224
ze86b5bb28472d01ba072fb258eaa455e47c7a3fad1086d423657039286bc591fbdc3d2f343c659
z3d5e13147b4cd5a9858e097c2593a21d75fe139446239d5b08b48937439b002b9cd226721105bb
z4b69c1c4a4d493becc3ca2122ebc5c614eef1d3f99d16716fc8aedfec471df83496373ca8d9d81
z32d8edb266ad4ca4fe9a1862c2bbab91c89b20d7f91fdc50a6dcb257ad3d9d685449ca4a700014
z291a78ed34741bf09128188829bfcd26ad671b47cdf6fa5f17d3dee3dce1a389a417924da90dac
ze97be9234103ba274a7caafbb153d6a69cacc1f928d15897d30e791fd0534c9e184ac812a0860f
zd669678221eebdc006431a2faadc86717d1f404d59c97838b07d40767dfd5663011c424b2f059c
z46a799456f02edeaac703029e9a0a3229b2684f13b31effcef29e83dc19e077ca983d29ac19005
zcc442935776871c974c730755365924066337791e84476fee936a78f894a5d61e701eae12da155
zedb70efbecc6082defca801c0c20875dd2eb412f3f5b4d50ea3ce162f742c9c50ff5e42b7fd363
z336df44a3a1012e608257509b4219c9283ce4d69000761aab0a16673353c7119ed12f4aafe54ec
zd608487513d1417cec2d1cacb5bcb3fb02a27bc68cf1fe2470a7e5b4c1a7d5bb6f764244e901f2
z98c8b7f219e8f761f1f1c5df76fceaace37e1709013350bf3ee3e5c331a1262e102876d2bb96e8
zeb0393408db53ecf7fcfc192d43d677ffce29e2a3d265ff0678fe3dbf28d26b531add5b0488ebc
zd0d2783313d9f3bef2c7fab107f92d83df02846589ad24a44f16fb96c8e32e0414dc2d0065617b
z2ab4e4aff1bd21e048c2fd4d268a4288c048c6780cf33b608ab96bc2b2e942b942c4fb116bbd9c
z7e5d6962eeb2832d015e1019360cbb8876c3d948187660bad2b13162597f27df3d18f582447f5e
z73904a87a28b6def32a0c7a86f0a2603720ad80c4376933c4662c598e033504444e65d69224720
z0c798eb6c75db38599704907241f0ec7dbfa8d49ff76d200166af6fdad713672c2bc947a1a0b45
z032ceb99092cc6c6b6644592478a59bc859a625d7d1fe390d3084041765da530ddf21c05b8606c
z7cf8e87f9536998691b32d21952c318924cff17b0656a60082ddedc1bc59af4321700f266b1e0c
z457f9eb0aaab315d64f5c180c81a5f0cf8eba9ce8e649a3dcb3314ebd6b4f42aedea1d843d3e99
z0406debdbe21aa0cf0962bc7081e7c2de1b52d073bff4435680a89964b01911a0ebe8f69e6e258
z2cedf29f169262a57f740990aba26fe6dc66aaa5a522a6bca80dd32f90aa09d80b9a2a94ee4e7d
z0724d9b4adb49eec0ea39352acff3140f0763da539abaa1af833cf0507e36f02e4367315074c62
za4776b2ee3724e49fa928eb5e3e31b7171f94c3bb67b7402e060ccabad61926e01bd019404bf77
z2be3e4d715384b8385269851742070b8e1000bff5f395be8c3428694ca5b6259a459cb89c470bb
z288a213a9fa64eed95418a283a49faf51f65545cce2cc2bdc61584d8f9752700d0ee809c2faada
z1247b0e080653d92bc7516bb34c696eee480bc540a742ed07ba1f9c91d1306c5141212279becf8
z67684d1b83879a66156fdc8ea7ab84a9104af7133285b81fd845592a379589a4726b66032ef4d8
zaa607ddd8c75757cd90c5c985fdaf77798169180eaaad2b69b984344dbc8e5148becc61fde5d9e
z83c65fabd17aea907873ad30d8c6a45a46f95e28b13ad75779cb16f8d64011ae9f3a7ffecee92b
z759cf9aa0a7a6779c108c39adb9e829471079573715373233abd362554ac127caa93b4d67e3a41
zae5fe4b533c5879d2ca0db22db4d9664551ebf90de6573abf1ae9af562dd0f24711dd9f7cef716
z9e37f86380a819b6f9178512e774bcc49582f95619ecbe92aa0dcd930a23944ef5ecc4bf54f86b
z5fb3a97b3cad1857c962c84248ef79ef3d79fa0190f903b7466e21c625a9a9957a1027333902e0
z813fd1a478b8e40b5cfdcf418efb1cdca81cd25f121ad8bd389023a54c2ecfbb82ca6a025a2caf
z27f9ced8cc29ad7b109dab3b069088f7563cf1998761b5f25b958f22b80db953161a1da7e8f7d2
za396a64a7b59a36100d606938781e6b80de79657aacf53eba0c045596dbeb0768fe471487ae1ec
zb8379c5224478eb88a17dbb9f863e11bffd1b98615630979221225b8354844e67415c87e3d50d3
z217cc8de5f63987376b31491dd0c5305221f4e9aba899ce548afa0d0250f489109253b969d404c
zb2c5e29c692dc9b7018b65882c94083a1febee11e64c78dc4edae08a8df74f4ab486c13ac4fa0b
z523ea9f72aa19921428ef278e0e99698b1b501c3c46722d95c9e61a11d7398031917662291bd5d
z1343cdf26b02ae637e40c8a693d00f554c0a0de0cfa766a71937f2fa9a2f8e5d65fe1a15cb6f92
z0a6d48c7463e2e692d63396349766a5e760447d9b6944220d8c55f4587d5081f83910a121a28dc
z4950d1e93381eeab6e37263fb87f5a0d5280af0d54f09943d978b6de429694700506f87afba318
z628210e196c4783f36ce36fbda333c1ac342da4d736fae8b60d9ad691ed2e98dc3dbf850390593
ze37e47d9c259d774595aa843532db6899b162e88cf69b2f20766196d98992a9db1366a9fdfb1d6
z8f8b9fe0f68081c277472c63d71ab59770f074d06bfa8ae5bff110c28cd839ddebdb2bab97e68a
z3dcf0730a759fcc8df673f629cfb65f3cd15f08923efa11d16b3d54801372b0549a2b7763a550a
zd238c84d535c935318987f580358fbefef36b183729d7b0942161bcf7572078b11d9babda7ba3a
z7bacb5ff457007cc2e94c823e07d2c718d2ee325a654e0bc7884ca9ec76da87036626dad453db3
z269b756fb8460702ba750932f730448dfbe4eb7834601096b935e5657d08db9a9e0bacdc5b9022
z6786340bb14a76d12552f56133856d906f5511f16c89507ac6adddad3a4c89809a17cc268857b0
zf913c3d18607b0db4364f2f9fadfadfa4a11260b1442a078bff40e6f1ce45ffc67cc006e37dd07
zbfe3a2abc1b73a0ad23442875e98a91f8a6618212b614148553607bc0d0d2b0f7b177ba00a0da8
ze9be6fe1ad539a98d5d0989e46fde3c050b835b79b7214bdd7c366edb384171aaabcc4a9dd1d59
z91eaaeac509d2bc068abf41e6e3375a5f97a2c9913ca2212fbcde6feb44bc4629f1b65feefff9a
z927f38f2b0e8774143f9f5ae386019dbf43e48b93efa276ee23a7782f1782c8b5959effbbdabc2
z79b250ec4080d4fa92b886685212d9d9a34b8a98839db996254b268c23f11af86ffb2fe87b31fb
z55fbf4eef5b01ff2f560b4ce858d656e8db69a564b3844380e9361d997f3f493504c4712dda8ec
zd4465e4621b61aaca935593a7a7114930e586aaa61ad9008b088de0ff12116a89a0f73fd1e7df8
z3f7dd5d4822bea41b3832b6bc1f6081f0df8af2c2bf35016078076134e8cd33371f151b534b4ab
z683be3841c9ddd9a6b49a45a64f5de2acfb7d50075e4a9cb584dbec41223905b444261bb719689
z259b7cf427778f24cf0cb5aebc281baa39f23bcf49460ae9b678454439c9338f852d72d5f32fae
z426a0531b24deef1a96511d23738b37cc1ba02cb2dda47f1e192032646aba7661655e4ae2ca99c
z55142d85d8b86547f7322882a370fa9191f23a89bf7d619b85dae3554bb840f99c9c7fb0445386
z5a7743d0509968823080504ee421ffd59013b8a556fe768cdb46e2b69513a256d1c3ec39173e3e
z0c35d4410f198111932f2d71993caa2962aa7029217687bc19bbad9c7766682ea281597301fbd5
zbed0db54d2b21a933bc786d050ea38f3d06a7790498761da71523c9a1b10da8101a478659d7f2e
zd7ca19332d04b044690da86597f5ef11fd834a3dccd2787817e7c098e9ae643abde22d5cb1cc5a
z699a9bfbb1f51cf372bb998cc7032bcb6ae06d9368e24024d67e9477dc200f634f1be4ebedd2b6
z6ca2e962177d997405420a60ae10918e82472a2e43d3efbce56fcb7a37cebb0ed6ddd07371e9f4
z168f2fae5ba1b143ed5a7bbf4d19603cb214c3fda037a3e9907c69dad2755655ec84dd76ec376b
z0ea4f94c343a653390ecf248f3b793e85b1a7227f1f0fdc0224c949b2a17a598425c4756d3136f
z081bf609370e76ef2f344e935f61dc901d164940faee64ea45f7bbec575fa833f6ca17b8960acb
za826b9127f380043f5b2e73a463e9083db7b15d2c698601adb39e437b2e51532572d4adfadcfa7
ze2a41038acdec1ffc9f216bee02f99f174a5ddb6a77e445729366b86c732e1116233e33bb8b3a4
z5a044bf6ddf2280b5950771cc9e2b0560e7f74525bfddfb88e79e71726a5a0609a8a21f75b8105
z58729e72bf20a36ddedf3e253f659c8335608898e78fc006c21d30060dd8c4430a650e689868f6
z5fa6ff01a58f8d45c5c7d3e5d491ba63ea71114946b21ade545103f41cbb21cbb6d2f18756015b
zcae9e83d4ef8265273eb6e1f6461c686c72a1838966fa445192098fb27df737f668cfa17d2eae8
z2402341a06873e1645ea82e53820744e8bb34a2da41d496afb9a61f5d91f1e04562cb2ba555df6
z4adf39896367bd3219070974a281c010016c15b4a023642428ca106fae9a64aee38e201f445fbd
ze4e3b72b3154d40dfeff40d5e50ac5d77fd1946d4c95e857ef936d4c132390ff0486f9bcc6f18f
z9ba967c1ae0b028706b066cc9fda88af059adaa164d5bb10204c6e9d88d8ea9cd1d13337df4b57
ze9d9f85c33bf40f282221ea23b7d23c901fdb8cd401871911b61ffd916deca7cc112abc86ae9a8
z2c2e0f8f6ce5eb77b8d3d90d40523b50bc5e1af62e3593e2c445dfeaf95bda8c5870140d4d2429
za6f823b280b48057e823ba1a48a62bc6006970deca80014f9446739854c9bbb7450a7ca6a25cd7
z8a3c7ab367601af8296cc2c8ec5307eeace2ff8058bac7a2ca03286706a65d5c675a75f77e4707
z44263fd673432baab782a2064ecf9da02b332cc33cd2aaf29184ad09441e31a69130d44af29ca3
z20c91f8d19c6e00834b950da8eef49a9e005c28c2d7fa886cbf0d07e9fbc3a896900a46425b172
z53019c228f19d3e5aff40d5d4de31fcf2e4d7f8ebb05c10e9a1937f45d5e8f1469fbde48bf0453
z2427977be5526401259ae36c8dc8bd23c5459ee857b8b580718943db9f31dbe79e298338ffe784
z15f13148078b774afe647e3d70c33fbd4b146fdfb74b06a2be4d3beee85e47a4f924fbc5cab7d4
zcd2f9abc45d57e399f6abdb87d42ec5d02bf613364055622c6c51ab64a1cd80d7569a1faae05e7
zc144e52cea8e2f72b5d49fb954e19d6077e78d6dc6bd8bc4c816ccf91cd554963c147330537bff
z88dd89dab289ca9fd8c25a5859fc6bbe8ce0759cd9f2d50b8f97ea3c859f4a61fdf376dd14cbb9
ze3444b47103d8899f99da0d373865da03e03f987bba7bffa497ca1ae99819d98106112b4278eb8
z311d2f39a8d9f1b4e5ccfecc5f927204a031fc234ef7310000be6ccb14c5f969eeeb5276799674
z5172617e81e27efb88dec9202eb43e7dc1b796b34d811014da8fd82b74414a52e1d0853d082f0e
ze1968393359c1bcb14221b8363fb087c7daf65e5eb95bb857988863e2361aa78525e3b4e3c104b
zfcaeb00636202d7e3600560efc1fe24f822e343ac7d83c4b92e4ec709bc99d467ed1c3de8b8c06
z226398f437db4d5b374a18d9d729229ac1200a08ec71e6459dc8709b7b682e615edcad43989850
z816392c99010fe8096ba6d154bdbce360915658c40e75d3250ada1e95765c695b0d010e88ec76b
z80b37dd2426736fe6f61c6451ff4389954b0d991779a3609875f5f82986302dd42f5592b1bdc8e
z5b58f874d3beb7d976600433a1801164140d6d8b4ce58b3ce6b3dbec6d16a6591a2ad37a75d748
z73e13289150c1f119e462f6978493e4fd0d5743c6c16a77e966b269ba462f0f3836efb33137f60
zfbbb54a6bbcdb58b947c9cdf68d88753aa853f0d4d592298e60aa2e81c37114d094b4cb1811d38
z210856e22ce54256dd8e6d6a2588f59e847c21cc3e85f9115fbe0695598654639887e72fba117a
zaa595a603694a2c1f0b769f031cdc2aa09ab4e6964ae2a2db9cccb1d498ff5f40985d4b3c113fb
z916a3ee3527b1fc66f550c41b41a67d29027115e3eb602c85655327d9aba8c198b9175b7e51c32
zfc38c19dee8d7a086092018818fd6c33773597ddd7cb2cbec8dd855cfd83f04381719ed1fcdc14
zc3ff725313f8b7bc50ed44967f85873fd92aa782790fc5b6394d5ab0ab427c9a2f4b853d3a84a4
z51b07495db6b953d811f99c755291668a810416e213de9bfbb5dc6e48d02e10fce742bda47e468
z7825323d5958a946a37ac7f0298a908ce02f022e81145e3103686651bb15f3f0c780040ada8257
z604f04468a6f6dd054cb0b1ec73e53c30771983e5cbaa672481b9e33951494053a7696c438542c
z4e62d67bbad0d0d393d113350db85b5199ca659259201121f510d6ef4020ea95693ab7b97ce799
z08036b8894d50d189d40da6cf922865b47f3ee64b45db41ae0cb0a9cc02606732ec1c0550000c1
ze71a6ae9dac351a477ddba60ad4fcaa8bcd7cee5633d2e4b90547500817301a96687a579effbc3
z0dd36dca501af1aabe466bef040811499b061c69f092f186f0e63a61c283a457b83bba589c5f8d
zbeba5306303972d8d4abd51463a67d0de291de9901041d3ddc34e4c448679bf7e9e93b40323ddb
z10fad313690005eae4469197718ddcecb5fc501b92b267517d63ef843371bca7ba7798f0961655
z9d1fac79b5ec3c726c3f77c0fcc10ea9aa9a9a9b344202c199a72743c39227a42fbd16241a6b34
z4bf2d6a5cd55dde45622986a13f72223f6b41cae4f535def1e2222bb4abe33d8a5d959e11f963c
z05c4273b6eb2bfbd6a2d5f05448c86cab1405740380c9b8da949737f6accb1984c955ac3f53d31
zafc7ea32cea2d04b1eb5b612c31a8da3572e520d9aca29533c765b2ae6751601274c3a1d1a57d1
z92de10ac938f422f8ae728105fe4c3057a1af8d4ca8ff0ceeaebaec58f22d435f4becd5e727ab5
z093243ce0ada11826a304327a506b57aa3d632d1bd18dc24d147b683bc27ec9d3d4b04193e93c5
zce7704fdbe7b8f729d1fcaa31af94e4ac18310670fb1cb4a2c2ec7eeb3bab768f1909532b8ac7c
z77daacc7af883b1959c28531f1680597a99e8cd3d98b3108f174c08210c25bb4c6a3e30474a269
z9472b7d20100f6a20a654368571cf4b9e332ead85e87390d10813b4897039f0b580889d97a4864
z943b90bb11d5e388f353d07a37cb746ea35b29a9e59e48bd2d05fbeea3f29cda221f2fc24e5ca2
zea622b057e0e66939c4c7254d505dc331c8513d5c64488eb1b114d695647db0eb31003f0924b41
z921e8fd91a51f79893f89483b146415cadd0789982fcadd7afba1123ffba4845731bd412d409da
z8955a4d95b5185a465ddd081d33b800d0b368385839e1ca6836bd5565650dd48c0523543e70c68
zb9a4a436dfc549112c4e939049ea6d6698c41b5a453bf50088e961350e221f1e5e2ce6c335e596
z958acee22300b48b4abf81b3b21a7bd1f7202a7fc82d8dfc736e27daa85cac5c10644ab54bb472
z76ce14ce62727f950b7d0a7739b8634ba8d57133f5b24b3bb4bf0f760de4a3b83d612fa38fa353
z01094a1d724b0b2ec1cee0f5a99a7b7c28841c9754893187f12c89c70574c49906f8148f99417f
z2ef3cb49290829d2f79795a637138fd91a5d25c39e6e252cbb778f2b4b66665bac0a8fa78964b3
z06cee88a526f6c6330660350c277a7cf80dcde4c19771bfc3544a8d93da5043d3e018c9d0b3ea2
z8b582b4b973d1c0912ef10b08d00377877bd5368a70779ef1604cd61b363bee30c34993c5c1ddb
z58b15880407eac2b2062cd58fe25f6e6ed4d189a5d6139650ca1e3cb5b6c816b16a792057aced0
zf53896b3bc8f2406098c531c1077a5c77e224f15c3a888e18da717441ddab51e4f681affaee763
zef892a290ac54fc9447b945d21d381e9afe8ea3ab0d50f43bbe3f9e741454cf8c1b919d6bf3aac
z254805818cc9af6e149115738108f9dcf82f60f4284acef5daaed8ff37ba617dbfee4b3431b670
z1b999147dafcdbfff5484bc4fa9f9aeed3c2ebaf41f7389139e01d71bfec3d2c7cdbef6f523932
z32da91be553ddf5451379a953ab8efe2a62d11269ee56eb2d0be8f915452e128ec501c3fa2ccf6
z604d4a49f58d11df3993fb3c4c21a5eab86f6f1b2f119b7dc36353ae02ca7c5e303bcd50464c3b
z67d081287f2446b505c88942cfbc768a3729f92e3fd83788684f83890110ecf1a86078071680ab
z5a6f2ab8445e280aa6473a71b8a07d3890f58e35b7c93c705a903ace3888fb27227e3f1627bc36
z7b61909eac0eb7c98db6afd256cba7a7e0ba38eba4e82a6813fc6f793ca611d41b036ea2e65691
zc48b2b09db29e8d2845355f781b3918ca21aa01d456b01938455c18cbb5777b06ce78901157d1c
z667816253aa87b46c44a854420a5b8d3dc88a26f10ad377e64603f9d7c2df57bdd37c0de8353f3
z74f8301a0188b4231c75e643efe3e1893092af17ce2381ca7984cdd8e059a48b84f8bb8eb65aa8
zcd057f355fed51ab8a50da898a74c95e1ba7fbc64af1b04f8300d5c9d238bbd8186da52a863759
zc94c7170a64a4fb5c5e2f2f57c124c200dd02f81e6d666cb27532ceb257b7c626cac6053daa3db
z79ce4537e3a70678db1650c2141b91b029e95d7cb952d22d217458244471bc0e1bb861700d5cd7
z9f1ef8b108348fab990fbe5249886e9382ba4394378a4bc54c76d153fa80320212e7e0234b345d
zbeaf97440fe103606d67982a09b54a87d3c9017b6d2d4c89446a64de000fe301df693654148bcc
zccedd75951350bf871aed9d6d4390050849ff34718abd656f7ad0fac36ca77e8f81e05fc780624
z6119bddabbff02133fb69a3aebf4db30b135514a3012f3fa4b33f995a1194a84eef6884c052234
za3664d80a831fa1c07af3974a440dc17ec6f749a0d3cd436205b27f174c7e5393061dbf03823d3
zefd93a267ad9961371536bce6d32ff5c81496f073b6d6d5fd7f591f9fcfe11869f03cc4d2e21cb
zd83c6fb69bc1508dd1e621f8ea8a56650d9c9e7de310789325040baa4261b780a604c544ebccc5
z1a0959b129b88d910e4a64f0d9c17da6c25423a7548150db02d87e3cc582f20463386d23c17442
z30973c0fe2d657d0d371574f2f81f35559b3b2a1328b645c46aa85c6e69ca42cbc51a1581b0862
z16793bcbd13255e24646525cfcc173d5cfd9702442367219f480857ee43c78ead53cea49069919
zd7d1dd2f80bccb9fb353e44247fd2641e9f8237fcc75b107fabf01a9f13c7b19c7da36cd5a47eb
z21498959177533a259db0ddcc542f6da45b534bfe1f69615f0bcbb3c07d45c842a118eadc7a37b
z35953d3e58e5c116fad858112437dfd537a745ca901ec7a5c94d583cc394d7b5cfec5d8482698b
zff2113e3f68ea037141394c3bde9fcdf1e562ff007be38ec7461463f34cd354483411cec3bc64e
za6ba8e64f8ed077afd933d228198b44b984f8316b45320590327abb8b9bda77d2ca7371e6c1e4b
z0bc613ef680a5e3a53c8e3342f963ea0f6cca6ab11de7a7b8fd549228160fc9e7c2da185ab7e0a
zca5746a7135c41e3effee90a28f3283087b6baf4f654d62f49747fe626c2f977178558b010a226
za947e282009bd122ea9ced9ae55b550dc7ea08061a7aa2d2a72e65d7f805d136aa356fdad0af34
z7d3f2558b5b8279789a11042717eee90271fd40ade82985cc6b57de3bb78920ebc7150310dc956
zc83da08a0573731799781b3762ec0f8968454b4a48d93a888d588c7bb500cfc2fe2a82d3bb4808
z670e4c4cf47676d2c13093afda92c5bad27d8c7d1bd073bd12269f40e1e44345f1467d93243bf0
z5b7493961254418bddf4cb979965736895ec466bb3fa0249dc1bcec3ac75e7e1b5af96f3c1f218
zf6dd9072941bd8a9c45f1a45eb1a00f27a50f534e6786ffc6a75c27f0ca0fd11c1530d54389cc8
z1012aeef798ee04df2435fa344e298a7555cadb7fa124ad8a4fe090aede10cba067f2173ef8279
zf0579309a25834cad8dd4cd7344fa539eae1105ded57df50f1abadfd5515f07daed23beaf77e73
zc99c30c3db65b6b317a3e86fff1a72699f5ed3c3b4b1488a6cf1066923e185ebeab0de6aa671db
z190d8c2f7ea7a387c6ad610b5f5f7d0e14b9b267e8c97118e03a76b33ab750bc9e8457c42d48bd
za90495ed150957e7e414a6b05c4cdf05b520a7745c6462ae49a17874cd6fa9d6f3c7fa64efec31
z10f1d386502f7cc4b7caae498b7ed4107207d4a78782ae65087bb7f4f1d2badc23e6c899637878
z840b4b0bf03c6b38bb1baf676067d7d8177ded074c682b21f1bcfadbdd8dd07f99c5a90a0a9324
z46907635c0ed0026a385fd281fc0e9438e4cabf5a44586ececd015bd96c5ac273e0fa8f56f9194
z034c06351a92a3a2f53c821e4a66e7e84647cd03997a9001cd4371a2f90644e2f6605169203b8f
zcee397ce3045fb0dca5fadc8de75282ae1f27569cb3d14ed8509217e26a7e1273f25a2b4ff2add
z09fa8e1ee09b076b68e3b83d6a26886beeda6598a75647c82907af1cb8a37c2c200f6ea86489fb
z26d4eb90c047e0a703c95841f7a8bc8f2757d0452629fdfacf1d4fd9ba38720530878306311bfa
z8ff4723954f6b70247717c34be36e8cd466f174ac157b4bb7222d2f8d323433987bbe6c2c1d98c
zf746c9468102712d9fa0b2605c26e45d90f6563d34c29f83efdf20d09070df40acddbece422972
zb94bc93733b1ddd1711fee5f3991324012eaded42624a44f48628c795a14ef7dda507404b6e19a
z105e9c7ed292775836564e0ff5c18608c2f91e7e9ba62334e31e2b162afb2b291bd56b8308c17d
z79b0a79eb0bd992afbb2a6d2043512eb72c750c78c76622e2e1899d72967937719fd5f44564a0f
z45bed22689b3672c2c3631ed36f20fff2ba1cc1cdcdaf7635cec4a6979c9adf5f9e8305c79d738
z082e2283054656c3b734942df5947617af9f4ba651c7f56891ca0516e34af01f6431a84b443290
zc1db9ea83fc8c870b94936c3bbefeea966b76fc2fdc41fc5858950ba69cfe5e3d206dd30b3073b
z623f804c7a0661febe06d67e5f7ff8bbd33ee8c09c451be69693fce26d2da519bdffe8f24d3a90
zca97f2c4f1f19482c10b690f5befa293f379928ae6aaaf1d9ae02dfc8680f1e0f4b0e19308912a
z39373fc7190981bdfe4c092467e9737b10d9246a3c0d7ff86cb40b8ddf423416b42937ca5632b0
za84f5151bc3c92f0b24f077946a1d69a0aae51e58b943c00b8b23f809551ca5a17fbbe7921bd9a
zd4793c56ae057947713d8a2a94954ebe1933ea2fe899ec5fc974d8448a3d0464c39bc43db52dbd
z5db1a94a9dde68ecc65bc542a1d3a40e1b0ffe181e548cfe68551a41fb7c0fb5ec46253e82e00b
z414f9f046def01c7a038307899ccd7cd6f4eb38056018d7b486b6241086708ea1ad896cc3f433a
za3a09a25a906910f76f5eb2900918120b7d0399c6f86c8df6aa5cc48968824c953228459ad5d4f
z9027063e16ca04f128699b4aa84ca04888c9d65fccab19b51667936493dce2a8a74f6d90e79b2f
zce9c3e956baa90f5e9f248abe27520cec7ecd0db026f1545429a35143cc1df2943711f38894be5
z64dd23370dc728d192d3d8d9ebaef4b7bb68e0cf40a75a4623fb918d41054a0e64fda04ca693f2
z694d9a49ac28bc70c4de7a65ab583e514e80986b9801be1408b63eaacadaeea6f88866474862d5
zf8dba7fe3f8981ff2d9bf17cb755ca878d722d23f6e4a9c10b9cfcbce9779917ca76d9a050aabd
z2f156ab015e1916f45231237c0534c5c532f56ab0fcea278b6c87d2381b5e4e757d84bd0fe8870
zf44e3b3a1b8c585e8f7c9789276ea362cb832334d516d018a915e2ed20713e3c6ef42a90c46868
z7f5dfbb93cb663bc207ad26cfb890e1c5cca1dba2bd38a78fec7048580ae9bfce5237d8de6b973
zca980fe0dd7379e26baa8df83ebe47fc8bbf5b5dd19ebc7ddc6303a39f0dd9c1ff2a9837dfe9e5
z88434b9ba8e6669cf273c82f87f6992b807a5561b30ba5709da106320145d647e63072da302529
zdb7dec9957b4a9d4a942cf8e6ad53866df9a456da2f0ee795c868b6e9a9173f78186207233c9b2
z4990f1e74652779b6021e862346a7b148229886adf947db831ea998ce5f7bd5a03fe707ef71f74
za60d02f26a80cc69d065ad692d55fdc40662a047d838d7e7db7cf2c6558d708799f68bdbcf7130
z349913b35acab25a64c2698fef47f37734d4663092704880eb7a3af777903e009388d6f3a37bd3
z9c4ecc8657eac5f6d6c84ecbbaefe2655de15023e24967c4086fe08a2cf5fedb4fe263df0a5f00
z15a80538c2f0b8772b4c0e560da9d3ca3ec3e93e9d26883bf55f5f2590037a8162388fc6f7bc6a
z21ac243d7dc959cc9cb6cfb7ba53b1db9778e4c783a723234abdb50a391f047452d787eca08018
zd64529b769bdbb0700967afdf04b83d44c41e1cbafec6f7f850c9d6dcc8ffa3d9e592d61d872cf
z0e5f9aea04a1a87c2b664110455a6432fe8a9531f7aecdbcb3e5e181de2a5f293a579bbdd810d0
z190c9e0c28a097cda4bf1c38fff4a7cb7ce60bd8133ce920a3977c2476292d4924d0d833fb14bf
z7311caf7dc97ca663c3d516f0b4f562fa6e22ca47a35f5bd44fb9c1fa84d78ad8344db273f46d9
z6a3f334e2e41a503cef1d32ea8944407ce45ff1f46bb5ebba905299597bd942e01c4c8141e4d20
zcee307e6c7c813a4a6a7086c69cccd619f4e28c15255d9b19be12399f4a5779dd3ccd9e8c582dd
zdc303f3a733bf22b581e8de9cd86798b6df20aaba3b19294da7cc39cdf5a5883f2b23a3df880f0
z4ff21a833dc5cd793787cd62d2c2b6fb0db9a4222aa3590344783143b730094ba2deaa4aafc5f9
z02afb7443b6ccecfd32b53aa7e367f01de258dea3271f41031c1dd027f6faaaa295cfb78bfc609
z4d729a0d1836e3e5d0c35e98532c2f590ea18d8a4a1ab771d4cd8cbc514a0f60cf4a3f91c64ff5
z818f6f4f1e3747bfbb2e0038e74a589f02c78b790f25334de1c6aaddccffa3453f283c4aadb633
z1b14901438222ceb0fb21aefd6b7f013f2965d320ccdddc9bdf8b08efa0cdacd67e0c082dcd6b8
zf629e1c71dea2f2db245b684fab3b27b022dbfe6e06df57fcdca1af9cbeb12cd4f1c1885c19752
z3988aeb779c42c704f9514fccade785a715204437a6f1eed26206de2b9736cdebf3ce09c1e0039
z8fcb0e5c267e8d646025b0d024f78e3138a5d5c8022e709dcfffd179173437884d5abcc9e4a93b
zb9ceab2599a2eabb0b2b7b4d69e7ecc35e50c83f0116ffd496ed4b395cbda85b35cf09748e2774
za9c3e852626fbd3a25eaf8a88d1d7990d1cd3c5f7c0adf4b16f0789c9a9141709f97f385867204
zc4e9c8e0275e892813ed3f6168eb656d2688edeef25deaa642c9cfc98495c853e771807b7b0a56
z30b130806aa298debef1f3f9ed4132dce6fb15fb7fb5607ff2480ce3d068f3eaeffd654febcaff
z03e6b4ef07cdd4c5f16775dcae6b80eec4eef6082d2220747bf35a8aa20b8d1a2c07430b31d4da
z97958d9ae70f04c27ac544551dcb247b9b5d1f228aa25f6eb3a977368915368b86e59d05b545be
z7d2161b16207a67148e5355fca1f90b66cc7bcc137b5405c7ed1d821b7ebe92f6c40eb929ba3b0
z82602fcedceeac507c06cad498c7a8ac72dcc55b325eed277bc5f696a22337e492ca51a7f140d0
z6ae649bd0cf496cce7e7da0a8ea21358ffee02dc445a9f4f4c04034d7d91b780f68eae5905a293
zbb026b3a035833269472ee5ef4227c8fcfc4c87e30c3440b06f47d7abc0317d3b0767e3983de24
z89b35406260b50d2ae1ab871e438be55b5604ca218d95d30866f8c9f8e45994532e9e1281547bf
zfaa529d664bb2a3cbc5a57571bd38d466e35f7a43a5df16eb3511d24b6d8e965c45156ddbec427
z0c9ee571270b2bdb263613bf4f93e03bed09336539bf19f674105e8aa034af70fdd537b80dbf73
z72ff7e7d3b29ba0e022a945eb0cb0b589c4fc21aadc98906d29d5a80c35f2aa2362a89af1a9e29
zcc8bef5194f738d6de377910bdb7c033f246b23e62cebdc8150393270910d7458efb3036cef988
z1d3ac033e96d49c3651fb4bd1f15cf67e07000cf9e16cda26adabef3224f3f97c0f41067291a42
z50fb659917ddc27b337af5687d7937dce1ca21c851886898a329b0a83f03709bef6dc2c7b821b5
z904d6e4a3fcb6dcedddbf45a04a12ff510e7529c93392427e80cadb4ce0c434e968608dda827db
z54fc34c20ece67cb0131adfcf0290799dd8c0b145ccf6c3d4b9c7bbbe9df38174e31f46430fe4e
zff53e981da1b8880a8ff25682bc5e7eb9cefba306751b5346a441575901c904fe36782a5dd4f48
zd91497ffeccfe288c925c73f68af0a4385b5c60452d1e344ac349af0be08f4c0987a8b1e3a4b3c
z6a2f34d4ae499e040c277f97015c47e3dbaa00e31f81f46f0ee5ce5a0e317ec6473feed045f104
z927a4a7ec44b7b7ea3241090d0243d447f2a75e52ad607eaf33023d697ad5f92c655a672dabfa8
z428cca027c04f362d3792aaa3ae5260b3eb8f80fe587e0f17971247e7c5f320d23ea380ae7b6d3
z36898364eb8d71a6fb86230e3ec34a245da976b311b2efbd5ba82d86dce3bd9c000dc7addc1727
z45be34e998960e426206aee37f57b0557b4e2ba5bfe66492c554148cb2e3feba894c76b15d3960
z955795f3eeabd902946833b9445ef6c7f0cd06b7e4c3fd3f05f1bff7fe6400083fb59259346e8e
zf18e65b4db8bd28805306baa4ebe3db8b88f9302a90d80c6a30120905f84d961087b345a498e7e
za0a65fc32a3cf40fc936ebb01f009734d8c92094fa3dd3afa083a26e824b52aa64f11a286800fa
z723889a28559d3016bcbcb4b9fb7111ed11fc63999f39912ea39621483ad619c6051eb942e0eac
z57b4214f8672634561f7be06e4a9fa1a8d060a836613bb070a093a78426fda14c2345660d241a6
z24ad3b098f4c1a8a291cfa3b459f0b14e7382b795c3b176867fb67212a6a0367758f35da70d65e
z742e3b692cd5dc8ab01196d4e568b1ec1e2432a875b038da5cb6e6be0238b82e0235ce11d42059
z61b1916b55edbe9ad3c26077bb955f92078b44353c9bd3465876a9a34dd0af1332553c567f37aa
zeab45f5778c810b5f02c2a23c055bfba1f10cb3a1c816f98176a70d28aecbbaf5ccb74f9afad5d
z3069cf7b7c1951b72e78239addf0c93a8588b879e01158bf39b1269798bbb24c3d8f96aab43cc0
z089674b36e53b15825d8272ac368986ad3868c429037106748e5e85e8e8bfb385a525178f6e9ec
zb93ba2199db81da4a0d9e2e2313df12648f402dcf410f74f08130510ab2a901a6e4cd362243059
z21866fe6f8e6ecd48cd98eb4cba38213f0d0aa7c75da6f15834c194943603072308d8ebe5e184b
ze4220d45569b4a679e5b939db5b11ab0564cfc3abaec86a49d4eecdf71abb19d8e8d9683985777
z412211655d2e59946b2858c4a062f3796cffbcdaa00a9dc4e6c711f63f1de5eb00124616191f7d
z4975107f34cb988c15846cc9b5785eec1a29a26a801bde921af089fdf531b9afdface5842ff855
z074c98d68b43b960a868dce9e1568ed04eb02840f263a9ea08de79d7304ada2d557bb07fff59a2
zaac66f0b4503e99b20a0b9aea6717ec628d3c068451f2ed5c007761e47881cfaeec910b4f0d2ef
z02f3d30552acf021f471e81788baa37b353ea8f5a4a3dbc9af2213229d30f2bcc7ef85f6c136a5
ze9700bdc7d1fac2f60cd0b23319f940c8ff5d8850a2f1f73fcba21bddd130efe1d0231f9c5406a
z19c69cef26d01168fcd9cbcce85b97d81a669518d91e4173cccecd0639fe8685b9645fbbda1ce3
z964f83f50800de8ccc2a98483dd967d69b35f91ea0d229b0cb69c8d1a0407be2e205cd5be3d904
zff42139a9b0a08ccceaeae644a81ede5c4a2da327d132100e620ef3d589b425fcd048c44f46607
zb5fab950a12836ac4da856ac185e11e7b9a6e4f831adb949df9187c9e36078a6fdb4fa7a0b9f35
zd7ec8a9fa96aa14d6bbe5fad307614b768bdb234d6638d722d019c3be110ecadbbb04872505bb9
zbc530627c320d651520b9f327029921f55b024f557b0ad767f1907e829cfb1ad2f8d6362637783
za18afea8d03277076de763079f52b64ec4abc72f25be628a7996a45d2fede0bdc078c51724d562
z56f46abcc9cb19505b900bed8d68dcf54858b8e3c9cf9b91ed8b868e38e72387f17ed9d8df667e
zd052abc02a97b51ddf85c33cc095cb2c05720e11548a0bab2ffce772740ee655a91e5f6322eb5f
z92207699ede2e8c93eb6645bdd7c70aab85d14a7161798bf57385fbf44e3ebb617789d77900368
zb6bf0f8302dd27999374a6560e827dcf7f651a421851f36cf5fbe9a1a1e70d74282288a5aaf45f
zb4f2cb8a5f05ee98db014626c2e0ad6bf54cb7b30caceac31d3475df962061323a7c5e0f33a2da
z07da0f01227263db6a2e124690f6c05d33104907a4dee6fd2508358973847feda41ca96039fb63
z652e228841bfddfd01246da6c9012c7e164ae8dbef54f1ca33c1317f3a276cac85662888c9ebdb
zac68c39fee3fae516711455c3b7b6d5fceabd4701fe90a80306cefc6b2bd43b9b4467cc236d558
zb40009d75c6a7e88d04fc84fcded1182f491b5b8af47813024db9fbdcdb1aee07ba3d6e1d127f2
z67d44fe87ff678f8d970ca0c752020cbaf1830f57acfa97ea21223cf93dd9ecfa52f1032c00ffe
zfd59e4ed6aecd04e962f3f8e767af5c75ee1a16ef79e041f33fd4365340f371acf5a8b07173865
z3b2b43afc5f14314bd5799c5d9c6f9a282104b2d38adde1075fb303b09e2c020ea160f9ff4c208
zeb913ffbc7fca8806b64f7ea2e90053c4b4f375c63b5dd559713c06cce222611f4088d880c7429
z84b762efd10fe5500a07eb635c83ba6f8dd628eae24e1059f9a57800dc302b9f6b68179c2f9c99
z8ba0c9ff580d3a6f7fb40984194bdd913747d6c0e2e30f291d842b3961fc95d3f3cc3f2419d1ea
z3c489eb95b4854fa6563b7397b549a81ceb8a9c0d8c57be272e71eae9c38a10930060ee2a1f418
z4fdc8182159e25541d7c4ecab821a1df270d3380e1e2b5d2bfef4e7fdc0e17ac7d4815b3f95d54
zfd04e4250bfe9ede86da0030d3db35bbc6d674d2eabd4ea01ada5338dd0a479317a2a905521137
z715cafb4679c7fc49c00fd09c3fc818992444478d3ef3c6c5288f476de81479da2bbae2b575102
z2f4d6115f76fefea1ff1bdeec2cd789c552d4dd3a76c718dd0527f6a65fb82966612e8eba4ccdf
zc430696303312313cf4298cdda05b45578fa179468bc367f7b79a61c44cf0f0b3133b236649119
zab7b524f3f780052f8acb5ba2d2709dbacab631f14268542a35476dc940c95fb93527134374357
zb0d01da3e537a73f52574b356aed5aba7d6f3c7b6d041d0198d2ee6e30d1750525f36c528f7713
zae6639961708578c873512f480326fa11cfa2b3d2c264cdbe40a83c8c3c39c4c1921d2e1c615b4
z8725c7881e879a7b3043a7360514a065a646b762f241d7282f3113941fb05d4ec38b7d6501c46e
z0344d50930395acf1d70c8421dcc986ad6241bed0ab86bc51161b6ee4d656524d944327c931baf
z3b85df47ef7d22fdc55bb01b9a6552b691014ac7a3671883928e5762bb4d29b64db2cc070664a7
z7624df8e5fb82bbf3343db9dc2b779ef677df1fbce41ad584127919bbbded5ce6eabb891f4c1b4
z2e758789e0c9f46ae3fc32c68cd5ebaff3d68608f571ca3eb9d757d0c400455dd1526d85062d76
z2cb4dcaa08e8232a22516d7d6b92b8fa19e287f7b7421ac2a68d13acf02b252ee1e12c1085e745
zd7a57cc2463c1c3ff4d3687477679c4e8c56443bc878abe45f4af06b703ef462f390af7abf2ddb
zc1951b68043ded369da7d0fbfbeefbf81f7bffddf3dd26c8f31fa61caaff45140c7ba7f82c7fd0
z9a8edb7954e3dc7f99442c7df692cc8ecaa761376d40fff64b9427385d82cafaa3f19bb9f5882f
z11a1573d548d51a77af44fa44d050411c9d78a6685a8ce9d7aa0a04c244baa0ba0c7fb1a99f6f0
zb6367fe39acbb6e02f8f04d08761010d5fa99818b4fc215bb3842bfd45a5a7821fe9740939f827
z7fe1360deaf60d8007b27c5bc3ac393fba90c9a31138649fdc8ec8783abfe212406fcda371c973
zc3f2966d04494690e3818058e125073f7c11425f87c2053091a08a535f85c50d7996809f96ab57
z294530b383507c7fbbd19fdfd54b061c31815165d27194938b44293271c02d51beb20f3989b504
z76d23ec53b0e56b3d361d436943f7b91be7cbe78d0a5ede2b81fb2262c2e6526fc37435d7826b2
zb64986dd1d0d607634c338defeb58c6406f812fb7bb67d044e9752fac709c0f0f5a4569b4c5af7
z2f876862843e71d4454ff4c5b51a7d819b46aa4860d9e54ccc9ffabafd56cd76c538aa0ff72787
zd37950bdcb148b5d52cf3cb574456d9ce6b9788a3b255c65ab31787edd1b69ab6c1197e1dd84cf
z9789ce85b35f35264cbb404f45c89cb36c3fd22aba4a9515a7d6e77c500b4282fc9653af8c8509
zca079f76d8d80df0b23c5b267bf2af0675c25c3e22ec99fc14d368c72e4591da5b3639c41d6182
zb3813a0525afb7d8ff7fcdb44d5d45a266c9be62d4c8be209c9804df4478eeb8bd928de8ad5a14
zd34f7f441b04e40c617983adaf40319e3e924bd38010b91b181ac029bc51653210eedfcc1800b2
z1c36ff24f0b2ed5e927bb767a7963eff05aa86d6005e2f27da5858b92dd6976998e5c89ced2f26
zf9517245c7ec17e4abd083f0e9582fda45a0bdcfb12fe271be5cf38b9a9c93245471436712abd8
z184955f9b2ea35941ec30c115b96aba5fe29de08c0e80da59d20e5f0702f122b13b6954b5b4224
zc0821b9b332e97c36c9d78dc283935a2b7d23b2e5a4291b49b4708ec3e6db35f35379151ffb76d
z77244eae0a07299f7b0201ac2eda3ecf905d1484d93f803f217faf067799feffe5f9b8aff30f72
z32da62439a08b8a2176e98a95980d4d51fc8dc9cd464dc4e0e9930ee9a794beb7d529eda506920
z0ce069be2e81e8eec91fe2037bb2057b7c883e502ce970cee147847690f5b83b7c847e67a9100d
z2913f57fd274a4e8529e6f82793579288350aa78733118d91f8efce48cbb1362ff9a872dec0324
zad1a03ea62ad9df6878ca0dabf5a9ede8a5c4416d5ea44393fcfe8a0c938fa92c0cc0d72dde45b
zf73b2ee9022c82fff916659936e20d6fa05d916665e2369587f167ddcfbc250375f152fbb166d5
z7d5b9c302c68da1d441004d5bdd18c3a4384bf35938737cfc750a28ac55014c673866edb832816
ze0d9066bcbbb8a07dd95c155f10e82ae9231421aa30ccbf942fcba195b03469ed3c1c91e650b4b
zbbbd6283ab63251cd77250d819fbec542dd4da90ec2d9ce87a537c576a88a5a1a76951e918505d
z2b20d9af87855b896645d3ac4c0fc703915fcf81395c14a1d07abdf1264818e8e912c4d0ccd68c
z462216ebf7df45fd323c769ed2fbc2ee6b82940775ec55e58f237f8959f51de39556ca7b26b971
zddeebfa3c93b80b9065efc834ae5231308ff8ffecc2624cb4722c7f4b5109c9bbca00796e4a621
z2eb5491d5aebb1b0113bdca1b46ebbbc36d522791e8f6bdfe1f34d00fd5976a41286e5b2ee63f4
zdaea9bcd336664daae24fae3242ebe65a16e8d62084d3ebd94f867a40841d93fcb67146579f40c
z1d06f38bd33b17b096c2cc12822b4183d357d5829ed4eef3ef3f5917aec9a4dd7c3f71ad21a66d
z5092e558da2061d60b7f9392e56793b0a47cbb5b5bf585c0df5109e545932a1b6d272c9a604025
z26c1db28277ecc238a0fd8b5f7ef0213003a0a4f260dff474e98d61e9edd24a0127c03e28ffb3b
zd8b5d88517f07ccb93d3568f63a6a2f25704b37836f45bc54436f2f5bfba838618b1e1268f43de
zea6e68736b89508ce7252556755df8acf5a5d9c3a44b06c627e5ae9c6a6abac6c5f7c9a6e16ae5
z58f1210d29ad9462f923cd060b970f4d9703ad514c073b9d438895a311f19ee124d145c794be02
zea0eb942323387a21cd62e55a37cec99f31131a923c2a5f410950ec76d129e9dad8ef9325ed991
z1b23bd69dff31f22382a54c0de9898d5a7667a50fa337dac6c5b5d1c2788e245d6d1ea1a248ffb
zafaefb570cacbdd4d3e286196342e01daecb6c4d684e0164cbad9ef79687e010a4e8dc2c0aa723
z7f1cd97edee790adeb8b18d086b846e679336a0a14ab385d3df0dc18735ebec265fd39f3ffcf08
z09bc3878b28ed09d93386386e541127fdcd0ad16a11229e0e53261796e961d1329ef72df0087e7
zd4fe3ba6a6b33a7ef8842b640f96f1cbdf791724f1833c2cedcac0d5afdc9f9ca1e0ba53fe3758
z71bdca4a43f6d67df093dfe569a5f3532ac4c657fd4c006c09fbb1a68b4b9ecbd161cef3e9711b
z5264a27d4c4e1b71ccb71ca66ec71fde28059795849322f7226f42c416b6895fc67ad8df7f7511
zccc71570a6a8cf1bf677d62dc380fa0128178e1ff764f766006ab306d2df0f60d82966a1e34803
zf55eae65d04d6e81ce23a500bd3c86fe47ffc7fcc952e1c6665838db310b1b1df45ebb4c5c3d1d
z6ffa2624e5ca0aa0441114ea50dd269bc9898a7e4dd325118b59fb24ac1f438a6416a2a03942d2
zece14e400c19994294cf98b9a17524657f6444901e9d92c22acb1aea80d6d5abfd6b510f4a851d
z12385a66d2639ab041ff1881e08164095c8230a10045f956a8b865cdefab8c6a27e0fad84173ef
z8b674f3ee095321ea82956236e214b28d8fc32476d9dea406440c53c896542e1ab8b60c3d1fac9
zdc58fd29e0114eb5d812b17042f17e4902024293c5f54cee109161624404ee2131d0ca6b438a86
z22884e208bb7ee8ce2188e8cc29b29b14888660fe1ff86e631ba7b140bcab1975bf539b8fdc4a9
zabe34a13f368e1929c30627510b8c288f7e79c705f7b1224157a9729c164ada8f6c180740fefaf
zbfe460476d716f2143c7727e66645116d4a8eabff825d84c143149c10039773a9a62d5e182059a
z4b324d4b238770144c31ed9f077ab800d342e92ec6d2261b168290bb63fb1ff2092c775e0ba33a
ze3a4c2a3ca2ce3d508c9929442e05dc2641892240cfe15cabc778fbbd3d92322e39f88202ed7e2
z7bd5b070b76964b15d89d686186e635bac53191ab85830e20c5cff09b79aadae7e656ab27be442
zb1698d39c0a2cca1870010f7bf3780be829b1d4da16bb6e8308a50f414101fb75f0b747696d032
z704b9bc010d74dafbbc9e46761af2356b2de8105b9ed9cd0d902c55132237c28cdd7f4e8ceb25c
z1cdfa0c1c1a57a70be69a9a936b33ed2ab0755ab375a0666e91e7c04589cfb876e1176d258cb60
z5392011d6e61e628e23089b0c1782ebb3413a07c74366303e555a6d6e8da900e889beaab626cbd
ze35569b22d33e9117b40fd8f8516bb0a638a6f2d8dab3744224c9c6b97c3752765a0f0a356fd41
z16813f8700bfc8e7d5c947b2d212b00981557fd7a54938df3d4614c2fef2c3b31408a51ad2f8d9
zc1332ba862b2a05a8aa032a311a7469ffe1ed78bb883899d4b59f41b584e2c784da4b6e45a3ac2
zb517351c7e922cfbbd0ca243366c1a1821a66f1bf7f15c9c4a2e45f6fa0886c3cabe47c98cbee0
z558fcb4624b21bdd0f9d36967559b927d296af272d3793743c127de8301478549a090615e023b5
zf39d1252637a02474919adfb0a4af9ce58f0227cc5fa7abe5cfa93646575e18ca340c2e709e20d
zee045dfe2d1b2970ae3f946497edeaf01ee806b837cf9b7361d0f51c732d5191ad720ebb7ca4e3
z55366f262616062c26468de95d6a10fd6e5826efe7889b3524a5d38fc0ef3064edab4f50ebaa86
z896c120f5c042a7ce4658413c7666d8eb52631a929632de5114511ba14c2bab10b682e62022c9b
z076f3e3488d3cd5563cd881752f3740ce1670962c873a3d13ae59d4980901678d5d9c57962b7cd
zc4801cea1520304ac95b36970c7396e1c00e844428fc17e3177312248fab15d97793e1c7679e67
z6a6375252aee60410821c52d77ac781eba279e99c54f6def32b808515f88a3d2e7e331254fd8b9
z7c963596585693f052275c4995dbbbd9e866bbcefd95191e3cbde603d8b7c5769cd7d42109895c
z2f6a6560333be2471e18c604a34fa8828c574534ee6b64038c1810297bca28d17413cf558102b5
z4adcd1208492cb4d10c0cf9817537707ee327d4f4fb5ed317c139d62e383b1515ea66261341ae6
z40de1b2e658d2d9e3cb54e8ab0f710344f835f00de4f7170471b1033bb5748636c8c684578f3cd
z54c2db05046cac36fe972a1f4edb58c318232cc9b63b7c97d8139d24365cae39709932079788c2
z077ad23d3d7618008333f1ee4a9bad814f66974c27eeff7dccfd3599763f9ec59b0884d638cefb
zf2f2af363835fc446532cae8409d49f8a20e999efbb784d49aaf4eda09d5a0e35473321e04168b
zfe83b8c59e7f26695a78a0a8207b6844cf543703e831aeb2280921849d36e096b56668d7d02500
zecbe692be4ec6b34a84e81dbdc94f701132911f824584d5df8b7b5036c701446df674c20326a0f
zaef96a944274677a081cae832992e60b6c4abbd702a9adde35acfe4fdb8608a17fbea04f111733
z9101c45758045cf8fb3cc9b5a681fc9b1895b8fdda485a6fcee8649044c653424ce3272745cbb2
z93d63ba38cec40fea7935cf5c6376baab5965aae8435b5d97ea81bcd81dabd577d96c7b8762d53
z6074403ad4a4c086ae6c70a8aa2f29cd98658808092bfd96118cb02a23e868cd8c9671d2535f00
zd04f55e989d470cdcf252793fa749258a9a4a8ec178ffa4065713d1c1ce7cc8b8fffe915385eb0
ze77def46790ccb9069924a5aff25085ee07274833d96075d7573974089692f29a2ff784c3982c9
z7c803f135b28fe468ee396464e25b977ffdd04048ffe65f9e434c9ad2b70d7d16de67ebfff6072
z7f2a362d406f84cafff1b1e485fe75ecde15de3db2454d52cce0374eaa1d661d6f2cefc618eac6
z5390027b3f4717e2be65122e5561b48c0483cb0bdb61779173920f3acb60ab04bd91d779ae3890
zb79e88a3bb8b2f6e87086d2ad4c52251828faced0b6406f69ef8d684bfd5790e04a73b76b0aae5
z402ccc53cd855540c141ae941ef772923f331848216ddf0612a7f031cf6395863853df6e3f7622
zc6b2bc702d79479aab944501f83d15e40bbde7b02b50030b1ce0d03f31d15ba2c90031d33c7790
z21e576d0ccc44cc109041eb8747e397a4235c20a008ee32851a92c92cc8335b138bcdaa5f8daf3
z25c956df900d25f6bdd5c014d682715a4493499dce1c55225d2390ab2b9e6a82f7ba7f1fd5ad64
zcd9e33978d79e103bb151e912c3f43809851bd98ffbd3fc4f9c264a9786ec3fcd4fefd8a3c2c78
z8ab62819ae2238d39d39fa36b874884103f41627ee9ccaa35eeacc66630ba162680c34a7b68b24
zd4d5dc9ede991db4d495d00efe446355e44376882f2cba7e95810726d21be86bbae5abb45018b6
ze75265f00b219a236bd08aae632b8d544555f42767f7212e370167c33cba2be6319bdfed3c7dd4
z49cf692b3f1054e7e6a0c48652f0a5fff06dbec2014e35a3bc8220ef2cb0124d53d816e012288e
zee9c4653d9b4c5ebc77ccbc6435896eafa2ad0c7c392e85902c3bd74478ddf49201e9ed644c046
z8fd73da93e25326e73c16ffbb27fd578b8e385d748dc31226b918c7f59c820320c03cf02e08a29
z6605508a0c3f3137f5bcd97f28663f540642724ab3b721ddb5c68654e9270bc3c214f091aaed4a
z3062d7b87d33f8c3bf66d75379ed58143f95da39b79d95cffa528d2b796bfb41e7ecf25d9bdba2
z9a6e45a46b6d4e2680c54c4a90a5dd5811f053bbcbcfcead2d282dbe29e90b1ccba91a02b55e1d
z331922f651a9914a4c975551c9d070499c3989afa7e3214308236e4283fbd605cda5ae3144f6bf
z64d316e9d43c0509b7424067069c31c6e4c55b32048671321edf1d51fe7f9dec7b30bc657a9eb9
z1ef720a1bc400ae648460894a30bb6694759f0bd49b8f70d777cb70fd738166f8a307f491ec048
zb98a2432fc9181810b6a60b0bdc75bd7cd9441de17bee86515e0bc430a29727050cdb13c7d3ce1
z872d738331d323647f953f80ca2c09f9707645dc845b466423eaa4298895702ef926eca337d13d
z20973fbfbb6542a485c5ecac1658446838d815aae387fd9c76692825309e1d1b90aad03d3d9537
zf4ab2544eaf0c866a29c9c090f2cb9a4ef2df23ae02a844f83f7b287a0ff77ead1b0696568b5bc
z09daea9a67dbfa6f9959866a9fbe4b8de6379183a30244732407b9462ca1e2a5519f06b278459b
z4cb4babe2ccc0d4d9117f7102940252f0f899f820512d09c25c130c53fc8806f0a482838c2ab1c
z2e8c0a27de7d73e1601e8647b04f6f6f47e1b6b55b7cb325cfb6043a06902cadb496c929787314
z91255d1932f87f6f4e9693caa42ebcef3a799506406f361e5dbe8655c5fb7c8b796548fca2f2b3
za0c4a5fb34372085fdbb6c9ad61550ea7c5e3f95856781f3427b49c79f19a28ffabbe8aab4f9f4
zaa7641c81e56ffc4db827ea4964a8b8dbdc0feb6ee3c9c41b01378db3808ed93a9781226143879
z1b603e6e938134c40254273bc3d738f163dc514731cc0988866e81c506eb6dececdd2468217507
ze5cae8929ab4eed942df7d04deca34e6a3fce906d44df5198f8f899c997ed72d3924f37d585d77
zcd8e365faf5f6cfe02d43e8edc7b955dd5de416d9b854a9040eddc76b84e2bb7fa2d5af13551ec
z940f7b522c09f15968b9b741a655cfda7346d921b559fd4b0e6672890939499311b991cd2fb303
zac5e52875c7e59061433acd47111044e2cce5b7cdfc4e3b4ae74492962124a80315ddcd128282d
zd71f2361b57efafae67af1b138b1cc1f2eef09e8a5f1640eca57d07d838e6a16d29a2a729ef761
z5def60bf3f975caefbe84e34ea41b0af3ae7c0bff67b1c3f0e6ce463acd8098ff52d0a4aed492c
z9300b40f027b32df74c968f037040094ad699cbff92df033ed66637311a21c7f0ce65fd1996f04
z91078c593301d8fdf9b47933e2be02df49b3efc59e2e2c897bb79cdfcb18ecd0ff8c76e0d3ef11
z35e123ffb3a6bd01949e5054a1481ec10d070e94f76124d4695fd69397db8f1ecc7d6e7d204f65
zdb0a004b671c6fed3266d68766ace8dba630804fb639264592725760660d154676cc7f890dee8c
z2bdfd311e697259046456499c78bbbb93271f51bd0871338c1606158205f5509eaa3241b8117d8
zc6c6024c999f5c1f50b9f9f0ab9d5bb8e3c74069475873babe9629cb79d1715bc2cc11f9317b00
z40b8c1b600c6d9269f84ca75fd10282e2ebefbd60e6529d096f4841ed3f54ddac8fecb35398868
z2513cdb34c9d263a4177094cbc5a34ee72099d371dec373059a3f948b112e2c4fb0454683d6634
z2f0cf11ec724822826cb39a5fbc811c439b615251c48aa5cd61defe0be0ce36d15cc58a373f172
z1723563b5da9f180d2402741ab07765433cd97b3483f83bd98c43e866566940943852d87eb4cef
z27441891708843833254b57ea3af03f78a91ed74f7ef3a2aff8b6920a469d47170b5a8aa8b86a8
zd778da5fd9e68c09861a78de99d8f39136ac89ce2669b0f5c0a02b4938f1b6c0792fd7de29c450
za285b16887e7f1cc8fda5654de59c56711fe153083faa1487ea6fb7aed7ecfc6fe7e0ab5cbadc8
zc87f3605b083490b719b330df6d4078435c1ee74f31ed0ecc7ed6903ba87bf2fe864583e834136
z7196fb903b3256989a711cd1fb7c80addbe042f16ec5101ef095a1994b6dc9695df5ccd46a3afc
za6e798ae4fdd3347e4c9ce42f0940f773dffcc055ca7e8b1d9f47c22a01d317f2f607ccd5269a7
za036527ef365f793857de213bcea08ea62218a285e8cab23f3266476cb671c223c2493286a9a3a
z2c0d2aa9b1d8d105b87cf7b652748bd8d346e0edef8d25ad49e1e8cab2ee71799a1bf3adcbb00b
z228f6d3e5432da4a2f31fc5b348d4c3d1f6ef048b2681848aa5cd61b8126247c8b0a297e62276d
z5e98bc8f0c6ef8f8ded3bd3de22f1c2d179f7e974a78b196562367bda45b9968f6827b5a8fec2a
z35ace8bff1df04ddb2620ecfeb6ce1cb2dcfd628114a09da71b56d322c50e1ffbed3de52af125e
zf91cbeacddb735fce0954b1c76e7dbbebb7201793b30386b4e69b1fb0e2291133d2988393713d6
zbdf5068eaee2f2c820e154836be17717166a5d0a51a87b34702858093123affb1282f8278b7d65
z7d2fa54f1411d58d4c84b2893ed6f6e86f0506a81ded9893a85387a4bda5550554bcdda7b077d9
z651c74d8d768def129fe6e34072bd4116246a0f4edd559f5d047e2446089deb4b1f08f55b4f67f
z801cc448d26a149d05f8880c3c9358298c2b5ec2dd3e7434d113e5d62370bd4d65cb86125851d6
z1392bf1b6ee15073b4f618267568235f7339fa9c1e20cf82c57015513724eb8cf50026c69c9a01
zba971f67145a6135f53974885d9dc674f27933d89e94e3c03e955cb51dc8e969a02541d81b9415
zd290124e0e22776b5ca81efaff528fcdca717c0c20a5ad7e396191204172c48016885b38222a9c
ze0997fc91641268d267a4d94cf99a196d992c49fa0e858a05f21d2ba9e828169971422504fd651
z598116fade6296ab047b390dd7c85cf4fe2a0475c89935b5c98fd2d6f670c0188a6d804b1ca8b6
zd75112a747956f6d7e6c7ac859e70f7f58e6860e7de0f617a966ec7efa6b3640db70cacd4e7aed
z75f5f8fb729ba9a0ee64608f760dd5937cd5be817c169ecee2b5d5cb86922057eb5a2f8622916c
z2d368f2e851ecd983fe957270ee378b094c9ee509e2f64dde4f119bed866c15db508406698c11a
z79aa159c28af36a69dd8e847d3c9d86480d5312d0f01ebd0c17fa92ada8020fdb1dd02b5dd28df
zd0e222d1be505f49ffa0105b8969ae82aaaebbdfe267e420ef1def5acfd1d2332cb6dbd36fbf16
zf304fe67df64c37e2d9791cd4ac8da6a8ed8b1376ba5e1fd52c0038305504b17dd9d9ea54c6d7a
za34948ec7885f3961c77d0a51f1b718e051ccfc0e86d64c4f0f4e7e6b56ec3af94bf6b0580c249
zd9643199cae93e690a8dca93c77fcda1fc1d3b40d6a8122290f3600e070f127860658ced7613cc
z617f3303ffb2021689a87e01c826cdb1e49c0b3497f0dce61aa15938eb61da49ee4ed60577b843
z26efc1c2d9d513e3cc43de174714e3172e9ab464cbffa95f500f2ce06577f79c305aff5ecbedc8
ze4a657f80fa6ddf8ee24c1e4a5edc0f391574b554471461f904cb1cda6ebef8bc035e9148c7bca
z94653f32b3d8698fc93aaa9ca602b8a5b671b7dbdedd807152f5b26a63c3e1e6a809b18d633f6a
zec0c1dc3b7118e8b5be04e9506db363c3a5a7fb2761195f22ce90b1f552ab40eb4a22052f044a3
zfa9f9d57dab9cf0968df7a448c6e1028ee8d3a105b8d6f2ff6b1b3c33298c9b4b7e210a5784f85
z8a766d4e364d99e6588f8c3af442360af73351d6e737a335ff5b906695ac42b44c803daad170c7
zbb2f80e166a68d914223b44ae3efe25bcc504d05b999e61159feb489f508bdaffe000d56256756
z0b10b5e6a603a26f270f3445d8d848664a6ba382d63b84ac492f0810da239335929ce4891c428f
z19c751cbc16bbf526bd36c28af29700f8624b1a7db93a7c30d543bc74b0df379e28a58edf379c4
z52dbe679888dfe54b14edb126b2b20982957a15296d1f5e7cb6cd18f4ac91d615d2e81ae19557a
zef3ad0cf4c72e1c1dbdc68c6d06d9b2f6c81926ff980bd6e36c28f792b624f710d935f2907f605
z5f2269af0ebb92047540e0f5a15edbf75a727a34f21d4f6716e2b1e4950c6fc02508f1f4026581
z09d19ef354c1b50124559e90bc8b09aff34809613162531c95801054a2c9c22cdfcb0a8fa9b4b7
zaef5468940cd073f22d37b1f22a190a4113fb0316044fc4e2c3960ac177dd7a5f1ca1b27b20a4c
z984820f6e39e15efb4e3b842625719f25303abd98f4bb99084d521317a7a4d03467aadcdc490c4
z66f67e23e9985ca374f71ff33f3ef65412f23352f84a73cbda1c6b17c9c55fbc483e9d339e28e1
z2754b485563504310f8885a077fb8b93baf3fe223911d952d53adb07d3de7cd033df72cdc0219c
z10e9d985db4f4184c13fd1130a485f028e907182f08e3db28dce0f201042f64be4112a8e34efe2
z6897483d1a62b7c2128085f6567a4364f11780b1e48b404decd93c0b87581e38193597700a412d
z8e06b72461123fc785f746ebe4aa6b9cfe4b7f5b62d6046b06a0ac03174137d1dcbaef52a4f1ac
z5c1a4957455959d3f56e1e1f0d2da6d57cf80e5a204ed22b6e18fd5f864203f5d975d42ae66d3d
za6a6707bae2b467128ac707f2edef38019d1f034fa88a0b75447ab29c06476bd4ec757a0e51233
za29a1ff4c686b25f5ebbb79cc0cafe725e92cd1313f02fe752b45e485cebd2d122a9f56af793a7
z7e6d2adbdc3a3ffe35fc76f46302054d49f706fcbeb122b8133115d639141f0602c6ef8f894900
zbff7298a68a10bfab9311796b66f12c7714e9a322612c4f7a431445add5e721fc9a3295e5fa0f2
z1ccef0cbe63f7a70df1739bf8cd08e0d1bbd60be71addc844a3e13dc0274d5755147a08b7feaf3
z2799ca58a5a31a73f576e172ee29e4037d9a89eba5a63ef2fff659c85ac2632f7d9e9056697d96
z559e0552e97e18fb40161c927d72366bd4f7923d707f9d3a82880e444fbbac90d8bf7c386fa50f
z0bb208b9d741127bf91348b37ac651067e5df82ebab38644d08b6d3a2c1344df275f5b81233c8b
z5f2fa027fae55c88779d7e11abc37861ed3540733ef5a9a85a64c42a1e974e1908ae6ea34a738a
zd7ca9b400b4b3bd468b09ef394d2b92d2e69eef855502ee9a94050b4fab8eb7ebc6731e2211a8b
zc83223400c9c80d3c9b60b3dc0a0c2562821d9b612a0bf2a82041afd566bf4d454bca05b04755e
z24e7ca41bc1b571a58f183ebe11369c33aa7f482cb9f0e99f73be4f629bcc817804ecb05419a5c
z7808b5aa44abd5273e44598ac2edecc6c76abdd29e653f801f83a152df8f10c5b40684581f99e5
z3e9f794a68e3a4f6d2cf3df68eb62684c5f5bbc4d68e4cecf6a5b04389779c6fcc7bb61c08dab9
zb01e7b5c7a97d9fcb97d5462da2b51a2e1dbe2600234a81922046f481d1dad33ee8adf5bbab09b
zd5f42df22233dee3ae386c6d3978e686471292135a4a902481be3beaa1bab0d22e7af1faff537a
zf8e0a1e3cd9b2ef3b0a537066983980ccc47041dfd060fd63e642a4c0d607cd13c2941247186e9
z89b1ff8da681e07dbc107eea84637475671d1e72a14fc27ac7f08bcda04a0ee277d6180b6954ba
zc42af46caa736c780289116a04d5206e0c27a551d2767850a16a779647a53395e2495231851d00
zc4b8fa031231b9d3891f77bd5d39d8f3e1297b8e72df286ab48f96bd9573cb124655ad445ad015
z8bda46ef13ebebb5365d634f55f4ee09230ffa4d9ba8ce9d9f421e81e9e39a662f91a466541690
z550f3934c76a02e8c57336f0277ceac320ac9daf76087df7e910832498f45cdbf514b403a6a4bd
z35a324ebcbb0682eff459502b5606d9e3783bc12cca1f11e2c5546b343a0ec2dc50defa7c34297
zbef50cb1518df31e52d4be6a37a5e4f2f19c2d9b231af0a8af2bdf95ddc064a59ae28043cbfcf3
z8253dee78a9a01d412c723720e2c627d60b5e6e4a42ff4851c862a82746c93b24660931e5e13db
z2d9e39978d75ec4b69773a1e3b585c458c22390b23de6938ddc93385f2c387fae9965eb4e8787c
z45e62891cd39399ae83e3935d532939188d25ce8a36a1b8fecd9a008b6605f9ff369ab87bdd20f
zdb0390ec5fab9456c747962f436861280a2271c457ec9733975691703cfb68f46c1545a2824afc
zaa0b6be73258865dba61756010490d7561c61dde44826f849329097e0456ef46fc7b0b05be35b1
zcbb8f957ca98987ae17aa293f77607e599f457247808d3e1f86bf97868bca03ed92879b6d135cf
z39856a1fd0716a74da26aae3c1ed50ed8e54184ab144ba41c35642f34047cb2ea2bd521d6eb4a8
z8c9b44414afe9750e4f2e2395bce9111141897d3bde36a864e8dc9d82a5d375c28a4dff7b3152f
z0aba2910c5ab508f189cb8daf07d3ac5e327ae8453972cfdb528a9f8cb7123a5957dd3c2aa8973
za1b501ec139126234c0dfc0291bcc9a89d9a13cddee9e3f4e2501d69106fdac386e64a6323b607
z399f0efbbc3dd91943dd1d8f7824317cbafad9ba51123f726de9ddfc949e3da3b70c0cffa0c74b
z73f648221e62d2291bbc635d45de3d4d4943dc1bb1fbd285f566f72d7b38a0f0b3dc74e78ec1e0
z84f0fad544df5b20aac56a701203d03a2edde02bff4fbef9433b612467b3c7db9e8b779c06a3eb
z95ab1d6c59738cb47fed09ab189f77cf62763691046ba596b8d08b9560613fb58ef9ad5b5a0b82
z9e6f4280a3c2f9b6dc8f020064b354f48f327f2bc613450c67b4c9c8ea2eaa8596c4b01f14b6cb
z317df44c16009f2fa738421c3900c023a186419d81a5df98ec5827fac8f1703258d8d9301cfb42
z8a244df1bc7930a8e54b27579471164857925fbd1bfc76fe989c6f91c5c0edb0e1900ed04e752f
zb600c2cd838730503a84752704b90fdc8bd3a150380cd68f301e0486a7c4502fdb381bdc3e41ca
z5d473258e9a9de84e33946c5e7d78c11db13aa3f07b38891b2b7bc20ebadb8a5fd94cbf27357d3
z4dd935525b71252c2dfcb72110cb75d3efb34b3085d15dfbfa3a1daef88262d007ac92badedbf7
z94c3fd7485e3d1b3a610b590fe4aac3d548001253a93d55bca5348532e776a892567544ba6d1a3
z9aff013828b78dfcb104bfd4c5eecf15772f3ebacc11a21caf495ac5c9a1e36351f7d1c135eb30
z6d187a5f3252fdfad59027c644c5b98b0b61ee0506efbcd26d1f216e5fa6f50a3f0aa07489f5c9
zeb5fcb49767582401df6c8985eb2ca1ba4d31b9bddb1af0efd445c92100b9bbd48cd93fec43cba
z8c1584c66f1792a7818cbabf479acc27a237e929bacf48c06de12935b3ec3eeb3b0f39db5643c3
z3d1980c5674e0a0115c9a2439455bac4d8b6ea73bc8d8e52aa81d470c3d51dcd9a36a209d36ee1
za5ce867c6786ae0332393aa02e2c58a3f9d3cfa6b80c751812ef3c76fd7f543ba65e5997f99f6a
zb94174f0972d85046b86bc22db90ac82f8ab6d25364e60df0bb9f2a6807198924ccd957d679381
z56a03d7ee06e49b59c365eedbe4b9e1184c7796706545b7be5186b01541f9c540a2777a866ca1a
za35343f09887e93521de9379b152d32f71906f8da1d5d1e4ccb662aafb0f5c2d724f9950977ac2
zb37d8cba662925a7d69855aba21ca6ab9ab3b4474c07ac8d24dfc7fdc95b7b20173f94dd2cbe08
z019b4a7b27a86baf9bc5831e307ce0a87353d8f6c9467437b0e880424af584b1194e9b1eb7dbbb
z74d88fcaea62cef36515ab741102681319f81b653d28d98e942331ea135607efbf2b26f11b2a14
z487c4a67b36a4076a65f62e9df22c672e34a57b16a337d1509af097f44eb71e512237f2492dd9a
za12828d19865484049c4ae3205497c648c0c33506378e9fce63b7ee55fd3d5050820b67caba4b8
z69e7c404ae77ecac89d6778d45cf2313195e489794cbf4eafe5f49784266232c7424af5924b990
z0958b07c0df9128c1b7cacc4acd35dbbbe7a4bad54deae8f2ad43ff6c9cf1e33821305c8f5dc52
zf24391a78d80612cbc4980e60b57bc565dd27b5665277a70c59b696b4ae35054c0653c6f4a3fb3
z4e41a20e5576b15be23c74cb5ceeb20b948130a57c8aced17a71a5d5788a02c6930c31f6c9a6aa
z80b1e9641d5fa0a42e0f82f90d6cbb94eb9dac7c87f36c00615f62a9e840647837102e1dd02010
z6eb7051172bdaf37b71452f9aa57ad0b1c18212303092ed4746dadd34d180cb4db827f2a2effed
ze25da4ce281d5ff091d5bb796b1838285bd40781fa74f0e1c1ed0fe610a15132dad5a381bd5799
za12f8ac732f49a474f49e7d4d909c7b281c90069b7a1be8eefce54c4f88ea3d98f6a15b62ddd2d
z0cc17a13fa24f0cdcf0265fe803b61a3d0e7ff54969d12c079fd97628e919fc4cc1e274e4f97ea
z45ffde66249a9c0dc1ad4603e773e839b5484f7859c61697cd9e697c5483dc8af591693dafc14b
zd8f1ceb47764c85ac19645d90062a848a8b034c00a7e5f6b817f3ec4e7c553b4471a75c70fbc82
z00883868a265aea1bb644469f2b2229e0a297749f977eb8b7ea1f39c71e780f95caa7ddf161dae
z03741027282b4d7c4742bc0c3f551418d1285d6483425ebfeea4d72023cb3a00383ded04b603cb
zd6464a12cb18edc9dfa30210ae7a814fdfe0530c14f731a5c389cd12ce23932197185ae153e13c
z075bab902701f237df8da8b8f462eed33b6aba29bc36e1a4db7ce103981adab8fed68a70a2ef5d
zd2751c8842e4821932600bcf0926b5056fc5b125a70b69631a340b01c98e34f54cb1c1c37b8af1
zc88fc6271c35b4976e46916fb0d47c9f78960a2d629d77559eb1dc21ffac46d358e76028955bed
zb51e241e8ec51fe6d4d7a4c8d304f3debf1cea4dc96c7cd5b0f59e02aa019930935fa401ca0b2d
z99a8324c88c8cfd11c91bab6f022a4dafce6e2a0d2aaa4a515a032d86295e2bde90fa814365045
z6e9ed873ebf15e7b0e815c29ae684067f31b83062bb821af6d433465d39bb32fec26635ee1be8a
zb152155127a1141ba0a12af3995cd08ec89b81243daee89d12b7705f13dc8ae636096d7fa95b43
z72d5a1da67ce74087323b5ec2413a7c2a3a31d5cee1570bb16dc438ad52646b269af4a3a79f3e3
z96bb8653dba66813a48570c6e20cac640655d9f95bddf4c7ba073c6d3697f4f741c8056148b26f
z243908957b8c42f84b0e8e9c3351d22b7430f0df202b8f3ba7f142fabe62130c6ff4eb52e540e1
z22d1583371a97f035fea4015fdea561d9142ad5c2a8fd176ed941998787247265a2bdfd16a669c
zc8ac891d7c6c96454302e458812778fd103f795273b9a1a057727b2decc8ed7bd4b83b26ad18df
zaf644e020b80e931801f987505487c16082aef14bc48c3ed0066b45215b84100629bab5693ffe2
z4b64a385c8c060a6a77d1b9b9261625b4e7523682adf296be58482b15b3605264cb91c8101d87f
zd94cd845cf2c52c6f290e4a2d8c610d2bf226835f802bb3abeb0f6fa3d18bd10cb1bedefce18db
z3de1a7e9c181fa6e618b671855465d7e202c3a04ee25e77ce7d576e72580285fe8aaabd0bee503
za81fc4297f6fbabf927da63ad2622e2a54f5921f0dbc0b8a032176bddf42b94352973ad724c9b5
zbdced7d82afeb11daa91b77dc337acd33597f29211c7645a0fbcbb7f2e2cadb3c559bdec96c30d
z34e1bc4662f9d64acc1bbb3ee74f5547ed4c6b175549657f53d0d3c6c71f9ee35fc601c494b554
zc9054e8456230db7a22d49fcaa91016845051f4f20047b32d041679a0cfa6ca9df63a0ef67c091
ze0f94eca3908481f8b8cc3af8784eb1aa8b44e52e4515bc387526dfa796b70c8da605881bcc784
z15e03482f18d0b7809b86f164a50dcad4c1860d9c0c260461763b787c7ebb044071070904adc48
z8c514dc1c548ac99a503a5c8103920b53aff518ab964e10591e0936f8edcdb5b00b03d909d98f9
z4631afb36fc65725b611d6e547ed21ab30518aefd3634f4c46de81ad6138eb2768eb650e59a4eb
z9a63540e4252a15f4786cd3e344f32b8d96c57c04179d172bf1a038869f111082ce1ff49e2d5fd
zbefa13270d9feafb8aaa378e1d87219f52e754fb3f188b98e7c19dfde94ed3a20ca6e6933a89af
z92fc42fddb37ce3c293e18f9626874bf8be9c1f10fc353f8e31e6ce1e966db4b6cb5e64fd3f1d0
z999cab69d2fffaaea2701b8b225e4a303c2a3d16cbe456f818dee877f4d5bc69243ca2e7cbb0eb
z5588835803ec93af9025f5c3c816828145dc0168b35031d110812ccf8012b3be797e9e33e7ac9c
z4fa681b35f46a7be22ca676288c901c0399a8d21545d69803cec200da2dd6cc14084830bc4f460
zaf39c8f7e62145b589cf4b6b0076bbcff094084b7cfe12fd5965537c0fb14b97efcce7918dbe13
z1db852ab14ac425546f54a9c01efda1a47da08186476cbb86c4be8291e4e94a8c001e81de5b5ed
z74099616b9a39cc43006e1060ed25f70c4ad7072867d4f9a950ad25cd2dcbcb1d1aa03d1eb57e2
zb1870dab2d68214830ae3eacf328cacc9ef9d3dc6c59ffe599464b24e2fa35b7561d6844ed9253
zb177101e30daca2071a3f24e3b01864d606679d9563291fef6cd809ea9010da08ba04f202f14ad
zf975b0e8e551777ff1671a5654ca54cae437a752f8104213bb2e4c3a4aa41836d3133d465ecfeb
z597120c462fb6681212e4bf24e62c2dc3667c142dcfd72c1c6ef4f56346ea24f06eb0f62bfb11e
z67d177c823a85b7ecbc9f43ead38818099aa996053ec8303800750cf0f2c34e75eb8edd79a8251
z940de8294236b97d9d5f96a3b4c473cf9284c95d0029e40953596b7b3c55a4b42f74faea5ed28c
z7c8c5bb67d28594c43df3bdfc1e4499f4c4ae6ddb046c71c9eddcc531a294540a32388e4aef6b8
zd52d168b1fa81b7400206ee2afda4ebfc53af5caee7469d2dd502ab45334c4d8d40364447ee7d8
zb87ff75740fec4b5a2b7e2e2b0f22e677d8f9979808ae066c31ff3aa59a34fdeac7ea16d4550f9
z3b6bc0e5fb197c1a16c368b56a82cd36f671191bf256ff54d080315ec10b8fec72b2f442a3f425
z46c96e0db06eb9de86462beac5b34dc1fe97cff04ef67c5b93f12707ce62b1b7f49f8692e6d2e7
zfb75bdb8e403981f6364afea2274c6a18e13271d93815f3f47006ce9bf312aa43c9421ba785cb9
z980b1127fc7c05905c54368cadbe3fcaec76b3852e170e8ac428b9badb66634f0b2a5e9595d52b
z29319516c795338e04f72c6880095f66a53967c8dc379a0388f5050ed5c74391dbe40918721e8a
zb501745f30665dc82cf588e6ec77192bb3ed91b2954e1584bf8d5e20b5e2db604d2a2cb6c27a20
z3fba36480307219c117eb7669f91c30884fee037846877a849b5108258afeee35530dd89d14a69
zc6d18a6cbd69354f503d0263e4b6e2f61c006986230bb41e37b9e356fca09dd130beaea66c0689
ze79a213edaf070a45e905ca3baeec8ae4a7087e069702ee349b10a805abfe9b82a7245e690a862
z574721b684133d031549dc53e51e10892e8690f291646f61b871b0bb7d170430a012d918b3d79d
zcb92cfb4d4c2d705859654ecfac5425f3a1b9ea63e1139df4317ed94e70ef0b7b98219ac49615d
z1c5ac39d58e36421373cc499f30c6c34ddee91f5a9967eb733e83be0e129529c4c98ad2029fcdf
z5cea562a60df3dda8dc65fcc93cc752e7870c6995b7b3da0302cd4bebfcb579ed599be26fe6877
za700f59aff350f7c5f013cc516893f0f26ecca5277db9cf1a3297cb9da14cd019e2217b01d13c5
z1faa4479c4c39ec09b694824414930612da30940246046d10ca400bc73d2cd53cd69994ff80b47
zfd057752f4992eb6f2ae1ec88f4165b160f1b6390292d00583416ed5c7fc7e633eceb9280366e1
zc41d1d45110af29e793d3b7607f2564c633dc3a2edad86169875ace19a5b1d5381481f76971a6c
zabf56bccc57933dd502ad0356d6ca1ca8f8b13e6fc3e1376140b4732550297819b1259d2bc77cf
z4ef9158f6d47bd6bf94c9e373bbaccf04993dd076a02f65236f1e444de767b19e4562513016c09
z9885f5d2235e0fa673ffc8b19067bab6df8da28b71cde51ba4e13f3922f3a2da9691f10820b576
za79c1a8c38e4fe750f06b6d3eef02c06f324c878bb68a6a1d340483897c572d4207bcb8d7952cd
zf140d4076b70b48e28d3bf632985a93dee3dc12a25e5ec765fad57b415f736f21c036d650dd8ed
ze1a8255f20c1ea4874110c018982951ed0cc4dfd79d5001bd90d9ea8baa54ed58d3844b1b3321a
zc75b3ff90c80c89ed23729402433b86b3496acd2eeb924b3aa678c17bf8bf4908ae11a6c8bdf8a
z00e937fd401e689d9421690c63037c5f228bd81799929b9d0f8a1098d0b5cca544c3f8f00d9b9e
z779e33d691e09a00b2693b1ed6ebee6fc1c359ba0400db070f598a5c588f640585ce187c4b5ff2
z8379ca2b2ce8046f84206069eecedc24cce5b7af8a37ffaad3f25634557cfb5db2d34a402e4972
zfd328b820a7c957239ff1d331647c5dbf6b2d7a908c305bec44c312bb32f5dcd266ee5ad474113
zb0581412baaac33d122f01f1fe0c2d67194a66f8a0a5e8abeaae52752acf130c42324902770f0b
z6b24600efe625a1d9ab235c26f40101a56204aa461b2395d80cd289b71407ba03ee15da60bc0f4
zc3b19ee9c7493323aece2fd50e7d6c511c220a64172efa21bdaa36299fac81097dd29a909f0802
zf3795221aa3c5414d61ccb914bfcff21b5755a99d6707d41e4fcdb9771615de356a890e999e744
zbd6f2cfd14ef3754edd2bbcd794b58a4231fcfc79fac30e56f0bbc744f117fcdb2bc038831b039
z92be9511bb5220229088341f23f122549adc851d7e2bf7b946f342d2d0f5ad7043a4cd19e730ed
z22aa38236813816efa80ccd087d735b4c5496b12e2f4b23e5ba08261caa7dadea0e09698010c1d
zd30686c110d120d4d52a5f2da9a6f218539e1bfa47151a48db08f4dbe7266e43388f350090d92c
z8f71df9e7dc3b06a7d2a703c956e03e8a5fafeef8a12eba21b9bb503f3855e10e99775109cc8b1
z25165a80ed9ab6aae70b6a7522b00425f3acebc9cfc6774c383666b7ca5d5485c65743d89f1d8e
z2914215f994216ea1a253ab79c51a530ebd99242dc6c3070992aa9467c5db5f9566b68ab690fee
z6f9fc13fcf424b5d31cbaebd06ba8659e303b2e937ea2848dc8f7863c803be4522b639a834431d
z249e23f3e255f9275914729421d321bab4bb8305fc82178d3be3acee54cb8fdd6bd0346cd925d1
z2075106a4cc764cdb9d6911423d304d179be210a3d09479a7148e9d2255eb0795668777c8da05b
z2b4e38630f0d05d4189160aa3b5b16fa21d518cad26303fd845a03ce8a6ba420eeb557343f866f
zebbfea4206d8e7ffb6570100f37da393f7388dfb6515e9a16c6850884cdbbd9951e51928a8eb16
ze3ee601559a0e8aed4664de8ee279106c08c8d855c77c2a39e2bf0668fcc012880a3184d5f5bbe
zb3ce76615d15a2d3e70f318a1aa0700dc88bab19aa186548038ad714aeb1c6a2927b7987dce8b0
z1995a80a887a6c85893e311e548820550732d6e52737b3c68cbb77b2281fcb863891a6cdea5e95
zde78f5a43e40e7656e2a3c98d79ce29ed14cc82387c08473c149b58a3ba54ec66b1e2eba482daf
zc7ac1e527a058b2108a1487c946b77188f5f192e8ab54643d0fda653cea97a4b0a2fff179b2b4d
za5a52dc15fcc3e0cd5676eaa9efeab9811a4e4c056a383cc1ca22c1c03a9e0bd684569f482aa0f
zd0ae07554e803e856508099e3b741cfa7056f09de14ae1d87ad6b30ed3816997e12510cf563546
z145f5850542784b50584065e2f87376718632c3f100957b29296b9a48773dd14d49c9a44847579
z5132471b0619644247a570d45b53f0595cf32b1cca4d26f7ec5a3875210dee559d30b43347e610
zfb569d329a1a435e136d8471934f57dbebbabec06f31fde674de25524b1fc1d7c0ff01c775614f
ze85fdccd5ad284d93d31e75120ed24749d3d16c2500ef35b89501004250de2eb1ce09c1b555b4f
z4489c86517d7ba71dcd2073ef775b00e003d67c67165d78d39cc0dd463ac5c0c70b3b1d9cbc697
zc4360863d8ae5e184cd6ee84a89dd329d320a426ed699b77027cfdc2baf5987e15e8f2c4c37b50
z0f5283dd5d91bcc938f8a35c377e119a2a9535ff1105b752ea2d28bd1e73c8cfd4250c393d6c45
z09320613b96899ee50647175a7147d2130ca52148dbbdec4e8bd47ccaf1500ad3d588fa0591aef
za3287e5828e3c4ef06b5979f8e31c2e55071ba738cf797aef8e7b9eea29c74803df6b13d8ccb7d
zc55d941d21fba12b9f1f27a9f878f2ae31758c32fc325bbf06a51422cba4138aa61091cb0fa0cd
z10e94de156db55615a6ed4cbab3c6e24b1266a398fa8f8eab7bf450114ff7e4da1d0892e3d4197
z97d0eaf62a5e5f422027caa42cde32335f453a3a392fb0a5a7a223a5a19315f84f44f6f80daa83
zf6e344d368d85fa10425566188743549d8a0b4d0a915d9c44801b6a479561124d3f357109891ea
z70eefda87bd95935c28fa20e08b68c740c2c364cf0048e5b21c5f9a4606b4c734360772b9a3384
z7a429ad3f25f45df832770e33666354c7d6c5d63f01c643519a2e7d90b90a0225d010b6d780940
z47899b65f6214729b124e46c3e3cc67aa95946de801bc8602eb3f915e4250ce43ab458cc699ba1
z445b31aa3bea2fbdaf9e3080bb87fb880b3eddb665a736f9715c29bfff6b54513176d1da50941a
zd654b79609970664d7f51db5d1f4f636f479b5f1342d236ad143034647dfc66ce08a6b110f7fa9
z25b8e0302de9674211dd718a478b4abb7e104385e27b43bf7b00d564191dc1503974a6d15c7209
z86f15530ffb114ecf35738c667589d7ba2281c9a6cd23c83191715032150123425309c9f818760
z4eacb50bf375350fe5ee05ffe4c8e06bd523270c39408c8261d0407eb5277cb45dd968800496c3
zd91d3062680add1587fb05a669c643ffc651fdee28b25a992a73ed94ccc936b4bfabb12e87a426
z788f85e4cc8d1f658ab120be8b7c97eb971597dda7238049ecec5d2efab58a2f191a9417f1c5ba
zb0f759ebaf7387d07ccf62beaf4d712dedbf33f40c52f77b70ae1aef3d88b69086ab7395b9f840
zbc9fba4cb935d06efd56c17c3cfaf5ec0d73a98661d3b8db9a412def875c167c9558532f7a52e2
zbaea76257969316d3e41bf3e446c89cc0f56f8aa125cbdd256f511befaca94ed078f8d7bb6bcd9
z33b8df36234da1393acd809f88b28a559991a85aaacf7458315d9049a68884a669726fc9b11303
zc15a00920e96049075bcf54304c1bfb418e9c7fed385e1d28092db86679ec18cc2d449592a1a10
z9d75413d246de60b271af21f498b96a0d0854010b8f9f835c57eaec056ae6889a253261520ed61
z28fea97c094918599556fe1ee62449d8424fdc3112c7abf80f3e17758d8287ac764413bd25f66a
zd9fefe5a132468db5f7f67791384c485e8f59062a9dadba29af333b05bd4f85d851aec4ac9e380
z07cf46bea28a7b99afe2455f3f9d13976204911d73ec00965a2dea40d813c6d62ecdc20ac1e481
zef8f0e9b944171b2678a44b076246aeb5807e7e691d5b4eb57aa51adfd87081379a8673d1fb48b
z1c25afc746c1a60232dfde0bff4845b041f522c1da0a6aa55a5d4f06d40a9bdd2db1f4c2af61a5
z191084f4c3ff4ab9a10f9361a5f97972aa5be63423f9fb35bffb44761fdf5618a958c8a9349eac
zdd7d6860ef8dc172ea5933ded86fa57029712135eb3a3b1c39a1d32a1c3d7901a8a82fe693ca82
z06a7576b39a7f7fc1718f050322f6677521fa5a1c0a7c95970481c291c783b7d2cc2a8168046d3
z067ac42e03b06a0134ecb8d8ea198e58b203d596b0cb610a18ccfa92da4e37f68452ca5ca5247d
z96c6f0e57b08ae227b2c93be38a282d13a265efe398503a4526aa57c885bbf006a3e0b8984ad8e
z2e65f14f8d05fe719b2db5461d85c740bd322b2eed3316eb79b48547cdbb3b35141aaf701f2bb4
z111887d482752ea6024701ee4266f4cbbdda7f73c7386d6017758581f21257009e61dd24e17f2c
zb291cdca37a05e8217d4a2acd28fd02bace7aad4e0e9b346b394d8e3b4dfe6611fe03c8c0b1973
z4de2548b315418a930225d2a65e51a9ec4b71deae664163161fb7baa7f7498d6a566f6d84f1cb2
zb19ce168c24896b354119032a3e0f9c0b3c0cbd781a9632ac7c540a0b12a711acb7bf92e607fbe
z30b001e57ec43adbd3a7ef1ae266d17942fa5d056cd96fe58ba60758f7c26dac1ae1fe8d890ab0
z985cda1ce308f158e4fc7022a1cf2f6a89a1a500e1475e832d6bea5f477db3b42dba1d11e252b2
z8cd9b0411ec0c61360c52b89f709453dc40808e2f8cb7781af59f1353cec8c5849fd7155e13c7a
zeecc94690628b099fca5e265c897437ac75ec269e934b0ef492f45bf66b14f330c10b30a37c54d
z05f346e342adc75f221489129d8d8649ed7763dd3aa65d91413b8147ff1dae22c7c150b8af6bda
z14e47665b81e74279e0844e466f36f7b53f764bf06b1e1174845bbcff9e09ac98311b21e5c9163
z79be83c05772149c3a787b885cad78bb2055302225b8655f41ce29fda0aeafb76355a9d30cbbfb
ze721ec4a7357b9a8aa0d0d26b0ea4872782a21f433303e6c2fe05b2c87cdf68fab1755a9ac150a
z36cfd38b89d2750fd2098ca7c5e0476d485b146bf486617db62843faf3a55ad9c7d3402422614f
zf902e2218a4e160ab38c5ff2aa029efb8c255c814f4f690f8fc202a484468976020ef35d8bb53d
zf7082c761d37d478a9d3c00efa9fbf0641d4135e9b47b40131761c199510a8724b2aae4f8f008b
z666b286f1ef9fb7a27bb15f9df8dabd1a51b798a238f9d74ee5e5ba14dec9c25c14719bb6e4a5e
z82ddf2bcf3bff6b437f6b8e9a5fb586eb0ce040292d600c0344761434274c35c9884367dd5a948
zfaf3bd78bee2a045d37024457a239a0fbce89d94c6ac90b4eea8859396350814f77121da674d39
zd9da66a1a29d314d03c76a1c3f62fc59db340e0359ee56af54a2b0c434e00e29f7ada7a7edc4e6
z757ccb6f9c9ada65ccfdaa4e56b910d156274f5a77612f491fcc1403894bae838cc8040c34ea8d
zcb3d0d475d4a8e372a2807b9269d2ab98f93fef16a608279c2ad51f31dea01875ba6fb2f269564
zc3bc8730b7d93bf537f3ebab6c6c81a0167946f6909909617637becc6e245fcb98651f217f7797
ze3cd2db3ad7af842bdc48975509125b1a5d68d39900748010fe8dc29347f44dc528d50fed1ce07
z46e17036f1c3e34a81749c046fb28f7c762be3204e00219d738a2c72c9e9e9b80ac2060c34e165
zbad9710a67e1c7e399a5e3ca1b80f0a4a6f93cb83e0772c44550749dbf723e1f671dfc03b4d44a
z61d96095624a29ab6b35c788b6ea44ee8697235e02d89d44e888032a0150a137f9bb9fe609e6d2
z271a96df1afe225d290943bb1ed32b918c40fee8237a07c14a6fec5a2da09bec2ac495782220e1
z0b59ad32a6f1e4ca87999d7e37a5205e74bc9d32b14899f15a5874c6fd96406f827daef362ccd0
z15476b13305eed4275ce41b41c444ed79a4ea6c03c2c40565dedd1426f64e2c79923d4852c0274
z4aa95a62bf1ac73829de8b6c248bf216d417a899cb3cfe780db579962d9221d0660e798e9491c5
z3231ff5c8ccbf794492d7e2aa586c81b942c1fb4e02343379c3f6b36a2e2c43ecccd2c1353dc1d
zf17163bd4c3069f197d83b21373039aff2d3ec8b8378e058a4ad6f08244ce01485d6600e428489
z0715be511017c63e18551dc0426daaae20df03463b137129fb1825e95dc3d4be50426dccad9e64
ze6ab27645f243846d25e05a429aa07fa7480689bab103eaefd49339b2efd66e5126ae15edb8aec
z89117474751d126f8b2afe83229e0b158cf1f917bd159c87d35e9c2e6914d4f6b30040be1d21af
za6127f1714d47f65641077fda39b5f4bb20429f1ebebe8fa76b01e14911f609e6ddca1df74599c
z600afc4147d91f613d9feccb07476590e1600a59cc5e8ee89c0fda263a1ad2969269f6e3fa2b26
z004125b3c9541e1fc31b3698292dfbee56507e4159af0581609d1c20b01195e7203ae708060766
zf1074c0c2e87cbe799f854255f3f2675629a4cbd53439d74a37e7f338a295985e6764b39cc4a1b
z9bec90b2e1bf12b0fec3d3825ff580ae36a62edada4461d94b2c2916ac6cd70cfb06167a481a9f
z73bd86d919aee11992513e2f7691433aa3dd8d7e9f3d3ce4a8104c1098eaf8a2611851675471d9
z689bfd44d6e12d77e30cc1f812261512cd9d82cc42e7e6f25dba9f882c50854b6446109edc7762
za3798ba56a95af9f32012c621c5cd8b2d5ad84647c3601e82ea4bdf4ae3fd41084a65407dbe865
za1a3c3f8a58ab034b9e41fd3cc1ff57459efdac9b32fdf70d1449f00eb68f4b83efcb8812e0466
z88b7a55ddd3bec8b583a62f0ef9a5e40ccf79d997a7ddce740cc6dad26b008dee0f0f56f9cb8d0
ze96e250379ccabcad3efbf5e5afd1ba881cd600ff623c7e825f6e45a7d492d525d067c2c330100
z4cd9783b692d2c2b2f80aae26605e425983cad7ce7e744dfcb2a025c2e41212f9d3fa679c04aec
z0a250eb1999ce740b9c4a5c18a6a3bf0e2b14d4f49055397900642525eb5d9b3d93d6acc0bad98
z6038b675850a1e5ec7300bcf96578a81625b36a06536058e49c167b204d6d03a8caeddbc7e3d03
z7604c007ad3dd1f5c7ea580f945e01bcaf059265a87cc3f648e331b8441b3d91cb37a663a23112
z9302829a706102ad9d286a99e93ed5919834615bb8cb2757220e83cf10772f07b43f3b74929448
z847d4d5a2912569544348e89f2b73b24837371ea1c5d4d3ea0faef352a42813e3697195cc80b1b
z333a31ceff973b9b1c9e964838c01cf84dffcf73e9dc3ccda1cf5e17440a92d69a5f3b25bb47f6
z374d5a853403880aeef0203711eedf4c904fb61f89d45767514d40aa7efc5c3369bdc07340ad4a
z09dc7a357e97b1c620bee6cde8481313d070017a37a13c8fd809152ea11beb33da8acff4e18445
zc5a33a6af871db21bcfa8d51ca6f0db35718dd009badc31163fba19b28bb291dc36d3702b52fcb
z83e7f83052dcbada850d6f66fa9cc74917a1cced8b5300ec2c8e4d4a9649446e2bfc08b56415a4
zd3f6e04aa981b88b2f9caae075d65822d4c60f79f0237270adea2dda1e712acfc7bc635c5fda72
zb52a22a9baef3101dd57bcdd7ca0c5a390fc6051ff4f7589d474d3f13fcabbb237ec724ce62cdc
z7980f44f61497906725d083e77c1e8a2febd75a9666be52c808d151c85516c9c9144a4b74bbc7e
z43f82f0b109810a2b6218dcf577b44be66c654ebf56c3a544435f50a7a0dc8077acc0fb156972c
z419616111a2ea068402fa6bd380c3e98812dbfa2ec37b3581a99ea423b93d9e610bc5d975a1609
z78afc0c3df5c7cf686e7cff82c650d7486d7383f3f1403f81d340a3876f38752b5563c11123e1d
z8e528bd27f1ab6211f1bd0600118806bfed6a5c73d41aacf342ec7fc08230cca277cb49e4932c3
z2878ad3bf174c8e025184402967104078a73bed224de65b39e1748d76ebb5a3309958621a4808c
ze8efc1463173605aacb52341a9ab37891949d43915dbc29e9da60d74bb9a2e406e8220079a4126
z5de12c9b885655a727b82f70578b6e83533f5a91deec6d179da023f4e88e86f5a0cfa31c36d515
zc502b154ffd4213c50a06368127dc90043fd4b25cb8016ac66f83310237c9140c73bf020533d6e
za5fc06ed19437609198d302c68d3c2c385999c34d8f0624651ca97569c0da303a4bf8385902084
zc3bd384559adf95be784444d81c104b410a85fbe450256c422dbeede250ad20de4599f22f1ffad
zd07bec79bb2715de35c6ac7191d048d0f6069b544d7915ced74b7aecbdaa0040506040c9de052b
zd7e1b412ac8a1ceb2168bf595e05e6f1b2ebdfde89b93ec5aeff0620f92804ca70fc7ebfb3f654
z7874d810810e6bca62476eb78092a67865bdeaa51b210386af8b83a5191d80e9a8a67cf06b91e9
zbe71486b2cd4845b391030196fde89f8c34c2839ec455260be2bbc64fe04c2140ac5cd16fca772
z29a1af01bd81c6b248aabe096a3a86ec877a410fc83404a545eeb9cc3fe84fda75fec9368ae803
z08519d9120dec4ca027ff45e2d789a504adf0cc3b68f7b18cef272676f6d0b9369bc94b3995029
z529702dab4731a4421c25f0d29f6454e6f523c231db978d55a9e39689ca5d42e3a1575cb1ff55e
zd3165777c977d3291f3613eb2a75d3324e56cb306ae4560e9eeb4f06d64e92fd8681d6ca097b13
z297268c4893faa896a76dd45366cdc74732776cb5542f589dbeeda8abb1692e34599fafe44bee3
z0e3bae7c3c0033c12501355c8551993dc93a9fe212e48f1328eaf64cb9089ed428bbb3cb8e698c
z5a02f7436c9ea8b0caada37d18e9c7d6612ff3804be8a8519e8cbbaf3adb735727431e8228c510
zbfcb51f4939ebce695295c82c7c2618611e068cf92c35c3e719267384c78f451892ea5be2504fc
z284197d613b0eab3a3e9bfb5e510b17cd36e0285b4968ae6fd02f3bc617aa23ef320b26e4765ce
z5bddb9c7695b256db63ae9874c35e7e98c13ba05db4c4e78be1242220160e6bfbb8b5261f57296
zce92212d2f1f02f75e5ce5a24851b143f9a7ef96719b3f8c174faffe5083900b30e2efb8c6ab49
z456e6b6c01cbee4e81efa597a9f5214e2db118ca2bf8d11f041d6e0e6db457cf2a9207efcb1a50
zf7c9856af7cf1de2072c581db811a67e36a1c1f3ad93b188279ac311c304a9e49e5f774e3bcc98
z8f1e8ee68ba97962743081f703771f1d258b3666c6384c2f1f50eb960523be859fbfdcbdd21d39
zb946c6a429544475dced74c065c8f0c45161810cc53dc222d2f944d16767a8f4921404379ebcb8
z62a127b24d10b91e1e319189ad9fc31422ef7fd5595551eb5f8df4ec29f0ad1fbc2f31421e30a9
z79189d5cb9ba384b37b37fb27a37f0956b4844a09bcc622f6d6c5283d965d05827e5feaee7e950
z45d11b98ed927b5515b45a6034345c0a079e60c71e3e761f01d41c71ad80b2c953be3ecb947182
z0923a038ab911ebb2555844307573e9945095340f390c1ceb83d6c327c232a4f4fec3dbce7773f
z498004da75c2acec6d7bd38d8f6646a6793d386171407697c8e30f62830452837680a6abb6dd6e
z784b25cc5e99209029bb90e2e05f1277164818fd7ccafc7ae6b1e9e3b8f6b751ab92a6d74c68f5
z102b26c550d433ae15d5031639c44c5549f63b70b1f7e803468922318e144758c54cacabd2e7de
z7033980dfe5e8133d5e421bf6c327ea3e8771e53d34f6e0e46c59a64afd906517a1ba508828678
zdf8c86fc7e958659d2aa2a1372b5802adec23440c1f797bde2cbcd5640841ca0a6bf52cd1ca089
zdfcc3e8585e3ff1e980ba10746a7389e925d101604af4222c24e62af93ab413274dc3865cf7671
z5c4627c10706612af418667297ebd7652ff9364dae1f064930cf5df6086bc533c867b776260973
z200c7b5c3593e69bc163d6f4b3473ca4c381d503f8f6c4f87d05c59faa7cd661e253b967b303ca
zbdcfd86df94ab05a12ac398d74180b9f520fe9856b84ffd7182697628f1979c2e7901163291a4a
zd223cf13a281a52677d9b84491ad60d1883d8380835a760145a6ef20205edac40e6fb9afaa69fe
z564a0309b06a57e930b5e54083377aa0a9aec54e04fe142b261d7833f837c1d5d6f386ad012ba7
z29bebfc98177398f85576ff873e8b2c0efd4f3705f3a4565ae189d9544a43ee97aaefef272f1dc
zfedace950a40840317b0e71382b9b32fc3c1e1af498b81d8995609499743d66ce37406cc443c21
z0cd5d8adb2bc344f32779004297627bd9d0298dc378dc7e020edb494dbdbc76d6a299ef9be8a1f
ze32b0f85c6929ac44792119dd388d407d071975a890c2edbe680dd10ba5f5e602a45b6ceb6b4d3
zfd676255a3a219f24225feb231e070866cb65a7e5b93adefc54403aff218be00f6b0c6dcb88e5c
z4da55cf07cc5d68e6daf525b2d22fde5c7772d37218b58c52d254f640958f8a3078c56fc08fee2
z94859103b5ab9f77fa1d01d02b070a82eb2a427f79cd666b6066929764188bf749610f9c584d80
z45d3e6dcd1d3ae2cca499718cfa3532d934b28a74ee8148948dcf9f4250bd70017924680a88c6d
z37ac7cda47110b4fe9c5eb605968bb0a1739bcede1025d6eb3de067b9687d0e92c6efa312f2048
zb5a606847729aa3dace30737edc4312f6a087b52eeed3b179b93ecb731b84581283a8529c717e7
z953a206f6b5d626f53996030daa0c3ee1c39f8496082f1f2ade8fd2cf79e1f8a27b46385d255d4
z69137fd4ad44d87629016acbbf01f4ec973fbfcf14a3ece14f77dd90275ba597feae956460e12f
zedf171c54bbf356555cfb7ecae04355353f87aeca50e5e2e78f21b5fa25bcd8702ce74fc42e01e
z6cddbc8539e8084807dfb3cdb333756bf90a7ea297e8034f4b2d867985a8dc98ecf4bef871adb6
zab40966aaddf442f43a43431aa38dd64309e372ec1fecbeb1fc47227cba545ee9d2ade8fb351d3
z6fc2c5430446b32518a1255894d9f7436efd96111e3a7a502de0745146837f22da80a1e91bfb8d
z67c1a11e60068e39b2badd7f33e342ea19b29eada02a36fc165d57bdf128b5a0f20df05d30d07c
z029138c4df24fc70f5a968e74c68b88e4f7f1c398a8f6c9deeddf64cb9d45b25bc38054e53b270
z10f7d2237e26f17221e05215807dbc31b5b27a72260f70c8633e0b4fcbce0d18b6bbfc3c82eb68
z9b743702c62b728d1c11db303221d7d3f316816a576e97d4f3992fafb7a8d7fb7fbfff1c46610e
zb2834b35a68887c917783b6b2d4b32b1ba0d9908d8b542dcbb0f87118ced60dedce8cb2f122648
z4881f53601fc75c5f5ce532b5ff57347751bef3c8f21a8dbcfeb1dfcbd7d2d07b1f6b4728eda6d
z3a3e5beb153798bdc582be050ced039f87930191fc7462c663faec3c0f7f454d1b9b13ec92b608
zbb9be9dedfbfbfd564d1c543480aa30c29c3263648d3ca96c33ae2d8a2b1f4d8454377b51631c6
zd7340bb69d7f1d79a2bd56482469b9b61974530a18fdee0f31e134071858270b083945837fec48
zbeaa55b8ed4e08ac89a8664d3927dc5ee74df035b17a925b17af56cbd7bee809dc78c7b2a9901b
z105d96e3e587fc1b26eb0bea74140f56c4264119d951a977048245988a052e0d2830fac88a1e25
zec66fc317a8c6f4d2b3aeeef1e59d4e03f4ba9b9612f7f3b4ee9554ebe08141832071becf49b94
zf725548c9a4be42e3ec810b3b1af144468a86c586382b42a8b3115b91d5344adacfa0f1faef01a
z16d28b75546a5cdac6ce957050a70dc388f88ad1962a9c755e075961df31870f53072bc0df047f
z16517fb12213fa2a3d3dac9ef4d4e7bd4dcbe7fa16ff678edc48994e148a3709dd1c168903c121
z4cd3926fa16fe19a8162fe5815939e97849717525f3e2cebe02ff105fdbbc322c8076d51c21e40
za606af8ddc1dc52d195adc7370b90566c3169c2bd4aea13f401919b4802e24a9fb9b3c6c0cdf36
zb9ce0d230105eebd2c568c798935ba130e635a075012093b8460f63f0fff7e21b51124aaf84fcf
zc52d5606f2db87e5708e9b35afaecede8fcf845c5d5aae258342b5650e893ac3388da7b7473201
z69554cdc607a0300e9672ce062ee66268371c56969b7e795fd7acc5c9c622ff959ec94d9ba06f8
z360349b534c63ecda0839b81791cc5afdda026c34b62514e3a113ebbf370b9a583eff97d96c471
z26824c57724144a76ec29e656d50058e9300e7d479034dcae13970273cb18cf41642fcd4fa9a06
zbaa267038d44f28242d30795394aa6f59537eb763c54ebce4745d440ab7211f66affc7eecb1e17
zaeb8dd024cfe14e56c8504c2fc8a152064693a8abc81addf375b93c9cfeb1d73a5f04d293698f5
z16a443e47550e80a53a6a3263294152c1bd9f451966331575568f3b73cf13bdc84300e220126cf
z85935123da50f2702eec44d70c07a04e28b0c549b263b0d83530258d8a2d687d8c30f48bb5e7d8
zabb4bf4f996cdfbcb50e423a434084aae88e322befab8fa63145c0a2b1261ac04d39694f14ff32
zb4cf9852c5408b22922c04e76d7d97d42d807df5326b3e4d7ef5acf73ed2958ea9e94ae15e09aa
zeaa6d52a146cc2bbab0272aa4be32b4696c5ad037749fcd35375ef2c12da2b4331305f3f6ad7b6
zeefdbc13f4612f5a4db23f91788b11424d7d0a84a51c458ff6f4b424afefafff0b1669117e9406
zbed8aeef3f3be0f395b0bf601ca14c20ee1f1c4a6436c3f40927b2eda16921f1fd70d1210897c0
ze6e616e9c3648a54616acd91c51969a592a734d40671640230b4eee036c45e5eda3de5869e3d31
zc929389c5bec663db34c46b27faa0d8e2c89a54a553543847df392ee3f54805def8651fbf42433
zda2bd59c930c4a1b50cf51c8f1c72f34cb6c90ed5159adb433e9bca7df3885ce8baf21bb2b08c7
z381d292118badcc8dd6068ffdb7c1bacdbaeecd51b916b57959143846beecaf51786f6ac9e5661
zd6e72d85e65b99be683ae91d8b1f004ffbb8f34fb9a2a047ae6006f3e96a45d9d0dcf8b811e65f
z789841f0b22e3c21f7e27d83d26e4db5085f5b30e7ff792b6db182e3f8ac957c88a395c5957fb4
zea39fd1432fd361b7edf045b0d0d266c6c3fe4d7e2d581573e3d96de2bb391c965e0ed42ac1e24
z1288622f631bf42c143c3cf81224eb78056b02ffb3810f147f254ac874324b6f3dc34daf8639b5
z2354870d2d41ea7e1db92f3ea88b66fe3b00aaa327eaadd23784326460038108cbd02ec1eb0629
z4adf34223cb27ca079aba7510c46a3c4a92a456bcf273f3db5fb864259da0b532de71b9dce459c
z1ccfaaa82970bd28190c8f5d93493f7a2649059c013b1d56a4b873333d3c4de8f54fc2e5b42d77
z0854589bea087f2b16cc28b80aad4f3f16440a5ad5fa24d18611f1b1f219adaa2866616d1930bf
zee3830aad339dff0143ebc5f19d291fa5e30ab090b22ef31c7d449fb9ef14f015b76556b1529c4
z94a0d1f78de116c672ab57836a5469e8f5d96988cf3216f186ec94d320a27fd1b69a3dddd262b8
zad1b5f800d498560dc8cf04145beebf5b971ee9d18ee7c5b3e96c91a47cc5aac164c929add3072
z4883cd240b48bfe1eeb6afbeb28538c9dd700b1f80e22599c0324c49b30ef8c5ed2fa42300d957
za393eb1a8f79cac83d25beb5e721fba4bff17f3bf759b3455dbb90bd1ecf5366177e1434c3677e
za4e1b4aa7468b677ded438a8d5f488b1848363e0cf184a438cba99a74d27e98b04b2af9ee19c41
z9eec9141c4392f1e454bd353d36e8545f86ee82663dc92382da664ac04714838c9b76cf8904062
z61def6fc4b5199fbc8b0cfcf8be87212325e951787abbceb29a5e0027004ec471d6eb5b8cfa4d2
zae24c08e13059dea7e4ceb3ee187f4b5c28ccba07c402eae786ab061ac9dfed8f7200221e4848b
zd96e5c5a0f6818a46c4a4a68e16cd661a7dd212234b5655783063cb8a3f8cf6df918a92fb90c00
z5a236c4a81bb471365bba961942cf373b33122a3502622b7be73e95713c61f78afee89095a948a
za42a73cee47ea871ef739a786a68e899accb3cf4a2024bba2aae42b7cfa3de44975bca41d7423a
z14855b8bd90d9b073d3495388b898b11fe95bd95153f422657d0dcc688040ef781b49ec16c85cd
ze7111df18764bba65624ba569a5634923dca70c93f075cd0d77e7c57ab92815ca876ffb264c95a
z17272f0e548bbcac8426f36c0e00f4cedcdfa89aae61f7d2d0f8842356d9fd86a813f1b4cf0d47
ze7ee48787bf7fbcc7223e707589bfb7e127e098f09b992506014f3836e19b4a73dd4242f3845bc
z67ff9eb98835999feb4ebf4bd5579beb12f1f61209fbe156b2e4e1d3d3a2d9df4ff079aee643ea
z38275a73d96527209845c457de2fa32860addb937694a4ebe494b45b7e934cade9d926d6ed5210
z31fc67c73dbd7c06e8d30b0f14166a4902cced59ccf5122b8731dcd571ae6e4c33e59352d86075
z66eb44b7632b2d11b6537860751f363e3d254ffc1d79a52d5ac05333ae7b28f31997f5da454670
z55d5e1cf4ea657131e2b619f23e6d400253dc6a8b336d0e59d65648991cee08781b317f5d54f68
z36326a58518ef6f9c1f95da00c1db803e2711f44d1d1464de25a499dfdc935ea3c5777b4a3b83d
z97533057a1bc85a186740c5548fc99c63b0d6926c7a15c34b789644f3b903fedeb621398266dd2
z0d88f6eb81df58bc61da70f83da9dd34363c0ad35c43f640f2edde7c534902eed120e082eae4d0
z301d7a47d1b341deb66f5d95c038ee00ff5d967bcec2a2f408c62cda617ef77cd4a7a17320b6dd
z9f95b46b6fc67c905b3f1845fcfc0baaf0a0852b38c4f5732b7dc5334e93141a483209acef5f8a
z4e24bd551a301f5911417fa54bb192ae0bc79f610a6d74ebc42a05722380ddf7b3c13ca5027f5d
z091b240e6dceb3253e63a49672167b211d47834793f80d13906cf97f21e9028ea1e03f0b38e6c0
za86482c882cbbc87d09df1ddc659a24e80c207c80793ad7c7c85fa61dea5c36cf675f0b3d7175a
z101ac434cb0bb4918ed59c55bb2af6e672d780828594ae6aabe27ae79f65b8d28c51eacca8af38
z1921781f6b4685704fd8989d1af79d2ecebac2285f3de38e752f173763a4a7c0a1f8d62d21a64e
z6842367a35f8df42e60585f89acbcfb0cca89577b4acbbdcb15282adf669bce2ea705f80692622
z91d5275be238dd64c09f48f42a766201284baa1a530500d5723a58e7d0bf5d5d6a17204faf0989
zd8ba6bef68357f3c29cc3090a1db7ed39fa27aab3c3a3f929a1e37641f5202a0f1325db2310163
z1a92313dc245ae5a67540ab175a2304b6a312e1d162c76c297ee41d0bad56874a21d46e647f410
z29951ed46e77a1239a993b8f15abadf0f0490b4fac8bcc7ddb73f24dea710676919f1852273272
zc55ec2bc77a9314b2d454576008a06de3ce14b36695e61359ee5418e97a35416ff8b04a47f7bc6
z567071aa063d01d1ed07e3a4f6daa53c7d5c1e263b765905f952d4a7c0da4276de029fa308a376
z64d7d63bf8e85c97d330145c5406463e4ef0aaf39e5992f96cd7974bd608bb2e8247a834a43004
z4bf07312f904dc5436dca27256188dc8f1b2e9f050699c0af0aba3e5c258211bfe5979b90cefa3
z0fa890eabec7782735641dc2ba4f692a50f4ce7e2b876e36e7a059a6445ec2c4d137c31eab43a9
z10e0a34458f73735079d5a3aecf2dfb7f6f5a58bc04cbf7650eef3e349802355783f55d7cdd63a
zaef57a62c25a215e69740f7ff00c8f3b02a74f075a535410455482dec3f6f00511635dca15cf81
zeeccf9dac8d148ed5c60064a9236a3673f4bfc33008835a6c328299127484e38e41df84b40936b
z8211c20066d4b0e6e9e25f56a0e6148207b57c32a83710044e0bb6d0f9369fe5ea489efd2de017
zcca9ea7721d2f0a7e8800a62d58ac8e7516cea428bad8cf94de7b16b06c3aefd771f7428a3b8e7
zd75337206845943d9d9d39935a028fd5f32cbe911614bc0ead6f6465bc02509b2020648033cbeb
z1ef7c1f73939b911f0493cbb6f9ac2d153487885e397f2caea2f97d84544f682917e63f0f17548
z720d353c4ce9a05e3f86ddfd834c9d2199109bf8964aa6e2c1e8ea274c9de5d8d8bfeeca92a98a
z646519607998871cba8d97e843fc47a8741a67e9b53237e7f10b8dbb2776fddb73adbe53552bac
z071d997731280096b03f1c2e9869c723a7a0a61660370a668f3622ef775e63f33610656f117b9a
z5de2fcaf8ebe67b62997df1085acec5c104f82d59f71d6bc49ca81662594a1794a39dedec3ee92
zbc8e2a53777df1ab6ba903a8b275de667bcd27fd18737e203939db42b23357495f91c1784f1bdb
ze50d2c570c9be5a514fcc7f51d65ff5ca35b7b4b7512a905bb85fa035e29c54f5971aa26495e5b
z9437a8f3e6f69d431792f730d19e81cbb5accaae05b00455e3a42417e862dd95d3f7716f5b3246
za9af6fbc1576d608c7cf00bbb504265c2e9dee9fae44f9071b422b1514fd5afc8bf0d3203a98a7
z95ad8276441857ae502e63384240362d1cf6d85edae01e24d5c1c6d6d036b9adf518296cc76316
z8686c1f3c67ae1a9923fa0d012ea9fba3dff301851ee54453cf317a741407165d3ae6aeec5cc92
zafb37107bc67afb5ed697b38806343d38080066f308b5fb57e84e0d3551de3dacc47994e10b0ca
z381f0af6894d227c1f8ca88870de7aa0502a58e95d3fa5cc44a72cb6a39b30971f1543f6615577
za08e8ca87cd27e8de15b2a8d8a875af2387cce2c197c23ee4c5e6e83d07ac9a9c73e13744fc95c
zc2748700138ffe8ede99c1bc30c8b7786293b8ff79e606b5bff26510683c14ef8d71621ec9c124
z2047af9c8b865733c570cbe084d7e2dac3b2cb1613f3a788693d77ca0f767fcf14e88f4fd561cb
zc246e786b93d7a9805018de9fbbf7c79fa773ec8a38bd8a4fdf7c8547f79bc421b14f62604caa5
z7e5850e6f64173269407607e68a16f03baad3ec93a0280b07ead2b506d16a8560e18e45e80800a
z60f1e716aa8cb10f3429a3ea14c2807123b981ce12d67df49cd69fd76b3c0b1fb0fae606cab999
zd72d23647c3ad4997be12ee6903a4ab2f9cbabd3e0e70be42dcd9eae476574ff4011daeacbe5e1
z38ff14955f1d7de66c12ea6457075d92555fbbe478db549c2fd58b7d7f9392899b5e64477164bc
z21fcc07235fe3e40b4717f27efeea5f122c85e842add198b3e4e34c4d8eaa64554ab6dfab95b78
zd30e7dbd20b579f88507d4ca2a5a601ab600439db17bdde34dc76fceb4da6352533a4b8488ec19
z689c365dbbc1a878ca0cc7033bbd15b290529d65f22972eba76c2052fc6a9f46cb0b3708756b99
z26a407a5eb0c299e3869002d843980302efe7e1f809bf2066034d9d56c9fad9e68a193b4ec6dd3
z638f609b28005b2c1fff0f60c73b09858a11171eed7c1b699f1c2250d8ed3b2c989407bcce5ccc
zd120154c2f8a62860b5887081cfe12fed4c182a38e012db649562c253f18de77dc40df7d17cb27
ze7f72e4d91a0ae99a1ee61f8ed40ddfb7439d77dfb9ba12c35f1735e5710b81b16c74ae5150b10
z851e33078ba2ed7817208fe0fd39cd7f7b1eace86e38ba3061893e8dca843506882f95c4a446c5
z546c3a127abccdc85725f5c975245a242e3d5213563369b30c06fe2a6e695f3559ce49a0a25868
z68bd17bc39d7d797061a5cc2763c2f30090073111247a0fdefc98192d0e59edf1c757b6db36259
zf2ee9a84d830706cdb40e156c1243dcd8e0203a596f832933ff73aa3ae8706330d1f5cfd64aa7b
z25a1482829d6b15c382c6e85328af81a4adba823b938bb3a41ede4ef25941d6e80de0c0a4d85ae
ze516130b926fd391c2cad1de8b11be9291f185c34ff1d2333013ccb79199e8e3d8818770db74d3
z90f7c4ca975e497129a28feac91e230ed3532e6b1d815e0edd8a3eaf173409dfae401121d88d60
zc54aedf7d49ceae9602131f123f34bcba8c81c8e14944e02c409466da8ac28801c4bf5c9f9dd76
ze9334cbcd427878afbe5546df7941c8c0c220e62dfdfd4e8c0aeae65e03d8bf7c5e172da12607e
z00a9773d1e26b54021d28780db40c7c1ab48612016a20c1a6bfa7c939fa0d09767d226f19e59fc
zf695ce8a58c2063820418a04aa101029bed4e2926015b5c4b90f30b4e1418ec48fd00feeab4ec2
zdf37952a16b05634cd1e7f500ee19f66286f63008514531b00b946bc525516d79d764d9f16b26c
z30a86d2255054a15594606f87dca1f84a49590952f5ffb758832befa5573ab47f482e5502ba21f
zd346711adcce6060ef9564638fe6e9d12ccd6797012e047041921b19c98e0b4bade59b16434b33
zd64015f82e7fb405a0a2a5a1056ca404362a03b4ef2f1d875bf3cb46b46a4ec25971219011ed89
z6e9430e864795c31b724d0bc40933499b0def455a5ce41248e34cc58f082ab8cea6f158ddfd223
zbb29cc2e7eb1b371b9a171ab355c3b67eb48f44cc91074b4b4e1c357981efecd73aa84d80b3701
z519d4641239ef58163240045a55761141eaaa730b1e08d2b6c8d9ef568964b07244cb1cfa9dee4
ze406cdefe0c9848c2960f7bd5171ff2bfbd067fe321bb6cb0f01e086d1b7693bb4804618654468
z5f95a4adf612cc081063530a80198b0dce1485396bd448cfb90fc4a496bd0beff3f143e2e85ccf
ze58db94207e8c4e29eaa28e8ba360562863b7a0d796f4f04bec7fb9ae4c9d636ac46292cbe40ad
zc687e7735b0e6d603bb69922482f741399030fa6ef0c80c028c4cbb4f664353ca25d8f46979d30
z5d440a6b3ba84507eb9c76ce74e55bce530e16600fbe92361283a8333a009bd2b2be10c70ca965
z137b2945aec0a7417eff8f1574d165cbdcc2b60f9e9d132ff431608320c579cb91bc83221f4426
z1d165b0d87f314bf670720b206fc76fd5620aa445bc61063e6192b8323a8dda43da60995dc8a70
z42da0d6199c5d024fbc1b88ae58f6a3f48bfe8414bea9346d397d3a459c8c6cdd8528e61fd39ef
z428194737a4a6062df3c9baa04d9cd18e80f8f351e62d0229a8aae6879bcd707bbe925acc47d95
zb35071dcfba63e67958e2c5a632552e8ebd0d79e28510e1603179aeb53e9c4617dd5da4c036590
z9511ef6ce92642f638ab64639c21379e503edf11b7a9489ca585cd2f98ce77e553cc9e4a0bf3fb
z531feba5d174dab50e381fc4b0feda6fd2ca5b66a9d9e18b631190b65ec7e1b53aef70c1289534
zaefe3186255ec219dfc0b87b747cdd43d94641887d666029b7bcea9b584b579279ae91dc11c13d
zf5f3d75a41466c8cdc513e391282d71a18623b8f406db3aa82ae8a0607440262e811b5e90c2b7a
z5642f8ea1c04223c37c8c8a4435f977188451be4d494727f82a0151796cfb2194f9cc391604fd8
z937072905a3667813ebbc8ad9b3699396ee934b84eaae47c8f670ffb20ec9fd285f66bde32af34
z3161a15b1417753bd9319c7bb7f243848e19803d41befcddb5b2783cd9d7757536057889963900
ze93adee07b5308f5747e7a65358e10c44d2660899ab0cca7082e5a3c1d18dc523e6a32e0b72734
z88c569290ffe4681c813f8eab70d8200dc2321d7791805b8dcb90dcd5418b034e831e9a2b3b989
z2300d4049c2667b1491209b1e590844c458b9ce870bd0807501732c2465e11b37f7118eff7c414
zda42f1a5751e8a4a5a8ca1b30d5bb34847e347ff5e6dcdd4598cda4814788ec3c40ff2593e7e9e
zd5f4dd894cc110ca3afc50788426ee5f0a231362a054d65756c91013a8ea6ea51adbaa05b1c12a
z10ef188bebcf1290b549c4b77cfc874eafe5439c6005fff2aca90cd073ea4ae9ecf813c3be8b7d
z5d2ab725ceb61d77211ef611d41228870ca746c413f0b287f53884510d529993c528017ffc8825
z8b1451d8a58f4b3a24dcd66b65a597789971db0a5a5510ead52d316f17602304ab882248fb4d49
z784fb132f941c779628a14890cb861438f4e0261682807ccc858695e16d60ec02d8b97b5c3bbb7
z7edbb46a6c219419a0a35b357906267e9cb0360e650e996893288dc09fbd77aff4ce6dd00da885
zeee3eb1ce7d74a968f0c72fdeef49c6190c473cd8f2b6f65725bf7b3e52ff7f6ac079efcd5ef4d
ze7b4192df5d7d92f11ebaa1b73955c3eb5b6c158324bb5050e1a5b933a0825352bae23b2a0fe9a
z10af59c7dc2997197678a96928ee03f9d66a3bc34e7ee9605b32263c845621d09456870b2e7090
z4e023cbb0ae3519af679c275c8060b9135e9154254afda50ca70d348ba0f1dbf0a4ff172a24397
zf73bcbd76aa12a0c9fa4f388e42f3281952922c944c62d8f16e98f4384a5f4b78f8ce5ce30ecc6
z0d8bd75d21d3049009dab676470a04f68b6c81a9c662f3cf9f7f92b89f2c05572941f5871f657f
z7eca177a4d9dee8dbb2370a6b6d3771c2221a68f189bcce58cb1451510cd3609214b481773033a
z57f9097190eeb8e9630108481e478a2e77922b820b365e3471175c00bf45a9bdf3d28a56f7e168
z4b8a8ba64a00df87ea1d856e669fd458f80276b7c45d307eba1ea1dbfdd5af712771eae259e5ca
z55351f6779d65f5fd189b8e4805d40a0de77bff56304093ed1e905d6efd99d5e76a7c89235c3a4
z04c0a3d6cc4a9b44999100d600645ea292146b6445b57251c40f53795bca11935ba1b758bacc31
z32f1eddb16ab94300ddef76dd77f922b68734fa3bfb1706306c4c9e8f21f383bfeef84232b5cc1
zfa1d6b1d0707aa17a763de5fd3fcf1cf0ed644e12d8c171dd3c3aa340f2451b0e7883d5844b61b
ze6650fd27be94e33113887ad8cb20e71e2adf45b64454023ffc6f85e52fc3e7371f6717923dcac
z94b31b05800620b803aa235c12e9d17beaee17d0d36e4ecee3042c9acbf001ce30620992f84b9b
zca778cfe71d6853a16e3fac95d838229c7e9ecb7cde51ae04ae8095b194cb8d8e18ec59bdf14e4
zac242ce13b938f823f715a58101c62aed400ccd4ff7777fa86434ebb33166f33b80c5ad3cb0757
z302765d1359a42c60538d471140c14846275d4ba33c9e3fd5bc446fcd565bcab6f7f4fb490b3b5
z9a0fc98ad0467e9cd219f74023d7fd7c84f628c7ed44da707f2ac9b639f8aef040dd494a15645a
zc86e8438058572c5e7a3d848e9871229d1681fbae3101ba02964ba867356b8048e4ee7bacb81f9
z33f9479617f8f16b8eaad769deed3b380f8a975eaa2c7d9c1cb60724aec4cde71553e22017e747
z3d77ebcfd4bcbad8677d6ac1b6e644f1bea3b9b2de859db577a39a143f3b0f2eb23ccb70f98d69
z0acedeb3623c4b28a7a733ac9c56d2486afad9d75df102de5255bbf4c95cfca20493b023dd57ed
z283591f0ea09054356b0db2a6fd4885be4da86be08221d38506bae46dd4b533e759c040e0a1491
zf47fbb06a78f9635f3a6d7d07354bedf0b67e8b83c135c049c91b0a790daa307f6c89d2d4c8f8a
ze71165d9866c766c0272c5ddaf7c88abc4e96510f136895feb10d45432fcac686bcb086b42f87c
z2decfac008fc55097e6cc6d0ac40cd3348a100812ded076601ad694985c52f27348eedce6b8c2b
zcc5b8ce269c4f320b2c2dbe67b857a86a0040828b4751e06afc50e13fe926c1da30fc1041992fc
z2c371375cbb9179555f1918dfbd9cddbc03745b5bb23630412f0a6229fed10fcaa207542268e09
z90b20ff84909d293be32aac51d1ada5c605fcf83fe454ee3f5b0c58ae89e4fb1dd00e65edaa2cd
z89fefd264fee6659a71ca20507e682632e3b435ced2c42c6050482accd3d53206cb64ab46db915
z0cb8ef9ad594e7babc8bc7632c9458f58dfcd8661262f9dced8edbbea2581b5cb09a9f620d5734
zfaec7f6dd3aeda868bf6120b232620db47195f188892e08449e8524a64267dd373366206c5ae40
z75c8066646efa8e7f533adcc531ff57d42ae96094fe2d0922b935957f2e3bef50ceaada4d5559e
zb2db7b9d13b8160d62eb1257650e17f06e36865e432f7b84520d339cc47c2e49e3aa1d7a45cab7
z4cd46cc88c881cfb7cef7cf8f8e3c992117fe981ae465b51fe63b194ce4862cc810440f9dc4a90
zb4d914fda6c6a043ca713469741aa3f528b8fc50b2467a52bef8645787d69818c8816b5b2bb2ee
ze6af56458fad7fb46ae72020487c3faa9e3fe3469a023e3689d5c5417a38375a1b98d8ebddfddd
z5cc170473c86333a74954eede8e149866dd761b2f2a632001b8bd87ebcd9bd22bc7b375ab40f70
zc8ff7f79db91eb8e72b240b0017438b5f8c4e0bb9583899ae78962414d6be3b78e2523f905bb4d
zcd14437270b10b39d83200bfd2581ea6f0f570314a4dd598f70cf2a15e9037c2e6594806a28b93
z324e80b9d35f59f7914625a28290b01454e7658e166ab12d8109e4775be5b5c7b905585b58f508
z330aaff284d26254b4328053b854ab05806ffb46670741823fb6f905981b0e5811a304ef80cc94
z5395cc92ff580f0e8c231be5958ff22fc0ed9d16ceba439262cf09fb9807af0c3861609ea2f785
z599449b958c15e91505486b7e847b545c76d7ad88a1a77cedc3b599594c4ccbaac81225bf65b59
z6d910c9b57756425d1fe7e12552cc9a435fd388af25f53bd4fb8872b01d5c01ef5b6dd3ee1f174
z4717798b5b02b514ce594b5a051edf0765598ee42771b42bf8788467ca07dedf5ce893b39c5f42
zcb27d9a4145e2af7d796f8c1ce9a8428990a6e88008cf260c8956bcfb90c179aa90eaebaa77200
z28a3535ac51d6524ac3debf634467de12143832bbff3913853ec4356e8a127fed57db015801993
zfb4355a67cff3ab392f96b5389707dd6ebccf5ac477485728bea55cc968748969e6ce7c92cb225
zb607970153feb1d80af2070dfa68bd4cecb5ee4b349fb3c0ffd5357c7eabdb7b2efc3d5a304f37
zc2c2f38803ccee4c4fb55a6aa160489861dbc917797cdaeff13c1584d83af7e1c8ba22d71ab063
z7d8db51de726e6373f0c9f2b20cad50cdfd8dad5efb03bf5729a1554567aea6acdfb0f51aaa519
z49dc36bb4386b478af31fa3178cf315098e5ccbb02219f9b46682ce79dcbe95dea72cb7246b206
z94f416a35d51e31abb9495faab260d9fb13d4fe332bc4f648d9bd0418f332b38a8c980adb44060
z451712d07f31a3bdcd9de76f3c1d574b63facfff413ed17d1e92276e00ac9de049d87a65c0b065
zbae646f7ce765d21a91ad7b27fb5d633e3cf70bd25c98382e11c6aad0fe7d0e07ed4e0bc7ffc7e
z595804d180259ea01a9f0955ad69beae2e207374d4f8ea3645e0e8ccd96e26eb1b8b9138968b58
zea47e548d09cd43d4dd6d597f4359216a75708572d674966bc3a70294be0f303267f56131ef71b
z001a89deb0361fe7d62765931f6d97c7c4b950cbce9141a9a2305147d571d7b4625d3371370e86
z93d93bcfff442fd66e92bc781747f341036c8be2ff9e5e829245485a433346260848e9ca25d067
zfff7541d1b83d0ce04afacfec22d992d229dbb13b6ccd9baa0a3441bcf815ae49ac7a7af0e4a11
z3dda96202d06050f7b9f573b5620b84b77d0e57beb217beec02b19b675cc7cc03e0c48767bde6d
zfbee9f9db58a1d4d429b012ac1a33fe34f348e22f6ac7184462cb45813c5f77035147ee5236cb1
z467457c3a8e650346a5374c8232a9a7fc52adc7666e650ce4d0cd7ba3b1c48ab18ea05c3b35ab5
ze3d922a935257c20b34b62a4c95aba0d5a180ac28c717966dfe7ebccf4cb1699ade7374ccb45d0
zebb75d9b66380b5cbb0b71da566cf6750f1b5859895d74c889e88b585fbbf14c4176ac26af11d9
z3359e8331ff71c163c86182954a329ca18073f4db1894274bc06731468542aec3ae301f82b7bff
zc0104dca9aed649dd074dca2f33907fc83a42a736df91b8adc5af880627f14859b121b0f6e7df5
ze8f083b022c9f69b42ad8b97d4b401beeacb05e4fdf69e5b6265fbcb42ce33c2d0534dff1818b5
z166ae05fe4c1fbb740c29a64abed23cb00b09f24ce24651f8392ee0288936ab2d7381a49134d5d
zf1ccace3ea06f44820d593037cedd6bc6a0ae22b47757d6e6adebd605ca5d85782e3995fcae18d
zec6a6fcc5318635792d1d6769da26cda0c479165b582c42850557bcec8f3c100e1d67d49ec4515
zd8acf9e7ea741865da5c9a937eafb46befc56fef1cdbcaf399200a9434e777b6b5df783fa9b13c
zf3eee26de5428502e6078a3896912bd73e4ca77445c091450f1a0052ab8d817512557f570e6d4b
z1c7918f5fc6b1d5919da78bce74abfc1b820fab5af0eef71c722a18d546eded86e028b58e413b4
z201e4739a18d12386f2b831685982c2c281d8e3c0a38183ef7bd124b519c61cde35d1aed83332f
zcd5061a4a7e2c02dee47e508ce1c0844f3b6f67fd493ca0ebcd964a9d27e58d1732e94b3635679
zc3032927ca7d95c5a342c219f0c1c0a89b53d1a9ed6e5520cf5c1f48c59d08b488a8276e8e383b
z79754a52719c398add07e1b0d99b85937b15c700ac8512fa74ff47fc469b2e059fabb98b948af5
zf0f67492631c2bbc4ec3d4ca8d8dca94b8375c9f02aae1624dcf2a73337b4c4d2b299c6535f72b
z9663501dcbf6f09e0ac495103d726a89b037bf0b281a9121ff5c7d48494831d96f96b846784073
z165cbb7df3156db74978b01e1847666aeb1144133223740824b455a15fbea477a1f203adc34a33
zc7d93b2d306a9d9e21c6ab551dcbb5f96091b263c6843966ed9f6141fef69a24f27a124dd9ee0d
z71b4449696e165cb08301c363aa84fa6ebf4e5cba9cf405f8acf8ae669220940042a9b26f17c89
z47614391a78d088e41c943da3384ac7d8e5518fd24622e38f043c6550244d92b6ed3e08f2a38fd
zbaf0c725101bf947f1ba7b02adc0d79b8cb81027688c2107fc59149d37be0c3e3ca104a80246f9
z56a7b9e1aff3d05a2d63525aa43acac758db4beb28906649e8e06be2432d048c8e6a66d0a55d3c
z04761ccac073d4fbd3ef5e569c5a93dc4ef09efa0c2103903d57a51fa9a55d9f9ebcef8514ddd3
z29ab082377d62410e3d90af90c7e215713f3cd4fe7f996b7bb075fa60e5b2933df48e03fff636a
za2d463e4ecb11c92d10b35cf582a017eeb041fcb5f45e4c9ccfa756e4ec9e4431fd56168537f9f
zb9212bbf6f52a08193eef0d7579b114594615692e018442dfb36b2227083d4886a895cb9a0e354
zdf0d3a85ad7899cb849bce939516777c91ba02eade0fac018565d78b3bb5a357d55a5a9b1b8bf2
zd5b0f1de8b756b3771c87536182127d71f9b75e59f0aa0c3625509ad68f3efb8d3fa1da7373b7f
zd81a73cb15df5ecabd3f75a65d8989249a930886614f12e1da9c5de4f29dd1f2aa36d5273549f0
zdda23a57b2d91853ce6c55ed32681a464b69cc811d8656f47a7ffee3fc1ca98c5165519c1b60d2
z7e5cd7bcce3a6fb1a0cd6c1dd71957ef5cf48367365775c01ef7b7866ac7056cd87f6d47404dfc
z8b2a3925874360dedce022d4b654a5d8eba1643b601cc95401b6453c974afc27e07eff10d776a0
ze4a898659a88c49bb7acba94e7820ab207aaf7cc6cdff36d1c2de05137150a7c1cff12c7b2a738
zba7c172c81cf0ace19add4837dc266472970cebc41887498c06fe0656c07c9e90635cd0963ecd7
z835ada9480be9010f06bacc8a528374bffd5dcddb6c91e7e93ea18a730ad32c282fad69cd0f272
z568c6d076387d87c3d5d1ebb2c89968be8033a83c6b200b0ebf06496b46759d26e6ed8deb5fcf1
zfad8c6def6ba8cb74cd2e7bec110244a3ff535d2f845a3b57de9cb207c832c51de46eb2d5af683
z0058a8feeb7c618698598d49ffea2b57217b53db8b314ccafff0d76766875fd08f1ac82b72c71b
z85c38d0ec2f21a4fdbd250c884f0e3b2448ca3190492dce140f70fa00aebfdd939d6d65e4b3c94
z9e67cb4c2fa549e22190130506142f4ca119da2a97677371ace081a1cab8bcd8cd6977c6a0aba6
zd0e94f9f65076fab53f431bed252354f04ebcaf4f31e8073093d4d8b6c7da24b695c7dc93630df
zaee3ef1d5600f8d86ab1f132f21585f742e3514c270079b47851869fb69e9c2679b13924a61bde
z9d67ea636a38c5118acfd0973645cc36a1dae26cc9a4e010c0d16eeef11f4738c56911ee6fb274
zfb420b20e9fe28b8c3bc07ace944d0a81c59b35b403ace2b2162ae61dc04be7e53d81ef3a2e42a
za4302c5850eec93a7f9eb0c9ba6ee92cb148f021e39273ed46d8be67e3c4fd560aeb8c2e5d1a9a
zd4c38cd43485e0f0ea0382896986f0d527894c028d3e778d5798aa7c3adc21ff6cd6fc2d514d51
zcd19373d768eeb8a3054f1053bcfd7e9946c49796152739ed661ffbf1d67c618a0de28233b60a6
z3992933cfd29cfde72b2e879d15cedc1c370ca49de02f01e1eaaddd02a52a98803019505add271
z7d69c6b360be6ebc271498334ca425eef10a799c4baebc5243510d4963ad29d2a280f6a8d3e065
zb95ea007113b02220c48e7a5052b60bd7430aa128e0ae8e6432cc26e1bcef2ce6f53ef8a3f3790
z50a81d66d31eb7aec7076974fef09fa2e076de2ce6792c9fa93147ff3a4eee059e9454d55dcb17
z45681ba99dc4a0b966514ae6ff8ce13d305946dbe7c563123601434b3e3c7e6f535484841b31bf
z035c0266971f889fbc281d176134bdfe4b484e9df014c9cc1b4036ff766af2441587dd5d2f9cd0
z9cae413b293f681e70bf7f508bb48180270dc2f1140dafe3d348e11d0796c0d1e02ce2de4544c3
z06ef76d6a92193b7c3417e38a4269eeb6c8d380b0986bb6f483c863337ab4167e2bfb32db779af
zf3522cd544001477e8bd9aff638da15e24ee8999b8825c5a46ee0a5e99974fd7577b484161240c
zfa34902d1e15beefe224493198a60d2a55ceb7840c099fc21bd74e0db5a15d303d2127fabbc99c
z30110e94f65daf0288549240b363c926eb848bff1be041dd3098be64560e924713079263f8a3f6
z22bc4484834eae0ff5c2d630284cf3e48c99
`end_protected_0in
`else
`ifdef MODEL_TECH
`include "qvl_decoder_8b10b_assertions.mti.svp"
`endif // MODEL_TECH
`endif // encrypted_0in
