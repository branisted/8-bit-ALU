`ifdef encrypted_0in
`protected_0in
ze74c34e226135848fe16db9ffd31815111b6d7fb642c521a3f628cf6da949865580b22efd062a7
ze90adae0e65e66a2c36a587d0a790699166942afea5fb71013544a379d857e14682c5236087669
za040f2dbccbac59e8bb4ed6e90703eabc5da3fcb4cf9f80aa1298f4671fac620329c218c100101
zed6f713217a0741641167633de77ed77c2548cf70b6855633c380db97da98ee96bd521e19fff10
z0742589f83f1287fb5cb27df129bff148aa01abee5ab49e22511170fd96dff46c42a2423cac1da
zc3ceb4384b5198832c65e6b94b52b05b4487b3c735d6a007f05a329d81de71f6f0af02300ad959
z820755ac3bb2b166d010bf8bfdb8726b6a10a3e54ae6e789051bf1b87e86ef94d66538aa03da6d
z872502dd8e5c09af1526748a380d58259c52a2be1417f2224eea7574e4c3cf7da76c52b788f57b
zfb0006c6b9e2aa4d0ab6c54bbad65e202aab8b9234163c184166307cd81ec7c0c1a26398143578
z7e9bee7f42df35c319af4183f5a400a074d386ac2e0a2bf8855f12bd8ccc8e257b87f740006eb6
z31549d1bb749767b40703a8042aa7c7809a76a73547ff90ea233355614d4ff499308e2426fd8bc
z5b9081418146cb08fe1110fa8732194ca48dd3a4031f6c21cb94cfe63bb55ad6c496dfcc40aa39
z89e81482736ef3c0a1734ba94ee246087bf865249cf443767f6552f970ea9f085c2469fce13d20
z6e350d6f9c9f3576f5c188c4f019264336747603027703b8dfdce13bee506ba006dc89e1dd4d5a
zbba345d8401c694d8b9dac30a70c9c6f52c876ed5aa163beaa790993fe30105b49505dae1f4e4b
z15079a4e2633582922fe8bc280d2045f3c503d8e0bee7b2109e98e3528c23e87edeb04cdab76ec
z8f686dfdcf6dbb3c7bb28d022ba9e5a9e75ef6635b9ae86b67e250514e0532390b3c9eeed54bce
zd1827415d801576d9cb4360e2a0535aa736256cf2eed3ac098a01825032bb1d1518e4418742b60
z49ba848f7853c632da6b710ab42991d0eb9d03018693d96177bd76ccae38c2d6e49aa2524b6fed
z48316682368a9c9474ca6536756717be61f896e67551fd7bc43fa3e0151006ed872c91ae89ba4e
z8d23f936b09184f38acb9bb08d2581826478068c4e69cf0b9b1f9b0b4ffd9a8a56fcbf73f694c1
z6241645c9af1feb42bbc04b3b5b70e02b62311a79612241cef056511532dfe57797c56624d93ae
ze48ec19686635c2e8f00467fa2541e617be9f8dca1f7fd7e69257d5f76996fcdb68e3b91c52dd3
z85a9a5fa439b6094df8410dfffb830b9a0945b30174cacc19a0a762af2e2a5f3595a9901fabdd7
z896ab8f7bd7348d9fafee65d9c311d65e258c0e281c1e701716719f5057861d0115e447dc50e74
zf91f0babd168ec37742d299dd1b36462e4537e10a6669b22e812e54b88cffca395f7c92f38ef12
zd474194038dbf47ad8049ce5ff25c14e2720cd260ae318057895b379e38236863ab3757f8d2e0d
z8525f7ef431e8aa2019ef4b71f1b27e82f497336c6b19ed4b52b5947f97eb585c7944b33c6cc33
zbf135d0d612e4f3d65ce524c7c37bc1b19342555596932993d28ac21738dcfe04acf5d1adc3a6e
zc7164db501b7c652be3e28aa09208400494f5a5db5b78e5e990d7e9fdef359e1b964ab0aacd792
zbb1ab33f266e798c1d7d380293eb2bcfc6a04dfe4836a2447c20d3500bf692de0ae8f50afe6c87
z36d3eddf789aeed346a10c5628a931bd5bbfc2b727fae0dbfd0818e78c457504138fc54c7267db
z7be362cd67adb9c6de23f849500f031755f3a600130b2caf520cf59b317978b2adbfa3fcf2d9a1
z0d09378efee194143cd6adb9c5c920eab472feb5b31012c5ff1d9ec35acdb594574c941f284b4e
z79810af85fa1ba374cf9597f5ba31ebfd3ce847108e5a86ff2d03e060b7c9e2c0e13287caa3a50
zd407de7259b3e5b502255e6ef5d7d138539fec262070e5384d41dc7e651897423e875b2a16c60b
zdbdf030617e9b1765643bfb4d1bb6d073148d933509c7319e8b2da96de302541dae1a4b0e81edb
ze71bd4b44949e7b7fb5c46a519801ad04ace6f431944b7efab9f09000d6a42c0e399409fc548e6
z71b857926f35211acbb50c02668f3581bb0936329c25d0643bb132d3e9e154702631f0d9121fc2
z2e746579148b6806765d0351b6868af10f0598dbe8e6a72ca2df59aa18acdf7f8bedb99d164dc4
z3bf50080a14504c54a41ec06b80eb14c498d3113a15bfafe9f0f7310346b2fd2503638a24d12d1
z03a21584bc205ef1c07075482e3ba08911305e68360f0baa0ee13f1082004428e2ae9f044d7cfc
za58f0c1a24e421d50a6d54a432bee8e1fd8d6b34757d307bd146d268f04fba977081a79a25649b
zd06d525a509135e97c13300d16e44315eff28761d6570f40fe301540776511743eb95a27aa325d
zb7c554eeb511eb16444783adba011377e51c9f6c98ef99d548324e35fe46bbcaf99f67aa6cac13
ze04c19bc76ed22c2075b805371c30e3002b7a8e4410154ce45553eadfdd820fff3b7dd777d0890
z5953e6d9d0a96adb679aac96c67e72708379d840658bce7f6eb22de34b65aed6ad6a5a7e02aebd
z32a321ac96e2cac2cb48315b8451d8ca9e0f33c741fc94ef3f094ec2b0f46b42a0846ef7c7eb60
zd1a54c1ebaba8fb991e386993a296453218ab99d4ee0abb0dbff07f04a71d74d5de689348cc6e7
z39af5f9525c2eadd3e668a7c16365ae4097b688007eef2aabe512663e66c4085fcfedd60bb98e9
z332f2e04a287aa52f50ad1b3016ba294901cdbf28317321edacd6e2ad0f4b54f7abb47ca776b5a
zeca13c1235d85d9ad36072e85cd2c5841c87cad4ee57dc3bb2f0083064bc925554cd4671ee8ab2
z5aae00895f4a0a8248e76e4ef3e9a044425b28f0628823e1cf727110d95b36e62adbcde18801e9
zd8a93680b1c12245d66d3fb7df63b30b81e5e7f0fa4dc97a4e182d41377095bd27a8fb24699423
ze1202be54f211264cf25f8e2a4f584299eaaa10ecfdc1acb31f8a461daa4490c6249ef06551831
za1e87213839084d7ec2eed41381a8c23dec85e518ae895004c1295b2e7ed3a6ce6d23ac6c91b81
za90623fe8094f5f0881d2e57e8b28008a56699068dbeb59b8ad509f5d9c3cce0adbb01e3e83f86
z386527734561b8d0d1397bde478ab217264dc52743b5c7ca3e36de6206e6dd0559eb0c4d3c6243
z0eb57e83b6457d744effc57b3cd073e317d69a2740e0a2fe61eef0a39fd2b7f64d936619fdb1a2
zd432d28333bf13152beff8205811f002ed477953c07b728b26a65f02aa9c2479c26e1e66189909
z53e6bdfa2404faab0d1747110c773562e6e64aaf91250527f537ec1230a9eec897926b8bbe75e1
z20eb33f1c21b67a26931e94c4e9158c8b5f9ef0fe1c060b117152e7cf5f74de6db2d29c5bf89f7
z88cbedaab7f9463859043d176930f9de4eae65e561affc6e16e537571d31c4ce235facf03709dd
za229d588aa9474e4e3c75fe45a84f8aea9ca42ac520d1f72373d61fcef30401ef1917f06d98c98
z7f08659ebffda8e28e71c679eea4fadafe55eddbf98dbe67304c3e0f40c9b7aa7af8d4309e56ed
zb0dc5764e36057bc9e0a472f55b17d6740aab5900383fe4c249dd1bb6756a59d36bb7a7d4ce1df
z17193eff022a4a17891f28eacedf93e3da72b0fd9ef38adc6539a6c52bf3565a6b504ae39d1d70
z69eb0790206e8ff0f54f04d3fc03f18cd131d0ae9c3a59cf84e0cef154906a4589d9c4c512a55f
zb550bde078a6e0f87094a62a9e7577b6394a3875cf6f9a6da760bf07a1ff499cf05adacb2b8b84
z2e7a8385c72f7712dc26e220b7a1f13aad53f97d4131d9d0175bbbe6d95b530e40c241696158a2
z74bb0df059627923e09322875e0b965359d385a64dea1d455866d55b3453446ed8b6397062be8e
z6c3924e3527ef4e0310ca2d6b4dc771ab8d360f061d9ecac093efe81f75806eaff682628a9efd8
z315cf80bcfca341ec104dcc03ae0e406bf8e88fb51d1736cc450a21325ef51ab59c30fb599029c
zfbab4bbb4f1171fe700075f65283b3a29f22945ba502470c758cd241ab9897a2fa22f1d8f6e156
z6101fad566a06484605ef241deb18724c71b29e075c827dea6684d658f7d3d2912d0adb8f5567a
z266351bfd79dc6a4037a1e7b54aca2e00990fcf780b38e4b36189c9c7dac80756231ec92243387
zfc88d983e789c2337857125c85374ef33cc3a2541451fe02964e74f61acd26c37574072accc3f9
zc02415f38c9d3b03f24fdb0e7709ed0c254588d63b38d834649a7a5b6b7dc8c111e5736e03cce4
z0a41b37349429382304d79771260ea35d684fed5cbfb2ec70085cd68899357022ee647b1114664
z6beceb1dd7cd4171af91948b891e0d786d94ac95660201aede2aedcbe040a350cabc24c29e5b07
z01859744924335c30b3a2eebe899a7faec787825f66c3604c1e89376aeb1c5f966e9240e83e890
z75b77293b5c2371923382fb3051ce2b419121accacf2844b420433f341fc3fcc9ad9239ef74253
z8ef3805912a237128fa8b0f2a4a0690f62902b77250b03d19480fe8a07af7138f87ea44d084674
z3d99e90f4c5e9a9e2f45117db13d6e537ce676f6befc342fe7b4a09505b598aaec32b06cafc088
zce455eea183edd6498a8cf64af188864fb726f020f4b838789ecb018d4acd129462f07812851e0
zc373721ebdb75c872bb90b0036eda2d000084cb33df3f9ae64d1c2c8a43839ed182483c362b451
zd7b9cfe26be8ae7e56a3e3045865b345b6818a2ef22fa2f5b4770bafceb5e2dee40fdebf889999
z687a62988b634bdcecb1e62e9466c0aad12e5a321ae57c0361fd9a66ab2174d6bf7b1b4ca24951
z56c45f4fd1b37c8e8a28e58290e60f744dfd0e1c8e81e2e7d56975ba7f0a69b36b23ec701adf82
zfb1d4c227caa7f14acb0284bd3ca4ad0cfff01f845f9ed411c21c1c61d804f0643ad106cce5193
zb22033d6d26111cd95578605aba1134584df1cb17d16dfe0aa44fce0beec95958914a35a7e895b
z2332371d7d1e35dc2a73df1791a5e34cc4dde073305d12bcac779f6ba432cd91df319c7bbcf462
z6206bfb707b67634c98ec45c570562bef164ada4a6ffcf329d5006e994d2ebb455ba9eeb722259
z8941191d33f01b1c06f138a843a33eb2a292064d5504d1669c553595ee4a2ea46754ef78efa70a
zcdc342a2f2eeb625d728863ca1d9415b78d71bc4bd806694eaa578af29ca8c0b6d23e20b6c5579
z3362ad43cb550981006fcb452e5c8e66abf93521496edae84e946ff078c14297da8e9e7cd4de9b
zcbd8b256c0366eefcc6ecc2a845fc6bd0761ec3c3cbf5e9ee45ba52745d6c946898b978eba8479
z81b2bfdf9128f8ae88a334ba5bc52a71086aa10e8db403ac6d8e6ae722787a67ac0683c930a8c4
z4185d2a45d9c493518ca3b622c0477a49907df5a0d2b47c8f6a75bed796ba7dbe16cbec0d4eee2
z04a07fc34fcea0e45e43c2310e38c8ae2b7e07eabd438bc5c3753ee3668edf995430154a0fdca1
z6bae7ef753ca7ca160f3c5e620d35fe04dace57f7e1ca5d411d8fa6b075262970c13d8775377f8
z23f30aba7854da658d311e6a3a1cdfa166892095232c93f1ba3f23322059bf63ed9af0cf3226e2
z6af17d68aa71cd368ed05aaed09e61895dc1551d3bb263b66e654586615556e76bc516d7e6cd50
z56db637f36634993e48ef572184a607f6e7a629926a2ec6795127a3c6f2d63cf16db3922b4c5ba
z23fd2d12847da5a428373401536526dbd160aad524945ba3f3ea865f2562f1c791f2544d55a55f
z82d19ab5e949a655bc781008c556a7a216cf69bd2b8f0c1ba44badd95189ade191ba54cb7ebf0e
z4d5b2f1e94773fa0e1a8c464aaaf284e80c12e0f0ae1d6e718c23c77a0d60da2de8c7e41e0bb77
z7b4eca214367648c05cd9b970c78be6a0a7e9e490ec9cca6c6cb2b6c7bf578ee5d307c3d4f59bb
zc2d885f38403e644f7458f138f576a1dd70630f05a80c1e1b56f8a951b9ab6010f4e55f1a59fff
z5c01ee92b11945ebc17180e8d4686d774222b17dd6d5e2f9c148d5b3990d45dcc037663e884472
ze1ecf961f71670462604a676ab1232efe701f2c08729bf09e8c717eb4268e71956bcda412217d3
z335b6f32964a234d075dda64e49d4a50668b6a548b93c8c0b085200b10ed0f330e3519317d0fe8
z731e22ebf25bd052459e393a4ce095949dff0170c5f9dff608a042029eca27e69a36c2eead12e8
z06c6f041f508bbfa98e723eebc96a847ec7650bb98d93e8a5308eacfe153d7cd9012bc6fd00418
z88450b446cb2eb65387e271380a7d326cbb52e517b2265fa78a033c3566dc5c9a74a622eba9a1e
zb161cb527f241a875a4d288383ddcbf74ad8bca5664f388574a40d07e93ee08d77a5892814bdff
ze9bd86e151ff1b66e3608f397266d280320f2fe5511aadfb3f9adae37ecaa2baf9d8140571d27d
z372eb2b03dfc7783b2f461e3ac9c40dd0db5156c2c874fd78b895a9c79295dcc924cf44afa56f1
zb9d99c679ee46eca4b091fa52fe08c14e6c4db8e3f05805be16dfb60580c37d954c5885674f336
z91ede230f94ab49d313a18a291887b69b40d3dc4eba135a0e8d4f6a3e805ef3f02d67e99e7f444
z69fb3024d8a0bc234075c8351688b9dfac6a9a4b48d65335ca13e2c0a0d41a2c421d143f381b5b
zefcd899904c4b4b42fa26fba7cb5c5d14dd855eb8337d4ad3c047063ec2a62622671296085d789
z293eba7344d91e61226c17e8e53bb6d06f7153cfaf5c4812c07a5e2c3aa0692b9bd44aec0ab291
zb4132ea1392d643ce0e57a3658ef2f0ff88e1f3a2d1846f115f6383c072b9ce29607d3700181be
zdc6e50f89e1c1727f79f000c7d421aeaf994ecabe2f254aee03dc63e37efb749a83d52a9012931
z5098fcf6e7440047d87c59771f5dff8bfa8afb8cf9e82a306f58795de434e99a0825baa9e41d07
zaab0d7e31ddfd727ab30ee3b5c3d0de6710583b4532d1682bc5fecc7c367a34e633b27b836f780
z18fa25b3a453e356f3afcfb023d1bd58fe276a5e6a01c95d5a54b91ba4ac18dcbb2b26cb4e6024
zc160381db735806b64e18b261dfd6b5a863de0824ca62367a098e0f2b7353252995f1560d52c7b
z50904b78502e22a34faf33a8fec9d2bb57dab354bed95be6fba10d87e48aceb11de832287ac5f9
zc52927bf1688f8b4d5c2efea22f75b2fabec7468808b305a2bf60b305a485779d67627973d3691
z8bdf823b546182ae9616c0267216f114c54673b82db58c8e5f42f52c25c28a9130561faa43ce97
z0544e4b8fce991fda4ed6f0b3449aa827156dde501d1f019ac811476aec2fd57c4af0633a4d251
zc0c8df2a9e7b0476703c85c2c464491a2a0676e2426989a05e253cb38a77f10203a169b3219382
zabeaeff7745923a9af558c6121cb4700c753f7fd545e5885ec59fff5294e269e9b1f498fce2a4f
z0a7c064d4a5ed879a7dc5129f683bc02f82c6498d59f56f78e61b98629a24724857a937b1ccacb
z28e412c85ca4a62ac11d8ba9b5bc882ecbe910d6b4e4b49d559472e20e93b3fe615b4072ee554a
zda347420176c1815b1992fab62c7d204b4f79dd6f72d5f921709ec493028cf8331cb54d6c9b459
zd3658626f6c68dc563c6719ec754ae22b0c2009bb5411a04e3f89f18c7d734a1d46aeb57118ccb
zc8eda0113f8db9cac54cf9f4cb07bb6d4b00f46196232d8ab074275f5bcf6df8ee8861cf097973
za1d67563710fce782a254f2b00c7782425052f9d9ff7d0c29e199d6bc2a60f1c62d6d4234c63e9
z0ea037eb1c7020c6d712823671f984b5d72bcfbd86e44b3b7f0f95ae8a4975bf56802299cde51a
z81c0f17bcd9dd4caf275eb0bccf9e43b94f380a78558fb358c41983575d32f7af3357b8f9e75a6
za271251fc6a41938b8e144ead1ef1aa0bad7664dae09685e04bd22100087be0c1ec39ce65812ce
za9fdcb202f1225413fac6e43a03e404444cb46497bf666294097003421c50a98a40c1f8da314c6
z730ff8a6b5585ca2da7ee936f8169563765a3362a2073a99b6ed44c43fd6091e33deac5b6fdae1
z6083fbe1189f6ea360790c3099a59991c1d379b5e915a80840bf69e6eb803913e56b3860300c88
z41d6f5e06cb5898fffde1327fe94e69f906afd11d9e94818e77c5f9afc490aafef06053e5e77cd
zcfd47e9dfb9fa9c9e055aed5a940db73bb676c3f96fe4a0fcc8515dcc0fae76a74a50463e5667d
zaa80591f297cb5d570e483881d003bc6d971b5dde0171fd4f68b338337d5a6dc6fcbc88c012862
z6011ba9d3952e57e18da51b598b16a6843b98cc914a9cc3f28347ab48398053e08b57ab1510b49
zaa2bf982be6050d2119a7691feecf9c2cb4f281852c8dff8b84d9664665be298481c31f3817bd2
z2f58dcdbddeca2327939960a24b12ca5e769daf00802bd72e519a40a5a9cb6986bad95f4a9abfe
z71f5091ef24c01d64332c1f079289f8229010f18cff7625842df7ac9170ee9f184d853b175e9dc
z6d1cf09122052dcc784d6dec030b04494dab416a4d0d598dfb58dfd5977bdeeeb7204efd004964
z3c979d0ae58591d3a8f6c2e563e8e8aa08e176b5fd775aaf9139db875c01aef43f2366aa8d7ef9
z852a803dffa29095de31064050e98d59abb7c908dc2c00cd1eb9460da777b2ea96e411c4716aca
z74a7a49137ad41150ca86020561fa7c8f2bd176d98bd9eda28f3857116563f9e09863ae7906beb
z46a879e48e402166499ee616afe5bbe8f3311383c64d3ca6b72ad21f7cb1ae1f7166423aac24fe
zf912062d7d8512c83ca1c94449c1bf477b99399b049c6978cfdbe1606d5b6516e6183555dc3c4e
zda3cb9df708498d4edd07256ca875efba654e90119dd09bd372a7eeeae3fe9b41da886178fcbe3
z4d80cedc4fe7dc4d8264389becd8757b83e78e3bd30903eaf02247f6dd7a8533327f458869c45f
z750622f91d4f87f7cbd5d61eaeda0eb1506d00410c17c83aadf504c77cc903af508e39dd7ffb3b
zcc6034b773af5e74cf002af5fb5a6f1f0b26f56910d1aea829f5937fb502b76664cb96e3410d53
zaae5d9d97abb35e8cef986b031a85afc162246734be1a3ac78bad3996113d56c725dcb98626c89
za4b7219dbd8666e88daf819eb394c5cf175c1259b073d3d8d4561156edcf68e46c5a65ccab0c7c
zbed449f4f83675002db2884ccb9ae5f6e91c6e1de121473e90d46543169331cbbefc1d0bb61988
zf19c62aa809e7cb52fa67984c504dc1c3e18792e80d168b4b92c26abca6ac7f0a44b85719a7f76
z2e710f6c95074f406916694c452458068df91566a86566b3930b4ad76a0b2a1ca6268f05d4e23a
zdf72f5b56d327a57d99a31a2511371712c05cf33134ff1c82ebf91ea9a02b8243e2a543f046e21
z33b133302f0c6118dc3aee8e2d1725ceabd1f1873d993e36058b1044555694cff52e95cb8242d4
z75a0055dc57dda4c279c1eb352c2a2172571cfd54beda030f1ec74d3639c7afcebd66771c8bb18
z43977b3cb59e7cae6b8e4ba14739f30f340daf3ab3041b8bc51651b3ef77c3e44aedbc17e3ea88
zf86ce80d50f815ec89ab73f3d89caa447c1e4139d908884f4e5806a2f1e42b36d6e737fac408d1
za5ca7f7176f55df1ebf751a16281fc7f2613ea8d893b2b0587bfd2882681900bc1a8cec53fd071
z17268d783f7f644e818d7a33bcd6badc67146b181de7d82950aa69001105b577f739c741142f60
z0c8b79e00708fbc0fdd391c41e81d416ed7bdff527dec2198a5b595a87c6fbd555f226dc4313a3
zb0427cb52c07e030b4432d0b693b08251cb1b86a9eb6b7bb3ce29e8a87cc39ed12aca9d9bd1979
zf74c15f3623cc8239209cae11a6fa5b06a03575339cf875e4bfd42662a07e8134015dadcdfc702
z7a059f4b23c07ea8f8c6ab50bbc1a62a88d34b20a0e498ddd14a1969a11c5dacf8cb2ae193232e
z19c202337bf364833ab9a727ffcaf0c808e095e9db45003226674c1e8ab3f9b2e80fff465b3fd9
z882355ce6998e3f8a039c47d8be4c791522efcea1e7b50d70fe57eae5d1d258fd82abe72c7fe75
zcd8fdba3bde4e4db300c71ea7abac75bf0cd2230c26dc0ffbb483391e6edf2decb0d9dd289d4a9
z88ca836abd3016134b16c45f32fd1f471c21f2775a9189a2f3a6560d4c12bd397ea8ea342f9466
zd5d7d75d858c0d1036f735a11647489a590190c609b2d8fcd09ab112e558de22e9c60061e5f488
z6e66ae5d92c801181b3808d16045a6d8c1561a2a2be70552abc5725ab71d8e58a7c07d1d876852
zd248139282275da2b70ad8031413819c65fcf09ff94444b86ffd4ae0ae4346905e8d3601080bbc
zff199a3d8ddde6fd7219081a35da89bbc73684c6ea146531f9667aa0cf352f0a299fec888cf7fa
zb119062a638010ff9da952294f72c6faebffaf30abc21269a32e03b917f3a04adfc4b0a6c1861c
z4b44319865fd76cd58bf500325b24978e4c966be1706a0bfd5f8ff2c173b0840551341ef2a5711
ze0e67bf1a4f32dd5fc1adc198609629e090f51ba05a78f185fddde8ae5edda75bb6590534b8630
z53bb1e36f0b6098434c88a850fab4d8b10f21f66b6bebdcc3ee1e7d90273e57575163ff93baf11
zc2ba4047f7eae1a703111542c9743a84af7946373957aabebecc2ed97c7324d5e79517f2027c4a
z2709cc336f3183313dc5df7d143d6d5148467f335a25617ef4c89ddbf2d67dc0c494ab63196e8c
z9a749479754372b276144b75066338192cbaae46b6b7849300860a5494bc18d1177fa297668766
z80ee430d02299b3dd3b548fd9950458b65027e812e38a204ca91a71a590b9d3345c2d2e6b39952
z8146fcae3107493ae6f4d95bc174bbdddb4f4a7f88bac51eead70dbda82e4ea99b350b46627bb6
z9e6916e205bdb7c5f9026e5cb4f0efcefed1b612c2f4b61046be35b4a2cc7fcbe21861134e741a
z43ab91f0b52c8d3b3cbeb3e571561041adcf7ce81caa5f54acfb6d5b74f3ca4e652f98901b1140
zd66282bb5416da8f74885d63cbf0e9bad4fb568627264051d7ef4a51e4302bcfaeb0a8ee1b52e1
z22149f3565a6706e641320e296328ac41f4a6d890ea28abbe942adfe684da37868a1845ccd9967
ze1c7049276cc10aeb19f9c160498e1846eef10c3d778dadc11391819724e592e2db2cc274d3211
zb46c042642b7e985a5f074c3bfce6a8eaf1c6c93a8e22676a5eba64d235aed1b6454cccfc6359a
z55fbe4a2e6a0e52a6edcc3a2dc06d23b01d9ac06dfca093ced3d9337897165f7bf78ae78bd8642
zd06968d254714e24789a8aff78d252e6b3ff79830a3f56e5e760962f4f36506989758f5e6875bc
zc73ac4128a20986f1532cd7180600eea1bc780a2539138255f530e7175aacc0177b41e112f4f60
z4ab6ef7648ebfa6d806a9962cf07ff51409f4a4b3aaedf4c65aef5f2a7a28398b7592881efe182
z50780a8895e188bbbcf5eb5256d15bbb426f51fb8036f05aa1345a9a89b789f52ab38970c95c41
z5608ef0ab00027d1ff9c6b7c9f32697989d27f56e79a4fd782c51690cd13d3f8948ecda2e32af3
zcedf04a752814da966af4a311e5bdd23d4aaf4a66d15d5cbba247f2b21237e8950517bb3cf4868
za2c8ab39674872b2f82164c0a79edd7eb83d661378f72d78a47a03ecdb103a9fb8783114759d04
z22a09cb3580196e1efe681ac691ae8395f8ba67d0a782ca51ed6deb04810a8a503aa4615057961
z8c3f974e8c68968508da8b00de56604309129397f088ecb7c9b5b4e100f2669e2dd4597ca57131
z81adc8ac9b0f219ed5583a16fa17293b9327fce23033104f51e6d0872b68b4d4af7997de49a5fb
zf5b2cfb4c6d74669dd5a293cc848b48ad890057f0db6f415d5e8f876712d06d876fa375e633265
z3e26eb723dd27b48db8069d7e2b9345f33285638d32c319e59f883fe2bef85d054398933fd5db0
z35270484cbe9790a43c31686aea9be9a4379c59cd69cdd177506d7569d0af3dd4f7a41fcff4bd8
z97a5d0fcfd525b67923444862e84ae12603a5cb95bd9f2705eaa584c7ebfb19bf52272deed0679
z3fa56c4c78f03b250482988a3f77dfee4e0ffb2e6e2e2bdd9afbb4951c64a2c2393d701651a51f
zabc7ec18ea9a968bd79380bf176561ff282e2d96f472a90196d36ebd77574a6cfa60c6b40d38f4
z247ff4760f0e397f50cc262777cc28ca50440a1c112f4a9381c2fb82c99885b8631367158fd66c
z2b7b8c4ba1beb9e06c88e8e392f13e00877f9b00d29f6cbeb055a9f8e0b29371b5943cfd018a82
zcf729c30b369bb20cea153a513a5ac18486fb42223a4b416b2a7c98a87f17920ac5bde3aca7d9d
z1a3957ca98728d2d95d71af396fe264a34df4c9b7d1216a89c477aa2bf4d9dbfa5704d2bea32c3
z7fb6799e343fa6fcb8d850f9ee224ca11d53084605d4c61232da30512590bb99fcb7ba67014c6b
z954797cd9e619af45f13554f00e077cd318a06130c12b417bf6b55d4ae84a8c3bfe7780219e568
z60587a960424c063259c8faef173062e4e558ef2d79fef73b36e3b7bbf3a74bde6c9df3051a141
z9009d3643dac2689a1dacd6a884f191aeb944bee2d5c458eff4151be2ef473dc6af9bf0d85d243
z7bb1b9afd3682237e87f1b0c6d15d6148a6dba79b236c8ea4f538ab05d513c4d727605882cd3f1
zd36988baadf2ab5d9c7e325cba7605d49c04972efd9ee0ab64e3874bd028d653ae368627c7ee6a
zbb8633f3dec2fb98aa8f905cc2e316fb81acc03c027c2af5b356d15411cf0025f4d4545f2bab6b
z7ec6bdb8b6ed97b20405ddcd0de6d32185767bf8b9a0db19f6dfdead3e54f098c77bbab8426a16
zadba57041e4d00b0b7f2de2b04ba019451c0b80822660ee996003c2bcd535d7ec251576e98a38b
zcea0fc6101966b85effdf97cc2e6e7cedc2b29db047f961b9fa38b1a578507af7ca907b06b9198
zebe24e86e0e2be5eea5b95cbbf8f702bafa5b8bf4afd1ac62deae21feeef759c2aa4df0c70a3d7
z9d0eb0bc7f24066fc7aba0880e075c7ec7136e02a16ead50cafb998628546e54fad3956ab5dcbe
zae95b23af2ea7b813f0221d7e7e0d767410f9aa105b33bfd8a736a4b2b05f3deb0ac747575f92a
z0e6bd88d7321a6a915ec7863444fb7af4da9f2c654575cdbe7e6fe323431940afc91dc74faa352
ze26a1d357401940e0c504dd160c4c24479ef847b1107fdab5649cecf25c1d997b0f785168becf3
zaf342757b993bb52585d257c4999fc637eec8ccf9671e1f6ac5f50eb979e38883946dff225d07b
z48d51d753540b9f5d2c9f3d0a81eec8ba8954932155c6019e80e3836043af8f5ea4bd6a959a4b2
z2b53de4483c26db3fcd2cbab7f8f0beb16f7817b833b371782edcb1b7419ae05b5692dbad0def2
zc46e034d591a9ab944ecbf5d80c28ba1e0ba2aa788ec3c2a9b8295f2c42b886d6a6aefde32d691
ze84224090bc67df0d7a40b0079cd4bce8cbeb0cdb7d45226e6c85985ba48260639872c0fb309ce
zb4f2fe3b067ea6c5be1135a207882826f7c84251dfa9d6e120e8676ebe507a5d97d136ecc11f58
zcda6808923bd0fec8dc9a309c2a0fb2ad708c9658b1928fddd542d72d08cae8cc3df8465106fd0
zacb47681018af45e2e30c6cf1e7a1737d5a16a1710966d17c73087f594c3d6861aeb23cd297987
z4bfd7a25ed0e788f44126845e480594b3133d0d4e6d3f095d4c7928801060558735b3ea8149298
z98089eb89de5a848b55ae5d18aebbb00cd81d7899b3e07da6444e4e8b4ac720afa00bd10e0a886
z7eee8c488d3baa3831d8230669401f7ccba7d1cc59b2578e5e254a19fa56bb9828adb80f917869
z3895b41aaa8a370ed48a48d922b6144334617718ea4c7273294aed798ecf9cda6e70a76b39395f
z91cf66724614f765694f1d77581a782456a26d45ff2a18dcc22a48b592dddb79792efdf1a67b51
z5d17468e82b20a5d1d83ac41ee40380620a4eead4002712d1b3eaf7494d4e0321a7f295921a80c
zbc6bf0696419bfdf50a0f5209bfc19417a7802bde02bb6e2223dc4c2c14e661c9cf007eb04063c
zb768a40ef4bac221ac65dc03554a68edc4f1feb2a8253befa0e20f1fd4799acbac8fc4c687ea3e
zf13035dd217649c942ec1bd07ff84af2b5e9486d25c31db6a80c07125bac0c9904607555f8506e
z53704145a9317cbc8a81ea6e765cec8efca8f4d4d0c7946748d8f5d26a75683873d69c59e6646b
z2bffe1ff80403cf746f0447aa3007366c14cb0157e546461b660db84e578af38f1716df6ca69a3
zc4438d6d9249373743837819111dc0971449132b54ae294b00f9228ad504bca418eaabf3b3edc7
z8de25a8f7b3b1c06304369bb44bd36e7c777e3064054c84e591e0f8ec3a05440a894143287c512
z4eaa9f0d70cdb81e27951fa1cda602db60b7ead05b42ba07e5dce868ebca3979607911f70dc020
zec469a1bb384dc8c0fd9fb0ef1c43b547b6f437a80fcbb747f943bd995177e0b1f776fbabecfe6
z92e86128492ff2c3631f3988bbdbb9c62a5c9120351d705a614c1e2b1e6ac86e916069ae9565d4
z9294f5b163f9dec85e83a691b1247a1d407591e2857fee50ea11ba2d02ef5d2e87e1d81987028c
z2af702d368876237fc28408fb8535fb63ca66034251fae3c876427f1b4891f215dcdea5c8b8d08
z648131330d7a93d594cec2a3799d7396cf68e8b167df810a61d0a9e1513d00527026c9578935fd
z94b3a962aaa6086a5bfd738ca02ebfbe3e0f2b445110ef3001ae7484616b800d296a049c61d589
zd81a63013baffa4ff7c3b02bb48a34fb79efdf2c08dd05add4342830794b3f985816896cf2b395
z44c306e0b3dfc5778b4cb44524a30191965c90fa313c1b217dc01042a92f97551fde6b5290d7d0
z95dd197def2f9c0549a3f7e88cd2d639da106b0f0460ef20725686e849d3208dbce467d3eaa1b2
zde94bce7d3989600a4354ebcb73097b656d72db28fc3f2761268c83844175a7e62d7577b594500
za421af91af3335fba6608740eda271a58987089b32f47265db94a65d74d9b2168eb7e1ab16a3e9
zdeab2a5c78ad0cf8c5b879dafca9d42e2dc0178abba7576e087a6c2f6574f97c478d06673543e4
z3219e08403f96cef8949bdb2e4658fa2a2a398f40556c4c3afc42208620a2d4802fb8e6d811269
z0ebcceb94d436cef8d0b78259d41b00425fe01bce2fa75a36f6b6bf711439927585364260edeff
zccd8d3de7d83f224dd6421e3c8c311b448a22d91a602c46f86bee3c071bb757a39f8b74ae12cab
z41bdedf77a7fd38f789bfedb7bb95f5d4d0ff0a6068ad77de2d6e351185c19f551eddaa949178e
z8f6e13904ee1030d66f7d30a6570cb5f4a367e0dfd248cdb18ff8473abc18c1d34e5efb49f18b0
z3ee855552e854eb5d3552c86453a832dd5f3201d0c180b13200b51b8001b6c9b8ac33519318e8e
z7f80f3726f44f3ab07db2fc36ed47e037b05305f81eecb007acf4d64e3acb9e5283b2b397d7bb7
z5c71d49071d44381119b7c4792683a289f9a6dac3619702ddb6a3985a53227e07ac013a7080e19
z652f3010e673809faeb0336e8f347318db7266fb9f6d27e1e04f576b6fbbd65aa895a469da89ee
z5cfa1affd5ff6c55a629e3f416f5ee6a1a608a7a3fcfb17960b41d22daac3e74161a48d27a0298
za8fba0e86991eaf79d3481e941c043ee0319b1632357f4eda88f671a06ee926d699e4dbe71dcb3
z1fad9c5f4fbd384a7b5950d0636dbe6609fe349e85e3bf4d69a410f6e00fb4603501091d4e1a7f
z8c305c5c04919c369f48c3777b93a83dba993923979910b05ba8ebe30f1e368274064d6643e408
zefdf963bc435101da5725752b4b2459bd743178b1c05b2d91411fd88162f516bd7911ac37a8a62
z08b8da7304b6361bb0ab5c13ecec4c911994b3b94e875ec71febcee40740aa666451240d0eec8a
z37d1c38040f40cc04a17485e05806f29fa9150d5a4797f2b98056eeb07bb6381df7c61a5613451
zc7b1237076aa618c3777d9c7b1d90ea65fd49ca44df23883c357d69d603bccaaf0ee17e02c121c
zcdba0d2242d3e75498459c6c073e657390c5756d3fec9ba68f745e10f3fcc19542290bf09568af
z6c281db6704a00674c7c3d1b728ccfa952c97ec0596e44e1002cd0519b3e64b8f0bcf970035ab1
zf05374042972df8c9602dc42222b4359f307fb71a5ba105ff738a817185265ce1456a14e5f3c29
z44d6b3c6869f95e612e57ae9896e31584c402245113b74c960bacb16fc746d6806fc5115272ab4
zb80970d66caf6e76bb33f69cb30a4765a64678fd72b017c23d6edccf092925311e1a79b7dd660c
zb75b649721e7e39e5a5dd966821ec712ccf95e5ed4b2c1573c889e6bee89209b30157769453645
z4b55e2af49e8f23f15460319d7520779fe7c14cc0c43901bb7dc9173bc363d86e06ff736eb9560
z548d1a07fd6b6fa14c89c0d138defe7c583f50b868540029ae395af896621d3f82077c01de0ab2
zcb875f9018a4a867979a8d7eb3be97a1bea4ee29cb5f2da17b186395d68632c49e51124734e1a9
z3b53fdbf13b9a110015096cfa806e25b3ef851da64e1010f733746d7113adf9a313952da4c2ffd
zd9415135c661bbf34cae875053db2ca4d1eafce657cff89927a590b658b55039d8b5082a194200
zb8457c01612000eae203bd7648e8f89187eef033eadd6c3056c1615d4dc63197fc314c8edfc8d7
za6310f220b482800d818f36ea4d8270ae060d8795ba969bc362947d12fec6f7caeb5e97259ebe3
z1cfa0ab6ed6a6cbfa31a279f3dbd65f2788fc46a1fe57e9bf1a19f27669460cdef3cf891bb0c3b
z62e9493b23a6d27068c6c05fc1b3531ce328c384b45b63a03bd90b2a8f8f16a7b9fdae1deb9a46
z12757dc420f5237260533e0e9ebcb3f3b94d7a6fd3f96299bd0fe418b3e71c894d25435374e49b
z68dfdd6e2edf3a4d651f7add7ce3cfb78d00471e70d94053619f8281d124f1a5bbe6d7156b003c
zd7222b57f92bc7607f7842aea4b91ba7c448e1fad19f3d09563523d9db1b7534c78686f55e02b5
zcad70a13e6d7054992d5c5991443acf304e211a6a668b468c86fd30d708c1b2613faee51ca1037
za45940c870596b44af8518211325c145cf6c3498eccdb8cd94baf0694639e7eebd6339725ac7e4
z78309b86df86180c274c9b2ae704db2c99b6689516d4399c7e605cc7f35bba0460a283af2e9582
z62b776b7c657b4a25c810ac76ddb30c0a15d67aec54fac393b4236bb22c67af230aaf4a35fbeb6
zbcadd937c4e128f73c67b6850dfb89e86567a031c543f49efa3de1e9596267fe0a97ee7b9ed605
zf5ae2307ebb6549a657b5f22bf0048c344c47544582f4c6f87ff06878acc43a8427a45369d91d4
ze68df040b8adf8f5336b68e72560b3da54506b204d3910dddb31e2d12442d6a748d2a9374fbafb
zbd61e070ea098a71ee2c49b0078e2c8376c8593e509266ab396fe6193cfde424d5884075cd5e05
zf4c9f0223ba826f9ded23835af7fbc3d0fab6977e51881e9b49e7197304ad1cbe2538ed8ad9409
z676574916245c0548b1ec3ccb5f25c67d3c444f646a419326a205515f8b5760b7963611499f2c6
z6139648615be8f068b97dc65bc6c54506a2aa29b886b6b5c2114b03e4871c2d62660355ca335fc
z7f137c32760b46c6668e9ccbc070462563ec0df5360b49c01fb31ac54766d6ce89c064b323b463
za2eea2040317cc37568aeebec77c8ec57114d1e8d78156f95505f896bb09b2f5d71fdf5ed866e9
z1bc4931d1c39853715e0dfb76a59442fa570a53d4deabd26f6d10466954e8c9cd05b7d46c74da5
zb9dfedd319ec9090a797ecae95c87ab025386894f5e1b3e4b237cc226f96e1fc5b045844328b07
z5ef09b9740b62b9383acbcb9ecc9f3b45d72b4fb62c67776f9479215a672aa7ad29f9fe653e983
z9ee71b28ee264014ef827a3b568d4fac68c43f9c2a2c2511bf6be04bbbb464ea139e2d5564c65c
zfc19171b3fa8295f4c6e2873ba6eec32c6e57308e0c27f284e7cd57fa48053cf1ddd4cfc263be6
z857f7c873fa8b55ecd725fa4cc37163f9219e202083e94e87f6e5cb4a604fa2a453d6c45ef554a
zae8cc0ada6f7ebfce2d0c511376199d3ae47248ba9174b34c24ab557e7afdaf3e3267b07f607d6
za6617d1f0c629741ae077029d4f04406aa4764d93ab48606c702706471bb237a8485d3db9a1991
z8ba94711653d32c242b33545689f0a86e49a8f54b8127a168632c34294730b454fc64924621126
z892a82cac674b408cb30b8ae4c76552efd99c3bae21479a3c71fe28517fc9097f730c7eb5b1c81
z045be9d005b53be5226d6fc79e69c85e5aa8c8831cf2e1a955adbc56dd79fd3d614cc8e4eb36e2
zaa81caeeb5e7b3600ba5b512562e0331a96482050c65d143130c0b562c06d20f5010d14ca08f3b
z7355c2c05a6d367bedd7f53b2997d93afa82c2103a4c67439d1dbe318cb851790a6a555926bc85
z0c7ad00c2da14b0ac2aad4c443a69158da8d4ccca5756152eae79f9b770d54d2eef732f55a3759
z4721d3d5e79e65c2232e026141e109b642e7f69b8f22188546467805e9350a5eb13c897f9f40cc
z077acaaa40e2af1180ddad51f8eadb215b01814224855b58d3e92c0c241b075b0e79dc9c2ca0af
zedbf4d90f8b3270b84f1dfd31749fe38444c9def7ea203aab3f166e10d0ff4581dc7fbe6aafd17
z61cbf4fee1018a504778e52fb408aaeb148d0fd31860d740d935c1564b592cf43b5c8ab5fcd9ed
zcf204e0db1c9b069f88cf0d546eb9784fb1b90749d34acc3370a98e1190138cf6de9aaf9e891cf
z8fd3ab51e5eb076999d5fa3d92abd2aad47364e01b16fdf77c3c18f0346e9de6a88a02171e0243
z3cf0ade22a1fdc3e4dd632f535fed168e99f85182fd89cb836797c2da56d17d2eb77c44e39967f
zd2a29295ecc27bdce83e912fa424ecb7d7620d68c86a3f83f24896ef47fab1df21d24309c0a745
z9c7ed35a160831044a8169c6d61be51a48922b524aa701018d6d8a1c901ba5c5cec720a9715c81
zc804ba2625717ce9b1bf85e6b451d66aa7b79680ba213188833a2618d49a400e484bd56551c410
z3beead6dd8a2e5301f13f19e3d84a3e262d8c90dbc751c8e1ef85ad49920c71e0f57023cfeba5c
zfb43dcab4f23e18cc5c7098b6c95a4101d9bb38504b8ca7a7c0c9a399cdd7902a9341e07f191d0
z47920312f8ae4100d5893f5048f94cf301a6bb87666f1b58c814bd8016535522e55d3b88195008
zc73c00b1a4666df22f405f8084b9982dd9134f9e39e260d5de7e6a71cfc5f03ebd59e96cfd4fe0
z79c2d522c2c29fd6bda2966a0ce3029ae67893806ba617da17ae48b9be07d005a96a610ab0f677
z55be917f6f787b278f784ad527c172805705b3ad7c9a1ab2c9741741d542e9d0f3bd45bceb744c
ze11eaf8b0b7223ad7323caa568c97b06a042fa5b037b1195ad41de8be288dd6ca254db87012ad0
zecdfeab054c9cce479ea2391264f0c120c2330a66e6d1277095932a16c2312b71f8d267aa5a9e8
z4450ad9daf31126550db4a66ed5dac2634471b2d927d93f6821cb353fb426e1b56be068f32e62c
zac4eac8a403d47e891864c8560a5d21ca428b3cf373d0df2cdfdd9dcfc615575980bbb8283095b
zb5020ef17c30980b7b90f4e43db3bd13414f4fa6c687bc1c84103615d786f535fd95eb6ff076f1
z773c87545eb5020b22c9b1d981d02af9105aa43c3ba7429d956c1eb80a543a073dab48cfbab57d
z73a0e43be8eb43c31180586fc837e0a147bd2c558a59df963daedd886d7bbc98cc42e7dcc45cdf
z0cec6c70c679a97672abe79923e8ce4314dabb3f685cd204c95a4dc303b97bb3d587edf78d8567
zfdc7ccd353f43fbe05d66c27d6eb9e10450cf7cc5f8829e35f4b2ecdf7394dc7ae61c36bc870c9
z471491bc6a33dc2d9b751dd3b0968a275b7dce3bb81f94170363b8af4dee5f5ba5009c4df28a8e
z3c557c300219772a276a8722afb7031d3bfbfd88b1f5292adb755835730005535f1286e40048bb
z83f9d16907a82ade0ab16224e73f62d1d92cedbb4b227790ef6f32cfef754f8567d773b6b201a3
z6dd28cb0bfdfd4a37d31d24556232619ec326d1f3c6c236cd852d24122e2b585cd35ed9b90f31e
zee17eb7514ae33978a40c8c3880e28c2b5952d21c987e8e7ba5cdd60fa01defb20c05ba5c77144
ze1055d85c5453afe5c00857934f01c1c28e6809d41a35c39a69f011ca44a74e08350a0235f3fec
z61de0c2032a81cff6029f24cae7b3746b9f20c59cae020b63c4e1cac7b75c54ba726e532b0e96b
zcb55130b5fbc28b56e9e32a1f3acdf7dd962d388777b05fefeb1ab021e64a022e5535406f276b8
z7aabe54828516ed15345870d82bf84563af262c8bd5699d7a8bb49f9360a947df84e89f80f31e9
z8efa5d54cf36ca2892ec8766d0eb1344969b3cdcd593787dc7f0e50452e9ae016ac014a9981eb3
z8ba22403e7ea7362293eefb882868072ce306327d8957b18018647ec5704622074f137821a81a9
z24a9eda683ade488e231c48866dc527e145070adbcb66c74312a34550ec87ab28db1abf5e76f9b
z56e043d1216d58070e7bfa567715f60d222cb81fca3cd1a3f3247838aa892cbd0edfbdd80d3f3f
z71568426e81fb5d5d42faf261efc0a8bd728489d01b61227c27d137c70668169906ce4fd5fef8a
z8ec95057e2ca3d65f0a50a5b6cc7a65ced050b04e54bef79b0e07a2380a4160c6b5e11acc24a96
z7d14b930c57ed25f8b893e49d935a5710480db9754ffe4054bd2c63fb40f66b480f3ceaf4e3237
z67cacd42bca01bbb7b4eeb601ff2e5bb920ef36079bee19d1e951a662e0524d5ece2904120e3a0
zcc038d12cfcbc764ca8d17cadbe46d95ab5a899d1102440332536a46bbfa723732508feb966a78
zce1c42d3ec6f8f8795fc5db218cde82cf85337bff2a37fa28a33e1e4da400a5d94e4916a5371f4
z39d38886d42bd089a19d05811353d6848431212c038dc782fbd15dca79c0f76ff5d734993bfed4
z77f11aeb4e27455f42288fb5f6fefa46dc77a80191607abdc159deafa5c1c2913451e8d8986c5c
z80775790aaa5f33bacc97e566281597a74902f8e981dea361d8c6e8e75b746e3a78f9e012504eb
z63311497defeb4c228f60bfcd39cbbf8dedb851a8eb86552d28888628f58437a09c741a8516918
zb2db808ad047b89e09faa421ac3eeac85d8bba61d6855458cb7fb5aab781bb4a5df3547845cd8d
z2395234ddec15141664487ccdcc78ab01af1d1240bad077af5f61f6e5c5c13197367fb79a724ed
zc09c94dcb0416027aa1a85c37aadb4691fcd07f3836ff2d544833d128bc472835b42166ac1a960
zbcbf0a817fa507865a2daaa57b53846c14648e01ab79dcc3646622d2e07d75bf32d90faafb8799
zcc76cc272f310edc3b32693f4609235e70aa7a6c356515e324907f7f04e333111e51a4825e9112
zeb7a721a18837d81296b7e4bc54b6f62ca9ad8737b6f1dc4c4b03adaef7e99baa2421983cb9e6e
z2bc1c7a6e5c74f23c90e69c84be1bc1075db0392c56b62d5e4e1184f57b10d7eb112db1e7c6747
zf4d51516dd26d92b01bf3d398484f74b491e6ac0744c8a2d9c017320a6a7c5e0d2bbb74ba86a58
zd212aa0841927bd5a740ea52732317e590b63c44be3b4a11e146e1a4d3ff05f513defc9da63ec2
z2d9310bef2f4929ecc1082399151953a2aa19197012654a01fd76ea03755380c2a009105928360
za7d7b2dcda5efce488b927b74fe6d9e10560e7abaf33d2631d3155fc8c6cc8beaa41f682a9bbaa
z7517e54e9dd2c00a68e29dfa71fd408aecd77484af238ab9584c0f599d2ec13322248d9724ceb8
zea3eb2b2ce89fdebf9f60486a5c06900879980326a599d5d9753991b2457021ca0d95913b6ca19
z7a768f2b48688420e08308608627b677a1adf1a01c439db65675b87c2185f6208a9709cb53e930
z46ccdb53b776e04196f9017c4c88053a49acfebd3fe6ad3ee39278a0c6448b608b137459b702d9
za0df67c08f3344b86e1d63f1a58e2b3d416bfed858939c3d3bab8da8562a9f66e7ffbc46e2286f
zf931da7d432265df1aec8ffbaad9dc12af2f1dc8ad81ce6cbc3d9e22a6ab6dd13162cfe0d660a4
z08f157b358519604600e202e0630a56c9908b916081636b92d572506c2236236b9846f36471231
z2a4a7f81961addd8059fb961245c0c294d25e9ef86047dd62061e9747badbfbb6860cffd682368
z6ae83230c593ac7adf16b3fdb52a9660bcdcbaa61c747d3bf33a2a6c05e7d880225b39b3de17e5
z1b3bd1a95e9b1c8620017ead580b31d145b3a006c20940dd5af60a5175547722c3a204b94e75a1
z30ef50d811770d561f67569f103a39cfc75b52fe412bbcc4782fc204c68a07b246ba73e27b0354
z26465f913a8d97eda7cad6ff5acf209c86d3aedcf5a07e0875148eea244ea95b6b14993ddf6247
z18e0487e40a1850ae74804d1624adca3b655b164609b8b682b8ddec5813f27785e0580f8b0e8f5
z4cbc380ea7fa9f96557d671094db38c2ffb4ebd121f0be264c6e02ad3aadc2f001e745808b0b54
z2840f533f29929bb040d63b87ac574d58c22d5ccb521aa7ba5f25bd459b58b0c19c6264d9d162c
za31dd026a72b70e1aa120017cbf39476453e21e5c8d0d7d6d396822e4a54fdcb52ed12b042f6d5
z25713877dc7a860bdea8886d831a0a02c0efa2c8c1a63a4bc3b8d76fb9ced97a66c310e6992db6
z9303bfe2b702fb9b0ba0cfebd10c813a31c1b53b401aa999faf500da30c61412e78f19fcd849db
z403577f8a076e1a779753cc909dcb4d672d0b0b3f0edc89cacaa5778eeaa1149f1a3c849be7e0b
z10f5fe4c1eed322f089959e6967c33eb411521b83a8834d070df32cd9204989ce6be7166a70ae3
z1c11d2ba483a808bd50d5c6a3595d2a9fe3d60f42a939d0f87c5596eaf7608ebaacc1ff2bdbc0a
zb9ced6c785096b13dd2a7e9dca7fa8666c38a02ab047a92c6c5d6d1f349c85c5da654075bba9a3
z553e45ebfca0b93f0580e21e19eb851a146395388459d125b8d7c7727bc5bfe0d93104132c3e0e
z15d4f6180f511d62f7f0eec4fa87ad881e3ad91c2514179b9b567c0ff419ff6ac51366bdd5136d
zb6d9759c6778dcc7f3d85f47db928edae3df90600dfd5479f4bd37f5e5a6ec4fcea63bab4019aa
z4d3f0512a1b66d7ff5f9a7c7788691f9f3ac2ed75404fd647bbc94d194b7a71d3e25cbbd755640
z4706037f0be61431cbedd8a636a5a02e28122b7a34f7f02c3551bfbf346952661eb3503ad1d85f
z9049d39f44cd7f28efc4613ca991c16ce82b7b16f7769992816b525b5298ce7d9a682088ed7f9f
zb9f5c81be38feb462c9fd745c3d21146fe7cf2e93d5898f980aa54568413dfdfff2cf1eae77fa2
z1336b6c41c3b378cb6ddd8983ccabb5972daa246e3ed66eaa9ff830e9f033dd9082154c61959e4
z85963996bc23f393dfd554258c5618f74d7bc7e61274a0f89a1f376ab7f8e521ee2b782d233388
z1f560506ba02e53d6bbbef9dbb60019c9865afb8f34d4fd43cca7ead89ea9c25aa52d8b767408e
z3d9d06df48f15f3a0e7fabed4e9b4206d42bf516261b1904e93b152d67e698fe999d2df12cb37f
zc60790c1da972b93c395ac6d9715c23ae7a40114b0260548c08a41537776ee19d34b4e19ec2b24
z97dff46a46112d198ea414967e2f5e5af7db48f0846fb806f020e643f7d1902fa2d5cec6497636
z589d86a3f4c712972a094f1837b3771befb017beb96238bb1d9efe16cd6644eb2abe5d9331ca2e
z47a4a397f4a1f9fac70f204cc26b0047ee52775c6e3b5c7631723abccd2a0a367d544930b5128f
z32d6e8b27c2fcf13b0ce568870cf8e536bdd8466b99ad7349e0b6cdb4dd5c4e8404df1c7940de9
z21c4985449de1c033c5177f16a564cb1f5185430d2e3b33b518596a086412c883c4775515c9314
zf54af084f9efc9618b573827c572db7c8d632c82e0461243109c57f77cbed4965aa35d2b553cad
z27ff518de176d22cc4fcc13b91cde50a5ee0d18e482a91246d0453652c30a0cc38bf1f9cfa6a0a
z026c0591b3d918ac0f7ba588ceaf79c010461e54f56e0679d1c6f2dce31db1cc65375e91f6ceb9
zd9c20d47f3cc8536213eb07e6cb845d42157ae9deb08bafca5492995a57150bcb4e62a2d3eaf3b
z5f27cd4286af270caf92ea616f555928daedca0f3e879e7fe79e441c0641a069fb564837ae5798
z044763d7321e4990dd2d429748375768c14e23bf8ea6ff77a50ddf527ff39418edc50712911660
zb8e9465c1853327c6e9c4f516175fa240e4ead8db41c1d73fb9a792e0d662fd35817f90c9b7833
z2918170344bd41e248ce5ef6924fca0f47716e0f53dd554aa6942fd633929581ecbc3a93998c66
z81f2cdc01021a17f4799f6d66e7f22a0cf5f7737d5cf4ab69b98c9e5eaea2c1f77f581f778bbb2
z4fa4f5890ab35685373f2f7b4d427488930525c24fd39dd1f30f14ecc438f44ab3da64d1f25510
z1d3594f4e00a9245b8f5854416f823676f08758b180fc2bf273e1f7c06e1db6ab2c1a76ebe0ba7
z30e853bf3f8753fd67782a8182e4138a8aa30d52d362dd417706c790a8b45cc32c80495e4b8088
z4fad3f0e71984c5699d51695cbf10daa1b4f46ae9cf3c07d511add1904a9405af5508b53565670
z144c1d1d408d30ba4423d08e28884c6ad0ae6080fa5f22f4c7b7e3f6bb47393f19b6e396a43d76
z38e814cbd5e7b97e247c6589fe8e8aaf299ab764c341a59b0a97d960eb371f676031b318d0787b
zef9ee3aafe6b3020c6cb952db65ffb348e5859c43740b9fcd90b892b24f1b079e663f1e27fd76c
z479f630b1cd0262c69b46511c11b4d8727ff0d292e0e4ff701207169615d82b70c831e813de46f
z95fa02d845f9ec39da8e8dbb45024d98e7873697454d3f0e839697b4bc220d5e8f7ab430606aae
z39b72a0d72ce20564389b9068821fb6ec9e7483ab6112c80509166391b84e25bf56bbaa7ae1e49
zc28e134038291d498ca93c91f31090b876a935dc81e8a5df3711df420b2808889eb4d166474837
zeee449d3b79734eab848e472b49f8fe9730addbcabb20fbec63d4a16d7af7c3ef58622ff55a78b
zf65ecf162f0fde5e5b7b88b064b8cdef7ba155664e173e897162a25575899c9efc704e9be3060b
z95043addbcaed2411e881016e5190b7f284ab81b25e9408a8facec198fd5de4ed37ccc06b5eaa3
zd40e0f4622801ad499187e392a6b04a2f2e9b73e5a8f4ff15b88fde83c961c2079952fdebcf6c7
z27fa6824d9235a6cfb2d92e6b2ca391ad9f7529fd33b511127d1e73230944421e81561fded44d2
zf799073f2985d7d1443ebcdaa8993bbc21f4514550adf2321b60bdba0c9652d70f8c7dc36469cc
z1583ad22316e1c1be0125998fb24ddf56b177dc0f007b7445c6b9b9775ef6b1284ea518c2bf862
z0f4db445aa8b60f936d1000e3bb51a8c2403651ae08706462acdf5fd86a7e0ee67bd23f305a044
z9ae5779d110e8e6d9b1df4efea88103684f857f73e59e5653445f7b6530a4ad05fa5a10c9ad0c5
z676d87e781fdb4c1fb4ca01d244547e656a286c66b27ec4625f13195f61116280c11923322071e
zfab0ff2437293d7dec6bf664da8c1f2bd7550ac9ee5fc52b7cd9898ad65cc6cfebf3a22b7549af
z8df1a15e02749da56fa2e1e4d74be12002e715a99a94f1cb49ce0a36e2710a56914cd15681c908
z8cb5c4b5f5d5e58ff6c391434095dc3c76069ba44de2b1b612767cee06100683c71669224bc27a
zac4d0d8ebfc90f0204e5f64c06af599b56d8563c766248f729147baf0df881af04b4735d302ef4
za455499889f9ae1084bf8ab8176c75c164726343e9ca27dd358de40d0f80dc8fafcd3fadd76cb3
zd454e7a9d9adcb089389e640b838424a20ba66f8a981fc016820c31b6072fbfee721a45de9b2f4
ze4142bd37eee96fc0d280024cfaa992bef8cd7722fab77320ec049226a12f6f4cbe4d8ca3844b2
zb63d7c159b3e6b20f0a97a2c1b61fe51233f3c3e5ea8032cace97491ba53e5647f57f2b7efee07
z03f583ece068133e8d7fc8134ffb2395e4d7427c7afa78e9e6c269433fb30616c2e6a7ecac68d3
za3cb0be68f641703f7c5053314b96d1593336f6a544546f758dba21046f3a09642f8585434d6bd
z00f38791fefc9417239f17bc3206f1a835900d92681d45db644398d80ec55873cc1962ccd8248a
z05a152cf90d33a40b29e44c42f555154751c067ede66c5c65cdae41e0351ee3b5e15860be7556c
z887f50cc71d920dfa76b8c4361523efb8497e718d98044671de66aefebd38c035a07529ef6cfa8
z4a59564822aa74da5890e770565a45cfc8fd38e8bf3ad4c15ae9d1dcffca3ca06ec650d83e4e6f
zf7bcfd49aaa4fa6437b9be4dad4d005af4612695eb6674be796be8751f8b977fd9a559e6425472
z202c92d288a8f395359571f2d4a7c9a61a1985767a729f05b8f2abb4a3ce515754f2f852e7ad93
z17c66c05b69b79c2e650d5a4a2919f0bcf9b6d05020f8d1343853eccdeb2dcba8bddd820d503ab
z977b6ea2cf4293988dacd8bf64c416191f27b11226d67535b9c0756de376d67bff52226fc3a3c1
zed0309fa183e4ac591a62e0bcfeb3c35ce7c38cdd069cb6af0052d81bd5892ea4b3aabad85d067
ze1be1ebbfb77a30ced1f41a53a7b7d22655e631dfd8f3195729e842dd7f61a0230a9b6a023f67d
zaf8c4dd70cd8ebd20154c6ed8d115e67d1b9686c2bac9a3f5984cdd790945b4e8203d2545bf2ee
zd617239c574bafc923ed27a5ac2974d94d5791bd0dd31658433df945b73e3f08292c93137c3f5e
zb40f6d6990671ef5d701c9e396ca9ab69bb7c3bbe89fd5bda0d194d6719567f7494e8ccd82597a
zd1c695924f01e8cb7b0c02ae4c6f21637581b2ef21f3919593d561dabeeba897b3ec04c8e1c954
z6e5665b23105c6559b09549083a2420a7bdcf5c8739b51ff2ccafac46f25db24ae958c38f9a2a2
z874398e381f569c71ff34b6bb03ed2f658e2874fa818fefc702b73ff32b2fae785c86845c96295
zf741fdf140000d3020505a7941f201b937db06c756408810619fdbbf435a299d312111893ada47
z32bafcce1e4adff618d8c939e57dc6fd4b435ac226f0c022145923bda0f99271ce892bdfbc09ce
zdac425666be70ec91a63ae90254c21cfa9fe12d75057c7c9173ebc4723f55918134b7f38622ee4
z6bae839c77be944c0d1694342bc7220d55e1cac8c311054801dbac01d9fe79c163152b4a29df64
za51f75de9b4b7c9b3c63d285e3f7c6ec040a631f2797b5b9453c2c711ae350762b523a9edc7d8a
z2617ee9ba17dd213989f984376abde0d6e87e007ca1432418a8dfeb212b7b1e6809e23a00d7eb1
z535eea00f1c382c11f38d0b41947d4c27a5c1c46415b2800216a3c3c7023d91a2fa4ed9026f9cc
z5038ad4ab435f7d37cce1f4e3e3662aecd6b2e65f643135b853f6689cac83acf08abc8ece7516d
z9099e308f1a25bb5731de200a396ef591d4d0c7ec7e15c2b5f3fb3ae5e09206794913f8b37d0eb
z3c2278b6695ae5de4ffbf3c52b4c7d1e363e633c1fd80d58021dcab21a6af0196f9167bc0b4dcc
zef65f906ffbd748350875df82f41ed41d46ceaa29d00d4a799b25d45cf48993dab6519bd1c4599
z384d2b2c0a15d2f7359bab3067899496f6d747d40e64ed9a200ea12d98b31fa9b254fd7b9dde88
z5f773d877f2876c0432a7eaca047e2ff67ac7b0417aa6f201816f52d65e4e68dcbb0ca2c361888
z172b33cc83addc9261ad2d42e5191e8c61f3574ff39df42c0d09d68d96d405b868dc35045418cb
z5195f82c6d880cb9fdcb4095566fc4c7f3aa77b75087f7a19c0b499c2db21d50dfb895d703a69e
za6b75cfe700935deb8d20d43043f4931e985a4f2bda104277835e0e5fc3c652208a8e817e1adc9
zdfafde03305ff4ddd932974f1170dc848784a9620d82da38d5c70c8d6325e6d52454f3968f84a0
zdc15854126f555659e50d456ca0c6291cb3a178c97de9a9a7f8b8bd90d6294f72a2221846cec59
z501839b91b4f6738dc483d445a347d15cd8168ff8fb6819b9f7c207f5188bebd8569dc1647705f
ze045b6a50717aabd752118c8bb5b15861a68a69fac0f112d7ab549d963559288136533c4af3820
z07d028316b7944791377225fd389deea904d8dbe059f48bf7f30bde0a3f0cd1ea8281f3d1b8867
z206ced22a222adc6f5dbfe341ad95ab9edacc869f861f2d0636901fd5f51a400fe8407cd5664e3
z47b18825ce85809a68c0db53e85f68f55d235b5e65e43d1d1bb3994615f74131e738f769fe70b9
zf6bc937348f469ae38c5b9bf0792503c9d39234ff3a809a102a8ebfbdd002cdc4b7923e8748382
z702c81d93fe1820dbb215274afb9a7a5afbb6d9223ae148250c6d0fd7e3bb377d52a8f24211c1e
z2d2969529d69dbbc6258bc45d81afe6b184b4ffd3899b6aa57787b490daa3a17b97297001411c9
z6010d241d2bb695f48021391ed6909ca397a18acba4a2699c7b78f5726d4d514dcf0cf100b5951
zf48446f0a9a94a9cbdfbbe43c35d60f70acb93e002a2b504a4e46df6b86af3c74ce0c75c46659a
z47f08741adb77ee696f522fc6daa9ef4f08cced0419cbdb7606e0e32af4eab376300d1a86cef50
z76816cf434c5ec4a674cc1a4f6ec61807a4f7d0df533f1dc66cd7f22cef017b43f5d2813cfe4ab
z5b411ef6a9e8c905c79795d4a54095f406b0b67d60e8a95379670e58a85b9daccb6f4978285963
zbcffc4204400bb77a32f48135ffacb710253eebdd9af3051c27748d41bbf65ab0e4e0581eafbad
z4cf7700e5fb162b107cb420ffd9e4c821e3578d7159ed7eee026d75eb9a01fc6a0d0642951d438
z477ba30c8153bacd2c987b457e8fb268bb9057d0b0c2c3f0860a765f81583013182159900f47fb
z077553cc640692e542179ca3d18834ac0d5e3fcb0d4ae0057aec08879ffd22ebb2843b4ccfa044
zc419b6fd5943f82e529ff60328cfc555142418d0429bf3045ec6e7f5a0ca9c5ac49f6497b881a4
z0067fbd2f71987db9392d5351dca073918f0c0cdd4b871b99f83e6d4d5f7ccc2d685722f7ae90c
z59c70e733375e311903ad713c401df3b6e9e789078c2f807b408910fa19524fdc1fc3aa0890351
z06f569da8c0cd2d9bb3c647b66239b9472e5312278b376a6a9a34f240fe9e134437653fac71c6d
zedd4990449b40ddb4a978ecf2c97a8d2e1bd5f4d0f6d59397a3bb2023b332a00f1df3e6e0f979c
zeb3b550a841dc09168a6ea6afa9399c08847974e93083a4df1847a920b4a0d21416746cc5d6a13
z4d6320130170ef9c060772ca22e9622833d5dbb1cb3e8f5dee75fb27e7d4520650af1156f7078b
z03f6b74f3adedc8dacf549271cee4771c32409b599daece13c88fe0712e086ac72f92d6b435cca
zd8b563a9f49cafebaec09237cb7f1ad8babe4ab7de0cb385767eccab99cd9b677ef3ae73490542
ze2ed870f7dd8c990628c533c0e85edbb6f9a4e06a6f3aeecb2b23ba59a26e0a9fefb589a465078
z1d8e41d7bff33473369d44c318360077afa67f76d1a0a8a4cfcf15f33ef0b2d9566dd6531e72cf
zb852df6fc75b57351824efa319d751a077caded4a6a8e48753cadfdc380becfe233051b3a6ba68
zbb05abae6a006bcfd747df8e85a457df5795e2a48a6a44ac526c1d644b0caff9e63306ba8549e5
z3e59b94b67292991ff2c3851bee96f4388d5b8d6390e0558496511a2da9269e130b8030f4328f7
z8678abe493db8cb2c5536f02d76e73a33cc8c5fb6b4ee44e91ec651b1c55752c8536e2806ebd84
z72ae3e5f9bc0a1933e0f70bbdb5dd22086bdde4f43e9d7a63f749614af0a4f53d42c8feb505388
z9c004ecdeb8adfbe37ecda7ed8850420f98f69a4bed1ef8eb259e054b9f8b39091fcec135180dd
z7a92b0642b0efaece8ac2ded11975eea52d1422e5f1ae9dc6ad3f3dcfb95d0038673a1839af38f
z91fa7ea9a4ffa609f27f258d290947c9a4cb316991c6d029ad1630644f22079aa17e5d780fabed
z909aa21dc110fc1a8efa020de2b6ff1da767e00b142121a5efd4a07507016a17810019562bc8b6
z30c9336d257a26dc811efa2603833530981d8da3aaa5b7d177e035dce8435aac1b8782748a1c47
zeffcfa225de1aacdd26329a8be9a3df81605d01f988c851046b697d13e155607bcc6b7f6a58b7a
z363ca1e0ce47a86a10405d15d018f72987fb77da3fd893c777db062a04bf76dd42d71ed7ea9ef6
z7f940476ccddec2f6ba8e0f5501928ec8690ca40f39940e54761282e0d1972b34125eccb35ec25
z74b709b899869af746ee8cce2974333da70534d8839d6494440012c91c311f387b3df65b093fd1
za654d6349ad0cc6b7505e986c788fce0ec077b0f901b0bb592ada8b02bc3e18198f8868c78a6a5
z807c8a5ff14202f4d72d33ea4e3d3f404b7ee37f80392708cffd9b0b8c7e6adb9c7a7af50f4c4b
zeec834f7e1503b12999c684b2c157b80422f3599d0933f76caa4527dcb58c0777368bb264bf2c6
ze0962491bb654e0c29a71f165989e819e22b3a4202351cee7bed61d88a033878912f114c703498
z82ef6e559745797f8556b5799c601478ebcf8a31ded00108d8222bce7bd9eeb325ac26837f216c
zf171178f51d33ac7cf0bcd94703fe101d4df27d9109fb2378ba8017e1a1dc116ff745bad2861bf
z2a5a2f831ca577f765311b1e231c1bb67f20f1441f59119f537a265633b0f75e1fecaf5efee2b7
z59ad40f99fd2daadb1e63df877e4f084d2354ad70f3df503550d611c5240d6aed0c5566d48cad9
zc753a7885ee88aa1c7660715a98e32370e3db15023d227cef062862c234de18b0c83e54d939976
z5dfe465cd35db4d066178a8440a09f88e5ae144e47770b329d132a27cbfeefde8115dc3f5cf6e1
z4f121de77375424dc456e32750f357289ad132265ed0c5960207d910b52eeaf9b7d5ca7020e837
z2ddc7b7fef482f14bb789322cdddcb2f920d65f9f86b0bc77793969851270e3b22a45c3c9807e5
zdcdb2b87fb81c58a452bb1c89466e9db475f947df5751b6f855031c511c23ddcf0db3042e0cdb1
za7134eb8d4e418d807f249febe2a14bf085ff2c2bd36d0efbadc1804376a007b2034204bff70b8
z83574cf595deb80f6ec4d40bc9eb9caa1805fbdd548e60c5716cf14417107a60d315e35832efc6
zef462d63a4f2595bcb27ea68c631255645db55052e0263d897d863c6733d0768387c508d7ea7ae
zb6fba8f37e66e1e5915832c45b99fc817650ae68b6d147ac30f24fdd7d990963471fa632f54852
z3875610ea8a8c386340743a819ce0a7643c71abe4be0aabb718b37b05ab489f479276dab2e00b5
zd0bd084bf65afbc3e2b2048edd9c1a633b32b2d10006a52229b553a8ad11c422149e61e88602af
zc5c87f10c88c433e7c95556d856bd65ec76039e5bfc1c9115cef6d31a91e2dd19b18d44c3d3fb4
zffe3d957acdf6df441570ad6b737b2f48bb548d2b8c930bbbbc465cc75728452dbc8959658e5d9
ze66c11702faa59e5060893f5818fc263788ad117252d17b7342a79647a0ac5e7d833539200f8d5
z5ea6feced0c0771e11a2822b153d175e830d7bc61ee50dc87335b1ee57dd482aa037b99ecc636d
z5fe14b6101df16279ee13b42e679d60769512b800c83f41e1682ad67129c6f11bfe00572db5e3e
z178e5b42f2b17b018818893323b32b6d791c5a853822d177cbe50fc824d5b4de49cabd9d934963
z921c431b2f955e4a1bbd83ac56cbb9cb7f004db960af0f65a0c699d81d77bd1317251cf1d7fe6d
z666710b4376075bfcee3868bbab3365816e2a06aca8bfc99316a7dc9d33c22b4696255ce0f906a
z119c194520f992636e65846308e2794ce86cf56b68b4dd912c374fb445a87240eee3d17c1adeac
zc3b2c87fa32ba2ce1adb0618243761bdc8b2f620a212c75ddb00f367e7b643a997fdf9e9e0bf46
z584396f150593cbc4e883fff5696740b82a4ec2be2a21c8489f5d5f279ded97167b3c20c54902e
z319ab3a3e18b2dc3e7c4d0bea959488ebf6da3fc01815b69b99b998992b5382d8d94e3fd592201
z0d5f9522af2cea1a84a1a90252bdb0d132d8a5c70e3e0625b93020d4daf3fb2ae28f4dfb494566
z6e7456fe88817d6a77775e103562fab6589883de36dd04a9946c366a81bf41c42d5f0583c28ae4
za0e8959cfa014a635cb3709d8b9caac9608daeb952337a9e598c71524faaea8282aff20170781e
z79afc932a73a666ef2e9477e78b43a6a1fb6dffa8cadf8a469bdd80d390d77c189a1ed6cc2e360
zaa94e2f37ccfa59bf0479803d41534e8f9be830806962fadca53a82cb387d2684a787972799580
z3251fd492728ffa645f79bc510c3ce299b4a49cc0c098e176e393b17929762280cc81e9add985f
zd16e40c3e55ef687caa02dce08e9830c56567d94c4c8dc14e206ee8cad3f933b462da908163581
z43dd8ec41285c32448a8a8aea491c7dbd998a1a5f536cca6f74025b46cc3513a48005e07bb792c
z5ca38c9ffdbd3d4e63589faf8d82b7108578ffa823ed98eb79660d015f3cb721c5dcab4c8ac6b6
z22e355635e2a7b884a8819fad12772340d9fc9bb5b6c679964b1fb8af17fea6d77c1c4f3e3b6df
z94c0584c56858d29e609a4c65e7776619f650958cad6d81e3ac37083e150bcb4cd05a07cdd928d
zd7bad21726f9ecaa41ff7b995dd26fa60f7a0a1178fa144bce2864c572422d9b135ce2411c8096
z71ac1d741753edb4c795920db5909fa64c9b3a2547e5476d78b75c7701169b9d6ee0beb5d39a50
zdad0dfa6a478766a62229d68485020216760f5c2dec0d34031ccd4eda5f1ed02235091f6155675
zbb12076faf64d4d0d79d73e352ba7e8cc496dd570b524cf5fedb9ea93c3813f1e3ab87d0552ca9
z7b90d84d327c1a69b7514f296aa237b6292728d90066e7a383341a6850b67e637caf7304817ac5
zca14fcfee19dd0bacdb4a866fd851a0e82af19f704d05449c6d1e59ff9cbb0e59e6ca5c99a680b
z85caf391d2e07e9401ea7ad5d663d20485347aec611d663f543c6c9f9445d1d7ac59a6be5aab80
z088c6fa3bb4f785147e1fb537682a7af585cea50465c5fc4cf8d56b89581c10be52ec49c0e4101
za0e077be1027a63d6222c438351b5d856be2cefb1982b0d1c5746e4388784bf00374e875dfcc3e
zf99efd5b107dba40d4d74b8fe5449c7c24a2bb301c7d0211b86b68a80d331a5a25ce66b5080036
z6b3e79897c73d6fc713b8b8c610a0eb75ce1b249c0ab641a557e4d072270d537746b660b424665
zf8b49317ec6c7c657a59427d781741340d76871cb12fa1cd54c15c98626485793858b7020599e4
z295ca78429909b8ecf8663ea5a0f34cf7e307d0c3d4af404595c906402bff33ea0a4bca7ffd0d1
z46e3dcf06bbbe198af6c664cd9398acf06b1b4006f1e9f698cf646b7654c35be3bee54ddcad55f
ze6eb17178347c2acf6291866a4c56f8bbefb72f76bddefba1d9eec458c07f4b9f5ca5543b95883
z18ca86995cce53686dccb3d8e933a01ba23e6d48039c7717f63b90c2e7e63d10d1aa46315e8617
z6f35d54c4d1ee685dd458c0f7a400dbff755409fb9d8a62aa2418786cdadf77e41da356863b1ea
zd8cd964583f8d49c8a1b3c5c648e509e90503047445fa8a1ab5aa76809e57491de671943c06916
zdc910724923b3a06da9ae0e83d9ff0decfe43d51143e378a64af3a2aa78bafc190b81319b6b8f6
z7198ff1e9ca5eb0f826e3756ee88c342f5c71b30fb067937f995d2bed190d87ae3fce6d76ac0ac
zadee3cf86ba020cc4c2ce595371d1ebcaee6bb298aed59de449e1d7ff21e1b1a93e5229c8520af
z34ed781dec506281f84ecb29b3ccbe084d3550af21361342a73fb2a240bace5263aaa5530c9921
z0115600529f74d68c2b50033f461a767447680367d6be23d679e1d1dca5d1e1622648269f65e42
z0f758f519dbb7b2524945b272c272736936c1df79a7d9900c9c40402f8d2232aec48977b52996e
zf8773de42f8b0e44cd1ca2642ffba37232b6b3eaa91fbc0daeaca10447069f27dc2e5821764236
zad6f459c7d49bea862a0557a65f078420999a54ff328efaf1d33fef7791450fa1fdbdc95490f35
zfb99a33b9183fe59a0016a21c1f9b5639c49556b41be2afb98fa2c3f7cd1c11a921a126135425f
zb15c17b16ccf1987396b7100fe27dbc6caa5dc6f605a5c6c1cbabe4d0aadae97e9a02f00ea28e4
zfaf19a6d7fab8090decaf9b5211affb1f5a018a3b716c0acdb18b7c9f5590a7f4fdc0760f87c37
z0d5a95c212cb2bc614e1e906b4f581ffb401318bfc871be1204e23532f86d474d87cf29de75049
zdf4be3c9e3496d0f1968bb513dc713774ce8f9644f23dca17d8a3f969e41cc1614c9a29be179de
z999119faacf9507de86668a3d60361c5e4de70bcde7fd25332c4af2f93a9a8ed80f0d31b0802a9
z0f8413f78e5112830c7e35411d636574c008365861c33a6dcaf1ce53ad0e08a4d76d755367ac62
zbb0b145d90a5e071db7b12936c705df5d40130d405056f70abb5051fc618aa24c948862479a005
z039b67f7dc2f53711a318bee288fe054718f7eafb41d0cea4b588aa4a12eb84f695f597e8caee4
z0de0f2716916c61772cabb27df10951e48993b31318f89f9ced3452aae6e27d101747a1f0ef93c
z826a50eaf6b04ca558b61572d337a053bf86254514844c72eba42a9c955ed6c322315258695162
z7685c5052343fed62913f6e142e1a6f50216b33dcbdec14d32fba39e85e5f7532a19bc991ace3a
z1e5ecd8ca7c8a50777912aa8254e45e64582ef125e3c2c1a3e666931268f7136ec953c33312a5f
z9e70df528dc953427eb7f7f2aaad5805fcdc074659ee21732f9f336f04ea64f13b0b7ac6986483
zd27dbb01efb53e90a4f3eab2729ffd32c402877acc3d853b154887fe4e288d5d47f261387b0f36
z728d3c1d8c79112f20ae07a4ab668da35a9447d44957f651ed6f3c8fadcf335351ff893f3544f2
zc03ad3cb000edef81360935a77a276a31cd976877ea8b4c33933699f25ed22c74206f8edcd8ee5
za1cd39417567f3244e731417c03a58a599f76a5a0706d8e4750dc93dda78cf8dd8c4a4bbd06e1c
z013351c9657a0aeda6793f8d4c30082efb57e5aa1652d979fd3b770e1890c5e1aad835f35d5202
z935a5798458ca446b97a40aae36b83c591c7d19f9714ea65328b209603a9066d1b9436992c4181
zdeac4535ec09b9fcd1842ba2a9b413930c5d4b0836c1abe6a9a55e617ae35e15e4d0889caedacd
z4c422d1b48ad46054f8c2dff45e7e0c2ff8d38fe4b18fe67ac9157c066923592c680cacc516097
z7597047858ed3200694338f76db43931839148a769c8eb0dfeebd02698ac2b9feee788e0a3575c
zf6f51662fd90be367b8afeb2c6b9e74af40b1ae35fcb78fb0c0e3379ceff8f344e67235f9b77c5
zddd3a6731943cade8524c0d62e5a7763c428de317587a1f6910385470f4d250b2d7a8937df748b
z0965e994c9e3448db6a47b5c3c604df7594749647c108d956948073ce70d99b1321d5caef1c484
z87437a253b7f80da020faf1d5b02173899f60e38c5b2c46e5d40e9e19c125e598a6b6a3a991f4f
z9f86a09aa3efb54238003a6b28fa928f2d1782edf7febb3a14e0b1b5fa161ce4ab962d81db7240
z358b48ad9ad17c79b4b3b9764bbed5c57dc9cb7ac2f0bdeeb8295da4c95cd88726a326c7bc5bb3
zea6e29f3b1792fed7d2bbfbedad1dd3d3d2149a69d5382ee74825a50ecf7196b54ea4c079e6efd
z0bcbf8f5b99776387ea6c3e0915242a10a2cf3d264acf2907f170eea859771bb0f36173f7df22d
z306e19fc7b64a3c4526f05931a7959642e6235f33d401a9248a4314f35d8c2e5953c8fe2c82d66
zc2626a7534fad06422ad416af43f205d251356528cbbedf2efed73c35c7b2e075484aeef65395f
z27db0e12c2a7a3ec677d0b1171bb7afa3b09e43e886434b2a9994b639552a8ca4ad488926b6d25
z5c9e038a229c63a0d88985e4cba4c4cca44b466ff4769a8442fa8cba1b6725caf021e10b93f785
ze6c79e0753765c6cd624d5b9912b38757796c088e897423f1efae1a1b7ae5f11aac74156989982
zacab61b0d9eb1bcd15ac49433adcafb47ec1f009f918db79a47c5db21ccafb1499c165a72a1c15
z5cb3f5edc31bd714918ad25350208bd4d973743b5cf86932e8b51cc18e1d3b6aacd7454e4eef12
zfc0b8889586c6502cfea723f5bdcae5c9a48d10d0adb6ec99b0cfde9f937b271b6ab222d29c3e0
z13b55e3bdb8fed231f8e36aea980db97d587ff53e432fbc297441497a27091c913dd061e305986
z7ed931ceeecba9ed33a70a4bd555ae1e864dc676d2dea2435fc87fbb896ffa2690fae51dfbd3b1
z5918dfb43d1afaa0852f81382d7360fe30736ca493318ca3fc75591df2a0ae8b2fd8cc04a28a90
zbdc7f0eddc3be9ec904f232cce18c2106b7b5f12db57ed05fd5d4290f2f398159a3ca7dc387ba7
z02ed22820a245da8d3a6e92973fd2843b3a41e5843db1467704ffce84f37f8b085cc1bb4ef19da
z9b72f1b7b79c8d44fdef6a20475dee8bd346756db200d112d592332bbf01bcf7b41bf1a978c732
zd52e0351ee9a9d1f26b3a751ffaa79f75b8555c3dd37bc4cf7833d9ce746e03167a02030a2b80d
z2e5572c526c0f90d3154d5e74c586e1badc59394da06044661790401767f527800ac6163b22e2a
z163a2b9c1af21019ab796b202967c2448820980f928f2ee7e2f99aa3a6aaba1ce63533ee7e3fad
ze74b954a1cd79c1c611ee05366ca662c6433e7be62660f7a197ab3ff218e8dfd0cc420444363dd
zc11d5089ec4d59d13d5a1f49e5b8f27eec74c651758b5f92b1c2fce9fbacdeb004e82b2fca63f0
z5205cf0734726efc1824ba9162703975342d6d1397ef1580a4ba4be3a345b0da2f21ff9862fc30
z71f7698c7b45652e209b0b2f1ce6db3666ac94bc2bf932d327436ff6d6c4e830d9f712cc21a2b3
z5f2f668fdbd0a28d357b9a902883c72d6d019d804b879628c1d6d8d73ab0cedc8b7362d4c8d298
z437cd4e6d1caf75655a3d8ea24b8b06a3ced7a9bd9161783ba9fd0408b501c3ec04110b1608ef9
z1121f26987a802e568c93229a08d10d774357305b0ce790635712acca35fd9eaf9273155dc9efb
z4d2f1758deac8434be26665d4510a89e93d9d8dbe44f9713108a6ac643e924e4d61e01f61309ad
z70ea5919bc09d169094a57c1288f1730d85b7000cc06c6f11c1732ad09580988ce4b65a9669c5f
ze7685e248102ce2cf2009aca42083d296b6c4fc8136aae5b5179db1ff34c3ee5fe6f6b3a5c3c03
z4ced8fb5225a146e658bbf044e7af0fbe80c28f6cd5749ba100f2ac1894d857f329f4201980bca
z266331bdcb1e8f85bff0f2cc0b3f01062d78559d7702c6db6a7093b3c4d6a93b7461a06908d4ce
zb798e1e8a60927617268dd05c84c228436cb3a477fa290b181561ebf6eb16679789b597b910a67
zf0d1a6ac0d5ded10ad5f26f548a33527b72f9d6be1aa82e55104c8e61394f03d6eaf359c06dca2
zc0810aef1d56bb7954d5e8d97c976d82b194ea156410980cf6e9b07504950c3920836932c7a02e
z103a4402e1f8e79c35ecac3f65777e2057909152455d8df991b1f181a030409da4a9ff8ff4948d
z4b5a4a3b004cd701013bbade433a53ddd6cad2aaa611254375b1e30ef3d551bbd42321e3d3ffe7
z8ab2c4f66b05e2e2f388c019be904f3df602b2d629a76f97e7d8c0b1abd5f420831074ad288e31
zd8eaef89c4a4a1e710026ed2138e4f7d4a525ffbdbe62b9a552c3b9ee6527df26d96697d8da1e9
z487568d3295df626cdbf3c57502f39ab87a2ca728c6581e569754c6926509487e7c70999bc483b
z04c5da21081f8547c7073e27b055a6dfeb30cb924f99a37d83b04b508ad58935d95ae5563c6ea1
z99a77b8deca94a2ec9de30d872f717a9e65edb4b97614d3965ac2dc61f5b53d9d768e3f911bf91
z391d1ca4eaa6992b6502c69af470eb4abcdc72f6c2228cfedd718aa16ed68c6d70393d4aaa9f1b
z217d15702d026d8768d508dc2f9445fcf26a33c97eb72dda70bb4668f57fe6dd9f48637adddabc
z812d29091defc04f6ececb8fa375d229fdd0f0749c074189593de7a2349e60fc1cf5407d9018d3
z0d7c29f63ae0962bd9a579efce78ed7ad540844c55b4860e7210d21114259e2afdf38a96044692
zc9333b0d4f021511eaec64ad3bc797e6989b6d4cca447ea174c52479e0bfc929591ac035fbf930
z245b5b5c54a1c0800b866c44190d85d53e7f1102ac7fefc73247eee9ae716417b7688aeb50312a
z29ee62c90d0ce32830beed88129ecde37d6df069a356a37703f107ae26bd0ba8c8ca1c0b499ebc
z6f2f1347eedc73098c75d17d3614ab5c7fd2291aed2d4150ef7eab6ab5c9d86029a235955ffc49
z23f1ef7fb47b322dfe936822d6403c0c0ea6f01946708937f47802000059bba4f71b2b61b716c5
z965c510f575276c219383acf4ecca7b107191d9a57f3f2eee7f5b6921c5878bf14c7d3287c122b
z51c270fcc9b4b34256afc9fcb88ed38472513ef8a82e834d74dd7a7db982d6c49fd12359c61724
z162df08f352ad2631c59e107440848eebfc99188acd36026a97ffa8c2ccf51628daab0bf526b0e
zb703f492adc7417a0bb482965fe51b398ae755b49f02a438bb00492d29d0f83a802bc8885df6dd
z2900d0dfc6c0d5d94e3e0cfd09509804f3bcae244614ac3fa45de87e452c63fadc1a559adeeb19
zd053802ad6af76f80197390843eeba1dbc170ce266e67993a99fb293433c857097693315e884c7
ze60cb31fa4b419b8c41742d563a29155b6e21cba262b3cd153a37aa5792d8bcfd83e4f3c419317
z2421f883235bffdd7478e33a37b0c08c7dc4be2cc08ea60237ec5566bbcd6edb1eba6a00aedb05
zfb0c4090dc8ef3fdb46797307d8544275097124295293a68a86dbb12bbde9c7ad4db52a218c589
z1a962bd061098f88a5fb9d8507462ed781641ecdda4deeb54017cf12ce3fb207dfe9af00782e25
z4bfa9870cf1f15d64d288fcc8d3f7344eb72684150c7d1c24b77dec2adea50ee23dd7839284a90
ze8edd655a846eb93177219f726b37c7cc5b9b53183ea9df099503d015df9b7c5b6bd27e8b5845a
z7d0758011a0f5941d1e96d624d1948306876bde6ef040233545858deda772bc5a4baaefefc473c
z6fead6ce0935844113cd9ea4c2250a7c14aebfe37462cff4949745c8fe223fe960f87180f9e9d8
z6f50fe92c544a75420b6b523cd7b997159888c50b0edcf9a5dc5546cfce4ee90dd6cf7be9afcc3
zf59c7254f9cd3680c9363b07c49c21709b3a941aac0fd987c2e487eaa376f8a7b140c5f53ed041
zdba53ffdafde09a848eb5061cdf902da1c9c788193f4f272b819a5e69cbdba10155905bf6bf09b
z01306c89421d94558d12330d85ad03e1b2e49ef8dfad336866925b2b25db4030452c74d2cba933
z93b9bbad94b47af776374b8c5cfd2aab3314443be5dee043923bbc237fbd0715f94f62f3813c66
za517dcc90992591f30be1da1f3a5625458669fa23a7563abb5d7bead249cc5372837231b709f91
z0bd3456cec7f0fb8cbaef56fb635f4edc2cdcf6dca82efa047c890b895bab6a075f9dff979304a
zd24cdc791da70400995dd1ef891a51228a0fe4d0cf014333148d355ff1ca889aa2039909604598
z01a3f01b7809091776d397b662f76e37cd1bb2bb410b1e875b2fcc058ae2d05d138aafc35e71e2
zffeae100856a838deab7e6c4c9a63354812485bd83b0e1dca51e3a56e51229cfbc282df7c4d440
zd86e7e61ace2948f4a7f9ed2b6925d85447439faccee88dd986634df31ef61577f7bc60fc7bef1
zc1193710a4f79e1fb8a47306b7a88400bc2fcdfb758a1b2c61431632ae1e1029f18102db16f422
z941b66a86ddb3f23b30c429fbeadb9d292544e54e433b106cc3b1c2795da127939ff79b3f5474f
z784c9a67a3f27849bd118a88d4f7745177af86d11b19033630f8ed3498fc861dda620b6639572d
z0939806218fa6fa1e29ec613cd0cd8b8174c277717455efe80ac60ff98fc52f6dd33f17c88cc6e
zfa8b5e59087818b2861cae340230edbf8f21cdcf877bbd84dbb088594ca51e8c4036adb39568c5
z642b1dbf6d66d07f95e082234926be8437d2df947c983b3198dd872a589760f72ea0d902ee455a
zcb849e53d7915bbd718b0a4a641648a9c7330ea2f68b6ab9fefc020c81f818a2132b17b4fee01b
zf0e72a94d18e7c860c4f077686dbaa5eee56ded5f82e2a85010ee4cad2a6715991fcb659510929
z5a6d76f2b789805aec23d91389286bbd056b54bae4ed61952ffbf66c2c0198f258ab5ba2156bb7
zc431fb6b9be84f351b7792a088212a08948bf66861814407123f39e1ea9163cf996254bd9e8447
z6acf158401c8e781440dd6593c42e1069fb4f3cd784fcf3553bdbabc37d881575063d17a326fa6
zc0274304489daaeb598ba2c694aeffa3dae0a2c98f8611e1a8f4b8dd1a0f4ec0b7246e5c0d2b99
z712cd54346c2d901ab4a15a3fa00f42f9db8834801dac28e0d14c9801f59ff464256552700cce2
z9a3f78fc6025bf54c0041468a5b813715b75ac4ea1a90788f838df6aea283111142318fa7655ef
ze59728a1cc226705c20ab9b29e0b408a6b77262c5b3857a6e624fc84bfcaadd0860cb191011fb1
z6f8af413158fe11a78c3f8bb6fad379d1bb256bd86ae4f6147f85558302355fa8ae911b5893f46
z1b5761966270a75c1addd77641cf4f9d9c048663630cff64a570364a825b519f3fd5eb21746845
z3fe5c69473a84d94a8c3c52e421204a0ec417601c1c9c4a8cbf261be8e00a27c4319f4774a087e
zf513ddaf196600ec2e0d2794c55854cddb8d5cdab6df87f477d04b1bf24b072bb23a8b712218f2
z3d8e0d755f5c68c8b940b5cb090539951e78f63c6d4f0c03044e05107fda74bdbffd6d1d7bedaa
z8b7db21dd757d7be265ff5215f06419de03bdf60840a0e14cd7319faddd44b2ad95b518497cd89
ze012ce1ba10d885f6b6ccdaebefc2866624a771d4d88ab6585e409b7198d9b8f118ba7969d286d
z75d3a9571a2cfcb6d2bcfe13e745ff3c4184f5ca8d5314caf45b2eabf11bb2b3e14200afcbb69b
z252977ab0ff339533dfc1a0f5352879a1154fc8c5b20be21a90db33c4920f9fd90eb0442a2117d
z69652c85576016b4710c38b134da013fad0fc7a862874bbba1a623521024bb5106bad48aebb731
zea7e375de03d029275ce7644a73c538cee15fd53a26ad683289256455e107753841713ba2733a2
z71b9ced998199b8af3bb2ab7861fe77234a245524324361cd7bd255e91b5e54b70b8c08a27a515
z021eae64289e2ae3ca12d6725b395d1eb673735968d5fb62d687205da44ab849d68de299779319
zda222695208f9f8287efb110b4
`end_protected_0in
`else
`ifdef MODEL_TECH
`include "qvl_pci_logic.mti.svp"
`endif // MODEL_TECH
`endif // encrypted_0in
