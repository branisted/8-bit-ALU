`ifdef encrypted_0in
`protected_0in
ze74c34e226135848fe16db9ffd31815111b6d7fb642c521a3f628cf6da949865580b22efd062a7
ze90adae0e65e66a2c36a587d0a790699161455169ed55a01f2084f11770a774ec4c588039b380f
z6de9c5084882a40b79a175f5c2114b2b6d78b070cb806e1c0aa9258297f4687ab308bc470f0040
zb0b1de382961eeeaf2e279e1462520fc31c119af8f2b214846f56c2b3cd2eadbe4099496abff18
z15cec83ec4a77b868344aa20ba7360908f5c0de2a79abf8b3534b883bb12180f68b5d4beb444cf
z3fba8f13afb0abfe8fcc4294810f75afe452434d2d0f1166236c82f76edf1e12979f04bc35693e
z32ae028996dd85737a8f5adc1ebb94f39c940246e887647b64782cd7ab429b0544c173176cede7
z01dfb26b1f73408344a52b7e1f117f12bb9c8077b34876c2e6fdc085981637012dc9754765e1a9
zc512ce062e0b8fb16a214591f5c81e1353b900a611fe1f4886b57940b41b7f2ce99a7b84b04b90
z916f717e73bd10589c81e207ed77ec660a8cbed5b487fa50acde1b055c8870bd8676023f21ddcf
z9c98cc47cfa2d654ff1365d1f45035a045a66c5dfa827905026201628cee5aae21fb892db766c4
zb5b1406e11aebfd6dfacc9da5ec03b70c276807a3eb15e28ec7ab1dddec42388b9424ea285623a
z248195c9f894b36317ca6e59c86f11031163f5f52d70922c037057ec65cf19cac58583b899d7e9
z5b165e80500bb14e47281dc3000df4f603e04a7828f6f0c74040d85c3c8ad036ef3bc1d66e3047
zcc69669174088ed23fe12190fcd63a31f35be060169de9e6dfcd8e2e136a521257e26238d47389
z9e12b9d8259ea711a62a19a8bf70c9dd32b0c623a9daa7936b9a056ab69c013ababfd847659ea1
z7c47d50e25dd7ee7d62f97d0be8df8df8e53a8df63bce8cbe1908d96440abfc02ed9b47103d61e
zfccce82318c6b8647b99c745ba86ac94af0b8aac10d0ecef801608d09c7d7ceee08e993f494a63
z155d6bbd0c1e854a8cd0992b5018499c802025b18f1133108aa46cf5580f2f6431c88711ef6fba
z654e5068776ed5e70847fd7742ce091dd78cb0c606e7c7e4c7ac905c8c3a2d05172090e697dcbd
z61bf0ee8d2f5e765e0bd94eb6cb5fbab6ecd9374fcd1ebaafdfbc33ab217a381f2276dc6b8c706
zce4696c087a5e29d74c9054ea11a41e569fd89134a599ce05298518c4507e34aa44a2f5345f32f
z0049d6cdc38b8bdab8efb0af6b69c43b5755c73f3ffd16f06d29833562641a205d580e68bd7cf1
z416c2c1a2245d61bb55cbce2e15303aa0cd0a077bb4f7d192a0d33de6bd409a2b9b74d21b2089b
zebbb1478d469da43b1341200dcf0dd069c10e87d05e068909977d0d80dad335cd0124f9c4fa9a3
zbb9db65f219ad01a2c83fe4d38e47604c666b68643a703d34b5f1965c29bc87098950f47c462f3
z070c01c49ae42ab029a3c6cd81cb7c8303f089cd28b99cb1c6805968df19184336f2ee176ce523
zb476a8a4262961ff659522edff7729c09c1d7ac9fe626fd9c4c89aab4ccd7961bb2cd8e9520813
zb7ae8de47db545644d02345f1d6db615f4d99e5213f0334b0e378714bc4b82a00cf812b43e5c06
z99e11087d3dd740ac1f83781c7e608553c372af49c072bdcc126a0c3e63bada73c5b743f809ecd
ze7c13e5e2ed99cd6dd711cfc8c88032b33b178fdea8e62b670ee25ef66c97b701e51199c48e633
zb6fc00640c1ef4127fe553875803c3f7b0080a643ebd118f77ebecfb40c0910fbe1812a1e4d35a
zef472631e2ae7c6964de6fa46ca39cf36483401e5542531533856e63ce8e749f32c6ee2fd4f589
zdeb77dfe80dfd34259c8613f6c2ebb86d6833d7ffb19e9b610d84586b230388ac5b697a04b6592
zc1c87ef34bcda47b352b25a7e461d72a1438b8c6c5e0087e1b7b586ab972b83d7732a51504d163
z86f84c06f7f206b38c5bf1f8a06090dc70bf0a0de97ea51664f059d76426f7f7847549c85b3397
z9c319f3486647e17c3d64792e4a5b7d0acd365a24200c726519ddd168d9481b1d26112db39afaa
z4bbed8ba581888cacd7b624fb7976ec7787cf170fb10428780f99444e0abfa53e0a3b29bd818ab
z2b8e07887fb4e77d5658afaf27025d81c446cd5eebcac567ff0268ef606cfc0d1d2f5244dd69e9
z3a7cfc4c6c6d1b73c467657acd1e11ef42a950ca3379341a1f8b52d7892118af595cae5bbc6626
z5f5a95ec8770cbefd39f3af719563e1f66a5d503ecde9a76fdbf0edfb0dcec52bd8a140ce93a0a
z0b1c2443b82c6efe5d772c23427c4925f447128daa869698110a922d5be71178c035125c71986f
zed4ea707094d24044c7dee2cafe64eaa26fd3abf2abb44deca1f6c8faa85eff1febcb87decc77a
z9d9ee715e5cf12e54c641232e889cc2fc137db2219e94f80060617ca6a743c1b8374744d1a3fa2
zfd021c5ca59bf7763b5eff8965a9a9f140acc93afa93007247ce974f3f62b35e7dbfdbd42482f1
z37cae883b56fcfb2426cf18d1228185ea5d1318d37c409d2b6ca523c4c8bcde679a98a6afcc92f
zdd201d36a72d7ccfdc4dade934a7aff50f71daffdaf17e4db79403193bdf3b0523d49b4509661c
zb356f18f409fe153d6af152ef9133b0652934cd062348bde10f97df2ca8f45cffb3cd180965c96
zb9a220bc9606aa76fb6072fd1beea31e7723234a74892c5114b2acba33e7da22bbb333e6f9ddfb
z886f185eea82d4a643d1629ebbe8d239497d48242ff9ae7261d70be5b7589b6d0a54a48a184d8d
z4438f90c22df844f379a38cec22d69d40ee84fa9e7a8ec32910e701213062e863a000ddea0f3b3
z1c84d2c95ad7854f5a4daf80ba5c364222f1931c82877f1ed6025958fbc88d8fdaf40adbfc503f
z46bcdedbd5441c98cd7465dce07a93ad89a3ef28bdf55c0a1f9602bb821e0089989d93dcf059dd
z6071ea5e4d53e2b449bef348562b757bbe91575c9c926170c7252396ebeb7610b1b9fb574aedb7
zc3bcc19d483073ae177328bce76cd2c8a83c95e876433c2350ca87d124ce19bc6fc778c9efbbf9
z50606c87c6dc28e9cdac9be9f14f569f2fab6c9cbb10bad5cf065478ce717decc45e20ef47f2cd
z97cafbd35c41a90127c2372ff7c48eba2058ab954324405f460450546fff8a9e303e3855dab2e8
z6b2ff4d77229945fd2176af99d9d1e86e966d17e9f7118edd35da7d2455380ddead2cb6ca07707
z9e8ccdaa30377c74ed2438a35710b9adcbefd80bc0dcb2ec23656240b9b89305d3796fe75dce8f
z07b5310915e5e268c430402b88ea03c46c18d7b5756a7032a6d5f5ab6d26f000aeb1885723fa07
zb2633806e8e9ccaddc3894f4d8d9ea98b5d04abdabd1c507c3521d0d93ea3350f4aaafb0992e0d
z18b03a5a54f06ad095b2865c30b76c29e559987fe3948ba45fbb57c38e15472102ac319685ef11
zc3112b9abf6bda90033ee1610525ddfe5ffe82ef5a13d1c5b07863658da888a4465a35f7ee9980
za6fddf71d0be7c71a1047688646f6e7f8111d86f6df010206fa0b7b3a771ab21bef2879c69185e
z735cd8e4ca9b773a1b3536e35d2bcc38275985eada54a87320a43935727dd9eca1f94263022a10
zbb5b82fb3d9a78b35b4e7d2cbd95ecd3a4207b1c2100f4a1ebe436818d0127f3a22507eb5995d5
z2cc985714b855fae3687fd3b26d4957c9232cc968cceefa2b2f2703b315e6ad0280fdd7c3ee4c6
zcc8202ceed6d6c79ff116aba023740f09aa30888a03bb8856a59cee28b2c4cdb8c8f3e603cf347
zfef8b607ccfc089d9632d60a1013ec48e361e36bef9ecf126911be05e0fdbf22ff4c9e73c4a756
z1ab0d6950e103c62eda9db0d35c5096c7fa831371c69574752ad4cd6454ebcf97f8548866b9837
ze69a7f03943e4bc274f399ea47917201d25fe1c6e2aec5cc1178b8ad7740d31051565ed08ae5a2
zbcb45610d3d38e673cb641312495c71ba29e6fa35ea5933259727333958c82cd6531535033acfa
zae247aad0532dac04920e9ab554dcfeab4f99b3c8b6ef4f6024c85191f91cfcaf07ab78e09e654
z4f88b0e23308b2cc34282103b24236056018f3669c8030cbc7295d498c0fe35f98bab75ab74ce0
z8055743d057013d407eba7d1a5178a673a80dd598abdf4ec3e015f670e62eeaec13e3b60d3d8fe
ze7ba6acb12fbb9ddde655ba49ba26564430d15e9f811e40b57830a5ec8fa9d3818a2cb06af4f41
z03261bba8ca8586493b8195cf69b561e956e7b11a9318f8ff1bb275a83c89e42fe5a625c854728
z0ed9ed72e783e68a454b419cb6a142b80e3e2ba7a697d311df415a6393c02e08665871fa7f1df8
zae8837240ca25f9fb1a9768b0d40570a093bee565e80b2db7550c5e6a092b0e803cf340eb0969d
z56bb8885c40428fcbc27ba0ceb1e930fce763f07b7d6110874567099167f52372abe0499c639bb
z86b137221531fa87695d72eb9ba568a72aa8f2cef0df97514821aeee15e69ef1590d0b6ef9e195
z07b54fd11fe50f182eab5d575c5835e54635c28595e3bfc68783ddf773cb8bae867eca51da1461
z7b89060619cdae2eee71dd645fff0f293e2990c436017444cfb15d86a591f306ddb71116f6efd9
ze2e2b82bd127da4f1f50feec15d7d5f00548971d14dfa86ef0862f2e35cca9bd234b37a769a086
ze60b6a8cbc5b392e53ea1ca8384edec0d009a0fae2787cca27e97a2fedbe7c6a26b05813dbc2b3
zd7df33c90515c397a0c3a349f781068a330aae24c79a22dcba3717cbbce8bd7b1bde5bfdd329a1
z2463be888b49da7c59026c1b5faa57b10869eafea52e42f35fa6b2bb313d9f6dca1f98b8643121
z5cd2569ff3a80337c2723f808031e63fb95fa7f013ebd857e0ae2280a1460833f951d87cda179e
z2afbf6813ae1cf103095e58519341f722b9db2e45282d5b091aecffd7c085135c1613357839c99
za96a192ce8dba710a3b120e976163109045299c9f0275dc7566a2c7af84110b0cff5c1f7f2d292
z8b39a4c6c59f4b80a0740ddba1a8b176ef4771151fd14d7331866d141542cc44d66cda3b6c593e
za87af1256d5e0e9a61ebbb565c0ac053dad8838982307f5c324562e4ea1f26f9b4341a70cf22b9
zf8f73d5c3669035e89ee502e18a62b2aeecfeabd08a9912de292917abf8d64b5402e8ebe8b8d21
zaea379708a34d6a22442c21fde87b5b51a2a670b7487a1dd9f804190d40795e32092427a1aec18
z2a94c6b049c9349fbe6c36e9ae94cc7df90e15acf716d13b985c01a9ab41e28d4f865e72b8a78d
z381ce1edc6cddde7eec80fd616deee08308988e5a98a6cb507f807da32ef3e7454b10788f5f074
z952ea749249821a1ed85b319641ac212c2c627072a370155d97a49664cdc8c1ffb14e973372b90
z2aa5c089802a3fa11c3381c8afc6eb0cb9765c5359f4f37a4bb8569c67ea98dea3c16004a2ee3f
z6dafc774719ba25ac026a3f44c260a6f7919c2fd390a429b8fc4e5a9a93ba2cc72eca84608c5a2
z37c230ab644ce20e1e9ca5c6a64c6c4a1bba31b31de5140ab047ebea718c368bb8f3a429361be8
z96f1465974e0253f2a3233bc7b59c1283b93deacf5458a1e4ae145da1903a52ad311d53d904402
z888170764f5b6fd85e37ba9f99e719055d8a4479a051f38461ff6948eaf6fdda4755ec56d5a807
z937d0ace325116f4179dc8699a5573d569a03b0a730d934d027e21b201310db25c40f1bceb2a12
zffe27fb1d388dcb1f4b6410d496d801e55e50b74a139797deba4f16815c76b72482b683cf0f1d6
z7bc38afe96331ec59d0ad1bf45b41a95078725ba5ca9d024ea3c0b6fef2d703f6135fb7d0e91f1
z7f3142c38c44bbc6a233348b1b7d4e772cd3e71bb313e631c4dd825d2e5c3e9665da9e6a7970ff
z987037a63957f37c23fe981b526cc1e406d73b89f4758da3ab859408749be4b8b353a2b3253d27
zad99ce71a0b49e575eb19a3a6f00a2a2b8399b80bcf5006164a73b171419b97cf63aa8147b30f7
z8c0a61adfcc53670b79582e7551b04598cad9866fa3c8ad0b5eb81904fa36f04b953bd7f84065f
z9e467ac565e07f65b9b62bc79199056564e23055153fc18223e1db38fb8881d438f34404566644
z452315d6957574e088bc26d9e8cf75fe7b2c8ec9865589293ec7b7d64325e97590425c6a86b6ed
z1d6ac87606ad79f68ab03ca7dd0f1f0963839cd7b47e4ddee03f9f028983489fe87486653ff6b8
zac6d3bb55b774408100ea8d49ad2ccfbd25b1d3126b6fc966b7648af46452627759d350ffa113b
zf9a63554bd71dd100d871730772682610373e27733a707deb0afd5258e01f066f98227b32cc229
z923ee9ff47c3e1df0f63228c1c77f27d15892b2b99c43a22fca441142b2373a6ed3cec2363aef3
zbcdc825b1da40564d5ceb8f0db2dd921aca0d36d66da5b7dc70931517d449184c52392449a9a30
z7d1fad30dd632018e4cda9b9f7c3128d6b284f8b714cef26c6538381bbf4809757fae3aa56e54b
z968d18cd4d13a266d3430b80cd498154c012f0437dab1b51675b9fbf5daa02284f35b25bd404f5
z8660ff306251cefab07797045387e67b226818e144ec88a0a00dea590f93f3acf231efe217a339
zcb7c2640ac074cca94aab5ea294632b6a59308a718c19fbfafa2edda5ef525e5084df2f62ea910
z94de1cc2ca893167b1ccb7ef29e091364e918c8065b50e009c2a166c5e17f8e8ea3df26fbaf0ee
ze725125269fc53aa7b71a7d5796e8c7571b83a9295193457791b010563a2d2a8cd36550b9bc66c
z46edb320e1f80ab4c667311522c66535ffdc3c09e1082203333ce5c3f154ff64e1c3c3d4911af4
z6832ad686274eec690422abe33a4ba76c8a12cd4f864e4558bef3efe94f91f0ceb45b9d858a426
z5ee6aaea3387c8da69ace8511d926d8de8f4b65ade1e2aed2dcddb629353b4ce058c9bd162c191
z20656c928b1480583a73acef28bf7a8ec0f9d94bfb5e8dae4633fd3ab8dff4d2936dbec3214498
z041fe81285064e519f14a7648c5686e5c3332dde9258b74e8a4f18b53a6938a717a6263f69a710
zb5781afc1f01a7073f7b9453857d6572b199e844d46bb5d410d23f3a9dbf9c143a37bf679c2e7b
z21f8dccb155469dca4283026c9ed1289760ed3eb532ef8b61eca42dc89353c4e3ba684fbc551f2
z0c15eb15514f1cd77024894821bbf2bc222e65b326826e8a27f88ce11a81d9122654ebbab93c54
z9fea91f734f80ef24bf963b9fc3266feb67e38b99e65578df3f22c50353f19eb9d1bc9591f186b
zef179504812b76509b0da1fe4f528c681c4833d2dc50d1cadfaa65376e348684d97443e65a4064
za8e7bfde4ddf9ad0173e75cb5c9323cbfd802feb8ea7ad271b9d8456ab0b64eeef47732b73dfd5
z9932aa067ace4dfc28c09fffc90618074c2e0c9c04b2ca0e0987c53ab63d319ef7784ac2c63ca7
zbd7bc2b4ca84958a9e111aa55bbde8b02bde8c8e2525a34896602675f10c28efb33953cf89a66d
z8fbe734fc42b685cad35a844b3cf0345c33bb8bca93b5519ed71b547b6492b2970e1f805ff668b
zfff5f5918a3ec3c538cc306a183583a3660b61353d3fae3c7a6217902977c2305a090b066df5dc
z90b0b4177d3eaac8122d30a77847c60d0d42b28bd8f093dfcc5d6974540dbcfa717939d03421b9
z6fcc3b26365273bf41587a6a23ee303f60138c28ab67aef9ae8b33731079008b9e94d739278cf6
zbb87cb11edb71e687f56c33367639f8a3dd2c882d89131bf991f7726b5308ac5c3343d43a20bb4
z4ca0a301a328a7def0b25949cc9f6370079f9d5346900f9a709326e1b0d836091da6b04520071f
zc8995d6523b4feae5269acf727b14034f480d5d40099a91151f9bc7eb174e00956d4a80b094388
zae8bb614732bd1e4520ef356f154f903402c79c425325f531e51f3e6e84de1e23a475c3a60f02a
zf7dafa88949409a1217ec287c02fff0136b2a084e25bcaea0f57eedf248e7fa0e3e07077a21586
zec839f9e54564e126d0b49c13dc6b9ddce5f86be9e59c4c1de600db73717f300a77713c1a7cb4d
z8b7087fb2711509577933782b0965d797aba3ac748a6094a644599ab51138e3e5c960c88be2339
z6e7897cd31d4ec01a5717a22d49704e2fe491b58da643ed0920573c5fc18e1a798a1b14caecd14
za449c763823b6b7cd2a205dafd980c3764bb5f9598d08c483d87a3c5a2b25bc6d5a980fb077d08
z7d04083072c851a035bd9316a2d9e56c92d0dc434be2511820b3d92f0a6259e9693637e85d0108
z963b45f408d040a112176fd25bc7e3bec995bbb69ce504cb658b82b390ba8a8fa8b899b71cf8ca
zf26d14a2826c022fc9b6b86a86f74a909218976f512f2c589070c56c887af31c3c0c4e2514eea6
zdc39fc8767c0a69d143c64b574730fc30e751784b76bcd740511ea8b44b01793f51b8d20c37a1f
z46b7a22f95509924559d763720d892fa8d1012738a5b15618b1579c9f27d03527d1e323f613f72
z92fa511c6ed3332213d5caf50be096cda2fd7b78fea71ca65aa8e21b03a2fd14933011a87bc744
zf5819ef624be85de56a92712604dc15b83e4c97d0939533bf1033c08536322e079648a54519323
z1a43180b0bc2f45d317268bf21636fd2747baf1de5fa0fab01b76771547a325b52cb86b1924b0d
z4c6bcedbd0976710e0bc8141ffe10daa3ffc4453639ad0a62ae1e79e3824512004514315492bf8
zdb4c6f15fe1aabde9698080552a268e3e1ce4d2f5eafe80c8b5c660bf9e48544efb6a1fab34d6c
zcbecb00307badd98c7db00bfb250a6c74d7e650789e3ec5c754ffa1cf7cb05b09b769f8d0a296c
z92fe53fb5c5d4f336ab7f88dfa9f6850cca354c5c3679801860fb51de9e935e7342fa2961a2190
z8d98926d0b0251f64c7eb98fa62546ba3e34bd5b713a9ce2c8185c4813d12fea55648674d2d642
z2f2cb1b3dbb55fcb68d125526ec3e502764de37619a9878776e07753e5b083a1f4c2a20e03ed4c
z5bd0d44ae898992e91598f22f3061ee07e3a2844d218ed8be1d7c5e6d09a8bd1d475cbf961b873
z1dd1ef0e1de91c518605d2a35cb8e7288105d6cca9c515c6839c5a15d0b3c4a2d72c5d00e6b5cb
z41ea0555c62530dc5bcaa682811ad010b943014071f13935fd4063fa26998cc4861121da07f800
z6be6a9181c28f3269e9a162648ca1cebf4d729dd1837ef9519a3d9f70df0ff970133b5c87a4a2b
z962b614570c9b38262c5f3e331129571a85f2e15fa1cc82aecd1ee3a2780f3fe1ce7e6f8ad1769
za3e533601c29da808ad1adc56a306436c36c818187392d159a0848478448a050f2d82d6db3e799
zcec69c7113590f73f68b102fc37646c7bb7d4bf56e65327eae936afc3d3c1d18697731af838882
z5389fec9b837bbf0dc4b28f5f1f563a4bc98f5fd37c663eaa2f8ca7eac26b93460a19403801710
z525ac0cfed3be811aea00161cc951ee1dcba7e0ff7230c1a93cbd0bcb6956c6ff7c7f829d55cfb
ze171c73995cf240a53bf71d382c11cc8eab3256ac2ad6df7da42e2724f1b85c2534f0d7e26a7c0
z0329715ee30a87f39fca923c11323632173fcfcf8887b5e0a720ab4958ae9e9868f9a0a3244204
z4c5f2e1fba675bfcfb203d06be04255203762283382819ec88bd2ac0329537cf46e1b6e24d3059
zbabdd2bab6a43a70369398bbeae77f0ef69d08b794fef399072c1505bd483e20c7eadae64102cb
z35a6bdd17996dc4451437bd941a9209542b453325aaa9cf561a83256b102b6b1767384ca5e16c3
z4d2f5a1d3cb2dd9710787ab3e1f223e55db0404f686860c8fec109a80a481a1414f4a1d6461cf2
zf67b86e3b51013640939339441e01973a575fa28d7b577e7d24a97d8f0ebb0b889d65406354468
z16b9722689de55e62d63c2864b539a309bb28f6dabcce26cfbc9ecba91e16cd342c6af2c5e4107
z57e068247d44d1c2ffaec8364aed2158d6eae28e5485308699814263d9832b9bf79ddd55e9b559
z1fef5e7848f1d547fa4d50ca79f0eadb24f6a4ed17114929c9a46b10d5201b971e4738f22b47e8
z91b9a245f0dda5c91d60b52c3c83582dd5ac28c19b12c0f26cbed201348fafd4b4cb1ccb238368
zaaf334907994b94647f2d7893aff4b789783aad86ce9df9e77be0ec8863fbc019586298778c1d5
z46ec8306c2771583be12d0957b5540d6281ebcdcd7a73c86bd6026cbf0e5c66272b41e7a8fddbd
z7892595948f676447741f2724fe3bb227cb649b4ddaee6ee7c3f9765037038b910a95878fe9776
zb847508a8353e4f023a7bbe30f4b3f12605f559777abd3323f5f0a3fac628457cd776b301bbf79
z0ef2ebf843ed647fde1bfdfe38c8d0851ee723e87a6ab551e1828a534ef973b99ab4b32dbbc737
z8a36bf858faea594f66d14f7e6b8a1cfb7d674914df1eaea8206dfdae4f9a4c4113e20da135cc6
zd633cc39da1551ebf762238e2209841767d04a7195f597f21a25aa7d40f889c34731aee97ba22e
z478cf25c60dc60a55bf044883ab30fe3122f3bbe1da6f4ac5e87202803748702a9a137d3bd049e
zc5d07213c2d3c4abb7fc45911b5bac57e06ea86c830a8027697aa4df34d7fe3fe36d8d7de1d587
zc507ef3aa1850561b49d5e063221226fd30099675861307ab7d55ddf42716624898b1866bc1f25
zd49c0cf5dda570bf4d16074eb6f4b0b1ed3643a6bcbb6d541833ff1cd2b9bc91cdfc3dd90316d2
z98c07cc784246ecec6c565c3281b51862a6d0af43f1a4f4a99ae92671d6fc2a3410b4b64bba6fb
zba530f209658938c998f6f1d8743411fbdd49b8fb1f127043526e4047f70edb637e7805e358750
z61a4626920c1f598414861628a313463fba7dbe846a34a1f7b3922cc669b439f4a28edeb705f10
z01275f4b3000bf1f63c5ff5b75f5af71ab762fbb2b0a52bb5149eb4784b04234be0bc814025d3a
z372f32e19569efc9ba07385068e024f9cd453be5bcff5ebabeea1a06a54f76e44463954418b339
zc92b475075a74d5c4f19d6d1c9a8a057b1ef07d2e59948f0c88d21ca290561cfab1deec5acd805
zd1ea631c32f786bbe6b96a60dd6c44279fcb3dd2fbca1145ccea2d2ab53302eeccd1f0ff5c38a9
z9af9546ce4d174f52eac665df1ad64d5d03db6beecf56fa86c62639dfc86d8a83daf235f42900a
z00bb25d3e3d011e5f73f8c926aa0bd4b639524be819b2d5b421f4e9f56eb53d6e8a8dc371ab8bd
ze9c1b1b3ae79223eaaf23cf1d500a59b31051a984d7e7aae898375e4ac5cc1dacf48199a915f96
za694de891264f0003e46b6178cf3c8ec24091b3fd954e7a67a51522cac2d41e54814b919a66694
zff5b4867338f18bc5e91317960fc437256ac8ad4e5891832f593d90d4bf806e67e6196a2fa4e12
z7f03801ba5be4910334cbd042185b0e62bf3dfaa43c56b5b4e28ea7ba6e02a999008fe6a675ef8
z7e22637c1daed5b9a27ab0db3121aba9f50f463a92efeb7dbec2edd0df69ba0326c02e082500ab
z9a7311cb218f0e819a25f671fe6a53a95094078430a06e8ddf267687eb999e778df83fb97a41e5
z88c84581ba9b30065fda6983bace531e2f83fd7b8308a5a4566ca20f35e204934090f4991e9771
za58e2d89ff67b4a686c779352b04045d91430ef1702bddd7f7f4d2be62b45461b6e2c844d6a7d9
ze4b1bb0cf3d18de08c37d78ac76dd334f46601212b53d2fb7f41d90a1c297102ad5766d54ec6df
ze8088315c6f6bf38333b4881675b57e426fea295475fbe97dc187cbaf0f50603558bc6cae87360
zb224d45650691cc59cd1efb8b5cceb43f587f25536bf7f85392fd3bc8f1753df08af42f8e6a87c
ze7a0ca4dab4ceeadc5a8a25977fff69b307a4e55510df9aef17f48108f6ba4f993c9d965e946b6
z90b10c6666f6404061ff2232c0c34e5f8cafe3b699d3452f122a0e7fa560eb95f42eed8c58bf91
ze5b871040f4d6db1f9c70947197be6ca8364fc25c6b02aecdd204362547ef830165b322fb83e83
z99cb05b324211c682ea4d47505b288274a35e88c83b134a59073c277aac0dfc7b41dcd6ac24333
z76eb4da01f45a9bbe72bba13715aecc8e3521787958c31ebb3414c063cfa179f050671c368dca1
z23dfe3eddc233ee7950c7078ca98ea8e7fd891fb0e2b7fabb87c596103e73d4c4c2dcf3bdf4e41
zd513b28ce2990eb2f270c9730fd0de936797432fce6171e528470cad75f8c13f7e2724988b08c1
z93cb35eed70edf9d09bbca43a179b559f0e3fb710c874f0484fffdae76377d96c0db425f4c4056
zd0e08e0e2741bd75b1c5ad121597a0a5def589732a762beaed1d2e6d9fbd6f28bdff840ae59109
zb6b7103ce84e4a12514ae93547bb0e081aa919abc03f2ef34a04816295cda2102ce26cdb341915
z095c202eabed570f3db61f491a81ca70e89ad3a92f4af6b083118879b410e4b7251052d4a47c23
zcdce3b0ae6a4063391ff1274901073e801505e7d62a379a6335fe01c7b861f16f18b52c2dab05d
z8fd84bcd4d18e7bfb836293d6d31e1f01243e3501cc6e34631bd153d4fc68c03e4abef2e469d7a
z94d74995d5b47bb1190b2a863869f38bbb0f0b21b7d0a1e6d968276a1a62e5a0d6f7cf16ae0211
z60b4d471066937c027b136426940b2b680dedde550da371511c8584e18d0e00b92acb9fa4d5ade
z7dc8667d92f74e373ac9d0c6af768bdbe91ebd879be5b06cba5b85fb943d4f4a25af485da7c77b
z4f234123d2dd110209c7c555fcf5ef064abc8add12e7bc359be69ab4efa06135932ef34add463f
z56d0a9545948b674ab5465b231b3fcb3d4b2a18a249cd9743bce46b3dca039d2c6a83cdffe107c
z6e59030e74313f7c7b7d626c10010db9612a68911ad68e35483b377c46a1a53422e45a27446d25
z969f75cfc6c97d4314f86eff205e390a3f74dd341f7d83966f5675796e4b9d0b369b72aaa27e74
zc66b19dfe4993e728629e09e36c41cd02142507c77fa67e1d8a2f88f9edc5e27681d603e0e11f8
z386804d0aa4eb972f2fe7a9c23ec03d2c19e12911c3fe43bcb5753e0397767f5247b72ca102b7c
zae6eb4ed727ad6f14daaad8e5e984bf97f45a7dd956373d53124b09fda48317a489d73a241a7c1
zc7fa17566be731728f013e43e9179165804585846211a718a4be9e280aa8af456a4c52af30367e
zc15479d8036d2066476ed04805e9dfe7112b55163ec5323282788fcdac016e36ce9b19d11659e3
z9d240e847bcaba4695dfdb06ad2203d42c8637b87c5aa6ec8539f4c4a7c2a267d305ee0db504d6
z94b0efbc842cc52fcf734177b7b28a68afaadcf4658a6c10177c0ec7b07e71064869daa373bb15
z7262f8d83ed2fcd53af3c6845aa3ced3871fca7cb29bbce22e12f15462c71332e2f641a89b48f1
z94ece85183b884e24b2d1ff032fb1a985e5e6d98ba1a19bcb7638e8e6dd2a8a0ab7a83d9cbbb03
zbf3c43f376a0bc59c7c63a08a878a9733e4691d7483eb46ab3025741340412b7f00bcbc220d2ad
zcb3bb5c14da1cf0f705c98ab3763ecc3583c8fcf811552caf4689d9847e3d3ae9347f4bc5bb1c7
z1aad4f85555f7ed4a8080f26ad167d851f02bedefefa0e3c089d0bca1e8daf54bfdcf581de1eba
zb029b14ac86f581e7f09ccfbf38ea78b4f6853fca46a7b6c504cafcf6520a6b317596e59e2a914
z935ce2a66126c24d27af43e982efab8918cdf5a854c9e764c23c5237feec97bf08a62523d95c01
z691d36fbf48a7c264b7f25678a4ba0fb0a6d840f9bdbc53f8c60382417ed196a5c27453c22508f
z7267c926015c69e9d391c43741b339b00c09b0b7b35660779b145c58ee68777324af6cd9e8b488
za7deda663cf673400f61daa061975875ca4114a08871b5db81ab29aebca4174cc3fb37ee691ea3
zd36bcad3d365de0138e2d57c7ff1a68a1e2d0a884c4b6a9b537c360d40945976cc4034851c5bf4
z543dbf47da5587397655c6a3ff368e4bd39ac6c96cee70aaf940b043a3097b0aa0fa17d80d2983
z786d1c0e548b72eb8113af1c5e15879c1568934c4c19a6e886c320bc9ae9136ef10182afd8d2d1
z2803c1a5f3353be4fc8e4ad44d3e73d6321f2d9b0d9366671908ac2871e656f8734f0137eec75b
z6a2a9eb69be211ab8fec07783cf4c90813474643438d0827e2593b75aebce40fc529869002f402
z6342b99cb715800b2caf42b0c5e7167cdeb2da2c824dc5c53bdf025d06e6abd15461ae33e12261
z17cc0ddbd1942e1d5b76deef5134ad86cc9e6e535e302b42ebdcb716e265df77ed1573ced2edcf
z12ea872d38c0333966965d208d9fffed4a84987ed8b76f79331ce1589e9b6e25291bc06d312f83
z4ab14e7a5e51b017e63237f665d08118062aa72f431332eafe0546967376c7e7a43f1d195d74ec
za7a8d97e6b598b7e64ca00938171ceb03adfcab74089cb1cbb0071ac14f4386b80a5b915b001f2
zebe31474a4ff90200a828e3a324739b838e3ea778c1a2312e9805ce976f10d6894b6c24b2d98f0
z98d50e6dbbfa79ca7a7b188f3b3f155a0a425007033abb97c9729dea0f623128656302f3de1920
z0dd520410fe1e0c4f057f64d3be8746bcc21df996c021c0e1dd0e46693b4b5ca92dc6afa0b876d
z379f1048b5389c795a3a25591f8d5303ffc57c9412683dbfe926e6c1d1966f73bd027e3cdc0aaa
zd01360fcd48386a74d07a6be68b1a87e37f0ed96f04af59b420d691a5d526219be1441a26ea656
z9cbfb05412e89cd06907aee440669954b62561e9ce005ef471722daea9ede5dc0901429f9f42bc
z8b856a9029455f2d23604959fb8ba3a3442ae5c8f7255acddb1f2e948b41eccfe7669f18a8a6a3
ze6a959067e1abbd7b85cdb528d226b60b2bac7f9b0a3a873d523e1b5711548313acca9edc2b357
zd24158aa192f9d56212785e7e7dd4336bb3f18f64f8505adc1ca7263a44290c00ab1ad91e9fb88
z2797dcdd03c1e2adccbe27714f4ce44666101634800326b9fad4ec7da0923613b92231925f8e72
z0df938f2c4903c0c28815a4ebfb369ab7c064216333f01116a24689659d8eacca86ea7c8d44498
zd494b5e3a7ba451c233b5be97f62e4a2ad19775441418eb28e1cc9e8de666383dd7b1bbcd1c84d
z5e96eeb27b4c6a591d9c3a22bf3cda7413639449a578e6deaa0dd68cfe263e4feafac4c50df6a2
z959a63f7913c864a502ea30e22e9c749cab7ba4bc22942b2d46a4919d8b48e7d5752943b5ea154
z7b1cd4283bfa8a5b7e28f9833469676cf653843509a203a6afa702d28ae3c01a295ad9d174ec67
z38230da53a9cc1fe6f4dcf5cbb661ba69aa3d4b58d62b4c2651933d029b22e63ff2f519c9bfccb
z79408bfbc8494a7e611128a75c9dd4ae2787eeecd999a0b82bb4d38d4179f00b792780a9388a3d
z6b0108aaeea1a5fdd56826ec054b7445114571284888ad468404af03d7baaf0de6fb14aef16b71
z16fa9321ecc3451ac69e736565cec32d3c3820048297fd695aff1dfa90a13653e37700e47aeee7
ze020beca180aa459562694f226d9d1a5ca822b2404389c56363354d259d2f7331526ca9078c28b
z47b93896a5f93d759c3a5efe84158cbfb3905babd89af2fc03786942de2cdacb9fdd7a867ec3e4
z414a87db27d5b52945cf297075825b2fe75ed498aa0f11dc8cbc7cffde41145d7474b79e75f89d
z78cc48056cc8dfbd8adc9ab9096788dd1c7021d47b5a971426c1930a0263b400240476e3c00392
zd4dd60008f17b785d9a02081a26d7de417ac7ae69997622ab419b38b0b4518906d5651e85a35a0
z5dedd13e3802d2a1ccba3524b723ec64311751c83787f0b4c59d4df1c33b95e18105e39f01818f
z7d3cbff883bc5844172a94e8c920ac5601fdc40ab14a569cad50d7b9d2f117d5a730ef472b5466
z85e60177de41d0eb518ccbb7936ad424d479611e07ecb1265f8a4c52f09897da2f7fbfdd37b97f
z126241171d4b170148f1a38020f1eb3f09ea337f34ab87c314635af671c5f18bf94e8868d50df1
z8cd10128329b8d80a4e706340d619d6ba7b4a6240f413b638603ee5259e65360b5f0237f3069af
z9c1b13f18c58d81df5ac967234921270cb364a3a6b6275874ed259765a9491b6c89c7fd91aeaf4
z9b0a072d83440588d7aa0d0e157dbd64c064c2df791d1b0cc0de286e8585dd70c4cba9bd8cbede
zf0a6049b926bc5606db12bd6a04a29c8c5869550254fc0a27c88d03b0683c14295fbc77561af03
zecc3b0ec3c3a552250df4fe109e162030795d8627c68dda2e55170b9edc25c04873c9c27590976
z4a0e0917de049668b9b6d3178efbcbba984168ef1f55dde57bb271eb47b5ccfe454d36433ce988
zffc42ed6f239588802b3569aeb7a13498a0854926eab634e9e11b1ae0c366114dc50fde65a3cf6
zeba993947a132811af4a721fdc6c0686cb3ac4a55d8e0caf1d72e35020272f095d60530e6b7375
z3da5f643035adeca3d379d2eea23515f7a602333caeadfcfbd39d5b631e0d90baa6036bc5f3b75
zd3900541f2b2029981df292413790983dce90b6b8e4a20d036299d7784e74161b69dabca30d8f2
z09d1533f504692eca680966e4b33f67a24d4b9262d21e4e6854056a32a3746f5ad93dbbccd13a0
z48c95b6fa8c22920ede095ef72d80110b7e5ac428ce2f2f9593f82bfefdbab7c49427a3d0a4a15
zf1c62bfeb57e64a99e80a7ade4bad8935108d50ac5015b92b059bf08db2fc3b5b97448e2536cf9
z0c1bcb53a11304259d7a8488cf4cc18a8c59b271ff6a5d023c4a2ee40705b0f38e28fd2c45a1c2
z02dcf127e6313d056b2ea8d3f96fae5062635ca35868435b0c955f4e6baa40cd2d340c163d9b57
zaf872f750233e869dea3f17a5312774dc8b0be7e7d3ad0705e7b61fb3a7b4a3d5205391e757b7a
zfa84f900080b6188abee9bbed8f6a0ec8ba57bd1233e4af442d8de94933d9c2daea2e669324011
z15c17c6a530ef71dcd43676a9cbba3590afb3320c3d126e9b0e4f1ea7fac2fd4faf0c18adf7e45
zb560a6e9a6fac8ef40ddda3464c99984ef63c5a5a8f000f9e860bf49a1f22dd6e1e8d51920b666
z146011006f68961d58d96324f17cc5b56910b0767db2034620b0dbfcac1b7f8d92da69977e6d44
z5c685ca9ddcd454db67592a8db3683a3a655ae3cd3780bfa6899465f85540f106b218ffc1e145e
zff2d2976fd7a92bf691055b9db27a7bc0c55fd38c3e063cc47c0956159491576e98797460877d5
z5fd027889b9445a6dcba5bbd7beda820ec142d27b70c8d225d38c107964d3bea41038c6d20d361
z013e260931cda9a2167c0cbcb0c21a7ba1ef53c69eeed142e18f2dc82e3528e457cc6296a71e1a
z0e39ffa6e715b080d7b12257e46beef8a96963da83b8e35b8000896d6ac12b1693c12174e8a397
z9cee63777787d695f7144bac9e1f366bd2c50bb1739cbf306c30ba02121246df57be25c3d134f9
zff3d2816d01e09bb314a4e04f67c578256db43450baf9b1041325ca992158913efb5e851addf8c
z23e326eee6c2e80f6a043f2e427db3219555e3f8ab18d127f2504f95fddbfd9c4104511a649374
z1bfa1537e7d319773a83135fc476a38f9acebda3ee9e6d115e83c64f8d7b79109999dfc14ffdc6
z0097c64c6cb43db808b10de576af7cccd1b8dac46ef32792f70a99875a343f8b75653707882be7
zf173b808de5cfb2c60ce648b5ffb82a70a3f4ce79ba10f075ffbef94a3e2425a45917804af08b1
ze9d2f5f18112445da0e45a13f82bd044b6eaed80eb648f4c9ca5ee11f137fce445a3eb545bac9a
z2e36d1f851af305bd7ceb0b4665fef98e344562c6352af3a102646810bdbf8772f73ba5947c96c
ze17c778d7556f1445e0ceb31682f4d6e24fd173e6ae0419bec2bb2af9e18586786621e3137ef75
z09045ed7abb6eb3e46623c0ae65b48510b469da96d56d32874c008015309a60565fecb7292f6b0
z27335b1cae919cb5ef725352faad92a145bcbf95d38500d70a179bf550f6f81081ad2d74dc7e69
zaa6bc059276679c7645f0423e1945316d292a42b6e36f0c7dff0dabf9fb03b8d1e1c3aa48293e6
z521b2b08c83de113c4a91bf8a44e7e55442d5d5e6858ab688bd19fa073ce11aeafb8ee599a69f3
ze0d0d814710234a48f631f59ada65d4c29604aa4f43ec252c6405dabd43990725057994dea21ad
z15eec707cf25100fadf4f502ca335a774bba57ec1927931226080eb1678c195e369996347748b2
z4cd29b61befbbae8f7b30ef51079b9de26fce0e16064386717fd8da937436f64cfde407c75b119
z72360c1f4e928d80e885c4fc0290da841ecd212dffa3dc1604ab7d1ebaf716e745f76017e44b3a
zbfbb01b0f4dd3bf71ef137fefbad495ca19679598fc4df4de0ebc32bf32504efebb39a9a8e466e
zd192951b57a04fd8c08f1a35a157aabbc17e4dfbd7550eac2b286c774fed5f511fda52593cb433
zf532fb0dba40fd0d7ae25c85b3cf5ece16826ea08ec727425aec049378ea1643887eba319da89c
zbac5fd71f9daf164ecaf699351293023fc0a78f2cae0e9482f83f43923a964028204cbe88e65a8
zfc498088cdb7ece9eea2606a6702fda682742de1b00a4d6454433c244fa166222e48b8d1f803a2
z21296603e018d686b59e1df032d9f83f8732d4af5a5991fa3cdfdaaaaa8a8ff6b5296b002d2c97
zcfbe7deffb220a6fcd2629ba9d5d756f55ee66ccc56e95accd30bce074b17d5fc548de206e357d
z1240196df9474fc80a0b4f02691d26a93c4ca3e1f9bd7d836ce6a67aa5fb41c2f8086fba38f9d5
z8ecc31add3080e6781b0546376e03329ec114d48e55f590435c61670350abe487da607ed39da38
z60eaad39c8207a179d386cf5c880ece5827ff309c6cbce647dcb4a4b2554b0ed2931b809e18f4d
ze6f3e7f2261e17e86cae4f2bee2c440c9e9b0580c471af04d86572b934482ceb5071ec0740839a
z58e50b1cf408ff97564256e945b329ebeac5201e923f91195a203ebfe0bb760439a9336acc3373
zb95f48948278ae008cf25d643a051408243eceedb71694e058302654c2aa107c3e221fe1d131e9
zff9883cacf7a1ff116ce08197abaf42b93357ae463d3ec1b387081441f817b4404a3997a5f651f
zabbeae63666cc15f8785c7cf6acebd003e143ba539b2bd748ae21af98791b9fed9b0752c53eaea
z1e2c79da005ecc856efe258ffc6a66fd5ff9b315c31f392765ffcca5431006fe0995d7d4a3a8b0
z24a9c974ea161016df7dd451affc1c593be9f9e13485f26cbc1c0d67d83bf00ee3db6a4801a088
z16b4a006c55cf7e2346742329d605016e87578fcb8d9b38e006bb553275ddd7d7672a0ee200c11
ze91eee871f8b9b9c100a9e98dc55caeca5dd675916b16b1096449113ad0e6e9ca8dcb2de241b2a
z93e49fa3bb322160c68a80e5786a46ae6a9669c33589021cb8911e494afef79e6fb21929080fb6
z57ffbd6df9e3b5a8bc7caf914ee0e65f28f73f60635a3a6438a929ab0c29ab1692be8f3a853424
zb46b05bd82f6c7a09cf439d72fed547aae58682e9bfd80f85f2cffcad9c4e833bb7dc0172663ef
z782654cc6cf2ef5d3ecec434582c8a3e80d19ebcfa3e39c2db970521b4d97dcf6d8d8e80c25bfa
z16ce4e5d8ade2519dd6060360799a5fdbf8f6064ba3fcd4578dcb96c80b2ec267a7536f728097b
z25c450d8a5eb92dd709a65213d3ec58930e5a53866e25f375365f22df3cc1503b7de2fd2b7cf02
zbe68d65234a2068d8c605b978dd3c0df07a6702ead22ccdf3b980b17d343c11355e8c6378d14e0
z288a7c2c2c0161b54a371416214ca405400393a50da2bb440c8f23f9ad07305089ebdf48d390db
z0bc353f178d67dd452be2858e51e25e51445493a4168549061a25e3082f8c21df4802d34520fdb
zf2654f1d487ee9056b4644f418f63c30a4bbc7f53201d110cdf053cb4643201300706932806aa6
z73f9d16adb9e058521471316232647c9acd2ae5a09d9a6535697de0ab9eb2468cafddd02775515
z92e6429918538caceb722748de9b885f4f710fcdf8ccd7d4e7e2ac2d25baf772b490664fc14e40
zc5cc7bdb027115af48f201b2059db9967fabbca7f561a244feb1e230da9f899d211b3be9f121e1
z0265cf1cfa1ebfde3b0625314ece3d7d30a030f4774c85f594358e5c01fd922099db8d7da78a0e
zb1d43b048adb03984a529841256d9f6231a758270c1a714439358966416bab81344b3a792c71c0
z902ad3d52b1f54b6c7241e2d7763c7b2963211d3509f17ee1e239ada79cb7c37ac76720e9bcf1b
ze34c620736a192d78e00ea10c907aa0458e78713cfe1ffcc66ba89be0d5565c5650e4f9b56fb53
z6785a689db12095161a9c51f96410362214b1d496042e1b7ca259daceebd7ee2f0f8880280c044
z664561587797e2c99c6941641b366b5a5bbcfabb0334fe9ba97612442f51d861002888984a6e73
z8b0037afbe9a398f37ac93438634159a5f3a5ae8e40ea3f5b8f1bf69bcc619cab3dcd8b66d1d2b
z1d30906cfa2a3c987b16bd3fa830d94331dc3045bfbacc7fad71af4b091aa739efb9ef50306da7
z3c3b0239d048d2a9840b6feac0a29115c5ffacd759cff1db830593136272b9da28d7873646ad80
z61c43ed691810be23c7bf9c4614b1f45b306767ee4bae2c6ba919fd6627fbae26aa1ef6dea230d
zcbe67fc11f35c4ef2cd8d0c2278df0217e92ebb2f84d902631ffa89ac85e3445a925f1e1973baf
z80079c8cd22d53d15553133e686b4830af13ee4d6353ec8fef80e2f9c0c26ad14f1838028cf47c
z7300f779484cbcfb47a41b20f5f659f9a6028ee2f44fd1d6a4f1373c6bf7825f8c0fd7268ccd6a
zc32290b1cb1f64398b17d520fcf3ee776ec784eb21590b5ae798ee722484d209ee52c5d7a14708
za86dc9dd66ee1c378565b02fab33c009abc935fe3712a12e9e97ca264f87cce1ebd7058faef0a9
z8c9d76609205d301c2c2f032aa1193c8037a087e27e9881e4bb7711de5b2e15c8688011e10e5aa
z9dbbcc46f6455fa6e87b6d03c86e25bc3143319825ec276fe30f6d603e35a56d4d32bc1ddb4b04
z5eae687c9077068bcc0f17433aabee19f450df51292d1cd7c721558c02206e7f4631df9ce0ae14
za9ecf9144bc5c30a17d5b08735d16b39d367b10420619453f172b55f7797e8f6649d5d49a8d419
zd50727cb181a8aba53c29220389a6d1d6bf5e2d9b160e70ec8904da0a861ec39add22d7917bf92
z13ede867d197939769c66bccdb805f3c9c1016d62998646ccd5f1a68f221f0832f8c1519d18f27
z762a7dd3f8c774ce5a21b9c378c4b0c5376f12a1bbf19d14893a1b08045806c5046a532ae4b06f
z71c5f2b7dad0e4f4e72e0cf95989c371537bad497bdc05489c0c2d68a1a4175a5f2b96448d7eb4
z9f49ba1104033c35afe8e14b579e56bbf3e60122a47b52fe49ab00aa07b15aee00426d61d98eba
z902310a2bc31b36dfc1e407d9ba2fd6bccf2b8e919477476ed6c6c6c9a70da6e47429d32840ce5
zcc226e7ec251c61682f1355a5bd3473d6239a0fa1fa81d3b57c4e7afe9ed1fbc440634460900d7
zdf8e82e30adfc8d99a612402b01ba5d6b7833327723a74f23837b26c9cdb298db2db7828f33c8e
zf444fa3bb5c1b924df873c12f2279a4b1fff9446c43d44bfc9b127def113bc19ee8a9d12dfce04
z8e3271f8758829fb2fb0c67a0917043ae9c5b4c8a60a1d643610eb5d753599f4fcf6b3e63b034c
z7e0a6468f538efe9a45b86924685dc89b6cf34fe54d5be7e42a80e1d8300b47dc4b8f883e79b90
zd56a0dfa548cfd29feea2c188d174e6bc0e2efaac1127b0b98eabf190d91e7650f76abbe90e4ec
zab3a2ff06d6f83146cafb80bb10154872e2d66abd7a2683ca5cdcf1f08afb1fea09a812549db80
zced8a6768750fae4420dc61cd7968e318fdd9f6df581bc195e8cf5ad03590199434b027b05a064
zf6096b5695f4c102b0f2859b93d27096ae8e020f967f6c37bfd89b0efbfeb74dfe10bb2a88d0eb
z8710ab15373088f6f590e2bb1f199022a0ade6392d82213f18247d935fff5a3df4f5422f45e661
z3d23970d626e0f00a45cf2a69cacf80b2d47f06ace4a80c41fd5e7bfa5bc4974b9637abc76c606
zf08aff4f091e38f93ba61e21ff0a7fe8b5e7034c782e530d4b03143790224a3aaeef856c01dd7e
z11211c50ab54850c4846fb4a8726b41542e42f199fa04825f846fcfb2fe1bf805ab0c94ccf82d6
z5b481bb145b8eedd85d1cebbb9a518dea08e37fab4ce7b2b5642ee1dc3aa45487bffe9d22f24e3
z33cd8ed78612afee36929789afe5ccc248e4aeb76a28e68030d15d77468ff1bfb5370e19b5d337
z43db59494fe1e7150d0caf4087f6eff9f30ff8e97c187ce70a574f40a364e9c1064036c933380c
z1f8142bb47055f0b3cf15047e6de4bd101911fe985b8cf249b81f100c4199b397a08ee9959b84f
z59d31ae685480de720ae56fdd6fc4704d072f1b4ed5b6a33f7d6b556388a33a498cc336fa34e10
z544247aef5e8f3b570db1bc0aaaa32c54180c4e40f4bd36e4ed52d25be4a215ac36d8265e2f5f1
zb778d154a46068688472e8c89c09159898d145fad187133790123971a1607bbf383e501df02ed2
z6b3ecf52dc95f14465d6f68a5e89c3a4bb6dab0682eb40e6692cf85feee5274978068c2c8cae7a
zde4f84a2a353323f009aaf6e31ed69f7d7390f254516063b485657ed59fedf233c40b01d2339a6
zf3122e2f325e8693ff653ab1772c4f32a4537013c5c6c6e093d3504ccf9f58171a6cca5061abd8
z5bc359e42c7df9872ccf9652573170b976383a41fbc5f01a05b6cd61b460598122a3504b520457
z1257aa156b473e0d76c3c8f5b574b31b235e38c11829aee7b574485dafd1924cc1f18184b41581
z22bcb9c9af693810452009a3539b995f24a629aeef159f4724c00fae6358edf9afcdf7f3b7dc3a
z20f357d9ac9c5a88016dd544965b2468cd3b96d7125ff4b58ce2712527e164cbf5f322119724de
z4dbbc647a2faab1fd0dce4aed0666ea3aa88da57b9709b1f183103018911a827f6a5f37efdbe6c
z158b1ce21b1cdc285d5fe9586042b47b0f2f630817e08107b6134832309af202514144d6f3c2f3
z1d3fc3f3f17cac8f7baf4e2c0767b9e8df457d1841d119838e3bc0f544bfd7ef61648a3a751dbc
z8c88af4bcc58e7d152f06feb15a3a4f2ec2228740fddb36d728669be9512cf1fd12b91f7655592
z46cdfda54cce0f83d2f8cf4b8cef89862e43c3f9763d29cd3f30e7eae5283b985d3fd9b46c6caf
z872adc0955cf72351c97c6a2724ff226996f82180e9fd4c9439f8fe39a618f571a87d0285cc03e
z95219b78ec8fd26b73c8ea8ed4724787d7baa44c49a5bb0f1824f5ddffae69ae6085ca66543621
z095c3879c90f57c404a68d49d5d7cc9085a1b6aeee84ad83ee1370366c4a84bef2a7d28b3cb5f7
z485af2bfccf7082f4bae64a744d5ca7116213c435e2251296ecd7eb0e4202a6588b155593bdf55
ze7af712254fec189860fee999e77369ac37a29c767f2f8e22f105dcd7ff21b7507b3b5a44742ff
z2d90449e575bf0c5e2bce96e812dd4553d3e9d2936cc153ae57bff0d63227bc695f3d6f6298150
ze60f861e9e372758549766cb2d1510a82c408b60d008603edec59fc4216b5a22bcc058e37faaad
zfe5e373a06b36b66c4b48e803cb607a90be0c1072e4953ad95341cff159a811dbe515ca6c53789
z1442bd5746d58ff4e919d56e3719f2f3c0793d2a681b0e7879371f2da8cc997d7463d26d93b3ae
zec808cb6db79fa801b8bddbd28e6139071cac51c66b986b2e489ece21f66540f02fee32d7907c7
z58d19ac3963076cef74dde51704ff6783f72379119e6dc23c56093bd10fb0b5509219abf89dc5a
z7e9e96486d3391c9bbc1f634805156910131ca3cf659d58f88a6983f9cdd757a086f295d6c2d0e
zb08de25826396c0597e1a803e57864ba3a03aa7c484ab563268f83303b933bec0b6df2d184ab91
z818f89f16cf4c75eea34e5f968181d2bd0909c2aa3adb42f9f26383ed96fe61a50f7f7fccc85c8
z7f24899bc6aab60ea3b537d49538721df893187399290728547921ca3e57d7b67197c8982bbd38
z03efae466db0b435ab0b0c3b7e915f7ae04728cada98be5ad83b040c69af2f7aab106b0e52d8bf
zc8b0d655830ce5f3ddecb9805d7b5550c749204423859231b2e927a8d51f14ac033a9c15bd8387
z1fcbdf9dfaeec851a119d86c35fdd9849557ad76dae958f124a0d4c1afe457ee49a49486254cb2
z525ae4970e5a8e5e47959b5f0adfee8f55a44c5054df814d2dc624f78b8fcd8847e0a1c9524f6f
z0598ea68147aba170d38d37323531dc572ccb9399d7918ba6e021013c5ce58d8ca12799d97fdf9
zec95b19c92d8c8c69ca9c402b80f70f100518e77c2f6e7835856b0c9c564f68cd2e319abd5371a
z54d06296e1488c708ee1745c319b7d038cebdd8e810c379304a0d63ad7e678620438ecc6b33b8f
z12499ca666b216105a93fed453d63c69162122af4113f01e5262ccb5f77dae5fe75bf9c2f68f5d
zc9f85b03243c8f2a36cc3e9cc3c008cc89fae8eaaca6f58d81b0bd84f17aedcb3bf360e0eb4356
zd27bf9c72ad7494eda6909eb772707832f8fc15278ac9da60028a9660167c1dd263bb8b0c1cb98
z54ee6834b5147c37a48f2a97a43839908273ac166ed7fc8ecc2a0b0d9ddde75d7938368c752e51
z55aee51f73e54c6eedee9765957c3ac9501f66c8e486d163df1b92bfdabbde8d55cccd3248d885
ze5e4ee60b12934bad55323ddba87a6688aa239bd15a5ed47ecaba066c374028fcb739b6ca85459
zc60d2ba82beb856634b7b72a679bc34df45b2d549217b9c71ade86a1a90a3e73d136a55e1daff4
z5b666216e065336fd4641210e7adf0649fd9ee1228fb1a428b74ab0df11c504ce3e5fbe8dfe1b2
z08a715bda88529995008218dd20da1a712555eb1b4d17ab0d1e123b89c580f1da8725916fa2805
z2bdcedf19909f991c2f772409a67eec91a33a44c6e3b14326a0c79624045ccf0488aeda0ce60f5
zd3703043fc995876eff1e5e99458e82c70d454acac44f4f617124989178393f22cb62a214f7834
z3bc98ee69b36324045e25a24635189de7cbfa5b5eeefc2de5905faff722c53d5e4447e71ee9a5b
z913289749aa78d1e074a2bfe51d8112266b245c08f9db32377961ea3106158bd88f3aab31aa0d9
zaa197f96b3f46c6c5dec908bd63636a6bd7e9e27c5dd90e13457e7da38303436dbfcccbf93bbd4
zadc26cbc26590c177d1745fa18fa129a709d2fc84ce4b6efe26a1ab97dce23a80d960ee6c0ad72
z516c0a1351acf5f9f988456eb87c1c28ed275b9704e59f7de9daa9a3264ffbf80a3466e6028c34
zffa03fba69dd857179a8b68c3200f59230e8d4bfc631b7e13ea7c47b2ddd43a8dba59bd417f692
zff6eab2cdda9ecb74436402c4ffa0708bd69fa15375a71a9e427d7326d17172f2017474b96700f
z0f40b93eb63de990500a5f013aa62c0668a2ffcc1134906565cb92feb99a4ea746b36be51fdcfc
z48870cd6488c4b14f81003e688a91b62a45e7767c26f737564dfe533179b85b8b23bf9456ee2a6
z03ad09666c8c488bdb25dade45cf5e37dc526b34cbf82c3db942d118ffbb5ad1d23c939c362acf
zc718049919236c5277032ba76e00a2b71a28afc4cd1415e05dc6a8326933f8116333c4f057c846
zd1d9dee961204d316cb1d44f014903e9017297830031b0ee41a63b3b79c6322b3e98b92b472bfe
z45dc0dd37716054256a8b68e533cfb68229c56052e3fb4fe097cf992ad5b1966816a9748ad0f09
z05a4916728f6157162b927fa9bee04577106f58707dcd4d24c46ddd0c9bb66fded22549af9375d
z4af11e92be1e17f6bb94b1977346bb4bd1c27d5649e39de4b2f5d6a41d5d5699b81f5c97b3237a
z43e7dda350ab328e222b3e3d1e58f527ea449557d89c6829b92ea3474a7825265bc9b3aaf65161
zc2955c96a9a94b46b0c46dd31c05e839d297e3fa2dc9bdfe1156b5114f19b8b30ace349803bdac
zf824b19cfcc632f903342029a36ba8804f4f6f3fe07108ccf03366d78217d8bb702d34ca530a18
ze06dfe33806721546c8993830e21f04f32d8c6f40c5c80651ec9372a5af54d65f63aa920bd4af9
za61f568b79dd486686f31379f2d26cd2b5a0c191b44e5454e5ed1906e2e45c0ece8fdec73646eb
zad5aee92a4600b0ec518585fc3b23ff36a99b1009bef6b07ded664e0b79c21f4eb408a146dacc7
ze1bf387b772f3545dcfc518bda6528a6751c31aa8f56afd0196187fff4702e048f2e84fd3b7bcd
z848eaf27b975ac9225e50ca3fcb99e0185e59363a3a199efbe4e57910e9205ed721f482d3cd80f
z64c0e6fb0f3e57ee00b2afdb6d83e6b184f81e8a5ea931425747bfde457913a3cab4c371d06149
ze7ff4638641e85ba6ee00c4784fe9b51063f430b6c4c2dda5fa71dd908be518711148e8078f482
zbd86f8f8647d05d9588417f2fe5688806f3cb05dbebadcd1d2aa4b7ef443f5d2dd295568e191ce
z9771eb37da12ca355afe7eb96c874d414b2a1f8f0aed661df367b453f035d1df1d5beaf6ffa3bd
ze812a4b1765f149dad2812ffe31a3fc2e55890378feab308118223a83401d16513db9403675aca
z8f8086523dd443903421b7509daa16cee51dcda646e5f77cd6dfa8522415d26698736c163d62a6
zfb630d634d65364d94fae53be833e78c72cef2261112a0e5a9b1accc5a1d4a0a6483e6ca90dfb7
zece3a2a0dce50126c7d21e9c6e160874ad36bf3e7ba5e780fecb0cb5109337b82950296df9b498
zd99d60c723c493ddc83d1702be56b9661d8ef7a06b6cf2cf349cd2fe18de87249265b6f7c0d8be
z2e351d0105618e2276df18dd4b8f3d90b96cadc5196684f4b02e4c05ac9aef5e7f257f72bea8cb
zf0113f454f1bdc18928f8e609023b9533a20e7a6fca763561bed265ad9bd951e1612a599b621e1
z5f4c02b2dee7754ff8227a12cb0a840ec9ff242920c1a6a5fb8b608aed00c08f122288303a6121
zb78b7c070c5898533652e2cd1400463e3c6d58306f34b20079ed5be39da5a40ee1073efaeff3ed
zb81aba2a0034d4d78433769a3cacf6ffbe9f5af0ee24fa818a3498cbbe875ac9455b3ad4d926b5
z4f0edfa02db169af4abf5a0c7dc6e0fbd3bca45b9cee2ac65a8973da47d5f938e85b0233f78624
z05384dce06e980d38335040b40a262fd5bcb84feb591cf483dfe6798a935f0c13f644eeb770aab
z382804aca719f786d8ce09fef25f65a245330afb2c278de074ea6442fbc7d0c157ac72a6745841
zf61b056d2888efeb2fcb32a64f852ed9af94202ddf17da423c153dfcc79b84dc13ffaba3b9c4e9
z24b45b10190f53649c8281468532fc5883f6bd9e05c51951234bd02937766e5071233e15f98cad
z2acbcfde2a7af14d4bc147818b8bca0aa66e60351c94bd08e733c72ac11656bcb775b658a0536d
z8b30ef1e1811b009d2696d4b2f483d879dfe34a9981b826e170c1b74cdeea2a4374926b78f48ca
z8ced9ba7555c5027361bb778d4eaeb4805338ed06898961ae957769331e08aacb7c0af1beda942
zdaa0beed5585e0d7ba3edcce357c6a798ebdb69e9cf07fd904f6ebaa276852d847834ec62288ee
zc33e0c3063185887294b46c8afa4d231108d74ad63b50787bc01214735e450ade5d6807da29ea7
z45b875d5b8870ecfad73bdbc8f232f32201d49cd5694d1774fc065a45189cbcde6b32ef4b2b249
z63a06e666a0de788c355c2006f6c2c66c5c215d6aea93c346f6eecc2f1c973c43cd87e5ed07578
z9e750e63394de707b06ebf8bafb6fbe5560d43a8a797c6b14366e9845e15b50b51f63f39f2cb40
z88e7a418138ec65586cd7e85bc7ed67b88a9d9c791ef04c843ad90d8e5814c295de26dc7805952
z7dfa789800400f9b5b79b1a39cb13346ee92ea3fa05139e008440c2751301a8fa3be90b442a2dc
z05163825ddc8c86e482a4ab980666322867cdb028e2f83adec9846c9e28970d286cd03a1d158e5
z374907a5f5b7027f9608103601e7077bb9249b3c12a6f3e2b13fbd51a4ecb047a064f318152df8
z51e5cebab3a23a2fe9b39563c5177cdc7f4ad89a52f59c60fc96d11f8cb00cac101f1665a4f571
zb74fe210bdf7da13962a31fce7356da89b14c845d58544bd1e8681d9c78d639d8f07e198d4571d
zd07511d4e7dcb6676d2df71296e453316119cd02077d7ce7038e544e628df84bf301af3ca8f078
z068f08a36797406fce7503fd5feb7ce6690c53860501f6bb1dbaac719df5e121c819e8f4fda0d5
z022bd833f5d59ce67ad85a1ab87ecf1050f6ec3c02bca640a258620563cdcc36e881eee8f16e7d
z2ccd90a73a6236c2e97a5341edbdda20f1a65da4ec433a9fd71bb4bdd08ae176aaded65046dec7
zcb73b87436655e81206bb822ab873d1f92ba39053645289f965ddd347a1f8012a71cc02cc052bc
za3dcffa6acd4cb391ca71d1b4b3148f5c983d28d366d6c2416ad0b705feb2135492975a975a930
z3819c5fd9150fe3ae30dd08fc7c4fd712e0116181a5989702a7c917b9d1c4d47fa3d7098b31a18
zdb946559debdf2d213dfd89c47c6ffb916a1f1d604070be9cadf5fd758d7f56d656f32aac04e8f
zea3246368435ae0de08e79416ec6463308658ed4b73b31ac950ed48de314d3e77ce070ef4d50f8
z1fcf6360771e63c38a0f13ed0e9477bdd766ff6ec0ad88c26aff69ee1f40ae010e1afb974c5ab5
ze823695949124c17f02084271ea6228ff8fb3e2064a5b4ed347b92c8ee4800516a2ba7fa4a5368
zc006010e447890f2670445d810a2a7a659ac526ceb840e2cd873706a85a67f4a4c6505d10ff31d
zed6a6fd23a3d03516e71f4726af1ee70abf99166ece4dfc4618b2e216a9f16a0015c39e18ea506
zb7bf6900ebc31955b5fc035be3cdc0640c2d88e6684a4ae8263eaed8461a3cd932f659028b4eb3
zd7a8f2ef1946ecc34e962d0ac3ea499c4f845a509d5ea641ba5ed3f10a4e09bbba1081c0f20eb5
zd7d790c282b3145ff6fd7ea392c6a49f16284354e0cedd853de6803a78d50b0ac0c3dc207d3adf
zf44452d0cba179af81ba510bd9a0b3daf310605eef255d5e2760d47bc7e36ac6504ca2f0b74cc9
z4fb14306092c7f2f9b30eaba9312db2e50d5fe54904b4057e5545e8f9a89d37120983d7dde5fca
z47c8daa74cc28211b68a0026c56fa59a403bbf4ec95aca258be147ac88fccd830d1bf6d54dec29
z355d530a918e66f83b3bda5d2957673613e01dae354930a1430b1b5b8e631f98d0ee7abf0558bb
zfef0f00964c55d66bc51a2afb2a3dfa9164ff36d8cfc916d07723208c6912d4a460a2941a17f3c
zb3aecbe10b8cd0c01746180fbaaa4642000aa08a2875175a21fa6aecbffe54cb9bf1695695b0ba
z62b9230044c3de5f9b8dac1bd8efd42b83cef8d16e4da677933a425d2e812068f172917375f502
z5c12a846163f30420d598d0436e115c1d322e67930df3a12d203bedefb573619358ec95070cd5e
z3fecbbaa526d8c05813cb34ee34ca9dcd3e9bef5b0daa5c4b6dc6e9b42e43b96ab967a0714742a
z5672a60e809e5fb536c572ad05a5eb082a058f75e69eb2c09b2da83b01a90a6d9e865bf85b575e
z2ed86a7fba9c6a8ce837aeae5f478a61cf4cda331fc1677e4e6c34858469034517aca1e64cad82
za0c07b1a9f811f4671a65c18b140025ccb52e7d8e042f309528d51cd32be29e1b0ef3be078ca1e
z9d0c0510f6c6dff7507f4ccce396b141758dec79dde293e866e6ec31bf2796935acb77fe5b85cc
z428085ac24698863eaeb3e6d948f3caa88b17121a9115293192d255050747c246c9dc92828a921
zebeedeec25c2ed29d6f5223eb62d177a64bb213401baf1e34c1209877fe1296f7c1d3e415a86ac
z712e2469273bd09d6b5ffed380b141ce3f51099a3a0f3dff66ca181661f435063ca9636f4c04b7
zef29954e6a5a439014c4c1062a8f4f15dfc166c430fc566400a889c2b197b52805fed407d30101
zd1a10cb92dc1b22ae7727b4c344674ba0e2f98b54c74ee97d26f2096b730e2d0cb816590e684de
zef3b8371750c3f2bb3b7da722f0e0c907de61722f800b3b0bbb88e17cd2d25ebc73c6e1afaa778
zd025e823cd011eb719cc76640d13519d505597c7960922de2027a1a7fca73dd4edc527b7d905c4
z18258d57ebf65b3f2d38a196ac91f19c006f22f0b8e67fbe58956e06af2822e88f0f6d91d70c18
za51ed52c0b0588e09fff5457930f9c0a7edb0eea10c007c9d07e9863cef4d57d95bfea81084335
z768a9dfa40fdb64b7542f07172895131d930fa1974f9ab0d00d6f70714837515586ad65a8b4e56
z9ea98e3926d5e003fb5d77b15128cfe9edacd24a47b726bcb3179040eacae3b2679d02a1313eb0
zfd6598d8d9196ae5912788b28cb6196fd628296b1709d730a2089eeeddf57951d93584ff0b6035
z1eeffb2577914271d9598018944cc308d276525ecb783f4e6bd3a444bd97fc56e361813da702ed
z2166daa4507481e3d344c52a4cb41d0c5115f0dd3d151e5a4982af3de4fa5a29b4cc97a7ed5b8b
z6fbb21ba43d55e05e6fe41999a0ed247aebf31dc8cf275e0ceb37ca987d91f1922a55c4bdf21bd
z7dd18079b374c3809d216560b4de9a249e0ed92b3eea968991f6a92858fd0cde9a0fb95cf26050
zbeae49065ff761864618c9f304fd7c8e5b528c67bdc114188acab59e8b70eea8c0d9189eb9b0ad
z455918a93777c972703410b7f08127ed0dfae5e547ba84fb49f481b3fff55271167d7d714f7567
z37c50390e24ca23c082d68e89061d54f18350287c49e31dadcce6a5ef53121684d21ab5d2c6341
zed5ee067973dbad1212c954c200bb058fc07b2255b123f1ec286e03e5c97eddbe924c92e9ada8c
z2d2c8a277ed6c3c303e7c7d871ee6dc4017d54546c2caaccaba226b52800525721fd502e6f18c9
z0639160c4947711a4bfcb1925599aaf268a93b446327e7ae758427761ccea89a588021f57f9d0e
zc30246aba89ba3ca8356529520f2433d0a2929db85f345aca597d2d289b286a0322ca29924a236
z00788f266a35631bac76ef18da21f35a91746a7240493664ffd93dd6db31c6f68787144d1927db
zff80f3d8aae65df44b269fb4a194d975dd2c2914eff954025355f7bef3cb88fa85c07d4249bda8
z3c3cb2a9c80fd9821ab2b3f51c457ef563f2f38d516b6840269a1fb48543f820aaccddf268e9f8
z855d83b4af7e70e11fe63b482251bab674f8153c4055441f0586f54a95c362da4c2cc89655764e
zd6bf270dce07e86a66486591eb114d5a72b8c1090df7f9669e0a08fd453ece0c16f408b958cdfc
zb3e372214cf0a3f3d1ab5cd1aa651a70f8c0bcd0b947832c90428e96ec287f7952799d821b60f3
zf207bb1a44793618a6daee732cf7ab5a0c544921570a1d6557701d2a33b373fbeaf358f5b8ec8b
z52bb49bdc202724f7b0223e30f21aca0319b204b45b25b26d835be0baf69a16ed3ef9dd60ff03d
za85af1d73dba2060bac7d1780e9e4aa27279cd2906303a059f23714565a1ddabc7c6faafbca252
z7aa8646fc21c0c6297098b13ed1a95c34171f14474fbe871d7c6c5ffbfa1253b04c32c0c515b60
ze718d25a4a0ff4d9cf5b95862ea1d063701964e6261302cc9042363a2272143cd64a0d08d3b205
z618dfc22d55ee1205b822bc3689f8218f37fe459f43d5dd1f2ad39ba1a0de586b4b2ca8917d663
zc08be4256a1d1f9fc43363ff64baa0e00187f910a5578a358f8a24467522a32649d6d184c31411
zc6203f7afc218e6bb5c95bca567a5c8aa3b9d0c60000aa02837008ca517ef58cf7582a52e4cb68
z5eafdb4e14701e3fb9b832eff21432bb2b614d6e60169237daaaa08a427d0e9268fcc1b0890872
za9dc6365f4b3f546cf837a8e40a9a4ee71a2c95c0916fb8c5e3a27c0d0ac3410f6cb699861d2b9
z8d4c0df26c397d20077f075fad4bfdcb7e3508d0b9862d2ad7f58bc78adf3e52f3e757a4621a1b
z3cbee16865e5222d61ed0bd23f1033d4c32e86c44d1733e5a18a0503d673d019900c866481301c
z0c36d05cc1c7c9f2215e1edc9d9e2b9ebcd66ffa46282328ee08622255b2525cf0503bf9ae8752
z7fd9258cd51ded43724ea9aee11c0f95053cd15ee3d69100111b289b5bda25d0899e01b846e989
z125b8c5a8cb3595c4cab9b1a4e8db0a639b8ad9fc746cb7834e20bccd3e260adba1e9e29eba7d9
za925662eba52eda960744d3402337d0c4262e89be66bab3f7f5b29617b18da36619d4ba16d078e
z5e5870c9274795f86e10ee15a3c2b7c6159f88c6820220c33145feade6bb3f26353a165b15eff6
z72ade09668b1896ba1e44d14b4d808e70c6b9efc802187819e82b86c6787385f41accb7b7435d8
zf65cb8a2874918e798fc92c2d1ee2b1f57d92ffbc8eb1b2f99ea0cf08777b06f0be81477a59404
zd12bb32b241207b65c79309c98438592e807ff0b9a58f591812d649c56f272f2fc377ecb7a3ec7
z9b33c13ec3642cbd8086705e2f4d3b754972b3abbac450c71802fbc3f61c212005d51421b0e619
z1e453fafca39b99e079ebfd700dfb715ef7cf552d6c7ec76b61bc4da59e366de9f14a8fd8a00c4
z3b1e277345fa669247eff481bc911f023ae9f3d615341598d25b0b5539d5f35cca592b9ef6c22d
z4385fa36e80159d5bb6577122c49af77d3b89ebf15f11d1d6ca1ca522f484f5424e00ef1a804ba
zae9d52d09d81ca88a4c36927e0aeb3b817551984a1c31bb05bcc0bdbeea68709a8c80e1b04a365
zb2e6bdaf04d85512beb5aaf1db6fb49f46026a8a30a982ac874009b16d073fe7e77429495dfb76
z48455f9e9b5927cfe232fb6c60f6e574d547bd6b095ef70e585fadd1186a8cc030fdb25c7b09c1
z67bfa00f4065ebdc7180fc68333eace031e3125aa220cd140c1e0317668d9cab7e691c2dacfd16
z1ddeca7f9a7a27259ab9cbc791fc28349ba003d4172abdd9dcb293e3c5ce76433dd88a34ab47fb
z098ba495cc3e07e489074dc5d8170614dfaea6a6d31a9e0ce77163f965d76accb14c082badeb6c
z6ebaaf3f8b268153fa365fbc199fa71057d2277ed1b9165022cb490af9f922284f8bd2ba51d078
z1a565ea2244d2034ff19bde0f2538832de0545ee10adf38b205dcee0f10d8b9debad3158833c73
z7da15719f4d5a90a21174541ea0dafa3e1f529dd53c13a3842a7f65a821cc2509ded555153925c
z5b37434677a1c9fc163807c3a95376ce8b06b0958ecda48d337c5be92a1acf9810f5c8c0fa2b88
zd0e915d57b3c08cb7b497a3075e8b523acd593872bdf550605917f3daf8c81f36b79f927471f81
zbeac3cb7a056029046dddd1e394757596190af969753e26c43d20dee9f4ddd0353ea45422e7f1a
z22bd73b43dfd301a67b4e367c422a269cda2ee736f57687036a3a183071cd90089c92e0940ea46
z43f22b9028209df0868d547f955d7c1c2e6b8f2489f8e2ac3412d8da9e3add45eea05b6ce6dfab
z765e35114d4401611dcb0953368c7180251bb66a6d025fc9108d22df004eeb02c0dba2b780f2ef
z05217c781b6f6d82dc369b97f0e167ec848fd237cdcfb77174b9147db03f485033e68710c591b1
z880d0263684eb78ce243afd458c3be3d37428531b6197118ed20e847064ad5e485c10ce4bc8495
zd214cea5ed45aa321e903f8cea5a6500ab0587512583528b022becfcf193a3ed8b68acf9f96684
z59decd0ae3e6fcee02c23201c97c83949a9bbb037a26f1adde32a6715cdab45a3292560f76f306
zbb4e81d662e501fa55fcae86348cb78fdccaa17a7c84a7067a1f57e010bb874dc19be1ed41412f
z639954e8aabf4544ff7ac601ebc359decc036e2f68f93f57a040013ddaa4e9c6e73fab322cfd95
zf889ec98d3973b0f7615de81f46d248a74e81479a2550feaf2f6b0cc7b60f5f361205975bda8a2
z2704af69997283e799531a895f102b040de26532d51c2e07305ee75cde29b189005a60f94cd93b
z939d62dfd4f26af0ae3b806be4582dfcd4558a912da467160382f55bc6fdc435133bc3df71c580
zdb072809c46816682793341880cd4dd81b6dd440790e2b06efafbcdb70fe4e58cd56938e58182f
zcd31b3c32f1a65ba8495ba968730b179dbcb1d92eda68b4ec3d7c33a95fba957193206e0fab5d4
z62d1eac9cc023a364edafe21e723dced81e2c15e07b5dc5cf0626b826eac8a97ca7031c23f1f60
z3113cd4ab254c8eeb329e80dd0e3a7ce6bebc09522b0bdb415a464ced2174e27852d3b456dafb5
z383256d6fc0b0102c2b25b4af2a5b6e49b3b6d34cef99a9fde86a64727f5de28ae31817ed00a5c
z3e5f2957265edeeae6dbf15027ea32ac4db2094cc776d171ad60d1f4617e29970961c437faa99e
zce2aafd776c9eb118b717fd02f24560a3baeac77d1c0b328de03eb73b77b6c428aecbdf73c5626
z277a154fdcf9a135fa2b9d8d8b9115067dce4d219894ffa2d21ab25163f7f6a12d8ba53599fccd
zc69818b97da7db2ea0443c0cffc6d87f07bd1c9402a5d4daea61df78105befae35ab656fc1c082
z929ea2a0726f66523cb0c6862478de62a48f25af6ec4f27fc95a1dcc89c32cced56a01b91f4cb5
z4a0ac3b1e547ce34c71c64bae612ed8c273af29efc1925513a266044cdba928efe7c65117dbd77
z2ebd0b88762d6fdec8f8d90939b6bd10c63abd22837a3993e2a16fc0ee7004a70a803621943e79
z208b2b719852f542465696aa93a807598c5b4fc9c8d877845bc7b6e6f97b90d30fcbefc49f79ea
z0f4250c5aa465e36d944082b174ec174ab71bd7ff8e13e27bbc1fd95422754b9e38e706ad8f58c
z1060d79bfe1690937dc4d4e7ac8a5899974ebd5ee453fb085bee21e0aa96652888f96ffd5d4bd4
z2235088f82577db1c03c9f452f8911f2765b5521e319652991c49116840f3f9355355b1ba9551b
ze6067363cec8f615061124816e10ae435ea1a5f78dec4de8841ce65cab934116578bcce42b2b7c
ze1e3fe0fabba5196496b9274c2ce587da2b6eceb8e5993afacbd99a80dc6169f673459fb8fdbb4
z0d7203e2878646f31b40137be15ef36cc28bc44feadcb1926b2bd07c50e730ec155e0449085417
zbed066f35b6096f2670e8fef4231efb95f4c1ab97b798385c61832565ad733b8a71824536d6daa
zc20d58516b6c9e21d22f5ca0a87bef628a87eac131771bca25765e4fe3129966ca93507b657345
z5fa44c589bdde85efa9887bc5dfd019d3b216b42f4eb13f574ecd8ccc12646b866a720783b4060
zf91a5f29f55254512db7ff2607d8710b899f40800d5491bb2d604629480b15ba949823b13fde4d
z47c6cfff5e9a9d9ddb9e355947455279d2abef3507becc192731785972aac67285ad3f2faa121d
z6fcb90570503ee65f2ae3bfc2d519464e076919a5b271c22665b14b327f896e3e6d90ab5471567
ze1b315c39be8c934b56e4943e6e7052bf40d0d59d1d33692ae1e7cdff785c9974c10424c937423
zbb1f97afcdc9b1b91c2f96c294f0c0bda4071843ed98a5cd3838311eb8aeb1c459d5ad26104933
z797a6b233c7dcc9ed550f6967e89b9428ab1ece4bbc76d3d8cb828fc2f3173130a33d9ce7b529c
zea328c3219137ac5279ed9beee08f53ed60fade5d6c6a6d543ae02d62084c7d8988c6150aee408
zd70ff7ccccc6bda186f6e1cf59b3a0c02dde39b91da958bf7633d8b6c3cf6235ae329cd1cf0f13
z9bef1bbf59cf72d9f35c0eb61c278561969f36621598d00f680eec4b61cdfc4b597ba026a65036
z52c36fa2fbe9e370c8f1f8d40b4a9a33cc01690080384dafb60a373820d6cc7f956f564843b19f
zfcc50569c5daa0c2b12ace53026c87993eeec04beb57926cdb93a409dedb1dd9acd312d6a9c807
z4e4d074fac5c4ba50b20e941a02f0084c232da068745c61f150afd3fb8f0a5dc1759ac6020bc75
z366ff4bc02a0bff79302d055497fff42874dc6aa9d7e22bb32d811b71462f0db82098c0f0aa569
z4d11429c2763b8468ee39a09f4faeefcfc51b7978bc6128dfa5465df3acac0a9d6f77fd4675c15
z7075beb25393911a0d11aeb31cbf46b39feec94021bf6264c4658d6372ded201a53dbf8c1d64c5
ze13c54fea8ce9e53fd5bbb26881ea02437ab882550f77c0db4f306060f428dd3dd9573ed61719a
z904ed986d5d42a7857f69f119bcf79156d08184ca31162ec86dcf9cf0b4a746b18e8e95ed90835
zdb6bd655e7ce004e0e81f309edbc78dd77869985cea724f92566ba26f93d4054c2a8704ebac888
z61f6238370911e829ff8160d95898da3de9ad3861222fe8ade93cc7c4d2f79e5e330afe56777ba
z9ef2e13166ed0ec6b185f4dab513df703a15047221ecad3105f602c1fb00e0bfd2f6bebc48f891
z95221851f9bf8cda0c0757b3db518a9efbbd810f99d0137a471cf5f9b62881efd882fe2a812de3
z617015aba36ae1b645e45a5b776321921038e19f65c885e039fce20725dd2f5d9a79a05659105c
z2ec26744d03c2385fcb312bb57c0f8255b4011814c71623369fb9b2bb3f7513418ff4729ed4943
z654b37a3428b1f08d4fd7b2a0cc35a4a283c9274f7043b695fcec0d78d3c39967daf1ff7bce6cd
za0f6b19e0c8245af22e1e95761dc14848196faea2aade8950fba904497527074f03d5c956ce435
z5d7abacc828e55ab34343294efcf8da8f0218af4b325ac10c27f820439d10658d28606556ac8d1
z2baee6d57c4f7a321efe543d51110167f1a079c2c7b264e78b426851b57a776f2f5759242cd7df
z9bb6311125cb082ae06068665b3e4f8f823f89288e0b259e16ff73ceeb692f0aec2e7be5a6670d
zdab9d11f6ecde5effc9f7c4bd4af7de55f8c59953b7354c6775d7625ae044bd9e427c45059b679
z07424d6700d533a0e6a24c85331137108d7adba3d1a92235014a329ac926afd782e1314eda7a1d
z1372197262fcdd575c2bfcd2e8c2c5b132b772155387a2cd323a43eaea67d00196316305f1a590
zf06f65fc20406b72a7eac2ef2d6569b4014744579222195cc95c9287d4ed5ec93d8265c8420c83
z9b5c90c13e311a73619898bc36451bd77b937ad8e9e611c45cf11b6fab6f3d570a279f112e9ca5
zdbcc442490f27c9d1810ec821d13342b3259a8aa944905e2b9cef1bba16a348d02e46057c41251
ze12878af1c1924d9d86cc660675ea753dc7df41771f19820e01095ab000babd05f5fe648adade5
zfb78de2ebc0a9d0ee9657fdd2f3b998376618c18ee1fbddbefa94234b643f7c09e606569edd5e3
z3551d2dafe4da5a80ee6bb180b7b1a4d2e0c107b3887e12ed8ed644b051815ffed03cf29137524
z55e2a0fdc528c2683b14907a344e822801b4c8009e52d940161353e0a49c61a50c69630ef03093
z72a1b93f4db75dd3f3b02d03eeb63f81bbc5ebcccf0084cf66ea4fdf0460bc208dcb8dd0bd8028
z390a5d0c1e437f9a063e4305db629202cbfda1f16539b6b374eb2b578efe4d6581c7ffe489254d
z2493a0f9d9f70c7a6ad4b38f95a19c3b7823fc8af40acf1701e3c364eea03a5ccc5382c9d7eaeb
z278f36b0cca5e0f2077d2f867bdad4fb921218e6f5fb443d8633c9c23911d9a95cf29320c20ba6
z22435463bbc10183f8a6dd1aad3f6a3f860e2fb48696344979dc275b7e9893220dba209e318662
zcda637b0d5f87490a0284ff4dc65ada09979ca5166dcddcff8477d9d886d5499f3d6be6e445425
ze10b6eea32c22e2b9bcfedefaadc5bf7df49e4ace6d717e34f5e92f995b6ad5a34ab882e846a70
zc2524713663e0da36e3b20f3aabe58049f20e4ec28d7e9395913ce4cf73847ccd84d046128316f
z3fe65f32ac54205d6b03cd7ec809d8c7e15afd5d7916af1a8e4078a2cf891b1b7f375c98424ae1
zae065f6ae55c806ae30b33493ed6eefc9122928265a7e85297f942b4e401a7753ab83968a7d64a
z2aec5fc56b8dcb914a1ffd1bebb3df5f0c377bd7683434cf5bb108519fcc6ce3deff7d706929dc
z82d9025174ce764b48ac0376c03fa5ff43f1aaf0b5280df2598d50bfbbd24e69b50155df915b8c
z7cba28a250b0e851dba1e5ef47af13fa8e02c98737047b0a2efd981063594f496f8fcd4a5ba62a
z4307f7fff84b9a4f6f6596f28ed2880248f9ba224400ec1083b49f539972723aadfd57c8203e46
z13bb2a3294428d4d56affbae4237c1b39c3cf85fae9326af457879bc523ba82116da10135ce82d
z997dbeb4a7108417fd39aa35e5a9540eab7d72f139420d687057f8efb86a5c1a3a71a7c3ebe97d
z3e08ed34c5933c4f769e8a0e89f5b2ae8ae5fb80b0e091102d76b67d00035b239ea6f4c95dfa12
z7f1d279e45650312e928a7ac0ceae828c2cc7b359c8af02eb8752f3280f999066504c275f21ea1
zc3e5fcd6e7caad01f5c490bcf2721bf44ff03312322c23b0659b4f4bd79fe60c589ad832f6d218
zec9edae14bb4d0643bb323a8c4a36e99ae8a3187717f4a39d5007a0fe4d9a2c26a920f37378520
z957e996f11f58639bbe3f811c6588659e0f19fcb0e833f4641aa6f4d06f7f8197b6254bfbbf173
z631d232e32c452fa6522391b8c775d0ffd339721ea0da97426cd22004a12900eeb45e0c1ceee9b
z95d11ad5e5bf2988c331240cc1dc51bd8932f028f973df24f146e2cb39c5f3f7a1ce8b20b5aed6
zef5f33aeeb8e36ba43db66f80b6810977b8631652eac1d72f15a450eb31d2175522e48e5b310f3
zd77bbb626d852f1eb3a132f2046cc486433653c35886d0f4223f36ebba84878c9062d6af3a6487
z8bc6cee264337bd1d8a84c2d12e112bea502dee75c7c903e744dcf817a440beff360f3cabdd1b8
z3da529b070e4b16b85ae918047393e1b98f18f15a69ccf4cdce0128f3b584f7eebcddd12ad48d1
z1c65b8bb14141d419e365fb3113001ed8e2c89dd1ec83a79877e4e50cd60bb27dfda5e0208bc1d
z42fde1b597e3fce3667b451d6bdda6761bc6423208f7d6b501218cb646151491926f6289457300
zc04fd82ae33a22ba6a5e0c992ef8c31b0455ce02ff2faaa884ef447c14ba85973cf8b6f095aba9
z53bb05f99dc3bfee81403a72ba6ec1346b1af5c6670551ff80585065cc5b804d11f2de5bc338f2
zdb53aa8d0b6607faa29fdfa5c7a3893de703969585bb0dcf140b2413a853051ad5b75a2a7a07b4
z6f83acfb6749d85b143d30066d4cb893cdf0a655dd498993c82127a8ce180ac4f2b9a635687b39
z20d9bb287eb55ab834779ca584022c95a8c23441a011171aa84f252c34a3780b6711ecad73a2d6
z93e08f60c5a4ef22d60430f010bb0424501190cfb669b55b12775570003de8be8c71bc9f1aec3a
zfdbc793fbc3ce2364ff9d2761fa87fe4337d113e1bb3fe4c65fe2ffc084d60ad256cd57a7b77a1
z16f25199a2c6b3a55c9f92c2ed1d2e9afde5a2499138e27d8b86c51b14ce2bc91d3a950c312ef8
z0c37beb5e8bfd2ef4672cc26383ff3c81f6172008d224aca929d39c8a2dc825d27cd07e4d7fbd3
zb49212ed42b87bef99c7a8828f1c471a077aa21f72185fddee78610acd80d5f2c89a97cc09461b
zbe98377af67407fb2bfc0c45ab674448f73e22d3749fc326c826f603519b46717e8013d5d718f4
z47542dea7d5628a704553a031d3e4fcf8dd9a97c97d4fb8775f53d56e89c4c826e3106d46a54d4
za0bf2cd7b1e768cbaf7b6a0119d2b9a7d8ee0e989d1c08199c9d71efb38cddbed00e5182d70590
z3caaeff01421570b3f5b8d6907c6e63e936953f86faae8e704209e61afe1bbe93a1e0253080caa
zf1c5d6bea85a560da823b74e416d8ccdcb4d35eaa3c3324aadb236026acd103bfa4d0d3f2b4631
z3ebc52d1c5171bbe3ada05eaa28d4f84a6cd6d5a34524e2e770dafc2f810730d3350e75ded2d0e
z40df4d4372ea72fbf3f16d6ae1aa8956b6dfcf7a0ef6ad9cd880b1dce68e83763b524502d300ef
z141d00ed4a5f482dafcaa5226c234c5de0164bf5e9c4d06dcdc970a202ae6c1ba84d96ad0917c7
z10481b1cc9f86e4bab03241645b5ddfe642a4a244796dc95e6e38a0806ab49c6f18be40fe79568
z4cf26229d94f333e0cbd97d62d82f87cdc02de167ad7dec66b40eec57b712f2415bc16130785aa
zc2f93c74da7ca430cce3c59b51ed88f3f068b9f58e1d3755afd50bffcca719eb86776cc6fcbd84
z77774510c410ad351c57101beed7c09412b43a80e2e73dea74cf741d3d3da54a34dc64ab6455e4
zd3be069c003d36a78d6712e0f4c9c1e267c5a40f06a916661af820c23503cc1210032300a2b20e
z48e161d764185922c84ef0a40856584d757bb33db40c23aa33ee4baee111ebbe0e7c3ceb0b29bc
zbadb9d2e4d3d707ed1f8813752ba209210473024dfe3cd30eab15daef0fb1b13b833eef0aad785
zdc3275faaa5f414c7186fff9608e1f7cc0897cec4cfa0fc47810d47a7c21c1769518d5fe25987b
z97b447100488ca1701c94f4e03e05af534fd8e1530da10b0d85c7a816ee7d33653cc41c2334cda
z824c9f9130b599df2bc5b9d2d13cee628afc0d1658da03a1ac58f35902cfebe0287ddbf0a016e0
zf2f1f8ccb4457a7899dc2221eb53d75186888030786b7c92bb48f4fe68b9d42ec29b7448e85fa8
z78a6ea940035c1102996b4121b324b8ab888cec07e2bfbd84429d28aa34dfa732b01736afa7088
z0bb53ae62714ab35c52c24814daa10652d10d9804358621ca264bdb0c7ee30b5695bb35838c627
z22a6094a27fb03bb9358978a5007b700a3697553d53d2637264f476201c67bc01b4c3bdcddc66c
zc14ed7688593ddf778d5a6d3f92044f2239f719199a4989ca97f1b859be6d7ccb5dc7922e098bb
zdb881c8fdbf08e27a36bf9bc7fccef2d5358b6461227f2387f6b428d164be6baea5c61bccdeb56
z29ebcc629718c075b6518d055394ada341760394ca1d3b632d3bf0cb66a74d903fcc089782770b
ze40c6857cc79faa3a4d87ab51fe6aaa1548e023750538b14e0d7d6757e1dfd3a375694bb03c5a1
z2b6eb806de85ce6567a907b9a85b62e534aebe49021609b7ce7a80670d1b072bfaa0c4dff2c5ed
zb1246fe26907332aaa824cdbdf8bb4933b983f0cc69c58e653acf2b06617002f99e15e179d3b68
z621597fc4bc063d7eea4e331f464d1357635fb0e7de4942baafd63f31908536c8205dfc704c07d
z747011ae3dc65e36f99017bacb18875abdc860181e4e203a1eb28fabb479218e144cd9faf933d4
zb9dd4caef51c7203fc98240af11830c08ca15e2c49bbe83626f6fe0d790249c8612e9ec4003adf
z86ca843304c9875897255ba61ca061cd0b91e02aeaafa6c322ec80312d95eef93c56f5bcbe3a11
za353dbab14fb87b34b60f3ae0e78766a4cfe60a3f10e8a137b7dd0f79fdd23c27c2ee5eeb92894
zf19bb3ac54f89c103d3d9f9d9c67b3320248514105980522ef58921619621f0a3d5ba6474e0207
zc8f7d4d5da6ed9d0d549be48798aa1c53ea37d9783c70622d0fd8e2b02b9a9b4ff4868b2c07e01
zcce9cdd0f04041f97423085f366b6a64980623d30e08a6c32f213a4dd4ed01cb3d7d16dfa74df5
z966448ceaddc66b4135a9162c01dd23f4e47f8db4384fa08165e610b94a2d661b748944bbce092
z2e5a77a10bbf3133ad122a2d424d1cc5bb43742df80fdb02a6d1e767f5741386e5bce76ede09e3
zb1be80391d5ff24935fb240a5c23f61b3c1b1798aa51ff1b3373b0863d488078520f3875486687
zafc3eec3a16023e066ddc873fc3144334a86003d51384796c55064867339e63a3fe61e413f3129
zaf1d1024a9768e4d292388cd69fc3ff74870cf674f32c368af75156964293ce83a8b5c76b553ea
z22cb5d949b365e58046967be548b9d42d899a33e454a81e6d315932421426f1e077d3ad794d5bb
z88e33e0a90eb43e07ea24e9b924ce97e9c11c4bb40219b833779f6faaa78735d556e31118f37ed
zf0fdada16a0e01a8e006f78865f4b0e6e79730b9b8aa6c54c315de3908580ef120689c20a0bb38
z85b4806de21feb3e0c71d90ab8ee483ee006ba565f55addfbda0c3d61d2d05127069cb050be7a3
zca7771ef59a6301d1e40c14e701c001d51ddd0b521dd446211eb38df6890b598d1f64f87ce813f
z068c37696697bb70fd12f9d41e675ec0b5269c6bec5afaddbe014f5fd636f582648388b0502edd
zaacd24e11abc53e274f03fbffd8efe4d8c7e1515fee6b4bea5b422bfbd10b3440672e6d0e4b58c
zab58df6b255206edde160169af063ead8600c691e9549c8641815ae087c93dc3b6195c6cae93c9
z1226183fab2fcb5fd4c76a40e6d2c4a7993651d60ec4e2424af697d2724f1bb4096900a9cf2eb4
z331902ddbbe1d8d066f6f67d14a679c5ffb437d6c3660f7c7b2fd318f56d8661f74e54b48f4624
z94d4bf965b8c1270596af4635c7ce32c3f1158f0dc7471f959d1f0d79ffb3610d45d7d9cfc0a39
zfa21575eb92993663956cf40777578414c3cf7aa40fd5ba3df5b7931c6dd7667e5e1bc6719cf5c
z935947dd22029c745765db1f25a6422226d35001e8dd933550e7a240b3f4aa78b77f64042b5eb4
zd55102ce00b879e8bf3f34546e113c4b0a9734597722f6ed879aeeabb25c0b5c0968f56da76323
z7cc7f4b522a22724264e59c86923640fc738fc4a55934f85a54f54d6fb22efaa9c0eb2908ca1a9
zce1b6226a8318420b8da42b4034f1fa3468013955ab1047f88e9cfad3ed9d823a1d0716edbfb45
z654bffedd4b2d7d2157ce5bb1065760094fe540e493ae96031d5a743c61dbd6abe00c46138277a
zb105da9b2be657e8d523276247300aca87fa243cb13b53785339245ab10a8904d453ecfcfb646a
z054a1468868be5c46be3ccffde1049850cc05a3fcdaade163007da8d85557debbfc281e08f1fdd
z3924095db612e512d559c29ff0b0c84692ba86c6c8c8dbddb006bf3eba5b9e89cd87ea5dd1eaaa
z8bf3f05b0c5b1fc0de26655d319f1f5f0ade408222dc7f8ffd6ab67d5d61fc1ca28d3a26ba8770
zb37fa42be41b718f33fb81e626d0657fe51442c14f06ba3415c4b330dd109c8887007f9953fa1a
z6a9ed6bf11e827ccdf59d629787703bb779ea8282061fa3a039c8cf00dd3bcee1a7a25849cbc1f
ze34931a7853408992569d6ab82ac0b8895618d45a5e63c0360568a9198f67bb718173c5c9e9fdb
z80feea59594891afe4fc9eb997cf77213e9eb2b8694d782e0e16e0c717493c30b687be3fe09a5d
z028a142086801fecc79890f418c389ae86295433b38a0dcca30464a0d3c2a4e793c6a63fdb7ae5
z9e4ec0ddcbe109249834eeed2642715b47c986ff7aaa6991b5dfb31870f9e4e6769e076a4514b6
ze26ac154ca5c59f933bf7d6bd128521e8bccbc76a612ba04bd167a67be2e1f51a7a0df0e699c0e
z3387220d2efa0c5b33a250f35120f963f2d9099d589dc8d32dca345bcfaf753bd2dc98ec68999d
z40979616e26b8e09d667923f2941e5670b864a66ccf8a32bf09ba5eb4a8d47ce3023a765478629
za4774b0c4de7d1fbcf6dd2d825a3d38f1f2e824353db45bd4d2c5e43134a2917ab21f4fa56149f
z728813ab7a9b2bfe18d9f5854e20a6640082ae2e0c846c0941a4adc2212ff1e221a57db3d23616
z1178e7b5dc1efba2ce18418e6ef1df1c9221b30015044930c182fd95d5008492206d59d30b03fe
zd303f3d063924c7bab4d8daa6636864d3190678a335c87cbb95e641fbb3d16bd513e3663b8222c
zded9e7d9d1e3ee73d73478891cfb9b762ac858004dad9aee65f787fc3d990782321b99c56881d1
z5bf162290e4f76dec805af2ca07b1d300ea300f453de7e8ea6b3ba7561a469a3fee311c5814182
z68da8f2c615b8225513f4c00f50494b8c63bfe0ae2354d0c64eb4f7035b28a288e105563923371
z304d52121f42024fc1fec21d511f575bd0c9199402d1b863dc8f4d63342b4ab86a4f7a14903882
zddeb1a7b90dee7f5c6e833cc8ebb0678e57f65b5b5052fc961204652de9aa8772852c4af7a79f3
z60dece6532f31951cc2dc1664f23a3e34832e7da005a0144f487274d2087a5bbe2e02833619c6d
z5e1e17d1c696e67f4081048fd2625478f5ef03697a13988b6a94444aab821f4c99ac9c886848c5
zab1372984f5906db95bb3c9be1159963421d150346aa241b9123502cc4637a238c7049a236fcf0
z92ab6a21728886b59df6af7b0550d4515e01ee60594477e867dce695d57a6ab1f14010eb0bae6e
z4602a37fc6d22d001e355e443759d051e9b8e779881e0e6ed49cd0fff0d45dbb15cf797921530c
z0f8e7891658b4814334d9d7c0405028146a00ac0daa24392320b42d92d5f7cb3b75f7ff08d3a47
zc4abd9ad38561647ddb760bacc4cadb74ffa7a9a25a3edaebe1a7b1fd405833e87311a00f92c14
z8d4f774ecfcb22a618386999563996f4bdcee352578f80b41c4e53456c8126d1f29865127e214c
zd94182e65533fe3e5997b77dfb995b2f6c478ec6811b9b70864e2e614a8ea3beecd26863ffdc38
z0fdba674107444ae6bb082d433965256c4bd14419b72859034a173f0799d86cb872ec861c05f85
z87155ce9b4b0b109c318b7ee5801da8e7ff4fdfd07b3117a23a7047b41bdb109677932106818a4
zc902ad53d3024029a8f0c9be80af202c7ded6b4d8566ac2ded23ed37678fe23a77639a3b51dbcd
ze57f66f1f99bb37b58493f0349fbf898186ee9a23f7959cbfbea63ef2615d62eb0989d38df1467
z8fa3216b0ab6bff6e925aa9627c8743ae73488f157184761a79e028ccb4177892a272d1b1c3936
z61048c67f0067618176826585a3258951710d9d0bf47fe2cf7c212692f81793efe7dc08b7cfd47
ze33cb84125933661c64a2312735ba3b2f544c1d6f43f8f81487f0cc2e0ea3c4c9c735e04db5bb3
z6eb1b4ab8f2bcba51d284e9c1974f6c172f98bac928f9b867e73891145b4cff8847f6b22b3628b
z646af02c945912ebc163d440b39833ca031459b055dd061acbd6cee80de9b1533ce341839ddfb8
z0410b2288e57e2fcb114cc7848f0097413d09c1459222d9d241f6d03e7b8f1257f6dd552124c26
z7d7e3491b69ce65bf23e84cba3d2d8dc26bdbf75a38ea7976fa64cdeb34cad6209f8a6d145b483
z238f48a845fedffe5c72d7b5aed0762843aa7e37c0ce4dfd91120c95e4727c672948f3110019bd
zf45b98cc2e19012078ee17b0d820c8387fd17dfba324bf296dcc7c8b4b6d411078eaf908dae45e
z9589d93f75e568c564f59ab433d22e740084ac06e926df20f7b07fa55c9d060d5c75f80ff3a435
z250478a7802ab2e88e7c1d2f59f96aa6d9fa07edad41fc5af77f363befaae849322dbb28c97d8c
z3af56b7e396d86360a389f2544326a64e7ac1453f31d160dde4ef8eda097896e64ab8192bdaf46
z71407533535b96a8ca34fe6855f74b780881a405cf9192e746cb3aaa08466da8b5d4a8df02a644
zbe0e9625007f47997950e9b1ffb253c1363a2d590168e918fa12c08ce73acff1c36b1ab97ebcb0
zd77f95c53df9700787a4672e65fb45fe4a1464035afa2ed0a50a9dbfd0c6ba92c3d41777c89527
zea8e7a6e3bea6eefce5318d3676b3a3a9c1450baca32d86b43fabb6c90bc74d47f9a46cc6bd910
z33e343c1f5eb3e22823b6d4ed4558ccaee654040fabecbdcddafa78f73f836c0feb613f6cd1d35
z9c37d03219f538ce6a0c7d583622a35a7f0dd933cac7489c3b178ecf558bf831f1ab461d880abb
zf66c4f5ff2b5e30f76072c215f259e6e2037aa06ad2eb6d6ceb8c69a9d4288887b527e0ddf9c9d
zbd7655929ef8889c993b09280db86c927a5ca6214608ae8f789b67008840a97e31b2f680223c04
zf13515bf4adbbdfb78beab9b19eb0a4d1186c7e7b1fa3c3fbf369975166b97adbfbc9f6f1689cf
z86708568ff2e135fb3125aa8230bb57e3d5c8b45aa0b6b216ac9a8789a2458fe146b19c162f207
zff0771a8e61f795091a41c0ffbc1b1c536f60fe319ff46e38e92d1fded28eb7a9b50915c208659
zb06cb0f5e6b44e0b766c03484516c07041d4a75fc022944e37ace993da84017d9ff8dc56a6318d
zec0c71415ef2f2f43e44d9ae16fbab61897fd72c13ba89d3d168bda4d5b5aa53f3e70b0655050b
z7b626389ff70826a20a13d93329295a92d0377e1243e9421126edad01aec5c63ee2b70baf61fd5
z40d590ea2dc52f6f61a3c7e593234db315f6afcf6c3ffd47fddb946a24143a7fd846dc75db7398
zb9d4b245df4a56dc8294005f4e77b25faf962da464c7c9bb87828de731fe29662013cd2a6f22ad
z61f3612c853f92e0ab333b79e2be5cb03873f1db197f1bcde28eff9912f6dc58eec8cc6478ebde
z663ea2069519611db5e70a80dd9b099b004e665c6e83d8c58adfd8cc8d67f85919b2fc907551f4
z1f7f0d41bafbcab61bf8659e5639efe849fca6eff4b3d79119de4cd9691c22d3561c1d161cb4e6
z50fb2b419d4defea2d5dc50661ffb0c465b1d095c89324658c97960a838cfd4cb4e5311d71c22b
zccc2224bcb37251b49dae02ac5138b3eceff3bb3a7b1d735cf5333453f52acdf113bec3b2400a5
z8d25b01fa3ecf0b8964ec0e9626dc855375552f0c12b7079577e30d103503be96154cc4c236d67
z2293a6b2a114f1621034e0117d74b7d7cdbd9a15fd585caff717a5fed78cef7311236df641e9fd
z4398de20bde104702cca31a58237811901803c6ae21692935f96a378dd698ae88840f5e19c6c2d
zf92a61c025bc7060a8079e3f05a2f860a04dbbfd124ec99a6299de5101473fa65bdaaec9424abb
z2a81132d3d2546b7a24f0e0c65b8821e083e174bbcc2185148f9f1c01db5f76049869e6f12f7e8
z267642c4721d33b4826781ce798c1d1eb973c39e3eb361a30c84a62eb3612ea68dd64eb5402cbc
zf9cb3a60a76c9971b3618859f661710f3c3de46be4a8c4eb5533038ab8047d2bda36665f2779dc
za9d1f29ad4c64daaa5d007ab670b9ed40d30c860bd7a2cb06faeace7efde2085e12e6771b30cc9
z2621c6813932fd64851e0a5ecfb7653fbe203669fb99081d73c885f0ada4c7cc71317e32d7df94
z57bce267fcc8894242b765f515b123efb05590e1543ef3c38c571fc7ffefa8ff3f4bce37487ba0
z8aa790af4589444e956f2485c4ab89dafa5fec59305efda2788dc694988cbeaa7490a6af1eb163
zaf3593cc9291e2044b93e788b59fb2b3da855dc2591a32d448f9d0c37160fdea23f41e0c84adaa
z346e8c619a79f6a41b051c680746b53f3a6caa4f7a6d3cd05cb67eaf72f2fc21acc9a0391519bc
zc8b668c068e43fa3c0f961fcba70b4f9f4b72ee28e76d16fb9e30312c95d0f9d432fd9d6e48198
z0811c88ddbf500fae9d5cdb2cb01a59ff09d79e907fa2065e8448c287ae0bbc78d8723396b737a
z67a1ed5871c0e82ccd4058022811ad9577185dec98db0f55393c88ee97e9359ac6f0252cc59251
zc785d321cb1f503bcdde55a81c522b0a4025d120534b529639795c84a5f582a5d36c96c0b89d7c
z2739a0d18de1098dc3429d8f32539ed0f6c481a0c2a73ec6bd78e0a1eb2b42f2ee7b50d125e564
zd04f9fcf1cf6f3f0a205c17da9395a7244b48af236a01ec37df7337f66eaf48aeed5c13d5fad2b
z723864bad4ce55fb8ceb641087bac97f23285f50a8420199e4b4a973ae25a84d150784797ab5f1
z451ea43e9f8f3fc223b11c31766d0ea354fbfd1c8dd01e45f6d6fb7c8d7535d57438db7f19d71d
z15ba79df67b0938afff821adcba7cfb6528053f803f27654b5be256acfe3ff234f7af32b13159e
z96341d88455c629cbe4f0f5d37922b0a410e7276a66d0097701ede403c4d21218c9019b144d289
z6237cfb0e4f27a7658258c71de9c7632c663dd410d3398ee6b38f0209efbe657663db05b8af462
z668f0632f21b4718097e30dfd2fa91cd0feff0ad8fbc5b677899974e7df2ca3ec3d075ae108e75
z77982cb3fc3a6441aaa7be26c7b957e46cfe0c6e6f4617528ba406e4b630fc7a6aabb14ec6cbbd
z5c3532902277709a7c5793a809718ad5f91214ab4da7518cd9ff7fa3d9db61956e02375eff8fd3
z7aef0c9c1a8571539c3af765b02c4c13a81de823e8b50c990758f0203e60a8c82a17718da15cf8
z590c4e6e6a330fa7c5ee2bc0525bb8921fe45733f7d2733fdd884d1247353bf5800488b8b76594
z3c555b01684cdc7af16b1a456413afd6704723dfe6049c23b26595164396c408e3e9caa9d60e21
z09f8b259918269a51a0c603bc94c5eeba12a1f274323ced6a040c2f8e3e09f604da1cd591f3bbf
z00f890a734618e01e0f06a2728a2a62e192af3e2a7ab2d054f7436426e7f2e46ccd328e999156c
z25aff59f66931dff3d4d371dea07de0724e90684930d1697e96ea44d0f1b337b79863b32bfe076
z7370beb73d7870e56c94da9a45ed432b94b6c253be8ad0c23a97b6cf65bf07dd48860d37198bc0
zbbdbf0ab904b533709d965cbb70e1ae70db8e55b71206bb8928284a9f340600bd0e430bbe10560
z3016365980d04ce318a7abda04ae5f8c9c42c911d7e4c30c6fe2b4ead320845a91410fbcb1225c
zb98045140a95632c99f8bc8784989b217e95cea196138c600601100f64860f74b3741cb8245914
z274f2ca7ea34098772955d8f46a9e141559a5c5c455f0d9cb39590ba61d8047f52e294cab4d2c1
z50fe674d4e9758bd7159e7563779afd2fa7f243d791f07982f5b039236178c743d8e6b8bc42db8
zb34ce49ea8c6d05374f53f5cebd89d455095646d082b722ace2a8702618cfd22eba5b983ffa203
zd7a9da879b48cb263fb7751e5f7c07b0c941d761436ca886f0d52ccbdea6043181848ab4838239
z2645e18b39c260f3c193c34ba2911f6bad3a3c8acece0fc13aeb1d76fe6cef1ed4f8c08aba3d98
zfc7508647afeaf30f2229756ac0828284a2b91493cc4e30f4f98451ddb2925055cfec8a02c2932
zdbffd3bcc560c919ae520a9765133078585b9b2c7cbeb34a233de5e76544fae3a9ce4d4cd1421d
z5c7db20e09950f7f0f5f9c189d65046972a9122ae2803c2658c559d486fd7a405d03f4bf9f96bf
z2691cf5de3d92498ef08539c24496cc4f81fb44f5995214993588647327a6130ec97510bf9d7f2
zc3117045968a77c0b243a64dd338e23fed8e4e08d3435ffef402e23c5bd3e03cff0100108f0bfd
z129f7401286cd15f65bed4115c7e652638f04907b0a8e9cb1a675376d597a3905fe9cee137e312
z6e3eee114e29d2915b8903b6b8e6c0e590690febff295726e5df09d0c7925bf208f86a02f16edc
z6f9d6eab563f246103cb43194a9add60510a771da6ff1259a8703c103980171355363fa3515de9
ze044a0dd34bd5c2dfda27995bad5de0b55d90d46ddbe0b6a0c55ef82ac4a6173f5f17657e06c2d
z09f6a387b2f7adf2eb27e50bdec660a639664e486ac26fdd2bedd67ce9e003a346efb6f3ce95f5
zc058119263a7024b04f9b48e210c217f1da76f25045ff65e77942410945e745e7a7056230b02f1
zdef2a71fd3b2e8e006182dcc82f5f55bedffd42a36e11ad926289c954b63b35a7e5cb1b8a0c46d
z39a6e2ad83f531bc81409beef0e0564a1ec4cdcf72769fb60acf2a4a0a0785ab5d7ebeb85a98ce
z00d1435c2794a6e9cef3819e60982190de324ba83f7a21259776561c481acb863f36f7d4e3a2a1
z600be61b15e3e90fc091efa6097e1ee3dc4e236f2cee12d64a1ce9015fc6103ce8e8a67b721a48
z26c74c48ce5f51a19f2ab88f43da2ffa4d7ca98fa03df0d82420b4fb84e7ea141bed3338559d47
z9adaddad8f44e1687e150605b845b711b3dad359da87f100a40bb47b12d0e6f48b2bbd95332c6b
z0b8ee7540c6c78b89ad55a0eccb9bbfa45ea5c352e63b7704087f12b11d433f9aa8f996d8d187f
z89722572d50395e84b01a51d3f90ffea0b15f5fdf39f16f2ca705a88d891b319cc16a99b5e43cf
z9b8b5b7488db7e6631141250a5098d7b6478f88c71c4cf3d2979f1452a1904ca6915d9aed060e2
z15422e55be1f0ae8bc7e4fe9e65ce1d0876b7517fd99576e2fd30b574782cc8aaae4af15d142ab
zfa97ebe51014325fdd552a80fe5d2ec0d97bfa5355dda142dd8a972d6d6d86168a2e208bb3905c
z7ee51848d4974a34bb4a6c682f0e19d3512f037a7a8c7dcf7024dade42e41b7d72b5fd28e9d270
zbc1f96f9fd7ee5ec7a1fa4b4d83499e357bc5642b4fef3988903e033482d1835efb6dc0a813309
zb582af536efd0885741989e8d2469912d6d9e8d246d575ffd3d65116850ab5519c5b2c43eac4ae
z2516f65db44bd71a65e1831affb80a0a37a74340c899411feaf11713932134f98442baee18a466
z78698e0159a5029eff9847556dafd0e4c10fca1a666c99447cf12b43d25109dd69c5e061c9085d
z023f42afc54227b3dada0c564fb196f35f1d2ec7076ac9500a44e597de7d7b0635920a385ab55a
zc596c8034d17fb1617348e05ac69c5262ead91ac14ee989eb2379abd38eb88cc4403a4d4b9d4ba
z0981d1e85e484d6a544ea68062988c7845fcc872867f936b218be516ba49754941c883d484e1e9
zf06ab17a940564a56a66bec7c77a22287650f675575d67811b5088afa160875ec50e83f84a7b63
z3dff2e6314c7c4541c0cf526ddb5f60ec503bc53393233311a6d8cb6d62dd8daadef5403b92f65
z4dbc4fc25b7496a0f70b86fe268a055506dc50ae9c351d80c955811b5fb464dfd9a3c69da226c3
z70954b027156c0062b78dcbe56eb12cc6e5b896af56f8ac45d00abbbf9df66a6c4f545655310c9
z123f0a6604c4e51a3a3c84a7e6f757d986b8cc333ac7bf6307d8895e2b27016f69599957a07777
zaa916859a3221abacc2e9529d43b65c68a747566f5fafe3c13e49c320f4081a3185bd6fe1daa14
z72d57baf274bd30756313400c9409506d4f0ab112a0b764db1c1ce64db4ff7c6ab5ee0719109cd
z0185e6be38a71dab12cf996375857f54caf0fef16edea5bf66458b02fecd8f719eeba26e918750
za96ffc9b675f3f3107a32663ee97bc4501af03bddecf27a2c7b84d3857f36f1febea09f7088fd0
z71c4765688978fccd8f1bbb801f3ca4d630ae152715bbc8314d86e6a3e39139aee6c295aa42891
z5a1b5b86b27e85e63917cf86b92094bf15f7567532286872dac254d6a59692c75b8838b609f993
z51cebf4efa9fd5ae279a8856df139c7664230a6c36414cb707200ed9829690fdf6db80c1a25dc4
z76e6f4c539a03a6a02565db8d63478a2804a7cfd2ca802602fe290dfed577248b1eba9fe83d48c
zf6f5988445cb431ecab079ecf8751affd15a91eebfdd97ce856cac3bfb71ffb083b4c790c6fa33
zdeb2cc387c42854a5a6d27cdd871bce90bac93f281bfb7fd9512be233404a7bc0a5fc479984c86
z2fe7c89233a867f2945cc2b116fddf6117e32001c380ef64afb7e3194dd7eb317c0fbfe622aa27
zbaf29bf6db29e99268f97655bcde8f86253ddaf00fa472f0a547d041dae11e5ed8792ef9741d5a
z397aeba3cc9ba09bdd1ef66c99a0295cc5b17b342e3e960c6dd0dc46a1eef1d7dfbd2193fe2f9a
z4046b6c1783933f2a318deadbefe935016470ef64daf543a40b9af97e5c770e0888300412be0e4
z81de567462b1b4ad2f0bd8e92ba72b7a57a6b4d5773cd9c83aa1a3cfa06a1708d7b5b6efab7667
z2d5a696b5e2444d3f35505be8e6317081b9c04603bc76e30cd8075b5b2300f7087e2a04e04356f
z507125b51120c057cfe1294f40b604d08f21de77e1f81213780022e7c922a8d6e5420aef0ab731
z85b80e3ff4071a15fd0009e690c2878855f9df2cc85c511e67bc3181b8406be674faa6782841f9
z19dc0a5c6ee69dda8065d78e4c88f2d0b8a58abc22957e82d34686ea076a7e6a31fa9b1a49674b
z2d0ff573e565fd7e0c25c2a50c794ac04b9d1eb786aae25e8ee1fb7ef6e56d4f0ed01c5bdcbf90
z83916edca1936022dcc170717b0374fd9be2d47784ff4329eeda2dd1e85bd6249bbc1043c9d97b
zdcab26aa20427f7f94262326317045dd1362e39aacaeab6c2dd608e136157e3d01301780a2f709
zedfec2781e3be6cc8646e4a5cc603844fb51adc87465a77231d31755b11d457271453c966dadc4
zf602c094cef225ba655f85c9caf639f76a97902f75ad9567cdb72b1bf90f888c621adcfaa8b095
ze4412da01f68233e1a0458bf289bd89f9c9f844eef73f47bea3ea9df22573345b40a6f497376b5
zc5809c51aa99ecfe5926dbc04ad20014d9696a49131d568594552037936cdcb7343c634437fcf6
z864835f0a17e7565433458202477b0c5c1ad14f1537865083f97c6ad5bb7e84e2197c1a99ed071
z369b703964eb7d0f5e3f674abec2e52c91451eafc0223f4d1f289f4d06d437af49688bfbcb4ba9
zbe9e79f119c815092965c3ec7b1ad47b0989acda71e171c6b60b20a7e90c55161cf6c760cce345
z41b97ca712e5d5eff493eb223c47d0c4f71d300e216c37aab73318b116a637556d6463ff7ae58f
z2af04df3514c97e1d6094dfff09963e255d222df22d5e4ed96137d79bb81e42f5f9b476e6690c6
zeb5973eea03a3c43e254d21784f4ff12296a86d9ac75ed7d2f2dca0d02321f3742acf24e01588b
z37890be8d55478c09f67b40a40e3e019b6f3b43566c62ef4ee3cccedea0a5aa4a58a9e68305944
zbf23ffce6611309da309092941f204b009923cfd0aca9e1f9ce98914862f7198369493bd95ddb5
zd60c893214538d34e616fb0e182cba25eac8bbf4e448e1b5d7c35b5688336ecfef8092089ca353
z1a1ed3d15e554fb5a27f7844919f71e308c7abafab2431258816056d04bacdb86ff13198b99cb8
zce7ac443d8abcadbc39172f370a15f3620205104355bbbd0412bf0df162109d366347cd3d69443
zff81e380587b4f4a0ffeebced21f04be8b1fd9160278db862c0427cf7dddc6403dac1abc308010
z2baa735e8477e2c241a994115b2198ec1deb840b82cd6193965e13f1798dd02b1e90fe6715dc8f
za192402af66552b9287a8c18f13953f211e36141f05b189f225c3579ff719b814969878ed0becd
z74e81a3de4aa1e548bcf2691d54eda4b1b4a568642f61c5cb11ce3626d3b230c3b05f1ff57ed8c
z100aa1482944aa55ae525957a560e3100780d4bd920b8cbf3df64aa680379a1eca64326266d3ba
z90e4c3fc86f6a36d2bcd98ba52e3a69b454e15deb6441a7603530bb9a7f4bf876a9440c4c3cdd2
z65ee83f6e4b9c4d5cc753142d0de9fdb3eadab11d9e43daf5120f1f56ba51f49ece49d06c41152
z3bbb01c6492f531a390d2c012f1bd108c975e9991194e16b570241294fcb68edabe565e393d3b6
zf8bf36f7f9bdbaae969d47f271796ae6d87ce525e9d6a0d8416355ad155f1379aa7aa24286087c
zee13d01eb07715a575f9ff2a302d0994dd069fc62d13319f8651dec13dee932311d35edc84784f
z19283827d58799c45e1a56387d4e1cb5808d46719ce33f6f352c61df6978742619c918ca7ce26b
za91b206c0499154dec2af08a5b442313b05e4fb66b541f9697f0aff55bb764c657e6d2a8c27917
zf3212d6ff3364f617e9aa64015b4bbd36dc85263661b8ac8ed71ac31cd294938a27cbeaeb4d867
zf694cd94cca3a0178edee8bc9164bb84bc3e482b5f7ff4e65f724b7ef29e44092c003e46a5c0d2
z892b967a0681c04cbdb562ec2cdd9e00b2ba98c21a50cecd988b2dcfacd08bb74912057433b0a1
z9710d538339bda85a227b4ae63d1b79a7309f65754e8923907f275960fdba69bb24eb582ba20c1
zf2f5d353fd4c862a51afdf474000fc3eecac03cdfeab435d0ed05c08fe04fc5315ef70a85b1eae
z9e4a8d1c3b5265f4491df977bea6d389530a6d834f86a7154f2757912363e00d463aaa745cb7fb
z62c705d2fdb03f2e86aa624edc9c3be745bc6044b3ed0126c781f0d6fc2518b1221a29fcfc1f3c
z820ee2682857668ccf672e34801e72382604418e615684d48a770676360a43424076078d160a77
z5c8a843888e0f348f90cf9ce0c0e9e6244bfc0ea802d30c830577d4f98abf74c53141d121ef170
z12aedc3533ede8734a70eb7ec62f4873dd01e52977a55a16c1d10f504eea504fa6eaadc5bb5ac9
z2ca5272b268b35dda5f65305aa813f58f568731a51550b0aee596613e00d95f5fd3717cf51d892
zfde5ae1e4c292e76f551bce62e5342d48f046f553195ff697e79365bd7412ebb7ca41aa71e32cc
z0abb02ec016d59fa72ef6f2c90ca580ca338828b447c2e92bdd055939783d87e684418b6afe319
zec33bea650c4f3239cf81c06fafde89b7303750caf4ede193075d6b9aad4e71c630211224fcc00
z07317fcef48c595532925f3d160cb1f776e1eb4e3c42128f6efe2702392267201ddf5b455de470
z524ac9a61e06036717e72e913f48f4d9d4af1be2ddbffc023739258134e872de0dbc5c2ffea85a
ze94f4a3541920546b14a941097d877755f9c414172ed1c956b5ce943a368329d871b3e0081b09b
z658ea71b99cd6aea5ab38142f70e48cc0fd1b4685ee81ffa4fa5e6aa648cee67ccfb88b95ab6a7
z37574cec139b1cb45ac5b4fb5b5dfc2775bedcf0ee20c9fb4991ec434815b1c0ed380af3d71c32
zb346afc63343b63044d1345953f7abc81aa516b5042231b3d4927799c7d161797feede5457c58e
z45d409bd1f20c71d4d5f3482a04829d881ddba0075b41f8e25493503cb61012e93d501180cfc32
z57c0d22bb24360b2436d3763a21ee7ab2f769e05047c6c8ee050464b4e542e9a62e0ac2846858d
za2648e8c81b3969297ceb6ef236fd8c35cf7470857945aaeb8ac672d47423930438cacaea0c58d
z80546d49a1f4ac0669973bf9704895a80306402e5858d1b497d54145263233de4cff7be6a95dcd
z3cb2694b071d486912c18f18ca7fd5a83b7b66bb0f438b18095f2078a4a53ff9d1b6c3726143d2
z5a80d993152f9d4208765a315a539a9277ff5c8921b2b68ad6f7ca01aa246c0bb038907f7256f8
z3b8cc57d44a5617654ac9dc21c83be7492e7a44450dd290256783fd05b40638d567cbc9fa5d855
zb5331c8e94867b82093380b825b2ad7c5368f473e539cb01585ce28ad4b225a7cfce9f69080697
z99eb986494316bc0caa3f47ada74f5c9531f1429c89149c360a02fd2bf984e537c3f177151513f
z8e0a982ea7b0f1764dea4bcce70c5c3764701ee499b600973f7cdf18b0559141644f1b893429eb
z6e5ca3a0064ab2a1b315de78f9818a9d41d53ec84e8e80e99e4d45d2a532d227b0e71fe29c3987
z7cb6991919e860c5841670d5e56307fcc8077c82c00d04a18132675a170c838aee6fa3a2456aef
z9e3c5949ae2e509dd4b1eb2188016e2fe6a09c8e67e743f6ffaf1fb04407b5170745d74f8bf964
z69f5f5ceba336a7542c0c258b93716ed26378d3ef75d7bea3dcf6741b85a7f7ccbcca30867d78d
zda53bf40748b8c23213aeb6fce517d990ba258df6899b50c783ff0532fb32c152d369f67a5d15e
z435df7e84bb6978be35669588366566fa084cc006d2c5043a8744ea93714765a60ceda37abc10a
ze9033f18a397fd959d5324f2a402ec3764b794b3aa34e1c783211356064ca0f7ab4b74585fc0a1
zfb455fcc75b9b50b2fa766ccebc3d6bcc1e7021801945b9d12fa8d67a1046700fac3f11b3ff4ab
z55144ffcace2c1a23787db235ea578e62019650337be8290298c933c257a0b2d890dd9583d9f59
z5096848cfb5414c4bea2f1a3a7b5e681ffc8ca1e0bf9b348c8e84b621a7510d2f44283bfa7fe40
z77ebbf1f41ba8e52fc04b6654b2b9ca0c215404cd4c8a0174b84b3fed932055abed783d9e025e9
za3e529e1b4558e42c1f7fb28bcbddf51f88fab8dddf439ab4f277f2543d5cf5adb6e70d0ba24e4
z6c2bb9073513bbf114b0420929fa9b96f86fc83bc87901f5962b048a81f5b53b5df698af9e0f95
zd58f43edd523bcbd196e3355c3e0aec59c20374934ac04ae96cabd842131f69cc0e848cebc611d
z10efbd5fbb62ca00d50cce9358ba9220fa6a055b21c1807b482571f4d8fa140bee2db9098903ff
zc6a189410baafeb426d5ecaa43c3aad38c8f17f1ff2576179751096bcc87ab7f5e31503409ebd2
ze35932fd5c2b84ec264feccae33fe7a6e45b18659b87557cb476b2f76740fd747379acf978ae8d
z8a79a7eed7dbdc3a9fbbe9bc1849f14764ca88a0274d2ae28c2e56205ff58034789f1a033af958
z8f1f2bcacb94f8097da0377bc2805564f31cf792ad082d062796ea8aff07194f258d02b92cf7a2
z65bb2afe0c2c8793d1f7057fc8c245f769910c9ca2338bab24e9080b1353c4310b879c4e973359
zfd0f0651e0f2b2f4ffb587fa4443f2ab9e85a889d9dce80589857333ab2465bbc97162221f85ec
z8db9af464a7df1709cf95dd8194d8d6cd127d318cf8b82969c0c542bbdafbce895e8f103685caf
z400653190bb6e82257c33163a794b072db77559ed07603f6ad64b9ef26b6c5cbafe49d3fa44d71
z0cd194cea53ce69a33e5d2c68a7375d349fb190f3144e6368b418b42b48bdcae21766882998984
z46610369b73511861dd7563a1149aca19a9f88182fb0ac54d24f24c04ff780f3af509f285684b7
za8531c72c506842687f59775dbed32f0f53d4209106096dc158c580850c9a8b284da427ca776cc
z3ee7b91fa4fbf846d4fd637355aee085bbc609915c1bc6914033f94af199375873b30f10ce634d
z77d6c7dac2292e0c4ca3eee27d66999d7ee43e32ce08877538774922f7cb4c7e28334e78727774
zd25510e98c92a7f6dcdcc0748de795efe756b3d6586d1d85583a7ad27cc90a1082ee56ae3dd400
z78fa91693125db69f25d0562c5df06ad6c3bd7cd8ebea5df5b646c4c20a9455b2f4d96d21cf47a
z1d2b8513ce0b184d2ceae1454fe51440679ffd86d32a2c39788a8e74e2f265f0e31fdf0905e2be
z939a23337b65cdd39ec20a0ecf969b73bd2ae7bebcaacb81d8f1e41ac2a2acbc3950fd6e1aa0c2
z004533a0617decd547f2ee4b60019af9cefa3c0ba7423a55a8e538696be3f4d62b5c9220bd6c6c
z339fa613a424d77ec395a71ad2a1c2815f6e68d25826adb739e8237eba31662fe4f68604e2da6c
z5e995f6197143ed8a37c0a3d714801c9db726a73e6a0d9aa3b365a844df1ea91eaaaf2d476d452
z8001e6d4eb92baab8b913be9e900fc190c719e4d5f97c873dc8ab4cb998cc53c91a6021c9d519c
z9c54cbb7142598a6b2861ff002d3fff6699a61b179f302537f6a824eb60540ad511deff95bc083
zb5270d2b7b25333372d7cc9efd7ad4552ccdea8efb53f63deb38017a5837eb062a163c2e1af76b
z59be89d00820c6fc5bd04e9cb0cf09ebb7a84a239b984427f60234b751dc45405c9f92835e9025
z28e13fccd3fb9db12396fdea5182b9ae8e776f3458d4054dfdbf5299757595e973f784eb9e0ea4
z5531623ea00659739162f49c97d5ca0ff452568f3b7eb83136629a9e0cb72f64fa9ec2595debc8
z0be32d6f229902a58e58f171fea065a93508fca92b7b74653d63b1d3ff684a7c08f93f38c5c589
zcb6d3c9210b5152fa3b6db99eaa7c80802a376db0640bfbc67d3b30898d1f1241b29df28c3d144
zd65066ac19f2c949cede414c8dee11d715c52929d5e8866c7e2842044ef4cd09fc868571cd54e8
za7fbf74894124e9011eb77d1cecc8fa1c6a233a0d8d5948eab5c3cb1e13b4a4aa08538fba7c006
zc3057caceb4965a44f111047513459d4436f68e0032cc12b1504789ab111b97be167753b8a4a73
z1658029e386aebfdcd26700b7203f15c76c2c9e82eafe87965abe2074ca8284a92a135fdbda0dd
z7b11cd99da89d2f63afdaaed0e23792c006c60478543886a446f0b72e759ffed4e25f2e22f67d1
z7fc0d3038be14af8ac1036d8803947c741d72a275485d17ba51c624f39bbb7b7a9b300c0134c8a
za873c473623bdcfdf5496a015c5680a28414749cdcac5ca7979c196ce4549839afa953f4f11777
z06a7faf318b0dfc2edce6ebcacafb6922c28b4d5ae44a9e5dcbebde77454c6c53a7ae7094a475e
z9cc73b5e910b87513f4691789ebd40f3e8e50cff028d8dbaa257bd3a8d33ed4ecc44e1c181e0fd
za62aaffb7c2a14371c712826b693b7584f1320f4956c4116eb7fed7e513ae301d78d12193c04a9
z9d28aa734714bb6d9042ae29d53e8af9ea9f1f2f796db9a76d720fac19a4525e26d5c1597688c8
z1b145403b651c9d2407582e3c96311929c81828fa775270c926d06b756c0a2a439a1589b94d17c
z1feb21ca595e41295c1f3162ea54eedca11280e7adedc52ee7332ff8fa7c017d7c8e02f2bb7d4c
zc7162e67cd326191d76cff6517cf7a7e0a8f156bcc29f95fdfdfb176e44e4dca5e9c4d285cea86
zfcb2484fd4d29074c280c80248c53facd375e03d075e64f40c2c08688b2ab4543be95d05a4a340
z342e07465a9c2aa60ef19ddf3c8c558967f0c1678e93efccb8dc221735fb054fb902e2fad4228f
z034b65a5599d904c2f2079719386d48d16ee2308483837814f6af938eb9e80ec54613d97ca34a9
z5e656d1054e89173c89a52e0bf411616d772387b0b82c269789aee0e7a8cd0de69b5c953570836
z9620a34c3ccc08bad539092e705ee5dd25486c43564ca4794a78bf01e948ce96976f43ef9bb3d9
z7b9ad1641c472ec1f5e6b091824ea12ed6f89497d69ff1af43114e073ece031c735c46937075cb
z8d7c01d8e0b586c80ed0d9a2b4b1287b09610eadeae941391f828362399d7739496e4d451770a9
zdc77851a61542fedfc638baaea8e3070ab5712ef7a155eaf0f5df31ea9a827a5f61c9ab1348b51
z445344165b0191ee1e332dc5a243c4037c30ce72c093899dfa715abeef92d89026233c14c88f79
ze6dabb79b40ec3a836b885f0241230ef47582955638d145d0df6919bcc7add93c554a6674490b0
z3fbdee6bcb1c67b5501373c73053b429d29c062d0643aba11575bbcf4a428de0d8335a23718978
z1d7622b746435dfdf5a3b507bd6b0c1359d307721f06dc1147a9cd507f45da19e0415c079b46f5
zea88d5f551cae0f07a2ffb08b730b70be5f18b0da762e9b5b26d711439b1c9b74c936c78b77cf0
z0e68d1664621b9aaba718dc20e31cca4f0ffdcf85f460f537b706f0d26264b13028e3370fcb039
z4187e75c675fa731a06aadb70a5991835d7c70d5c2ea8c5564b7065031329f0d3af6c484294322
z7a74847eeebf1388cd0d643cecd536b3dcac8bce2bb3aa10d147c5db42791e4d631c4b83e08bfd
zf024db7e223f59a4f1729564e46a30bb7bc1245218a41c9d5c35fff21dbd59e581f4b8006a4168
zc762e70f5f010948ef2a40895ed7f352eb26e74ede6a7a55747f4b313628721bd7b18a123a5730
z9aed264c6641edc110344db50bdc0d02448a6e3970476297c146bef6c3c2a9d81d61a419a8aede
zcfe20d68e3bfab85f390fc3cbdc9a2cf0f8ab9a7afa148ec5a64422f462e4432edc0ec9fa0b233
zbb01fc7b4dffa4dd04b2e269381270a975ec7f5d59080d7e5a427c29b2fe69d5160965c29fa569
z53b65fb9b9f4a61dbd61daabe7222b71c04b663c8bf8fd844cb88bf1fd94ecdf9c48ec7e471f75
z5fbebc7be7aa9c87cbf2be2bf89e25b80da28e91208acb8eb89f49400e4ae73f0c02cbdaec039f
zc862c2a3ad33b1cc754c530abf9cce36aa3a0f4d4241d60884f23276ccb6ef0b026d8abcfb694b
z5e476bbd9f2bad64a0b0350ab837ffb779ce786e6706f438bd49680e84540e97af03ee8c97f033
z3fc373065c2a185216c9542f7f31b93768376e44d1b73737ff6f5105d92c52cf30dff3502d4d44
zd37e17e713718b56a7b5ca2e59081c597b054b35c109d880153a817f2844725023400a95e18298
z82847fca70571415aac6baaa88e1fadb16578d82d895cf366751d10248c73638cc62b05887f6f6
z572c4ad1b77c57a6a585c26fb4f8381d1d6fc8276e5b8f2fbc488b28d27f29062757556020985e
zcf96875ea2998f754f72af2828325b8839e82127335cb2261cac899ed2aaca7151945d31629c40
ze15ed4488e13b86ad4bc9b34dd91a6549307bbd89fe8285ed9f8090c8c817c0f0a83fce7acc264
z1f74bbf7c5f3fac852971047fb680677bebeb7775937ff775978f59ac413eae7d7dd42a19b8d86
zcf7042f45d17ad154a57de48e59d16fac3456a342cfad65a8efd5d3a6b0eccc0096eb361fee148
z92744a9735ded5d09bf4e80c3373ad594217d08361aff711c9320768649ea237d20a424eeb44f5
z1c06bab7d4afa7ee6ef65df36c352669966023a2b8b4d1a1ce7729d5ad5d773a900edc18e074a6
z7117e1aea793eae47aba078521c94fce10806cd405ef012625078e435e50e6a4fcb75b0f5ad31b
z9cca844193daf4e61be1327e226029a8c5fcd890a9938b90968b5256765845ecae8bfbe500d785
zdfdd8687960931598539d24691734c470d1520a9c89479393a00c801f851e88c8d2f8843f78781
z4666a5026b147a4caa6d11da2e2114d3b4b02bc4deb69682f1566e64ed664c6b58d642afc6f16f
z413fc1671c2ea2ecd087a1595499a96a1614f6b9044d227b49792212e9464d671836eb0d56d6f9
zf6fc3f3325f2300145510e4e56f1d61a56b73665dae9d2b45c3dc66cafa1ab4bd6d62208a89d9c
zbd60fc61761521b1630b2cd0a49354ec44668ba5f26ac203656cc63de011f6f4888afc255a179b
zb899754a8967217ad3ee1c2a5fc1e23653523c44edfd52835d1e79773433cfc231542c8dd1efef
zfc1069b42fd865a475a756c93b3ddddf0ed95fb89ec3b313384794ee8645747da7c3dbb478e440
z5dc4ab9eb8517b62e3c2b67b0ab5bbe2b5d07fc9c3e5cd95ffa62f31387e290169d0392854a7f3
z2e9a0c9f50469e90067e75ded0e8469ca2b4d24c190fec94b6c2110f57c7c19b862233d55da8a5
zcea8d9c96761479d0b5957d87a2631330e33967f528bf18a990fdf4fe5d9714610d30da72cf0d5
z26aa91a4133fc1b16ac9328812b386419c7fb8d5716c196ee8a78bec625c1b4892f2363e93dd75
z0503ba245d4433bd5738cfbd2553dd08745b1d3efb51e6465a2572acbc2a0844dc9a685132dec3
zdaa208ea987913fab4c5ca77ee4e755c60d9632f0677ed9cd711e1455e6c369eb6a35b97a30a83
z14a6c85a6e080d5bc3254341eb669b0a056d584d2d7341bc87e4ff43f4b15cd7dfd9b8018d7724
z4e91b58530fe68cf810bf814cbf91f66ef950f8d38d8ef4e043d872c39fd3408fa89c6ee89ba4b
ze30003266b052581769f2d129482ed90b2aa8ca43ce7e897921c121cabecb9c135349070f7d43e
z0f50b9c1e250ed6d7d260a51dfccb89c26da6c7f5a616f9e973d1e1cb4ac3432f41f7bf92a1a0a
z539068120ce4cd830f2a2652ccbfaa8105c462b6cb20cc45cab4c9986de189acf6141cc2058caf
zfd00089e841931dfeccb2d9b565c2b682ec0fa4e515f6f7bd07a7dbc6979ffd626b0f46dbdcc63
z51ffbdaa19dadba8b2a4d92e56f1eb64b7125216c1fdfa8943d378d16d390cdb087efd5c098f44
z9f957acbb555a5952b9e192c4c4784ead246a51997b8cfbb4f957262a4106f527e06a951f136a8
z9c5dfc508f65f4d7fef35dac06a87ee14029ce413b5d38cdf9458a57e9ce929699906d2fa2c2f7
z34eea22669c44f36d195b9c23e3efe26b44afefdefcd0591aa46d19a70d3498fd947ef979365f4
z2514728faf2fe127c5509337076e711b2b7d65168d2d432ff64be8b10aea768c7582fad76b6de5
zc053b70ed176fd4d8d3cb784f5004e8a310e739c4d9a72bb885052ddec0b3d9f76e96e7e42d5d8
z3bda90454ac905c83b1f773d45f6c5ef13af80c416bd0966647e97e40520bdd664e37eee967038
zc02a2d5fd88c3f4da9554be930894398481fdfba1e239528cdcddf7a190d43933d91f306e02663
zbccf52f5d923856e6aeb117f30caa820208805d9801f6d0f08c5c74f124d1927fe8c2361b6877f
z29fa025437968c1e524252ab81109bdae9558a728355d0a5e8ff975664e229211810f393e3652b
z3b813a0c69ec384e9a5f20c10ba252ddf5e9c4270caa5907d508a1cfbfd9ad013089c1288902e0
z96250bc8b283554d3f87f8151e85bc63330d20e63133c693b208973e64c454e40d1b7b7bd5f9d3
z789f9af1ba206eb7dca34cd655968eb367c118f8fd958c684bdfc0be880755e6eb6b440512ee7a
za1aacbc674ace0a22ba921aac8582c0298c2e70617a33363e574a2810303570b7c55b52b8e4814
zc2004dbcd9104e50acbade4389b9d32267d5dd3347a6ae78a63a2781818ed460e06a0936eaf9c5
z2339c0823606f532ede13d09d28a956046578622ac613c7b0d07e531561ad7d3e9604bdfa6653b
z5b260e0334090c3089aac22d5b13dc3a951c93201ec4e38e472a70877ca7db3b564a738f05ae99
zb620ac10edd245dc780a18a209c6a79187b91da2d2f03e0b2bcdebb880249178a33b7bdf758ed6
zf6ca19447b59bf159eb7ea06b3d6085f1f43b7897f616480391ca8f0b2cc21d22cd69112571c2c
z7b9b9e45ed2c01ba8cb3dcec4fafcd20ddde32ffeed95dde419f7f20a6f9f7776bccfc01c18065
z01de82e0d75f52ed403dab2f43168e7ab238284d92420140b5d6986b26ae3fdc41de3bd9c0d657
z0a5e90f278f1fafcac9d9054fc304ea99c4b4e217377c55f708f9904da836eee4f013d8f51a36a
z9bb7ffb603a5ccc4a3725f77b0db88f4d8ee2557d91454c70f6645324ff3256a0a502acdea3aa7
ze8d40a613dc868f10250606ac4424f4f051590af1fd1a7e4f06a2c34420f90bda7c5c3b7197b9c
z3f361b703aaac684eb121dae4e4d11bd8460b0d37822154fd348158f6fad8c61fbc3c52ee83cb9
zaef9b064f69431fd7583c0f32f40144927a4524c9e07c5f4ec0c7d9464d15ecd5df225a2ed5bdd
z75ca4278d67fa5ecb1d672b8a574267947a7174867dd7d9f1f3b34d0426a4bc0e51b5c84ad8990
zf3f399e355c08c0cb8b69c3664e0a4a768023d3547ed1deaf1e1c9055a4e028e871d87a85175e2
zf7ab8a50700c7b07c18807d40462cc96ceff44ef4808ce9b56b96df6df92569eb76d3401dec5b1
z8f398b649b0a178107b1b73b1966d99b1c6ebe7bab52c254481c4888a2015283cfa29e5ca68500
z3a1893d3c76207ab2bd6c97a9fdb9e8b83acebb662446808dcc773ae015d62aed73f4263a717dd
z99ed28f3a8feb35f12dd29c712c1fd41f876ed38cc5a78e0110dfa89b1d284fb57c5796059a02a
zf2f7d6c91a003a20248a89534c0a4e7c02721035aadfc0254232c6a6b9c0cb2cc69619e964d9bf
z39a045e35f4f2eb3805248b4d351d37db6253d78725dbf0cecd11802743b3bf2d7de61a2e58435
z4dc018994124a00c66dfdc2a0e6519313d2c9083beb3952243a987c236459d732a2317bd15e420
za542fe2097521169880bb678d09e0f1ef28289d843d668fc5980f3db5b7ecdcf3a0cbaaca8dcfe
zee8586d5c29c7c8533287ab3bae2c169944ec969471ea5d52a1c96df089eba983a48e66d2999e5
z8f52c54ac05716b799f5250949a7cd44007e9787ff577b85e1fd81b99b613da1cb23614ab9f83a
ze59e67b7dd7bd699ab0fffa7211978925b4e2c31f184ca82c5752695c789f54b77ad66a4fa9c36
z99a89cc4809822d35555dd5ce4338ae73d93e55dc4766129da61a2a8c0e7e55840aac7a4cd9254
zac7eff3672eac103d8ffbc53cc33ebd606ad6ac7d101bacea92600dd76d1fba85dfda9d2c76abf
za16efbd4f9a7a8f925caefab236303d79c22a95723461440dd41bc23b5678bdbcf752e05a9edd7
z2cbce33975ae7cb5050c0f0c5f725a48ec7f7609782288a1cec05859cc34e82eb12419d9787a04
zf8161b351fd441ba94b54226802136f2ac1e5721812e13be4f1125393e37ef3b4a5fa99ad267a6
zbcf32a97e2757174c2f9e8c310f4e098daa6534aec58712e558f00a4704666bd6d63e5b047037b
zde4fab749561ea02c06875c0f2b214fca77a5a13b004d1395602f47a7f849909708b0d25bf2668
z43f719e81a9d85268409dba64d063cc74891c702b871ff3a74d9f3c28427cca22b3084e0b1ef7b
zc2b9d069edc771e5f4880983acecc98e8400452b1c4f84394e4bdb913d5f6af8c08fa371443fa5
zf482950c688e06b9e900f006aae42b5b581b06276ed60189d5f74c04ec3e514a3dd6e3fb8270ca
za9f4adcc8bc3a51568128bfcb1b1e6ca829838e3fa53c71d4135378607defbbf7290e23b90e424
z9e54420b1ef2bf6a1c013c72ed140681ebc20fb4b5a8f0394addb9042e85709068eee9f397cc09
za43b411e3b017939279e49f72f2b09d0b7e983e17ef0d302457332478f15c8704b29e7266ea447
z84a3af9d8ff0c5ddfdc02f28da6cf7c65b6f41e9714a53e8ffd20519a8895c07d5c7829a943b96
z62fc8afc0381f35b53deb0a99a0ac964041210461611a0b439eb97da58b0145bc46019e1bb8453
z7875a8fb1d689884d34870912e6f4c64fb2942951087b33eda378ac53c0647267b3aa393ca9b05
z82b8bbc94ba635326ba3f9a5299f63abf42c62147d52b69e10c4f7cbdf519467b8cd3b9ca221b6
z9987bec0f369de98af0cfddac7f7aa9cd040ad710480e98104f8ffda27bbe633c1d8e3a22e8aa5
zff9227039daff8c8f2e7f2da4ce51b5a74ffebd316e25ffd7fe2f65d8360a96b73d43432fdf801
z42f886dabaa798667a320ef5af640247abba8bd613b8a776b460565eaca7459ff7474ffcb8cfb1
z1e2747fe104dc1bb2d039cab0a898cf1016f85cc514598e73619b4f1f37c7ae9faa999aabaa02e
ze4712a70d01190ad58f462a784e9f55ce36e52a80416a8c3ed73a6a14e9609d25b2ad316accf20
z0e90483df7e8a152ad1ec303d7f42fd94f1fd255a1846a0536361d7b1ec1018e5d93bc69772cf6
z9bda5d8f7f6e0c24939de1d315356cb53f08f27e0cbda36881f26e04eeb0c5d2579c7f64736e01
ze73077d89f3ca87e8f1dc77c2b56bdc24d549797f212d66445d62466c09135bb9f940524368451
z68b1f78eb7940592eef6eed47f5ab8671850e1b21c4a41a2c7c85d36cfe539323ee4cf8e9be521
z371536f09e95b433e8a98de23db0e6fbaae13ea7ba97c25fbb033669072f926af14760c6ffa7dc
zd423c4c012db69b414380fc33a83df158913d61b92d4eec8caea58d44ace4bad5c96a9056ecc79
z0aad1056eb68677eff7d72fb1727f78b37ac33a92b62499b83c64dfeab53df4048cfaf6448eccf
z1e04e373302bc1425fd4d54b834fc8d35a48a05b31ade01e7edddd68c2878c5610050c5e398d70
zabeb52d5afc642e8c53e5f53745753f5fa624e4a396a8148f093e0308199f5173dda391538af3a
zf86f5ce222de84645520ff67db10189851fdb705bda28197f9890452a7d02572c9f70d2ff0f1f9
z24b0f2cd4148ad8478f3a75da9c6870019e63962c7c7228db740a61d34e008a510676dda458053
z2bb09e865ef18858a21559a3f08807f930aae9f73860ccbeccb3a82e513b7318eaa9125257840e
z386c6c7e6e62f0570d8da27075307693a69db9539d041b5d72bdb0debb25dfebf408788510f00f
z725986a5a1f40d36d1525ee53e533518c79146b746642c1aaffdd32cce94d5c81e04e5b50689a1
z9aed1a5084d328b71825482cfe04050324e692a32052545f2f95b7bff0f16b779344bb3ca19fc4
z30a2e65dd536bf76f94f6ed11c63fef7723d140c4852bc2cc2829308902a5dc924aa50625bde0a
ze62be19c93e794e1c196c3565d564a69e72828f3e325bb9ec9d112df6e9085ca1080eccf00bb3c
z579fbd39dbea099a04f74452cc7ad8bf650dbe52c4987990e71cd2772687171ae7c83ca5030442
ze0272ea5c6546dc4b5f1d9630cd520ee00973aa5c73187b57ee6e1c9f790f8aeee0c75fcc5d1f8
z521a511e9e8ed30608bb75538a597c1580fa97e36b17eef545a6788a61896710fe0c8bf8899dd4
zc704f1c9608af6230192b2b1e2e465f199bf86305344675ae7a51b0fbdbbd51ceb879e4f7d700f
z35d420a79e0a869fec3e3534c9e03d666da00868f64bbbd77d41204554ae42d4f2eb0ac089c655
z62220e64369e718ba24684c8ab3b22b1ff35766c5f93a13ff23e50c7e89f95ec75cf3814dcda9a
z459cb1365bb70b667e1e45566dd26a2a6ae76f6362a3fed738b626b7b1924e7ebc464fff514fed
zcb1d1b27ca4267f7746c6f4aebd276924d86d043f8eb7e91bc260c29c6586c678013e38ce0114b
z95eb538cb3d0e16978579c27bdf3510c435c78333066abb6b161e8e438c7268f1547e9206b895e
zc130211604c0949ee9ab798858062bf1096a1a4f486731852367a6fbf9e71dc9db0f82e985c9c1
zf60a8d6569fd4e6ad766f708c308740e52626455cb80e8ede31165d1f44d4ca87542fb1fd07584
zb266cda4060838912910f705317192fdcab16161631d235d40c8f5435118e149e3e4d1331782f1
z8dfac2dcfa16d2180e4daab4e0b7483acc5592d038d4a4e1ed87b619ac71097b12f2aa012e12dc
z036304f5fca5dc6b0f9310bf44aa04cd059599e8ad14e0c187ed841c0cced6733575e33b63f157
z99c096e15d9d128e2f224ecf23aa0d36ccdb99319c17c0af198bc1aaa274859854f64eb9e77e84
zca8dc0882ce3ef9e5dd1f61e90ae43d21410f0d322f2a749688258ce8f5773b75623a400b131e0
ze7713cfe4fb3d4e9210df81f9d21173205b29168b565e70cdfe3b087d47e11c61b56e887e1486b
z9c9a69ee4b431835aca55a3ba6dd3ce54e508bf9982e76adbcab1057013e1def5b515a097f724c
zfe9c5952ad4ecb907c0f6e709da3ee0d18a3bfc4cffe8aff8bcf89b4e741c466f7238cc70124d5
z3f9678cc3988e0c6b2f6587d783c64367311765db728f8df13bb1f3676eb1e2432a970dbdfb974
zbcd1525cfe59f1344105ea2d55d11f74e48b3777fc7e22309cb25a07ea76907ef2a0d4deee1da7
z625cd98d36273d28666ee4d22a3b1c997c37041da9081bd14085629f9c47db45f7e3079d04a8a6
z17b877bca6daaa298e89ede7fe452b2256d0131fe19d770b1dbf25897190675117c36794a8c3ea
z32abff9f8ac40b357b145a53f2d70c27d877a4375a0f4e0171f445d7fb23758e68e50f45950865
zd95d32c1347d0610568dbe3a0e4ff68a97df0a87afdb1f170a2ec05a0800ed420db066d5637523
z6e22d04a41a1882242947654e76970f6bfebc20416e5c3f5cbd40344157d4adf4fff61527da86e
zfa1fb40c32282da3d5e84104ce6696756dc7b14a0a8070d56015d2163fe73028d5d27181c9146b
zd7af105a692d0a2a87f63ad674363f4610dfcf0468a5bfa91144075cb2c17a26ecdab17cc8977b
z151c5cd5f9b9f08e866d978a66f4d8a2688ade7e5619904a33e33907fceb2fe61de1c4a1840bfe
z412354e2dfe4200a2c93742ddb97c250a34a364dadc98e3411a5e29de6a62b9de7bf5a33ebbf7f
z714db84feea6349bd4132acea64a47ae6a37481be619c5ff45ae922e6981e78eb673dd1bfc0c93
z1047393a0da567d036f47a43fe2e2d3675da8c65661c7b93d50ca7981e9d3bbebf4072e2849fbc
z29d86486c6ac2217efef4e742ccb9cc9a86bced5a4071eb2efcd126213487fd8c07d17ec70022b
zb36dc97c6bb221f74a266338a9e9da4923c20f94cca49791e04b2d90eafe263fd5876f1f4d3d02
ze659727d4fc521f91379473c0c24190c1b1c06bd5b583ff95b0028c2e3ea595c56bdd65265a6ae
z27a5009acfe7734fb444ae49b7462d139a40e9de1d1b73ece264e743bcaf7b51642196b411a109
zb0f808871cf749ee9489eb463116fe7a2c0770f6b88809d406d19414ed3f65f90173724ed18486
za35c2d2711838c8f7067b8af3f8e8cc2215af3c7ad5e4ad66a299970254e3da56bfdf41c1b8ff9
z3c7f6b519b57cc74461d5769423b2d5ab67d43b857236ceac7704aacfd85ae4fd914ba33ad76f4
z06cd828ef1b364f6d6bad1c6df527c8f3c10972c5fafff822cb09063ae7f9f50140102e33b08a7
z01cb5de47854ed2b5f1aa3714d19729590e6ab426c0403f3dc0f10adb328e53c3c8082b56c29f5
zce52d25a8905ce029cba2adc94fafceb88d9144aaeb0c2e6991eb340a8c37837f88b13d8e67b6d
z5ee90e9eb6156f81fe648e666b7699b0cff4b0dab41c0651a6866470468d7c2485c96f7f0393e3
z7248e563b65e78644f76b00980ed2714170f1cf24f1b25ea3a4bd4d8b82f1c0e59b3a035ff4215
z1de57313c0e5623124897fcc12017c0a58ac68edd3eeff6b317399d5cdca294272b2b23101e019
zee18ce1bb4c06b1f9e24e12cf1d685159881235024eac528e31de2b3737f44d8bc27b1843a7dae
z59a1cade4911e9ae9a4c853aafcfdc5a5772c17604ed77f718c894f6cc02cd3adb8a258b9c94ac
z7f660b73df6179f2a62a99ddb2356af79b7b64eadf09b52ae1f702d467ab14fe60f536da536de0
z082e8d53337f205c18b92ecaaaf6b2491943d6d298d511b221d61254acd7d4b63677fbec3b04da
z94c68815bf4747d95075394877b28cc6815bc38aa89ea504d2a54d352f772b161772faba05f0b2
z05342b71e133c1378b6ba13a1c0067904b6056922f242eecac21dc4017f215dec545d91c6af62d
zcd7c6fa3fd077dd00eaa37c44cdd5b7ef1d11ca7242ae4854630b10e51e6ab5d2c2ba6f0d02ba5
ze92ac3740b23daaa6ff9fd9afb8e4774a652675a71b9b4d1ad242225297b684263466293dea935
z4eea21d94ecc07d6cbaab85ee4309a4c776f8dbacdb1f99a5c92b5b709dc317446aa81620f8d1d
zae8e1733a580ea9158e976bc557bca3abc1913cf30910367beccbc4d26cc9d5513996515b1a992
za39a148a3266a9c5187d99c5afb0c50abd81127555c0c20f0145b68ac62720cbce763845b7f269
zbbbd66aafdcf3861dc31b2b10531feb60604046c81d09ef1202a9ada02e644ea07cbf94f2deea0
zabd459f5a4184483d83f710615b0c882a52b94e008192e808f960a6848256361dd08933e46b426
z1a46fa0c725d228b370d72ff83b1f0c8d93ecd045a5084684c11e9c809667ecd467a83372a5bf0
z778048eba7b531e505c296d0d27240444ee88d54b4a94d5059d9d285e9215337a7603163145fc9
z37be46b48bc50b3adbff5183fbec0d6d6f51c76b12698679bbea6e5ac8248b5b143592d7dc162e
z5f64f24f98c2c30a4f4ada4f778095cf87ae7a1cf9aa2b2db05623d4f4a772eeeb8a9a068c7a37
zc33c2dff3a4061f62a4b72b2a7fc5d3fdff9832062e8ee775b63ee1a902ed2c5aa7f9c0ffdb958
z3082eba2e208e40c0d12e110ee68d7a846b6f477ba67c977d2e74584b836f85c527b9745f6b06e
z7e168030071f8f3b8f322fe16a93e9ae8ba43fab3ff001320a6c2ecadaaef357100c60b57bff40
z9a5f9d5f7e9a6e899b97e7ec10e55d164eaa1362789461f4ff6a5660c6654c21f148199cbb03bc
z37142ab5bd37233e2c7b1e727c71c58470ec87a417990ba31c7b09b2fd35acc3fce81adde8e456
z8103e3d69b5e5ebd59f940a2b429cebeac7941ad8316dd830ca9c29aceb60d3792f9455997175b
ze9bfe2d5fddf41da8fb682053ae4d97dad10c4f33dea00d52261b252f72bb4c94d139f7a02e3a4
z75bd7e82fd6bbf85d2593e16b79ab0b31f1bc5ec42ed6d8d2f86f749bde3a21cfda7dd18ea19a2
z1a660b1c397a83df0584cef4b7d12e36c98244ea3a0c5233ea93fbc56318576cdf1793f4b4bf68
z2ae695f71c87001f656c61329e37e2d0fd49b5072b82ccda3c340625e231c8c6f2516097ec669c
za70d88d6733516175f3aff31f7cc1a20fbd49064078e32e0a47f086bfd629fb2e56dc1b5b1de31
z521fa7d7aab7fc1343f209e7293e9388d4614e708edf548700251495ac3142bac6c726a77390ef
zd8e049506a58b3e502cda93691d928346660c875167eab74c6d8bd42f6f6c9b8a1fd2e1745d5ee
z6b290a716030eb15e44ac0ca3d9133f96e7684bde603b8bdd3d52fbe7e3bdb017b4a0a0f8e4443
za4fcc733350d46af5aa215ebdae6813b9aadf8382451e20cddc631074bf8f63104c889c03a0fa1
z2e5a77346666f491ae44bbdfa0d2fda0cc9dc8debb1dafbcd347170a89138d10cfe71a5a95de7b
zaaf30e17b4898ce70c935d921f882096e6b9cfd6b984e6a98298ffb9e000b72cd9f5d6a1db4034
zc344b5fc25b2c6302aac1b5c7aeec714f31fe2ae7c2e4fa9f7daa51fbbc4cae8ca322f95de7beb
zbfefc70e5b1b113ce4a2cb4ed4a8b74a3c35bc397679b3cb630109a6fc60cf1e1f6d55878e7510
zd45924017d1ac158b654107fe1f20c586d6d87618b35bf7859b604d64d0b00910dc203796dc773
z0ec06cc3fbd2e9333ec8d729469a793350b58b96071b96dd91173876bb40c74cdba580985b640b
z46db887d56aecbf970143f48442cf94ffc1c36c6d352456dffb19fa0af0c8cc2d9081960a5875a
zed97d4b3d0d34b8bb82b763382fdcdc0416aca4075bdf42dfaf9540c7b199795a1b8fe2978239b
zd6deaf8c474d135b1e2470dde3cc00355ec2fe4cfa6a86ebd015bdc44e12d7bdc9851f67f933a9
z3729b3a40492226a30ea91634c5ad85dd242fffa7c973e869cd3a3d5413dc2f424e6820b4d2975
zeec137f4a9ccb7a73002f74cead6e7bcceb743be46f8a1ef106c423697f9799098b298325511b6
z3d56ebc79ce56d8a36f63af089230ac6de1074e575cf304119e8c43c8462f1ed9f2789204973ac
z2de5335b8cdf900ad864490d5a3254eb52865e95813149fa19e2644123d2db48102a602bcb46da
z90bbb76860d1e3529fbc0060da699b9c6fe894369afab5c6ca5eab410acd3e2fe65496d9d43f8d
z2be300fe97232bf294820513298291bc2fa21d5408ae9b2e09425fa4ceb25eda4c8f8e6acc0c8b
zf1537b054f4d272a000ed093d45092050ade5b57049fd6e18ca9d49a2dc81b6d9d3add43776537
z075d73b3b60b4a837985074ba114d45107a5b722c633f7d338779dae5d15b4f9959781735373a0
z94a3329ed3aaec80a3003d19f6eb1322d27d9c7100e9bf1b685f285819cbbbf39a47ed62e8baa8
z73406fb497595464f6249d666404ee67db76ee8f370c7bba549f346e250525e7e867d9a5db878b
z35b8caab9605b861db57395f70fd2aafe3faf62bb0d26d3f6d05479d31c89c997c4d7c78302068
zb58fbe4f3497305c33a54dd3399fc6f47c2170f169aed273ae0fcaa11185bf333f17562294c80a
z19d84902c977b5a8a4edd83adb79d011ef24cac49ff77b2ccfb497c0f097d5ec5018a738c102f6
ze6e1cee6f1d09632d61a5ed940bf14ba65589da64669f1daa9caef8e893eff5fd93a5d87be9b1d
zc9e609089114709b67adbfa4e67528a571f6da1470fe58e49ee182bc0920fbe06ac504dd744974
z167d972a5b56c3e09590ab75ec3a80ef760d9c3d4eeedf349221aaa422b4ab1f421ec0b1100dec
z2b67125585cf4bb7ec27ac642ce96c9c7c49fd56f354f64ebd1e804aa1abf35ffbf4d6859fa0d8
z10c044e9d3e21f0abd35a5894aeeb7e3fd2307428eb25690810b1724faf47ee5b2ded2b1cf0cc8
z0a700a12d9b35c325b3f4d7eee8bdb2dae4315f629b7fc38beb76d9db4eb63fb8e12d5dac9f1b3
zab69641a76f0ad2e2030b26701e260271aacbe32d349811147f09ee8465e02b454a7152ec7cef3
z2572a8b059e9d7aa46b0f2f3b1a660d1b73c03bf27a0d89aa93f3616b5a9e0036e907a66cdee80
zffc2ed29d9cf00d0b32b8e33343b13bb1d1c632b16f73409eba65c1dd2acd0ac0460011538c1d3
z87be110ece3c8b4afa921613ec00133cf7f5280ad8244d4e9291be78b6951c6ecf9783e5969fb0
z7e3b66ff854cb3a68eb72a44f3639c42846ed6d0938eb3ae4e9cfbc419ee7344f844d181fa1ae9
z0318e3cd215945f65dc9eb007de77ca8c37cf9d9ae99b9f2a280e7bfec1c90f02c8795d57d4e88
z1fdf9d95e8d0ad92b0751ac851c437d4074f74d35faef0322cedf3145cbffeb40b439bdf8013bb
z976de911c5b465ef605304d5c698b10830a312c581dc49fadd01940328b2d7c02da36d0c20b068
z84a5409c7e7b3514577c1250a710f6cd54c9a7f1591c9972237555a8af5d45d408677614478e2f
zec47559f4e0323d887bcc9411ea74012509e55e0fa49800c6148b832a48ed5dddb489a4fb4b160
za030c275e365e2c09bc925d74a24bd1ad03dd818931d8e0706326d90ca814f3ed9b5cd109bc6fd
z9a195b97eb6aa1aed30708ba86e53322751e9abd7c670ea8d2f53c11642f4eb23fba2a22725487
zc187cf449109ba18fd1ad0a291819c05be82e670d5cf85494da67916b2d2091b7d679d7d3f3fec
z630b0c753c1d6a244ffb23da687d88b02bb099564070b8b1e8e0e11a12f7a4c094fb2169407f3e
zb2899ea3acfd7eb6aad02dbf2038086194cb32c2ac3f4069598d7fbad63bc5887fd9b3552931a3
z961506a1023538fc5a20919838e7008d2548ec9e9e48d01e7a85ae0df75c8d410f416824da249b
zd3efbe43734f038a6542d4ea6ac969d34c626e57a7f186fe1b791e877afd59f4215ba31d003d64
z9fe8c435f294962aa8d4ed3237aac9aa00b8e18b09e5751b060cca3287215c29b89e86549af687
z9aa2abad77b2fe79063a544c41233dd373b8c3ea804d6b3ee646bf4827949ce58b7c922a195798
z5f8fd909ca8e382753148d020311b59027b4ccc15dcfd587d6d952c6c6f248f8d4f9b27bb979aa
zcfc0d21774fc6cc7d1d1344f297bd99a7501ceffe791126ccbabd0fe004defb7c2f1378c576270
zb84c531ba120f8a3ff1d1830b75b5f6d2a0391202aa6856989e41a296d47ad0ef7097cc4eaa1df
z442468a2fcd56d3f7007cb30816ecc91818bcd3c65bc368c004e9a19c1e4d1a642de316ca69c1a
z6c226a377b992fc2e9f73baedbf5cb5d6fe7cb111db5de6578a7ddf86b8c286a8a136563f77637
z947c8215434f79b00ee42d810c4a088f03333f7bd2bcb0c86a718f5dc403222edaefdcdc49c67c
z5043c1cdb1403f7e3ed769ba4e6cdd6b623168026925084beac83909bb972e1a1d68b598f631fc
z24e1f8df4f23a6b35921186eefe81c534e57d9a3f8a1c0eee7b0aeae8c5a63a096fa4c73bbad50
z5e306252c2d8f244a7fc8ee3953d017f10e072c5ae0a724a79521f8ee3043a875fbda592d0096d
z27124cb75233f1519b4027d746a40f093b6c49cfe8851a160626daecdb434a885ba160f9259815
z53db3e6ddfce232c1306ebeb7efbd8045183bb2066c6b42c653ba85e8700d4da2a94016c20f7ec
z74bfcaae21e81a2eeaf0537779f6d28f87a65c94bbe6f57e227df8e23f27c932edfd96057d978f
z0ca798ef5f346b65cd7038f0bf0071749f00b755fb635010234ce38275845cf67227f682959a3b
z7215f5c9967c48024a4c34d333eacacfd22cf7001fc6d74579a9208cf11efe73ad032da5a03ddd
z6b7277331ce07626aeaad4ba8ec9ecb5cba8f8da1e310fb75355ba7481becbde5c738fd3b65e88
zfb438fee0608acd5af19be292b1e21aa9da58bcfb90e245c507cdcc30b1ea680816d9227431a69
z9a3b2e869e6e8bc13542d41604b87bef2e5748a450614a46bf333ba9aa76dcefa7024940fac590
z8172234e6629fa4e3d590a80b7a7aca48ba5e31bd4dde3d4f121e04195efa1723e082a86225c52
z4be07cb65b3c8a059c7d5810486c9eb92ec05683cda119743fc3b7c9c8f087d5ea11bf6cf3db0c
z6525f794c5a062932bcff1226af0e60167e6ecdb3275bd5d97ce7921f97b89e92eddf0efb2bbf6
zdb21f496a0e7d7e56300a338e8d5cffd6ae25be2a579900b789b513975bb99d0637589efee4332
z09ab3277d12257e192bbd5e9d3ffee113a0a4fa32c708d91192a47155f4eb7ab0602f45e26fb56
z42b6a6d2d149473fcdf371e62d4cb4eabd5f8b7f23a0acb3a8cb7a38b7560922f2643b7350f422
z0d1f200f0d6d121b33160edd5866947cdfb491c6fe5b2204802303636705dc458c2a8d08e1a25a
zafbb35156ae55f72243a4dfb9c163bc8950d777f9334fd3620cc6ba594b742347bf247d11fc31f
z61bd9d9484177039f34e8ad48fb12815c720e4d79db9215df8f7c8c29c291bfea0c16ab2ce6ea6
z01edef8b644b60c4dfa5f27beac7d549ad92409b5e8b09abcfac1da89834c12be260b19a1c1125
ze09b20b2e30f962249ce7816a0bf2ba4d6514651fab8fe504889e572df6e5c54491111656a19da
z6998aa20c1fd0c6152acabf4906a2019b3909d67382b5ae810a5b3bf7a28fd8adad0fab6d329cd
z65e7655e86ffd3312170fb1fbedbc1b7fc4c275e73885aa54952de74d426ee91516f630c31483b
zf6fef38d6d64ccb8936a11bbc520ea27def1bf682b67a71b35fbdee04c0a868e05779404af7e64
z0542e96e64afebd5528068a0bfd3589e108d7f8fcc60eede4dada0508300585296bd09e6e6107f
zb950aa13734bcd9529e9902868e84d47833b3f7e7aaabd53944c25e85c49e97892a1fc79c75bbe
za873d72582082b622eb04feae929a95e5d36ccd7255f62a2a2fd5075646467045c7c4e59798d6f
z281ce6c4f6ff19aca0e71517d2b7bdf8464de4263625e71c8010b4b73b1b5ecd54f54a91cb7faa
za154cd9fc87bd5b4d73beba527c497b70c27c2aaadb17b0d71b5190d040bb3ed8a13ae73279b08
z59961bcdd252ec1f836b9a1c66abb314395cdd615b4a2a590294439974482719248230681ba3b7
z6d930c97b0fb3dad92d1f470df368904821dc8344a5d7182ab2767e73a1637b799a42869cbfac1
z6c50261f2ab8a5148f698ff5b8dec4817b41de8e88141337c86264a1517c9f451e5141cfb1cc07
z923af6ca51e0e89baa7b32955a2860497e08ad466746c131e95c30cdc9ba9eaaaeee4e31171192
zab38c748b079f13351c56915f94ea5731f7abc6f3c937528f53d792a86283ff0805e51750a0860
z7a2c7b7a18c0bc00e30e05fa44a0a68fc555403de0e79c6c6f6983c8fee0c38aa9cb8c81dada8b
zb65fe1ba71b87cafe7a8263f3af5cf94db40a4da304fcb480a8ba7aa1ef0eb113c0592f70ab393
zfb146a4f9219f81d54773b4d96e13fb2739dbefff16e88c591940efdd8b448c0ae1fabd19dac25
z89faeddef2a1e9c4b893ac499dd8153b20105aff41bbb8308a53e98455002e864244e73454d809
zb5d6b220d1518964c0894489ab562b337faff6fa25e04d081144b0f0c15fa65599d1e4dd38406c
zbe10580f2a0f04955b04166f3143f0ae98cc2cbe655ec3ffb4d902af095a1bb6dbf08fb069449b
z4edb7daa2a34129ef590ca686a71f918b14adcf2e2045fff12ff177cfdfdde367b5ff52798bc4c
z49a5d1f810eab7c0cccf0718598fd565f6f7b504708e63c0362605c679cc7aaf0539c5ec2a3274
zb1e05094a8efc566339b67e2dffcbfa1c06e812deee4d1b67e631a0c4f56a331c4feb97facd751
z86e3133603103a2360b061d1df4c2af2fbb437ffb1458ad06dcddfd0e4462cabe932cdda5c4681
z661745de86c19c1b7adf5b07be735bba6b87c33c432e24494287502e1515f9bfe68c381d00ad8c
zd2021c00d68e6b40f06e655a37e4b9c06d678cc55a32f15e08b2f9e3b38d51507558d91be800fd
z11c60aadb6c97e70e8d6b6d5db3123cf06ae186afc9d9009b08bf9bf2cf674230584fd0ec492b7
z056d1ec6381697c5c6ab15eaeb46e71f10ecac9e8b937b29e278544bfb54b218134f5bd1ae2e82
zbbbaa9c7e133a0e546827ddbd915be0e9a4200f801b2a8ab0a24d6ab5ee7ff3673e66266684412
zc6ac413bfc4fe3463083d75e9d7bcac36c5c081e9a71865aa284ccb650a94455da57fa0b0c290a
zea70964fcf9622d24372080ad2d2acc14fa77f5f72d4e320c63762bb847563420005404af497d0
zfba0d96e54de930c1da8e96ebefcda11abce7b4e716e369e97d2738a582c13d9783b504365ef41
z1d19894bad722e3adcf35fff2c2b3b3465092df8bdd6d80c21de6a01ad03038c5d23b8a138597d
z9c1a36c8dec31e5f9306961688468aec6b469951f48a71692ab3e3b668c71ee9342a4280ee1696
zd2a0437a046bf294901a964e5ec14c86224e887aa0326b15463038b09ddde0e0ccb7f65507ab38
z0e1b83ecc3672bf33fa1c2a0decb652c00a704b061f9f4563051f94584577039cd95ea9a21780d
zc105b2cacf558ff7d18f19dea25d416b7834aed63a3176e69ed1bdfe5102c51a4c9fbdcb7d34e1
z80e3a46ee1bbc75e99d22b704ef8d17a2005389baa0d121ac0fabcdb03d30231e7c30055700678
zc8b5221b6b12f171bd8c2963ae3e8da81e8c06b7e4d2ada05d5b64a42555d6ce3a87f3ac1f266b
zf14e4204c12721401444541eaf93c1edf57e4459371596d657d281ead9c725c27739998e87e436
z2a1b6e6f47c067d4813622e17596b87946540d789743d439d16cece014a12a7880f34ec9b03e91
z57e59bc232f24b3d106f22db2d0a03ae958afd01e114affdd6f80e0abeb14aba08dac98c497296
z3e03d0a3a9e5d7e55f434673e01b4795a6c30e9e5be5036ebfc8ad18a5aefbb4a9cc9db39862e5
z53614d237b4f2bfa1e5ee151acbfe0d95088a9dbbce1af63131a045226feff1f7b797b8ddeb8f4
z9ac6ce8d44f163f6e777f340d29f9e38ad8c457f5e04c5f720bc4b4380adc9401c88990b884b10
z8a99dcee86df874e6938b3debcf54fc4a88d0eeaae4a14f4a537f2b42f172c2f153f69143fcebf
z1171ea47e52289abdc67678635f683177798f9c7cb0ed840e97dcd4e6d0aa6fcaef47a68264c7f
z00f553ed132ea3bc798491f1f963e7d79d03c99701f1cd49cd1518a1fe60bfc0d7c9c5b571a6c7
z7634dbf780ade27193ce8dad333a0fa8a0d41b163ac0d4ed7d9cc07499b576d628705c5f08af97
z96a231c34b498a2248a58a4d8617fedfbbdc917d7d4fa68b7ff8485d16b04af1c0786952dd4b0c
ze9c8a6c8d5133d1848d97365f1ca7ab34f5a5f405665b13e3b1894d8bf2b6e4c3e3a621bd78366
z05bcfe56601d926b97c65190e4e7923c27468d73fd029a22b9b51cb6978b3391f69decb4298590
zcb127f2f61d5b230447c09f358e5de334c06cdf6abb5378fb39872623e14da72c36baf8311c151
zd45f8f29c87a1cdb8749c33a717864b465b44a3a3ed47268bd4225414a63a148678c4e58d29914
z02b0e5787ea7183575a86f0fede4a80b89776d8af8dd50e842feb30c9203e530732c0fece4ab66
zab921633d2bef81679aa1b649ef75c1fa0df828e7d0c2dd6e6db3a1a4c42ed0d1121c51f6fa2aa
zbe381c12ea8fcf09a80f16ab82475676da9e98948f56a6da09ec5897ed87fe0e13b7c1ac8f34d3
zc021adc62d62c4f3b139ca8bfb102bfdde90e9fa1c64fc0458c3da9885d57df9bcc61246a80d3a
z9ccb8beaa21f128e49a8493e5bcc60ffa9ee8a941dc2bc9bc8a4cc6c036fab1bb11dc4029cc2ab
z68857046207d278dca317d4d527d52364f424ffce095464c952ff5613e8457729de33e64493adc
z301f5803234a0081b452b7a895e62c3326e6bddde417c7de9cf67beae44047543f2cff51d9143a
z81481a1183ae78e674de3c1bc9ff5f7afced46b17f64feb7865630d5dbdb986cbadaf354c10f82
z38d627051773d281ad4182b9a23df88ab6dd19a5a12dd35164703daadd64fd8dda82e63f9ea7d5
z948fedaa99cf74d3acbc5ea2419a49b97b32d826747fb4d052067f11e4783c9de5bec5e48fcae0
zf0a164d5bbfb40e9744a35528e53084fa83331a451f2e1f7ec99dadccef65aa191e785caee40db
z8399d249213f181c2d0227abd325ca0cac2dbcb365ddd0009c66b72b5915e12d95882785d4b7ac
z278fe5a111e7b0e7ad0439f298735f2f62723e5e483e9dc01b869175b224db8ad90e02b9e42a65
z768f2c4612cb5e2b8351cfe6a5ab6a17bc3cb57ffaf1ce902f43ada4a02aa9e3ad0b43a0ed6c6e
zbeaf28ff98ecd17f1aed10db36a33fbdb97d21c90c9b507ebabedd74ef0a8d2dc3adf94fc42df8
z48f9993f737742e577f065700a1b84f55eef55566dc1d06ac1590555c22452a47b7d7d96a5e820
zd7114f655a6a5de5d7a607695ff242bbca24100e67194de0de1eb953cf6ad4f75e93bc2ddfcf34
z8813078467f606ffde8fb5f90de3046c7d8f00d3556b0aa194f7cde499a61cd266a2a82406dc13
z140f41228f347c7844c8c7814596bcfea48d14cd7e93adefe581a02964e66737805dddc6a43e25
z249203d4abf92b69c9008f9d4c78f9c4bf0fc845c6b3cef2f4a34a5e3c2060d2a1c35ba182ec11
zce8a57e7d63a1b356eaeeac914d5bc96cb90c344512fe9394d7dae7707046c89abab1c90c11400
z55630194a1f7e46de9f7b9b1898b1bb29f9b35d26e093acd3c2978355e3b6281ddb6c78b93d066
z63812050326c73e09fdcb946c22f9b7e85ab5a5d792743de7238201e674e9e7105203413b6b55e
z355166d3ffd7bf20dc350f657d97a65f07e90322c94ab98a69f2d12039af78f476c30e48d68803
zabf18299b2ee9756e0712dfc9b864350e144e9d263544f22e6ef07f59af67f74ab62029b5f2e2c
zbb63d1a8583d3a2d5417385bedad824f2d912c62914eb8d01e858cd635292592d79fd85c27bc6e
z8d86a86debf66fcc790a4e21f0ccc1398d39672a944fdcc36d29586faa1897b47a7db7ae58d256
z0677a8036b10740e056ddfb69426cca7cdf3d83f0e0830c5b0adc953394938155f561d8b94d4ba
z1da5286763426ab31b147000ca8d7a2fc299752ec1d09584ce1c78d7f612c92b56e67b2224aa3a
z523568cd05e5935cfdbe9dd53c3aaf31b0a9bf79d2bf9d8faca1d30be16af9a48c6261553ec61d
zc79df5e3809366bf16ecfb3f53e9b3bf4812e7735b1c8826a9a95ae1bce7aff2a399e2778adb36
z49600b8565b98656c1b02abfcbf3e08f540d1738194b41480dc5e7ca5817279daf3c957e46ad9f
za773fdef568925d55ec123312bd2a979d85b6d44bee438dea14ad4a1b9ac8df58e7e9d521a971b
zb21e36f5d70fcb085e1a78ad41cf7f978c799674dfa79bbbde3b2451fb5e836a459539c9802396
zcf96d0e660946f1b8ee524cc1b6372bf6ad14bcd91fd98f29dea1dd79e17dc25b9544c4c94d91f
zad695af46ebf3396ac66a155137b2d35d66834eae64207640f6bc528e80063e9739fd7c6fa0700
z6ed3370192bc72f31a1a9286513af0830753abc48c2ab1884586d0ceb30ee6598bf91042ea77a0
zee29a9caaa91e5577ee293fec64f967181a4d3b15455b8ccd733a7ecb20a9ddb8e10feaee67d78
z00138cccbe26b9acc1c803a8f3bb47980bc18f3f1ee318eeffc7548f4899ec3f506f590247da35
ze27d9f05aaf341433e189291ddb1e6108d12386ba364db14ab52d070ee6641bd228450cfb90d13
zf7911574dcedb0ec23cb72d5c475181f5a09af4700b1facb95314a888154ccce7f855b31715703
zfad8051d3a684f2ea6ea708adeb0eeb1c692eb55c21483baac0e1c4256d54bd1294a9699cb8c14
z7ab840ebd22b0e60cc7b76b6ba296a70f859e3406fdd78f7744a61a5bda51278eb6c9af32c2e47
za6929f1a123a46fb2de919e5c0f671b5e095f628c78a227b2fe01c5a0f669deb6c04d330663f7f
z91a8669f8f84c954e20ff202e26475ade27df2cff1a1c0680f4538b4cab94e9f53c20635d6c533
zdd6d8f470fef1ddfc9fc3bbbebac07368aa0eb661700025a617e24957c02d9d4d2ec69bb663687
z3f8847ff635e7d8c8bcee4d3f494651524ee0b3dd70d3ef26ca7ad8b228589e5a49cd2c987da61
z9209756fdb47a88b2649f4f78f197025024bebb1c51f5bfd6618194991af666f473b34592883b7
zcbf76bdfff50421ce855def5dd655cd3d64245fa928619209beee8c6649282f19185bf0d6ea786
zf280404f34aad20bf6c92f84e3c02e770ad06bbbb76658c4d054a77b98a060eaf1326490b34cbd
za628a8aa068aa8c07d9fadaebadf46222e28e0a6a0f5d7fc64ce928266b050b963666b6fdbc904
z121810cb84242bbacc37d32d0b613372818bf954b3d2290765805a0b5422a06a6a33205157c73f
ze1e7972ab65365dbc5031a9c2b27fb73a4f4faf839ed18bdfcd79c4c2b84a68f0d2b7f3a63218f
z68462ff5421fb334799cf6081c06047b5c94b92814d2686ed2b829eab75e9b2bbf2ec64cbfd9d8
z2c177eadf7738e1e2421cc01b1b5504928ff02d430a71fd81ff71ccb2fde8064b40bafab7ddeb2
z2f25116a4d94d456746410e69fcc0d65381c2c32759a439eb25e2356a5b14f5802c0aedf6657c6
zf3dbfb515b935d6e00caa19d6d091167af9baad33b6a85703e5e693ec009f142f256a8653ef001
za7aad40f28db684a9b1bafc58ebc8a53b6017b3ccd2feb0771dd3dd43dcabb71b50ab8bddddf05
ze3d2c60520ebd65263365b771d0027e06e5b40e6d5b784be5e41f17f383bb6daaa150a2dd5713b
z4b73366313ffaa2ce82e55b5ecab8d71d70f7f7ac7aa0d2c3c69a92a1326cd5d9c28adede93246
zf9e639cc3493e1789060871ce1fb50d1660fe3e4a47aa2fbfc3797448ca772658145272721eff4
z08905b7bd3e65050df55226b0f7dffe84bf91b59be0e2c8b5de255068a1ee70a6b1ba3695c97a2
z98f661a556759a37a98fd5c5a08022a135bfcf47da47c13c0b2f1d48203185b02d42f08b437276
z201d7ed9d26746b1fe170ef2148a094a04483c5e2f0bc6b06c88f78ae45258820cf817fe590dd3
z8d748bd158fc216f8d89d2eff14130b30341cc9439f8707cf4f60a08998163ff9caa2fef941839
z7a056b67e6e76e70a5411c00dcc53d5bc896e897d1171e0128c301dedc1253ea8df2f3b2d6465a
zc49bda91765647bb9eea6dd305dcc56ac10227313de9682346e29b3948152c1249f2f2202ef317
zc149468339237068d95f2421426160d393e2fa091feb2641c4263be43f8a20ae4281eac6de6c75
zbe9f646c7c0d48064b498e4f1c0d02c040cd2aeb05c0a2468da0341fee9c60d44715be9ebfd723
z85ba732096ef292ecc1dc3e12c2b1976d4a0340c18fc48962244f3696e6174b677130bb6af88e2
z6804507e7e5da5ab3e8b2e04f3e4f76d39bd74a2d681118627a359bb58098653e5ec460f5a28bc
za9faa9154f08f43e74af6358f98755af7d57f390360d6383cc6479b61df815d2b158c512d8ff4a
z944761fc19e0f06e4a386ca31867c5ea4961f8c939082184fbcfa9412f976a87a200ca95e49323
z8edda34d8a66b1d652fe5d582613b6e2a1936e0bf8e95110e874e70c1249b222f39ec200b8152f
za4d5b2345f3a5569a173e424f089927d50bdc50d149dd3d8d07b2f187c3335967300fc7cfedffd
z3b299bb3e9c63b266c249623ee801fb6b3526dc6fe26bb45c5c2ad0c9fc27d13bb4bafd8627c7c
ze963c68358a0319c3ee6b87d5cbbc09038cc0e8f6f95e7c327b32a99b30648de4e04df45202783
z231a3b5f30054a19d4e13ef6920524ccd4ef0b4dc3e7da9178085a75dc696467d4594fc3725f88
z8faac33f0650974b6ea0a4201f0845e2d1f62ca6d71b76ee76262688f2d3c1fbb06cb0afdd6a81
zf4a37f18acbe7fbf2af6b0d92ec06e0cc83965d5aa3d26d96e8adcb048f90d9227e59077e7c188
zeb26abe5d2f10cd3e3e242b511ef34e6d6a20a32d2b8f68b5153dcc68978c81f056dde24ecf9ca
z7ddb2a4288f6e872b457ff3d1a0a94482271a3a0dbec65b0a43988b7745a455d2a72f770eb23ba
zc6381a19c9d64b2849a51387581c92d8a4879499a1758e554f3aa3ec63b7c2a0af58dfe1c578d1
zfd8a685e54e56672c92c67b0e98f445c76ec9c235a634a37a29f92a1fb839db0124e11e9134bae
zc2f650488df1ec0760d28fbaab473e113f1ccf6dee18753a044f64fa7a16629a89bd0b6208da52
z6d188fba81e780da76db21eeb102370f008638782b534bcf97c4489a43532373ce0f7ccaaaadd5
z3c5e782093038250cf46293fefbd11c0e06ab4070c5cf15d056eb95d59223ebc6999c024b00e18
z85aed088f0509c39e48b9cbad74370292edda82919c033462d7a78e6d5f9382ba2870c909a9a28
z56b42b86ce3f65e4b884acc48bb4b2b53ea8d458de77e5a0225981e429ba945d485912f6a1cf25
z7bf93c0d3f9d1985052ba3a5de7ed2eb1a66ebeb8703e9bede7de11c435856192651821019cdff
z6172b691d198afeaf2252f928a5a6c3c8f49a900fc7cf0a6352fc6e7987800e8dfb83207f705df
z460f150aafda6fb065541fb58c28c04a9a91a87d554f572849d290973a808b9c1b3bcd0492fe7c
z7aa7ba9b5b0c9d6631853e017ffa45fb68df4609160e86b01257e09e890eeefb006c7a7972a037
z0949a09de849e915d34ae1c4e7e5b3d63913d3cc18f7ade9d90e181c71aed5b944454deb4d8787
z331ce9e5619e7926e3667ad589ab7498049d64222917aaa4b294aff3847a1a6ff1b33fd9164b96
z6397bc0776f0cf4aad156108d36749bfa4bc73687047b84e6a743a3a17da9243a0adfb535c661d
zba18631484838a3ea5e20ffc78d758f8d8e68d30f06d6d60a4ecb9051735b7f938f18154097d62
zd0dca8be8fbeab413143f99c8002c2eb4f22357618f1ca8f8d289b4102f307b7860029a44cd134
zbd4b7c2f3ceb4e86740c8fc6cb4ceae0e5015c364d32fcff874f0faf224e3f07d174b7da0b916f
z85c71782acec3064d3a038377f82e85a6eca9bdc3d080f93ce8d6a387d75ae23e0b2681074dda7
zb7c7ab735084730a8ce5203e7004dcaa5b48c1798e7e755f5d65125ffed7e4446230ed03a60d30
z99c7308bb99a6837adb9a507678c7ead80f26a8238f81b6dae1b09847c6d5ad4c4f15ed456b371
zf43b91f5c2ac6aa4c118c68d5caa69835ef035e4476666f9510a0863152623a73cae6ef107b023
z6a866545653fb36c3a88ab87508e52120a01cab37043fde5a54488026973695024fdc45c28aa1b
z4103ce4ba8fe0e0b8e63954d9dc1c702c21428950f28c9564393e988c96151c80671e59e83b424
za9cd43fc7d48a41d763ded012339c4bf9955f0dbbda617baf1dc4dd27bd8bba462a04b9804fb58
z8d236074974f2c5635d2912d0be80cfb64459e18edd101c95c1fc11cb362025aa7fb46ed80f1f1
z52bb89abcfd593c1633882ff8485153e9ae95949d079f39a4b39b02623bc9cdd6171761455e812
zddae7763c4fd65d11a457d51bf9cd1210c1c38abbae7cd706389209fa4c9de72757e68ae22c08a
z0c2b8279f2c9e965d868c5d48e70480be0fdd1c6c800c502ab5504c1c2a0e90c2ba173baea7d39
z9819fd66528ce727fe87fa23fa0040a4c8928b76416392884d4263582e6cd3ca080fcd62af5e8b
z24a16d09ad94e00686dc4aac8bc65a0cec8f1e6c0711bc2db7282d8f91778bd3bbc973f6742e14
zffd41ac87e939c3d93b791de983c8e6e6204fd1ce9705e03f919b20776e9880767de93186374a8
z347e67854a7b019a1d198b8d698ae4a1c3ade6780b61d15a7446e774057ec6c754e87c5ff7dfba
z12a3cdea2aa7cc78ce84c5ceddd7a282d7b11cca134b5e30c8f3bb2118255004ba4bc127ee362d
zedd9218f490aca922802a26f1c907d1d7618ed17fbf18c3a4f1f9e7519385b91fc670784b925ed
z8fcd5a5ca9c8425b27d8af4ffb1f243d2619fd9c38cd584f0839c0129b95bea1d46c4f88bedcbb
z908b02b6ddb49f30d6bfb5548713d60775e39d73f16cc79104246d56d0720c4fdab995889f8f5d
z3e7341e9cc6ac97f955529fe259a9996daaf8385330fbe999ade44dc224be181693c5d42e5dd3c
za6c9387f193a9f975bcab0aa0525c43954ec85eb84ba87e8089a51025d1bfb929ac8d360f2b71d
z6d6a19c2dbae92c5954b8b4d11a3b5752b713c752d4a8ef9aac825bd6bea002d9b903b73a5efcf
z3d4845f9efad4d5faffd97af472092871f32737c598d6b7a8fc9e7b87f8c19c6c90b27e7d3d2a8
z51660b13c2c3ebc4bece48e8abbd5a4d56362582e519fb3173c58d1123d14431d094f1eb1f3a47
z8a29d3843aae2be5840a671c7d401b8842d8742a459f7e33e32f16a04330e46b43b1ded5e10ba8
zc93c42f4b2d91ab81f06690143f9cbbe8b7c7ab52762b16336110271c6a58747ab7d102d2de817
zd302bfbbd2d6ba9788e2aab298c0bc6f846303d05eab3481a0d5f1fc6c0c519cf1075ad8a7958f
z8ae05b5502971112dfbed9d5602c8d6d7b6548c1f636ca39df512807ba2c27af30bd0baba49d19
za2bd858578b2745325151ded08eba2d3bef6d5eb2ef98138239db249ae63017e6651500ffa78ad
zff142c413d9eaffa59758eb025e20471adf05877795ddd0c1f066d0fcdd2c80faefa6e82ec4490
zc6791172751e0b7a3850980d1a900ddb7b24af5dc204dc6fe65326e9db8fc0387bf7c1393b5ccc
z57de6f79becea73d3858fcfba88790c39448744149e80f275208f3af4907d69136f480f142bb13
z006dac94bf7759bd762a1b455a19d0741e83aeb168a94aacff207a1d18600d338694ca556abd11
z9f2b49185543dc7dc5dbdb06494148665a22c74f1f93e0881f4834b06c6992f13fc3fa2fec5c27
z74f381c5cda979109710e34248d5eaf851bc789d19a1034f4504fd3d0247ca8da348d0b67a95ea
za440753fbf64440a9efdb66a69d8d2717d528b15d16ff3f4c603f4d7db4eef65b6f3b9e3b02357
z256e60b0b10e7524fc3a289880d84d0804e61f26abe541c8999533addb45bd413341c3ebdbd47b
zed48a6f04e7fed7a714c7b84031e0e2e4529e9649ebdd95b5ca9be35458757e199906c053ebbce
zbab04104729277c16f4f48b3445d3b0dce3bca4c3583d605c5063bbe90c95a93dd4e54d06e80cd
z708ca7418eebb192e7831aea5f4815b0a1aab6936b355065ea8492062e72d7af192efd9e21869a
z7ec63c52807fb3ed17c5dd2d1d8e7d0f7bee606bc6058febc9603318af50b2d2871930bc5eedc5
z1bb563b8c872ae0345a601f4b429eaadf122485dc6053e34dcf9e81cc77aae8c70e9f3910c3814
z94394d3f57ea6ab99d4e7a4b4b49a33012caa02d36bed5701c51027b710b5d86b8ba4a853458cb
zc3a32a9375e013aa41e187691388ffa10168b3e41146cb79153259e467f441450a9d9be63b0ca9
z6742a444e4d088b3d6b0116f028ca79bef8f67fbd55dfa76e47b39c45a439faadf1f762b22beef
zfd7f33c59979a6c192edbca4fe2087575d9d57a24046156ee6998c96ac53141e9b9a53329b6a29
z50cad956aa1b3fe961192ad6f4463af883d43f58ce3d5cedeceaa20f1442fb93eb834566e62160
z0e1ea4d97c9959364d1280b39939cc9d2181b6cdddce4262e8af08693025fa5d4889b08a8d1db6
z3aa281070eaec8705a0218041a5275ba9c18741d74d8179713517d2481f7f626b4df4cf79873b5
z8ed229f3952630a341578cacf51532c8b8ca34158d9742737380f53ff85869864cb7621cea2a54
za094342e83d27a8f68d8241dcd3413051525fdb42bb9d0457fedfb70c86af457c6e5c67f789172
zcde7d9d94c4e03952801b6dd3c011d8ef8c53d8fec2fe204a8c17372dbb00ddb84e20d9734edf6
z5c1ebd457f7642b2bef558f4b93533a5efb46f6c31ca7a3b28b0d464fa39f9b1eb33c5fc3db22e
z7e01b645bff90a21422318479322ce8e05874d7b2b97e8831c72786a1e915dca07d8464111a560
zb188dc64ad302b1129eb2a88fb30b4757f6a3bce31b096a5a7145180e5ab490de6d79bc992e323
za12bb755c6eb5dd42a6a9164ccde18c803af7dd79925d2ec143cb9e250e98418ab33bd6a510d50
zcb33bd9143dcf840ea872d7ac506136213a8df3c2c6f086dab09fc6aace244e1268b80deb2f671
z7395e2a48861a8059509706cbda5814fdfd932aa44f1a704c82c936bd3dd4768232331fdaf9eaf
z6a3c037c8f7b96196214d98b365f70b9e1e2cca6430d7514070a1f5b05627ca65a928ed2c47b2f
zea01854b225f26e79961d0870089ab2a5f3489b5cd727d12a0f435e31d567330405665f67540a7
z9e20129d9aaeefde0d9f005689ccead8ad6da92b457068829392ff5a2bf5b00ff7c5b8bee102a6
z152c54dd909a1c4db8993d07536f5591655b9dd0b98d6b5aac01e05f0f3234254204cc97addea4
z1115a7c1f28e73b6f062dca675babaa790183bea4af9442bc5b90257243bd359938cfc413080cc
z391f1aea4206c82fd915298d646f5a0f749c653be8b886176141897b99fc798421ca3311895449
zf86628b2d2c2cf4fdcc341dbafad21f898b0dc54e59f9b14fc2b9380cd19ef82c11affc428b531
ze490d857fe26f08809dfde95c70452105981554809216c80a08adb6fd8125fef17353668a142fe
z723a354f7601dc7696652eaab736256e77a9aa32edc987250a65f3af5e9cba87d08727647dedb7
z62b20bcc9196a355feee393078f94a465ec03146c08efc421d5a3ececd1eae73d8162a60606836
z3bb2fdc9d2d6379fa9468ec8d8414546ffdb5c25f15bb30219f1adeab1923891353bcd76e075d0
z563f8e4225c720c3552e017e7222434d6355412ca12d4d95b23c03c15cfe563b376dfd9f1c9f59
zcc49b986bf9b1c50c4fa625c57da5571f595e248afd8e3a822f06dce42bb5cac7f633e8a8ded08
z8eb591c82ba01f0a88067eab343eaf1f00b6152bd18d6953419c0fa9ec9e4fc840b97ff24ad153
z08febf119b11edd4a52a0319fdbc2156390bf571961f1f3b3a9cdd774f41107ab59ffa31d564ae
ze687e97da9f53786f11dc60b9159987120ca71afda4e1738bb0e567f4419f5743df00955c30eee
zd5555b5b99cbd8d733143e778a2816355e5b9cb0033fa3506e7ae997d7895b14e84d094cc86742
zb49bba4bed1b369e49b8cbd0fe19dd9aa97136de5d85eec2cfc77764f3e6e7116a8b76aef3ee62
z5354039a9abae010a2ec8fef52857f5b188a1e0713a0bb15a8d5327d0a12f357c4f0c8b7d6d93d
z27bba98ec7268b214285f2d51738af25f1b354fa772d51ae2c5bf9a42bd03f5e75b5b08dfa2fc4
zcd92b894b0b41ab2f496a955e11f9e223a2b24abf1f1b99351486663bb6c660cad7a7548b2fba2
z0dbf20ff41a8dc1e27e134e57228165b88a22c5f94e127264b94ee73e03ec895e92ba43f2c0b9c
zb59be3be807f9c28c603f913a3267004528802faa00b3a236afe6ccbe1da4fb4f93fd10fa67ed4
z479c91d46e62e8cc461e1da7f63120f570d9f385293790050d793e3c245b0386a43fdddb170671
z0a6e3062e78ed1dc5f61a9007ec53eea0d9496494e7b7dc434b47b7d5de1d7562b1604dcee4276
ze47e26fc5513a4e55fdff9df0b349be8e41828b8c194d14191d728dd5ded6c82c49969cbe7c651
z7d2614f08c68d7676ddc1bd8dece87c2e71a402397ea888481483a4e20a3b9cbb04910bc4e0532
z076c648670205df30a574db5a8db31167796bcd069cd003699751bb0cacd0a056e04723ee6681b
z7b92a555a7fd6e3648037a6e622ee2162071c4b680bea7abb672c81f113e8e5cb1cd6f4358eaa3
zd6ab6f51828ccf72fa273fdf1716aacf6ea59592c9a072e2495aaf83b5217d19df5854b10d6d4d
z3cdaf5a19d6970e3eaed0d7eb7a07d2bfdd09d7ff010ec7c4cbbcadb54e9ac3b4da7f29d9bfbf8
za99b9857c9e8d4433174e2da20770f45daa9e5c94f50f77415ce1a67930a3017993adf9f3e8324
z8bd7a2724200f367de772849d545fe285eb05f8955cfd46d95e2cfdbd1a76a2abe37583732b8d2
z7b75d8ca0f45ae0041c25903491c13e7274c14fe5e3131b16268b994db3574af7f979b75a2e2cd
z3385fdbc71e57e77c49facf6f0723460edae2ea5c940e3a432642995441c2083c0cc56f5f10450
zea55a132c0a1b174fe8aa2fbc0ba14a57118338d1445b04402be848a2e76d8bef576c64033efdc
z119b39021f1307981cc030e835d6562bd20ff1458717a0011e39d5ace341fc5a6859c469778cb7
z88058112b1ee7f38e44abaeb471c292b6df97a8e99a774f1b03497791cd2f1b47e7053a971b28c
zb992cea0b9c0a227535dcae2553871984c5c275220a0d0ec9c31880a665f160a6c037ca2163fd8
z61c95d5808510e06e9975ebc99f62affa8c9249d02f03ff41535ee54bdc449ca9d0fed632662c8
zbdcab8be4cccd2c65069852475313b90dd5be0449dc0b7bc44d87de75784c8e3f7c2093fc86245
z2f29c91ef06ee472afb4f096cca0033e12d6f1c70ad506ed6f34addae4c9c21cda9825acd8df20
z8b6c6044530152af330c624f3fff7180628f20a15a2825d366be12d22a3cce2d55b16a76ec0474
z476967ecbae682672b9ada00e39009e62663db7081f0c2e693f5d8f9c1545b55e129bd6120b9ca
zc36377a4ffb9483e5a92ab04e160edae62c8b66d1b891913a5b613f3a02f70e2a5f6e13929c278
z1a2599a99474ee59ec8d86eb92889b195aa6eb6be3ec465f01cc197ea9e290d20665446a6db36d
z4c7456fdec6d760249e63ad92bc74d726ac1de10fee0c13ac272f0ab6d50244944b65931da5bfd
z35763925f0cd2723f4447d0cd0d84e3510fd99359e6622f39b944f27591322176fe0e4324d3d8d
z46cadeedd092fdf77f056ca40d76b70266a58e0f02dfd39a62b4aed0db1b4bcfb337df6bfd8841
z48befeec0c4ed841f132014245a2d8d7266013e144a059763baeeb1ae17a2db11de1ad1911c89a
z7d9c66688c8a384a3bcbb75eac890efe2e1ed6cbc207766fc2ac75cce8cb5609ed8971ddba6883
za20ded0c4962295e18c2bd20f6121a8920fe82bfe50b002a51ef0acc35b70e74408a63d104e1ed
z802fc42c9170d47a8b22717c565f6f10f9fbf47a43f0c945a2242f3b5328fc47728de80de040ae
z1530e4f674eec746a12a79fbf0664720fec408651488616e8d308a1e872b4128d0405c32ef2919
z1a27d22c0c0dde03d995fe374c13b17b3d76b1109359f137aa01886179434e0754a62ea205b534
zd173dfa01004d9f466528d2e6586d674d44c391de8bb2a86dcc50251cc028287d14e12a69ac2a3
zf1c1fd3ef849c81a13a15053b5888592f18d3ec6e03596b9de65357c92dee00f842d749a27adb3
zac68d26ffa6b6cd403182d8d605c843f44e11880fdd8654e9967d65c1b27b651777c0fcc1714bf
z84ee0454dd2b8647d775cc9cc32d1e5631b692c74a9d321cfa56f8aa039d3f472fc8fb6aa0667b
z35e88f9dca79b7af8caf6e18bc1f3f3b91c3803fccac463c4f00a0441a8a8825ee552636d982d0
z1cbe8cdd03ea735dc458ac469857f2f9b2914bf3e27e0c59b8ba28959b138f2196c8d189534a6f
z72c8ac6eddbed2be9ba6a7e9d769fd33a46efb4798b608a5f1b10b933326f90e1748aa0aab6f9b
z280e2739c6316699acd25629fe09998978d433329ebda6a4f99455cc7dd0ee81ce59c8125d36f2
z78838089ed0684651a1be8c36e418e753b0d3112bd3d761cc7d59b9118724c2398b45c5d724eae
z122132f6c179f95c13ff825ea525c6c759984bb3a1c4987dce70bb9b06503871e4393b299024cf
z21c7931f2f872492a27b8b06081105c16a869ff7d01e5b96714efa08d6788a9a42b5d69c7daf82
z09704acd0002bd128c4fd52f57b676f8605673d157c9083a4d9c4ad6a4c9afb7571229419f521a
zf277c1fd2f2950737a2e3750090482d589a1e69bd67d00cfe3401e1667c4655e9f5b8ede3633ce
zfa82eb7fb74852ac883c8087623564c32a124bd8aa0b13a0b74eb05e5e4b5c2c62beb09d81f574
z0a5cb6edc666d28b7bdc6f38a5aff91f8292655cf1a4593a2022ef48ece60639d640dcb2434c1c
z5ca8523c870dd87d83b7439fb9b54f10e07953e739dc4cf6c6e498791877615a27b8cc7e7cf9ef
za6d8c82d7230f9f3178e5e5632f86bdd43f487eab0449bd45fc0db6b9f603180fc757723de1ee8
z38330c192b80683b8a3099794df345fba0e9b728102bbbfe35c2e8a7e8dd66c14054a738ab967e
z5adfcbdd98cd4205e2060024c4e6b8bd59fa081a6e4222cb9f663df0c4f082b6abef683a47b52f
zc71e6f4ad971f304c6f2f7fd326fafe14954ccf591e7d010bd114473878820094f9f9d5a1098f3
z0a24f7f0dec457488d457c190a466569b002dc8eb8c68a254817a609e33d118612efe9ecb38986
z9c303ef94d73f4d2a4faedb6496915da7e7064ac5c6dfc1ea5bae2b5a8109d7f0378242deb45f8
z1327b53f7b9b70011ee9f33b25fb2196d1a3c2916f45b3094aba2fcb6bb3aa5799106e24371f2d
ze6b56eee0e6b6c2d424ec8aae99b13a27f7ba64dc83f752a9edfd76a910d095144a9b1c4ab4978
zbf38dcfc64dc47a5b746fc63c264e0a5c15ac52962a0b3931971e574caba374a59f256f86e48b7
z0ce6fd80ec7bfc0ba8632bef68c0cb1bb66e2469f1a4299a999cdcb2ad0875ec5128b30ae5e30c
zf6608354b89efc1418507e08b8dcecfd18c994542e5a739194d5238b1805ec60690d5ab859588d
zc15440d08cb8ef93f2f5885cdcc3b5efc290ee94bdbe413e4e7c5322e3c890bac96cefb1af8ca4
z0d2fb2e5f388c01d796dfc6c4206353f215129bd63aab40fe318d74874fe0d1537b023ef772021
z1ef0d5856142f3440583cbbaf6b50ed72da73a7dc8abed58526b075bd488e82d215e07048c1241
z39249469f7d1b60f07c7fa0fd9b01eff7b007442c3106824f5b09371c55712673f984ccb75c311
z5159364d862aa1ba207f0a11d84d51bfdc7c7baec6da2df51b1d7bb63ef7b0a533e2ea5f4af8b4
z5ec893c89f293f0f522e34fed28a4e2abd982b910303fc120b433000528f5915eca8f641735849
z323f9360a1a41844c27f2b624ecd5bc547cf3087222b64f498988b20c7778c64a0d5d8456840dd
zb67474affb12408ea5c4cf3731088bd840fe93407837f323eeed6c10b2fef20347b0ef19186544
ze6639e285584e838b61a66d1ff9920498a3e7aa7a7172e801ad27cce141469be2f2394eb8547da
z086c1039bae5a96b333d312e26d71a85434cad0034c8e96545bfbf35bcd2838a1c8c5cd524ed28
z68b92e367eea52055be4b9c5189f99ddd4d05ba52eae3615256c8fd14363bc1a01e717141dac39
zeb205913e4e8f18b3fbdfefdf77516985818dafe1d93451b0abeb2ce07e3d9374dc92e1abae6d6
zb2252a56b1f38b8699dd9f2531043289f2260233a014f2d64fc177f6a52204b487dee9bab98565
zed7e3d21c6703f58eb4b402c2d87cce32f21bccc1958678c58aa4a4532b33e82e0f40c011df6c0
zbb4a253014fed1117a7d05242c5dd2fc2dc75943e73f0137b199741b31c19d84e0a0eed4930ff7
z2494b7ec5e10e4260bfc48cd538223179d86a8808ad0ebcd8ecdc43793d311e85bcbd1f188f924
z676ed633e43299f8b0fc31732ed6b08cea4d86e1316a46336eadb0cdcd4734613e0c7a44c00e95
z1ce31116a5616150196e91c251d0bf172c4a38d5f6a1ae0a41cf5108d27ad4668a3b7de3716ce4
z92c941a5e5f111fe33dc3725e444d73d7bfe78a100148594c422c1d068445b521dde31324882ba
zdd41fa11c2f5dbccd21b3439553e5802db763980ac3837146e26295913d40b5bd09ea3e7887a1d
zfcab5a42d0c69f910b1dc57db82db29a006acfbd86151337f11d0cf8dc39b8932ac7674bfc80bb
z5f5c510478a6a344d5a2a516167dd0cdb3cc31749b22cf9e35056b2a58e2cde108671d62baaed3
zb06a529f2363345332213b21bfa5a1d1e2ee482260c5b130602421b0780e25f4d4455129f09c23
z6ec551a96ee5cbf62b8243cb8505e6e5eb7de9c37d25c860339d2f486bf6c70c36b59cfeed965b
z70800ca39befff9d4ca66675f9c732cbbf11978f61041c306fb94a92ae66cbe570d3c58270b577
zb7be341344446add80577baad298ff9d909c691a7c71be6a95754d12ab2f11e63701ebed9ce66b
z63fb8d37cbdb2dad936ba1af4d584d9302359a2646f4ca9e36e3f64bd77730830c3973b39bb6fc
z196f271c7825096c306cfe8df6f20e42a9a259fa1947fedfb9282362d8598e362d11ac4db7d4ee
z80ed4af354eb63dd00257b50fc465b07498cbe4ffffc3edecf474280a89eb6ed5f37855014570b
z6b364a20d18d9a58c65641920d7e8e25f8145178d818fbd6eebf1726785ce40f3368c9bfdd0992
zcc1f219716ba6f7e19db54afe74f5df640c3f4efcce9dc34ff49d6fc2672965d5f51d269c10bae
z0610bf1b1e3ecc8c0ad4ac84ae877889d72ed4e49b918e0a7760f7b7fed9d3adb0405f27bc0b5f
z2eb5bfda787946319da6c50bb4554f1d107fb9e95024e67f1d11e9e6c224816446d03e0b960915
z2e3fb389c8a1be1de3f11200cc79462787b54faca7c35dffb9d12e156f60aa44feddc641b2e998
z097a1f9cfbf6784bf66eef0c28b9681cb6fdc62a28ed50b7759b2a3f9bca2460ff1e1d6cb2f869
z05a15a4b8902c89a01441d10d3c662b6be7bd4a290dae181771fefdd1a3a68e23bab43c0dcaa4e
zabac1f0d098992c4f803854e20767593f4f194954dc308ff0774a4661d26d204bfeecfa7292972
z783300b29c34a9b529ec3a8b691a820a8e00af122c753995647da51cb61d51fe3b5187e0f937d3
z405daedf75ead9273d2dc75d4e4b9d50481e94d072a346cceb867443a2bf9c9bb27eb109533e65
zae7813b9a8a9e157dc365e5676ba8a9fc2349854d6cfc8345bbd60baa9e10b9f562dfe51f2329d
z03ec0bf4ca1c3cd5f5d13eedefa106bbbfbb6b698cdda4a25e0644683f85d4ae83133596b71c1e
za77d8ce852bda678bee566b6d4ead83b25a4fa84ce22716f7baa1c0ad742329736c87452757287
z1a30ad0f1a39097ff58893181da5653f9045b3a1135b37875be822c99138fa63946c382cc16b1c
z74eed8175751edbe9688aeefbac860f5d46a0e5ef4b23044dbe0656b5741b481efa6eecaae1158
z7e46598c2a93fc5828dbd9cb36e54b31c662daeaededea44907c31968abba2e1400f4b224b3268
z2cf7740bf6bee6de335e8a4ed478df827dc1c43b28c003a9320f47a61020b17a940325d9b2bb6a
z8d5e4a816c292039ee6dee9bd4763314463b3b546771f3f34ad5c9a4d79cad486ee6f1c8cfc99a
z67fd3cf4d7975bdb91683c39ba2d3bf5f9f1664561cd4c2507516614fecf078d498c200eba3576
zaed6ed289e8630cfe82435747e5cc67318fb0bcb80b7317d9c0b7f3b549d4b9aad724b6d8afc34
zcaf302ea16cd7282ba646b3bd3c2c63e491aade876c79d74b2ed1afec35c36d46f7f640643c91a
za88adb922fe8ed9d3afaf5881f80090302cca33ebba0a02f01f388048b3c6ac155c5712a0ba291
z717ca261b3d71184b65c5ec2f3892027f2cae5bd09bab49dc97342250dcca9752a52e5230d0404
z721c2c28d1cda2b9008e8179cbb86e2064aa63a3d411a2d4635a3ac4391a6169bfc1e0d4bddbaa
ze13d2e7b576e2c3beb4414585b61fd24083d329aaa3ea8df7aa57d853af2226a2ac0390fb5f9d8
z753f8030bf0cc4de8a768f874fc12717519c910c711c217041559435f47f07f4dde6ea4e06b80a
ze58ca304f695008aab586b72f7f222e7ad8763772baee0b0b3712b939cee00d2643b0764df7af9
ze883e8e627add10e33d541b9ad625825a351e22d9db57be5f5f64d872aac704bf7061ff5b4141c
zd648de03d8062b89dd4abfe095cc7d2cbdb9d74cf83522521bbf446a293e02811add77680027ef
zbc6bee8b51f0e7d00f262c8aeae1ddbe647bf2450f7b0f19e62a401d4d39c3a1a07f15daf2302c
z271ad92a89df7870496e349bc57452f9f9bf8f6a3442eb35aed72a9b7553f66187cc9e539d54ee
z06df46dfe4bb1ecaeae3c8f8ea20d7baa2c85cb21c19e5be0fe01192a37b0f42a348c8b0e2d125
z12df2e59f8fb16d9496fe973dd24c0cf895c919a9914f430a4d67e46833b65e6f0400861cdd183
z4a6eca3dd94596b673fcc035a4578625fed9c07aeb6485f7692068d86c55fad67b66ede66c72fe
z5039f5f298d45732b12b96ecd547c96473c43b62349d065a0fe27185af1f842f4829d1f871d357
z7af3bc51f10f518fe8d0a4f8326ab79a55a188bf8a081e7e582fe4b336c49212305e3926f63450
z6510341cdd5735abc5f07b83dbf6985edfabcfd298c2d8c11cba4e4726831bd337a09060c375de
zf3ff0880f961bba6dfa16a12dc7c16ff4aa62090c57ffb44973ba9001e85337e0a7844e3188a2b
z70796da4afb76aa175b403981b6572c6188c4bf0a24d1589940360dfd15dd7ebf6d178c8599743
zd65e98299ba5b8acf3361f149aa459b38e93c264955ceb3c55f850159a4c932a2a8cda9cd861c9
z93663170e677f27aab69c38161994bdb99c3720711b0d814c8a225ceaa437c717293f13656586c
z3f2589a4b7fb59c78569372cd86b26e87aa57ace42ff905fa725e8b0cc6bd13efed18da11bdcbf
z05a8c49367f1133565d155c575533713be03d45f5bd295a7c9499fb9883030011086c5b20286bc
zfcdfed157de458387be56df49b474f0352cb5b532670ad46dc317ba4406d94d9856ee7d920f7ec
zae97be0c76c7757d29127a0200a753820ce872d7024977f70886b900e4d4332ad1d21b514566f1
zd3a3a19c761809d4b2f699991c6a543ed91588aca1cdcaace34e2b9745da32183d5cb50889ab85
z0bbd9005fc81718cc89e77964af1f245fb61d4846f50732613f6818d789aacfe4f1fb90feeca98
z2c4061acd22b9d20864dc36093321807e134d43c5604e2b306c678cf855a1802307c9b20772646
z23157a2b93e3e2a343bbdebff06d7903160538becee2be2639ced6d5da8977e91027095e96e1a9
zdcd1efd79a29ef1bc27b7bfb948473640b29e08650a2c8f8a07baed9b4092979c56bb086afa7d2
z8901955d4ef7626d59c574a8ccd8db608d04fda5d5824e2ba704ca5732c903dc560a467a0268f4
ze80646cf0e707308800a45c763b2db066960bfd2ce8fe6be84987e661c1cfea4414eb31c27e07b
z9d9872bb1b2312cce898e3d45ecaee4ece6a102a24ac4358bbfca4635ac9640d06af49291d734f
z6bbcb8c54ab2d05eace4e1d34a622a133521846cad1eb0beb37397448cfa05dd1911b02b99e802
z54049e1cb54c601e0d0b0a7c6dadf57a2d2a6ee47db9055734ac7bf602215acf9d8f97a53c11eb
z270951b96f6d8f01970cd07e8198fd7f40fbb3dac7df7438a59f8b87fe3a8fb90466bb3754b297
z358a6b84e2a84a0ae2c62601446a9a6bc5d82b35d783cb0ca49ca0a51027f9409538e1888cf12a
z2a5eff0e61c8cd76586523a6c91dfff9200936cd628cd2414892a99dbe4c38ef324e4268439e44
z6e24d7cb8609bb8c2679f1a63e87ba6f3ecec23f122cf24c092379baa6f0e90ec6cbef42163988
z27dc87996154c8c1ffab0d422d8558c9f34196f0e82dfbce4c07693b8a827a9ef79f23ee6249e8
z1a518f247468b97642fd7c465365bf5845e7ab59f76b5f2674c3a4d9627dc87a5ac27b746712ec
za1abf2d085367549509b14d3af1f31cd410b221a785e8f59176f19c42ca4a7f1ddea81e773c35f
z14b79f475948bba93993d1b70b786299b93249b8a9c929aa0b83936a4fa201acc58258b63bacac
z7a0f2263cce9b74236af0352b1342816b68a8454b65fe42f78e6d38169f4e861024e2c28f72b1e
z2c98fa6dcafe8cb36fc7bca067512135c04e2de9a97297257f12a86caa67d159df1a58f98b5a90
z3b2b1619ae9b90ecdbfe4c5dac872c5c945fdd80fb3c3f165f22d2ce0e1c1e89372cacba6a18b1
zc52760a2888cdd93628c6b7212b4ca51085f61a5e7d65b82e2897a5e7b21f77ef18df1d0f4c379
z0642f32aef30463a6c81a82e057b93bc844412fc8f2fe161ee0c340402b51a0b65e3178c428b6e
zdf5f39aa00f9e3b6ccccdc0bfdcb5af65ba299edf82caa6e0a71bedef1f38926351e175a60ad4f
zd3a701fcbc0cc2fe18be261720bfe580f90926a39bb9fbc45376a78f0f87cd0e5f1e6f29a87503
ze02426300503fff092f0619b058e7926070769dbf13ce3aa30633756e067cf9bf129fea89077b8
z4b1e696f3a04245d3eaf161aeda2893c9203954f1a05675b184d1d8cd8179626d2da1a87d52698
z9150b065ef768c7ff9ec61b1379c682f931459daeb3e2f9be2751807aa4ce4973ef38e8a8bd752
z8b3d4484f4b2021a072f05c8f016ba652ca29ca40ed6f79747ccf2b1ffea527e50534d9a95f8b9
z6203c304286da9db26428b755a71c6cfd22c42b1dd82d4fb257cf488d57fc6468c028729dcb31d
z0b28ff73d831bbd06a0c45a2b1fc5771dbdd9d437ee66ed250cac08c53a46b5382228902aef320
zecc027268385a5ba0b175b25623831a0674ccd7e4dfb1d1efe3f85b190f73d7c09603c11545d1e
z5006c44d03ed2531c4b84bb8c96724e836e58c2fd1b6e6ff3194a7d813b0c05d3d364559dbe1c3
z09bc74b5e6f128d3ce5e2dc37875af1e1ac79c2152595f4744419ded567812d040dc9096607ba0
zb6d72ec4d18eebc03ffe07a8d2b859a5e19208f53213e2cdba7d325c64a57f12707ceb52b800d3
zdf03e28c8f0eb345881fbd17132ba24078805187752d15d2373bdb3c9130948e378c889db56090
zf13783cfefc2f48521a0aebaf762cce3574c62ce2132b7a6b94bcc15ae96b25aa26a7ce4df5c77
z503078cedb86072f1afc2704eab968867e5e9ba8a56ecce02287eb21b3db6ba0352c14efc7ccd5
zb4e65604d2577da177e8c21048d73f2460d2b97b4b9e5d95bacdcadcf3e1663123ce417e880bea
z942b8bf9984881c6cb8c96e2903a600a3c0c72eee2e616ca58f657123e7100f03094b776d9c7e4
z18cb6f9cd54a377baf27d9b6bd6036459c96f30a12f1f94eb17524c11699de85e62663258abed7
z0bfe95f78be2eb085005af25815765429a5546a324860a371dd927238bd795575045c6539c5b6b
z1e2f7f19de1384dbfbb390d15e1e8e51cea4f33791ff93cb5b53b260cb187dee173ad684d87644
zb361054e67df2382b3b222cbb1f98b94adf0eb41384f618709ea6b239f00efeaca0ee74354da4f
zb1c070a5cc9274c5f9feb2c743da7ab788b1ca10324b8153d5900782430607433451bc9e7e8331
z5552fe05734fa98e423cc43bcfb38d3ee626447124a7c60c953b9c21e44b2835106110d2333929
z1229932d35bd09e52cecb6c8d7c3d6ab361a15243501a99b4b2b8a8c37c8b8a68ce3dff8c4a16f
z98f1d8356c65961558f36561be5c78322952ce4e4f9b0147cb51d6d39c4f1deed170d5ac82ec77
z381fd6fd2fe684d0678e9b66e8765c9b581f5e773ea7bc7f27ee9eb89328a4edcbdb705e602067
z7755d9d0dab1cb9b3a9497f84cb04fa3c98fbb970aa28770d5baf138add41233e92e3a5c41fa5c
zebada58d35422b421f38075691732824327c792791c8f0e1724a778c3968cf005c99bb5a220090
zf36001ae5340d20c4d420aea469bf62f7d8425bf749cf7c98b3cdd8f681fedf7b12a1ccb965d85
zb8e4d32c6245958465e506ece5cb0680ea698ba02fabd5d6a577a9c31bf3d7c254b9ca37530c6d
zce97afc9ae78b6c9362c7718ab8266c279b4488a2e88e6199ac3c3f573e8bea5f7249ae744d5f8
z75e52f231467f28d617d9927246804333c8e3c8975965a2ec4e7ec0dbd9edd5d44a13904d94499
z1cae20dc81c585b014139a88f034448d09a8c5da9bf76df0e8677d0260f4737943b351b36ef2e6
ze0ebd8310f768f7db6edcc3f516dd30395cde8e51b45dffa47245723d415491c9347908f5ac08e
z0d1327f90cd2dc0684650d06f347429d1e52ae18ef54ef401c19ac3f63cec338c9876ab8090fda
zdcb637cd1995a51b887a529f88c53b62b881ddcc1ecb15b1c7294cf8a9939725574a8dc0c167ab
z14dd24913f7187c0aae0b234a5c41d0daf5ecdae268cb8501a2d9f0b6f131c5f791ce21c27c423
z2a5da1fda013f1ffe8b2a0fa5b54b70936e10aeb7e908a56aebcddbde40a2b5d6da389d9ada0c8
zd0ab300b4413ef86cb7d999e71355695ef8ec91f0e1bf643649f17e132cf6b366294c3b9722552
z2954d869cf35e14f6e42e6c5a156ec326e16bf58a3b00439a25cc152a410dd36dc7320e7a095de
ze41072d9f666edc3afefc43912e05ae2293c0f2f2f21fda236f5e8550ddf9f6c0e27d8b8f6ce42
z5643f2a23f876c42d18e5f95400f40a6223977ab6adfc79cb7bb6b9e46c68dded34dec11681234
z22aa9da9b84b9709c4db583a9e1b551dedf24d70c291ec8bf7381013c0f425b48073fcfe8c8c8b
z09ab64f6774b125be6a408c227299578d2111be51edd42f73f8704da1315589d2e7ba47e58f5de
z3d956350c05679ae197c6f399f4e7fab2fa2fd6666e236551db202e032c6e5d35e1809ceec8ed5
z3bda1a1978bea476641cb7a49d01d915dccf8dd842528c67ee97c8146ed4383cd914aff003d2a1
ze0a68e6565d834d32ffb3326bf04be63fbc527ca0f66680268564ffcc1b0ee745a17325e4c9ed2
ze6fc857e7b2a0f412a8fbd465c0cf3b7825d46b9b4d5d7f852774553d4bc0f0b5aac76fd4bb5e9
z089b7895121a52c2165b694695cbb96f1620c1a1ba9e2227696dee95a5de88940dd35211610c4b
zdfd5477280d7dbb0b81fdefaf0ffd7cd6cd013de7bd691768cf66d8a098009ee5f036c6ff25bdc
zfbf60dd0ea086df66cf487cd352ef515dd0acab168fc05f7e77be9931ac9eca8b7ab26c5dc330a
z19eb1e4251ef02b489990d56fbb910277bea409599c14f51cf69da0c9324c510aacd63779b1111
z3119dd7eaafd1f8631e546c452326301469428459d5d147673f2a5dec459a947068020f907a2aa
ze6ffc31b486167a72bd2f8d9250dd0d971047b71913bf656235405f5d1c21d9a7f8d4936aac7f6
z58f51f96fa43f28c78dcc3141faebf498630dcb0e7761384dd48c921a4f8fa6c1dff957d406c07
z5a89f053b0f0b2f1f53b25f1882b658afc0ef0e75e8bc2d9352660f73ca136602e36232bd97b7f
z67f861f7f1ec48b236739e1bc72c3046105720a690158249d0335ef47433f58ca76d162a761597
z9d791afe937af59342cb9430d61254457a8a2a07a9550f110e7daf89d24f3af10457f50d8ff14b
ze8f4f138d63ff83fd4717f4596c14895a2dbf4c54cdea1f361d10b4aafedc5eddf921c8d7170fc
za6a8d586d9cc3130b09ec998da25f4708b7c98af39e5e165ecd576d6884dc00ba8f775df837365
z393f1c9fc2a9fa76c7074229de7daa6562f19d3ec94d8c861083dd0b14f85c8e3a31b734e6df2c
z846f0c8147d6dce0ea9cce20de51c8a1ad5e55f87b113c0dfaca00d2874ba53f81665ebb5ffbdc
z5f608245d9c8feac8a95ee4969a486aad16f1c5ad00ab82550d3d80114a0336d657365157d197a
z1301abd399d5720a0d8c4021bc6369261aa53d79b3d316b8d1664c66edaef58b930ce5960ddad3
ze687b157d7cad08cd6e90317282b146c55232b3ecb63cc59beb80394037082246b6a2ef6963c9a
z7634b06502ef5e4440a97a7121581e166ed6a4cd830ed086727ab5c2069437bdc74ee7f5be9584
z280ecc4f7d91efa5d5dcac3d9f1643cd1a32e1e58f0a637a96ef21dc1184012df0b90b6e7cf630
z39f211f458d26990a6904c966711cb619f655e1b9ef9b3f063ba083ad2a14cb59b2e5843034e61
z39b686413fa7b95e5dbdfb3be07a23d3f1309eef33a9eeecfbf73d5e1e9a4da9a83c81399a442a
z882199bade8a4afb4b7589233bfbc2096ba7a6765bda0ba38a5f14040ed1d0554163f5030636e5
zaac45f511ab42d2f7398b6df09c20b462af4a1e15ceefc6dad4fb9b75b5a5e7015bae5a12e8848
z128759a236b653a4a11aecdb48e19d1726d283a406903520dce74d76de61fb5e8b6d91b7e77c89
za6f64bc22c85e3ac45310787b4df7e9427cb34017d4d1eec50353978d1e39510e7d051e243a22e
zdefdf5a49672db869ac4b35494ffcccf0e2e619ffecfb57793a34fa904982d5d57f60a0a35d18a
zd4c0aaa6d94235bc2c707e2736a8118299ba6e58af15c2066230a203c0df7b2b4c3d4df2aa1876
z41ef3544e6aea7c8f3c3d4b53c31ae5b787c881bee1537db4ead8b5a355f184d908973500dc457
zbac9814904bb2662cba0e8cfc5a5f657d0d91e1f7a28c97925984b13e23a18e74dba5d224f6b2a
z21b112eb1a043f6c3d44f82fae16ffbf0af628e955eebbc4db04e62223a37a1cbeaf6eaab3d0df
ze73c442aeab5c22d95e6c59c9b31b9fc36b8396a1dde8e060aa5f1d26a36eac3b2ca722112c305
z921cfd224f563643659d81908878c7ff17c56baa4527ab4e9a2aebf8036d83f654db3fe4a91ede
ze473b90c8b246dccdc949076a804059490f9aee763c8bb211f284b63ceaafaac9603ca9fb18f77
z3930f7dacdb64c2aa41dc422903b81a4e55b4a4b059bb8ebe1e53c138bf5942030866617268e4a
z0887e4ab71063cc2a3c8ef73c23eb3f76e0bb12e106849d98e00bf514954a74678df4779d8c9de
z3844b88445540cc8f5821301a0966a769e891c73ef94382442585d4b46ebe38d6fef5c5ea5a83b
z43f350edd580b8355f1f0b6f5981e29949465c4eb487b71fbb8d6a406d90992094a2379999cb04
z206ad6efa0313b9849b963026dd98e334b5c180838c744cd075277e6ae309e3ffea3cacdd54d20
z7a11bb017bdfa97c6f70051a806aa79273e862c0b504d3c403c3039b846d5d8547931eb352eb67
z702a7c5b657a7e0bf0bf6a6d46429b0d19bd01c8b0a46da4cf1c332fef3379f5a1b7edb3cbc811
z4d28f025145b72a36066e86b89d4cf9df38658994c1b986f4abb2478f20f9eb51486d6f6bf0559
z96c3ca7fe0e6b59ed1951bc1fbc8dc42ee1a68812e8d786e47bbd7ae31c53175abe18500853e3d
zd898f832a2bba298bcc897125b4a7bbaed7c3faa5308af89601159d6b0a9ea06a74fe8d57c50f4
z5b50f4777b22228388b080f53f39f9b2d390ba507b4534dbb927ef29baa144d5a1c960902b9635
z238428c14facf4f5be197ffe41185f58a6c4251ae63c357450e32439383963d80daf731e266cbc
z00081eee7728ab0640ce035d1d3dd2a715955f1a0d87259249594ae3388ec42cbbd2d179e51732
z29ffa63bbaac2bce6e2cff1802986ed1184d4545ee70ea4beaea7b5e26c6e8234301e92d55d171
za3f5dd0e4eacdcb7a07132266ca9c0dbe90fff0822f53a36a194059db1ee591e17516b28e67641
z062a11b69fdc7cc55384bb6d9098a2a274578719dd5cf49877d7f21cb38cca4cec4decdda1561f
ze135e1ef43a68d80b21525b51956b15ccae965e4cb20cf375a118dcf5b1b99dfd6e4ac1d18fc70
zd6c8c6dd6f0167a0240afd4e4c248badfeb3c9bb1258ac39339bcb73478e5845078d130d5daf4a
z30db95515ccd884b1b17599beef776c57fc0c441a1b7e661fa08dbfa769e6f1c34fd3dbfce0aae
zd5b5c3583e1eb4efb4369b80e1f442166eb0b775a3c1f1e38876aaff2ef8258f3e4e7d36ccecc5
z0bb84995aabc16ef7976183c61014743d00159c6f4de04b09c8dbd24b09ca1cdb857c9aba8e87e
z01d05696b6447e4a1cae94c966ba7de671d0a03b8b8b7af827f892e74b984a184cac5a88881188
zc31be974a6dc0f24e27999bdfa6e7936f2ef7d561a117dfa1c0e93c254cc03a9ff613c8a804a47
z8eb3c551ffbd27dba8ee8d8f93b326d7d663efb426c7df2e5eab523839c9aed1d113ba3bfcf98d
z74a309cc50849ada0bc0ff0273933635097dad3590900284e8601288179563f25ed0093da53c2e
zcdd430eeb96ce3a2a07d17ce6c88f29689715357f0ba17c97bdbbd693b3079a326b4ec88fd46c3
z4e6184b3b9aaba88f69a8b7cc3f2ae10c75fcf929b6d4f156b4bbb2d393c5f5edced9008fcff3c
z308f9554dc38b812394e92a75579b0b55fe772e9a5b77ad0e29c257d6982ab103a81282a32cf0e
z600fcb6b23e1df247ff898bf3caee2cd67062276b4f2b46ffe8c35fa4e9f3844ef1eccc74c1a30
z8846641faa2f720699b908e2a42bb2ea8e0381b22cc8071520969a3f7cda0d935694d42b1f8a79
z43e0da591732c38f8e27acf29582de0bce8798aabbb81561525d140501df1c3ecd10672e6e93dc
z6d256fc946ed8cce10e1fd306ef67c10d761256137f7c27d65c1d36609e4607c3c44b845e5f540
z79233555e5c1b72d0c4e3e33bd6aba3d8664195852386cce1893ac9b6b6542f084aa10b5a457a1
z83d6d8babee40bc931dff8c4639aeac9f56260d6014c51b6ea0a0e9bd5d4198ab898d821457cca
zffb1b7c6c49dc1fd514fee8019611a05616ec9a2315f9139c9a5191651a99d508659ea0b9a7073
z8d6317a31464cdec57f013cf5b1ade4ff18ba231753467b341390764ac7c01918716dd5a10790b
zceb37ae94c7d690c525447f81fe210c8ddb5f97ac031a82510887cb752b7506a5534df941a32be
zcf9cac991435c12f64465daa97812a9bf87f441bbdf021152f157fd49927b6d48e76d32155795f
zf3101ef9ea176c3bf47c01f9e79ed3bd630cff980f206d2f46434a2bbc6ca108164e6a9ceb906b
zdae2360f0d2e7aeb88adb573f33bd4a8d51f0212e91654b3787514af3b33573304c464946a5fc6
zbf996aae5150e59d72fcdfe9852a2c47565c1dc2449ea141639544d1b6e8e53d5432efa0e2e7f3
z9ae2a4371711459d221dab57465d6cd500b4ced4fd6f6df938c3cee8b0fa17d34830280c4c9cb8
z802837cf8c82346d0d2fc02bbad1ae419f9b5d1078cf727c967d050876c38c7c815d123f8a8c76
z5bf3808cb7c87b1cd47292274c3563f83f248964ca3e3d3118fb7f8a86a37b522289ab92e65438
z66a63854f1d5184bb3334ffa910995484a7178fe3e9ed9d59031d5ce9fefd8f7d7c2279e9bc249
zcd6a9619d93b6390e0e4a71dc47bfd5ebae37dc27c83caa2042fc0bedf2ccc772f240419cb601b
z1ca846ab7df083f143da6626f78a9e8f2a0327df69ddc54c48c5910a39ba5a6b449a7b4f4ddcee
z0d55f32bfb9f09fa26488acc8b67eff30d458b0dbb68e36a3aedaabae1215aa291fb78890f6079
z26b584a0b05e9ae727c49c51ee5ad51ff02453b4e7a68b01435b3fe1a6ac07e00a1d5fdc1e4ba9
z2354a5ddd491820744c7c469631f915d8672ca1ae2812ad1e85cfb0aabcd1d37e9cf8ae04a0bdb
z8e0bfba66fd1b006f5f636b20a4cd79318c2a22a053965787cf19b76ab147a0a7766b57719867e
zee70b0d40708c7a2e796a8d671f641a064902f38f44c34f96edd1c3b3b388c1cbb0853cd0b1e67
z9c736a4d6bd7d9ba9d625ffd8e207bdf9410d093f7e65a8be04d792175904ed16f29797bffd5ae
z42cf1813aa7009c7cbe0d553364979849941eb49bfc15efa1e8d05ff7d2539cebd7d8d4b28486a
z49406c78b40dd560a6b81900f99b2144e4b975fad0128548eb0cb9313fcb3bef3bb47f9db922de
zc63beff2f439355843ffe565d3495cd63ff74ce8cdab14757f1df0e8edd88d7e986450d0618e46
z55ed7e17e3658406ce08b54fa433722e81f9978edc3670e35af9139db056eca58f87eada2f5151
z2d90da53e54917ab29d73818b12979ad66589651f2df70087c525a417c89a6ec17ba257b48e476
z651366b1f0889c74c074cecf3dcda82876b63f92562832a6340f7c09b93df2803ef245575c8d2a
z4691d1ab7fbefedd14477a6e994640ba4ed95e3fed0c33871de433ee03eef8f763fb9c22f76ffd
z14a4c1f57489fbc8a4a6b89a915324eb8a00ebec1d298974a8f39c6242bd835a14ce1e242e866d
zf2b6509d8322ce55398247df4cccc8218f8d4ec1cda662763cb680691d9db613b7ce7b550698fd
z09826b4976a13a07f54b932c745a073207a2c509fd08c4418f17d850732044eaa45c7f0ab1c219
z046ad642d578da91faeca6637d57cd607dd9528e01d58692c812a600f4defa8dd4af22321bc066
z6f8ea825a07ebb354fb3022abfbf99e4b38f108b14545cf3003ed8e5541da567b423169f9b50ce
z7cd732afa67c1dcd5cfb51aad24dac0820cb89887d4a145bb89d9186f684a1ef9d4fb15dc84467
zaab07216a3fb674bd5673faa3e71d191545ed1e29635cb9bf5b19692d611dbd6438d81e8cd357f
z96b4fde6cafe8304c7adbcff3439b7de4320843b9470197c32c5f44dfb1a846583c52a829dc85a
zacd626feb2bf5240b146204a60c1d7c33c0e1bd544436839d8427e3a2f60850e35775eb9835550
zfd46d99f97a5012f7ba9afb5851797989c5458ee3f8056f4d8d97584a38ee4037178a1943fd5f1
ze11a390fd53943a66842013d64d60eb064821111b3518e1ea88c918cb16ed716e4c677b3695375
z6d29ea29a81359794822641965fb4c0fb01b30b5f9de56e0bff485ccf11be2b3c2d2ae0267ebba
za1958eba8e240349a45ff293fbf217a11f9c8c9734fd623fade60754f451881ee41da2cfeb3cf8
zdd8459ec04e4df075ca9a3e389c293768a922aeeec993b56c0146ced4107efe489c6adfc71a921
z42eba2270545aa4df6ca6134c3441aad2e6eaf23f6876d733f4e75db0609c3ff6673df142bf3b3
zb0f3f861180d43382c41101e32872b616ccfdf6a8f2fff5df4fc9a19942f08dc87e0bdb0114eba
ze21751eeeb14fdd35a651daad558ffc3744060f41df3ef2227301b47fb095aa80872eb0856d20b
z204030f019238d615364f9e43bb24e86cf8b14e0e7333addc572cfbc81acb1d577467a69aea4c8
zb523b2b854612216f013347d5624f8f2570d02e505bb5ff8e8d20bd45bf5a59413d2a67ef5310e
z0da89201295e01c6c005e4b50d52b686b26e7576f2292631bb082fde3ffa5d7f776f498f109dac
z1f8c6901f214d7fcd7922093fca5b4f6eeaf2af5e9015c805dc2581c82a9b45eb4c929a898758b
zaa23cbac6a978010bade513d7abee2cc548ab6bd05274e5f3580b72997183fc680830132d54e5f
z571cbdf60b9ed5d8d5a0d4f4a6efe66cfe5dd88ebf0707796a6b35e9f9601572baaf33c9609ca2
z6a9985fa153858c8f6c525912b75e38446a9cf19104b57c6723fbc223270965b2296ff0fe8f7d0
zee250458a9ea4550c6abc64b5d6829b52485a343664de3c25ffc44d1f3c99609debc80015a8707
z82e15fabc53057923579977396754c4d7f8e98a10354fd8dd0ebe6fed74dd1bdae85c8b6d7cba4
z9b5e878e53459406fd105e6b6040289802cb5068ae7d4490c84490242ec1e03540bba1712625e8
z790e636cede402d74505cdb8c0355bf263e72882c2331c7c120f9f3db15a0b0d7bbc9f3c70d89f
ze0b90756b57980e841793fb129c56aa5120989aa4741f0af31cc318d09b4bce27f23f813825456
z887b9292b843d3a5e3115cb60c90e1eb3d32fa891b1f2a0b7df8d60748467afa0d41f643edb9b7
z99beee4e2aa1f3a8c9ebfbc66ec55c24690e006c4a8bcf1cefe0dc7ea050c49dddb99a881ddea6
z4aeaf23bbc5dea6dd98cba1f304ad4c3081d4c8b8ee0372b5be959fe3ecc1901d54a2cde849c37
zc1c968425d97d84824c675ab4fb7e689699b2daef3763c86efdc72b21ebfefc4f2fa4f581b9835
zcbebff9ffab8ec2a2f34b9c9a141f6e02bde934288444fca4116fbe5d084e3415e92c5f0a18a06
z330810aa27f409dea76ecbb080a638792ea1c6c49f38ee4b872cdbe74d0a9e027cfea1398722fc
zef843092afd51785a69d7de7877546ba3a0bc88e99213ce8e98c76d23d74fe93cb630398bdc568
zad8a17725a1193f31e5e050bb924de783b46f1617ce93e3e9068bc4a8c69242bcbc0a0461b1a35
z530ff5ddfd4bffc64d9c64bddd35eaab809c077c45817deec6997634df5cb4ff9330be65f84f5b
zd33b3a739766eb3a9c7fae7d20c8e99b5316649b6481492176f434a865e88f30797b05c2913d32
z4bb3b13080bcb6177f8e20837aadacf180727cb19cf873e3164c595803e57a085cec5102ead01f
zb63211ec3a4842ed0d78ab48230351aca1313167ada95b4cb31a725fa478c330e4a10f520a102e
z249d9e8c3ffca6196894c84187d5c952b8ef016ecf09338a0f8c980276cf75a32a031a803f9402
z9e60735ab93bb9b7c1aa114f1061496ed57966b8a0766d2484f524320d94e2cab49e8e8bffc28c
zfd2dfa06823dffc10653b870fa96b2db2750cc51c07ab63d51b7de6818ba0c0480d972bbb9c2f0
z88f83abf416c03a420ff735d21a3763e79e793651b41e500f498beb890dde88fe9ccc7fec64ac6
z9cbcb3fd04833698e75a172201b879f404e56e60cb4479e8a9e6ed2587353bead622793cccb7ed
ze9701822418f3495082e9d600f118dfeea554a765a2426815711f399f94131a9b59d96baca285a
z14f381c902d40cc105448549547964aa772a6eff6ffca6f4e37c98fdd2ec2ace2358b8bccf52bf
ze5014db0b139c2b229b195fc9b2d5726247323beaf05718eaaa91930a33d2445e4e119af96ad86
za83c093f43c25c7eb97dbf3b076ac184362baef47634dcfc054cbe8a4d74374c0ec627d6993773
z8e4be79ae870e0bfa44e8e79be290df8e895b1f77c25dbc6509fede5c91153d20833506bab3f2b
z677de0180002c561cfd29d785c9b01cb193707702402dc1f0d06ebf07107e4ba914ee415739c7d
z4b4074a8a1ae5f330ca67314ce1425bb7201601c2a695d5ebab8893097ed7b2f7c55a75290061b
z549c0107636511e466930d7cc86bf15e42eaf92e5084203d22327931d7d16204fd5830cd5d989c
z6b83e4e8ca316a0aea45414234d14a7570fb4a98b46f59c3feb556ed1948f3841e5a03ea51913e
z2f58129a6610d9022c8e0b6d018075e86994ca4dfae74c521d7be9295f046d3248edbf9d5b7042
z5b3f30a6efd2ec8a1c65583124e7f9baca19cee525d3e25d0ff42b64c4a9ab7db76a9338ecab35
zb6fcf0be3dede1ebca4a9c22a0bd81a244d7bf8f41f3dff7445c5bacfc0e0f7cf8e509e98a8397
zbff76f14c3a7e1dddd8ffd5aedd629d96de33fd237c5ff64093ae96db43b367675135ffb679a60
z39432336f5bd2427afc1f6397b8964f761d879d65678297f1c8f40afbe1747c4bbb50fba5e1e5f
z0a3cdb19a7eef63a55addbbe4f216f4c77c930231fff5778725d231ce20d78bc2d6eb4622eaa26
z9a0318605ffcf0ec6f6528b15193f67112afa8f299bc539116247ba40464ba56cc4f44013e359b
zd136ce659537f0b3b0f3eba0a4712d591d2183dbb9e3d4d37442059b48415b68f3135dea3da913
z86db30c2ec332a859f27ed13cafc9cb944a959552c28c3a5e5972b6447e1822947a33cb4e40db6
z58af1409ec50085b78606c94d240a89c2dfcf3011fe3b9a5dfa69b823d6ea14ba03fdcfec9b38d
z13a8f7c2bcbdba6e6ba14258f25d25cb7426de20624f823434281524a85cfbf5243132aa179187
z3639826cbe723b0776982ebd8824bd03593ff939cd2041e4bfbc6c4081120ea48b7f89f973dc62
z70a8b63a6f66ac4619a27c08b9dd5e162f2243ee102b4f7bc80fe9c3b6fabf9f2fad6aae0886ea
z1f4fafe02959f153f817a870d3294c1b4fbd101d7fb2233bca0befc46ebe2c314b3b23d5d046fb
zffd4d9441d57b406853c580fba0938e0d73769709a988b33f5db33ceac6033b1a4f1a74e62fe8a
zc68c4eebcbd0e1d7bdd29d16f16bc46232db37b96796c2cc28d32e336f13fa6412dea342bffb77
zd94db8d2b6e3272ed44142d5f156abb5bdb851a115483171952e3fe1ec81d1175ba55cfebb428f
z798c4664f36ab3b3b0b0b80d54752379aa135054838c821002dc0769e97269cd67f0f25c5b773d
z6281bc42b497b2e6c12208253bd0f257537291a1497bec9f8f2eb5d1a931240278e8914a0574e4
ze0f71712b1764179efd118e9fac5f945941ce2850670a5fa49c5cb9b665a9e44c63d56c90de1cb
zdf5adedcd58051c15a797ae5685aeac97e34ff1755718e7a628a63883e138a439c652eedc32f7b
za6040a13bc0ee9795e647adf6b62df4b31ecdde3582f48306cb597b38e42c8b765925aafcd9fcb
z1c38ea4d7493851185b4d8f5c9637c972eeb5552e2278105b5896eafd5954fefe0ea70afeea02c
zcc71f10e7004eb206dbc41332ca9b218d5d016ca6524d20be4b4502887cc28e0c60272f9fe2724
zfac0aa4c2f416f8042d14af65fe1b0e520572ead610225c22960f497b1ddf2a3be0b84c66024ea
z392c4c0b58452787ec09eabab14253e33a388c795e407d9f052a8a11fe1714d02e2076e480e69f
zcc662fcb64d893b1b8e71f2019ce4cb3eec56b3667ee175af0c3d67ddbd6e898903e1816206bd0
z731bfa4acb95827aa526615ff1cc51c386b340fa682769168e21c4ce9bbb9fc9894e57c5be9782
zd77d986f3e4db6f96e2655353cfe20d5b29c1b8e69e1797901dfbb0e538a8f0db5f69c744d84e4
z3e83a205917fbd14c05660e19a36fc3b4526f46180fd60a713587c093efe19a80344e86660e1d2
z3eae0093bcb96f2534607681b93fe884606e8c288bc2c918f925cac0d037c2577259fab48b650a
z34532428476c073167ccc43bcfa03ca4782b3b263188aa6c9eb7568b38197e0d169deb4feadfd5
z5bfe801177b7faaa03c68cff359c3e01390f0a6d9b4bed4fab99d5673d6d812f6de95bba1914ae
z9ca01223e593600c690b20aef2a890cf91943b50ad13021c05491723842357c9f4940231681217
z73b1a2fb8992ffe297f753a43af467bc2c972e8feebb8b0831dac247cb83118ddade3a7e99ef75
z34b67046ba9d6beee51e75aa7e8add05f1db729edd31fae3b51d27a3930b5c1b5dd0bdd9746198
z4bc109ed999b181ad74565c30af2b33d8fd3ea535e6ad7cc9a2a0ff8ebef7e62980274a3380f61
zcbf26d1a8459a09d5ad5afcc6ac89cded639346a3ac638cf1de3e2849c2e9d022f2a119cfb841d
z883e69ad390f610c66e38e6c9942cae696b3d9fc89fe384f471c3ad2f4a937ace829054d28a2f8
zd01a74edf05ab101592ff71a5048c33cc6e02e28aaca36c0a6195973bc9f77e1a1b1f07b5dc978
za92b4fa2e584eec1ec9540da34a345169bb6d5641abd454fe750619739d21028b63c7a8a20b218
zc349a5fbbb309b8a1e020e5bb2850eaf9b6b1d47a74bc4d05336b1be0da1e45d52aa216878d2af
z58bf6d0de4ca8a05378e87123047363f306948dfac47f6ddcfb043b7769313104c3b3bca13bd31
z4be36a57b07ee477eb0352720c5fa8c6df8b96f454d1268534d6457fc4339f6157d78d0dd47209
z0eac10efa216a68183f91ea16638b3db6503d4e24dd8626cadac84319c861afbe72cb8f1e7f649
z1fe324739423bcc79759b3c0256df629965355d4b5259f332fa7ae7385f9e24214b29a3901ffc1
zda3500c9b708f2813efe78870724684b5a927bdaa2d9a418af8aafce56eec6a1c126543439c3ff
z271e2455c6ceb753bfc4d9d90d51be78a8f4dcaea9233cbeb59ffea936d47c29510c28bd02f92f
za536d6df64a5037b4680583b47322cd084d171e5c367487d675e3413b184a1068379c46ac7bea9
z6debfa1973720c7c5a78d574424dc38983b4437247da61d56ffbdc1cc2af881282d526cd03fa62
z376bb00c81ab4de93d6628427ae982aa75b2e18c66ceb54bd3462ba1f08af5f5bd687856996178
ze5c3dccaade418a49a5f127a489d2b1b1a6fdf4d8959a752a317b353d705a9050dc78a6503c5aa
z86f2fe34a35813cae5bec53586d6fba6c52d0150b317fa27da4fdcd9668e80f3143370bd71b297
zbb806846989151e06ee4e636a86ffd2da04658e490ddfe05a93e734b741548dff90cab71628077
zb4024b54a4f8f2d264ed4cb502f3fa4196f14a41f1f7e1d95b7759aa9866a2b514f3a5c898cc27
z0e67d689f8eaa222f1f834f3e94e4a936997edb76b75ab18ee187a8c494700d045e6a778185a3e
zcd104c865e2940e4a23e957658a0b5c35c3a1ceff1da4b14124a43264deb2ed22d2726c5392e62
z0104e5695b706302563f955405a4057cfa024a0fe969dc6983159ce451769e3bf6ec9e61f1edf8
za5a07621074afca4abff777b8810d843432426695c740a228b3399885e327583b9dec91dac491d
z486c4e8afc574c4813fbcf625e4209d1a8f4c07f8d45854ff12131f44b2a00a87ac1036b6e97c8
z7b305156ffb67b148110b48a2d2cee4601f1531dd39e9bdbfe7f231bb166adfd645667b6521a00
zf104bba18e39d7ca7c9e9af4cbc986acd67da39853731ae58f69abee9049bb7f8b8cc3d1744d0a
z75861eb87a4558af0b99edeb091af171e30d7a317db2a80339525f72fb2e883fd9a929fdea9a97
zbb44febf85875e06dfba2badd0b94f9f1dab65458fc0e2729da38ebd143e6fdbb8a7e430d51406
z5d68e91a678c776e25b20a5d07ccb2aaa1eb7038ee92785e08159bb1ffd6f677d777b95a3867e0
z75a7de94fca4038ff2215d4866d4e321f8fb092d3bffa9215a7c0e038920f77dd430e98818fbe3
z7a41e53e6c21db067ab3753093bef7511f2abe2c6ebb060cb5d431d01ac8a62b63e8b5bce8cdbd
za38bf664e18a076185ec247ad50398c90360e37f64d4dad0919932dce7a0c8421cb6c80f510148
z9df40bb8ce02866e017249adfe836af59ed7c3e3007be6f4d36ec702e82711fce9e44e2be1c729
z8fe9ef10e37481ceae9b3a1393bbfb61ae576675e79735b00db40f1f6f7eb289bf478ace06c5f7
zc5e61cfab1626e710260c30d8b2378a41ea456e896cb2d6b43ab9adefe247c7ce9ee9276e9bc59
z75f798388db44766cb0e1c075d0f765a482acd7943f80e2ab9d8e8fa3574d690b241b463934d22
zd353a9e866784b60b38540faecef448cc8091bf976b3ccba806600684a1308c29973b33c4cba1c
z223baaee971d30d94ebbfb87a4d5d09dba1c92aba030698ed3c31a7acea5ded2e8007e6b0910b9
zbf311469189a6e49e891704eb257289be81b0ab79fd5e09d43da198b3c419eb7accc9c219969f4
z1d150fbe50f94ef9f5c8c93b02168d64dc4fc10bed4dc6d86c5bdf9e2e4c3ea3cc2c193fc3d7fd
z863f23c6a4ab35811da2d5656767e5a2efbb2bcab529950c857ccab1f7c24cfc6e3016d5ca026c
z39b9c6373e4023a48e05d76eb6cfa9636d62a94d46a2d4a86fdd04252021193c1fcf18325be973
zdfe4b4d76d5b10b29ede98e38b74210433e1b4e0cd0ed1e15226454f42c65e82c0c960a8c0d5ed
z5c422cfa9f0a26a2ba74dd1dedc0c2bd18407ba889ca667c2ef68e411f72c35be9d980a5060996
z82f865969a997c432d5122f67bdff6682f81d24c7887837e10ae6069201517ba3bce08f603d557
zd61b7edd4221a8cd0d2a7ad4beb74d94f17e51cd7cfab7c48d14d0a69858bb6d6fda508a0b5548
z14a80aa635ac2fe5dacaea7ab949b4846889c204350832bc7866596934cc23fdd2cc5c6915e79c
z6e62591b5754e7a541f0134795a60e721171b9f18c7c7630a86262cbe282a9d72f5ee6e5b395ea
zc4a2dfc7678fe65ac9ae3df95de23e50cf4da32ef23ec652eb18f1dfe72b4847664227e4bf2b93
zf354d9ae7be4029de57f34dda54ec49330f9fb84ffbef7841f98e781694545ea4f1f9166f2c22b
zf8608c553373dfeb230cc149ca3143e927251c201991f02bdab3abd0bf6e65c7d6b04549f3774e
z7ef9b10dfaa5d33fc13ce07fafe43d17d3e69afa6b0f90c1a824e18aaae0b4cb3783f95ade8055
zb1b33c941151bec1ebc48a0e25382a89318a2c71971f90f1b05f6c9eb6d85747abde22376950ec
z21865d3c195a679c8723f11af2055201ef996bb2d630d8a5dd824f5f08b881e3aa8385924b4cf5
zd12da40b13c3f68aedb36f842fcadd18935c95b45371d26f57ca4a42800141fcc27f3161fe4eff
zc8397cb126c29eb042218214d27d7156cd614487500fbcce496ae0377700d082bbabb58c984fc2
zccba2d507b6491f9dc1662e2f8bca65d06acbd3c91f4599a18052fd4225f118d1749f3411b3ed9
z1dd884d67c8a12bb802e947f70cff3713d7f377759e4926d5c5858ffe22f472fc657df834515e4
z53ad71ef008776d4d4bd10211163d7131726f61580fd312d6dd561b3d33b20bbc8ce501225845d
z4ddb124d4cdeef4483290de1e2244b5b395e78690fd3d626c4dd9e5ae5782c2f7f9588629f8791
zb47e6ff93a9f98ad00f52296b547b82aad4fcadd5bed85e9da010c0a1ca40c29aaddce84a99ca1
zaf8864530b81b9324162d3d753728586b42c47f3220ad9051260370351c710023c1fca26cd90af
z306f952046937b03911eeb646af7b2bfc72b1f4cd26c576c127b74c6e59df484db21f525a9224a
z826d412adf562010bfb1d1e2e915b3c069ec22bb2e071f5297d9ddad8dde8051e035fc762c2425
z89ede964ce96b79813bc4f53277f52e2d2526d61353b06a4c03efd37bd1944bdccc03c70553a0c
z855aa32fd377baca46028568fbb6f2936c8cce21cb2da885e56e75a4bd9e916bf5836c25844176
zcf171a902844b35fb9b2abd03f0ab626a3c38d822aed49f504e8fcc7f5f9cdcd0b4b5eb092059d
z1e34e987d1d0fcadceac3c66855af268ba294853f2f3b44d3346a5a94643b912a6172a85611cb4
zb4dbcde878f0f90013cdcc5dc6739d7f988b5dcd99b6cecd6978494c660142deea7281808bb3ef
zf6b71e1fb61ff55d9c8d51d284d9f4cfb58858a4a892eac768f25b91d009ad6bb1223742b9da9d
zb7a5a04c6b37163d9a75bb24106d474ea0847983d8d3b0e46e3e4286eb4c642d8fd0510e2eb0c1
z3d213fd36853abd319b371ba850b72dee53a877c5254ddfed46aab7e1678b4d69490e98f6cbddb
zaaacc40ac46a74b48bac7fda0f53e795fdc438f4666997b12d07f57d8f05309af9cb795b51655d
z7fa0291c34216502f2775754df65c8647ac8143cf6debafedab7494680d5e46d88a64f74b501d0
z75d196ff94213e8c8dafdae89478bc491964b26a1f5f868a75c202360928cab5a32887a43f01db
z82070525ce779d808d7554a533b4dd7ede613567cf66484d2ebbddf31829a96541eb488537e290
z31b7d9f3000710d8bbc368b2370f97ffd9e5161a577e4e683565bd8754181e6d922ece3aa6f9a8
z6a64ed6813835b49367402630c8ad52e218287572036fabfe07aae88554e716929a2b31b182a19
zb1d50f400cc9923988c3054f19b1a078e000026deac4eb958760aa14ed75aeee0f27d473ebc753
zd7fa8df5de5b67db4c66d240646b971b18f13485b4619a519277bf76671b286387fb8bf7800e7f
z5806b84f01acbea4226c40afc6e7a69b4bf9b2c1af0a3d71d28dcc65433cd51a31177f32eb74f3
zfca9c43be4ef62284b79b3c3b3878ccfdd2cac4caa819c8522371f5384a464a3aff17dc0cd6f76
zccae35f1bce42cc51ac438bfe6c246536aea60f47cc04d44300a76ed7fc6d52bf749883450f269
zb95139fd5c66f9994c1e32d64baee9bc6abdd6b83b590b2cdd3c342327f8a574f69403eceb05b4
z964881f212d8d5f521f55890fd36b97a107eb14e2cf0c5b4f57b885be85a3ef63da41a10823acb
z61f20d1ad64e15ad20e5f2a830ed1444f89044eb720ad689a208f71f14d78780b0404461b4b66b
z939f9dfa5a743ca9ab9b8fe544b8ab84c3047c5ea5fc4b8f886e4fa5d2ffd20859491130aab8d3
zd73a81560f898ef552a3cbb5b6a62b9e43b4d9e21630c49a9af3d86693aabe36234226fd0e48dd
z9ab383c6c71b57f461d1a6d22eebc6c6101f00ace91bd01279a72a00f1d23729aa68d66eded77c
z64ead77d1ea206268d22000ac1fd377d757e16b48a4d2a4d5d9f9f9961ed173083120f86bea69e
z3ac6e2a7c778bfe05e30de93f18560cae691b329d637204d73d7792962d5c51bc43b416db46de2
zce666b319b6d086c16336d0d5b4b33d50e8a0f57a1752063ab78d2e74b76647e21de6427b03d27
z7f313e6becd3e8fe059f77682c73084423acab16bc6a3211777de7fe848f07694247bdebb4bc9a
zcefc46ec0413f6644a97a14138ef781b0f134cfd38231ed023735ebf28f1585680967a4146d3b5
z00b861fd6b0f187d180aaa05727309c7355c81149657b7d82233585c3055221ec4ab7958c82598
zb1ff14f612d43db880a8d0f805eb3f778ccfd38d0f0bbc86c44e36ced5aa260187220aa95383f0
z4c51abd876e53ab625132f5089d6066193aed763d56d67f2ba1987efaec2e88464ce8a14dab289
z7a2bcd541f8251caa73f4cefbca82e425837350bf3026a6aede4f6e83b5afd1580cd7e9da59bd2
zcb6ad08b0300d9d70c594037fa5be87494bd5528d6f6d3d6f36733448b878206901dad2b2d19ba
z372cd8614ac21a6f4ac78c7750ab4d31e2ff47403bdb222c11cb20d9f855b93ec10182ef405ded
zb0e7679dbdcf97912f0d1e409f6b7f51f22cf533da1c5ae3ed0397e5c59dfbf686d1a6ef1354a3
z2265df26375c17714cd18bd2170708a923ff7f35126fd029b17bbdf94b1d4ce6dc56ce7311b811
zf2bf07505e4cbd1f8f8bbb6fa7e1d950ddbc442a437f95f6686e8f43a808bc28c11ece7e6c302e
z8c5e8725816ed3ef70266d29a41a538a0f65256f4b607163b238e8f14c665cc5208c56bd501ddc
ze9aeda63779a253dd63f9007bb54dd1daf20bb51f2b85fe666297d3c91a8c95ebaf66d9c01335c
z3bb5fa22a8d66c582cb1578450aad711e78f2324bb257e7be576ce1f7316ad1038d367312aa4ee
z05229fb8a71691aae7bde99d17ca1287a700ae49a76c565cdc6707073bf709f0661c192da9fd04
z46cbb7d8e1116faa21e4ca7c6de42377866c8fe9676091b87ef3702bdf739b62fc23d778e246f7
z50edb11e6b03f4fa1b9db9362997145f19eb0c92f49be84644f3428d139047c1cb18e2c36eed05
z10cde2f9404ab1e4b159f202d4184c7997d17942499e9b11e52c16cc347e505db97deeedf1afbf
z0eeb9a6d0e3c9ff5523482278134a760340f5f89aef61f04cd0d7a8c9dea57ae59e95c82c187ae
z05d32319b309b89a6926a2cf2dda230c1c3c0add71b900324162a5689427bb1ba9fbc0e6b5f982
z83f0efcc6e59cb47eec5fe1fceb3c18aecd5d2ebbcf9bea1a997ffa81219d620f5b2e8eacb5681
zf49912ca6b3e24c6db69da946be35c9e2b3045b96894a0daf39a36c1564cd94cdbc24e3a7f6ba6
zfb9726545e5a59e9f0bfbda63681e30cc34523eb927b8942a9264fa954eaf0bbc637f6e8fc16bc
zf3199b56ac021a00c1b7324e3d3219b710463969e555d5b6c1107c276c8614f8a4aa5ca5663dd6
z1013078eb6469a2e684f8afbf01a2239eda93eb15f26bd8f2bd12002cfd11180083c250c0b11ed
z3702493d0e621acb38e1511c2bfcdd97126d25aeab8bd628872d55dc96dfae36750e8a20549fc0
zbb4de8f391ee0bb11f32ce986526424a21d3618a2c2447ecc790510dcdb1ed5051dca576f6a83a
z2b053b045b875a388792787b1a86dc948c86d8d156f155d676ff9de8887930d450babee290125e
z758eac058fd9f14b17e17633c9328d5d96845cf271c374eb55ba0735c58df10e1f6593d80c08b2
z6f91fd5143a3a1f230c20840a0d7cb23a776b07d4e65e39c613110e149f57598ae13999915a79b
z27b6583ff01bba0181384f8200ba60af842a1aa75401ea319d987c87e0f017be02399629d6f088
z2e22ddbe443e0be2fdbd54f1a2734c695f665af308b77bc4e3c2ab56234c90bc5f3382515ed3e4
z162b16be4c21f54afed801e7d143cf3270dc4e1781277d844c6fed4704b2c17c3b4de402a4f6cd
z45c193120a16b5febd69933c3a97be0688c23ff3697c2fb1903581920ede364c42eedf4d194f35
z61652bd02ea2bdd991f38be7d7d53b41fc01244537feba7967be683a669e73bb1a3c3b53eee3c4
z5425e0e9d022768ef2d9a6103bf51e5c3b435f42d3c32b368bf99f617841132fe4a09690d799a6
zbfc865b59efd65bd2ae660405f328040beeb57797bee22fb27759feab42a7cba5762b2771785e2
z8c49dae2d168c74fc041008d3c878d2c6761fef9d790f05053d42022a85ebd9e60a0754a0f3f24
zfeccea5ff508f05267e3d4420a11a54951aeef47df85e82feb850325efe339c54f0e494477addc
za032f6590ac1b2c956a62fde7a05cb55ec111f151e75056645b4bc853097196c16d6978ff17b47
z0bc8a954f4edb9e3170ab7cff1ad08ca0868ffe0353e97790be885855ef363b4a16f0a74127495
z40b04a3dd497d9b269e565bfb483a6a843feac7be9722485698b8aba751b513eac8bd3cf672035
z49931e648b47e0bd29d767648d6f989064b4f1f7dda9066fefdb0266179cdf01bb75850a3ce06f
za1e1a50794585bf2bdb7cdcfa1dd255b7a71c178f24c026502406a6c7e9ceb5a4ed0b9bc04ca52
zb694a8ad9fff53b1f0c3fe85ad818f5dee83f80ec51921556d4c6ed26f3262491ba184387ce5c7
z28ac393f023e6653c02d6acfcd9297335af826fa09fe7bbabd2f2fbd0eacdb23b8383942f41d5f
zb54d74d9a004eee95b1f5eb54a0e3ca6cd6c574eda4553c7cf7a7451b627797b0a84a060b89e58
z959dc81ba67a3404bdb1ce18761debad53e335e8d695ef093e425390d27d555c0ae17aeda732f8
zd1cc92eb6422980e4c74027cbf7687a90070b96fe62956f7458103388fa7d52246c14beaafc9e2
z5362d6bc272d7c77cab160f6616b96e7ef12aa9e8171e3bf237b1c3f8b7ee0181c8527808e700a
z53da989acd85f95deab46d67f3cf5ffcee0f1b2190d6acc94f599cf6305fc82ae88b999eef3887
z681b987b87629614f4df1274e53da3d417a907ffda54e3ee87129bcc68133c940eef5b1b3bc383
zd09f53c509eca729470cd9d795ee147643cab7ca7f8f4059ac087d1f5d1218cb762f71a12cb12d
z0d734807a2e783242f4efbba2f5a483e4e55fc0b7f69c97aa259c2c4b0b272ee8f50c63e32b41a
z8aa9d3cf1518b8f75994c5ce3c51867cab01c1fadc6b17f2ea3779739430cbe2bfa609145ed174
zc50614fe143aa2723dbcefc7f118a966d3b73c85bc4c220ee29f5897056ba59d763f7292024549
za68d8b9826e5cfe520cc43249c56cfadf29e3a3b1607cd34b12f451d50d089d656ad1f59c6c4f7
zd7afed976bedd3f049db9f876ece4c8e4b21051e058f66dbd9ef5759ab5969396c804a3f39ee73
ze8913054f34c235d823f56fe76dc02af9cda9bda07b9854a31ad54d8693feb68cdc07b18161d4b
z5683c8d4ef09672685df7388a3b497f9c27e6e8da70b68aa2a8146d229d1152f8c4860a2a00d98
zb4a34de7165b2cc89951208e2e4f93620c5dcb3b7e05f973978a34759db0b74443c87bd8152712
zcec8be4b336ed4ac0e9bfb3ab6dfbb8fd6ec6c0bad492a46f859dc711cc6186b8fbe835595edf8
z3adbd4e92edc717f474a560413059ad0f3cc92603abe8720ce931798f944000c0b70e76e128467
za67ccf86085055c11d04fafb1a37933e7f8009a71dd14769216545fb59563f4791852fedf5ae2a
zd0bf9fde5ef56c17af48900435fd78850e2dc23a3dd8f74457e06ed8d24d6f75743d11454b9d18
z1b5e7a0ff95932f45cdc0b598dfc565ff86419b80fd7e67fcef19eb2a75b1acca49c0a903fe5ac
zf39e92967c9d7ac5cfc3c7fcf9a54075d6151b486585412c57bc70fe21db9ff736b5c032fcbd6d
zadbaf9831dc793b14a03ba8cbd9ca5d19ed62828c1aa05a5ca01d99c04eeea02b8115089e9f5d6
z95706f36bb842c6403c664975c4cde8d8d70de2b0ad364144045da21a963733956447bd034abc0
z109fc85f3123d909edc6e9589899595a9b6a194abdeac63f9771577acff2cad9937bb28dd17b03
z4bc7be3f70dd6c36b99279bdc16454ad2d3a7f10c4b186ea6a3fca414e268d0b440c013add174d
zc4ddf26099b365c4056aaec0ed9dcebdbdb4113270f20429e9b1943ec66799f968037a850fb1f0
zc785f7e4d1e59a1e213201d0ea121e427a11fd664942080ac73b1b94f07d3d8018b8c0c422549a
z142d4ab0cd07bda39e3a61a04881eb34b81ac22bd533ad10de00621e4ce4241be21d8e627d5d26
z86d239f1a037408a5667e0e29f6714ca52525ff3c3536503b5a9b0ea08638ed73d5a3db9e9ad44
z79164c39536cd8088e8384c050eed7849155f038626594d4ec27d72c4281bace97e9a6caa08310
z1aaaaf5001e15c86688c0fa4e68d6408e386dc874a43d26d8fea1870420811311a09c31171df3d
z59a5ccd6912059285c1897ffa41a7d677e15a20c311e4c9408eefb370658802858815e567bd78f
zcde8245c6336416277f7832f0fe1c57ec0092c233f11cd0cd3ee3b2a398e47775b898786fba2a3
z2cf9321d689ba7fa5d11fa079b2a625b33eb72ea649774b1122490d976d4d694dbadd5c4aabbc6
z62e3dc75e7949753a072c847689d0e1ccbce88f023fe07cdb3abc486b6e27bcdbb322c58894417
ze6151a2dc21976a3423871b7f6bc85be2deb4a2cc6712939fb3d876bfdc563a96354ed5c55d6f3
z5d6beef3bf0f7d0b4414c465414f2d0d1353d2a1ae191bfb470ac2533107a0eb6833806a229a01
z9d7ec144b9068c5384d790bb33799aa47348a919423b698e29687ad9ea3cf36a3607c031cc316c
z410512bc1de38a023b349a0056654383c18022281ebebfc02433ed1305bb9d49660ff70047ffef
z1bed160ce6a4efdaa259a1da715b78ce13894adec5937e1d68b8a1db2d6c2f7b2fdaad6b07e574
zbca61bbbc6444d7897ecc42319612c2adaeb84005b371b6396866aff1adb4845d76b2c5d2ccc0a
zd37da86b66bc62315eee0563cbd4f435a83db10c61fd3bf4c57bb13295e3aa8f3d9dd1beb0febd
z59091848c9ed769c4bd0da04ff790b03f8021ff9c607df9b312894d96732d06ed6cc14d0cd3061
zdac384ee0769cd0f0df15b2f8c08def19c94e616d2159014d6152f34b46087ab9a98e8afee362d
zd203c70a8d4c3e65f01746094b2f991c78050ea75fc1be1927ff74522302b00c7decc1bbb22bac
zb65794b058737627d395a985b4fac202e650dd302b678bd8118871e26944f83dea7dba6e619a4f
zace726d3f1cb6d83e5d1d0067362fc56f3c77548708ad66c65b4c2e66e08e83b6eec06decc619a
zf589761f4c3492b34a651d975b0258a0ba7dd33369dd9cc5b3461cc2f7db80ca8765eb79cd7cd3
z32f95ed8a0f693c4164cf1d37b8d0bcb7246e19502de13fc89a400b125ab9bdf0363168e6c59d1
zdb0710a9987d7480e1745de3e6b7ef6633e0c58a585051c336b708eb20de3292f2668bad8bec4d
z61295c86a4e00a68468a3e69ba75c54bd67ef7c56b711205309deedf28482371ecc1102361f319
z5d7923e0ef3dce8ff73f79bb0d3c445f94046f11b65396f0bd9d0361599b9d7a2e87efc362b086
z62f9662a377d54d04d87604460c63068d1582548df5ac8c9564b5dfff54f30c66aa51c3256511e
z455a5d64d14a0816321812b51797d21467a51c4a55ab405c316d844fc2a52d83bd79b148d3a6c0
za3cdb7439bdebd5add96141a38709de04710a8e4161bb3c96499bc9d5eaa43ed14fc4ce2971542
zecf09d8974c263a8afcf541650bfc470b441ea992a7e3753bda197df3e1f6dac4c44eed7ebfc45
z5b81c33bd0d903c6425b8c0db6075f9bdaf775f619202be199b7117a673f7f695a7062918a297a
z03bd8e416a950d3108c8a4c5e2607a644e04384dce549dd95a5ba6479a66679884363c2a9faefd
z52d9622c757023f76fdad1f7d3d5aac2e36713265a4ed42c78316d81aabb207ff4c0264fb6b3ea
zd2e7a92ca7b85757790cda3971fd4e894820be70fea5e791db0dbce5295be9b354d4b6eb996ba4
z905aa503bd0565949a7fdf617766c05d10d8d467d7198c9adfe77537823c0eb0e7a3ad8dad9537
z987cdd498f2fbe786622247e6659e7be079afaad98e0ecf5042690463e30824125fcabca43cb07
z5b825453ceb9b61b17a5f4fbbb63e0d94824758efb0831863c213fdda9f430308c7913ed78c897
z2c9a01f68030b1da19c918971962a4a7bd746c7a3e6861332c39697b4199fd46c720e3ea2d657b
z3896e950e94d96f43813a8a0426b9ae7336b014ab0297968105376d11749b8256ad0ff90fc3f8a
zd2b5ed10417f32257048e98acf617f16717d06164e05f6b2fa2aae4a9bf3eebda2f6dfb48a3d69
z0ae7a0558f1d245afc89afff3124a7f909a6736f5015b9762721076537b348b2ca1112a160ce1a
z73088e542784861e0aed2eb4e04e5cb51ab4f3cd7c1d1862400040e243a959fd02bd8d28346db0
z67806f189ca95e72378a626903f3eda0a7ce2483d5c4be5bf0b3036d65ea0dde71cba74fbaa5fe
z351916885bfcda61c0611aa96ef5305d41d72b7c32d34e3b0ba8d952274de60b865a1e4e4364d4
zca0581c0f6fe0e19a268d59659d59ea16c6101bec1f3cd9c91b8a73833de2974bffff6ff79508f
zc95abfc85a35953d73f58a7392236887592758152e2d179c7af94b91642119c38bc28d1c076d8c
zd6f06929c506e32d6ede864678c785a17863ccb2c7b38dc4efc39fd6d890e20588dd1b3ed6ab28
z4172c4c94323c8491ebfa3b353dc05bd54eb9ba9a90c45d789820dc295e01d738620e40fc54182
z99b9eec30dd4c7ca15a0a0c42f7a7c692a057e621e34341d4892f07f4c164d5ddf2ee5faeafe12
z95418a7188f8bd92db62e58728418f06ef3f97a1eb47ffc0100493ad63dc3b1426524fab65ec8c
z4cc44d75d8d38ea412397b3623a64544e2494a764ad6711d1fb09c6cbbb9c650853760706f9a60
z5807e96cd1ed6b55c5e5796570e13b4d88dbcb3d0b0fbcd16a5d43adf55f73f6c7fb401cc9a91b
z5359c3ecca3d2c3bb799ae260c73f1b1c11bd220dd2dfc4be72ee7eeddb279b84e0b7231c7e21c
z0e75f0a93072095d08564a312512adf660a30b565fb69a9df526648a152b11e972fdbafe81fad6
zf9b8ec7fafd7ba4d192acf699c9e54d3be40ec0017b3dc31b8f843db4d7adec2f67aa8d0bdd55f
z01d5d4f5cd927e13c896b25a22b742a0bf98c1a194a80696b887bef8bceb755a09addd7cf81c7e
zeb7c9a41bb2c0420e6bfc111c7ad377a41c8de6f1af4e077752e6eca3ca4553719d02efe5710fa
zcd683af5a60fec53a212560df5b79551c55958b2152726a30026c6085b5161f76fd5ad043589dc
z3dd139e8922213496cb08d910376adaaa06bee335c740ac7b655775bc50146a37e8f72b8951506
z8117ecdbdb2d663fb82f408893e4727ef9d21bdb6fcb915c8d2e60a982b7d4ef640923ac3b4d9e
z4c6632cc367ad8959f00dd8dcbd118a0727a7e66d3c82d243e925e743401c86f2c778d83ed196b
z931261faef0651ca9c8b9622250e96c423afdd4407333ba9c52adc3757a0697b9510a424956277
za7c9c7ccc033cb6b4643eefea603554cf98deec9f142f55a6a7753354d05f0ea3aeff7bc043f9d
zf5f69e5c55c17932e88dc8eb1f17a6858e40823ffa79e0151fc836ade907f3e1974d659794c455
z8dea95bc70bdb2c068cb557b52d0bf2ebe2e1fe64787732322e6d2b2a71e98e3554e4e5f81c120
za9a3ef4ae97f59db075cb4019e0790ddd534563ffbbf360310ec33416d0c8af8a8051c87cde35a
z54079bd04390d51e661ba35aa72f9231ddfbed03d8fc4f66002f0ca423055a49300874fb8f38a3
zf5a5c6e72b9b3a7ed1bedbf161c6b2e80dbf811b40bd1f0135f7fff8e60bbb6be776d20c949f66
zeeaaabc2c8abb1133bd1056e91485efdea55ba825c857cdf619c0c3a8ffa043b940d6c2e45e3e9
zbfb2f15d9e10796e2f97293cfbb8fdb124e38c3cdd4a1a73c76db191c10e933a8154f9d8eeedc6
z051a99480417e6e26a3062b27ee256f9b025ee7554bd4607f67536228565b0448e7df721c2f3fa
z634acd68e807ac5594cdabdbf471126541747693893a7ef87140f341805d205965f4032f0151dc
z39410d8a1b389b46d6ec823c5902fd8b11cc2a36862577a5f4ac75d808440ddf67a76cbd26e651
zdb6c106a82982c0ed6f279993687f21eeb1b5919a920541f46abd0c91730ac69dca56708d4674c
zff43dfb2f39b70e93d81641ac4c530297d108056be08d2cb10b9063190b977af4a1ba9a6e5f5ab
z09a5b025a82f2bdda7475c636336f34825f02bf1110502a2fd3ad7c21f00df84a643a4d94d1ac1
z6f5a6feb7a55d15e816c880e7539309eaedcaa9a15dd687d0057db950547f4190b7ca8a8f3c981
z6ae2703a636095d6ede1fa8b7ce62ccd1fdb6ed52aadee10b656658493cef76ba1a2d156d6a18d
zd4d0b993bce30bbf1d4cd352950972ca9ddf50099fd584393c68b440ec5b2f356ef0c1f8e2fad3
z25e7598b0700d1001113a7dca1a507d1d32dcd14b9126678f3f0c7b5d1e3780b317c7f9c4a7186
z7724d899d084488b944979a0e419c06b089155815f06c1fe268e8321a2931ea0217e3853bbad16
zb5f767aa97a49cabe97537f9de6fa2a20a7a4991769635109708d33619189d722aa010284cd042
zd8393f307eea220f0b7fbb6e31c60406a361b374c907b04f924259aa8f5684f6c8717e0ec64fbf
zd8eb0ea9f102aa71a4ae884fe56944750d4cb7d5abec7cccfeece34b60e6403c88e996a1c3d21e
z62b656914c24153fb4377f02aaf5c93164250a44e7289f79f8298c53ac18facfbcc5defc12aa7e
zc0f43087d2a2fd12b542f74c6493c3daabe0e5e414d75b7087853335b0aeb51f4ca8bff736264b
zfd075e3bfd8565c27197ecb8db18455911430008c38965d6f3e81f563a160a0bc8ce51cda2d348
z78bdbd0bc4053879f1ec0db2cd03cced75b4740c65ccab3833ee945ada1d7943765dda9cd92d31
z6d4ff2d9822fee95ce260b9e09303014731dea206d97e2955f02c6334c50bcd124e33eb8f1fb02
z7fed2529e6414bff410324d96500c4f4221f0471a8c6700c6666e997027a69362ca1ac6c6a5619
z91c18a6a5d81848a86f2b1a2ffe43d1cbd4f5926b5c403fa9c070134983c9c73057eb853d8d32a
z8b0293c59699396fef90c8a61fef2b089187fa63ec1999dfabf0feaf22122bbc3167c646f17bbb
zdbe905526eb813492273746e9ff0bdd154e4650b1e2cc0514fb6e85cb7415f856d51bb262e23c1
z6256cd7369f45d11d7b4640962a0a1b4dbe4921d3cbadce75dec664068ef269196a7808bd168cd
z8a28d87e254fdc4c0e44df6d0afc3e9fac309f98267a54fc7d36842eac7e5c191b6f38249b2b27
z6b43a7d30962e5f1a1a9181f5e78aede7187e41852f120c7f2937773e524fc01666dae99c3f162
zdcf5303adaca8df8642f49868f8f13ccc66e98ce5aa20f1a3fdd0fc25f02740336c41a669cf459
zc134848ee99466659549f87f3897cf96100f0da173272c3a1227291ac6d69f37dd12968650492c
z8bb7b5df8a18ccf2b4eeef65b5569e1343e0507983c0185c3eac643191078531015b2a304ebaaa
z9b6bdd64f39fff170d818d976ac520ce6bb20a1e92ca8fe41acc4a65b71168b53871510afbdde1
z7068506f42dc057ffc0da8c3454fa59d5cf1242007b9778044271258268ea18ba13c91423c41a4
z3203b1620a1ad3b3ee7fb7e1ada7006e648be46080076d68e619f841e4a54c5b8f6ce995438ea1
ze6f19c15bec1093d2c27e92f17f36ec06b314abacfafab7d699139c3e255764dfd3a4ae197fb53
zed4321556769eaf83ddd21439de7879184e72e4a3cab5feab47cb6f6cd7daaf2fda7813c18300a
z9dad9c9b36338cffa82558b033e39e1718bbeee222b67c31a0e87861c95438a4dadc4b4c04dcce
zee10942d6665c22cfd66b493c1bd04d27c4886c7c9c165a627c3439d52baf9eb6ed4814e268bac
z986e6487c63d0a72871c02b701b2aaf59f7217fa5d71d125732961aa348765f7c4fc338d40be6b
z4bb485a3b73ad616ee932ab062c4e965947dbce57c4735f53c037469c89cd1f65b71fcd611114f
z57accc411a8b565f65586d85620d489d35bac87e0c96306699f5bee12de5fa9d3fe62da9be5d13
zeb60764f8d4e3b9cd0bf49bfaba4e86de9e58eb4acb0a81ac429b91517e3946c320a65edd45c56
zef86d7911745ba30b48c5453fe9758ddcf8cf4f935997cc76a1b6636767154094ef70da24c3618
z11ab8b33011656745ff149492509fd1fbeb4570f10cd616339baa812fd7139175dc10ee0cf2001
zf3f85df13da22d47c031c2f204fee51335079093723e786be3fdfd9a62d1f09178e7d3630f2b41
z8f7d284eddb264d953910e44dc065c438d02c3f00bcc33add2123c2bfb06134224ed5d12c65c3d
zd27f8d3a37aba15d709d39d1c52e4257eb9bbb6115e373f34ec71b8c7fc894a6a1cdbd36e5a5ab
zd370a74e033dbb83d6139d24d39449bb326cf080dae9b6ddb6259a9a050fd1fe3157405b488182
z38bd777ac71b38aebbc46a38c115ca638ee688f8a349768a7aaa5b5b2b11019653023161b04823
z71665d46230fad5b4a621e49652d1845ba4155b654b93c411ee75b54aedefcdfdcf73b524bfd79
z79652a07a8061ee26b90d535c9c4208d39f223a0b68027bd81b17451eca207ded066bcb858321e
z47ad878391cf93ce9f26f43f4627f4f58613209b1fd8dea821274dc8f873bdf8563fad67fd16fe
z36eef67db037c315c88a7700056dd3f111b5de6bb87e11f3eca42485e13eea9fe9ae5c6f278c59
zf94dcf90964d2a0d53fb8be1201e350fe83a8ddd5d29d73f4bcf37e5b0c3ef136fbefffb121973
zf6129e04d3661b9cec91f0c9ee79b160e1386b7edf0db68bbe118ddc82273decef350f0bd1e555
z4f7c839dd526f3a6f1fda872ddfa5a494d1103cefa9b4211695277679af5caa8e700d8cdaba931
z3d4044aecf4223aa1ef993c2eb05af4bdbb8adf3d3221c9bb2825ba369b960deda4f75939e041d
z7de1af6e68c8c4dcbeb55f5d4b18192097117fc09edf0492c80f412f1d3cb6e4b3d622ca85008d
z0b619ec8752fc07a0378ccceeaaf29256488d5b816609b733473edb3005452b67fcd8c83bba4fd
z5837a5e7b348ac0197c229c193db4ccdeed5f1afec98e764dc62578c6d231bf485b75d744c3fa9
z138b03bdf29a556d78722280c6533f967afb13d2c650e05976e98aa2759349040763bb6c707d4a
z534e4c3b10ac5d4dee0e09284be1ff39a7172b81ed1f7f73531ac7e2163d462e90bb2fc170a313
zeface1fe3d248a7dee52a91c0bd69303091fb7aa60acdacfe9997448b71eb79a72973905478806
z4b9aadad5dcda498cbd14d3d9d4dd8a527373d703f2708f705a2826859bf1988fd124083998062
z032162384bc4b148d7a62abafe310812fa768d0ce6ff462aba66f57608aa28aed5ce0c5b541cd7
zab0c3b6168f892ada1a7cf7d09fff7aa3c0f01ae79283efc27783cfd13b85e32953a52a1ca1277
z095a61a03da3912f4faa8018ed6f640fc8efbe94d2b5fc0115bca2630a40fef5186b667aab3b55
z938b52dce18cc22d9f4d5a5ed013877926bf8a1396f9631081001ed1318bad50c0e4980f89d671
zdb96920043e96d13acd420de4e2fd5611ee1f42f655e24fb3a66fab51869597adb7766ea8eee6c
z3e6558ba49a725df751ae8fa08a480de8402f1367de6a7dd64a96e02baa89848435027b22348be
z0443f35af83d183786e3e41a7bde1bc312dead30decf5261aeb632fe1539a7074bbe414ea167d7
z361cb517dcbea61aceaa1c6e49bc7a82d0d36c7e00ae373e84fcc6c370dd2712f805c9600665a3
zfcaed95a1f77feb81d385c1f8089bd60f8c04fcd67a95e693f78e0dbbeffb608972513119a42cb
z24186fe6ab0c12dc7469233e6a02445569958586950257a643422be3a343463cb56c438baeae6d
z2675c7fbb1c36824cda56cfa64fd855df67d874d0bd96d0285e97e85575eb97d8a99ba37f5d25b
zfd223fbcbf1ce90d3bd4badaa484375194cefa4e15943bd7f37656ab88e0baaeda65f947bbb97f
z8f1c5793a78c984cb620a67881e54938fcc18c1e869889e70dd175eaaaf0690081cb83e8901c32
z4cc193441c3e55bf991dcc791d11ee48222239e98ed7aef276f273abc28b054d179bef929ad075
zb6afba91a20a5e5f9d35763bf0ae59f1737300c323a4cebe57c2535a1e451b001f2d67663a7cda
z8b144e066f34f93815020b8b58d7077fbdfa6921e40a64b1e8cd4057ce82f547e3e293fa7dc3f2
z455ad3d24282d5fa0ed83d5dd2614a718614b595a3ea9da4e58fcd6ea22b6c99780dab96d487fe
z981f86a8b23cad79e4de92ab45a6ce0a7a602f18ebbe9200e3389d8e650e35904f0bad18c54d0e
z194eb7ace6ed5d5f9348588bd14f1d86350135851c0cb5c052c6d57db2f2510c6f6e0aad09fe46
z4105504b783e0c47a3a3e9592feb25edc40b994a1e025b477123893fbd340e3d0624b45c68af2b
z85a4c3ed773050a705af83f819b91aeb6eddf680c64572220d32f5699f1d75fed69445b6f5bc8c
z3086ef377c192b16598aea8db1c74e72b1c00c90244977486580e12049fbf53b1420b3b5c5b775
z77d095c7645304c4df861e54cd1d6c5d5d8037f878fae42271ba0221c0d57559ac00d8486ffd72
z061e62bbd48d37372932d6eab8a5817717c5435796ace08811da8bcbb6b92ba5ec2cea43372b81
zc25d1763ebb91caac9ece800a6c8eb2d66734348b98553788595f46b44ddb70d79e6bfe0584f48
z5aed6a8529abbfc399fe18aa5049387a5c4fe9639aa910c7eef300f1feaf4b8f752684d44c92ac
zdb33b93fde53d88367d953186cf2f94927ab24f2446074639c1e66579a4a78c3971b1732673cbb
z5aa7db0cdb7e41e90efc5df679fef8c99559cd10e057711a6d915dafb6280cddbf03023e273f3b
zb17431d09d1699e0f847a7921cb930835de7dbdbfc35239947894ae2d808ef1a8d2398993b7a33
zfafa47377dfbb253a5d9de2975ee81be85c72472e78db1d91ad12668910e8daeb227b7517eecf5
z86e5dbd9371ab635fdb02a7f4fb30e25fcad98f89c425c41f47115b2f582bd5fb5f70721bb4899
z6730bc9edc1ca46f18eccbb960c1ce914f4683cd0784c5702e941fb6fbf2f818f93ad23e4d970e
z5b9d07b3b32fac03c86e3a9c184f70e3779ce66e670b5de750a928f93952a29e1d0f0e90341b38
zab5b00800fa9a23b29d5f37f95cfbb14ddfb2fd71db5484ba86f6f65c6b3158bf1b5910aa6e549
z48304a8f9e1d4d08b2fa2b96e902d43042a25eec7031064c1c8232286132a6f7b0e9c21c79aff9
z848c3d1826c5954b404329641b230a4292d2f40b5165c3bdbc01b894690ffbe92adfba8fdd97c7
z641954acef4ae79f7542518c28ce29e430ff3ae8329efef89ec156c1291676ff24fc84d247190f
zc4f514979d1dd80a0f3c2269f0a65e0805bcd2204e09a9165a9ec545ca7c842b57266158b47c57
zf09a37c94bac86e8d3eceab30f3ad4203a036c8992a3b32ca7644366f8f0b93670ef40c6b0be7e
zfb385c0adff31698441fc67f7800b222ab35af0de56e45d6e651ce2c99de5fb05a05e953a22038
z8bf4adf9b67cd4e021c5e6b8f1cebfd5ea10e2d00d75570c8a2a9830ba963ddbfe579644fd3e9c
z5f3fc8263cd09fb69effcd471d077bebf8d3b1d8e0190d76edc9461884dbfe8b58bb32cbce8a4d
z678dc636763e606e096c24fbbea008d517c4e764e356dc828a91e43d939f9d42d724972d4b4ac7
z5524d5f6485733c7869468fde0b1a1fa7b6f21b8549cc02003d95be12b4b2e2bf120a165f95b20
z3e42d474446431134763eb1f6d756bff4acf4bbfba073ac71e707b90224e71a8947531e2d9afbb
z4cb0c80a304289067366ebad6c5c92edead3a9aa3042edcd58f9a3ea042063e9a60c3a4679efd3
z61ae6fef86ddc6efc57f249cad8fc5a136f110cb435089e401f7dfa9de6c26244734f2cb857df3
z26f92f89448666e23073cc189723582c5e510c7f244ac0c701ad4983cb0515d02e32bdfe847799
z493c3e16ddc42663407ee15e64130389850f391b58aad837c2db4d8cc5c475aefe76c1a8b46c6b
z913fbcaf348ef3ba5ba2710292b618870f80b18d6d3688f37cc403d3042e9b71a6d8c7517dbf90
z23bc5da7153e8622e13a22a0952c68046fe043e0325a69896e7f96fa45b0986b9cc1a3a072f9c3
z3f27a40dc122debe7888ee7cea759c5892e9d932bdd5abebb19ebd9f6382c0a23a2dc9c7a9cfc7
z94f7203b4ddd238d2be1f9bba06903a4d110df46f38a142f9d0149f5592031e5bfe9fb29bc8c5f
z24fd12ccbd559e2c47b10a4869cca591378fd0e329f408a67304da8fb16de69d2094643d693534
za97ec97b930e66e020b45134620d8057f10de7a14f09640af54ebd5c73abe303a2791b03314398
zf12a65c27610269e2c08b5776c547f5cd4df83e1c713bfaf9054e12fb12248c706912134bb4a4c
z5570a70c3335435f547d26379d6ca819c94e30d75e0eb9dc94ca25cb98e6ecfedfd18b03e7147f
zf6889a2fc76d488353d7ec232f6a84bfb0f4e95f3fa9b55e812143ebd2a01f198931e7f339a488
za0e3f55c13897be6d38b1d47658b6987ad18ef6430388ef6510c1c9a66e1a713126b125d946db7
z903c51a2ab3ecf5525899a30a3bbe79c0c315c357c4016c751c460808f26df87a7b3ccca096a13
zbd22fa1f2ad4df00085238a5fdf764c7498584b2fb67282b3c4c30b3e6693cce4b1d2a9858c90a
z24178dcd54a3d7141590c77f26a5e6ad605f7abe609cfe31fdef5b16dbb534e9e976dba78adfac
z7bb9fba1ddd1d90a7b640a2c71a1a3daa11a8b96de66a5222030984b00eba7b14ffaffa8f61ed8
z9089ec554354f89fdf5143021e8acb685e43eb0b1644dfa135624e5f9360d3076d305b09fdc307
z959c68992a419fd9a2771b87fdd6872379096b56561f65707f83a8912d1f9d414a67c375878a4e
zfe3c13c425039806817e9a676212d96772f7e8510a441aaee7fa5b38df9915dff26721e9106234
za061de27538c723b300e54903d0055e7f065910b7451139ad8f778ec6b02365b7c5b83ed04a40e
zdfeabafb76d221f5dd1bcd0441ba6172657568dbbdf415a0310d21c31c2f1305d7d95d95d11778
zfd574694a1746a684805ad7b2b54d719f9a5d2bca8e637df26de47ebd35ec9604aaef61dc93c99
z80c12ac05bb073e2878857d1e345a0b11252fbe186098a56fd13ee52cc06e0a24868a66b77a2f9
z0694fd13eaddf2d908f2a54f9344de98f2b8479621e9a4709e903bc0d455911a5d1988cf4adea4
z6d645c9e41c72cd4bde77d7361b011f096389a9058ae777c95f477a695ea05bc31e792313e3b02
z2c71efac42f97f956cfbee4227b4286eb0ffbf3c9968d94468a669b84dd9120e166780e2badc56
zb508b8fc4219f979ecb64dd6cc4398dfef415ae286066ec0b226a73d9918cc8556342cd463f8e8
zdc5f281bbba26b15dc0577c26d0f94a738b1765c0e2e5bb187f1fbc085fa1241e52512930c22b8
z9d7343de59c727bb93b798ba57b7faffebd19f05db74073afde6cbf7ba78f81cebb587729017a3
za433610ef72bd3eab1e7fff7f6c555d4b4872df5cb6246d4f7aa428d8148e80389fa7c444d1fbf
zb83ca777530e51bc47bfb060602bd5c4d22552ccb531513ce0d166fb8a1b4ff67d28b1333d2ba9
z144cd3b0b245f76599edf7d00e7d66f5d474257a958e9be2405a20eded63b5a39def631a874b06
z81f0615965721f3e39a7098208fffba2791ed09c79d090663af34c86fbe666ec5191558edd5563
z68d32ae5037f66c691f49f815e52cbae788c460af3fad1f3764f94a0c3aae39edc8190728b81b9
z63111e835b36fdc8b48fe4c1233c6621ac94c9af56f0e8b8729402c0682c83518cfae02a7cd070
zf05396f35df245e7262536958d344cf431029bf5f3908ab8a56fba11c498d23a316d688e64893f
zc9f82fdbbf27d842edb644d34a2539d5b7ab4bd956d00f9c073199e37a45580981a931c6455920
zb4941df322ff865e66e7968157584bb384250e40cc7607259d104e8ffb6ad4523bbea56ff8f24f
z44b98edaed4b85bcba864a1433867489b0cd6199f40ee516681d5c6096421f4aa5b9311cae7a31
z96550561f7b46c608b4af0d03155d72728cc87533d2d17c088f6d85338f850e92fef0411af4cef
z358f1d1def28b9b46a86c344ba8033b75de0e5cd9abf6937e323570d53d5e895689150ade42df1
z5180f78de4794f9c00e1d31388642df36fb4e42ec2ff7f4096341bb26642b857a04fd8ca46b2ad
z34749cf0542f0b9265b71399eb258dcbb0809b6685feb2ac57c6ff5784b3439c847fb371dd82b7
z53cd990689d85f3ba0b09093634c170455ab87a3b757a173a1c6304e9669afae66649e32277317
z3b0d17585dcf04da021fc328f872e50ad33508cd167de0a7173e5e1efadaa39b3bc2b6be7a4829
z73056e95eda2af70bf1a04fe8e366c9c5cb2de10bf3b6d97c0a8f5f8cf6480a6ed3e69d1688087
z416cd262841cfcb557da7aee7268f803d144bd2e78bceb0cbfced42d14234b5678467488bdb26a
z0a25d92ef8000379062c0aa350332275e3e1ee8c82fef8ec99d330fac644c503153ec6a354c672
zb4132736a4cf55e8be9affba7b513fe2195069b9d57f2f7ffc2c5dfe35c5b9237e728b716eac25
z737f41241b6130508c054ad619b80bd94c4e18475aeeef022da75b66f5df122236273964a54ab7
z35382cff19a2d931f6f37e86dc4c63396f46718e70f7d8666e0f851631a9570a6054aaeba1f381
z313f25fe69f3fe0e5759822f4f0159333c827f9a70448d25d8c58cf95610920db44cf3c1ff9e0b
z65fa4469ba424fea2caae66ebcb764b7ec421afa0e7bbe6d6db522e1472a25fda583359fb9f97b
za252b29d167378f0ade269fb4208df0fd44cb397eaf5051ec54c6ade1bd877fbe70c9954feee73
z76540009bf4a9f081991c82410e32083ecacf2746f093580af40a963dc5e8d0a858d01a6629d83
z00be4ddb845458ec6f0616865149566068e9400cabb2977daed8973eb96bed63a9552cd37fbde9
z5463be75928866b81f9856474a0ba5e915fdaefdccb0a5d57c634a852f064a7ddabe55ce5271bb
zf6d21d17eb71b0a1dfafb7432401f2e336628124cabddaa363a8cac8ff9568173a3866752235da
z64e88a51ed2d1c6cd9e9920df249eb104643d1d7ba9be7b0b787cdd961c952b9a963c7b071ef4c
zae7d8118fa6e98a66041a0f2576a36d6212ab6f383dec1a24da9c2c4dc28bca1afcb5873d8edf6
zf62d5a824543a8b65cf89737306a4ccbf5cf4e3a8c135b86f65dbe4903f7e513a9d2571de49ede
z56e474b80619c0c98597b0c0308191fe6058364f7f72ff303bfe31905f02a6232856ecb1da0a65
z669946e0d0aa3b9114cc0af62a0564fb74863a4b7a77b5a4ccd83dc83adcb5aa6d47217747a80b
z2a198aebbe75c92649c5b7d1c7d4d81e94236b62cb44a09ccb57b71bff57c8255804c7c1153bc5
z284a8d538fa2b1ef7378f33560fe5a6b2b154a69afe9e51d777dec7aa5621ecd48de750fa74efb
z47cb479a6dcaba79f3ffa12daa26618c3346fde029b456c5a87a88b1eeff4d52f873b63af02c47
z5061df0d13dccc65290ee6ec677dc403716b7120e579322816985a2b14b10db16e15bf0969f82c
zf5c581e0da5bc72f5b03466c4b65193ca7bef45f883f4595244f439a4a6a62d0a5b83f6eb8a488
z04dcb1213345b2edbeeb67f7846d03c25449058f9ccfbe5bc26297f641e1eed449e8fd64b17ed6
za182dcd85ecc7d4d0b3ad36cfee18f3da404f18029b2810d893c0dc13562f4c10002c9bc6e9645
z82b6202c7fe83d8f7476f6d22d183543dd8dae71d055a2642ecc10c2fb0b67c356986a3d957063
zca5ef75482f1a27b5ce83bcbcdf49090821b32df79361047a5b0ef9fa1c76a1979dc96cfa08e50
zb28fd7a78da1639093f6df312dfb1882b6c9d3c175f6a46357ca1e2be12abf5e33c34dcc5f1aa9
z682a7d0142602bfef7aba1d3e31636e26d7aeb17dcd0ada1f8b8c234738066ac31855cf40ce904
z54b9f938e5827e7419663f9199b415888c104b83003c7089824891816bf1c00db427c72a0869e7
z1d226ef5f88e237c1706ab123459b8aa1eb16197b343d1a180b4c47d0df62db7c487c7d196e3c3
za0bd59ee926b7adaf5ec6dc8e8a5ac7e739bb66f45e073f70292025ff70c2101cf151a83055439
z045f866a5a0d3216ac30479ac1d93a084b4cb7898b17d9e79fbdf35a37a3eb4f050e74529cbb81
zd117605b1dfd62aba208181c05efb5c0d825775c5707682ef5801003909158b7b1fdc370a51ee7
zfafdc69fa3328d30c99aee2caa5c05ed556dda4949a9b2960dc1bc517b5cb00dc4c6e2be62b8fd
z4131fe549c7aa8890f6c64e993182c7a19f022d7b138f31f7bbb40ca3f77461f5bc5e6ebc93db8
zbe251c5efb686fb4db22d85ba0916fb0b8a41a84191413d4ce13fd51b4ed18b61b5a0069d5223a
zfd74659748aa199e27d32863a772cf90dbc32edae218345363ae55adcba6b035fb779c21f6b18d
zac7d7433475ad8a74699f02dc661ca445b3c1a472ca89a7795973fd643add4268e8294bfabeea5
ze24130118506cc3e6969e8fc3acf6485345f1590cba34115b8c4051659d906da12d258bd1ef612
zeec19e5f1f024a97206b59d2af1dd3e5fbec74d0e801920689acd6707f5662b4b368290537c9ad
zdb66d63e7df3a02af12cf5506ad89e6705ce345dd7ae03f31a942f7e2fe6f920adcd07739c9d06
zefa96021199e58c04825ca48af77d46ad14993a72dd486c3cd766087029f74263060f01c1d88ee
z0f3f1d0c5b768dff90c0a6f6af898e6dd4d99a6d412f6c4c04619b69e19e804e97a393fe46459a
z190a0a352d5fbcac2aa3d76a6af6c4ad662da298f8e8d0d71aaf51541eaf02753295bcd220ce5a
z66c0dc86109e3543b0ef6e30370d687f8a874182b1433342ceef532146fc835b5b28ea1eef1e0b
zc8e38826f4ab7d9b16695f565540e36b7b1dbab3ecc28b264f791a8eef80f9283d28d291b98203
z545a2a22cab9eab32461b28dea52a1d8d01571a426751c178845fb6af5dab582ceb60aecfb9409
zae8a0e11db068e7ce5c1324a45891d9205c0a3dd87c87a4267eea500d88771129c355e65af1800
z2502f1d70f96cd9f88986cf74a451b7c202c6002677da2bca7265bd1b4395035bbb551d23ca179
ze9011b44942f0c246ce5bc5a3e3a4f300d94535c33aa4424a24cf5dd244e7ee8d695af056f0d56
zcdc7bfdb87294e2340ec18465f17412bfb15dfaaa2cc7be6d7f8859fa6eefafd0d8f7a89cee60f
z25e928b3d1237d9920d4249be298569ff3f3ab460ec059ae7bd712c7375fe88379813e2fb7600d
z661d3dbcb7029818f467e78f1b9361be17f2c83186029b642067a84eb20f3b607f4360255ee00e
z3d4af6cd691bbc29d86bd4ec866f8e63312eee37004183984ae6ddeee15600bf2e2c38ebcf4679
z1840f1c2b4774dfcbd0c9449d7b21dd359947bbdb8ef2e178465505d82bf4af86501394d655fbc
zccd829a13227cda5a9bb216953733b4086dcfa65f0834ee0b0ad2572448786df99ae924b20cb53
z368023668de9dbc714bc6cde08cbe3cf18aa00168da1774ebb265c691504ce466e29b8945b4924
ze78702eb6de65c1d0e88fb8a20f99cc0ad42ecbdbf122ee8e4e5c880ca520cad983c337133afcb
z1e7125efb8235b059fa66f716fce1e767dc6e3b625bdf07fa35043f9c9a1cbe964ec491a8633fa
z1d8fd154ab7f3bb15c687568a96e669da1b4d86e1fe0f418af83c3b44dcec004a8d9cc60326953
z51c3037c71bd1f3ce1990bacf85cad8659822a267f9d4d2c297f1a2a9ac19cae51fdf01ce35e8d
za0551ebe693f90430f95369c4fa421c7c648481dcd5496981815d5936d64e8c218c1ea12f15b91
zfce2b65de52ea65f756d17e3138115e287436664883ecdc8bc17b44c5a1c3e2fe1074a1b9018e1
z64804aa5c0b699baf8a4c10bd763addd200e519f8b891e502db63c7df29f5e194a16e787fd803b
zd598d89b7b9adb7c41e0977616dd9303bee266b0fd29a0949b37fcd7253a3de23f648ee16bc3d3
z8c322da3fbfd84938bf5e3d84448cea37ee1d2f9344a5e1f2646652b7d939f740719a46b704e7b
z7e0356d500668738f1a3542144d08f44626b26b0da867bd09ba8436b9dcf974e55e871be074fc9
z8dd5086537f97f589b5f84a4bb7ec731c39809ffd0d1a3592899dd8d08686d83458082b06dfe57
z3b074ab73c7471d07e345761dd203d77225d4fd6077bb2c0fa7ed672d7aa9b6568f14f46a5e768
z86984e9e3d1cc8bd6a40023434eef6e7c5da7c0d4de2f410ed56d6492b89926b609b22b0a4cf49
zd8c4ac7008e249f13e6a26e99d1f607ef82cbc6f8a89521696bb62ef67a9822967a66f04df0fe4
z30c1f02bde0e64318c7688467658e2e9bd8f414ef7465e2d0db93693def827b37ef1c2c8e44e57
z51d1480cd12330311a3146a4488a70617fb12f470e055b9b6beab7cd9147bb390c639f7181a0e0
z825d963a792a5aed41277575e62df4e666962dbabca45bca45758c47b3ee5fc24c131d9a6d9aa2
zc19a352771498139837fc2e0835e1e56935bf81e71d75fc2777e1535882d7d87d2ebe339cb7135
zc6120752bb670d2c62d02a29a708f42e20e33b5a0d30e54761d57f7fa2e8f67d02568ab3ce4fbc
zf9dfd975dd1e4c25ba8e53ec515b5467835bd5be3c8e80629f343072b155ffd537a336489db44d
z977d7323cd9572158de9623b259394374f43870b5bde257d29b68238c6d464b48f6a10192a7e67
zced3cc60e2a3d19a9254b1ae5397593480c27723d702a1eb29421b3548fa2b98142ca8d15a68ca
za62e2e4abd320db4c8b11176e9de348df6c281ce741b1f631e785bffc408278734da58db9d9deb
z4f4bd853f24db68a9bdbe8709b5688a31e91e5714b70a463524b991b61b3063ac29dacefc2eb83
zea2ad7077af10e97bdf924753f607b8f83b5af11e9df7a2bb19327710c4ddce129d3b9422f62cd
z27c7f0050237872f90d860177aa1af52756e14c457e818d6f53143a7b55307704b1991d222c7ee
z9c013d8caa89027cb33fcf4254b9e94d442d0eabc47344623a7ef35879927736721605e3e12ce1
zbc76335df3fad33a2fe8f39cd3353c33b3b9c9385f3c1bc3cb1620670dee9424df0a031fef2b93
z890c5ba3d669c64a0d541b8fd42d815004a1f8923741971b8ffa34af91ff5a233c59768b222f11
z433d6584e98c8b6e5606631d9ade461e1c0c62298c485de460a6e2dc03ae25701b8f79425aa261
za5fb9579fcfbc1fcb9a168798afbca2c2010c5e02655d1e0828a85ab33cb6e3efc2acfcb613360
z7e6bf83e985cc6fdfbef98bc8ceccedb742d358e267aa6d39143bdc2d29f0baa4d5637b71eabd1
zcab650fd54c14208fc0313d5cc46d06386e94a62b8f610eeeb0d780f1aa02aa2dadea54ea6116f
z8bd89758d463d75def1aa7ff55c9f9b3417c79a03eb7998cb6a17928403de80f475b7a4eb2fab4
z356b1a42cb2c48cf7611d11bde552750abd1eb2e4d010ea3cf17d9114aeafc775b4dc6891d269b
zd43e2d7b148bdc5728161133aee4f4defeb3022ddfa662052adb57b35087a58f0bc5dd37228534
z9e74bb2c15ef30ee2f5a2256a51746bec5e623c29e2f754bebe3da610cfe953b86adfc016b725f
zd91dac4aeff884c631369ed643ca4bfefcc7e3a2990f37ab3cf677edf4fea180f5f88bfdaae7d7
zf9478591409af8d288ef48901fa44c6d5c6fdbb0aa0397db40c892137f4c8a4f17eab58620bd5c
z2b59c84b5fc1bf2f1ed5cbc1ae6ffa29771e50fd346307d53ecdac9746195bb8bd7a273e66a622
z1ab039d20a7c9509fdcb4403a7215a405158730bc68cdd4bd7c09b01f7836a4eba23d7f4ae8ef8
zad3b915ea5f3bee0a4fc21bf4f4665dc7c6b64dbb2c5868a07d9bbe5775d82c35891f164ab0680
ze29fa01e2dabc037df8ced6feed53e690099ce4c655951c8b487fbbc484ed90c0c06f13b833ee6
ze0d9d81c7be3174fadc498e245042648d70e30e99275311b2ea1dcce8c9fa7ba0a8d1030c9889b
z52d86accbe7d1982684921783620e955e0520fb13864f8c054f57e34ddcd4c7380b84ae856a01c
z29681a1255db70f58592c6d9e0bb2b5fe2e324a2c4e2fa9c5ac9b985e5944c1a2a352a769cd75b
z67cde300de7a3999b92c0d78202618342eaec84fcf13e73c1075711a50f16bf01629543b2ec9da
z51fcaddc5b1e717abb6818a633038f9737c2f056fbe19a479b8de32411990e85a68986b33234f8
z300a2851e94329e2a22060b1f451688083ee3820780cb57375e855ef619d17e7845340e4ea8cca
z5d8c069ed88d8789cc95ce2711b15966d6e6f2cc724218ad41d2acb94c91004cfdb1a7b9ec72ca
zc35e718b3ad689a8739543b67f1e5f0cb85ffa144f069b35e653839374f0681b3f4ee31f21db0b
z9c792759de0b0d9a8be5f6f39e843f1ae04279b749fb9e49a73bb944b679447aa898d25dd2ca4c
zc68ab6ad24b873dfd2a3eceadcf9d9b533be1133887aab459c0aaa587d1a0254dd5c1cb2d55ba7
za8cf29e517c8c4615bd45c8a1bc51342a6e3f594f888a274b6136177b94b42a6f27a7f83d74fa3
z4864a13886d3cd12e46cfd3cc5beb1e28615fadba366bbaa32badf2600abf5dead68af9c2490af
z30b178efb1e7253a1f2df12bf873efe120566788f920fb3387577a5c62bcbb7540ebac6154e7ff
z177b889c506d565db892fc7fc707fdefbeb4f21d048f8d85e044d14310d08563713ee0043d0d4f
z3dc240272480d6b333949760661427b9497253ec0f764212dcfb28bd2bd86c1819469f555cbccd
zac8cb0e80653a2a37463df866cb4828e6b30d982fd08a29024086465bedf8b80262ac9c9504858
z76286acd64ed0868ee85484e461a1a97d445152d1a0ab3d40a81d01cbf64b15d4d21823fb70e8e
z961d529dfd7f23218e68c58672442c3e472ab4c577bed66397f1c7d267c6f2d02fe0ef06ee9c26
z4d2daf8ca6c142c33747e0d0feaa5cff1747ca98e29f3747f5bf70105e7dd3952c796eb3680fb8
z17d9f3bdad404d419bf880f4e6266818810aec86d296444fb968813a494b3797dbeec8a0583dfc
zf2d1b1e76ec72384aa9dfb318594c22e133ad2b679af7079c0ded29c2322a19712e8d9abd45ba6
z1543105c40d42ee36c624f32f86be925c3a3230ba6ef876f8764173c09da024782d8c41d9efd46
zc4c44b2e9d02ac085c637c16c6673a8110b413dfb682a9fad6345515afcab71df7c2c418ef9f23
zbbee6b14f267e4327c55d398e2f8c4962eb1840d5fb5ad95ce436d85ee9f6e8f8998cab7dca1af
z7ebbf0d14e19ce68beda0475ad45081e37adb7167876e6adb8bed41b39184a51df2b8ccdb1c4f8
zebd82b26f894163186dc1d91818b76e64a93b42d11709eadb4f335c438ae0b7d59db27d72a4e7b
z8280c63b332052fccb6148b53a815a12888810c0597af9d23408f308e262e0189888de933d25fc
z4ee9ceff5e174ca28e21088857fb924311f4bebb7362d355f05999f4b143bd58bb9fb4f7a4df95
z8ffc48f53d57cfd42fe3d77d363957fb55d20873f3a247bdc207e01d0e723c7ae231c538c86afc
z02033d1526b27c1302215ea8c47d9bdf5b79fd13accc60d81125e3d2ae23f0fdc95ea87029c751
z70f65dff1625766ec96a3636ce0695d3e0ec75ea67e035f9d831b83709e004bd04e0453936aeaa
z2070ec8eb131f75ad06dfeed8505ee9b651d9d9521166d38f6dce866a2a948d5e330cda5161c51
z94fb731ea6da1901f6cba097933631c10a51e91187336d2108cbe2985e5bda9d0e57fd557a087b
ze0512b937ca5d0cd1a150d07488e3513c4bbccc8318786ab754b3d2811d3b71353a6c83d3f3154
z8ed30a565e35cfecf4e43061182d9d49450e6e2053492445ac15bd754c50aebf6ef9c9c95a7dba
z05f6b87c866b986a146d5dc9d6167df5fc2e376ec28e6aac6a77ed60d81827855b10a400905f3f
zc85073f3d50702ddd84cd3a58e2fe2deccc6be7c6437b26651b4ca5082e3d2d3fdbbfae67df631
z01a783f3d41171fa7c685e685ce9bbc48dc30265345b013b759efc5c0b40df4f2cbf4ce5706d51
z71ed1b59c99f4a6eb3ae0a2e46a305c656f58fbec2fd6a59dbf3135ec0cfb02b89e56eccd5e9a5
z4e1fd3722d2324fc9a9dee4128c8f3e8670c949658610e436387ef651aab3274b22a21d3005f50
z17866aaafb96fddac5442383b685f61f9d16c933fc5fce687b94038036ed4db5e1a704b08323ef
z8d1b44465a1b685dba83c6e6d975adf5c5315c777fc673ae5d89264c2dc2dc663d3a81e0b6f1ef
z2bab43f750269c37ef10fd2298de3c2994ebbfca1108ea1118e3346543b2d9121125c8c82d3b5e
z3baf9562477b13797f7f93e03ac073d4941afe3342fefaccbce7ab30ed813b8bac285f5838f1b9
zaf27aca3bb8111f427029a7fc9f59e7e3ddd4b7845b63dffe54574fc9621bb766a01cc8c4839f6
z546510b3a37bdedd6ceaa388f71a490cf6ef956c05bbdcb27f26c4be2faf06fe7a2c6bbf50331d
ze4951bfa15c22ec2165a02ee66f741cadd780342f52a99be11cc48386a8a54c6b2d2bc0cdf71f0
za574611d066d162e1e22d955d7956d365100a2eed9720e1f98d2ccbcbea1cfd037a9d8b01dc125
zd588dba2d2ba4a1cd39e11d4bbccdbabf6a80a7c97553c7d243917b8c72bde08e72cac163f20a7
zfe39142fafa8402d39e808a874fc9dfd3a7c62a76cfd98d8022ff74527282961cb3d900da5353a
z48d0d70e511f55016eb9cf61cad15c64f2ce750af40908602d3de4664af984eff6c79edad45c91
z3c50fef86a4d030c681c633834040bb83833616ea773b992f87b55c1c39c6c2fad7b96dfc722cf
z13d09c1606dd08d67394c6fac5468fc475b8fffd603086d8cadbd0f7c78562aea73ae30a09b023
z237c19ed46bb1cbf0125dc2198d980cd183542778e15739ed51bd78b2e9d9b52ac37cce977f432
z813cad006d27a5143ed2e54dc29ba62b915bb68f1dd6402f5ff1fc6cbd8fa7d7ba94c8aca09154
zb8e313117a6a6630570a48fe9e8823f291d2122a178529f47a54c2dd17a662bb7f00f256f8e09e
z8a654a99a7e34bfc6e08febe7f4ee2882b9c3cf544f85d1f283b15aabca653d5ddfde84a39bff4
z3a3cbf6e36e6e80399fb6cd89719680792a3db04dc27da75b3288c63651e0db7f962bce345131c
z12bc21b050de6278a99590fdb715281e32258e37586d34d136c39398919098a81d17007a410ab7
zfd210d37d42abb2e29d9f86f0253daf6e4ce173db53ce565910091fa7a32f8a42db958c997317a
z47f7ffed966660025040be6710f66aa9d7ea8b8ccf60142c80b32c5a826f55b2b88e95bf077e84
z773e993b9b96cc1dacabcd649e60edbb8483abb51a9289c7446072097872bbaf15227dfd99e71b
z68dfc6efc96d79f87e6708a57a77ba1917ee8cf8445ce99a72ab04a26f3ecb12db7469caed85d7
z274205d690a2ea24de6c6b0287259bf244a1a1aeba044799ae6edc281acce37913540f36157805
zccba1d8a92fd397366e667a8eb91b5028cd25a1ea64670b334255c5f3e463e9f9ef2b739b96ff5
z697378616180d5ecd40e06d000376d7e85f20f80b88e6b785d0d8d189e1fa5063193696cc6f3a3
zed545892ca5f9f316a84b6d1577ff2f6cf442129d3f4e8f972f09aadb7cd2604b69ac4cbead230
ze3cb9068c36e5d6f4108bfc4ca65ff7ca1aefc1a5e1c0197af68c0400b1e68fa5c646d59230f38
z11fdcb5194da5e73ce02a0dbf8c4edf85fc1646f807946eb78cafcca4697153a5f850a3670a681
zd04dcdba1250cbb429d887c94e0c179e59383d685fc9445fabce6aba7d3e627b2df4534a25b244
z86cb26bd2ed59934723eb1f621c4dce4539ced60ca95503727139c2beed61b74b97d8e07765c9e
z346b84e423f2be173a6fadf702d3467ec630546bba838ab62743f1b1cf02abfdaea89c86692c0d
z6732eb6b15d810964fedc379c67616ef42203b5ab3d9c198817244068f40a7080db986cec67a74
zc535e6893e2b3e7cdaf8188f2ff3439e6b4ff96cf1ea5be81332a4d059781f53933a9474915d04
z98355f04fea46d8cfa148b4de544d7ee38ae4301c1de95fcb4c83e80833895a28743a588bbb062
z19122935da6b5bad0142493bfaa248fcb977e9a445173990a9c22c5bfd88b9d78650f14d303398
zd188352bf0b1623597ec00d56defd5866b616e59afb7ca0704615a3e01520f8b6668590014d41d
zba813446d10ba9f3e206bfbc77f5aa89ab920f0c07db19260b7d97f62f5f70c769c9523ca6f1b2
zac350a875e7a3690137fd01a16193964204136e638112426ebb7238d9cbce422c7645bd93ce059
z2ce3468820f737314f7c49ce1197909f5175dd0508480def8553b3c7ec35e3143ca99af83bf778
z75408e9145de47616a31c5b9d51231c060c38db1de8a98f92600debc671e40262e81adeebc5811
zf7feb0e57be303d6a9995300dd7558be57bfcc8547ff03d2cc2b3fa5b73b080849449191947e6f
z603f26a08989befa67775e33a9ab0c04c5550d4f638575569bc566fd0ceaa13c2b375572399115
ze02b2a04a36b5f371a92f78cf74a75023d173b6b1750887d055d157e8f32caaef102d0c9dc97a6
z7479eeb8a054cf61e64bb6e6bb779adb419d85a1195eb729096341c9096d3d291bd1eee7d5dbf5
zd416ce4ac64341b9e99c4ffbe4cd537e94e43741ac4eec4418de168107bd3d061c3a938c2b34e7
z6b0f3daa0edd000cbd18f546f6e51781a7c41ed4bbd2456b14305519cb4cce03f4edd7febad6b1
zc1031dd1fabb854f489b0ae5b6325b125ddd30cec6b671c3bd29a62ad319befbfc3c0f3da28c94
z1cb02bb74cf8518b988ff50d2510fbec3e2b31ebeda6aa42372b79f6a49369daf81d8c9b46222c
z8fd3ac31502efb865ebb0f2b3609e82aac25f4e9f81f0243a420c73f1dffa1ebd05398c6c777b7
z8d082a989c85469671370dd03523512a5c5119639f18c8c862f358ae30b9f9f83bfca7b755c26d
z8c4b2fa44ffca22744a4413d0607541f23f5564fe9738d12491f95f5286636aa67dc9b60cb8ea2
z6f8602c3ad9683e91c3ed313e6b0680def9194d10226cc331bec1e4ed53558742f8fc984978c71
zecd65a21d8a0e4983b877f2121794d02cb4a7e0252984890cf0d6d92e9f50ab3ab7a3ffffeecdd
z23202b468d9afa6b639c158ee3c2bfc18b3713c89a98eee18739806514fd48d68604ec6ac3f56e
zadfb7a112f97853dbdd68a69373aabcb1391976a9098bdff8108ef36deb67ed2044f82ec56a37a
z1f1bbd19d06b28be40f7f2fdbd9c21810e49c0c55093992a86a0c9ccc91408cfbc0eb9a698e4ee
z48e04833ce84b46d45ebb69838b6e7a97a32e85ff96222841b419d6e69245b0c015d0cc85ca9a9
z5759e13ce2881be481b544e7d0c9380752bae79d33305b221c50115686eb673c78750085b50374
z711858cc917249b05d69e9d9a81c8f4d7829fbe720d4c3156ab9dcf0582717c20b4c69f674a418
z9ab7871558f3b9db7a6a34a47547de85935bbf88367d9ef731b33243a029d14d888edcb5fb260a
zdf2356cdb71d31c677a1cd020f208d52f92d7fffc671c9b51ef967ab0953338472a479cbf82b13
zca6d113fbd4648f16c3b89dd71839016d098c03c31f6ae6af6ac1351f8dcd251dafcfd182a50d6
z9b2b76a70b6836ad6519f67e0bec1e6aecb5f90f43a118a2e9b4c4eddeb15879603b3f58ea18c1
z809c7880c424f2493e294e9d5492fa6785f9c9b1caf709b8f09412a98bb06ce43e063bd00411ab
z3bf3597912a81b5b2efba5018f7543324be9992403db825ad35523d7c8dc9bff9606dadb9d00c8
z07698deac3b02c216ffbd0293b6679ff7cde48ab04cacf1cf332a1684bc25704ba1e095325287a
z9ce6f50d4eaf8f3f3aa7c416dd742df7494d92fd3a1993d445bd5062b0483f987276e09939e1c0
z4fefcc1cb3d9e9413d230b5b434d932adab5e4c810d55f7946b2789dc6ef6776bde544cdc1f86b
z7b3f6d99454d80f653939e1e6dec10c47f3065008db4de59e69acea031754dcd95e0a084559bbe
zdcda3dbc6a18472ee0736be13cb795049b99cb36b05124b6bc3c07dfc70f9255d7b331da6602bf
z3f0e19041c80c34733df3ec91be6975dfbc1daf69f81f26f213a6a1b8fc254649e130edbfd7d8a
z17b9ee930330d6bc9c22aaa34d6f988a1705a4fcc72f42cab28078c277a467cb4c6e37aadb0c55
z080dcc8b4e03033afbd27fd96f1dc2c5a35d0f02947a5bf66e56c2de9bc8b7a5aad1b3f2869b05
z41cc99071b9a5ebc18709fc567bd8acea9a4a94c285af9bb79b781523eab68b2eb4b8aa1db5e8a
z146ba1393ae9732e2b6b66bb7a980f80ca3e4bd64da7a28dcfd359690cb5a339fbb31b78fb3598
za9fc8d0576a63398b3ebc5624d86f78cc2b89a3157095cce88627940064665ce0deef7f2624f5c
z2dc8a03b34afba07a3358c260f7a0b9dac0e8065b3408c511eab1f9f0f2a578fa721e10247818f
z5caecd232c87154012e13ee2ec347b348910e85da11ac78f9c7cdbe807e7d451890264411dc027
z41410c15c617a10e65c47470faad54a4284d9b330d771f2a3b6ddc4543aa8da12a6a9e44325102
z15dce33a6b83029e1de7db06ca1c0c7de8912303dff3c3e3e6c0db749506558af94991ccbd5523
z3a2973cb54d1a18a8457d05d562cdbe85c43315b97bdf2faaf29cf7534bfca29351fc65e25d98a
z68a0db85c3ac8549a96fd7d0da1f6ad6b3064573127a943b73e71db632f3f0f21f400164a2fa9b
zc4e1761134556ece2b24ee7abc4d22fd5b46cfb54781a8089b43f1268f0fcde79f22a0c3765231
z4e69986896520b623ffde4399ad3ccdcabc04ac949088d036438ba7cc3b40383eace965499af19
zf81030ca0c11a5dd0f988c14d1f26a331430ae23e68d27a20086008c070a92aac35fd99583a513
zabf00234fd4814adeaaffe24c45796e2cf53169faac54c1c0c4dd1f4dc9640a867eaffad64803c
zc93f199b4f25e83a1d260399376a009002142c738694ffa149a3c7659a1e0df824abd2ce5f83d3
z49f133a58c4354a163a657bb14550806c8b997f9ea093a4c335cb74382e08c3b836b23dbd2ce2b
z49b0c006a5ab6f3910eb14b27794d5143d778f74e2e754c3f44074a0feac1271bd679a9f76febd
z6748ca57ad03ae664cfba2b0457c5804caf1bc84bed9ea9a784543c548b5841ae8b287445a672a
zb05ff51d5dd439d939a8149a00f36318ebbb4917be1017d685c4fc0fa283046f85596a91c8d0ce
z41974af4ac797f5da173a87bdfb92bbbd1e5f020b25649f19e82ee1fe5a6658a670a133e0edb48
zdda5892e08dd3b9d6bffd43613a4e69ffb638ac747d74ddb98bdeeed869729367a87a3e133c7ca
zdee35890d14419579a339cf1fc2cfb5af45b770540a8aa8875e0e4854a89572969cd45af61f72f
z69ef9c8be7447973846daabe5a46527c540131db865cd2eb9b37e0acd0e50b0fa15a033d9fc486
z86e8b80c3a17dcca2b9b5afbf945965a11f479a2460418a1a373198d5d221b1e506e87d7255cb8
z90380881bc42860cf16f7713cbaf3da58f6cab9b12809db8a0cad44e5e9b2a2eb238b88fbce50e
zab5d78cd01c846b12d113b53757f13d03253cf8f3271a01af9add37cb45244a30898a24dae0290
z2e71bf89182817b2e1252914abe08e6f7bdffed3761ae89863557d992b6df523b6f3077fb2a9ca
z6d5f402e6f02504cabb99c7675f71b069adc356e995f0ad1c9dfe4e2334d159634f370174584e5
z676e6ca5954363f810ea7f71a834e256fe3c18cca95cfb54d26fd9134ed1058d5e8f6abc2d44c8
zff8dfb393882ec5e3bb9cf716350906045ed6f29da8fb037ced80e5f3be9db07fbbd167b9164cd
zd79dc12a3565abdfd3de8ed867fda5292f1f747f35d7ea25e7194c01838541ae3309ea1f11847c
z37756e39a5e5fa8f5cbc65cd7589a519982d5ed8163ed2dee9c4f58a2504d1a772faaaf641b296
z1b6c9490479e18a8d5873eac8265427a540f9766c4febd704cb1c7f32f96c9dd257c0e21f3a672
z3c4ef39fd2536fd25b371dff089bafbcc8f79aef00bc82f9ed46c815a23c440b9fb041dc8123fd
z0fc67610aa25ce706b80f036ef123868c543a0a85d591babe38d5aa9243ecd41e0cdc6bec045c7
z34e9978066abedc2984a4f28805cd24b91e03fedc930d32ebb55bdce91140757043cccae265420
z32f19db3b36ecf8d8ddd31839e5e446c618ce548bb6aa9991a37de56bd2efd4b14ca0b99281a03
z58d159a4aa3defdfd5d286c5fd268f43c44f136c9c95f2014fed1c1d5bc723d362a5e887cd16e2
z6243da7978a580a0ca4f145acda449b1248664116a9f035612d80f9ad646a8e47b915216e85707
z5d35079896ae0e3917f5a112ecfe394ae981c774d95e1c5992ef6a5d1cdb953aba632cc998c4a2
zcf0177362389cf2d06622bb5a8c7f89af0c6683a2d7b8882667166ee37b6e2d062c182073c315b
z0cd5871d459e12b7f2f180461754f74a7deb283e81a69e65d4742e1a4f37b86fd1418bacc08b1f
z35005ba21dd926d6df3ba782cd9a230fad79ddc6a5c24d6c1c470634f50ea24dc22a7fa8fb31f5
zca4aae7ff3426944bdd4555b7670aaa43e6f6905da13c800e1c58b6df9b972648b793455751e4e
zeedcc7620f7626746a2bb6f5170909e8f6991a3732ec1fd4839a843a6e2d5a6764f8b2ad0b17a0
z3a935655c7e2f17acdbb06d525549c0e318633af757712ce99b0cb99df98406d112a354100871d
z490b074b9a411f10aa753014b75ae45fc70ef148cacbf5d4e5e43057a04d1ce55fa000c0d9e559
z2919919d3412f3c6617f7dc00972c9917f123359a71ecbb31a9cbe4ec73ff8bde75b854b8ae0f8
z3bff1d9be35bd5105f02ee2dcc7dad389e6e958b4c48c1ae08665ce425c0a663c093e30fdca626
z67b3e8d7d1beb16243cf94bff723f330b87f1fc175136adbed15e0e3ff7e4eaedf31611e42dedf
zd362b87aa633e333d56ebb70c2bc988c34d5524f2144ed471ed1a0215e11b13b0f4c6a5caecac0
z567775b37faf57d1c5323ed1d40a3413924e7bb9060d0fcf6d8b850f372ed5c49a640a3f6677d9
z23412a6a4be492b162342a1efbf3111eea617321a73baef0f84ebf7ab046642a90f16ea71dfd59
z29ad314c0c66e9004899e93cc5db26eb5299de1a00cfb1a4eeebaa4d2bd25109d669c2b6f00777
z857778ac7f02ac9a4fc017aff233ef5e2018c885ec8b3798ef5c92d5e52bd4afea44649054c0a9
za4238a1ab3d830282e39fc35cd532000af9c0652275d08f05cee2c345525a7410e14a93cc6614f
z48ff065b2655b7e587a37c6763f8e5d24e9fa5f895846baffa779ee100b5adcaf1939237965c07
z907165b9b9b400eb2d9f7107e796b55af365aacbed897fb60c6e1d39fe23c101c06007959946f9
z790f0ba5726e77f39f15a28d168c8086fd51f74f9ee401b147e1cad53963ae487326cf2ce2e033
z5dec495e8bbc5048493347b80852b5b798b349a18f34a98920712966f082157eff6b4259c0563b
z098c5d078281989503964068fa09aa3343f35877ec995c414c4607b70bf7931f6f7711e425c488
z9b54edddd20f2c8bc3634e9cb40b958f95d574696e73282ad711c87202e9fb149adfb150fb9276
za2141d1499aa79f1b5544f7f096857d8c7965668b7dfe8419dbaf5fa7059bf8a204ee2284df4c8
z7a049af24faee5c387c1a71c38a8efd9d0e0ef096ef3a0dcf7d34c4b9e11dff7ded34493dd55e5
zd702977a44eeeaee10190b3b244722b1794bdcbc1dadaf210d316b2ed241acb7cdc13bbc05aedd
zb8f35068db5b1938c04709b7172f0a37fb9de4e52c41c30c5e04c9738f984fae417cbda375db78
zfdca4ec5506de2a5b84ea2a1470cd0077faa17c2467093bf3953d371b8e42f61c8f1563175e587
z95b8da13b585d0483735bac43273c8fd1e7612900a28ea1f91bdcfa6c5e567254775fd81ae73b1
zc6e23f40c48bede370ebbedc7686a57e9779d1d87d2d5a7044f94fffd68cde6756280b1140bc17
z496001873dcde9ca9d77cbaa5adaed3be39ff005d3a111a0eaf8a8d4f89d1e20c475a2f2dcd614
z10d80baaac6120ba52d857de84f33ba97ae5ddab245bf1c10ecd7efce0efab70c98ec6b7b45c9e
zec967112d51674b0e2a47f4214493e5f1c81dabb0e193859a8a294c88c0c255bb647213815a8de
z71b7c8232f99191b144df77d4ae8ee0061976c7b44d37e3f90cb04218566a6d2f358e8170ec924
z6b8b34a6171ccfc597757a5a9f1297b139509100ac5391e2142437287a61bab9ad5f8349041d18
z9f8911700046722aee9660429a926409e7b0c755522f1c79ffb1abed8280f8fe7afa144345b6cd
z25a9f3c309842de2068143e69c2e7d0a4d0882075c1423c03d77c9ffedca722dd672047682ee4d
zc73baaacde5cd5e9e08b95b3d9ddb412e814c70ce88e42c0076b5e7ddf9381cc40dbd55454ca67
z51a7d7bbd87f670c0c03febc0675b96a8e3ca01409c9a4bfcd33457fa33ea1fb41d6c210cb4093
z1d28c3708e1ccce08409d726a1dba259da06c66d5ee65fa0d0a3195439182f95eb7b02574a9f80
z8e523a7540f7b9097752954482276632176f6858d7d11c0f37cfbc7e699ba30b66415f402336dd
z97d2c992b4c1805be04be84032a694e73bca6956207760066e69413d18a86f0ff14d80e8099769
zdf982bcc722986fd2181a0011b9d7795d4a0c4c60fecaef69b1d8d5f24512a85b07c2be1024755
z0edc87d04809f97f0c3ac230c8fc58eccb192b3a488e6df41ecd289de00f5c6246b371f792f141
z4317df1f691f62e1a5e0a37a57db1494ea8311e30c958ba684c886d021ced617fd09763c9fa47e
zf9ddaa74785a2335093e3e0c2a9c31c7e2bde0c4c5e27454225d8bb1aa651c1b5f2fe0d28e09ec
ze2793cede830fd6d3d133df9e88136ebe42375847e9aba47f1f9ca12447174374e33f6da24dd4d
ze1622dd5b284f0e56935f294e47f7333f2aa77a7f8f56f54a5565e894d905f7b0c5141910e25f6
z31b4e3e6a885279834e8b3e7611b2c7ef75a8859ac98f682e8cc6de09605c673b49e073d698260
zbb56f5428dc661d085256ec59c09686825baee59f7d97aa4fdc5cc9d174a65073ef5593984e430
za0fa31bf51fffbd7a82f84e62c671704faa25a9dd55ef319dc17d6ea4b423da59359d05b606a46
z22ff132aae61f821377f6083e7b4b2354c9bdd84db58e961e364573eac3a981777a7988225a8b4
zedc22b90beecd7faba0a3d253d56cd94e106818e683bb95f16d66da4400d2f2b3949c1f2ed5668
z4087627882e023d4e13a4c65d47eb3ada63eb5df5444d0c6a7873ea1bd9bed80cfbfe86ae59fd6
z8a19c4fdf05be3ef48c19e6deb89623aecf9e287352b44c17d9f49c9c8254e5e86fdc3b54390ce
ze2c8cfde051ff600463c96e20f2ae4936d9a6e07f8744fcf8d98304a16edb4719c075ae93e06ce
z382a05849a6c386d144a201e1532696f808fcdf6626634cb942c3bc5c3053b2bf6dcd82d748b9b
z17ae3de11a3d5c09162cf51f137e5e1bd0d43e730c76a90d48926ac5e872592e1a713d96d9e185
zbf2999efceaeec79518dfc6630839b429918df82b7fa5ede407acd0fc7237f58508c82a743850a
z86acaa62c3d1d72b58cb3600206837fda7a27ffb75f63119a5f71197425acfb3b4f9343ea052da
z2839267c0d6b52d2eaf9cd0a02b50899ae439d264f93dc9635f25adc8f8918099a2bb0e8ca5412
z5b4e3675e274c45720c358f0b1639ed80a5d4b6a914eb605b9c35ac96fb80bf90777120fce605d
ze96dd0d9695c31a4c3dc74c06a79c34d26416414b0243aa70a5f91ea7684f68272658ff78e454d
z25c63f295d55f21f860c1c4a357c9e20ca2a684f458bf3c9737f5e833b13011b9f8f44a24d9c01
zc90347d366885ad535fc6d84c350d90b8477103f49dcf0b9d99f007150b3d6cf992cf94d8e1e92
z393393ab6f723be6d4b287d8248a694bc96860cd7f2d500c59bb269406e309e21581e2ab770861
z243dd808be9f0691d1d47a7195fe7ffd0522e27d98345ccb51aaf39fb6206cf9bd4ea2d3d523b5
z789aacad55590063de3cb93aca2de9f8a494521fa6ea356c310c4bf3da5f4c794df93f7c0813a1
z0a71ac50e1f032f02cc89be616f4984008fb104cc2a7f19ebc6f0bb34b2f482e13dd36da08926f
za966b2d4e4e878393d7fdc577bee37f3f95f9a0f459a32fff6a7e9544010971ece300bb3a34b29
z3a60f04f53914a61c6476b88c92988981177536a543353a63f17b2ca9c22028eeabe385cde62b2
zfb74759ca19ac0b3f393c75c44cc57417aa1aa02491b46a71353e498abae368e75fbc2415745e4
z5929b9f653fc1f79f851fdf3758a6dbfb5c03ef84203f6fbcaae1c0622ef568531d8b62cadee3a
za4c95100194c35d17175abf4a2c2f01dc9efd8942422b1cf594358760a4423008cab8ebf1c4986
z26b17704d6d1ad4213db76b909b143d490c8660e9e74bae0d5182e86f3b3f7b9e16b50c083382f
z5fb2b294f2748b6c64e6c142661a8671036d21f58410096a1bb2282cc57c095743fa42667e11b8
z27b95d637a65cb45929b88c47646f8234a1875899a3ad184b5848d07b18364ea02bc6fcd5202f5
z17fb7c90d0aab232e843aa2ec5bf270f244fc20f0365d26f3cc973fbee24b1002276129bb3c237
z8ea641b418e9c922223a482064062050c95a2e53b19a6c6fe4dde37e7e9a61f1eddd0531a61f3f
z202dcec0932261c70a73804992cae9af330f36ec81c454650c885bdeabbe19c315552051d4ceb1
zc7a4c35bf4cc9a8471bef945a2847d15f708d16d4d148245b1941bd3a6df7aa2c2413c4b7d1ce4
z61a37604ac671e48aac3873110c741861885778a41a55ba7822ace6d0ab9a02d35d99a2077078b
z98df065e20f786348571f9b5743037669a760b11611a7f315259d6fe7247497467112a4980389d
zc513d7e3ec7526aca7e23be688c4b6b05c0b297cc0dfd64d4c6c82f7477bab8b1f1b589f58f7d7
z6259fe6fea6e4feadd387435102580f480c17e4835c65fb03fd7140fef04ec5ae0565a6ac8e90c
z717dbaa985289e4532eee2f59cc64a10f853f36cd6e6bf6f5dc4384a0b7900c81b223b5c78d184
zc4d025d9f096a7065062adf785a706371b32f1783ada79e898cd04cef4ed349e1109489ff6cfe8
z90ae142e3c8e09b2738c6e0f485336b9cb2748a501ff4b5f41b67881038f3e3672b56c887b697f
zf408378887b399c0cffb6e1097d5991c654313e62d3b1d6f25d59c802b4fa891a4564effd2e47d
z1f24f3d025e9002b5426cc940c9ea20352ce6ca8e60478ca0b1fed752283f618e119ebc9b92342
z6955e6e2c15c3b4bfea17794026ab6d4cd6964e5720789a096e42d15c29523180ca1124fd82fef
z3bf19c804d35f2901864b59f9b89f349766679cef414ae355d983120fa84e1a35fd7163a8bd4e7
z686d21871220fe2d1dc7afd2acf9f1036d502c4db7f9def7f00d20bfe63d06fe52a9363f5d359c
z90da15dfc28fcce8a50c9ee812cf0030061b29c5fb8e1d9a468c86a7ec8dfbce298b3735530df3
z31873e3a4ed0ba46a040ac899e8f989661d708d9bc5e03e4013e2e980b4f36abaffb795551802c
zd2aca8273af049e13f853a4b47d65f7127de0b5762d0a39efe58eb389f29e2c98c54388c207ca3
za208c1c28c9f1434d618e5b350817f93cdc2f9701245540f01ecccd372943358d01ee630cd51ac
z3a8221b4b3a725d197f87b1562e0b4361967c965ebc30dc38aeaedd1815c352eed2d3cecb70902
z667dff73bb7870bb41c7ee164ffa0cc85341b355973893db62282782a6f992aa8002030fdf0a52
z80899b4a13c798b281a6eecdafd230caab2a193da1a9762b54c745c8ed96bd6d243b94dc5dc829
z5a362748c3d0b6ddeb9ae2db0c159898726fc924cde51ee0f69687d60b16a01b3f3219db007f5a
zf814a4dff99d68633cdab15ad31ea51075c02c5dac4aa95359c31964f4c1cee7c95ed3d2be4ee7
z7373d0fbe36ba1b3a6b040402cb4042ce41d4555d12d873a7e42bc39cad3286654ff3acccb0d16
z7c0aba252f215f8fe2350b0639748191fa7562312a642905a5edeffa9a307c112d973ddf9c02fd
zc3346e3770e558e35644f1a3691a489b792f68bec9b3f93465e7f1de75d8659672c5bf91b59322
z488b733391d08cfe9c4f19314d8908ea00914f620265678b183f1a7daa0ae29ce9cf3fdeeb4c94
z00344ccfad3c19800c6a3211e154ad21d1193caf93d94ed93c5e0ec08792d835506d5c302cb75a
z1dde67e38cab5e5c146d0a7480b685f7a7cfcbfc64a7236125e678a12219fb89e8344008bdcfa5
zd3abadaaa392e30fc47d65b6c9e5baecaab94e2f9144920aa38995e0ffa9a63182ca2b6528146d
z22225e06907cc08405cfb161b02ac446185ceba37ba971423e06c9565a10d780fed3c341cb9611
zbec4aa17d56c2a613d8fb7d0aa4cfa494462c5268f5fb8fb6708fde9e77db3221b4092148ef929
z6695086cdf3787f8d624a45108276faa5498d082b98c209716b12604825f078e28d8e180e43276
zda2138b5ef08deff948b95fb25e69226564ac42c793e24e965877e09046afffece35ec23143350
z794311856c78b8ccfa42ace83c3ad21fd3475e9daa75d8b6d8bd050edd5eb5b8c2ebe58c156b90
z0800e5adec3845e8272421e361cdfb2fe37bf537aac48ab7c8f12ecdd433779a2401a026fbdb93
zd50f3f73ba126a3589be28412311d5a91b680c9d852696f71d21613ae61b88958fdf892dafcdda
z8a20bd69df2cf465b40842e363cc1b6d4eedeb3ca4db03ab0d9189e9d9d07bdfba6f70c8ee6396
zc9fbac54fead7a7b8cf13841d3639c9a5138f2b82109a74c57f85b24515fb7df292db6225cc45f
za8503eaa3715d780bc01383a67983324ab0161ca97c1ca9024f3bed77b1b61af855a869eccda71
zd6704f84262526de0a583aa06d15018912cdc74c170cabad356901236da06bd3a76ca5b309c73c
zec74a742af7889553f890b8b90efb8fb1a32f99e76eca90a2fe0286ca5661593baf5d6a5deae14
z0e12e04bc3aa2acfcb88737fc26351e12415d85d22bc42eee5fb0ae7b3b02d67cb235e64aac91b
za1f45b2bc8f190faf91461c85e23a87030ce9ad8a8e9b3ed4ef25d6159b14251c2df5050aa0e6c
z4709cfe2d7e2a39e6ba190f9422e239b6839a8d0b1acab56f73f7fa0f51fc4d380a51091cdf0a9
z1f989b07a3a5db03dbd284e4c84626dfade4f7b98933df4c73584d29776e87ac6a00a7b7fc98bc
ze641bd2001b4533c24d09c3fb663254288ef1b07c418185a6b529de17284f1d247ded7fa5159d8
z48fa7d13fb5bc3c52d740a19a47de16aa5b47ac12ab5cbfc8139ab229743c652566e1323ab8f66
z565c45f1ce9fa8b78aca58ee8788f2707977f1329ff25361cb1548ae04a37f57c0669dc488d8e4
z379b4640985c3532b20ce97ab794403ec480d3cdc3c58b4042273b3d3052cce28b2cfb242d1771
z5005ce4c9bb570322cb90736a9acb58a75a38dbe467dbb74eb8645d682001fbd373be385c2632a
z17dabf9f5243049e31dae85454696d88f129a7fe2c29237e3a2ed954cae94dc385776a2107703d
z9b375f71242cff28860cc7012f710e2e7bdf3df88d257b1ca44a4edaf909ae9739095fdc43f667
z115473ccd17dd0583eeed851877af70b89a8c79d1abf66a6fa4ae7b5027701719c1778f626e65b
z8e698dba7c947d9b91f50e832c658649a833b72fec359e523df9aa20fe564795b3ff0ad875082f
zc010cbdb1b55c82c450b86ba0888c343f6f3831fca0465159957e8b7e7c4dc53761cf106747e2c
z7260e51c0e4f530bb2f5a171a8cd36e03b25ed003c694979b9b13c4dc8332020c4c145728d8b12
z2ff5f411546517af6b2b8e20cf32fca79a16cc9a0b708aad96c1b148f8f8f902114535a315c0af
z2c648b0fbb35fe5d47ba8c42f740af9bfc3fcc1f25a0aff3a65acc035fd690a88c638e91ef562a
zdbc31361da93d02ad4013263a4facea60f25e30bbd32fbb0bb5bd90611564c50aac02797c3577a
z3a6f70c55a7e207e8edd63ca03cda749485a3f0bf3d39291d234bf44a5b4ed0dbe5b4e247225e4
z223c473e007c8078a43c26f63867979f50d4e3af762effde511a1f7e85c4aa6a01b020788ff6fd
z81e45341a78f5cca11f9ff9501f018e62e7082021bd71948fac575ce0283dd5eb85ffc30d965d5
zfbef0a868dc23d0f355151afeb2dcf00c08df8389b05c34628345e2377727dd6bfcddaf772d4a3
z8b3b56c8f98780757f8a6f4c0d519f764a5d117324ba3e67eba8e486430b79641939a52401960d
zc5d9df1e5e04531b17f207c2d48964e714b93ae985db0d771ffc8161ff65db8da87a4ae859d088
z70973f8fa546be9753b65096670165494b504d9d782e6ca858b20b2803a755e7db6d3ad9ef456e
z825c925723e3a60fb48c6b073a23f0d7fd2c655fa94ea6e1ad0edbc036695844473f4311797ac2
ze1925e783d23acf2645d51299445a0036eb88d490d98ab5cc07f3c4e757f00a7e24b7255fd153c
z41fb4d9e8cb69f86dbd12681da39f6a679f3d2b9cd159c2ef4a607f42f7665a0b932c295894518
z7c2792cb57dca6e0360878be678e11a808e8fcf2f8e3256b6506d5f6c90144c7cd88595b483a6f
zb82c482f189ba7b46aac1d9a37558c30ebcd67a85ac87d9b34ad98fe5882c1f668ddeacb180d52
z769914e821045909990e54ff8d84aeb3ce56d900ac784faa91e69e00cf4a86542c2fc665bdcf6d
ze5ffe94d3352f94640f76a21b9f97022feb542d861dea1c4e4618f43c9e51abbd16c52263379ee
z1b37f47ed43b720630dee2d49a6673c2ee04cd52106af12f4f47267941a2ef97f9a1fffbd0c14d
z508e4f662dadf6817573b104820fa57164f20fce6a41a0be2ad868ae1bb9d34470d5c07214b4ff
z095660f2bb2affc0552fa9458dc0a947777cbf9c2b814fe0f6c2c13bfb52aba3bfff7772f3ddeb
z5677c02556e2e4c3fcba66908e52fceab4f3886d920f3d344808b961505431e0abe7e486d333c9
zf72304cf5ad86ad8a76193e77e0902b76d8f56678dcbaa3f861acd2241c301eef3456c800e8793
zcc05ec8913b7a14a03fbe2f094e740e94632937acedae064eebe2774ae3659f6feaf8a5fab1259
zb0defc5b0da3d86a6218894d84f5fbe6ebd93b995b79acc04ad6b0a66a5c3885da8d6dd2b3ec61
z3c4d27328e64a108270cead1ceb4daf9dc8b4cf05cacb55006959c19a15aabc21b90773e54efe0
za9e7d4e8222763ef9c4f62cc5e7c33be2f50bc986c8e8f55817f7ebfb43c96006b0cfbda132672
z88a7370010d8eb6de2888bb416a5df786931d5a060f90566b3a8adb1933fc259662e3f6d7b5c06
z4de90d59bb6c1ff2522bcca8eddae3526d60a1e750c3903ab40af321333855b8c1108a73bf1278
zcd2a7b803ae89fb1e97afdf4eca4932fa8beb391cafd560b82b4f3be39bd306ca748339761c87d
z798e15240e59f1833bf02e0d2c2533d0d1e68341f5694be16f1d8b96fbbba90cf2d4b6e94ed151
z9a0ff8e8562695ffacb334b475fea0d3e42e3d602b20aaaac2f711c6b30961b8e515f12082112c
z1a09914c5ebebde8e0515d26719876930d1b53c247c8c072dbc982bc191315f034d122c93d4b7c
zdb4053e9d9c820b4c79a8c17bdecfb2e4d153c0c618c6674b0ec12423b433874e03eb95b965bf1
z84df169ceedec925aa10a918a43a6c5e8ca3da6801a7378be5dacf5aff1b19762f12d77f713fc5
zbde2a024e1bc4c765f85b3a2f24c1fa26ef9d3ff5b421589a98dcef2a54fca97021acfe08c2d8f
z47dbfbf0a87afa1cb3c10f8e154814e5c93cccbc9f545a066da289ebb2da41d0bcaf7f423bb6a5
z36946e59ed17213b49f84948fd6dbf8d622c9ab00dbece1f00825f85c14f32bfb6c346ed1a550e
ze0d29b4be27df97d21d70dc238ad6d977e20eaf4fe79901e44239af50885fdf255ccc0fefc0285
z6e7c58dc1106391e0511d6abb0997e57968b630e1e74b28420b7099ba5832a2591b7ce53aea5ac
z38c828d41415aac93ec9ef395c67f19bde3bb46d60d30ddd1150b3bb1256f04c78d825ad76afc2
z22a7840737dfd659748587911b478fb45f4b485aaf9df182e855f8d0feb4d280b0597d18afce22
z92b694a1093365afb0fc0554017ad55e490cb0621b0a98abef949bf0dd48af2c06a607e41927d7
ze32316c0ca49443f6267d1e754a2f3dd8790a326fa25ac20a1a2b31e31f2ca29dbf8aa90f87560
z2e20b0a8449a823af456b0affd21b56279c64ac431274b642930bade1e191b59e09fac22711ea5
z949d5643b51727dc5406d10f569a7a30d44f01c58e98f9220469053800f90c115a8cddbc0354a7
z9a87596384d6614441bd5d331bf68513b5dbc578fa25ba0994fd726fee979fc3c4b8f996371416
z32df03fa51b2b26560e52ca686074a8c134392679001fc26bcbb92f4e64a34a2718a77a6c53f1a
z95d31bdb670c972428d6de1208c28c13942c3d654d5242f41f36fce6fc9eb6428848917c444a79
z5480fbb63a6e3ae7af898fae2c1fdc846bb6a6f44a4267252cfb9099312758fb26fa2c3129d84e
z6e79bc419980c23755c0ed9da1add1eb70bf7a9e3aa353fad6bfbce51559ed2f308f4522514193
zd71a3ed9a7f9493ae98a319d43ec72657d0f68dbab55acbc696f1c5ee7272f36415266a16e3163
z6439b532f68864241ac1624a76bbf75adc50349c380039d5d2d41916d7102db719501d8775ba49
zea9e1101b393428b8d6eceddcc4c8208f66b91ff0f7641bb5c217df99e7d1c7edc1df652fdd3ca
z14fd4e2676ae847024fcd461a195ad9e8b23286526294bbd22d933636759872ef55e5bdf9d6e1f
ze11ca47d72cbcdb1708f5eacce608c779c3d1b6ec96160ede796529073378a40e12e764428ca1b
z9497860b74a4eba83fa69cd1f741e6775935b894b3f0cfc5231bd14263432653aee4e7f1c105c7
zc9e9561f374c84c8ff99e8823441cc5e3f4f6d3cb0cd1f5cd708e9cf967a458396871589203e50
z4e52e1117620cb4a4a3f4772e3a13905609e4230f20f2305fa0c865ae0c9805e0d2ed3ea2c607e
z90b64bec5084f925e46878ea1e6135a58c2b9ed61bf3a37e234cc645cc092c2abc9e6bb370bc59
zc340bcbb3bc30473c4688072c960492fe3962df368de0eeab594f3781e4573c97b2930048b3d24
zabf26bc168b02289a10df77f6ccdf543e8ef7094659d69a69d45ee2e47eee8bb0fab1fb8fe3a4a
zf2862c22f4c6ae90130f61c639179141e877251c29671440bda57c543207da47de6e82fee49b10
z604455b4171f9c2167b4db10b0d6a0b08cb89473fa03a2e0b2d60da2f7b05e0800601bfb2cc3cc
z931d74ec491d7fbf81a352cab1f043b1d501813b3cde6ae30d7a7968981d0de7260e760251393c
z3e379941c5f0fc3d74ed6b61ba513c80f7d109eb281df6ade912b113051746deca3f69cc342bf4
zd2f5cee5ec7339fa8a5d4bb7d75974a4dc046201bf6e74fb6f22b5a69a51153d0ea93dd6f92984
z17028c70e7110e5aa8f776ed3df1942b0fdafbc6009f59cea28e668e0ae2d362061b0aed873e2e
zd7d801942718c8f6dd1e7a85979c79b897d12a4a8880320af68063d482b4887b1d81297a2d9ade
z75cae0b1e1409807e5a5f68eeaf253b5f98a6f336054a31d70d23404e0bc8023dceeda0319e698
z572826a45e335c8e122677868fa452a4b24110b5d5c71eb6521f408b6805b2e288ffb0d57fdcc7
z7712bdbc6948c9a755977a5bceeab3269989f7a8b7d2953fc35de177caa1d117db5a432002397e
ze7c49fb04c8cbdff30c6349bada78f0505c913b06b40b8a8da57eeb4e6d7c8ae13ed74a4cc20fa
zcda9002ad113447a0d249b5400eae2282502cbdff1d4e6a671bf74ed3ffe3893d6319dab67d150
zd5bbe8eca236a1f0429e085e8c606d9be908e3d30f838e8240969c92171de3e6e36b23e0426bd2
zf62b88ab0dee7cf326b419b606bd9afea7fcfa5f05b48e3d6d53161e9f90c048a17ba0e556de04
z227a4a74fa56d739b9cc290497aab3ed64ba4f732fc1064e78401eff367713994734d073f27356
z5e77e13ffe4e205d122bd7066f80e70979490dbcfca168b76edde3e28cfd96283f1463426ab4ec
zccae2e6c38c12a00368c7e8867620322bcea9c624fb34c766a577ed1c94c72de7e05bb1afbcda9
z7cc6496b68b3f868624c8c984048eb95333cfb525a639fee2f223824f4d73a6a2fbd46aed4342c
zd043d51449b6d226bb7108de8de5e02da7422d0ee2d5b50c45fcc24fa7d27939d886694991a4f4
zb1d081efbf2d929f7f0907e7ccaea4d4413d80f22db91761072f2f8b42fc8c0e38c821082c5031
zae37723c21592e815c65b5f197a57bf5a7775fe56664887fb87d885658b5efe69fb805e4388105
z40c079a997426a9a8a4e682913cbbe104d311ca101370b65aa1f8c9a4da92e874e632fce9086bf
z9a2302b09989cfe2b3f0e5ffa5ffcd8a3464523bfd546b0b7bf5984e343c43747bc934cb1bf0bc
z3a4f72fca282a107a111a5dc59ea9875876623cf363242b25658bb462463009365e2ddb4eb9448
zffc02bff64891a8ae552b133aa5a77dc1290541563d0e344f9297247815fd098ba70c24d3d018b
z8e6d5d91d6fa3de3283944358007a650331922e626fd2fde36bea13eac06a975f12b3e879f0ab7
za533568f07e976a2d86c5352ff54e21d84da692497ccdf4317d3966902ecf95636750c052af71f
z6aa3b5ce4e26e88c5babac085269cc788a2beceab325d005d75210a24323548c3b588883665066
z40f159473b2b297bd6dec918aa1c6ee5e98da51104352873e0bc207bdf8a24c105c5d221142a68
ze243088bc54cc9321a815b154e66cefcad29304d403765a25882e96542ec13699ffbc47d6d6411
zb122a7474f39ac3911356b9f4aa11fa4f2f0450ecb0a28f7a44397bb56b746c8b767486864561d
za9137f44d7daaefeaacbbd9fa7757f84002b191bacca010205f82d120732627147be409d00c221
z38c50cccf83aeded9e1cc7bb88913cd4590d21af80a6ac76a98fcaa9c7a633361f417a9a599251
z23a8bc736a55c55c98b84e270b1acc7255587853d8398b932adf4eacc204ceb43cd11f3624dc46
zad2f49a333299580ab29991dccd23894db32a7dcbd8e272400360f419ab94f80d47818bb194602
zd544a62fcd720c563c68cd6cfef79dd0dd6e25cb0ebd41cbb3277195bada6879ccba754712deee
zd39bd859e747e9bad223194d403b4ff8437b16ef325f21f8c6470b1580b9bd572cc2585ccbde07
zcdf3fa5aefe80bf900df3323d5cfab03fd28073e75c708d9a887bd0faf8331a77ff1714c907fad
z9139e5dc1b1d0156489f53de7f96ad2961bb46dbe65e93535ea67bcfd2e8676819104bdbd8f1c1
za9afa5a4b6d800efb09799c84245d3f47d49a77dd5ec067b523ec5b9775ba794d261f56b44571e
zbd3fcff4b6e8420cff39466eb3b5bb987caeada865f30fad96ba1f116718263a5cfb8bdaf7138e
z4bed59227a8d8897f5dcc064e2de6fa866a56e882c2290c79cc658969a263ff864442a4077ecd7
zc471e545c1c746d159bd032e970116bf49615f96ec5b8f1bba22b51085be2b8b8f3b0ae7e92ac3
z91488eb7a160ecc4b74df16bf6a8864cdaa57cafb9a016d01dbe123d9835f972f7b3636aacbb5c
z0dacc151b2f9070f08701dca68fc76637326f4012e8f515f334269f52caf7c296989f17ef9d7e6
z1e06404484ece7e44bff0d338169ef869a382537384e598333fe97ebb38b32c6229e0c3e93b6a2
z1e47ee9b6452db48d35199d7de18e355e59316720d47aa322d413a948cce15714a68e36af1d7d0
z37b02a1a8fbec962210b2a69ce7e4c6fe6f023513e8c718607d1599a8809924b022a38d4d48a22
zd37a107998a8b0def60bc86be11e56759397d4543147770503052cebfd4bbf0ef7ed7f81d1d2c6
zf580270d4e984651da6ebfbe8733f8320e1b79fac4d0965bafca2ab701412b39966443793f0a28
z801389f171601ea16e129d008171593ee0363fdef9fb29913221a454154339bf40c5e7f8ec6a95
z5d4fbb3bce7f523904a37cc3ef687bf7aaf835283705f744c67418b562bf799e2c0a7ddfa7e611
z01fa21826dad19376226715a68983f9974922adeea1048941546b8db880bc5941959e1bb4db926
z1a9b9fcd350eff416a9b2347061d58e87d865bc20f1456990933c72cd0ba147bd1a2678ac89ea1
zd12e1b1ef38a3df69f46fee4f6e4fa690bce3016eecedd3895f56b57b9d2b9edfae06a90e2f0fd
zd88d1a43da2a35ac50f3fe53bb1783778e70a73e89d02fdf1fb97de9145b40bcd70da1910c3507
zf1be81b0e31a741ea539e671dc63c4c801d1c88e0f42b4d52769b50594175f93a26c8cb24094ee
z78f02c7ae5e6d84ea6ca2066b4ff541a7909ba5f0e7f5923780ed0b99413a49271f2ce6f9e4a4f
z2506ad0bfa73da17f78adbee7a1b757bf64f0b8047cd6823c3144fc03c321606926b31bed540d6
z6294366b5abc94257caec477c5584caa479d19f4eb597d17a8c4e835ec463f379b83e3f28d72b4
z3bc5665ff2a4e8ebd6419e0f8fe5e53991d8c48f197b4012dcc5919fee6b1f47b981dd4e685554
z173a6e46c7a7a2432830debd5d7ff0b87646e3c3268ddd42a8a2dccb9bc72acaf7dc81597195db
z83aa029c7c5affad71e45e640d77ad09ffd28c3f6240fdac4a808325748ec7eeda30c2fc5fa153
z1449c31c1af87c47bd8e95d5edca6a6b9d598dea34f086b4ff64f1502092f11af12d678f9ead78
zb6acb1e864862579402261e4d67a2ae9e10bb1abf079d21d26da8b5ba1fa0aaa7c7aab728bb4e8
zd908748ba83703a2a70694dfbd51a2e983bd74dac0b5cf48e20e34ae31b098950f971f31931d81
z567617f85165bfe96d57a2574c0b2e101fd4f6d4ee8c72984804ec8bd19bbe47f0131674b572d3
zf3a6dafbea597627e08356a1484e5fb771dd260bddf36ce62b07bd9d9518445d193ee94fbb7720
z621cfa475cd5959b7c15c59b8b30af68fedb0394819b617ea39f79b8d864e2f08d5ca5ebedd97f
z466e76a0ac5e499ca73c5dbb95988c05133cbc43ca4ef00a2a043c7968ae5c8a11a8be7746d77f
z1c9952d5ee22694dd69ae57fbea5656dfd345e1def0d83e5836e813dac0337c195c11d9dc7d82a
z00bc405d931720800a5b1f483b24247adc82453ced61012e0c5127c5cc25efca4e8c7c2ffb1d96
ze98cc9f9ccbdf12207943b76617923365957d09a04956c29ed8c71c3794f7a92b8b73b55b72d29
z4b4c90db0edc51ff24d46b1e94d4c3e886a9014d9dc6a64171248424d3f6939657e7c7ae1c5f99
zea6acd5355d195cbdd683a3faaa06d467fab87f64de43a053bf697330cb456da080d1553dd31a8
zaf3370c38f81a1b607aeeab3ab2fe6bae64132ff03b11d8afa8685de034c9aec657975954b19fc
zaa0a501607adbf16de3eeb4cb45832401703a4234e341ce292409f68eb48e4d5fc86e39e55126e
z5e8dea9adeb630e7601b40dfd67b0aac42d1ff0d157564335b91f2753c716b82855f416591967b
z2bdfe5d178c402b96e1dc2cea094b7a72cae77de1012d525cbff9af6b4e44e3349069a78076f0e
zfe99867af736f23e31ed248a3daebf3ed6793a06692f9c2cdbaf46105f17f4f2cdaad471e8caac
z429ba40e2837d577ca5b97456eddd01aef3487b33c135dddb9fcb10ce39578dda125f00dea0cf3
z9de0d5c6052ecdca00bf143b4775a996acff889b5f5c192a4c3982f65e935d9c6cbea939feb8f4
zad76e4c8a56c323dbfdc99e6b7db62ea2c9c786a11c923f19fff596344e4e69a29c83b089ad6a3
za71f392b61b47f03d3fff24642fb1949961cd3233a5158a89565b6055f679d09ba0cf273b69476
z565900b671ba8bd8f5e854838f1643bce8d44eec8653bc971eac10f9c9f009b70b4dc49c7276b3
z91775617dd266c19317ca0e1c4bfc4bfd01e560f13bd855a88f42888d74645284a837652d0b486
z24551a2010ee5aacdb033401501a0c1912a8213e93f1f1cb2d86b2ea4d5db98b3db4aa8dff2854
z149798f101bc0c96a6b67818c02b1500801944e6099ca237ccc027773255c41419bf0eeb8dc3ab
zf628f807c16f6395f862555b46ff621f5db3af3e51c16fab409bd87aac28b3fc56f21c6cbe5680
zb9911ed0964910d125e2a962e454603aef67e20d48d1eed240662166b1467bd08a0611e50a805f
z32eb422e7393f9e953d4ff0cfb246051648b5b35236b1ed7e3ad4de8ab5330ce73a65128cd69c0
z2e07870e7f21efae159cc826b5ac735c3d9690ecaafe3e7a717e813ee2af51ffb73b046d61451e
z9ec1d37fdc4ffe05775701916c1c89ab47c8ea683b91b4c40cd7317bca7109bd12804129b8f975
zdc428224c9c517af8625325f18c63757e89bc783cba92acfb8fa4e81db460ceef552c5caff73fc
z338ff7bc13851b6d202ea123edd2913bbfb89b55f65523fc818ce1630e745a2f3dce363096b842
z70cba84b81c21a8bfa32c662f82ce9ae18f41a666f896747d6c11bfa25b1c5933dd3a7e56f350e
z024a1543aca9238eb8d6a4e8197da0156e02f69d60e2252951d5c6b49aefad907eb0539f9cd961
z35060519d1538605d5d3f5ecfe42e727a9d6bf61d1b7e479170fde458755555fc1f365b87020ab
z884c35b831e530899d0af0b7daaf1bd9bef039df5dec59d8f71098ab0a29414068b5b5c3ffe69e
zc1bba1b2fecce3c1ef36dbc43583027d37886e81e2ed1d9436d4fb433358e434cd179426abd7dd
zb4c38974d1f3a1a3dfc22fdb0fe910333630c00bd81d42b80b98f829730c809ad993aeb6eb813d
z5a6b297b5df863dabf28a12f774acdcb1985e191c19fe6df1490bce4601a56d9af4bfef944205b
z9db3e459ea3f53f36f0533861bd75cde3d9ff0618c4b3dbb469a1eaf75cf8f82e13ceb118b42f2
z8f2af82bd01a806c74f7bb73a994c5858bacb713441d67e99705337f0907e2ff4006eabad54cc7
z10cfa02c6655a4d9cbc73836023b451788f667246399affe066c75d87741521c8284ec4fa47e3e
z0811e888e0d40dcf20e5f34d2aac0772bce67cad27740a641af7dff9c83733ebb27b79eef74dc6
zed447bf87c4d2c206bb1665043d8d12a9903151bcaa0a8e9cdcdd7dcc5b9c62a6f76bc4a9c98aa
z718dd8b4ab38f9dfa80617f0afe4a4b61ae398c0929bcbf35110b0250eabe6eea74af80068a3e5
z9723bceb3f96ddac0ffd6b82781666e0453ffd696dff80701cbc89d4168587901e6ae74a5b7932
z7dc84eaa69309090b67563ede158bd78a2b78291312f8e98f6ab661af65d1535fd7025a3a69505
z71ba6a41066062e3bf13b76ceecc449b6ffd83c489da03591608946a4943dd8ea6a33cd0ff48cb
z398289290bc6b2827983e832e2cc17c2165e23f58c520db23880d4d014169676f991eb373cc9da
z2efec7db746f9c192467d9dc0d0e099d26417d3c56f8b619be9c6e7b106058bd00c303f13303b7
zad09b1bba1fb2e3104a233540292e4e2f7faf8b2663d5441b548e81108d77025d19750ab9f90f8
z02f4dd9b2ba4d65070b8afe8b712babb8ec9c06efbd2784530c51a1078b0541c37b31702cad93b
zb34caf86658c52a57d2b1357838caaa86be8772f5bb2dbb156c97a808cd9ae398427c5cd503e90
z1c18195b8cdc18aebff868a0ef97578dbdd3a558adc0e0b81d2a9d894402625240ed1aac3d9dc6
z5dae6dad81e889af0b595dd812ee4a02875161d2f59d1bce8fef987206af432779f8bd6eb64667
z5e7f1c530045230040777be874148ec1d56b65e3fd9a696146dd72bcc6249b5de691562d0da8b6
zd397147669ac1f2b8131653c86ad0e08bfa6a6b6cb5f32e0142ee2b603edef66b24e09a3037963
zc50be84c7a96462f7d1922489696b1b88e2346a3602dbdbe1ed3dfdff1db0239fb25c96a78adb3
z52b46b3b325157d3ba63b3dd701924dbf7b76befb9532a5bf4e40e3bc47d25d986ac5d2c51ac9c
z8221938eeb5a6ca4e0155b3bea2833174323a782570ac1a9d901a86d4ab3a7947fdb60b5549e18
z5d59f72b7a6024b35b0fa36ba89f3f89c556636778bfdeaeade9e41883d8d65c60f6f89eafaca4
z5d2574d4813822f130ab2299a86871e24aff42bbb66606c6a51a4f30886fcb1571c1cf1b81b536
ze938ddfd29d58ac81887ccced6da6829a98772f07bf2bafe6a40194bd528574043e802f479935d
z8c17fbceaba2163311b65c6c8e69ab7e341c42548b041c1f1376e542e8e425481556095bc83c1f
zbcb8e1940cf84522f443a677497a76d52a374cd5e67ec472b2324c2cb23b5b992ef7964a0cfda5
z20377a360de0a115b0334b304e5bfc7aaa56492170329923a573fcab52b7ff29b7dfed6a9eec93
z6352ce22c476f870078ab855d20c791fc9325ea176f9d27dfbe5451a3ba498c65f7c32c0924d55
z783fa4c6ecf79d48f780be83b8f426bcb1c2c83b2448c0f17fe28dc58569608dd17089fc77833a
zec4ef1c27f73be2b060ce8573ee37f3251b0853288f686771d8879780e56f9a708cdc2af0d677f
z2839e07cde85ca3a1a51bee06462cb252bf9bb5bf6644120133f75aa3e414a18190000518ec42b
z84cd7d0f4e19cc44eeb9fe03f9b76ee9b9e2f67e0e6b56e438d0a0878f7d1ae4deda55a10a38cc
z24addcb43a42e1c9178796a15d813fc9fa8d432c9c06179007dabdf26a218c3848942174670079
z36c02863b22fb28a895fa4232e70ee11a25237aa0542b8aea4d920bc108d9cb1f299eca7d373ec
zd22cb85304b5926592b6de16585d4a99ac2a65d61d206fd3c15b09f974c9d3cec316cf211c6503
z1530b25aead61fe387150ddb5651f61b5cc55dcfbc13b9957313207796b1aa57c79e697d2162d5
zbde70c602ad6cfa632274e59539a114a492659ab2a1c68bfbee19f5b080a4da2de4d79d948d9b8
zd19150ec56b85219f2a683fe974a0d5b50f2d8518f6808d98384f00220be4aba1d7e81fe02a83c
z0e1e6b0258240d37f46397585645bd73356cc357cc0afe5558bdde89e9082306c076fa2718d9c7
zbc42089fad95ce5e9ad0dc7157df6e04b685390fadea6b12fafdbeaa019be4d693cb1e911efb14
zad5f1ae1793cd43f86fac9b64bf577ebb6d149c04079751e65adb05692632c7d3897d201ed4323
zf2336a2159f4affbb4c00da2e3fd4056adc93e16a90bf9fd27d510bb9a0a8ac58b1ff0ea124c15
z178d4fe7e1a65fdc6f511861723ed0770a1589e2ce9b503c21838eb1c36d117777f76d85bdb21e
z45f7538221c671ad68ddab1952d99b0d3eb1689628f4af8989220366ab9fbe2d51236f6b82bf3a
z4b50895bde3867f5e1940fa21ce9a8bc461f10c72cc59dec08da7f14c41d21f867bbf3958c8a31
z59297c6d6949aeafb43fbf86bc4dfd656147925515b341c4c1abad465a8b74031fdac333fcabe3
z7ba2704e19ebe616c18c6e7daa7170d9484f9fe7b35560a347be9200bd12a2a7d2b562a8c7ff3d
za3a1049fdbaf739b56e38c63080a91ff2bc03d396f0318dccdb1feec5c372e4311d50e7dbfd024
z52eaf710ff9094f46f0a095e3a8ede05dd958ddc09ff76efd9df36a6383430bd4b36823debcd4f
z335612b3ea1f82bca5169a915ce24a5c0aff3f0c765aefe59d10f9cb0afcf283d7c8126e9950d1
zafc36d8385c4a9e3433754052b7212342a1dd862e5145f4dd234868747e59053c8efc2d120478e
z877f731fd8d025635fc1bb8545e96eb990346d761c1ac4c729e7aa6b1efde3e90f4a7b57b494e6
zde9066593964b948ebedfbce681027074ab9850e09b3da0f6dce7dc0d252c8663628b3c636da09
z5d1fc3450b7a82751b920891bb5c8cd482530f98cf4a5ad0662232b91153313cd3a96cc806b7f0
zfc81ad9fa5763877e2fca266816b9c8ef1369bbac53d56f7b56d48d142e3ca42b023d1b0e0a081
zb7546ee915df4836d076356e845c73cede130427db06e1bce8a5c6c0630b884410cf95cccb95e8
zc25f232f2333bed3b2b7c6e5638a52a4cf509507daa0034d48e5eff84205f7232028b603bf5e03
zb65bf23b5b2b04e487cbaedf3270657443d68a8769a2e7407bc4fc78df590a3da66de25500c9b1
zeee3c941eb91b584ba654320c3b8eda29c5483759388cad390ae1520484208bba32c232ad2dfa4
z012016087d51f946fa49845ab8bd0e10f292542cf34307a9b15094d25d1801c82c606002751b4f
zc76707fc8c2133e9e333f0c9f92c67acf2421d8fbd33039f42328c2fdfe5d392d46eb5f5879f28
z4fc393b5ffe8c843a34bf5621f4ac8e4487bcdc27459720784dae22350d598fa34bd704418498d
ze058227d23a96fd25b622afe79f9f8f201d202023c5ca2f70271c63114b48af7530d79d40ec472
zfca615950d6ace05a4dbe4d0db8b14c3ee641f9edee0aea59003ce7bc88dfd747b005885efee90
z1971efdffdfdae4f62b7b0f6bc7afb4a10971a95bc5485eef3983913258aa524ed53c496c9374b
z996db1b76d0aedd6dc771534dcac61bcf1e2b41fb85c60bf9831c37e466a51be43d5ba9c04be87
z127fe5d1e2d13524e7a8c65cb17199b339ec01a968ceb12dc2f3ab2c370652db596938fee43f5c
z975fd4c43e982f1ecffdac149463f48cc9828f0ed0f22cb46b91b3717a767b5779735d404ef825
ze81d93905ba5645598798173762cdca3bacf96301e36736da3a987596ad240befa285d70e008f9
zcaac0aeb8434ae17d93625a976ba0bc79981787461fab78890c5268dcd416bc75d6308013bab1d
z8c6cc6c1d8dbb441a1bcf602b2a0f5f8f886d86e8674c7879f0dfed4889abb14bdbddd17be56e5
zc04ff08551d354cfcffa22ac6df67184fc75fafbca2895380637370d992cccba9c8fcae97fca84
z14d86003d11511fdecb5f8e8695a681f4a13258d15dc38633f11fe6e9b5c0eb57c5e9046c58079
z125d690bcd3c8e3cdf68cfe8507b84882fcfbe60e09feb9b907a707452962e15206d835177f42a
z40271eb5587887b5e96b453a2e2ce412b21a5e4a12d63f1937b14bdea357adf450d0ea23359d7a
zf001e3f70610cbd4f4dd1943879b8cf2fef0f26e96d8432ef08a7a9c1a09a6c994ba95b089c0f3
z9a8ed1904a853f3702f0a222427e4f44c3764e5b07d7c4fccc238dfc2398c70f0b3da467ba5431
z22b2db88930054e5bf7cc7b95917c031382f7c0c2678ab1a13a0db2bf981a94f98d2b90728d761
zb582eb4fb51e1050c99be51ce93c4038f42b05609c6105adf9812558acc67ca37fcfcfa2b64e93
zc2499f171b22b2a0ec34695d0d55bbdb77c7ad3bda867a4a2e537f7a4c218e3da2109d29653ae1
zf67110ca0a0acebfaa32564356d2548526c21b5985063234c261d71ad39df7ae5ddb1e7ea5d524
zdbf57a62ae314c6ddf442dd4e62d7e4e1b595fd98301c99e8ba31eb9655c2ff7aed7be3d9285da
z0d4869cb0ad10dbc40125364b1354260557021e5b937d0574b6ee3c5edaffa02062afe98d6f965
z80ee58a9fa7922b6a82e0fa9e8ef0657ee4a7abb0648618dbe77e9bcd63e67e18b6547dd8cea82
z382c4079f6288978e858f990ae2a466807ece70370a7a085e9ad0771210cf192f29129983a2ef9
z608db8ab43934d270e9b0ed3f682ac5e5940fd3a7d27399469664a30b6a94fb0dd135fb8effe61
z1b471c7d6ecb205440a0cfb233d86fc986a56ff18594727ab3b57ab74a03dc0b6dc2c40349e672
z86d39d6d26243f6ad0ac2a29401b72c604b5bbe543e19cd3501f3a88b0e5bfabc0d6311214b0a8
zc8910c1e2687e0b7ed98d1c8fe98e18561fe6a08099f4b92ee819fd547773e93008bb7a3f68c53
z09613d925c5a3fefdda41ed69e22d52c861f5cc6ddc83c5bc4e305a6ad0adaf2b493ffe42f7776
z9c3e994e51f0b074ea75c330eaeaa4ca8fa55e3410f9a4c2150d47942d62777ce29d0ad0f1f993
zac30fbe3a9bb2182a03301dc3328291a6ff151edefa563e9ede871396bf7ff623cc7180edc76ca
z5999531433cb97148cbd5a6cfd94d5da6e5d8582bfae5063d20bb9214b775cb9a083c5c49be62c
zc406c6ef9f0090c4ed6c5fe2c2d687c0100592e41120bdebdcec860d28ec337b4b5720675dd2ec
ze619eca49b7d327a2a8f4b08677c42027f56c34efcc72911ee7ff3554e92bb48d21fcfaabb7c49
zb1e0bdf9746967d5254159bab5ab3c6f9cf98aa645fe44ea0fb0c24ba9cbf05a3581e9753abc99
zcb26a73d5fb7282fabeadf38677686a774d849cc99bbf7e9e4aa03169335d7bf700b5b4a1f45ee
zc65db3f5fca58cba23793cda488a5452979a931363af66e519740920f84f7adf09cf4e623acbe7
z3a43c7baf945d924fb3c2b3d00f85718cd0daf65b2660e551dfcc0396e39a4f7eb24efb156898a
z5e0a599a7a2bac16df6af2f1551ad719827632b1497810842d353f37b22ee747d55749298a7df2
za6e4fa26f29423aacc0aa796857c1cdfb163a3bbe206aba3826ee7e6d375c9d3520ba3da1f1d05
za610d199e6f02a8013fb023d47479206ddb1c4d235a64fa3301d853bf6c9c205bd71dc156d4580
z5146e39d4dc39028674969d084bf5cca914b659fea335ab57f3f59429006f963504785180e3f98
ze178e0df6f29171234ce78ea3c556cd85ae2940755335ddf9662d04976ff4edab70fdaa5ee2b84
ze5557af803057b378a4d2f95bfcb5d684980fbd4df50cc27ab043d8b88a08f204280d5d42170ab
zc61fdccc01d98a48cb78fa73037625c29fa2d0c7edfe8ae23c059c7159b22be423e8138d4d7cab
z4d29ef8c38c8d62a630e09a70056f816d0dce52329575513afa0f817baf9b6fecd94d01e936545
zbab46d92ccb5f47110762b8de7a86fd13005d37cc139ed526234d83cb6b1d250928ac1754b460b
z610b887ddf0eb7d50ead853e6bb43adb032dd9098d4b63d2572a8729bbfc3c0cd7e1f76148a459
z4ab675ff40059202910a12dc1d376023f198b717eed9086637867b06d089e2d3eb7b51bfbfb6be
z91df146c5c1edcf78823c326e2ee24fc10cfec5967b58c3fd26e57a1e6b5c10acdeb4bd912f944
z7974c5398e2a848a8ca8772df219aebc864c1f994bbb86bb0648c2fb5ef7c10c93765b7a6dcdc7
ze4ef45ac061ceefb9e36a6ec558a8952f192d0b9aee9550ce368c88613430d70ca66cddf7f10a3
zf32e0b982b73df59069ded94bbcf8e043d2cb0dc605a754adac7b45a692085e9e37259ba17b9eb
z11a2ec5e1b7864caabc72d5b751fe94d60d1918c630bff50d3b5de5666c63e298cfcae7d305cf1
z019440090f24443f7b702aa0d4e78062e4964f3ca3335e5784647bd43969820a33a7aaa66bcd02
z0e275b3b7c7c937c3ba1350840ee5bbdccce6be156897586e2e6d9bfe234848a9c18bfbe6951ff
z2b4a30e7ffc58fc6a122c6b7d7b1df91440ab3e151735350b33adb51a3c7e5ce1625e0eb79d6c7
z913e2ecca021dcc5be15614d2a640edc127d3a7f826f0a8d1dc0024c06081e6c62be241934c341
z8ffd08959eaa2102808e855672d7ed78b06779773df1a3091c0250770a9aac71462c625061163a
zdb86e0a4213f66c0b4863a1a207276f77f1fc929e048b1af7ec51b7b6176cf1488b3fdaa580e1e
ze20f96e90cb5e635082ef8024e91e6791af14b3af0c75639cb027469fd978869fa790f4c9a451f
zf807a601627a66db368a270ac0d9aebc2cfab452f10430cf79e746a4dd45e1d0693acf376b124b
zde49a453966c7ad09bf88ac52eb6d2ed82fbd7c176adadcee3dad166f5bb2914fff8263e2b535a
zd1063fc8bff640ae018d68202789a2f338bc6ebfc17f4bfea8d6bc374a6ccc89582394591136c1
z3f61cd5f3425d6562177040893b7cf99224dbbd39cc0eed44f206f9691c3c7ff7371e2aa4615ce
zeda552b9df9e83558fb74f5a806a96dfef2a7613052bb93f713b0563a11d7dee68cf1429969343
za9f611345b3f5576ff57a6f4e54232031c445e115036d40092f2854aaccd8255ab855bc2959b9c
z5097660c32f90e3d3430b0fb53d4fbfe43d79f51d041ba315931f3327fd12d2a07cfdaeb98ec35
z2b53c4713857d69965df0698e3de740fc44493d7c9fc8c031c285ce8d75bbd548124c747d9f7e7
z4fed64927c0a398eb67912c9a2e2ee471b564f77072989ba5d04fbd54359f6995799506f4c83aa
z56b5ed81112f52d3eb976ab09d43051acfb02e377d9da37bd471df37f5b75373104a1664cb1de2
z8216e645fea2649fc2c1c9d245c013fa2824feb87e0b2d4659ef6f26696bf20aca3b176ab01844
z4cefafcc2380c4fff3b45ebcc0f91e8818e4f0f4546a47b3907026dca6b51b77815e581d66b50e
z711aeffb93f0e08670e30de221ca0cfb98576fc0b4ccb4db100b306997a5168f91baf16979f417
zeb24a57f3a22a47179a9cb59cd76c8e1ef41e694226b10d52c15296d268028938d2e859ddb441a
zf80cc519cf76a8490977b64e4bb3400c13c9aec4032437e9266e61979d56f59866dec543a63990
zefe2daf3c88512a6f3bd7ce711d975b8c4c4d6a9eac1ce8a51139349e09b0e824c626abc1c9df0
zb0b342ddaa91e69173e2f96ca08ae2f88e5f40ff224026a8cc059c830c775d1d1c1e08ef19026e
zdf1c1bb06300c043fce53a11a05c9fab0566364d60edbaf72f0c66abcd4f8b2473b79c3b3378ae
zed442123f0b64de169b9f7589d4df5b61319c08ad01e4a0bfef0df737ea4ebd51fcdd3dc8c0cd6
z18feb117d176c4ef84fd1a0175de581e33c5c7e0d4c8287586c55fb6919bc82c96404554343334
z0db75216efd24886d8897582692430da7c0da2c6ba5ae7315e28feaac8db5c7333beeb976da874
z3d0aac37048cf9c7d2fc56804e641f1e222b9bb1b53e404b14622f9a800ee9fada86eaeb6ef027
z11d0aef7674486a4ba538cc4a0bcbdd08593bc950c1f2c05908079546c84d7bf142eb59890e0aa
zba38b1438fd89bb7764169af96022e2362be4d9f28214952b625df18d248dc458d86308c328ebb
z83cb49667ecddcbc67854633885541431fbfbf0a5af23892d059e9b4ee5b8aae13600f44205695
zc87bb2df1bb039e2e12d4078a655a779e19454bfe918a8d494134cbd5f41a229b2f959510f5e7e
z0e44a3fb1a09887a822aeba3f0e375e10c7b3fe745a2d6d725c1983aeb686df983829f040dbd55
z126671c9e0e729b955cc8b2bf1ac3077fdf5531944dde0dda043ce6743ca39905f855cde72572d
zca1727a53d215e587f0409e6b2d71a7833fdcadbb21168fae05ad43b7d7061e97d7d4610ac9224
z8fc6c332dd489bcc1725bebe6616339595b7c106f162721a804ae6a35f2a91cb63dc079b7eb9d5
z935632af7c5c23bcd15ae588c427ec97ede2e6f64114b0cbebe350719979bfc56cff181818d149
ze82b6a6d852d653b94b6036a18986b9ba780adcd7e97543d56c8002dc6f54e5bd39e4832c79126
z47c922f9a16c9869b77a0a3b768bc906f1488dd02723e6da283b913f1cf1cca94cad15d2e78d69
z300e1e6b2b623790fdd853289ab47b15426b74442046c0aaf904fe41fb86183724be4a7a8d9b9f
z6bb9225481c31853550f8680c5210bc609119c4abfef82e6c2eab32b39f94b4dd74d47e13f8637
z77585d140e5351069ea575465a53ee230c7c212ef13876e05a1cf3e3264c2fbf8f4f8bb176258b
z60532c1349d6675c526b0f13d15f2a0377d381eb2dad65ed39e105c817328722e2b240c3ec6e50
z3ddf40b4b346f4eac8bdb01bc723bbb131c46c6a80707d62325d280183888dbc6ff054365d3492
zb263dff03bb9c96f8df5cba9f4a23b4ffd9e5d8d0ced7a0d3450785899006627bc74c8ec2649d6
zbce942ca7c8f462935b7f26c7a3baaf61a49d77a337607a817fcdbfd824e823c6a175bcc5c3cbb
z07c4287c1667dbdc3d20569db3fd72c0386ec7446b22da584454111e08b4d9b4b2cb7925c468d6
z20aabceaba24cb8f23591fcefca2f61c3c0a37a522207b5bea8785100755f556df502d48b1b90d
ze6d1fbd340aa73ff4bd90726449b2559ede699540b253f27e950523ad5301ff8ffd7e471ac0079
z526e7685802bae4564a7b4bdb57ab4f215ba742c5d539b70df6db2b5299e8dde7ca51393698521
z4a9fa486ef061f80329f302f11dbb7ceeb9a88476b49c24e323c77fe3688380134ff09965d010c
z470df3a90ae2c8c83e5ed732ec640e83ae11a6878bbf547d1ef92e6f523b47d867fe3a9187b103
zfdecf87be78b689e31207697043062c318406758fc35f27a6a5aa3ca179df38340104d289f854c
zbf3000eddcfba576b628a64b25204f3f81e17a82d2e7d512f1426fe9e3970a7d01fbc240d2b196
z2c2de33c221c8c2444efdc08932e8aaed4adb0daf633ca950e68d20a22c8457583bab43a4b946f
z8faf507cb47c559db07f446c1a51255654b49fe8ca3ea416e1621cf14d7d759465cedcb669c8f3
z18ea2e2f56ec767754aabaf138ff38b3b05669b368509c6bcdc548da5cdbfe33a59b0dd8543211
z691ed795b243cc00ad9d933086921fc27355e7cb637cf7be67883532ece27c0dd05223312c6743
za3b9a53f581de6174741cdacf9faddaf3381b6939eda47aa859b64fb6fd3ed1065bf33bb5b2ced
z57c38e1f37617507d69bffa7b082b6c13d805da8c3d32aa9d682639e06274c025ae7e9865f5086
zad4c369c876a77c495c5c16cfa2cf95414db9f5760ee3f469a685e3807129767f2c20f74badfa9
z910e53b96b5f3e07ee3ec875710666fe18ef268c82bd6e0df9250da1ecc3fdec351a418ec6ae10
zace459a520f9cccff401f0c1880ab603236ec224011fcfdf0af648d357369cc2afb36a72c1923a
ze3dced633ea9da5a9a7f4ed9594cc7e958eeb939f12e099127557dac63382d12aab9ae52ff56fa
zca55cf3dcec3ef828e433b7580c9fac8ce7d187b088f700e9e83c15fa834ebb242b2bc8897ab2f
zcfbe65f8e7aa99fa040e74c9b2fe2d17812fb6409f2ceaae534bc6255af49b7e0e0462a17bf81a
z393ee5862b881c96cab0967017e7c7e31f3699c25316dc0637228f9b86fc7fd60c96ee90f613e1
z85881d20b09d34bee35a52a0dd6d02d4cb3462ffb2d8f4ee2a1fc65fba3739ca05a2cb5841bb9a
zf1fc368e1a6a6dd8afe7eed617ddb4c80771f29a690e24932cb961ab07e08cb0ce35e51afb8ec2
z0dcf36ee85a374185e89e32a1b3509c457fb6748cf3098215132bfb6686c96f233c2cf3384775a
z4b76ec426072d453b9d1ecf53be0ab0d9e111e4ca43991a2afc2e9393b55178412a5ecdb97563e
z9149f3ffb9912a19cc20a6f01f97733717ecfab9394e347a5ed5226818a72b3ac7335c440947e3
z55d3442dcf8d97d89b4bb90b70e589ffcfb7ebbcd7c2e153e0c85b132e909b13bef59061fa884d
zdb05373e5b020a583fedff81d51d7f16fe40558ca3f5b41f770b79bf880577a25e1d75fa4d9111
z0e5f74d2379bbaf5720136539c848db493b95d255a43ba10559474f80e07de152727297c2939ed
z679b670cd92c4bf9ad9d504956f6111fa67f54ca40239f4eb788d618513da80b8b3b22378a0ade
z7f627ae3c75b5d7e954b3d80609488b9735796fc20c91045b9c1da5ba9c5f77a393bcad4d0bc3d
z8be5a5a7aaba9ac8de9bd75e180ebcff699040b25f76afbe1f33a013c18fea48b94518f0a73431
z8b2ffabbed0d1a84e36ab49d97e8dafe23e73985cd907558400026efdc8ba3fea96d64a2a60c3c
zcf0957a109575c61488fd37a819213cfc85450c8eb815769dada52a7966d2db5780032fe92a87a
z16b49404cab72a00dd540df678a1100c87b0f551285773f55e4f0ba7e9443dfc66b1e14fe37178
z317ae3efc3b52aa2f652377e465061a0e0f337d134a22a518b66a316b5e0ec8b34a40814f8d2aa
z263521ec5840eb15925ccb17484b60158b1aeba700edf0660ae4d103aa9a28afb883ad43076683
z9981c9b3b706f0f74e310e5d39f5cdc75c0ddcf9f86754376a5b15252ed8fd3da68ca81513967e
z58c253466a2dc396bf0e0c60d9e4979510ab0b31d1f6a78a35530de0750065c5b0acc08ef01a0b
z5856a184280b5ccc0c73b1d6a33d0d4588f51a3ff0f047fde1b7022eb346e968d7cd4f1da8101b
zf9890983beaa80cd9a4880e3d0ebc9320e9980d14d88cfb32916356d7f8537ced8bda24714ed51
z46376ced68a4226f56adb475d63c3e6a55b2fe9946c771c096f9a5134193f45d1a23c222ffd86c
ze1e435de53e525882ee107cbd673a31c255244344e7d2edc4a1983c490edf61c75a706030451a9
ze8d7f11320d00ebc9839d504c7fba3dbcee1043850c182d417c76e111f2e74fc1a9fb9ddcd4a60
z454ef5ce7cec7b757f9bf6ee122d53ada9675c9d6692fdd7824584b9904496c4b781aea7c0a130
zdfff3d87202caad2b986769a0732a1b00b116e9bfd653af0791283ac3e55b0c83764e34adc316a
zec870df5d06e2389007c8b43f31e0fa2ef872f7364c7a2ee46d161367c2b7a7c403b0cba10663c
z2b6a38a2a676040051375a43c8d7318f5828baafdac57df26c1b2f9dbbaedbbef0667893a394bd
z3734ef7179734543db6af9a808a6f81b500d399c7e7fc6c6b38808d7a085003b1baf3b94c065f0
z9940784a728f9cd4be3b5afde37b375735428a9a8f5edeaf051753efbafe8c0e6b1fc4e13a8fa8
z942477184f2a868b4ed61bbc164b03af6716b09b314a3566500be97c936cd9ac87c2234e18e85d
z2d8dae0f04ae3f7eac1f6af75e1bd483a3a6faeeaa83b00a698f3c03383c7b2f3cac92a7c9f97c
zc19352388acf29a783bf12ed1a09f8e453450f872b77ebd75e513206f9f46d7a8d58ddce9f11bf
za7573ec5ba2c5e22d2e8fb7f1a95ec2c0e0b14603516c4668964650e62766db846fbc9dbb39095
z31985a1a78918fdfc8e3c58eb770a3f904f077dc794164f06dc2ebb261cb555d92ce8af74fa608
z3342682bc98a38970f8060438e6362fef99373a58c871ba02c739ef77d7c7ae01302db6561c311
z92fee0e86e71d68845d2a142eabc6ccfd4a6f044d37023aaba37af9197e75ecf4541ba455d7c0d
z75e3da26000e45b9971fc05f13ebfc7eb5c30cdf0a2c4f176300d2def6646e72bd4bce95582cbc
z09ead11a08bba7e7a6d2087ae8924b61ded9a647084782aa28bf9828ffc1a327ead20348a7e009
z5364f4bc2ea6afe73419d115a99a4a0e81fb9da829dc3d8f880cb3825b164eea8fdb434364dc85
z51f987e7b4dd5227f4ac05c6f8b7eabd310d09ad1dbe0c071cc9f59e392972a5095dd5850aa2a8
zd51b5ed2e0912802a17a22aff5ccc4bd5e4603eda1830c74e8dee081102ee5a8e9f30d741595ee
zf2154c11da294ff87130637b258316ea4e8d622993090f9b5f36c62c0080b7e3aac95f8848996c
z8d0255acef4b4175dc9c869d8d4211621c2d54dd2f474d78e06d465b2341ff11b450fa965e2075
z779ebbb0f866b29b4b67fb194cbe85b25ac65f64e11abadb0ce2b768fd2c155454e76bed510beb
z8df5192f0c546b9d684b37270f92f88c75f185d74d8b340ec7f43656dba916e66f2f42f43b3365
zaeccacdf48d7d0912c7374bfa8b715e0eab05220066b74093cc19ca1dfb9e3acb22c6c8bf0349c
z3d7c09cd2102c8d3c8361ffd292afc2c4c62efdb88d487b5800da319b3b28562ec4cc92c5e21df
z667d787eabf722b077729308293e8e63a097323af19a6c164c13b09b450497ee08bf8581b08560
z6be7ceece0af611864ce3cd7ef2009ac9890d2f9c63c32f36b06e7127a63655aecda90185e1228
z22ce264e6475ef2e2ef784484b239621f7b8a85410bc0e74de1fc3d2d3b7d16641a8f24f9a24fe
zdf3274a31032af23e3b1bfc23d894a36fd8328acf03436d3e06b29a300b2688049a5306e48c171
za2b3c11143ceb705f79e551f4128134bcae5100905206677c57cd0338d89ef0ecca541867d2c2e
z1e3a37ee1646425f03b4fd0e42872eb97fae98a8ed6f70d8f66275e2a3e0b3fc167a856d1260a6
za059d9138118e168b307fc3bc6f8b7a91a2d1c0d93a1f2baaf5e342e164f44c7e144019c32a8ed
z1b2cfda6b028e11db9a4e05aceac9cedc3ccbdff224dd1247b45b5f86021659b28c27e4d4ee0fb
z3080cfaa37bbd0bcb7fca97717632f8eb4d7fcd6b26ba43876cef2003dca565a1bc968e3d4191f
z6a4ebcb43d72e46a111665fbee5b8491b95d56c0520e350d131bd3ca2d3777217aa3a1193da5f3
z91cc0d11a1f46afe76fb5c8e1874ee5c8be39ac84b0ceb18bd15bcb65b5bbd45fd928e89ab05a2
z5de711da24338c015381da1773d3cb1bf9d27b78f735f52c23543fe05aed63b212a93e7b0c7653
z33e6f651c999a9e9234ef4c629a9db42de65d80b1fec139b1c7b758e366ae5c783ab27f4a7e2fe
z5cbcbf79155fcd10bce3d92e9c39b77e9eaa73ba80daaf592179a46afa2566d0013ba2c48e2b9d
z42231f6a1b8880e6b49077ad411df3f69bab857f83e049eac2d713fc2c5b3114212f02549f8872
z66d5e5f71475c80a237b07854feaf023750ddb9f086ad6e48995939df945bb0ef22ea122f551dc
zd7097adf1e428484c384541a83026c9f50ffad12ee4cd10dc0e937efad6753bb960a91bd32630c
z2c34a20e9996236eedbaa72e7bb32dcddeb7e50736a47651a84b9bd6f12b0f18e29594022968c1
z265108e01f12be5474bb0dfb017efa56602b3ad2d8f077e573723b7af46a45988e91d023ade043
zecb310b8186841191dd935f166e7d86f3a82ded43657726dd6a27ca1483f656e2a85b59bf2c071
za9b1e0ddea17b8402992c0150e4f555ae5dd2c2e4aa3c8e38a551eb4f67f418059aa1f83200c57
ze2fea64c3ff40dda0b50266e4da3c66309409be7440683cdd0d72625c30ed2873651a8d510f4bc
z83fc499ce4662d60a8e89d148489b2d0a35add17792f17ea00d3c5721c824eb6af254e5bb000a6
z052d6b17e066e05ae9396e8e4de8666a8f776262b7672cf17f8c65d30d9805841e77046ed3daf2
z2b3dcd231a945b1c44f765e5e0eebf649cf67cc252ea0046a8eee34e8fac853c904e2518caf7c1
z99470c81dcdee2f879012ca75c82d8f3063dc23ff842f9806e4532d4273c46db842bcf06b1a3ba
z91576398cb05ebafa5656cfb03dc27ca4e802ce86cb05f6a9568bb3fa6b46fe8cf86871bc8587e
zfe17d38ca3ca6e3f90b1e4d442d625da8c85e980566dae5f0011f19e720273535aa751fc8e14ea
z3b97a19c423f0d1b7433012c9775ee95553a237f8582d4967238199fd69c701741c1599ba40d3e
zdb949638345f0e640a86097ad668cc30fed4abeb57ebacde41bd233a8ca757ce6260c98e41d4dc
zcdf8adbc835b6e54f9b8b75843f767fae5eb656ab8f3518dbaafecdf2c2a3f4f8342688b635b80
z789f66427f5ca6d330621cdafb1e78df72d69612c6153eded3f06cae78bbaef3b4da35ff4ba947
z64c1cfcd6b1901f1bc5e9c63d23204e54d29b29f782e7c409eca1903f2fbcee041378eaa6ff952
z4eda0428fda3b94ebceed83c7d690f31a3fcd4ec01bea3b601b1820d0c414b968a2759625e9dd7
z7bc65ef560b5c110a235f8e6aafed1bb3e38b3b8dd27bcad57cb8dc4e0224bee7dc0cb6e7fe876
z2cc3e50f51cc5e4514f51ec2e66322e90eb683480e9c55dcbfd3579450e8068f69922837b6aef5
z4c7ca154fac8d89a0aa10e95a3ed9b915ff392d7990588a1ef130f6b0fa9b6ba38cf10befb83a5
z059dad82b19c2fed3202c3529c14fd17594eb883988a3ab1a90d5f18e2b3080965156ae3e6c9f3
za6ee40afdaad08a0aa2913c418472a9955417fc3ac6be4d78d451302044e8ea0a731152c6e782e
z07380d8e6d2dfc5568701d43b89e78a6b5d7ff33caee3991223eab302c94c10d98f6734077a461
zf5ef42d64cd07f5c5916ada66f251e45709f536b0a6e63d25bb5028eceb9099adb6b2b9a49079e
zaab09922395179d04a0ceeff090c8dd59d09206317c746557a07b68d2e0524c5ae0fca4240d989
z2d7eed1645812483ce681358529bdc72ea2d88a3bb6b9c0cd6b7e5ee08fcfbe559ee389a4519c8
z066c58b8254614e50f079c2ef4bae2c1e82500a403214af9c42026d31bb3dc4924a4d52f60d736
z9880364987c233bbb460218f84c0a8d2741471c57cf429a6df1b2c0192ee25455e860259e6c94c
z253b360dfd3846099ab4cc73da96216a692d1212bf73a14b5ade97b60873c363fece160f65d926
ze15ca60cd0fa60a9627304dfac225aabd5c2a7b7b89b876b5b8f94ee738fed9fbeb8dc0eb842c0
z7c05e67ba918f010ce211deaec7be009af5c1fc51704b8165298ab2474e3a7c18a5811e81a80bb
z32301b463c3f30e1f942e3b657319d3cfa73172f9f538dacf4ca4f914a5cb9e8f7455c6ea1836a
z6aced4d7a37c8315abca5c53c6b7c95b6a2304795d508575ea7a26ee093a96178026bbc71480c6
ze1ce538f62248c85d5f6237d183c1d8de37167758c3fec757d04c70f52736ecc59d456ab2c64d0
zc1441e5992e7249ea188185267920d1d7186e156f6dc062bda880f60ff3c887cf9617932c4a0a7
zcb4b15f48be81c906ee026df53fd06dbb5d13a60d719b9413300be28be6278a39d0b44c182e648
z80bf7c08dcab9a918cea28c7f7f084f020e3c86d7fe28bfce3fc45dae54ac38ac99c63f84ed4f8
z8f848e1bd93a93b17d47235ba76c48842c8598a336cf8ee04a65da727ce484b540e386fcab2729
z0d4ae8cc74ef0f50e97c6199a74fbbaa2cdb132203e6ca180dd3eb220ac049d45c12cbf0790c7d
z22168778e8a4019cbf187ac6fffba28699b98c2bcc3343cf1107d0166b5961184076f8f39fe65a
zfa930aa21a8ba5d2460765a0fc8daf81f3e96681d0b66ba44dda15cf701cd33e870801f5f976ea
z2fc490db16f937bc0091b69e8afc564c1802c2693b5e4b0b03c83d2c40d012f6c595444aac9805
zd5be21f2c4f97d1b8e7c5d534429d572ad9ba119f8a846b515607ee4567b2f4ca38aea22fef79c
zcb3158a4ab03d5fd0ea4d958bd55366b0999c3113783fb003191ade353fd6ec9869c75a4967bca
z7cf0222fa5fbe316d5c9b13e3f83e1845c8d1eb38a8e4e66e6968d51b70dbd19cb884e1d0c9c4e
z6a69d6f2209a70599eb012e7be1d07c30a0dcfb18f66ad1beef21b4bd9356cea91ee4140ce4185
z533b09ebe0e9e5b1d4654059a8230392949c0d47d0f297472b6533c504c7a06f971b74fdda38d1
zcfbe4fa0cf6ec739f0764c6b091269c3d18c9d8bfb60910bc14f5dad1d34061c3e5ae76704203c
z835e3d1233114d24dd3ddf2037136bf705cd9dd4844a09c8d62a2842fdc432305371491ccdae89
zfda1caefa8bd48a0f9f39d96cc280663f18b54d8c2ac359f7fe3d2e205533ca7fdf8e56d4ebb39
zc35984169b4406e2bee104225fe6b1d908f4c7586ed414ccca03084dfed67c68d2dbf8fe6d6365
z4b1bab7b34169bea1491e68e8cfd0c5ddd0bd0be7aa8bd08c9d124091120e757eef3bb3f30cb26
z564e54781d2cc471cd3689de1b8e10851597271574234d5ccbcb64a17fdf05b40531891fad0f2a
zeea274b68e030df2a04ba84431ec2ddbf87702d8b3ccd754982fb5b4959aa2471bd80c89ed31cc
z54ec1393eb1b9800bd989c93d7a6715c304a68381fc98fdd02201db8faff8aeb2c15effaf1627b
z3b2a862664730416114479bbc9b283200e1311147b109010c9c9f9a512e5c1d170e2a28ec15699
z5c42f63f1207f2571200b74fc66919839a04bdfc725f048a0dbab46a02967fcffb93c7d723f30e
z9f37d32e7748a9bfaf612bf2b906ff9bc1e67634aa7048d6892e89c6faa9420230f0b2986e7307
zde872d8ea08a053b55017641dbe0597eab370a2edef960c2c4634a469cf384dd46ce8f1ada7b78
z767d0d9f71536bb82ba7f6b0e6690226c3628da2d3cfb12dc0f98f919d52756433c313d91f15c8
z7095ae6a85c4c90140b9beaeecd48186676015eb6d04ecc7c725c877eef29270b70b208b40b8f6
ze0f89a7ad6ef59cb1f579ba071bf81756e84b608443cafe6b919421004ba7190f61462310e002e
z464de8657414b82bd6ba744bc0e59d8ff046525f431c0914cca5b1556894f5b053f893d0fb2186
z125010580be58572e287b28adf163a02d6135d727e3fd04882d95a9fd49bfcb582d1c9078fd2cc
ze6563b96872388908156c12005be6e175f7b59e15a8e5b8e54b1d826c3cae137e732ea1d76bef8
z570214b5c329b2519dca5447cf5c8d837b278528fea63b4c8f017b76acd49c74dd4b1b2171e9e9
zeddb8073b987b7be8df13f6d8861cb6c6d69932f67a26e76dde1e34e9425b62258d4e1e44dac41
z80c0def2ec0616d2458d74eded6e9fa555e1227a4207c56580c2f20088f96e7ef6c249c5752224
ze35ff18a0bec6812ff881d1590b57e0c43ea3c2a913cdad81f4b4e59a595564b006e95cc65581c
z38f655c34bc99617d57fff1184b3eea4500694f82839f3490399e1d79ff9fcc4476ee9be2b8a6c
zd4256ec9a8e5feb1602704788ff055c64ce3ab53c57ae7af4670f7fb4941a672623a665a3a5dc0
z410813c865d572d84778470a2095ed7e696274679842a5a5a384df2f2a06e8b681ecd8c88bc4a7
z1a88d5374c2f277c2bcc1b6ab842d5a6e32b546f4abe009c9c0ed2b898d185d46223cb6ef8135d
z979611c9e115ce0beb2f8b17cc5308bcab5a2b01a7039d89fea4dc13d8d990dc50f3180518e8aa
zfaef674d6130fb9e88739f27241495bc999a139a8801d6a8b9a279dac4c08dbaeba16e7c0a3057
zfb0432acbcc45638a8ece07b5a8b2961e6bd3a8a18170b98a4e356894cb4c8e64f536b865afcb8
z7f5add4aff57634494a91189fc16acaf3a2eaa1b62e5a0bdc24bfe6ac797c282dee38e00a5b15d
za90ad6d811fe0c2e687c0fadc7e100fe852f4db9df104f9f5636d06fb02f18da41ab718c21b93a
za8dee429d0fdf87f1cc08a0a7412d67dd0fe729ae72f4cac678e4c2f17b5f66b657355288e819a
z9fd9ce28e0507a3db3ee8ec62bba7965a03274889812955c05886af3b7bbb02f860ccdc2d6b186
za605369c76e82572eae68a485f1309dc37d5b27063dfb1ff77296000387b8cc836947ad6156d26
zb6037f5cf0d1b121293080855b1b480569bec5a9e8e3fd4682f6eaa8e8ce094a68d529eec9cc73
za7dacdcb8b41d92d5cb6b337a99281ef65fd09f34e330140cfd72831125f02cf552b7a08b319b9
zae0b6de51a4ab7606dd7acc6e2c1e907f12c17dcf4a9b75012f76f2617caedc3bc0fa23a5bdd04
z8771c4ba2d0ce609cb02fc2e9602733ac2fa5a3d7083814f9b829d22eb0096d38d0f6f48f5db70
zb5a0f78dac62c79c04c324deb768e630f09296a7d4c9f7b6959fc80d38bb65851714129a84e6a2
zda14b38de5eeb2bfbc6043a74a5f433cf7c506d22ffabda03ea5b21d44d6bf404950caa75cea61
z0da13853bb5cdc8013609617667142e0d2cce0abb90a5013621e87744ccfc0fab02e7687a9cd9a
zfa628564cd3652e418e4c58a1197d1e088d6e72faa2e78094bf2655f45d07aec5c1fa0713cc56a
zc164933e2c8e929559ce1922c284ca8142062c63159a8e295ff84d6208dcc7a8d75295363ab4b3
zc4cce5c2be9a17da6c5ccb654f18286debd1b5e21d33510f774e007b48a9cc94728832794bb21d
zf5cce2fc25607ff9fb2cde89bf3599b256ab586441080b356480104e099782908de9925d271f28
zf0fc23e59cee6f9d3ec0fff128a6d7da8425f9ca0fb9c081d92f9c96c7930484310f3cdc9e1a3d
z8c6bb620f020116fd6d14b8ad431082a07ffb84e2d483c5dd44fd83ebd4f1339124ab36a6437fc
z006d7049f046d5261372219a70834dc9f7b5a37fa3ede3eb7e8ad58ec0e5ca35a6ebdaf55d5971
z403a698a03bc0f8abefca553a43935edf0f77759e2cbb53e5663c4710d22b2a3de31584dfa16dc
zb812ac63f2d1de0bddb920b2294eafdf992cf69249c04eb77472af399d08fc8d2c7e16904a29fe
ze8dad21fb7dbe95f9c30a6923e6c43f79544972457bd5d514345a7d02b66113034a149230d167e
zcedff6c5e5f170b18b7b3ea4c388a925ade92c1ed46061a66b69acdf4f85a4a85167b490526918
z00f59472682de4c6f981d030f88b5829fa101d03c4e2cb931a606fcb8c8b2b7b04ce0987856c48
z4187d2f8c9fd9107cb9c3d9a388bdc1fbf79228cfc3527cc6d17d5a50225c26c3a0e002c3670f3
z3adee411c3fb389e1e79a63b8ab03e2b90dcf0d1d9bee8e6d2d6e30dd03db3689808ed16d64f16
z8fe5712e03d4dba906e80a7d3aa2f09a9b39e44579b6f25c728bb08d841a2d40fef3481d776d0b
zf509358fc8d0e6bc9003b277adc10cf77d354acb52a46f32a608315479c445238c17e2e4a9d46e
z1b52ba254184f8ed97b9c0d0611a4dc276881a1cefca03455b572ca2faf05caaee0931b3280c28
z6d3c9c5c1eb470f67ecff0d0a4a6ca705874989bea485821ebbf5afcf54c649ac72735e1307579
z17f34792c12147ce868360e6028f2efed9fe422ac5f5e7810e11766ee5e2d1a4efc4bc5ed60a0d
zf40dc610ec32c36d5e520c40a482a9de38ce86a5e547f3664f18e5ce316e50b3f582e00ff92f0c
z151c9581cad5cdb22852ba0e92f4496beb700e6d4d603f15dcf0183f3c007ed9d261abfed7a7aa
zeb21d65886485923aa552b791be6c437732626498e99913784ab08955d4a5fd59966fe4ea196f6
z33f4442de1bfce04e6cfc45b13b807deeeace1b9a2f032bacb3b871b06e4e0bd853ecc24f15007
zbd4e9024d297c6f6d1c555bdb0d65196ae5fe662f2d8b699fefee7ffcdf04a0da9bbf3b8fc11c8
ze89f833148f18237f2dd9f3c7bac9d96b05d5c00bb8fa7aec6621b378d8612227c6f1f18f589f4
ze4b814e61579b32f10e600da773f1568c381de003683cb2c4a674abb70fb5b49c6e9d3c4b4e11e
z8aa62d811237213a9745cd39ab855204d1227b5a9089bb438b04e6792194aa2ba98243148f6c8e
z84236bbc95510883860c210a329bf0af0b804601e990dc95c5451d4ddac737abc3ace539bff0e0
zc6e8c22363acb59d40afb40c8a9569e6ea6d1665a2b66beade755669657593534e9dadb7d6aa92
z6d5fb185d1a35bdc38c405180e6842df330696cb28b370dccb103a735c32171d774c7742d6769d
z7c25f638aa78a7359e7a634fb85d8472283309f7b5b351b483fd3fb24594b5505d4b4e4ba14d77
z1d0d55c279131e84fa5e2131b8a0160e3ee1d95441f69de7728317ba7c32200e59f023869fd9e0
zdd274bc7b05796082c0a555b76515272be20c68fd912a660fd3fe79f4a9396bcbfd47f05f9ab1f
zd41867b0e3ec74f5de3c3bbd33152e0d6c29614debda8bd6116ab8875f3ff318b806470ccd2e78
z3ff837286907dbb3d1eb5df3d2f53566bb70798ebbefd2c2bffd8be89f79255e48fd4b9c15b3b9
z2ea20da56315926850adab22ef986c5ddf5d57ac21d14a59b244c9db578b7fbd0e27711236f3ce
zd969ed2b777ad1c99ca04cee76a9a9609489929c3637c412594c61d40f7fc50b87aee96e069f19
zbf1d92d28e64898d28806eb64f98bdf7346b9bd083e40bec2da973138ef9dfc26e38c66d96668c
z7263d317c91f13e271f6ba3e5cc93be4ea6c819a34216d944063ff1af4173f48a2e8681f6ee65e
z9bab7ebd49ffbd1374a656b18f3a2b81bf984e89ca0e7e89fa11aeedbcb79bd08e2ab6084622ec
zd179a8b761e3fe0838d9e957fb4a0cc8d68550c20164b06c36d428e2cbcd0dccf23759fe51d470
z1a636b98b352622cf9c6245b44296d8cf4a81a300400314f7bf9d686fdd5a7d6555b0d11762ee8
z22e7ab532bdcaec962dc06fe4c2f32f1c972c38f5513b0d4614d7d6edd51085b99f842cd15366c
z4ae503587c8fc3e058b6b93936a7ac354e35fe37dc2f7f414269390f83a41198d950c55d89903f
zf3e3a9ebc24403b0be6907c5ae7843712546605d451a4a1d92d14c1b85cce6c07222163ff89495
zb26876e26df2039bb58bc035fbb95a25a26a49cd8c8c18a2b998fc712916273f1dffd20e5aa69a
z57cd3e3a07d8c934502a000caeadbb180bf66c95658583289fbb0f9526514a689dc26d090101c3
z87f9f81f5634b10d8589079e62dd90207baf5b788234a0741a1f9fd70eda60dce68a9b08fcde08
z094281e1dc0b7c0ddb09ac97902c103e56963838f5de03f5b5a0d269079dc33387d3cf861ea3fa
zfb5861d4ec487952ddafc2ddd9f95da3c02a15828ef1461db3e781eb5196edd8f5b8d7317e8548
z6f96db4cc916bad2e8ca7e6e7396cb96ca76b30c6d0a92ce23cb16fd92c0412168a7dd6b93613b
z4a27a3516a291ffd498993efbc5a594a1095a40514f9b3a95050c18e70b286329f34e1d03dcbf1
z11eb9140519afc33997e7fa117907c28f64e682fa0934e16952c2f4763be6f7608400fbc522952
zf8848c9e31e66b9deb0a10eb32afec9640578661471d12b51476d6d9f51815890048b129557a62
zd43baccacf1515fc51e9e0d8c866e56c3d10a1284f017e2008ef587bdf833106f9c7a9d9d8204b
z8ad12c26039909cb2fcd0b57ae5be8f17e26db810e564cfa9c61091b31f758cab18d5e53a3cf01
z9179e40da246b4e3786c74ecafa75e9ef54a29f61af6045761979495bfda8f0347558c63ad8f08
z088419ff19adce2c76005218d3c7c60f1b5f93919e6187ac5b8eb5a39970ccf593220b07341726
zfedca2d5e8437ca10aac6c1583f5664f9e92810ec43e357254df14ca25915d7fdf8530f40fedf9
zcc153abc1181e652429cbc7ac0befcd0fec55c5f92dfe833b9031480f6ec7413c1e769b65ad9ff
z120427b43c3422d554b9409db1176d50838e323f2cd3bac6f949fbf013722d5b04ea35f5a69f90
z8d269e1c9a921ca0ee92bfe229c4fef8705a85ff5b364c898c0486282606b29cbe407f9bfcc6b9
z18a4df2035843676fd5ce13480a7c67350553a0c70482b61415a7c5b0362ad3d25cdd4611f4606
zef874dc34f0eccc0c95051930825e76fdde5e602e5633a986d0120ea2ee808545ca2794497bd76
z3a56b6a5a2405e6e1315b1d136e83e2a1aefc7dd8fe44c4059652087f18c89458ed41b0837adb4
z4e8ef641d668e344121ebda69726fba8a3ef07ff77942958dabe11f716ed9ccea06af6fc4db616
zea5233543b7ce0a42c4ff8e6c97bbc7c02ca5e23b4d88e7254f2cda0ef4ae0f5e3dc9eb171a2de
zc4b6da54a31ed0c4d576645dceb8ecb681cebec03c29c4525eb3b77e42085f1b6fd280623a8b10
zc8f976e8132ddee898f1e494e90f8fc9c22bac37a50de0a84c56a8f5ae724444f50863f75faf87
z323f6097647e1af9a5ffea44a0d6e9d219b4bc65122163abc48b220c7c54049bc6d04c21703b5b
z46fc74f86f48300aa6c614261b88890f5ab108e226f9d0b6a818c9f805631f608540ed3c21c7a7
ze2faae28977180992c2f439be5ed21f76eca29b872438670169bf60bf93a757de5182a64be09ba
z8e54c127035a6ae0a2e8f7daa016b15f5fe51c66037ce488c10bb7f8cf840ec35c2bf8581f7700
z11177387f729da4928d1d529bfb31b50bbaccc2fc70efb63a6bf78c1afa7be648deac07989235d
zed50c0bb07b8c9263617b9c15dff174c14fd9a9415d62a205c66a5ffa56f984ab0295ff1110245
zfbd46dd6503141635410b62adbf21580b13cd21a4798896e0a6560a8017b4d1145175eb2d63a57
z33d8c58ebca653bf230913106a3f36f4619f41bafa949045c6d66d26875b7942930fc4273b3ba2
zfbd3077fcc9a8915b1c5db20c9a7f80772d0ffc7dfd2785af0021d34737cb5e6e6395fdd8766d8
z9a4ff06d71eb9aa7aeeb1459318bf0610d00af09ef629fd4c93cf251d70e4c6bfc4f8951e558bd
zfe00519fb31a0766d65bf87c131ead5969550021efc3351e238edb5ade50a1c4f980ea0985d257
z7ff3e15cbfc4854d268239d6986925ad0cf9c894594ee6ff44e1f7b7fa2319491b430e2e6f75c1
zedad64c43b59387bbe273c53233e887d4bfcd943e4e5d36643649ec6bf6ce3748a9baa5bd5fdd9
zaea8e18697b43933014149f0ebf9f52ee0a071260e93326c551a3d0c1140465b134f000ef204ae
z5e41f1aa4888397764499b58264e072baae51094119eee1ef7726ed7bef61e08b76b1245faea87
z1157e4d3a15d2d238e57de6860724cc9aa802e84233fab5e727b3a3ba70853933437aa80f83461
z1286b64d22723536c243c2190d3fa1d4b8e1280f9cca91b4ea4d441c1e7996a2526773ce176a88
zdcf6fab3a3c7cf7597255bffa13d550e2cffd05714fae86df9f8dbfe7617a7234fff7bac77466a
z075a4d9373ab6c713e1f544eca6fc9ad2d5acbf56f0f4111641dd9c9a989f974e3a2cfb169ea24
z12b8ef88ec012ac9a012f3abd15b8571cf540ded3342107b93c6e465c209813c3a8e3dcd0fa4fd
zb7fb674f6ea04fcc517551e2e272096617c3a618a2242cc327a0c04c90581f737f34640f49f7a9
zdc25e407162e8554005fc1c91b3796309a3b95e0b854e44c154177a26dec75379b5873644a30ba
zb98adb8fe509173bed5adab790a8684476a873bf77ed94d96eedc49307483b9094b814e6d8f818
z41ad3411696939eada0c2ffc7f54d7c7a9cbca1ad5718b7a5c2d6c0a831a968f20da49df819a3e
zca67152d693f79754043e31d7d56ce3664146df4b8a26643edbd18ce3ff95335d137544e585345
zce3f941b1f236b007d0b1fa9ee63ca9dd43857c2aead968accabafe4dbc54f86d41ab99d5a58b0
z02eacae5ba242f5798bd1ca14d371ebc193a910f04c59076a365481d41da52bba0dc81e7836d64
zdd17a84e5d712b02a10e4a9f8baedbbbb04af2b3f9305c93d2f5e94dc9f824da31556a52ae8a08
zb87e5ce92bdcb1441a336d180bca246f27716588a978b93c25d90a8fbc15345072adc97b89a6cc
z0252ff45de99d0daace5ce525741a90bc549598b778c766853a45cb124158e8eeec0d4cf3e9436
zd8fe0d46e29fe78eef6e3a4afdc3cc644e2ce67b41ac071af0a672f74a8bb32f409b66e9263ebd
z1d658f9cfa0cf2ca32cdac2d4001e0bacb6f97da50ae4092182f5f48bc48f04b6ab4bf9a874594
z9546358f8b1ff96cb1944fbabc236968cd47f98a7a3dad9e3ecbf8f5f4f2ac8c786bfb37818c4f
z1358ef092cf76f0640d38cb09a23552ea9ca8ea1215d3a9ee4ca9659714eef3908687eb08384a9
z27b4ae03dc2ce4631a1ccd4329bc107913837a49716037b292116afe247c186efb4d031b8803e1
z0c4e78c60ed9816dc8e060bb1abb03f7985a9a6703aa5c8bcf6801fb8e02fe456e8798c5515d8a
z399c7267627a9181df3373090178b692405e000b170bd2d4d31db81def119c880cb17d398a5eed
z45aecc0f7126be909bf8ab6cf81ce1551b5bf82afba0372b94be21b9754b6e521dd644427991d9
z33ede3c7a23239a948cf9463a8c2472c006a91224fdf12993e2874a92a7c05ccd623b184839766
z7c29853d9b7afb12422037bf1913918e5005c248b6d8a081d1ca5b9e0adcaf68769d631630fb1a
z3d2c4200ae67059b9cb399ebd516e53fddcb44cda9b3bbcbf6016a0e4e807d2acb8a23cf1d6d57
za01b7eeee7be4ab1a17d474df3a611f9fbfda384ed8382baccb84d0faccef2292a5cf2f9f93e8b
z280f83236dab0d2c2689b197df04722f2460a09a6e5d2ecc87bf6eba71b0a09a8f6a37a5e59e59
z15f77befa871f584c34f31e6cfd7e84ed51c1394e6cac67dc9bc1cb12a2fa06aa9f3fbb35d9cf2
z7e06a35631f31be3c45e988320b5542ce681ece17d535d09c2b32d18676b8c3d28f4e2c6445d9c
z74c7290fc6e584ad2c7288f0cf133a1f2fd3c91739dab1f53781bd29b12d57ec03eac624a1ab99
z207829f2f06fdccb0a83041f4807fe31d279b07e9995cec4fe6bdce9b653503ade337905d6034e
z16c49614f8b8ed8a3d7068f8a2b92cf6cfffcd64fce7f06f619fdba13809ebb06def243caa7efc
z755bf7219b0417dbe63f190fa867637ae23d26f1a82fd7061319a8c37e54f00e2e90fdedd5bd25
zf8e43b0ad3d6bc9fe55dd86d8a20ac18ee0c8eda5466cf62ff76c8a9b47ca1632004d5284d5a0a
z0d6010d1fff2180bc418a52ff1b579f571dc12a800f6e6d9aa9f810caa81507d56c018099219c5
zb6287ed96be300746d54fb4c0ab2eee0cece7558c65c4fc144a5523853892eab857932057602cb
z30c4ba30208c4d92d2e478e463985734a2252493b8c40599b8d270f580e4837277afe888ef2922
z079403a5065f6282982799c79812d5db1c2c477dc4e701efb53387c3da7b29a50c9636caafe532
za5c91a332adbfe7f76d3d7bf193c1b0395deb3090fc216358dad9bb652b43371d216b19edcef01
z0af235bd85f1d32ed7d0a34f7fa8a90fdc286f6595545acb1e4c77ca15f7b02b2c936c567d3d13
zb1d4835fc32cfb7e8c508857c208c568421b5836e31e6a133ae637dd7c7d48d3607d2c7d9c1fb1
zb3b51f0349f6b17618896bab470431f3ba1b85e91fdd893f75291f2841cc195ae572ebc69b0f49
z46461b493dd8bf175ec65938a8b323391715801e69d7793302010bea4cda539961eda764e92314
zc4690fc2558359c200e91b96e6c38067d42261dc97d44166179f9a0f28998e3788ed678351e535
zdfd8d03106aff0136b04d830f8095b90a58b910bf2286dbf3d447bf3470456ead488c4d2449e79
zfb1026062f3c8207f3b144f41e55a040674c909fcc425563fd03d242b229201327c90e66d2821a
z3444d6f58703d383efa2a0f0be861ca6b7f653019ea80f5cc16b9b42029da3448d969a2704023f
zc0b61b18ce16a360ac2c0783b41cc5232dae879a0e98ce361cd61271d1d50f8c70428f7ee182d6
z8203de03f94ce9e09b8ea62d4b70ed73ab873eb4e23b14f7bc099bcb59fbe6ea3281c0b3d626ac
z060583295cc6f59514b0c937a37e5fafba364041b587fe6759ceb87f77440757ee47d4c2749590
z71e5075990f3da57f8078cf64668eda54562d9c887fe7208467933191709c2dde6c5f187024ba2
z01effc9ceab456f1df93de53e33536495d65f5a1291e5df110e9eba4a9abcf88521cbd4154ff9a
z4812abe7985833a7d331153ad56d3f367f74a72001094ab1cdb5345814d31ec65bcb3b3cdcdaa5
z01a13a97b05d03ee6a233df569d00231df6f5c57d23dfb7e69828c5c63f13fe7ca969fefc8219e
za2e85a2b49e6f888a936ba5887a899ef137468e3f62e1cd3812d914bc0e1774c9fb0a0f64d29ff
zf3395b3c71aaf585117b4a53183389b7ab191483e8752f6e7705566267db38395d0eec0d75b3ae
z5f385e7131f0d39360eec3c4ba52db34ecef9e260fe9931fe4983e4e2c957f7d4a133ddd4a0012
zd10cad2c685af85a9a5ae5392a4999484a76eb2ab47206b43c47ebe902f81f49e3c563575beec7
z9b0593718b36d55e49da1102f875ad8ad6bff5fc7ac49ae4507e87b52584fddd8cb7150ddfdf27
z8e36c77b4fb1c666385e8ccbde59dc78f772dbaa8be70fd7c6470b7e61bb82e045a24200be4411
z7cc216da2fa8e7b8e91030f167ebd91ae8e06d390faa4c19fd572c700e71e4f7752b32ca71a3f4
z4a190f5cdcbe0bee5b0f6f6bab2212381e0e7ee300e011e48b4742027bd900d8067bcb58ebd4cb
z909aca5188b5af0783d8437d18d514e2bfbd7d6119ddb871c4aae4491bd986c04af4bb1c16e648
zeb9022b64384dfebfb50cf8dd1c8193b9c015a4881cd706eac2f2f61df9af36f4fe1dbba525cd8
ze321d5fde8f11bdeacb9045e71ffac00deba8b9c57c15454f1c354ae8b3501b0a7ff5df3e14851
zef8da976af1fa4dac457715399363cf8bcd0ab8c16726cdf6b60c7adc1e75ee317bce3a9e31376
z38dfaef8694ebba87c7eaeacfe9fde48ac7b949a3751f75a0874c424fc9e06463e6b53bcbc66be
ze8e07a3613fd374368bb1e9903083066689d0b21a9b544f670ddf905c9c32ebf07efbdb3c9e384
z9c41a2a38a5592305844c4c670b9c77ccaee4b01fe46ed8fd5aa22c923d0172984990ba51e8e1d
zdfebeb075dce26fbdf1cec20d18321550f274e6df1e6e92980e5753b8c108f4873fc7ef09846a3
za82c41b3d3712f0931825ea71740a4973d247fb17bcf22e97091f13ec1bd44be14f4e9597e5308
z36e92b062e4c9c3b15bd1b81b480fa1d6640438eadaa94432e90870aa0da15568008bf0e13c890
z7a4d1824579ebe496d8664327cf43836a6c4901a7e387a33b5998be508a1a938a1d7c4bd001685
z527e36ce2e4d451707a448265dcbc1a69c9dde159ee5974c9c0de4e2d4ffd9d3e1cfce51fef8c3
ze3505acb1aa8cf9c7613734ca462dfb95127028ef32196e3b7f19f80bc616155301eccfc9d3204
z4561410837c26452fe16beb29570781bd6866c567527ac0bed19f7d6cd45983c4454fffe30463a
z605230471106a05786386d1c524d1aa6f01e194800309e90c8ee4ec768a1481415f686f57ca7ad
z6b358fee650bd6544257692fe583e8c4a2f283c6db8af46a6a6e0b026282cfb902aa1ac330221c
ze41aa5765d49fdbae9a75144a2469e6ac06f528a7e11435c5fc2845df7034dfb9b56a8097af776
zc6dd7ba5264d0f4d8789211f5a6ef2ea1740586edc147c1a535a07bb5a45d149a910468e523205
zea7bc0eec5c3dd6ce5783bff11e0acef77b755762f05d8783e47d08b5cda9393ee4e1be94cdb49
zaca1911a519481152936b4e90a1b4b662618399160f95e24127f4a9cc83c14141b380dd84c46f8
z531713a2a7303921b580a62b22a4487f96f9064a6159a3cf9594afb7bfcb6d10730edae3d9abee
z64c34261cf3f064d4fc83c5719ebebb80094e9c2cbd24e64fab07535a1ec6657063d4b364cf86c
z6862bc21e96ed238f4370662526125f53e211956e3cbe4cca06a45535a00eb6ae5ef3f93a04f6d
zd989e5df8d616f765af768f908139874aa3dd580cf6ce8bec9be5ec98379e8130a5c4e5371179e
z7084ba0bfc83905b36c8e03f463629660aaedec634caa50d9fa4531167ed7dfb77840b1b410cd5
z15d583bd2dafd207387212360db097d21525af3415ac9d85c4144c7f57c51390adcc4862c81d26
z5d89358828e4eebb6b3d60028afc2f64887c7ccf58d5b7593880fa7e3482ecbfbb3b964930d9fb
z4e53112320333e05d8fc4b0478c71c795939b3a327e718eab68a866057ca37dc0846cde7b24738
z557eab355510b610cef2f87505fd88289f66540e3e779cbfffb4ca73df775de9cb6110873f7ff1
z8d60adde5514274d2038a9d57cf0ed207a8e61ad457be8cb2ecf2582b63b03f93c56be4c847ccb
z77dda445acf232f806117c10e2e27c080201b702fe15099fae7294a0d801adfcb865c58b0f4786
z0b29d85a58142d823a45e16c6c86eaca5b0c992edf16e1fee719cb4ff8f5aa27a6910f0d65639f
z3de364a0f23bc3c78835eceb08daff2d6ecf2a6d055aad72cf3d7bf0ef6af988d769528e92ef67
z31e9b98cda33cef146a79d53f861b82c87029b4693d5bc0fcbdfbaef3418e06c7b60e7ec5233dc
za3257939277d4a8520e1739705d377ef139ee7f4ce2fd5a4d9707cb0c1996b6e506a0f5e8497ac
z0e05e99e8db62f3cabfb0129a189b16455f59cf9961302283fddbeeadb5ddd39e575a174cde77d
zbdacd3be7ba9076443b0adc0fef08598cfdf9dc3910279d0f2c3ae96001b6339bac9d6de892269
zf82bce1665165ce04c55cd5334ffd1c7a445d1490e4e29fcbeddc5ae5e94e749ae2fc1734108cb
zdb98ca6d3db92d6d9a527b1efe9e1157c03efbc265a8c8eb0a156243601c9350241ca00e233093
z2f678399380ea88cfc35913a4c335e688d58a269c36f6577f13184e48c088d0b3ff938384898c4
zd55119e942165fd4cbf420ca7323ea95cd0d822e3980ab489184e7f1fa275d71b36b38e7d0c1d7
zc6dc2b0a25a28613801a7a45a5abca9221462b9ca1ade2526737d5c7c0b9fb8c98620809f4ad06
z72f05383ff8ba6dcb5f89407b46c9dae37980e3166dc01cec6a8714e75c67a668cc575b9a254b7
zd8a1eeafeaaedb66fc142af4a160b9a13e7fd10921611f8413a98e89239a605eac4d8d929bbc75
zb84c2c2203743fcd61e2725ce5a92bb7089b082d00cef1de5e6c5af2fc278a8309f23298986a94
z9950a38319cabb12062efc505e8244dc6b8961aa5b0e4a730097bd6e4624f1c53a72583ffe1496
z723ccc1a85a1e2051faf44399ce0eacee8fea06fc64c0ffe1ee545d64d7cb3929deb35204d0832
z78d8fcef2b89686896f590ec22c9aff8d8507163216ba5c1ab1715933f0b64f48f9d8957e71dc7
z0b6febac075860530d62ba17bc379e66f179cb227dd8329cb28b387bcd8b4c89d7b6284fd3c5c5
z580fbec4c6103f0575e9d10152db0ab2e97309df6f7b8b5199823ab4c8159e1872bafe73a3d784
z165a3d7ada90bc656c5c2bf42e9938d92a24c00f1680f513abc1ba8f2d6c04e01d301fc3d94ca0
zd16f43cfd5a8cdb3e9a28a3a7a1051a77636b7fc10e78e976515b0884885ca516c202e2478f2aa
z53c9a1f0f72238693ffe8aa6459ddcb544dd5df0cdb8576861e3932643754c8aac6cf17ba9fe1c
z13f02713362c30ead49f0bf06687734c399252ab8cb506ebd6e898c81245109b5094e9019c16ca
z676ccd0797b29110f91b23aef8b775a50b8f871d717111880c766de125a15d1995daacfc64e377
zba85ca3218411a33ad99fa5e1026770feca6d6a4e9e943f56720583ddd2a055075fd224a83173d
z195915cc830edd66c6d5eec6adb459d65d37f3530460467b5bd3e8901143484a00eab8d81cdf0b
z462cfb661794a86195da9ed7aa6686084188c03abdfeef49c53ac819d2fdd0d9e28beabf567eb0
z973dc64c5f4c8eadf1464a2848bc54b6ca81989d2fedfeadc0187ec7c1023a236228b409d1a9d8
z196ac1e6a925a6c9669167e5a9011820232c6a07d718e8a31ee1de73d23675c2b0d1ffeb363f82
zb83595c590000d2ecfa5f7408c5daee4cdb580412f5e9e5213cebbabcead43217138fdde5b9cc9
zf962ffc814ef48385c8fe1f82c58e514e991f17cf3661cf6cc6903c21f898b260d38dc50df3fe3
z99203328a375672e680d2de10864d49ac1c9b9737a128169363bf2db1274e999b30997e97b66f9
z10cc76a7d98fbc04d11eaae339d7c6d99ce18c26b7856d5f835dc4f1e77b8a4d9e8602a1f72ad9
ze4cc00d157ed67f4059dc6c17fe4c4e4cb562fafbf04135e1c0eddaa23426bd31155afc3899ab5
zcba870c6decb7763d9937b08abbee268e0f9d3e2a172c49f38b1a5338dc6bcb04a5c0bb115d10a
za0b47e9402068df617a034d4cce01dfa3b9911fb3c002f230c1cf21a4c13850502421de26d0ee9
z2f4cdf952f7b67b5bf792bd7d8fbc7ed0fd166d931daad8f17b905ca007f8e668d736feaa16b49
z9e747d40418e3123411ecaa09fb8de6738e5231776b1921655c8eeb21948dcb5b61bb0ed7612b7
z6b01f7bea3cd20f3f12525f7de073a5132ba6b81966105e0956309baf3b8222defbae6002dc6db
z326294a41a1958885b85d399728fd08897fd4cd4e38865d237781aa632ecb63da9e8e47787fbe4
z49a49dd1d1c73729bc86962d649466914361ebfb72602e88d163d33ca9e8ff78972ef06646c43e
z4cfab285eafbb2a35f869db824b2ce47ac5b382952bb020d7b08500fc7ec32b6210634497aa48f
z1d3d9064de61a381bc47b74c3f4bc9644910ef834753d5348116e16bb1dd25bf529da828bc5e88
z3459995cc0bc6e8803a330b95423d99288187b8a4f10f57ad6e81ba1cc8fa9e8331e76d458fa8e
z972230b512f11c35d878f47e1d9cb0b225b836d23b2e110c0e90cb289bc5af23ffa0ed37b7e4e9
z5a44f751e0d18bda152612e94a10058b47701898c573af101a31b4a579f0b1e296d0393656f1b6
z4e9ada085e23a1e329932f2f0091513885c1d5b3d281b51436de4dbdd8453f71030437dd1c28c9
ze63ff5cb0168a7db6b7f8c59a065abe394878d748e23ef62da568938fb4a3285cc6432a5b9a16e
z1464f9fb29154054a91b2ca332ca05df4c04f0e6cbb4c6bae091fc622d0c0d838c3a02ba476945
z19a893f00d89e4144fde8111ab247960a6bc6dcd5083abf43a86413103180cbc5d1968ecbadb94
z52cc44dd8061e2ae994d9f65c65cbd7c7f299458d470a40988963f8b033de07f8dd8980c8f24e6
z2bf6eac886b63d6d5ee5ed63edc3b59cebd1a02d5ad06da2f9aa7061250cf801730f2734ed0282
z3eeafc5062823c6b565f9499e45b16e1691624b4c29afd7d47bac111e7c11ec73be116c9e105cf
z5c3e4708952d293be8e77829ac69506374298721ab7a9aa298885c9061274f4deb0d3f710dc95e
z815f058d710e480d084632c41e716cb92302b85373be329d3a4f268698af32a1436ba20c5a8f58
z475b2a8679dd68676a48f5c9713753f8d71fafe630921abc4b96ebd5756b4f2bc84f0808d7b62e
ze9015872d190decfc9f3c7f81b917def7c616926b894938bc20e93697891dfc6880add94a9a04e
z9d8bb3df98a19ad31f83a20840fb0142dddf71ccfbf843ac11f5bceb8931ae427d606426aa57d1
z1eae81ef7600d14a597564562ec15b4b44abc03996a3f0382a30ef8f268fd82d750019e1af472b
z31273b93560f88d2d21728d8bc98fff7cfd66499cc3071f07dc53092790678a87a51ba55a72724
za796cc627c17423c999c160c78e02ff7ece25174c451ba53a236b2656ed15b228446068bc41d30
za5b15bd39aab17931ddf605cba0f0db716afca6b28ffa1e6f68d372b86bbedcf0b1f9f952c2aad
z848d66acb1811efa7b14c0a8c40bfd10164e9fb34834863bdcc7dceaf2301d79231caf30d3ce20
z89c60b016e58aa8cbd7d67576a302ba83a65ccb0db1e9208b2a347710e3147a892af49ad234f5c
z19e1e28ea6aa13497babc53cca9cbbf0b88b77bb3474b8c2d8771688e1aeb19c65d42d24e2c0b7
zeb89223a3fcaf2b99a3e753b04eb1f7f6ae1628c503f5d0ddbfc3dbf17a08d22800112d126f24f
z73bdb57a026f010ef0af7a73ce4da6c6ed872599df39baff6860ff87f7d8e9ab8c28fbb47d727f
zeb964725d218b19969de0ed96044a5f3ff2867c42ea5679022b77570bf4fe9732f8924448ca37a
zb6b800622b6661a1dcf693eda49ab5a9aba01b07f0af1778d24474c0dba5f1f0c994888caf2f33
zbf22be10d30a37f0134f3453f61102755d113923055681274d02459d0425e598e85210cd69af17
zfe5ed7c22bc31c482f65f6e6262fde4dd0286f472b3df02b218ffd20b78419f102223bcc94f504
zbdee4a0fd078413cf245613905b416b4559db2d0b783c3466adc3c6e46f5698ba6aeeb84a766dc
z93ff9c7a205738103b4df0b1e8d0f4aa0257d6e628b063f40dc4f1c653e77e4d46b2c9bf96494f
z97d66abcf24ce753552bf2e6542dbcc2ab1a00a7a022daf4530aaaccee9b9785171fd13bc974b3
z076769bacacfebf04d90f67e7ffa0f05321280fddd13341e98faa71540a7230e7d097c51b10230
zd78e67990f9785b333446cf6dbb61798bfe5d81de485b1a81837f86506176dda58d5d8c50c7a45
z37dd607e43bfa4c3772a86ac027bfb6f2e6dc35d36598eb4fe267592a20d2012f5596f4625f772
z00aff2f7cb577b0cbbcc244f9e8b1c0ac23309462661aa137658f07ec6ae7e5eec2e23363f1edd
z1ce005c62da72bb1dba93e8b73dfc1b04ee09655629abedabb2d6c30747c9fd1ee112091bb7ce9
z878a4c949228093bbfc981a537bd6dd93185f984e10a1a3eafc332e9ead2fd3dcc4ce53ab4576a
z14505b721f66333f88083b0f01ce3ec257aa9ffaa5067dfe15b9a96a29cdac495ec9bea3ec35fd
zd3fd731258a3182f65812e7edf8d156492bfd4954510641ae12d74fbb4fc941ae58081187eebb5
z59ff9a8fac33dd72aa49313a38fab2fde8e8001fa8809ffd01734ee888623051a62acb7331f63c
zbebe6260143a399e63b8f4d8f95b6bd8f815293d0684dd8d11c4a769438a4b1f1cd6373782bb35
z0a61317a8d92b658918068c5efa8a45eee3c882eb2c25a1178da7e16f511dde613d65bc786c5f8
z465519b53ae05d60f0a1631149381797b88f4a9a4a11f4dc78df4cea700bc958c859b96e7c5d09
z1142dcd2f8ae431926aeff9bf7fb16f0ef730cbbde8e70fef1cc1e1fe162dce339dac6d61368bf
zd7d58bec775f0bd5ee59b2f6c4cda20f40bc884273bb5c9620ee08ecbda6f3844c0566ce5d3479
z465ce3594edaeee356572228f0f123ae53adb61f2fd6a94d8ae4ff2f52e71baa4fa335dac32cff
z5cd8577adcdd1045e3d636acaeebfa93b05463a19170e88030a431878159a0218d2d177f4ec2a2
zb75178038716ff78aacc9c01b756c110b7a279999352876d87e2dd7dbc5e616cf046a2fa9d1b14
za70751fb5b59993c99db81fbc35934204cbb7f25c988c23d951ffc0d22fedace2c521c18f74133
z816cc10591d442fb705b5495bdc76569d55eefea797a10c99b4b272a81b33874b91b6532b9514f
z1afb349542dac7cba2b957f54dd4a20b992dd62ca89eab086f08ea912414ffaa2e61668f2bb628
zac945b2ecb3fb1730bd7b0bc4e535d885dc0341da2f7449bda719811aea6f66fe3c13da02ad4d0
zeaafd3bf73aaf61c1440b32a3610ddad05d17291ec57109951ae73f2f2af354778acd1f0913ae9
zcc55462ca834169e1c809b43096b60a4a772e1000ebd96198bf1de32d07ffe6d8cfa845b567d01
ze90afd7d7fe6226b77f756382629a8329bb4676884f5f493fb4b6bb392e0d81a52957e373cf157
z888230b806e5cf7d8cc16d0296199800acfef138e5b1216e9c86baa32865f3ee1b52f3a29041fe
z53eef1927c1c645327ca36cd2b6f37150b484ac824e22990147493cc242aecfa5e948d40720d44
zd65db665bc3904f05d8fc959f37b78afc6646b1d6b89ea7ab4a7fab0b8b75e01506c0883930f08
zc824b08578630d7ea5e39bd115d0ae05a40006a5eeda7e2ffd58a346e90e8d9839a108951c944a
zb4e0bade2dab9cfc97877891b9e956b3a4c238c78b389cac16653736c7cf46b703ab2f07575501
z316129aa3e9d7589c222773e92b0d53b71b728e5210c292e1950a1fa28e6520cd3205d5c75dc4f
zf3233365475e38cd35ca59fbbde78f972c10e32903e2cc2862600c0055735bf61768b733f9b40a
z468521749aff7f155ae78d2f328ac632a0404aca33412217e437b7ddfd13017783acf2862c043a
z79f4821a86019374729a2130c25a6110f1cbe4bcbabfc56bdbafb14dbbdac5c9bd837125d9e9fe
z12ccacd8cfc55a4080fff91ad824565014bc713a0bf7155c33c0f25130f7df693c8073d31bb77d
zddd822c6e458109179ed7f134d8c0ad33a423a201f26da1d25a0d42e6ff605fe210b32d45957ae
zb936cb3c981fe6bed7c0a5cb5d92c3b4e3d85a72c766c8e6dde56bbc30e2628fd4c6f8d1c9499b
ze84909ee851d7255a6821af5182d964550060b97119530ca5bb393b3cfd096520bcd170bae59e9
z8596c086a8433d0e72d8b4abc68663b8c40c16af5ebab44045ac2f58db52fc49dec75dd5b2d2c6
zd7928493823055c60cbb1ce5d71fe3b5d1c69626081958d17e101093013f43a303efc982459d07
z01c5e74f2b6f2e1c0c2e8764a34e45626d8488de8732c35ccc55a059e4dbbba4227ec98ea2ba8f
zed143cc0a43c8d389cd9e5200f249cbda2bee0e03bc44f75919dc2136ee9f2b321e9a0d604f2da
zcc1207700696b9df8534abe835c00a0aa1bc686e96dd2db9a8e75d184210387eff1873cb7537b8
z14ee5a8969c090b583f22f9ffea13c10e0bdc8279d02403ef52460c2f1b9cb2afe51d70c54dec8
z9cb201381130fd2c476a035af19a47bbeb0d85c351bae236661f1bad02b407e9389ba7a05d4de4
zf62834137293ff489dc44b0dbaf8af52864b1c81b7937f4ece9d96f44fcfb6acd65183975ec962
zad6428d6c8d71a6cfc910ed72974e217c204adf3e7a0c12f981030bf7b12f57db2370b9c1136b5
z783b333c8b200c18de262137aabff81433432868797ebe39976c7c8434da4c51a4ddb92525e21b
zd63af8f3f855ac2b7e43b652e662eceff4839459a106a2326443d94e2ab2eb04482bd4f8284583
zce06039ec448d32a50c084c76f066c0c7c34e4346f45434df5458660c2cb9ad89898baa2c69511
z9dfbb32913f91ea9c53b9ee23d4c62280680c1a01834c5934a97b246e57b1afd8824616496b164
z24927990a1863e3aed5222845333317888ebf4f97d677f0fea54c91d503a0f42dc2f59d69f2df9
z14294ce19aa792ceafd3f824409575292e51b52c8da155bdebd1e67f61d0e8bfd1782a24d9b346
zdebe1af824bcc9133e356a133146cdde6b3966ef60f6e6c6108069af76e9d99a51d65a61e3850e
zb03ae673d2d17141d75531a14f19ae2a4733d4ec2bdc09739662ec080cb65f8bf619621cc76e9c
z1d84209bfbffe7fbd365ff8ac72b166b5e8fe3847575540013833a2387008232733faadac28374
z76d274dbc80d2d3f2bedb0dd24f30c73cd7b68697e1e713b914c7006833c56cb9c9312d1556783
z4cd84dfcf17645f7dc52a108cad79efc2e66a2c47edb046fd6cf48718f51de8ca8ab58946d722b
z8ae95bfaa2a3e8ca1c88d7d3c0c6ab8131a468e2ac7b6a06231ae5cc621c4d6d67d44de46c42d4
z8b8e666af33373e7d726c7b4cb6fc7bd9dc22ed56ec2e29f69901f4a5ae1766d0511bdab54d9f7
zc8ecd59f1cd3fa7016ed56293e78c3f64d37d7a823b5d5523701caaacf2512eab3147a031d2422
z659174bd42eade75383f25f7110faaf33828314886baf8d4110b02fff562c0b85095f8e861ed59
z000e802d501a17fd1a62995cd4ceb832c3089a8b4a6420be855101e54050e8804aef3c7b1d4d7c
ze2bb188a05c4766e91ff88e35fd0c6bcf1e2ed7c36844cb0be3af2d18fdf354556d690333d46fa
z8c81a8bf8302bac9c92d340d3336d0b886743e3770ac201a0e1269e9b1504200d71ce22dbd6172
zce80557ebd9a8380f2be5da5259afec9df06f1a16827723aa8d43d16a61f39e4bd7ed65ad03190
zebe47337d8fb208e30cc5b8482c251ad781a06bdfb17ca7bcee25de05bc6768795821297c4d0a1
z2329f81ca15ac84138dd97a3aef90c58774d5050d3823b7c506a954202f8ce2c5dbcfbf5f5826f
z8cc2a8641e143044bb6abd7c47179ace942b36d999e2957d76ebbdc8cd9d5c505d235a4a351a47
z437b4605fb5cf79399e41e6cc72149e5b63cc063304c151af5d51bbc04140f870a5446a93bc572
zdc94c9a20e0b3a86c9d9c701b72a03878930a99a9dd140183ff0a8ff36d0a8595bd99006c95d51
z50377967f648cdcb2f04765b240a4593ba70d21af27c58c4b0967740032698875484285f8d5b0e
zd06167a23650049c57035586c41a7f07d26b021f1e2ed5cdeeb59c0694774a72dca3c1ed818a3b
z889f19b1a371a51c8588eeface02081a5ddf09444e55c2e400cc69544e4cace3593a6fafaa92e8
z25211fd64f90283112a1cc525bae3741ba1ad55c48a2818e80277573148c72af36116580072ce0
zd76d434167c146626ac5d545959f7d9d31e67e62a1aec1658aaae8f530cdee6080d5e34fdcb8d3
z4c6619eb163477d94585d21953c50b67186ae4a71f037bb6bb4481b03096f84268bf2a5ed0bc5e
zfd75f60e764152699a6ecde78f66b5909b00e448432d5eaff5979758198d9d6bdca7e165a74508
zab907a1a01ff5e3704a61159c9fd8fdbdb13bb256e18fab4bf62da81e59514558f45abb979585b
z72462d2ebc72f8f69d8de8dc03e061a10c8df0eba58e8038831be31f8ae43a3cb3975c3bf7ebc5
z348c925ddb0707117224885938140afbad2402eaa5dad6f120a5da388fcdb2100d7f61d0f6d3b2
zbffe7c3edb9c89d9ed3cfbfbd7befb4956daefd8f0dd3a3d90374f2e88cc51224b3acf98c52485
z183fb487bbe226c936a8f5202e29d2b68bb09c1c004302631fb20aea5bd66a3b8d1b75f9172fd5
zfd98759bb949ddb6e5419e7c6dd2fa91c1870efdbd2871c665af0a8ea28ba7509135beb1e2b09b
zddbd9f10524f5f3ef198f02e29b91c41ceb6dd8c6ad36064cc44db5f8ee32a468d314e2807fad0
z9dea2b76e216b56bd8aa623d86af6aa1741572a259b4678854f20df6abb8f15ea1f45f0d2e53b8
z73a58191204dad250b7350d70bc31026d19e1d7435caec4e39fa6cb4915c4f8ad35ccae82b23a6
z082b5a638634644e723264e6af2247c0c209ebc609ca1859477543885e37c8abb0d66c27979fbd
z9b969fc8294c9f497417122c6f13695afee287c2b12c5f02ebe643c9600d11fddf4c6dbb756826
z12d3a9ef07765e383cc26f709fd04066e0290dc0c689cb0f242f451e0f6f0b4343373b0c1e742b
z68ec90255a00ca4d393652159731532aaefa4c0b3c838261be5d2360eb99cf951a4556e0805cb0
z0f6311e9c431e6ac2d09deead73eab19b5ca4451c70eaf697b836a129bb9dd50d77746a2caa11b
zd8649ca295d8485f61e5dd7efd3a01569407c761f0f6ba016a12582a84a078a2b1fc6f9fcc4299
z2f7e21ca9e3461f9601a9790d989b825fb1236600717892ff0037610e2026ad472d8450be243e8
z58874a61e616f88d2fbcb6a1bef6c82bdf8ab50881ec6906a04e51f91d487c004af56b1de6561a
z44450ee042ef1c7057ef556087d4620e4d810f6b10ef7663eb12f7c3cef9343afecc181d8600ad
ze5445c03ac06d8443a2602ca8f790a0acb3d2c17ff7b3729e5cd109a1fb561265d18217b2e81a3
za126abf58d04267a7ebbf9caa43a1d5ee6f8554bbf4d077a1414cfce9e7e195dd8dbc7fbc2f242
zedc9db3effa0155791a6665024c5f9e8a0f3e8fbfb78f6fd33d3a3687e6820b57877b59a7bffb7
zcf9a834e113a4c756a1e9b0cd80135b67b0157aad3f26d0c0eba3fee4492cc716d6c45b7368485
zd473a97c8366280cfda375398b08d14a32047c57aa80b7fdddf56a9fe0ce4f94c26f273f4b0ed2
z7afaf25560fdd5f6f6a9eea810fe8b336651e09643692a247e4c0504f4899b5fd3c312e3e36633
zb087a98f227fc85ca0af22347a0f543149d2ff27e8d035dd3cfd213100f419357198c6cc6849eb
z65d0fd3404ad1c6fae65b2978631a0938a0fce4b8fe1bff3f39e4739d7ccddd4bfaf48e07e13ee
z7288e6b63ea89bf7f745d2fc4e5dd5cac27aaa52fba2513aac176d72f201f70d9321f36ef04e19
z95a142d129bc59e38d1b149ca45717c50b0132286bb73518281670fc396d0f9d2e0bb924859a6c
z2217549a58281f234b6164baff6f17d171e311c566d4548b672bde62258e297f4e51496008d2e1
zf6f179943de4ddd9fbca7d9cd8bde9e90a1b1f61c0120a63df735e46c891a3f88005b2bcfe1142
z2220461d23c5bead6d63ffe7bb0e75214b065c6b8fd06231dc3ccb62dc91e5c54aa0bac28fa1f1
zab56562e43bb32b9bd403533e500777ea2d79992172c59112476c6ee19e330a834521162def773
z2b6d3ef630268867acd29eba18b9034ab5ba7829503fcdb295034e8973121b981eccc8f4ddff1a
zda86f0a2b5734c7a669f686bead1bee8efc0ae921d4716aebc6bb3c5d75447ca8c8db87928657e
z1159061d7f88122fe391ef8eff0109b119bcc7a8f3298d899e7fa14e22016cc72cede51dff5917
z24295f09613ddb628f8e6ba5645f8af7464aeae894fdb150c0c69a1cbebaf5efe317cf3fea4089
ze4e51f2417e11a0a5c9f202b702268714dea928d7f16d5814db2bf245d213eb0ca397736fd7431
zb566fd9a21f536c21ff406d10728ae4ff454d8e3adec64e65ae8898977902f478a6cd43f52f87e
zf949467ab4c2ab0a0a2830a0adca64a755e4b5d5cdb52f7260ae0558adf72a3c60367a23488b09
z3af50a6ef2f6060104710e48794ffe9645b03e3ffe1e41fc601a1d417c316df7fe58013df9849e
z064678c328a47e227359cb74d19eb7cf279bc2c5f86fa225f15e81afea87d4a3c4bc7ebf8c59e4
z5bf1ee957d62127afcc975ac9f62ec9c54fab4043f2466fbac150bf96c14284c796462ee46e7d8
z1560a234de30c68ee610c38a5ea2ee5d62ddc6d05e187e4da090e46afa91731c70bc90115f760c
z3a2949ed0213e2a8052b527e5f5a8019ebde5a7568021f65c168f766db4685a66cc7fbf0ca468a
zf4e2a0d0078f6abe57668cab11669d8d8603c2aecc9ed5bbd10f0f4cff12bc6c37ddfbb5c1e994
z88d3677926bbdcb8113b3c08afc715470e77ff5c6360c32ec01d2144a5d2d3ca3d6dbb0f6239d8
z8e6050367959b4dfe6c8a4f9616d337ca9d46becd3a8df6faf9d58080330f3c6fb34915a2ceab7
zbd77828db7c140414fcc66af1ba553bbc7e7088fb7e1407cd939d2bc3d0fe340c934c00044c81f
z6302f9558c33da2cf3ab9a1da7370fd85d4f353724a36419b7de48227783471e09c198fca07026
zaa0105de175d3d94773337a656bd66dbb6debfea48edb9057a56ac29479dcdcac8a81b0a3bdae8
zb04a102046286d3c28bdb8b36492d262ae47a503a0e3b1d0c61c41e662a894264b7cde087f323d
z3761e1e1f9fe90bdfc1fb1e2ccaff31e2dc5dbb33a0fc1f5984cdcad5a159e85296488d5634a05
z215adf4f64ee64cffa764971e3a65599a072517e2f78bc39651402e5cf6b03636dc77a02d5bbfc
z8040232b24270fea7fbc171398bba30c6a54830d039be9599e47a023cdb32f0f3e79580ce4a4ae
z525afb14cf0eb5192725bbfe975c26fb40c6771ad48cc67ae27b588dba8ad2b56a857a10a49393
z39910ed055e0acbc74c504d7785554bc5d5901e115d24b790a0d253ce427d53366d43cef80c70b
z0da89fa678df838fbde306ee8362dda17c9271e9933cf651d5fe8726ddd37096967b9613f44a9f
zd35d7ef4173fa562afbfb49cd9bedaa31ac3de4cc60735e6d2b3d777d90148db36827df90eb059
z9cbde8d6e62346344986f05bfe26c5c4c7e8b8c7111a7bd89fd9ed8073cb010fb46259f7cf4da6
z801092c6aea02465e0d30d7555c63ebecdd503f381a9e6ea034bc738a755e286c658f53f8542ec
zba52c08fb4dc55cdb7a6b6c00dd2dcd61e74c1f84fd3e8f1433ded8f27a2622d42b0877ae02449
za09f63e9f29dbcfa444c62bff56532e8f28cac872dc795a064096cabffc0a79647615b96ddb171
z14ef90230d3fb4d8685125a791258876e56ad4f7be887acf958d0c362af3159cfb734a0e70ba28
z06db3d5957a30f6a3e2ae34a55205a8db6243f0e7356be9261798f2ca90af6a015105333b4deca
z10abeba2d9ebf453e5675a40394813be3050016e108cd26a5472b78e84742047041e54911da48e
z00a6cf0a6c933da497c64749bc257c05b647e69dfb0324928db03f3ee989f65fe8b2f68bff793a
z25d48451410f1b0ffdbdd4077763f547b07dec4b420c1000f2693c7e97f17a47c32d405ac8905c
z91d84b7cbb736c42da415422b16e869081a91ffb44b0b3fd28651b9c5b5a10e2f857a998d08919
zb8445e1bda0246dd453f4f074e96dabdd7066f585844426355d6b4d73d9aa92aacaff9a6c5e46c
z7d4f7ed9c72ebe0dea720dbfde11e2659bbe07cf8e15de331dbca25c27421041c9234fff1bafb7
z13e4354f0b7ba17bf9c032a84ddd0bea89a113ff750e7b92cf60d8a8d9b6d98e2b6c9c977f7a81
za35a6108abb5d0f1382ed4584704ae42dc91d9b9b746a3bf3435f6845a54200027181eb263c3aa
zbcdd19f05a969881e328aace170fd7f7e78efa8d5f6209decce88bae47482f8c46e317f17c0cf1
z209055679e5931fbbb62f5f5032210d34f72ce05c87919b3a4ee2b73558af797f4314d7572105e
z3bb6d0ced3b6072d8291bebb9525c1db0a48e48b1b63d02158fd4c493ef5e05afefebe3a571309
z105fa48f4c47fd36e4d02bcd4d3efc2aa215055248247ea93d5fa7e427481919673ef4b82e80b1
ze50d8c4ee3006656fc4a921b24c3328304166b2964050f03c4d12ad6b36ec93dd957c185bf610e
z0d0d4875de36302c6a177822516f41f457a0fd3e02f71ed7276b8d02fa263142b4b71af67c08a9
z4ddd54905851dac782482c73b7ce84a9476a7e3d903896de24df710739995cb6c37bcba434d005
z38568469391b3720159ba1a226f05e7a6c198a8d88de6e3d26b1b6b1e30f2ea521fa0db2fe470c
ze15c69ba8dd4fa1ecc46b1c84778db471bbb216fdb3954c284dd70dae68d8fba5e0665fb86e93e
z016835cf29d2b024ee60eb2d0642ef93d4efbd3b6b24d446062d982fa1c6cf7a82e59d7b3901a4
zd8c32241cda62a3648f90b43adb07e5de512695219f43474eef276449d11060362b07a6fbf3e2a
z36a668dd60f7ca2e0273a7615b1d14c6c235fee2a20b03f1a16422a80d0f457dca8e1a36e0b9ca
zeb7a175310631ad555462a69ea122da08482e69547f83a8f829b4c9fa23d96a5f869defed95334
z38674a717f74deacfc7d066904e4bc0b58833c0179005fe753885f93a8571e1df4b9caf514a878
z5e0e8df276769e35d3bd8e7ccc85c1ba709802da2137f80430d337b5bbceeb3cb02fde8dc7e3f7
z1a396fc40ea3526e2c6eee486e3aa40c24111912228a6ce6095735936348d084fb0e8e5951178f
z72e7ea25f24b51063e87222c48877e66be9f45adb2cf0a73c31335bc4f328c22ad90de4ef53996
z6a62f14c395c920c5e80e668887d10bf6287fecc5c36efa7eec0268163c160164477b24494ef12
z48a5cb2b929d38291a8a4e306abdff3d82c97a8a262913714afbba376263251e7c4b511f2bba19
z37f39f50e80e09662bce285c901278561769a42be934cf10c3e7fb1d6f0f687b454a366d6a07af
z6c1182a7b4996271de00d0f32bd126cc75f1bdbc2969ab46e31d1c037607b9428c5b9370bba70d
z851ff02502230810899545d3f59d71faaa664bf55814b54640c94f19c3cbff3da740a6c0dd03a0
zf9da685723287a53e5d9ae98e12edb640609977fc7823f9d4d9486bb5b65643ddd54b82eac4e08
z9035daaf88bdb246a58d8aa586d6da0836eff0c3fbdb74744824b3ea7b7afb5d1cfb11b550b19c
z99cd1ae598e1a83cea91cf1e5e0e9535d310c5e5fae246c2643ed29c2d9fa80e6be744e103956d
z955b724a0c0f009406349330e2eacebd472287258bbdf52451a9ce3ec8ff2179b1ae707c2063fa
z15a7e96210535deb6a9ef03952fefca0de935669666ba535221c59a101932d8e8667f4535ad3b2
zeac805b93acd6b64c543f0571a0b270cebbb92979fbc4a0156969c88464b696f442e2f7cb12bdb
z3071463323d881dafeb76a4bdbdcdfe606ec823d1ed38d866b32672072d8a4b8e0d1a631d31e44
z76bc6b90b40589da4beb6fa6936673be76d78c2756e7616c07b324c708b7636c070ae468b0f62b
z7d066602f0483ab48c15d6c6239f57824696b68492b6e9bb4136aff9bb1280633665695ed2f44a
z5794b6e9c7139a4227f3b5062fca3bf7117a846e6a2540dfb4864318bfdff5d00e840ba432638a
z7f6ca15263978ae87df35513ba3870f59a3d6d8f1e937e6aef6a2ed181dbd4c2e263a07167a07b
z84be00716e17ce39873e154b460c3c34ce7b600dde8733b7a22159f8c6e8e7b6cd10387329dacc
z7b66753d1ced7b978545a033d12bd62bad0a435a1de62e3a03949718d6a70cd12092bdbb0f5da9
zbb8157a849368b62bc60ad4a743dfa69e76272f7fd6d8a4c9e5bbf33850ace3c07758b83f0fc8f
z17e6e8c347d03a090cdb0413349757ce558e86c5643b51ddb30e135c2788c236f4137eeda15fe9
z5b017aaaea3fe78849ddb9ab7900ae44e61e020a120a65d4f4da5db53bf79b3aa88da12f453c17
z883b7400b219e7b1e62e7da70fc5e10e5e28813bb091c3329670b173e3a81fff3d2c4f5ec9c3d2
z3c08c7840824dbca96918a6b9d31f0b625e7280d7103281d21765b0f38c543eb484f32434ff979
z48097be6cafddcef175340fa3e6b2bfaafbeefbce16fe2220bdec9574788468323513ae2f3e5fa
z78f2437a6e37cf459f8082d0c77b958bbc1339b4a24debb7b5dcafaf7e06842d94d13659f295d4
z4dd8ce92a47ed51a097b3825c5847bb6950b5130a93253440dbccd755e5c5ee745660b71e17d11
z48ad5368720d3fb936e38e04fc1e41b6d8d58ed011649bd6fba7fad8b029c7b9da7566d4efbcb6
z9e530dd081d9b207a38ffbdb903de1b36234e105af91f863a71f69f312e895b1686a1dca91a504
za71f78c20da3f07c1feb24f208f279a7d61bca2a87ab79ed4dc0940fdfbfe5f52e67c87a094cc9
zaf66eed80111e1e42cd63896431f61cb7027e11fbc0ffca67dfe93364dc334e6075a533b10265b
z967b9db873560b28223f6281bb590cfe2d490086d9f44d7c87b87932a16d30fad76b4fd522831e
z5357b372f0f4d367416fae9935dea91a500384fecc930e4cc30689c8d6a51bdf45886e0d4c748b
z7f81c47a121df8a89e1848e2dc50c0e7f03ce07c4be09b7c325e2b11e07cf26e27e4a9c01d8b7c
z9c6e32ff28534d57de00fc395ab09efc1deb62e06ca29802aea0d6b3b6f2de7734161709859cb2
z5fa7b729030ccf9ba60b035e5273487d347c3624e37d0060f563984525f598e1dda00a52b021aa
z149c93777003b0f434bdfc2b330b90cf69ce43551ee63bbcbe382addf634d59913c4f651e46db3
z70ac8f801fb346d77467174e74385c8c9968111be231d804280636128423f2846bd505b0b302e6
z496cc11c43a83c29a22d7520158b10979d121bba54780b3e8df7e706bc00c814292c65291e0488
za7e50399884fea7d27c730c71a56f8934bc7ee9b855a099c151a40c602e3b4422d300d556ef6ef
z81e4c76c818d6bfcda65f832cfa3e03a0c508b4c576c95b12c6e604bbce13916bfcebb1bf89ac7
z857b493007a2ef06a211373710138e6142d6bbc09396e61290c0bb874a37a5de74556bb32ef571
z585d9c74ea83aea17fea0c93a1cd04c0f81b5acf01971b77cd20d02d2a1ee7df7d994f6033b693
ze89adbae7e64ec43cf739e8641bd2255fd85cf890db92b9502c9927cd28faa1e297dfd1fe5a380
zf0bde2e55008dd24c81ffc5d697877e4e9cde31e77f66951f8e94e28902a45a21f48c597c170cd
z0691c1091298114a1b5fb86348a3913d5d7a4b4380481bd8aab2d60afb121f337dbc62783ea429
zb9b473f7f16df64979e1c482fcb137ac215572d1a0ca14ecf86fc9b6fa34824de7fbd5bc638566
z091c7526c5deaefbaa9a9caf74d2fbc43bb8f723e567aa57b0824cf9380cb138c6623f4d40e2ff
z0db9f5ee70306e0ed118cfabefbbf8251ffb98e9f95763d59ffa2a9db9b4652a9fc8629d8985c9
z6a43d65c4bbddc0633aa5f61b56c98666c41a0f41c8a2f27b8696442c4d215bdf09df276a42c27
z0240b763697417d131153e3db2c4759d5c91b2aa1fbca1d00abaa02e36e6384089f2750d92f9b4
z082398a3a5f967e707cf6c1084c0f4b3c2630e1431433ff54b824190c34fd077d80c94dd2da03b
z8070b4e0c954799da5b12860cd8c6fb89f19b776b16c542d0eb7e3347ae06071f7972af30dec4d
z11d525118ac8ff7d85cd3cfaeff63bd7774fcaaed820d0fa84ce4db1278ce8f6ccc12cec51fa09
zd1664465b5354229565f08b6d91279dfeea53a56d7fb34b04e9103cfa5d72801dfea9267f3bfcc
ze70ed6cce05eaf6a51422f4247c668de5892d3bbd7d0235bb21fb9f8412336af0b58f0893acb30
zaa18df41e34a655344fbcba3235bbfe32c2762c8a6e2169f155a0b09af9f7e6d1abf01f427c459
z9afdbdebcfd111e90de5fb953d61065da18d18f38921f01a366ee4473ae9b3acfbdc2e05294b7e
z2c48eae90bd7108e43907432e3f3f402b22c7476f0e72b4ade5168f0d525662332fa32b1ef23c7
z2214e3e587fecc36b319e96de998f20136158bc6fb14b59c78a2c1077830950653f8f1639c9dd9
z0dce2437fe859f8bdae5be53ac504fc6a303ad23674aa4ee9c45a6ac60b27886158e5afec188c8
ze8863842f0b68347f6bf3dc86ce4e4e7d6b98be0141758bdc0c74fcd4cf3facaedb479cba39b39
zffa0593aa62106d337f6eb7e861959363f5b21ebeed82499a86cdec9c9e9ea509cc67406c0f795
zab4738d93e582704bb541dff1eba3dbfbe72080e377772e495727597a77905083bb82c7f08e063
zdb0955e326d343ce48217a8f3829198e5b6ea5e20e694d1af1285c94f1c82714a2d70bdc2edb97
zd295f330b18bde2053cfc366991a9b91ae4ad993d4e6c0596d279f8c81dd9ca5b1c4ca43eef458
z14080c120f1f521d1247c5978cdd2fb314d64d56a5be49139811e4e9b30cc56e3baefcf96ef06a
zc3a40427b973a1e880e2ecd028d79e82028c3895af395e7658596c17ba7a0b91efbdf96b167deb
zf3fa34d1c3fcb0f8618ec98fb461bab8028886348024a4b4c8f83c3878789bec22bf965df64b39
zc9e3c40b0212876fb85164206b126ce4b79bcf3604827fe783fc2a3a0054f422098861a0ef6cae
z279fec803d8dbbcab0f3ecb1a55fab55c19c191e8af533987a728f1e699fae5b769ba522200f83
za17eeb7c2c40be03a2d699cf34a81001ff243327d3bfd0792b3c983936ba740d8c6658e55f5aba
zce942555e70cdffef4400a32fcb72f464d417683e5dab03eab61384a047d3b5d0b98905b676b02
z25c967ee1430977e5eedacdb67bec8bca576e028b146acb11f8aff4ba9b82b49b559dab5a17348
z77109fff3df58e8b159e8d4019b2a72f428b22c2af362f52618ee6fa018eb42ac526646ba3ad35
zf4fe42ffec1dadd1b4cf236eefd3fc3792c8208f3e866883aae82b19e11efc124fb0cdce6e95d9
z8aba2dd1ef9f9f8273f72d38b1ce0c7eb0eb1359450e850680dd3bdb09dab757faf857b313331a
ze7ca4d06d2fa47bead34e3ffa32591554d82f280f7dad1480f2554b1a9d5ee6eced4d1ef1ec229
ze80359ad8bc8048f7f3d42cac6a01b1404e0673f0ec52dd6fff76b403082d2c76e387f16327f33
z0358b297da3f0bffda83878d6fe6be80024e06ea69f6d74dab910f7c941267023b53ae229bb2f5
z04233f05fe2b261b2407a2db2d73b6ca0e0b05318b02142bea8cfe23ea535a7ed42d89e65b2238
z03464a047d4029863f9f597292f6e75342170e64adb41c1ca9b6e4bd2e8c7aec0afa1cf7257e47
z1491088667459eb596ea5d4accefb65d05a6426bd19ba02a13c5ac415607c48a2178b6ca410fbb
z8d72e3ed2eaa0f81e24951cae7c59d6e8dc63938b377d0573776d8f23255bb7e0193c5ab876eba
z6dea1e5af50555988c9e05baada7dcb095de31ff732c7ecd3c939d32ddff743a9a068246dda86c
zd197c10bf2cb35e3050557ecba6841b260a5a0b355312bb597d0eea4c743bca1546028b926b62f
z846b83e10f64427fa2e4bd8ec5fdffb94a5ee672e8099d829c7fa97f8cb7bd64fd1cab88fdb88d
zfc114e138d65c1ad6fa3f1faeecf4ffe34f88496bccf4b4f0ec7ec275b898eeaa70bdb08549310
z3d696797c7ddd3054e7b0ace41fa48be6c6bb8ae209e24253d9e958020f8ddeba36f692940129d
zd48ecae5d2b8a41066c652e29118ecc8b545eabe99cd4ee99b1684ae464447b3a5fede6a680fef
z82db43adfde9ddd61e8c11484f69eb1954b983d5b186e3e1fbc9d1e68a8af53c31dd9c4127fe72
zaddee5c8d17584f4f10866bc2ac625da3f7c6c6b009022638490270eeb8062a83bfd5991a4060e
z3612e29b9a8b86402c5d8d324f6e4e70bc00a3392b631261cb5363409023247767e31aa97ab82b
z5edea7aaf3f27aeab408e7dc6cc6fc7aba886948d83ca6b9b65433dd024d98ad283ae8eee36cb5
zfd97f018f8cefb26e291252a2a5f16afd7d6012586d4fe82512058d2770c340f2f82b95c3da99c
za6f4bc74a2945ccea6d818fdefada1a6273b0bf82e38104f47bf2bc83d0173aa285b9afc04534e
z4f7e553eab2dce0d13ec4ea742164f81e516f8d9b01f2b1916b216253c5ce795039291325b4e4d
zbb4723eaca01819d0dd7111adb8fcacaf41ec90d3ca0bb35e2ddc2eece01132a12e285c70977d7
z19c032259dfeb51de453eb2db827b47735e99e1cea2a39ef36b3e5484aba9e724ac421f9740a8d
z199977737db0b4592dfef0edf683afe3a4ef6cce38a9312388b74e49176c251a5c12dd98c82619
z2960588a9a0dbc15c4bf99eed4fac6bf0e90c2dc5a6360e057debdda659c920b2a814d53bb62a5
z9612b3d77c0676a07be7b296df206140fcad86bd8e645e54315589dde589d7cf5adc3e3aa5f958
z54898d79294866ccf0599f64ec056368fdefe545c757080724aa8a4ec09c59c8b3364d2ca86d13
z73f8d4fd502ff4dba08f9045cc0f08e9bfed75d8032478756fa334b582ce68d291b931a5637e8f
z35cde95fe9fb61bea7d26ca95ee9aaf2ffe3fa224c44df496e6c9e249eb01c0a3c221bcb802dff
z615e2f626c8048a3430fff42b2b1fbeacab3a73602fa67bdd53dba7c1bc1e8c6fa9dbe27fb9339
z2d094d280f1b4848eb5755aedba107a71e0c357ec7dbf9e5187a50b395c7a3d1c54ebba53da28f
z3a13f3c17a1672495c2e3fcf629623b5442c15476bc869fede455f28f72e2dcbcd84fa5efe6f68
zb232a6a2d36c6764c70a73f519541b5d6eeb2e4f5c348bcca363348230338a536f46cde441d4a6
z60764b478468cf246bdbf53d05f0dda0d70f7dfed73c7b93983bd65d4bf1a093c4fc34fb4424ab
z51c01620de8dc8bc68cd99e9348daf113ce48b11febe0a9eb36fb39f0adbef20dc2e76a8d535be
zab1b331ee48fb3407c3a454b9f805bbf8e3bead518c69a947b4fc016589899d585e261a07e74e4
z0e6192d5dc0d6e66502662ddcebd34fe832cc2ffb7cbe17dd5e01be7d7ff4beeae72c915e33978
ze111c5ef9d6fb030f975e14f50b483da0b8d07083e8fc5695bf34e88691b3c7df502e02ef33e65
z9e017a7101a2e66a6046ad120f5ba5d5f8b533820ba4fd55082618a49aa50748b6c5fb40e94cae
zc2fe9f41b39d0af82b3ee484f3659c9f0396682be225e55d6b9cce88ad249dedb86f7e927e2365
zc029638ed5ff542c7ebd7e9882f6a7fa98ec8dcd5eed1c38831215c8cbf00231383eeb0501928c
z6d4182fa4ddef250c13acaaccadbf573d4b6ec0c71f4363f406fc8bb44d75c24b3edab04811f48
zae3fe7c294dd24e26feb4569bae96595e8b694a0a45fc26dc59dc4dc556c83c60e12725b4c9d82
zdfab97f956aaa2691de59b8a1e48e0fc163c3580f35c13eca1499fb4f0096e673806d5d07cfc77
ze648849dbf368111f61bbaae1a9ec83969519f6b9d9d9aa6244f9604fa86985dc5f7641e12fc63
zf2322f5b674b732659b9804b16364bd17a9854cd9ee6a47be12246944be93b489f1199765d8822
zc65a9368b01ffbb3cc964f961266fbd9d7f282ba7086d13c7b929bf5e31c2e942a8aaf6c92db1e
z43c7a775f5485491f97bf65a8c681c0b889b58a90099d101faf10a45bc27e0bd91f8aeb9931f53
zc838422e827f9f43383ce877a16e89485dbd3752b4ff04e2654bb7c9b65b419f9f448917e6433b
zf2a06b30cd6994f67fd2137d949f4f3dffd9266b0d0106bf721424d748f31618ab0248ecdaeba4
zf66c3c4ab3a2e9febdba6f13f9251e718f24e81047a6a773ec5f8cab0756d9590165200e2d3de2
z81f254263d544323494d82ec12f90438ac41de899f66d0cbee3ed5aef6f4a76a40b3b12d30bd26
z1de28cf5f4d84d4450b12f4d71c097aa1646ea3670c9db62acbcdc128c9f67d061416b82e24980
zf0be0b1988eeea2f682dcf33b9e75ee01422c0b5438fbac4bc765778326dd8524cd67d4071c98a
z4e92aa471db2c2b1b61d2b3733aa97fc6628f8fed46dfc63da7ee8bcf01ce6c145d344a9e28abd
zb545d0888d5637b0602ce8a2391274847edf69156e3c1d9eb1a4889398099d3613cd447e4163b5
za4fb92687389291b9303e9855c9a859ebd9444b1d1521d84474d1c6df4b866538be4856856962a
z273c0086be200eda5473a180a2d97a5508cf17d551664d04c1eab7981dc0e8179218f04c077c55
z2dd64a56d1003684f688ab0d40e4bdff97a8bdcbe978de146cb258923564bdb692d9d7c180082a
ze22947c563dbd4187189407da55f5703a99b699dcfb0bbba8b0ae50d20015858f28da9feac9f85
z925364598969f1772704c5790332b11bdacb648dcebcc3214364bf30085922e7d77e9aafdfc44d
ze50f744e7eb41993344e94cd2834949cc8f505d4245254a597572193876013ae0fc80b354bdd40
z1ccff1ef198ee8e175da13c4d62d0f2eca56181b242a96f084533cce713383b5cf3a83554ba383
z862701a074e12500541a8ff170cab10b7c2bb7903b9a17d70a8b05227de54479e0d153b3632081
z6b08a02defaaeb2e2294dbe81bcd66b4bdca3d12a01cc6b52815e6afb47d8ce617488e01466b67
z1e01c2c349b020aa345bdcfd31acea31c304ca3e763f6a0cd6007ba7a3cfa3b9ac3039e50bf7f7
z560eca8c76ab03eb6fd9738ea0a6e24620a13304373949745df504157593ddc51f4bc0ad31e01d
z09d908b6440bffec346c146fca04ec8c91f7dae4ed5f53c2ada8d5091293309ee162e6330629cc
z1ff33ce64b2278c2ed67cee289f0d52d1389f957dd2a7626ce8599bcc3975ddf7064c7e5a55923
zfa6981770604dbc19ded318b1b6cf9519c20237b71441aec2d1db3eaa9274fd55868e97d008642
z2e9bd6de9997aae9146e989e4031d1acf0afd42c8d686ee35e045c19324a0225ffe5f3f14bb6a4
zdb0d4132ae1d5c5e328372c454380b4f36644fecb09d779a353710f45d8886b07e9f45a61fdcd0
ze37c0bb49bac8ebd1ff7560f832e25cd25d196b744ff0a7efdc6d8896dbbac3bf4118fbda3975f
z67e35868f3008f63e3089fa4751ac64ce19143190fa17250379e46d440eee5bff6b3cb7fe6c5cc
z08aa82fc680a4f886ae3e22414a7c84ad2ff4547e32d2b22a5873ec7c27bd19c5e7a8bfa073a63
zb74b33cdc9aa301caf62a8d57901e3cb55b30ec393619844f03d1da516f70be8d3d09e6f68a4f1
zaba0aa65de90897194bd534f1b98db0b50172ef55f38cadb79464c277fa9c946ef6709ebc8d003
z2608a50c03e8e6376835ca135ea38d79dc846405ac85b9d71ef1a83c50282cb01b3b21244d99da
zfee37112a172f2e2b90e730fdbf34d695424676cb465ee53139eda59f6c0ff07e4cc3797559ce6
z09e4b747a07e8b75b3f27fecf321843d12b5422002e36eaafedb599ac6548731fd3cb43cad3cae
z424c738ee110777f00d72f91f5851ae785d393bda3524ece41fcde8794d02b4544921213705912
z52f540c1c38cecaeaa0620850fa0edb1f41af41f947e3d937196070f8e9626ff0e424ccb3f3116
zc3bda2e3dd09b4dba2a1af88959ef19e8e3481d25dd369b823b1d18e7c11f7cd0f82c1ae3883ad
z25646e7d70d686d5e26327e82a2a01a4657857d0e12ecb91d1a940b3d0b02cb1a891d1e74681cc
zcfca68367355d4e01a6260632e5665cef58d33e6a0b783a38879e17cb7e64223794acafeaceefa
zfaaf07cb547cfeacf64f9e6cbfad7900f45067a30696856768485d7fff14d5f69eba47d54dd2d3
z15539c96c2bd27b73291f05a163b52df2464b163cf1d2707d1cd35afb4a8baa710eba11ba8a6d6
z48ea29a72aca7defe7ad0e4de28fc20859501b7d35cb81a0aa3689759d302a0c957aa0ce20702f
zab717598a12f437231b322df427ad85daf3db3994c0d0628f80ecaf86b5bce1b02f7dcea75d369
zda7a2c2909bf9388ccb97862c65ad3e448a978f4761b5f9798e6290df551cec7560022748e7132
z53112f3a025e10f5b4989f2123c8f6a78869164652a8c42d7a880ab57c6a290014d069b4e70296
z3b7699d4726eb8518b6ae9dfb12f69b2b1aa3c172cb144ba021a0bd169e9278d80f1d7543b1b60
ze448197eec7d7d0c4df1a3e0540999bc1044cb6b4c30a49d158181929a4b8eb91f8d3fa605d4b1
za027febebe51f752ee393aaf060fa8b2261da1dc349dd4b735960a7ed25934822f43b8cf234429
z04d7f0727c64d26c63506785534802df669e468cdc9c35d986e9c68229dcc0a953e4543b699c56
zf5396717907ac871f57c00f2580a3bbd8eda0eeaeff77b38d12dab9cf522d738b37751cdf39e55
z3290ca01be292bc4a02b48bfa214b09c1b16ca288a3db1357042c18c33fcc8472f14bd491e77d9
zf137da6ed218ca3dbce9c15af1cc318bcf36b7ed4da3d07d6036b53ea631675e64b7eac36d2fb4
z3f1d4551281979969ca8667cead7da9556294895850472ba5199a969f9b0f854c356e15ead7a23
z12ad14398b0af153601aa068837cc8e16be2ddb33784a16fcc3d3969718c036accbf84fbd17a85
zaf70486f38087698dedf8ec5e6eb47239e3d2e38cf57c9080ef761d31e1e68cb128ec96117aaa6
zcc440817d1ef9cfb8265d567c3f70149e3a48cfe15402a035ef7c5c41628c3cd97deabf61beb74
z28e6cd6643194226e7a4e75eba8a29b25a0c5d2aaa1ac7cd56d4d06e5f42fb3fd73b09d6c32f50
z8f685349765a067de33c690f899f053f45db9eccd690d1e2520ab13ce6fb532f7232cc1e5e1aec
z1b1740e3b9126a351bda95502c7e3946240b72c06a06fcd7182ddfcb43157ffa24f1e880b992ae
zaa1238c708a3610a6583bfa4a20c96218fa3df547306ba359e8f29b37fb46a7bdb95ec3eaf455e
z08f11bb5baf86b0303863d5d28360afa033613ee7fc86bf698432e26d6956b7ecf1845c7598d43
z7491d349ded092a693fdad541f7be50e14bbdcd7ac69dbec425762cf4232f5bde544a184a87d45
z5835c9b10aa411cad9ba34a293036b224ba8f12fd00aa343b5a8d75cb92450986caf494b88fd48
zcd9afd15acd776a928b1a21ac2a6a515f982b60dcc43470119e88bfe3d56cea62ba406e2caac4e
z4e13dfb0608ccbb9a02d120ddc7e5bb41ca80ae20a543ec5a0c9aaed5a456d577ad43beaeed94b
zb28d15053c02828082b66b4e1b777600272ea56fb1aa6f0dd7935f156240a454056ed458c819a1
z3f50b68504966990384e326819dc674a0e3b718ffcce36dedc59fbbdaee5adc3b54217e06d6ff7
z3c84d291f554e7fdadf46177d711e17583ebb42ac10f213d3d7559c1a6365d66141b22904ca13f
z83f2c6b1b37dca2c7105aa292718a6d47496fd69aec7f88e4f248b90b4fbe58526d2f2baa7fcfc
zde6dfd7b6f1346203eeead528eda4e88c67bb144b617f48a5cce27a96deca262e46e746abda4ab
z775aaba0135fb3e90876269c224b7fc943a75b64cc4ac066fbcf847b8088067d9e54d6ed7a1a9d
z2b4e4fb8885447c005b814cb770cba9f405d350f32cd2dd1a9b91e15b122038b5f555eea618f0c
z0e36edebb04981b7577332d93679c6e74fdc6599c1b2ead90605464cbbc55fca118cece30dae03
zf84d35c0a77ba5092c0bf56c878d17ddaf5aa2e509ef6ea2076fe02673f821d4198f5b1f656d73
z41fe57bfc8773f112e1cb9e4a63c731ebad1b7bddcbcbfd31325b029b9ef4d8155c85e2f435af6
z035180bb371a9be61b7f8ba44addfcf6c31b866eaea014137a6d1e2a04903267204e0629485b39
z21db5b639f33deff101d23782880629fff46b1d311b6c773588da30141a4cd63d37a13f34ef1d9
z8db9681ab97891452b192aa9af0340410fe847498d4474d1f4e2b62dc948768499c8dcd64c6867
zad12f1376efec2d631bcf37b25d0ba5bed3ac47cf3710bbb717537f2cd239541a0caa601ee6ca8
z972d1d4feba50a390ffd1307ada66fc77477dc486833059f60554967c93cdfc0b7f12611f91ab3
z8b9c9f7b938fde9fd8d9ccf09eed0eaa2bffe62a1d3b5b0cd5689512023e2a7a749b0f540423dc
zbd3feb0ccc8b9ce274be37d80d6be725ff9ecd9e83fae0b5cd967e909467f4260fae6cb4071a39
ze3f7dce98651b06df43224886b6814350f1b13b53b18d02d5c8e8eb451c5f4ab7125b647843bde
z9043451786feff517134b614f7f514c1022896fd6be68a594eb6959efd96e71cac7ce6d65a2135
z2b926e158c3666b510b8baf7a1c0e2ecf829441f707d9aa057b41573d8534cbc20a67ea4fcbdc7
zfbf06a7087240a9ef804fbd7c91847df0e013daca21bd761c48be13a815a22b9da5e671fdada4d
z0d4bf6c81caa8d6b49af4eacc407908f5b707ff8289d11c887a2bd006e12d0f9f17168bbe20eed
zf959facdfe3403d5910b311b116f4741e6f0ef78ad3cb1b4fcbe785f9911640d31a8298c20659d
z1da4dc5290fc36fcb4531bffccfabba3b34ac88ee679bb7b06e666da4b7040395df259e0f70f4d
z8a56903c916ed434501a0092d87301f49db3f5d602cbe3257bc9a4faeff73c78038d93764aa64e
zdbeb6e9fc4e58faec47b9a8516cd2d678737118c17b3a1d5860f7899fd94680589851f1b0e6b35
ze2cc8dfd435c5cebe680fb4dec6c355754349cf4fd52eda4fdfa7aeab4ac8ed836e809bd9c6405
z2a7ec4f7dc03150e4e4a2e485aa45be405fb9dd65a79f7a0f82b00cc5f394bac37c1f8a908858d
zef19a031ec867400fa7ddad8724679c3aab79226186e20250c04031949b2bf215a5d1222cb186d
z991ad6fa5b94c02db7c9aad04544154c2616a34f58fad0945d8ce171a08efa1950465e67119a29
z4cb60043568a96d083175360ed35595811b09ed9d5542542f565eda87090d4d3a3bcc7a2fb40e2
z57a762a06c8164158f4f3f0f7a8ba3d3ba888790f12b34d0a33f7d507240d6ae7ad6a30b513285
zd1c32d768e74a034ea191b36fe5d1d3fe511b520547eb9af303097b1469769544e878d3df5cc0c
z239df46f1463db0c09fdeac12349c360bb3149fdaacface8179ce3ce583a10703854584374bc81
z98e67f3f9a5470e99aba5199ff9e5f945a97f008820cccf956853bfce36b4b7db69e0771fff6ee
z86f1675383875d334368c04a4d55ff6eb96e0af185e253f6a5ee10c1aa63f5664eac3875c74481
zfd15e60105e3ce7db633800b01cd7313bd947f2782ffc2a83cfd7c0a4372b5f9d38c93dec3e96f
z1e3987afa16b7537780c5c8db65649e0cb9861ba238f9982a32d761e1a03a49bd1ed2d873b3776
z3cbf839c47fd31a19a380a0bd20b69e6b0bb670885c3924d9a0b87d36b421ac5e220ca33fb9f0c
z805efb872a2d814fb4dfdb255796280cd47fc31743ee26d3438a80f579ae48a4d55f30d5726248
zb9839988b10a601e5cf0f579d32c5760106ac0e28858bb09bcbf12cac4fe49aec9c0be4a69fa6e
za1d0d1f11cfeb479f32e5faa342177dacc38e6895dbb9d969bf5dff40b27662c8befe30b9ca3c3
z0c116226ed9f712e0b63b8a1885547aa9e383125dffa5c3f2443541a72e8a7fe6420e1d9d82c07
zbd0a318a9365d733c818eba161a74f22e48b341cce17c7681b6d057defeb512a461b5cc5860eae
z7dc1765de4882b7b1b8c346114f7891275ff08fd0f042ba3f7a4422f0ee7c0de1f43439bc63aa6
z0347640a628c15f264d7f8aa2fad3fd85321cac27481e9c968816124b7584cfe2de0d9084ff01b
z07c521f9b8eb3755ccf0e00747f2a6b4dabda62d159eb9597a9b0e35cbbc0fe6a673d45c45ced9
z3d3383a82a25c997935d2c5bff5dc2b394a494eeee3a4d0cf452d1b9ae4fc6e0eb3cf025942dce
zd5416c292c72396e69891afd75a005e6e25d600550393e2f22e7a69b0170ec54b2b987a5da96b6
z40434d758bc8b6cccca731efe643361ce06d4ee8d565c6a28b0f165bad0257f8459127434ef0ac
z222066926fa06d117e5bf2fdd85b67904b853e02ecb8c371bcf7299c2a6bdbc23701f18d1577c7
za748b5bf39fe25d2d4bed3615eebdcc6c306cc88b703a6a6bcf19bb44ddaa7de7ac8f73834b4cb
z6cac99e50d89cbeb4ce8380c31513e6b5bf3e7f0eb7eb54d03fde637b69c542c987379f540f878
z3f11c8ad9c50051684733c595ef954bb5f138e366954a2b64e2f9e4a82ae807ade8c1807d54a1a
za9a014f7ed13aa2afba0e71d0ed7d9c421386014f6f6a23f682a2e874d0d6c7c82315bb32e08c0
zcb6008fd18987bf9e9c2622ab811d5f0743d0a2476c09fcf6790ab4ce5a0b7583acf8ad04f300c
zae14296809f1b7b2f4bf1d6864f344afafc68041d6f7143e16efa3703cba090d6688de3148924e
z1a6a9af985b4d57b9ab015f4348c4c3ef60e857e2a7fb31d1374badb8197bccdf6a51b21027a6f
z11a9203b764dac7ee6f195defce8e9dd9261908c853bedc9f01e7de511300e33aa2fd80d4b7995
zc0d7f9159242a92f41baccfa13bb642f9ae43dc0cad63b2d26abb8446aaff6675bd86b7ec56f6b
zaacf33ce3a7845d43894a4213c53b0162c93e6e8eb06554577b276adf68781663eb8d1ff1a8b6c
zb7a1fa5261dfeee7ef9f9a5421d5f3b5b83f077e57fc5102de6604ca44a0c7b05ca4663b124c55
z64c6ef8152c5a9243437ccde9435003c9ccae71ca7ad9e3c520a8ce20ed7951e31b10921f5e36c
zef2b721535a34cec4fed15613c0cdc14b01255501e4a977daf6f2623d71d2ba4de0aa1a9dd08aa
zdd442ea0bc00a7d4bf513938cd7d4325be93317a060db6cdc0aed1e81da457cce91851402f698f
z9abf35a84b5eecda8024a0980ba76e284e7e6088a2c89291c02ca96c51e9450a2c8447ee0ebafc
z8e0dfb8addf7123152b9ffe5e83ce7ce1e44d870e7f154e9e468a4c2747e944c14c0888eed831b
z7e973f1df61e3d025d7426ecfebe786a2f92edbbf0f8513c78ec7a742a55d2afbd2a935587e16f
za5cf28091ad2c5cf974fc8f16458415e1395a4f4c536fde8b948018113bfadd5bb7aef95fa9b7e
zf2fe8a7cc5e02856d9005c9cd74e1be758ea07fbaa3143d04260a6746810e2ec8bce766585ebdd
z0fff82e60d5b842a56f5d807bd9d0ffd2009758a951bc4c545d7ea5ed54f8d14e5e62420bf427c
zc8eb9417e5374a3ba545f8f733ed8bcb115d83f435336a058efec13ccda0cbf4a09f914fcaf364
z22254b6dd747c09a0a95028fb4ba773d8740c73875619697faec8e2c8f48c9bf0fe767990fc0c3
z637dc5b26bccafa41d8457f295c792578e131f25442bbb7944dc1266ba9ab9fcc7b30bdd7f0783
zc465cde1e22b3c9b56a2ed5d881e3749ec8aade80a7cc654af9efae9013240978235ca7006df50
z0671e435293659fec78308719f8984f77b998816115e87977983c10ab38192bb43a71cf47133ec
z7046e82aa11ce8c8fde7851b10b9541d7b0636da4b0be072adfff5239b1f61d1e4c5cf722961f9
z0043aa7daa2016257aa5270b21870df245bdf5daa2a2a78213de1762e7dee2dd63d33db1bdf3ab
za91ddde1316b6224c209b05d5a2dfdfbcc71a8f32c217cda23c9b4775742f37fe1ecda8c6341da
zcbd05b1bb0508cec1e52b06cb7c4ebcc1ded72286e5ffdab4311fa5254695f3d45e7711c3c4b28
zb346dce4c7087770bad4ec0588d8806534baaa23a6b22cd2d630e5f1f57d20f6200c652c4153cc
zdb1ca77fcd3d7d5387b8e9f516015e611550cf4106433fa7e162b343398111fe7405c8663ca5f1
z41c3b233a7b04a96aa01b6083b737667c5fbba3935fcc9d1eb8212309344d7dafce0211ba27f59
ze347df355c0ff0d6ef01b8fb9eb0fa96e39e76a153f8b918d72f8fa85daaceaeba111e8a4226fc
z8367cc3484c835b4c81eb1810636b59485e29035a2d0e7da9323e068d50d1c579bd1ce783fe79b
zc0d05158b5149d85a4edd97e4925398e38dd749f4d0b50c5de5834dbb2359fd6a12779ce2edb29
zf520df23faa4447a4e462ae00e013b4926125c08f11737d21a926898d73be1dc561b814558343f
z81fad31dbaa5cfc76d102a1dfc4ae6f0857c6bde8f30865b1d91ab2d2fb3363dbc5f1b327a0bda
z81d8e9cb97d1a9a351ac8711aa2ed072bf4fe7bf9a9d3c7e8e1ae1a2c0e7a3fa4874fa5f6ee5f7
z7db92504c60ebde68d633baec71a25849956cb5faac74010bf48550add0c56403d16c33a2855d7
z83f71fc05ed34281957269d3ec81a8a5994babad7348f9df7544289f42cd03a27be6eb2773dcdd
z3b873f247c2cc18d8ac6d5405d7a45dd0c8484e432eac615cd5df078c05b3bfc50330d93b1fab6
z8cd18493d22b2f84b1b5c55b34a65f219aa848bc699a8f4c589ee6ed65a1aa9955633b2878ff47
z9ef7f64c0d15ea89eb388c1e2c8bdb6b2803b738e95229261899cbb26b069cf7853b1df1315e2c
za4d3d22a85aeaf0089d7aaf40faf8eca8f3a69a2874d62d8d5bbe8408b0af7d70c4c096dca5e74
z820e812553097384f39eb2a28c218625d3768c2ab152eccca818fc8431d6731447cbb979d231f0
zf52bceed82c23b03304d50d02cd4af039d5256f693e4a3c7a137560768bc9f88763331ccff26c1
zbe38f0c9501379e2dfdc40ae06cc544f6c27246a97d97df5e04f5efe21a4a97fe56e14c043971c
z52c74597e92515524236bf41ba9efc29ce6f4ac6c49adb22115b2923edbc7e183395b0048f5807
z0e69a54136b7d7f132bb919326c4b6aa3e0ca8bfe18e030bfd1ddcacf21d46697c0fc51b4f8f87
zbdf7a890cc60fed1dbdcd8d3c2bd23081322e270f57074d97ffb6e09811e083d906d1a0540ff14
z39ee8e7748f9248ecb9f48322552d74c4047abdfa22d263029bfb7d778b99af4ca96f996f3622c
z9a4d7827403ac25bfa8ccadbfb5f24a830b6a5708f51633478c1a942b0e4ee04c10105fd4cf251
z836c616a56c5fc38e374789b4bb38e36d4200ea797336784282fd4600b48f281e48bca2c6fbd81
z6e3077927668d30ca69f52f98a7616cbe5c386e13ea12c36b5457fa0b6b69877293f11b24a2c97
zd3b54715acdad43f72afbdb6aaf6b87e9dddfe87b4788a5d29513131a225faf2e3f057865d3099
z457d1cfa351f669f6008f6d474b1acf7f4bda08117a04fc4b9c515a5d96e801eb54ebcab6a3ac7
zdb206ffd60d69908c771b1224884581e773d0f322cd78a265852f53c7b483b6c8abd188cb616a9
z16815677c5278e4b6727b74c4314aedfa4308d596cc86033693d6c5aacbe2110c0bd0844641f65
ze963cabf2dc8b9cede2d5d5aac520a0ab348eeb37b8aa71ba247d8d3410296a966ac3e88fd1c55
z59c46577b643ecce1b37c9e28b0089c76081280bb58f8abaad813b898dbd9c0d405932a2dca273
z2744277b74e1706d8ccbf325a3fd27942ab5a21beb64b57cb0c3fdb0e99b687919b34ec1f0f31f
zb14d008e651b510f607604203088c0defd5e23e8a1b12c8cbfb06d195914b9c413654aa5650082
z651f24b6dffe91f4ff65ddb8add9259978fc5a589ea824f8206a4a0bfcc2052fca3b45306ebd03
zff8d6794445309f61604d96da49781aa4eebcc8107f082c5b6b04fd18155c74faf01dc5f729c6f
za71a7d5f7ff0268f0881d790239dc73e9e7a431cebcad5600c8677f8adecfc028e3a2a59609182
ze911d9bffda67f2e686c233ed0fc59552be7995cbd0dbcbc8a42c018a972b031cd9bdd7594e812
z0ff32d54ff8f58c30d26054044779443a0de63fb495cb96a4fec201e3ee5080e368cbb7080eb4c
z6f814095b8817df334c77c6061243c2bcd941d8eaf2422eb247662df5b822794b3c9b1371ceabc
zf63cfcf9be16511ce2dc38abbb97216bbdf2bed3f7b839d8d8abd7bde6802ee7594966dbe05c8f
z653bce57658996b7dccf8f3610c12dcad87746bb887ee5906ec5fddcb603c917308e394a3566ed
z94b17579b9380210542ab3b31c157ad2f7174d804be170a64bf876847d059698b47c84a41d26c1
z6ced1a09e6060f12f4a75018cabaf753e2ec9a33e8edc39e7214f487b01f8899c638792e47f5be
z918bb040220321c1513bafe6643bff6b8d3229d4dc9144b15fab9b5ec81bc93a91395ddf32ca28
z1014bf703f3cecbcd7827c80d74ca47fb57044e10b9f067186fa1abe720dad16afdf72d1a15a2b
zb72cc77ef81ca3b2be7e8bfc3b260063d2529267e3be21177ac2bca650232b36162a8014f4cd34
z22bc08cfafff426aaafa0230dc587e5bb1af18809bece832524c81767d8210002d1368a327289f
z14b34d4abc6b238767e38faa3ad42de1d478b893b4f4bddf793454db4aaa9098eebadfd4cfb56f
z1016f4dbda7b3bc613d11d5e0f72cdf626e55dfd1dba5579f8d3e3909dcbc8b46d287c33c91a42
z0533959a8cfa194606479940db49da448e2d5353ac0fc517984acfc1dac82e2e178e18a7b45b6c
z0fa0d0a1adbe76e5e615b10a56356238039b9869f1170239c26de53fd276065a27bc86be558540
zc4b09ac936e7f430eb2e26b8608840535a9ef2594bd21006a47132740bdc24653defa173e415da
z45c7ca9b6e4bf81ad62394ff868cb58b6fa006752ba14b5a3dfb938a5bce8a3cf8c82bb73d6559
zc52432d6fc9994bb22f51c6db9972c937f93a6b2103a280a8c604b99f2643705213d3de0bf8c91
z7156f4ca2159715d2ea8542376edbfafd02a7cd1d9e665422328ce53f05c15a92b1ea151fb8dda
zd1039cac6060ae2f398168f757a5608d896cef38810d91c7c948c5fbd1a833f8f4dec8467a2fee
zdd75c581e160306b46221fa5bf479904648bfc3c164e7f8c2116f103fc1f5750f950294db2ba7a
z1b49802d2bfceb6361d737b1e04a79813bf2c63995dcc2b029f30100f4e048d735918f3f188485
zc12881ac88263c63db1c9cfa13db1f76ec879abd84c465e2964474910eab7dec984a2060b8be05
zdcbad190ca932b1eaac134581caa9bd929430b98b9eb48ecd65a35430879c9405bb24a30a3b76c
z86613e8e09c267e3008fb261cc3ce9a818aadb690ce215cfb9b0d8ae5b5a7881c61bdfa4422559
zba130d015facb80acea47c425aec68fd5bba37ab1d39ca8294beb7b7967db33cae541d5238444e
z245b331acf85efaf404f84ae7e8ade14d789427f7708923461f4ffd6ada96974665e1fd7afaf53
z2e307a653dd06d337ad11b1be2203e03f3b76f17ba7e7f855eb6a297508d91eb9fc6be36e2a81b
zf5081424d2ffdcd363bbf7e84b35ce46c973657e3a6e7a31d6de582f9bd5fe9e8f77ba0a53908b
z8203f2a5af03af5124bb9d4b7e6c49668583d5d1d7fe42294f209dbc2161ad5e68aff42fe9b957
z146049d696cf2fe720acf08eedbca4db734b7e464701de83284d138c7c31e6e16385216f77e5ae
zfefa754c3015772efecceac27fa9eb227308dd2bc1abf9eeee4bb8b0821a7d7dd747e721e71b50
z02fd5267a247ee0321416f043da675d1cdebe03f4e80f31379707d86d6d7eb413d333a72dd7f3b
z8bfc673676e2454d917afe9a1cda6f7e64979af940fe6b09249411d3c48c98afa61c4de8dc3998
z12dfbeac7cb99b7c3ef730d3cb1bda80c01744fd051a5bc4160d89f66b73e3dc0fc8cbc5a4b0ae
zce9e4288da625e44efdde0d15d9531f71e14bc7df1ae67be33240bb0b5bd42e270d7875ff00c2b
z222a764f88518bd1b712b117651af48b8a397c76503e4e73ef7d87388099c917fc82d9f05d8552
zbb8a0164000d04a296b3e328b77a19d1bd4c9fb6059536a9ce9e121b59236ea040f726be1607dd
z1d8cc57d53b9ab724071f42bc50379eed6e44457d5cf0b749c888e6ccfe675ab97f8277ee32bc9
z5ca10cfd99380b27c439d33b3fdf0063a1665355df89866613abc4d304e8fb261948452a408315
z18b052a9d54adcb577b9cbc403414118c3c72c6f92a78f51737f51cda2cff78d34dfeaacf4e468
z4d23d589fbd275248f830d3213cf6b471eb56bdadc8033674260d35b494d92d9b598b1b62cf0a5
zac21482ba6d1a7bc4caf7f306c67e3f8e41c80744d9f78f08f831995dc058ff797d58f3d482550
z5e0625f271c6df5d6e18c24282249cb338d7cb969dc8b2ece85ce1b662c7345cadc0d5a20894ad
zcee96723f3af1a16eba62e153610a3706a49b811ad0cad9f1f1b5db9cb80da4d8e91c527adb4ed
z1674faff212e62318cd450b559bea5d89e0904f8939474ede9978dfde440d5fdab0f589f54dc6a
z2cae01001451c0dc4198065f28a06501271ba21e129c6e1d21aae6c551c96ae222bedcebe52817
zc65f36b295061d6fc8ffda19c47ad28768ee230e87167c12268348f9dd975071980e1328d70f50
z24bd1d4319f3ab9a6aa4ca9e0e1ea5ca03303cf55c80c1df9c185a851add5b4e66c461a575bf36
z85fac5555488be615b407351622766bf755cd5b59fca4968ea9be475e11ac0e9ed367f08f9d8cf
zae81081ce329e3ae82315f73001121002b81d75218f32d918c60b3049aef710258d996c706cdab
zeead5fdd9fb3950e69b63df4529165fa3a62c3b02d9a7f900f44b3c1df80845de8417f90d8ac75
z1f4cc146709963216e85922a96effce50d0d5a4e73127dd7f636799fed2b6a6ee72ce198eb8524
z53bde0cf7db997068f0fdd45669112196563a510a0b7e7c6de0d7392ded0ccbc4b4e3905dbbb7b
z97d32b87195fd308109c2c36e6acd7dff13cc002e54f1d7bba502680f26f448ea152c0a9b25772
zb53d782d1de7f7fe0dfaceb9b0590560e37bbeeac006672f30481d7c15e35a461f7a2266154b29
z27825474c196c9b97691519f11a388ffd42e709847c8879f08d34140b75918f0831df6df02dc25
z06955b3ee4cea1834546248003e1af07b933aff6876e21b205649e5bd863cc7097283743e3996c
z305c284e77d3cd6705aac403e7862a4f6dc4aa2eb32fc47ffb3958a1cefeddd08ff221475b3c86
zd830d323347a390c48894975585de0bd5aa5e72f5d530c0dc5901ed1009a618e6443b701d53fd8
zbff144db1b37c16355e8b9f0f62e2116237c4cf154db6cb18565d5832e98602232aa7ed05c575e
z542aca9c56afc65164b87980206e64c4a88cc3ed47817cf2001e4d7b6cc224c56d5ce29acba25d
z33604e1c9db9682b1c5f000ca4c76254e3bf2269615361e2c2b7bca85d4c40e9c69545255afdf2
z8599fa0efeb12b64533af0076a3a2ab04a726b15086c4b47119454028f60d9110c7f758e7e3860
z07f04c8c9eabfdc50ef948c7816cb80c1d66071e31ea19224824a2442428c7c9c4d52547e82983
ze202921135305c0b9cf891e56060cd76020bfced6865a06f8aa79c5ff3c7619c3eb70985a17894
ze5a36f3295206cc918a834eb21457aca4b2f7265d45846f97b641077fc8f68f4d6937bb28437e0
z38ffce5b298a84c9a910211152f54e47ea696911a1443a625ec4c5bf27acea0143b76ffae7fe87
zaaa5d16cc88af2197a9f1472105f87aa82bbbd8da53f440ca2034c924b6348eb779ef87c123c4d
zc7f037083eac36ef508619d19ccf9ce54e9e4198b80ec461ed891f9d3104ca190e75113a007add
z5fd7de4e2eeac5838dc5cd100a994a6c3068d2e49de6862250665558cf67df32d52f6f12e89957
z211f92c1fe2c467ca49b5b1c73ff9e14a26c5c86801e5c2ae51098de52fa41efe49c22b800f032
z9835dbe03480a996f6e759c9a7fdfcd825ff9da08bf3c6ebeff0f6ab2e8d99e533599cae24dbc7
z4d4b13df97f404edf332e06d5f9925c7e81f61af05322764abbcf64184a57411b2c7ad485260fd
zfe8aa71b95a3eab2d0c179466629ee2ed8b0ef549551e57eef124ab067b39ab25ed39a45f553ae
zaa412cff1a033156920372775b0ac8979cbd872814ea510b81953cf8697f46466d6c8a835cf60f
zaf242822d30289e29e9e8b3fc6cea44c7e98ba0114f8f66aac450e604a5678349c7922de9812b2
z31dc17b53af8ab2fffe0520ce5febb1b9cb85eacc8721fea65caf7622ea8d19eb37770cb859e39
z8d438417cd95b354da42715126e5189fb05afe1d1d90800cf9797775d7dd1fdfe0a6ee94b5c3f6
z8877b9532496fd5f4c3eb311c8f213a293ebe04a0836c281fffdfc5c156b58020b1a81dae12c2b
zc243f390a57d48de167a39f9e7b86520c8d98611dba06f87165c82608e0e54a7427b3e31d6585e
ze722ec0a7e8d5f33b57f1fe2c99eb1722ff2366ba299cb456b3e40850cf2c0df0325c6f704c92f
z73ca6284527c9ae2a49ad2b1b1c7285ad882b1a37a9dd2007767befd15c1b4f193fead9da0d90e
zde7621953cf5eebba0ccdc4db3f87557bc04e241dcd6591826256470de21c10cfe6b45ce10b2a6
z2860584f0a9e49494f292df9a84dcb111e301d9f41fc02c601db4019c6aa8f97808ba01314587d
zea3a498f0112b891bdbab811156565d6dec110de80a45c43c7637f21cb94dad4eac5608037eadd
z989f02207827ef431231c61ab20e2a14d2de7c0438cc2fb64cd4b47acff0e5828b95f84f911e81
z3d582de281902e29d87d7626123b865522219ee126ce0d40e05792247a8bd4352de039f7ea45f6
zb565ed209e727d8384c3b7acfec9dcc344153df67aa63adad20ad56cccb470e813d161f0ade471
zb9262f1dd10b298803341f48c1f9f1e5d738d85e18a88c8dc61edcd250df29556d513282819f28
z75bc377490442c5a6b7cec2035b927f4033d13d0c8bda3d4b381c051ae2b7622c52e811674ce12
z19eaed8d4de51e8c754e484407364e8386a890181a257ee554b101b65ad712b94f1e262959aac1
z03efabce6721c51f21dd45f1bf536f2b23cc1319646695516655b4f4d25970e7e8ca633e1ef0ee
z972c32f20369b0496bdc7bc50123e765b82299354753c5acdd13ec5c782bad38975ac0735c17e5
z554dc99831f3dd87262e138adf63f202c5992353e0b0df7b78d6d7a1d3cdcb515e2d3aea2e3e58
z9aa8120d259e365eb7972aae9a2823af52639cd47e462cc95609237e5d877e8270c2532d84a2b4
za825320369269d0965e3b4e9b305088db1d6b0d530fe1f687786d7b91c11634533ed7c14c2d457
z3ddc1b746d19f13b9399a159be1d045f6e5633b0079c95337d0ab24059dd281245f84428ed6e76
z61494738a000cf724471807ebc0116b5c078ccaa4a5485c0f60490d83becb94e1a68f53e81e710
z36cf81a7eb99f3bd458d5223dccf0ab83b907f107230d74ff1a449894baaf9771190129ec00edb
zba969638f01a33afa34e39ad367086a31acbeb9638613d324ff32fdb4b8dccb89ad47541defe62
z51146322daa16b9fd0fe7d9a3a6928297bafa1915f012fcf6d6f0f482e782d8c98e47e01e2ea46
zf992aac904f998e70167df6246dbaaf7f9406248d70d13ab0cbccf9859191a3d26f89f47433959
z114599921da5f4c857abd945e0888632819723767ccef8b4505a0742516eb2b03cfdfeebd28bab
z8830ddf6b4e114b2dba5cf26131ef8aaf9be0d1d4fd2e4cc01e930612c0c6c127caaba0acf09c8
zafcf44c9d2004d7ad597f6d8813dcaf63e1d84c7290a62d11ef0e88cfe8b4641ee13a1bd4c0d64
z6f5e7ecae656f51c639d87d35ca0b2b3f7e7fbd54a7393057bb510abef6c4562a1dac0e94dc1a9
zffd48716c657eb41b08df99bbcf6db3672b50b454a2c134be9d97940e7a30c87bdfd9ec9ed7dfd
zdf98bcb83dcd0eac5bc74443aa0d6e3d36bfc9db7aac206fa6b2b0fb272bb796687ce51f5adc62
zb01eb15b0f502db810f5665583237791440d15e4b9822927b63bb454190fa141b516851b67dc3a
zdb40e2be551877dac1971133d8929a6a22ebef730f5a325cf72b7ec19739534f3c49708fdc8d0c
z48e91f43332ec9fd677fba09e82f4614961d36cfb4a7e7c21fe36af014c34a41cc33fa2859917e
z53b7c5f955f46623b5435cc7933e9989ce83b82ad2866ea48d2cff84897fb3fe9d97d89baffc9a
z85d68fc90fd5694d24f472916dd5e9a193e26f8935ed0facc53d13ebb27033e2c04d5a78cf7118
ze906c9daa6d0889831608e764c4d427de4017ba09b3f55d1c505a2f28bce3400c78f99ee6df124
zd9afafccc42521ef9b67d8d389a7201f840b4a02bcdc049efa0b412d059f5aa21a0051277c9ecc
ze64bb3b655415ed9daa55d0336a0fa8149402b41b88ec4138ac1fc475593fe186ca5d28008e2a8
z48493de86e95e2fccd81b595b782203b9dc191792d16aeb37762adce05c5e40e27180ccca5f5d6
zc4242fb12631d527827aac51363868d491e5373873cfb14c9b031a0ce5237132c1e99f87c92bc7
z63018f6de15cc3602a0f56987f44471acab536c62761f126e394e5e5f265d89f0302bea60f3457
zb770160b7e7cac51cbf5c4cbe833156ad57466189e0c71ea09a8646ecbe809f44b4df177cd487a
z9c8e29a61644c0fd843c734a4e5cac597811d90d457d3b6e651065d0fb7e6ac9fedec6e95f88be
zf454ec11259dcda93c5f721619d156035d94ffb39269ac4ca51576154f78057287083a76a6d5a0
zf1edb7d06c71a8881502689b0e03a4dfeb5514025dcd9ee26af6eb7abdf3d74c30519e67b06769
z87185b4e3855e5bdf7bd3d2d05dc3e4121e7dced2098be24ad7a0d3fda20d0e0dfc52f7f10a762
z807ee0c1603f8dbfa78dd23cf08e67287da819641d7d8d00b9311b0902d85a761dc9456b248745
z49b8bb11db1c542139ea660e518516873f1c7fddb71bdb55482a5857942dac4cf1a4ce998d86b2
z0b7d6e4ca241942643bb7d533fbafab2fae23500e9e46c0ab892296e674d142687ea0a0528c8bb
z65646570719553eb752514dbe8c70595f252e3214feb6fa5323734affe7615f0c7a8d0235e4b59
z8b64c732542d9d05961797a96beb2f6360709df618aece8629db121f71b85878471e8b22790e35
z05f4c726d3fba6569b2a9a61f1b5a337018bc4f34ed0d83a98bfa09db5bb32f214fdda525b7329
z59476a82d89d8a27b82e72246c45ed4502ff017118bdd41f32defd2b9eb232695277966cffbe20
za11c27af1f5957c927ef058b5f5639d3ccf7b830e35ffa98f5c5626ca04b89674189926dfd056f
zfaa1df31eac1d8f73d2cad0e21b116c357dc76897ca11ca7ac82763e089fbf2973ccbf766af1d0
z192b511e8f27b36246aba76fac96eabceb5865220cfabd6c2e2dd073bff27d90d2ae3f91eea537
z271223844286222a2dfe83c4c37fa0c10c06159b8e645507b32509097d6eb24a31294136100b36
z139ba6e3314dab18037249c6ab5933e2a3dd4dca273004d6a24be9ee73cf8e99de64002ff8e81a
zc5ac3619dc8508abce7cc09ca7a840e24e626e63b1cda2a0c38244c99720a0ff687b840ac29fcd
z9bc134c52d6c005f98f52f915f61b8de2e2ff6521b1439fa08ecfe99c82ea022bd38ee4603418d
za029fc166cdd29d3d11c6bf99aafdc9a02e0c8b3d3361ca05069efc52899f25a309452337a600d
za9472ad4463a9f8cb5bf1f743a4d3b44361fd4921a8e82e173a1af81628be1836a4daa187ecb10
za10ed100cdefc2144de71a5082f522083a106baf35d5bcb0b7324922d5b204f93ba7558b294875
z7c7366b8290db04508e793408c5193b4a2a6754b224543031dbb4a5b786e648bf294989ce3925f
z2869e0369aa2dc8e3a9677606f31dd0bcf37e932b0977ab00ef0c85a6034421e21ac6d3dfe9dc6
zbc264eea4de44e887a49918d03eb1670dd685568896a5ff5bb4d0599a6a486ce50b31e3a7fbb7a
z441ab9fa39d3d710a45c3d3736a050013697487ddb4b59744880e2eec1f4966287f47aceefd443
za6e4a417ae7f2542ad3dbf723639e98ae22b8ecd84d607c8e27f466706c0f2a00e5ef11262b57c
z33c7f4ff1f0a48de8f9ee500c6f8ecc6dbcdc344e218a56634c077220c2597607daa722d1b1e63
z758cd8a566435c621204cee4ccdd61cdd96938fe3d1bd6f316b99ddcb324dadc5af9ce20cff95f
z65484db68f540b6f232ee7922ff7ccb51dfdb48b5f00084d7bee6c478dde889fe389e9fdde80d5
z1fdc8d6c9a3858442eb5858df761ceec7a240e61336d9faa70fc8f1b92be87a8abd30f0f4d1e5c
zf404e65dc6dd2bdc718ccb2117db4243a402fc6dbb5fad6d7baac889450dba3847e86cb6a2e989
z6c6ef6f011745c029dbf95d17e51237458e20ca8b5e69e6f2f6070f6cf907039b21781e3a10835
z4190d283d465d8e5695d7c506047275329e307e4c9ee7d7d70c1f8f528c2f44ceadabf767d5bfb
zf1df5d3cd93bc1ba4d0cd67a0d5d06f418beaf9795a7cdfc1d2c7331da0a216054a10da4dbd9d5
zccae6c462c5ddfe95aaea62d715dcbd677767afc14d7a3d68b28c962d9252d2b27e64ddd6b9701
zfa2101e258e8bcac26791fca2fa21f1e00d493c40c97aed418c0a0406bd04ddba86decccb810a8
zf25b92605db115d8e7785d961a19534822b4587b351453b64ccdeb94daa68d6cb7cc6c24a1dc94
zf2a8a717ad76f32fc0e7947f46a9c518b1ea14149b0847d8088ad5ea2887859c0153b06a9d2ade
zd2520b7c2bb886cb3db0c5cdee53dd05f59fa364b97d5b3c611ef528e4374dd89b058ef010c18d
z90e4564164b1bcf03e2148f3c0562bcf9f0cf5877aa298a396fa843d8917b119575770cc7d6100
z29d8dfaf94c2e80d865825f5d8323530c4c2d39184ec88dd0e464e8bcbc412f9327e2b33100d5d
z1b87bb03bac6dd02ebbc0b660b2b359bb8d89a2e4cde49d35c328276506e38dcda418763e56cf5
z515b2c2525760f4e6a4eec6115c9455bc9bdad45064c2c0345ee330916e80fc488a776db208d2b
zbf1bdcaf63852375e9ca6ed94ad1565967933614c8be1928e4096cc61ce35d84f93ee765d12d3e
zd82b7192a0ccd25642527c88f2844682a45a5acecf3b02745566517df422ce5e554845bf2676ee
z107336bc1840366ca82a65f37100762b92b34b03723d3adce12350db1e85b07a28f11dc75b7994
z04c889adc70f6fc1b509b6ef1907168b0a99edb809c848dab2f96f927c58bae47d50cff1c209b9
z16abff78b371def8e7f4a480f3ebc1943a5846fc3d3f4b312b7e7276521cb12a6080f1abd01318
zad5b93a856a40c69abc732c2abe241d5e21892b9d03db78cda3566bd87d3299ba6950a42abc218
z92a5040e87b56f0a746f07f6efbfccc72fe6b1c5251030f2e2c54eb760817c602d1d4f02bf480e
z1e52e4d6598be74e48218289c57f4e49557924180d41c58806ead56a33b84229d0497076e0414a
z64e128c8e68008b7f90e61113221bc4bfc0324404c47fe365f2a5658c277bc34e56a88984149bc
z981416abc92e4390fb14d96f71438723f529fa0937524b3a332565d1267ebe5aa5c35a0ec8221b
z58101bbb4363c528bfa6f6a734cb5a75e1ba3509dc84e4b70510a3a7345277b618874907215dea
za5c150904d80c8162c48385eeff7a386fb2af251c41f9906d453689404051f08d7561b3e12cee2
z08e4bbbd58ffbe4357e4d7edafc39bf7b14bf9d71b79b44efec1895ca2fce32acb05072e63de63
zf10e55d6a80db9db2ff24e810773911e12a3a2d5f80aa5839cec8c1e2207ed1a6e9922a53435ba
z66c3796bbe54f80855ba8c55ea9facb605911b38f2deefbcc55ded8e5d7bc4e3e1dd4464a30c56
ze8a8cdc2a20892eb690bb995e1cfadaa8bef044b5ff8af15772d68e4a50fe2d95a046c5bcc7e05
zae763da94ebdc54d58a02f954be6676d8e5722098a1e3d4e4bc93047a064667edc369d016cf4e3
za04c94ee13275b951c7e9566951b63b6dd3b2ddf773463ac380cfc2984ef05c419fdd42c988e1f
zfdf6528df0e00cb087985d33426a7862ba73696ebe8a42a20cea0ad37b77e4c3f4563a34c6e62e
zf7300a1abec91bdc515a2a93775c886786fa54265f21ae9edc9338a468c5510aff65e7a6abc6c0
z4518af8dcd239161d353a61d552d60550d94b48bbf2051d1dab19282883b300299aa1473b43643
z20cc4349a0c312b3c355f20d6508c435435d2beaae86a794df19aa5bf4f9dc38e56d4433a92e46
z3208bdc1cb76e9756db22a265efb23210ba37a68e0d0469a84e72ffd2acb85fc2fe289e94fe0d6
z61705a7040577595ab4db16581d7190b44e1855b0becc841b7b8fc77447b315ecc31ad18209c42
z1cb15ea5be47ce393030809cd9e778f723b354d96d1bc08d80667dedfadb371f12d7ba604409fc
z93d0276d5c382967742c84bd3993059ab5bc0e97685b871f81374614606e52166a2595c7fe516f
z5b9d17bae88bf62efb7ac37b8615dd73b737f77381dc29a3ba63ced5d1335cee80292af4df5875
z44a4eaeb4a6a6f32bbbc4309bd6f9c1feb4cc0f0beaa7e252aa3588540e639c9e6978d227bf4ab
z595859ad3d1d91b289b6784070b6321887e58206aab25010f410d93e3e75af5a583fef52f45bf9
z8f2bcb063c12fa6d2ddb2eaec0f31a5604c989bb313349e5404934316eb96648b1f16caee6e59d
z2565b97e1e6c7416d5f6ca8048369ed2e1a235f36f2ebcc9bb8cbbf20d5178dc54b43a4b1f309d
z3e790f1e12f4d9b25bcd3a59a1f4d31e336ff7f176f33b090ae31de3310081c846bc457e9eab87
z0fccd692ac009cac1cecf76d955133800dc2fb6fc6ba641fc460df96a42f5c224fa3b2093bfc28
ze984681c4be0ff73c5d22a0352c8a1b469700d51333e2560ecd3378685654d3e35169ca8f9b946
z9b70e64753a4e6ec8a6d5954d1fa8649a27e524a516735d8518cbb762e9e9a4913698a8f1ee1fc
z4afaa837e974c4d9741310eba8f7f2139c907005b633e5121efc4e70115b33d2956de9d9cd7398
z08da023527c765bcbde837204fc8e1f75c2c68ef1de3d1a2328321285b7372c36a511027db2969
z932d359ea98b3899902c1e3d37f5e3f9648de126631cd13c9ddf23f8615f6b8e2e0b5152e69591
zbb0b8ee23601f96d17c1f5e8a4296cdba24c0645394fc0df42de76347a86ebfd452424de88f86d
ze3e6ba50661740c80da1ac85b88056d0d999d03f0f9ae3b809ebb83d4becd113af49681e7b4ab7
z7447849f97a20507b84443fd48dde8659d2127e76255baf6962ccb23c52dc46e9b31bfac39d5f5
z0a82a65dab6347c716124354d71cc589f68eaa0bad879f7eb37a3708511d7d99a2d8f3114476de
zec2426dbff31758893d5922373219b17966f0945ebe9e9b63b83e94edc85e909c3a6bea0133726
z4610f6f7e22ecc016d
`end_protected_0in
`else
`ifdef MODEL_TECH
`include "qvl_ddr_sdram_2_0_logic.mti.svp"
`endif // MODEL_TECH
`endif // encrypted_0in
