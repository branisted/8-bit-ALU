`ifdef encrypted_0in
`protected_0in
ze74c34e226135848fe16db9ffd31815111b6d7fb642c521a3f628cf6da949865580b22efd062a7
ze90adae0e65e66a2c36a587d0a790699161455169ed55a01f2084f11770a774ec4c588039b380f
z6de9c5084882a40b79a175f5c2114b2b6d78b070cb806e1c0aa9258297f4687ab308bc470f0040
zb0b1de382961eeeaf2e279e1462520fc31c119af8f2b214846f56c2b3cd2eadbe4099496abff18
z15cec83ec4a77b868344aa20ba7360908f5c0de2a79abf8b3534b883bb12180f68b5d4beb444cf
z3fba8f13afb0abfe8fcc4294810f75afe452434d2d0f1166236c82f76edf1e12979f04bc35693e
z32ae028996dd85737a8f5adc1ebb94f39c940246e887647b64782cd7ab429b0544c173176cede7
z01dfb26b1f73408344a52b7e1f117f12bb9c8077b34876c2e6fdc085981637012dc9754765e1a9
zc512ce062e0b8fb16a214591f5c81e1353b900a611fe1f4886b57940b41b7f2ce99a7b84b04b90
z916f717e73bd10589c81e207ed77ec660a8cbed5b487fa50acde1b055c8870bd8676023f21ddcf
z9c98cc47cfa2d654ff1365d1f45035a045a66c5dfa82790502623b57a3af03bf0f0c0d35b51558
zb8b5f2d29acf03737a9ca2a053b7a8f06800d50b465c41b30eb585f62f3d0c2c5a43bc337624e9
z8dcac249110d9d254b0bbfa98b07e9626524f0cb9385477931294148de8f9d4f776e2574949a4d
z351b61ae8c8b909229ae5d638664f396414d080174af55041c7abcf2568bc1f30322a5798e9561
z9ba8a19ed48e77858cdf7af180512d15d205a7ceb8018c94ced893e8ccf8e7a349abefe5bd1b77
z5ea92042a386bd26ea3f545e5d21cd8e0d9ed817adda04b62775e4fba2cb865f13995f0b08fcaf
z520f41e138a864c59c12307758dab92e31a9cd6de816f9770f2f7554b1b0d8c70f616fae9f4891
z408226c56412cfa618c1f4bed02ebfa0131086fa120048570241ae18315c3c1ddd27c86412173f
z3114e0c9cd54f3531efa139dae0e0e8e335bd16c9944887ea653c23d79b4cec332b6f697dd9817
z825208370ce9a157bfcb0238125c6e1edb44a21ff273e7443af2f1730c36c52f8a079fc2a6cf77
zd6d27d42303aa3702e88276acbe46825f394f0c6f6fd70acbff3c9a57f34c72df1164aea9f1a30
z8e4307869b3ff3a10dc460047e60c5b73d9663b982a69a925938c1b5f2ddc91a0ea67ac3b7a7c9
z57d194417a0ffb37dc4235a7d79e31f307bfcfa5aca8afc1a4a12eff9d2d9c6d441959e88b3359
ze72678a581cfacb2ee8a655a132b1d38e1b8360bb431a18818683d57fbfa8ceaac0da3e9ee7c51
ze2c7370a26759b0cd5f58112a450b1d6cf2afa684c050de6f14cfbe7d61006f2167a08a2ef2fa8
zaedc49306b1b6ede159b08e20bfaa312c496375739a7ed57eeaf4c36260cc1a9343e164b43d40b
zdd51bda7ca60207872c56b7a92419eaf837527f3332095c9df7ca22a7c2e740350319db67ddd2a
zfa7b60448101792d75ee452d46bc937dfff12dceb97faf13f74f36e01c98d78354fd7280b39e79
zfa03149cb661d3d108a64411aff17c37d29e4b20e05dbe886f4f84aba85e8857bf5d301767d902
z80d4231500435b136d1483f45a544757ee7fd9ebe9981604b6f6e504f97acd860eab10ba669e0a
z5f2c47ba2fa2f83d98f2786ec2aa23351f7e6254a4be9a82b4bc20bf052c9f7d5d2c2dad0e69af
z54e0aa8d4ee2495c2fb68318f90b41d97537fd797ac44a7dfb120051a20d8f5e3670a9ca365f62
z75b3b881e9aa34b2518e1a47c88eddf03d4ffa9fbcff4682da7364a47552802e119125ac1cc357
z0f8b04a0180c962edb2c96df27e21d364fc9d08f52072933eee99cadff66c7ae67d3061df334e6
z94820e917031a6b1b53179e5d0b8c96634ae7947b7e83380a7764af81bb163f334757c667015ec
z1c0ef47fd36f15a08299c549361dfff63acf122e4f91efaee682b0905e2d168795ff136ba022f8
zf9cdf01f9c25150f58458531068920fb1054b125f9cf0c1996aa1b1762b3bf7397534fdaf53017
zbfc18813cef99fe625c8cb9abebdbe46b80da755e045c73bde61f94063ef6e813264e2abed2180
z6eada8a480ca10b18d032c43b019df6c3437807ce0e16a958f971d3e4eb8d49f9b9ec21e21a478
z881f2a6a5478a40f39b93fe0f0a25025480d534daef7f5e12a97c4abc4a48a941f4a6955fd0c99
z2b1729b1ea5efa95cc4502b4dea69513c85f57b9844ae497fc36ed5ef9cb624daf89dcf6fbe87d
z36acb134190a035c508b3f5eaca6e75b827edbc598e0692ee50098e0141cd6212576149908392b
z6e7ab12ae4d76feac6fa3f96766ffca860e12fc7c24c401ee3db06f1fe5d559af7ab33f892fb97
z75a248ab7e5d7583f4ddded85df2a846a651bc4cd6b0556ec4b3415c63d2e0c6c97af1bd77cb89
zea08519c10b8820278233c8468cfb9e5a0e4e16159a0e59d81cf568d66b6682cbca843f0aab53a
z46ba422481870f760a815752a2cb0bf43b1c20875b5478ef034ee065819a71e02125112d7c509e
z0c05f9b6c8fdbf2fd4d13c4533b07d10c757325bf7f5e1a6c3fb0cb40fb20f5a1d03a9f93d7b50
z968ef97d9699640a49963809e63efe1ae7b96f88360d322fed893fc3e7d809af0a6c0e74a98cf6
z291670880b6b456b4541c9aa49a9a33b8f98d118190658b730748136e22f87804e1aa0a1ca2818
z82989381e814b6d4a99c556907b2e156f92c7d21906e2e11b6485fd78398d63914102c579994d8
z9f6860bc91ea249702eef98964382177e5f70b92dac24073c37b2bb2ed71188e4fdd3f180cd9c9
z2b9420c556ea93ffb4348c6cbd1cd2d531da9515e47a25aca8f9f9039da74656401e0bb808c277
z6ccc22f5c0406db2c42643de7a69a9aa8fce25e20c6fe45019cbc493ca7bc27bb456a8f3299cc2
z4d908b0b42ffd3f1c3191ac0249a195ed3be001b8cc9bb9133704ee2682889471b2efc318b6c9b
z571d40b391413ec04db6ffaef81aee6a4b8ff28f4e2f19bca7472fbfc54c41926f5ed4a9f3eb54
z06097c84c9844e8077b56d5c0d330bc59d1c4878ef72951f4c3d66dbb5aaa32bec881c84714962
zdcfb7d0a6472db91bc8a5f03e8746bfc118cf5244b1c26a06686c1c6a3086ae512d3a2dd667a01
z90b8ddf822502ee54df0ef44b7a1f2ccf9106163fd71e926bba7f3fc2801d366a093b1c9c0f470
zc78736733542a26f52655662639e5f1ba842f990844a67384baf67350d6bb3bdebc879b1251bea
z30490cd4b92027043338c6ea1af30e7b136548ab3341a99655b8b245393f8c089e6f3eb0f2c414
z9b3cf952bd5a06d23f1d6e6d59725211841a343895f9d85022cd997e08f877dabc043a503eea5f
z2de499e6c0ada9911e8cce715879a79780b5f863489fb318677f1ddca51566288fb3d9d3c19acd
z3bbfb2c515b3da9d2ed38c565d6e07322bfb71dcbb82b599f7d0907eb68ea1e452199d659a8252
z2bf4c1059380c4a064c75972c3fd75531b63b108b4aa47a9d74500aaa30a8b893ebe9c0df92eca
z4e1cd026251554e2bcd1ec5c2855ad9d0831cf18ddfac8f88e7a93c186cce1e6a2eea281ea65df
zb0cd0634c282cf5bad7ef0f25c1dae5bde1951b6f350469f00c465b7077e5825fd9d43ffb45740
z1ba2b40b1b2a546166e84d189aa758884a08b9ef158b1b8b938ebb36a34a1674c719e6296ef71f
z9ae6089340cb4648c46760833ddb6efc85cc21632811f69500a70a8a702f4c26814a29f3e25c8c
zd908a381a7cb9eb3a8dd1ebdf4672641294d74fb01e452eac2b07b2a7b00d7063fd56f98b00f96
z3801e58ed1b9abbcbbe71af805b39682f3fb3893e018a4757ee7cd757b4c613598d108e4cde930
z7133e898c47b91a675093696d7142e4282bb50e546963ec10f5dac51ae1123b9c600281106017d
zdf7cd426fc629ce3fcb1ef6666c7489f521a05cb23cfee91a9ea7fc0df2760545d1d6bd2caec8c
zdc210cc6ce8185e40b03f250d68df39fbe5cd374d98927f198f4153aea24ebb26b219d25fadfa8
z5e6c5bc484f699aac79ccc1cf19d660cca52e7d20cebee0cc24788a7bb9a17edc65cb7676c0e60
z1937d034d29ab585641c791117061596bff0f86c2b1e46f44055a756b94219d9055e0f2c9de483
z7fbe885af3306f94616a6be378c3f95cc84c32fefb49a7927a13da6850f22b77e81471b649a258
z557e237fad4cbcbceafa627dfe1b375cbab96b4cf0345026b147e3490b587072ea1f87f3b22c94
z60bb30922683353e9ae058451c674c79cf844267fcf57c773f5155c40312e920fc49ab106d82ce
z6383778c8e77952b330897f8a2e7ac054eda201c83adb19c807b5bc5fa4e44643efaebce099aef
z14cf44768d36d13f5f077ad5e7b1e6ea152e4f0c686255190f080bb7a091df6583c262ec01f3a0
z65b618bb6f6bf52f784afbcc9802d637e6c0948b655ecbb562080a7037ad77c3bf777de2d76fc8
z2aa123b79a860b4cbd15a52a3f0a3f3c52e159a2a2f8ec0d06ef0c0df4dbfc51d0abe77f1908d8
zbf134ab63e04d5ad0b715ce8e14e37b772fbcbd19f0fbf81eb7f81d048cc2fc32234228b15d825
z1a4f5730b615d72a1f739da2dcb63f6fa080351db77e3aae48bffbcce93fab2afe7e41f94bfcf2
z84dc670aa12e32e5a351302c46576f9445055f5a265ff380aebe6491713312c37512d41a91ceeb
z528de1c5413175afa3ec561b60a6060d3c68e97e9fcdae019e3a344663ff5541267de3e9336f98
za24afa35ae1baf247cb2800d610e61f28e69b9d118a91a36286cc39eaed0587e0a4aef2a9f6f68
zdcaf9df47e14914530b4e0a854291631449d435fd6bfb04842124644f1356b34171bcbf8eb3796
z8cfa88a6e43cafbf8f908193265c14d2db3ffa35b29de0cfcc0608299d2c24b2b88c9385c72de6
ze3538be23acfb554eb35591af52d25516697d94c2b89b091daa29e3bb189505c5ba699990d8a0e
z71d828cca1aed16f8c66dd3c8244b9c784b15a214c50925dd326d5e89eff5bb480e08651dadd82
z06d467612dea049ea4bc3f83e1501d83c39b6b24128e2d174584423ad429dacaad7e8cef0aab7c
zdac02122136a874eac821e190e889c83bdb8e7243b585cac061f9d8efa2bcf82db7b597d4a971b
z5633c3f1e6929103406e9c508826b80e17cf2daec8267fa4ef65feb376d908c4bd54aca0902676
zbea93c2a848e2a585aed5fb8ee991d5f1a80576d29f817e2298ddce2e1137db4fbb76059eefe68
zd6fd46852fa6d338e812ceb9850cdd1072af737aebc5a49bfad4286e280b528f28f2ae80b2e14a
zc8aabe6b056401692f74f95a0ee891309327d7d20d387e052c484c622fb2a0997ab6a4b0bffb75
z3059226d8fb664ffcf817f46173af6e566017397f8c8f577fc45ca2ee58e2e063b6af33febf78f
ze84a9de1777b58ecdc462350ea7d34b121d3ae6e1cb81ae0ff44c890bbf48ee74076aa2f5a2357
zd78c15d2deebe68bb25e668b001cca194a1e2fc6486546196ac7dc7047de4d8a42f00371eee331
z24e91662232ea5f670aa09baaa6986b466fefe43b020d37d3d79016e0749e2fdcf4b8594f35705
zc1d392fff474e3a2fbdbc239ec9416f235efd5ce8ca36f78b439605ede4566e05f56cf397790da
zf073ee22045cb96850ebdf14d39696499cd14e02cad560efe889d9ffa4981446b0634eb04f3f2b
z043af7ee76ba052309942cfdf4d7530f5baa61199e24332c334d6d9b8aecfbe3339721568dac54
z11924a312b84e675080af74ae84fc2d9b2b432fc2f9f63e9e9134fe9516f9f47b1723fa6dc1dca
zf863fea4b440094b31714170196d68fabef3404a3f3d18778218ffa05f6b9e3a251d80d637bfbc
z62b512d257a59c6b09372f04e874d5f9acce8d94621f673ac5183d6f70264fb67bc2f8fe69a134
zc3e52585ed23a931f4b5c0fe366670576a02e837f74da1aa6dde60a03be5979bd6c6fa5a76cca0
zc5a35bf07bb8858d75931f4d3c696aba96e6742eb455b79cd7be4b20b230f904eb447f85623f57
zdeebff5fbdf49b57b46304c54e358f58f509a7d547754dabeebc6af764fcf73b0138fb22fc0580
z12caefe407aab23f75cc009b93a614a8255bc90bf5142b98f6bac833bf77a308ce05548d0657ca
z1da1a42e6af8b12539ecaea8798da520f8582f44d48a288e020552c0bf3d481b83ca5a1f9fa8c8
z2343208bdceacd6fc516fafdbaf98983b62c1b199f5fa9e4e6bac5fd54bc87505e6c26bdbd0770
z0889e6cee27f89259ccff77409bd77dff759ece8daa3c7dee108184ec659d9f5844a8dadba5581
z1bd1478766f562824c2a21780c23fa5afece8e2f3147869705befa314d8d177936e5fcffd08517
z0ac1e743c3c2ee760e0798a37ae5d0f0bb54752950ab896b47a49b6efde1f09cf864bf9f0a89e7
z197034e6501fb5440efc28072647450685aaed044a79dd12e450bb61610eec4349c000fc38684f
z42a73730630c0a907a25ab49c2b8d0572532a7d72d8e1a811ee58d0349dd15234ea915db1e8404
zf02cbdc3166caeef4ea461295227b4d3a68b9646be3a70f787203ff4afbde0033548e1d052e732
z7d7489960c6880643856fbc84cd4756a1f860a17e3fc9e7a81f78f01289ac8a55d0f9b44f1d17b
z4ad2d5224656d5d24a213b3c421c9e27a1f17405360b2eb37efb85941db471af9f6808a5d18424
z8f300c33314406fce347962f0d8a9a4f74fb5d2d30e0b0bd1b780c1ced7fc33172cf7453d6084f
z59a22c421b18152b7afc5f14ad170ecb75cd18d139a69d15f8a5f2b9b248377951cacc8c9d2a41
z67ea02061983ac1df916bba08eed8bfd4c6c0e6dbed591ec424e2e05b02c1845c83666a766fae9
zdc057a7e99552d33adf37c2f0edd6296690e6c9e1b067f6397befae5837395d7d5f850fb2ef871
zac0a532e84ddec71a0e4d27ebed9d1de481003fd02deeb8e90b15497b385d7537eed884951b846
zba5cf9f1ea53ab37c77fab53bdbb4ac4fdf902cb8f0d69f9b6514d9ccb23cd0f594d772b469e75
zc533b53ae1a74d33853612e310ad1839f2d25ba40448be5b4db9b8edee64751da512b01c58cfb4
z7478b4c5e49a6f2bc2dfe9f0d453b3950bce1a9422bdc28da7a94a7f1dcaf6ccf9c6538e1c933e
zafea98e048264ddbe5136e05ebfac6242debfdc1b9a38498fc36c00d3f2422827c418c8646c4de
za0303afeb6743a7006f968eb698f89e840c092b7b268c2223c378e47f1d4a812f3458de266a9de
z476efe82704683f68d2a1a9d83ea9fc4a16fcbceec601deebe1f61eed140314de38e2a6bb4f2c3
z4c739c2ec169285e2e31e2a66b216cdd53a4f129100f6d04a2cf8fd62b0a9254db315a97e8d810
zdcac028221b46df4caa96264bc801c3307f07bd834d7e27de0065b30a1ea580817580be7fa867d
zd3db2db44ff17a721afc09eebd595251fd7269a4d56bad3c3fbf344cfb2f5918f235f68992891d
ze91c51ca3bd1f87a30b7486a5762bfe75c2a3d8854c63e9abd2b3e533e89e5213bd07b8ceca71b
ze3837124b8d8966ddac1eda3b8108e84edf0f800f59331f4dc63f8a3d4490c7bc4bb1f341bbc72
z807f201c41f9b6e6a64c3a0a087835397084e78e18b0b156325acd024d7f82d2b827356e529e25
z2118fd188b89e21194326f9f286fe59f26d56e6d34c8b414da5c534e0db8e99f1cb8c7f70a94db
z8bee1571acc297e344375ab3a262c8a8c6c6e2e338b2095b85cd25dd555bfe073dd0af7aafbe43
z719d1abc2bd09cb060f438a7740c6387ae641daa42ec6bf692b2c7a5b4149e0449c161ab485ecb
z8de1d23a759ab654071a5162fe25c546f388a238c8f8af9ab551e82b9e0f2032972d7fc5779d47
z8358ccb59324f07adca0c6b109d579482d6a2f5d252449d6bca2d542c05000a5b05e707410c07a
za29b0f47ebf2f4877197af7d5323054dbeccc0ad5d5bea428063b896714006e7861f67bb9aed02
z6b2eb28d33b428e0422afc2a76e208a243c530d40e2c733d81643965f5b821715d542e969fcbd7
z7e36b1b9b67b6a477c1e5c84c0811e1fbd2b4590245f3da8fc054a4773cf87791fc3fcb711d895
z96daed41bf4f37e03a7925324beab6028c508d9040f0c96e026f2a4757ec4cc6daaad64ec4d508
z39cd9ea760456828899fdea276dd1ac1bae16e75b32bc8b2e920e119fb26b1d91fd6a932aac880
z0f784c7317b572124795f0220880ad1d324b63815de848ba01674c44e7e8943908e5c442e8c3da
z00c01db62c66b209bc3e017c91d10028f6f37a3a6332d62d5089fe1938dbd9dcf3738b20e3486e
zd5b083305fb083493f62dc9443270e9c494a9709339b0d1b94806e577985d8116f92737c5720c5
z81eae5179a074540ccdc9f6b37c4bc738772db9ffc081e170b2f658d14ff18b7dd8d0ae9d3978d
z4788f325aa1c6e13b0363834736cec8c065f5fb500112cd59090936aa0a7f3ce2eac0c730ede9d
z1f50db3880888a8e6e50dfd3d2bfbb5c28a0fb15b55ab879e7b172646b193243037804c3cbad9d
ze33609c082d308cb919b10484d9c1f2cda8ca538abf5ff0bddfd919eb57dc2f1f68aa970d1b0a3
z72b0b184b5e94a9db4613355a1e33f8f999573dd9d4e6a890571843fdb789043fb8774fc95149c
zc0748a8cd2c35eedc3638cb8cd05f8416744895959a82f1adc8c9de525a1ee1ad298d489a96d5e
z8ecfd03fedfa9a6918bf538373209e7df04516ec5f08667c912e2172fdda61a959761add2e64b4
z00de72e9d0ce777307cbb2aad7b6a6f1456ad0992945a576e55a5da86a8d02fbab72c3c4f3254d
z64f3c6cbbabc8c58b0399f8b9f554e820c18c4dfa543ce89c23317c4c9f816267c4b6bafe04c52
zc9533305ae5765842ddc2d9ce966bd5cfd1e4f98215049b107528cdda8cca1b341fd9bc625b11f
z2b9f87d8f73104b6e6788e4767492a1f6f3b5ae4dbfd5554c643e9aee1c3fd4cb8606c451de32f
z8d4209c4a41faa0c6ae4cc334cbd1af07710ac6b85c60f8c572bb50b3ef854465c6950f9b7552d
z39bdbc3710e2d7ff318bad83e243df635e6daf10f60a441996640dd4f5b068363334c5c0a391ed
zcea8616c7518a4d7de3467dbe81428304e76d183b4744e56781a13ac4005d33b3dcd8410a31b26
z8d36455b4b9d174d049793e84b78e7721a180bf97e136b88f7d1bfc8f23cc1359418f789cbc91c
z12c5897fc1d3d6f92aa563eeaf53f73412b92c3f9f82d424572b843c458153130001034e7d4eef
z44163891e45cfb9a88048ddef52edae544a83dee0da2b505dd23a71d3fc7062ffb8a2da1b8203a
z05c4343b486041d8f967e734666f91c70f562e5fdb7502e10a5d0ddcdc097df69c10290794b33f
z44577fc8f799c19d92d3a6075d4763cc25b675929249280078b8ee176d97874ad2bdcc94635658
z533d27b570ddaa3035da1be3e5e532bce43b71e49e7e09f0075d8169256cbab45176a1001a30b1
z12590ddc393878122506312b2487bc142ec1ddcee528b9752e5904c04c9c36ed2e1be6b709790d
z6715a2a2c402327acfe6d69abd65fc71975c0cf6d94b240ede55d1a70dd14cc4ccd3f9b0371c0d
zc12a52e1cdc2700067d7aaefdad42f86be1b74d5a78edd83434df2356c9e5a0fc24833fb6d2799
z3824386575d1fc15460490a18f6a9629784218861b965b03f72e4fa0241d0732f05a2ec071271f
zd508dc2bf65d9a998957027bbf675b13c0e4d16ac7acd8e90a93863d25f3ca33d32b3463042f71
zad231ab46e5d38fddcf028a997cbeb14711fdbefdc6de0456696fa036bcd1ad106e8151ea45caf
z995ee2c1ea653e8ecc3bc20bc01ebfb666d77afcaab796cb0f335478a50894590a7570aabcb7ed
zfa26688725833d464a19f0f744d66f7888af2961ec7644f41016163383705e9ae2c1e7df2c05b7
z08eacb08d3c75aa6171b1759e2835986e10f269a6a00f600a250d37fb657ae04832e999cee5526
z2eab2e56960ef6a80c001e57100b19c5b473bb033e76d73e8b3968f2556d01181fba47a8cca7b5
z23411925dc903c5b43f2d91725c9b53fdf7fe38bd52d682ee49f6d04cbe86c7f8b73634417cba4
ze93daf83563d1ab775728ea7ca01fbf4b3905864ecc6c7137d29f5746562cb0b65bc49a84a1f89
zdb579add018dc3b95800a9c40ecf38399428b5deda1e93f8d60bc4a02abffe8485a16a37f5be1d
z95285e5eea0c3dd3b891aa23a788ee9649b803d07e072444f5a460abbeea02515ab223a529e4a1
z08179dd6874002f4664d84631b797b5b51f3d7fe1ccc7e05ed3bd789b2982c85482d71ead303ee
zd94ff8950c17e0142932f496cb6296f637d566e128e0337790a64495b77e00db2add7ce1d375ac
z4d2d145028ec3a72f98b16715be7086ad4bce755c1c9a949e4883ab07846d564ae14c2825ab536
z45d9c2e5cd5626104864270e0867db0aa541c39d1f840b69d584929b64b2d514ee9c33e35fdc83
z4ddfc736b805df349fcfebac04c0efb3cdc45a81a2ba815f03142f797a2c2d773ded785b2e38b1
z5ec7064696e6bfe8e26000e3faf4f9ac4b518b6e8b060e95c1cdae0d4588cb6dfd11b3ee958e47
zacf24a00390f8e070567c4e9596515e804a74f93fc665f562d4ba30f7fea4ad2aa4161ed1c6a46
z18afc305468ccbd79d1a9db4b65d6287b2cfc268026a4ff3d43289cb2b83f756928e744e5a72ce
z08d502254426d06f03dc59cfe3c35341eceefe053a122644208469902a454f414f1752ebdea4ed
zf37d63c0e96f445d22bca2dd8afc3c234f622658d9dae2c5d59d49d6e057414785d798e00ebccc
z0dd866bf9bd1980d22a7c31db873ca9c14f946da04e08d074639cbd893d47a0ad1f422651db22c
zdca725f7a13111515c02ca04e261366f917eb86dd4091a169d64c3e6e2a393462bf7608e5e87a9
z97a81c9a669574b03e5bb4685f5a7a27bd29cb41b504c231d344f88a10955c0cdabdc9c3a8c249
zd5dd0d2bcd0a9d8f7a4730762dc4253fe964e9b3ca8ac9965df86a03b20f155be6e324266ac41b
z83124206113e3350469bc87ce621541b43f4c128558a873d4bc56dd9cce8b28505522a3eb4ee9c
zd9f96c4b0c9087c65b20695b319f2bad4c3fc134204f4e46051edaea8ec71d409b8f2677c62844
z841e010d30ec2c1891ad1492fc2dba970ba9eb785689c9b4494ef4c788d1c400ead893d1fc47f1
z0a3dceb06faaf8965f21cb1d58a40c89c99861d60a76a5001cd0a97e3352442fbffd00cd731831
z5df3063ef61712cc39123ed38bcfd7286030723ed425447a4df1a133ea21ee24bcea6d75383c6b
z335ff216f6ea9de4b1c3f428286bba27232511d3186f3a89875b90a3721cdceb3a3e876748fcf9
zd7adecb629fc691168538c1a9d77dd9181eac4d83cfd56c60a92c77e58d363ae05c888301bc4bc
ze3f562bd6cd5a80ca88534d562618ffee539098b09359f0306fb7e5153d0c378c57cdbef06604d
zfdff7476151cbc662d10aad63e6fdda3d9ecb94f49a1c34eacd1c2f7e5989fd84b5ec449c9d15f
z152ca336d56f3febd04b2fc0d32ae5a3ef157c2a6825b4774074618d6b03c17ea245552b7bd92a
zc9b4499801542f4fc10fb57198cf804b155c2f74ea6e987361efebcfef879b1ac3680e3a36a6b5
za63c6ca931787a54396283ef449688252be3d4cec75fccc39b6e18432b3e0b3eee97ec786dc9a1
z5b046674f0ac2a4a6b5b8178bba721ff32e4bf81bfdbf4276fee00d632de035395581948e0a07e
z4a3fcec8de2b4fb2bcf4991ad482526bb910fce34ffb4f06a3a26cb180adc9926ea774cb66c866
ze200cfe15084966ce4f69936dce5fa7404d57785292bd24a29cd1b0206411da47024832e954c23
zd0603640ed9d3729f1f320be0df511e6f9d0d70e6d4e9d529325add2f63aa1d7d6a77d7945db4b
z1e5bcca00c11d6e6c332407e09b93caf4c1e1e524872df87c0e85cca52943e1fcd77513b34c3e5
z0193a30b5c936acd7d11b1f02f3207013f42cb74881a403f77ecfb2ec7f98d808bf1136f33401e
za19f03a369f685658cd0b287559a9cedb302adabd3743b69c8ccccdbed18feecdc1646d67b4ed8
z36777500b342226735cca3387e5c7a986aee72f0c8b81a642468c3c85c8974bbcc09f3f17e83b1
z6b6965c767046ed9e40960ce900716af70904147b883873987155efc2f51a0072edf0e9e8534d8
zd05337906bb45f5d09cb3074842f531281b8d18199ff8189d02b40ae86bc307f6d5baeee9a8f63
zf928058e567cf50fa7b98b02a9840e1f21cf764016b86d01dc6c0fd38c010fb24aab59ca59966c
z5c612e54d433ba9059f41a770d8a9f86c5eda2e6c4f8f1b14534282adaa6993f6e990710fd6c95
z75d45e184cb3ef077472464bb8c1039327677c46da67e8b328912b8cc95b05c1a8d75a6e6432d9
z111f90fd7afea4e5c443da44f663382c282f06d226ed4ddbc6291ad84770d44d023187a4616fcf
z2b0fbc5256de058ce23c62f594741eb1a3681e09f0a7088973800845e436f99326a374e78cfee7
z7932fcc65b81e522aafdd8d6553415c39c17516c252a44769db8383f5b8b20c6f2325e579c666a
ze01e21c9009606be869ad3a13b8715ba0e6fe32c746645242c8bdabcd837311df8c24c586e2d44
z7fd7b99c7d7c1dc789ab19adc8fbfa7a46bc5ab632ebc5799d996e8db703568d727b2f403e1e61
z7a0cec84934e58d9c637628476b36e603b74cd716b4a7cc646109e1e0234203077ded4e0ed6b16
zbd81768e20672d78aaa9ff99db543ea13f20b3333aeaf0a8d41214dc9bc26fdf4b3fafa77e5c3f
zcf8cd6ff5e075d1d06daf46d51b8a60530bda9ac989d866ee94ccc07e2eab1f6c5129ee39477ea
z129abf05d1603cb661b8a04d140c1d78df8b696dcaa6e82fa3164ad609f915efe317bd97e6edff
z3e34d8613a8b2bd739ce412794172f2e040d8f95bc335b93da79c6cf9e91e26f25ebac39cf74a9
zdb0a99ab83e54d8062b348ebc8097169accddaa0c2ff192b224ed950ec922250585d1fee858518
z06c9a51f8e00accda230bf2140a0cda6aa712fb948b85b934dab9826fabc9816f6586e137eaa69
z5eac2623ccd21ef57155cb13625d3e56f7b635a5da610be6208daccfb290297b67e31a2dff014f
z2969845cb565dccf25668f6c72844e030a63d25d5628ccfb93dd1bccc8d2043ef294d358f2903d
z1f4625f7abaae1bf65aaccc6e94c438923109db1a8e0d6d9bc802f17a7bdea25eb48f210cb9b6a
zac405700feae3defbde6234222d59ee31320f6752880f108152296243d4ad0c98e9d710e10baf3
zeed9acbe650771146d53bf1a3f9f404a6e432b997a01b6b70718582df951ae6708c74d39b7f6b6
z97e9323a0de2eb01d230d63aa77c07aee9cfad027e770c29493a64ed5a92c09736ef171a467cc5
zfcf97fa3f7598da65c2647edbbd5a80cfa66df54a6a84debc740b871bd2f74b20d2513c41a956a
zf3b786a0651c48087633b2da1e6a21332ec293ba09d984a04d7e30f0ea279cd79555f8f8178261
z8fd3abdae1068cffecb9950abb7acdbaf3b84f8f1214db365adf01a17b02db9f02d0c382cbe198
z8975839cd434b2e1e276c50eca3b222e496e3936d31e0155b9a80b110e7129eb3d60a5871272f5
zd71fe4775ebce5d539b90a87b6bd78486d6d444021563a5398c92e879b73d683115db2b86d5f18
z6f7fde9c05802620a041302bcc8f783e2cf613b6f76d76e986dc559f3611bccae7c6dcd9244621
z6a9863d409286df17f1b09b1dae95738c25eae50d42362fb698061204bfd96062809481ad94423
zac8d2b9e86ebe8704c00ff255a8206ca22221b069cd0437dad5955bbe6a25ab8da4539d48c7afc
z066c179a3a703724f319bb2ff7c93e4bf1080b10d02d754cadc2de2e77ce59cd0ac183ac81ecbd
zbd44e76ed4ab6799fb31619b3fa9f3de35c8d4de6cde214207a7cc29e6837407af6d646ba7dc14
z712018a528803a321e4e6b7d877e1b2b53a217096ec977db4607530c165c8362364b7ab9bec770
z06eb59434b1ef60d28c08940b7e29ee5115bbc7e6629d66d9d469ef7770328ebb2d19b5fd4ca5f
zd9e0a96ba4d9d9458738022f4e1067e0dd1989d22b941d65bd09730333445f11d287fc28e0a3fd
zfd36002b54577351380837c186676da8e5dd49ca0ac8a9f6d7041bb7506dcf6b41c333f60bcef3
z1d40385ba0324fe66a5641be3f628803bedbad08f0e2c05a2b65d25617ce9161ad389296edbb56
z598c5d89248f95d1bac870d86a9a29c87fe45097a796f1b3347894f65d88c28f9ada959dddaf86
zf650d8db6a9167d87c889fdcac8e64a986fa4a923febe9919c2f0438156a2720f6979abd55a6b2
z83d94f3fc9fac4e387f59b916956d6a8a71a5f72d463a2d810c80ad138609ba51743e385ef28d7
z8353edd0ac7fd5228cacfcb74c293cdf109346c2dd4c6c0fd06809eefa6d55d995e5ea9d08ba2a
z9a626eddad90660244d29f2ea3d389a5f56b534628d7d2c17f5bd5916b994ae1509c225ba2bcc7
z0bd42263ef0ceb09a65ef08f7012643eb8df72ed761610fd13529e20c1705b293f3915676d2fa5
zff711a3e0637ef76c30fc82340f9bd8275ab60a6db56046cb85495aff8b9446e8beef69a5c9b9f
zbc1dd2cb4870cbd8410072590e51b771dc8a6e73d6b292beb492ee50b7bf348e4539f736aedd11
z0b4c814bb67e3def23f0c9fdcba962d5740000aec3a0b41ca725eedf41b0b3772e4e5f0e883a45
z45ec51138d6c4590ca8af90cf0470a2a49c1cad692ad37c984148e539ca24fd4469949b4cd05f8
z98520bceb9254b1f820a6411a6684bc5efead7aee35db2db1ebc9a8cb3dea76fa451f9d179aa9d
z320234a3cd5b7013b16e48b1e231217ceb939b5b9d4a9cc86f5b075ffbebe577dbae3d786c6603
ze35246e151428638fc65bc4f23dcf39b27cf0052dbec36bee149bb1a7df7823c5c0ae05ede1173
z7fb59b91d58618f3dea2bb567109d5ae87f206a12358e0b73c13a648ddd2b0e22a829f0057b124
zc1ee90796c313ffc8f21077c6dbdadcdb549f0c18c2406f8463204942096f620b26684729ebbd1
z746990423a606e83288f947a1409d52b95094de07c480fc50242d5f52baade3753982f2daa12e7
zfd4f688a59c00c2e32e0b665e7fbc8afa555add98381ea489623bbd3fdedc90248ca9695d83568
z917ddc314cfe5ed5f903dd9619f85265b658ee5857bf81d0659415b9d7854310203f869cd0d581
zd80124db66758c6ae5be3933d708831b104548987f187a7eb2514671bf3ab121b666486a5b46c3
z533cbd99871e07372557389a1a72131a281daaddb59eadd0ff9a04f26ca0d393f50755edee0e87
z85a4db492f74f64fc13a6b3df67386d4adb1513c7668195785a689866a33b555296e4423f12ee4
z276cbab97fe08bfb073656d74ccddeca4e7bf5b1ea6095c7fe3d3adfd42559162ed8fa3ea0c043
zf3788d2efd5a9865a2c42d80613cba9b373ac99dfba8af7345821e229ccaacf8d324fbbfa3b87a
zc1dbe9e8c016ed490648ebc77ea1f9cb4c8dc708aeac77e788232ad8bc423947611b606068f41f
z3dfc64c9352c4b9d360c0a598c880bf6706dd168f61b54494800a35b2074d42e55489d31614d86
zb88dd849f9715d311ca43d590d729be5bc45783870286236565cd75bf9502edf0d730893c90ebc
z62ccb70df3b340bf3e5a0814e18f34779839169fd55d06ff14793388e917bbc7780fadf794f9cb
zd3380b58e70fbc6ae5b471ed44c0e038843f52d3965f89bbe01aba3e7576637b17a520747e6436
z578e648b0a1cfe0b7a1765f4dec6cc7b24fe482106e6c6e11d9ed594d3c2f3cfd41c417b46b4c8
z439e31f6b12fc9863efe3dd0b1daf30e6e24b5c79209570cd000ecf5c7e3dbb79b3cdcc9510c24
z9bd4b818c73327e9487bbe943f1563e16c056a731ccc1d785877b08bbb31767fc73da1473d9f07
z7efec6cfc144d7eca51d4dee9f247b15402370d0594c5d7ce7e9f5fddf5d82e6a12f13c4a0f1ad
z15954cb8f3565291e958b7066e2cf03a484b677b69397293eb78193c63c766174ed43e0ff47379
zc520d321bf81d1778a493196fca91d6f200c5b9e0a2468162860046b35874bbd02f936638647c1
z8eefaa5881e3a44927cc106e15408833d42b12a4f464f97797b96a2534826392c21fffb05a4165
ze9cafc0c4ad4385be0b7ffd67b381e1e847c94b223917b9440b46a1fc1a21cfc02efa819f91f52
zfaf028041b195bf01f27f4a13dec1f91497c68332b1f99e5f8180ac4982fcfec01570d3c3a64b8
z998e89dd9368f18d5a83c9043fd80578342544ff16d7101c0927e5b2a9593818e1ca7fcdae9f22
zb645c7b9f6ca2891e2b699325f70a79ffb4e3b122a49b8e126dffe194dc87a39a78d7449112f74
z1cb1e9408e016d82200a2ca7d8d2f07e7cf05ac1e7b4eb64a1156b1e0247f17218b3ca7773fcc7
z12ecdf93d2591325a352e491122011fdf437cc91721d4ad02132fcde393b52364b589c853763bb
ze620e04507872e791c1742386165fd6c7d9057773aab03bd32af728acaaa71e5e6a0e91e0e737f
z885a61b6c12becafbf53b4467cacc3418597710095a6ec35cf8fa42bf8336af7c141e4a25848d4
z533455ed8f2433279a7c2bd44cd250963d3e57a91d0fcdb9d5dfe26dd58317f56acf8777fb02ca
z2aaba271e6bae3847c807c3f3e18d3d7612756dc5c43872279f9af82e168ae5b7844b529ed1e07
z5e42db4d47236540f0011a434d2a6cabd1babddebb0d8f04f451d96b1f5fa9e0b96c88f790fb87
zaed803f3008d8f27432a5b89f55f706e5a2eb2128a55c644b5f64dea26ac21b0581d488e6e1443
zab7a33a07e575c5829970794ebd99075ede975c992d604bff822eeba8cb3f5f934e6a7116aa0b8
zf464e8fe31b496977c7e411fc40d3ab9849f17da409e1b9e32991afa8e9d8848ab0162ad319f12
ze2f225e5dd3f970a9d037d05e25f8fb35e77beca72a9bfa78d1a39343c9e4f02efe61f1000fc81
z5c396fd4434b0beff21a64b0c930c2923aee1a1fe0697e11837863dc61a2b9034555ca268fe193
zd695ff4106cc72f96b862c8798dfdb3391a5d24dbfbcb3d9cce2b983aaf2286fbf103378da6a59
zcceeab77577200c8c2f558777553dea75adbd9e17aad51c822143abae124d22489556f70e38e9f
za27269c707c189e9796dace61de34dd1eed912b2ea3860a24b232c3002ce265439aefd53c3357b
zd9649a56272e4fdcb15d1ba024c462f9f686e6bdf0d2296d08cb366b38a640b50af9d13fde8c62
zee831e7835f5f426f4a8c7e7d0b1448354dc2b797a961b6198b57595ff512e9e698bb7fb06aa78
z6dff4ca5d27c153a346fca56581263f6813963281caa41edc11e4b99944606ba7bafb6730dc81a
z8805f019f83886baf7dff9b7cbf9bd253f1c3623822eccd1fa6d76b8ef579d28360c6a2710ae3b
z0379ef68f980f00ee6b9457596785650aa4ae3c4ca0566c139ad7e9748c48833daf22082e3620b
zdafe45e7ab6bd561ca2f8c0872554866f86e1630831fcdc0a39a5bd52659864b654682da96924f
z855a4933233d2c81083d46d9868c35b96e623291f94b17ae6c0bc14936993cfbda29e4b2f9f164
z677208b0dd5b076c97b4e7eaea1c03d7fab703eb3651726e9f89d25098398b3b998ab18aac389b
z36206132d91dcdf10783e90576f667523296b40a24c0654002497b3f96ae04da850c41de55c5bb
zc8dab91cf0309fa1ed0deb0a9c08579fd95e5526e8fee0a0df4b08dffcddc5311e1f35a40f389b
zd506b8c211912c34200237f0316039edc91e52ff7087fdee45569adf78a15eac15b9570b01888a
z1bbd59557192ce7406a27e494427617e5a5d081da5f7a357dc9b47446be6a611bbc4c8f9dc5d63
z113d28eb886b35a131d2245b0bf4b1c691f7e13446007a02f0d63c7384ba3d3efbb4a140a56f75
z69a6b4f4746e486989cef32bb7801b31a37477bc469d156c244dd3f2cb5a9c336190e3c56c1a59
z33c6c59d6b238092b8d84e60957a53545957f9cc6789ef538998871b833b9cbae5a00c4d191bb8
z2f8bab54e1e8a22ba4841a9d16d88d6119893599390a556b67e9aa70797a19a61fc42deee905de
z29e1b1746cb9f8bd38c8b24b613843d7d08ba592b036f62ff923c6e5805b75b95c9b87386c320f
zdb587fb3854e07dd4fd733db745d664df456da93920ee62cfcafd11aad2d4af36bf5c94a0826b2
zc2d56a66eae766e6b923f60737cd60e529cf2c33403dba15136aeb1c745a8473f6f3b9e2eb1028
ze2fcc47029a85a95b390208dd1b2c856fb561a9bbe0604b61d01a9436b479ca3f432ffde777930
za877a3632b42327e693743ab8042ad64800739f2b0df7d6aeedf4f4dad9cb1382eaf37f3010cc7
zbff0fbaf5bd3e333fd85f0c9fbf4f5b43a4ef4fed7ed2f0cb059ea2ea607b28dbbbb7e8f96603c
z1bab8bfc70f55621890dbbe099c8c9fa32f95152e6413f5f3c07cd65c6bb81361ed100e5435b48
zf0c12ec116422ac49c95ca2e72b431f190d49eba09cc562750ddb04f6914ba0448ddd3b4bd288b
za1cc0d6a835dc30ccd9b6fd15cba2cd0246147e4bcbbd31a6b4f8b106f9e855f3f2b91b629f099
zf8ae844af0fef892db9aeb615559cdc3b8c4819270ba30476dfd064e9ce2186423859e5b495461
z659d69636791910a1aeb4e27cb6c38ba584024c1b745237613a59aa23821207d4ba577552aa81a
za75358cea23fde003ca9e45898ff120bfd92d1d062504e67709e98f6ca22cdecae589ceec55ad6
zc06c43f367aed98a8375533c16793332688e68410caba65c8d7d03f37ed2954bd35f26aaa2b8ee
z82e48b8e772a911161cca02960615337a65ada79c978cb01a6ec371c0b7fc0b883786f1a72646d
z0198cc740a20aa6c89b951469efea3042fdef584d8930ea37b04a5859259d4f0e13ee6d2218771
z33b44fd730ada26c1967e06b95a7f3a21e6f58fb99743327eae9a6b7e99fefd30f2da76c16d72e
z310f104ba2f1cd47a38392c6b4be0f89fceed59edf71586ac8deff1d5962740edbd60223fc6983
z5f0257c99a74adccdb51c0d863656379a9434c7aa8d27fc83a7fb5d6d43179bd676b388b612ca6
z2475b396cf785b9a51d62cbdaed9cdd8c7acc9dbd298a7f3f3b9edb2968652201be5a0a251c2fe
zdc0a0d348dcf8caec8a45bd8eefa47110342cfdf2a9e7f4320344dc9c4d017daead077ee2e882e
zd72105437313a0c4508443a3962e5428c5eafd5d8b43db4efad581be7019597b7dcaecfa1f0383
z0c5dbf866c67317ae940b9229115f3e195d993439f76a8a996b5df2fcb2a481594e2c5e531c4c8
z09bca81a47b5214145776a54e8b25de76a0bf46d2bd76d6770a7e6250bfb928a525ebe3d47e7aa
z2439b01e3da68de87f6af433a23cd5479c333b3185d6d594c26d9376b1d233f280d51c3245e4d2
zcab5ba933106f245660d9510afba26d961046e822fa85a766bc63e55db008d0e4a8d4f018aaef2
zf7c1bb6c9799557420d4c310f7eb32c224b417baae4f4ac39cc7a45eda5e5089db7d9c2419f706
zabca460904575dc9c87465e99a90d239e2e849a8e82f8502425130fc30a07dad7df37660a0539d
z745fce83ceb03a8ef0775fc3a59a288ece60037db38317ef1a31541e4c5b1ef542a4655dd1fc0b
z5457575e44156ee3a4425495cab155a27e10a41a87c4a1e2e981e6ec7f9634bd483a83e241aa1e
z697fe19ee1998720a4c27e56b44edf8aefe0a0a8a65d8b7bcde10fb90b8366a9054aa34c02c550
z475723355164315e0dd3f1dec8f883462ba647d1ce1b067323468615a9945ca3a2418afb8d7415
z316f172a578eadb81ec8645e9528ab166e8b0c676232c9fdf079c92d94898dbe53879ff1f07e7e
z26c2cd95272f83e0b5ead06726185b25c96315af565259b4c09509171dae97e9a5619dbb228329
z14e5f5dff55041d500199b2e8beca0a2e14f7b1e4a126ff2d786ee14eb570b484c3874c324c45d
z8b7d0b9ecc08efcfe0d88e5a581a81c6e67a73c528122ae3a70ab9f5e0e46704a9f75deb08a637
z1e4fcacbed6d160331903c1dc3abf743111a6d2038b9f6c8a775198311bf884d83e8c32ebf87af
z2f6b4cf27b0d0f3c87e0fbe62867f3be31709f1d61fb03f9d729a9c8a5d75d751da45208bb4373
z66ce4bc6c98ecf58e0ee98cc8e709b93b934f2779dc6da9f7638b088ea1f5c36eac432435e0481
zcbfe4c7f12d457a9636f2adc7a4d1ea9db4659e82b9c0a6253be06108f23ce0578445cb5eccba1
z03c8075f8ea2b72fe9b51afaad3001e3bb742f7b6c7e067c95dc69f0f810bddf94f6aee94fb867
z4755692eeef544b59d57c86f7e9d13e1b0faa634d98776ff9830c18c96bffb610245222ab04128
z8471d05ffa04b50ba4d1c99e3994a35ffdb8fe6967a2aa7736b3b0b768c25be75926a8ba859b7f
z477ff50285f08a877757efd738dfcc40cf7c1c8d00d363ec2b0d8946e4b3a9ff055aa2bcfffde7
zcf266ceeffa29faf189aa1dd023577884c5a8dccf8a11d3eec6a3b1c7743f3d3e3bcfe3aa5c629
z2a09330a0015c54c3edc084d95364e6ec181baa6dbad7812d7a17fe8177d2e675a1d6c0361a080
z235d59e26c4a0b06e5288dc1561ec79973de2fe2683ca688c0b1121f4aa2ccd5ce45b0b78e0b73
z85604aac0c13e2f189303763376b847248cdc3ece15a12c36689c2eb29ea092b0b176e0beae381
za3aae14ee16c825fcfd6dc82cf4aeed02e5b4fb00c5cfa3c705eb22cbd1fc8e2633eea8f2a8211
zed0c064df3f8ea6e4cb2bf9489e0221874921be7e6234abf851e32eb738a545fe68a54dbf5124d
z69aff05a23ba71e22e50e711ac1bcf3804a62c533aae319d2c32eedb006f269c2044045809f4d6
zd5ca671729b8af8b6f9e0f8f56f3943a1cf659489121bae016a2bb2c637b81c9f776a706f3ad36
z28c5ded16d590119b46963f90187b347efee4821a387435562cd59fe54287691d02bc4aa8df5a2
z4c25525d0d92dd0787654a270d08e8f7ba09fe896ddccf27b0ebf7c2227cc06be93e246e030d4a
z2077b8e3b9f5765781b7d01d6be0e2fd9e4eec91298bd60c219e8802aa1b76792189d487e0eacb
z6b1c5b4255f4820ddee78de0bb162a42e0e2b1abcd1438fad4593dbdde2b6b500738fd53e9f0d1
zd4e9dd2caaac562be02721600145d7c7c3c0d9bfb5861814484dbe6d50bc9a009ede46e4e9b368
z6852dbf08a9e23fb8a0bbdb22f50f83e546c50d89e3082335fba8d3dac384be8ff750a19b03947
z8221884ead5f826a8090c00b9bfb28f052c695b9054151af5e889f427ba8b973d993f4f30bb074
z94fb42be4072ea6879796aaea4ecf6f81c1b7b5d7eb6c8df21b4174d4bc4c31e5cc099fd694665
z7f439b529d1c634c7cf14b04bfaba2c9f065c145d2b87336d17dd47fcc65f493c2fe0fc07e5cb8
z1e93271bd12502f6d00bde59c481d213b708fc7ea9b3a4d68773a4d66162eb28f5a85424f20e89
z2fdad004dc40830813ee831424e45c949402c1aad6e16441f89712957c82a5e95b24e68e563504
z8531e1e88ade40c6d5dae3e5d5434e0c384e4ba73077619679ce01246bf7de06afae5f2eb482d0
z7a3e0e6eadbb6429b18d98af5fa217736656e35fe597b50506d3ba5e63c24e76bd7d4f92dc88da
z433fb161cd1189395d194e31146f116da0f14a2a934b86d11adf990b41b5fa613c893cda736ce7
z63ed61648897f7bf926cb5156b946bd6c0b2dae49883d61db61e3a6e7f437eb042e9ccc092f2e9
z1ed2542cd5e4a5ad0247a9d8b02f1c53de266e48034247e558317174ad3fd9493cc42840ec5b93
z336006b9071e92940a0ed628c6a703009ca5dfd24d9134f283e8108f1be4c236b5ff7085b50d57
zadc4eb2a5263658ef4258d9f2c0f717232e7dcd854a580a87ec04b60074b3b7c2636495fbe0d0d
z02686449b6519584d010079e6e319fce1539694da5310bf4c265669b794cfd258af5d296e79b93
zd7479910037d34e5b6cf313a887b61c3399830dd8eca3ff6f1fa5850cbc2b06176255a02a8c475
z3a6732b4c7c3b1e2d3326b1496f33513d32dbc905563fa410f125a1bf78609ee5470c6d9c430d8
z45a0a21265171725507abd691d32b4db4667c25c1107f566b23b284a35a6836981656d8f959b09
zbd3894f6a97ba454d6eb89b549b70897204375d841a0fcfba669510deb031594dec546f0a16ed5
z6e40ffb8caf8653a1418886782cec6ac5d870845b77cc58612a7641852b6542fa5d7a6aa84d4c0
z58eb3ade463dfd4cb326e05d6d9a8d4939a8f7e2651f775c13362b59cabf09c01b5bce83dab572
zab67e5a8306eba9a7eb2c96d3f67e1cfb9028b47765ebe21d0e5b9025945602505cce71eda8ed0
zfbc2b5a66aa1f8db068d25b8b4cc7ce248e5dce714388776b04178bdcbdc1ff8d8557c5c5c3455
z0ae2f7436f2d16a0c1992a99af190572a07337130a7c110ce5c9d3be2713831fc7355d6d7ecc87
zcd5bb4be84696eb0c4d351081d3c37860fd22547d549e9f4feecd04603b7c4d0125ca7a65a165b
ze232104cac48fcaf1561171f4eacd4e67c984ad992fd13afbdcd2016c5f30dfdba97b4da0355db
zba7463b081fd93e0cb4b42f6a21ef15d0d8669ec37b83f28d0e040ae27bbdb3a0afbefc0949dee
zb8196973f34b513055d5f2697aa39a8e86b885881abf631e6198db24bbdab40661f559a5893ae0
zc24bf9a2a0438bb1e7a77aaf84f53f0ae216961fa5e08492bb25a890511f2ed63c80055d00ac98
z232b278acc3f32b09b1bca43ca04ae10a9eee12ae799c679e8069cf3b15305fe9f8adea87cf2c9
z8e478d270b54a32f163bbeb7b3eff023bf0121088ee355bc5a99bd80fad6b59fff14e3fcff1f50
z4f7395e28ef9613a3d78516394cc72baa1e4ed825369017ce9346b2481d1b02c236163f4f79345
z90d4bcdd65ae8834477a23da95383390574e3f123c59848c9c614f775dcc422ff5367495b87785
zc0f208828ff14a42bb2a7fa1497e0c897cfca9b1cac52d0c70e4b7227e692ea06630fe80513c55
z3be2a06138e20c88e6fca9d8247da78ae3840b4db0293860e0f719df68664cc25312f00134d818
z280f0c500b6883efd2d3742a717788ec22fa849ba3035ab966bfefed37922d351e4f490512e764
z08e9de31d48edf0b79c194a7fe5a05fb02e10926426534df5daea4b9249b2f08d828cc0e0a103e
z9cb07f575d366c5550c38fc187a1b77641d6d7254072ece9223b00ec28ea2ab3c64e40795f622e
z75c95b6c741d07c3d7990f22a549e35be19b2608471875bd68a2887c350c9aaa3589803690cfa7
z5ab673a9f526b3f9d99fa25d7209f9a93ccdeda2a21c0c35f16ad9dbbc46512d45eaf475d049c6
zb0e5244b6391a9014827dbd33b03786d64f52dd46f972f9dce902149e54518d94b60387f510250
z136d5298db1f495be410f2f4d24292a0d15571dd7a716b29e5cc29d0e31f2b8ed4edfa0979d198
z2d5e8c2c75611e843d136538436778ca525e0d35c52c8d68c0f8da9bd85476d4cceafbd1ec070d
z55d443f702dfb30eb68262bf0025c1392af8035d9797460abe0bd7b43726722264f41d1b763f8b
z6647af8dc344626d3184811a36c6553264233efdf5f86fec9b9fcbd16401b38f52f51ca54d1593
za46c2d4794fd0658abaa4a67132862bf4ff183de1bd1b801fe341bf7228af2b9047696161a09a1
z62afd867a982226a273f8593fa5fff3d3bfd0faa735eb8603c89bf06f2da95167a41804e2b6aff
z4101e88681f85f21599866c603c641883cf5e71adfee65f69b705fc8285164147a7a6372ccb473
zaa2c3066ff7f542168f82cc4d1b73ea18dcfcf5381d3128cd4857e10c7a96499c50b296fca2c9f
zaa7933f46835e1ba6bc90f600d0c4b7158f5afc837554b371d0952cdc693c1c7a1a3762024eb46
z203a4e4f626658f17f45418f96d711edef2eb3bd80943b5bc7b1556a61e52c2b5f4b6932006f7c
zfd200c7556a5711c66cd0d484a4a1bb7df3e3ddbbfa485a4a0d2867f46bc83d8920f196af802c1
z30fc139fcbb455fbbf6da739f323bad3a7d373a64c3471c88457e525448348fa66e9ffc85fd002
zff91943c5053b14f929250df0ca9731ea19e498145eecdc6d370acf793276d5f3ba8f5252f1678
zd1ef6193085688ef914fe4cbafa6a0f190fbe6c431072c0ca0162f9a4719db16fe7d92004fe200
z44a4258a8bc46186b7f142c98ba7e7f888b02fa51c536a09627a4f0188a19009ab927fdb853acc
z66be17da2c4017bd9ca4ae6822d5def349248c656d6da07f3b8b6caa0ed8331b25f21248c33f7f
z9dc8920ca3de82848e59ba9172e9dcca48a3434567423305f9217620b9580372b99e7398dbf3ac
za519adf93ccd6a33ec6ba8a5c504fb98cab3eae055e93bf446dcb9eeaf487067306bca269b95c4
za2302480ec356d92ce80cbbe4fe9d13bbe98613c9355b0b4b65d32398a9d99521e972696768a55
z3567d27a0b120477f69b0d2a16f96bce5468e2b86805c25a8d99ad997e1295d954263aa7cbab5c
z21b8edd84f3b51ffcf817b7b2f994d236efedd60b41b0ffa66c65ab99ea7faf0afed33bfba83ce
z9c63f6e529984d91c16eae1566f64c12bbc924a06ef5ea6aae8a9f1e674428a4856b02b80c9005
z6a65a7833e7fffdfc30982cb9fa83d201d55c955d58080f799e09060dd8633416cbc3c606b90a5
z9bc610bf79d23f34bfcfb1683d9da00ccff3fa3b475b82d5c1120caf618fe661d76c8befc99803
z135abb0458628d3b365b0ad5cf7bb7645c8ff7a8adc54bb3f007d1e1553117df9a8f7505ed76b7
z0a2afce3109a09afda75336d8769f1b60191b7d508717e7c628668a245bcda8cd3b6f3597ebfee
zc185bc979774ce8bc5fb98c87409e2ca4812903f524998bfe91a25c22e2de5897db1a07072e477
zea8fd0a3139bb418b1b24897a14437bf0fc94f4d2f7921cbc22bfca79d252eb1ad7438221ffcda
z44ce3cafb4c8b3648b9fc80dae5472df4b20378497d0f760be00d60d9cfc4b62578c29e6d7b68c
za32ce0ab11eb2763c9d6b13bb8259cac468eb5df6d5cd1748b371329c164217c696c7a764446bc
ze43c600203801bd80ff24951eb252bf5b7faaf62d5e7947f392f346176eb53b023ac24382e6462
z19b585841a2f477867c7558f5f9a441ec86105bc230dd79b369caf2f4d13679177545118f9b987
z69e48b7c454b05c441ed6a31da27b1aafca4684e6ba564424aafd28f9eba8ecc06c39d82765487
zb199d74ff5ebfc75b00c2d911b1c20d34450881c167759fd1942cdd35cf8f28ef814d184b2eabc
z827398e6b8a5c71846ce46475316500c8ee75fea8d4dc242ea8d5b659975bbaac9e3bdbdf600ae
zf3b6ce950d86823e983d484e19ee14fbe92f951f5626e36dd810683443e7e16d3082ea9ec27944
z66a272679ea020f6fc8695d0695a837602031b8b0fa1914a76f478207066fcd64060ae4015fbd3
zd428234c4d500739b398c9909ed85d6d8e1509f742553d7549268e3d7ad3a686f2031e30855759
zeb9baadf24dc8b268544ac86542e5ad44904a7db59ce7b5e8503f92a685a585c6884270b81dd9b
z8e1a7f0d51eda32ace090a74877e22da0db3d30e462ff49e9ad955ef643e980038aab05862b9bf
z7d62bb41b03fbc4527627e4b8c3e0b52de6c1c632d02f3d5427f492ea4a14ae7d447817f6edd5a
z86a643614dd34f722d530ecedaff887f21fbd1125c2cb8421efd30581ab6c63f40dcbce13b0116
zed4df65e7cf8d2b3d8adc0cc948b1da0bb34c9d0df34dc969c88a9f570cf107ab2ffbb477f44c6
zb04c5dab226ea8c65ff8712ccf994b45a3da140089a049dff0117ca7fd8b0858f5adfcc865057a
z6930a799261bd74ddaf5b69d40d8cbf70e8ae5b48c25fefaf0d25892aff9eb9b29c0f890020b28
z8c65b3c8b811f17d838f248a6aef15b77bd1c18bb0876e90a0be5eae2a561a57f176bea720f826
zed48bccdcda408030df70fa90f28aafb2247fec2445adc109a5f7d63d1bbeeed30deec6d0def58
z76f9a7ca009f8633ecee3df378f0900b02ab9322ab8348b2c52e7abf7f325c2ffd0a81fd7ac970
z25134eb19bd45945ce7bf24b5c809fab09de3ee45a9215af7e48847736de55b55aa228be3ddcaa
z48c88478cd5c49f3f79e117a6dd0ee67d5cea4420a47dab38e9216392b4333ca688d16564d3a63
z909898b60f9202ef936f982b21056b680c0b8d893cecaf851b386f55447cd44e6d9c98b3d5082e
z028942845dbb9c2edc2858290b81da04f91cc297fa146a696dd777d00083fa6ecd81e919b81bca
zb573ea34c9156fb1e1dfc965b39398c48f2c725a253e0d2d6538b098e0d1369e593980ce1629fe
zb732c4578879304eadf74ef31065c75c15a8ef592970a9ba9a97495014b364d6d5a9510c23d297
z04b250991a150948c22b49f8e2d157003cb27ea6c45620635ae46e686aad383bae0d34f020e601
z7ec1628bf2607177f1d90240065fcc692447d2040e7d35c0767b227a5d41dd2a59a88220580a8e
z079addf2312f727d775449cb412189f4079a2817537af8c41b544e2c3f4365bb221430e655d159
z66aa381ed3a0a8770c80fae33ccc16d125517ee7d841b7822d1f9094a12d84fe8454e42065710a
zf398181eff682a7c2f5c059572bf315eda041b1976ed6d8693fa450fff4dfe86cd6b14a445f37b
za9f2a91be2fa178189ae93b48d9a01cd25356f6925cc5e93e10b404804a359a811f3963195cb97
z3407ec2be35cf8f0b2e8d26f8588e3392284fa3c28781514e0e5ea413d969a120afa3159cf05be
zcef76ae1800bcf0c623aabb785ae42aa91a5eb25e5ea9cdd3db6b78b79f0cc3e330f01c87eea3a
z0a3ac98d9c56715aa0f10dc66c102596aa5268e6054a6254734a0dd7f7f74533e8025eeb20a833
z07a2001254ae72ccc7f0f028efee2c169d8974583a49bda583a67c769496a5082434a3021e0caa
z2957d59ebf62b55e889e28d8ea67e9d03ed71d70f5880dc01a9a66acdcbbda4e05b4e3f221773c
z7bcfff83286ab65d4adcc66bb83d486873ce9dfcfe57da4ef5c9e306735261060f514cd807302b
z1635811fcb918cf81b17d4617d525cf98821e10fee1979126129f27da0c83d0167af3819444cad
zd9b6a90da5670417c61ffe51516a3d5578fe69c7aa8f1db2e2b25b798573e088dc5590b744d76f
z16f3c354d00f152fd41a46bec33322fc55f1d7548dd0cffdc9205d26821ff3ae9ad14478410936
z2ae2b296d6e340b9d575416cfdcd7beb9b2f7cde3d08466e0496c18e3ce6c8ff8e0ae6c9cd414f
z337b07a8dba7eece3a4070b8511c5a328c422caf8d451adce618293b297c503f4746f66b5fc05a
z1abc69686912716dedc160b5eafd3f12c59ae4dee489cf9c6dcf95ada1bf6537875ba70b69a519
zfb4f04b85632ed9d6d0da7773394db4b5333867d982abd158f6e70e280b5b5c51870fb8a7addf5
z9b839b1a696d401047556eaef66e00b3a989344d65092cd2048b74588b4c99fc94abc5d39f4bc4
z58adaaf0c847724ea71fe3c82c50ebd47c498996e2c7cf5edaeb755b72705b2c13787bb2eb67ea
zd9438c69097d7e7e429f758a9126a6517bb4b18b5fbdc5224a516c91ab96cf1f77b7c074699b42
zadef903572273a72b30725c0b74d19eb88ecd4e5ba73d3ca495f2be537d25c28c605876ee41920
z78d126ee477db787f77c747d9a5a76a57124ef733971e523b5ae1a9eacb4bf89307fec9d775d8a
zda53d5352939f768322866e63b6b8d61fdbc7433313d0797e267f0b6653a464e0cbbe9eb2af7af
z088e406f17bc3194d58eae6595e9bd9f88a6b154c4c9e1e6d758a7549fd34429d08abd06b2f808
z9e7da741c3c987fe16f2b4be8ba13ac870e56e1269aefccd2d706d73f06d33e11ddf075b3213e0
z84b3acf99d0099b99f9e8d3c4ebc7cc8ff3424e318a51f5030dd1a7084171c8cc2d9265534eb8a
zabf42bf9a38951ca7078514d04b29814474b609b78b4d3dd3ed4be20b41ed45ab99f335099067a
zb0b4b369336bb9f3b5a680fe2e64437d3797d5ea447707d5169f56c78fa152dd2bff24ae199d4a
z0aa196f81dd2c198d01945201118d7136b3fbe312930b9fcb8871d41bdf2541236bc868c61d09d
z5c0de6f2cefb6bef66f3fbf91c59e16f2b61dc4553f843341861c6ce4950ec10e05da01dc049a3
zd0ba57ea292e6752e4d67c721bbd35b3bcaafe8b57d71a8f49e31de1d278252c535b3935a70f52
zbf6cc3cebc28e286ac2bc3a0521f6868c28e1f03bac3328c0ac6268653b25e1a1ff471b6ead7e7
zdf9a311e17deb9410ba7fd4df55653824cc60c4a68aa09ecfd8db6f33bc6f8b5e1bef6729a04a7
z5e02357a803c8e69f72ba673390a8590cf9b092ea54b976765cd24c2b1b9f4d5eb68d62d5e7f94
z0e8c5fd9eda9524091d070caeaaad6500bb9391a75558f226ed0d6aae1b1c8f5c5f7994871c6dd
zebd5cc49ac23f21290927d20ececfb12639d831465ccc87529432f7daf729ee06320055d142259
z6e8e585ce9786e871fad5169f19f343a2302a851c1fc4592a0dc4a3bb7f5e773474e499ea93276
z97be3d44a370ad19aa68809a2c5c7fd8b977348907a821a70da1c223331ba5162f53e7fd250e4e
z4b0172928bfa8072848b53e4adb2641a7a73e3e758908bf6ff3421ef01a155912258760fce5c58
z502980748bf474abfc84cef383b829db1d44ec58e0a858888eed717ca5115ff8a522963c16dc6a
z4e8d70c9f9bca210d5eeb63f2518e6504ac118c86365b5599c89f2ddab0ebf2fa3bd2cc38dfc5a
z930dc0a5e91dc8582420e7658aec59405b0594998c0d19a4eafb2111c8b5ec2478772dbf5a2ade
zfc44f04490775e47404358bfd367ae647b14707ee158604c99b80478f67dc099f70ba67e2b6a23
zdbb38a09aa279efee9e8aca582b75422cca72251f3b4788de03833b5044f7a674774813997d2ae
z3daec42bc0a696d53b98cc09cdf4c04b78845cd771dca3d4e988bdad2a7fd3632c1229e074a668
za6485b7ada5168f6225a90f38b5bd3552405030d932b73f1415ad196db1fd54f0163f1295e5e17
z8ddc9a0757a1e9b6ccdbd62adde1064190320cb5d1a88063402d66b8c5116151c09e9a59748a3a
z5df4cc888420258a7a6947d122a09d6c54e93da54ebed12fbde572c8e02ffcdb55937ee23c3195
z4181a101d9ec908d08ab9db3069e9e28dba6a38b21ee3f40932a0a9c6f519c682460160f77543c
z1544c847f17ab9037cdf6b4546308811d19f3e7959f130aef9b15aa59e38048fec62b04b16404a
z85e884141ef6b94c67e6c5957103bbded287e15fba5d23cefc2b402cafac8de54f089d932f0a8b
z845010692c5e8658e2ef4e169df1797881d7216a165da402c5067b3a9335e329e8e36a796498bf
z8fa957ef9d362dd0b60368dba5ffb79e536a58dcd35104671a7811331256c5740189d06a02d3a8
z4c2555c1afa15b75b62b63e9c66c42b52ad3ec947fc172241b2e37852d52419275606fd0cd8720
zb86235e1e8f758fcfde6e6e103eed0e706327b7018b95084b236261df2f6e708cea5ca4b353d33
z1e01035bbc2f83840899b0ea3730c242cdccd7c9d6e25e74889fb2b75595cb1ca3c85570daeab7
z9f176baefea81f23bac06396f6195403a7d9ebdb6da125e054d76af8ef1cc17d2a3921037478dd
z9a94302d26a917c1e8a17b4514f1a9a1a703120f87950edc4e7f5c7ae9354fe2cf7bae6b33dcf2
z35788b33ed6b6a3b1b76d786805fa4732a9205f38cb283d3d7d881c22f131da1f48ad68730c7e2
z6e7ea9c384f406aba6137fce413c9104303950a6f8853a13fdfb906e70e0e28ee8f0ee0ce3b6b3
z55d94a6eda87e36b0af511038c3edb90dd90587191e788f4870d9ade57c91a5e50b849d070e02f
z08b947f0946ddc7855963e984b3ca4f68e110109676eac80bd897e64fcb270d1ecdd6a47474939
z7aa1aff1c10fe1266d19c9772e39d9b8fff7ae0189bbbba0db35e832d9d7d22ac95284d7b436ee
z1095aa1fc247afb87d14d10c887625cbb64071310642c93b75aaaff5f3393844b4640d723842c2
z9f34521a0b823c5dde22be2c124b40ebc177c5162f6cc1a5305da7706f0123ec9bce2ac56586d6
zb9ce03e79c0784d063f6bd4059f6a1520a6bf4c2c0dafe4d890a233c67a294504d53f105c6629c
z2d09bf428796c54a8c6ce0de168144bd9e6f584de659ca77efded24b60307ed436c3f6668bc78c
zbfef96417b4a4a33a6c999b41407376b6e5b8cb006026c33c8fb7036ea0b60154c62b35e10210b
z4fff0b41d26aaa1624c1ad4d7b6d45554dd3487d77b8c8bdc41a165710a5bf05f01b577a0e8f90
z102332e77178d6fc766f793f082515d0c645fc257b4f680c2036869dcba2b01ec893a1369bf4a1
z83ca137f27bc389cd0b444b2ab0cdc081fd3a1629e2dd4b8715675ae4be0eeadf1b010710c2be2
z7feee477d3348772d8e15df74276d84df1d1eb327e917ba1e6504f747ccdb05f748d5721620655
z1505e90bb34358dbaf8e90ded84457899dd3ca193555ac507ffe0d3bc4f6a113033c2db69d6d9f
z91367ff7b5cf3f5c9f155fdee77af9cd1335c52a4675b66c5f989868c0125079354aa27b8fbadb
z6576a71b4badd0b59b14dfb4a340efdfdfd5d48af3bb426fb559589d80693baf28f371ae3f05f7
z4ce0e882149545a7331e4ee2dbe8b7567610ef4e8428ae86da00c9c47e5522f795fe1ce2682a5d
z8d3c8b9541760a5bee1ba9059b198c1f121585563f65374fbd90b583f4a7ba8af5a7058e8046fe
ze906c145ac6f17e4c21f39d5f9fc4d4622cd05c03c6106b83606825e5795c465a206a7877ea804
z97af7b315252d37d1ff419f733089cfafa582678a13726e68b83608286c5cf8ef71ad0e8e1ef2c
z454a9842eb00eb5c575118ff2f8de470d129d8a6da18cb5585279a5118241f7dde73133d638f2e
z36ac920fbfb5ad69784643fc2b07c116a743582ea1c6fd3370674384f7d5765b54ae9ab1e3d86f
z1c6e8626651f67960b09274d5e366cd3168af408ee7d5f1558e1e8d4e777e9030e840adeee3346
zc8d854279b48994c810923c8d7f236f1795f1105d8c0b477655400802d226ba28a115ee869c790
zc232cf93c5d4b67fe9f46469a042af7ceac1e7ff1ba3c9e137a31d080067411f0e504ca87145d9
zbe79c0d3a1e9b79e2cfaa12e2ba13658ed9b87f85162de3bc7c23f57b323b92dc5e20e8211352d
z6cebdd0c5fec7464b4f0a5e67830bb8449588768cf32163065f0c0d8ce9b245ab3679aa950198b
z9f9ea938bd1d4968b3b8abaec06b5ead1aaf017cf679d09d4b498134054648b96c341268e6d22a
zcfa546701482f9aff2905dca4baa02b663ea186b07b250bc1c1603c19246f54127983d29782ef2
z647ba7cd74b9ed8fff31f730846de03d2110b8803d0cc63b57aa647742ced6a6643db2c39c739c
z0f2335f689d03402f5ea600dd64b48a164e92ed5bb260d40ff7007c7cd6b912b8ab271f6e5242a
z8633a58e5e5ea22d52d0876bd1b913e88ef9b3374288e927ea6df7c9f2ab4c523572b603576585
z0b0130142bafa275c30ef27bf49a27ff6049ebb77d6114686b49bf1457ff8f9ca81c5f9bbe19a2
zcdc237d450401b4e67a2e688178b8a90f45bb2b95d9ae17c7a65d220023333fb30b4d31e5484be
zd65491224f0f43a83d9c9eeb8e79fbad6664cba74efb60e39bb8585f48fc203da63aa5a571b485
z683f545cc0205c2b26cb0293e8c47e7a109afe4aa94278c96160deefff865405934ab92a60214e
zc88fe89d6904341cb54a1f66b277c15a0acae1e5a5ec5094596997c78a4ef9cb089f02b808b53c
zbdd0f2c55d414a2b6f90bc615411d07a56ce70489291e9ac9176aa71b061ab77ab40c890196a10
z465941eef415b9db093d7585c41c3af3ed4a86a44fa2da1bf59b03e11649b26f70308139223dae
z239753116438a2408b53fd41ae792dd3f558491464ece53d7cf5ec9eaa83451b46d1aee3185be8
zf49e579ea34528ab54522f563dd711e6e5e43f914b5ab30ea3cfa3529cf1a8d93fc9a6c1962cf9
ze96475a6e4fc1ed58e7099f9df3b48121ac14410b0560cd81576b493cb63a338a74a9f4bd68f77
z0caea11d63667193482fdada977536a600f5949e1980318cf8a3d03337277346108328ff5751bf
z8bda1cf8ebf902905aa92661c2fe6c88550f3cc731f7af5486cfc76064136d6e6de4772ca12e0d
z0047a1d0ef159b0c3c9e09dae6e007588ff35de24ad9936ffa2c7cec73b0106f0730856c226915
ze4324944630def9f9633a3b5ae6020e6fd5be2998115a7d5497fff7566cb602ede08fd56036858
ze779eff06c3be020b9bb8bc7f026fccb627a777be6a0937f4ccf19250763429f106882214616d6
z249f963bd32556570a11776b59f49cf17bb4a3e4f1c22c65930424c39b0884cf3d7374a0f005b2
zc4f4866366d1da61a5cf191e4c1e7f09591effa12c7d82f40e5499136e3a1a1f071a6a985c67f4
z44fa6bf97bda0345b8f389b08bb0e3964d58db66f217818d41898a931649cc3b783d4df9877043
zcd26b98aad0ca30577471c572f67d2b3fee030cd5ee89ad02bf890117a6cea3637e2896b94c0a8
z496a67a604ca8e1f87535193e5e0cf75368434c1537502fb13a1a07de3d1bb3ce35e0f12f8eb3e
z07bc3ecee3c0a231ace76ef6e3451c596d9e6facd3606d20b1af3fa1ab0696adf14af1a6e32cab
z168a1f1c3d8de5c6eb19201598eefb12188125f1defc47aff4f04c36c21a72df1a54bbd510df15
zd258f544974ae1781a7dab5b4b74c7b2740489ddd6150167fb75b5571b2c04f8186626742e5a2b
z45a1e3a9bc678acea885573d771fd08581792177d82d5f62aa2718d972a81fdc50640852676b15
ze9976cdda7d1cfbd21394acad9e1b10d313da13595b160b03864637f8024f1b8727ef0063eb678
zed58dd0ebf2b81d050c2af0cdcf011a147210be81c05d2d251c410fdb3386e80fc5f58682fb598
zc8ed2967d8c89156c70e8e8b2d1802e985152d7dfc9ef50a5dd2a79be13b554565acb4b0a95ffd
z1b83c3f3826cf0696be6d14790b78e3c2cc7397a7e00b44d50ac85256b278a641954d2d64d8801
zf9b46bbbc6230e52cb91b895a1b3a7a59ab47305a9c602fe84c88fe348de3854ba896e1d6e360f
z913c7ff7bc451168ab106758417080329e4e43a4cb2d5041afe535da6e2787d1edb54cbc77558c
z04a3702207a0f85bc5895cf2fbac6b8fd4749e0281552cda363b02518afcb19e725d64f00778d0
z3f74485d8e9f2af5563845d842a77e07e082cf8e399c429bdbf2627a91ff6ab430d5348157d27b
zd130c7647c10b0bcaefed821ff5bbacbec90a212a82afc8f6e2cc4df97794af24ccc4ddcf6c03b
zf656a7bc5f8082951a34e8fbff7ed21f791458912f17fc0bb03b7ff548c8185f5a5af0ca565d23
z63e6632e026ebe2f419c3dbdf2527602c691fcdc3398f00afd35bbc53ac3ed8a684e9ddf25b2f8
z2ca1d9e0a8a320fa2559db6df7f7f3d8ae93f5e1733f1beb8e9e2f00c3b13b0c4a078347727cee
z1414043b91b4d2fe991aea3f4dd698c9023a414da459b553c7be963d10cc3695f9ec56c00717a2
zedfbf0d200bbab87439d813135a3a307168bd88995f7a49950cc7f4e2a8b68612501c67659bf0b
zad98e25ef80a036e769900600127b92218f37bb4d1cda0abbe01a1ab2857ef8c42ab7f256458e0
z948d65e027d5f0d6240ab5da76192e32206e48c6bf50966d19be7677ce50fbec7c37543bac5840
zc83502afff8c2b8faa693bdc24999983bc5f4abfdaf5c75b55faea05665658cd5c0a24f229bc5f
z4777cf0edb6591bf7d5e2665a6ae328cd886d1133441ae2c9f8d8f5f41461631c9b00f57b9e929
z7cd4a77d4b4c985239b4d7266e08f297c3c130b1c2b057775c77b6f3bdf9fb7e3b1172bdc6c9a2
z2b22dc729ec7946e6bac651c56ecdcda2ab0d47f5f1ba8a3ba505302385185dfe535a04c8b3fde
z1365994e9f878c3ed0c0bc9cbf5a7522e98730ca00a6d24e2ee4c32f932785e07174caa9f71400
zf0e00595458df945c66addb81a1748095b48b211df217e6c1b25932807e55640d83313a95968b5
zadd5d898c6cab13278e5f7d9e219c2a5adfe7cb6c4dd6bfeef7363fb48423209519e920771aeff
ze2894b892fb2fffd63ed74593d573c593a491da0542b4c1085d98ff2208d8d3d420c2241447e5d
z73ce3bee24c040ff46e6e7e1d5e9c41edb67724d8872e6ef5202ea4871c8e6d00dad78ecaf53db
za6c1d40f38bbe803d3c126d30472eab614fe60409f7af1529b2a8c24bffbd9fe276c9d31313dac
z83585fe25420eb23447bf1d59fee942aee63346745812dfbe9b309c7846644c9600fcd1289cdb8
za159f85138c23a5ec4143d861f1a9af500a09d5b9692527bf924e2bab8cca4c2ee1758a6c3fe11
z2f33d1c2d7cb29fabd6ba88eed2b9bda7e629d70949a17b8462990b3a60b92c2a51faae7df3fbc
za00cfab366f447e54acc52919cb7c0d33f986275f5831da3f9a245f7b851c57b9d51c76986760e
zdd044790bef25a92ed96e6482be382ae59e395894308b2f52a89a19ba98750f0063f7ed014d39a
z0f91a5367c6bfcbf8494b489641b01b1f8e8ee3e2a8dfa413eaa52d9336d01c13826f0c0c74ef5
z7e7107faf2046e0c0124de509ffc24718619108916462c19cca9489b1ddfd34c1f38cde84bb512
z16bdc657310d70ceabb2d4d7d4b3fd672392daaa802fab22b26f673d718130fe5ed3a29ef3ad67
zd628d596e8150f5bb026124793cc2f0b81ef3caceff7c174bc75ca16a595fc71628fd83535c762
z99ad8e97ab8f83215c260a209e98689f5fadbd9d86bc5fcbe87226edbac294d6a77260adfbf64f
z4774e3d658f74da67727442790d04b49667190455880513cde2a82687d40c485a82e144e5892e6
z09d5d658d8d08b1bb430ea3ac4e04e93effcdeabebf8b2805098e7541added7659e8480b0ccc1f
z59c0ccb342cad6fd46282e366af41f731248f9ee934fff97ac3dc9eb280d74596d17265c7c1de4
z2bc02574f4add66438f12b1b0668245ef897e4a5db183aefd74af68fb7746cf2dcb6677df66b12
z618bb41b3263db126fe95f4c23f255e1f3705702b66ec0bf3bbc682b9bdca565962bd70494499a
zf48160ed0fa667adf4c9792b2b87a021242d063519f562182d102bd2dd8f6c624e2e213bcb6191
z890579c31e9c285d1e41a76f5dfb86728a450281bb33b30eef83f776cab322c6f665f46348a18a
z6349592258869904f39b726fa48f401837e657aff64fb9245aa384a8cf9d43f7a45bcfb3d7f048
z21f9e3da444e7e6af314a7c25b12e2ce6c99d5b6c9d1efd1ebebcaecfbfa14dcbd3137b2241812
zeee4dfd4796707c1020246a654a32c982c327646a301b75e4c845c56cb41051957a514483bf5b8
za70867fb351944c3ef92a4948393a394c0a42ce69afd6e3b4ffebb758d7d71262eb74555ea9451
z1c4ac25fb86012830d1643788f5453ed425955b382927419eb094f4032463b6eef1e4ee2f9dd75
z161f758cca0dec9c71607f460c30c4718897e749a2fd5e79d4c1bd61304f0661b7e7712ea65c91
z836f665ffa9d18068afb031039ddb1cbf2776897351de9cede1b577f073632c7098796a1451888
za6d260fb592db19a3559dc05b30ba56967bef964a9cebf66669a79e917dcd144e8a9a3bc86b486
z1cef14df3e572676cbc185509c97c277bb7c339dbd6ea04510ddc2b7f69d5ed6309fb8369b7303
z5c0a9c1e6f22ceb2af8945efbae8ed437535e26026008ccb954fbd5e991572b35a9befc8e25ab0
z9e18a8c78cb1e43d24f58afce13a8c04f439c1e92518501a1c791739198274ecba1a6735386d0f
zf7ffd4596f1f43bad0ece20060537e39cec3db97892047e1502de427f042870e90f4108b1adf2e
z8daee208c855e302be3e1b2e1702778829e903b6bb8ea3e1244c5cd53beacc34e10ef0949838ff
z05b0a8461cfe1226062f18700d2679dbb5a5bddca494189c16c8e0a3b79e2201c990f183ca133c
za2cb845e8661eb21906fbfd4388f09f242000d2e3c6a62ea18403b89e6b97a08eac8aa1832c6b1
zb08f6cbe37bdbc2f3e07b910fe288d39210f60cb86acbc436af417c5aaf810d6b425a5def1b6f2
z9e7f401e28e57b946e76a4fe78f2faf70efb750a7e53333ce35847f074d6b22c83908204201e47
z42f5eecf9d9df9ae6020b1053f242c2937c93a7ca5f5bda1c791a8ba5c873e4c12b4ca1484d498
z70aca63ed8045d0bf68f5d6b5da77f7cbcc9ed28bff5bfb6a6363d5787f959ad245844747c4eae
z4154b724b74a5e0d898208c1eebad65968ae31f59ed1d00265802acf9ea90545ec739d657d19ab
z89d0ff7a2a297ca2910edc0657bdd02acaa21ae9ebf1b571f8ed83f96acbdafe4eaca47dc9eea8
zbdd8d360e0f2b3cf0135674538292bf5703d5c83faa4fc6165f90c261fb6d22aa75b64c685fe41
z3466697c3db0f890b4f1d98d45a66d3ab9e200d1188d998dc9f2269cd7905e4033ca0fc83b96c5
zc2a5dc8f7f8000e546cf7289c1f2857e3bd141d3ebd78af784d454a60f01e0776dc92526bcb438
ze9ed921c3bafadaf627c681c2d7379f4f057dd63b071615fcc7f04b9d1c10c77c20387809fabf9
z1bb0782a6fd1aaf887e16b4053ac0f8c229238ff9d5e1d6e6d8fc09d3b42b9ac189d4fc712bacb
z2db2f4903f2a9b22bbb9ac7f8492cb2cf66836067f945dae50bac92f8ca9c4c76e7963306d0cf3
z2a49fea8c52431411becd34b2b21a486f95ba3330f1bc012877314909c3a40530443e3ce9332c1
z0220f3414ee2e5a25164a21bd60fad262f7acb2e198b832f46b7404c43a28be1792f7b16846318
z1562d9eebaf17e404ff2c70a425e73c77bd7c3cca1332d1d64abd3beac0dacfc60b7576be10125
zbd9337758a451a407f88fe8c36ba9dc7ff5514d64d18bcee7d311f9cafa16db39a38d989da7b6a
z71b55441f219f00bc34c98b953d2ab3806eb957bf642e71746b81f395e798c9a274e2b52d6fcbe
zb7f865452ec37d706ee90462d9d42656526ce1fe2c28d505148f12ac2340cd448bc837f1d68d32
z34bb472a8ae5a9808326845f0d70293f6ab5da6eeb45ab324411f6f9b5a01183b80386ff6eb290
z86080f6022185e54c0eff0f69891b99618413bc749cab9f09e32582f870d6e1f3409da4ed66221
za6fe8d128a02d696c84cb8a0cb3159eed2300419872481e4b42976fb219bb1a394b3dae1494250
z2485ffacbb7de02eff03d3d7ae32cdffbffc020d8747feeb26b5d97c4009b162a893e3ace27385
zeb271a304adffb34648130479932a21c2e11d8094ddfaa4f7968296be6ce7aea5c04f7e4bf066a
za48d2298c52ce0fb300140f0ee5122ee1103bee74fac516782550c247fac765bf943f2618c2367
zafd063a0d8ddb9fdb2ba4a3c177e31701fd4494da041c2440d243fecee7fe0a161893e7f28eb88
z050501d698de1b725206b8be8f3a822539f89f9eddb0d79ecc67501687f3fef7bedcd70c8f73d6
za8ce4895b33077d38ae7987a85549a9b20cd28cf2fb27037c3c202bcc2a4e2aea618d94bf2b7ad
zd0033e1395db83849496e92f8044618055e175e09ce9d7c67e1e9e75e80c2dfcefcaffdcc66a3a
z1d3c1e6cb4f8151d0978e97d27ebf510387ae75fcd167169dd957bbda54f81dc1d6bbdfa48acab
z74c121d33ea6a3885002ef8d0e6dc2f4f813154cb0f2aacb0501ab3eb9522c04ec85ba2ca8e721
zbf286489d87409fc783cf57682a0e62bb7067a64d06576ee81bc3180dc1cfadcc272dc46ae3e2d
z3e3018aba92c569b1a59731f591347b257dab5edc53324800f0a6f7d1c402ba259d1b5deb6c265
z8670f697366fa8eef73f8291a6928e95f23b43919d58a360b5a227e1bdc66a79ec2035dc27aa19
zedc0262cb8378defcdda97dbab34cdab38c80dbaed426d7bbf3a3266d5caa95def2e17a7efd1a3
zc42330e9a2809a188dcc30077938b1259821aade4596e72004e3999a0fe384f6752744fac4e06d
zedb27dd38da281834ee770b898c7a74ec828c2b6d622eb0907fe3827d294c41d227e2bd17f9af6
z2068e1aa1009d173d61127e20c490f689befff9a453e75427eabfe7f9f119afbe1e59ab9a15596
z975fb2dae21bc842022afff654c9b3af40a9bd155786d14b5f585ce0c7212a3b1084c5e7475063
z2ed297dcf8e83c3423051b732a50a8fd05783e84ef51d0c850f7833dec0a3584393669e442f9e2
zefc948d507d0ae8f3b5f32d31ad8aa224df85cebfb0add00340773544c86e154793cef96928181
z4ef2bd6227720ac8a9b177004f79816b5dda3935ce1ed0204a46f7618a57d6ba92ba2ceccdd2cc
z3a6f25367b6a3f282604c8b32e975cc6fee977d4edd9ec63e8729a1d22f3e8ef0d95a9ca6041c9
z45dab4c53a72a0e7595de4cbd9c1eaabcf9d135d875ab9931402f92c942abf6396c8604493a363
ze42eee74f4929186b080a0aa119f07c948b764240c65def3208789054c4f421d245c6b3be00f26
zae660fbe664c40bf85ab0407b3ea8849a17b9781e462cf31b361894c3a6bb36ada05faf5b860cc
z6328dd5b113e9091c8869adf11a441c0c2f4930149ef9c7de36b1fb25760fe8ff4c8f33adead47
z997488dfa1f58a880133ad3a1c688c2b1cef75c99885ba457f2b8d45940fe2c8e2bc4fff1cd912
z9aaf002e2019173aef522b159013b2ba6c81ef8f3387b2bf6b55c37e15e1bd522a8680b952928e
zc05db4611fe47c4668f6005403d84642e0933cd3848f6942ce11ea61aa787566453449c9bfe7e5
z018f0437b9d75a78733d200880b2ef64e82396e9769a8097dcf1cf9c6cb20c76f0ce8b46d45833
z1102420368d7c3e1d52624f3d434259bd37069f4052d0acd85423b8280038e19875b96df58bce7
z096caef945d4a53204a6c0027545cb3f0baeac96bf3ce4fab09172919da5ef6bd83e9deeba4771
z83c9289c99b53627baaeeee75825333a094881a1de92e1ae117b2debb651d08849d5cc4ee6d4b3
z26acffa2149797f20ad59418c476b43bc35a1d37ca2f2c7eefa8ad28ab65e823ad3ae4efff06b1
z8b21b1574c1a97052dbafcb797e4aa97f791592c718e4946f4bff2174ba6edd2f3e821183104e5
zf0ac1996c04847a645c7fda62a02510d9f2ebbcb2b4d52f6abd87e1074b66fe3f5b0364bd6cfe1
zc6a0e5e3b7f37e060d4da659228d346aa0ae74a4bb1058c27d7e2b82e46c2b1ddf7057a050cb32
zb0e35c2343cc20dc8bae5cf0000cbbc5dbdf98458d2a7f328703769f4dacad025dcafd243bcc60
z6da1c90d7a2c8b1f37f4a05b8e7063549294bb4372cd37a004f4ab765eb9b86f91b0ac7954c9c1
z634cf969c87694904812250bf3085b6be7cb69d3d65d9cf1dff824ae98cbf8f531ba339bf793da
z099bcaa3b64f7f4229b25f541fdd3f9423970aa7a973aaf9657af6c6c794ffc71df77db65779d8
z075b1bb70d53af47f3ec17ca7808ba2a096c9c0e8649ca5177f37309e7299e90bcb794f4c48087
z22f34e00f71975d5392a10dfd1d2fc2aff9d5eaf2aebc14f156516bb0790aba2528ea6d5e629b2
z1c115fba757fc6da65a3818d2f96abd7af7700398e95544ed3e83515c72c46456372c5101754cf
z92b4121e384033bf41328f078775cceb02e5b773d3832e99547119258d3951654cc707bcc76b4b
ze57d58e0d0d4936acfe4992d36117c1f8e0f2d3562db97d739f1b8e41cffcb6024d65e511e8281
z802e581a58081de99d762f13e7a6ca238d6ff0dc1f56a191b313e6fca07377a708e2e9260ca9fd
z8a1f1448933ffbb7f0c19104720ebb037150322fe15c325806a03664dc5ce6408abb6093fb65bc
zcf0bf67a13a3e8a4f9ba4c3985c2f66e4e5c4b4e862108035349c77fcfafe61c0da8614dde6732
z3c7e3cb0d7c8d7176a9a47cc267c4a9fe01133342118de41db98bef6c7b0a0b5502c269ed929d8
z77cb7a96ba87f615fccdf8f03b931181b896f307ed5dafd04d4889e29e4365c592fb10785a23ea
z0ec5019796923228a66ba026abcd15e63b8f88388158007038754240f5da52542cc61be1f9993a
z88566523adc754fccee6655ffd9932516f6fec9a59e916bbbd4a4441232087fc25458ae946f559
z4429a9f9e732443774424e4a17517eb709072deeb367fc8c689088691846dc3d5f5556e52a923a
zc8362b4eb136787e67348bb309701438b08bfe263aeeb6e78f6f6b5e135960a73d66bcdd842688
z2f133237b93ddc94d75bc2812b1b86a358d630b39fa06d79b9af1fcebe83c6aab8d306e3d40f34
zff0fa74d7ecf80f640b8f6db32508cd039acc191fc06921a742e17a4dc4d52953df83694311c09
zef5063855a9dcd34f01c66b9132b37d9935c0c9d2c5dbe9c2d32f0746adfe061eb7fada5939d94
z57eb39ffd100c08dab6d3811dbaf027e971807f5498a10d1ef7278da3aca1daafbe02a4dd8c7dd
z1e9ea344944b9e23b2c358d7ea4d85b9b5089a08062dff84393b6b695f1bb5f4df34383c8618c3
zd0bcf75bc0454572886f8f5167f80bc70281f7c9eab5fe638ba5df8948496ca9d8e2f00cb0b69d
z7c0f7d0acf484ac5cc355d382f8659d73a170a64f0958c81496db5ff232b4cbbc38e04ff7e73c5
z0fc6130aff59244a98699f6d1585f0165770b7716ffc30897a59db8745b93bd0c6de22d9c00881
z2e4520ec2a108c61ddd331d69b9fa5d6824dc56b975535a84c8e320340889e6d8eb87508ca3f04
z103e0661a899dfc874479d4c03dc9c6cd815f685f31cc4bbc8262feb4b325d1e70102ab38dbc35
zf64277b329b99e4b739be35ba24dad75a62a7ca59e06f79b7e3cf736c156f65325cafc2af4b25c
z75c282b51ee7c7f96f4c2e4cc00cad07a2ff56e2b046a7bac72b8c37044e1e117e1df3b9f330b2
zf19804725a133ca195db27b6ae5320e32e738bb772572430fa6ff17e58170b86acf51602d2e230
z52cba135f9d6eef61870830b882231ca4f183d3b09cb9d4325b2cc618b7b5eae22c005288bb5ec
z443e25cea1641032b14aebf587fd7c8d7e4ff6cce80ebe61f89fc7f622655c25f081109b081738
z0cd3be0d0d6ed0d29e6e55c6435dd55f5a82153784d190f23ce9aea32e59844b012abb8ba61159
z9ba66bae457760ca0691a20a3260dc0c68ea509a170e813b73a414b70d1ccd514136ddade3842c
z76e9c0119c5ede3e434e223386c14bb17852585c998af44c213c637e3a08202d9303e0c577bfa4
z425d03a8a048c19a0db890a313908aeb6bd16d716a7774c27971ce3fc82200df0db0b260b34203
z2a3577ce247ed181f0993b3097d6c8db5d6e0c3b3eadcd99fc7c006f846f8645580db530a5f93e
zed86a039ff158e74b6a5e62f6fad84ac5511ab12bf075660220343a997b473f0aed90159e61333
z5a1d4eca75198eaf4147ac90877ca0e6227f05a6961fb4203ecdfa5eceac19bac424f54cdd2769
z926b33c9eb4352b9e442edffe32dad026839dd991157979ec742ebf30ec72220bdbec4df16efd0
z24b202a066200157e3b5c35fb989f3442a4526ef92b671ecb25c67a0609fbad46d12222407e68b
zf14cee59be91aa39e99ee593e7c8466f31b30f5572b0fb8d050a64eb350a0740b0cdcb1b52af96
z348ed26b1a37f9f8fc590e89b6b475f3dc71ba5a2bf79f8c198cc4adc1268ed6e795093aa9d125
z8d58688f4e06a0867e53a4ae7e43facb6e8dcc60ffc1a7608dad55b183436a3f428a37f94a1555
zd2ab1ca72d4b20c94700928751e9953592e52ce4fa14900ca4d41919dc4107fd8c9b99dd807df2
z31c995874f6d3d4252f77f838cd560e9e9307611723ca44a67dfc2f22617ebd8d31c063ba7be77
z6c0e6bb85944b29ad1adb0f5faa898387597a88641d87974322b7aa3dd3b5fc295fc487dd09c4a
zebc9e10dc69969dd450259eac8c75ad31069dbaa76eb5d0899535f25367af1f12bf0eecda267ee
z0bf454af99d05e4c6bc0113a7304a21c7a945c11a023c85f8bdef84f9fe1524a24fbb5df0f7987
z1d01ad81f45b75aad24890aed40c416ce19e7c8f37917514c1358ecb04561eb9cf3e34cf2c7ae7
zbc3d9659c591e226da724e403a92ddd8d6befda3394c69aba07e490abff665dea54b6a16bbdcc0
z2d315b351230b233981ee5a24b63a77f1814880aac62deb46fb7d1cc949fc67d2f180cf44fc7a8
zc0c4859fe648b196477fe2ecbb643f96bfd5aa6ffb3f79f231bf14689150d054e2dfd016b5cc57
z71b72026360319dbe4196e9110d135da9ddd2254bfbf0263f4fc3368adcf29d7b315dac9121dea
z42eabaf3ace1b366d507e3dadb6e1e14a7bfa14361c10409240abee51f3bcd0611f79eeb2473de
zafb9b461e74fc05ae0026f15c839c2f2d571f23638d9c306f3ae4a0411af276b41177a2ab90916
z06bc40e6b153a1666eb2229a98a3d911afe6bb706f480b82f1664a2d6da7b8be6389b51b4d2ba2
z3f101a272f48bc0ac6e69847d8c7bc2122355b34d3b0fad83e370bae18ca0a60e29ff7221d186f
z1acca91317e0d57705b4091e0e87b9615fff53a901acbf76cedcd22fb85a649b25399cdcf105a8
z0e85efac701c8cf21a2633b9f06bbba87118066f763199dfb27fc600ae1fb42f2dc135bdd341ea
z19c3919728928d14ec7430db9aff6b24d2c8a68d9c54a78fd9f9c41c947eb7c2b171e66b095394
ze98d9e09c3a255602a52b5d958c81ab67a09b8b9c103248dd070219595b16abc23f9ad4f88bd1d
z1a5befd48d319ea2b93bcac466104f598a74f51539d799c88c04d33000c6c0c13d56a215720f75
z13b7fa5f2268439f1625740fd61acf73675f70b7c7e55920c8e7becb1784aac4fffe8988475e64
zbb191e894ae381f57ac7607e1acc52efbde21fc112cb8ec71cc40756ae4004c1b45fd7326e5c10
ze31cc95c00981e1e50a2b76de671514ae01f1a435fbe44a4c1ccde94250ec2d50db8b35fd70054
zf485d91521dde2673e3d5cd7908ab9be0e0ba19b17ed0a141dca911f5e2f32a166d9db10cd6038
z03010d2d0d5fbb97920edd9aeee62308fd5567742817575e0f5bbc5f252ede8b40fadd8e0cbbbb
zd7070ad8a100724782c727324ccc7d84e12a08e926f8c328a88a082c4fa9e725539c98492cefd5
z76ff9a38c1aaa78c1376e65d3e15a0c8e094867a73b7549bb27bc7013f18eabb2e362a1c6c77be
z5db4b927112473cbef2f0dcca6c44934dc0e53a65442dd19e727b9b2b58225e88310e2c82804e4
z4a4c11393e908b048481bbddc914a53f07698f98b5e52a376754485b4bdcb400d29e5bb842d8ee
z69e003400c4e8c28be665d11cf59e38d8b735036eb4f7aa53112e0edd999f59bd4ded58760585c
z18631d5ee3710868e57a550cc4ef4657d392730fc809082768b1cb4b744859475eb07a8ea7f7fd
z0c585857b3664744952c1632202a2eb065c15036b1f42d65e75c8020657d92939bdc1a1e3445f2
z7cdbc5dc17361b60292d2973cf0e5113360ba4f1b4d0bc7ba97bbf9be00164478650c95fc239fc
z69c05d5bed67380a6ce2f4a9d64d5fa50c013e170aa08641268157d9cc6e60bebbb5ef4245c7b3
zf53bf51f691ac11c7743c157409a94ed189cb09d8675135ad2b8d082d30d045b32c8ee5b53e8a3
z231f56bb44b39f4803f7000b67bb547395dcf79677757cc8561289ba7a78f7d54b0e2807b579fd
z5858761424747d3a6f626867c6720090e60071a01e590bc344677c6e180b37448612378ca628e3
za8e6eeae1ec0e9d9652dfea5f7826b7f7979e2515254c3a511f61fcd154d59ead037aa478e834f
z59004fe127707ef62ff470d204588d6691333b411e17c25fe99ec7df1cec4e1ed98cc3ca109b3f
zf19a767b1a137e77d065f2913ac8b930833752583bc896eadaadb521bb0a2c476828bb449191dd
z2b5ac39a22a67c3910feeb287e51605c0ea9cc147317a79abb02c64f2d9377a4732666f6f94f04
z107744a09c30d1a356aeb0dc3b86813e151c01214a623a305c732e34dd1d44af9f770ad8be1c47
zb8fb3fbd98cec9788c87dd6dc613221ce2a3477608de7bb8fba46c393550fe0112660cb922fa13
z2c01ef69fe79244881fcc08f255ff57f4040e29389f6072a3dddc343e8b9942b74169869ffd2e2
zb1298b4c9c892cf77485f94f12dd3f755aef9d036eb0af7eacb72c8ef5af8611c9c607ae897e7c
zeb939a099534a1af5b9c3cb965bb16d84086a1a15d3618adb743493c0fee8adad3bb593c90c56c
ze2c539c767476d193847d5b65c4d3f35361eecaa3d033d0330868a11f363cf2aa74b2c1d3cd5e9
z3d7d43d316208367629fd4df9b05fe30bf8d2cfddc815deb323bd58a4b494d6b4ba7e1894cf56e
z90f949116c0a9251f1d2e95e16948aea71d16ac603eb31eca5028db1ff44255f3b7628bbff67a4
z401bcb666d058b69eb1443a7d597ce7940f0030dd58a9f355550efb3a7540557acbe650e44274c
z3ca5e5dc8ff245802f2fe49b98c9bd215004c43cb3c216b314ac71c56eae2b7443ecb1ed481762
za2cf9aa77fbbcc261f7859a326f9fce091c93914dee69ec3f862f62a49c6e78651f5d88b50b559
zd5f86d6ec0913450edd02cb420fd74af2276f8f44ce26d0b6c1a8821d3895dbeb158db179f6794
z3c0d5fa762f8b1f2f047cac55ed0fbae3f6db4e8fd113d5d6bae9c77782c7256b5f9042894c18b
z356b31b2ddd98e06b7ac35278fbfc57e4db592a9aca46d3c7d115cf9897b8fb16df4732f3ed183
z2a87dc7b2dae34664d402e1e01d63a8c7c10ec0f189922c5d3e3bec2e12f437e6d460a71d873f7
z0da4a7213027737bdcea3097a58ba390790038899291f08b61e938e67667f80bdc1ff0e4cf8b9b
z5527f905347a2c269bbd835d9c31055048b6d12f7fddfff7c997f82e4098648baf275da2863ca5
zd4885da3caee2c6554ffab027c77f2b1f97c2862a0a5df54b53ac2717503e535251d1c3935b342
z850bc6a6d36b8ea2b21329152e16199e6413f4ae6e78d3573f752f44ce06af02a97c1c08cd63d8
z48fb85fa7f88ff930c1513ed47fab70935deac3c71a198ee2dda996ce5cca3f89a5761903990fe
zaa02aff19b11bf707e0178195b835bfd42ecb09676c5317d4e2a09c6872fc63aeb9a534538f4f6
zc229850ca157df1d526830fb58f86a3482d9cc1460180a3872d8cdebd5ad8a3579cb69894a7500
z291931b4b444c6d9134b14b277cac35431cc7542046932f27ebae4ef29179156663f2a3838ea3d
z04078b7ebac7628cb741812709ce6efafe7c77d947f93bba91568845e8dab2d48a0eb0736132e7
zc182921ce7c6454dd0c5903729d4c049bdbcf21093a813eb6dcc78af308c26ff80ac42ede9f0b0
z531a20d5722ce2482784af5de93053ad20b6dc4552ec7b297f38f81b6cf26ce7d92e43fdb81bf9
z9fafe6c62839e5e8df5cabf5be7c32d4f0e4201e5a683279afadeeae2a524b5a1da004af48f1b7
z54e312203c3dedb205c63ba685364030846ad9f3a0cb39846d213fbca44863673ca741cd30a64f
zc091504f15e2ac74d85d03c5de82bbfcdae2921abd8b45de56a50b091b210cb43e7acfd4473fe3
zf160e39931041150312c133432527eddc9aa2f6185c4cae9a66907dd8319e8b25fc0644830552d
z57bbf048305690460e691cfeb51c1bd4dc55e6cb24e8bbbd8dc1181d0b0f5e2fd8aee16142e772
zbb79e48b9d29ea0026b1d8cebf5ddbec17ff1c853426b56a7fefda5e44a81940395a18916352eb
z6488b215060ba81d25aa79c94b617d44dc68df5b1ad5b72f5133f22331e78dcf64bcdeaefd58a7
zc9235c5ef3c5bfb440ced210b8b890af5697b4893fec3b1ebb4d72cca23c266a5f00ca2047519e
z2a0db7507aaf8cb8dc581794c32adff46c0a13eae113a009e4bee52e595924b8860f9304cef69a
ze94c9376e110bf72a161f053ac8976cc6c0f49a8e6bbc01fecd305e4f18112cf625a272139a01a
z15daaf9c5d24936f579b48b1375b55f6fa439eadad512f74579d6c7dbcaed2a66fe5cb49b988c9
zd04171e48ae43653335e67fa0e85760bb44d0f1d813f2a334e247daca2c4349d903057347c26d8
zce610ef5217a46d66f6e6308b18634177d01f10b7c4d3ff7c8a7974969192660942ea3b003f740
z7e66af31198c2c792cb39a7c3d028760737a6979835f4e731594bea4c5082f0bd202ba162ec6c2
z6dd38b9f823c93bb8ac63255c4a77f06badb7cb8fbef7396617c491c55d06d359505ee858df0e4
z1d98b61c54b3620cb246040d702be0bbe61cb4eeaf754a04ab8eff69b6a0f9ca148753230bf676
z2973bcac6eda4e22a75240974a95defebefe4422c037d34a57e2dfad44602cc132481528bf6ce5
z6ca930dd07aaf2ca6215f2bb964dd2ea0c84160e0633d03d8d1420363fcea0f22713b376655907
zee1760018eaa3c4506f176e17c8b28bb766bc20af3ae540b58d6db3669669efb50c9d1cb106221
zb1f624698a7d1924dbd3b686be6b51c476253e082e17cd9f2ad5ab876dbe4a64595a17efd6cfd3
z32ceba848a3834a5bc49b707f49cc01583cc99402797e1ab94287453bde03a3b264b70a26ad4a9
z03e725626f7f2ba83a1ed23baf8594ef5d554ecd1a742b762ad60ac72b0d6821000ebbaf9823a6
z587f78efd98ad761bcdd056d0e83481a174726d3f362ccfab5f42059aab80180e727c4ac3f15b8
z725481266a728d0762535cb2ece9d6700135ae7579fc64ad8214d51061b386cfda3202f7a31af6
zaab874f983fe028fbe14fa6bc3b8c024a6efd85fa68c0d59b6ae4f5ccceec892a497ed0ef63264
zf506c8774a8f9dcf4a6f3c65e7ef453a97ef06d7be842f6e2007cc592b2a0c7142b84ec8762351
z2e4d7ffae577d2eba89f853739b38a5e4937bf234205cfeb31d8f021c4144f03527f9ecfd3a9d9
zf370a7a3a669352a35c0e3d765c1667641a94abd0d62995d97da88c9990776fe52625d3fdadfc0
ze077e7f6f77bec9332003b26b51abb90216bdc7847d230424337416fe8dc3284ec35b0ec8fbe56
z5f7cee49d9c73b20b8e3e3ae66d42ef286293a4c43964eac6824b755dc47f6501475ca43576585
z0377451ca4090a06d5cb931de73f0a31fff16cb2dd8c98b6bc97b941361085b945d2b9455b92e5
zc6092387bfcc3575d3eddcca38a0935eaa5c0eb9e5488282a2b1f38a4787be7ef1fdfb6d6456a4
z0133bce041c328c073ec99ce1a05866ece6ba0cdb73e29d61b51890ec06bd37a6d22c78cc3e4e0
z6aa4e1a9122efe9616e437743b03911a0c5816efa596cc3f4c9a5c74c5ae1ad8ea754e9552625d
z6397bdd574104e890a9605ecb4b8e3c308fd898c58de4c4916a33796e810f8951b49c6686929ec
z62022f667f8790c4cd5e4b940195468bf270487f307cfbc5db8bf0ba90a9b6625c9bcf422a9e39
zae178a4a190602c45201152b1281fd7f0864b7a8560d89e96e11c8f6bfceea16fb83ca7a1dd3d0
z01b1ca14f3dd7e0c910b268bb211b67be9e888691a4880525f718f9f45673f389d2a9f3b11a746
z93c1a6b1825cf9143e2c3e82273a58f75859e145e18369e007f4453cce38dd7795c76dabf8317f
zdb291dacbad1bf492f9b7fedc432067cfddef07a0fa76e627da7c62fee22cfccc95798954bc5be
z36e9d7196f81652df849eeb610e0672a81c118aef9b25d4919faa0fd9a222222be083a28c5d4b7
zb47356d56b2471daadab218be74bec3821f87743e9b46a8defbd29acfe198ba725684f6dd91157
z2f20c5df6b6ca55d440b1f261b75526c74dfdf59985057f1d2209092cdecd1db2d4873452ee806
zc9e40a951b6283746f602cb1d3ff4f7119f34278515764eccba917e9b26aff923b1562ec1c4faf
z3112ae0cddba6101e344bf1f4e56e5c76c75c42f1c27d0bc52fd31f96d52a8b6574a025741cacc
zcc694f7ee7c675ca0a43b473eaec480d57f280cb873e8ef26364bca1f770d454dbb40af08834db
z0ab78d8a0dfc3f6e199ee1b37b8afb210713a2557f49745a638bcd0d108872b83f40a54c780d53
zf5a5242b2d8e369f3ccaa28b5ac5b1b397fc0175db712792de3ffa56b9bf050bc0ee3d5bb43f7d
z08e294841b6fe735c2fab75d73ac274e8e6aaccf12729b034ffc00745805b837b90a3853882ad1
zfae8619451a6431f48fd2f5872b422a85185717191274fc365383f459098743e0712b5e4bcf458
z7567ec091c40d1b53774de68d925db546fc7e3c1c920cfcfe9136a12c1d71e07b485a749a968d2
z2a3ecd5c8f2f5bfa6e5ed750e70847b5b45542817214b0ac13270b1338be41caf80144b4a5c963
zb77c4f340f2b6ce61bbf8f5b4b6408dd3b2acb86b040fd9b32a8b7d331ac96f9bc23f78e28a8e8
zba94e6c2f16b49251f3e7759c618aa36cba634e0ac8473f6c05bce6094e0d7283696a8a3904521
z7feee9b1f3f9c8f2307a2ebc6adf650717178d7725725f318a1e1e8c83b94014f30a42bca00dd3
z82494e4c1d9ff83f0d18bf176e174f4a877425bc10b393f9b190c9a9082585326aa229c26a05e1
z4cde63a69147afd9ffdbf89ee6942554ce8d2cfe353bf04e8d8ab2fc1783dc094ebe9e32fc95be
za5e3350028f7400ce27213a8f2ed4b4c303d8fc58af91394b825e24ee41332f9570fdd2d71b8ab
z923520f7bba05d9c19c9f38852a961b83f487a02a997691c576c768c5f438015977789b3701502
z991302fa6d4809f579f6388c2848bb9fd7f40c191d3d91121e8f8f3b8752f4737006e9cbbda0a4
z7fa953053111873ed63a418626bbab06a080e8285b9bb5d74c0cae7541886d6fccdd761b9a5d24
z844c23592a6fc372bc11c8a3e403ee1d5d97b0baeea8e6587f081e6bf2c75d86fb0d9022083f32
z34b6f8cb072082acd1046901680266540c99bbbdd6ccb81b0f33513f1dfda9f52ad9cd37b1f434
z3b650106f54e9eda2b7c65cc7f5653c87015b4bc7ed494bb65a87225891d0f2b33b9a949c568a8
zbbafd6e09681fd48de6ff843f120a9b8574cddd78d41c08ad0c4a7a83a99e5d9b3c1cd464598f5
z605f989787e60f7bee10022826ba45f917d74c81b1095ca9c296a55493e7e3870d702b54d65a4b
z2120cebc8e691a0c30ed5ee6be45e869aa44f07ca0936a3cb4dc3d3ebd4b7fbf313319eba5b721
z72b83c0b11a1a60787f0d84145507bf0cf824e5b371422d688f7f64f251165b60e62a475ab31c5
z0308dcc71c63644a366bcd585896bec20d01ab3b9df46236629506033f68e460a5930436251517
z977dc5661fb47245b5caf06b2ae20d060605d165d1f81e1899b23035e8a9ade3403edf08f7f41f
z4b7c6276d2c4654919cad9fe86dca65c9159fef1ab6d30b3e170ba700e29f74e0f9b4d5d64d104
z2a014af7e93a4c84516ef792987b2df4e41b33fb66dfdef89ebef897ba18623402561cb6dc58d3
z999fe94fbf182c8faae981bc58559bfb934163baed5565603a8a53025883d658e0f2f999138c42
zcc2217cbd8e8f6e23d51a96528f4cf99d5584710caf00368fe1dabb0c0a6a67995032aa68310fe
z717598c93dbbdb03eab5bb0120e2c95e65e64ba0ca21fe128dbd064cf3cce81f3b432a263eb672
z742a9dd2b8372ed7105b53b6fe7161b181d28b2c9604516e0a2dbffc050f4c87bcbe2dd7bc5503
z92f0af8f772157b4515bc3af3bc28b173a3246a1778ed5ebf588a9818619b7c61cf6cefc88efff
ze21890659a423f474ee38346881c2d50e5fdaee813fa23e262bbceaafa92366be9e4715e75e85a
z231f8f538ad23d6c0a0f598fb48e5a07543fc3c68dc242dfe56eb77d364366239dcc97e3d022ce
z8ee3b6643e72f1bfed2f4946a498b8d13e5a103662fe3e7f011c413be735575e714e9231115ed5
z9907b15424a8340c954e88e0e6800abfdab17d69557b94c2ce36bace582a7e925ad42dfdf6771c
zb7d7da52696653e20a773ea94c764f2458c74f5115a59465057c424d308b28646dc060baf1b6fa
zecc4f0ac0253cbf4afb0dd1ab3d4414f7244be0b13040e7bb5e5c0d3ff52a750b3a197732332f3
z9e3e0c43b904ee4a04b1bbd5e05541b504c587c1c9d5d7212cecf980649e0c0dd0b6f215989702
z723a41a88216f8a5abd0297506a78447770fb0ca409c8a8cfead86667ab445262ab2d4e4ad5b20
z6859ebc300ed632ff61c099c5bd48ba80024ee5840be53c40ca2239521389d46801b66b6bdcc0f
z38468f477eb5da15a5ddd0b2afb81f7fff7256e0f3c260cb7ba480fcb189f5bd99600c1f60ff87
zb67d3cb5ae8227d27a156b6db1c4b9c005091fb72daf11e6647c0b88a1bad40d805d3f818011f3
z2bcc7ed25ac275c3f86e7e5b9f1cbf41c89740ecb6741c98a25691968b494cb5aaf89db4d99948
z8d46121e2d90a98f3fe9dcb64aa6eb9751a7b2002f9800982680a3effebfedc030782dc0b70727
z26c2d37f99d9b243644af1f9271c30503613bc3cf4db0a1f5de966181137f38e82ce149c787a3c
z91da59d4dc26dca7949dc1a2b892040db308458ee5e8a3a1ba6ee8da1e290f12256d0c0fa95214
zfff98a6001d1ae18443f6afdab1f7414ca18e49fbf19602ffafcdbd090c9b82e66f34c2992ed9d
ze04b6164ec6298f4fdeb19e1d5154db8aa03f5dcd21a4fb73f7d6b16dc87ff444ce383a5ad36f2
zd7a639676e9de791d9d0835f71c5389679facc6067b8d6679192e0745b8b32e263dc93318b9061
z7fc436480621ed2aa1109515829382ffcc103c1544992233ddd39524181a15238743988cf61d7c
zd029a72642e7e29d670c53a5f6935bf20e64fecf17ff9251b17028c059b5ca348b31825411cfb5
z4f708a0e6c21eb9d57fa18a9da98bcdb89c4df19ee211e459cec2ecbcc278476e0ac23e9a06b30
z147aa7bba1eebed599aa599b29f1532e9ba13e16460f6d91f69fb7060557d02b4d0323269046a0
z385edc50b7859b5e848cdf6ba68cf8330d7e4bea583b370b917104fe45d8ab090a3d8c74579913
z41f22a403f5a8ab7966de400193903e6e85fe2e48b2071a3914430a00942dce573bec989e18f3b
z4d7b6cb4b2d6a9bc5d2066118719981df7928d34c277333815f3ef34490502bfdda31680e7ee4e
zf29e5c3124fe49bf8327520daf360f3a47190752737382b3401b7b69d93321cbe6cb20750e8268
z8a4c8a332ac258d78147513f1ed3df0905ab44ca301aba576ec7c6e3c149700af95f78ad4feb48
zbcd957450b08329df44864a0c3d8ab6fb3b6db6dad93272965a61cd7ad68ce37d6823e6a73e6fa
z4e3d731d8f3de010c00bdbaf58a4ce2b3a5878681e627c3bef15c2b91ca5aa509087e7a2c316f7
z9f75ece4ac5aa7e62c4f74d093a787f458399d2f4110c7996dbf1db62fbac3c0745b800a67f912
zcfa01962e2088a770702c779f4ee57919cd3c28fa44615b8dcc711bf4491123fbd39c02981e1ab
zc87b714e3a3325213b4903ee7837da0c28578c979d70473109f1761c140ac5159fbaa9226b6c8a
z715795ed73d72ff61e8c5db9c3eeb4e787031df88f8cdf7be30bd31160dd049c77d295a90d6a21
z0739985dde4a992661e66f7d3e3666ba32ff15753261bc1b24d228166422eedd15c25025829cde
z129a188643cd420e1d4bada9cf8c482df2cb16bc9103eadf9977c4fa7d39f79663bc007d780492
ze430f3704aad20ffb6fad6f931fd9b8e8586e4e9dfc86cc185e23df772ffcd28abce65370cc18a
z34d29e065d01bcabac8378de58edc622bb580aa7703e98e717f83078c25c631edf93a88f779a56
z89460c9d3f0b285de6514a47a7a747caf538ea474d9b7c5b949aa4c50b3759663ef43a291c2fac
z86e3ec50914f16649e549eb783303b20436c170f74930971f905c128e453c7ea264f948a885eff
za2f651ba601d4bee748dfeeee98c8a105a22929a9a0c7a92d8681d4ee72ea374a108effd4ce9a1
zbf21e68b24297c427fd3644b2ce6cf8e7444c41d240f60880d7f354805e452cb8044981d058ff9
zc18b90e35b6b0403085bf41b6c57f4828bf4f7f6b6a84e48d0d25d4de12906d3794eaa54274c8e
ze6d0b828b33fbe11df35ac2aa9ef8fc4b10bad46893edace0d48260e5c03c6e22173fa28442383
z7f2372be7d5af0303a2aaaf585d80e3eb2c40630b89e86298dd0d475c4d0fccd91513dc6bc8e2b
z99644a6e029ab777111d9b787b51374b98d26fa9b6c37f221ac4f93617e0e749b46c130e3ee82e
zc8a1f3fe3c6fe90d213fc09cbd6c55e328b80cf91bcf1107aef407e1d02345d52b5d675c1eaae3
z8d18997a3f4cd0c9c281e7c965786c3eeafaffe6bdb91f3b924e49f730a84f102644b9c1a6fe9f
z91caa6c962f7d982d0e75ba8f3f4370f02d13d9fcbe16aad9fd918ef82004b759f2fd8f615a054
z11eaeb46ce9fec4624b7e3cba3fe41acd1c753695a6cf71f7db5dd533be3d1209b84318eb411ce
zeff9576887ac11a7c2161fcdcf6d1806d55a6719f93e8658cbe78eb6c5c432779712ea9eb99a96
z7bb61486b6c8db1bf3bb20e4ac74c0d3e5be6deb8fdebe6ab9a839bcd37719d89846e26f638047
z26bc5cbf5585e7717d6083f8f3fd151db56ac097f83808a4244f6d9e89965421f54a2ee00381c1
zc0f979bce62fe747c37194efe0157cebc55f633effe4883e9bf59958a2a7882e0e32964801c6c4
z3366066f9ecd2ea2808a724b095f47329fd4a531af9eb1f57d1db219e6c5a15f14c1dbcb51db38
z26246ac416ddb165e1e9402ad7d93a84a675b2c8bc78e9df269ffb4836be4c77382fb494343136
z23c582a4dde6996441d249be296d06fe86bca847a4369db36eb2e0b7e805f29bfceba3ab0b9b73
z2fb67f546baa38bbd7aa4fd24eb9c9b40b8d20ac8aae577367218b7eaed148fdbbf205c924a9f0
zd5be1fbfda4add30ec7bac79317350225fbf058e64bde08838b1c2c52dbce8d9138fc01cc969c1
zfd3be4cbbc9270bf714af69569a82da8c2ddef5658bbb5f62da85b2a739fb45a267c1ff1262283
ze65db8ee4a19bdb06cddac14e9e69ba02179d82619b9e54b5b7a67a4c3175a36deef26b5adc75a
z0a065a93e66affa593e8d8c7217f085fe130b3b60b23e8d8c1fd47ff76deffb0a5fc431cde8273
z3c2c34411f01c383a287f93c920c87af15a74a4229cdb2e4c6715804cb7b25d73ec737ea6622b9
zc7e0d80de0d4bea3e1acddab000f4d383fe981db0da771ab02f9249020f774f2c30bb50dd22b10
zf464b4dfa9af4e797509e884b961de538ede6b9f67a6e5f940123cf76242adc78884d361cba55f
z97e921c4f4e04ea83c90c18d097d3ef4abc5dd4a34588b0ee0aa86403ebf0ae8902c5209f427e2
z635e009fa8baf501cf219f54c315eb4e14c7467d195d4e10c34b0c1d0b924e14eb4644ce6353ca
z07aa524e991be00dfff52047e929d8201cdc45cebd8dce0c9d1c4e67e775533a26c701f1c5397e
z1df2e6751e6fe4af72e363cdc921bb28e663da108361b9468d8e95be9daf8f11b65be2c2801180
zac3771b75daead9de42b5dfb46fade61d9513fc3ecbec17b6ef66e037f10a8c5c9d5559848658e
za525e12b2ecb90bec347cc01651f00cd9b88f4368873e21fc31718f16757ca9d10c1fa0b1c7270
zb7ea0802588280467002c20e0d7dcfb06af49359e2f06f165c755e5760c6f83d966882458d1c82
z7074948fa5d919f6ca9b5faa6736d5de49b18e0ee3959ab5909fa916168ed4ec4dc60647d99fa0
z2fc61eb1da0bc5eed992924455eb9f1e097a74d0c777c6af26fa3d20f607f6655fcd408d573e75
zf02055e2a4d99be1e111cf97fdde6198276040c18b587b244d2aa8403607fb9503d25281b78e40
z4a21ff69549d137fcfa01ac55c0ebd495e18e16503f6c67a0ac29df74e2bdffe476a7421cde505
z48ce7e74ebf5c7f8bc43249e391798b75cd58040f951322e6ff1239236951f57db1479829f5591
z62f9838e892ba107ddee0844d46b57fc2a044d2215c1c2b671bce194ee05fa85a174a79093b431
z5afa63bc996afa0b2b39550c134961739a3ff5ce18a48fa9e0d541615eb68930ebe50a5a79d8c1
z6a61ddb7deb070a7c5cf8a3547b4950d30c9d3d2cef9441548de9e5b61139cb4fb4423fdfba467
zf02aea638cd9fce929dfcbfe70d20296c67555e2565940f9c19454f84bd669c52b619497da455d
zd766f98807d5d39cce5d12dc405b82a1e03136134056a7428642650493b37d40006dd115be2276
z195e94c911ddde3836a3774cce7ac4776c71d34aea51fbac54a7b7571be8438505d2c2b0f2441d
zd2ac22275b56c515c4a479bbb9af5aedc19d88782f4636cffe156d5413e56b237fe5c534ebcb52
za8ded5c13fcc53886886adc55dd4b1c60e5de3e67b2c556fc8ce3c7ac7453b5f67437c2f27636d
z23ffc53e55b883c0103b7933482bf2813b4bbf11af20ee7c7e4f9b4aa16d068204c98b6e5d4123
z44b45e92b037554b425b973c484ef0e06401de412fd10caf0573c6c9a38cbd488bb973f2448608
zf94b870673e1e25ac974688a2a602e44f717b882d0692c22a0edc5b5d88da447d1865bff23f5e5
za62ad6d228b9099089266e4ad27becf015ec551874f3912dd95dea421b3cdb14c4823b6f9d2681
zc5f64c8141b8c3f2c96bea94b6da9bece10646e9b15f96f5471bc45782149a6296099541dfed06
z838db810af339df39abb72f70065e854594264baab6cc3c230f3ec9cb509e3173a8ec3b6be28d7
z85541a4fc48bb034dd941700d5cc964af000d190117925f360d8ef9f2c39efe06de6eddf90c274
z42ac3c1bd4d8be164a8cee05ae1491aa639a9389e1e1160c26c257db83beb9e0bc055030882e36
zc9672a1a7f9afcc5f2547170269409291edd29e4dca9a52c5f662a245b2537bc62a955d6bd4f61
z671f4aad747b9c13068c2b3f0096032442f70df56fa2da56e42893729604e78bee91c5081578a3
z9f29de10942d5e010b6f638d2e0aeff4630d04541891702851d7c6b734c80878e1db5053c40981
z8157ae2b7a3b6c6ae1edd387716fd09db178512db6a6c9664f14b9499215565c72025e24b46563
z8cf44c1dbd650056b3c04ff31e0f1503ade07008228a7aff178bcb1cb83e65993e44b1fd80dec6
za2b2077f78531f0da8887329a27a60fdb3babeaaa4d98fa6d9898d5c912b20eab7fc34eb973353
z302d651de7799d182b63c3ee177c08545dd2adacf79be52232a1f4a25ca3c51755c09f17c4db6e
zd28d60913a554277638e6427846783581889a9cd12429f099d3c150abfae0b0cbfdb22d419d020
zf5604f80f9a99910430f73792944de7825b67a9677d8671a65aed9dbcb491de453962915801238
z150a1651c6cf16c6874726dec6b021d6544b33e8dbd1636552e32bf3a73255743d8684b9216d10
z456c6a0078e1ac2ff6d444bfb83aa1a32f2fea68f9745c2f4d869e7e984c626fa2451a57410d85
z8921b31999766d01357a254643276f34f9c81bec3ddb4adc43bc1b41b59f95bd4dbd770bf42183
z262f4ed383f161ec887d9765c625a02b271814c4d22b175f381b2dd025b1d6ef505096d019f4f1
z06d02de292a57e76e8705bc58ec06289008250f8879ae3eece7b86f0c3527fb667692023a4b5cf
zd260816a6efe0ac56a5e8d2f9deaab85c2d48839cfbf061dcbc3cff325a05e73f0c847a25140db
zcc72e73f170c641fa9235bed326f66a802fcc49f65c4ee7f4bdd8744575f9aad82f19b8d9885a6
z8d8ea290a74ddb3f40573bbde3388e4b6ef06a2b36e2b8c315c4a945b255e3cec82fd1cb17311f
z8a41d9fe7b07ca973aa99f4a4fffc3529a059ee099f8527a85e7ded01f15463b2adfd62ba17a34
z1928b627cb8ff4def1f1448b6cc74c5ced15d731e990cabafcec94d5ee7bb57be942d8c2af98e3
zfe0171643e34bc59f057165a5f2fae4269f4faeb7888b0706244d5a568eb071550ec60eef7ea3c
z6be510ae700b7f7203db5beffd1e5a78e58643b62435f1a9799cc6bb3e6a5a7958b4a1246fd2dc
z5268d4605f16b5dc0ac0a9357d666f47d4145621b241c8b7a1d662f50d0d76a24f55616e42dce9
zb5d45211c4bf533422e55b0d2c163aa21fb70ce12055875767e39e86e2f950e42660395a7d6dfd
zed89cafd96cca2539f4297924f92f09341ea96a02c999f028ea5805184dcb1bee02b33d472f880
z70c0a3cf6ff59698410ae9d3a549c20b0132ddfdf658da0331696c53d1d8cb9f832e39d8303c9e
zf00d21442b2070bf7edcfacc7b58bb6716ba098dfa917e208ac5a420fc234106c8f4f7b78d99d7
z1dcfd3df60a5a47a1a65ce3999a1e924a918390da6e6cc3f2f74cde50586c0df3c52632e8e115a
z5a6d0fda61a2043eb2e3ec816a60414ddfa73430028b9f690db2ebb34dbe73e5ba65bc5768b43f
z22d291f1f9a4226c5883ac69a76f09a4701137c411cda03edd610403c144d780bd15ccce38a46e
z696c0241b926e950c3467bb5c488348cdbec4a28d077912169ba1b80360cd61683640301305e7f
z8d03d9b8626839aca442542ce195bcaa9a368c79f42d2ca14e7dc416f27317e9b6218b0437c187
z5300361bbab384c82252dd563f5ba0cc99a4e256b23f122588d1218062e4d4a74d5c427b29e615
ze4bd6df351a93224ed31c277a80162d5396e19e294b23e7ef3f4625ef18931e7b9573dbdbab06c
zd5fe2edcbce143099507009a99c6b55741d75af6b76a1305517925d811005bd70cc70d6354d333
za98364430c53da5c85cb1c342b9116caf1e52d9bbeea7aff81abd1ed62faa5bf9819d3b774654f
zbb3f6ff02986ed3afc07b481dffd8759facb634bcbefe4f69345a9553e7c401f3c08d4f66d3039
z07bb615209bc1669693a6b6b76cd1b8d53ce86f2bb0c97eeea2d7fa1e82ce653c70d06d87cec11
z552b76418a931ee816ebd579e69a44eba18a08b2cca95d7eb83d13b318bb3788c2d2a3ccbc0b1d
z86b17d5db93fda78b8200563b52f71f656eab78050a76944478f442e9fbeb5a74f2134ad35c776
z79bcdcdfc3e8d95f0baba37cd739a562c658c566de0ddd22157f62078f9f2913b65d92af6c341b
zb12842411aae428bb3b22f8ad595b512f39274a91c5e9b7e709bd8ab48bdd072b11321da42ee77
z2ec99698e637a74500499ffa1556de7dfa6a99b192e083a59b6540dc81b5c436567856f572f832
zf60e396502b6c369446be4e22bcfc715cdfbbc3de21cb28d09aeab4ac5bf65e59103ef6a67c1a9
zb4a8dafb9c0b0d4beaf8987bf73951174a1bc9f95529e7a2629234738312736badd457990293ee
z60585f1b152563388828e47cf153e3528ea991d45d87dc79c2613fde3b3d10fe6f0284ddc92bf7
z3079cca989a326696ceb2a5da6ee8a9a8500277135c92db3ac49cca872074626050a48bbc21a0f
z6888a3e2d5dc678974c403b2459cb6b0c1427c97ae7891741fc2729927c39f51eb84cdb132d5ff
zf46bea3ddf4da8e5051b54e5c2ebecfd9061cdf4b881723d9f7bb9d33ff81814d3e96f2cd92c11
z1a160cc93c38703af55d59709dc387c9de4cd7323245c33aa3bb7c230eef822faae891c7378433
z5b3198d5335a9ccd216bd55437a69bb30bd243143b8438907aa4fab9441e4ece5717186b5a5af7
zdfdfcee204a07bbf10138c80f89ac5b13e0977e41ab88d723702b46491b9b4477f263d98d7006a
z32e18c81932fb24f29073b4eb4bc9b165949e38320ea6086f183f2d7ec02b7fc4dde5b1917c14d
zf9d19922a8e517fc7558bb7dcf0687b862ed4c6e4b50054c9f0a5623491675defda59fc6d0abca
z32cfdaf7a5960607f92707f0bd5cb1994272acd1a9951aab79d1dd68bb18d9637140d1ebe8df16
zb8778da009f7506672fe0bc04171f35a13645224b607fcacdb2249980ea51a7114e13e6988711b
z53c38e372210140a693a8e7ddfcd44b3917f72097a2ce32d97bfcdc082abb5683f45b434d2b634
ze28b559a0d65f76b1a0d2b1325adbb548dd2f73f1a92b3a02222371360710925299a25068d1c4d
zc64ca91b4dcf34a3b5247e45deeb1241fdd9c51e2ba40a1ab870140f49bb7a5d56737032ac8080
z059ed360663dba93875cf8c3bd117616e155dba0aba001103e013f0c11caef0fa0de17ffe15f42
z1fbb8c91db2371daa131aa3d951ade2ddafdd1e0edc26f0123edd3f71f79e8887352e0f76919f1
zc2b7f84f43ee4ffeae9ceb6d2ac78a7176c2162a0fe1680f78997027915ab00ded8c51117458ad
z041dd19356cc6ec8ff32975a743fd8728c5a378e65c3794537ad7670d7369f0f3639227aa7e042
z8018104c8c823288f45306cc036e6f28e773eb7b85eae54774ffaca9f19d181d82d3877ad66913
z3ea94ba46fbdb3d1b67b07869c4ba7fb49af2af0b31bd467d54ac73f7e7564660e7832937816c8
zbeb883ee7e11680e644d959fc31f4c996ad3de1c5c2a37212e0e8ed8acac199d290de790b0e011
zdcf1f4f870deaaaf8219057fcf8e497fbcb2842dc2f0679baf71f7c01657db5c0f86c8f2f5b419
z961ecfef8a4c971bc9c08a02829d6b5fe62cd860ecaed2b38bd8a63d270d47d87b6278be0082e0
z55f0e65329cb27e918150d6008557b6326f4a234d93c4a5afa28ef8eb0b3a708e8a7539b256433
zebf88b6c2dd3c46cd1b04eacd24230466def29f09b347a7174a67f8916b71461c1c8ee190ae1a6
zb3875f334114c2263d35c1c3f39cf82914b409a3b10b82e7154d503439fea6bbf068d6b41bac3e
zdebd1aa0540b99611df6ff6b50edb80aab5d165d5ca16f0b61426f56d8229361cdc7c21fe91a13
za5a5f84e2024327029417536ba7d6111fbd54c43e1a53081065d5b235a4ff4c0144215321ac8d3
ze8fa1f177d5bf13759daddcba339629f0cc90d239bc59174c6e8d139360deda7ca3fc26b51b47e
zc13d9d1f2dbf1df1d75fa237c7e7a54e37505d82d26949e47e618df2dd5e72a6d0840a13e05d62
z699ccb8f667c6c5c1c2de165918e015b81b6531fd0b6aa5aee2b65abac38357ca2e14d9c06e0ba
zb818c7439b5278e4a81395330e1bc9e429de824ae168ca9d1976f6d149c64b2f6c8b8107a5c656
z7f7b6b2b071e4e41daba999b955ee467ec02b987c0393695f5ee0033f4f9b2b341b6ae32215b00
z48a16e588a3a719b2e48a276cc77be81f9b3763de219437b77c1ede28dab219e050cc1e91caa8e
z385a0463e55352e0fcb29bd2db0bdc49ba93dcb9303b462bfdf5be2a96941bf57f1a5c29088aa8
z6899ad745825cc92d04fadba7af67bcabc6d6f3150d7af2d31a2397a3e431de2463446a93109cf
z15f7ff05c559096a83c9bc5e9e322c05cb988b4a71c5ee7b04b098536427691d1e68617f4498e8
z426911560d557b1d4bc027a5266b45a8fe6e83f69b70565a6ea7440aa51d513765dde33c3863b2
z6ff9934458d0574d966f2e70e6e24cd8986122952cc4be0ba51cb3b475d39ee4264740f082abfe
z743d1ef81c77a316a8d6f66731687c9fe6e42bda6bf6c83adc99c676d6b60af7e21da2d577e8e6
z4cb99efb567577c3712c29d54fc5a3ec3675d80cd4440582e423f480902ab295c44382a135c01b
z91d7e0d3282564261dd92b6a95feccdcc41203bff9221f7ea52e02dfaacf931ee7d62a7b1acc39
zf94deb12b699ca776d4228dd6b9f15bb87c1b0e80d95d9779e8fc86be035cd8c58ae17fc9145cf
zc384c59514db166d394c90f48a129cea9ec334de820ab12f6198de17ff3de188091c76a7a499ee
zfb6a88c040799a0f7a9dbd484b6c00981f19d47a0add4e3d06aca0bacce1f8bb62f7ec3213fe6a
z14f5b869f64c24c73ddea2139ec42d34e6610fe88bf29b6f31ddf406e278a069fe46a43d093e19
zc2c4ad988a5d462fabfbc2059c9ca7ddaccc10330a80e8f25cdcfdb802e60399830a6ebbe38846
z6707ebf2adc85ca9a719b6f685b4f13a60f383447c6509d90091814f3c70887b4c7a0d9184bbef
z22003b975d6256ff52080ff5830b65e949186eca1fa89112effb70a4e510202dffbc4c61bac148
ze128c85d0e0ff3f06052afceaae45da5d1519fd6e338d57e1a4d594703b6b6462f7399c39f3a8a
z51c40dc4f7b51e5c969199d4dfb3f46c2ae538123c89ce176cebb1e422613e8fe3200bbe17c5b7
z1415f96ff36b2d93aeb62d255376c0ddfe0881f436ec45b16e6c0c8502a2e000a781ff2e4543ab
z3d4788c57637a1794a4e4e66e2f1b4f10b4f62a2df2ff60715fb67f679ff02b897b42860e4c225
z30e1af364326e5aad6b7052636b15573fecb1402cd548ddb0fb1bbae66533803010897ace09142
zddaeeee3178bb89e190971c98819f841d5ce6ce72e557484d7a497f41ed675e17104d551b15e53
z45b5a118df3fadf34ff6edfc63a3c1483b979ad9a75ab2e7702521cc20e4609973c572817d8fd7
z0ac0806cc402e6ec783943a4ddeed76fd2807a66472ab3ad0da021a3aa48e8b8f36e83d6012ae4
zb30938c6d649471357eeda2402015d7ffd601f284cba8eec4968c6a93375b1b3b587f97dcc59a4
z0c5bcf5cd1d56099ddfbddfd199a0d6931c1ea2e69b2c7fc32e96cf146cf3110ab3297c3f7d05d
z470892f7517e26576e5392b0c0c85bda880104d0a77e32f72556a0354052eca93e4f35d59f8872
zf2e4db2fad240a024c4935e3ee19e4e3da8f50b5b86547d31983792d497a9d23e62e7922395ee1
z81da96b5d3fc40d9a5b6c76713fb149c2c6811bb20ceb265ffd465a308f6254059360fc0d82e70
z95925b59d4f8a282676ee5ecad79a093e5b17ab9171c39325a3a9849b0a3a184845c1a44b689f2
za29caa84560d9d9a1c713fd6210a568eb8fdd3c91be38f8192413b30d5e42932bf9daebb5b1f36
zb9d89a9dd398c0579c9c8ca7962c6c0c568e0c001fc08808f0286137b858347d2522d9ec346187
z5ea1866f1efd0fd89a6a97015cd3107f33aa05980244e68efa6e00c8e33f3cbce6a2cfefbcce07
zff20237d7af2a9d52ef847b58b59936afa5c045b8a8bea54eb8d823c913aa60e36a91d75737af5
zcdeab64fd51aa48c972570d21cc5b500957dc5822bca47febf8c15bb07e5c0c904250ae2d6d28f
zcf657b33b7a38f13cbd5f978a068516e71461e40f1c99ed447e1a8624cabf5673fe995e894cdb6
z9be93259ea3598ab6a19f735d0e86f5949054aa31f44dbc4d33c5898a215ae583e064f387a14f0
zd4cc14198e840c524364bf22b1202955406106674c03ca27708d9c33ffba41c4a65e1831a4abd8
z4956b30ef833f2c57dbf56b2016bd04440582f21ca7073e33f097ddcb1bc8072dd3572f38f486d
z3924d000d4b4d94de1b45c8fdbb021f53e5bb2f774fa372c622106eef7d13bcaf025582cd3824d
z5e2df72642873f7e976f56e4afe04c08a32dc637a5c83a620e14a5c33acbc56449e56f8bea0ce3
z2d207e608fd86f3803a42a9b1eda0e361750d894efadb85eb81f2a78c992b04f85f24b02bc4be8
z1a6c9495e738555f0b2523edc48a12d975d2ab04c31f4d9c85fd9cfabf63c17360eb23ee00c1dd
z643006d3bb33b7eacfdf08c107a14d43b971f4edf28d70cebb0ec0527037d249934b9129e4bbdb
ze74d92e4b2647b722289ef4eeef7f64c702525b8cd7a449e6d236656080b5c6153ff8bafc399ff
z7d58295eba66d70b76f8f227cb704acda610d4611b91009d6f8c7e1509729d652aa94bf0598097
z02e497583f0264e5d607b835655f1c95d84a97636455ea71ee78daa39c9a5f64f6afc056c5bdf5
z8226f3b9503b7eb96a4a9f9f837d6d53c47fd62372e98aa0ceaf65420579e17a594e81fa158a0b
zf3b7dc13bba5a6a12d0a65b40fe7e2d7842c590a85a12767f3b8b7febfcec6a935659e9869e7e9
zdb4a0f0e93431f62c80c1779808362ff2e0818b035c722f1a79b3e6d328e909112ac09e90b3a79
z1275a8cebba57c0b127b6a484a767c6196f59a543ed7f932839751abc4b8bc692f2b6e0c1b51a0
zb03e51ad18bb480b03dd54dead8cdde1aeff0b0b2d0daca48259a386b9600bb3f518faeb39f2eb
z08bb0a021f0a4686a00221b1199a807f0ea9c59a55ec2f27419d96ced59dbb89c317939c28a4e2
zdc57ad2e22e149c0a71929fe6f17447a8a500e0c8ff9866d4ec242400d709c0c14e10d7e69fa1f
zbce2659c2ca40e2e7966bb769892d607fb02652c7464ada214107fa41c47a57e930d750cb3bcc9
zc7df31873f787bb270da5c5daf09a6513ea20915704b7b310ede9905b5745b65c8f0fd2fa2654c
z3339a7376e237d821ed717e68311993ece3d64d033ab1d132350ddae3d17fb523f014411dad1a5
z4cef5a09905f6800bcd5da546d66b97e8e35f510ce3f47579f80316362ea68708e56f0d086db70
z52dd933baf1ad8772e29f4cd9d261f4af8534335881137e775ebf6627c485920aa598620983480
ze322325994a66fa74d97ee287ec073960e0183206963b23bbcc939457e431ee8ca4943fa1f375f
z4caa1004aaf8637608e072c60ef2e54ec9fee6c5282c42a133630597017b4424f16e2103553043
z99d5113589a0b1e47f3aa32e0a6fb4b9e67c09586f91c25421621f9c8333ec06bee1a7436d6d9f
z1f5e2def3251c81ddf071c99b731ed24bb3b9e22ca8cc9d849627078809e60574a58b80dcc54f1
z97379aa62f920ed006fa43f129f9fbd0f340df439d07d40fbf318ea27517fd55990c880dad7b37
z3ec5c999e3376e5c814b1bc31ebabfd6c742bdd778f2418b83e51f95e94d0047b90d0ed508b535
z35b93517fd1ba7e0e84e51a8d31f61a75129c7fb0c66c661eae7a5ba9d008ba8989987152c539d
z06d26de55236c3bd7c469e0efb7532a0e88db3afd79cd6a32b46e38e06dffeb6a023797a35888d
zc61ce782a970cab7005238e47556832b7a7ef2d056324b497fd5deacdae83e3a5e6d8c61d32106
ze233d9d72c49c038dfd581c9d0c5b9d563450aede9512d1bc44dd1496bea954a5ae1ebeaf05a40
z7ea1b07686ba882cbffc4ff7a2be2cd0f01bc21a855fc8b3cc7e9970d87bd31571e9d9e326d399
z2ab1687cd9c5319d168801e2fcce41df394477530a766af0564779b293c1c810d61b95e161a550
z7ca22c10f7d0a6ec56ab3eb735ab75088ecc0e2c25d16e901deb90e8b8c704a1baff341c583ca9
z9b9c215d2f986ac12afd4b5756d135f3f2a438d446f0aa05928a2d489e19d326119fea59be1a02
zcefe1242ade15f477906855cf3245e93d22dd09e300d1710efb04a532c5d8b1d2904e0e4e21aa5
z0d1cc75d3aae8bc871dcc2cfc15d5b2dc077ea836b943cbe81b8396df5cd34f6e6a868479278c3
z689b5b90204aebb0454db4f4dd3c9cf0fc4a909c4550a0c2035600f588ba5bd061b2da5ba891c4
z2d7ce76ec71c0c58945e15778207e0881eb312cb05e5b037ec4dac7b7ec321ac652acb7d83391b
z24f52b9a68007e4a383bf61d68bfebf09d17550b6b5e68e81830ca395ab1a8bd7fe39890b2b78a
z2b11b62e1e47cef85ff881a553351ba7ff636e6a92964040d138037af822cb8b89400cd9920173
zb11bff2d0acd8115828fe25e5e3a60ceed73deb415d1b29bd64ac3efb8e1b0727bea5af0b08b7f
z7ef3f8000868e6633427854c77e7ce7645cba6fdd7ecfd74407124bdcb3f05ea293fd2bb2c59aa
zb700f0632e3a39a7d837aa07f3aa1cecba0206ab8ecfee7ae565ec59f55d10f7b6e6292b0a12a5
z75b096a174771f7a961bd583296b0818db96d033ae4dcfc964dbdd60db213a6cd5b9bfa19cbfe6
z9c5f94e7562775ae2c556886ccd0f646824073d78589e5461fdaeab9ad6c14112e5a8067d0cbf6
z07af4adc3fd1b176ba91c81a0f7a55ef257947649d875e23d6ba875a3e07bed5d5fd3945822b25
zbcf5852dae2e6199e15b4fb62ec0f5dfd105ec33a87f3fe687a39b15553c45bd04f0dc64ac3f20
z04d825627453bb6df06d9038b52a816188f5c9fcb058e23abf32ca25f18b6e87fe74f7170dca8a
z28deefed0cb14f27561cceaefc29c82ab460ae13c3e2c83670edcd042efa09c338f45eb6b35bf6
z8ebee078c06cfdbefd8710aca2d3ad308aa58aff0397f938427fce489b9f0bf6fac2fb7b37356f
z14883a6830e6151f08ad76a8b4b8592e0c2812b9a16ba89cd56438958586d8aa4b1234603bcd32
z074916c66a7e0a52856faf8ba1b887901fb55594c8d7239f10e9141b0d3adc332aede3a2b16692
zb93139bcce902e9063675dfaef43f63e34338faae80f144c87609edf0e19c99d0b7382bbd3a52f
z4c07f4a78c1989750d49d417b90dec7af65557b8fe879d9d78f1bb11cc91e9a66bae64b158e399
zda45dd13eafd2e5a1b9c29df80d08067e355ce9cfb4b1ea8ff7ac76da5dbd939a62b84ee94cb27
z42f692bf25529fa2e0fe4c44db3c873f794a9fce7ca797c01fdc0b337775b381e73ba191ffaa88
zed9a5f20cb3ba6f28930dcd8281eecf29794d59110d01916879f0fa24592bd076412921891137e
z7f7168de1c158bcd8131c9749ac6a99a35f871eb95c8129b1966109903e8d1c87d436a2a02eaee
zc975bfd6b3029822d44773c9387f21fd999d22e237bc3a91260a51333e2c6ec1f6475652abeed8
za94bd33dfafedaf2991190d757a89f102866cf4f4443afcb423f843d82210d56365513a011aa40
zb688cc0a999af10acc21da096de6a220646c5fd439e2bc4d4abfa861b0faeb756a236d1ea11274
zb869585f5b510db2944850ab7a1f24b57f5d16039f7c110982ab9c67ba0b06b47e9d5a704e247c
z55695b1bcd00f13a20bc0e0dcea0d693263c35efebfe91c9002bbc884d8f36c6da537b9aee344c
z6f2a5e56bfd7476bd69f917dd3b968f54965c0701c39f2de202ce1edb39ed08eaca2ef4db18b10
zb224a75dacbff993d4380b54db2ae4c65758189e281921622349a240d70ef6336177116e0971c1
z4aa1d3b7135054f614c209b2c303b89719796cdcd63e623daca7b4dce3067c6a5de971b97c8cb7
zbb8a77c3dbd3875f2724136c99c7cf8c9995919d4368b794c97f01c569b75d13c5de6d8750fefb
z5862f03ca915b583c630e6b67608ea4e033f1c69ef6c6af9900e573cfd038e6b75a1a72894ea6a
z2a99f95aaafd48e983fa74f776e05654889d85462ca59a909e0b42bd958596f08f0647cbd6874d
zd7a604704b81a87effadec4b9e5172ceda57ae28d8986286e1c8b7e82e9ec3bd8d18445dcca207
ze8ad498fe8f541d94df13d2c2e617575c47a5739b810d1d67c310f230b1e3577e0f45dbe3ca636
zd67447e57d891fe9ac19cda1e97199074083283ea19c61ae4a9a6975e1b72ceac52d8693bf58db
z646cc5fed0b8bdf7a04de3ed61faa2dfb2f690f80b82f3eec0623d1540a965637bcb512b567d32
zb14eb0128751e935a2992178bae9119b2b65f7a580d4d4f05cc575ad15a86dd1d78da210065448
z890bebe1a76f40890d70924b53f742f2f6489e0156784cd121bad457a8e832e2127eeeda120929
z3eb2287513900dc258bf787f3be23b3fa5840327e083b901618954047483fe36fec5478013f4df
z62a962f0d4292451d8c2c531dbd1830b252eca118128d229d7468b0af2a292f8e2a2c13affce2c
zd638993ecfae36fdc4df45d53426dd0b2e3903cf193e31fda594e19608e06a010c2768e4811672
z78ad787ac550e3da477c4283ec20758238fafe4c6ba7d6d6c4411549531e0cd27072cc871bd10e
z557f9d3f4de0bfd62cd46fd7812ba72e3d98cc7883a0b73741e19e0cb670c25b95fa889105fcb3
z9ecbcc058b6ec7aecd2ae2a03cf25982841ca19c8177013c813d68d4537904d34570ba0bd224d4
zf11dca4a45a1638f49df7f5a917709458a411e0513576f9eed1a1d17dc3906da3d8d6e02096e5a
zb6c4cda99659163ae744f07d82cedad5f315bf8ea08a0151c325e0d46c14095ec627c9b15ba445
z09f912d313aa4fa022fa6558e12f93b94b8e9a82a49218b8d03ce586fbcd4cdca76037a50e16b9
zfe6d8876d0cf48f49a47933fd9bc71ae9c9399bddac739d23d28af4d7f0c76f809bf9f8f1059c8
zcb570dc50f3b348e855443bfd74dca120aaf10848bee1946b01ba5ecaab2bdb6e96dbf61eb4358
z42352c0c3cde3e3f3ba1e4edfc8197c292e5c5a93882edb07f18ae8028b5dd571bdff6c1624371
z4bedda9fe0b090d768d1fc5cb930e4017ec9ea6f35b0fb2669f5d5e02406ff083c06f20ae5b8f7
z3481cf5e2ba7ad2ce40c72b23bec4c80c9384136e8b6e32b6cbdf3fb85db4d5890697c4572aee0
z5352853c4f300b237c205e58f1cd74962dd6a778d35bb30e08f0da628abcb980ffae904f32dc0f
z64ebf4dd2fce492d841fda78d5150f392956cd97c74d6ca4d9aef1ef62062ec14904bb550d756a
z6053b0f3fcc334a24b84036d5e6627f79eb7dc1837b7847c6769be3d5a030084e284dc0f9c97ca
zaa9e61da298773d2d9bdc0acb0aba2d6820ff7ffb588c2f7c737dcef455defaeb451ace7966a76
z8401c3000e6813b1a43c6f46a167dc1136047d1bb255c1992462772d66b860d277f0df4de41da2
z52d97aab8462b439d41f1545ca0f1fd4be3dd13b6ff1ca33be23418bff677ff25975dfb277516e
zfd5671720c62ce8f8569c9707ac21603fa8c4456cbccbca1e9426f84c37d19d37a160a071216ba
z3706e63f727583b9b007e18533789f27dbcbd1ac3f6a75b48913c0b9d495251afc6deed1811673
z127b26fe26bac73566636806b219aa097ac8a7df0c7c49b7cd3c873b1812a777095d5f45421047
z25e50e7015d4416c604b6b268a686eb14afbf3917b264514f6ffe36174ab7a55f1bee38078e463
zf60d2369b083a5e9a2410662134103fcd1a491477ac5120c684c93ef6797a107096f179dd7259f
z5b8add5aedf8141922c119ea2e6649b5e05a01e328bdbeb24097a87d9f1ba85301685273b7246d
za38a1d2eb59ecd1e2964d821ea76fe25cb694ef25d1d1457712035f7e4118b6821b34da9a45289
z5b131bec6a267b4332d80c886dff214fc2fd0ffe8a16b7747403bea1a48ed9c943775753a3fb7e
za6a94a0dbc690ae1e029c206ee0abec7a5120f395d6f778dc2da34623b352b25aca7a52eddb9e3
zbb18b222aea494fac96aade28da9c43c3b60afb65b479d2f7c0ecd3c360385e6793af85e59bd02
za18df219c13dcca319c81e7117a96edf01c6eda59c40c9a8ea6d913549adb76bfbb50e146489ee
z469bbcaaa810e2b9aa08a4a42e2e04c103bbe5bd24841f2b69a7c87a70771bb1e76dd3810d086d
z450ac7e600c13fa86e24b598e064dd8e5c9e299d4a32ae0c80ebcb4364b712852f9ea15707ae6e
zfae05dc35b147802d3b711a9bfc1a2d1738322e267f4281ed002c5020e249aed17a5f4ec0a2357
z8c632f8a32eb840f8c5df6248bc86839673e4c36545da71e5002ee9ce930d2ffdc995946f79861
z1f83221e4c6b948539cc3e7c969f2528d26e4abcba218cd6d3eaf62a66521df67d0a916b09333f
z9f09f7dfa3e71ff1992c1d46823fb80691f3159f2f87bb1c12d47ecd6b5179c94d4ca668aa0978
zd5b648057875a6d37e3a34a96136f02e28df2befc7f29711fac06c04c1a60e2b57044424cb03bf
zda31447d31a39fa34f9171d3408151b107cf1dd9366772c2839f3827698338e24858c0522d46b8
ze82f74ed65e33e9ce4142beab5310c61d65dd0fe7667a6ac8777294e6e04529eb6db29a7d9e096
zd651ffde9360bc89da24ce4f6719922eb972bfd7c59855f522bb695cc2df642478ebb2ae6d2c29
zc9bdbdab340bf4dec8c50e4a5145d3253e0ca71dd2695ffbc68c61919c7d193c0215eb82deb2e8
z717d93fc5860569ffcf888cb1997a856fd8d7554f5db7003eab797c68a7ff2306dfcf2e70df82f
zf9f7326a5e46d7f3b7a21270a884030e21df59ccaf0f608443d834f46794c86e1f75114564f474
z712d14f2d9ed282382bc1b54633fadf4f685b5da84e039ebcdc9f3e5edf18739b8741726322ca9
ze02e326fc80e84a05870f184deded90b7a7e6033480a68f148d946877201766306f9aa1a66c4e4
z0c257b0ac1e3cac83e7dc3226bf73d71bb2405c97a186c32ade6cf58211c5f1ceeb505990a04f5
z8924734ef30abe4721f9c25a5c720d721db4695cea39d9eae58aab029b0d9c7efdfa2b6e83f0a6
zdc7fa156f0e1a5c7b2d909ce68770935cab1dd245757856df250052a76b29841e6774f55f7ceb9
zebedd42b5de50e35ec3161ce93e9d4b6902b99405b5287b7e8f773aaf1e746f6971bf68d76502b
zf7e9440b1acc283ecc4134118a6a06e3a74e0140b527833c347cb8f744b184750c50b805547aff
z71404967798cd7a1366aa1f285331314f1c38140d38ac8eb4e7f2876b728a876bf9833b6da9190
ze521738926556bdd5800fb393eac413296ba26cd71fe26dfbf9ae0d643112af62bc45044debaf1
z8f2ed6e2f184b76327cb9100a45a9f4e28284ffcfa549fe3de72dd9f9978f49b30a9a677da79be
zf74023403b172c1dfa26cfcac8c6378deb927cc41817409df89d7a1fd1b14720bca4c56952dbe2
zae581ce8a511cb830bbf0c4300d707ed4b5c26231600e6f223848252839a4fd541556f596e69ec
z57d536ab4a08c42eb7529ee3407d925a23b5c98dfa93d79f4974f54dd2333ab7860783693e4078
z64f28d2ec0be4f0cc45d80810a08c4ec508a8248a407a1c1cebd0ac5cdc99e26a9231778bd49b4
z34de483bdb13f7019abd0cdabd18f83898b965baa98f8806343a0513e0269bb05c37791f1bdc91
zdd7067237c1920fa49c590dea488d58434f603cae14c6cf903b6aeacd42003ff90a4a0f961c4f6
z604c85c2c224c40b6847383642eabe044bcb69708726c58665da692535c27b632b80734ea90c86
ze918ca267857f55a9806111177e2940ea91748d9141ec20cec5c98250123eba2370812bf71cda3
zc90d9517b05d0d679f1345466f2b7b9f5ececb09765c0c96d623d37985d86473a1dc428b2d1a46
zbe6d40fb22fcf6fe64a6eb87f77ec1e1b8ed94b49c112edc8bf300172df4e1c7cf5654eec5bf34
zefc7a559de1f6c8a88ce6da7f780b5c97bc8ad02f3d02fc06da6d07e8d03927b4dbaa4f171917a
z9653daa31d9ef5c9cfc09bebf22681285fc9e153ed4c136b7851895e2b7ac0b22e078b3bb80a73
z4c4f7e76db264ce3a9c9594b6b142c33f0d49484ae8db65e570c1cb43aacdbcecec727377b5101
z4c5b873ed16c69312e5ab4ecb1e81e098569794f452d5c3eef3ed4db5488778d11d3fe20e2c7b8
za65b1762ce86afb21cdb942b28e821d13b2b802f28bb2aa843b57f6770c34b2c8c705694da2d10
zbd5fa9c201af39597e921be967290387ad02cbf43a40ccbba3a69f6f9bdbbf84760d9983f5d686
z21af7bb0fea1f2f72f31a2623ea82ebf637026b3db8260cc9c48ac627a57aae6668884a5cc45c8
z7871fe55dfa3a0eadb640263e3488aa3ca315ffd358e2fd44fb8ae0646d08783850b3c84311ce4
za2dc85010d0c3e127a828ffc8eb48856835f99bedc30787d9e32f93025b080f3262634a6ec1c4b
zf201b9acbedf9cc68e131c3f4023c805ef43b62ba2ab300736a48cc4cd4ad2c3d57bbe437addc6
z1d607ac1a1226ec880346b80e505b83852893e7f04a106d6a87eef62c249ecd2526752f90c9678
z0e6a71979c26b237c88d38b7b238e0bddd16d04ab187df919918544d1b6285387895e938bdfd04
z8a8b82af00b6e79d7e30ccf8c9c961543aaf48f7459ca5d017f8ccaf4c1149aca79c5900f216ee
z502519af6b0bdb932cdbcab6f6b70f76a3d90814747cb7bd2d494369a47db23e5a4b92655275f1
za10d97ab93989848c856348c2e9d5791d72b772e9ee3e99f68dd62547a351c750f90a1582ae550
z20afb360b9fbd793353b82f4b2315b1e4b5857ea1ee1fefd505f0dc6f722ca30b7361fc845aa44
ze8e9540daed7db31c09d73cb41d420ae452e52b5f1b07ae566bd9486f1f03ee5e7674817303c1d
za908dfd232e183be25bfd9f10ea53cfd9d2c00c687f2c08347239581a0ef230f140fe7159ade99
z3fb812cf9cba90e67c75f9cdbddafd98e8fda4176623395cf47b968955cc0ac4de956757936c61
zc447eedf7ad1482d34e29fc76f249c536d8dd35066928227634cbdc49ec5065cd7c6ae2f474a2f
zc8ec70ba9d64f2ce3cc61f4e2efd1e431f0d862abace1d9d940dd769a530e1f7742bc74314e8a7
zebf6b4eff92fcaa4cc4e46dc3d21b0cda270a7494ed196bd1f7a97a273577dee6ecb21a26ad7fe
z523a137850ec42a528ac539c2da74cc8d2266a0ce17417ab22b1282f28e08d82a29e99a33893cc
zf25b203ebaccf9c5f01782ce015fdbd14cd488b347377d957a73b065f1f9858c02ea4d62fce7b2
z5b1d1feaa0695625072917a64d2dcc5ef313fbbb7729e561e2b9a01cb7b3c7f7a97aae7179e6e2
z644b80d662a0d1f3b7887cfd241cee1e2544c05777c2e0567f3f74b0245acf8c014e0bc49efa35
z761218723f5fe675be194c9b295c72907854b3cce04a239a5332ef16c43e5bd62d09f1e89f2633
z76275e9e056535c62be21e22c2ab1a3dfb14c8edec6bd13c58633d6df8e80c16b7017775ff1aa3
z363767aa9b154a84f7bd391c5419b31f78e25ec3164e93379666164ce01ba2cb5c134697fff898
zb700d4d47d5656b6b1ffd56fcd3496ad625b103a3f2a224c7b921839aa537f8b49808411b6b3e3
z858e1c180587de3efae475ea6559cc7c046c7708b846a7fb980a676d27da5b37609addb48d950e
zc12886c420ba1caac4bfec5b38bcedbe3f2eb12c5e8779b06ddeb38a8d7b2b4aee62dd418a5877
zadbd8f5c8de926823af7488a7193d246b45b3608abec86da1190212eda8c88eef29ab492cce38b
zb6f3d0c265699f66565712614ef77a668868937b1dadfb5f692346daa372fb8bad194916f149e5
z7b5cce3031c239e1416267661765b5efcb13ad32ee84b36a677046ed6401d2c6f14c3015bbdfbf
z120ba3d8a9358daf9f8f56526645fe67814a8a1c2a29af1f54b33156e4ee97cd58ecac89c02af4
z3e2026ec4fbc76adee76cd09f9e1ef585bdde33e4abcb0b24f6b50c35829606d1f0dfa78277384
ze09babcdd4b28ce200e26a2a1201860f5e0912021526de26da2c43876962ed4f8b71bd4b3ffde7
z4bab18d92483e0c5a445e92d5e4b1657cc0cc9d9d8c4c7628675be05820f7477191240f6024b3b
zcce08c339289bf512feebf8aa93a0dae85cc80d84863f2248ad41c55e5cb9715f94b11750d88ec
zcf70ab72b592326c8cd6403363341fb5aba56b5ae427dadb8661a7fb39244f68f9e953c872ed42
z4a91b4372d067cdf2192b6d705a270c3208a2ef12b1474d538f6aedaf22efe6125cc4cd217d0fc
z798ec74cd7233157aac9e3c6e7ae2fdbdfcb2d6a284e160e060a0aa4134e61c40ee2c144be3e1b
z3665ac21661a9039105468d4df7bdfc5c5715d21d65b3e9dce3ecd4dcfee120d013935829a7c4b
z4b4a6a96fa98103e3fa3107154b7a1b886a3a344b8f75d4f2135bac6e7caef0f2746d2c25cb901
zf38933c2ac09e0f575cfe1f78dc930cba6bab6c973a380b38412ee062a16d52b8c17b393f389f4
z9107901aa65f9493beabfe98883788b77b9cd150133e6044f7f5bc76a02d1f0f19c7c30dca8192
z26398603ff1ecaa66e6ffe1094f7ee641fcd75bbfaa431c6517b9cfb443a960eececc0eb823fbe
z6a14ed62f3d0f565503d72c0194b06d36a15a9b25a7b063ef36cff4eb8abea4eef48e915081510
ze7dc69fac8f9929385f10133f80b58852fc461f9a2938b069fab3ed4a0762ed22bd59baa159d15
zc41ca00047cf4d44ae2ce9a9788735cd521bd330b8c9cd89273aa2c4ecbdb7cd13647ad0c87741
z3958498ba70cb981184d3b8817961718b8680a7966362d0aed3d2b3d55cfec582448a310fd3c4e
zba691de0e146b833e2509bd5e96d74cc685f98d2bd0422d6195fc39869002a89cf783cde6e6750
z75d10eddaf7e03194264cb95d4caa05cf22bac9a9b57b276ed037113ce79424a9c8991e7ee155a
z6bb4c8c7b303cb48b7a5ecd2997aa03fe7e33c01fe8d937a0208616adf974c2fd1edfd544fb3ce
z6d91d520bf353574b6c7288e3e158cbb83ed51dafd5b1f9164087ea06ed6fffc718d22d54f7613
zceb0a9579eb2cc20178edb1cb6c8ea765dee2c072cc3ea7c40c1d1156554d8c6f03dc37fc58e71
z2f4ce99cc8da00fa82b17ad24f3831d3da763df11f97ada19edaff9f40a9b2670f8681ca1018a1
zdd82982b4c427bbcf498d0093b407f32aa78c27ec3cc068060d15f25476f03cc4e11deef0d323a
z0faa6d1ab15e533cb7d9f16db95b89f9c929ef67b2a0fef8165e6e32ffd791c740418b559ca13d
z7dc4c2560183ed7a7b8d9b25d079f7f82baa8af60d331844df70bc2cf7227f9438ef55ca38eec2
zebda1b4d17f9a5dfeaaf875d2142b96f76aecdd4572c28317efb52ef23780389b5ac3dcbf3fa6a
z1c1872deed902d173cc71bac7202f30c14927831307532597e2a97c26b1e3beb992de92b82fc62
zfe26a34bbcc09878979fd510cb79c4a9fd7cd90dda331d0c56cbee0f3d04bcc53957febf76ebcc
z2c1664fa10bb28ca7d3be55ce37edc77e5904f5122d51ce55d3470786484f65e4b0228b1268412
zbc7d4a38000178c90784e86a01785f6e24157d1047f88db5e93f3ead0cc5327c3fc458517c8509
z4c19d2c333ea780de1cd7c0d1c084f6a970d3af493df7bd33cdf27e0f88b880e4c361257540d02
z3bf753581ac2aa7dd9924670a6b9eae64455cc76b30e350ae96e0cb21dd4814bd80802e4da7116
zc0a45d6755bb6a801f436157f5a4aae1696dee7ea92d1ac664f181ebfbf502d3c3f9ed2598402f
z606a268d47e2ab8ed8b939a48911f0289cc4f22b04264f42a17fc18b9a42069b57f3dabff16113
zb930512508ea5306789f992835f3dc78dab029578472a75415978257ca1613fd4774523817e8dd
z6f1bac9b3afa3beb9c4bf1117e0db19be9660f2c4288d158e96387232007fcf32daed4de98de2a
z6ac1a66f31bbf745786754bf95a7dd7e4a2e24e680e4fad05c95a53c16fdd476bd1b6fcc5d16fd
z5d40bf276ea72b084de1511f770bd58036fffe336949f9ea063e9ecbc66d4df0b034cec4c2e5c9
z1b6df0b8d092634babcb0dc03b8d095e32fd78ffa3094fe72ee800d4c8cf29d4f1fdd6983fe5f8
zb7c6f234668d94370869d4a70a378ecd9f9ae32469172f50fc02df637cc948fb5fba829a40aba1
z858d554edafc8a43a9da772dfd17d1f31c78dab13e05aa18dedbe7e301e6e5b8c97e3e89959e63
z0d18d47b1e55b60c50e7f4100a3294fb03bbcc783c86f18f7df37c3071046bab4cdcb480a8b32d
z4b3d17e29112bea3b0eb745d1d2ade7b3be556c0996a2e10b47bfa67a915a58324a4415c360334
zeeb0ebcbf8253edb5dd6f6eb84982c2fae1cdd46e2d1c2e95ecbe0328b3744c94df49fc7b7060c
z601a637860810a69be5b2e746869e9893fcadac7ebe64635344857d9a514a22492a05823309428
zb408293f7ad0df8f827f2836862cda49f1548688d4b2d004dd6893b7821a63b2d265c59dade6fe
z8ee788ac5e2ab3dca9b63bff31fa71955be434738ef6a53462c6835c189f4681256cd7f1664938
ze458321ea0e97bc40a1e4419c58dcdff3ea046507c629c8b0cffe6c90f238d98296b86424f5bc6
z80ad1d4c35a199fe244e66afca23b1ee7a490611321554d6b99b9bc5f8d54c13d0af88dc5810b7
z7af3a276b05383b42e904bc378803b28c8fe6bfd0366d9561291a9689ac056610f8ba1e6d92b41
z3f82f7c094ee6bd20771633be848021bdf7487f024fcc6a61d6f32e9dcbb522c240aa75aa8fa66
z88aff5e4e8628958240eb95494f1254a80c82acc6ce8354e9b40e6d31a518a8c2faf6bf9fa43f8
z300f370cfa0873ed7644a193ad6bf8eb5a9b6d717e1c43c137cc7be47122250d77c4dc9b34cd7b
z697f11c80456e141c17cd2ec260b28159eeda60a1dc0383de0941608a9ec1407a3a868d7cf861c
z47a819cca709edafce522516d652c084e2744bc14915a3fbe53106d8ba0ab4f30fdd3848138795
za49a7aafd680a67c2987016ab8090bb869b710d1d68382246035538781a5e9827dd390df62d044
z6c30054ea0cd072f8d17173ec904e1d786b1b0535659b56ddd1e9c3cba70271ced0fef3f320ba6
z0e0529416bf167e1d361fa7651501654c0e2e93c9e0989104f4b38dfe27cc7a613b3fe514122c3
z14e5335cb39023af96aaa5c0ab46f2fb3323ade7277822d2c0ae72a4e4c3ef93d2853939612fa4
zc61f1fab5efc1f0f12727ee093b2061d0e5089ce6e690ac595d5c70acd46499dd751fc96772b0b
zd61d51d0e05870e8e066275a668637fd0022694aa19d65ef4b823665054ad83626942d654d080d
z56cca3fbcd28dd3d4869da7c4341402e7d22988869a6d0bb316a6ecb80ae5f1dd51b5b5f782d29
zda30f6eb26dd7a3713157dceb9e62fa1107c2a764c01ea30165a5a312557f79a568e73566f9677
z71fe49dce0e10c61b12100817d6efafc7e559063b636d6000af4cac6ae9f6fb0cc1046ab322359
z583804eec945e6967ae326766bb207e25ae7bbac5defff8a5162c1c69d20767d2e5ffff73ede1e
zeed5933c1229f5c8bc298ab6eb695a733ea55f1f6720bed6799966eb5babc380f74668c3eba5e3
z41e5de0d9112bd17a04c0424cd6e85d951c66d88c593a7897977e266cfb56d8d80f2f37e3670bb
z41df151d6b25b987e03d29c2a2de14b2a0d0a9beb1e6e6a7af3291e5ca7e20061d205b76f2053f
z45a0a10a93b44aec7109a9443f00683ac223516f2a2f9304c0c81b0a1f4ab373be3a1f453cde20
z351f03e09772502b22c255dcc28b7aec8a1aed3948f48ce61be4591e514908336fa986ef7dcd71
zba3debf7d4a659e0df54611b6114ac3dea8ea522efa2d11a34bfcef84eafb794d2f67fae2cf3af
zee551d69b0baeda2a0e64f8e8a47cb6ef07de7772331f6ed92a0e133a11686f7afd1ed58d0a36e
zf5549c7f1ef3abe0564e0cac9a4b6c7b794d05418ec24e950d7bf2641ac8fb438d850acb74f9e4
z61f246380f6a840e64e0382b94b254121f8e0606b55bcb385b8dd9c39aaf3316f1b1cd66254816
zb60ead8681da3e12fc655f77ef9e760fbdac49902ffe1c45e93d5d8dd61e67ae3b21054b2e640e
z74b088daf75b1b56cf2272cd15fe40a7d97d43281a7203721c99cad96a92d0820a8d2a580703e5
zc3bb8ea235dbe51bd340fdcf9093113cb9ba9de220509e4e95b9e37ac0d249847a617270f42c96
z609c2054d3a7e396fe3a8ce763654f9e9c6b6666052d9fadd1e2d89cef946e6746bb6e86319120
z6555bd65fbb7b1a38766997296416c803c3b3baab494865f2238dccff9c8a676a052d787dfd65f
z214faf5aa9b0e996249aa10817f5df8ec5e21b9a3e7edb1c4943efff03070a3cf5143ca5f3a552
z6d11ab204a49333203849eb8235ee996e6301a603ff0f2b7122d794a3bd644a8d1777474783d8f
z5d572c10290206200d965072735a04f2105d358f1d4918cd11414e6016879e9a4e46866c5b781c
z095758093259a156b3bb6abd840f1496f679a6e88ef97d3d19c9d47f9d455a11525370892ee5b9
za1b34d2a7de229149ce98bb06128c4f1a54739fd6e13f8bb9dcade791b54b52523f01cb433a099
z6017064b4c30caf3eb3123b53b1c8b53c98d2eee37a173c2820f9f5a07ac1db128bb5d59b44dae
z4f9bdd7719afe64671ba1fc5e623b01bb645b2f8f63cfe3c11f324ecf34b99aa6b9aaba72f1268
zcf887ac8e0533a51e5d62a7a342fb9043648047375fd3e0d062da347b26326110581bc245db396
z87e016bec394b7f8fdd69bbbdfd9042f00f9da0d2de3ded464af52b08c173fefcbdfcd331745cb
z3f3320cd19fa1427caa0113c193d88a6c68d21741b2f2c00c28c1e4f386798d7dcfdd8cfc58a07
z3d6bf3117a6cf6e8534d32661150afb9b691de87550ec8fc0e080118b7bc4278a7eaf0fa9317b5
z8aed19859aeac281f784171f77f630fc80cc387d46153e939070b0e0078156ced390aca5aaa6e2
z38145b6381ef440ecef7b8c49a7eb1ad54b6c1db896350ca98ced8f5560a265319f802eaa045ed
z5015c7eb1f5eadaa99617d44ce954afe5ad7b112f07c39f294e4629226cd99a0217fb9fb12d875
z1acf18aa2e369bec6cd4fd1251ab65e184ace98610465d97cfb78307af60888c1330da9fb54260
z6d912bf58aa81e90e1d9cf71b3bee348664b3026bd1bbeddce61bf48c285023f45118b2bacc81a
z5f02ce261e0d8bc7da413a69c092dbd40062a4612f93435498ffb28ae2b5ed149953d960ba6b30
zf7a3dc73d2569b675b46f9b4624c3062e26d4516e12d181a75ce3af915c5e353d095d520b72f3b
z758271c1c4637057d58b19be9e37b1efd8c98f615b129a35540a89b71e4577ec73caf1e0cf60b4
zbae98ac09618e8492ec12e5da6334b72dbb8038be9b9b856ba788178d9704f9ad4c46317702c14
zf782a420c7443378162641a647456fb5d40a5237cb5a9e0446ff925d478ce499c1e572f8a0d372
zee8e0133d2981b9535466aa12672ec88f9fdfa52ca280199adbf28d2c9492dac19a2178801b66f
z80f5d1fccdec165350ca95caff15ad707cd3364466edb5027d2fe69b3f7379326dc60158c97632
zfb0677a5ebc5b098b8c420f9413c9d74981eff3b635857fa19db9b3dff0835344e71d14a474ab1
z7697b95ccd91cb510fc663eaa6387dbbb83d9eb1d36101d445ed0b008805c41ccb9a43cbe0e076
zed03af9cba523c4ba09e6ff0c7df3c54c8c2c533f614fe8468c5d7c947bfbba934e7d31805717f
z1c329abca4578b1a438f248e36b69a30d302285e62b8667d2aa739ea1d8df4dba2b687123f7d68
z56197977a3282bf11f89a3731a943e110b618b360d70c53eddcda27e24449f79156788cc7829c5
za537c62fcf6ef56755b58803ed641a375e913110f9af918faa009ebe0676d17c59b9b224fa14ff
zc0a598c035655c8fd612a2161a9ecf3c7de2d4dd8dd8f265335a62454c37d691bdfddc46a23565
ze3d36618994550bf9ed6ade668b00c4d847c19699850ca0571c1ba076894b44795e653c0e7ad39
z8092ce746015612d05fac806f8d09c26da1995008a9ffc0acf2da23a118617c4a527cd2aaee2ef
zbd6c8af3c8a4c24257cf4fa4197ecb8c5b4f842fc4b881e36f54712b6157ffab766c8ff4eca527
zdac8fac2fc9da3463b9ab219b0891c936b753e51fa2c408a1b7d1b1ccea947f95cd968dba6d47f
zd17e69878762d937cbd2ad76bcfd1c6a9e10c0ffc7f2579ebf4fcebb0a0e25e209bf22ab045c41
z4280845a558a77debe543ca4850916206e01f2c85cc6fe7e7f06ab0a8ab959516005c7b25f1d6e
zac530f4f5bd5410d0f4ab04371fc15353b042561f5cd4a9a2355fdf9c97ef8e8f26f7927e6d3c8
z672e73cf5acf7e082b532253b5c87e0c071ccace2e2c90d5ed4191066fbd069161df46144f344f
zc84583473fbac8d1af382b4485bfd4239a8d6f14c0134328a50a7d6b2b5e4c60610d5cd6085705
z75a11cb710f90ab9f4ca2251fbdd2320c9ee64ab46d79d5ee03305295691b2fb80f87f8cc48654
z0589dbbc8e17c22eeddf2ae4e47cf26af8e36d5cc2e6dbddb3afc1229e73674ff26050da57df53
zb7c8fc49a2d9b62fa03aca9cb1c9dadf883854e55ae1f983cdc127c758f663eafc6bbd448842a7
z14e027681cbc911b5eb7aa812b3e6162a5eeae5aa072fe7347f6248178fb1edd73464c0377db4e
zcf33d15a9f4d4c05b9fdf87e1fe870fc1e1daf078554de8ef8128a34a02bd5973ef39471ed9503
z2aec5e4f2c63ed2703e4a99f6c25db3590f07e335737dd0c0462766507c6b0c9e30032b55b4c19
z697f5c41670129ab63dd7619ddb2cf4cb57feebcb5c702d726cd87d83edb5b5b681b82936f61f9
z6422f037c04af820ddae69c951e4bf85faba076837c51bc9b93db5c2d33c67e69dc4594101eb3c
z999f78647a69dc5d6fd0c4a3a7dda24f32b4c38b4b555f9320bc86cc045634ae5a61fa2b7563dd
z6eefd120331da69fb7dc6d3f894a1434c0fac2969b5b58fb8da810dd65979bbe2077c35578fea2
zf5634315d9004eb9475f631edcac22ffdba2853b1d3396168394eae4f2037e0733cb7df12d823b
z48a4385755b7e5d721d5a2a00ed361b1a986768bfdb910a850b859afc2630069a18149f529804c
z87e440e5684bb4b3bddc1c386d70c58337147b882d3ad43ec8724fe98a6f0f051d38ee0591ba6e
zfbea3ec319509f95bf0d594398c7b90accf7a3680672709b3fb3cebedd5d1d9d26cd7ec65d0a4d
z6576eaaa0441193e57f9b863b8aa57e2778a8504ee76e6de93a863ab5401c18191d12f00825fc9
z863369ea2e612163030d537d9bcb8536e285ac1b493138a980890f282cc304377f349b88aeaeee
zcf33d0f09e8abeff3cf808eb8c884f6d335630dd81283025cf9ebbfca615c92de15eb5a9c34d0a
zfec46ac049c592d6599dcbbc51c824a92be3955db0a83c285c6dcc00c7416e5b77995ecd3c572e
z7434a0d797c9ba186e144fe00e4def7f55a80b2f550e13d4f91f87e4ce362ad6c77cbd8e9103a0
z3fd2f29b7fca7206f4ee7195c265b3b3066228b3e6d58062f6cbfb1a322783dfbdd01d60d38e6e
z4383100eadbe983c5f1dab352ca68ce67dd511931b477008e74a0bcdc9dbee251355176b12e34b
z9f50fd998d2a5cce9250b77eb31bc8bc1dc5f666e727dc3f76f84ebe017e5285734dd08978fe44
z335e049b92d69217ba320426dde8e425ed6be9122c79019dca0d08970c0c95b23bf312d4f2aacb
z50f3b77cfe856d51f54a37f9ead4abed51a32b972c189d5f15887eb9833d7a5e14889c14d82d09
z8b8ee07ce853b1486d9585cb54d5953d5a8db816e01c5d800437f236c6f65fbff64a9e4fc5699c
z4b0faa82b7fce6fc1c060ecc3e96706eadbe39f8bfcaf75aac6d4f28eed40a9dc3c852c8695452
zaecd5038153cda887e5f6edae2fdfd7b08f0d59ab78b0a0427e674256f02894d79b33027c23c4e
zaf851acee36c1f8110e9da7b4daff2a3409909fea60f59f17070dcf43569d87bf9e036e6fa3a4e
zbab4e13fbfdcaf7d16b713d141cd35cbcc49f124e2bc182315969ee16a75f2a46c35b3d021b45f
zb005573ebeb941d44b44a5767df3fb9b79a58c0466c05404d608f5a2a75eded907b4c66524d8de
ze2b61c771a28c5ee1e6e68b02f74062f277167ebc738928eb7619a775b20bcd2bdd5eb81178bb6
zcefd1a5e32f6e1123c4f5e7d7188c55053154e6b731562c2fa3af48ceb419b108a0c87244461ea
z2948c361774fac93bd8e558a401de4e7ffd534c5c079b506eb8b006360b0950ddca41bffb39582
z6f8df83e3a733519c9cceabd6a54c6f360f126b20ef5e90c58120b1429ffdae061b38e5f73b5be
z8e8a8de69cd7fbed3b27806558a86b4acf43d4ad68f37e5f4b7d375ad3316b555c5f1fd22dc304
z92370efcfdc30cdf11024027c63297b3f41f1495ef2f03c4e8c642312801f36bff39ec1963c5a2
zd0a0bd4e320ab72e2093a769067fa6c4ba723309563d1d1fb966a85a774e9abbb4b79d26092399
zd7b148032819f84bc44b8e36c1223fa3a0c62ef60abd92cce24819c371cdca3c88c9beba7308d7
z3fc256e12318266471b2f7b32f5dda9ae685ba4af88e94bcfb6e48ba770eb36c97bd4d4bf35809
z1a815b6ec659abc32c54eb0be0f2a1785ee3854a228243babdedc100f59356dc30258361e40795
z52111e2eab29f30a44af25c9af07a4ec144b7a505cfbe0310fae511b79614f5b21353917698999
zc4130a11d90775fb9065b6b0c83591b868d51cc8b7ec01015c928d06628e3f07bca97bf6dd48e7
z7562d85899d78a6de6db6689df8b7716515b13d6e8b47a9904f835608e95643c43e276301bd982
z091d67b436d43a3402f18d13320715511cea51b44911cab02b696c3163e775769d08484b2c43db
zcdbf055474cb7ab8883a0bbebbb9913bea40ccb441068f9574de7791bec9daef75f7221a6f4481
zb0912cbd7fa5288b005dddc1d5e1c7b63a438dd1bfd42a71950ce1cb71bd7d5a927ed840a19fbc
z9e8c1253c3b0dfd4d86c5924dc5ab2a296337a34e342401d966d618b6cef61df74b8113d2e8436
za480dd41dc25dfdbd8b953d98b2107e72ca72c37a322254e1328ec5ce329b931f79d8afedd8d06
z6cac2246f0314db1e5502d4b5fd2045bd4f032b215431c54e711abc5eb84f909fa58d340b3accc
z6fe18548a5fe82647cf1c166d32471a73710d4caff2268c581d98f7e080ba89875a3fb80e29f5e
z26515aeb45927977dc97919fc3f951a911b5c397c379d795b2810972a434c09e176415bb5d3f20
zc50699ab64f59135c3e8586985aeda029eb8a11a6ff4eca8534900145da7605868b53ffd346fb9
z511c7af1e3094b2583d1998d41a8e2f9799bdf69e86a26eee8ce2c3c893615d10825f7fbb9d53b
ze91f5e1879a344ea1f1adc67671c8326481d3e43b6a7ac62d7a9b97928995f178521a2e3602084
z94a23a0273c060ace49d442b787c6d73f9df0e064e2049fba68cd3995f1c4458f66698e489e21c
z7ffc0680a88a7c69f8746c75e00d0f0d96e2fc433676e5a2362ea898244606f851e2c0418b1bbc
z0bce72a25beb5a9d4ab4122e8d6487e902691e98ebafa7b41330fd467f1968fa06b242d4473acb
ze4da866ad7c7f2233c89c63582d4818228986c698d369c37cce201f59f2f31b0f12a1c36ac8f7a
z8d8b35ad831d84a17541f0058b05a0cde7ccdc48155889e918adb792c11981023d1374164d6e9e
z63193bc020d421629b7da73985965eaed55c4be3186313e2d9c4bd851599a157c7e0e1dde5c9f3
z5839b20b506498c5ff947d62d17a331ecb19ff89ef8aa71394443d11e2c6da84bcdbccbd352558
z9eecb03bcdce03afb24f0fda0bbf742a8c3648eb5620c7f947660474c7916b9373e8bd775914e8
za1a261ad6b025767bbd28693e4036cd0ca962408b4436dadb5fdb25bbf534e6d2ec37250e1dd4d
z7e71517dfd11fcdf0fec887337823bb591becc008e015f3a7bc92e41be0e80e4239ebd1fe4bd02
z09e66162a9c8793c69dd785b39bedd4644bc8302394b7c3e66bc5ab986c85beb0173beeb16a905
z7a0f3244110509a70d65d28b9d0cec97e4c70d19369b3c208cede0bd50c9fd39299dd0acd15a76
z19b86c37389520d2964d34c282c30400b5e205701ca050a54bc1b09aa197312fa78ddadf1fa3c9
zfbdb50f618840d088970884560fa3dbe0b53681d590a7d2d7e646cc0e01099c366c6453ed4a0f4
z4f2cc51a95d95764f729f790e007a5f2e151852f804a2d5881a2cfa0c3e0683f16da6997592df4
za3e3418314df11e3018ea14a3df7fcd45eca0543f251514818daf00b4069ab09bfb1815f50ec73
z2ee110f04f6ce863bfd692680543fa9f4d9af1c03d917a3343e99933d7d4c2bea1366e4bdc7b1f
z0404df976c8c97eed0cd8e1da609fd73d67a7a624eaf3faebb870995ff4186a45d901007c78a6e
z13859b8e98cad78c9451661fb89719564c9fa4bf5269b3cd37f03c6afcee8696882bd6fe2f4cb2
zd05c5d2d7b10a463b9c874c78dafa56a366afd063b697a03b3020bd1f4400e6c5a25c5cbcad23e
z58d712f153059abd93bece1f60557c3329f54ee5366e89d7f4763255d88cc7c2b9516f67f5f334
zc79568ec268217bac358a43dacfd4033ce6934d4d4e78dbee0bda9ea4c988423aaa2fd6fb19367
z8a419fc35eeadd47d3bc7745b290e0f87d3f4dc286f619a786c64a52836d4a986edd08a6a352b8
z981faa1646ca5cb1b58cfe433288806e1194b87198ccb168499761800ca5cc590be80b2b042288
z0dfcd30413870b53ae88155ab0672043501fe7407069224eec92d8252fd62b7fcc849bd31ab987
z08acc7428dd7acd8eebb083e935cd85bb035e1e492dd28a1be24ba944109f7f8591b9ed5d9fbda
z46169d1f8ccd6847b9795ac1d73e39d6f125ad2886f38547110eb210619279ddc7c7d244fb8f92
z7d0ca94e1e4355db4fd8fcb9d7c656e5b8abb66bbc80229a159143ef51f764782a510bf7c93c38
zb0352f477b59a4a9e0010c30f971c0324e706cf9bfc3a18922eb63b7b8485fe6c0a1763786b7f2
zd5e50dd11c2c172e4cbe888b0d927e0f482951d0b28141a87e4bc32aa1c71b7430a5273af7ba75
z961fc46908c50f7ab6debf4a1dc63419ca63ef9926a4634889a1cb2f2a8f809bd904bee5018efa
z0b60dba6113d3a32d06b67676cd868efd2eff90dfcbab4d678ada18d7cbc58b1927676c251c5d2
z572b640a91d637b104441198566864a2e0c600ee32dde78733427cd48419d955fccd4e2c42cfd8
z955aad73d49e428eac447a2884d189f9ab3244376d6ccd702e026f3ee5c534ebe2447edea00e4c
z30c1081ab645d237ad60a5dd26039173e2b469e0693ef3bd03b3f00f17547aa1d493d4f92a09c2
za3df66e219293cf2157b1083ad669b16ec706479b3853f2757afc5bbf495ea15cd0c46cebbf878
zb9cca4c25c1e62acd67b93aae2fe9e716e9fbc9520d4325ad770ad2d26dde39ac1f2cbe72f9c65
zccf5c54e8a39100188b80a5b49221e22244cd13146925d916a1b3d63eae3906775fd6c86ff1cc2
zdc833ce7554d2cc80c8f02b6330f76f9e37d0e999c6f3a78762eeef98c769fb0cd2d7bd7377d15
z424394b1356ad9b37ed0c053e3ddc816e00e5027591fe6a46cfec4f8e54efbdab342b803f7ff2a
z10488ed003bfa052722089b863110abee22d19d6842445e5fc169e87eae4c58994c3832b1d741b
zeb174b3156b463a8978465724edc018e2ce0be75858ed47a05bd5ae98c18780958978188fd02fa
zd73892c4a226b7f4f3e8fd9b631bb7acf00f18c90d2781a528dfa5a9e751f40af7d87bd78ca04a
zd0df60c83feede1cf551a9d00bc203236cd66345503c548590cfb033c02c9ee311e6d7266e1ee2
z6bb9b15e16dfb46dcfeba3626c5e3a9c02a9f941b306d9b051ed1d9c753b6fb8b25d996ff7cd18
zd264b3f3a3e117bd4efed98bdf3f5887da06cebc7d5c8e8642094e6be23a11aa0095add668b5da
za6e4216848b6c0c20ade2cbfb21a28a0ee75ed72aac69796beba179ab7ab72fbd0c8c7dae4735f
z1c35c3d435249e99bbe58365ba49287a583a93c95488eab08a8b84621a8952287f7f6c5f84bb35
z8aa3f4a8be19c3d1b579bfd2e2307b8576ddbbfc6b6ce2b971a5b2f084a63e3301d4b6b14b77f3
z664843aa7ae6c3c611504c7ebbc9b5dc347a5a0fea7b37c3a05b560111d6e742835f86951d8410
zb86c62f7c322e355ecbb4358c47adc92c0024d30d5982851aa0bb0d493c24181514c3a4fe2ddcc
z7111006d965954daa51922e61a5303b7b10ae37060f01e1d002bf7074efab3c34d8df7055809f5
z131903eccde381598073e291336165365fbbc8146cdcb721ea9b7e2d298f450036c2f9c1f830cd
z8fffc5df1bd3aef5d69a5e85b11c9fca2b6d41450d5dd9bc2e097d320168cacd491e8c9d584d0c
z279c0c9d331db265ed647c32b8844160bd6058a90d064d3484f202cff4fee0410509c00ff7cc42
z582cefd0ad6fbc515e743cb07ce328bcd05bd457f57afeb6d36db800ab7f6428a9f21361fb2df6
zcac4c90dbe6ff7c3ddefbd335c7981b2918b89095ad4aa653d779a612f13d952da37d4f0a945f0
zec62207e67e7958e0be10aebfe5abab0927416865395f713e61dfc7bc3e3a63ba8f47a37ee907b
zcadc711887b3ad67c6113adce82c9103147228eb1d2c382517c396095cf19fcae61020565ab236
zd67ee07c9104c14f6792f3eb744c8411e2da36b6c78239ad4f7fed44421a30482819c2fab11686
z9a9f8d2c54441f56bda9c42de42658e034689b9924d7fba04864c3c3ab494c50c842b1d4cdf1a7
z6ce7ec53f1cdeebda6c01451d30a09bcfd61b1326072417b50ba92ba1bb020b1ef0808e0c62446
z64b703d82c924468c302f04ff3fd142191c2453ec793741b39e5de2251fb6a643366984fcab790
zca1da10191179d92ca7b34a825d22a54ccfe5b5848bac780b702b63d65da8df3e99a81df12cf9a
ze9f9fbd195298eb690d789830eb2056876d2d3d41f43aae277d78e2d4c4c1dfda6c5957c010507
z29b6d104b5dc9f3419c014edc0dff656ec209ae773a6bd6bd83d3e7f57667d6099626a5c5a2120
z924b3f0b123b0db23fe66d694e7d1afa05fc9394489c0f487f7c68e2d33a93bec4b04a951784ea
z786eef9a83982e08128d1f65e892188293d9674240b4789e404ca7384ad383af5c628525b0787e
z7e7a3068a910a21411a294178db18b3a40c6cde7f089a6762b35e24b87b330df0be42ce5e430fd
z5e2b9c641a6e321dba39986aeb5f396fdbb4ec3a87617e782bdcde4fea13895005863b650f8d1f
z6c07bf22b40c92a0c652055167a0e781b0bf1eb98d8fa018bef8c0e712795b4b55821dba99ff17
z9fad32f97cedc12ef30d7425fcdb149621318613dacab1d1d9316d4590c0133494d084030f986b
zd5a748702ad49158071a4183f52f981478082571315c7ea99eb4eecfc956d6f0ee5090c7f8323d
z3085d12404987a4f45af9aa2704e68773922232912f74a724f6c8783f13ed65fc843da00fc02b1
ze37a3336d963af7f1531c49f2de8b6e729f510b397e90b14345c9ad7eb9328164d00e1cb5788a6
zfa1a5eae615e30137345d18602feacad83781fc2f2deec639b3442c44e5e5396067bbfc3c4ed74
ze6fc6773a7f7f1d89399e820f110628ea62fa86f84546aa9d9e5f908211898b4efc2f7f733dad2
z84010d5b677d7e9efaec004110fdf0dd4be18763fb85cbf5c4ad721c4d5c259c9fde984fb2db78
z9cd5fbe138e252578a542ff5d59c3adf88a252ea54839ac224044cb25f7a28c5acff7c4c9ec642
z80995921324b40df1681c63a33ed24992b8e1fa7b09435d9210079c680796646f067033cd66d76
z21805e500e6513f92255c8d64466e02b7b0d3d632c00f00dff8740ee21c2d28a732f5e9e58802e
z735e98a0f3fd3890259fe6ef87deec258c86670ac913693a014bdafb77e2b6f0de6c691e19e064
z0b4bd248b44992d5f507f3135003b486e945db9d2744f1f6079caaf0c48e3c117d012851123889
z836da0cd304789a95bf8e1329c580fe662b5a073527c34c4eb683f89738a8a0490c7cba0333b44
z2df05bca904bb2153fb35685576c2a515fa3ac415fc0475535cbf0c22fae404bac7aca8b30a0b8
z21e8b3e2f33ffabd30b93f348ea079a9a45b0f6fedf6adef648ec6789389af6b551c4db5772754
z71ed6b0453fcda0b38aa9982e9525bc3939a367de2f1478b416002cc0809424f3e4fb205affd42
z6304ece46b4d583292bb6527c9c5768fae6df6263134746e572978e0b0c81934e2c71707c40d39
ze39913096f24487a14256da4ee4ef24e4854293b812573a3d46fb7befa4aed9a794c56e2d6b50a
zc421874c293fff5e8be7db45e36547b275485642bd1223936c3d6b14607923fca36b97e96115d1
z7b1921698d39e11554b57e8104bdd1b06cd24a2e792e19f52cc7ad1bcbc20b7c6f9a8e091191f8
zf81454abb591e09c22b95f8269d17f763363437bfc8bc9f9cb5ea1ab4e77fe77e7da2708844619
z711925e7abd59ca9af66780990753e32e57856e246a2bb3387350f3e0fb011182d6ec164ea91d3
z29c1d889ad444dfa27c1546fba8569bdfdc8331ef76e1cad8f3c96acf3756e2726c18c6ec73355
z2bd046f81120e31e8f58321bc398e02ba42d3443981c5cb530cc673ab304f2c0193158b60ff9d5
z5af9277d18968d657164c0f656b85591cd2a61d7890800cfaff6d090d87259df7adedb52ef1872
zaba8249c5bcc1036f3ab7ffca12fb8e1fe97886428079c03c288441ba1de79ca10c3008bcb6a7f
z31a8343c88840f04084478c8b1e2efff285b3d423cc92410a4afe6647b173a9721ebd3c3b2d57a
z974763737d1e33cd954a6f9054b41575cb5f9b91b2f916590418caa25686671e844737068e7f9d
za81c5057ee96b15f61b5534b62c4f1e02a6d3029011a331300f9e5889c08b0dbb50c2e107596bb
z4415fefa97d4d51abbc92673de5b59e6a3861dd91be49ad44d1980eb6ce11561dd7e5f9c44f830
z659c7edcbcc509d288949f421f2eedc27372c30816def27386f8fdabc74506ddeb02eb8a9e597c
zc6ba7202a8e41864519d49727503dead7bc39c7fc47c0f26693929f30d9a4af9e085372fa2a08f
za913f7e0dd46d86130e2e3d5252d69223368abda35f6f76644e1c8da97ff4c00fde7757f49019b
z5ca0ff67d6fb5c58af516d65b9510f68719ec8393cb73ce1fea6d6fb310925c7d503f0bca46ab6
z5280f5f80b836363f34fa349aa7a1de791366233641557eb9d1058d93558f88187a721b12f6e03
z9f7180011330191a4bcc3157953a89ccd4b0b3602058e7ded1a0e569a613aa23c84822ea9629ef
za8951b1dd38bebbbffd8d0afc5cfe5a225dac8d7bd73e09bc4424cc9381b39498160e11fe2705d
ze5a6d07821f1747cb1975ff41b04df641fee28a4783037e6d9d7782d088988c7a526ff70551c1f
z8f81110dc0dd5913f0e078b7518ea2cd25bcf0a0aa59dc14459610f61ed1ef030338039bd5406b
z50a8a836dbe18dd5da0c7bc915b490ea683e092585256539ca2b7f5ffa1d863c8017ae2eb383e8
z572975b401fa9998c0f257558a8140a3519c5fb8e4e48aec6bd2544c78850c44bca7cdfb1db12b
z5d91f5179f15044636dc566344b7c5a3fa08b172f7ef58f3d8f1986f90a055adc99d0654506a09
z19c41ab7c5c8816d4b6fcf3722b8b2c05c55b5fe6ace7550ec9e3be716b5526dc219d58907c3c6
zc9314419e8ae5d91c913b264154cef87bdefb71efa2e8af49d16f3e45be95185be9ac3991de743
z99c1afa1f37630cfedb7a0fe4b05eb98ef154b983a13c40b59cddebcbb0ce2a6a20e43bf2682a6
za76918df43d0236aaabcb7123e729ca6a5f0caa153253a9837b517ba3050bce7263f54e8dba9c6
ze8a30b50566b2c08d21b28ffd85c785bc861ae67385fb35a1b628794ce47df164b060c12d6abbd
z2944db00d1d751a7f104ce4d06bd347fe1140e619fd59a4412290379fd07727c44083001196587
z87a830cd2fd8a93d0280c6351a30c986556818cf721a408dbf51dd93e139d5cd0e3366c6230cec
z8e24432d35b41725aface1687fe28dcb877c9cc841d7b249726e538de1f31350380fbf2bd4873b
z44ad2a249b5283c55dda5ce48368cf3a0e04f0552194307dd162b6306bcf8bf08dee7b83d12d72
z78625d7ec41553d648dcdc444710ff270cb58be813097a9c35df38b61e8b0cc9355705a823f833
z954096d3a80e66b45518cc61a86e3585012fb4a483b73022025bdb41aa9d56cf14d3d07d537cec
z2804212c53ee282ca0932324650c87ee2385e8b16ca0913324b71d8f310c2b44a107dc3a57ce4d
z067f769a72c56695b12717c700da99003537f9476f134953ff65158a958e07e20538ec6fea318d
z376f9b10e34830a75f4af886f0b936024f460033c0cba28392c9ac0d14f222dfccb0d7f4e0dac8
z120e1826a4e28e01eea2b65dadd54aeadfc0978fb16ce86bbad00b66ea85ffe906a2746e421d32
zcfbf18b0e3e726aa84fdcbb9ffc9eb3abb4fcf84506793cfa59a5cac30c73382bf15a40d7f9d4f
zc40ee7f3e4ca86288cadf66d5096d72ad46ba082833a1abd8b03a1097f96650149f305458c264b
zb9f42480ab70187dea69a8d7e34b32e27aa4db4831e9b34af9b5549d5598c88e2e92f939c5e621
z4ab34306bb5071a5fb11305a08af41fd1e733539d8637252bb2076865917e5803df13df5364057
z2faf3f2287d4c517993088ab053ca18ebd75dd5654966fdb5192bf348d82cb586d2a1b7b1676e7
z6df640de177da07a4199aac8f77b9c74eac31c383d6e9565c0804600a29d4bb8bf7d76470bfbf1
zdab23f8f2fed85e20e667f1e1c460e77f8d12e293c011ac937d89b77010c69d404b4241db8ae72
z73a5431e8105cb01f47e30e5b17545fd78fa1a3651e78fb96c6dd411f8f505e493967a19ffbe72
z578af55620a4cf1b213e654f088ab644c54516709ff0ab48e457494fda5b8f505a2a1dd5cdc18f
z6321497a839584d60c99933a199e23909c7854800997456fae44001889ce20de85e76d33ab24e6
zb80cce2b9e2c3be41ab22e2da06fdf9278709a8f485d300a104ebd0bd2b6136ec609df6b0e3436
z1c75f6339fabba81fb19af40e1a07db2915df905bc75b5ff88bb9924653814e30adac6ac92175d
zce0719b41644ef84696a292dbe44df56eb287b601c6c59ad9d11d14d0e60294e046b6cd16bf683
zbd58c350b091eb951aec30fe02a3c19d4e384b6475bde4e47aad58b9e208422dfb3114fe527418
zb17965c952fd2c35dfc017ff3ee656b3f6f48835c9ca4064e71e7a6bdd22134dc6874df7fc5533
z96a8258fd3cae8c55a5945e8907977a28f03f0343c65979be469a5158688c8c122710746ad43eb
z68865907ca5343cf1fd8c1a91e93f5ff3eb54e7cad2327f1df49253e9414b07a4f0db202f1f2d7
z0edbd2d93ba405e7063ca0487a3c4ad1148290f55887b1ec3d1dd986d2d98a45a9419b4e12034b
z88c9df4e6b23e22858bd6852bb61dc152808ad1aa24ef420ef10afbc6f4bdcb8b5dbd7ace5201b
za81833401f7e543e50bf7ce79e51b728aca54a69d6e97d894000039155bb44ee6891cb9b0b4bee
z1c225bbaecfb4dba424f44bd0a3341b857709b1e2ee4a40a0c516408b10ddd283e6cf7bb4557bd
ze29f75ade018fc83d3c8589c10b6cb862a68e48b78efdf3ccc3cd767bf7a8b2f1af91aaef32900
z9626c81930525a5464fa75323747b902276e72d9035903065da02b3e57ef98124c5310ece0f8fc
za3c5ce14ee87813e022338915d129656663ef136be8a971151666ce81cf66b078136e179d825d9
z3992170043518bce2022ef0a6a843f30c075f987c5d866f89d2f7100201d78404fce0de2d10d62
z023999f1a82dbb813126e82132bc52f93a2fa7c1865266049941e2be0febf73901ae18a8a05d48
z75737b28043ec9ef89b8a521d14c0f45a44174e57dd500e47089bae0dcc6d0e42c3b2acb5d76e9
z21330a2630896c1a042a49722fc94f7e4e1f8af0e9ca2690ddd967e1afb745f1b006765533b1ea
z4e008e97c1caec8e2d378769a184d06591b1114036b49fe1f0c4b0d8443f567b9fbe558d0ebe52
z41f936c30ba7afb61a8b71abd91619895026647ea7d86c53183fa0eac265469f20ebd449b56c22
z75eea4a850b680c6681c5d6951fd70f8656250a9a5b54b5a240ce4e35033d7974b6ee5c9a7701f
zf6072e33164b9f237e498afe7a3accffd72c3a0dbd952635ae091d5f70b62b868792ed47325c30
z2cc34a48554f2ef6aa112d3d3b4208db234f987a80be72dbd0af27fc0df0a580aa319d8c50a73b
z4c965719ff9dd91d533ed7ec5e8311d1c18b7dde52eeb50010e442ffac5eecc0d6844b3eb25855
zfc1d1cfaf182116e32819b7594a1600521e511be7fc8d4d4978c6c9401b369f516872dfe4319cf
zd03c69cf71e1ea4760d0f0f232e90e3471da9372d0c9c4fee8a2ca89b40ee7ee9ea74715adcab4
za033a18dcc7e45e169987ea4c3b20ad9a98741a06cf5c3fc6edcca59e14a530b3e7e143927c55f
zd47dba63570bfbfd24f9973f576494675b49ffbd4bed2ce0b3cc8475c67494c5d9e0a38bdbc598
z74107a79ce59e467c84052c651845a44edd7db813fbe3f7c47f392f42bbbd0f7d9a2ed1aec5edc
za300959fcee8518fd28aebbc3358473e06a60b0dd56152d8ba82d469a3b94491bda268d2975b26
z37033458d5a7ad8fadb69f1493865385fea896a34910be1ecdace01d2acb3eb49c30f9b12e8597
z5c3a6683fd6b5738c67273ec2cdf4d183248334a52a35dcacb2c0440fda44d709640898fc7a202
zfdd579ea32c619f20e6471904e4e42ba2bc6c7c7d3d94958dfe6235a5824e562607cec461e1e43
z41e1ed085153b65d0ff748b41b766979dd56cc932db03bdc7272b722726977c9d9aa27b23faa7a
z273db7c229eef6b47fa84a66b83e514d13883b5558007a5885c40c9c14ff5db14bbca08fb7b998
z1ebae8caf3f7a9b6f6a73aacfd28bcfb19f7907fc9962971a71f83cab27a6033fe8a2d1ca27f57
zc837469c775f444ab5f9403d59f1677286adc06f55f4f6e9115a526c70810034fa0573677c3859
z2ae3c2b7e1a40d5b5d1f79b41e1179dfe94824ecacfb2c32fb6d0396520ac00f93d9bda8c0f214
z82d0d660ececf3356a92a6826761b468199806c558c014735ad775ab58d1bcc24cbc2784863da1
z5e4b8f2bcd867cfc09f0e84046238fb2639b29685e1bd471ea1d6e1818e657f8f1f28155e36778
z1ed05ec315ab58bcf47d1af3d963909968dc9963e0548a3c590965f74771173a8ce6fb64ef319e
zf7c2ee71dca833053543357e44170e8b727bb31b9bb59d9c37f3991b6f1d6eaf2b3225f1bb2643
ze3cf7b1662308b9d178329ab8e4f70cfaeb06b0e58f37331993709e6e23e76ecc44d2ea27dd92a
z45b7ad6fd918f2bffb8fc04f4e45077665e99c700fe775df814536e9d7902c388b82da6ef33d0f
ze8839e27aa198d3465414b7fab0591ccc6617cd1a65982ddeb347c2bd22f337a08e46d27ffe5c2
zcd671f480b155ece63c4fbe6aef896f154dc2925925bddbe4e826e5861a52a74fcbf405b54f597
z4590e0d1245302b8b58c92dc9fcde3cb87dc8cb751a7b31f69cf0a97b00326f693d6bb8b2b1b32
zf0ab30993ba389f28ed94ba40ecaa826d15451bf760d58bab9327b6651f7685b39ba6ffb4b4cc2
z0f8bdd553b136287ec27bb7331fa9702e3c3e5e31f6e76acff30d991998057c50c5ecd28458db9
z1956309dbee4432f74d08f7750726678703a71b1b6cdc20401d0f970fb2b50a3e774dd929ea175
z69eaa5b6f77bd13c63029b19398dbb61f47a42e5b64763ae462a3ffa56e505a771728554395452
zf72426fc3b000e9d37142c6fda5300e49283f77864bc3ab598625eef1392eecf19d240aa6f7c1b
ze162561740b0ba17aa48a5ae531867d78ef202a0ae8d2403ca6d313aaa63c8ee3334275c2ee760
zcdb1d6c7ded4d7b2b2afddcd92d42a5dec5555874896d5ad6ba167f8253c357704dd03aad18acb
z44025522debd2b6b8dbce641cc22556419acbbe1f79e61a8c982bf3727a437765e7295630ab9ac
z5d91ceae9daee4a56c061bd6fd9dccf9abd35c9f6e3e2fd1005ad4a7cb1df8d1e7756cbd0fa6f3
za7d30b8725d60a42ced3ebb26be08ec1d0353c6f98674d1e25479b01104fbbd441b74a1b708360
z5f10edccff889df8c04a05b598546054578a7d2fac9c4e85f331d6d3757621cb178d3b98b0a3ba
zc18ef9fca99939857edeb9a04dcd3927e1e8fde8d25558b67f10970410f9e2fb1fd9db91c8084b
z2a5b3f465c209f5c4069fc5de8d4407b94517f611ca2cd070cd1aa141db2f6ab47ad4b6a3a3fb7
z707037bbf7167ff83940d7bd03b7beb7094507a9a366a4cd2175d5b6d3aa9b54917b2a0623ddc0
z5528354817fe4182f48150f74f8922fd8ceac01ca5ca9946120923f7b8001d6b44479a9a400ae0
z628a192daf2d9da5fc5b9b338485b0d965a0f895d11e3db6246f7d36e2f4b032239ca2e53adc60
z29662d242f4e4f4a9130dc23a386b76e5b5f0d098835e3436a19f23435a8aae5cbc0398fd6390f
z1bfeac188bf37e1f1fb0603ce0704c1307352c3444a29c1fd87531fb721f1d60325aef4e4de1c5
z1cbcd0ca64a38bbd8e72e0de838cfcb9b6545cbc886c3ce0c085426a1a7b8b100b87174b6c08cc
zac6704e020314471d55208706abcb8d241ee407fd0eb2c79c90f9274df412bc4aa547a7af1e95f
zb169b0a04d59f202ced23f10ad39ef30d7ba71d28997bd38cc79ad6e475d26af84011ffc8df04b
z67be4fbaf51f16d5756efb6182ae3e684b74fe82eb357e045ebf34d9d5e493a506da80e8a2960d
z5956e4a1a0be7e829ae84faa93afa2e580d16e5488f75bbf0838192319a57a23e6dafe986a75a4
zb43f9c4124ca72acb6509e7391f696c41c2a5a0293f2a95f589fb8a1326c73448812623e992ada
zfc03da4bbe95605ce6d44c816a2c0ae31cea2fe30786efe04e008e560337f75656e6f5de02c4a4
zabb7df38fa04bf3f2ae91c98b5732445c1f05e3853cfe191ed9a090cea6f1566a41667fd5d5832
z42d14d4176e50e62e16b3a35959dbf37e7381076611783196ad6b25f276ccfbc4966b0d0bb8d12
z8b5e483accc19bb2f66cc64ff8deaa5721d3b222e44f08defadc18505d335d2c86d881cd1204f0
z46c31bc1f5411346db04df4870f71beb2f73dcc16c2159080958b39c41220b94ba37b7b65dafbc
zc050fda47e549e090a81012a5456b782c2da94be6f7a4167cff54942a4b34fd00b16801ecee885
z178aa020d2a7e83c450d55407359b636218df3dd8d789ecf6071e447f6c733cf6ae8ec9da9b51a
zb53a6207d8c86da14141f92c41e44c6c7a29d54219aadd9a6868095b2bc9bdc687ac60019e8a84
z3f3a87689ab78a5180bbfd8a14a6745ab446b9dd2e0c73d4d9434e50426fe990f2f6858742a7b6
zdd8450d911cc2b042579b565bcea6dd08969829f6c6d4229fe4dfb6a891a6fdac1e2e1e8c64c92
z0c04c77dce0d6c7056fd99d03f56b4212b27944684a8e6b053e56c3a98aed361d58e587a5be46c
zf1001a682505197085f2a619583861c245313c5d5ba1580cffca3c1fd2d050a3c75215732d5848
zf00383db06d41a4485a54b83319cf052d37a436acd5f64e8d80ec505122551b9b6ee265ff5ded0
z0fb1da631f6ce21a3a5d8ca9b2b164ecdb12b63f1fcf0314d6be76e8e9f04378ca62b0b8147048
zb60d02c49ae5c3635a6e1a9452da05fda7a2415124748f76316f7c393f0708678a44865509f8ad
zd9693bdea5d8c8e7987c8fd8de1e25780bb9aa5a4021b08cf6c4acb4252c60e40513fcd6be26dc
zeba7ddf4554cab29433e9b5c3d27aa24986315954140595a3e7daae31496732ce847800ddddcf9
z035b0e2cfe6087ed6220531eda29c25097e37a8377543c580a93bddb38f706a8e0d943df0eb8e0
zda5e157a6ae3915101d22b1d95dd502249fe9956548bed4011a559ad2a9211e54071b58ccb7f0a
z6684f768231508792c0bba18456353f4f22f3abe2a13c4bd5aa3947ecf495831f605fd4ee88ed9
z6e501be3b7fab3948cad696910419144588016a16a0de39784781d125f69a4309d68f7f59416ae
zf376ca449e590f33ac4fbafe4649ddd54d8d1dd224566b4d8f5ba8c9b40100c3609bc564239de2
z26f3834a493f3f85ac3113af8c76ca39bf36a7e426c930c072ee55f06046782136ebc084c1b727
zf48fb84c8e6c3ee4f151cd9124a6d3e5eeb9e1afdabdfefea56d7d9a66d58789e9a219f0db034d
zf83a9ac57fe4da67a62c95d38ab44b96e4bd605854455091cc064511b37c178722811d7ba0be00
z654ae7a77b894ef5cba57df93baea6e3d2ebb76a1f885b838a6224b98f934f8bbe956020386241
z4ee19efb9ab0ac31fc96ebfcfe65a29ce255b0c2969644763dc6927fcfe08366f1c103ccffe889
za31f0c65579326fafa9eb7291fb876f96a6805afaad64526b34f7d4be3a569d6d88c55d4943a37
z9238edd0d6810eea53bfe4c80bbe9b817f7d14e05e52cc6451659989f941f730e1acef639acd5a
z786b64a652419a70e2657c9bff0ed01d82676c5e40344298b01a21c3efa68d4fad6529f50794ab
z59f3d3fd481d9ae88de0106cf258d2d04d880f77f1bd288e032f07e013cf3606f0c7be374a2a08
zeb6408f0385e724c2d1c4a64fef292f1cb444a71934a39ba3e4ba25fcbce7b152f93192ad30eb3
z7389c5a6eed5faf4acf75cfa6976c4fb8c3e5e85bb330c6631ad4ddcf7ebe1024361918b564708
zfd981a74fef619fe67f0fa5d94acf0ad680e0f6ac19f2e4a53b833db26880578aa552b9109002e
zca88dd9f08e35e96953f18e1fda7f9f04782f76a513789be401bc9bee6fdbf8acb022ac45b7ffd
z97c1da578ac7c05b9850f266a759484c80f158a208eb6c28c7f4ca5ad3ef19a5440476cddf8e42
z1e86050fb94ee7ea788431bb9083d08d5bb9a176bd5d62ba9a9ac204b4250210e157d899a6a46f
zd8d166250d68e91a3fe429983260f7754ecb17be28418ee54d7bf4ce0b364459d9c646e67e714e
z4f630f0c3a9c58d6c1aef7ed29cc8bbcd564a63518f842ef4fd8313199750aca07c12af5b43b42
zf04340aeac6f4ed958916cec6b5617a8af9be5f2bfd6bfdb1090987f17a03160fdd640e29fce84
z049db8f486da4c862011331f159156e4d2e6789af056e330a7829c8bf1d229e675f6ce824da3c4
zae9d5e070f07f38c94773e2c7d2b7c5d90dde9111391d707b367b88323362ee67bb551cb1801bd
z286925c5622e9667800854ab373f601cb0021ae41e0503e1bf06ab4bad19b80b705b54b0f9de79
z14d36b578d3902d7fd5ccc39aa038500ca416b8e9e65c55de81c281566ad1e735c48f34855824c
z30c6f76dfdaed1e0e062dcfbd0a01805e116b7359d8c11118d3c2ba9daffcb8cf816be1723c7a2
z2f3df8a19161e6b58be247dcfb93557cb78068397284e5614fce7c4658d8871e54062a8d803760
z59ead8387f4ce085d68ef082478697437710405554b26b641236440ce0dce34d7130ee6e4fe567
z3b0017ae32fe5e1f9eb8aa9d748eaa1a6cb85992db8724dbffa6d2140fe7a15d53e70f99d8ab7e
z2ae422455b6a9da7ad66b303af1d6aa5294c9940dadfb81fd1fdbd3b50044a9652241157d88168
z25defdb8ac006dd6fefda119e062b6a3061d6e2d1819f2a5a4390355cef9ae43e860592a4fd82f
z4ce986b180d8a1c36e0e4cd83bd5b2309d10a74b03a769627446464931b1671cb8e652c8f02612
z8d5853a30ae3af71782f8a4909583aac5873d54af510f166b3115224492296fd94c11d70378148
z2ecc79651af41e116dd0392f3ccf9928e2275c8bd6034386a29306cafa8a4bcf158113dec00014
z7a7a831b4fa8a8eb49b8ad870b5e1bd4856374f5a1c4db204439d47e0f247f067a57ea91a3c0c9
zbee2acc76f33caed66567d0df963b4c69fb6979ae03f40d0eb7cc84efee9da20eb01ee00eca9d5
z2ca751f73ff6d81a320dab1a05e2039bfd689261307391d71f7b9b918471a53bbd8056f1075f96
z37992a5dc01255bc8ac07f270f9ad86f0f84170283c31df28ed1e1162523e3197382ed668bda10
zad90886aa692bfa7c0fdd7d886d11f88fe2f410569dee1f497d8c1b67d19c7610ab4cad4dfc252
zbf11b4471b9c2fc0cf76c8ed76ff3066ba0725a11890c62abfcdb8d651ee996c8ee5b154010f9c
z915c21ccff85a4dcc9da73aa426aa191b65f03e02cb0fc749131e6f48d752356faac7145aa55eb
zedef8941b6b72eb3aaf8b485eaa10eff88412ae0cbc7496e0aaadd491e458d39af6452bdd46627
z68b996c8086d8ddef12b371d3a72b563b40f8ddc58dd7d969b5a3bf422efd1a1506f6db41f00d3
za736371a5ddf88c108d64fe4180b3656621d2d6b9a021858bade631aaa9fed95dbb4cf54fe676a
z1eddffb7bbd5d47d466c49fb15753a517e198b28cf7bee98ceae39a941997a6ea2d8a826ec0d02
z7704712dc58d25972d85091bebbe8e95a4862248509c3286c1740df8095b888cb6522c3c167d61
z94ab6bc64ea8acbccc6524d78832b38df9279e4a563e00cc7653fb2e13c66572d07fca84ea760f
zc491b32809f00e2e574ac3a0bb2a41815a7f7026b9b590c4f27d2c60bc89ec526d1ce594b23057
z11e0b9d2c7dad1b5af3b486679e5d7140350bdf5b4f3e8bfd027d2e9683de011a5d916afba1602
z8f365f87a9df63bd06ba0e42f67035891df085b0d87a2af1e3b848fbe51a9a0d668d909bc48ee8
zfd6f52461c33669b5b0f5212e0daec5156100ad1f260c77f3f023cc5e8f4752aa0452d978505cb
zbe942af7dfa49f68d79b77a4266732a663a5a20ae3cfa259ab2df5f49d58a4ebe25660053a521d
z89539ea7b217cfb4d706239c29c60fb14c74b1a14d5a7dac448577b2f713742b8f96ca4ad899fa
ze02226ce130451ece0f2956aad2452c8c0cf7098b321d17187e4796b4f3600db84e798afa918b9
z21cf5b0d617d32f36d4b5422ba2af9646faa2e0b4b651b6c5775f2f0e07bb15d8df42ecd54ca1a
z13db64b89d6050308cfa923b9c77f32e7379bba54bee04869cb9475bd467c702418e9329b82459
z8650d9885b56a477025ac335a4956da2ced3b298677ae7e5d1388bf7329b7e97b0ac69aa69d015
zc7a50635173d835649c08148199842fea84d25c96364e9bb69139b731b52ac4b414ab9bb9a0728
z715c36f60f5e3fae6ca9b1caca56c991a7ab9b4379354282a85ad8e4d481e5b97ba55107ec0c55
z43c9747525d5953e5720539b4d2021d32973895523cbe10c688bd99bdfea7ae439553ce1b72795
z219003fd32a0c5c90e411982720ea511e93b57273ee05e0630dd02cfe0f7252f21b60c59c493cf
z9fcccb517d622b9c8f1b5ff7b0677f00d055759908ec9060dcd875e9eb42d549558b11d012d730
zfa0725c48e1302d34e10aaa0ff8d74572fbe739b7bdd54fd1c241cf9936add2295b7669b680333
zb3504c81238f9f32c88e478a0428badb607cbdc82b4d38da4e818294c591a119cb7bf0de035cd2
z618418dbe8e7249894583207628b3ee66b98231bc8d0499ef0bab36e39976311677f7814999ae9
z146ec40564a18482187a02bf90e8896c0b7593177fc09f82bae7e3c62555eb07aad6c8f82d58f6
z559c98777c885f183728c99a61d3d154a7f23add9ab804e20f96c998d3915116ed54a34feffb0a
z5513c011b4f54ee2258f18b8be10fc20a00d642c8bc24b61473072bc370cf1a00ca916797ac23c
z3d6ee8fd0a88c988c9e098cd3bc90c397a41256209b47600d2166e7d1a3a2d3f242520b3f47f6f
zdbcad84f615298d1b4cab2f722c8d2a2cb846bdd0b615fefb426a9b050210be4d54eda518f34bc
z1867f4f6c7d83aea38627fa77e46f06803b95c0872efe37779e4d0809d3c991d76e44d7bad01d0
zd37e65cac860e36f7f85c8f4ba12ceebceb3a74de010bc2f77bb996ecf92d98ba08dfb3425937c
zc9cb8baa95849628668d44ad015421bf9197b772ec041b8400f97bcc1a4198013239df25d27a56
z7c1b803c95ffdc6825cfd7b892ded0999f227f4ebadd87521ebbcd6c20c3b5023c3ddf7a6c9a52
z634fea808dce8ddfebc2f7fc8bdca1ac209f464f198147ad72d17163419e4fe0a98625b0a62a78
zf50444341f3da195e17a19ae13cf55858821330e71aa4eae8cb2e7b3141922429ec017d3c2de69
z96ebda57f06d500d47d745a8e7c77fba52184c91967d080ad78c03641320a7066cd6004aae637d
z1d436de3a4ffad12aedfcea162abe2550b4fce3ccf2a6cf01cbd2bd967b3d2a558bf62d73fba8f
za45bf119ba2303ba033316f74b363315d449ebbc9db22c374bc77d8f4b5fd808c1ce9ef97f41f9
z7d5105341071ca3d9dd35d3cc52a09108e374c387668cddceadcdeb265c567ea4f4adaec11154a
z93568038519de795d3356a8c0a08de971fd84f5be93f85897d07bcc543a20b5d07135796a8cc3b
z33fce25d177e49b117ea86ecaa6ec810e8dd64a7f9220feca499b25ae8776a0167430fd9a65fbd
ze229f2ccb8d2f5ce470d23deb6d8b5d35c391c75efb15c35d9299745a24c660ceb8f5eb012dbc3
z70abde58ee919add447994409dd7d481e4852a8d40e958b0f45fb7ea16e9a3d5931487a6c62abf
zb314b86e1407bb4856edcbe2deae394c5a0161d81de13d6212330354572f8904171c371d000888
z367f8cef5126612ac07dd39464932b7b8f547d6fec51da4bd6f289e9f88149a7a2c7c3e18b63c1
z3426dc328b04876a794e6d46abb359822436fcd591f320b7001fccd93f62c5e6b26df7e369a5e4
z73d67cc077ba4eae44f860fea20db77052bcd1d2e3a7ac63f06014d1a55ec78a2898d8351a11f3
zd21c05269a5ee01219799dce19d6157c1cd1b398341ab35ca4670890499bc137a46647c49aff5c
ze282d39b86d3406c1431a60750e7dac81257a6ad34080d325e3c0ee238ce6fd5fb3be3fd608647
z6fa19d76a19d2ece67337a37a6433ce36aa51988bc28a3d3f7de530892a371b35eaf9ee4ef52a8
z51be81786f08cfc9b9b31d1c8f0219452ef1c06c225acefbef5c3320581a4f3b50dc425d8bcffa
z1a02c730ff6a03a95acd30af5a072c2af2cfc107365c4663ddbc312c1905dfe43751072084cd46
z0c03da2d84e9d1bf2445fe181b942e8656d50566f7001b854cef4ad7d8a8a80cdbf5b40fffbe11
z05a9ec61e6b2e8f7f67d664759f63b72d3ed37c2e6e580caabea3323fd9634169ac95ab23539f4
zcaff07af3c9f77312afaa90d14e92dfe783073352fa762ddf5843c2369dcea296f195425df330f
z12cff25622e7703e56354177b68e72fd5e145ddcced66cb123488d5fd779067276d47edca7ec33
zb0ec9e41d1932b853a4b1ef5c75764b40366cf687557bd9fdea66ca714d3cd67d2024f2106371c
z5471b17f20d02ce7d07ca9f2d393ede287d7ae1e82417adbf88a56807a94032c39f2162a0f929f
z591c17505f62e68c8795b7290b22c1756bad85c3cddba3f79adec141399e37a9f17c62b7c0710a
z6de0f24a54be4ef51a87a1c43f01c20805ec2b8f230d746391f6e0cf3014566c78a8203ed2817a
z72488594d1de80b668bd0a670fd5eb6806a02ee8e446ade84a870eb72e9f0ffc1d0f2a8b7c69aa
zfb44f9d5ab70a32f9fefbdd7811a75726a008b4545fe5e567878fd27dc5c476065aeb2456ee35a
z04a51f4ce31d253072cec22ecf056d3612079bde6c26e9b89ba30923e2bb5002c9e2054fa44a2c
zb2a974c7c0c64a68a9f9b4487a1e1f4f57c66fdde3ebe846a0301c5d1cb0846c3a008fe4875ccb
z14fed1c3acb3faa509ae83e4216e74c9ecb1025c429aade58e95082e0bc29bedea87e0e4628eef
zfaa191a6ee0a99b788608beb91ae646d03c64bff848efcb58c42218892500270c4e81188e8c07e
z6c2cc4f9b47ee09632612e8d29f44d641ac399875094cebb7f131979723716c9e50d400017df9e
za0eda20a9b325735634d6a958315518973b6e33f725989f51b3e74aba31455170b18af753b1040
zf3e0cf3f13ff1a8be8e2656a7c7edfbe5e222d6285e126eebe5e545ee54d7b7e09dce14be4ff88
z3201ee8c1ba3d7e79eaeb75686eaff8b0f7dfbd7115c6563a0326eca7e9fa0d36e712e650684c3
z8478a56f4b55ed3fbe5b91c37b2387005c6d6d81b75ceef2b5f0a47f3084e9bde1715ef45d2c49
zda272d96bd940c1c3b1362f4cc4894a52371c8071436e99ea0c51c16f6a7bd1f022f24b1643d23
z9150b561c3edf4c9e30bb28be2f652e042cf350da98e9b1dcfdfea62d27d30f121e802c3f5cdc2
z3c48845c3584072ebccd91a6b323ce084fa2b84793d4273796081b32bc631a5b30406df600ebf7
ze5ec11490dde806108fe45c677a87b697cf557a0d442c0e37ccebce5d3c41171e51129e92c0b84
z74276c5741d81daa70635c5722295659278fb3eab9c3b3ba12bf12805887e674e62a6bd8268a1c
z6b80afa139636e50314a4fac039e3127272c0c1731bde84d03d8e23569a6f1c9a65f29eafd01b1
z64565f750f3bec7962188ad03ec9faa7799d78a1e7712138ff184f57ab32a40fc2164d2bb1a9e4
z48b3bc009e34138702ba3f33fe0d43392ce8c66c93ad82060a9fb3868d41130508421d03d6e944
z403d18862258d457e5c7af0f5e1980804aedddb098982a09d159357330896ff540bc33eec31601
zc06721637e5dcb9cb69eeab6c20b42c968afdd4f42ef5fa84221596ecdd446c2b09090caf25519
z9feb910e175f2ccd00075ef787f643e602914dcbf372acdd13a9fa2f94fe453c4f92a388f2657d
zc7d9e9fd8e56de556c8e31ee4bac7c5a6ee4637295c2684fddacdbf807e2b72022c7c40ec5ff1f
z824ed8f8c30b504214ab467038c8a0dde24a8d9a8ed188debf73cc3c3a1aa1ef5acadab4e8fd0c
zfcce5c5edfe516f98c3a540bcd55f5c28bc16b225c8a80e91d4dc596d43073ae1064ab1d4a3ea6
zc1b0fd4f8bd8804de08d501c3ee78e77dd9f0ecf104e2bd564fc65b8e94a85bf8c60ba8402b35c
zb16af178ca2d5f1d410c917f96807a665a3b7740ba8c9659085d86a0c6451b64eefe77176a7e0b
z1ea743f6a345cf7942434903d462df2685821f463fefbed97a544760c8c54d3f1b84f45fd299f2
z45c1919e5304b56cea40cfbf21bd5438ff7a1f487631ecde836f2db204a883b2bb121ca2e94cd3
ze59854fd9d50a64547814aa79050fd6c457289025a0be527193be27509ef4219ca99c1dbdfee15
z8786c9e820ba4c44f155b8f46bcedf2975a5d9ab0fbc1a4d75a24762b58277b98846b85089b34c
ze07c6d8b7cdbfda488921f3795d096bf4eaf47d5f84d3c71b0ca725d66d21d993b8b46f279362d
z2bd70de71811ea6c42d9e6299eada423185032379f2cd144430b38afddbf8e2a8b695e38c5ebee
z53975e097d00c852f7f60049809f56b1f0811174fb185f6addeceb3e7524b5bf1c199258174e3c
z2c24fb4f8d049d34cf8f8f8d635ea883f79d0ae8e8870ddcc676d9e6ea2040c919b1724aa3b729
zc01a5877fcdc04081c9357a6ceba0ed5fce0eccd5db8ee9203f0682e6c46905417da01bc28d034
z9cc944f41ef3a5ddf96209ddab8a46cc0460887475df56fb5a67a1a05da1f6987031ebcb8963bd
z9bf35da750d2262c6cb3789288d94695ef4f778b9fdee63c52f3d63aea7b0c665402808a975fc7
z28462b99311f469b0ac089107cb80d95dbbb9903e1d27288670cf36ba96029ee537b0e43daf73a
zcc0e465e30ba7f8f5501cd1548bcb088934ba218a6064e59019ca907c1e4b14805e869b6ec6534
z9e6b49d08851ea6348794f7bd3a0efd1dfe9a3bdf96735c61fc0721741f239bfb71de214ce9c38
zd630af4bc6da0cea0b49c1ae7eadda3d5714dd5adee2d953c14be0af96430f2becf919aa1d6a0f
za88bf16b6064f891a0b6a1672a16a0fd1e3ae644bdf4bf914cd801c68a338c43c0212680d69502
z711c221b293972d0c9576c6b28891a6b23ca58603be95e26d90e7cae5ad9966bee0d2864592859
z4dae45b8ff70d1948c4b10c61c9c3862f788da139ce79d3415f0cc6d1c34656c48ca99d19be4b0
z22bdc78aa60cad7e5cb8ea3105eab7d659f0a9c7d95fbb614a8cd2ab7ffeefb1717894a566a5cc
z9861f685b2be348bea048d7b19ec18c8366440a2babb1c82089027cfa0a4a3c5e914dc66d99257
z81ae30ee2d97874ef3c86e1ebea27ee37537b0421d4fe77fb316cf0cd92e9755f5419113c03ea9
z5af1dc7e444e7f5c53ac69c806f1e211ca64dec3f483f4fbe65e0a6f6da20daaf48acf2ed5f826
z67ef2b87230ae78742a82817fb66538ae2f762a8ab32b13d0aad84eb9c841b393fc02e66900002
z9322a8fc4c70a7e6dcdef5b13e38b97a5a85c7615eda0aa5d56912f32afc037a096ec96dd58de8
z6d22fb6ab8cc4042e5e6e1e8bce3685629943384b99e10ce74d13457e4f3c86e908c61f4ea14a6
z183f6b867d44dc2d85d7871e1c34287b58cd3b2dd78a481097b2f03fb4ee2ee78a08489d0149aa
zf459d3a2d25351f5af4e2ea7a1e6362403601736254b104e605e3d03e06741b49cee8e2555c0f9
z4f5c5ac15248572b50abc02de37e5ef127a11ae63eb88dd84677d551896789fdc8b482df14352e
z223f4e2daa8951a3344d15691447b05fa05767ad87123f3ce144ab2046d3053587edb3f38197be
zc3f8d6e06bd9332b8cc114a8e43e11d5005f16b933497fc91b9a17af1446f31ffac082ccc49d60
zb5d636580e44286b3ec0cef69baed9778b10d326b63470d79eedfd24709740b1f37d806eb1cb8a
z4d8092b2d8189b7efa10fe7a1b4887b35f8bb7e856e8345c9f2b7b77a7aa5059f776a80180e08e
z7be72bab8679ab75e07d7268d77222c49145bea2cdf400d5570a0ba2b659f8d67cd92cb7341613
z87461b04d0c8b636a887d263061e1bf6e6477706e0c662ddbfe34a496b3ad852de00a8c1f979ca
z14b6a0d95b7396611aa5c528ff112133fb543407582c2971ffe2a4af0eb6eb0032752f01a728ac
zbc7dbda0233dd39c771ce2ca8121c121e319c26dc8c9f9422361970288d4a432cb00cf8f48cebf
z04c6a5d940b30fcf5d754097a9394361bfce9f8f8266ec27705fdfd6b608eb6263786ea8e8c0c0
z88a4a960479a79e20c8480f3fd68365222344d831aaf01f17a06c0cf42d92482ecb4c6eb24b908
z51fe108f0cb73fda63876dabca16629f4115194835e4d0a46ff1fa6e9aa4e8fe1f6e9b1f4534c2
zd4a07f68fbd23e4dbbd369a62465059dbc97a661a658dd05c039f27dfe000be4cb9495cd3616fd
z1aa2acb02ad26eb1091c81a1b94170ed44b9cb08766f569d8283739f661c0ceed12e1243de8934
z8e74102c3cdc6371da07f92aabfa47bc8595439dc4fe6b085c7bdf63214c801b64f72c558bb3ba
zf1d532a1f74d23aa50fd99193f3b3cf6f81931c60a93bd71e4f34cbe77f1a9de708b3f06b2322b
z1a5e4d8fce124266b4b1a7c45cca36855b09900a69bb44e0868c655cf1f00249c2aa65498f5d6c
z42ee61d1f364ad13533fcf3a7b24c373622438388518f18565cd89ce052c49152e4710cf447359
zd42fb80fe4d18a0a8b13ab864173ace15ac2646f0c232401408e2453fefb187ed3fb7cedc2b6fd
zabbdb054c4c7e340806550633ebc7f3f1cb548566ba4e9db7102479d6d11970f04173951042f2f
z28f839ef4205ce03296f249a67c8785fe394092805d4dbc17ff5331dc94413942ffc8485a263db
z3ac4c40e600968fc0a38a68d2b3b120f47d36388947e3a9d0ed5d6e1054088ef0951f449ecd9fe
z69899303af6d9b432d15af71d50fc35ba8560a08430c8ea2f01e5773cfc8d28dcc4999bc36f47c
z432e5b168b55e2e859baf6864baa49de5fcbf0d61037f589c7ffeee6595723d7ccb3a3dad96b02
z98461336fd8beee8b50e40f6da8ac2ded2ad80a697af4027e75eb75adf8f29a510e7830501ca24
z0690cf793aaef5b1293ca16e0d0ccaaba99c72b59d90ff251f1782756d00dc6a7932f96a1720d0
z2c2c3832e92c30386a97e420d9df5abaad6867f97d43087f11b3bc7bb5fe822874397104fa6d13
zf1a410b087fb99c29a77314ad7c844ee29c1162aaac76f79634a4cbe1a558c31a9835b6a58c4fd
z3d8b766104a1a2c1845cd90d9e16926d9495ab96c5a2002d6722ec936366f3c8937210ac5f8d6a
zba77705dc505c0810f7ebfdbffc3b1e4f8fd15937ac90872fd16e50739dfaea9136f2514592612
z6a14a60d1049bbe7f29c8a2f215ea0d7652d5bae5077393ae401119e1996fc3662d5ab012f247c
z1b5f6ccff57cd4598b2faed397078e491c9a6b4a00c76ff5451449b2f43fc5f09604c2cc455d3e
zf0e8b3d5d9c3f5932dba6ffe11d0ff100bd94050395eded22fa1849d8077780f957b9b66539134
zc79094ddfaec582a41ee6940ac40180b01e089092bed2936fb67d877bf08753a5004a17803b5ca
z23c67e392dbbb7b2af5eee158de9518b692398a911bc4e31006491577679a9196462e3cd286e24
zfa4e4e2b7c50d53a0b029a75ef9e16146d4422202b65a4015fe7dd93073e1fc474df425851bf43
zd1a36a5dfbdb473d89737f609caf583b8b0ed9630f8fdf7eb71e1d5a65a6c10dca83f8940ebf7c
z65d222294a5eeacadcde54870ea8cb92772412c8198d9f8e05df8f76c743b4ad173fd8e97329f0
z7e00af77a14e6ffbfe0078c49e403e9eb3ad4fefa4601d9f2ec872d47e06c39222d04b96c29960
z3d86b28b13d4b0af078eb920e3e1a10e8d99e240205212e8d91eb24ab0505ee59c2131a1f9024b
z224c828599f5d075c4a10c6d73a1a4a7a45c060b4e163332d9faa3fb9ef0c220ea74c0c0232ce6
z7655f6f67deb58bf79598927a37ce9e626e6697be306219e96df415c1dcb48d0c5dabd76ab56ad
z3fd5973849f53b36498b58d51fc283cc3bf27e4e50ad46bbbf5758a3657f86d65728c889619b7f
z8439f94672a5d39cb1022857022f5aa50c388e2c36329e7842cd14751078e02149d292a9d59cc4
z1fa66f043d5a734cd0d162faa558b89c32f31dbc1139df6e841cbd4e21a120235b8ff141701d07
z7012986a152edfd470ebc8ef229e055435fcf7eff6a6a1f72cef8635c38151ad7043cfaa2d0a02
zaf0e5d9c308cd72384c7f94a66ff53aeab7fb8375a55625b489ff58fec16145f051c8b35447726
z47175842d3e128b898441a0e785b425456f818408e021aec9b1dcbe07dec00d8e44d5c824c7f1c
z7f05eede5fac91ada3d6994c6cbb756d9cc3202a0b8c9aa81838a14e05ae09ab00b25a1740315f
z2cadbd9badebf4c8e18aa4daa51137f6c2690789ac6a1e3778cf6e74be5949f17fb21e0fc328bf
z90a9370b67e88e35664d7344cd53534b4363b55dc9a19f16dd7751f186a4a1060a7d0c46deaddd
z390932d6d82c7493f2afb7634a1e4f66b18d474a64bd1c96a2729e019af6c2c6a59459f04528b1
z636cc5ae56e55bc762a10fdb00c32113bd4b375f411b6fbccc4212daeba34c1d4378a1222b5a56
z5d22a72f7f0c45ef00386b492f5b3e84f41176b2c008785e6edeb5978b1308203d5b09e2eed3c8
zeb0977432b9d76b9cb6aece81ecbe9f1f62cb1c55f5238cd48192d93b17f6473670bba488c71b3
zb2acab7630a88c2ddf17a6ff07b8efc25d8879784c72d6b8de68f32d35b2c5b354f6f46b2e62c5
z4c5cfb1f458625acedb0cd2dfadc2f02162b13331e89cca7c028831c8aed7b708ddcea4e3c33f7
zeb66434dd0b6dc5139ef764491d2b8664b506c4b59053a4d78b96f25c28a6327bdca18d774775b
za2f1a64ef914e4af42414bb1f51417985ab95f9d505a8f79fd8f54aac27169c47b1847c13512e4
z5f8f7d1ba98be92a719eec0667215bd59fc398c0f2ae88285b64dfe5b894fa86b6d4d6f8311590
z2c697e9b6a70f3c5b98d8aece9a0ef5d23f47dd12824ccb0e0bce093887f39da9bb0fbc5413323
z282e1cc7e4fd3a2b07506332d49846629cce51ec56513a5c2901c4b5b70cbee9ed8e19f311a84f
zff487ade538b7f714ec284ed930ad0bb66a54bc4d69b3499d10f9c2b41da8d6b92f2bbf78f1033
z65cb8849c588c0b5e4c4a1c6dc8daf3af689efaabf16ac04029ced3c631948a761e7f3a029af3b
zabddd31cd56c58283b707549ed76e9dcbaf06aa520c69d17a04f8c3478729fc95c7305dd557c25
zb1ebbbbdbce78f4ab0e86a9328ef97d3b8b41d2d5325b98720435437491264583a322c7c79bb24
zdf0187cb048bf420aa5242bed9cb100f349fa9fc1ae9df1c0735bd978e47e3895523b6a16684bc
z52021fb9e23d49c8a9985b975f8952c5fde6ac832188498510a1039a28125b13fb460439337359
z87424700691e00f2d899ab32dc88a1714c3f35a275210ee6129110a6553bc94af0cd962c10b277
zd8e53b427e2d3eb2cc2f68435e5f3e73a14a6267d6b35b6da8598fcefaa4780610a6b4c5293696
z2f1917cae277a5b5800f4a0dcbb29fda8d9779544e05c1ca94f5c4cd8762885584478bd106f6cc
z30afbcec4b04f41477fef9cdbc8d2605c41fd69e14051135dd4896d555af2087ca1badeffcc802
zdb2be32bcf388a79bdf90e21e2900e541cd404ecda55ae0a1c0b61d6f765a6e30c0df92733630b
z4ded82e2b6537169ea89b39d1da2d095804be8948eaed9e50b464d0d49a5c6a1b2506eb98023e4
z4e018e0526bdfcc2738a3799a81618c24f81343426c2c22c9104763415c36eee6b5b94cc388abf
z285c83f831c45c8c39fb14c45650111b07f177305d135a2e2a84bf339e993394b62308ed08809f
zefd85fa283183613952a3035826f482d343a624c197aa76d3ccd62a8e4baff52bac26935a868b4
z6f04c2c0626fa0cbb9913c8ed9120702d957189563ab0ee7607a0f006f6f739d529d6eb3f4b1ef
z4bf59bc5e953a6524fc0263f90d247e9e24d32b972d4e18445cbdde9dd619df1b2cc4ea3a173d1
zb13335342a53e4be232c823ebc2e45cd5e3fd1fc42620087741433a92bc8b5cbf88c49ca9d6a0c
zd630e7f9a1b261b768c71faa2e383bf0ec919360552614794ad761a620bf6812c5ea123b5903b0
z0ae2f6e33f955a089475a97d8bc5eba0a55aa901f027e3cee11e9ed14770bd106141d2ac7cb656
z7ba97ed2579307500d891f007e4661b28ebc5b8a7655c85b9bf9d1653fe84075a1dbe12d7552d6
z262a8f9b37597331eefffd9a2d45c554f5de8432d4200e4091e4eff90c9b0bb5c0adc62ef38f78
z02b2eafd73dd9167d40fd4d9c97ba4e752759bdb4c3aef434fa31d545460c6f84c7695688d84a3
zaa9e2006ff6cab486a24f0a2f59d5df1c43ca0f50f27ea1feefd2b7f02f437b6dd610809892af7
z2242c0f5b1ae1f5405f5a9d1e364f90c469a734751637e50ed061e97d5c23ba3384d8dd0e8b625
z86a0754c45855e4e99d08138031204d86963526f919cb1177634211d13c37717abb1456581f6b0
zc58e33221b109dc9950e4c4f9e30c2941f1f36475f17c13b43caab51b04bda7b317c7de37822b0
z9a95326613d4346de8cbf03e3bc2d29a69b8171d930ace558edb1b920c5c824fefa9327d308cd7
z4b279a4dc5530a23f2e34a8ce3e79d2bde765b9a58604fe5d11811c47ae57f2ed0943cc8fd7e73
z435a6446f424e1307328d62a06645f191455289771c917eaa682b1200efad5ec20f71aff2f6e64
z4c5ebacbce13367ff5649b1e1fbe90f98fe9838c892183ad70be697d9023834adb8506aff5e94d
z15b2156d54ae5e73b54bea45497c0a26995910ea4f9a0fcb19512fca8eaef676bdc882f6b2a916
zd5638ac8ec9d3c01ce206419d75872de7670916b2358592b186385926d801dc853c0b3616ea88d
z6204550725687635d541538d27531e4d39f62294f37a1361b84bc9fbda85dd7f86bb06408d4f22
zdfd726404f8f2a745d5c970da82221e45c957e5516160c842a2d1247efc64d08a5153b88b784e9
z6a25a7ac5f9feedd40f1996e98e2ccdad396d77470f4bf6b779d4aeea579f27a5bf768f1ff21b5
ze61e775299bf0d5df6e2b9bbf0f1a42e195dc62d807c5bb809787139c7a4838f6da59e00b1c3e4
zd1c6f6ecbdc0a2159ebe1ac2f01f86f75743edda3fa7c830fc49cf6c8a6766bf79ff8d550da8d9
zaefb2c5c12250f8ed6d625db0799f01ed0e883298452aa143be454970aa1d1fdf51d62bbdc688a
zee4f811e84f4714d44b5f8dcbbf5c568c12280f55dbffb465ca051a8f2c29374a125e12c1c3815
zdda2e62de73610bcb057bac0430a9bfa81583295b04c163ffcf4d73cdb312fc1066d81b37a0417
zc5cb61e37e84d1b93594eaf1785d973c536e919877b57cf292447c4660cce44edd7d0b9e6e6786
zc8400809acb67ae678f50e0ab2b28818789691f1b0ec94545e61b4b10daa12b293a053e035f584
z1833fa769baa18ae3d3c5293e95636a1c39a4c67b05ac6bf105ba711ba2560c705380534f98678
z4b501bce30e4ce74b94493d5d1375d8e58f0688588f10406686f00cc605dee7055b0bf63f5ba83
z051e1532cfa56f4790ee0583e2169e4b1ca75c4a024ddf67c034588a2c6eb7a4dd3e208b6f1ac4
z65745dd9a8b3f869f4df0999a2a226e10d4c86e98ec100ef6fd735584fb904af5ad79e53ea9922
z5b050358e2bafd9a42c9e626c8a4cfbd360aebe01da2ab013ef9132bb1323fbf1854eccb3b6850
zbac9a5168da8d558f48af029e2d49e1db0133d0af956eb5b66b17247ef380e7ea3b2f79c5ff467
zd1684eec2e8ae2cd9bedb1537cef893ff00e7b0b23356f909741d0669fa6c180ff494584b1dc88
z9afbe6d38d48494f40b879b266c19b0f46d7b69b14a9b6cd8eae6b0eaa91e3f77af77503b26e1c
zca08044ef2679cb02620333793997e2a4742baa616923b74f844cb930d98f4692f39f25ba04a80
z32a22272c58e8abf1dd10d3a58254fbedf8e367f527e1ddbe5b6b656faf041157108e1e09c5bb6
zc049587e93288e12474499de0a92f3c34220a5999bafdd43dde0d0702cff7d38591fa1a5824138
z5ae68633c2a729a134b2a308185b58028d153bfb61728d0841d418a6c55f80a19b573ff478f68d
z36f7367e2de550441630f185ed380bd989f4f7612040b02e7650ee2d97c09b4b8d574195310066
z55fa437b32c9eccf6bc85bd3835909c767627ed4b519025d8fba3f275c6b23cec99de055d6934a
z0744f8902fb4c0c5488e99d864ec962567e0e9121cbd6199aef4cf65a7f87792dd83eb23e2b6af
z46da36145fd1f520cabeac73f65e3dcf1bcbe5cba9db066ff638e4080bd612811cc8aa1088672f
zcf8e27a42555949bbdde202069883b78c5bb1cabd4b884de00c90c37066d8c3defaeb48888a482
zb268bb350c5a919cb8bc3acbbb76cb10686a11110971b264f931107f20d3875ee4a6577ad77d14
z011cdd119c3ce40da8dda5cfc3425d6154736ad2dbf0f77122338f60135b064539e41930db3dbb
zc0b277af7f7aa237db556d8011613f44f2f19bb0d752877144efb22e6eff2da1e692d6aca4936b
z4e41817cae945b119ced2bd07c0e1a372cf120f91fb8bba3ad8953ea7ce15f98275dfa7a66bf4e
zfa3cbf57db2b6de977e138bf2c084b0b4ed28669e2792943815ec40b5ee6a82c0b921454ed15a4
z9f42445d2ce9349b21450f3330401194eac2abc8640b8880a80258274f6b1f379a2da925bfeeaf
z4988759661750eadb175b2cd1a27e3c3aa058080da98d5da64da3f7d077f016c708ab3c8dad4dc
z8fb215211de036a9e791479bf968166395c532f99c7a7d1f04f3e0043ca4a7dc3332b66516d478
zff87b5afcfc859babea05f9f8864beac7a31845df5ec949cc5d6e8f41f886c05f52dd17592d218
z80e4b902fef79bbb027065bb694125747719aafb6c2531d9b829958b7efcc0b574cab8d0408579
zb595df5af2ad1371e22d4ed700ce148831ddb95089301f46d79106c25a09569726f6996fff3d79
z22b10528eb77173310b4973a7572659ba88fcc629d2c9aa2e8fd8789f858df67328d2794dcf98b
z2dd3f37e658a8abbb43e0fbb0564b5373e314a87047e7e5c0dbede9cb5d2f62e88dd4e66c1927b
z1d3cc29c9da1318fd8a50feabb8e20f30548b2aed9301c2917fc106180f0fda03d9d29978100df
z57838d29b5f40c8551045bd0b8eb15c92ac214ccab8bc2a348c7e3e0d9b503603cf0d2e81115b7
zb3fa49eb39794938f256caaa3b6007dbd29e4fbd4594f9b3047ebbc7a1ea34510a69064867a5db
zbee0584114969618e70422e5bdc36f408839cdde965e76ff2bd919d4466604dbb96328872c8eda
z090fea392796e675e188045b0750816dbbb1b7045d5d1caa421ad9395e7de30c753aeecccfe652
zbd4afcfe3b77f866f2bcc1cc30f23d93b993c1c1ab70c75bed4b93ae8e3e076869f5d9bc318841
zeb1035004d3d90b035a2cfe7fdb639b66fe412b190a4f83ce7751e5a65e6931ad15bfae792d10d
za3df0b2afa91ad3404b694c868bff9239639045ef7bdadedfcb5dc3c959ecf237bbb34671034e6
z8a0ee80a5212ec044aaea57cd96958c6979870f528936be72de2fc7c26c3a8767edb3bbb1ddde1
z38f88fc3d59ef9a993cb92b70b79caf8415394baf60efb255e38b44ba11eaa43df9c2dbaf704e8
z4a8e66f80f79881f79289dc1f9af7e5a9f19533c87d86585ccfde83b2422169edda382cd750ed6
z9d8a69be6c3ca6d7826ca0fbb00d7c6b55ed733aca7aef1e2f31eda17319fadc104a5d2e156f5a
z44e3f7e8d994e95fdf01d68e342eb6ae4c392bc9a071abdd27a718025aa5d09a29c2e3037a994c
z6ec85da64bbf30a919d9c3bb8baa5312e664e31800154105daf0ecb56da40d2e42b2ca692844c2
z7a4bf1152f72174dc86eba733eac6d211d1255927719e84b2f3f3ab00226532fa0291b3787364f
z4a5d4f57025bd8a9c592d58073c023770fa6f9b89d8392735a89a0a13a451ce6baed2c0630b129
z48160cf18104ff8ab68734a10d3c39785682eef40519c5b5bf8682130061fcedd89f83a647b899
z4e44f18c8e142cdd0c44da62a19e330716fbf827ec2b3c0ad4326a21319ba986c901c64269593a
z94919b664bf787745e8c942fc94e9c80a3265d4d1a18e794c66bab2db96a8745ec4671499bd214
z4b3929db0c5f8a0562fc3a51157ec2196e8390568d2aa8722c6532bcdf9c218f1cb1e0dd386d37
z1bbb255e0564a55ab46b8498ae0b8e9fd4852e5db25c4ed60a9a80a7a53f39b5378812e73c9077
z951a933e59e144754613cb3cb35286581857595cbe30eeb9c9e9fd105b59a3792d321c4b6fc229
z007d526abe1c79b868c38b8f8a84ae9aa674f56f5e2e39e5dd2cc65b923629c024faa78f41088a
ze5d521f7affacb6dd6686c638ae821f238c53a1b9182af77b28d9d326dad1071786195784db6e8
z5ea1db9d1d85e0b51cf76bf8548b5fd1aa4eceda8cad68165f319236618038532d21ee97224952
z3640e532c6b2a3b02f923bbe2e0e9df1580bb09b14634ccb0532266a3bb5515e503eeed1146708
z958170efa31da523963d4294448bb858d94a9400323d1c7a1144588df6342acb1ee5e36c982d46
z3c9925274d4e3d49f6230fd2e227a6bea7b8904f4564540a3ea2f81f8e7ed87ca5b5fa41b9eac4
z86797390e797f002d1ea06a9e59ee45c5eecad90cf00065e8398986d215db537deac39ce5c55b5
z9ca70b6d1e0358db925e8501ea7b0702affc6d8005138c4ecb645b0bec1ce1aff530a266972613
z85e659f2f1d5c121c4cb84ecd64cd74e70c09d425cccf421681de725c479bc229c4497d1a21d0a
z9d3ebb585a4b51ccb459ad8e34acf2e70c295bed5be640b4b64544d4c3d47c0362bbe085a7508a
z6535711b14ebe4f47f818a41a0a9193e7e82dd6db23f0603fb75e0b997553152366ffeb986a1ad
zfd3d4a89c2f87310d317a210a24e130d62d2e94346d2d44fece53a013cdeeeadfb8aa048f48e86
z75fdc3b9463d56e260bbba1d194af4d31d5f9e4b14650a9738e55e51a40a5834e9f73938c01438
z813a9a804233199245951fa04c9bf65ae5520c35c5d86e30e545190c4149ddc594dd6a42d24c58
zf0edf2d1ea191e57fdd06c4c9fe6a75ff2b51d17d3238c3f2b731ad4536e5d7993a1715e7bedf4
zafd09dd9a5d5d524371d2ef901ff6f17d8780079364cf8350ee8f5062600d772bc253ae0434423
z150a442a854809201c82254ce03c550fbb11c365896bdbdfc3e22c8e1059d83991fba2b4ed470f
z263314cf058165ba49d97ad25de985e33290e7ce20875fefccafc40d3e30f59c469ea94ba53c1b
zc68acb1a7cb98cfa7abdf94de640a3df8c130b9d91eef9b2d6168e2a9dededc8e7a5b0f56c79a3
z91881a34493aa475cd90309a97499a48508f813a457bce2ba23018c280ae36295be8c7d37392b0
zce475c715d6a2f2ae09ac653b8110662edd739cffe2216ae4471910845603e744aa99513620f37
z36ec18d54d885c56717208d57c05d51a8c5748c31c850d8210a201e71a6cf30e8d6a964f50d283
zf656c623f274d844206d6f117a983762749937e2de28a55196cb4c4c12ea1df353e8bf04f8d8af
z7be9cbbfb7c945a883af715d4759fea445f9e31e40ee3c5fdd0aeda59510387100ae5ae7dd1ec3
z9aaa77635c06e54f510921d960e6d1593532153f7073d69d77d98a39bac07e80532e5541cfa1ff
zaf085f3564891e73664bc6a5732a6611c22c7444e47d3351c65a7633a8baa58b8bf32a4a13e008
z84896e1b3e7b820a941373f07bb2bd8d67af6e4b0bf57a866457165f05d8f6c0eaeff669c60c4c
z9e8b0537ac1d23406df98cdd6d070a2e441f29d45a762951216871d9419ad928c8fb29a07cbb37
zb52ec7f3e9e92820d34da9987e7b99b362e36b66dffb12b30124e92b3f60b43a2662a5db17eee7
z065b5a72951bb5d08751f9bd692e4cca51b784c84bbd25ec33ce41877e9dab22722d08345ebe87
z54e23a45287459399159e17a22233bd9b019cda545e32a9d1fc885fc3e7e9f7dae577cec5416a9
z2b48502e44e1226ff6955bb0ae8fa2d9ce72340c479277abc7b73209cb6653bef815f5908345ac
zdadb6677396606da6897c4f32d2c09c986d7c4081ea324f0cbd657df5a7fa2031969ef689bf8fa
zad4be7cc5ff3f9b3baeae63d449abca633767785da64450757a8e10f6b9729d2c25ff22842b3a4
zf3dabd7095f0f7587f7c269cb5ab97402166c443cc32703db2442653312082e0bb4d2f89c34c20
z640332d8b339ff1cd93af7269d60d44abfc9913c849931059abd9f6d15c3b1a6b376366ef3c73f
z054ede9f779beae1a3be068c684d3a319dd4acd4a36da2a1164fe6a5b859d6452dcca33624b147
zd084b48fc25061f911dfe32fbe31ce9179edcf5a46fc65b29e260eba3817dca986a7faab2c6cd5
z5deefb4bf76ddf5e1a6fde010d9f23cde5f32a1d6bc0a2385aa4bdbf8624f74b03f2327d141a71
z8637aa2e35f68fbb088f8fc4f9ae4079ec6a9ecddc923a5c290b1baddf036e53fc62ce29cbe42b
za3aad250fd370664891d22730879c87a16f21046a8532451ede02283b777b4c1244ea96f58dd2c
z793b82c5e875121bc272b3c620056eb38a0bee825a995cfcad59eae8b85225ce38c4c3d2a6ebb7
zcc79efb5424ea4895e423ffe3497f26b9f7c83eddcccb57fb278b7e02c78efa5ce3383df9cab81
zd5242784fecb0c2e22d222db854840449003503a4bfd6e57c276b13b73a8d2dc05c1438563e2a7
z5892270f7c18ad5bc8939c8db74588aca2d5f3c700f5a5dbfd743d3607948614eb86881f9cbd89
z69a3a045341232d6079f918c611e6028a646b4ee5616bd9c284c34ed3435232becbd1735d54e07
z628dc110b8508bce58cb685be9e571b7fcd5e99d6c59475b78d326e9f05c6d2a624d7ff325c2a6
zf542d7299d92e5552bcf0b7848bfc177b6d39e8922adb7f73f883e6eb8c926c313df87a13d5e17
z2666a82dc50e5561d4fd8d22dbcf61d46e15115a1a5b697b325dc3c2d259ec2f39a9352b1f224e
z0d23844b1ac28fb5bc29cc03d01463696359265463ce4da61bf9cb40d2c6fd7874e54e29e7fc2b
z8bb848f8346cf1ed1845f654c1b66d8247b8bf84556c473a51e8c6ad86f7be9cede8a3b05e0a27
ze2958d5c3a0faec052f372bf8c56b0fcbd9bbaaf71e727793ec5e345d892c14d1a4e983b4fe4be
z1990031908b0476a1735e63219800c577af3c6b430bc6c1fea3db84a328dd837451e8966a8e50e
z0df0341541eb06bdd5f75894add210ec172cae0ec8540f63cb7dad36a02ccf0ecd92d8eb458d49
z42e45e847f5cda4e2080c2debe9cea1e3c29e2013dafb4c5aaab9aba4aee6fbe96022b8f19d806
z41f0f868ee48eb726b30d01afddcb139798eb7aaf5007bf1a490fd90fb6538e390f4d967dcdbe0
z80ef8e465d3aa903cc4aa31618fb521fd9e702a2dea1c52d216de755eb5dddd34e9ebf1f318dde
za76fef0b5a07a7762db1e8a90c60b1ffbb36cd16d07228e959e64f3ba54711a5273958b74c9ca4
zedc8bb8241c87a23622511cedac674908cf9dd7af14c17c5fd5b2e7731d16e34f4503809324988
z0cf37182e32a409a83e908d8181906fb2047884bf9cf8276bfffc3744c515c28b19f1ef8e63ea2
zbcf180618f0eaf9c53b01abc02dea3771dff5463f4c30aee6e1d7e8411913915ad2bb8d4459ebc
zd86ecbb6245bb954befce37a15ab591db829f58f48aa88ff556370dd865440002329d1786e576c
zc1bede246c3bbce340eeece8a603e7a03ba323d237325ed852566a55c840a07530e3ebbe8ef75d
zcd5c157e14212fc8d03f631cb697ce8914378b92c35ee88af556ed131996148ff8c53a8f8ce40d
z7fcec1c0735ff6f31dd9067398ff305d01e06556dc0b048969605080219a7bed57d14b2edd44e0
z2eb60e62e6d3f183442f74e3ff3061ac9b4641720c17864423c071a20c2e1752757163c6ed3150
za3b5008f4a0b145f78ed0678d1bf587a83e84f90b82b48f012dfdbac42548e19f284a19c5dbd65
z9127572cb30f6849b691fdf0d071685f7489cf04be1389d9a426ccef559f650c4b3a48426ba511
z14fb7913c9ea6cab79e83e8a02023f149eedbdce3e5b69b2225eeea812a88c284fa9d6205a48fd
z5e6b94b8f87a38c08b30c0a4ae665430415e49b88306e1b98ccf8ebd9577e7594f11e0847ce76a
z42d6d4b737c29edeebe88812962bb122e22bb78b07309bfb16736b9f8726760b1b7c7f93818152
z671543291edef59eda34bdab37db7b2e698fe846b036310bfce889ff8a5df5e92580d9fe848458
zf246e14f1d8a43e2898e2fa6813012962745f96ff76238fa9e0802b18bc47631db115e080caec7
z5506691e0c6ff3b9caaa53931b738da8c565db7378210266446dea3fadfa9410150dd10eddd1be
z5d3434bcacdf3cdc8859ec7f9879a175e929d1575ad25ed5755c6f030d9195c06129f0c102952c
z4581b3a2a4fccebd1995876569918eb041d9a9c17984d584cf82e162673021e045279308128b78
z2d442d6eed374a169be53435b3872b78f6906651ca5d050d37c52fd3073242bc8dc4be3b1452c0
z079ebf415d46c52913c45f55a6050506e0de98ee3e45c205093147138aa8f30999ad07d60cf56e
z794dd037874272e9204ab8d903a8537bd9e6aacda4ae96618bf687814f304d863c7e9b52b2ca05
z88ddd967d8e801246d335917e6c9486045e5267d0d3471a954c0cf73c351a65215ae91c0c128ab
zd0043cedccd6f89b07e35c551e6dcbd6887abbb0f9df437f5e669a9edb17852353a04b2a48969e
z9d893f6302082b6de1732c6d68fe031416378ca134e29e03fe0b7fa993c7f2bf187dfda79d2575
z21e80385132d636cf7e1c40f5db50e521db84358db6ab505d8ea090289d76e7cde37256050fd37
z193f9f4e6369daf0f1c1fd725d8213db3cc4a0f9100490d5627d89093c1eb3138b14b3d20db4eb
za4fa49c30eb7ba805e3b990cf7a7fb96c99e39220b1b3b9d67868a34168a492e3e9425023bf2c9
zfe7cfcf58ea934b6ef5918a22b91ad37a261dd8ac627a67ce1ac44b1722f535aa620d5d0fefe13
z9bf88535bc5eedd32a5ca1c4575214afc7c212ca4424c7651ee04c63ee37c099603653b3b5046c
z4ee808f1654ed0ef7d0d16d3ad2cb7a53b066c2571d5f9e96e27f0c2553d09bce239e03ed54c4b
zbfca7c497381f5e5811e28c6dfe1d2d36496dd29af77530d994bbd633542e5540b5c38c55128ea
z4088aac5dc2c947caa9a688988e519f2a3aa7e089fe4b9a8606bf65189a3c2338c6b6a30d9abda
zd37b8073f3c6849425ad5bc2a74ae7fc35fd3a0a1623d3e8b26b4901d48d974c0bb949cb93e150
z73ca69fd3ef87679ccc46198ddf54c1f3b54108145b5267f84a249355a3bbbcd24750364985f62
z2809fc38056fab98641b2b3ae64f12a7d09cff5ca915b0616349a38f036a7c3e27cb7ebdf07fb3
zdfaab3e088531367aaed9b050228af34de394a65e3fe59b9ec0ce686b93a7dd72655680758e3ab
z453e810c04cff9fed00f23d0f8651397a4c187d74cb3ac65922189e9fb4759d2a49ac59dae0c55
zc7286836f226c2282382e5adeaf70e87e237d2a6bad50f473f67e7e31f4bd4a76d7ab6a4b66fe3
z3d1af0b138fc2b3ee57a7519785cce37f02c42bca6fe8a571016a54426d1460b213f244fb09f5f
z231592951f1208a3944a15cb1bf49ec75af1c7c08108d953c761ce3ae5e9859897bca61a07b622
z7c86b8bf31a9c33d3c9921d2a7c5d926c1c22bf8e9d88230b2844a947eaccea13d85943834dd6b
z855e611c5c2ebb009d1d898b45d6a13310a6227f4853dc91590a444820909d40772cf4154d1db6
z53fdff69c4e2d146034038490a29653a3bcff2655a9a0755c017702e918761a6b66d57f0dc1c24
z7fd786cea2f927c3658550b99bdfaedd34149d35c0c129edf5438fcf8a806d3dc9fbf7f35b471c
z15711629d0a7762a787bf60b3d7605ab2655b2afe6c02ec5cd607da818654bc0b454d9cf478981
z24d9c79f7d9aa2e21cb5a2fc60c6f4e9099fb214191b8fb19622bc53b0ec3b47c3bcd4bbfcad2d
zd0de2d7fe971b4f0c1e9a19c807f0d9a932b436df61cf30935bb11c6e805f6b8d4039d0bf6979a
z124237cdbd987b1f2e193629c465be2da3f7ba02a8dafad1631a8ba39aeb34817d04aa06d43c0b
zf144717cbdb8bb20c7eb6f0939657d311d65978ec93963bf18f8530aa01999e3f68e8e289bd7f0
zf55083f36185c322f9992463ff6f809d7d34fb30a0f42eaf018635e11f96abc499f418576d3fad
zfee1e3da94e0cebfede95de90ff278a5beaf0f63856a1951efb10cf61383ba18189937e9a76689
zaf20bf206018890d79d716887ffb10d5cf6df4f4e9b07293f64820e07a0f2bca157bcd7ad99b82
zf635f653323dc2e0e7a13a9e2abadfdac39b448a5b368d07c167669ddfb99948759b48995e2c66
z5c649318fd11cce8394a9867d80e043041489c1c0fc68a52efe4f45f90373004ecbc876719fa73
z51706aed0e191c874a03462b35bfc3402cebdf8afb2f88d2dbf44a91910c3fa232bbf7719d512d
zf4d1657e33ea3287ae89254e46e2d4e1c49e72b02e10b14474cc1232638bcd78a190403c8a2d61
z8dc355df073225761bd52d8d0abb40c22ae104cf6f4e8b52f2ce4d00973098c61834cb20ad157f
z708febe87ab12b6531c3e65443f703be948ae5c1e5e60df6e93df98157e6499b7514d007733336
z9c0238c9bc294b5b19be0603d3e3fce39ab32552e1aec5c0cb92cd2488724ea5066062a34b24d4
zfa3fdb08be7021fd13e927b048fb59aeba446fbbf160db8eb8d0aa1d07b4d0a4f732ac1440043f
z143ca7ae858099b9b47df6dca7a6ec3524259cddc8bb5148933b614b45b94fa382f0a1b18e2179
z31bce505397a80f83374b7fe800077547e6b874ea1e1133ed2626b591e705bcc4946fe37fd707a
z84b24c66249624241a69bd4dc94c95e71c86d41449c2469719c4a41dae79a01f357e4a917a812c
zcc770975578f0e7bcc4de022e69bf53c011088e807aca86b0c463234c754059ab5ebe46e63e9ea
zd7b174e5a7b72d1fec3873fb77318e50dcfb8c0e036c5e5c8c610c302a8da8013c557346f3fcab
ze2e5c16bf8259ef1b8225fd94cc91e8ed952c3e153e45a6a931c51cb801fd347921a5a58578aa6
z21963aaf2eb2a360c9530d6d885c4ccc099bd3de6ef1406e1d786cdc8c32c9d6df0e5bc798608b
z866b47470f46d5dd994530a82e1f4d37b331c1413e16341ec4ed0146afeb6685f67194938cf09f
ze61b92131d47e7f8c381f2f0d4ea67112d3b84b32e91f14b358acf8f083f681a807bb47168fb99
zd35e6a2485a5e1a5c11ec7508ea4bd9f1bb22d4c8369383ac64af13207b31c9b49a59d015b69be
z97bb39d81d0204fa91652cfca6802c2bff64f333d941a8f5a1adfa61f9eee77a685346b09c2716
zd77c415f51fb3529e751d7073af6fb314776566f3c627a518bae5cdfe343ef9e50f93348a574f2
ze59c2094cb080dfd45eb15fddf2d9e7d8ea1a450a74493cbd008274578345c19c6da7854feef09
z474135f3c997d75e2c4b634aa34130de14e38fd7b92990db9c87f0da1ea7b652c24aed0c3de614
za56f8049c1a5c50a7dd7699f167366965ed05917425161bbb8e9270f3e4e2a343bff3cec4f775f
z6032d805e33e658049af504ca6997549b34e4732c4cb2dffcad71d5bf48d23d6fb6a4e011f6a58
z827a6fa2eab2bcb1d8e0cb53ee5530263d8fdba34daa4ff1e38ad96368e3859fd6eb5b8270f48e
z567955f26f9fb51514d040ee610b42484aee5c206f117bdd49b644a75dd430d9965aeda7c3be30
z293e4944e3aa5eb2c1f8764dd1ff527ace24a51fd53a9c75bba3efad9130251113dfb556702a36
ze5cf7adfe6657f3916dada02ba12c06f9c304ba0cf4029acb8aacff7550c98a4e702a13e08064a
zae9736a257b469bb287b1fc3bf2a37928649300ac6792248e21eff4968bb8717d10f9261b6ddb0
zdae687f194105a0a17714b7c5d2edd9a67ec6fa9dbeb19d6e1e1bdf97671f25bea957240ac08c6
z36b8ca3ccb9736d236423b7e2d7815eaf5f0bb2429500bed402bf00aaa21a9d6dad18dcd4a3c1b
zed99f280b26b9829547d7504d9cb641361735d02426c926274b8e438cd8ed13728f9fa4201ae3b
zde57c344e7ce724fcb5e5a4e1dbe559886b01577ddfbfa35689646e50355482935349c2d4ebdbd
z9efb20db6574a17b87f53e6143f4a628ff31e79ff995ab260e45c19efe249d89a302838ad93b05
za8f1fcd740a3de575fc15539ea224212fc2efac42ce580e11b7d0100ffea689d07d6d4157d6105
z61fe035735b4b50cf46a421b166c1b2386c11077df3da38d0044be31804d672278d01611a66a45
z6f13bab402efbd26cf164a4a1a14520313c6f5038e8fbed9314d1846b8142dd0affdbcbf1e0334
z31f491281760c0a51d00f4cb36d16820ac419db9655715b7f31e03826660c7b5f3242219eb33a8
z0fbe34815ce7796587d3faf221f1925ddc8f10041c71d5b3705469bf9ba95b1cc23472fa06da03
z5a64497695ce4d5df07b28fe08228aba41209a14848597d3eb29c7fedaa876ee7e0bad2809b136
z6e3a91c1da4ee0d1560e92cbd9ca1ec082f0ef1b3480382813162324b4182f1eda8b5d8351a4ce
zbb68718945e90b52cf071a46e0d34c1f187a15f5941a36971da2dadbb9a889d2640cb68b63e602
z719eeed74e5729861403598df200ed9851cbbf234864172b16040479a9381e9669016f9195584e
zcb9449578cb48dd6f7c767034af2fc7cd279c0aa31cecb8491cf8c97ca5de931164a31d4f11a08
z0204c5d27f8e6c6c9f772db4f5fb4bb53b047c4c518beeabb2509c9b9a445348c5addd3de05733
zab90c3849aabbcd84de5d902c753f85217914be9886399c041daab7d6f1b3c6a56de6025ba0958
z0c338397fdb973808e78d7b7d12364e10607149056f360d590e58a40918d8ad848796dc198425e
z20956ad3e19a82059e539c61899f678b75319a76f3c90c3913dd3fec480e46e7198bb1bf73cf69
z40b7f0b83bb1275c844ab72413f82287c1243c11313baa5a94dd6bd17db8492961ab4a2afeb78e
z17b0e806033b19a7853c007325a5d9909078fa04ceee00f909c340c4fc7bd0cc3e276b2f3811e6
z596d79a70f12951c29998af245ed9e43e0909d7b1fbf731fb5beb9f44e57cc61e521944c8d03cd
z4bdb0e646d7fe04142b9b661d20a1c57e82e9a830abeaf39abc8213259b8ae1093045b49bbc3f4
ze5fd8a7800af7752acd6c79ce535f8016a573557b505335fa19ac3963472c20bc2f7cbbfb104da
zc31200774a64c2482379ea86b0555e154cfb6aa9f9cac89e1ddb31fdff90b0b3d50914b5432b9c
zb7fb295a129d86c5f550601ded503c94d6d1fc135983d31d2d485b129a7bbe49ac270b50a53be5
zba73bf07ed677c4bee8ff9cb78776dd66b1d0f9384190738b20e155c4e182fe5a1d31b9469f393
z9d4472637c04570c908a911ac6a9a96faa2600e544b433015d28100b986d331a758a25c2041c65
za3ad99e9b118c6c6386aab4616e7e20a16fc3a4d912ef0611a18327921b8c56029cc56e231ff36
zd617d104eb92e8fd11f6eb720572da8a30638b40c0409c9a6e8e33a176054668e593ea9bec5661
ze8ac32a1d26250066ac1a681d18b8917d3daa35918a774acbd1747a3985ade16af02cf6c8a323d
z8f9e7f62b6be56c4e4ddef17b2f6abe86a03d203daca3567d2d8c05ba7bb56b93bbee3922514d4
zfaf9849d988d0d66115b7c6f660794712fd282a1619f6bdbf2b7e28c119f562b917cd1b1fa0726
z963016c81b77364f3919f9411eb7083d51c1a4d82b0572d2f5849155f341377691ed048bfbf13e
z47f77800f1e58c51b8d9f8ad224995154f2a8b5c81dd26f49e4115a7e21dd7728d2fc1d5dc1406
zd71bc5a42d67023be2903a445355a7cf53854893560f6e1b347bcd245f3776067a6e5bbb56f649
z1127c0f74aacf4805d1aebd99c8c6d83576146fdefa12bc8e41f34c89849810d8c51c27f95b10c
zaf973faa0129aee09eaa471d7cf44523b86e04ab16953d07f98f084681e532cca75256a4b94133
z9946b10ed9da6e64f6404f280bf6f4d5d14d6a8e3e1362f6ffc8004e4fcef715e4d89c61d7e254
z9e09925c26c569dd9b5c0defb29a0f123ddfb7e4e4b93fef869fae3e88483363ef3fbddaf5e7bd
z6e7f94dcc56f14179bbc3af52309b86643d2fc52655ed3e5ff16e729c8e076fc61055e2ca96ac4
z820ccf1fdf5c1953ed2300e6e723a77ea4d19fe5aac92e97ee702c06f6f46ab69eb888ab96efe3
z240d143b58abe6ef8ee8617976c84b678b80947a34a84560d370e8fe822d9ef77622ec3f37ecf7
za9913b465d16cabf107216310438edb1b3688bfd2b466fa2299f181bf329e868df61d3f89fe32e
z7e3a64d209fd44b79feaafa8617a41508cc92ee747bb400cd03f348f620fc91d29fb76faa6be85
zdbc8a2c598716efbfc0dabde324fbf7800cca876d9c664f73e268c185f217205977565fae48912
zebecf67a28432571a6842dda5a9c805030225120ae2f269339363a4731640d1eb4f14941fab542
z34faa08f78becc8ea45c19cd3d0a179621c189b1825d0b0a128a91a4c2e78ba4aca37ac27cd2ad
z27525cbe82d301239963b0659fbbdbcc59776b2daaf70608628dde90d1a36e732c5947f77b4328
z6526876582b9e1db6b4e2af762f63a28a6e36f5d728968de6e5858566bec5e2a6765fd57b6783e
zccb90ac660f795896e45b939456fcd7a3fad2931ed97d18c4f837ccbc4e29dd363f280647914c2
z6acfda2de7550904be68ae4b36ee40a525a7b8341b2a3e0193f01332858ef45923c2aebdd8c312
z96665ae8800110b3a3dff6fe2436efc70fa426e8c0102cc32c54053793504f5173c010a052831c
z57b74f93e716eea6d0ca82cb71df895be472e625585a8fb4a6d931ebe91b27c851f6fe005c8d78
z9e46029e264b78b0ff94aa25a9f1d9df1133dc277d5e11d8ed14f73f0b446352d177d71f835d75
z839ed19f47ceaaf9cfb4c8ae79b31ecf269e9306dbb6fbf25278646dcd7cc3e5179d42ed6a29be
zc1af5dd5e0d52682190fe51f0bd9d1dd353ceb1e773702ffb8a98c96e3fc96cbcf7c1199c80bad
z55eec2e31218311f6e33397a4a08e0301b173b1bee4393672bc066c730218c36837b7b2b3f9eca
zb6daf828c99f5ca3572cc7b650eca105bfd79d9677e6f6eb2725a38590478331080426141294e2
z52f1ca729bf4545c9c45811c0d1ed965b5cb691417bad040e239f87b4c7c988bf9fb9d2623fae3
zadfced5990dddd124a313b0eba09707a14447f295597967b254f105eee903f2bd913f08771849b
z620e48c82e2d1431b496a994f01d8258b87a41948694f7bb4f4bb92c32f5e68c7e46290150db3a
z0db5abf7cf788edcbfe4b09ed19f4b810279cab71852c2ded19f3fdcd7c54daa669554f50bc3bf
z03478ae5df8b947a6bb559486c6a62069ab92b77a3f082d3d390f49ecd28aa27ff83b1d0e7115d
z3c655380e6f4ec12d789bd477d272198783dc37e884d41b5a23daf1865be4d8599528f76995f52
z1bcd4b5b701807d5cfe76f1a0bd65bfee5a605185046738b2190989db88cce6f7a22f4d5b5b866
z72b3b8dcc36c22ac28efb46ead51e4d9ee6b1738b6a3ceb97042f3e6fe10baab5440268e88858b
z2277a8b4aaf18963633e21d334864f1133ed27e520028d3b14a6509efe07f0598764fac734cdb9
z307aac8768200479ab386b10bbbb7d75011318dad6bcfdb6eec8ba0a02b0e20472e009228924af
zb270fb2777ff1e65dbec926ba77abdea33bb3385d6f36c8c4d8a2c7ac1c785e4f3bfb2e8225e93
zf2d8f41518b0447f32e5a5e22576339ae3c6a2baf254d91739de108dfb5ad74d8a39183055f0ac
z0e8c47f6442b5e5aab7ec4116ea1ff1e768b09e1d34d43f37bfa629a0c61ccb628a329c0bd93a0
z44426fdc8ee835701419dc1562af24fdb521cd9c8b37c85a6d07ec14a91fd232cb4d12a1573064
z7f88585956868e04f2ea7db8f07dd4a3b331c705327dda55ce859778be1488825d441c38c26f10
z79195342746d601f9e78b8e11e6bda0207abcaa5dc19f12a9edef09f4f8c8b86583e081c2d36ad
z07b85bb49d4aa0173090394c1bdde6c1af0bbe95fe7d5ebb966bc5aeff68fbd758a75906e8cae0
z871e717ff312d5a51ab3b13588c3d60a822ec0c66a8cafd28bab0f32af8b58f401755ef2ac560d
z5a44ca0d2c723e54ed008bff8ddf9ad62ef657c5a2c3fe78909a458a02feebf78fd0cb1d9ffe36
z18dc94c1e6f6759af1abcb0d473651ebbee2435b7358f40113f33457664cbf42dd3c9e4f47a308
zbc9294e45192459afa36263015030fd9934435d4c74770396c05ec7e87dd26d1a5528d80e2a731
zfc9396f9ee7ac444c21bc3c76ac56ad747b2cbaf3c2c94f1cfb6da33e5c3d1117cf38e3d9b4b8a
z6392985c44a008f1ddb5535b2a6fa2593bdb5bbc7b6fda0cbad9f6ee3a7b94354997ca56bed4e7
z7d3cb59af1726f2d79f1b93dadc6820b2a74733d8cf162d4b75904e11fd62f9fe286dc29dfb5e8
z06cee58f71317ec315f0dbc3c7bf40d30acd350a2d6e13673a9d9e19034515b0a5f943cfed9ee1
zace4038bb49ff2db695adf469f95a64291905b19d1ddd116a6d0a51ce8fb7701e89dcc326d23d7
zae830e8a061e77c4ba532bf1442bf421e0b8b58096c47cfc9dfeff871700641957de24794ae61c
z8510a68f82fb800b5083acaa89442af43ab0ef87b958f6439baa04e0db3f62c17eebd39c599581
zf3e747377faede68018ccecbbc59da7c16e82acb496e62f7a8d60c8c6bc70fcfbc4bda05d3ccc9
zc5a3478b749ad4cf8c9864caeef0f085a7c3ac52bc0e4b54ec2adf56327b938c895e2c08c6e4dd
z615cb9b4826ddf42e99192286328b8956b18b39ad0a5a1c7827cd02360aeb5e18f2cbd32401c23
z857708d2f7c9c2fee2a90810aed437f12928dee8ca0e47daa76779a5770fc4801a1f036165ece7
z54d3f6dbcb5ff066deed4ea0cef59502894435d4a3add2998e8e6d6cc37c1bf1447eeef542b541
zbaf5f2e2e9fe1ed0f94607c9d1944af6625e48dcc35e87247bf439dbb0bd8d4aec124f07dfea7e
zd20656c6086c2c25ea4f51f8bb847dbcb38c0f306c88882e37a9eb5714a867eb8e3e2cb5ca6902
z0ee997fed43933fea3197dcdd244a35839f62269e2eaf0a8ad20f04d34c7f85abebf76c67f25a9
zbadf66e7290d2937e832c826993d8dac9278b0c7b71c7976b7203c2a31bc06753fec37c00e194e
z64f81e71472f7be06c5287b9e282a974e1a3d18029df130e14056d82ad2ea4bceeeceb00c4e096
zecc8c8f2c1a11cd0ac7ab530162531e7db098003662a43f7aa0223ad5239a71de9fdc28716d47c
zcd8652038fb7e48f33df1587d9ae44897bbcb8aa04d2589020472af0ce5f2484ee2eaa14fddbd7
ze545e81e54574d46c41bc6e34a7145766c77c6975bdf483b096f54e09f4fb579a7a79792bc8173
z6fbeda37c7f2af9da0b7886cb1778745085316de902a8ea7e861b6f4d7c0bd61d389759905fcc4
zb32fd287685a191032001a64f6f22cf8b9434adfc544f86f1c6d1edf00fc7fa743e65e8a1cf39d
ze4b75657f5ac91bf1c850afec594281e3a4e107d789c5738e59fbd88c78faed66a50fa4a437566
zf1e80d03163e96cc7c6937b0a541d290a11634aee18bc9d77a9fb1992ff0a7a5e286ed5183c76c
z769b70af0928939f7eb1bc5a61bd1d9fe14a788923719f652ec38ab779fa1e569815ff0cd10d6e
z6d7e1ec1decec508ecde4b7f2d74e61908e8bc6066de6d3a1c8161343504afc6209e2808017671
zabfe0d8313bd16ab7c0c62d5d5840016dbd91474ec4d6beee9ec4837e97d60a77727798afe8d51
z808015e0b76a3e552db5c87841b35418db661c822a5ac59719dfa6ce6f004b8c278ccbfcbc95ae
z6eaf6dd79da8bd8b6a2f8bb29f5830e8521b7082da9c01d9411a950e41565eab1ca58667fabdda
z59df85a7e130af6a241d69216dd8593c509859d49aa9580ddc0465f81e5b977f5d9461c6946666
z5191fea4a192909877e0bcb34265bfa1e8fb9d9e837325f04d779fe83048aa453617a8c49f84b5
z81d05e8b2c2b9ee24b1e90e34d480893e908ca874bfb8d899317eff616e06a1a5fa0ca82ca1c35
zc5f3ec8090a73af358b3b85e172e605eb2f710310cd35fc25991d10ba6134ce687f42232538676
zf5f748d588a015b4bf2283a6b3a03ae8525ec46b9556b79c2729faec6146ced80a2f9d5dad9cb3
z0a37dc00a60525538c8b6bf700f3228b4397994124c10326cd97ee1ec5bc8ee7eae4f373aa4058
zc36380ff5153da7125d2eddda794d0718bb68c3613e2755bf0f0a2933e2f47c6c6b4a8de47f033
z71b41a9f44b5c624578ccfd3eef21bbdef76c69392b5b75cb746f4fa1538eaa3a88074985018b2
z11578b52d04513bfc6c15c024c75c7ec64b114ca3e4afb279c91a4088c665e14d1513bcdd938e5
zc6dbdfe5255bc2b36a5c239e2d30d302898fbdbc7db1f540a0373f6d189b657ee9263d179021cc
ze7476cb5171eee8f19adba2c3a810fd2f520ef7d74f52fba47d7abc945cc5ec62b5780af8b18e5
z94749293fc4615573aefee6bb1c6a2f44777109f9b0c392195c92281fb741fda84ffa5290cd7f9
z9cd6d872ae946f8d4db423f1b9997b415675cbfae570e8c5edeefdf4df144b0b1e9e956ba30416
z096e69983826be79032fea6d1d6077898789325ccdc9b7cc509751f1c171053f758f6a0ef11983
z678835b6083065e98153e9df2264896599b1b24d81cf35b674bf003c338bfc2029c50fec77aab6
z29f08a37b36eb8825d101bf7f31d5b2efc215477781f37b84cb94acd0f649328e3ec7da5dcdd59
zd0a700e6872274a4cdc932a407316a593e19ec0a2732e336fa91b81aab8aef1f0d3f497d296386
z42107a73e712f899e18057ee4415400bc8d7f242b06f4bbbe4116202f2f37655e5e750efffb9bb
zacfeb5a3173fe5edd9e9f107ba0f6178ce638592dd60d40750c669e1b6a62651d8e3756570c762
z30a1a48c7e8e9a22926a4fed4c68970b0b86f0ed3b3848e34e7bba3879cf065c7d8323cc88af37
z710254a6f9f1ca5461bcded0988e729dfd95e313e6eff5d3a48a82b7232f216325156a835d4bf2
za13b12c57b0a508571134093a3b6e56648f12d9534d8cbb021ecd28661ea104ad4a9dee33822b1
z9ec4c781e9e6569a6e0977d03c39bb887be3e785f330a1dc29e37cbc8dad1ef8c5e86a26a88f47
zb6aeb82e527bda8c7b7dc46824705eb77eb0e096e9f167a63352a08d01ab2e003098f84c5f2f77
z8e554f22d84e4895dfd8df088d676494f91cb5b82268e992a737bd8808a70189986735e17898d3
z79e668c9a312610d9e1a756c9ef1b4e9d9d59ea01e564f5f9f444f103a5477f569ff1fe8a6e471
z3f2ba5a83af6858bff20adb15c1b664975d8f5aba46e272bdadac02748d60902a041ed67faef2c
zbba964c7da3e1cdec563168f03fa60c8ff9e14fa44384c49ff493c8792631f0e1457d869138a26
ze91fa01a0cee89a46e807314300957247cea686e35449152b98853fdedf19dc2874317142ae96f
zdbbba2769dd165ce96ffe0e1e03bbea801baf6c186df2c603f4b268f2671dc8e76f6f24e75739e
z43b5bf84b014de1bd784a1857c8662f39716779018ed16fa654cac89b3fe7c049d08b37aa760d3
zcb2c1405b16dc2421c42d492b13e6889428db1c0b308f47c1c94d49b904288c70889626714b448
z6bdc00031cb1378cc420ccbbd806eb89bd42270d4cf97cbbb9c335f2344a89859e52694c08cdff
z8752dfb352fb1a98ebb70708aa1936c55a7433fffd0faa957b4db85cacaaf7122aeaca9d3a5d8a
z132cd237f87052a57ea1f56b55596f9f946e2c9a0dd1ce64d3cde684e509e789cc911107d8f4a1
zc1a0f71a68652369a6d05b5412faa031592ca4f4f51c546458c78465b5954577a179935f035356
z45b25958c98baf239a6160eac2219b6bb5fc9fff0244b019a2a0a472f627c43841a8c74a958785
zfe89905182844f8ddc5b5cb7752318062f171ddc3c57cca722202fa5d2b493c7995a4891d18164
z89b7a9f84687cb54eadfbb9799d3aef12558525071d4d6bc4ceaa0a3389a1cf22f880c8c3f2ec9
z90374f8be29bb7a84d095aff230887c4f57e963989612635b16ff9561e39ce6698a72bc70b627f
z81e5602fa0f3d3ac3a715c741334768830c81c92e4296ba44c8be75ff02c64841b5aeadc471159
zabc5a9cb866f0257d9236c8ff99629e1084c9ecdc77b8c898bf949e6fc461063e94dc80c6afeda
zb40543c045e6523e086751902e9aa8b15063e251f72538fe13ee60be3365f12044782234e36607
z0d5ce77677a6a96c16fe71df0d02fb1aaad91037bd2c3fd8cabb875e832992c6a81268eeabd753
z2d56f7ef7d2f898f8394058d8e2c332a0776fac6fb7dff6b29965802cefa2db287e98c9e882e55
z19a12069d841363eec323756da88423fc618d59dfec413f2edc52bfc22a748e83e164cbbadf0c4
z5a3b4161ff491eaa233e037a5390273e6e3649e0da229ce9c4b27b89a38ce4542fec9b0bc36b72
z6d34d309687fbd3ed0f57df3746a5329d83961ccb2acc923d03d1a38587c9875f2335d01e498f5
z0fa386497fff2acc9532d9f34cd13efa70bb2a7591577275ea9638f8403d3bcc83bd58844354ef
z2cdffd49873ef9e44f397f8a0607e94e6b30947b5b435491040612e18a7a2c777a674a7a6097e2
z2e647afb1b98c923f82338a3c3aa790e440db06899fa28e8b6c022d7fc65697e0d557009fa7c26
z9f41049bc3b12952cf0f0a0a6699f419ea78d7253fdc75cdd86f34f00290acc0d4d2d42cd57ad9
z90ba0f1b645777969f2cd2a193c95dbc27850e806578aa43ceeb75a70530fc04ad12b728cdd43b
zd54498025652583b196ce291e986ef4a42ff333c15385f83ea100885453be412277f5a3606ec43
z75cdd22c8d8c3b36efaaa116dd23e6c255982da3a0403a54cce8469d64474eef991590c6afe61a
zcaa676f624bea0fe8816a4d4ad5cead8cc65ffcc29dc9c05189ad6fc9a4e5638642237d89d31f7
zd768ab6ad42d17bb808c7287c69e674aac7097a5ffa9b350f3a95d37bc89268b981a637d08bce8
z196feaa049a782575a58471113fa2155ce50500e5064e39a6a3a87f44c2d4e20fda1f2b5f5395b
zb4e6472e1b4d3421d595e766fff8a226864e42244a11d23385c04eb44c26794f2f07b15c0db06e
zef9a9fbc3421e38c01139baa4138c1c331750085fd726448d75cb340a9d76a089d635ec85bc8ea
z46b0385756e81dae9239daaa150326bcdf695f8a9fb18bf0bddc24622a3aabd2c436d3f2b7a097
zca1ab3712288e9899506f4a59a426cc2d8cbab0ce769dc8a1cc5a782690d9efbf94f5fe9451e49
z296f5f4b1623bee97cb722b7f4e2761515de3249f5a203f7580482100669ea318ec4421d49f4e3
z860f28d78d37776457b0b2bf7d334bed0539ec85bb43242b99b6c99adf54af5893813bea191209
zc96b7f50158a12e066de0d490a12793c976c242da4602a7b78ec3a2878beff67e2c6c5d1e8c1a5
z3748215be336d7be6083fcd8f83c63d55570b0d104a7b747fb19d3854962590bd1cd98bdd0f84d
z9fa0ecc23021ed20498a908c429f5d2f050629e9bc0139df21caee80e9d661c2d47ba473e663ac
z36681cf632f7ebc5d759d49f67080ff947d2a558b193d9171f98eec7dce214c0db8e71324eb4b8
z77bb4d659e49a977e933c3569aded4a0fd11d24f37ebc1595855b538ee97d491ae56cd072f74cb
z9db97d853cc3bc4192013a7235aa0db0e437ac3d2075befaae3d0533da375c5ed0fd19dd137821
z4a8c8c142f4dd41bb173350857d045e2b18c9dcae9f26d0c036385161502ff41ca89e6dacc462b
z1b1ca4d029144dd6142d5a5392cf30aebdd8357467d1dbb177616d650ca6dbdfee7c6faae7d5d9
zd3d44a309d1cc8863354ad6be5f6f8cb43b581f8aae917276dce7546632b31871b0ea41d3c4f53
z4d9c42674556c7a99bccec845fb6e4c6bfe70ea0468f3d6697ddc7a948449fcd009065ff2565de
zb5379be79c9270f9a309efb58531e1ee210caaedc6017ac28fcda53fb0134a240d21ae4c5e3cf4
z2af51ff1249d7814357091c5ca05b5c52b78595e4671ff1f23e04517bd26d44df9751a494a66cc
zb0779adae552ebe67eda19640c653cee759abf35d732ecfa859fa7f1bd09826c31977a4c349ea2
zb2b641dec1688a612410fa8aedd3ddce624974f8972f44bce93ca40279d41a2d8ef4756d436b13
zf108bee3ac256e0cc0d2a5af561b3e89c60c763eea126b6ebae0ee9e43f2f6e9a69f454276b39d
z45d2ef5b426296216547fa00e652f02c722ad4dfb76518515d0e191182e4b1cf6221d14cc8a0d5
z0bb2c52724f658b08a9df0368a34e0f44b873b1f88dea438dc24e3baafd55c9cbc6156488d3068
z62fa3ee773c8de1077d7c250ecd241099f43db2e9b9a694a9b22f6774410be7e3ac19d00467ebb
z15c63095077b75ee07f57810769594bda3bd7230baa0829c26ad2f36266d8bb1b43921ba4fb859
z27f6219acc18b295bcd7a7fead2629ab11f9f9a313fb885c44908ba6ba11a76065af183369dd87
zf587d530f550ec615578b3a08ccb6f0b4ee1909f90f2af6edd650f451105a66a3e9096b36962e8
zca676e3f63d9106eb9b9020f374f7b916f56b694aacc35209a88288eb31223217a39a0c51a7ea2
z31bac100e718182a72846fed2cd230f38870fc99257e9a3f2f9ab57ace476378243a4d7de6e438
ze4efaaaab2ab3c108f2c4249feb4eebc8325effa76a9ab29d9672b5fb0e8703716f601f46eb733
z7ac04b7d0da184f8084d4a5a5e940bae2e39cd17f1627df4fa35fb7862a489bbbc7b1a5e4b47bc
z93189d9d795d4a4f23a2d051e8e9423ec667273aba4a3acd180d3d87bb172b687ede000fe069db
zafcdfc55b1eb827932abcd897ac84ebdbeadb245d2cbf1892a50acaf30fe89e5a5ea9c6de49f91
z9ffadb99b6d5e195efd77ec2f6e4baea04e7f96423deb294ffbd192ce9ebb20514ce15492c593a
z7812226fff9a607b7083de1ee62d7ea4019436849cedecd5454a3fa1adb6a0a5837f4be266b13f
za7cab8589a8577ccb9b0fbcae0279c7415330f63dd9d886567360dd09d33387cc8e4da89ce5deb
z45274080dba42b3ff9ac5962c4b3fb82d4b89cea91e3b45bfdab73e89d5e85a15144fd7a529ed2
z113b81deb5788b9a0dfe8728e77d3830d14d6850ab8dd8f63c6b57a7ddbc2353f331b050f24545
z7daba74073cb7965f6db5fbc4208a9572156c0defd3105c88f56c1eadfeeae74638bc25543c6f3
z73b5245b0098d8abcbddc5a73478e6cfeb8cd838f28bf079106446c4d0e36d3d0906fd83b88ea0
zb911b0e47ef732d4f01d12316b87bfe5bc3f86abb3007ac06578e3ffb7af566ee5ae609766082b
z4e6242eaed28ac17f03e9a06c63d222cdbbb614ac285e5069a0d8d3d13782214ef9fb3dfccecd4
z015e86ad5d545cf8cdc472ec2c72a1b7c7a98bf609e96a851e0c46535f65ffae126754e01eaeb0
z458dc79775752cebe2317b1a45dc54a830fbee92393e8165d123b7b064dbb7e3e73da32553895a
z7a7f8d0201787b1d7e5dd2773be6463b8b38f23d21bac6349d92629342c60b68dae75f5fd1a20a
z1160606df60001f437357e9763e29e6ddc898a6730d961956405ad690cb6124e640324b5963bb5
z59a4f1e251327c3964d7e208eb2e2163b6a8e8c46ae5acb1747383f5ace22481d2ad8ba3e584c8
za2f6e34cb785382c8bf1d8182f4f318678c413e6e95af51ba3b9ea1c9f00920a3f9fd8cb3dc5f9
z9e8c73eedd4c2d518901a8b2c30eaf14dcdb442822ee294d7d6c14b84c378711001333fdc04bcb
z214fc9cb291f72fe3658cc7e429139016923604442645d29f3bbb2c7e8b3931071dbf881b22d74
z98870e3dc47f71a28798715fddac93a01c174c702cd9545a89658b95e3c079f329cb3678134dba
zcdde24c344662dfaa96665c9eaeb54a64ae0de76474972a3ca24ee4033a2f8be1077d5d268ee9b
zf93f52d774bb7f48ae42b7d04df53721e18914afdca3c37c91d38053709b7a90b026773556563a
z5291ae798b24e7701926ab3b53073f253fc76b9db2c84870901a297dc7d4f70a9812be5d20cbe8
z39027963c51d4f1522ba1cb2152cd28564c805b2c271c0a93c9b13a47d63694b1b41b3544b28c0
zc0e3c1aef0133b8aa3eaca2f65b0635718f5d5eba14d6b622b76964ed480e89bceb7f8478bddda
zdf9b4f808b8cc1805ba34a076489fc7ed5534f1ebfeb2696dbfee4f18a4e1ae23b7754945b3178
z193b53ab0a6c49257814ba7b44fb454dd689811079a2d62c4e46e35b37e99c605e3bd187771d99
zcf08a5a1fa3f85cacf1e248747459fe1ea5cd8fea3c7c53c85de0b47b141931038fea5507da746
ze56d3e0c11e56387ffc83ba133c5b1f46a7036e0b842bd22045db061a7ea04ac3453a9bfbbf664
z386a2d25b4e228dfb9bbcecb40ecaa6eaaa7c64001ff74580e25ae15224821397711469a1085e7
z3437f071528605e224c5a39c649aac609b46e00139dea5cce8c09d5c0953754b1ceb9052bdf9ca
z13220b69e1a40f2736c36342c08b5b2d484882ff3bf820eb7b0d2551e9a97e29d9f8df0f4f54cc
z70f1cfe9017156d019cd9941e30d386582f47d4cabebf31584ee9acd3ae5c3418d230bf573e460
z6d4561b5bd693be3e082e4be46ac1bc0fbf69d26e62486b07049866e7063b708c41c58de5b4c33
z675a3bec28c522a9e50e1cf557053dcf703901a201fa60bb34d93a61b2efd2292f6e51e50bd6f2
zb708e42d005509203d3c30e66d2bfd81f158be9e2287afde48fb179724ef8052186ee885dad802
z05ada1478d5c396b5f447dd549f93827da086baaae4a2927f275a9b533b49922f1fac5d3ec2d10
z519353463f554acdd107dc7c1d3dd4aa8b704c68b4904e62493ad2780a625a837fbd026796cc64
zb29c28901f25fc879e44c0f3518e634b5c5d679ae02525eca930b4191bb1afd452e42cd19b9378
za5a743fa0fb8df9992e8842ad6da3ea517e5b027f993ac4ff788b9d339d20c7c735a514e0ff496
zb854c3426f3bbf8593c39ebc3f6d499cfd79ff19548e91db4d9788e61a546af0b0f14933fe8af7
zb072dcb29216a2dc62e46078fe681dfc6750d59188771beeb585fb0e70c299ff1739cc3f0b5835
zd1cd438cc50b7a3b34881c0afaa69274d08fff51316320bba25cbd1a733ff8259adb32d09e613c
z022a2d550b3a2eb35317167505b1223db030b4b8f13bca93cee44a9666089c4b7fecdbf4130b4b
z2203b15329d706043976498ec005a74d72cab29c29d156f6fb90d90b2a6ab0724524f1d2f974f9
z964a4bc3a1785a45a2aadb2302dcf9d0488f5403a4909693c0b6a7fb0eed4d5349e50efccda37e
z9efc4f21d015dd2fced13d85f99b02f0dd3a83c5ef540052a2a544a72411737deb7540c71f584d
z32156c90210abc2c83dc3aaad2c0e8004a6bde686b5e5d913a9906312258f370031d6a3d375cd1
z0fba1b2d76e08f4a198538def6868f61545117039358dbe52796aa3337eeb0477c6d6206757c33
z182ba17864187c9901afa366b9e0521f4952bccc374b2355cc2099e6bc44dcdbba1ab94c32270c
z2f8a62240a6b97a0d834351dd8899f6618f1c1db5ade85d121fb29575177a8a83d3e77dca2fc48
zfb9db5cf5f1b2736f03f52f78e3c3c3a4a5c76187a307c22da8be32eb679578ada95e820b2d576
zd58da5a0c19df4f7315118251da2075e8a8e3ef7acb770c2f0bf82be05ee5b275048aa14f342d6
z931e28003e5b00e6d85c2be7f7e637957ea7aa2c6c774eed28abb128b0c49ed9873ee3e666f322
zbd4a63043485cd124e8ed2db794adb16eca9daf333ee9793fb47095dff0f9ea16c0f6fe0162ebb
z28de99e21dcf28ac9aea552fb6a6bd6c68b2af134250b20ed66a758d13b19982495e4e924d7bed
z81153f05846d00d4d02312a02ff0f1951c9265b249c66ffea76b7f5ff1b0d8ba4c80932e5b3db9
z7e1024e523893e845611f8e672d43c610d411a80b165a765f0c2e4c2ab030210d4fbceac76f63f
z8257d7b3716c4b4a8684c16ac4154511d216a4087b8171a89b81d96854890950dc16c1dd407d68
z72d8b62a20212dfab00e022963619d31e1d2bedb6d6811e84674399ce57df4e139a3b9b45b6f75
z44d2fcf2f3c3423809ee8e5d35078e544e262edae371909453e29919eef1ac7bb7a9d9252cc96e
zeb779e32755ddaf2b3fce646d828011e14e97df17ce7ad6fb6b7b37cdc7ebc140811923bff59b2
z70dfcf80d7182e7bd3888f1d81053916db671cf06ae66d328f42f7c9dc4a503a3ca2144d72ada4
z2aa38c4dd3db1d9c54ee399b51d385649ff39a8ad6b00aacbbec180eb7bff7ffef6fb55a04ca08
z6718c6823d59e7ea68e7acecb53790f95c242b26fdde7532f6fb6bb3c3b5e9668dc9c6c658d2aa
z57a67dfe6412b03f049bbeb3c0996cb40b63f5dc05768bda86ae9ddce2cf5a356d770551d92a1b
z0ab696744cbe6f33a0ce2d329c1d50067756ca823bb841729124c5f1ac4d4944160be6d523c90b
z0606c224fda9c81caa2d42147686d510e32f788a48a4032f61c459b40ad796b650ef04a022c9f4
zf429ae9b187dc8b32d0de230c07f3cc229d41d1c96
`end_protected_0in
`else
`ifdef MODEL_TECH
`include "qvl_scoreboard_assertions.mti.svp"
`endif // MODEL_TECH
`endif // encrypted_0in
