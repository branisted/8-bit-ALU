`ifdef encrypted_0in
`protected_0in
ze74c34e226135848fe16db9ffd31815111b6d7fb642c521a3f628cf6da949865580b22efd062a7
ze90adae0e65e66a2c36a587d0a790699161455169ed55a01f2084f11770a774ec4c588039b380f
z6de9c5084882a40b79a175f5c2114b2b6d78b070cb806e1c0aa9258297f4687ab308bc470f0040
zb0b1de382961eeeaf2e279e1462520fc31c119af8f2b214846f56c2b3cd2eadbe4099496abff18
z15cec83ec4a77b868344aa20ba7360908f5c0de2a79abf8b3534b883bb12180f68b5d4beb444cf
z3fba8f13afb0abfe8fcc4294810f75afe452434d2d0f1166236c82f76edf1e12979f04bc35693e
z32ae028996dd85737a8f5adc1ebb94f39c940246e887647b64782cd7ab429b0544c173176cede7
z01dfb26b1f73408344a52b7e1f117f12bb9c8077b34876c2e6fdc085981637012dc9754765e1a9
zc512ce062e0b8fb16a214591f5c81e1353b900a611fe1f4886b57940b41b7f2ce99a7b84b04b90
z916f717e73bd10589c81e207ed77ec660a8cbed5b487fa50acde1b055c8870bd8676023f21ddcf
z9c98cc47cfa2d654ff1365d1f45035a045a66c5dfa8279050262529d2cac9e64fd27d9c7de62a7
z731bc808811ded9016570962244887f98fe5440167bd0088f2f049df882af501358497c3b28776
zcdc5426c7f52a851c35106bb93e16fff98478405cb2c034d92a13b05dd6952355a8276837fe1ec
z31ed579935d1f03c8aed1f61cb6f74edabb0b099810d7bc07560d8599c00d4ed4049381a6e2b8d
z86a7f6abb625239b7bba7d5cbfc5666e6b305ffb196abdc98f050cd1496e9e7a9b8bd29150791e
z328fa776ec981c1023a4a6b0b906d95d57e23d8183faaea82947c6a546574dc633563b721366d8
z282bf630835b168718286369a63bf7cc0c40b1d089917cb1f1af9ea18d48edf68b793358042a72
za32361b89fca7ed7e1db604dd37903e9f4fd587a9ff097a1b7e30822142d15cdbe595876a7fec3
z6b09d9b556be001d1a3426a11438de3cdb5b691cff32ccd5a632b884f86ea1b8d2be153f7a8bad
zd62eeb99691cce09ac48e8b75b0f4c085bd6c2df6be22bf9f2903980aee22a7fbd3c6264ff436c
z5ac914e75034810168d0ae609a433be67781cf78ff39a94d1f5924c85a2b4d1cb39ef047c039d1
z1f0a1b1cab662c6464e8066934e4bcc8ead51a123f370bfc5d96adbb4937f548eac50f43fd485f
z9b2288c38315812439e842be36a605c5916336da6c8ba595c206bdc7abbdc3a918f8f00928d7de
z51d98636c196366cb9caa2aba245d19b3912538cd8096cb4f36aeecabed0d15817712fc02ffdc1
z08f8b425db1e6194ce163ab83b616c5d70a78db2fddcceb5d3c5a3b3ba8a18041b0f0af7ef67f3
z4f2b3f0e0b2942d485b82c7b86af0ca80859e3128376bd4fd14cf000e7528d309a7480bb2b5d1c
zfaf06fcae634c6a8a5608783015423c60587c8ab7ce160c7f7dfe38fe98a3590c8e1a7ef693d51
z58e1f00c7d7ff8730b4b6539211f62490e4b8591e9fce7dffdbfc32571ada0884416bd36fda93a
zae6b589a53c8c43934179f4017dadc050d36c86990f2a2325939b531d7658f06de3b85ef4f1a39
zc1cf40c0758faf84a26d9880f2715d8391c6d84b48e4f7e7ef695bf9e34bc2f201a671bd9846e0
z662a5451aaf28a6d09c9898e1ed46db9548331dbfbe3826f2edbc6ae4851bde6438db61ec2fe9a
zaa5be9ec49802b817b3abf65b0e14e71cea0fd667f95e4fe7744bf9f1d482dd01c96bf10454356
z093c9dbbfa998ff65fd4c746f2c442d64e9c58023a710701322e15b07e94354ed048871d95818b
zb6a5fc078d0d37b389d01092793a6f1c77d07faf4a3a7230f2da4b37171793812b36ff4e06ff72
zca526dcaab306fa07bb7d00b9cc43dd373c587a812a52cbfdc4550591eb5f059e70e8f2a051334
z71d49f60571bf83c2663835ec475e40fe526a05ca1dea4e566d82d4943b7d59e7d39ca0bbe1709
z0ed083e11ad2138e865d7d054567efa85f56872ed138a8b65f84a77c237924e343c9468941682d
zd264418ca3047118de6c2f1123beb0f4a21b5816e58377949fbc3a0fa40c6ceb3628f500409b12
z9f215d82acf678ef1a1abd5a91b03d6d6dabae04d37e1a9c84cca3397aeb53b935d42ec60726b7
z412b424e7b491c17a38715292bd4a9e3ac80a0fc7fccee64b132d64d9d8d5257847792783e2702
zeb5a21bf494eb342f27a13d623391285babf4590ab8b6097974bf0b068da8fb660b016f9b1d3b0
zccf1b1326e0344c4026de8a23aecfc38f5a8b9882be757b8dd035084eca9b65f2a4fe555cd84a7
z1f6e7ebe9c0e78c60649950275688cc4f9951dd8d7230fcc59590c14973b52c8ee108192135d78
z1f71a165aa67ac24dda893364dd792ef72c21da8fa89650a4f25f37554c727fc2a826e4c6db8b7
ze2ff2d96cc6734ac2e9df14b6c801fd39e225f1c963299705ea0d6a419bd5f96e0f52fbc76c74a
zb7ec076a2ce607887f7d5d45b3f5196c27ded06122b7efbfb74c878457abdeb43020cf6f4160ac
zd30444c9de406d44b3461b4ce220728cc403ee2b34ffb72f7662a19f393add3e99664a509a9230
z549535b75ceaaa337508d10e2ba9607842c36effaf9267f1f21d2fd62a5201d92e5a5bb64e021b
z0cb9a733066a2d454176d094ce6d1d855145795e1b137c4418cd2f1b933b31357ea3df74f322c1
z271fa855cb8cf99826a9af8c62fb4c9a1eddfefb967fbe4707ded081ebbb9379e139530d1970a4
z3635f3251a502b38ca7c89841131b7d83a478473f879372a6fa3178aceb35db86e91359bd7e7fa
z3be35b14ad0ea1feef11522ec2720edf98f79f7661f0767c6f4e19fc3a59580b635abe2ee766d9
zfe6c907e90793b766cc651d859df2450022630758b501cfb0b6542a9fb4b37333393a8e21dc507
zfedab22cc7710c09a44121781e6e614ec4e6d126a34bbe05ce5eb0eb01095df87dcdd4d71adc34
z62a25d08c09893feaf0489f289f6dde9a3ba8d7053dfbea24fc365c5eea79fb7782beb706a2be8
ze8f89a6dbf09161c4efcf1d71eda220dffb783b0a948f2e72e09d3880d58944a2cd358b63c0a73
z1f88dc302b7a1840aff69add841aa679d1b9db3245bb7e2b099c288992736c7e645ce4a52eccce
z6a9a4f8eccb0b0c7b6deea318505d5d9154140529e959d1db80c9596cd08983d372641ff1ddbda
zfe83078c63dcdce47c58be18f8b778202708f605ec371b2a1b33efdf147ad1446d84c1cc40ac5f
ze2b39df521435c47f57e56f32ba1997368e14a1355475b008e07caa9c96fa62a7eb5b39851f593
zf1f8c0e688b14ac77070aa559eb6ad7a306837c272a0d19179e0c55786b39aec46d10632f4d094
z0ef262f8319fa477a21ba4f65b0971948c6c8771297ef56b585b33e59e10b4bfd81d0bdc6910f3
z9f6784ad1a8dd424d4e56af9d292df5ddb6bbb8a793d4b6a954bba02cd873bba654ece89042233
zd9f2286493b698292abb87b30df32e1c8c500dcc787a0e69cff11f08b71e8d8e45f057839ebf76
z0046dbafa3e4c989e23122066986f8bb250499fae8e8546e1a5d50c23cf6803f7813f13e5a2900
z6bcb9983df96d22f3cd608ab074c6c5c28882dc786e0f4bc50167345eb8b76076ae87c08c5779b
zb5fbb84fe1ed1158a4d3b0cd0a92ed0eb40059003644819cac4d578a63382a93a3dcac90bb694a
z84e67df357b6b3be36c833334492b06a5f5e3d266d3c9b111c7f808ef07bd004d24eca6a0f33b8
z5498249c88e5009077a5bbbf1018b32c6d82f21518ed8bd90932d192744d6cf4c3c71b55f91d6e
zeb03b8176d9e744040ab2cbea02d0e710b6d69f7123b3aea0c3f2028d67bdd476d25992a17420b
z108adb4d457f724b5415d8fbac942ddcef9a3188eb68997054e5f5699da4bb0337fc8c1e0961a2
z6366068c41d4eac826562a97d9624729034282d7efcbf02f508ab6afe9005c44fd7917a8226247
z71f130b25903d8b83797b1f223baf641410c1d945c4b0fc166399a3945760bc3183d4d404dc731
z245ea251c97757aa157daa76e41d2f1db018dd885d6003477fe324b8fc9553b1410a65e41cb12d
z48cf1c3f6409e1fe8faf6bbdc50dc5f92718fa11e1ce961a59a96649e68913af183bc3adc23346
zbaeecb8c2335de0003f10db8b18775889e7fcfd8429fb67526f38d251893728844f88b88d9502a
zc1b0346638fe1da6c14669073db9101ac72dfc2acb084619c109abf86b4620803c5b182c72fc3b
z9ba36eebbd43f3e689a136245e2434eea6dbfe5c1a99138932553546d818ce12838c1d26dcc462
zc83bd33154917c648e6ae0f9977263d8ba15ebbd0e517f949d7fbe484ac7a283f4d2c56aba1123
za44f1196e0ce5e13f7f2588e7cf3ce1c0a3475e8f3a2cbb1d83bb844751365f37ab902974c778b
z6137f6e2b9304d741ade0c5a4d58d2680daabd9ba5915735a4c2a3e12ec142c9bc24042a50daab
z0aae85629025d5356158786ad2b5e8fbe65dc5c25f09dc2febc75420110f2e020876a0cfbd4ea1
z18f9097c5633a0653647a4d1ed64f77f9ee55c00889d4df0b2fb5c4198719c70ca33f4ccc90304
zfefb3a225280392f4a13feda29c6d8953724bc6a3d7c03754b5edd3177adfc800ae16933d8a54d
z15208e4fe0d32e10b80c031871724f5845c9abbb98489d7a7d6cdbfbf5d6feab4aaff4fcdff50a
z1e9ba0647fcc296ddf326f817ba2ade98b1b072907ef7012c8ff7bc8b819d2e503dd51a81568d3
z7f7d5db9087f9dc1466b3253df59c0fa7506ea4e4bc369a71a165215a22e208680ceb0592560ed
zd3ea8d53f8c89f265393b5c2e6ce683bea8da6d6728c5317e981ee05d36c2fe8e83db5a3cd7d2e
z0a981ffe004280af4da2f17766be975ffa0fb845e456056eb8ee52cb852dbf5bc781a5c4ded27c
z6355b4743384152336dd5c04889f8d946958f6f1fc78b77aac403f3332f3594ca6af81e9b2f153
z2a274352f45acd858e8c2f81ea4cb05d365b3ac0f344c453fac1d1899cdc54b11fcd94dbadac65
z66d09303b35762b1e3044287c0e047a509419d0049fc5f3a51600e580133627ad540babfced7b1
z5d012ee6bcf43a9128ab4ce3d0f6b475fefaefe31efc8b564dcd85718584e804ae36002a3c3149
z3e72d7f16a59001d8ebaea0ece60d81c02ac3b69d4b76857c8c871920d70f9a58afef5e827e1d6
zeec9e55887c716a2f256bdb8aab109c8b9bee61331a8adb6c7a2b3efdeebd6a142798cac243400
z2528b4c200f6ebef27401a22eb702569159758c53d5432edb816456628b79e23c2eb4af8ae5563
zd5c279b7a1d5db88877c11d078edf5795c4f851a5e3be90becfdaa9a3c0d26483bacbf9d4c313b
z4ed9d0feef3c62e7b7783528b67469ba960ee4d436f4586c53da267d5a070322fba01f6726e4d7
ze4aebcbdeaa2da24685085bd33961ef8a0c013dd84d50b0283b789ed6872bd42a0c05ffb6a0c8d
zd387951c0c97419eb56a3aff5610c977b7541202269176b1491589bc95eca6a1022270c10f655f
z67ab248a2143ed09ad1c4f78d83d972e463f2df8a467fd82c4252114a48b98e84bcb438fff58f0
z7209cbffa68389b84d427b485e64233f6b02772afdf5fea25469e06d3957e98497a5f725be9e7c
z23c033f258013ad81975e1c9fb9852e4d0315e4f54ff8592577d783caa1a8e11a68dc264e0802b
zb057758176f69af8236e949d78c740501cd7669744a336c41ecff8d39c851b2af7323f2d2ad8f2
zcf0c6e8cb213888a6d77be36f593abc7642d112f579f77b12f4d1e169cf91aaca5e42990854971
zb30742b33cab0b77b4970da4f4d48b8ffa05a753a98f948df46bbc5af4156dc7e83051cf25d8d0
zc14ca4c2eb36c5f8852db91fc67fa85d6bd78849e693254018efdf1b503c6be0c0a4741e3975f3
z67692787140534a3b105c7d3819a750094652890dc721d6eafb49f1410c7adc3a0f45e8096afcf
z1dbc74e3e5ea205a9633ba9ea48286d3de59327e3f4fe812dce29db516022797a715b4fe0e65b2
zfd01e95865f2ee458d676693d69d02b031795030974e20e4197592d535317c2690cdf9a6d5dfcd
zfdec075e21aac4a8a2d28d504b9ab71a39810641386a7914cb08ccdf25565c46c6f01d5e9ecaaf
z82ff35dfaa97ab8aae9c7714c94875d4340fbd28864ea5c20c08e638c4c960e96bbd08eeeea350
z66a34055b1b388b49742f2571f44b37feac640fd695854e612b11fc6ccbfaf297ca54b81241a42
z2209cb30eaf6319ff2c4f92630f132685cafc301598fa2fc7c5944e1d5bc34865e388794b41e8b
zf59f4850b2a2d30d03d39a3581d4c356748f053b9bfe9409cd43b900ce5305e4a58c7b769c7e50
z25ee755100684bf75edb25883f1a1aa4466a40d3b75933b602c9590fa86dc576022e428a00fb5f
zfa76a59fdcd3bb02673d45c63dbbf742e48ad24374c541a12a47b09492872d6546d467bd128fc6
ze6d39b12162621a9fa58252baec007c783fbbf8b1298335ceafeda700514cf10e993129e617a8a
zb630ba1bc8afc99ecb0cc04e5a903e71780b3e27a588a58f03cfcf953c8eb06933e63bea0308a5
zfc0fc6dbd50aee666456f091571c6eb7b11e567a93578cd0ed98e486b2a527ac511b098437cdce
z0d0d46375f0613cfe37a1613fb599cf00fe9ed73acc351e80914d762942905cba1bde9e88a7c80
z803d1414de1c32475e630de8abadb0add268b42a04a18428c8bad48cdae269482338259f5ecc41
z5a86f39c678de376d007219ae74982b1a16a0f76b4e85192bb767198c312d0fc974fb39ff3e992
zf7dd141e23d26e03fac7a5cf3fb5d0cc6142596e52b9adc6ff68386f0913d459b88f79f5cf1876
z82dd685cc6ec39c25d4129fd934f190583b8d24421cad4490e00430fa9914fdbb7f371c2fe2803
zce56accfe0ad545d3c1315ae2a5d951687f815cea32a9ae3e9082f336360fa08b528456d7f322c
z66c3d3aad543fbe0809d175e4442291168274c50e98c7b9adc6cd93969f8224d2fc78839c658bd
zb7f066025743878aea3e37b3ae2318105af524a1794322a8d79d3b1ac4cd7d9670424ac2a3a376
zacd8f39edfb4a0b2ebab39b04e554929fc30eee48e045bdabfe1b80f91ebf229f0730070e098b9
z7cd56faae028a37143011742f594d2c5325ed5cbbbbe62f1452da9ca69186b11642d262300673a
ze1d771bc55e3ec8afc7126aea426b0ae08baef9faf53f249625d314eec2ef655af7633b25ed130
z8f5d0d675a66673e4ff421154eea5a14711ced2c29ed223fa0fbbde0688cf6fc5cfd4767b72bee
za472a106ca6290cdd391c4598a742274716a543a49298d0727687a64921cdd907ca056a7b45084
z8899a313d506082922862313a412e9d82518c4f65652b90ef6877806f103e80830f3662b42c44b
zc56fd32df763e0fe40aea09010977f9839ed6453800bfc0277864b1a3655152e0755d9e3b23d72
z79586c595d48834635f238cc9b360f81f8505c7aa8a2db394def95e8473087231388daa08e0595
zf74a0374aa020d7b8424365f50947a67f04d6405167b47293b2799d4780e8f7c7c1461c0e543d0
z3f77a7c8a67497191a183fa48b9abaaac8f131d9bbff5bd1a2499a6375e655ba7a889007a6e7a9
z92676c13a93822a9cf33a44635d126a06aa004348eff759de4188554ea11e286fdb5a487c5ea8c
zeb7664818d63a57e20047634dc358656a7c4ac1cb32d96e90c55c4df35c59765ef8c3186a9d5f7
zfb6bd8f32bbaaf1e52f7f621ddd6ae8610eb8eb4271eaba1e6773338729b0202705474b3645144
z4d954a5a0e1cfd53bd7aae1ddc59f53901fe4c818c0bc792f77b2af80ee3070e4b5be2b1827455
ze5813f4555297f69fc8a1927af4db0e014d2e9fa9a0b23b8c6c3ea5772216a3b496571f6da899a
z6055444570cf4ec7f3da7eeb0683988c68bdacbe897e4c9c5023ed4ea42dd610468a6c8e567a9d
z28c1bd1a1aa7e42692b596ed3ce38e2e1c17b050124aed9afef237a481ed6eececf94f6f758ada
z49f32fc38fb72b64e871c73524596825ab97af7c4b7fe8ae5c436affc957173c3c5f1537509243
z384ec9573f60e502d6d3d7db5ad369390d8f478ce46771944ba3a54866cb4c8caa36008f2337a3
z6817858825cf9ea548aab665fb7fd816ec4c2dc46d8745349dac93e578298855e775e2935f783a
z30187a69200bf057fac6803e806cb4c7a73eae0875930a7925c01643d015b0ea9b753c25dcf208
zb44abb32bf6ad8692ced2ba16c29051e302bf2f0f70c2589e499358dd0ebb5df58b0de65c21ebb
z0967072b954778f28d0d458600703f4a7c9bc3fd2c8765f57bbbde02f7b965f76fb217e079eded
zc2d42bf21c5060522244aafe7f8a5cc20394c34a90af1d163589f7e33667717b2e4b19f5c41937
z5649c022b4de0abd095117a20ded951f43ee802163d506af7e86e11cbf23a3585102eb1b60387c
z3e34622ab1163484ce1e89261f00b8ff88ba9077da2df591cca178ce3a4547df5376c164756d65
z1c02f2a120e9855ae761b47cb949677a99610adfc069a97119eaad5543b4259f4828491f2f8e67
za549859827a84eb1bbd03bc74761e3bd7cc36f775ee8783c67abb81b5ac5c542bea3607f91a63e
z7f1e80790f51b8edbaa9c95a3c51e7fc2c834400d79e37c31389eaf03a8279f2a49605e76b2867
zcb961d57c7b9dbdc6c327953303231305760c1c744550d3ba20f95b3e2e22b49376357a3797c2f
z6b8fd261047f6d4a7ecf9d8d46ea402826f01ac70c30e672dcfdb812d2b5db890d9b9d761fbd97
z0b5658087c025de0103e9051adba744bd3913f21c401936536a45677e260be0bb90cc4326aa526
z8e83d82cdb689a7b2889267522302344fca8665f85bff4cbdbdc3c763ea33def3f0a531990c0be
z385682c7563659cc682ba00d47140443ec899abbe4ec745e541e67f0ab5ca29da87a5905f014d1
z4e12d82a42c8527746794fbec5464edc34b31fe6eb9f8e3c4b072485b1be352e6635321fe538b8
z7cad0f693764b649325925c1a4769aea42a9d17609064922f2c170b244e42558598c0f8d37a7a7
z8fa745f63aa4b23bdc572bea0a66723faefd2c9d599737d9559c97c3c9408cadc0e6a5d35d328f
za1ade492cdc8da3f3bce7a6c8f774b2edac6e5841ecc99191507da4f25a57f0216542f6915ab6f
z9a892e317aa69ee7bed3161de54b43964c43a7087231da7ad17188cc49c2196607040e8b5f2e05
zd434fc4131dc0cc657214859389f47c31c0122986245977008160ede8e1ff404aea775e03e99c3
z2402c6073c6ef8a359e897c33defed53d374a70e6d7de22ed7658828d9597768779f2b72713cab
z74db5cf77905e34951b84c6539539b709c317e56f7599dfa1e6d04b4b9838021d1b68a828b3003
zf6976f5163851949bf3ca7d34d20f71bb80c1fd5d614441ca467c490aa5763663e25cf1bfa03ff
zd623258873b45628a1d7e83a9742ac0c16a42a085dc5356cab068e29d90c1eed426020da1f040f
z198d3f120d7825778d5daf6367bcba8015292e9261767333badf790cce5b51433275025458a7da
z7149b802fea519fab8048b4c9b14a912aa1e8d6d9c08e6bf153d559aaf8f205b0ee97c4bfcd4f3
zce880e0c2b3489258b162828ad36898c115b1704c4a06d68eb7288cb342579d5077224db623888
z8c5ad275cb71330ad01938844c62ccc2a2e5d491ef43d15bd315c52b226a9826364cbe58c48689
z81bbbe85b35d6cae17a33784a87323760ca0e9d528fe17e1e4a1207cc13b3dd8b09a3f7cf5e5cf
z099059f9b5990914fa7f23a287f3f45e418883390d9b7888c5858032b3bd51118bd7af90b9ece7
z458108a9d4cf0a083e074840b3e7432f8be040eb9462a9c89febaf9ddd10e3f6a1e63846f70a78
z51e31a9d901a2046594103d2c67d37f7b5538be09318f1929b73c51963f8848f29107675c515b0
z720b6b7dc4d85438114a60f1d4b687b143e21704a0aee988ace4e52081565a0efc73d2d0415830
z72ca3cae509f937bb58f1ec7ffa019340a3dc6801a2d5d5b1fa5e2ffb27ef419dd9a32496d3fc5
z6ed65177e42d6d52d70773fd6b701e463c8a62944fb5cd5259ec7308c0f09e5f006bd85a60e01e
z73aed78f7ec9200919fe8780ae7e1abce9a75caf7d70891efe0fc9763b78b0f8c5715b58e01727
za0ad8ccb1066a567986af7041dd8a2a70e12283f3c05d235dc047081f427747747fe423f2be0f2
z6c3e40467663f833f7ecef745fac4dd959175539132c315c5ef663e97614361fa06f1d67796bcd
z0e04bcebe1a0cdda49f8b4800e0d55989789c92161ed6c3f80381f7569bcef20be23e83201bee8
z84196cbdc6b4162c541d3b2f94cbaf8c49cef60481cac1b8d0b5bb05de8b707937a5da1e137167
z4f10810cf2d5f67c1652035708ce7bdbea6408b32ba3b99673728d6b5e59199203b7a0aefe8d54
z6865b34259864d08f2c52932d14708705a7c4f6351b4600fa1e98df9e0038cd93bb3654e48fd8a
z10934d6f9cb00f633819779a3a2c1a66f97ae239437330f71792680956e260f3126e38d7dd95f9
z0185069fcd3c288df435d4edea03ebee5618d44623fb95d37aacb6796cf8abcf6ba29cb2e36f45
z5077eb7b7019707df6f2d3885398e24b017b70e366d1b81a72bee87d06af38117c0cb98f49510c
z256b5fa22031e24a66a631b4d3e11f00d72153635c728cc989f921035e063aa6d52f98196c1d8b
z9c2f4c0ad850f80fa4660bb620e096fc04ea48be5099f9cd31bf80f854ec73db2dc9e3c50ea720
zb7bb11b13e6bc3c4112fdaf2f40ad36170e96095b16645524ac1b2b09a439805c2eee7011e2c5e
zfe8a1ce91add807ab5ee85d5117976ef53b162d59cf1769faef4bfaacc7eeb037301d380533c7d
z462035f36e68fff9867d9034531497760264496929c3cc93e079925e725139dd97a17d8031d832
z6b3398ee47d2d411649e8a1755cdb9afe59b21bc1574bbbbd304644dbf832291fdcd099ef6e2d6
z518fd02e6018e7e3710ed940aacf027feb40072b7573691675932bf53de222bcd7971e404a2b3c
z64da0c996cbb23184f8140f911fc913036d2770fd6a6cc6bc3640d44a00219d3bfc2dd73647d78
z14f12078fb66495a937eede3a3a288bc695b8102d0390bed84d5646220ec435f92802dea93b323
z4266459ec7e309abe7e6236d187096bb9d5981b9d3b7da3bf01723ddab01e0716ca805ee7c80e1
zc9b22ee53d05d6dc45ca3684c8a54cdf129019c8e50dad37956e0d421ea4125498dad34e7f7cbd
z33031e77f62888bd96df78306d95feab1227964279d8c316f3997f21f3b02ad3afb719edf2661b
z43f464ebc7c0e1c3623b6b650578ee1a8b6627eeb1b531368856a25109df7efb86cd3ccb637786
z830d12a77f6b239362fe60c37ed2756eb07210b17907ace08cc680faab1f907eb0d9934cb7045f
zb5321562b87474c0cc57bdfec074fbb97b033f03886b1ffe4e01ca4b8879d42a7db3d53f11127b
z882ef89ee46b728bb5e60c09497e828fe443556358a8f2b211b7fc5e58dee537cd277ba42d9e98
z4fba74c81646d087719613df1734fd39502f201cd67c4fcf472220f80323de411bb9f224b0298a
zd7af3e7256f2d32f3478357900ddae3cd4c57d7bf26f38bab3f9641333fd825cebb542c5ed7958
z9724b920de950d5a51fb47a53f40998e27839ca3e3f26fa5196e4c8d7e50653f6ed0fd06987d02
zc54d8f2776a003b3f67ed7c73ccc295b516df9a763d058a2b65674b946828a6c42234b72d20127
z771b150a290ed8bc2cf85b7eb421478f7f4fce82aab3c7ed0aae166bcd7a5ad759af77a29c15a1
z66f596dfb7263d1a4b0f8e2b907253d9b6a18042e12cae12e651e9834fcabf23e2cecd8c146f36
z121664c266838da7ae9dd5c38f0182d722c17ec0011d47a91cd08f97a3628869d63c8938f7acea
zdc671a5feb15668df8a2b0731b90aa3991f04dd9232fa2377612d7d2f46c07bcf69974fe490c7f
z13c9e0f59df592b87581d2d726dc18360a10b6bd7c0866465aca08592445dd0f0228ee54344264
z9aee3e336e9c59fbc65212552178ec2e388eb11012f56580d53377fb5692f94bfe5dab08114338
z27c015d3b19f414c0789bdaa791252bf00bb52d98c5043c65bd0ea012af3174e0ba988234e6d32
zbdef1f7e24c42c1ecf838aa92d524fdbcbf05835839f083d7eda6658fc801358a136eed5865ceb
z3e771f8de2410bfff4737cc78fc94b09a8c0a733b1620acda17fbeac7115709cbad036b3e8a30e
ze3c17caa203736c3129f3330867f77232a36f847b4e804ffaa7c5a08a9a9a5abef8e04fff7c178
z0a49c08ba2dcca4cf499c0e3dd1bc8cb1f559367e689b85644d47d95f5fb6cdc38e086154f4796
z3d51fde9a5f360412d4617b20a7fa3bc6a540596fcefe2f3acdebe5591de40947c72a665574367
z3820db79d1637ac3117e4eb23d14587b77649f2543df0f70e531acb600ba316cb0ed4b582083a8
ze573a426bbee750985092a20c64ed97419f0dcfbf7efb41e8df5f27b1fda442939a525a9c9a891
zac35109a37d68e1834043f6b070a7c943035f12e06b90cbd84e87661f6470983f873c39f75301d
zd8242a353c66d2639d2f30484a5564282a5bc1efb50829858fe824b42d3a582d868c4b25cf52bd
z9204a76cd4e9a1fc67aafa6a7b01c43d6301d010c8e93a6d0ab3d1a0096bd396447cce16478d95
z182284d4bda73b3cb463b2f0107ecbcf55d4a6d956d1e8f55290465295713452fdd72b51e7f266
z78021f1cb7ab8aa9cfc12d1ba4060e9db746259d45b5f3bf06e0f2f2fca3c570c98c08c3c4dbd5
z7f6bc4b2b5b7f335ea7dffb5ef17db672e9980e2c1ea9cb7b6d1691d60e2bca08ca61a83663b89
z3d8b933af3a2be8502e13a313d9c10aa68e4399be03b931d145cac8cdb64c2f5dee3a9038c2aa2
z4a08c74c3d3d75298f805f4764308d630879c7f125ef5a7e0c1e893aa81279f352debc0bb0ec6c
zbb398cf89fb80c9c299b9f09b60015ce877d2d36ae74eba5bba5b06b1197f408a1a205b818f376
z03f4dcb5e55ab2221371ed66659a2d03ce1be30ba5d59447a6d93532cdf3df88d1398f2f9aff66
z7b26c2cd2ee57e87a9e370c0e2cc820970d0e685189316c1efcde513a98097ab431a9eff1fa852
zc964bfe6fae19c9ebe45b16ccb7984494c51c4efe781fc127515298814b0ed3834da876054534c
z3ea474029557e2aa713db04fc03852c4e7d9e6fca0e417e5b8ff1d06e7bc6c325cd277a9974267
z409fb4feb2636744144e2464b5dc383d42426b0b9db17ab52abebab758f31aacbad166f42f5d66
z7785e796587efc94f37831695581e2d43fc728678277f599bec22ee5ae96ee7b077b54cf464c8d
z05e36513a1688b94e4e7821e5633d0e7dcac20a4b9fdc5a0403a472555ef6675acfb7d14e9c9ef
z85d0690e13a9da748cd1c577a40666c4e9483e765516d213703f316ad718e5df831384c926a63c
z4e4c23bb28b6be703ca8621c9466b4626f26b5b7af3437b761cbfc432d265628c8692888e043c1
zf88b3b498f2b724fea9a4684e17c4983ca6b33f3a7627c33957a0ca03ab3e9cdeb6429a2d124ff
zc2f705ec003f9eb377cdba07c642a523dbefc3852421ca06e7e554f35299db0a6d331313f210ab
zb31706ab78c4bac8ba5d6be6469a93010d7d953c6a04c404d79e15013e9856c5e3b2b95371d63c
zf786ceeceb1e7164375efeb214d53ebcbd3dc72b9fa132a025664d7f7cd8cfc965a7b036176dcd
z41e023008ad7808c2c48fa94c1de9f999981143a234f1e93bf5311b980ae6f7d702aaf6967a913
z5996125e6b8d931fb739922914394ddaeb8ed3e66f6341f17530648b6fb9db713cced4fc1a5aba
zc27bc1ba89a6f4bc695962f8262bb86780476b221c06c534799e5d8f1329d0ff8a33073d19d547
z39b17fac5c9415a7ec60a8d68c02c33354db0c2f8b0e21caac44faa85a51c5e7dcda2416133a79
zde639418c32c7b5688772ea8b763bc57f2470193adddd1ce2dcd7f92b7e535007e873c1acc7c0f
z2aa82a4bd3fe2ee764b5fed29dd3de6a67cf2081f1c9380121f8eb3b324258cc74c5441df3d4fe
z0b12d008b6fd716f0e054e508eb85a025d3f72a7a9ef9767a82c636a382def4539de75487c2ae8
z7bfe21e23eebb6d9fe6a0c9af5f19a87c6d3b29bf35e31664bafe0d0ac001b8f78aabc8cb23013
z06407df7ee498325d01ebec545cdacf2b9ed4a75e2524b79aefac4c9d3c4af583c781abb83cd53
zc779c9494724b6cf67afb3197bbf53fa216118e60326677e717d2a58d214dae991e92fc42e0b25
z46936298c44486e1d8dc1d79b6a878e9ff774252c05e29cf152d3816b7b5b62644afe40e208608
zd31c7a7cb92c32eb305f35540cb7d45537fa6271b8cae5351ae6590520e0d1f5b93b03154903d6
ze2c35f0312887e33f2be03e514eb1cc1578dad53965cd0c475463ef5e0e01a2e41882703799ced
z9d58f21dfb783b5d10a3b5eb6c241b313b1254d64805e0eb0093e362e46bb980a2f9690e8ba704
z84da2506d04d42f47b4ced943a81bd0337ca166b3324116ec45e672c1e854c9ff9d8eef65df7d1
z7afca15d71f92a1eccd52adc5428aa8b053e59167399ed9fdb388472c9ba394f92c635571ad3db
z1a05e0e2025dbe5d0bb4a8edda53700b54c8e6f3346354f827e13ce229bf98f0ed218a463b59db
z5c40527d5b1f0cd4f91f7dea26ed290110326441cd2dfca3929da03170972a562cae1e95971907
z548f7756b78e7ba3bc3d0f30fbe64f8260df77578e6b0dd75795b3283fde8eaf67e3885ec0ab87
z89d845584dd2479d9c22c9ad820900824e9b66919ee3699a963efec54d973423d94a38e1fde4ee
z3e841fedc7ef97461ee89c50afd9bbf14ddb8befb7afeb2f6c02ec69cceb0e99b8792c14bb3b16
zcd3f4861d2e2e98c8d232b352a7dd28e392ceef669e5acf6cc1c758035f42d70c66c94bbef5a1e
z57a0b06edd59aefaa6af3afba6a45f670b1d2b00f807b25d9e9863027226062c5817a25b3bfd33
z7aef4c8de2ddaff020fd7227d49b39068f1b196f5f5815e1d34ad2cb337935bbe47fd93f1663a8
z5b7fa8ad4c0c0c0789e53e8cdfd52d1404b90abaf5b25ab0443f32e97cd80292e214240c708fd1
z977e00b5ffbc289258fe386eefb4f37b88789f298866691e0325d09a5ec10b350a82dd8c4f7e27
z79c007755256633081375f2ad5d1482c3a9ad90942471dbea9f7d1191bae25a50ade6f65aecacd
z6cf2d2f4df3fca4e947b74fc063819a9defbd9adfb7d5d7d1348f6b59dc067729066e7c9b1baa1
zc3b8a19102f9533edbaea94f882252db413b5667832f086b47f72391e2732a1e1e9af259a1322b
z9d937ba3a93adc7b19108870b3f222811ebf8a8cad3be5eddb73df4618c7d73698c452b67247d0
zb0d59ae8661270a0c022cfeef27492b2f98e9973b541f899cbacbb568b37479062c8d06e127f12
z6eb22c0b98af53f58ecd49a1db719a8460f02c8537b4f99b902d76a160df8d59bfbbbb47f734d8
zdcf406c794b072350deb1d6603c222f33d5a39cfe56879f29c9f1d5592f37da23701f85dea779f
z24e2ef4ae391cd15837ccc216e1db9f52bc7c6fda4e3a23f87f6f9a42b7dcc9c587961d46047e5
z2a73df2559baff9d8f6f2a04373de6b931fef1816748722c56ec5506f78d7ea1d54050ad347853
z00e1a33aba8e686b31a5c61626adcebb63b9d481c8e3a55c8a274b0b67c9f6b7d20f5d3bc13cf7
za7261190bdb64738dddf7b4784893b3450fa8b3e028c2480689db46220717063f4608525288585
zef2cde1e819b296aa87440b3f31cb64d044f897a18ec1c325f5a1aab4b9807cf86a1b8566e8f55
z4ee5b4fc9c51f7c72b44e500b863f45d1658b5a7f75cd5650f1cbfc605899fc0616362536c0748
z73942dfcb4f91ce339baf13ee5002d97f2779b95f4c9b711717eaaae1f0c9ab2a035ea3834a377
z2c69cd9ceba15584de969116c2c81493ad93a1d47fe0144c976725ac02154b8cdf6dfb0e283bca
zb7f4f8e1a91be6e22b6ddf48c5deb8fb9bd1be6ec665bd12c7033cf5a27bff4e9249ee2e1c5563
zee718d12d2fd17daa9de17457fe3d06c2bdddb920266264ab2adbd21473bb7752d54cdbcfa87bc
z7deb5bd0d1b508bd0e9e0b0c27de21bfa78bbf571a51193747b62569f4d53c4a093200a2d224ba
z7bf33faba92a6d1f22991069c71e392c5e8ef30ffaef8fb77873d30b86e1ee41876cddd0e1b97a
z799b031f24d5313416d79f6b220b35ddc49cc9b505a7bef902ab9d06bd39aa70c779e8533582c7
z7f7a348fb0a785b4025089c84dd028ca27bd40a57cd2b9306ce79c050a027c8afe8197b52cb0d2
z9cad6317ab36b3ad0b4d224d5cd9eb3ac434471868bceb4a1e04170d5e209e9f06e465ddc698aa
z0c73dde6991362693a906581d3fa350826039708d26eefd0d3d708dcb1d531752d193fe561d7ea
za4b6e496938977b262f08c3130edbeaa1bfe9054dfc435ca914e2dd4df87abb6975ae0fb4e6114
z09b6ac04afb903d02a6369224afff09508aaba3ea32819214d1e9878a8269f30d4163f264fba1e
zf1cf42613bc8be5cdc38065602a9734d74e364bd867bfcc8219247e0e03f1883ffefea70cf7f98
zaa20d645bd0c0b7abf21ebcca9a914c5440cb5c7f7ab53140aab6f57230fb6ed4992c9074710ba
z4703f2451a45ebbf8e60800545301805b5b9fc277b6646d9457b6b68b69354aefbda3eafc24458
z7d2e32985eca38f8b5bd092b5633998217b1383228339d23eeb60bc957aee8e8d5f6ddeb6888a6
z7b84f72c3f5560c6151943f22f0f7301830f0cecf0dfd8ca685408fc6ab538f73f6968cf5b36c3
z74b18aec035fb499a0138cc113ad6789a9c7b0989ba5c3485bbcfa02ea5ef5a50eabecb3035d13
zd116a1a36c752232f679e418c3defd6d7fe4d811468854ba1f467c419c92aebe3dcd3a38c579fd
z8ec6541c553de663759e57923d909c109f3421db5bd991f41a36ac8531bde9c8eafac1e4fe7538
z3d2c0ee143182c7f3fdb3b35bf169967b3f491924d4494dfd11cf1a23a1d5ad15b9f7cb2daf027
zf41ee1066f2b433cc134f8dc68afdbca35844728dda32b24b1c9d02268add48658bee3eb2cad80
z20f06c60c51d2dedad87a88676d9cfd0d403a7265c103d140fd0072c8e753428cda3548aa1a5ad
z5760f50b4f330dea07417d6966f549abfb5d6dce49e2081290da78589eda05d9b96c31a8b7905b
zdab7b6a951fdb59d09e87a4128e9ca07e2662f92fc5342ed224e06e1d267e1b2b1b0b7d5b68e19
zcd48c078f12404f33d5397b726010af430cb10006ffa26275c9a94277b5a1755461cc3ff777cff
zfbdc341562c0032c984a1a1a0838d58d174f1b1f696e6347d029028304b156d07d4a5d4bcec3d6
zd83dc9f2dc3d4ebe1bacd9be7e6ac146d48f1f4f29167d3c80349d88b75e147a51811fdc2ae8e9
ze8f65c77d21e71320819e94c450da5fbc66fdba7714aa849b6ef4edf3e2188d8d13dccda63e4eb
z0827b54310e5915a3e7cbc75a3a61f53752243d057c6e1b697ca0ea6faee6732102a2898c7a4e6
z2004031668d55936449adfe04e930dcb0b0e444f591fbfb5f89216f072b3f0231e61a4317fd730
z89b724022fccb4ea6784c99dc2e6f27999442344fd5cb0b2e2ad53c6ab68e2af1d6dc902fba2a9
z72de79b39da84de719009186afd299de01c3cc2caf90ab178d09937946cb1504c81603c0edbac3
z5c364e787e6934249ba5fc2a467e50bc54c7cc58c7c91c3f3e4ff4861cccb9adaa1e039d865ef7
zb7925e1ee3ef17ac2798ef957bcabb63e01443c5c14596687cd12b4a27caccad0e64b3467a7b2d
z54cf7ab983f723e629ec6a182230527b4fc8f1b27af90f1cfb888c1c9806d70e1402c6bcc13967
zf3cdba38a0f3423c992938dac92299ed39f4f3c62bcf9393fc9f175bf19ab8bbc864a759ab42c5
zd6bc5d07e73b37fba6c0cff7178e65ac06629feac309aed9cc49f86ef1b461774e0a55c3c6059e
zd462d04b173405fc744d7f65d4871cc623b753ed9b3bf6c6be6da168d6df59d562f8dd2cdf315a
zdf89a27d59d34044fb079001e1f09cb1a2a44d63741322b4ef6035a2e3a956cded79ac341ffa3b
z9a6bb34753ae9648d8e56546aec75d0c0415cba76d2d6069b2e86908be249952f8df73f4106ef5
zf0027dac44d7a0ad4b88783e34961e5ec2f323e0874469959d1ff060ae65e23470279de967692c
z5e4043bb88121960acf0f2f2ac0728c877f50278a15622d1aaf926bb30132b22c64edf544f1e7d
z630713c59a7354ab4ab93d756ec76ebd3b96b4e91edc2797eab0dc3e3e93730492ab4f3252f996
z5491f1fa6d6e1f67d33d62621bd538f26e3445da6b07a1c170344fd7210420bfdcb06aaff42af8
z2d65e9666464cb1da123e4d6bd41660bab6aae1335f22ed7a822f57a16ea8cf2c6c9f879dac677
z1e895e47028d324cce161cc75423d5cbc3fdefd11c66dcce832a596eb8492890fc9a4412077bc0
z108435494462c789dc688182195ef0aa7a362369e0f8324304f8fd9941cf0d6896265ca4942498
zf31a4be3abb019841913582fa730834ea0d5ed494ab795be0cf4703f9eeb27e41039c1ee448dc8
z312027799bccb82973010e8776ffc6b0078ea170990e9189af4c762915907886c4e4e189929980
z9b5e525441498a3819461d171d31dbf5ee3db4a267629490cbb26244b8fe6ed0ffd4907d0b6cc1
z2df9c12172f8c5fd3b2ebd7f6b594b35e863e8e1df469e932c2e8feb49b31bbb09fa31f08df0c6
zca4ad1aed69353f1bfe9c86bf92e761f4db04a8d84482292977f69151d56eb560316dec8b33006
zd7a34471de66f92c45b62bc1ce8dcd98e6c3cd7877f4279a82aa62c24351fdce7d179d62540715
z4b1ee54de0ca04c8ce91bb6cc1f56026522da5f4f156cf403750e7b222fdd4f2e9d2fbc5c1cfa6
z7799905d216c6830bd909b0eb981258a393144acdb6ebd5052851c302af00e429e76fcda28ec2b
z521ac86cbdeda19c8f2381c52fb1225787cfce7fc34b90713f5022613957f7f83ed2bbdfe800a8
z4a0e8f3fcb6ccb4221602bb16239788753ad99ee52e3bb09ad14fa1a8eec08542785b9b97ab76b
z4e85b2d2f917218340bbd2b0e46fe0159836475b447d4f1bf0e7302843b0616d3e3dd9d27b7e35
zd9ce50a4377ebeda3b68dea26faec07a9c4b4279e256ee56da41129a3cd15a6cf9425862a1ab58
zb28eb285bddc45f023be7bd6eb0f2d031a73e32078e195689c12e70f74a804a6e9c33e1e2868e9
z28508eecb832a5a3a01bd268892c52c468da9b45db7c58f604807903ebf1ebc001b8db9dc19746
z4f69d76f4a2ee81b73bbb4e3fc6bdc16b58c56e4caaac22ceef79a9b6845a0caa395b8148a6611
z49a7d6ce3cebc603d2de24af8d952be95a8a01f390d29fdf5763bb442d0472ba35a2f103de0efc
z921620843303e071f890f9a8cb62132cfa200fa76598892052592beb3b6c1b01c8c3d8af0dd94f
z9c863ba7cac5913577e30c06a0ff600faca61f73788e4dcc7aca16630833fd1cf1454afea7b30f
zfe699a6b0fa9f45d058dab8c4728c8227daef5a28a049f76715ccb84ffba14831df31dde3d4f11
z6ae668dfac29d976939ddb851136b381e6489c84d7530113005db441bedf5222b17a5429999a74
z68969d66a77793cc85e8d0fbcc76e3ddebc5cef2f5f488105b26958786175fff1afa658597179d
zde67a8f0507a1c5553d84578e531cab6bcb86be6a1e8eb07382969dd300bab4273156ff359315d
ze8533f6c6442d7f1043b43188776295ae057dd0f930306b5cd36739a1cd787d3f87aef60c68a52
za468d7ced143d09ffbbab2d33ffe9e5448d03ed11faa607eb895c9813d78786aec5d09f24247b2
z2f09c12c168d924c978eab918846b8102bbeaefed13172bd04f7e3476338178f8e5f04efcd16cf
zcbc330fe14e595f72bbddbf4b3370ea288c00ecbffaa4b7fb5e8e95681ce2af305cff912a6910b
z5e381d39b7c3c9b4b0a884948a733adae9b0d4978373c34c88c4b5be97fa2aaddbdc2148d801ec
zd167693a33704d0b8a1f190034c62b13d4b1dd13910ad8eeaba03463622053e1cfd9f442a4d96a
z419adb535d2574c560f2340ab8c2f1ba877b478da772fdbb3cc495fffb00dbf07d29e7d7405730
z7dec7dcf5e2d4188e62d1d0699cb72a8d395388a6d829aff87e8d4492880fdba16dd87309ce43d
zd172d8f6dd69407ec99e7c5442cd938a90c090db8d566c808e3ada53290f4ff9a0a0ff503cb3fb
zad7d964573355e9bc247ac91f40c78488b97809b1500382abfed356872732d54f6e6fef6a65ac8
ze093a854a95341e53e6e6182e5d69dcc33f0bc1b5467304add08fbf6b5b33f42790e78ef2c8ef3
zfa27058f41335bfb05c1ab2d1a32f72bb219f21b820f8c1dd1cc4a12303790d81a5b9e3ff69381
z3df99e6aabf27626eacfed465849ccea780bbf3247dff063904c446a47c6334753ae67826e7adc
z6b9c3eecd32417023e34a3ba227a00100ecc849ba5a41760de5239fef40cc4fd01f1696a5e3420
z41494553bc11e70de05f02f361e834350d997f1719fdd1e4b970e9beaaa37fe02f4b8ed985b9bf
zdf5b4f8e5c5df3f3d156fb428b532bffc8af03df1f23d1dab0448254945567c0374ed48cd2f47c
z90c8fb6221129d9fb61aa1a188db2087539e71056970d138d8e9b9a825188aad413a2685b53d14
z6ff0999c4c20efdb0f6f56ac592547d36afa4482904b0cdbdab1b3576cc8794986bce9757f7dac
zace0872e5f734e94bcb55232f8921719425ef33ac120822ebf31ab46429e0c676dba8032ebd515
z38b738866e5bee1347944ef232a3755c1df5c48de1fa36a5d96a11b1cd4100110e6b88cbc93344
zf3893102d283896fa5d8390028798d355d19d2ff4b4db0bcf3fb5915a586c21b191cf7d138f7af
zc1f3c146b55598a46b5631cac589550076bc5364e1560cf65d0c631f19bbc2d0c220105d149875
z91fc6965e65d1deb64a0b9a32f81fa4b27f86dc691356376d45b1dd475a884047b4085daa3d24a
za58b7a3909f6718457d971e730b4ef62b7f6fc8fdf2d901f1efb4f3dbbf6bf12d8289c3d3a5600
zd9b1b63fe7057384ebe44022272950ad760f5d4b3db0f0850ec796cf573a67125452860ab58d32
z5e4501a01aab253fe3ccfdc75cf0d1beffe1dc4ba8684596f3b8bb5e827b5f40afc16e7045f56c
zc8e60bdce099e50f45e39982d01caccc57098aaa11d744574c61ef92130a03575dfc23de7cd18d
z5f84e432159a0671b6f32539fe6b8a5e57d09cc941f51d2b01865f7a85bbdf25007283785296b5
za6f82e2f51959a5a479f62816dea5aa555f9263e8172aadec4a9b2c154bb9423ec10b543bc4a32
z41c09599a96949405c8074863d4cd609b5471e856de56eaa72b132ddff9390253fca10bdf2c675
z057509031579444466d2a2a1c3a8cd826dcac6992c154bc7aad31616d44adaf73a93078cf3376e
zb69b22ce823c144fab204a3edf90e159140eb056b4612c335995f55764802c4482446874daf518
zc517935bc59ef9856860bce4800432409fc4f78924e14f6d8a2788dd5729e5b69a30dfe369165c
z5da23ca74158227edbb246d65d2944e7748e956a3cb6521743fd6e8ebe38c75e663a91c6de0ca4
z95d4e71d6eed60ee6763ad65f644f2dbc909c9cf0d9c2d98c8d072d544225d3059db43541f9ef1
z0f31723fd34936f22d1426b20e2e232683b0ce87def9bcfcdab062aa24c812007c23c1c903d934
z848777d93ff3f0e1917fe95217d3bd8b8709232ff66688178a3929d0163c99e95577df5ad616f3
z27e9df3143393c361a1fe642b2e481d91d1daad0e54315cdd0f3b6bf0c45c8b5a7f5242172885b
z04ff9eba9b7afc02d14ac16b2bf08ec1de16220f1d16b43cd0cbe9b35b707fc8c5303e7af31f90
zb9254aa71f59bb623190c837a896f491e7f93ea41f1ea7af253facdf61c90e546db75fa6a14455
z2de2c0ae1bce367c8695c9cb6ed419f64c54cef07abaea2c5cf1453377a0dac249e485d9b55931
zf3bb64b8f125369496bb91fc70399a932aa7b446221fd87e538fd06afca5961d90850581a606dd
zfc63f8bf64f65140103d0c773cbdde3dfc88886db02d3eb6adb1c8045fb9df308887dc3e418da8
z271f612f87b4895d60846cef2f2a5e3c7d215b1a3c2f77e7f7384d3be59e6902d133ab9dbe660f
z333741dabc0c8c5143b1657c9a026d7fbcec05daf496b7002b138b5108663eafd9681b11db29fe
z698a987a05e56bec6b373518de8cb3cdb89e826cab09a8df73fce9dafe46f714a9d94b4cb2d4f7
zbf9e0b4b4d9403cee3ba29ffc6cc6cedd29db71e35c1c1d2dd813cfdc1222673be5714404d00aa
zc623c991d7e6b69ff6a7e8ca051fe56bf8aaa301dd0ead6b22bf593a8a529ef3f260dfc4c8f7bc
z01cb071911bb74a80829cf2cbb481288f2c235ec3ea2fbca6c90d775839ed8cb4b2d574512b7a4
z92f63763cce5028509736fe27a65bc08630b0aa07aa4f0d01d66afbe40489dae0425c45133197b
z30f2a49be0acc62229238dcc5fbd31abc4a9f90261c8fd7be3ef9b9b46dc57a7b0bcc21be15a08
z35ae33221003d54838badb31929370fb7c16a49cea23d3b57ed223c69293202bb2fa7cb7c28ab7
z019b1d6e0ad1c4de6767f2eaf96dc2a3bd643edad8b34ba5c782c11fa086318b2e29ea2fc8d8b5
zfcb9d893e49eb0417663a480004883b67fbbed801a6c5f0abfb2a3fff3b38d4a5a0079bcea6274
z4aec0cdbaffda43e5b3be140282c672ab8531ff9331d6047cf9a36e0ac2e19ab56a693ef167dee
z812a7a695f57f1a599a0a835014c93a2849d36b5c3eec7f7cbf5f2ab04d0edbf78032064426116
zcadc76acb115c480e32aa984116dfdfb444767ccfec0da4f4331b13f672c1351dccc79fcfc35d8
z3f0f8b97c6e46e7766fd35aa74bc2c003cf792daa7d83d1ec42a0a3cb4e68054c4e11030a6a77e
z6031d0a67c64df6709677b0aef6c8d1afd03b70dab15dfa21088f4a5f192eab4ad65882f2bc8cb
z9aa8bd22ff264ac308903b884be87ab5c9e272081c5588e7a20e1564ec73ef1321c6d1cdc13f9e
zbfbcdb252cd6bef03611e8f866e1e1e17309c06f2341a0e0ee4dcf88188be8fbc084b12dfcdf5a
z78139b65f5cb6e0afd7d5e23ad28a66b08ba59a6ae2887b8b489ecda9ae47d96b7d536324be01d
ze0841cb91097bbff972268cf2e52c24189bb36c93ec457cbc6500b0421c0a09c6af28f33483c9f
zfa357173a85e628f1ac62d1398460dc02b864374e05d4739cb29a3e842a5cb66a02a1abf5ea3a7
zd7897f560b07e79a736739c6d4b5c56340e7bc6f7c8af8b5d816e1a95583fcbc83d547f0a40b8d
z2e7a615708ca210d9157819a391a44e51b55d96bc6ecf5f1f4a8ec9385be7f64e934a97181256e
zf59185b99e3dd3622e5e4bfa21b6d2dd8cbb81db7e8b133c9f27828b53df30e84eea3dad9f1631
z07390748ebb4c7528d929fb8d8c5535c7753ba4961a0709431b3a3fe35429141d5a8b3afbf1c27
z794227fdae42d1a7d4aefbab4e8834790a2308ea12be3bf7a3dbe617e45b3195f34e889c1d9d9e
zc6da5bcc430d5e6bb3314fcc65fcc51e1f010f808a9b6182ac685628f3e50eccb1c536581195ca
zfca0a09df1f8522bcf6ddcaaf410aaa7e7daaab135fa34055308723e7d37204070ad98491be370
z273c1ef3bb7c91ce989f7a2933a869fff8ead21fd5225075c9126adb1d3faedeadd2766f0cc7ef
zb77702daafc6eec2a92e647174790983b90d98c2739440de64204240df57d49d1ef07765349a98
z1bbf5d3b5d47da1b88cd18fd00762809fcf21575da227e5e45ac6000225d09563a6f8f84e85345
ze5512d2a8bb96c239ed7a7d1251fe0ec955027a913f5d47aa082a71b088710529f7670e5ec83bd
z14955e21f4258c8f29eecef712e5c304ce2c8c6f4b2edeb0b3175e80257a40d103df818b83f3a3
z078f90d52587cdf2a539555623ed374617e6f69b8c5635afcfb4a8d91859387325c1791d10fba2
z2bce2b98c607eb4a47a24c815bfa6b891f767e69fae27010d2017d15e0a0e42a11aef3d2eda47b
zb67e62ac4978c6431944c15037ed72420a41abf664af5c342324a54244e9f5e6dbe801e09ba20c
z9dc7d948809bc688257e87e3d819e721f6b7a1603c6f8f438173ff45d239e6919898210aeeda21
zf4b825756dfdcbd1ca83ce4f3d8d9c51793eabbc506389b91f4eac386c3c77e5c0099ff703e8cc
z2e87baafa78002f01ff395517b396320d3dca517ff6e5805a26d076b5024c33eae812f86e18a2e
zbf1ec4f1698d56c24a2e892e33ca83ed4b761553a4152fde2fbc0395a54a7997fbd2007859051c
z91bb57e1ca4c0f664f895a2b863c47c54ec3e7187a35de163712b23328c2b5f0a4b22d4eb597f8
z6b7a646be9e0a1d649c1a0b4a456d929c0f32282d77fefc68a1aee52f0a78c31649d9fb2dbed10
za9be21e6f3ee535b4841461a8d361bc64bf740c8b1c4bab2240ee11919244acba39b7ad8d3c578
z836f448a64e6b5b89faac5b7d673e8527c49907b243d23a7b0e5d1ea4cfbc59ead1714ef79cb26
zed39b8c1c4c935d69a2ad09bc42795b34717124f22c74239b1398ff33e6b81dc4e83ef81ed9304
z6dcbbae8a052a0e1dea2a665f0773e07d2fb90f8c6526fca42cbeb5250d51f06f4737953d293b3
z8b959f37666df15151b243064b19c191571d92152df30fd0bffa5ab20543e7211d06a12b1c695e
z46893890760b223e364c1e48ee4eb224c39b3c01758d0eb94752460707d06820401504e9954f2f
z31e791c958e2d758ff8098fedd2ca7850c79feb2ca93dce3862a7513f52a40f0597f14600ffff5
zcd4f2085d5f8d1ed9ce85ef9b4e83ae0eb039ae2543a629a990dfe871b4ff9cc0a7512dc6c9a75
z68010f71407e5a4ce7fc80539339a354f17df3e24f7a3c7be869064844e191ef5148ffe41c11d9
zeb0203f194d7edc112eb495b9619db3b583d0cc70803cca8072b28a5a21ba6fdc16eb65b54b35f
z3b50c839ab3cf083a38b0b0509e77cf7593e74ed0fc2f728fe531628b359883c73a4cbf432bf53
zdf80415910496006efda5b24266db6516016f7d1d9e6c6dda0a41eea4288c684aeb3143b7c2a80
z5c6016ea702f882fbdce2b2510eaf1719c451caef4f9ee1e22c72ccb6259ff6ecc4b77171254ee
z58f15437d2dcda92ce694692b0f5dcafbf48db7ae8e404847933f2111e87b602d1fae0be6cc701
z576681b793dad266a9c34c2517d6fe1b53d45ba3876cf4dee6e342031afdecf2fc1fc7db2903f3
zade6c450f4a4624eca8c7f818e7ab1168b2d92f890a5b21f2a8c3b4abe18869420130c6b62138f
zc0f753195e09ecdf6446b3990c58e0c12179907f20d41d13d4dd8be02c27b12f8bb08b8f57f0b5
z3691b1db772c4c541f335a1d207f98c0af88344a9202372ddc3114af6e009a1e072410f7521280
zb343bb5fda5c3cdfd7ab9dcee602d5284ecfaea54207c6f53c0fe335d1e60bdfc6463b09288a8d
z018bf63326079dc57dbc8119d10b84e3c0ae86fcf8a93cb75cc58c32b94003567c33d0f2f1d9de
z75a63cddc038f4245665217ba7adb1e0817c76ee4ec699093586b9106eb8a7de0030048c4998f3
z039ed94d69723c05312908e7f10cbfc1728403153180b36b356496549734f41af1a362ce327a98
z0a306905b8187df8ea679fcc48764ce16f965505b9a351ea302d56f1c28e25673285be9fcc713c
z946c63b24aeb6cbc270ee30e4be29329858eb26a0377e15c186dbf60857e364ec18caa4e75b130
z5fd966a019a87137189975db708f2f84f5150b353be3160754fa39db5586e36960fbd6b9f96356
z86aecb6f3bb3678dcc5554be6d2d81ffd57a3b0e633c10d8f0b17ce72a2d85a653d6920d99abdf
ze7c4ea68072a2d7a0802d502eb7b486c2ce9791b46ecfa9476542aafcb335eebb638da7999d043
za6f29b41bc0d3acba040dfbb8524da2569061e62143215b547db8acac09ae92db374cb5eb52e4b
zfaf6f9d15e8ab7dd2a785a501edb9f36a7a19e53cf560b5796586e10cc0ce16c158efa8a2d002a
z69ba12d4d3b171ba358b1a81a9e87d06b3fcdaac03d8b08ac86c0be8638063a3ff15f26b6aa14a
zb4f07f45216b567c80ecd33891a4a280f778dcff8c5a308908f170f99b7b21c0b3e555ffee4c2f
z66c0c67879b7cc6d2f222cb6ebbaa993cfa803960af2dc4e95f01c93e892541b361c9ccd0a41d7
z03b2eb534788a9a64b1c9888d68f8ffe219ae0346e4adb43481ad2ae1d023cf5ce908e25415415
z732f6cc861d82bab44309fcd7f87fd12f6f7edfd0da412d6412f312a7fc11ee5889065724cb393
zda5c82bd64f6267717709521e843bb6cd6794587180dcdeeb42fede7e72549db80f384345c8194
z654a7adb5de1ee50151384d1bf324b28329c8384c7884c89a8100e7a67e14fca3caaca4833ed42
z046f36e07eeb9e8df6e496ae23c143421e7f2c5df25c42f5ae672725a2a03c150f6c41d3b63585
z20748847c14e02ee26a026380af2b0e04fc1561994922ff79c6ea3b569f1c147ad8b7c16fbcdb5
zaecebe57199287533ebb55446a23fbdc72d94a91f32e725ffc1591aef2b2bf37510593309b0990
za90ea5dfc2ea840ad20013d4c6fe04a30bd3e5453f165972fa8ad4fcf93df90744a0872f1e57a1
z28abb7891f3b3bd945e7d133a0439e6d6216f92fb2fbfe7200068163ed41e948b5b26ccb55edf0
z12e8cef2b4b65f4686f210a55b0211e999d7a4211f74fcc74c38465187733b6d8961924657b9a9
z7d0cddee1c4c3993a862fd913d03b708389a50ed031756cb4aa94d8d7a4cd38c100f69bcea3d6c
z68bfa4e940110b500c5696a22f3b9751e965d5afc47e42fe542a8c84ac7b095d69b2244f4e5e62
zb055fb81b01b1aadc0c419a0710d0106623e4432b5e87277ca833df9408958ba88304805966a54
z32483a2970c73fa4731e466857f4653254b1c9e06fa4694007aae29fc6d3d6f96e42a6b69475a0
z826be85a168b06e5884acd97f3fb771a04392a5772ab19668344a7b8a14b3050b9bae19d44626b
z96dbea3cef249ef5b689173cb1090f465b87e17a5c3d52e172345ec46c1a8de6ef7cdc160afb00
zfddf72dcbd5d8e44ba2a8584bd31960568007342d4f697a2571a7f42cff32f5fcf888363574b56
z55fb80758bbeb76b8e08b4bfa878c0a07c6ee0b13d82149e6aa7bd6bf91f1be4bb5c614f33fe80
z5aa5aec19bf9d817cd3df32e1f471502842414a1424a23350860727925dff9d4e94d7d0c7c8074
z4bbfca3da3f7892a59c91f0dde1278113f4047cb2d5f894b18493e574c56cd90f4513fe8ba6a97
zb1da5671b31df30031954151767c8a862615773923236cca6788e53960fc32a831dc811c344f45
z2b2e3e3cca8dccd51702adbb0f4ef09eb5f25b371ea5ec761a4dd0affc59bede0eaa53801be817
z5a6ca785ad563d8e593f0f2ebf8beb07b241218236f1d55d5c83d5c291d4cc040359227c079e8c
zd4cde834dedff69721ed7f67846384e903bcd45f1f1a8c706dcd4ba3ec67cdc43dfa800a783f39
zd09e871b7c9412c5389793694e206faaa20406ef74c05b14be6dcb95a7b82f2c531289161d7e1c
za1d9c074d6bc63546e43faf13057ef841a5395aa3a24605cb5c91a981e5aa8de090900736af017
z7b72e567bc4133f5f12e7c4550ffc32eab654ced0d78b3e8fcb845b50f240a6a84e85c028727c7
zfede5ce598ab3cf0a247013236ccbc80a15c9c70c237d01d3c837372e6dc415bac7b893a25615e
zfb2a83b8e87f1f960ef69b7bcbd64f01cd2cde260c16b9afa9a8e3d01d5e49408fd6381427ce8b
z25ec76b1ef0aeb778725394fa27518767bd73293aaaf599ae14892fd204077da2f3db91581dc35
z5ae9061042a59ad8927b6e0e244ea6fe566508078f8f2155c2667bddcf4881c7837dd5ce07a00f
zfbfeed3ecfc3ae1634270041a603c226bbec2a25a6e4062fd00bfbe5375c1f15c7178fb495e604
zd158fad97e959615c7ed4e42c660972d62959d1c06ce16c796bc14cac73a2ff04cbf7e50405837
zff391486f84b615ba3831763bd0c290bc7078591aa56f9bc2c53f7b608f9eb12cbb7925bf6d67b
z737ad91f9867f95731512d7d816d15c94746df60b9a3d126112f80164e8728f5f1a8955c22aaa5
z4a8bdb399aed621ec080f53ee3e7ce63880738768b86f0cd43930e5b42467b330e697d2cea131c
z2e3d025d093f90ab40a5f70c72dd4827af7f1d005538e254dab0c6acad1d78f4929a62cf764bff
z512b1852a51bf839715d65b6c9026b691ef4f373f9bf5a2f55a8e97886aab42ec5d9ee511c47c5
zc235a2f7c3c080caf4cc83e825a8cd687ab7fc7b413aabbd905b985849392c1b21647e21fdc087
zeeda95ab9d49658aa362b3d1f2efcfadbfc94f093f0405efd74a6453c8c8892d691765523d03b4
zda0f20dc4d10c38e90e0235ce7aebbc1234baedea3ac1cd0c5539995ae9a627e790af5fbbc1a09
z3967d8710f64cabde32e613aed6e1b528c376e00df95eadf125a71d716d2ec4e8f5170a141ef97
z2fc1b9c709c7a7046d824b52a6996f45a2f6a7b43465514aa2ce31541446ec5b12f8f4bfd045cf
zcad969479f2ea23e1d06b9fc7bffe95fc51ab13fc446e5bc985de0d172102a2d5ef6a127cb1f95
z08bc64626a797c0c1205fff55d012dee6100d97b492d884d62f8c7e04dc0bef7a64b99763c6941
zf4cb9e3cedba52e999782479b6fc3b2f95580b9c72f2fff054cb0f50cb347584eeb4457c3b63af
zdfceeb071af8f44426692569f7678150af565c39c69a4ad2fc91fd5848d886366a8174d10c3b42
z2ce67bf04e954f7e4f1c67d6d6ff8c4e8ea5969e892be3d324da61d478f72b248c4c9753d6c9ee
z7fbf74aeb1ce8327d9f4cc23800be20790a46b2c8898fa3dddc9e2439f95b214615051a7f8ee46
z50f4453f3668be77a96a1185b8736d1e870ce82f58e02555950e157382c0a4724f9ce57d710ea3
zb2108f1624704cc731d9c80a8402d40923ce8845363608e43644aef4ea2de4fd0f4128478de614
z0409e4339ee8f9b1778d5e2c9a3cddb515290c6afa51d5addf93d0691036c456c65f1ac11d3bf9
z7248a21782e35ed769856381b790fc03aa8c28a02edf11aafc6a5a34249171d3ec541fb0837bba
z230f5a2aa3ddc59a71f342949586fec913806b972d815ebf16c2abf0c1ee321c5d146b4e5dae70
z242153a084c0434a1a86075d5b68f61df7d6034344634e2d098a7b0693e248b1b8900c6772e947
z4f2d94d9ff48f252dda710eff12d5316ab67cbe9c85f7a8580c920057a10cce5661651b1fff04a
z404838df19cb9929c15706ecef6c4efed5214b3ab48d020445edb38cc86ef3ef6b614594200286
ze36ce4a032463ebb5b7783f81bb3edd038d68f412ac9519304b9baa019f048c8af7b2148208a6e
ze9bdd1a85c63d5529d219806bb74f441e2bde98b11a63358b08a363ff65c3376e1861762062469
z60bd10e164ee33d424eb8e91d78237fdcb681debfb91c1d3fc47e01ad1a2ce358c3cf639a400ad
z8a92c1db032cb92681a388c14eb00f4dbe055c027111b52f7ef4dcab2926ea736bcd662196fe66
z2af800ff0374e85ee36276c4f48f22b9c294dc58949486ffa68369fbbda72e6fbb2df023232a0a
za33cf1a167e608be4b4be299c2457df3691a61105bcbcbe44277c426411cc2609600b6e618120b
zfdc6a5f26b051ccc43a2fa3e0c9c80d63b1d2b03f93860a5ace536207b7a3b99406d05d0de549b
z648bd033b407dccfebf39b593167cbcfa41eebb30f65682b572a6354c5ab4772271acd4c4910bb
z39fc82117ed837910f7b8fe6e8d9f175ac7d503bbd8065189730c6402959b4804271531b991adb
z2aa97273a576b5894378032c2082270a10645c45086dda3167f2d4e91bdf01b02cbcdea4e5e8ee
zc59679ab943a41dc6a4e8bc457cafd1becbfb98e4b79ab1fced3c2be8e81c939df6deadae09e8e
z5febc71799ebe02396df1fae1357c3adbb50b211c3a089e89afca1fae06d02eb66aa8535fd8862
z79f7c584d1e8628636f8774c4b82d8e162e99df8a39b55bbfd3f6c8d5229ca238dbee55b451923
zfbd2be41ffbc9c3c4693287204acb119312b691c2b2fcd4e329db5d21446273918d627a1b641a1
z3e2c985e363fb93452dd49cb2b9c128cb6c756b61c7ad5ebd092943c712bea2a2d15df871e8217
z199fe008abbeec09684ee57db04baefa9a505e7347ac144f00d19ffb06499fc964672d743f93ba
z8aa44c6131635b940a1e343d66ea344019e5893b61a9b162ec6b2472f3308029c0e09cd41c70a5
z80881555ebe1a6b121918312b7df449578d9936ec3d5255a386b677b60379cdd06a16c4f72d1ff
z27710957117dd3882fd5c811445624a4beecbff58b3d25bd57957639abf71d756b3da59c0bf19c
z6b29abfea03be87bc357a32c3c66ffd54937b5184ef1afb1de362fb36251c1d13c1db10e1ee3a3
z1751b0a3e53bafdaa5f172e6ac67f6dd1bc88e29755fa47c235e28cacce2dab6c44bc68d78aacb
z5d1f8dca0c5711c2f68ab5d36876c2335d5707f2a23536bb871a85006340b1aeb6b39cda0387b6
z0fe0c80deeada0055d844a33489badd0759b5a88f2be84bdb716d3a7da82d0b5c172de86360d69
z1e59cbd74ea2425cb7db1b46a217cea43e41809dbf63c9e509f521846b04f83ee0a1c7114de062
z14b96a4168e1a03a2c0486b5e410caa33b435916a2f74c370b6734c5350bc4dd71cb3e4692b12e
za8b62fad87d9336ae9bd015a80ffcd248403c648433ab0e94122fb791bb008421269384126ddbc
zbf709641b7dbf781c97834cc27712b12069b8cfeac33a70a10ef8e1f0958fac3e01e9ce2d377e2
z6c425a12af9344bd4ac56ba7737b8b52707fdedbdb0123609a44fbd3eaa6be2e0fca3c738fe075
zd95b8cbe52865e7a4c0ed6befac3684827ff9cae63adc9bd245d9157d30357dc6a8f4d3d1cbe42
z4fbf2471ea39e45148fb4844c3aeb64952cd2ff5dc11f03de10da7ca82651a82419171eb4ae7b7
ze8af54987de2e398053bfa08d0ed0725ff8cda7e4b54a2169b8a202421c0455f144916a01bd7b7
z3433f85f2012a66e020f879bc06599fffcf5b577fc1ba5fbbf2b4f38b567a53147ea0aef80e0ef
z5eb5f8b02e7ec3d98e5266910045f84eb643068734168bc2b4d46e2cd22b109cf15946823a8496
zcaad96dc44f8183d54b3476e103af30a94cd5bd66f5b6c86e0fe330b37a207b550124c6d9b2de1
z32644df7c1f2c59a3e19893ae433b14f8f3dadcffdc0980ac6774f48b28a8477a1d06c4fee97d6
z44b1684ff67f7069046bd3e7d1f3737ef7c328456817c66959b03c3c06bc5bf118ffe8d7144b49
z3a0711c9f5a3de408962b6d51646c881d652d26a608a507728aa973d8091afc4644f10d7f1e2ba
z29308ba634802f63f8bfa48feb247b58d350da1f48e04dcefea1cf395a46bb8129008f1ae2aff0
z44f5121759200c06492cfbd0dcafdc910e2a7774afd8d37fa25e250e58fb4c8c65e706e4226a98
z630d78ea57328e515e794b5f1302859b92758042698c1bfbd9a7ac699df2a0f75f2c158a91911c
za4e0dd9331dec0b64e9d93d2a895ac44302deaa3c01e9a19d0aa7ab18a8d00c4cef312222cb3cc
zd326f7ddd0d5bee81f1378c2bc3b718b4aa61dd99c59b6d7d9b75f851b6a470df2e15f30ad1cba
z9b24df783c1cf02c54301469d79f3b854fcf27b91f2e957bdaf731c34db62f7b327b3352161a4c
za4913667904b69ed798c1c7a3b4c7efd7adad6e1141499742680a2613f0c0ffe3213cb0e66fc56
z2151fe9b24ab57c441175b0d140ca937cd0efb4a797ce638f88201cafcbc82493e77221cf85e46
z37465026a4eabc3ad0adfc300934b6f3ba43cd072c53bdbc03e07ca91f700e52e94924ae1fc77a
z7e6e3c1d9e0ff916018672468ac207920b62d2ee0c189b7092e6cb9ef9134371b6d535e8eca317
z256987e96e17bbefdebb5599f164dc3bda85c7227abec7f3d08905c243e4a90f46bdaec9322efc
zd9b8902345c3a535b2359e51e485413231b770ccb191ec309ab048f2742447c0cc52489e996f68
z2d4bec99654235b0e5cb54642d1c59c7be7904512675fee1f7dc62458f7bc765d8e66b491494c5
zf9b3119ada9253e6f0d9c5efeea261de6c206e427603838a7edbb3f588f650fcbff085f3ced568
zb25182d12cc4c113a1475d13127275ff1146b490d6a1cb8edeb1e4d31f08c11195cc6cce8616d0
zd787f06f5c8b9fe3d37557332b375a0ce1c6a377e22e845ddefc434e598daa1d37ae2cfbe5e304
z7f08a73207ff329207f496988825dfdd6cf105db9aaa34def932727ca37be8fbcf04c166db844f
zeddf321d83653a87b66977a4d43b3aee38543bf75537fea08c3f4f13828b4ae004fc66ed996fe1
zce15f659e9c22c6025e7db922d5c75e12f6923ac13f3272489535b8672940bdc73ac93e23825f1
zb7cdddb1f4bacbe21d45e4ecc3755515dfafd2c59de86cb2c091bb18da766330d8519ccc6beaed
z01c755e837c2e826f6f62b030aba750aa926ce0dc9b5567e1db9156c895beddff61633bd8e7dcc
zadaf2b2756d42470ecd7fd85cfcf1e5bf5fdfdbda8a5d7265999478af45ba183ecf4d5fc60beed
z23ef420efa3ff4fe16b70b548f896450915f7017905f86c75e6bc3f5887b724e64c88c024c6384
zcdceb989fdcc8f414709406cb6ea9c71869f62aee34c046bdf9959dd55611d19eabe7a6bfc6e0f
ze418a04f34756e6835e16d3d75e02674cf23a13577b3da9bdf6ae691bbdabd49c53af99f54b307
z2718b1ba5c012c876065632ac5fe70d57af212b9085d1b75123eedf87ed0f0d9beb7c59af76193
zca775482ca90a564e6e76176dd1a23c2b33d6bda1fb4e901c012e50509bffc57f843351c82c639
z59b0a00563f20ec8c0a4f1137ee773aaa4f571ba0940a95ae27aaf6750a9bf49b56ed8779e3699
z66b69c48a6409e61e3c853ca4254b514c07c510996c5edb0c980d0f983c2a28a4defeeba2c45e4
z4a83495b38790e9d1e8aec65bbc0e461e48988674d6b07cc58da7c4a42ab27fb0ae1bc948f8eb9
za78ad08259139f695abb8814e03598e30230f25e1644fef8366cfe30de934bbcb0fb91436e2629
zd8af810666597ac2b069a7c95baaca3b6a81e525771a053db9cfa5c0673d6bf47acf3a754e8365
z0c87dfe6321d759de2adadbae9e02eed953b974b51e2568c96645673c5df07bae1d98aa0f8176d
z837662b5a58ac8720fe37dea1ec2bdf2ee4a8f86806cd88314857e4555f84e88a1ed0635de3d6f
zfb773436cbadab67fddc3d23176aaf77664e965b35c73e99bddd9dd8d25566c4e9846d4eaf1bad
z3ead8cda2b0aacd6525a107fd3c3ebf7c7d99e77367504b516983b8ccc41f4b050e8ae9b09293d
za6fd67a10891aefa1f20af9ca1fcec0fac0fc3e2eb88aae05ed00c0813c6223b811a81a9b7f49b
z9b9a994acbe190fa2ffa66cf7c95e75766f9e26eb3ce656e712c99191f5d9167bf7b27d133abd3
z4cc36973af742b00ae993685386bdb281080467a2d2419baea0f29d16a09d4c190b24c408b8267
za06da8ef38b12d576cd1d398075d51a734e78abf7a3e76f02b9a30ee76d4c49257f967c1c54ef3
z13144071941e2d02595f577da53094680d305e748a2c8802d8172d8d09f083e01ec8e433053276
z5722495d8e7204801d17ed0f73e582a37ce7756dd4e8d31687f9c0aee753362c186037b648aedb
zfb06d5f98d9cc2919ab129638effcb9d7d57da9ab74e28def898d46337f68d1accadea8ad15755
z0a6e9a8c93dcf1bbd61a9ef67336c9580247edc36234d8db235133abf1823ac1dedb3cad14d761
z826b77e60a44ce3087c5699ccd1e01812ca78ba0ec8f24e90b055f1f6d7159444ecae12693c500
z641f7fcf16dccf75fc7d09e1d1b95d898fca21766195202c5c72612ed91b9636ac6f65f7674a5d
zd6d171fc96ef45462b1d272f862fc4f4e795dce8ec471a929dfa43186e648dbfbff37ac5a54ffb
ze15054a53d0d432d38aca2560412326eb207645ba28655ef57749334231d4fbaab1b986431d5f6
z574700e58b1996b64dfed99cd8cf8dbca39ced2c60fb39b905bebb22aca08a872d4d01828484c4
z955b2fdb74929b0f44017b44ea91fbba062a5a5e58de37d8045cf6fd29f8ad140dfd6479d19c3a
z2cea71e1bf5308e83054e3af153a9d3a4a084b15e11e639236dba056fb81f26900974556109676
zc302fe7bf456eee2e00c02bc3ec483b574b5c4bd350a0c2c949ff661bd86ba0aa8d8db1cf037b0
za61a4d826b2026f7d7bc38cefbee98fbf12ad5ff833f355be9836b83edb0ea672af52903f310d1
ze4963f57a2783dd151dfc700efcc94dfa4e315a75d922afe871841a53dfff39bf69686692b8bcf
za3935bb6b4bff38c2ef443c12b130c502e3b16a2655218f56202a71a1e1910147cd19a6e24a48e
z4292da573e1987f6cd9deebd167b98919b8a8a555e7337c7ac63eeb5dbfe23f50c6ffe0499a9ca
zd574613439149fffe21f6a60f4b534ba42cc34b976379666dd72a77fabff0994ed54166d3a54d0
z3640470361f97a45764727351832721ac4d7a071cf50005425163e70df2cf370b72e3a5162f3b9
z3c3cceda0e99110416b68b9c8164bbe4460289fea878bd6a046d872e6315eed9f9bd24a74a1160
zc14990eddb38cfad869a158ebf7d832aaf89e2d43490f84be26bcee087e718f2f3d3ca7eb5597b
z21347bb3caaf3050ba3ece2006929e8ee61171b127c08740270115bab6ddd60b0338ca633e4ef1
z7976ae2afc4b74e7b621538f23bda3da9d88a6752d3bc7098f0392ab6b26bf3ffa131ed4187239
z8217f459a92a46652812ddffd7594025acb0bfc386b480dbd7a72aa2cb9b74857d5a3306875429
z2b0aeb3f37387e6f45d52f5572f56aaab9af00f47a7d51a0abb738bdce7de8e8b56a5099f97227
z26759ae8053f14f0034a48b093e2b37e235b8d7cda12e1d0679cfba79fbf65dc867dfb84f58d42
z690156026f6eeace08920efc3259e3833e6ef3ad732ebfaf659dfa76123af465f52dcad3833db9
z38cad63e12d43913988ffff9e4a282ba3c79e3f44d2428a8f88d300aaa8b9d7ef902931f031a9f
zdb5765d3af17a9c22833c4c3dee80017c84011a80b657daddc2fa656cdc94e179b15c1ab03db73
zf9005be9c64040f6598895bf15a3b243f9989f872cfa0af25b958c799b2c44e24e49035a2e2e38
z235c7a2d658d42982b36f3a45accc73d5458104b90b9d0bd6ad9ad3756058abe6802fc7c67335a
zaa9f5d2fe353d37a1127739843710f67cf42f362059a0b029497631443de71b8b88a0ac5c61dc8
zc7a8e122d478ff49d93c447abf6ec6cf19b5ce55e581c3008ef1ec0e5ff3d5c67ecea541545f8d
z7094e9292e8e5d18c447b692d2ede47fa410551ec2214a06a5c05265d5318cb3fb92bdb53de832
z47ed6005c17d4b94628b77aff4ef88f325220d9ad1aca9dcf5553f9cb3505b104c636834307552
z931aca2063f47a844d117f952a4998192f658551f6c9a8fe1f9c38733231526ceb5f5ea2676c60
zc69336bc8e39ca79353a905798e5924b647937ba362657c8d4f3e2e847cefc8b1a4be91f8d0372
z2e4ce0afee2a16caf94e33297737bc0da5b9b5bf6d6c9ef5fc5efe50f5c5144d310995f3310def
zbce6bf9e59983c55a9ef6cd100609af842227bf34f9b81da899be06248d58c44834f16e0c679b5
z363c89a7568348cabc0ac0a5e37932c3238c6bdf265c21c599952a14fe1c122bf20d2d1b99e500
zd9b858fbde1bdcf8943f9f4d851453437fcb3aeb5f3e8f4f14e2e92da1e4c7bfcbf23afdd1e059
z4dec8b0b51d1ddfa9828787a09e1f9da7627e0ad7b18392d4c588669593774e477a1355e4ffaef
z02c1d0dd60c6e892f9cb808846032f6b6f500ea1bb9ccc97b61ead138ed6d81aa7762a05bf1160
z5ea7abb98b3c4ae03de7974b99ffecc28b2f3307fd107711fee54a310a290f5d6e70014582d928
z8faf2a13200d816637f501dcf598a029a4a33f47bd6ab54835c61bc71dcb2cad2f4e755e4f8213
z3248d71f6155c8807299bc995f2f5a2c7f63d2800a91892add82fb4e7d9cf86677337ba860a24c
z84072d491a62cb3028af8204df0463d7a7a968e805f93765f33b80d239c62c003df09edc650833
z87512c85c38e79d206630a5ff03c39436d4241ec1a103dd84d568b728a9893bdbe756882dd9188
z92394fd0998961569bfd9d119a3d6f6eaa8a8ce217b179c81a10e81acec5eb5cd99057fbb0f07d
z653189f1a8f571943c8b022a5cb48e8cc839e922f994d7df9af30822994ec854853b9033d5da53
zbca14df6e42212d9625683e8d13064f51587c1708a08e121ef521474557ca1a19b9e15ccfe73bf
z33f226b2b1e0bb62fbbf988007edf85f32238ce1d7ab21fe34f916ac7cc6dc5422b906a79758c5
za8c727de86441e8a9fe58e8d0f3ae33297cd9298b6d42088d49774d1dbfc972e1c7531c0a7ee5e
z0d3f1ea8462029abfba95339b53d0535ab543f60df19ec271ddc3f82730cf78e45316909772c0e
ze2ae8200db371afd9d5510344a262e02cccadeeb5f8fe74022cc6a82b196f11a40624ffbb27b85
z2faefbdf6bc6e5db14001bf7b0d3b064b3cecb1afa1c974fba19f96dfaf78f4439cfaaf08cd0dd
za92cfde371d5c6c194dee4e9c03021a4333d4e8f91eac3c037665ac80c7eac471c790e9c950eb7
z196e23b7e89004741e32f305fa12f7f54489ead383561ec6951b1d1d8472d586878590b66dda3a
ze00e9b5cccdeb2cd89ca501c2035fcb70db3c5af8b1b47ea85e085b6d4ccbfcf2eb810bf80d23a
z7ec070bcf204fa0fd5d2a8e3c36c7412f290e6473e92ba0884ed23a8b62fd6e1ada1098141a90f
z4c73202959e946100cf3a21db951c5b4eed1949d510b75ad665811c068bc42a157699bb78e7a65
z69c7bb2d3b29844ca5f1e8b7055cc086b221b46af949c91335ab39844137d260a585a86f6cb13f
ze3dd98040f85e283acceb7a5cef74d67b16dc9ce7144009bf76bb2e1d90bb95ef62f4c3b29e0ed
z6d937affb385ea1a7503b7b0ab7de608a231b2821c8e0445b57e04d0a9bf9c2f4aeee420aca223
ze84af22fdbb7b22a071e195310a3c6ab6f4fb60bdb5ae22916dd2db26cf650c98bd783788080d5
z31f85b597cf48fa46108508dcf80eb0064cdf49f3776d4610aec3f56cc3a304d43a4217f227a7e
z4f869bd8f0c8914dbb1786f22d50a0eccee3694afc4926bd0450ae12a8c267fade1fc7ca897208
z0d453f255fc3f7ef640d1824f76c5b9547fc66f85fb389d1827d5e6af8053073176a38e183b66e
z918fa1e5dac70155f69caf73f46e7e6afccacbe890693fce25816e30fcf836c06add8e321a4a5c
z96694fe8f47d7a9068748d23756265d5868192a4f49385872a2ef8417a43075af1cfda4976568e
zf0713aa381daf30efb612c524c7876e768a50b1a9ee50f7bb598947b56838ec40f4c3ac2304080
z45faf26eb37526e56e2690ef0f2311ff385f128fa254ae35fd1c446adf401875cf22cd266d5994
zfec08feff26d4c70d02aef5f22e69db786f83924ce76561a2dd8e465e7f981ac67ce0ac74a7b42
z6809b75b40c7a9db26b042a6bc9b9ca52cacfa51cd70d4a555c19762d792e8c6b301475b8632d0
z210fd2db100aef396d9af1944a74f540d121780a7a31fd6aed9a2353324020f4554e2688d55cd2
zbc95dafe7b8f535de83d661023e3777932adf2d8b283360320fc6ac46c087f31cf64581bd4c769
z620066af84d853b59c10bf66b0c420584963c60fe0a96006076816f5e965966e5b777cbb6ca7dd
z58c98407e6e352e9e2f9de0cb2aa27d76448522dce3fc381ff86e744f2198d5f33ff222273df2f
zd4f8ade5d7ef6ba6c0c60ba4cd875da2ad83667600f9c6d367e3fbcf4bebb8e0d1fd87d8b500be
zd84bb22f2e2b5b8377c945362a39ee2ee75eff8a41f6e4ee2c92407e14c46d91b083f04a2ba5cc
zd4847cbb846784fd35b8d0078f1a78c3f46bb9830028303ef698adc0a666b534e3c120601e260a
z90504e87a0daac4bf61f9c94a70f60273c2b674878f32aae7dca0890b583b5c95f626cbafa17ad
z3fc73d043085b00ae6ca03c787d439a2e93d140ca10b5857d50acc6f78cbbd6f55995d5e0bd51c
z841c360d7c530fab38a22441338d6ee1ea3a4293b006f58126060e767a91dd3525e908566269c5
ze141f793966dea493d8b05489b215a81919db15dd4f3ad42ed77c985019959bebed3ae616c8cb3
z853263b2225db294b1837eb8120cb93de57506b2cf5e920c3abec4042ec756a9d7276752eeb3c3
ze83c25376db736b36d6359743147788979952c7ced9dfc93b3635470313c717df5db918261bbc0
zee52f27ff2f59f840b93b2883deb78024f9c6f2688bb8e77869adab661efcaeaf2beaf635837fe
z1d9a419d00fafbb68b55ed984a3513b908ed78c5fd0b3e88e52af918296a595b36f61de1dc085b
ze378c7d78f0924aafabf249bc2dba668608a3117e295732828e28e94fae36e724329f21f1ef55d
zd1e97f432d5f2c567e86d5376b02ed80323ee768b6cfa7599f63573de4b0143cd452904696ea92
za766309f44005d4aaf3c35d231ac4b29e76c6efac28a0d0d7a347ac938d7e12f1ff8b34a1f05b0
z674d896b164ef00d05ef42d15ae97358526dd1f3493d3fa554130a12c446bda9825c033a94548f
zc25e94486f82e7be4dc2287a3d9837750b246d19da109e76a7a6e54e5fc3df5820ab019af8ca49
z2ec0ff7e63c2205665055d3619a55ac8ee128cec95d9e59e9898ca90cbfb2091d50de0c0b19df6
zb05a68c3083f1fbef9066f4da25e357160bfdf6ae09c77f27b5061b04c7519265f01cf63b0fdef
z084bceb6a9ae288a306a38f07f3b67a232f4593d3d84ab2fb3d6d40ddd45f4e7a266d0d90cb6f5
z809e2b66994bae5959ec0f945b1a2d5dedf2fb0658ef2dea69464d05ba1e25837fd7bb830341ec
z84252da589634d336c7df96de772508b2bc372a3876d74195dc0ffd616e3313e5b66538aa6b46e
z89142103e0446a9a1af14fd59def76dc4ad51a412b0c858a3ee2f60633fec30ec21502433c73de
z633cef9b5181931f62fe0524c42cafb09a613df94410e14c3c77d4bad67c7e9a2baff794bcc097
z82591b9a9058da95c9ba8e288061775e2648e728f22917e2a07609c51f1e35ed83dab24a23b480
za0adbe4d0d8baadfb891a6e4cc678d297cde01e3fd49a667424a9fd38f985800ea651630a0fed9
za1f788099ba8a1ae3c855849c7549316075b1f6b971e6b65c1398ee88af65afd818be942f79e65
z0669fff4b96a2772c23f63f5584e8bd9139a6eaee1f7b0168799e57f31725ec13a2634934d75cc
z645f8527c2b1241dbe95cb73d7067e3d3f32916f7e3834269310d7d0fa5a046ec87dd7ce89cf44
zfa5c74ede16a65bfd9e421b9918de46030af03725f5e44654dc76e037c5c365216e7d26593721c
z5e8093aa33c5d95354774c6a124ea412d196902bb2e6f9ce2638e904ab68fdcab8d7ca1af9c1dd
z40f751641afffb8a5878f28f4f6cf80e6905f64118e2896723aa5abde4806fa8c561fcbd57e921
zd5379005ec54aa072896837ac21a22f67122f52761fd9e5ae84839a8b045f36ed1e06e3d26b3de
z8d4e70557645ed42848fd4d88950f4521296b57d0179363124a545c444a78d7106053443cf16c0
zddf642adb2f257d9d0fe4a7bf3fa0e0d66c8aeb6cc85d0ae36335643726b64957aae8bd2c5232a
z47ceca1a3f129734375520eb5f47b46129366d9360373536f87f76de2287b683116faf915e6438
zab076918fe4d1704da875c996b93fcd792bbd1111c31a14c2b0967a07a43fe4ad41e22bbe1ec71
z023d429ea424c39c6dc67beb30e5a859950758ec20507cc48c004494e188000c889c2502afa0d6
z63e823a0e8a67ec3282fd1de59008c1304755449bad962bb2a3fe2dc2f1707e1d7747856be2d46
z51b20490739442194e680c6f29cbdb4dbdfaff076146203318e3cdbe3ef01f8b30fbd008b7d907
zcaf83f2b7a8a0c926a01d506ab8bb51c11140d6900d33e2a613426bfbe983217d281c5881f9ea9
z6355cfb7277da4936c6102c3954ff7ed8888a8d7a5369d8171d9c64afc13bb10fd86f190cdebea
z925cd61914e39a4c34625185b9cab6d0b184e6f835d32f6e208ea2dd39b9143d806b21847788bb
zca8259f528ac7fa3e9cf921ecc894dcf13964ec8ab7906b1c4b1e98b4de016f1c46ed1f1e7eae1
za14f8dbccd0863d143a5ad6fa65aca3d1da2b5cc31837ec53c337f47cf7ddf55a2c1e4216d747e
z48f9d3122562ee615d5df5a23442250f50f98368c5146b41cf2d7f1709a1d4de8b7c0e3542adad
za925ea298344dc6855d64699cfd83c2fe51c96ac590abe3d912f953e3b1ae3eb325c843397455d
zfd062028c8fd336670181399a0d319928d12b4fe585bc5350f594074f6fc42d696688d8db892a8
z86fb49ba287073df1c6b6771b06423641875315e12c5597a97b52d5dbb8ad00b33ba358a5b94e1
zc4a0813470f04b8452c2cef15b776e799231f5d3ad2b4d292eb164bc6ad01086b70185c7ecdbdf
z0bf15bef4a8d4ec3acac793d02ba7d3bdfb1013ebf44954ecea467f5d951bcec8ef2a6763c8922
ze7f78399a95d30a061691a169ede522a09aa3e3e33311942576e50a161307606f971b410c87b8c
z64e1602b4ed84b452f01c011fc5b9895056a001862a69b1b9bbc3211f84c0d719d155ac8ea9b1a
z62820e28dafe50ce3174fe41ce8a14573f97cef2ad719966f7ca6678a707a4526a8cae4d2ede0e
z08a7b5f01cf28da6ca0d70326a4111aeffa4c06c747c3b7479e2c8a2a69d507e695f8d58c92ce9
z9999f1ecbf998b1a4ed418ea45d97f0eb67b1caeab754d7aed4a6dc681b2708711d6da1c845cd1
zc28a115e71667a17f383612c9a365f54a999a5f5e3db3e5a3920e2777f1126a47e0499ba24bc21
z7b0306e1eb7d903b9df8a403ab16151004739d8178963fb3621c08c5e0770008e0a1a4611391e2
z07814e710679ed69ce33acbe930548adbbef1d68953340dbff03b7fb4962dd516137ca27a9ec53
z388b8c1ab0c8137872ea260b26e9029ee02d507cdb22593be7ef93156db703e42b9bee435c4db4
zb2f1805c6ca61c604ad5cef84e27bacd46ce3332d3c0581a3428c3943b33015a2d40ffb60899c3
zd3b9fcff877c287552e1e2af4c464cc7606e94c5b834ed6ba0fec8b6fdd7cebcf6379789eb6a17
z85f2cac3b22e0930449613a46f65f528a69f682616cb58e7f37760e2ebff5eda3f72fa83011a0d
zb7e4ec0f6a385d397b06c4d0e3e478fc57a4c4d0c9a342d7815ed6df5b4d05ec592751bd3b1ea3
z1343ac2bb1206b72ba0355ee36e69decec12e25c9245970878e68066fc74b4944b5dff92c8920c
zdd7bc2dba1417a384e92f9e5c08c83d0cd74ea2bc91103d96124a301670d150b7d899f4262fc34
zba1e30d2d5c1df82365493ed0714b6c46762e91eb1afff019819c2ead9ca804fe0382b5a52a98d
z28d0ff7e0b43cf5e7a394b6e6b5685f0101dd23f02be17465a80615db351585f307dda6673887b
z5fb88b03445d9ef21bf4fe1a7a9f56d7d6a95dcffcb3f3dbf66c6f37213b8f2e64925bede480cd
zbecd582907b71704eb8f0bbb562c2afa9442f2c492970e343eeef4e691ea1c445b7061878314b4
z5313ec7533b69d646779effe86c0a3271f76507d6267c478b076485eac0ef4db56993a5ceda5f3
z9958d349cc395965c8958e9fc5fc474072b592951158231985496808dc1f9655d68156d37ed8dc
zf62c254caa02aa573b90b2492f49c4d4597f726fee6ac779e5967316153f2f126eaa2ac8546ce1
z5b2cd717b5a727e8147beb46a594ed912eb226b1d24eaa3453a5bea34dbc7246519095362db017
z520b7d54593518bbe94af986470f3ca7e2e008434830e352b6a7087ffaa27b2c072563e8a0cad9
z71942992a09c16bf667ad6763c537bf2303a649a0b6c13e5d1cd756a80bcdd00ec65ec04777eb1
z53cc520a62fb39d7bbe444dde2a59fa62cbac5ca84ebe9499a25a3d7bd731746ac76a0ba59a8e8
zec2e661baf53cdf6f233da67c2d14ba5bb518885f6f163e659bb5f011b7f25218cf5799c0423ee
z3873317467be1108bbc24955305ed09f6611eeb0a23b0c100a243314a772d08d2ffc192a58abb3
z9b1e4f9ed36430d02c2496a3229f245090d9bb4a1d3251d68c3ef9a82d17c6f43227d2e87a3f11
z9f0b9051afeef6fe55a1ae0964009c94f7d9ad19e639509070598d3876085f60af77669b089dd1
z58324a63ffe865093b25393fb906fc76f3b5c8bc60bab3b22f3502dfedc070374702566fb2fcb2
z5fd1c9a5277e074081ba9a3be255eb9bd7acf1afab3df38f6cae3efb924e19734e69c2cf67dd22
zdb5741d9ba49bee2884faaffa7fd916e1da9a2381fdb15b21d620aa01fae4ce151a0f8ef0de7bd
za7c568af426524ffde1b01a1966d737f9b6958d75dc9073ddecc36d8205e8fa05b0a0f890749de
z6b516ee250195d1013a2fab07e3cd00ed46ecf402cb214bde684a14b5050924dd81b4e97153609
zc64e9a364e23d415e10634c48079dcf5dbb36dc6425f56fead5fd70bed85365cc2acdfe66e74db
zf6215cc05fe2240a101fe047aed2a4b000ebea76277c7229e49474e1a7651ad052f607c24ff515
z5caa4889a3c4c8906dcdf5d160df193ddd1739ef39842f5b64a56d06b8b761b0b78a5c9222d6be
z5adea3cdbcb1570188d7856542b25c503bda7f0dc57869e91f2119a173603384272af56d5a321e
z58285c643a61f20923e1af432eec8fceb32c3aba9ecc014c270742f647b4ff7a10115f284e8881
z2b1a7dab681594deb5f9143ffa5ded6f4e6e2e156ecd3017ac051df0cdddcabb1b556fde1b30bd
zeba39580e6072a7ec9bf4bd6b09a0339607949feb75a881bbcfc43756ff967455c5b8aeae8d43e
z19f1fb88a942ae8c34a417360fdf30698be0e68f17fb7e320de7d1f9fb69b9752d175248f49199
zf37f1388a199f637480aaae492b4f421087c135b99411ea720b8a43169d5f685662ff95d746f3a
z62f7a2075440476e5cc89057e2f5a187abc8e14530209ad3720d3decae3cace18afbc05accc8fb
zb74f1900ba9d9605f491c0ec4672066787c2f3550b89a1a7ce78349cefa9be7400a7fce284843a
zd9cdff2e0dad5a6ceabe9ccf742026a5c986c47c8b9abc7f9fe7f6ec152f78eac3645b4783cb40
za7d1aabd407d482c5cb3fec4cad384f4a23da1da1b6c777be66c89c65b3e0918cfd61b324b5dc8
zdaec7e106f7a6bb23b66b4a4b6ca7fd342789b017dae8f3d0a1ac1f5d83e3025c3ba3fae0b96c1
z5ed1cdcf995be7c9dc64499c166ec4c0061dec5f0eabed37a33efb3fffa9302bb06bb0d3ab5e6d
zee2ed130d45b8e17233bcff522250d688db048ebdfbb395e55aacaf550c813df00deb9d63d8fcf
z1fdce8c5e082bb634961eb285e1dacee01210b632fe53a541fa4d6f3a6ddeda67ec6cf64eb4d7d
z0ce01a9c9874d1006724fd5d5910fa8f3910f0f5fe9fec98dcdc5aec06d20954da514df5bc0b70
z77239529725b0def7a98ba7cd984592f01c241facd1b3cef3c51019099b4c69adf8e5820518323
za56b36054d4f30fff6a2f0ec8c313f66449e27084ad846fc09d5ab0436e79b8b3c320fd1dbcb67
zffef831ec7bc784be33658e044ae1ac9a42751b62dadb2c0a19b4d1621d304741261a258994375
z32272f766352756badc8967b8940cb00139af1c55e8a8876bd27d59302c9d256afd10b69ca37d6
zef083b7899af78508c7870b4c5c28ff4eb81eb2ef082c1a0f886e3a3dc83e481dbf219e63341bb
zcc3ced4d2ae293b0bc3cb0e98cb19800056d3140877dcba35fdc8b54bef995132f9c6e007d8436
ze88513631e2e2f63b9045d5e657de1bc077f1bc56cfcd15c92f1ed03d2158963875dc863ad1d6e
z3196ecc528d018fe9e4e7ad11c0f5c3e0cd26e6516e3c87c9995f277fea31221ee72b4c867d090
z9b24d3ebebb03837cbff5c91d1abf2c90dfa1565c9ae455317bc364d36733280b8d3f867d1d5c6
z3950ea51a60caa797f1ebe12f9a5f5d7434b07d4c031ccf94836da0e76a360fbe8ad66c1a57573
z6bd47e3329baf69ee9daad62a9b04f2599a81c21cc430350d41eabd6ca2f4ec3509508369543fa
z825c9601d56991a90fac8cf569c742d0b287446dfcf27cbede35cb4c3defb0295cefc27a10e8cc
z8c2b2f5e78a2ede3aee5f80409690b90681cd9ee02d34e521b28720eb4e36bbe6eb234c0bec6f9
z5846f69c605fc003d1455a651a1b365826246026923d06903fffdcf7a80e24cc97db281e22dea9
zba2eaf57bc231166d8af4091fe170a4fa9be7e942e38d27686ac7ddd8740e0525fb6b21808f600
ze5949d3ffd86506021801f0ad70d56d3ffcfb4861615f88e9b795ef70c3cb8087d1d00e78e0ca0
zfb04c475082fc115b307b58c8b2f33d00fa3e9650f03091ac249404b8b89178e9dd195502a29bc
z969a19e2ea873b8afb1c74d70a5ed76ba4fe679cdf10a06e5971504824a0e2fe111859e6fd1ba0
z5849bae66517ff2ac4a6c62460812695f581f7db9f071fa3a2453aac8b78753653eacea63b478c
zb335594e52c91529bef9afeeb8cd9a6dac24ad880a472514b879ed4b58630107ced7f4675ef32a
z11bfa916ff37506e918e358c80ab3e0512a69a233a3286f34619367a0f1a8c7c4b7fc5104e0633
z61d262aed5a66fd3a8bfaa9d2c27b21073ad5cc8008208ce1e00367b1b642ab02cf5718faa7d69
zce345fb5b84e84149f972a9bdfc9b4c66c347e512e1e620c6857390cff5bd233d56d742b0475b9
z17bf0f04690f260396e735fd5885b67367ae0acd70bbd8e53bb3083f1743bcb521a8993dd3197d
z870d84899bd29fee6ae41e19ce4a19e58978998a3c42a717b4b1c0f0d16eadb8a7443608eb39f6
z38788d5359b704acaf92c44229d6b8a3301b8e908555430c3beb02c18403cb6bff960efaf6fb12
zc1b64af230a350ac3681346d954a1ca78d02af688ee3f048a5c394ec8ae1d39279949d97be8df8
z8602fc6338c6afcf53723f37b5785fc7aebf1e97ff269f25bbf2057659d79dd4b1969651d508ab
ze0e7a76aba4c6002286e38b62303e3ed445b35085868841d5bd2f39639a7578053fdacfdeb895d
z56d114e01d1da1391c58a8576920390b797bf456fc2c4a888fdb55983b03892a00b2b92801e439
z3ae9d6f33aeeedea366fecbbb5a27026680e2bf63d2f3f21193e417315231962224a06d5947b6c
z2f243b15a259c52390ba0687ee06994bc1c044dcc92c03cf2a428e57e57f69f1c0c8035bdf0df4
za3b5f5ed9674af88b54882d669ba28f1306d630aa37e41ae13445c316833e7565063965834a746
z2caff753ad04b6a049d7239b1c55535ad7d36f44b0d6f7594ec4993293d971c760e6a7a40fe8c3
z625e781e4454609b9e1b70ec479f5f070fd4ee228ba19a5a13ba4286e255f5e8072cda483bcffa
z83c2d00601de6766612386a5d9f9eca483351cb9e4721db4d07b97290d587398eb6f06c9f477d9
z70c6c4ff72bff6504d4018bbfb392bc5fdb43bb84e359ea16a91dfdca0ce710a9135ee29596453
za7c83c6f67eefdcfe6881d3f04734f0639cd1b93e960b7f0489bddd05d7e92eb845de0ba0bb02a
z156098d7c965c7536876fd12d027845f3737b5371fcd0bc29de8f6ecb92ce480ed7809db3ebc4e
zf006752774f1de585ae022e2a0903116fdc589e74ac0e161440d07ffa75a81e25eb11057c4548f
z7cea97f696c7711cecffb9cad8d639a8e067540c4beba3b371de946078f5a44150abeaa983af8b
z6592d2d4d091fa8e984c52cd9858039b93f274c8d043403b80c195006a030dd85fb77a652805a4
z98cf89a1357150f5b6cf32b466f07b6c1f0a5e87f81d7ce0f74f33b0aefb089b5b5c8a30270d1e
zdece02cb79874740d79baef69aca4bf4afbc38c615437484f298beb9f2e1c46ac189dc582aee09
z98f8e57e707983b484b49367a5e8d9a029b4bdbd7f1627e4955bdb3596674755ab231420a9d04d
z53ef107f1286d12c6cf0e0d58a140277339503f6f3ee8372c4af2dda4b137affd7c44111321b6f
z6e5777a26d4fee59cce9675f44e40db20ff8a8cf13c815fc274139dac496cb227de413fced41a8
za8365799b83fc451befcacd3149cd26fd6f0b60e398603f37ffd86d22d2483b852f881c96e8454
z397dbb9224e8e93dec422e9f18bb898d8681ca8be6119bf407259290fe34d5aadfbb0b5e52dc8d
zf4b1fa7a3d9a79ce4f1d30018ea00235642504982c49cb048e31218f789662a4ab6db50809aa33
zfd03b9e7a56e5f59e0832d1ab67cd940d8bb1087743e6e16ad4a9a5f9ef03f00435ce392209767
zdb31aa76ddaa05f46303dc75e4ecd0509b80447686632604a1c7f5e864a7acc7d9cd3c3dbe28c3
z9b7ab11a081fe420e62b630ca8616cde50f50a9053666cd916a5e53632483f4e52b9d539f0e1b3
zacbd950eab24e973d49e4f27c749413c8285bee9adc500bf6cc0bf898beebd8221a690c5ea6fc4
zf38abf67d229f3fb22de73787195fcc17ad487f1f38470a65f61032056a47c3650899e50123f4c
z71e88237f981ec7fa2a87a300209cc7f41ba31018964ad36d4906497205572ca9aa8618d6b6f17
zfce616128462cdcf99949a4caa38437d2e1e3c075035bcafa2e3e74968ad5605e239547f4071c7
z53a5a9fa8c7ebb3f60ee5cd65d59c970c2f6031a78c1d4c32395145f24a8c7a460545e46a1d7ab
z16ea7705e4dcd5477fa0347f62fa4eeacd9196dc7f7693574671b597c3205576aff13bb8af5aa1
z04295d28be07bd1c7bca31920d7b8b3e96e564234a5b8695366333b2f034ea4ee7dcaa288c199c
zc420e935e8a345a17b8f657266c9f02a1e683f6cab2b001e33bb449ab919f757ba4e46ed974f4b
z5489e98618802f7b45290c118ae8c8162e541bcde3ff5f8e0bea9e05325e5af503d9000abe8895
z3a1bb8e658102510cea9eb032ff98b8ab2ab9e4cc7e9cbdafc0531008eeca837ac88242f11f547
z26a9bdbdad4f2beb27b8154a082726ffdc7990d18def638328caabe600b5913cb77bdcae823dfe
z341658136fef1ede518abff5a4ab60ac5203681b098848638811367277c28b117660ee390cc908
zbea77f957da3266a789d0ced7a135f81ce4d0128d80ec62938f42c383ade15be93844aa1e0319b
z3895ad829b70a32dde0b530d81bbe6e084acd2149bf36035ac401ec4c06905adc1b017f5164346
za7e31d8f87fcae99243aabad5ed82d7d4237732742489afe8af406c9dbea438c2fda7261672887
zd4bb6b33009affa6d2144aab9d37408486d17aef817f3296193d6606004e3dba9979c5178beb70
zceeb4ff7c4ad21c0efb403d5709052ccd02c9ff3d8945c5ae473daf7178086604cb179362e611d
z9a721dccc5ade7f6a82257ddaebed2d8094311bdcf40476bfdfcd823c8fcf0bf498e0c64fef632
z2f2567c4721bfa9b04dbb36112ae39be69ec69143f33c89a97e622f9f4677d27576bcd91e3d546
z2c0b147719ed6132c47c9467c921a709c5119754e4ed86e202031907b77ebe6978474a2325e385
zc286d363bd3f19dc649a7fb14bc5b8d4248a663ea1cb434144224e90fc2963a7bacd756f1274e4
z5e4e7c33d435e4463e5dfa7f7e934b57b326ed7222f5389030c31722bfa1ab8489a02c276d6a1d
z60cf39908898a03c37fba5a3d375c130e7450db62ec5a82b6ecc4fe461e7cb27952ffae97583ad
zea882e566e0de66efef5ddbb5d12cb5a59d3a44ede17207fa6ec4fa6486b2593cc06bc6845cba2
z8427be62131cb9f33b9903cb40310160fb928d02cf8acb5700845dab484b27fff9c2d0abbbecf8
z7ef67450bc46fd61ebb51240c389dffbdf9f7473ad18df00a4094a49e07948b34d9bddd05c9e3f
zc0b75d58757c70196675d7eff253800d37e2bd3af5b05688202fba9c81a6cdf76ae45d4d347840
zd9ae7982fec678ec8f670b7726c941ac5f611619361ab5ced113158907bb178fcb2365c355e772
z60092a32c06f6aa7a4a5079b52befc4739918c678963e06959ef26d7dd9087961dfbdbe8c94bcd
zeed1086154a901cfe38863ea76905f67ad7a874c23cdd78671fb7a0972cf3197887ac07f165119
z7d71addea217fceee7e63bbab99f5bd9748ec90afaf6c9e790a75bf211bebd8378e2427545e844
z9d842381cb42c9beb387115a70d03860408a46467533350f20f3d732c852ac7b47cbeae73146b6
zf7aaf7d05c0afcfce671b4a417dd9069d24b208b885e974dd55c4ca8361ece07fe65e5781c7aac
zd950b76d82bedb66c36caa280352660ced9f09a72ca0b9763f489b02ad731dffbf6701f7b5627a
zcfddb9560e4039f119d2003719abfc216de4db1a0f47f15d0e3e6525f96d956d8075dc7b35c424
z101c6faa5517849ef97b0b32df7861bcc453c0bf4f56c17d1190128f7bd334910bdfb1f2f9c00a
zd4847bc1a5a02c837fa4f8937b3639fbfe638c4bf8974a935b7ca63b58d995c1620cdecdfcbe18
zf12d749aa529c811212dad61927591a34aa01a14818da69a73423d5a47c4a701a1922881f790ad
z9fbf81ff86f022bb8618f0712e95417934426f0fabcb14602b1b81d874cefe8ebbc4929c1dfdcd
z831ee9b7eee43554607d3fc9ebff6d49c8b1c0c965b91b01910a39b15c1d31ae18c9b56f18a48c
z89b2f35b4da7614c39706cdcd044aeca261c0dcca6f413278311adc928c120df0e7ab3cb23bd7e
z4fd679541c7041be925779696a2094519a7ad40be3c9a389747338d7f41a058b2f83d1b1817416
zcdc51fb640e35c01c0c36b15a03dc60d57478fc01222e28258299e65072e3035a9caa48f0c2de3
z783caf7ead7b7fa025c75fc51919c57d6e5c1e1ddc1ccce7d7ee154c36d96de6cfe682dd188989
zdacf49e3de33e5fbff6f04075ab80e3bafddd4482cc49c558aa262f44d0343fd26869bbd09107e
z1f8eba477bad9eaa194bdd966bc259b87eab708251130b6879642cad3032a7a5969ef789dd3fe4
za93546e4498b2d96aa6bd40e3ab0f03c4f8e2e59350c0a3868ca675accc01e4632c5df1180a0de
z6f2caaa7e1eedb21ee0340ddfca9667fc17a0ff731641d4c1f12787289c4019ac8e93029724729
zdc407040c32cad4cf469bc77a5cc3a3740558f26ef3b9eaf34e9955851fe6de874c0f2604a8096
z507f804c27ee6617137ef70b10e28a9ac0b81abaea3e4932eccbd89ac7bc1e912f51318e169fb2
z4e8d9b6f130fdbc92c22aeec3fdd4e3a6ca64e262dac7e2b4dab629ed06f7c741b7099fa8b3e95
z76e4e146fd12a681d915e5a98f6f002837a39c161ce4d3e26fc09d7fb4dc74574dd3dda7471da6
z9f4667c82cbd09d91cd8a2f8800e6d00370418556e359c79f14fc7f5918509c1579f8481d96e53
z33873facd8408a113bd38718062a6fbfc20c373dd5d7839454f548ce54207b88c3f5b679ab0f24
z32de655242b07e381a3b0d9db219b78ce73bde7684fe180a7f51272c5f8cc0c7b82833b33cc6d1
z68f98aa7c97317b2d53fd990aa53ad55362e65d7a2b9b2df9f0b7e63549b445a6dafb58ffaca71
zdc5770515af6789b3925305e8490588a0b017d4ebb208381a5d7ea40dfedb92589fae96b8bc798
z9d3e666beadbbacc57ae8b617c062806cc515e074d55439e8c7984c905e4fc294c843ff784ba2b
ze352f229f181854553d7fa937e592995cb10314ea3f8a27f755ddfb7928dfa15ea591d670e847e
zfc3870980394514daf61bee1051230d7da6a3eec5a99a28e9b3dc14b1de82d5d7bede76438f2f6
za61413785b1a4be51147d2cf4b74a7de6814a43ae87fe5931b5269e58ee05c838059d94b224289
zc26a5fd58419467661e104844851ede510e750e7e9773a45756e9e664693f3aaeebb19f2de5218
zb3a24261f95ac54f712dd4f16cb0d5bf93bfef63db5e68c8698de16ed211e8397fc6ac40016c05
zb8b5d74d20a41eaf1d2ff6f3fb6ef84ff93c009a17ce2fcdd2934def287fcff8c28bcb6a8f1983
z4f413a5ef3a9df8c7f71d22abf4403f65288f1936c1783f2d414db6c411611d568f0437b3ec6a5
zfe143af4a2948e311b1e54dc16453adcf7d02b52c7d1842dce14caad9747b4a253e303eade1730
zb0594d4339f876f99a94d7f2b075eb70ef43e2d155ac7b219b0a79d1c9bb9f4b238b97945aa5db
za7f8a08f40383c582ae6eeb09f098b5f8cc53a166b5b6affa7de7341400e2b56a866a59f266d78
z6725f7ece227b515d3fb3d5f3d1e42b8b50663166c2d2116a6d717be399b30dd105078b26b465a
z5d3e588ae31365190f007614b5469d4dd77785a723a75c0eed5b3b2690a044674002efd2549bc2
z5abb3d1e6c39e7e4d1181cf4801eaf9c7551fb612b6c40769efae7d4ba995afc60fb5f6466f20b
z8d981bec5b185ac36025743dd449a41466cdfc1e5f83dc4af95950464c737d7b9bcceaacac1a0f
zf6f3e3362ffe6b151d1c6ef76300e24fe462f3a39198081b4219201c34231ee18625b1b20e5882
zf3109079d0796925b9599fb4c02fbdee8a9651a7024900354a8f77f1186c858e799a7dbe8ff1a3
zee24a66a2ea9bd810677ebde8aefc3f50eef1a45ed204241b8417ddf450300129fb090cba8af54
z2b68fc5f52ecc11060c02abaa4b5f98b5e88519ac14cda107a2ffb4df4bdc270a4405e601e24c0
zc7eb82d43a7f12304cd319b61ed3f47762a168568bae3d243e2bd3fb4d4db4b38893261e003216
z0e6c0a45365268149ea083fe9375608c7085e48bd8e84214fd3bb39519a23e8ed3bdc5184f6e04
z29f65e9a7953630edad3d69ae4661eaf584c4f86f8d8f639903b3afba47a93b041cdde28d74148
z4327c1242281a70e9701b66a27718631937c2b47968e81539e891a1a41d294c0a0625f81ae2f6b
za7e8d0050ce630c3ad40f9457b61b8825a1a0f904bf6267b215c16068e2785dd2c25f348752fda
zbb6c7b3a6e49d730b4a39338e1e42447a8aa778187be94bbd61fe10dbec7ce8361704a7c22f347
zf8bd1ade7d86efce9f0c2df1e266cf36ef6f73550f4fc95ece99dc8fce45f69aa44d102ab257c2
z3d209afeeb1f8685eec444029c98a845cbde6ecf7925f2b2ab38f2a62476514e18fe3bf08a24fd
zcb6685971996df90a28fb2a6fa38b7b0e345ec11b880a9ae05b36ae5ebe1d42fee6c3c9b786157
z18741cbcb3c67c54e19bbbad7a49a686df12ebf5ffd894c23b1172102cbeeb07954af9f54c1668
zf869baa6311da6c0b1421f68d632dbc774b1fd6666de25514ca000004d1a44dfaa92f29c844fea
zae233668ed5ca4028a8cec441e98beeb29b99986a311fe6763cf7c58bbff097faf22e944a02b74
ze717e7da51d00564638a051f53e8027308fa9293778efdacb3deffef6f3931047002d5f576cb84
z1f697f287a13c0d6c4ae465f84d4376adadc87bd463040ab7abf1b835f31fd5a8017b2724b125e
zb42dc0c8606088980666c3a32b260d7c64a90e4791006ad7470a9ca33e20660f9a8ddafac56c5b
zc64f76a962ac010b344561860f257203c11a2ecd3826484eb160e5939290d7207353986a07a897
z1965a346e14cfe979272725fa855e9a204b855a203c18cce7810c0f42299b5eab261a94cf80064
z9b005eea25f703c8504a3ce5c5c245ced921f96fb9b63aa03f736e02492746eb1c0193bf6ea0e0
z55a6a5ecc2c467023696a627ad302c2f4a66eb4547a88931c3516099a46bc0a45cbc0c40664584
z79d8f6b2889d6d5abdec05db53e6d81d8bda98a99d7f6a7a8fd5b57dba4e0e6bf3053408dc7a71
z45f6915db08522533d47104cfcbc7fec08af59099bf403cecb8b74f7a383f0944e14d68846e945
zd0c6d231ed97662e2b29d821b0571d44a33359ea34d113d3d0c4998f5c6362d538771b5a3d57dc
za618ba9785cdd60c1135c806319853e5e90b53f733763589a2efb7ead75dff7a6c52f93a0032f4
z5c10438f93faf42ff4ff1b595da622ef9ab143fb241df7d2ec0286d04fb526cf03ad756208ffa4
z369dbf2aa5cf25d342790f8fa722e22634475077abf7d741c603f80e0ba2486f5e8e4db71f40e0
z073aee920ae2d1623c5f62560c2de5728495c99d450f5772d0a7ae4ba393eb55bf7f64834206bc
zba7d52e0e2a367ff1d8efb62c42f2ab0521f87a97afa5785d942786af5e167c1fda808d4a6fc8a
zac3d06a8ffb58c9b4b48f079a7c53bd76d9dc95977132dc5974ad8d7783afaef11eb4a3d59b3bf
zbcf9cc56aeae4a89b47d91cbc5263edaab966200a784cfe973724310884e1d5c7b389104211530
z156d47f5c03473f14f6ef71104a2d747cb6ab2ecf7d433e5e2ce9367e48b35bece12fa22af42fb
z78ee872b89df9a3bb3857dd112f8866c6eb2d84e257aeb6fd51178a9f1bbca6a8dcefe988f0f93
zc4919d815ca93f088cd52702cedbadd1144938b9ed1a5111be1e9afff2b24494d642064f5f143a
z3e8aee176dde88918e912ac4ea9e9eb97a95975200a26385e0cd678a6865c09d8292b1efc190bb
zd65e8ad8b94e98e7d0d532863ba63e2ff6b238e87cc7d8ba2808c848858ba2a194daf488f41e74
z30e2a098eb90a3b4e5f1fef7994f0d7e7268f545a957911eccefda41782deccbe1bc430cabb2ec
z06b7dcfce793eba0e23413c0a6288de7392b0dccbde6b560eee7f06ffe527df8a88c0320356a9a
zc0404516ddd2095733227d2e255cd773452a2c8c0e6f8ed0e561db4cf32dc11f470c016281b689
zfd40e516699e967e022861c1f9da9512f4c1a554cdce5a539270f01985d08199fc3fb6699960dd
zb479e5192f60e280daa8ba2dae9cc24588ac488ff0219d1282790fec92d9d2197dbc90e1f93bc2
zc173e724f0c72f79f84ccae636826a0c6a45b557f77d6ad31765c334ae65ca9650bd5a57bf897c
z428fce0b1766402125643a4975fae6febae248adf1aabbebe8b9cf19240ea41fa2a8ccc33c76e2
zdea055f075c126bda772bb53dc24dce866334c2a0b19ecd704992b6f62c3640663c20a2b49e2ce
z50eba5c76244cc63ef56a6c2cc318982ad88eb998fc6438b30f1372257196f079a150bfbc0bd2e
z02462da8076fa60a53e30de3c00968109394b80a1eb46df0593dcdbd50c8aaad3f1fc76fa55905
z0484e8f4dd29cda3915d66e00f05c8abb012bfa1968bccde70666f9cf1eae24d68332380c26f7c
za0b4b1f5eb98e65f1e77f7aa926e2bb6175e1b40c697a5ab0aeb26238ddbe191b7dd4c4b51d58c
z5c6c7b0b7dc3a1c22be046c5a910d039860c625610f21294b6e7d3ce1ca8cb2a0104c9ff6302d2
z357fa5820917a443ac579e9fdb1937ad5ce7ba32b5b426328671a50ba5916f8c10df77a7eecabc
z87cee288ddc95e58a10d431d7432e8e89fbe85a384b8d9ae6ca095b9fbeeffc64f11b65f637bdc
z517555b6960bbbe2265542437f75ef5053149b24140975c4958071f3266b008248bea2c02062f7
z6b3633687124047234f23beec950a20f4a8a6442f5d1e64b5d9cf48c3e2d3b6553e3386caa987b
ze6a92ccc37c15567c087a58e83c4258d748c3f9e79d06eae80d79dd3e52a37cf66d0342164de2f
zf7dafea76c0eaff72dd7137061d17f47a59c1767377d3bbdfbf64c5905d879a3d76afb3d4dbee1
z77b80c054d56ee2dba292e745eefc61cf0f5dba80c770065171f8a37b597056eb80016c7e4a505
z00c59b8e41adea3da69860f46c4ed905fe8dfccc30791fdbf0c8e423d92768cd09a1581749ebdd
z006941554cc883e67cd9ed9959fa52fe18de6beb8dd56e0edf277e912d3f581c3f49d37ef0cbc7
zcd41a131e377a49940c0045cbb3750a0bba96cf13ec750be80f168230efef23f88f0e246d90e0f
zef05918f1cb6c6f7d1667f035b65b0eb63b0d0145badcf1d27044453696d14657444a707433f3c
z86b7b1b7dfef8cf1c744813274bfdb1ad3dd81f746c6e5cd354e0248b464a28be4e64b962425f5
z1631de5f9407dc7c48befb85ed3e31dd5772aa220e7aba730cf2d6bb1f2a5d45e5c274ae6e95f6
ze531048869f34c0cd589d56a7b9d00db0a7575e58a3bb66ffb95cf3057a4b28d10ae6c4f28fa27
z393f01d22923ad4b2478d140d8f5a46f1f32d0aa062a31f5c1e57e5b86851d2c11dfcf3db5d71f
z77ca6eef5a54419bcce5b0b089b05b1897ebe718b02ba03286fe5f200bb19f7fe243e66ff50f97
z7ab0792273e5a59da9e22f0d00f3bfaeffa6bfbce29b562375122994bc9f1e91377268c6fc56d1
zaf5c41484e40f88914527c31706bdb7ec0223f0a0f24e9c715597024c59fe57e5649ab2a77a7ec
z9621d2cebe7827ab76b5639a7e39ac0b0545dbd776b6e406015af5dc845ea69963c3f207d3e56e
z933fd65c1e35fb821dadabfb8c70c3d44aa9492c01e95f7a33aa2d29a77a06b97865ebcbe8841c
z55f7c38e7d6f7cb740b20c210382142bdbe2651dcd5b4b9ccb33ddf5a5aa7dc808a076b1a9403b
z33f47b2ddb97df1b705b89668f420e6ca452d96d2d52afe528e1874f01613fc432a55e6daf0d44
z213f218196bd343749d9e8fc1b3d206826a208f3be1d9bba1d1fca5d59982eceb9b6bdf2e371a9
zb44f2ba65b6b939ce3dafb0c5da544d888eda317cb2670a9f2444fa207332ec095bf9c8bd85d24
z470d59569c343ee617f9e5946d9ccc263fea9a95b2467e411c95ae3398d6587b706747bbc5edd2
z13e54c7b1fb197c93867fc65d9fa8587dc735fb6276097468839e44e375338b8001ae2e6db874f
zf47eb6d54e0aced13460a37aa438c706933c2548091bb39f3885c24a5ccc9eac62abe4500fccda
zed734172c062a9c4d7e794fd9369933f47939b22055efe00391e8bdd48421ea6b88314a12e49d7
ze2763a68f4e5b0ccb6c26137a570fc88d634c2d822f04efdf39b7a681c16b091ced84e5335437a
z610d77b24af01e17c8a546ad5ea27a31f7c4632c486a5c165110ebbb7585af43698a924e4bb4f2
zc7b9dce70eba0a71efc631ec38fd7e1e1016deeca2dfbaff48482f0e15cc7420a1a2b4ab1c3a1c
z59909ecd68df7d9112ed2d9ffcee93b9940451a1f8bfcd73ac4392ee1e132963791fe1ca508337
zac437a8ba68650a0f7ae9f58adb5ad21e048d8e70f554cd289ce41362496ea0ce998206fa13ae9
zc43595c6db32e842ce1e8a47ff0b6fb1e93fcb5e034ed3c130e78df6a6a9fceeb864d677aba865
z2a49cd50bf89e963621937f815ae2a6903faadb4a62e60571d86fdee6ed6a8d7e483f18f68cebd
z4eeaaa5ecabacf06c4aa3e4d291cb7760a357483373dd84de86cacda360eb327fe5bd46fa39789
ze417e7d3dd374928da37ffa2c481a3e3a319d21245de16e5ab606db65cf3e167ccf488faaa4cf6
za99d4092b6a4bd57d43d618b7e50a11deeec00808da11b9dbc0742e82af3cb2d45bc7f469dbad9
z1c28f4163917d58e6cea6474b29926cb198e44ff7a4b348a29bbabdd22229678309c16ecc76f1a
zd0a5c11549b7cb27a6525188b6bfc9144048ffa06327b130cc9bb33e22e7cba92de9a1c55d15c5
z043274cb229250662686dec64b86a4fe2e5b062996c4ef65b5261392f069f6492fa0400e8ffb15
zfdb06fdf2a170171588682520fbd476b56a31ff88926ed3e3be84292b2ba39ce169fc64099f3ad
z97c88487851a78914080a4f15f7c196540621aa62bf59e6a20b899c81757998559d73b3ff29309
z40eb9568c52c5d03fb860c2197595d98f9e07e0c6ab6fef7ef9093260e16bafe78fa5667da3587
z6c8a52418f728e741452b20d7e117cdd6980b8bba578779ea124559754b2a71aafb4d0dc6b85c7
ze1f8a4ee682b846e4f1367299972025346407a272c4366d84ecfb90a8e496ca5c8b6f89df05804
zb6e2ef0702d346471011f12415a12d518be56b111bb3242bc136ec0cb13c22d7dfac0a3743dddf
z87b244daaf264303228670b867f7079590ed1faf2aaa3638df7225f6309668beec7c1f53140552
z07c64735d00710b7cdb9e3a7ef0ae2c68be5ecd55e50a4c8d1339a68411928b133f53bd4ec1be2
zf211819029f7db20dd57fe7c1064d9d10eaa6a2c329f8a945dcd8c3d04200711edd053622f5991
z4bb55e0f124cd6026713aae719d22ea3f3c9cdb1abff97be292d47a5e24fa4a82d774edcc9bfa8
z0b4fe7b57c3a85ec6c6aa6b6794b2806924eafe71dca2f49083a999c7d45d214199d675fe93f94
z1cb560f0bd0b29008150ef9304e0177a1e3dab98943a178dfc01e89787517d39810d43eedeb700
zd40107fa3c555fe596e572ce02b56c807591016b934dff0d9e7addf6f549c4041635a61f37caed
zc66a2ae4c2bf7b5f89212cfdd999b51aaf4d0dd96f78fb1c0d9f674b983e98328ea449926711bf
zad85587863c63a3d112c8d0154586887bad7197256860280dfec03b4f98e26b2fdf0d5bf451466
z0337b9ac757edf9156ccbcb8bd80332cf92afeb33dfc7b84a8490d8b12939e3b699bb5df301b2d
z9e96c8e3b94d85f13c6a3d565c0da8cd1c6534be4b05406380d6beeb1bcb0118bbd554797655ee
z2b994d863b6b45bddc35def53e2f669ee1b43f259bbfed2f6ef2ff38ae299bda6ee327924fbbce
zb5a073fcb4edac0820eab5fcb555b2c62d8cdfa0d8a4dec54815aa973825b316bf6e001d5760e1
z629c82ee1720d1c1a72f204e0dd8207131d774a0137dc5472d6c610612620d741d31be183a1e4d
z12f9f6abd815cc2cce21f1d52d6ad85708121999feeeafbc51a027e142c14bdc9c85222e00e9ba
z368d26b691aea52e62b241efacf364ce4f09e83e7aa3464547fc0e947e10d26b6798fee5bd83f5
z616adecb0f04fffcdda9e82bba4f9cc5ed1ec4b2539094ae562fc5ca846e5cea8c625b3a615d56
z544d83e7d9da54f79a4f399eb09f79703e49554066c82007e6cda2b859c1946f1eab7ba08c5482
z8571e1e7c5ee4e1dcf316b96492d033aa5c5c73cd3494a41edb79d9acb1ec4c10037d1e594402b
z1a01b20bdd1b61526023f5555188d40639b0214706ffc2ad6a0f11af0babf3a6ebdac3bb7422c0
zfd4075ac00fca91e0c75bb2202a4316aed13303b054e89a2d2c2716391c93cb5e66d8f9f27fa67
za44c5ca9d950883b2345bc1bd1ce8a727ff7cde9f64b414cbe214e5f1908e1365226a27a7e54fa
zdc8d2557088d4f5024d906732619715d9f4dca1bc097d970b43462614493ae5db9b6f7a9016c76
z7ed36d029ca663edb2b4fd8ebdb8e1f882f8a397b820d0231222b0b80861891f0bc50a157f4c75
zcb3cc4ba585d4a0efb71a09dffb60777f6dd77e22749de093d1477f9582222721defc291a8297f
zf5499d1ce0dade85a43648ba0804b7c48aeb0088435aa04a4dd8eae38e311f5e84b128b77c6fdc
z010c0cf196e1e098bd7f824347c8d517e16f502f970c32c6f8216464e524f96e1354b4d853896c
zd21fd34e66a00604cadb1b3b66e5fa42b215d29e155840d3f5340f16ba41fdbc614361958fdc12
z0b580b801ba8b2b07feadfbaa42a2fce8827c68f45db0cb2c2ab490b99bf945931fb3e27c7af50
ze38b94d109d89aaa0337a6d6f66752f28238c25ad1dd76d0b82a85e145b6f35804a164a21c39cb
zc149957ab1e1d688232841afdb6c49a7a4cb0e826c9ccba6f719b4484207d4f3b6f14d9e0dea05
z3973a614922a12c9e3b4bff382093e6bd80f7e4bbaf7893b2892f6d7ebd31ef9016c035dbbe0a5
za19599d8e72840c4b935b11e193e20b89eaf86bae22fd7f9ae7f242a3ced9780f083a39a7494b6
z7c3e37321be633311bfda2d216633cbd54845c13ad5cd8fa31b1672ed889e957ea6d62a1cc915c
z45d99d2e1cbbe92dbcc830f9690bc40edec554ea399b405c9e33de494e3e8b09e690d03c9e1de4
z05e1d56deedf0cbe4debba1ed138841475abb2ec5436ed3431e5134952c7e8861daba3bca8fcd7
zf21cc55028953d4046f6dc651dc63f86959bfe50a308e621869930c12b80a63e1b2066c2b3d805
z9b26eb296513a41cf112269b690e7c1f97a6d8b6c9a8bd1fb37b5929b7e22c1541e59ed800c5b3
zee9016b380e6dbd1d976586f22200154d44fc53db30e060d8fdf4f04ddefefd311113d1d851f8e
zc8d366d22a31ea91807c9b1aebc1dc413ace03177ab147899a9785daa8a32b361c1b8fe09254c0
z9ede6162243a1dfdd5417d00a755a4bba07e041a7122ba70443413c793c2553929fdde4ab16903
zf0d1621a3baafbf822a87cb57c1d462e3138d911a2d439c54bdeb20a38fd592bea3b1a065c3add
z08485ebdcff2c17ca7f100c77770ee4ead75d9bd1584fffb2177d3a676a7aae401dd0b559738fe
zca76b9260788b451412f9117b1982262a84690af4dc0d088d8ef448f52d2255e2d4a45cfd960ee
z0b3d736417e43af5ab491d13124a135786c3294926595a831412aec42bc874e5dbe476920af342
z52efca2ed8a4712cb7c8a9414a4461b4555716ec34da4ba59641a668c83b157422d9b66d22032b
z97a8164cd647c5e0724938241100b5d22f783e84ffdda7ffc4a70b0c6aa0760d7434c35180603e
z89497ffd411fdf6269d71968758640bf2e0a80105b0baab692178ea34b49c7c9ed8274b77b2ae1
z865bd75392ed0ac6c434d121a6472a4857e5da404ed575602995187971d24a6c02604659b3daf8
z0ebcae31f57185e664b6acc50d7f6b113b65a1112998a6dd93872f63b658d405c6228380be2685
z4dd7510d217585cc707bbea35695f4bf16bcbd324b1bfc3101a265a5762454b061f368e0946cb1
z6cf7691dfa53c1690cbfbf864fc968b82914df9119af9741f50ca12c75c74f718446381701f8b0
z789ea5133ab84c842709c5c614817047c546e3adf9429f49da34670ace606beba4b53bcce696e3
zf0b56c4d0851c59cd5d973a6c68cd45b7865c81ba725102b2e47b8f0e70fb35d3a60a528414d39
za615567211bcd2229fa721f6fdb542336305933928414615fceb36a10bd478bd17d2ef03d90ca5
z971336e12fab0601f961445d5e2d7da4d05c234cdffd61e254e4ed39ef68da916eed3d7aebc2d2
zd9bffa78efd956c261deb0617a7e154e83ae36a1ced7d626529ed3f7e75608ac74037bcfa07bb4
z0ac017480bf42138a83f80ae18f04a8481ca6c069e8fcfd5f32e528c1a86de48aa061e9b011e4e
z20c1ff0e36c9656b12e59d963fabba1c06140eca9ab889b952358f2e9e4adc773833a9470ec7e9
z94b5c14ed77a8e0e908b1eff194ec538658a0800ddfa705202cdf80a1eb78358b62a511b80a132
zfaf43cc92df9cf26d933602e1ecc90a31adb674520a2454a23ad159caaa5c0e1d17e2247321c6e
z53ac0c6a73136021c66cb9f64d18ecc2db372c3c472090275bfa3e0637d24569d9ce8bc75d377d
zb2d2800fc659158ba43704c5c6a4dcdee5866a8f5522474b03ed8afc403689f2cd6d11aa2405f5
z95020b29f1dc81e5e42d0334e556a6294d175719f3c0febb5e505cf671043dae6308a5eca92986
z3229775eaa7e4f6654ce5819e050684d8ce66d8f67025cd2acdc9dcc62658c1bc4541ac9d9304a
z1b393666ab5690e03565a4301283b429803d6e04e6b7b10e4c790f991c4212de788de1510bb199
zde99850559f09815c5945952b92a71bfa9e79eb63b0ad2808480d7425bd5bb476657ddafe61f9b
zde437b2aaa881b8116f51002ddd28c62719ce522f29c909db039b191ec37e05dd7c66a08a1e681
zcfbe61dbd7803596a2c119a0ffb1814ac81758ceb6943e71be3164dd81e3a8120ad1427f75ed30
z27a0b2758d4b182b9b5d0878a007b2a6c34651603923192de03e7a547e3c18aca4b6bbbb8065c8
z57a2a82adf6eed9164f19396c1eb5690063239deb34c83a890e8d466db7cb130bc58f02fc361ea
zf544334b623652d10eda340c9d3f468460bef939089f38695319089eb066c420074ab18007ee00
zcd036b664f50392b5cf896feeb713307e80c6ceecb0cdff992fcc1bba8ceb4fe66807d240e77af
z00162d2f9c0d33c83a4825ab7c0d27c21da4cc9032071b095f85d2a0b70659e2bb85e8efa38a1c
zc67b1c55b38352b2f1ca18c47e9b0919bd3a48595f2f610f38240d3c9816797201406ebe6a4767
ze10d31dd69cf885843fc2c18ad87f922ed88fe09f134a441fcd23298570d3e2baf99a232107a3b
z8878a10c8d3611f710164f451175770eb96271575a532ccacf17e9c55720e3cf8b526b7d17f46a
z39fc0b1b5bf7fafcf01b4d0062245f478f4bd656d4088a46913d0617792cf9c31352d5a3b6712d
z6162aa8c6e7841d678d279438c8f6a18e0c493d344d397ad78a50c46ca6c10952e403a4bba3c47
z43a70dd08ecb71ae9eefd3b7bd6dd2e9987eb03ae134ef58e5de56b42f49637682c22d6830c5bd
z4fe420edcb590e285e5236129d7c926a57b2e21c02760d3662dcefc180a614f000f1c813b4343d
zb4c0ed1a119c314350fa4ace73a1d737552de4203a241666a1048b165ad389d5eef0d60f7d9d09
zfe01616a9fa2d2e4049340f88f912d2f86a7609819a1262978f974db06fd7faaf2cb657302692e
z48d40c2c547871eef34234788e2fc057b3720c4a6dfa0e014ac806a0e756240476103efc3fbe69
z00d86b06786e4a680ab0908a87d7b505909908948ef982fbc1364e417e8ea93a5aa2df55230189
z1aa635c5bdc577e438a09ab1168a2c4d37cee5da7700aceeabcfff981e3d62d8edd63ef4afd408
ze88bfdde77ab35c7748fdafea3e741e6bbce1b7e0f2d90f0961a62560301423c19427b7c08a92a
za714ff5afe130412b6adf8bdb07f77ed3a9fd373ed08e9c37590955c1f6484cefbdf5c15a87592
z83a317d80af04e64629430803c0252267902739e39d60ec3cb224622dd0c64680e9ae0aaa9519f
z9c6824384850e35815cc0973c8cd30905fca3d4a5b2278e4ccaed4e09473683d0493eed51033a6
z3173fca73f94980a7c481805c1b97906f40bc43ee569ce8cde7ac3074b5503af712b5b0d4de806
z7cac8f982d73a49305cd155257090067d22489cb7777d7f801b6e6440a1d7a2ce58c66fceee04b
zb3e4f4a2f0ec132886368ca07d4b63e5f4efc4ba0af41aca3d61843a78752f2b604a3c7a5c106c
z547aa932b269db8e80c1af94c1602075dcf4825e00aae355335ab47f26b7c3df67a9ae68c003b4
z0b13cff8aa630b99698bd6fbcd520677ad991e1b599471292be040a6603ebb1afbe4b7fc8b4a9b
zebbecc4d2add40ee71db2519a91de3beb0ebb14f391669a84bec01d2b8818a99f2e4e2ad8eff05
z08a6cdbcceb753146e289e78b6cbdfbde82110dbf9a5010a62b21459b0ecc5f7e36f693a21dea4
zf6a5b8cea3b323aec7539ee53ebb93c885e57f56e9a8ef1c8aa3664b2ee7bc06f95a208a795cfb
z317d544b137d0b2477c620db8ac1f7d90d4d16a85b3e93ac89bbec671b207159b2db1c32ce4ca5
zaf602c95e16ea52cc43e6e40e0d8373b93de645079fde6c7a3bcfd1c93e3f74be59b788dea4768
zd4763ec0b9b67bade281b1d701b243b97dd9256ba24af7c9df45dd3c72db536f633fc8961acca8
z6c3bb6922c7142897ca9886aba7b819a610207f81d2c20ad0cd29e9839869abadb847555c80459
ze9bb9511ecfe5ef14e1938975ebbf713fb35cfea6d7ca23eddb0b5975ce61c3b475b0b6b76c0fa
z5844154a374a1d24f2e5d7087f6954a72b8c007e81dbb75de340ce53056c4d4d8048c06b09927c
z05a2205d21bded0e99cf5b85af59c012cc8b6aa8bd92b68f174a4e093cda93893638c007d5c94c
zb94c81a4475807432f034dbe7117a2d7c9328c7e15a210fb2ca5a7b00695641c47d370a761bd19
zee045b439b02a582d791b1cdc195971696513e050b5134c063cdfb99657e8017f8bcf47e899d49
zfaa8d15919b77e6658eba2a9ae0fbabf84351b2aa871f56850159301b5a9d4184378b1bd1fa793
z5ded1ffb3f944bd5341ba31eff77c92e479d276def2179a1a2021526700b26769bfbc666d1116e
z4c26d0dfe14257e940a927b1a35abb0141f09daac227382feab423ba64dbc7b3f2032a5b9af091
z4e2deae97b1592bf1e3ced2955ed7d0b90e40416421adb3f98abe738d729f248f1e892448ed4ba
z57a6407cfe7652e477b003fd0842b806c63a9e811e78a8d2341f6b27e08f5b1f6cb4f51b2efa6d
zecdbae835bfd6373c24b5d95f3676026c2faef1843b5933f1a47985b20d11cc653ef7644493118
z2d1c243ababfe5e901254ad7fc7f86c3d5522694bba45078b910a238389c5e6f5c7ce6dac27839
zc70f92f56a2fa6386211a3d954161eb001fa04c4866b4f6da2f4d86501959697174196ed656077
zf3b62edf0680fae95d7c8185fd464c00cc5a122d5d06bb77a9563684261d206835f3734657d520
z29441a0cec370dccde878e459e9163da1877213bb166659795f542e68562591edc9f2cb0da3872
z44b60dd3eb6fdc8c0400b0cd1939af541b176293fd19d271ea351849d664308460c427b8d67e81
zeee656d436b446f861561ec65e9b28cd92ec6d31f42bf46a3dfd848d9ed66425efb177cead3c66
zdf33cd24cff840c3fa6e07fa617aa536a29b8586ea6a52af692e68081d1d23c5f53d582f39fc14
z81774c7760e6c86b155748a3155693cc78cb0c2fc5f26533fb6e85dc33094141da945be38c972a
zd7fe975b272ad06db8dbcbc96cb71e3711bb0db2c2776e656630a7ef5a4d37720c9a3119c29fab
z0c3ecaa24a28ec58a94c9f2e1cec98340802187de6e9634d061d9e038ea590b7f2f261a71ba083
z5bed1105195ccd8aef55048e50374601215a4a5776848959a906fa5a0408551eb9f5543f7fb940
z63e28c77ad54f985e0fa8c5e264673941ec6c7da2147c3143acc0771f95174a472f485fdef6f8f
zeee06bef21c477929db7afbbb48f3ece7c6dca274d2f16037ecae98694e398c1571345d9f22f51
z60c5cb2eb62e5e8182623855060ba435aa5a3438ff286be9072655cd7920d008965af7dfb0f013
zaa8584ad9c012fbadc7470ff1d622d3b77abe93711b1c1d6c2d37bc3e88e1e61f4ef0b5dbbb153
z148c3429a9bae373a7bbf3140d8b42fc71bce7acb430483cb24c1a9e7da156a10036ca1eecaee7
z045b091958efb9d6c3bfcbf6d2ad675dd455992b4ce4f21fb2a49a45a019fbed3ee85246edb44a
zf5d37a07730dcd8f3e1a33c9bf5b230e949d218b92f32d04a57bf66f2b84a9597c787299815204
z92a4e7c07509f93456a46a349a19e5ff6d014af2e0f2e96016f0b47b5941128013d1d7d2d8c187
zbfbd6485d91ca87e6fc51bea6fd70bfacacf3becf6e97a3025e54b28b798fe689cc39dfb808208
za0cfab64f2b5d03b57199bc73afcce529ee6db9fc43b21c498712e4d210f7fbef66c89f56a7952
z8e221063894524c22efaa4040232949366519eabc442f7b2a83cddb4532a9e4c4d84538f998d81
zb44184c9fcc272be01c8c089e33f09c981999596c05f02229b6c9d3a11e8a8c22726658ac5fdce
zd1c35b579ed440fc19ff4908e76a02bce4ea99d156dc1759ef426615eea7e79eae30424cb96858
z68f840c8a59c97a77c54fd4aff90ba68ace1fca8a01eba1d4856589a392da7fb9926cfe6cd4f25
zfdc50d1808f8d9cc6894c738be00d8a837c01dd020f41acd94d90392e5a979e20f849f12be3388
z5efc9a99a03a0f1843ff3912126c1bd78da56e5f6d804befc2d250e9616ef07c902411695ffc29
zc45904d80a4a09efbb2b7e98d3394160eb8f122b0c12a0e95f5c2f8579124cfa71824df2f504d8
z24c0674a317c5f89d4a01287f7cca6e45edef37396c295b3e0f3463fe82d643a8cba4032288c42
z2158cb3163ac6c7101cb95d57ae8e679ce8682b4875892d8494c249e051bbf52dc40d61ada09c6
z1d70d815bd4edcdc39a3a48c545b87abd202b356c456356d93405ed5f7fd654ec261ca699fc4db
zec7e1822051d1309c3d6ec868383f61da6040fb5385209150ae4764f0468df7a4cb544a8a233e3
z8068b9d2ad3f921d370d89d6f8d82e58c12f796b22729e04f83612ba30468c37c96102ad7919ba
z01529567cfd5ef27c59fa7130601e37f04d3812e3cc01a33873b325af349cf6257d31172dd5a00
z94c5d7afd8d780c12e7120909f85c54a9ed9eeadd02e924b6e692b6be90ce886ed6a9a1d1bc5bf
z908167d663b8af7c9a2c0fce6bd1801f48b45c39ae35f6a01947c196c8f7e54ed3954a28ed4d4a
z4917eac172d9f4114b9b8f8618d9bf45da46e692dda74658fd2a0b00b91939ea676810850743d1
z203af1e7386b04c7977c028fd111382a8c2503387e7a7e31dc8e99e7160676841b1b0934875c18
zc7d9d863c89d1e68966224bec8a5b20b462d0fb293a30044f92a5026589e5df95a6b9e55eec09c
z61d82d44f32b673c5246479d02b7290e41b09f1dc008e898e70877f92469aadf41b5bd460e6999
z06b074caaa823b1f9d008c84d6baa2abe282f5cf3e81a270770f8cf982e9c374fe155457845b25
z5764deef017715bdb49b9804c0ca04f1303507c89a2e2d1b57299ee37d886c11a27f15e23caed3
zdf7fe2b7a2fba029702027490a93a59d2facc3d47c952116d75d6610bb507b9ffc999cd238be0d
z0ee5b9a954277f399e29f40ec1a826c349bcd8802ff406ac6f77ddb93a6d638e881080c280c199
zc34c5dbbb814e2f711161bd779dc3f9a12df206b1fcd92029f489e05e941edcdf3800c1b4c8e64
z6f12a9c62afe826b6bb39572bdd823c35abd8e554f2e13bfd17c68d4ac88950d479126b0c1d635
z75721523dbc999608b97ef5845f8adaf078d3fb84121b6422ca8a213d90384980a83b40516b485
zcc0864863a01faab045eed63d9c056a3fed10f0baaf6e8652ecd7e78db0d1f0e5a756d91baf067
z5ab68f8724523b62699340a89fa01a7c6f5e757970140841c659418930e0280bef45cf7492ac6f
zcb7418a2dbd65c77ac26d68daec4d524422c81fc3becf1a98d410f4f2bd6245d040885d6022b0b
z53a24c54b7e9349fa05d140905ed38ede1d98f24e2050a06b9b5b562861a736d607b4ce715e478
ze5372348d69bc6b7091aef034399957c7d1f67c146d01caf83645f73daf4806f0242130222cb54
z49c5bdf053cd07e5cc4d28ec3a14f9644a4580e5f52234db1d56cb82c8fbd8ab366a29ba44d9c9
z1d8016f1cd9f0ee80a5e8a706db7ab1ca308530e1d19fd8f5615b4604f79937e86a1bdc1b35d5a
z1a63f5d503322cbcde02520c27c5bbe3f60df1aec1a61dcac43d9bb2f6053094964972283ae861
za30d823f306df3a199dd6d8793a8d29fcce7b2e12083529d543489be1573c12fcb24103cf99a22
z6ec306a7880446b14d656aba8b53b3c4bd9daf25801527e458cb942395bd4aabe33b58e3cb9a1a
z776e06c64b50f15dcf8a04df5be5f7498c934a465f48e96e76af5201fb23470e1fc07c9b7a9797
z25089eac291d9234a7bb21c4f787a423ce69afa8147343ad4d638fa349bd98097d0336f6134a34
zdbe9a20d2c43d329e114f03bef58ec3da464212c6e789bcd28060da70e8494f64a8d19590e426d
z07424cc3352fde767d925c1aa627b579659e3bda32958c07f81c57dd08e74ec221145a7f23da0f
z2ff9e1e5ce89e2598a6f57b881f719dcbc1ae878e62d85b966fa56503da287c975bd6cd9c1cdc2
z00ba6b9c56ce9e0e7efeb74adfa175c05d6ee4c0cfea30a89201fb93a82c6b533f82f6938a0db2
ze06348d4bcc665e2edede4fcc6a8d8b986db41cdc157de9d357b61208e880d406f54aa8f9d3275
z248b618cca3a0237341bb4817c919d0e6f606918715360dfdf59c823f8dbf46e0f886bb040f02f
z6c8907ba475f7a348589484b1c9a5858a7036b655fa19161ed0383f05c6f8d3868fe60b60d3cfb
z0cb38e1363dd0654eb3eac219a1acebcb2c962f25b5f02f26b161aef9fc6ba31343af28965efef
z40b812bfd8523892fcc6bbe75f20716ba68d23f3f6f3c0f0baa37f77fe0d241eacfcbddec1b963
z067e2592182381f40d62627b440debf684608e9ffe10b4c434cc94ece4ff46b62aeb80d23970d3
ze9292678e059119f5e0ead514c5c25a77e3e866ef45a5cc1b7bdabf342769e0c5e1cb05c995e98
zaf8504b2c5b712749b83f119ba9adcdf17af44eb6ee7ac0fc89075b3d0bb5ff2f43e41937b6c1e
zf9e290f7242eeb394cebb3a7e024e37a6adf79f8e2bf7f6f1bca3814e9f303edcf27c2b60c6d85
z01c8b316d9d1bda3cb651d7cea1d12fdaf03e942d9e52f161c4cee1f3921a116c13ba0997a1eec
zef09563ad35f96422da16c45bd9a49856c461e860120bca9a84cbdacabe5600c0b0963c5b93f98
z2f5f54a22c10930ee3358b3c169976f5044eb24b8deb42a5217f33dc0462217e16e16e17777ba0
z11028a465810c17cae1eebcc42a6804f6ac44fbc056c75e18f3e9426a4f3950dd3a6313b7777c8
zd2cf971795b29cc50723dacf9e6211b06955d6014b279eb24684952dcfe9f72a9123d4c6aa3648
zb02e85c9e8c05aebf0bee197630eae2b4b52d524323737ee91aae21bdab26795edf1151b5b7cab
ze490d8c6756278fdd6fab51e1a79bf8a080813608f9b0f249c5a95647c65aaf80e24ee22a3b942
zf714fd347fd0603741f4cb4f56bc41d92da5b0c76053faff793d73d75874344df62de5dde37776
z3242129adbe8562111c86f52bd533fab8a3f52b21949162a6c4031c719134b14f2ca55f24946a4
zefcc4c6a01ec3503fd893f10fbc61e1ea1b9f69f53b42798903eb9afa5babb7ac144f97a230a0c
z13833e06eccf1501cd8fc3574b7ba79c1c7bfea3a845e2759ee29722c884626cc200ebbef72a3b
z1c206bc4e15e81a0736a4184c1bde28fb8a993d56e2b4de5c8dfccfee370a3889c23459814018f
zeeaee609cdf1ada315659e27af2ca1c37999525c9063363ca63597b631843dfcc48c0330af68b2
z9403b71cb439a6f4b4c93087e256ef216e3eef6b171584dd4f27f3c8a186007b9da6a3c5b146cc
za99332fde7d83466022daa41cf33ede10fc7d4b759e8697f073316352ca175b8a23a8e40643c6c
z132060470eed44b44529f206b3d6a3fb35c2f7b6cd26eb1a90840d94d5fcaf9d2325205b6fb64b
z82354849ffd8dd9f0705c0f41d6df0c22eb30509f9a67b468cf7b13ebc4715778b24b8c956670c
z8075dc664bca8d5ba38cc2698c5ecde4eaed28d7b381f79e5c0c7e4b203b28ed132174ebbcb097
za70c9105c7aa7dc2e71ef45b045c07ca794e35e1ef215e6c29dbb56b19e45027c436d547628542
z09a2871e6560d74e4fa6ceb54012cf0cc0f1e291088eb1e13274d75314f9b29216a95365c10ae7
z7c6183015a41a1063f00230abbea70f5c4e1f24f332f42f812bf04855d484cc7886de14e6e9045
z8cc778d80a38f66a6ab8eff9898eb3ae41853daaa2650a67021e978fde5a1b5a2112fcf0b3e2bf
z178ded1becdee3d52a062cb86ed0db39ab6cc0259d1005cf1447342bec48c8334b7318dffb98e6
z90792915d1c0dfb82efdb07b8c1bdc94a160b68c972e859682d3ce2b9bcd9206746ca1ed40eedc
z561032ed5382144dd57bff0f0ce0b3d4c67d52ccc468f7c0b02744e76df8ef125ae04d9dde53f1
z1088a8c86caf25b94f0b1232d23eb49c4c1faad5c4db1283cf22c757c3e975370757298f1f9339
z7bc702c7c3cf2d6a9573a1789d04f2f200c39205b7885d8df57a2c4171c5d3add5ebf8d1101805
z9aed17ea7e2a91f24a35536e2fbf48a101f30ed0b220e0c9414390d7adfb3413bf40bdfbad662f
zdcdc35b6b452b6da5df3754b1eb0d28b09345f63f12d65eecc7ac8ea4eccd403cbaaca10fa5a50
z2758677368cad7e982c62e946337ae43f431267c4f995a647b0b13ea98238a298ac251b3c9917c
zabd2e19285160af5771419aa037283e938d6185f7711a88a27920fe9fcff0ef5954f666924cd4a
zb547dbd405d197ae2399e2dfbcb7706d4033bb210dfc2250c12ae28188f223a1e5e07f99f1ff37
zf1eefd84e79620a9cb088e184978ea45b8cb2ebd4631d6af797ae1a2eda434d16ba83b20ad8c52
z725d5be4466f261fc18b226416be69898810dff534598226c9333ad6974f068ada2f1b2b90aac2
z5fb7caaa4775efed052b51a7295cde46445a475acf008e186b539e4c5f44397ca6b6e0f37daf2a
zb78cb6502e2a59fd8e5f091049a10e7ae5ff5995ddeab5c325a87fc6df8095577d1306f88ff85b
z2c7d72fe3ad3a59bf2794e3b2640503d7f1b533526b56766893d0b75ad48b59af1b0432b11f515
ze0bb7143cde1beee6986108b5f986b74de7850706d535fa6e9537d3da859434336eb7cbfbd552c
zed13c1b4940c5e4cef671ae72d1c0c5addbfe48d9a0a593a1d0e3a0b9a2d48e68adb883372e671
z27c33dc993c1c06ea972ac81ad0ccab64477bd61146d400827df09e195996158e329e28f277d54
z8355e2a35564bf0508ec9de8cde81701625fa053f2a8b93c6ab63d694b16bf4d9b80c2dbce3d42
z938475f2b02ad4cf55cfe81d639a4fded0fcc45db7591871ee71bd88a1c5378dba37841e76c13b
z1c8813a0683677f318c5db86e37cf01e71f3240c83e29c5948c5edb5594b241eb7b7e0cd931730
zd8aa308c47a809d76f0252d117a190653a10cbf1b4c1156381249f8ff45fce341b9c1214aaecd9
z218baf2fe591ad01d845a8eb58509aa5072616bebca2ef6f1396f09024b3585f73d0e06650c7c4
z18fa94037188f5ac286f553cb7994322772e2e453244051182e090557ce2226b52c419a74eecec
zed5597477130c75c5e0dde57f901387c49416263e895bab9486f77c486dc86bc4c7c2a7afc24ff
z69781b43028cbf7c4f97357e4fee1f8c49fd44aee04ad22b69cb7c51828718a7bf8f4b4c9dff21
z90e5ad7fd992616fafdfa5e646d46003a9d8992eeb6f10ccc19edd3e9ecafc65fa14c3221e86eb
z6b3553dad9d61cc0a2fc028698bd220b3cae0bcf1be10385d595bf4d466b6bc30efebb385d3eac
zb5723db5e31b0b88f716c816540a0d1fad98b295963434bf7f88dd2bb7335be8e1b3b59632174e
z9d46b6f54af236ace5a84db604e483ad2cf652f412de2eb6e929b1d501ab59a3ccc44c0f1463d0
z800f769d112ac5ef4f849d45bfd155a3fd82e20cc6c1b8160b08427dd88cf98bf8d42fdd031f31
z628ed70c123987ec7b760c4baf5edc347afe7b49cef82333789abc0099e6f67788b68f41de299e
z8b3ad907e9bab41e1f904784e574e4ecce6c4a4c7c64ad0680eb80df7ee332281bcfe0e75cfb3c
z32a658a73b74a489059c504190bc2ad02a5b66497882856a94eec4cf2484324a130b629d2d775f
zd89d45ff534642acda16b723625c432089a046c2251ad7adf96728c146897366087662261a6989
z785b8ba0d5136b687ff1465afbc4eeab8841d427579e4983535dc9814b5b33dae9993da4b20d70
z541711a2387d2f4387348fdaf00b76eaca1b9c878c6132611f458c1e4c314ebb18f1755c777d09
z37de0420abec12a5b68762374096a8b68331310df18288ebe7d25c7542f3d861d1a6017210187d
z84866d342071564fbc982342b3d31360125dae02cb258bc1f9ae44ff9759bf78d1b885811b7ddf
zf98b6d92d380ed32a0c282abee4d33bc4e765f400b16ee3c1b0b7169bb73825e54b432862ebcbe
zd7cc0e7329952edcaac6bc3616cbcecaa3f0bf0416e1742cc322ee6abef985931546190278031d
zcb6a5186075370776c3875266cf2ad92959fdffac31429990df1d0e664e614e4fa8331726f351f
zbf7b5e63095088cc89b500a5242922f169c00fb7f98cf7deba96bbfeed95b208e91c9a745c30fb
z24984599ae8f76c658a14988f883c80afb8e683bdf9ae9fe511e52b8ef2ad0f1f70a818f245c93
zb449aad268d4ae9093b5d5efd4411225ee567df193694170182e383ce8396b8268b01d6ae7fa39
z34347821947d955763997bd813485ef09e7428ed515948d6ae93290283ccc818a5724836d24c19
z23cc0e29a3f83f4223c8ce24e52659dcdcb6b9f4f467cdd1f50d0bb501fdf76bf3138a61954b48
zf6058f3d9f1beacf1ca0770c86b37a182fa022078cdff5da4e3291dbbe4ca7e7f0fa4789fd93e5
ze771269b2e8aca8a1861c010423ed67f3b11057867bb4f04fe179e9eb2596e97680c5519aff189
z0dada28396a3db5e77d18235424dcfde7bb955164aab76bb3f772a251560f5d1b372d9cffd885f
z5b725b4711c1a4087c937ece6c74ffe857398337503b9bd9ee960ddb493ad3ec1b102bd5b80089
z52c5b57467f6cdcba8daf57c717c3da6502fdd70634025b2061a1f83b0f79ee3a993c80bce3c66
z5b4da794c9a71fc41c14e7fc4f8bd98ddc8b7a8046835b742a8e9eff1b2e2ede31dbffb7dc9d8d
zae6dff38d53dec0cd95090c2671c6b44563f7dba705800b457d49f3327b4311517f05c006d29d6
z99bbd4c3f13a2f7021a064c8fb2a1571a5ae6025b6e85fe259911ce3ec4fb2f8859d44b53adf81
z4ee238771d4d8703ed4b0ffc3a6375e15c4446ae8d4b2238d94265baf8b924ba2a2ca5ddf20bd4
z4cd46d54ae61fdfa95f4f1dfd636a0a495f8af477f48de9f799ab8e5be1fcb34a86c7a1aaa772b
zafc92bc14913ec5668d20be08771d42b966f4da821e9e91dc5089d17a093ae41fb89ac165948cd
zdf69db3baff311c9e4eca1dbb95e56dbdd4d8f06b010912518e405c73db516269a2c4881fb7416
ze6124458af75c52da524f262a15a170d21590aee81300adc0d28e09f3c70f9648c454cc1d3bbb8
zd23e20b6c890a8427c24f1f20b37c7ee9871a25969b23358e9f69b79d996ce5decfb216ec78f26
z1c8f3fd18dac91fb3efa5059310ca43db7e3fc42cb9aeaaaede7ba8146a7d5bf32f4bc1303a9fb
z69f2b0dc37c0a1e11bbc7c2e78fed96daf7c5dc627532e66ae84022fe2df18a53dc92e62216718
ze53c6a6d31963520d131b4580ee61ee47807795d294434d2636293748b2a2db2e658fa52f64ed3
zea619128bd550e58e49a4547a2fc4df575e5abae65eba4796b73c1a8ac94b1513ca760fdbfbebf
zec38331c3ab1b74183157122ad478bd2ab2a3be52a781c1e01ffa3f67ae040d59b9c3c21b0a928
ze423b2bb7667eccc471eb1ac068d461238eb0fa64386f9bb38e4fc8fae2c3cfce73053cda4c19f
zc1ffacab782cbb2de9e922c76f25c3af21f00f449fb011528fe9d49d5b2141a71fd7a04acf5f00
zf959c9d17cf4cc354624dd10038f5edd13ca47873490492ae7a5bc395e435236e8f63079ecb4bd
zad71fb695bfc9daae0169c8a5cadc233884f6808712e94d83bee6fc6de4552e2be5d329b92227a
z4bb4b07c2497d1553f48983412a5e81356e340f3e9df68740fc8680ab5added1c4ba0e543842f6
z2b34bff65b1eb8f15274b0f71fefe3aaca597d9a0d29ab38fe50457b7d6011973c4a0a3291f7d5
z88838b29864029988450998fc81ad96c3c06250fa6c06911ab821c8e47078460b9cd2d2ec1cbe0
z82f04dfe6326bc9bacaf038467c720a236066e34e7270a7c9958b13046ee49df652bd2bd60e381
z8feae340634d8f81ba152b41dd8f89e3e38647f89334ce2b3b74bff609fa3267dfe55fe89b08dc
z5a9d66a08205ca81b3c7a86885515c95210814568487251972bee8d2aeb1d59f95a7f99b5e07e8
z886ddab80ae4a0bace58ef3997726e2697b38dbea13892a8da624e9d15afccf8efe9698c0116df
zf8c10da5dc44ec62c09847c875af5957ef0967af4f21c6f1966c7037d4d1d6e929de2fb9c93e90
z32a15093b587eeb517c8eaa8970583419d37148486c95fc189a188b552b837406d241fdab55125
zff9f520899510acd01fead8e8d37d4e9f245e31679bf2b2505d5a8bf49b843ad6f382970c650a6
z690440f8aba79dfbb1f2bc6fa9ee19bfb13c080585d640c9705afbe073665c46f422fa2c866125
z3b9349c8557b21b7c8633f24b56504de3f9b632b09b4e599341f4e60dd95de2bfec7d043e501f3
zb712786198109e6faf7612c1595e9fb2a69d46b28055ce02c6f4f21d433bd03a679c091a585633
ze180648b60fe9db1e8cba61a1a713ef08fdc337d7248a2f690221e8b67ec94785d5e2b44ba1f0a
z4ac44b165ae3a5efb2cee6f5656bdc2f389520c4b19f04693bf20b980d43f679f36836886b5904
z560edf3fdfa478a4b46c6785c4f9b3774d35df6ce75dca165e536701803512967c0bdd1c625eb1
zff3c4cb0012a38c34281c425afbaf8693406591a843a405e19b28d219b374ab8ee3946bd5ecd84
z449444c840fdea3330ddfd8b10556def956ff618f6509bcb81e2aa85134b103618fbf573d206da
zdde191ab6c2a9d4bedb2e6e002725705400d51bd1c733810eff7ecb75c32dabbd60323d9e7d28b
z37862b97867cc3aa0e2f450142ed62c3ebf9b47c5428bd6796a54c905ab073adbd61aad7716a11
zb7e69fe91eebd9e8838180d764c3d69241aac7e9e9db7cf5ce485a7e728117fc5ff54caa45fc4a
z8d3745f52beb84f118b38a5ecf25e6a8950551f8422f88ce0f16f9c32da005db9f6f1b90951917
z2ca7624e2f7a8dd94439778d41aa36f8435ec64103ce1afac21adb3544eb451d3da536e2cfc281
z1f6bb53fd3d1d799e73db93da8049c70064af04f6b7c99509c707ffda3166d34a4ada57e5dce08
zcd8c19b129314bdc09880adf5eafd13a2833eb2ca6f127a863ab44ab1692dfca3ec1671d488334
z756fdbbb93d09f42726bd56e996a9a44a63bca2f6c323168fa8c49ce10dc59cc409231a6080054
z2e8cf2e45d703c042e43e066d6099acb79228913ee99e89bf07c1a8af2bc94837d173fad309c59
z5c3c49315388950f56b9bd383f0089cd1e3c9d4cd73d4a1b2ebece292bddc936fdd31288334b90
z1df8696f03b3b5e3897671856fbd9dd4e02f3340cdfa2ebd23be02dc0879f5c5ff0a54e5ccfdbe
z5a6c42efe00105374e098df87cc94e99ec899a236b3302ec73f075fb14e65bc3412b8c1f5e3915
z6d663c42ff3fa5673e956acc7b5455d1eb774938cdb74e3cecb50db7df598856d25ed7197bf80c
z86aa191549bd4a7ffced6b79f71bba2287ea4c035f3dca1d0ca62f02b191b3ec01291c939d1a0c
z6b685ebe3cbb0abc7d003762f0504f16b8bcdb0021128e40dc94b7ce4ef0851882bdf39340e214
z2999e37e0a8f8b2881d0b43781c92a459ef850488ab895678e0c18f62f5c7a1126323b9ae2809b
z44f89da8f5bfcfe116d9c76d67d823420b5948059e472385586614fb498455abc53eaefdd76c14
za4d8183cfb72ac7c82920202a031cc4a269b95423e91d10e864dce596e17e0bf314566d61b0d3e
z3f900b4670bf7d9a42cd3930de21d9174bc287fe20584ddc09f2dfee0cb234c641d8abec23883e
z78ec232fb64896f22ac0a2f196597082edde9c6fc0166c31b60e93c40418c07a6cedb0d128d5c4
zde235185de48a5645250a9ce5e1fac5f655253ffcb03b0fd9c67d907403b0c8c274ca62d1c6d28
zc722c1e0f0aac517f294b55ac2fc15c4724f0c295d6c29906b2b865f3ce9eab635748baa76fb4e
z4af1d9743a9786ea3abfba45b9552e501e630befb8b7b2cfc43404fbfebce700a51a1d88478cd7
z0d8f013cec9409fb34cac895cbdfaca2f4b01900090aaa1566e1d48e8ff8185e5643bf42faf6d1
z3a6e3def7128101f95693160363863ffcc87b671f157d2074b11c69f540cd2af005d400a67f772
z32b4733336fca92ea17696b8bc70191ff376f006a833c7a7e4a637d92102a602d97dbd811440d3
zc3580a06232900176154d16ea2719415730dd13b8905cb9dc7ec10918df72012de4fbc62d83c7f
za5d5945ce85fba455baa26b2af8a44e22d6c07d78f26d3468685aa92b3ac3b234efc1da7285037
ze94fcff06ae8243b7a43afe211ca2c3f1d17a52e3ac7f62edb66868f607d649a517e5d067f791d
z949b647285abdbe5d48d6c4c8315ca2ad808d70f56da7e9e5354e17268d0a2c2b4dce6c234fa6f
zf87fffeabd7c8b60a760a0ad87806046116429631e29b5b532a6df4e71164583881d0f10fa342f
z16abe91a12d8e91a81236136c21bb3fffc51455a2dc1853e559812f32073631aa2664271f708b6
ze8dc35095104cf9f365357c0550431ed06322939a770869c7378be158db9c9e463523c67baeb46
z49cd79b41f86c23cabf3257d0767c8ab67e4f839461955242211768712c948a5de86b79625ed04
zbc80070fca86c75e07dd151e518f1283974dc3ad303ec4394b7da99a106cdf2658bd99b7a9ab28
z3c863d69c6989dcb8719e76091cc5ed831ee5e657d92a9fe6307f70f5d677b79d29fc7c3341765
z3bc87438a58cc1346e3d499bdd6314cc94a60671a4812d6a078527e30e9c93e61240d3676710fd
z63babd83a084b7de1fae5fb2d689f9c36605f97d29bc0fcce9789109efbb0a32d6e1f82abbb7f7
z1f79d0a84e6a99580eb901119ab321b0690e1576d63c8e47300eb1329ec9e67e6cef7e9c7cf04d
z8823644a746e44f24465979420edefd11ab48e0eee9172e34d49430f34933a20c1a528216c2575
z1497b91c21887e104cd97faecd2ce5c646cbdeeac16658cbafc7a811806838ded843c21ed867c6
z10d793344f402aeb55cb580d42f5aa7f2163ba38ac53e68948f324a8adbb9fc90128c29b142403
z9f046005c78ffa720cfc40a5295f2f4269f4439ce789e7254e5c25598abc58e6884d0d488467f3
zc13079ab4ea890127be345f18511b884da14b73f1bc2896f6c6962af34d00cd8b4a13310f30be9
z62663abd2629502a03371ee44e05fe4d2b1e106b95af862013b755a36ed9cf65c2b1c5ba3b320f
z8bcc96c2251a10c2fab86a942aafe9e9efaa9a918055e4572886e72175cb8abebc162c285d3884
zf283566a608e1de32e1b34eafcd030697ff09ed83d3026587dae9c21b8cbd1cc1a35f0cca36d3f
z7a3aac8ed01a05a608a3dc2304a2df09157f575b35337e4fd6deb2a119b25b36a1bd702cb3030b
zcd523120821a801801f5f9dddeedd536d970130a87908f10f7d98ebff7bf648d23f7bd1d1ce216
zbfb41a185cf746fbbcd36cf378ba046112c486c315f4f15f47290c5b56cfa47c8e6f4565e9aae2
zea40570d1da120149d161e7aff3bc626df37d808046e7f88b230a0636a0a5c9fb167e1c03ad01b
z6d04df75d8e5600806c87ba7694edc9c6e011f9bd233134d85ed8b5adbdb211319b13d9e8c846d
z3dc42abdc2560439f98f83a2f433d8dd3de93170d80099085e85f8ee9f607a8aec0c01bd1f10e8
za3b509415b919afb7439acfd8ca5cbb28003c85f1f2959de9b0e3db1dd0ab927426b9b0b1bdca1
ze577b61480fbd9137cfcbc74ce874dfddbc7f08c962a07f391f7973c2aef05b03eaf5b7c30331e
z38e48ed75238d63b16c92166cdeacb8bdc0e05ccffa9831ea763e8531812971d3c3fe403b76b29
zfeb31dd6056672a50f9ae39438ea38cc976968da92b3007a63cc476d70ec1683113bfd166ce07c
z14e0e9ab2e54e72f8827a0f43ec3b7b1b951d1d7553b0b6cdee3629ec45e0f4770db8cb6ed67e0
z16ccd3785c8a21d674379e4818e34f248dfb87e7163c389efb56865557c9ede1a951c7d1ab7373
zc7466e5a941cacda834d1fbbcf41c987568e4eea96b9ba0803efcfb7484f82be23c36c25a2ce52
z6f8117c39f85c5ea012f95f2007634de9ade9177b104671de1b08b163f43b1138d3769f3d7192d
zcd191748c024a11f85ec3b75d866e2f14d9dd5ffac17b3203af35381450745a704090eaa948c1e
zb6d5a0c466d5b874a3e47664052debec97467e4f56cbb5cef0f81b97be91dea7b9bb951fcf97a5
z4a5f1c8b5eea374c64e0da18cad5c4071b54fb01db099a34902d5595e6b7a6e6f9913bf3fb5b01
z518b5b4d125d0c51e626ab229f48d126feda8099e411044cd024b78215ded74c51d53cd34aff09
z997c538e0a62f881cf949f20dee4d3a725cfd695ac5e8c694dcefbd83cc897de05868df98fc244
z0492dcb508a5eff406ceab0bda353017a9a82c96cf30ebe3d3261c4945df1387b437dfcd134eb9
zaf997381cc20dfbccdd6d328ea28d6e9ac9d3e0d979dcb1350a5a501e4832acdb1a0371bef18fa
z24debf3c07a2c6a2831f49ee749d666a72aa209def300b767b53fbd56401f1aac4d4caa3b6732d
z30ada376ba1f267ceae3302caa528d65631d367f0ce3c542d91957fc255d92742551eea267d4c6
z3fafdc78ce4ec6de7bdf7b9e55ee9b2a7ba500076b732b285316940030f10d497613326f28a936
za6c7be02c08a1e23f2f3e26cf37ca872585eb213c0a5423a1938b9d4985b4e20dcaa79595b91b7
z27b5c4122e820cc08147e70edf660f6fec0935a9c780d4571f865badd749703d8c1016154d9310
zff2bb57126370097c79a1422f574fc5d46bab61f7c1cee00d6372e80f6c5ac740691ac58bbc08d
z6bba0fbcb8a1bbd0cce487c62f6a2a6900717056774b777f8255735988fed1b097b41799ece937
z136607bc2f6138713fb8c8f47c8cbbc8f2fe18d0d5d49d14712caff6775cd75010387d5b29834b
zeeab1c688ba38afa86d097b5cd7c89cf90c957eac46eec7b30a6c80fcfe509d7c03810cd17eab9
z8bffd35434ae9c6aad814d4cca62b771be177bb04a24e54ac4cdf78ad9e45f2b7e611dd77ef559
z400b290b57c7510578a6316ed44fed4ca790e1e8ac84027710c7febfaac864f8c1281c959d6916
z8a69bff6b40880afb3f75e78a16fee29421fa253adb678e9fbe345cea31d320eebfdb7f2010a8e
zcb2164d8b685510823834f2850ad868b176eedc29a652658d5e4edca11c5b0654e5e0b27996e53
z3fef0739e61ac675aab6bc4da2029e81aa7e57eec5b1219b033bd406e970524a75612b16349a75
zde5dde758483d43a5fb4a62e6bb34db16ddaad7928d9b5fe599ee1fe07125214f0fdf91b3ef37e
z50f15920a288100f63e2c2c3ba0850486ad1e3fef0702b05bd279b24685baeb86cfacf1a1d5755
zb49753810dd1f38c3915de81aaa88ab54076f0963c6e6e85f21c8035bbd0f64b3b249676d1de6c
z0aa1870aa85685898eaea36a8e104f255fe608f74f6983bc3835f80d8718cd71f7b16241001f10
z5905b5cdcd9d4fedbbf5d9231d0428f5b01bd56f9124ccaae6a5109ea30882c82ef261790edca8
z79678e15cb82bfda24f7b597ada545f671a04bf2d030672622012d4161095c7ad9d6db88029ebd
z71c1f8a93ffec0347dec03151f23127dfaf20c40e5cd36daa3e23d7556b376ea8ea4fe49968fb4
z7702f99826e5e430d2406c8fb5726eac3d540a0602c4c3b885477157553f1fb5c111f0cdc16f35
z4930bfe75b080868bcc85baa129e687426723d04da81381e78618ca130b373b50e8550ccf247a9
zb1c261e8efc237ea31157e23ac2abc5eb76f0e2b66558e586d8e91238bef78ab13c5cfbfc9f819
z9c0e95b65ae90690c918a0481cc62b7e5e0a7e0a3afd159e2f6d01a54a234cfbf12b0c6500ceaf
zc49db6900842a2a939b6ac2e484a5cd7c4410ef3c26e1a75ae732ea97c0eaec065f09b587988a9
z4a44c78b8158d4240f100872b6c7477a0cb4b491ecaca92463c0a47a154f33e1f47edff5c796ac
zef6f4a3b54748cc61d8bbfdd3ea97194b152b72dfa9aef9a39b6ca952854d441aa71457eccc0ab
z3a8f31e141e9c7aecc8db55c7b25bb7ad03fed30425d54e3ed8ac0c3b63a006fcb3144255a05cb
zadaa4487a649e045f1440716ea59a01d7b420292c10d9e69b8bfd90cf0b4e9128e0e3d264ee662
zcf6aeb2b967be237d6d28201f1edf70b2608c504fe296d27f6dce0fc5cbb2ae58d6ff46ab54bbe
z0dd9fabae450e228ad5b64c152849f944317c0357aa5bc3320a6a26ed16402b0bf6e5d56a3a647
zb0d0c4033922007cb7395a67ed0fcdd28736cdd6195e1cc9e5b0d83e6bda4631c377b3edb10a09
z19ff25953a596d4dfd853a64b7bee0f45bbb82656cecb3b0688cf114978120c344ab54e683824b
z4a2bf72d25826993a4f43a825dc7f6cf78372c88ce4060ea452389301ea4b8af6071f65178e752
z0cb472f99bc84b76ca0c28019b1a158c72cdd1fa109ac271faf2233cd2a1ed43a6b7f5bc14aa86
z382a58320d3c19618ee260060ca0867faebc2feb75f9ab36a784e0590ecf68dd357968d4436b34
zff0eecca290e3e1f726cc3493724888cafbe64181ebf57f02aec91f5732f6a9987a6547b6d708a
z42030f7c34414b41b26577832cd784e7511036787f86f47b359bc316ddb915e78350aa5288311e
zc796d9fb9b46949bad30c54a79dd0fe10dfcab17ad7e769805f4396e4b5c3efcdee08a9a3964c8
z80eba6a37218af7f2abdbcab3619b428586d7bedb09a1d70dda074ff552411b319db9e45090e8f
zc4d6080fe5247dc63d98bef0ffa71f017088179cc49b4eb4617a61cd792cfabbf921a984c5432b
zf6bdd2e6cbfc439dbe1bfae5920c5a47dd6189e0a326a99517cfafd1aedbc6dbf9a52c420cee22
z3958836d32642cdcae0d667921d33fa3f018639d6b9548a2b8dfb6a6f7fe8f90d817bd162ff7e7
ze66525e769e0cf912d239194250ad78b2d97837b205616a750efe222a695580c418fe3fb086c58
z44c5d328af2c88637f851616767298eb6c64c2d7356db9ad8cc362996ae47b65535d061619efae
zbcab8a3267f2bda06bceac8301c00ba8896c5c6a1aa3e288b76ee510c2e79710c99ad4db3ecc7d
z95babeacc3d811b1641fce8c9d8c4467aec1b16d523a83dbd85208ccdbe1907b15809aeebbc6d6
za6a6a2411857aef835430d16aa6aa5c0172cc2c2ff1f773acecd6a0a9a2d10c19fa92aeee1dfe7
z53c27049b5f9ce5150ad4f434b9cd1e5bcd8274afd9a1a1140daa35c375cd599f0c80f195f356a
zbd4f923533043dd342b7d9503ec55ed69839c61c76a97a002a34267c7d1da7ed6d80473789ba9b
z6d736168a6cc40dc1d73281f2cee666e0815286f12489e3ec2e4484dee52d117d4d50abe6927a2
za72c05168958bb001fd0bd9c31137585fdc59b82bf74e88b21f875ddfe77c879f51b445d488f6e
zc029fc27d6338a0c7ff44f3a4491d034f38d12390360b11b85344e5b7759ae2970a8659e3aa75b
ze1edae4360136ba51e2cb1ce650e740fe037a4c702112135ffdcd873ab4fb6dcda67f8997a0177
zda545d5fe24bb00f0a5a70d0af71294d60d109df27f43c180f5534a09e8497454ee22f1829da10
z3c0b40c583bdbc937eb43ad4e08ab42de2670c38502d9a7f155e20aacb539817bdedd885a1e789
z92aa5940f8eea374675b83d726df5b264548a45ec46d0b9289ca75af8886683314ef9854d317b1
zb9cbae6b9f8d1fc9c1731148e5b0ae6794fdb37c264eb469d33981b50ac609ab34882412d8ff16
zc5073bbf68f531157d72060450bc7e1d47a212ae384e646fd9b8faddf7dcdb7166b281efabe0be
z4a8a7e5e974908b9f508efeacd2274c5a1d920f9c9a88d2b9d60a13f3258f7f2c1959e9bc6077d
zdf869dd03e6237418045f1f0ae1c725d6a93f6755b514d5c94cd926c7e8e52e4c9d4b84ee7d4b3
za06ad1bd30672e41ce2b68f6131c8e6cdaacde3e4883e31ce97b5d874143cb266482ba4df81cd4
zfc1f6d75be94d17422f5da0682dd763ebc9dda050251bc7bccdb0d300d6c437ed495561d2d4224
z4aa3b732784efa6a8c9a8c11ccb9048a7397aa00f2df8c35721f608d960a280b2d2bb10db55df8
zaee5d45f897a5608d90b8f1ab25b3c8350cfe224823ed1d440b93cbe96521d0352f75db6383cb7
z18e0d3f7700d344c9d0fcc9f14343ac63a407024fcf596407e6f5b0df78a75796a1761fd1d0996
z95de474fbced39b02d16258ccb84c09c28f4463a8bdd732d2f640a7e033ce52cc16c648b130be5
zab7aba39f98d002fc087b1d8e558a0d7e0e570aefcaee59569ad14cf31deed56ade76b75339936
z1743a047718093b8a96269ba96bf246a52ea7de23afa674ad7559835b1f2a34018fe5ec274690a
z05258b5436c729e0155998cd78f25e7caad4fda8190329e874c42586070830008cbc53e16d4945
z4743e36d60b3cef4224c40212e275a1ea1135e1438fff5e10d4af455513b24368da08adcde5083
zf730217c28785e325226b27e1699f48f3704fe6a5d461134689c2fa5fe4111c6b39ca5894b5a4c
zc3b84820a696f782d5f44655b2fa9b385c2be7ecf1940f4dccd243f462e7d94ae55531865c5a50
za553b1cec75be79c59403488ca633f154a6a1951e41d4f15cc22ea1529bcce21e5ed86f3ee9429
z466ad2fbf75ab0826cc97623101386800ab348fee21b923c8736a7915db43cd97917992f6132c2
z690b18bd139f8292ff16473ff055bfc2ca159dc0e663c66c8bbbcf12d2af8105f4bb696da45a47
zfc18233eeb104328f864687c79e3c3c6dcf6a790ff92915933ed4d2028bcda61f53edfe24e72ce
z046a5bdba72a5f48096ebe01f8e0c3ca115e07f4064c0d28bb50ddec7ea52a87b25d2d8a1d4ac8
z8e22e2e8f52eec459231ca5e0d5529e6b562ecc4d4daf8a1a368c6b182680d7e6ad85f70f5b35b
z35106347c99dbcd4231870cdf0a3eff24c28080a3f96e1efa933346029c383ff23a2e3ece3036b
z0e794b8348164f3ebc817ec2c294fcf98e5131b6f5d6ddee909236e540024b546c028e4eedd3ba
zc9b636b52e7fff625d2ee76d6094aac280e52289cfcbb727ef3fe75e6c0d60261b526353c07011
z58c8b569e3cfabdbd8807f31e8502e5eb65bccb8dab1274129b333d06fcaa558ecff75caa77b94
z4fb7e4dcb7e3650a6736fcb4e026cd598e7d48690ae21c333b168751982022b6157bddf2b48811
z3908b1b709fd7d8bb9917a96a791490450524b77d72c59095b70dffb423565906cb2b199d07903
z00fb859b1c8cb212b494f2d6f3da5c9bc8012da71430bbadac65824df99010abed3bf8dd28b553
zb5143f837386e2ea32e78c2245a6d0c12392c69312e2029dec5a42b419d06cafb734b82f26b0f7
z89d791147cbc5f50a51b8fc379d29d5ef963c08e2fc40da571175a083046037e955954d6971e82
zd776567b8a29751610a7592ae49abb11cd36afc9009cdb94e25ac5da210752a8dd7bc42d81be93
za102fec7eac6ac9c200c65798e029639f5f4668f852638e9be01b4a9a73d0617b1b2aae68fb691
za6a51320e181b3f5696ccf85d5eb288db53de0733ad3aaa4dea0232254980e80b15a78c700beaa
z7419395967c2415fc2020b49cc3ea6ac29ce103c2b19d125eb906ed200578e0d5e0dbee5dda531
zac2fea7d49335144ee03d6aa01b14bade416f8af52c30a4916ffab7d9f340931eaec7c369fb366
z8dde9630872db6a421b92170756094adcf53ffdb8da5c67dae2d58ffd8d2362ff25945ff611c02
ze2f21edbbce42f5d913141364a83023daf2c8ad7b52fbafc0663c3c6069b6a075feb87ba4e506a
zfea9f9a7389b309d2ae475192985faa43a7828d42b200be9da02c58bb1c25f68f8a2afa552b2b1
z9f4fbd50b07d253e638efcb1123322068e362fa50608c7f0abfbfd30222c2a38405c78ad8f46b0
zc6f7a6275f77d5f2c716187711fa1986fe73611d118e4f13de4805ae2873d0f4eaf1cee10bd97a
z569622ee1b3798e50c008640b4f58c9890c307ff9154c5d8b949110294563f76022cdec3cb72c6
za04318befc3007e67b0693ab5b197f0dfbcae7f32b972b7de6ea3a600f68caa0051e27f03b5796
zd021d1448cb02091c68d679fe7f26b34d13704d121b25db9707c3d2e2bf403ba440fdb826d2a01
zefc09d9d0506667a91893e93ba684212f0b38510c0a43915d9c2e7227f9d64604f96b76a334cd9
zef7ed87beac4bd36aadead108120d7dc25868f2f14430a57fe3790978d02e3f909b37f594b95f7
z46a12ca60b3f9da6cdaff211b477cfa28014465c9ccf7faebb9a4443110366073ad4b63b91293b
z3a8c34839960c06883815f1b5f95d6282814e4ac418b1d10116000de910104bb725cd020ed77e8
zc610da6659e31c80ace474fd0c9d777773fea8b49b679c25e11600dccf7a9a29dc00b4135abec8
z38d8f92665c5f595d87f2802f660184986d81d4e466e6b9b6ea69c78a4b6146ef3bf426bbac0e6
z3efce843591dfcde3e8df46a24e84f640465d7e7cb94d1925b3d9d83edb79487f1c8258baadf36
zf48ad5148be5b3e7f48c13401c671c211598f77e80669967d0c6a1fdb20aa8ec561b31849b69be
z26e51cf41e077b488183b1597b67564493dca32e960d19712b6f19031aa4ec05e518d9eeca78c8
z81ec2169f7077f785be2bc1504c27f857a34fe9f820edabf3b8d9478b7ebf8e195caf8ab9cb9a1
z1428c04d33f51e60815256605f7591bc3249a30c23c9fd8a0dadac61dd027ef78de9258a8dbc27
z8063c8857bf75f7e104caee3bdd67c738846c2527f4f5e4c2a9fdda7beea326ad9acf3c1fbe599
z04a6985546a9cadeb8003ea52d3f3dd41835f499b0f24b0a17c81e97911bc58ea7309023447f0b
za3ae8f03cf5f7d55535f2dc6b92c35221bc07c9127d8f744531d46951507ab0fd234c2216baf5c
z85c04bc32b7cf44423d0a6f921bcb18be531c86bb64390cb798c965f25dde59578f124176a2416
z4d94d6e304c9c824d65acca2b773fa2558e9b45b4975bd270828a9eef7a2a3d85ce6df4d7b7f0c
z5d1a6a2383dd614c3b4c1a012ab4034df978ad38d526c181b50e11365fc61582caf883dd4cfbc3
z290e16c460d8309825079a36ed7f4c59e0fcaf962b10581e36195e05593058ac1e51961025f188
z85cc811acefbe423f630aeb506663dfb737775cd8e2eb49760f3a3ce67077aef34d718ad16d943
z71257561d14fa11ec85ba20cdb9cfe975d82567140905fead9352ed4df1eac23daad36afac2d83
z5c7af53f6c9d30b75fd0fd74e6b86ecb10190cd258af131fb2f31e4b944e24706c23e5a9b921a9
z40756c2d801a41e5d13aefa309af85a9776201a7430f01d1f61c297cbf34393e324ecbd50926b8
z2ce6a06a6e3101587d65f0a63dabad5c74d2cccae88a56778485d81d6e087278d0ae14cf426853
ze0f03c9e412621213483c71a9500e0e538912c62547ee2688dfabee5c1abe7c0c9c1dd599e7774
z0c1f60ccd8d17b02885e45ca9517c8a18b7d17c6342e7eeac41b947bee45b68e1a3f57f7b36420
zb091c888d4c74869874cad64183b5d9ef7a48699f3ccc188fc3c8e973430ffb98f4cc832accb35
zd73be95def6b9a45806d836d2b6f5a031994f69a71bdd0c568ed74dd1dbfd497eea2626e8fb490
z364e9e20b1db63f5fffbcc033fb2ac897969f483887908adedff42046d553ebfd874a27bc192da
z392158072445115ea677fb2c0fb9b64b51ac0aeea3caedb8f77e99d4aa04096a8e8eb3cd5c9206
z5b9ea3509244e3080be6f3e592306fc2680b5ac54285f1e66af8a8deacfdc00960a7ce9b48f00b
z64d689aac03e60f5af715926ef9fe564eec8d3cc66bb6f44eba33c3e70ef08bd7c689fd0711cd9
z1ff31c47dd1b42fe0cecc6e86b666fae9af74fcbde201ddcc26ae242d39c29ef65f5e6542ad471
zfb7dc959f1d85c55340e6cfe76c43d3ec80e628572637437413dd510c30081ee82c2d5f7c0d479
za46b97fd00192e7758eb607926a3f1cc82f5a773864e0c7646a0bc7ec338ff5d6033078c5fb85c
zda6945c01daba2cf989f6e61633756a7a6142d8d5cd14ade41e2e293abb87266a74eb19dbdf604
z57c1314be920f0f58c5771e2330f1efcec76d54e9fd1a505f1cf3a99260fc25daf964690b6ae9a
z3e2728fe35ed1823bb27e49f5f3747ff05bb8c38fbe4c8fcc3562614d0fd6909df86fac168d437
z0ac282e24f8db0a5a6ab1c3d3277f3057cf0404a41b76af59a4ba362fc9d3a3bfaf3a8e9d0cdc9
z35107a4c914a86fafa21c395b3c95e431b5c6aa4fefdb10b36594624fb44737a509bb25f0b7a6c
z94c509c05ba227e93427c3975ae8c5d36d85ff6376a87974b9742d2619c652adb68bec16d88644
za26805783dee88fea49079de391b4c2e1bee409aa4d5c24a393ca9c2122e94d3d1ce2ff28dd2e5
z2c505cedac8ed039d3221c99f7bbb3a83ec506002a2eee673aa891f44f515cb45f55ae7fba0d60
z88b13f66067d28f2f4fbfb2bb6ba1e7e64307e6f7eace97c8bddb45f5d8ff461d2a271bc818d8d
zb22020e13461773641f95c32e7108dd8cbc23a7bb3d8dafc6fb100256140116e27bab17fb1d269
zb3eeed4f77dcbd34a8885b3189c7cec8c77ae02b508886a73c6bf9634c1663eaaef3752225758b
zcd56700b59547ed5abfd61acba19e74bcf6f22ef51fd637cf2543a487d76ad79c05b8fc42c75fe
z8ed4d74615e190a82c2eb5d53ba7aa9c5cfff1c545c4b852abcd119b655f9b98ff2ca95093cb8a
z9ef509a25f78ab95e8ce91b3d60ff965e799d043452979c950f4003e571d3afb6026dee0fff907
za5557e3690142f80e25de0d3255f2c7100173e4bd976dbf297208301133a4cba880fa294b492ba
zd4c79d8dbbad811cc5d46d1a3491739811c72a7d3edea4878c4cdf6255b62ff53e0ac02da5bd27
z25d63e98a79ec0935028a86e91375d5a2d11e52b568678a6d2136e883ca80829e32ad4b3bd6449
z2034384bb5406b880c83e73743848f05a7a86f216a7a0d1c9c4d568ca51f2f3df574da82b26105
zfd90e7e5972d2968b647694eb1c13173f2432ce7a353ab995a75900d244ad7fa9e8065cc9fd076
zfa06248fb3d4abc916a480f0b611bce5e332797430d64bbcd7a3b4255b964b1a3845f9bacaf9dd
zc7cdc44479f01bdf181de6c4974d4ae75a0259af0d05dd880dfc4c7a07011ad4468ffd27186528
ze0e79bd32e1c0a82e9bd5b2fa1d46ac2746329b6eb31909daf21d367909cb7c3024298198f702a
zc2ae96011cf4918069fe631a1a7a246457f2ca452351753e0ace6fcb0033b11cff6354caf14917
ze2825bfe81a282052328a0911b2ed6e70f91d2a6f3b4c8314e8c891c607e8145378d9cc39647aa
ze50183a31d61834179e2d00904c23c4b5c479228ac5e1c12a1c1109ebb9ec4abba75f6587d4543
za75c9e47ab59147993762967316577e7bc8ecd19826ef90b3b75ff0f23bfdfc060af47a043667b
z4db31e45d80b4d4af7c8293a2345ca42fc060c8e8d28969c7eb17d0b59af858b15af81ad1758e6
z8e0fdaa6697e01fb75bb14ccaf86213f2b1aab972e6700260ac896858009cea9ddf8fdb9973b46
z8b58165a0241547cb34b2078a132ad83de3f8cdd911e90b5c7f49b07027ac1439aba749cfdbf40
za91e1c34f7658bf27463af7a5e268da70bec20103b09b92d398b6644aebaa950f1b55f9b635512
ze5aaa3d55d342a50d2cbded964d69ab03a8353e2b192ec1d9fa5e3cc46bfa0dbb1622001a7c2de
z1b029459c5df97a65974bb6df86e855f7bccd6da195cc07a743275a350d6f060fdcff109dd2421
z7ee7b7743df48f45d52b10cd2f1fbad73d516b826e4482d3b11d93738bc8f1f1a2213b5ccd2b4a
z5d025e7840e0886e83b45d161b3ecf4418d4aed710f1e8a535f796749be6b0c595742d5270ac91
z20aa62f226a819b7b7f6b6f28524eb67e2eee42cf82c59359fcc5e94f347481763446974b64699
zaf0a58586d78a9dd23f4433a61663bc094be3d8ed15aeb2c131b867549ec4895ee138b49890f2c
zcce36e0d1ca97b5956488258e3b9b6146795e8c2f8a3df4df7bc61200f90a11afbff97d5955b1b
zcef88e1232f852764cb7c477f1157c2a4e35d1ff0d78e1149b0cf306e3edae63bd1e76c2b5a677
z750b419e6fe2cb255ce0585a29cdccb806faa7680eb3352a59ac34fa846be23de9eb8a65413135
z1bba795b5923962751e1b15d9a404d9c6ed2b5c9e8089a612ad4696c37610e8f2c88cd87f9285b
z9158754141f030121caf4e109180754bf9606f8c499407f47a465293bf99168c1accdcaecbfde1
z068536d337d6c0187a092c96422675d1e230a826b6e0adae59b2ea4a14e2e53a27baa4afe0b9cd
z912da5148f28d551a5d0e9af8137469ec615b0f55167d0fb1547d698aa5e5e852355f87918ce8a
z92291c4231e8fe83201a77659dd341f236c8df2eef534ec932279c1ee70f5bf0c677f1484df96d
z11daaaa05d787c791fa954d455f319e51fb963c1912d3bd684aacdc9ebfc6b8d4581e5eb43192f
z7df6a08a4decfafc67aa201c347d5e2e08406160e25cc61d62bbb67400349ebd8c6ab766d4bc9d
z8a136ea717d519834ef57f69023621808a35d454cb80cdd5e3dea1813b1b0c27ecd0119d898ce4
zc249e3d76d3da201cc3d9ef25f01731990a7a34f37e18bc1f49236ace31bae769385b50b8b8551
z4822688eb1ef0514d9284083a8ae91f7016a7909d2a5474f3f28748a2a88dcdcd90aa5b9485886
za21a6264d6c1aec4f6f5c813e8fb6c3fa52266a1d1aad8b21003250fca0583d5be2dafe7d88a92
z40ee59c5b14662bb1893657d76a867f4b319444951c20ba94d07738821a20efd26188bacafe87a
z4f1c863b4c4fca121a7ea7c72a6e65c2827a3edb23452ed0c990ea0080edd66b69d235a91a5b47
zb5117e5473c6f49ce91d9d1757c1d3e99b754cb2a09439a8fd93f87ae7e5ad361e12c4f6a1dd62
z2ee89e81c76e2e2925a25aab34ca51e92a3a098dbc3b5f5f55abf8d1705e0f97ecf36ecee15205
zce34df15f6b544d381d20c07e87b39f4418398a60ccb80572eb90551df3be2c398f1ce8a2ccef3
z7e80c48d7dde652c419e1e15054c8a89e2aef421ba26885802bbdcb142271900eb9b604165a6a6
zf5035c01a94dd4166bf9d58c018b2133796f239d90f380ab7d70bdb121b934a5c45d77c05f184d
z31898acf243c9a8d72585f256eb45c915f617c88f29e776bda543441259e21e501935cdccd4a0e
z62649efd2f930c5e5256229415ae127102c8b23937a853caba2a3d36215d783b447eafe6656afa
z1c30f2104bfc819c79c73c131bfa0e0274c2c9b39d6d51c390186e6cc57bc58ac1186140754c36
z23605ffb725a6ef54629d18c4b7ac8098a6dd8e4fb98db1a1e31a8ae938a57c43b4cddddf05b8c
z1e3ddd5bfc8f2db1ecce3c9ff3fabd63db8a36fe738b39b020668904f72f4ebdada7b4aa455988
z8f4f575baa81e7658350f5a783ba90d811865eebe2fbb95a651e8031c2433250f0fa230a3eba25
z85d8b94e5daa2490b49041ef547ea21a41f90d3dc6389f145ef66a10ff0a4b4fba2e412fb35dd4
zd2f98d5c5bbca0966e76bbba537a49c24ad4062b02f7cb8232133ae88fa00085b68beb43a1c5d9
ze24c5e0b28fd3c720f86522f06077a3463b50144e1f708f3f43240f610dc734608420a1981354f
zc7a05a312d5b3d976476273a482cce8edeaa987514bec7a20ad210daa0b403598b5485f7deaee1
z17a21da25b1e08d0d4087e9938eab2d198e461b62b5978e56ea7c789aee39f24bb8ef9ea15b126
z8de0633a58a733bf6aa4ae52fe04feac0b1224c314f4c9757f24bde801b9d10f3b88267514a548
za9a56598abf494f5d35ac4c8ac715fa1eae8b8b84f6e8950857859313788e10d7278c54367f5f6
zc7a6550bbc2e734215cdedd5111f5f831ae71562eafd9e417f925f371322634ba03e4dee7a93c5
zc43075a0b22f8e059aa0e09664c14e3f0e05da6cd8574208336a9e1c74acf8ba01740b65aeaff3
ze83f057691d1a05931e2a6b5ce837da40746c8709e44fde2060386f4013b6dd0a6a1f490b87875
za719d60dcd85f90fe4aeb2f6c63fe858e84ab84b236234d89aaf4f78b7c2bf0c5a0c7846d18191
z08c73e1006d8ccf6d86d20281a0e9e920f33b1f74000d2206125b737512a4489c27ee341ca376a
z5bd4708e840694d4ec6b1baf69159fc797dc8babae9de717c3b840cbbcf189dbec4d80770e5ce3
z144ce0dfea617c1ffb2facedaf0a78ebad66c3600e0b9765dc2e41fbbc163a9412ac4daa37928f
zb55c5fd3790da164d2777fc777ff3de875c221639a1c8cf0f297354d0761f9d47ec719676cf2ba
z15146d53778e19f3da043fabc95277aa306fc907a057d4b1019ccf61730ca136ecf6b29568f526
z4cbf4fdd0b5fc4ec5cc7f7706b625e3b4484f0cbd131102cecf876423334ab9587db3967cd5303
z3df8640c4d8dfedddb998852bf209345655eb141693932ed1353cd27653225e1d469e429c1cde7
za3150858493d11e4f5a8a0e1c7ccbedfa0d9c4dea6d2f75e55b7ad04fdbfe4ca78eafe2d62e783
ze9c4ea856750df24857be2cd0272f91bf000cab7e8479c6ff6aa9d42bcebd2ead98941ed262f48
z8b4f2d53f5c500a4b2bda4185ddc6ef26d23108334609081376eb4d448604dae43473208408014
z2e8a8a1b482a2ae411ed82dc8ef4513d1ebe2b9e493a748ad6d0671cb0c61b05b670345e513ee3
zaf048acf9f7be2205182df0566e410d77b98f9f594556290ee25178c0ce39fb315b71fc52200d2
z161c7377747afdb74581206f862de880c25c7d924959139ad62b0a5782e7157c5af44bd7ef5581
z04bed724844e6d4d7bc02328c10280d5cc6d3f2ec95b193866f3edb2df51ffa187dd9f6fcf02e0
z038e40be8301e19d051e774f35d12103b42b757f4f371eb87ac8f7be34c5c10a08fe7b635eb6e9
z67dc0d7c24e55291f2247a484a51260a78ee025b9abdea0615096b31bbe2dd0b2aed75dc0c9da3
zd3317c6c090e69f5760d6d2df3728ae871fb126c0ffe979111a2dfc0eff1c6b660917c6ee30f9a
zb0223f9d6c9a2387310548685e281ca011f874afa675801e84ca35a5ab94d69be0a4efecd50f76
z60f2d925a56a288135c8ffedc8a098a89f475b158d1d54099b2c08d0b9abdc8f3d9bbfda700f66
z884c6e5e749972b7d246af015a1a2f1290c241e95ec72f7e5e57d0c7dc2c56837d0e28d4ee451b
za90393af6b534cc0f55291ea99387b4b0e9f5a3c626d6f452c8faeb619e7c7345e984b32ba9a39
zc50bb1fb6d90566483891b4f33a338dbc8a8c5a12d48d01b2407a13ef399d2272c0e7e29d92056
zb56c778e300e77539c1ff055dbcc890ca7a018793ff763e53b24c578583a9eb53947368b5872d5
z6a6a824b982ae3aa9a5dcd4c5fa6bd96083d2130f6ed2c86ea963b5c46f423a50f6ef9f7b44f94
z50984f665bf1609007abd76365c946e22507f5f43f39690fe1829542f73c022e1dc00b2405cae3
z7370a635e43384e6abad23e2a5516bcf03d4d2c1170cff35fdf13074e3a16e651044a61b979b70
z7947e17b9be6dd2ca45ceeeab08c79cc62befc390aa67f751f410eb7cb0faf6de07440e0d1384d
zcb0949b3c07e1b8eb99d60f9a515496be6c86e7eb17acb0bfca5b2bc3a3ad4c80fcedf3a52479f
z3fec7adfbb93bb6dce34796c864b0f88c41ec495de9a6d56cbb80edc78d4f3ae1184963d0bdeb8
zb971f2dddbe3e02123bf612913765feee184da369ccd7155eff0e716a0a5bf401a577233a8406c
z851b3428025a301f3602d51310a48c645117469e87c977281c4178314140679596d528853f08d3
zb0e5c93aa19f0958d2ea0027ce97026fe3d20a5925c16817ce654a2dc0de757585872317ccb404
z73353edca6ab0ee6ed1f1425de9b69dbafc77974cd8a468b843435ebb16d23c376c6c461f37353
z630209996be2342575690b981deee032a289851bfab8e762a02801815ee1316760cafd93a6cd3c
z1cc4150c4091ddccffe6b743511c7ce89c26596e8267f747ce59af8e21b44471ccd60dfbf50f5a
zdc9adfef8853e4e0232206cde4b1e7e4f9e31ef1f3244a73e8e51f21ffdb3817618b8b8c22e18c
zad4438cb2b39a150200be2c01a1969bb4912511cf8b21a5f0814db8440aa58ddb66514a5b0d52c
zd5888135f7342620d4bac401c2bed1b7fa19f63e403e6308bbdb0c74b2253af2bd97a727dd71a4
z6b0dadfe5e11efb9a7a97b421af6e2136e71a44419cc2d2ca020c0fb37dbf4bded3e4c3c63a385
zc7c5a87cb514bd1fb9675fb1d98187d9ca46087397773e7469b72f1e709490d6356f32fea9c0b6
z20be9d0d0579227fda675b3997327c63179a9141affdb8d3291a79fedb17a40400b539e7364702
z349786cb987c91244c1822c855b35b0fc0c396c30e09bafa0a3c478e5a88a45fd9d6082146e10b
zf9c896776ba3e26c26096818f636d3afbac54fa981c2814141199a1a699038896216cc1fe09471
z5c14d1b565bf206a5f6bd93200158c79d4cd6f49ac609c0bc9ff527e80e958a9e44057fd289144
z0107e785c81eeadec296934ea3ef0a589077e598e01bee8bde7378b73195c904d7bf74086b1ecd
z8a196b47750c894f99efccd95f598b095d28640bfeb1788288aaa70ef73d544d5977df3a2684c2
z119e804b197980e17a7f1e320af68095e2feb56252fe69283e6326f6cfd6887677accd8591ad5d
z9fc60ef87d471ca9484b2311a0d060f5aaa31223f17679da361a73539b6f962281eee421f94a8b
z2fa7f474ae14f9ae413da0f1ec37d9c28976909803115a4065f2c991f1db9a0e9ef61cfa12f702
zd63dc2707904f508f47a4c6bc135394db6e8c6ee8657478a0739b6cef3c93de39b9a25abf83f11
z45967d8fbd240185714fb0d0f1482e0083bbede488f2dd4e10a6300220503d003ebdcce77a47be
z2e17a6db6358943af80a9c0c7083eeee75d1f6c2d798524a43baf002fe302640bfee418fa5bc72
z87e02ad66a1c67ce27cab1aae24036a1f25c81cf0a502fb7d7efc42dd48a98b2fe4c81663228ba
zea6143c9ee61024a4cf6aa4fa5f444a1e83bd24b027bab2d3cf76fde463922f89a2b2a4151c4b4
z51922441d3b482b140465f0a9f577916788496c96dd74abad4e7b0b4c58feb757a0dbe5f92a30f
z911a01d65476e403f22f09a65e955a11720d11b8a68c6f0354407383a00abc61d52d0871edc74a
zd0ad6fd5f45db1da8285d2e85ee553fc83ea38a9cf7934d5c477dcb448cc21b7ca535406dcff9a
z36f728c55668f5444180932ae15bf79b16245c258fbe07029c8063a57b7bf52fd814d4ba6ab7b1
z785075bf99a756f0e32f7e0f340edd7cd5586da1dd540aeb065cfedb47dd8e8b9ea47d4796e101
zb5a234f3c6d282e9ed8da983848d60d033361f1a178cd123b3dc08f6a1e1598d2a9f53ad3f8db9
zc1b6309c2a143e5b9f2e4ed35a6e9122e8f78170ced380a6db2ffad10d29b0832f11ff7b4d8be0
z1420a0aea90904314f1bb2206129187d3adc856415733877c1fb2912ca36e984cd84c1d043ded3
z13ca96bc5127cfc69a23dfc734a149557dad2a746b4eea44e842fa66357e0665b6e1f74ef16bd6
z105677664ec3f5afacafd2f50b555a00f7bca155c8e4c983cb0046a12915bb89c6fa358b0f1fca
z02a6cb314dd5fc105b5674707838a930e40b586f4fba4d9cf268d6dc4ca0096a935d3fc21459d9
z45a9d3284aace0b4be7cf053bcbc1d986f41504583057f3cb9584106d710e3aa2eb1aeb43a2d79
z2031cbb12e7009b47f8d8fdab750f96496f6036014ba87915478a89fe00b72c7a094a20455cbd1
z8f4fe802c2d02625a79f9311a6dea6fc3e9e2ef82d84502aa9852195aad0210d4773a0bd2a0d38
z3cb744dc88a388125b06e3114ae9a9d14dc8b6e7824b005225e05e7fe69b36d23b1f042117aef5
z24eeb8f1741c28a785aa5aa2ae4a0ee462f0e1f94417e47e76bfdd67aba1292bd57dd43bbb6479
z9c57d0d51e59d22936477284fd8fd4ad0f1ec06a501ad087c96ec8b7db2ff3dc8ec3cc233647f1
z7734ceed9a0b483981c8bd1bec86e357194a2344ca33a951bed4326334aedd4a038a85635a1255
zc24a6fc4e78de7a213b9e0748bd2754ed914025f0ce63f68ff2188301736e953be1e9a421897dc
z2feeb325d6d388348d70f40719af13a0acd195f2bd9b874313a741aed886114eccd0037b24b10d
zb8468e478c918a47afcce0aa9f62b0c69f877fa3840ab8753b2ddb283c7ebbbc9034eb064d6b05
zd69592c6ef01de139ae3bf42bdc22b5fc166a0466136091e509c94804d96b0828a8a945f8f6fa6
z3eff6de3cd91bdb65ca95992ffc83e86e8b4dd3c53e782a94fca536463bb8b660ce93b86700701
zea35f6d8637cf1ee096bc5f4cd1a81bcc72f2972c28277a4fbba0f7022f2cd18951ea5b1540f9f
zea8f9bfa411f0848cc2bdb898c8aa3ef41b4bcfbf88bad78fec9a2c9d4c6b62053c026d2781d89
z091942964af06d2bd846a233254cdb532ce993325d99b78acb1bd1f2d1aa4c84d80e472b5c8340
z384337f9aadea0fa0397485de6980e19bbcbcf5bbd64e4321351d999d4e469b5b919e3bb3edde7
z1cbcd71bf57d3044c5100eefbca52e26d23f25e490cac30cd90529011ef356d80edcddf1df3e16
z6e58eeee26391265b2b5acc65cbb5ea1935eedc58bc936d0b3b497d7b1708442de40d6923897a7
zcf3f681b590e8daf402315a47db9d5cac420f7fbb15e53a6b4fd052c8a63f6810b55745f6a1825
za1c7ea5dcc0644f65db8cee42b54a5e9d7d0cf9882f9234381a07e687d59bc0b0573bd9eb5ec52
z738b02335fe6f1e37da194775eca754bb8f6c067879d63a29873ec09ed3415c7bf29c3836b61b6
z83ea6f3fc50dd79e49043e6bf02ffcbe467ae72713219c2a742f3e7c79180975900ac2a595eab8
zae15e29bd9c2b4823f18cb32dc0aef33272ade79f19bde075884c80cb3ba78ac8c02b9417ea5dc
z30710b06687cc8542f832261794277311183c8a18682a3ce3e402fbf0b2f1937c2addb947156f1
z84fcc6d0e6ea58773327ff1d50a78f1eb5a17a41f510617322c9d1cc855e8bab60230438a3cd57
z993352f85fe4714aa8f89b73e665a2f8a51e164b2d925e0ba5397b065983c2bbe8eee24f5fe675
z58005d26880a68e79f6dcdb49a97bff11cbc0567189107ad2fa5f0072144974592c0bad4f6af36
za43ab0e502dc6d7729a924d4c48820dcfa7087f145538b7071ea218a1d06012baba5c6a9e0907d
z0ccee892b8796a7b6af0f7efa3fa629a3485a0931e524f97d995d64aba65f4cadf6c6797ad2f0c
zf46e9de33f3a686f4eeb281a47c0ae264faf4e0f8fc7b41aaa7b9e52fe6081b46637ec8c0ef150
z58ab080b60703b1344f6b664da72e64c55c7411aee48eafe2d28514498eeb625db2bb2fa9516d0
z1b97d1eba9bb64a9ac916946f8dbe08bca1cb1e35bebf039f8479d7e68793f877294335bddcd9f
ze1fd51ca037cccc25d560f00e031c49cda873963afd0b4e22edf158c7dc454681b02d7e32346de
ze135f503b3eb62ed997d54dfbe8e67800e009fe0bf5d9c0b6b7de94ced07ef3b294f04ba5b0dfe
za95c89a9907a21e4ba01427b80fa6cb09896116701a2fb65125e4963c9ebabd40e6b664549c820
z55147cb1141a5032264f100fe874780bdaa92ab7128b1fb153d0100e274261592f47a74bea3cfd
z1e66f778f3d138cf1a0f9e0c884c8c804c8b24ae35ac2441e836ee67555a5b0992e2fff630a33f
zb0b9ad75cdcb8cbca237f61f34b29078a7fb894850e25924b288a32921464d07eb2432d3e168c6
z7e167b60b5047d64f35bbc1f7bfe9b1001add48956cf1215c6845133acf31bde807cb633edfa91
ze4e1ac97267a502e98fbd89a8eb76b5728a4cb080d174f0e76120f4b93a225d4d57325ba88d484
z4b660a88cbd89dbc6f9087de61cf25401f99996a02f6f40b39fc1dd9adc09a7970c2c06d7cbf7a
zc3d17c4c1002fee6d4dcf8d25d928c9b018375af88dce4bd9286237e921e28d9ae5da0abe4223b
z744cff55defbf70acc9adff3e3052f2743e0199e8f56c3c44a5758716817a9fbb0ea4429ad40e2
z07c7b2253043056f43f4a1ae6f14ee3dc577d9afc38ffce97738aa3557f5df099d76109a92d4b1
z7ba3bd147feae10414a115a0e918e8de8d001941636beaad79e092989206d1c8b292b67bfe9e74
z649685e818b13fb987f63b743771ee34fe74714850dffdaddafba93c887a548ac3a626055bebd4
za15be77fb44ca040e35d567f540027473e31d1ff512676c14077ce8ef6d6f41ea79fed8e9f1de0
z70ea48613c0531e37589cf80d43ed2e1446146ced36849a344db428a79f75bbdc521072b9495c7
z57c46b62271d200beb5c9d852921d2f9f1261a07634bac146449bb22107e1d8485d228a0d2f263
zca030c77b3c8d9f64ed4ba49a68b19c1ec24b9c02b3411b1d110af1611390affcacbf043331fe8
z0cd81dd92b75d673e743ca25408ec2a91507c0d8728ec79ac7b04c01ebce87f37ec9a987985ecb
z6afd3ea687beca6cbf5017f08c7429cc7bc192c859713ac9663cf8ab08d959bb421b43f4ee7464
zce2489ca267b98592f7f9c5d117be53b6b6677a67f6f1301ab20d305a6656d452f3990fe826882
z45dcfa51651982f00966c18673f96aeffc467b8b4e572587ce8cb3fdaa21782491b824b628bf35
zf390c8aeb48ce0f1147216266019f95be6ebb26a2d98b9c1a02436054d190bda95a09debff1de3
z15837647dc3b2a23e27be5a466e2a2b76df0364d921482129c9cebca8e49ea92f68892710d180b
zfe3fd88276c0d9be2e37d2dd1a3362eda64b4c94714f5699cb53ebbabab71d997f9083e54e6434
z92808b6f6970cccd127a5ca9528bd8151c96dea51a711c00dad84f9192e9b699114c9f065ed479
z0e1fba648b9ade58c2f43a3e7a771c727807d5d1340d4c2ae4e92641de7a1b3ba9481d857f5c7a
zf98e6e7312a7a49dd64000cd6efa173b475b10534ffb804d11226462ae67faa0fdbc875662e2c0
z5cf937a0cecbfbd2eab6fd0ee5961cf5830165f1bbf6ef10cb913725e362fa56f049bf53decff5
z7e766d552fde0d5744fee66d55ee5c87d572185c9dc3002b5be6f1564a5396292a158ce94856af
z173fb6bded6f8076118cb7d7b4d605f1fb4e415549c08fb04b4c92cff56944f6131845776343b2
z32e1238e15242619ade23f0d54135cc26201f710a53302a0f5202af9d00a1d7d451500cbb6405b
z9cdf40a34df4a1358c56d30cea9f8982a6d46fa44fd80311705b0ae1bf1d4b62eb10eef8a2f8a5
z8ae55c9f0ca5f939aa9386d25d08ea8fab33fa5942ee75e9abe0ca11719369ecf22384d3c76265
zb4653a39cbd59ad33917c1dfbf1ced886d52ae8dce4f50978a2a70b5bb7cedc7d8a629081a184b
zd5815423c77a20dfd9f4ea9acd91b873fd7bf5b32fa207b0b48d3bb3c2625ce6bc528d2c74685f
z82eaf13b772637bdbf3a20a805aec26a601eba0204986d4fec3eebe6990791f9dbfdf9202b9f90
z02e33931d59658ed1999254cf85eb6ec0aa4959267562565c30e9f8c4732bca9c39489d02e192d
z7c50899c63ce90863fb7de6ce38299a1b8dd8bd243f3253dbb03a6a00c21ad3792a4b11f81d051
za7ea2f58bf054aa59878043b56ea5749746808f9a50f7fa4143297b44225e4191c940f4e71829f
z72cb1b245a86a387c4bf351bcd5ea2473159599a70ebbb71cbd46853826c50510c7018d6cdc581
za52cc19dec2be4b6d1e74ed643656fe9ee0e685fdf1dbd7cd903317901f1d1fd3e1e0db2cee86e
z92a85648ad22f75942a0f16cc04b2caf2ded995b7f1030ffd2c72c5a0ef4cf1230b349ae5dba47
z86e981bcfb8970b6630c1b18337abd2aaf86a77ec8a49aaaea266f50c302325256fbd76f86a08e
zac291fab776396a9718f49652e80c7912fc61d42665ffef3f5b6b093b329ec508f9f3c3f061164
z3ba8d06b67d4beb4d390e7fd63d33f8f6a90d581051a10f53d253e00f11d2782bed9386b35255c
z13e4d978fffce7504f3b431c206a68a5c941fa0dbcdd49c6b9f2c81ca0634d61bdd2b5ac01245f
z04c40dd2af14aaae67e74905c1bd13b5eae040de4ca98d9a93e0494511dfc8be23b922825a375f
z59b4026b6eef713b6ddfa10737ddb1305328a0e67b5914c38683827f4bcb25b482f358d7335636
z63a254ce5b0949f802f0fcb44fadd80b4aaafe9e55cf7b795ebc8ece83334cfa3afd4d5dd45889
zc72c1a05df12ad5dbdd06b1ab44c000ba4475978f63f7bd992b0415a095dfbeddea72035949d0e
z6c7251aff6d572d874fc7002028aebb669b63bd36893e0a0062c76809e7ef9a359c25d3bc8d949
z40ea448d0ec981b79487d8f76b7ae50101da5c44c21a50480b5c3bbeaf533fce295cc4d322d51b
z8d49e056640e100576e0a2d04a4c76d60c026e6dfacf50cdc5623b219764fb642a4e5706eec944
z0166511d0d0c0ed1f9bad4de83240fc7cc6ffd4d66856fbe0aa2d454b3adf7716d9ed9eb4dc9bb
zf5bce1af23dea737043204f2b1bef72c17ae39a48edc5261dfa20e1ee2c7a809c7321ce6a83702
z598c399248b481be7881aaa5d5ae208b34f43c1c0924a57f2e6c2c9cd2bf3ede3054881e788bd0
zcfaacbe8ce3eeb6322ec73d932f270209b4bf89b4bb3e64cd7381088e96a0a24725b947cf43704
zc1e1f2b3630c60a2317a1b588c398ebd6f6977088320a4203b02c6fa5ab8a10cde79539b96a48e
z437c791335c60a98bd628870bcd2ebe4161e4a5447f14fe305a8b8e851c2dea81da16b0f5aba9d
zf31d4fb9da35b03f28347c7143b750a00ef13af9037b4aeb9de21f3bd5203555af24d5cdf5318a
z089f818fd75d9d6f829c27ba424f6a449b58a4b9e5ec4fedbc5cbb00cd2ce3629a16ef2178d67b
z19ececbcea48b8d66fd1a34166b0311d454f7ca2341c2e8487f9bd0105d45f42d631d9b01d9ba1
z5a15eb705697a62f530e26bf5cd35dabe29158800a77143372b7961e2eb3c1f30801193e5506a0
z8491b4c3a5a9cdbb61b5594684e9ad76505d896301c6e4c3f1b52ae663e6b12642fc2698008560
z1ab072d9c657a455c8fb2e3b74d29d39169d48896eb9328ffcd3005ca6321e1efc2ba0821935d7
z133b7e23caf7faf975a65a2119b4881c93964b1c65ad8a85c4d6c45d1baea95157ebdd7b01f0b9
zfb86d3a848d2ba6a4d8b4980b866925801f16429471ef095a7243b5a9e089dc76d2e1658c62204
z8f893a1d620a9932d1081fa3bef04d126c2f46d41035286b0e00a016af96e5e8a335e37837c1c6
zcd73af6ab121777b46dc8655466b812efa3c3e002f2dbaa281e0bfa49dffb64e71032f0ef2ee5a
zd8b8e1531e9da60903c3a7cd3e75a536036c4d5075e52f61871d20eb7711e7d1c82342ba4cb7eb
z7ec01d8310470e44f751345cd7bfff8757cbc24f306a9a2f0d5c707d1bcacb083f4d5de261e8f8
z23fb9b6b47418ed1279a419400d572d95798571bd97f7ac1a294d9ec5c72dbd49815860dcf2242
z7a4edad8f98ab098500b47afd81d584e23bec7ccb9e80381707fb6ba3cbf9a933e5a5f403f2ee6
z7263d73dc4e1808b528fb78b467a87ed3fe1254466995195eafab768d0c5c879d2ece1dec449f4
zb0013dcda65876ff5b94f54a0c12e1aafc3f4736ffcdb21eaf620705f51124d32114734cb51409
z1cc9d3c03fb49185453a6d7a0303466f9fa205a505d138bfa6630c644d4a129a31aa48602ea9a7
z8d2c78d38ee11a90367f8a2474823db032ab106f48c156c4782a32e35c9310aec960a928f04ac3
z105690a125c1148139cf839c7859e33eb63fc2183d27ce913edf3e81837d3d1de148d5435ce896
z376e3de42717c3c9449f44efd3ed60e11160c0e6d0ff9bac2c179a614c29ec682eed45c977c0e7
z04030347549c0b9ce2a02c18962a4dc10e0eb6a75e7acc5671e6ba5457252df2110d4efa7854a6
z93c750e8af5cb800db8396fd8439d97fac255f6cc04f84c9102467f72880b52892437ebb3e6b64
zf5de0761d03f4103d40c578a85eeb908ffaabd4d68c91b44b14bf0511c871233dcedbef3dd770f
zc2a37828f7244f9e9dcf584e603528e8fce0b91ee0496686242358fffd87629e2b2c6295074d8a
z8dba868678b5207c45955f742cced530d4048753dc46d0c01f769260a36bf89db35c142779d7b4
z81278811e3269c110b567183302607a73d96161f7e1dbc4cd4135134ed8850811e2793dee64463
z41970d6c3da0be74e08b91578a2288d7a035115a66b465ce25795e9c097f14fa1fc597fc60601d
z3d538c3e04ae6c9791642613c2267321f035c4d9605468534bc03a29c8dca3713579396b1798f2
z26d2aa6b8138dfca6c268ee63463d1a198eeedb3230dfd6ba4627726cd62780cdf583f6267dd49
z1c6375aeb4ae58a4d74edb096ab3f019653829f1994bf1c98b899e605763fbf4ed73094f24937f
z9017998d9db23737327431a9bb59041bbd6597bbcbc97103a5049f76a384529c2bf6184cfc72f9
zd4d784a141920a7877342b843e2f2bd83ebdef92ba7b582c924165a8d0a8aee0b4461fcf9cf8c9
z1d842159d93cda3704d9c12ef17dd234fb52e3f73100fec11cbff5f14c169928378a580fbfd635
z229f7acbf5f372622185fbd2eaaa9e5947e114f2022d754fe4a5806f569d1bf239f514c1b9718b
z732d1da9493e6214eac5b0b02c70292cae0ad0b3c5a03c4431c6922cb9d611d23f1539330ba86e
zcfe6118324046a8692df183fcf1e83faf71efdbcf404a002c4df015df586a30e72486b79991817
z73d23567461a250a2db6846bea812043bbebea080a04ee010f08a9f67a3b1eec888950bb12dd77
z52940b9df9ac300b0ec822b4be1038a9fff208f4be7046cbd0c8b6cdb0311958e139742a52509d
z0335f1b5c13e90c099ddd77d0180d4ef331513aa507f1bf27cdc30f81fe3a9d1d8f4c2c1e2e827
zbf405954266092158592966053553698dda179057cec20dca7f95776ea7f65ed4165c4f85a266b
zcaf52c212ae810a183e2bf913a7ee869b5b57a2abfaba0f49b5326cd81095959de2a05dfeae511
z26fe2a3cb50803c76468c9c43c73c2d57229c9bd1c43bb3b9dc6ae9ed1c1ecae5f0ef17ff44c49
z1a875b3add6e2b76f29063bcb81b6faffe6b27014270d60a54bf2c08f1b5b634561cb250c9d9b0
zb261664cd678a3464e111c6004a572003073db92c667026884e1f0ff0126063216d36b74f185b8
zefca7ea7fe3f9b70804904cdd19e174ae9232116d7dbe51137ad5432db2c0bf87304db9c2c5f15
z2e716bfe51012a4002a00347cba327df4f0759b8796d4736273c63c6eddb5764b7d21addc77b7a
zf0de23439f7fc4acea3a3409d645478da15edf1ab5fcec6101df87ba295f349654a742d65b209e
zbf7a9edcd4839ce3979ec2f2eb5bd98009576bda1dba1e761fd2e4cfc62214068352c0dea4aee0
z767f7ce60190021946c71a8a2de13adbc41603ca06978ca385f53bdaa024fce15f83e7b395c7b0
zdd55712db655435ce040e54108c612f77d9cddde5b43d906693fa52683c77fc9b73d5f85c25d31
zc127060a8dd431086e342ae4b896e7635eccd99513dae22318d655b10d5c550c62464163fd548a
z0b61039a88646d654aa6261544d7bb650bb81a58886ddbbe44abb9482ef7ed53869be44f494d4e
zc42d41fb401e44ec8908b257811600ca369750d49422c89bb41ca125161245ea37532c52052614
z64cad1bc1478965d954510621e55f05c84e532037618992b292a2f3d2cd63e166cdff1011cb8e2
ze00b412b4f86fce65c4248e90e2479969aabc84350ebcf8b05d08e82d2b52b828b53d63e0fa956
zfcb68e89ce784d4723bd1eddf1b0c45b53f68376959c8f4cf30662b6537dc48a82a040402ff925
z8ed0b1af61999438187ba9c6b8f02e81a7bc15613c4b4b8eac9c6149157f4c7865af242e2581b9
zfe94bdfc3b69c3c1db90fe76e54cdee33c3bf7f6c335d43bafacf53144b38162ae87cc58e016b0
z9c6d6f483310772f34a48090a5491cf33c269925b60ad365467eadcac2deeb7377cf432f455cce
z9f47d5397f3eaca2f62435ab4df7588f17fe3e8637777c76e073b8a668a3295832276607d38c46
zf28f9a9ff800ae3da585b6edeb079349bba4f631a5b355ee7c7fb4d2245127e6e037d17f811dcc
z7b946f062d201eaa274ed6537deb45a5b594aa89fefde5a19b413bacefedefa4a242daa56ef6a0
z86254376bc254e8feae88e33ae4b07a844a4369b32699a06ac917e477ab0f17d8c29bfca711d52
z3195d6bd97b4dda04527816ece8a5c21e5f79b5ef30d6257e2a4e4743dafb40c1d0275736ab137
z350ad8dee93ca4532a28244eb2db57ada0f6086d644deeac21c900379c850a3c4861be6d976cd4
zf90633087556b4869781b5c464295d72b3022ae7f2097c85fffc8c15d9c923bc72d2e31c9066ae
z22a173c27b55bb26e04cccb677e816790b7dd0537901296d19388509665d2f908755da7056a3e9
zb9a2755acf1ee8f64a069f360a4e4f581e6e53890d2c1b760757248e9364c38951f3579e3018cf
z146ae53bbe4e7e49710a522159054d22c657fee121f586ebd6b55541ab86e0a5830aefa3ce2f1c
zd8c2182dd9f8ed19fcd14971f56237cc5488e60e5f8edf727cbe20adbce75b72a580772cb0ac7f
zd2ff44f3c70ae81232f23d6005ae7d797d235a3749e16d3a7363e6f4bb6f3e1f52ec9e290f76c1
z784116b3fb4284c98f82f4f3962909b6499dc57d342bff90782ebbe48b4a9e1124e43f3b1eefbb
z67439d0fc7035fef16d810e4be38e01d0b9b4d77c24e43fee4bcfb81a965ccc724b76507babe5c
z05c934f310626ef3c88d987a27e0dd23a744846570164c7bc913d25ee2240cefcef775003a9f23
z8bc75525de4fe7ca1d07cbfa1d16d3c1048d3341d3be9d83418fd300621398351120068ce377f6
z08ce65baff59ed8dca371a6f715f6b81a82e3e03e73c14e9e6d942549bcd2224bb7b2c5b0ff0a6
z4a8c3d52366ec471026baba41755f3b629f2acabb2709f170e10ecb979c8e0a87f81e3bf6ebd61
zde7f4a2689bdbaa0e8513d6d893b46ea4ae357806e7c68de4c3c407c4921d01b69ced7fe600185
z9ecfc2b4a69924a2bedb8110a4eb51e94a809654ea676922b66c8afd76bc43e5e16d1c81c1005b
z8dbac93886709c3216903001a6bc480219fd52f9403b7138eda3f4166cc7c7b0e09be6ffc5040c
zcaada17314a35406b4eb3d04411bf122b93dc0c5091c5e282dec8efa69b37811f95a76eeeaf80a
z258df68f5ea4f123593094fd77719f5a01c8828aef8952e17b2277e9b1c7d4ac1353f92f7579bc
z00819b6c4849deb7a602d574121411ab0b1efdfe757ec1c2a258d7698d1e8490b9c5ae137a0874
z8418d18b0ee0461bfd15315117a0046465d6f54d0cfb44db9cd67de280e61f20b4c414201e101d
z6ed60321ea6969dedd2ef63ffb176fa7acb505037ebf545fc71493b5c5264a278914bfbecdc1bc
z8df646ac1f462d65e661a520b415146f4e5049b38f382c2c7778c3f6557c67a5beec19dcde633c
z1ee5da9eb501b29ea6b89e6b5b4815c4c77d55e0a2bea234fe79b388e6c76cd3a53ceb481559d2
z754fa980029b08de69c632c3c6301be64979549edc0db41544807e5397c66ad2c7d306a87bf813
z6fe5fa131e03e455f27729c915d3eadb7449db2eb1f70e632e4ff9c4ac2b5ad27271f315159ae1
zce9f50823fbaac7e1ba6d99e7f78ccda7e70a06af56a33d027fcda794a30933027d0aa1242f3ff
z031343ce96591e8c950d50ca92f50f42ad7f2efda3ac0f621021e0792d04b63d0c508e6bc11290
zc4eac0bcb5343057e33529573bd1d0c79ca228cd0f4d8d74b637abd513f58f87c9907298bc0e83
z9a80ef072785d364ede06f5d1a4513adcebee00e0960d35cad3bcdd33e15be6c1f18ccec74948b
z62b0e9cff1a5865d77d40c95202e5bc82cce20bec38a1ffb5b7e0c3e2e7ac43ea22c74cba0d010
zfbe5edb460963dee20f289971f02ad87e89844bae73cab4c6b7f9c57c0a03ee4650fb9270ae101
zfe5aaa6ff93cfa20e117bd41cea395e041852dfc625188437f6c4ff321d0224f6f83366e4bca38
zdf63b135c88b2c687e5d02c3e43a1629778c8070f57a8b296e1d861fa67945300bd89d232f3daf
zc1ada3bd47fd47bf625c2cda3b75f613daa219b212442abc1fe947f24ea571f3e7eaeb827741e8
z83acf5b341f10508c7bc9e7dda65255634d3a16d3079dff7eee7ef6aff9233440ad784c9113c91
z1f85ab22ca5613cf947d97af1b2d6a0f56f6f2b63790b8df90ee5a42c13e1c02d140552a68a149
zb997e9d48bb62db26aac297ec71d99aa7592e7d695773402e7b5e3995e73a5cee9b0c7ac476d85
zee4859c3d46673545a61bd083b9adcc06ca236f70c80784003a30af6438be22e7b4379923643dd
z0c792bc7fc6fe435340943303f7255d429200df27fa92dbbb49cc6c678a3820f684fd955b1fcdb
z50232b8f8dcbd2ea0550dc3be456c5ef50bd0fb8ffdd86d57b465c8a86e518d14f69bbd1436410
zd8a34884d4503e336d11b72d04a414078d892b13185dc03396284b9ccff0f2c3701738ca27334c
z0fd2999780a05a204d95b9c10b31fb0af8b97c65d03b37999775433da00bb5306b11e9bb40c159
z4c507dd201c5a0246846d9d313b8d30b86f2d6ff6b10ff91b6601ae9d2e9667980eac26ae1aa94
ze73524492afdabf764ac5e80b36d74889068983c57da5724891b712aba98efab367f743ddf364a
z0eab94f7fa4111d590711426549b98119b957aad6b5a167b42e83df8ff7ad6f6cc0c7d8c775007
z7125d8ec5fbb778911e24a8b766806f641749a7ecbcf96c9d605dd208f422cff064d7ba9083bbd
z329339e932e46436c2e00a3c1be8c4704317fa5e4a73b54dff29656132c7a12e7b4964236c9cc7
z2c6bee5bea492b16a7d3cd2f5b4ab565aa9aaa5d0b326ac9f3041046976f51ffa7aa587171647a
z0e46e9900fc50953f447069533c4ded2a9830afad4aeee66bf1e4bc9d7eb8546705384736cd2bb
zdbba568772a4bf1758aeebc0a89ef59502f037d598136be6e7b4724494bc8f0b1d2a02f1a6bb6b
z69fe3ef5040445bcc9e9f2c9b3fbfc77c7e4914ec5b009f4e17dc9a932c9fc59d7c26c32210fbf
ze87a7ebdf75d767ef4528bcfcc025920d2e09074b96394fbfa196eb5485242c619b7e01d387742
zb5e143297c1436e35393a9ceb4657f10c520cb3541318e7a186dc5b1f9159334104073d404ad2e
z97950597e65cbd74ded5fdebf1519d6f02cc286ca714100557b710dcaa650563b47e59d274909e
zb76f4694bc65e92ce7f6274cae8d5049fb111fa28258a75480738c7a29dd706584833b36c76574
zdb91bd88b315e8591b01a2388b2f077bcefc2ceea84af6fdf8442aa6a06d15c601335854f409e9
zce5229473e4f810aed22304146a84d99333b00e9e1a53147f67d2238c9adde28d81835e3e18e3a
zaa974e2501f607e0cae34355f07f5a831375b34f1431b3c1cf510ed854e690aea4842e7167d02f
zb7426f4687233a8e05f44d75e1b59ee3e22b4518a43fa8b3145adb7b94455ab65e68f30a299ad1
z720c7fc6da60cf199a9fdb7df020601e7b41fbe6cc6801e1aeb61d0a128d1ec486c5cd780f2f95
z7b32061db6352bdfeee0848c36cdc6452dcb3281a4591c7783a6804a03d896ea07d4b21df17760
zf664270fa335e4aa25a69e7699731a4339be4764465042f5806bcd90a26d6d1628238f69f37165
z0c074fb706bb35f60a41f9358c13b1689301d43073b3e6abd73b30ecb7e09fb62d1d0ab40cefc6
z76e95c78b2c0c4d7e84668d8d99455b734065e9a6df722f5339e5d3cb2b065c0b24c498870a8f1
zee7aa9105420658e0ce3496e628f75fb142a55868c3fd10a75f5ed3501b8bdcab57e0a8fed850c
z303b7aaed76eb53fed2dee5b0325e1b326625c803f7d1d01c0f4306836ad83dedb978bf0c295f8
ze1bd10afbed8446239b36635a8bac3904a0aa9698637257f0547305c86c7b8d34ab30dace0baaa
zd7197f3ca504391a29ad550933f9a61d4a8b40d11d464be89a50c0d24758cc53a158bb745eefa3
zf979ccb998717979307396f790461e32bf5b3f47f4ba0b722f0110d80256fe73d957f9456d0aa5
zac64e9f061ac317b8a96149ed0b000d9a151a866647b1e69bfd62a5a81853bde0fba0e58ae332d
z2e01615ca28e8edac2679302b66a205b7bda67a67cacfb96aaec9019517b5109c420706038d1d7
z0111a0ac1971fa912b180c1b12d17693c67cd8f5cfc188278c3967d225a85dbdefa8e8e9a5a121
z6db2484eb9c21a04725402d553b3125369a85ee6e6358cbdc4ad3509af9d0f5ab443c2b5907671
zdbfe966e3aa11dd335cc959b8ef368d904e4908d3e62615838ee5e019d75816f42c46333887826
zdeb2a3b4e2056542b9a2ddb9b9022eb24d674ec0a67475478c32feff3a959dffee882f81c95fa4
z52c92ceffa4b4b922720153df1f4ee2808f170ca89f37a6c022c77827acd802a9e323e2424b983
z1c3ee1957680476d8107e2e32cf7ee44d169ffecbcd877bbbbc4a48e432f96071d33f7cc109ccb
z510da0db10828985980e323d3806ee7b65c1868c41c8a82b63f62b4eba124ad259164224ce663f
z5cd8918468036e5906ed1a37829b130d01e0c16211f190e333a9cd9283ad9e4b7178147ea8377d
zca8694d21c7d641492445a2806fe389af01e8589e2a23f52d6442e3ac3a0f6fcfb42038b099999
zca07f381954eef8c5efef47b8646d7428b2e42e592c02586b5bbe984b201f7ac82e4344ce5b1e9
z7735ca5b48d450343a394a1c4d6b1997eb12407629ae4deae0fb65d4afef50950043c8e0192964
z05fd6c08cfdf640354bb7ddcc3d9bb308cc798d936dc2aa5e6022af3ab1530f87e249048d8bb0e
z5f26077f5182de67b445bcef50cb15e88fa5c8b99a2a3586bf3e3188e547fdfaef28009db3a2f9
zcf3d3eb4dcc5f54334b796bad2e76be58c528970c517a9d28961042d380c9b3b0073184d36eb4a
z804ad5d3f18f7940372653aac63552ed006a0264d454602701d4974a023e2fa7d6a7f169995de1
z977e97b0e040898f2b99745c606813ebd673689d6006b07626d867b6449ff7e211985b75bb62d1
zab0017ad7bdb2e87757f0746d3aca71696a0205c683b967bb3eb41a3cf5a50ba6e1cc51e81aa62
z39bc04552115b1910d959419169d9a8c5ae89cba76f79e5f2eb93f18ef137421498f095073c3e9
zfaaddec381f131e416041e91be9871c8548cebec052d3f725330bda80335617cb99a9719916f43
z1c8a5cd5247c1445f04e2f0c43c5b18905cbe79d8d5eec79b82a98446d92557c8e0eaa59df6b14
zbc9eaede17add5408f21306bb41ea241675ed854f2074cab69954f529934d7c28225cecad3fdd1
za0ecc16222139ac44efa87f632ba9fcc35a0b221de138a0bc83d99763bb1178d45504cab96e9b0
zb35770146509a36f9c59fa48cd57b9c49251c1c27d93971a73cc1fc13792b355c31e58c770af2e
z7a09c48d757213ae0251d2e137473eeb240e79f735dc767ecee1093e1ba536d4e67e843e9f8716
zccdec306fc5aef44bc6b0f5edeaf9a597f5f3e30af1d3cda68e16262bf2f966d396dbdd2ec8fa2
z4e3632c40fe067097ef824a60eb860bdc530c6731c3eac1c9e5480b6ae581a5db8a2aeb864ee3e
z3e4064f87d1a8b80a3b140e182e39f00176bf15dd4f0973d82b247ce7f4af9ef1eb173199f82b2
z2557626729cdc4e9a371c2766489d804ce62bec2033d006c82a4ac0215985748643f2c2d2eb337
z3180abda83a73f9111ec447713c4b5a595405d0d8643df9111bf3c460885445adf3bffb3dc2169
z381da688bbf97a8ae153dfd6766f5dc5aec3b030fb26be98adbc7ea24bd0c38ab2ddec98cc0394
ze82ff04dbaaa3c03a3aa307afd59ae1dd0e178a2b047866188f7302aafc55bdda0d173a3397d9d
za30c171424938dc0531b76e9b3852c3156d817629315e3f3f45a4926c0041f3e4a9490fbc13822
z4f329bf1b71d35c62da91e785dc6549580db54c9b16b443349c61ecf3040a266d97a6a04a006f4
ze97192791c33d3bac8cc28a9f235de53a0430c18c0ca6899eb973e851308a65c6a00f2faf540e0
z8328762f5048c32aa34b5a3d5508e3539c3b277de329398d99b5f6bcb89febb7b2c7494c417c66
z9271841e26c816b673bd0a192b2e26b306e08482e9ccdc96c072c0e2313c7e065f3342fee60663
z6f163c7e1080fbe2eaba786c543d0520ee9d71a6c487be46816e3c2d1544b3725ec1e9c969edf5
zd1ef0c3f124ab2020378f400760bfc518dfdac1dc81689a56ababc4b2b70153656b993bb230338
zadd2c38df98be8be80e7ea4946e4f7d1ca530abdd3e886a91b382ca7353f740bb377ad646521cd
z21dd261db4cf5528658d844cc6fbec1e06dddd2446fec11c34bdf6a07ec125189965708ad7ca03
z7e7d3269125581a80525212f254374d5f0e4bbe1b3034e2d48892c6988554c2bfce3a1c2dfd98e
z0eeefd1534e28885d5e06771e2682a3ca158a573e28c325de36caf3a787c93c28a2010987c99cd
z27dd103726da54ff475e5276cc885a9092c3032bad9a690e4a0c413742b6dfbcc36f11049501e1
zf58b26abca90acc3fb2f96a2ae2507e537ffd676f1dfc26b598e89fd5f69328727afbf3a8bd3ff
z2ac39653b0ed5916d8f7d1f104d2d785ddf9be1a447b9a6b6c1a4f80c0ef170da2685d38a22145
ze609938d77e4fc8368d36898f705ac8755507286470609e106fcebb4eba520753249a4aa6946a4
z6c0c8f720aedc04837f40f0fce745eb7af558c376d7ee712a46847ec2d468793cc313926e2735e
zd08e084d75a7c817923b1d14eec39ababd4bd3f3b7782a9c9a2696fd2f8b536a5f97778965dafd
zd2801931d93f1595c2956f9087d983be40c7c97b6a53ead64ed2c7105d88da4c6ed2ab4acac91e
zc3f4d2e3e32f5b16fd62808088ef62f5025482eb6d2a60dae7964ab44f691fc5c8cc41d2bff91a
zfc7bf7cbfb74a1e62941b8cdc98c22fd5d045b23ce031236563ae2a58adb3162dc40f1a389a31c
zff4010df73512bda1cea414094b5c88a3cb7ea9f34bddfbb6b1d5e27b2f01d51a40d5f987919d8
z477a71f1d780c03d5b0896601b785dea69b9db521780aaed6cf8203f9a84cc390712076218054e
z3da16f21f4a697aa33fa9ee121a46952defa7686af11abd315ff06888ab99059b57ba0ccceb06a
ze03201114aa95bb2e5bef3be36aa1275b2f0232dd2fa5022579d59fe51a73a4aaa48c1f9ca9487
z4418559f32b3ee30f805cce4635c35c067294951ac1b7de95069ecf2cc3f4bf55e611ec2df0a26
z5ff59188db8d1317904b81e0aa84e0d3b2c53c0deb5148a0df47448b0ed76520bcb392f11228cb
zec7943cfea35dd8afc451916c96307850ee30ab93f1ea1e18fbecaa01574a4684e0a384109f353
z4239812df91e02838d84aae572f37c3c9dd43ae74e41221f23984475ddad2b96289581a18bc4f9
z4db02bca60a86540c166e5e9b6be02455303002fb9f8a6ba2bef30b7c96eba0a346a93da81a69c
z742599ba548616cdc3450ae853b4c697e24f4b6b9b6ba095cc28cb8efb8a0c89d2b0474032055a
zf5775fc7eb0e97265bee532238b7f539b51dc2bd95f2c8fc4d8f8715a9642c282a120c9133cbc0
zd078f021597a72b9cb4af49ffd3296df62a5bff3a00eea79aae50f5cef0c9490b4630dfb067b68
z848d373c589f5fe80709d66051ebce9ad769bf547a096033b15f04402f4454051b70bfb246d748
zb23ec5d520a6b50ff7a46b6cee09f4651e4e80a8b329ccccfddc573d0ed8b0f074db5fd4ad5152
zaff94a4aea0d05d69092142d42b12710e1b59ffd0b95cc2084c145eb7d82f5db3584a94f3ac071
z10e628110af93d6fb2386a44efa30e6af5a889ee457b33943d05fddb32d25e6ca87a39eca56ca8
z6cf777a13fa8632d564ebf34eef6e3253e395eebc05507f5650af76ccc5a76719812fca994a902
z5df14e61944f919912d25d30202cd869696459a834ddfd6420a14fa4bba8c2815b90e314f4838b
ze7e718b801dcd106e9e0565ac9c343efebeefaa2fcbeec2a170c9560917654344248470a93d38b
z99e4af65beb228009905a57ab5edc0d16fce5ad3d08b804bb5636a778b202c1aaf828a9e8577c7
ze53420c563c564afae12d6fee6ef98b0b16da2cbdc125612622e4ce07d9cd016c4133a20199d69
z03b4c5903f3bb6ba1722cf2f16dcf430613504dcdbe5dd2b9d7d69145691c62757303d0c9df6df
z3234da303a6c7239ac2a71bf9de7f37a2a4cad8dd6329065cef32a1af60b1446cacbc73b762036
zeb02d1d78f5c60df2ae08ec01e25efc03e2e7ba27f326bcb15301dd2b05f1ea350797c199c9b3f
z50858f494cfac9c4c8488bf3feaf33682e90d5382ff610d82261e54c8e8bb0fdf4341626b354cf
zd0340cd8e3712d72cb98e31817b4311daf9b5693ed45d0d9551f1631b7770f62b5468204edaf44
z076111f86b15c56a60d9151535edc19fa7d76fa378f83fdcd78bdfb033ba518a812befa787de14
z68cf749ce4765181526a180baa182960ab60488aaee69a6970f93ebb08369c414b87fd55cc3748
z0289311b2a05c1097d90f0a1863a7024110b84b260319d5f9343a46789aa3a91d6c78c99c5e456
z790ba35b7eeab7e76f691ee9d99ac121e42182fc21a3ebd2926d9193f4f6640fe74f9969322a76
z183021eef4d31ad1417944fa2541f7f0a7c2ee5240039352735d0d5f75aa300ecc7437cb7511a1
z7a855143a08def3f10342da3c88ee9a20a37dbbe4786a212c63b3e41edddd130bf6a7b28eb582c
zdc962f013fcac58c531127b7954e15b5f56a255a63f67ad053c1b025b54852f5516ec2bc6f7691
z68b425f26c5372397658fae86b36ecaf28029f67e5f5f17a651d920c47e628f298d95cabddaf86
z9bf6222c6828cb6cc500d8fbd7bea4ae280f61cc2bcc834aae6bb8ea2fc1521e820cec13038b86
z2fe1adfefa9bbabd97ca692d46154f2c49187daf9709d418b5557844416c66db33939fd9c10bfb
z82b9a85f7952f7eb3443bf5d2c99a2036aa3c4400c1c2e501e53dcc2557c494c38d9a29209b418
z3ab22e8d0f5a5175ff063a497a90d85cf6ef5195b6c02076634805809734e661cbaef425103c27
z2c0908aa1467041758a4f3d3f4c12003a1aac84262f29a6ec00f455a51805d2b956b6b1414ced4
za2ffa5b5fa5ac8b37eb7ed08a8a270416196162ed35e492bc47dbbb01a9288df761dc89a17e34a
z01361e675b01b6bed1e90c7c19550de0a68b3a575bf5b1b2d0e9ff8fbc1b9df81f3da4d7d7b6be
z35b267c77d37a6e776fc205e657762b98c2e2dfd2802ebd1efa00b3523433a7c54a4df753c08a6
z1a13961c20d95ac9a980fdeea5eb8d31130bee253ccf2f44acd97bdff6cde475e3074c30f90c9f
z215c3f81c7f7273f52fc2bdab32b3604c09dab2f4c14de5a19563f6e52e53ebd92659f5a0c7343
ze7a538a550c2324a843825886450f5a1796c683ded76de99acb4734dc3cee28e192fd807f8e5d5
z19b30e2c76749228066b57934c298aee38e9452c05d2f13849e14615fe2e2d3c44e2449582f4db
z37d0aa864dc2b31c9af751f592d99e0285967f2f72fe1c2ee1cbafc0190e8fe6957fd6142577e9
z77755d0115cda79760d439db8f9b0f129f2435c168ed8e0ccf66ff9a2a9e5aa09d817fa7edcb0c
zee1016e2d71305ef5158ffcb9a515108ab85b3997c08fd64cb254ce4af242d7f7f85eba0909e42
zd1b747fd22f499ec97b37532598179d80e0e4d52175e846cbfec2fa7fc050600d0941314d76cc0
zb4afcdfe81dd5789f897d764531c84dda1c3062c9f0374ca54ef9b1980a2ad9dca242883b5ac33
zeacb39be6a7470bee048153bf7be383d6760eee96b4bff279ac6e157f6c40066fa214bc870db48
z47d34ccee33a5019115025a96e6388ddd3e866cb3729b5e0896f293a4c31c70690c83cba0d839e
z2ed472776d2a6868d2a5b021be2bc6933661cb59ad51ce34b8b7b15e449fb551bdeb16e54e44f8
zaca6489b87c114ad0159ed53a1dfe7b1bfa0ce171ef9c12b9ec3a6d5c90c04225ef7b4c58112ba
zf36d9c168f1d43c3975746d477ffa8db8434309ff8a199e7b331cf09f2814d6fd44f4f88a778ea
z9dd7a1ff28459e389d2a27bca7d49c84ff98caba3703ee725730ee8ad511f235f097e4d89f330f
z292453dbc98c45b265e9eac0ad9a13e9ad52368decf092461403731301c49c12785a3ce5245b41
zb905d06522f794ce76db7f18891dbb791f195c3ac3cbdb8fd6fb4721fdfbadfc341ce79c66da6a
z04f09b25d655ccf721af2b21b5b665cf9985287af6d01aea9fa457edab2e0c360ccb951f3d280c
z74d7ce33cf015c59c41236cc4f5392034d9a04d66e39fc0c9f5398af799220e3b6edb26754cbc3
z44bec68b7f1d17ea79188d4327b03e31ff4093ca1f0e9d6efd62420ebb4c6673af644f23ac448f
z7d416c423c51a30736d42ecd0e6019fb72f48ce96d7890ac7afefff6b7caa04505ad20bf305059
zfaa79f778ae51748f05c3f6ea7cfbd6024ef96c77c7ee81582bbe6124b18722ed82264b9acdd68
z784cea81561172c0eb644f7e7278506d7edf65c42e1950a0dc062da2124a4bf59981423713f04f
zec621497154a38b53095911de06aa50a814d7ea12d42b3ee234797184345c3507e8fd44e328abe
z0f9a1b37dbdc2c1030b0dc88bccc1d2bf37f0ddd4728ca6bbf394e7190e48adba794836d2d3889
z00449d8d7902bf8d7902961a1362cca36365bbf55a7f7fde3a2a9528506eff9e0244da1230dd6c
z55e787868b2d35bba33515f36cfc7cd3afccc00eee432c76b4674425525a4fcf61304a971ba99d
z0ad550b4c42f826eaed5e33b30f00bc64231e1229d77c6b2420e1a19fb04fa17edb8451f99d988
z4a21d1a39fdf4f91cf872d665c244775c5a263b02f1110688989c45a1c93164373d061ae05cc64
z72e01ae14b958dc8105b1f8dfd3e046d87535a5a4dfb5fcb82a0105491bd81be701600d27c11ea
z61a0f4a16546ad6e97fbf5c394ded4e3eb5936e7686c34e6922c06013d7f5e67bcf00a08ecf8c3
z7df32c847da75d0580005bcf9f9912117be616af7694fa50017285e6cb7ac75e42eed139acace2
z3d5651ca02e9f8223820ef04071c3bb3fb8ba8e8b505c3f7c314c2a6c9a4944856a2ae7fccefbb
zb740711e31f57218d8b788a513cf4022393d0f0ec1d49698a4571393caa6ac55caef9702bd8522
zcd2f111423c45aa37b498cd505a8f1256a0ab4ba565152fc6798acad0474d19f1aad38188bd8b1
zc158e4b64e4b79fff89a47a5fd2b94ca0dca592b7b94b80290993ede8c2b7756e3edd8d620e49c
z547a03c7c08dacfed6a5e5a3f356abe4959b7dde774a5a03f4442a02c7b87f7dcfb28ab5514e5c
z5030e5d9bf5d2b4ccd32e5a0f180283d6d4cb117f94bf4874007ed83f8b4e163ce9902da549d91
z5c1611c4d9c87330a7f34f484f47fe1c4eb2cb436a799decc6bbf8ede237ec6553897fbede3645
zcb7f5d417d80751370c1f09b46402c933644662a7f0be0e30c7502b52282993f6d2b807fe93e74
zd59f42568f5f9ed82866df0521e752c26e61fce25250280ac9a6302e7904cd3f85c84513b178f1
zafb32eed224dc18a3e9e1badac417b1e871c5baa2121adba64a847bc48d05ee0b2390a8a362aae
z26b49ec65ceaf3d96151a324a99ad310da3cf9c9c9ebbd4fc6bd072b0e8820861c030685b81bdb
z3ad4ab1394986b7f9cec0a9a4deaff02b9a65dd9310b64545c4bd9d9127ed39404334b8e9bdec7
z43509dd89a57bf3572839bbce9d95e8cbbf97c3b6f6749c6a6afc82e3e9cc07bf57c6d2cdbaa7b
z0bb17cef497313f95ef80ce65b16ae6ea0b32538f9d1bb0e30c95f7b7ee7e51148c201cbd81354
z52ac88e14db4c9d54377ed7e5068139b8fe5f069ee7a577ce83b5a850c9161d67bca03aea362c1
z8630519853fd08dfa5e669cf6138a7cab64414e4911454bd07888dd343940469981c9693df0089
z31550e639adc37ec2ab740b8e15b613870580059582e5430efc8430a695f228f82329f215301a8
zc90fab368ba1c4b98bebf8034c789a6c4b874ba5049e31bcc6e295430f4224f69dd653cf36d360
zb811d3ad2df222ddf3067d65ff79ea390f4828b07a0c862451c0a5e581fe36f97b06711f25a417
z3b1e35e47cae2bb5ded338975c7c7752e99ba8e974bd5fd0cbc5a7ffc6fe217d29fc24706d0e99
z67f17f100b281e6a8c7b97e80d36f1f353e8e99a649862f38fbd2bc880d9b7a139b27c73896757
z779c2df205bbcec6cd7373ba2c82d3ad2b96d00a8b37e2ced1ed2e5c0ce5c4253d392fddc15de9
zebf226c8db2965d2ed151e1dcf92e9b3beb7138ad95de202b9e9d541e9ca15c0ccf61e385fa8f9
z6897d5dbe93c55d1bbbd6f4a0fee24801f0b39b8df4a3998941c78f5022992093d26eb42d07b6f
z7a999ed04498d6fda5c6af30a97154c5070be2e995f69a652e62ef4f03c2bae6c03cb3f3533e9e
ze33cfee416f63b2475dadeff81424852f821e887d7e111eead6d18fd9e839e22a729a7fa537d8c
z7c1a0611033074ccc993070d1fd59562ace15a1fc832f96913d26bea40b1fb6fe6cc47f52e10fc
z011ed9e879673116e93cb9b4b11093895ec4a5102d201b6e518d61b02f4a779dca439cdbbb1262
z9209e1fc2046b032b94d2eb6c250ed5cf5cd0abf784c31de8bd20dcba14d606289ce394e8c726a
z1a9241b3041d224dc37ed633f8884c026b33d6684c78cd1df3a8f351ed7c10cea766c0ff562073
z53b7eb7ea09d66608c4ed2ca021b44b077930ea241d48947f58b5782083c60258d17dfbeefacb6
z13dd6936d9d2609d419a1bba485065481cfd6a1cd9e3d5c197a5ef52cda4d53c1334168dd19704
zed683de959e79b09d7f8d59b89bdbaa2aef44ab9e8175a28cc6cbf8bb52b856d18051cb8be01de
z13cafef4801483391469bdca2c42bbc923fbf5bd2d040d48ae3dab10c513da4cde7f39f34dcee7
zb040e51a7023fc4c1198727d003688893613b36a561e17bcb362a99b850deab6367db2b1634240
ze808061654c742d95cbb4d0cb8cd5861e88671c92b49a2c613a8eacb87da413ab921b98d791b78
z7ca701d047b5de25e61c6f46a3d0f51307576cd836d2235b96b2f599b6432b2c08e234e14c1729
ze934efd822761a068ab83792264270c9d9aae59baa0ebab39389f842c12aa9bd2c49ad8f3b6ae3
ze177dae20b33526c1ce1e99c7508e9d8a045f4067e710022cc5b823b04bc76ac411a6b5f8ed5b4
z8f938633ec01bf55ab8e87743d451ff6d838a84b8358c5d64471d2a0791aaae2cc70f5dcd89420
z893594a1087fbcdc193bc736518a97062c710d93386922bc1fc2fad5e2617d359aa35333f40452
zccc8093caa90d8763fa5b29f0451dad58bf55b1181017ac3f82941cfc1060de8f6d53afe4dea58
z81bf503ebcd65d3240ce76415940a49fb2d69aa0e170444827c1dd54c225ecf6225a223748881a
z243ff74b7c0abb970eb42315994f8fb44fa2b7da262e1eff24ede4275d71c831363a62e3121cd7
z5e88b8cda933cae9c95aca2f020555fce75b82f38f31093281dc5fd062dfcf812f628dfa4a6a8c
z8249646b1ccd8e5efc5acb595255fba3f48ddb261a63bb519450e04c250ac8cdae451f395b3f3b
z20ec48b4680a2d1c6a0e0256165c67e79e47eaed328e7ed40ebb957e05492a0f449576997d57f8
zd5908fe18077764dfd35735fadd84fa40525721ca87d71dc884de0f1d81516173785daed278f8b
z1fe39f35cd7b172a382d39e1408e045c36683c46d5d0305d5b711a8cd5c97c555969f121985792
z8ec422c6f79748b67949383e7800e64702db9384de75df5dd24a3bec0c30649c40d69b2779b95f
z11bebcd1bd6b4cf6de6cddbab779bf1174f41a92485a6b9eb8e509161bf999eb9f5d65a44ba3c7
z669398bfe4c48fdd4175e360943e2df592817dacd6b1d17bcfe4937b3dcce0553b8506aff032dd
z7fdb265b15b56aa8c85eba3fe6dba2aca546d3ae408c0203276ec6e4b6c39fb77f9cc910db1ca6
z179cc3d2602b71728743a2e9df634ff6309eb65c4c3d410245e7c8000669216988387b519b9236
z8943fcf8341a6974f28b39308a31a6c4653638cd1eaa3f887432853db3cbaa85ad5ef3f5762498
z0abef53ad84b3cf92487857780143553dff0583c0713ec113c28bb6272977399c8e4ec6b87e256
z315f0ae63b8e74727a7338901783cb0705c45ed7097ecf0b66e76cc8c4ea09b047ed6639644169
z68465bb138302f3b8c90efc73ac2090bb7879de0f6ec077f0e096bdfbe80885dac7a85746c2846
zbe61ec50dd23f3d4656bdbf0c18a532b08c264855a0437360c64b0e06631f7a7c18509f937cb31
z5d935e65af817f2dff1e479410505d1ecf2186a279840af09f8e249ce3dd060654a14fb5155d54
z9acedf500ff2fdf579cec106769e26b038f51e5e7ca71831879386d4ac44b0a0fa50653b0f08d7
z7dff86c3180e35fa451d49d5ba0f03b79a9c6066d1c6a00f419357eb61c62599abebc7410c7ae9
z28c945ad7b41f7578a5a5709ebf047eee35ca3158940df07127f71d06315057546339b0e34c163
z9ae8392ea9ea1c220de4a2f8eb8c2ed0b8276aeab36d1f005cd9d1f3f80c2403a18733c73d28c6
z8075bba4bb42b73b65ae38eda2d6388d68089407952bcff206a00d3eeb32258ee230d92552a6f0
z60bcabe5d65693094934ea723584dbfdeee7547f5308976dd118236fb753caa705bd45b91bedca
z67e3cc70cb9a295bc0bf91bf3f8c7e7698785a9bdf1cb36596edc9bfd87b2f4ff9281ff76b83aa
z4c06895ca5d01fa36461c9e895a2220bd6cf53d25df1986d50b3de16b06d2f67e8be3f21843cdd
z1258b02a0f2ea94e9dc7def847c376aa0349e40c99e97f6fb3676592e4c2efbe34cdf575a60ccf
z98bc8c10387382f520949711c7a57b3211b4500eaddb1237767c5b9752e9ea84bf590ae688d875
z9136166a6c5aee961bcdb4579fb1f91e4203345b19080d87851a9df6af252c0a9c0b1094a760a9
z7834565a094c0548637d4f0b4cfd458839c5b58d75264de1c6b6f08cddc8c099711ef4ea147380
z464368f9de59d25330656d6cd03c5245098aaaa99efdd224bde5e6be9e099ad6619f7d39d334dc
z3a6678d459f98d09f44449783c4c013215ddd2ca626ef03b218af7552941dd41e5912e1c343477
z28becd40dff2379f77bc7cd0c51babf383ce4dbffd32b575a80ba7e696c346c48be59f11e556a1
z65dad46597f35cbdf9cba79a19fd9b75c1eb9f43643b527a9b46440ebbe186ef93a390e2e3b36f
z4d6e36e5bbc1be8800d04178b324f22c3bee4dfe88e2dcaa075cb11d3d795767711d1b988f9163
z81dfe2e264444a836fe65cc724be045da6acf33acbb8e308eacb199cbfb9e9dc85d604a3a17874
z3bf9a7ae7f3c4018b9aa17dc6e6c706830b0af201819363ae179863722bdcfaacd45c913634f6d
z171397b4431bc34e2748e41a87f80c315cb3e8260765496e756b61c0a6666e7209b9d8e43c8698
z5423d2b3f698a98833213ce758f861a393c87b3dc0eccdb24cff5442a6f91ff58339427d7475c5
zd6efdf3738437741308ff54956ab81fea590329b96f73f6fa0d18ab63a0cabb67a87abddaf2dd6
z22e7834bc19d56f1136088a80e5b5d71b1a035962608a3258a0c30cee8d939c26ea2cab0473420
z90b6bb79fc19d632d7f602965759745b0ba430eb6095ff5fa1762d1024fc07396a3e1e6dcabc72
zae5b04c4dd7c1f32003b22a03fea1d691238c6921db3b8c2a25aca24d760c0b033aaf8e27c96b6
z0d6e58f527bdc53db60f9e02e0f0337882e610e0cf95b423fe0cba006738780f76857bb2b50ba3
zc7cccab8e8fe8d14ad586e935a65b6b82bd380b5f66000ba17c311816d61187be4635035aa7fa9
z27019bb183d854ff6401ebff7c5d9ef2fa45e2eaf6d3933af7723437b4334c880084f9865e0369
z39340f8aedb93ac9fd49c061ed5cc1bb9c59cc0484c8f6114bafc31ced08a8fc0c63bc615f2c7e
z8ca511e71381130d420aa60fb918c3ee730d9a6fe2bbbc3bcba52330d7fdd95fe649d6ab5cafad
z517b6f4310e32a7129bab924a4ccc1bb979da4b6238a07b8283068df59be733360ddb00f568ee8
zb000a5e6cbb0faa23422f0881f85d6d35580b334b886b2bcc4a4deb30695ce523dd9a68ffa242e
z3cdfb4036cbeacabb39832c52603ec3f9e90e4cefd49df1a08513db1362fcb93af0603255a4dd7
z04a9c0dd23e8e063ca452a8043b7bed8e379acde2b18f1ae146e88627b8e77ba3c23f778aab208
z5393ac215afe835ae3bd5da7ba7d209b46929690727e4ebec280dd8ff83621f519470758804815
zbda3d66c24d59ec48035c89b98b0c1106963eb3269352f03b4f83a1c23f3385c2471368b02a953
z99604e38ec2f5fdc6e2a23e8b1e6ce72239762dddb925c8e2ccb565178fa01739a26af2bcec2d7
zaac1223cd87015bcf333513ec0779e4d08fcbd918245c5e4d87ef84a4c1a0d04df6ea77e7c733d
zb7f9da812b0d88a8786be9ffc7caf88a299b9bc9c080038226c731b8769392cd09f5a6cbb0ee89
z1bc47a1af06596b94520e8547d819135173da16fb2019a1b40dbff27e21b9d7a73f5bb26a15468
z45599e19f2e7a5a00945ddb9f371f1736f52c9269078b5f4ffe610c5449d659cdbe4d1e000f706
z6020a2f85b3a7926391db496cdceb19a9b3dc2b49ff3cb2c410d123d14edb4f34ab9e8610a2c77
z98ac06d626396420dcde43ca8c224498de2ec811753b54c374e73dbfba0ab50165a6aa4a4ee9eb
z7a2885675f0a10fffec674e11a0331eb5dddd29642e50365bc951b8e709db238ffd12ea6278bc7
zad8911ed88617aedc916ba5d2e888e536f70b902b7a4748b88fb9d91fd97390c9dd039874a2b23
z5466b4072397ffdbf4d3a0c8a62186bb1df1dd260302222bef69fee522fb85cbc890923f6c9dfa
z37353e505c976287c2746076b0dc31dbca196c650e653385e128f8be04d0a4e08252a86f8d6cc9
z9cb5cbd60e0ad60b016e00849971b034d9d9166d2acdcd911cff22538acd31d2a57c253444ae5b
z666df1992e06ed8b8697a645715e630e8fc1acca8b58bf965908c90b93aae4c22a823490919566
z0629e2e857fe0c7ddb8efed785fa03d6988c57399953d91562513f1dff8e08d7d29301d559fde1
z62e5f68783bc6f915f5e5bcbb24cea62854bbba0b796a5c07b0e0ba3374af26071c88813078363
z9ce9f67cd56b5d48e31fdda278f477e5fbba9a62ac70b0365790df095ef77b427baaeaf0ebe63f
z32776247d497698ce1702240ef9a56c57956841f91f7b2dbfc328db72ac558a21ca8e2af261022
z0675150b331a5671bc429e8618dd1184ae342b07d16eda029304865949cdc2cbb5de1e777a1b4e
zab7dee8f5f4dd0ebc23ad5a9eabfd27d51f30a2cfb11358173a049c7e30648140a96889734bd6a
z532b3e764a83ff3843b06d7410a5dbef5b0d3e73d9a799075566c059f83f4c2db04768eda7d96d
zf8189fe0cb03ddf8b674316f42750a888562a1f56ad2aefae8322df879ae924e881b2b88fd25ad
z4f941503dfd16598d5ed71a6382756510dc464f25f08a9bcef283c384274619cf1fcdaeee647dd
zc2084567deb3bb2ad238ea02465a183f4b98c78236287a0ab511705ede870cf0ceb3c40284d232
zc197b09ea24965403c3d8334d10627ff1f0f7ca6ab5ca114fd5cf53b43b3499d453339778c2290
z476e31098915c2d1d85b235bda8478399d42a337607233b42e5069d9168528201193ad8d8d4ce6
z86e04376b1ed271d360c6fbbddee78d2d849c33a524db9a34af94361563d2a9ccf79ba7ec74981
z53e6e0ba95cc8927eac325db0315fa2ec982d8cd663307bbfca135700c85d8b1c363712fccbc62
zbd6bdec88b7f95e46e157621d7f48029f4e297a9165b26fc7a0dcd85323c04b405d18646013926
z7013ad0d2044f92f983457a1c0822cc441d74ea4c6abf33bdd5761e39bb7ae205378b1daa151ab
zaf4168d7eafeaaf11338a31a0ac6b9c6105bf0baa003423b30f8d2ff2e01ad428705ef110d0320
z8c83751f7d62bb7e5fd74dec6c865e8af7b6759fedcba740ed626bff050d90efb938b3cedc7325
zbaae87d3d2902ff603b07226ae3692b487d268b079883788b368b46428d2f1d61e54e5897cd5ed
zb46e8951348b83f9cd4a9aaf879ed1e9050ad5c2745b1ef5e2206fddabfd0f29f5340e2c9c15db
z7c312fa1999cfb5c858b5c1a54503f38da401a890b78283f4f1ffda18d8264bfeb1443509dc793
z3259f7242c4ba1303402ea21c2f63520df4ce4f06a1af3b59745cb602383486f2019cb2c86d81b
z339f859c26fa6dd0c5b951b9325626a83f419d2e8e50caebc977b9c8a7b8e4216d60401eeb5ede
z9b130fa5beaa23da7052e0b6a0baccc1b175c25ef2c171151425c4328b71ae991b9c54674152fe
zf530d08cf629bcbc834fccd5b8c84109249a9deabc03cd249d9d8f257d9c514d74da8d65b66c28
z1a04622120d055f44db0362c0e68509d0ecd23c8cc65ad9fb80bd22f74ce3ea6baa2b70b3ce3c2
z919a817840b3b5979ca09293bbdabb823d4cf6ca14842fcd05879ad2e0caf2bb497b05ac1018a4
zdaea9c7eb187df2e87194a9452ebf8174454f160a58ac5cd339a8b042cb07577edcdec31b81a35
z28bccc96a84a086a63bff829d331efb86718d3c678b5e6081f01897b03412ffe0407ca955bcfe6
z18b77ac907490f4c154d85c035fe709e2659d7c3148a9291a92d9373ec65c7ad971fbfe0670b58
z6220c3cc7570d722ddc0ec61fa01e007b30ecd17e4290a622c7d73d33bbc78ef3f7417125c8385
zd8edcc6f89982aa1b383dd6ae5da2709ab430631866ef8c540647827110d3d8dc66d359e2d42b1
z3fdb028904625582784a08149369e2bb0b905cbfd0c4075e4521af077273141b4522fc9cd99038
z1f97a423cbebeebc09086ff84c16c52ffe0b887f83369f49398f125e86d9681e1b047b36dd226f
z1cee44891b8c920b4514d198f3e95da1561e3242de3a828dcd54aa21f55ee977852cc2bb482f53
zb52435f5df40a04f855b9bfe9c3820362ce8a3727d097f4629170e3f0c0ef4dfecb0d4bb678408
z98e2f805cb7830f74666e722f1757ecfeb107ff2c620b9a35646549fd1acd3cb25eafc03958e0d
z2cbe7bb8a49691138e580352e6478fae91c116ad74ec1746fe4025f572f671c51baaf13a646448
zaf6adfb8cd3318ebf8fd32166310b60b8984ae06164ddb7481b0ce2f061757091ef64020c405de
z569f7d9a8f9400a84d380dd08b46b68df47a3f028ea390dd4481b465c88653efeaf474119e9356
z350b82b8d5b6f17a9f4a8f2d0e462d6684f220318f210cf1511bf3313e9fc992becececb0e8517
z5f3ecb9e0ad2a4ce352dad7d17589b059f4d3d6cbfe3af8d4eedddf50798c32e68a945fa31205d
z6b390b4170e62eceef62055ab4398d65065d936e86c77dbd4ec261abe95f822c62570953fa78d0
z8386b1b36bff901fa4928aa6a8681590b18825cd94e823037beb91404cbc79b3bcbec593315094
zb3a3db5aa5261373a39b3300d3a532ba5aff5b053eef7351b2ff2d8ffab12f5266d911dfdae992
z95c7d71b0dab73f1430038110a3c0e16f78f8e92e48163819694319817837450716eb3f22c7340
zcca84a78dad47036b751ec007e07d2329ce6f52739ecf13f7f1769223aca880e8b34ead6c12ef1
z3db8e31c73bc8e640396464f7afc138c27224208fcf6db582dd6c44fb704f243523c68a92a0c2b
z1cb3a4d45cfadd03c340d12f8e5d2ea98c26084e7d2d85153a4b4e05d8160154ad72ae7c55a9e3
z005a67743547d71b53315c20e49ad3e937769a5aed7e3616fe47d629bffc864528e77e94fb58d9
za32620779a3743ba715d3d79304904b8bf6317e9402a0ae87dba89e1bd455e4ebf2883a79e313b
zb94f7aa084a2824b50f9b8fc6d08b948153aae0f0a4f615cfd8b79c880e041a07191897a587d32
zd7c84625830bf2b7263cc3aa32f8d90c7908d6b26150ce0f0aa668b5535c9d0265fb0b3ae391c7
zb7efb9aa6e730a83820148c8c9cec7f963444d32af0e8f822eb1c40f040a24096d46d02c10491a
z789c7dc5e2bb65c0f4bac011b0eb206033c9444751e9e6cd6ce7ac14552436292336bd890f8ad4
z43b780446ef51d2c4e3c61382a9f0ddceb01909a50032e761930d99965d8a49fcf1c3e9b8f32a2
zd285766daf48ccfadf66a30205e4b77852de23a344570fdf652b6458e66cd47489fdecf45b2d2c
z1408e59e929763bd198b012440371c590155b8f8636deae9dacd48675ede72a51b978796641843
z57bbef9326ccba707a4ec58264fa9745b3afcec0ee63ebd2a7307f7d3efce423d4ed6531deb809
z06e69bc98b80e3f71ed5fc342afa814834c523f7516187a46928af1b22c2b0e5224030fdd5f740
z385b3c4ca83021357ea451eebfd350a13b444fa7e82a2b8b45f69c6d2eb47bf19a8309eb1c0a4d
z7795876e16963e729d67296788dbb2191ffdfdacf65e31e889905ce0f3d9391d67624c00ec7f49
z9045530746e9fb7ca6cee62d080845f82d6a8fb4b88fb45c83f72e11361f3f91003410084bf1bd
z9ccf5d28cb6f88d82be2699b35cdfed3dd959d9ef4422954352a14a9de108865f3d1e4eabe7926
zf7ff7db69d3f5a2cc8f2a987a8eb8f0c97484efe78215603b091d11e6c78d7cf1a3bad672e9273
z753fbd0b7b2046a2d64bb3fd3fcc3810acac504d3bf312577e16a81a4461e3435309a21971a2fd
z7f5fd7ec6c1a05a7880dd9ff0b5cb0bb11f99ec3e6c0a6498c2f25c7aefec3a137cf14d359e950
zcdce1a35183ad9a035550e89d9dcefd005047054aeb84036ad9159192838f8380974e8b1c47254
z1d39179e905ff94452b555a1935fde10ec9d9b8378b8cc2bb5659bb6f1050ab6c0748cc0d6980f
zdba5ceb62905de4cdabd6f3941691a0e939dd2c6a3c3f05a012d58755c810c60a271e62f5be637
z6e4dea9effe0db3eaa1bc7c3a8fd22a041097c62f272602b0ddc39a6a55bf4d32c0369508439ef
zf42cc10c1a1890352c614806fdab71ae3315108301373244cc6e075bc46aeb7973d104b74c3468
z3d4f8ec538f48c1159c0662a760d00d3cde2beaaa5a5f2d9d6a7299e2a9eb6fbab09aada28d26c
zc853b2b1891abe534cca45a07289b9eb94f1813e6684b2f2d14d1adcc53fb4d325f9fe4f73d4d8
z674e09668a3f2f1210dcfd892fe41bd02f18c58050a800f9121ecdb1625b8e61f7f9b3b458a62d
zdce4ef7c031bc38768eb4441c8989932cedb0fb7138f62fbc182184d94e8c7035ab6f61a2c6392
z55052b9deb2e79cedb2dd7c85b03fbaae5d6238f4e2223599b63cf7c4b7f6048f89e4ae15cc1e4
zd853ac68b652236bae0843c5a2c20d50e570611f61a4c9adaaa0c1baea39e7da7b896cd8424490
z0ca7060ff67e221a091ce202d87286f22976d7b02131fa121ee9a124b12191a9e858d092f58ec7
z6110e41b5d74221a648c2a69b5622567bded0a45af45e285b8b1ed058ba6ec06f59b2216909eca
z5fa352f29e70d3909ad432f85bb5e69a63bec87ae771c6e63cb9d1b0c0f2421a15ebc9ff84a739
z604b67f4c3c4b36b0f95f2b92b29881751a1ff7f945fdfdf1abccd9108f23dbcae28ad951fc6e4
z4e9563db00dc57ffd89e9f09fd5194928f93937b5295e1c10331b3e50b36a5d5882736053b7bab
zb4072a65923dd22c979835e42393ba42ca16afe48e1ac3caeade482396cf4104212ac4de763ac7
z82902fd1a973db5bd5476bf766bfd04ed3d0aa7ca4dfed91a6b260f285b47ac9447e3f0b3a65c3
zfc8387f9663ca7ca5e4607f468205fc1fceca00c8bc68285c0ac0c27218018635a159747e22e35
z5b06e8ae36a457e69f6b9199ea7cc44fbc3f5d6863d140ae3a1e5a0607e8eefa4847b250d31f77
z9ccd117d1c19fbdeae089a54533220e1a0410ff02bdfe5b9c6e136c2e5c9233ab3099d1ceb3bc7
zc6a1ad0fa7d09e3576f10ce29610b7fedc12e56ac2ef38b01703d681a73edc0688f17180663010
za2b860ef339c2bd9010d836e5ac5f8bed44f1f7cddb4b1543561d906651960302a6f0b7b468000
z5eb2039043e56867b8a13f5e47b1b2e5e800386a5eb2971bc4e71f4f58a9d01ed7672a70c6637b
z571d33212301914329fac2c488da15dee84da7718844c0ca452a086107b39111f308a0afc22f58
zc19d34d28b7c7023a8993251c90f761f5b457bb28726fd0a01d80a72b54a3b256a7c2a61a22567
z942515a20b6da789b21478e7782dae29f26119443e23a022fdf36b6de4852ad1365cc87e56c5f7
z4718b041ac773dc527ad8bcd8c4f75130237bf599555e055b8df19215067b91a35eaefbd1df6c3
z951269c430226d606ac678bcd6f52deb5338b54ce4354673dcff2becc83da26b3bcdac2cc34c1d
zf684a2e8c378df2b259e709e087e0ac7156d48a817861c032005dbfef3898e361ba6eae259d698
z748ae275e396a0ff8d5a201e1fbacdea466f2acbcd24114c63cc48a28224b2e07d2de8c741a542
z11f21924dcf67c435875a527029631efef8b26cc44922e652567979b78fea809c124a5a5a33049
z54ab0750e227e986a4a902ccbe336e730a1ac6f7c5c0c0cfc6da25f46030b9dfe1c9fb5ff3fabe
zc33c21e983df3904eca6e86fdc53de51fd6e0970fff26ed401ec6cacfd696f080cfb21a2bfa8b0
z1668abbc961391b5825526344259f806d953f7e9069a1e4b32ce3ecc0ed0b37260a188c7645919
z4e9363ac02fb7eb11d80fd3f621cb9444c6c1bbcb5155fb98c2fc1391e974a80fc9269b08dc31e
za713d5a924531bddb72a8502b303af703a16e7274917d90e34e1b8296f6d5aa8a5c54a2b5d7473
z092bccf9bf3e4b0893578e5795d72a369d779581c941e98e798f80679919f820cb4057cc23998f
z648952d56d5aae9e4378936d88427940c7cc69776cce1dcce3b0beb13e07d0c9f01a199a7318c9
z559ff398f132ac199538e4ed725ede7b17988ead321ec050051bef06a6739dc47bd3556ff1efe9
zb0d6e05d7db2166649cd910f28cda5f61661d108e26727f3b00b0b2df18e5ed441b3f98f2aea53
z9df371574494a5756ff93e22acea6ff61f7de958c337ddffd8192046d14cb43bf071fef48eddf0
ze389441b20ac66d33713d8a606f67086c5565baa602110ac85b8cad597b43510eac3834b253fe5
z51531c8291782d505d3ac044f33a15f7098ae85efc88ef6c8dd65549a65a38add4e487b92fae5a
z7c6d9440b8c2425adc08d030e14f2a0a0ddba1396c4a0cc668d8b6867b72a26dfe1886a1704e12
zcfa4e8a9fc54a2269415c7339b7f441d30dcb5a783f8d08c0cc68a6ad2153bc4de5adb2cce83b7
z2855cde36cedb91c0fdcd3dc59aa308185806dc3b0e3e6fc1a5906f50b3461dc295f3896f4e39e
z6d7740b2234697b577ff6fdfa109ae94dd5fd58ba1f889c3366ca28b4a77fd9702f7a1027f9932
zc9fe2aa7d177da21a1a442bc938b90831677399ed443f452fc0728066f4e57933a57bbc5eae480
z1248e929ab02b060099f40c579926e67a2e1c32d330ad23d5cfeef8a9987fdef7a5bd97cc5658d
z854e1a3c69e492168294a0747157ff0c48e09775f67aa523fc70d2c00dc3186efb07d70433dc32
z48c02d57050ef4531f8bf612b3d50c03b42790594e7a1ff81337ec9bb5de63bf57875211040a56
z48116e51156880955144ce3f933d960c92cc86611261a82e10763b16c45257ebdfc17a1c303bad
zb5f47d2046b56375b76c98ba173f986f7d8ce2b13ceeda58651091123895e74a3af0ce14297d75
zd600c7331d96dc47dcc63ae669fbccb03372fc65809393bdf302051acbfe7cbade7932117ef76e
zb79ff393c4b1dfd7cd0cbf2615936c1d12eeed8082ff1a3e67f999020a5171e3ea16216b2361cb
z9dff7cd8ba094acf076de3670a24900385859a3f426a81aa15e43671fda70244fb9044b3b7239d
z618bc84cfbdc1066618373c7bbd36ce083afa985ebde76f676a89d344ead6d55d67db7452a7cfe
z4f971f037c86a3f6757ff87d167764de1ee113666ce4952e500438d200883c334ded4f1591da30
zfd328bd90dc66da76a26a8fc11d30bb9b5d0564464b6bc93e0ed490a868350d041f4b76878c42e
zaa72279c83e3ddbb1ce13578cb2d1a942cb22157a9533e0a542448b01cf936e09c416b6b7e680e
z1722929bbd538e87279149fe9efc547982bacfa951f12e12388fe335fefbdd9708b2a3c138ff7e
zf94141e17fcde38318fb5fc0bcd0379b5028101f069b30f331ba45fa0c8c3ad926905b1a151467
zbe33e9bd7370b46cd1965a1d9da31d3cefffe853417da4cfaf208457d4c7c4751585527624e095
z9af862b38bdba2e45c40edfe252c6c778072c8db44dd1d7ef5f34110cebb8c5236418965c04e57
zbdfba9297c74cefa43a76f215234e72b3a7865a629f06eba9eb62dc7c2f7813441d325e9347a91
z0baf86f2b6a52e0e12e696e041fdbcc051efafe7201472376aa60029934a8fcb9b36175707c080
z12e229c8ec4177fe15b6ee8c577fad2774740de231c870e25c7e240cc0f9ed64aeabac7063be55
zc6ed160aaff69310e6519f2285c16d86e125e06d0625209a7e24bb209452555aa22098417e0e5b
z3683a1b088cfe7e9ff7abb819f2fbacfa81b1fd90d59f30be8069e7c76f099539668dc70701755
za33353a62420cdeef1ce2f9255c2cfebcc0e11e59ea8fde7770d0b1c965e8358ebfb3ed06fb393
ze5e68a3d9e507a115ba9841006182af0448558b8821c8b89de1a393ad42423881d22b021f37990
zdd910a83a3c36913bb87c68c2747e418a7b01aca6e4693c4eee1c65f6603b2ba93228584f0b5fe
z5234cf81ccfed2f57f3d268bbd68b7285ea6382812e09da457fc1da5123a6c9d1a60c67d9bbcc6
z2035422a0f27812b64fe541dae81e68a52b3e601d20046c1230b0df8dfe4a3c451245af700d304
z046cff5863646a3f4c0e62c6e70dc0d15b273ca1dc1a0f16b2e5adf52ba970fdd3871847d10364
z5dd04466670b7562998e28f789abe54a980cad6330386860a97e0c2ab4c4aaf651c5568b2e8113
z53684df6caf446dd4480281421cf92be76cda4909e573b9a81fe908d940ca572727650e886d024
z7186e602e1180f6d08e2ddaf51b6e471d1ca22a5a2cdcbc4747f7a379dabbc295379fde59d5745
z447dd0c873c844aee26cf8754b8cb151feab0b6a987a08f1f435a152bd5d6a04330385e65c9e50
z58e8ff48e838ad4b5dc75e098adb30c4e08d77a20386f70e23bc3233dad67938d2c44088fbca33
zb3cf17b5e859f826b9edee0f108e7b4ad474c298c104747145392d342c3999ac21f68a26e927ee
za16840ed33bfe3115f19fefcf266e1e7fe19cd6b6b9fb0ca771fbc264bd607cd05a48b31287305
z0019ef3e32d3227b4758d4494aabf325cd6d057a7e88c5355249ddd2f045871f42559460384aa0
zaafa9dfdc1ce532bf8243e9c565569b0aadd2a6fd067d01b7b25587e4efe50ee5cfc03fa8cf05b
z2f400a379153288699d62452c4c56c149275219b0253c68c1b97ceb22d0a9d0b47cbbbd2d3b100
ze94b24dc47921fdb29cbfd159340b6f98ed8b40d8af789b525b05885e9a14876fd3162d9949e95
z97b7a4fb159269a1470109609c6f2eb322891ccba14b1b48b09aeea62c7ad7961368b82450818e
z20c54e95bd8c58b785eb3f0a26d7defb9a13117293a36e9cd3a42faa2d2e968ce281ec88b076b5
z7f6fe220ea5adcbd09d03883b0af95c77f3385dd434da0c9c6b6fea03fab3081f7c1e47498b5e1
z730a8345c9d4513569d7d67b18a3d2c15a91cec04bd41a2f73741dc1d9da05f121f614ee5fde84
z7a7cf97831aee9fef85308bb46b6aa995a3edd69c47f7dc3a3bf9a2921a14b4c14eaaf9acc11f6
z79dd2482c1be4e87a1994d7b40cfb9a6d2df978e63c95e0ae52f54632350e11701adf2cb5881d4
zb853a0fce84747396b7779609cf9c91ed3a3203f821e965096a48b054a24ef7de85e2c4ae44c75
z168c9f405c35d9450b57ee017873f33a8c404bd2491303bb98da822eeef397c5b8171af613a586
z0a14915af2dad77e86380f2513820e17a653116414d464d2bd2ad501dc81451caceb4e41b98f76
z4b27a2cbeee546fd2caa12782874759ee0db2d51c1855c99cf9a38c1c46630c0f60fe6602e0df2
zf68cf6b3e8b56a86d2570b905fd254ac112a10a391addffa625b40741365aa372896642615a822
z02d4cfd54bf0a1885749b11f4855fdc00ca26693bf15c871f88b7d4682cdecba81d2e5c2643e23
zad6356bbe5e4b143c10b5d627220bb394fe1039f332e02f7b867337fc3aed82b35591832b1fefc
z85fdd692e666fb5c2575bb99d7c3160578588fe9eec127952c952aeed4fca80435ad949914c109
z4e22962b9c1506486c0401b7d957b0c0008c433eef86f040d758c42e8c19c048f2c2e0b6dc2c61
z3b0734cb6f206fcb9dca1f495c031317477548b02678f0fcaad1f9a082572e7d99af8e797ec355
z8425c7b70b2f601e87b1c599bb94b12cc61c3e08f3b1502d6be9d0ca2e64a3622c935af49778b2
zd6ba4e46c9c1949ff56de95ca2e4ff884231ad57d9a2771558d7c913bcf099ce13b2503cf6a706
z83d0821e1eb415ab180bdd36fc35cf837ff4981075f418d73be35715016c59d52055d14a24d637
zd6db6acad33645ff610275767fbb9df4c918523f468af971ffee8f687b44b8f6a242eb71fdb05c
ze2495723c0f161687c3759e5f12974cf002d551418d5ffbb9e5a0d0ebcb4e9dbbe008b68522313
zadebfbf9db1987824b1bdc33d8966427ca03151b18f9a3ec41b1bd4100447f67e9026c0b5df2f3
z4670f226e76da08730480e60c939af22fd44641528b171f2ed60a54986a1653757cb334161ab6b
z8de198e030174200d8648e5cab2e9923a9ffac44b058e315c3067080cbbf75dd4ae6b16424780b
za0c0c0722bf8467754f715b9845ddd567ebd34ea4ef10d50401878dddf5a82e99aef5768baa7b8
zb2c033435ca5c6d1efdcb631a9569269046901882547a74604bace263ac7b0c9e20a0d19bb4a64
z26723d136d121c7d9a9913053e17fb702c38a66dee43133f58805d0cf47de870ddcce5858cc7c5
zaeb6b2f3c8723b203b8f0f9056f96d054e88e05540dc8458903a9baf740516eadb9773f302ec21
z2352597730cf369b323ae1b32f44d53751b1041324e7df7f0ea03fd973cdf0231251d178ad0f9e
z906d7f79faca5b2d9be3d1c1e2d2c5265b73db38232add636b5464906471881cbb9f0aca811da8
zb18b25ac850423684a029050264943cd62b0e847d151a155d5c6c928306e597ec4478223da985e
z286a2280f884ffbc1d5a79e24c509462236d2577b235972172dbc67160b4c2f484baa31b148ecb
zb704c141524dec1eb8f6b468a29d3412e494753e30a47437168467a521cd35ca676b0977bed3d1
z2c631d213e348893e0e610fcd1690bd78b86c0ffa3c16cc0245f1ea071aed44e5fde609115a2b4
zd1f35e50b892be306f2b0d9cd3d64ab95cbcb3ffebc260e6746ad74be51eb18ee72c4dd08f8bce
zd196a61b248bda32f00479f0bb94548bffda04b305692a815cbd7c8c440014e1b660c2bc561e77
ze5e7881c793b5505370224cbae2866f59a151d77d1ac6db07e073d15238ba7449758fddc404bd9
z07f7149709cbff82a7f84f6627fc3a3c6b1fc9432ed9140cad482f78790116e1726d744998516d
zf1311c2d3257000a1bbe6e69bd964cc77bc3e93eb3636553dc1b814621907633fc29ba629a50a7
z3f7287291325d917cdc24cbe4267be36bc8210b1cac03929e80b028c00e26596210e52eb73729a
zc2543a2a4685cde84c7376ca62babc49283f89450018197a19197a13a0317e4f88f75985d14bb8
zf598c97600e8832dad4dac38531b23a9d3fc4c15c230baf5e74e5638d1aeca959aead56efb005d
z8da399f9896728c7dab26c3da72517de0705e6188bacc75dfe66f44577641112c5f7dbdcc1f451
zb441a3faa873f21fbb1311ba0027b7888a5edf385e2fecda6286ba979c8b1b503fb4dc3312f083
z26abc8125ba1669c642adc915a7654bc377fa33d29565ff5213cb213992cccf84b367b63f91fab
z49eb1648844dc0754a6e9b152f654f96f1588833113b06463d04cdac59c2c4ccb5a320debbe8af
z75603d78720a54c2fee54f40c04f970b25128c67a37847690143ee569af677a004e5984e7f62f1
zec77bbf391493e1605e03ea40732671cb64045180623d47a73c96e7ba0b3a90b0bc40a31999c9b
zc9a67a8bf03ab837e56e2138213c0a4c9c2f604e252573917c86866bdd463c601535e58fe18b8b
za5fe947bfca9ff7a9b58ad072cf983037a5b6d0690444db68ee02a2d812167bc3ad0f41ae59de0
z2e6bf7fdf14ee7d3e680a451e1c2dfe4b765105363f864a144c49c760cdbcfb7e56e612c1afad6
zd7b83a7567cf82781d851f081e197278280520868bef4c189f76e5ed7552f9f6f38c543fe8da23
ze8d1a8ca23676027db904dd69b5da6e8e78afec51558576b24341f456960b9460c434481a5e0c8
zf35f666db991c78b6df52363cbabba0e464b2507ed3a2ec067ad1e97db98a6237c3661ffe8a244
z9522d39779020addf88437125b0c73ab8f0ecefc5a4c4c0c39004f096d1df3e08b58e396934573
z1ae67400da41b702ab70dea8b5f709df562a013e91fa253cfd083e13d27f86cc89972cbfdc31ef
z35fabc4baf723e9b1f301bd0f5ee19169c483e1a2da2a1cf3ff63a87129e0576ab9412f3c6869a
zca7ff3da839be49a573491a6ca0296751f6b40a9eb2ad92590478082964c5fa451887c2efe52e6
zf33d50755cbce26860bdc17f84a87a8c8764fedaf316cecd75256f5cf2d83f4eb1e9a424d1a56c
za1c19dfcc89b7c50d0fa11942187f344411239de56b0734086a3a32f3665e23a3beb9b55063244
z944b3e2eac92c764c7c7784bb654cea290ae0f86a9f9db0788c01caed54a9c06e68c6f2f69b0b0
zd95a12bc88b44bcb392fbc0e89c3302b922a82cbfd8e5280b27224d0b96a48210edd44609a3d44
z8b3029b85731061d0b34ba4a55db2c6b5ac1c9d47a4d00e32d1508aef01cd46211bb9eaf22ed0d
z9b3519e05eb39a3731d4ec968f321fe24b2bfab839772cd7a09b0adddbd378767ca4c68edf77fa
z132db4f36ecd95b20066e938c626c448d5c630d343386e6e6921360eb0a81cb7d024e245a6e7cd
z592152c93330fc433b7a1db82ef7a9b1e2902113678efb34d15c45c1ce9bb68a0cf8422f184eb8
z3733855d5ac40ed0e6d306e4374d19267ac9ba941480bc3e7a4a8099ef24172beb26d1cbc9c913
z147946a6f079fcbdcf5921dd3f1cd69d8897df737565db777ac75202ce7ef9335f612412d0d822
z9497dc5f3d77381a235e441e7fe8db680c0ba63d6d3aa544d463474fce31634bbd20624e988a63
z0814e600813870f599cff93a5bb6f4dd8463490e336bbcf3ec8092856ab09052e0e58fedc97061
zdf48d549b4833b244814904daf74588217305ed4f2d533933c885db2f9c8c07a611f61e6d22caa
z4cee9ec4d469c4a2dc90b93cf8a4e9fddff9f6e3d77fdbe56bb14854f7e10332f2639bc594977c
zd4b7e403902f9df1a21f531fbaea46d15300ade93e69b39370548467a7e99a60a8c5afd1bb3567
z415b60786764983261c9d682cad0ffd9647f7a09c2cf8d097d5b73696557dc4a1effe18b642541
zde8fbb5aef921793bbcada56384a8d8e5328ea8fe64ec6eb5fb25da738595cde3ea05056312852
zca05a74e2b838bfa23844f9bad30d07bb05fa41dcf8b949a4cc183c56d2b05908081a428c8b3ad
z60f05b99bacb6bbd5d6716ce0d364c7b6e1d1193ba277e1f651c75d75ff171253b977fe3f1dc46
z12b77ee4f0ecb9e8c167525416129c690dd3710ed82a314a30636b20cf8a7ddf73b80d73b2292f
z03191c07b0eca49413570eca93d3acf2bb908c48a7adc5e2b192d695bf488c45cb108b31e4e0ce
z7d9cd111565de30abc5160e1a3ec98e70d8b8653abe8f17bcabef68ae545dcba558ea4cac7eb9f
z20f433598c7fb47975490a25b493ffde9f89ddf78f1c16e498a715d48b3702f5045eeda3f867c0
z9ee6b783a9389cc5811c206e68209ad7da9b1dc497729c59e4fc20579fb3ff069bdfaf413fe10a
z2376d19b50b2c6ee9b7f0c2883d084e8bd7fd80dedacc8bc79e90b39f869ba803478857b7fd115
z2cd4a6119361a59ffaa2e1652479882d9a2c352ff531449e247a2b8c141638ce42b020679474b4
z24fec6aedccbd6c85d20888343211beb835bffc5a9a1a2c518730e0a14b3bac2748e18c13f904c
zd062d61fc67a3c881ac36fee08d809b68eb02201666878af538fba7636f475527b6d141fe2a12e
z9ad02d73bc1d9dec58c50df9815b69271d959b9b7e28ac0018ea3fa5399f41773396ffca4c32bc
zfff093b95fc2b63337454fc6f32474d51a590da1ffa0e74cd2f4c0aea7424f6a76f463aca87287
z9bd223a452ac3958dc0847536a18d78097aef0a26f12394773691f4210c7c64f3c99e5dae1f9e7
zdceaca833ccf48ce8f9c83f2de978bfb42d96b5a7d2de3316bf7906782fdb557259f95aa97823c
ze8853c7fb6aca442d9ab02c1db6201901e9c81c4825807d973ce6bd9609cdbfde1ced206e0cfee
z8ddf457cd5e9cf40b70c564938e348186f86146331e3798b70128fab63dd8d6d522262f3b666ed
z9ade8772d09b1984b5e09fd2963557078382fca0895939b70fc48f967b1b5911ff18bd26f9606e
z979443172e004473da56de0c25f47f2eeffd81ffe091081e595ba788ed919e00179cd9b5950509
z85f0e601e1462ac06f36135c8f50b185cfa902bc8d649de470e4f062e48e1a31c2e59c112b3ed0
za697ab6e708a0d1e09f63b149bd7b904a1de70ba6ad06b251b8953049372b7c269a123e08e629f
z21a523eaf0705f4185b17eb976a1233b3c3ae6a8413c90a79cd9c8d61e179f9100940893b46393
z3eeae46df6a80fc5be583314b4a5a979a2a5272f322c5abe7a31e8b281c18a3b2069e75a34d49c
z5dddbd539a1de9e2a4f7f85d7256c2ac8bc502eb520f227f4f61cbc86486518014b03d1a992ef2
z047a362ca424b3fb2e5be49fdc1b7c353787cb3e4411bc70ac3230096b88a294aaebd64ce5d4b8
z6e5a3503518661f92a69c6de6739b245ad25b4472c75733f86cc4d3864d048bce3baa4952f103c
ze002daf72af7ccedfb42eec6c867411f7d598074e74da1bf1041eaba4acf7baa9226f12dee39b0
zd4adae57452b7bf1e811e97f0d3f7020de2c02470e87765ac119fb800d13cbf88abeae07c66360
z55045964d8fe2d0370b634ae0372494c7c72de364df06744f6a82c53ee4e350fc185f49542c2e8
z116e3bd87c1025290c805437911bb6d1f3dcb3934375e7e29d407614c88d6e84aa6999b9b7a2e3
z5c28928bc32debe276c52fe299f2ee0c0a85283446d8aa20c752860bb441ee306fec10d854f49e
zcd49bf5105b956133ec40c24761425234078556f63755fcdea41f8326302d84148e8bbb04dea2a
z35d55931585c66b7ada4a506effc82943bbef4110c5a0942f49fb0f9ed2432bf2f6ea879135526
z19be1d790eff7e2f3470fc3470e4f8153411a6c66c800924e9099155a44a6c69aced44b05ed1f8
z504a1cc9868fefa773e7de2f3d7bfc364cd6769e5957df4d46eb62244bfdb4e8a65cc7363d9fe4
zc392b8a4df0adbd9ead407d0e976ebc2a74a2cef0cde802541328e44a9633ca517e0351074660a
z0279270e7991e49669307cc3d8d247dd18518b66468a798c10aa5c5b8be09f8af1e9fd1af6208e
z26823e2a467c4f6adbe8a6b205f60e88149ebba374ce643bd839f9d2683d0601d2eebac2b2d866
z6690957d2cafbbee0531cdd93e44cb3cb2b2ced3f5a8e76e7077d655b2b3688ab80398a54973b2
z2a5142ee453639abafb9f4802adf75c03868410ac705d529db44a7ea57651bf453565f2ec0073d
z2a646f1bb4ed70a276fc20cbd656aa4695af51ecbaaf8cccad5a6887cdcc859710d44045e533da
z01ff47d7b6623a2f7d8e527866984ac0d600567980a1478b18d53ea4591d874bc635221a66c62d
zbd2d5e192a04d2ef2a9a3053d31b1b59a6570b89010cb77eddd149704642acf57cc26aa2f78c24
z097b2e9dfc760253607ce6df92fe63361ca73f12df162e2bbd4a2f8c21f16ccb3f58284b252128
z4393f1a1fbd06eb055253db72ad2fa36af565eb80038743f2ee640a0846888f90e453944770340
z79006a9162faeb1244902f714969efbebe8534efc9e09800c7facd2a340d2573f62122ba39241d
z1bd772e1d12a614f9d4c230ec7c6d52103e9717d5092f8206246af0fafb5761cea137a7dc0e789
z732d456e45f8a75c685a5506bc889797dde86f44ce1266ac924990a04569de1a4264bbddcfa7f9
zaa09b1b8240bdedc743c716f5bf4b950236fcf179c5f545737e17349268d60c03f444c672e5b43
z3e9ead5abb2c4c21ccb3bc2e9f254be0eed360c38ce19dbe52c495c38d0c25b5981205149cf089
z89b082bf870d9baf6278ac4ba6874cc7ffc37114d95fc0cc373318a60d349932e01624f427da7d
z6d838ab54397852d3684d54ea646dd1692b0422e41b5814238e0048dff5da17f7175430b5a018f
zcdf05caf34c966cb3e531b47862fa6739499337192ba4067283a50534ce53f0cbf0f1669250827
zf113d51b3a9c3f2f8f69e02bbced7db7626984ffeba143a37f892b562d503f9a4674eae37aea71
zd3967c694dc2b61b3f68aa67af1606243154031337ac7f95d43ac071fef647aca202eec547b41c
zab13f953e2f02d1657e989a57361a00838a429d38dd100b0c25a5c10007d8dbaf2b2b54664c731
z63eb07533570397b95e6e94d17ab6e6613214569e2a981ea15cc68b1956cc3ee5e15ac3ec74991
z1425d6d813512c2044fd5796ca60b747237d87f5809c7b23952649986839344aa408ad752841d3
z40161c7e44c32629950bdda509052abddc3e6ab10ceee6ece096e260f24f8713b875a07264ab42
z2d6be6196782ff1d3080850ef7d2b0f2ae964d930e6cea35448102fd3c18f91c23fbda0de4a109
z19442498427a4af4f4d057c32d719c83c9f601550d11cf157581c9ee363e71c64ca48f5cb1343a
z9053e6cc91e7af95d5fa84b237bc825f5ed742134bde568788456292a4f7e2645c843bea052c13
z30590be2a77a540f9c0d6149854b6f3c3385d5df1ea4ea37e3129e8ad3893f517c85c254a315ae
zbde6296664df82ad79d1f86f9068237dbfab8b07e449115b16153f867d2180d5fe50649500d9e9
z0bca2f66961790df945d30162b74430a83952d8344f83a2c7f4ef137a092824d6ba964a2407ea8
z054439b9f8aa2ef92655307beae0338b040d75b934e43107436d3966aae65015c2eb1ec413631c
z1a2fbdba8765195508fcb565e00ef13f9e424693a09a45e82d2b20de3db157044c8898223c5122
zf7ffd8ffbfe955d48a34a593054ef4275131435a01497d3fb58c8c491dcc994635a78a5c86d644
zc29e04cb1ab0a41a586cd1643573f8e9a2eed65409702b418ae7250749f7d666212b3743f8764b
z14b1f9f1ef2aebc2b2e1204f561d859be540e81b24eb8143b97050e4947713618e7c16f9a433e6
zcd1da86b3928677e773ee04deabc0e7af2548761f9eba8f6142bb3daea033639f02bd57265e197
z78531a67823b7dc7543a27d252dab6538fc6562de20c1b317458d8bc805a193c85df71c016549f
z43271941cabc95e8f3e3c4ed292ec1de0a3e8376c62777d553210d5428042845dab7ab3bdc176c
zcb34a999604ce24eff01e5166271dea7bb83f26fdc7e89e6390ef502d9288b3e8e10550740def4
zb15c543a271363006a41c306141ec141583c090f536584a02aca3755a75c2c709f8db5ccb067c6
zf5e866d90c96a03c13f7c31c482f52d4f54ae3547df67a3bc306b6020006ac86880d8efd08ac7f
z6ab1ab013fdacdf75b276f5b9d5ed749dbae88377640b2a7d5768c071f6028d8f65afa2ed610d1
z7f85699ed2f551d2bfb8dcb4013c682ce55a976078eeeee06ec74d91b17c6753f2480cfee5abdb
ze5a2cb46283a3134edc7ddb3df78ef803023fb853499e0f6d4249efba5642699e5a69147f014b8
za37c3be72295b342d8ad71efa933a49b32fa1fe7cd511f846671be44dfeeaa0a579326923cbe17
z52798105b5b5ebd01103ab7af08224dd2bebe9023b6c446e648ca3a201e640cc808aae5fa97b91
z46dfe8fdff8e77730a421d12b5419bca81ee02bc825d1b5bfa6f045942c899a0251ba255ebac62
z93d7fcbee3cdf7f8a63e1d7e5a53da871c4d6dddab9a5c4aac414c9c4727c1c6151a2fa89fb931
z20f0d74fb652e00808919c73731a6ca6aa532fbb34679b20ff0887ef7d5c2dfe5a3795fa875366
z1b5632c75b3aadb0479ab0f3202899590cf44a0e94b5eaf499f72f6b6e29124d1578e275248f46
zf67009c0c441e31d0ee2696912646f2d8f72f6f8f0dfbf1d6bbe401b7ee96c63ef7e285cd9b743
zcfe6da498f34dda8e9d6ac6c9e580abeb9e10e711a225a229e5983cd243d2fcc72ea82a38416bf
ze3e1e963c7610d028fcb272cdcde77655dfd3659c8a542bc1bdb65776acaf59156eebe3a2c59ce
zb0d9d3928c8c8be95a0b438e6c5770d7e87f164ada2fb6900e3264dc6be12aaa47c158721140b1
z5bd6e370342d85fbdd1e2d28567ac196c5f9a0dab2f5fc9676e12e7b5326c0641f29b59f5da54f
z50cefcb56d01a6069a6c37c8877b3e0fe8fdccf475fc8c15fbf6ad84a965d778923cac1f632ea8
z0a0b361153162b7af6eeb260675a82dce066e6bbb9cd907b5aaaed2989738ec0a70bfed4277603
z522b1f1d77c083677994fe57dedfbdd91ee81d44f1598ac98d1d1e153d36d5426e16ff413f4326
z9f7d6ac9651438b018961d28fe14ea40a987f7106eb6902219abc2fe964acbb9ab418a1f85537a
z4fc85ed6f22a604ef13e13fb15fdb674180dd859aaa69bb45bf1f9d359b2dbaae5fb1741a90310
zc9a6b90d0b31c57033acd6eabda42a7134bf6b4515545cf9f98c2359b0c32cee5c0327c5c679a1
zf56d0f0b26f1bfcd604330ab7107beb4f4568d88ebcfc3893a796769689ede3496821cba36b007
zb1aa5f8a4df24312812a9a74d87a01decf87b1db9a9d1798a9f210d9302bdd50f5c75dbee5fc2d
zf803d4061707813af73bdd62881547ff8ae75b03b83fb5de12ce57ffb511247e4803a40c60dcee
z14d518e337a20b45070dc4caa89c6266260e1a8c56177160ca303b95f39bfc4fe8ca49c0f1d346
zc823b423d62dd7e7cba5b7c605fe097fff77ebb491b75cfacb13930e97bf0dbec9550e904c0ac9
zc5438cb243b3784cda77087483fabe6c375de44d71e3350aafb02d92030c0bccd0c57937b6fe3d
z3800d94401a24f02c7da19f081b200c6385ad85647f54d764a1ae51f4f9e86ddd2ad4639ff4f31
z12caf604a2a50bb3667ca03ef6b409599e0c8ddc9f218225fa1f8c33d12708ee5c1b78e6b74eab
z56c5d61b5d7156b6893b250aa3e582c437af192e5c212e34663320dc25baddf5f706f83674ed52
z200a47a5d6ad0c53d44d5bfc7a1bf0732895e59e3e36de9c7f385b10c429a1f364fba747ed121a
zeaa99c39b2247e6061b18d756031c700cdc673be891b0d7a5a575651b45465d5e54073a8abd930
z4b5a0477b24da8f6da7642123030156cc7de8d7714da554165bec10cb7939b3712b1af060731e2
z9c4334c161e0c8956c9f6f7501d1ba6d7918284e79584d3ad312aa0a7f7c58e348c48585a93a8f
zbf23e839d980d490236d7bfcdd1257510b791198549f1f786fd30f7215d53bf12f163176889524
z2e41e8fcc99157d43b6f2b2193e47d2803b653cb37c393c9bf7c056b1192316b5ab5af1f65058c
zaa52b5f255fb20c11b1da944a8a41827e78f097f495dbe20b54e99d4b3b2dae2dfb5aecb654dc3
z2d2243c045d3ac66d3e195db3e104e309e475a70c106ed9073a432d406a7d0db9d75f81bfeca44
zefa083c169e0e32ec4d0f35c9b9ee88e067f4f570672a6b992851df992e2f2876050ef52d82bce
z46a4dca313708f17e2f142c34b7c266a122b8642741f9a9b208ccddb9027e3019752ad84fefbab
z0a660dabdda53b7e37805b302fdeae9b7d0434ddc06a0bdf8e136f6a666954408885403ed71f04
z698e11592fc3f18b8136fd53a3bac2721f9ce2141a20094d803aa8646a5c9273e277df34b5f4c1
z691ae84aa14e5152c86b598a53a59b06e46eb79f8ca8ac395cbb113f1de12f32ad358f4f54a546
zee5573149c9b0b5bbabf8288b899b1083099e85c63251b39b76cf5f58f41db22017c88de8b9a17
zf5c6d3daa509661d51b94162270f74043225a5d3cd9e65d99a230f9ae2ec9595699602f3f0871c
zcaf2e1ce5f14597910cd38dbcd9ebe0cb07be46f87fb3a906303d14ad06f244c6a2855bb463d7e
z777e8b9bfe40a65f485aae02e060150bb44c90b12242deb084242961ae2d94dd3a8abf49bf0cbb
z087c06de40cbbae58cfe57484e49595fa2439bfb737d5a1ce8230a52f7e739647110b6728c4a2c
z138ceb16e706c0cdf15bfefa67cedfa63615f91fa8530fa1b2dd547927964dc4ebbd135da9a831
za5048bb58df8c36fdf16b1d9a859b07af0d7913fdaea96839e1a1ab28f7b5ea907e972c34ef211
zfac92425bc5b4d907018ab7df09ae0c9c56c14a422af8a6a47b01bd0079380db9e53e28c5415d8
z6eb6d00b8cb553fa6347678d04c036eea2f56e0758c35ec44850545ebc9d35a5ba5db223f8bbc2
z7906620afa2b8063d0165745220500f76015cbd5aa5b70f276a42c21825e48c71955c2ebe2fcff
z053f826d6ac23e2adc9b1019b76bd1ba65cbf4b184e3d4e8298ffb73b85f3e730ee0bdd0669646
za192033c11ec07675f92af94667fda0f82771471df5d67b1b473b5f27fe57c2bf80238d0edccce
zdd8bbb0d0ac226ed1061d315d81711a44d9fb7431f3c3704c23768fbbfefa32a57875a1d43cc4e
ze82106c2bccb1882587eafb9519de7940d7d5ad3801ad7819c7c5bf256672a810769aafb9dafe8
z19cb54b205cd18eeac811b3e18c4f8f6c922cb41476de41a14a077d3f9d2deb8725b12d44331c8
z5a8c277dc30c0f76bbddc9de967910712419fba9bfccd5c5898112be780f86604a60d208ec540d
z09952f0eb03db8590241eef226a46852f5b612e25bbcaa1354ce5a3795b80c62c79146aec2487f
z6f027ea47dc811995d5199a16080060b4c691bd81017a43f6945f036ddb011ea69dc2190c838e4
z4a301c8312bdad839aba6b8cbe870bb795f5c6df1a402a65a25ac2b2e4be3676440a13265dce80
z800f0ea3077ddc0e8fbdbc67bd0f0ebf308850b6ccc98a684f102d1583bf28d54821f6aba62b28
z1a7dc82d4456454d89fb903e86919114e441c9784df224c038f5245a1270915d2afca88dade2b0
z6d09db1e541752b46cd6ab25ab46bafd6b5bd104d63cc30d4eba99b45744059d0a5e70cf21aaba
z745518df1d28ea5bd2d233bd129b6cf5091b7af9bff47926b049896ede336f8c691b8d71081052
z864c22dba044589e64aedeac07f1a281b5beaeba3bb6f6a57a6dea70f7656f6980663bc0ec3741
z473198822aebf6d9160faf46c275ed539c98a35feff516909c5bd2953ea55c2db6026152ed2992
zbda936ff7784e43415c057c7c7b9dfc0f0d59b6bd213a98fabf21c428239f93f800fcd1fb728e7
z257595c2fb690bda221a6c0f2d4eda41e8cb83dcc92bd4fff0876e339d9f38219af93aa230935b
z5a03b52a5d8de91c3293986d03a7e44691a2e9f41c41a080dfdab1bf9fed6c5e5a8ff0494bf141
z0b1003e03597efe072fd40aa0f37370e06ead62c7fb724ba82b72b12abde76fc3234f987d90f2f
zaa227edaccc2bb83d2dde1270a4886be91f88e2a2d2f934979d586ef11abb1e68e108d71c98038
zb7744eb797e425f662e24489f3f27e4ab575ce3288e17c60a96d9e0e241a539bdf7b9a984bacee
z06f4452ce9395774c4ba117d2a5b1d95b5ed25406c5c8ced0dc9bc3878e95fdfdee38db4b1008e
z0ba9d41b1453849bc21311ae1163ecb34505f704da80bada1d0ebd00543a4b8935574a4349e3c9
zbd7d84b7511e6f5cb814123d5f21d66e3929947b168edad49dc96d324c90ed5fd14034e9030c9e
zb040218f3c3f254e02e055e2c09e26d0b3752e2f5a17c24b0d17eac1dad017f91feacfd5e87834
z4090d29363f252e3e747df0ea415e1c679e2a290cc918e783121c21b5a9304a61d6c94baf8a605
z28c3f2f6fd94ce8d828e2b524a82fb441f8af5305267d5a851dbc5f1a7bc8593677b59cc6896dd
z33d0ce3c13f878f7e5ce3cd91110f0ad89b10dd6d530b528a267664331d8ec6265082b568fb1ac
z81d31748e4daeee53e9e859137a7169ad68958e0e24132161c11046a74ef8c7fde12b4736ecf0c
z98d9be002eadf5c6a398b31939592572d02963a72f0fdd8c51fbb48ccb75d3897858691b5e5e95
ze162ebd5470d3e491216ca7f47fa2932ead6a964222351b98e281b833b2024e69f54b1367ded11
zdc8a7247bf38b9502be43a0fd8e9f050f80f5647a17ec9ca34b3d7d5c3434dbb31e4115ec550e1
z29d0885ee8ad74a11902c3ae2db283a85eda5c4dafae413b5c90331f27b9938ce86ab0af8b157d
z8aa7e02a625830d4e550f14b272eaea891f43d999e628c9ff0eaba19eca6d70a8d409f7d235631
z7150de98747fdee64fc3aaa04da7508fad08d816d1e10ee22e0110f3be5a9cb127a36abd7d023a
z8c25e73dbe1822a2c31af384bde233a64fef943b05a4e7abe360b1f8003c65e4ebe937d6bda633
z2f6c1f036bbeb7cee6e19a5b90538c6919d5a937a4b80d550f4d020735bf275f88d8c0efbb0c00
z50e89043576dfd29d27eace48b44a5cea0cc936668be7f5b7f55f58af66b2c250b0789c27ca762
z3201ef3c454bb79fd050bd31e7dffbbb18efd158178ae38a61a5c7693e08f7ac812124d303e0e0
z49df8a81223bad86e6b9d521d668f3bf48fe8cb3b869fe70ab649d650aae33e4b76fe2461e0b7b
zc951d6d3bc87ffab24c2c866a5861d7d3bfcdf6ce34cecb68815d5790c913c30c6f84411b9841b
z36f558670e9bd7aa15905b3e1b1790f658899940c5e1398f685cd4c96caf3cde9b6f11d6520348
zef0eb982db34bcc1a01500df2edbd48f2b8d5f11200b00fcb1d111a1e02b1452ed78d14f28f20c
zb8255f8efce300c6a43f8be579efe2728fa7548c97a0b8e675caa4d5e0d7ea60fadd45aa144632
ze9330977fed311167913d54ee4ec301b30bfa664e728c5592bf9ef0da34370f98fc8d7299b8725
z9b3b06d9452ada571112da501ab087cdab69e3ac0fcf0b9f33fb996089533b20902a62bd1e2148
z5216e445fb915c93aab1159d1f9b7b749b549759ddad6f5e5d0b5c5291cf3e84072ba87af2ea0b
z6e0dc1b13d3cbe6a03c3836646cb8c6d707120a087df82b6d111f400e61cf3111dd2742567184a
z77b6e507840fda5532de35c5d9ac719930194e8d1d18b5bf12e73b10306ccb1765f082204f63bb
z01266dcd7d0e7ef0e25f4fdd27ac5ea4a9d212626ed4c0c87685095197f72f172eedde483e1e0c
z43f67aa41ed1360c3ce31f846013fb21675e958af21b3ba5fb197bff719447766e6be546223149
z513b7a416033dfbc5afc4ab1904b4a830d84cb3a3aabb3dd363b6ff8b525d0569e5ec716bb1079
z005d5d130d8411d89a4de86881511be98c3c4aa489f671377f9c75c009f3ae70da96e9b1090cbb
zb51d772f25c1175022d275c9fa5213b202f1220b84a28ed2c9612b110e169b49851301c94df34e
z31531b09b377b3b6331dbe1e31de96f447ecc24b5e9f4ef3d12e3c8d52896fca23959823dca2b8
z58ef9b31706f91062914b57e2163e56d92c287754b0a7e037b29739ece26771dc4a1171dfd867b
z0f15b77a7b43ccca9f9a8e56a852c3d58b6f9571d173117e6c7c5cc3f39deff8f4b410fc333901
zfd5214bf182acf3dda9f45699c647ce69a9f3a347f42943f581cf22af0bacb8ef476c362f6f69c
zdfc95ab706947d33bdf099b6a62a4b3dce3515eb082804e80bf6dbb51072a087db37fba6e60e8c
zc48580cc643b6a4ff2bf44abe558ae60bf8559869112ed0e3c64307483fef865d1e9277239bc0e
z454e730d68cc8ff3df315e4ddb9ceee299dc35a2c0a591946a756ca8339a477fdfaba4106a5eb3
z6b71479c98d8283795daf207a60ed064b9d26bee0c1c08c952130213347cdc308667bed92e7022
z78d4f5208e3bff43d5fc54770106216ccdb6d5fa355d645afd3d0325d561b1318875ccfd284624
zaf9af82789eb69ad0c98fc841c1d2552ccce32baf34b511992ae0e4e6a3f9084a9ec294d29629c
zd57e8043f318f761e455bc352e13fd6aae069c8df97bc083e306422706e088ccf0ff35e47d2c54
z193589e10f2e81f5d505c41a8702c7536435ad58f78a7da9f2e1a381f953cdd2b34969d52d1b36
z3612f8db71361e370e917842100b78bbb72dceae410649ef23cd482a1383831a925d699e2a5871
z393f6f08a598ef58e34c833db388438002db997914fa62f44e7e961e84921d054ea5126cdedbf3
z3a29831ee60824a1172e5681c297fe000233445952468b9a027842b5613ebfb31d32100783da94
z85ee9f53a5effe2e84f4efdc2f21196351119b3a105227f1d97eddee1e381f0a7fae3b77f70ae2
zde29d0c5ff58009ee6be5ecaeeb1634c9bf7aad2c8862a101ef091b599a96a81c0c0c73d0fbb37
z1e8297b9a330865578c88ae5879e3d987c61299ad6302dde0290186601cc289c57e2be0d3421e0
z5934ef77ed65629b8d4f33985cb711654e550b697279ca13503fbfdd190f79a4954452e86b7396
z47cd00e6ddd16cf1d5ff152600233dfefdc1f225f996f5fdbfb7ea752cf48a969144467d9bb20f
z401e2cbe8c4cbdc3195cb76ba176122b014d3b081136b24a810ecf93818a1d45e64261a07cfcf5
z75b7712a5abf2fe93e133c002dd86dd856269172bfa644412bc0264bac2baa96b7f46f2ee8ea5d
z2e36355f35136143dc52495fc0d11f424c5cca48a1dd785444f915a02350017fc24313723909f8
zb35d53e1d9ca6ea96f77eacdccdfc58b14911846ebf7e50c4888d7269660c8b248d4ee9d1b54a4
za148c4ae00b4341fff20dd78050d0a04d84e1da53948a6b59caebeaefba10e4fb7caae484f8ea4
z39621a415b5b63989100ffca4c6f2a9c9b6d63f1c79c91b1b67a790db598a31efbee865418dc17
z97824dff31c8ebf434338c03231ae1321a75d47bc1f420811a1d5660e010116a65c00f9d20f952
z373a58e46e72b65d38078e5dc63e93e0c5d9f8b216a56b4b8a417853f6a51c04ca5c036f549697
z1a14894462050ea0a0e1072445ca640d18dafb62ac8ab18e6a837e34af13635fb05eed80608a2d
z4b19169be07cb4b6ecfb16358f444ac0a3b1f9b547ff605fc4ade8eee9202b03c4cc614c455692
z3846416b1de13bae7d42fccf3f5c432e4656a204b72f3476f04781259ab038a33a11223ff16331
zff659ecdd2b77871b8aa8bd2e61e2810d060fa0688ec1f2603914d10467f86c080481004a651df
z9a4718fe4afa976fe1886b7fda4770733b82255caab49e4d66aa056ac57bae5e4192540e7f0f60
z46c8daa4bd30ea0dfcff9f4c986f01f70cc9d3e25911c9094a7ccebac17ff2cd6077018f7bbee7
z8454826fa1c13ce2d2eef5a5d3e08f005dfe7feeff151781aac8c1b016ac5248ec73ed1410c6ec
zfd0cb249b22f0278f9349ed54ecbbaf1cc85b15b1995f2b5349675c349318a1b62eafed6ee812c
zd472cd4509ead5427fa63d25418b3fcb0aaaec5a0f24f00829ae83fb9f567fab890b21d9fa1c8e
zdb75a2d1ed117f03f1c0bed7eb7a0c4b7bd65e250b353c9e45b80d80f9906bb07396c704d04e51
za2ef626f37d20ecd06d96b232a840b855475116df1e8b30f6b45a70b89fbd2eb43f0648e4c129b
zf5b865469341a82295358b17228ddce2b7f5ca36d782c4eb29d78591488b7e8b97fe966e46f487
zfa3cd8d3165bc1e5b38efec4cde4ebfb39a40553623e10659d081d4de0e4244712587fd2f1231c
zaa915e8c002baa5b72b7d430710233bf2231e882068d60389e50aeb2940345ad16318aeb3d0f94
z852f509cf24ee292daa531414925d510fc0054cabbde9118912d9a9b25858645df0316acfddb8b
z90c4dcec450e4b3aabce6dbbf30c711aa59898a99852fc805d6e7113dcd7639e05ed6c29f8d792
zeee535a11be4597190426da3e920fcb048a21703ddcf623a6ca33760410234ad6ea128b6f01e09
z7376868bc4412f4ce121211b929d300450e6fb1dec3981b97d2fc165af703bb5c88d637d8366ef
z076bb9d4459aaeceae6bf8943c2358f965ce5f58c225937177b6a1fe6879411325f547837cdac4
z73adf22dbe5eb7f36f872e958c515f0a1bca6633c99ec9f16070682d29d06eb0a163b3f8403843
z719a23e59612bf3cd636fbca7181dee4d051c3f9601319c97f21d201dcb216eeb50639b879b1eb
zd5eecfb92a857c61d6f58f7a9d84ca71c94963317ea49871c904fb75128443dc63fc2340ee9560
z4cd661464f545b75d65d1b74be8d383caed0bd1a2253888e2fd27b6037050c5cd3891b4b0af833
zc8569fe9d9fd27b4647b0ee7139eaaf36125d425fba20824446162e2e64c2164fab9976659866f
zd5709e0e721d4f78413775ee098756e75ba212cccfed9d5f3e9222a147a81b602409525020ed91
z71dae4e589823925252435be058165b513cdad17e3d28a1a4b5cbfbb8ea0c8f5c92bcfbd9ec4ee
z48f8a8fbc36d39dbd4cbcafd6ddb652b927cfead0323ab95036753f856bd0eaeb4458606a5abdc
z2ae2eafe47cd2e7bbbb667d1bb6bc5925adc8332df0338486611c534402e7c038093a3372b065e
z6129b0559d2c48a248417508346966c737a962dfb8a24a2fce354d64b0add50b94ac1e912cbb24
z142b13e2da8479e5a65f9f5f9313dd18a8601d3d5684b1fc7924a7a2b92f01e7d98f16dc9f00fe
z3621f6ec3d86514778ddfbc960488f23104deca7845838635605a1a170afc52de95be97ab64275
z6a5a5d5ceb8a8069df5cec9eae1540cb872c079ec182f0e250de96fc33514ee94ec371948ad3b0
z2faadf3bc77a77840e3fc548c5d367c9e5050cb91a4eaf51974b750f42d2c01e0665faf6da11ed
za4829a9022bce79fc43e0de61c8ac8ea8dbad48b4b1402f4cc6a84ef1681c3d1e81974fb023917
z9ae36ada654c76c0c2d3bdd083f919db8a8163e56a4895d4a13e3c0ef9d53ae3e8443b342f6bd8
z00aa61b7fc66d8a8cda31e56298247a79ee01e4a4c057531e72368a0c6d0beb309d9a2ff9b57b7
zccd2258bfe8c840e63922efbb4d6911b943041b0f10419e553668de993eda6385c133ff76969ab
zff3773470b3617d67e9ee9820f59d7fc150ad01a708837b7d84e325ebf673844f614f2325d0028
z3f820cec72cda33352c80f5470a70ba18168c0d9fa3278fb81284b79738ac00b1763e9fcb34905
z5bc901ac0caa73fbf1e94851f312958b4913ec9767f712e8403f2c8813b4c8355539b7d77cce71
z80b812567fd4d772062115b9155334b35983cb9e4fa5621edeb139ac57259419367f879bf549fc
zd6068ce4d26b25a0d45e77059d3c212cbadffc6ec885a8c09867185d038aa106f8a7dd19ce301b
zbdaa7ca8693613a0a43d5ef70c3d2cee01b29871ab4246e3964a0785919484aba1397108b5ffb4
z5a01655cdd0edf68846e32eea7d6327b3a3b71fd886ad4fbb2985adc8201544d10a301e48492b6
z751ba38b60e44b0bbc6a5bf4a322ef47b033e870fc0d7b8cbaf3cb853ad7643fdc29b07e5d80e4
z1ae7712fb898e3e97e5c352e5d1cde8dad425b91a3e76a7adff7ae31af0058f633b013769fb4da
z3339df7ccdac17141488ca82fd5a9071eb21c725aa69f4c562a09ec9f0352af51adc972db614d4
z53f1b61b46d84d1ddd5fb96fbf8c69dd70af4cd4c4c16a620f854780f15887a3cbc13d9fafaf1a
zd78aaf588e5acd1ca6aac08192ed75ff964a19c2a8b29edfef304c9c37b9c1f5d8a11b31ab7632
z53dedc731e6c457c3b09e4722a2f54bf28156ea4e0b705c6049184af589ce6fec86fe87d0d4440
z746012056e5279f91d55f10165be6f40d91097bb0233ab36b6636cb6d8ccf4df26f5bf2c3100b2
z3a2702d30e36f4858858c4dc748fe5f6f9edb52d8cd3ce81c33d20e3560c6402070d2f8f60951d
z170d2733368c719b667cf3cb90672e4835a6875926cd9c7f1746d50f57ad5e43c70d1f3e0605fe
z16534feb8ec41e6e84e8aaf9fe2c746558ce395d8b61e703b2e36b70e78873dac9bf072ef85433
ze61d0c3cee1d40e5c862a788fc610eb1cd731e1e70f3202d11e370a9aa5222aae647d5ed08cdd1
z268b1f40ce4a9680ad71c2565f172b95b909a1e70f0edce194d76479303850adcb9ed1e546f9c7
z7361eac70de0d5f0f0e949656102b579c8412b189c9cea4fc62b77027143848fcb12617dfd1945
z1e885a7473edd9cf4f477df84c2cc33b5153310f57bd58493e1ebd67b2f895beb55d3930b28d9a
z244587b77e0adaabf2385ed2ab8b4ddf9def50e402f74ad3eae319369c5b45c663f9302ad376e0
zaa1a9fa5efdcf36f28bf6ab30f6eb3e26bef68383d0479bf43c1d10de694b2d0c09d7895d4b8cc
z105adcab279e3ff736b1184599d49c0667ab71ffdd0da10afaea35017b5c6eb7d5f449956acd2b
ze085cc262522dd2584f8955df7ff289b350a08bb1673c8ae3caeee4a32dfe529a3ff5e64029e4c
z598ad33e669bdf12859883d504532223f0ca248e4e221217375802e018949dee5a5155fcb0029e
z3da911cb34f0eac72a4d2621b8e5ed5d6321d19ef2deeec95591db46188f21e07591a7e0d07d1d
zd82b414b29b01e78033f30d0dd7df23938acaa9ab02e9a3a34787ae954d0d284b25de8aa4c319c
z54f9ce7d1997bc4177d1b1ff18cb69bc39ca284c79896cf62afdedda820a966f00e8548b8b9b59
ze564442d891042edb7db890cbe4702df5ac483d43c770708c10c82165f47bc7bc0204212890005
z6301eb2cbc6244a649d9e189c2b01d1e471e865a625353e10b836647be8c49e3550cd8b35118da
z40d472f66f66699040715cffecb7a9da929810d76baad2c88e10f02f80c5b93ab9a99c09f41402
zae20ce3575ef2bc2f93e3ccd0f39bfb0c6aecc7de455b59851ff9d258349003947d254a1b5e4a7
z93314f007463bbb4ac2f3041b757e9eca39270ff0d21e354cd41c275e3bc808b9a96395dd6cdf3
z03e0d8002f2e4db3d0e6dd2be3b7533150ca26f6c640d07f3e0002216773e7e671a661415fec8f
zfffd3b09e26cb22deab7eabc3a4c14eb1ad8222a40e54d56f26ea50cb4eb15ea77da2b6af53d65
za19d220f078cadb56ff26cb0196fe8451c1d197f57984f64d4b26afdd09ae720d9f758e5d56b2e
zf4afea12bc256d3f5cdd0c702acf0c3d88270fac85a0fcf13e4397c51db533cf56574b4b4aaec7
z815adb00dec9ef211e2ac90e18113a72b745d24ab14e91bd0918ea2f808991ef2c8f4f740d42cf
zcd7d829dfd8ed7a35cbd33171d97e38bc7efb1acbf8c09abfa2f8017543035b5d7e94c44107ad3
z6d45c20cab5722fb3c84ba03ac7003519d43dc367f9f63236f04d57294ca59fb91570f207264a8
z94789b87cdf24f9b1a27e2d50414f76ff241560fcfaf67071207314bb348534352d39d185a2560
z8ac4b4e1077efbf6b24a5f92313f978365669c1e46bbeb2978902927314c698b24663fb71849e0
zc526255538e1a0ca83b07b59eb93b4fcfbf9a1feba79ffa79e2f39040feb00558759f373d1b7df
z1b2854f9e5b7b7d42c70dfe13566a0a8df504a53629e03f4df5d1f39e942bee3e22ff2c9de60d9
z63d04776d51ea93c57c98014b0fe6d579286ef5f72ff9a47a2cce6e29b24bd7e466994b89e6cc8
za28651461b48e9abb0803c1a07aa3dca509007be44c86f904dc1bbe249115504e5ffd4d89d4f3b
z205f23712b5838360601bd605ae431a3efcca0e2278a29c849d5f3f05761be687b05306dc28e1e
zddb689dd5b982f69117ca298aed7eabe6f2ec5cd579ab2180d20658182e660387d8adfe384d0cf
zb5b4e60afec83d3c435f17a6af4f122ecdd21a6d4216bf6c642d522f4716899d199af1ae7cf6cd
za53eaa00f0e63e5acf9986fd992da323e412828cf5ad835a0cf13d0944efc24a826b5e596f9864
z5f514e23debfd7ceb227025d8680a7f011e7ac8fda9888b020a1e058c4df08031296defe8493ec
zea79e4a068505610f15cceb2c6b570a4ddf33af2cb83ae600da081eb0487b9f361f9827e9b6e35
za2cbffd721a436e6c07c1a902fdf9fa650af6dc489ae465b7f7af143860b6a51df2068c638e7a2
z24b09f0bd208d708edaa5c231bd05a96bba5bc2e3ce7c13738865bbcdf112b5bbe8e34351229ad
z02ab46a24669c44286a5ccab372b2cedd0d43f69ee0d0b68970c8ece74b505d8256c76ba140d7e
z7b42224db3b94c6a4fb5c47f5e7a228744d4b962fec48271f59d56a8434048ad536a5b3758e0fb
zc50ecfab930343f728eb6df3a72594841bc65ddadb75d41493ffb9f5202e2e404b6a37ba25bb44
zb6a61c9de6694ece2f6941452cfd0f3527ce5f756e3f84f424a951b28e345d82f0189902c466dd
z74a2cde4240edf920b7e5d91b5ff41a2377cdda65c48c6c3783d67639162aa054a814ea85238e7
z03ea5c2477b0252e254f4cfea521c0c359e63c4504a91492eaf801d7d5b17ad25cf90f499e16db
zf0c424f57d99c72f123b807adfffd0dd34d6db834c06124eab9ab3e879da43e13c7ff3b2baa3cf
z33bc34206eaa2f4d429adb390b49d2293a040df39c637c8bf0cb8bab2d10b09b7d5c71777a4c5a
za7899d0d56c4c3022f670a99a62f1e724248233e70390f3d373194faeef329d7ef02ab9279160c
z751546ef7b12857b9d6aece6bdad985a680c3d7dea90c1ce71e0710654c1cf6cae4e9f39921d77
za2234ed004c80647a8f994244940a4f97314bb9cdbfd8b1b7f53d44470e6ae9678ec86f83bb346
za954d1ec9e6f258903a6f1165bf7528ce1459584c7e9f66b2802681e337cc0320f8a7c4e5cd825
ze993066871dd91c459b418185f4516698d98e2ff284beb4c6abf315f91da4d0d2bcbb99023fe81
z82027da8d5dec4dc5e270d216f0d384a1e7d70f6db53e92d0e953a0635a1d0c8c96fd8fb1c989f
z95f530807952972a4f9b773ebbcafb663b78e0189608d2f19eb61b837f7143155a2b8d8eaa07eb
z99fccc5b26e0bee2acef56d2bf36fc31ad9e656f3af92b99402e3686037b32696caa10d5938042
z4e3331354113cee1c8bff510c58de4b8c14fa8c614c8f0c2412fa8540f07d5b9f3f8b01da21956
zbb18fe81b469f5d565bf8d241a06d89099ee6ee610408c8b05474a80948d34db0434c639c5dfc7
zea4090b1da90e40b63aa00ff8c06d19d5eac3a9efef8e0a1e1621267f47033cc96f8cf263c1ea9
z06a0a3021bea58f0c8a401f41e6076da9457096ff9b2edad338952f9e637a5da44d5557e1a1559
z820808cfb6cf88a7512610e60eaeeb2d3cdb9d14d52b1c31e90a840edae183cad7eb5707db4bb8
z7ed29bf788da4c2bec4d47d57df28f9adbe2bd49ae95c22a7238eabbaf05925f8047c33d1e5dec
z8762e2d7821bfe610624d6d6f179d599dd5fe4347f5da2cf720d314fc7d9252146e2e1022ce0ab
za95425a4111b24a2a8e7702a7b9721dd3636098187b0949af90dfe4dd8ec66de6050b6f81ad200
za48d33e7af2eab5244f4a98339097a9e109fb244b031eb286b694ecc1f8a8b965252789bfe743f
z05e5f0044410365cc55c6d9fa36a17c64d31bf36851f5d5253216b98a457ec904a480a63921b78
z9e93c5ee31bf09da22ffd74f15141ae70fbaaba222bff2bd5c582d2c07556852b66210577aeff2
z2cd9549062b1bd98ab17cac3cfa87ffea7752223865dea49b3796301dbfe32bafe4c2bad6716e3
z79f0e51fa7a7910b95a05e10fb6183644cf9e8aa9ddd1cdac0f1878d940c89f20cce427c83030e
z58da74b81540b30bd8c839372be904f970715638d74628e52c0c41f51b56eb67eb7c995a2b431c
zf1f2c43af2f2e63643971c5782b16ecabc53d88bbe25439095f6df0e69814ca69108e22c913bcf
z8e7bbde2b484f81ff0a0ed9674e060beb748f7a8a7e7ba52671d89fdc0bf52be6292d518544cf7
z61f163861f3aa0b9c203bb20132c9ff0ccd2c0007ee5cf94eca3bfd6e72e9297d7d44a1feaca2e
z779616dcceedfb23f7b0a6fb746c53da8b6917932d324cda47cc53b3acd7ec5b39abe0dec631b1
z99c7bfac003604383a16139e6234c0491a79799a2a557434c7094c39ad9292487cc97b20c91ee9
zd6ae1538574cb74b430571686f5444d0504a0e9c7e08187e6dfb162bb81476dcf40b7879a6892e
zd60b56a03896ac7d808a7fb112a979df1d4ec807369403d3da4d9d17b0358d88ec2e33fa8faf09
ze8ea3ed1ffa4b691633f489435bedede4b970867516ef3072098c435547d482bfaef688d5f429d
z9408a9b01e05c73e811525693cb336562d3659d791a69e72ed4703fbc70d0383a3e13cc7528c5d
z6d7ca64abe7791e600690d2493f3baa77b7fd4d45712acd19df9f3fdabbcfa46d17fca35254652
z80266d008de449addd4b259aeb42d75fcb6aadc13cbfa94f5c40b3897d4cd57c180d5361245505
z6027a1ea4ba3a5ddc1ff0d311236ad196d1d4fa4a2da5d2426392b18a5c210e990f3c8719b07fe
zaee49b604ca09d02dbb586b5fc2c3111b68f8f799fb3c79d056767fd5071b5b287b08d9cd55ae7
z251e362533fddf298ccf49874970e6ec6bc56810ff386b4c4d5d4791f4a6bea33f4fd8867bd3da
zb4c786072e443a7a042253a24f08a842f173c4cf49f718e00e1be8169ad16572069d0629618863
zd6a63a293c3c08c4829dacb863042c35a89036c540de9b8cb71f887590d8a0c582394fd16676e9
z1bb6006540cb1241f3830813c38d09af56f6301d46eefc7786449f6ba44f083b43e86244547687
z2d112e11bd46c02dcc3ebcd7035c45d73531c95b9b59b1e289b69dbafdd75ca5effe25b35e170d
zd1dcc4e7b488ee3517b6e5e1f1e6da3ec89248232a060c4650923129d89070bd6a3af99976b478
zacbba68b84e7ee836ad4581144a8c3f585e4c56cd919d510d0af394cee493c5f5d2b9f52c9951c
za95d68fc9b2fda2817518dcd261965716a0c70ffc1e3642705788c0464a0e200ed12f876cd50e9
zc3e9370ea4f52b134271bb0ab5a6c05a4f60e365c9af1816392469cef756b3bd51d422c44d7a6a
z771578964df8d9b5ca467d2837973d7bbb29abd9a076c2b55133866330326c5c31bc5f58b1de5e
zbf96f208102938ec4a87e688ea4a48d3a7bdce7da5cfd87ac5a5c843df82b4d92ba9799e57511c
z989d951b1ae8cc2830401a671b5a90c49a685c57eb5d8e94fc1b5c6ac3fa9bfec080155ba212d9
za5e825562edb7647848c530da62ad6fd7c65a12a8b98a14c3277e786fe0b9e11c395f08f16ca92
z4413ef34414dda7e425a232db46edfc7e8609700c44e6795b1328fac176e8ac7b64ba5be401601
zcc147c39863cf55e9da07f356ca680b5b70eba75072f57b73d317fe493bd31846bc1a6715af235
z68004fe99d6ded64be8ba62aa1517ef699becaba6105a8a998d2fac6e6ec420eeb5e1ced223772
zdb2106c21a3c512f0579fb430875c796fbe977ef908be18f7feb6805cbd83593178dec06a08491
zbfd5cb27107d73cf4b23f8f16da6b1d3860ef8ca0cfc404c21ab0a023394fb3aca8e48761bd4ec
zb7df18026e122d3dc58fa579f3ff4f75d17bb99a9d5bf028a785c8c475d220d53c7bef6e32baa7
z55d43a113dea1e101b96ffa0e4cac4752aac79abeb25e4cb02c8ec19a9bf66e60b7ad1d69ce58f
z097f570e665da8703ed676fac66e3e9a033c64113570b059dcf2e63748e4ed948c03d23b355da8
z65aeba4a0c7d690bf836c88a540f4394e90d24792084d04120217dc89d600ed05b4931b999be8b
z7fbbe929684f35b0bb162f830a2253227bf12e181e0a828f676d9d5ec61dd753484b46229ff094
zdb4d1a143b8d58cd85d04d923e24152e8f07ee091dffacf672565a33ed0b31db6d705e173c451c
z730363e6692f41d9c9e765e28e067e0e610958b62e5951344fe5e6336aa2bc0456fb57f7e46a75
zf8f140c705c49333e903f4a1609fd432d401c404fe4dfac83da57c3b571dd9aacf786eb3c2dd4c
z229e18d67b876b9c38938688df7b1c5267e53e2e0b53b83b9e1406b1a53ef73383c6356dfa9be7
zd379f56e12fe1defe9ffb6393c696e02a83bf02696469a41b6a00a11c41f9775b5a93531e84160
ze8f0ce4d5551e38e368c3c9cb94a045943e8af611c7a084de95c767b43ad1a82c83d05449bf52c
zdf80208ceb7a03c81c23060c220229bfcfe4f9d85f2b554f76f879256feb5b7d0af9b66faca520
zab394532f26baef4cd40df50ee8e5fcdcd6077fb7cf218f46e1a0d9595d2a9d4cbcf8e10aa2d1e
z2afc5ee6e06245d5795c8f89e99b6f733de19c5bd909496060f094f0d7b0eaa55f7f149d4ce19e
z6c7607c825a83a34698d17406b976ff763b1c0a1df70f7394edd54d2348a6cd1b62e2235727e54
zf928abb1fbf8ab9284d48373e094562771fd6adc61753b768d8e9202f7f1b6dc077f1860d70d60
zef09139955c9c56f652324f2885eafa046e2bc2584a8ac744b7fb4d4255ff306834457bba0de05
z0f2dc8a7f1498637eb2aad4d4f54d3c36d6a79de39f59fdb0dc579653f93fe29e78ef2d153f4aa
z4387d174185d86fa75fb075c98242e97cab235c25b5bd9e2e743565bd039f09e3fa77047890829
z47b4958de0076c2eeac9f852510714ae268321457f95c4b4a833a53a5b12f8ba5c1fcf486ddbc6
z2ad3ededcc870759e67cc51fb4c1f483c238f11f9b90353b663cf959a7702b49c10d8b88cb5d16
z30645f9edec62c3631ab9ad8d645162d14cc20083ac889231eb39bd7b41ddfb7b83833956c8585
zb92a020bcbaf09a44855e82696bd1fb9f6dfd78f7e870938cd8519d50c22053963ba2e0fdfb599
z96ed8f06082ff5f6f80877b287fe1f2e3e213eefb72cfc8dda0183cf76135cf5d4ad8d1866f235
z91103a097425a6c6b8aa6ca51c9f3e832933e23028f881fa8992a8bbc7a876270061b98a7ad8d6
zce48727b96165a524eec219d37a09137a1d0aff4f9a5bd543ebded5ccf44941bb9411c05b94157
z5be6add021d5123616ffc2fb66359314d4ba31148f8327b0909848012f4ba837ed5ca705b09b25
z19db9f3d20fb8aeec3cbcb1b685c6d556e1eff030fbebfc97d83e791f08fd64b627cc2f7cd99cd
z530841452aa32550663890f97b48581a2a38a1c0d849b5fa7c97f4edc84c7ca0bfa70c03fc3a69
z53ff8a9494c509900f67beb1d1b95f68b0964bb339c4fce3011b227db6a20e9a1237a6605e8a58
z70fa03fccb1c9c777bcca9c3de158e4364ce3fea67803193e6b0114b51ab8352711e2d39f7375f
zb37743e845393d103dac64104924893aa89050aa384d784ee794d946a033b2f8159c2684d81bde
z13f4149d635e9a0d2116861384cb6ed2e9adddcafd0129954a74905cb1718eed737764414ee28f
z68dfa69f026aae6e505ee58279e55749f858df0579b4fd75ed07092827b7a243ec63320a490f70
zf789c571b90500c07eb49278216f599572ec5784561f49a2219f88db9bd9f130dc9ae1b7c6c4b0
z6c5547d77d0aeb606c21ffca98d0a3e440b0b5681d1e8b1770a9c1188a77470a05d46bb1ee5620
z281a0027adb9f2f6e5d73e2657df86f40dd2649431ce30e9b6572acac66fe17d8525f14c725745
z678f390581593bfc5ba206ef723745d3f76dfb6f1f74bc4d080f9ae9f27bef7eeb9c00191c9fd3
z7bedfbad69afe2b443ef46d967e7fc124743911a415a4ace522f64f731103d1ae89361748ac09b
z42621c39d16f4fb06ab18e9f9899f4354b56c7caaf6cd643dae2765956cc71121e4058d14e4864
zaba67b1c2a5a1ca9a572031f37bae64553862bbcddd0dd57a3674ae492725257d420ede4fd9bc0
z0c1e05ac38835f0bf0253561826d8458c4571608bbfaf3c4d5227af6ed797975433079caeff444
zb1a542aa15ea709ddbe449f51c03abce53517cd0800a5671124c71d269e77a04a75e5e1d751d86
z0da90cbd5699d6bffa19e6ade35d858d0779066312cbf0d2378d6e97d5c0a2ae4cb58f11853e86
z89beefb99e04f362081489c9a6796fefb9b1384a4d0c1da0b98863aacfb2e0653daba0ab2016d0
z1f3b9569d93e0b4eff28c6c23782b0b66b93f81bb44e466e3a10f963333fb628f2c211d04b759a
ze026a5dd701e343923622ee3a068d45d4a13191cc35362f1bd30a44b9e8f0fb1b169d1a5674387
zf3fb255e2a2effa58c41cddec98806cc340e750d6ce76221ed3e012bd06d4706caa694d94f6f0e
zc68dfc0d4f7b30d153892f5b85ccfa0f1eaa4c8b972d2dd1fb20eccc1d58fafda84ce9bd0e08cb
z6f24ad1e914be57b401a3b4459a41a62a8f9644f5ba83d8c2e2445e9bfd19d15074a5ec41f79d4
z9f9e4e17098cacdbaf16c09c7ead2f9acb6f1b9ec3d99321d7be33a0467b17a0c5820b23b3fbeb
z36f3b708c9abb0448090d656413d87edb9d0d0957b810b26c4d6cd8f883eda041f353b0b7a36d0
z8edc38ca5e3bdd692a7511a6174cce09eb3003747b47ff79b88e899cfd479bae878ccd63ef08c2
z9658f1ca7d12c8ddeff118178416c3b8d0dddcc68f78f957f7f3e2dbf3d9298d3c2af32835230d
zcfc2908d31c7f5da851ae5a5911fac9d81fd4803cfd5deee880da573549b2f77193674dacfe176
z025cfb10a4fc8f1d25d9e98f9d4aa491aa49e4684b167cef201d3df4a8a41d8ec31b1d62f034b8
z4f82dc4cf1b9f6b0df8b6620af188b47a1d1e7e8c8d42aedd2f3356dc0b8adbc323d97ad88507a
z385bc31a54e7058053bcfed2e12289ffe3ddcdf3760dd1fc5e50db4454e1c98cc04ceb911cf41a
z82d58007401a4a1d6205253e9051bc3f2bf6d3d10165659330fe42c54a9b7e78519eb0ed90ac1c
zbdc5a4dd3a0405a5acbdd07607ee642deead431070590b9cd6099f9f7edd77a031b4a04bcd6307
z1ca452b2b6442da7a01f0fa7c44987eb00851f0602f2632056a8c545696a8aa7cadc2deff3a98a
zd700ba3e1ded9680ea0776ea5f913fe8ff6707dfe0fb92504c14a66b87d49a5d36d280f31c140a
zed5cd868a2ad8243e30964ecfc86b45660956c0d83c0162e4ae099079b0c6cd73938575997e1f4
z06aba8f239c919fbd26b92113ce7fe345ef792a48a801e5835e17b984773e83792dab67cd532bf
zfb2e84865882c6783c6aa33c912f844a0487e5b84796678ad05034366a9c76ad879290515eaf0e
z42f00d3854558967919f42252ffbe075b9847293b84333087af6061825f83e42833414d2e194a8
z82dac060b330753f56671a0a4ac356acd6bae42b292c57335d8aec22b6cc007f4d2bc2b11bdeb3
zdccb1e7a7cb7ba8b386d03e56b473ba56f571aa66e97c2ffc65a986ece7a0d4ca8862270b8a6c7
z5689e09c85c33bb9bfb4ae55b89acb4751d4f36df49e9bec1ff1641893dcb68a3079412c27488b
zc3d587d013e7f2c12120f28bbc5bd82c802252b84632f6b8a67338b8af62b468f41fd4bbe70061
z7a16d912254ce786df33f452a3fe00b3bcec4b23525a1ecf5a7c5aa9d10d276779f30d4922358b
zf3f7fe63e8fd0b51ec6e6fce5e6b4ad54a3fb4b220be776790bca53d10c914db0f92425f607c00
zd43a0eebfbbc773d9ca5f1fa89c9877ea170846529439ed9664f3c2689f84f566cd62a70a7c907
z5cd8fd7df6a11a55eb467d9b928911237ef91ac0b5440f9f40edcd976de76b42a9ab501fcab6a3
z10553f7baf3cc463a147f1d442e3c27323717709f87e3ac68ffa9591996dc69fa70cbf0f6f3f67
z58376423ddc782ead7e73695591b0cf3c14751b10a7c1cb272d5fdcf92db4d39e6c21a74577dfd
z24098a8a44e7c31d443a12abfb2db2a6bffd7e1c4629e29a0c832efb714f0f2288bab1b23f3850
z266c733ae8604f6c06b32bfc0a2baee21bfbd25062c3a60c88ec43eb982c8d7a4fc11cfd001f7e
z2a2aa3565cf6bb29ed263efba0f36981089c40e8e9f4f3820f6528fdd85222b123ef2bec95d8da
ze89bb48d86e990d5d17ae591cba6a49ce2da6951e9181f53b310b3dc0662a541071a4685077e52
z7cb4c07a52e408e7bb469428e21cd38f452ce7842e7aeb0dfb0478d2ad6ae509ee750c651de589
z2c74bcb6ae8712e18c4e783dc2267ebc2b70f36cda59130843a863de6cef337909b439f3ddcf84
zd53c713249c17c05add9f51a93944c7d70923c59444fc66056877460f8ce9358a9218ed187d3ce
z0e02464ce1530205ba376bfbc681f38fe6113f2efa0be21894e1eacac401551b69c19f60e8b7d0
z583b68a58c31b2ca621be1fe971af6c62759db007a8c5349ad6ff1a45d96e9282739388b5d1cdc
z0ca81907ec6f9aef443d666e4e174087e831e17e18c39b5b83d6fafb8b1eecfb21cc88890fd8bf
zc081754023c7ca856bc6c73de732e9cfa8c100a06a69ed85c8972d8c9c192f97c5d5ac4f5eb349
z52ad7a9f16d9ec7b021491c46dd95cfc314a2fc3d57f974029988201cfa15fdd97e3b477aa288c
zc5851bb6ef5a2e825bebc520fbf1abb6f44c8e160b4e8d8213700a84a17f5f5864aad35c624874
z7f30bb67ee28d5c159fbb6b57885100a3b394bae6bc580d0ad3476e46652cf29e1c56cc2a0b72e
z4c3262a4d587ffb7a4fe253f632273a0d5c051bbdf39dce55afe1e5524cc86d323288614119609
z563125973a7e22a2e0d7b72b463838ae7bce30860a5c905a7c64241868d260184df0d9a6c4beea
z5b3bba972e8733ff1e0b816bba3e890b726cd74be1156ed1c7b991a7c60f06c838174f296e2deb
zf7f12d9017a4e8cfe39453b0239db437a12363d02ce5e136f41ba4b71a8d6b701d88121662bd7e
zb0a5739d18b1670775462128d24e1065c1bb6a2d8bbbd091c1f826b16f75d809e9cadec8ec834b
z3222cecf3b91162c3d5a3aa62b636405002468e9067a326583d33cd5bca0eef12968e7dab65689
zfade697104739e25a4c85d6a156bb7f4ff0a6be17708017c04f7dd48d00c7b13dd78edf2dc434c
z367b6c5def11688f91d3159aaba26403b8d9ec1f132771caad98a9de71195b795411f7dd501950
z1e2fd9fb9ec69aa6f59536620732b79d01c8143f5c7b35f51af98d7a908b6baf9e6dfdd6238752
z2861610c9eed7854d3e109711cc6f22aebcfd302a075dc6246738d9a5d575baaa47c6d39707545
z29ecfde28d3dcae3b0a9f14ab046651ede9d8e6933c29ab2a7ebe871d1862172aa394647037cb4
z359755cfa341d2b0eba1b39bab3d6a94593ec563563225d9d8b5324fd893ffac63366169869f67
z500da18762597b56fb9bff93746480e953e4042b9cff4d15167d8d7a5ee5825b5b35618552a526
z3834b80ace0b4adc29fb03b6c0fb74e8df360d219a5a41c7b54dfe6b6ca14f86508b03b73d35c7
z68f83e0ea49d258eef09d73e7a31d72b9895c6e034461169ad784e385436f73d806c3581adc73a
z9af6007472a9ac85fe0406ccc614e1261b03ea1600e47f7bc462d457a962c01c7c2567ce5088a5
z6948c37959754a89b0e5e7237d1633bf7cad002adaa72463df238b1436fcb5848908d9ee74baa8
z5e5df04beb2d29c82a899282f15c3c1228db0bbd1d9429c8a45ae333396aa8bfe8e9ede1ca525b
zd6d458e4bbb97125cc386b820be3100afb36853178178875530b2c5a6e57e4959d853388317051
zd4ff39647db4a458556f5b0656fa9f81af8e7d1838d6191c7410397d5ed39af5b89d999cbf6c58
zaa19c0bb7bbf1fc38f6809203b3383f8a8d1766e56909074c6d44d1a53a24d2363911c7174c2d1
zebb5b72628785e7d79f7548fd24153423b4c6e030541241fa4c98c511f3d16ff948b9516281908
z47a221ce5ca4a89aba448488c31f1f2a9eebdfdd3f62e226d01b850efcd9d621d80efb3f0517ec
zdc2126a9907b1cadd560e1fcaec4f3d502a3a95a3ba2d011bd7c5e51d7e22777eae9470862518e
z92d49e3fdf8241feee73df930f7cf74a3b77995c22ba31bf540d688980b76fffb9acb3b2ce744e
z573653d034c2550abe60cb5a37c67aae8d1ed7680bb13ba76aa203c186c700fad20106e2ff27fb
zf6dae7d02c8310b1d358b9392b87d3c2f635d6b98b1741805af6f13c7e4caf0d48da980b563717
zb9b1c6d64ee3b6087db024610bf18bffbd3e5b2404eb57ba458256838347c0cc80ba82367803cd
z54043da313816287cc69adb9bcfd022d30c7644706e28143c205f3afb7859cc4a8668f4994af53
z503740d630f7e8a127e4fe84f05a38ebe04c50db7c920641e38e2f1af10d97a77584a08ea8a477
z063ee97d17e6e00c995a63838220d014941d3b8a36366ea17ab9e5c396baebcb6d060253a4ec4f
z76a05dff9718b6efc129a5ba7f02a38683f493191151d3475c9f8a66a941b64ecf5e8c68ac8d2c
z8c16dde4ac4cf42cf55a31d745274ec4971d16a19aae23e6997038a39c6011cd246ac12ea06201
z8bb9e2237ad95dba60feea7c94272b0416f7103fc85fc5c93bc1f8d70f6ddf682fdf08c0fed1a8
zcb2d4002562c2fee484c9b2b71a7b51016e2a470e584b7d4fa124a3aae79bf7d20b66a3c482940
z92db52e42f8cec96488554550a0114026aae5d5f728dc2460b6ad188c048e60d09c5b2c90b6492
za5641b7185f0209ac89a275d613be6c347181cfbc3345bb89e8a6e1e8bdd6d3beed4954ae7196e
z55932559a926cf499f3549d0db94cec628b4d524898face1c4e9d1307bd639a09910609f89dc89
z1eeeb3af5c67a1c2689355321de0e68ee7d2d30d347ca5fe9eac9c4cd6c39feaf5b9a2f20fb4b6
z72441181b945b58e9db989c2afc83be4911a79ba1eb987019810db2399118bd0a8e25316667a07
z3d6b1d69eeaca18e2a5c342a68d61ce951e8da281e83d8d03a4f70b6e003bcfd606bb3cd4d58df
z1f4931df53061fd048bc418d3c2ab7a91381711131dbac6d1abe41880c3d4cdfa48db4dff78141
zd6f4dd0ded964eaa65a76e47dc3406fd64cea623ac86db60cf9d323e00510dcd520282bfe165b4
z6498da49b43da0fc7027f00cd4d0ee27d423b45a16304d8e63d9f4beea449a7a82850b552c6fdb
z094e57a6944d615b4b2ce2c2c8e25b7f7e40f0fb5049292bd2c871e61da5d7a6f26eb90f700b95
z5a9440ef709350df151e330ecc2268edf437f5848e2a8b8f597740826354fc04d79329cd0cf7c2
z82ace128c2a62e6987c3a8ae815dc0cda5c66525c0477d0450d8d0360a5f83e6ec26a809767cfc
z4c77850a49e5ccdbd230978862451fed2c33aaf60be0cff1f48968c5d281da913f47ad64d6dbf8
zce3b4a11315e2be8923cc6d5e5a2404cb1ca2ab53c64d121e4982429ca3c2e021a38c6e5f4e7fb
z8c1e8f53ad61c33da9a907755f4ddafc18c1e4076e103c7d8d60ee899ce89fcd26d8c9976c1802
zce8948022078dc627fbbc39b1dbb536bda107d9a9c4e83c07d4d1fb5fe9f7d0c2960912e295bae
zeeb26b486a37ffabc9d559ddab2d83439a7de2d19e8bffca7f6c330f3c9306b9e3f94bb7ed39eb
zc225bc23e4468dc3a13a1413e5ba798e3ae94bb1c6862af3cb04fb1748a7f33cb3c03110aa684a
z9fd9b9f88db8abb19d3c9b2b9b67a56f344ce647591aaa9bfb37a2085d47051e672d8b29aaf353
z0b4c4b3d07180b107ce241af7ae40a557f5e535e302987d6131a21ba6c8718405813a14c2732e0
zd9f131c4fb3c37ebb6c00580c0bf5e8b07e202474ef1ddb8c0ea529221689af87db15a91a1e848
zae44e86ae8b0bcb2ef87435b250fb0fba15b2c31e4f2c2992b0f334a8a5632aeaad1d4da4cbca3
z4c76d1ec6194feeb01777233f3b732bf6d52ab28c156b244fe89fc95d896f311cdb3c7cd9adb6f
z425cc161b728f79598cf50bd56879a1839f2e42aa2cdeb777396a853392030d8ac6a33308e5ea9
za1e4321c0beaeb981fb88bc0e189036bdf3ad084d9e18356c99ec9ec043ddf8507b73df68b6ac9
zc081c0cb75314fd8c125b90dd4058eaa5d6936dfdf9eec94e7063e01ecbeb595498c4c977e22fb
z7f48782acd25b9aef9875ee6643d596ef83e8fabd8e8c34e8be3fb0dd48fa525b5a68b5d81d645
zc783f317041286a3e4f9e1e2e9a07f402c98004155d2ddf5016174ea0d0a44b780b0b82c87fbfe
z2f2cd5210dabbef934865b204d83803fe76c5491d952c1759f8df10c77ea49eed21a456d55f01b
zfa0a87fe8d9b6296a68e9fb9b6e0340762a77a385cabffd5470f587718b347bb1ef41c16170962
zd7097f740432914068ca056e337d0567774b6198b94c2161d5f29b37122b8804f11018a2785381
z9122a9ffc1742d9e88fa22ddb0ceefbd24e58560c21148e94c0c64982e22a8dd88d667696432d0
z3739cf148814d43db08e00d6be7745f8b59a4bcb940c799a3c9501a62c14392820203584d5f3f8
zddafdf7a9ec3aa364e6847d2bf2594a88e450042e74c16ea8190b2f1386003cdc756852acf09d8
z3ae71dee0a55c3d1d65efbdb1e19b3a4b95e3edfa1489d1af89cebe956659c98815dd7cdb6744b
z7e12410040c33f851288830c03918c14257642d32dda15f8c6aeb430dc745129f8cb54775811cb
zce1019f0b0889230b49a927bb0fbe532edd5fe1650422cefbe7f0891cfafc96be8270f4796e352
z4d13c8e1accd91526a6a15e284d6f4a6763c9974cba897564fe4c59441f18d9151ab6303979a6f
zaa8cc6efe0dd8a93bafb364fd467256d3456454ecb64812252730a10c1fe868499b324611b88fd
za72ecc6d6c3d4b261cfb70757516a1455921c18ad445c89ea4f2a87eee4dbab7efc7cc7ee796ca
z1f93a7af1d864001c7498582b6044d4b80d1dc7f3459f0eccd24e5f5306b4a699e1fe4e056b988
z21a539e8d0e31dbac9b115d47b69e39862762331c9a34ddd28ee2b910a637a972aef5e26194ba1
z09740544e5558cc66c0b93f43701e0cab71bc1228fd30bf967137801ba3d3121fa00b4c7b564e6
z2f3620117a1574d092b6414bc2a05d91db61a56716f3851b57f734f79679d90f390bbbc60b2f94
za24fd4ca267b70913edc0f95836c52143ccd77e18f4677917916b4f6abd55e46626fb6e6cd8595
zbe98541a144b82760943e000cb2f715e43b205a68b62b10592aeee2e70c95ea699b9d091a32201
zedbd446915c508b0265330e5c207f6f3eb0f2346250df033fb9671b8ebf0e8c3a28f66295da06e
z7eff53050e753ed26dddbd4fd7b69383d66026fc8e1e89bc59d66df5112c5a83fe55f71127c9d1
zca917f276f4aff994c7f48cf3875c86185a6dfccb043ed81fcc75630431ce78bd75c4238aa3018
z87417d597b3cc7870e8434fb1bc5d8761361aadee4ae828dc2f26ed719238ad4e1a68cb8e8be9b
z47f5dda49bdb577dac1c66d56a86a9daffde1307f45619355499ca467aa229dc4dca723799d1f6
ze555796fa8c2dfa6162392d1d5882d307865e20bbca57cdf69ccdb5a25c817ecce36c28c2a1c86
z994ff760e4cfae3bfae3aa438936c1a70d4dc5f8f64921c87804b4a22d49b938a53e4afb7bd3f8
z827ef5714a57a5ac93bf25bcd059ad84881950555614f8bc8811c0d25a5e551404ae44c741e89b
z01e48790f70761b2f0011d0cb92b73c956510e95779e63cf265450e48960b8c6403fb15947c6f2
z5ad51e873f66a74e20102f624ccf6c2571c81f1028934d87c4733f15c26966213315b785d94f86
zaabfb15df2b46a97639db5ca042143d6bd20b6924b55f9f19c4f199d468fca6ca95edb041075e5
z32784799d5b2a85eca6024567fa25638241e5b9c9092c840a1dee0d2e38f57f259503b2f3303da
zcb75b442ed54fc804c898ecb637cfec7b56a1c9669e3d9976c751db81d5863d87300730972611c
ze4b59fc23594f175a00ca55b47e887c4329eecaf8a21a21d7d5d3ab8492d597d44969cddb89769
z656cc9352f597c00a78491380e60f21643abebdc78926b8c8dd759a020ecb328e65ccaa0004bd3
z75a3dceef5e9626023edb39d976133afbf53daa204729593a129f8f00637d78f805ebf46be0b96
z107f7cafd3ba84ffd71be7b3669f036f0b9d653e3dca6c38cba9ea5582fce72b400d1aa457cb85
z729b3f1f870630e1b402bcefb08101a8adb2ae4c76af2ff3c0dc94df0f9ab3d16557538a806e1d
z19e0a893fde712c2d489517723b3136826158c3d9cc9c3bb7e41c467f81bbc8198c1fbc397b072
z537b5fe56032bcd4da8cb5c96cb009511d8373bbf32505dbd05c6d392328bfa5715496e0ba42eb
z60617ff44dcaf97cd1800d862310f915591a6470653975b0fb96a2db83aa66b151299900379724
z89b3310c86e5f3615d3319bfe96648a01546f50f83ce119eda7d2dd06fcbf0ca3bb6c609f4bd36
z705c45ee545b7a1db898add93f166bd646c30baaf93b750751ef62e300c46b7dc5784c49d4e2aa
z0aa2ce83ace0f33257d86dc7426723bf731dae3990ad2557046c9740de1142adb87dc22ae316fb
z0a80329f745648307967360d2aff9f1334badad1061f1e041565a787279bedea1494494da91bbb
za8e986bf91aeedf0781384d45c52dac2699759445fec727ff7a2082f26505a11c02622f764f522
z206d8604b6a42d705cad766a1e8414f5a3ccecdf767b745f8562dced6e1060f6e050e46a7c08a6
zcf5801f389be516669f7e8a617cd75b25928e62c9ccb1bbd8708c79b73c25eb97b381f223d0b53
z81c93f7f5d1d3aac22bf209a6d95bfff1888f38fd6f8d20b726f0393ea322c1a71caab4f6d8e82
zf1c55136d4e0ef7bc1491de04c78b86f142ff19dfda4396616347493d3b840bc69cf8cc7c9e412
z9d86f714117972be53a5ad0c4ed328dcd291fec1b8cc436d06bda41e4d3de04def65125af6c0d9
z49dd3c7d52b318bef5dbbb1971657a1fc330b76b561a80f2c418933ff58be10a6b56f3e8639f9c
z4dbdc3084b93d5c0082a858cd3811688b882e9b3b3b0e2cc74380849a9b922a2b6e2014039d279
z19dacbe996a64fd5e9e4ac4952125e4558de25dac590918528d9c5e3fba5918b6480813456310c
z7a9aab647c6fa34110feb355e5a81ecac3cb14873f80e59a0addcb44c305889b98414145015bc8
z8e836c0ba2f81a4f2aab1558cf70ab8011de749d14558d8a18e8aed5a3d42f2d492c81618d9282
z6004f28228dc089184cbed9e3382791289f64d4dcfbdd35e1b941080a9a94f0abe4e432d3f0ca4
zd297f35305312c602c8a69c3d99dcac371fa4b090dff3d79f33333332aac77b54ef1c0439821d2
zdd9b1942ad2a6b8c34fc0829138ccf72b62614dafb12376f460308a7184e9d5630f6d57834630a
ze5153f0ff8f9927760c201f9909cb40bbaf141c362af4b36104216ab2a0f89e344069d29751d1d
zb09a4fec5b31505164f347d67b690104c197e338fe99720de12895bcb1e1ec0cf681659c41472c
z44621956ed1a503a212b05a34c463d864fe10086ee88034da36a893944c82297a316b03d02bd29
z571f6c698cc6fe441b8e6b8582d88edb524176b78eb1fe472aedcc13e86658b6f760a92964027c
za048e2269e09b76c6d3f501cab50db641732a07fbd373fa16485a12e4c278fc0429e5a04969fcb
z581df9206796c8f17814f790a4f91b5c3985c9984495bb7ffe2e152d1c276e427123ba4fe725c4
z607cb53ffefb59ac42af00079cf8ded7c012445753eb1650dfac1a101e13ae9d46812b213de8e1
z572e728611778b8d906c065e63a3e93feba373499fe96854b559cbcb59a53d4e1d1ece866a6da8
z69619faef0d9c5873c80555b2fcb62096a49c59f93d854b4f898ede9c5d081c3b5f48e6ca29f67
zf2994720791ac72512881df0770d6e244d3f4f48a53e7ad11b77feb81953b2ed766c61a74e1fbf
z738ce961d8433c1a4ad63004ade5dd5e5b1913da04e6cb026caf42ee364836e655c4c12f2c35dc
zfff5ff4c9dbdb6860c7b657a72cb5afc5af6a85eafa5cdad5a59916534ef01c8e205ee89ae5044
z00d3ada84672b7725a987b91a9803e81056b0c975da99d265d1547807ff0333806408153bbb9cc
z7acf6fea78e40ed615d5971aec177a7af93e2eb7b5204f774c9c2ae0b17e8bb6e9e0f0777a789e
z67e19fc486bf08298a88e19834af1013cd9181e187923c6103dfc376b74935050857b38fa69478
z95868eb0faa82858c61fb5de1fd0851e82b6184b146fb54b8dd86f35b77fb47139bd9b4a7d2711
z7d3c4ad60e19dbe98ce48726e7917efd32c1e16436c53d82576c7c8696f6effaf797c1bd0d8b96
z38c6a46c95dc183366838dce0eb7815ba4b4d496657deb107d6834085e3630c733d9c3fee61406
z87250fca6297083a3df1d018dc8a48acb8858f301d99267d8cd369d7bccb36958574d7ca5833e2
z76f834fb834c49a87444922867d580a66ecaa6de44a5ae9a19355ae85e0e4b07e95a7dbaafdc8a
zacfcc3dfba243a7b00a77ad9355f3ace758c1710bca0e92b2af721a9f324e361efea74abd2ee8e
ze5995aa12fce2da3d6ac35cf30ea2678f734aef04e67ca1a21ff12fe296ecaa81c131b07c8da60
zeb60bfe14a55564d9b3b7c39316e9fcebaa027734a018cdcf1b5d70c5e398f45c27cbf25e007a1
zc53f217ccc395af2475427f696f54241eea7193d27d8103b64be8ed3d17de1cf1ef736e4968645
zc58540ded5ff3e5eed3b73fdeb2c686ced50b768c8d037f4ab7f44e57d7726b58982bce3ba1991
z86dc826811b1cc4cfaaae7df16f5b1e0a12bf15be113617f8c3f554f7e301d4e7d92f78e3f7c4e
zbf1685f2864cd62cdb04e0a7ac6e6de8102ca75128c5e7f770145304b35e264895d886c374a6e3
z5c2f4d0615c7b9de7993ef8ac943d257b11c28653eeb8075ecc5325b99a03151948df1595dcea0
zd6ec5ca0bb82dc2ff8e67fd4351ebc9cc3a8e7f75f01731cb0a1c8c36cfbc66e4bd64a9a9b25fd
zebf96a79f6516bf6ed87c442f1c6a8357bedcf3f681ad968de7fa2b1bee2dbdad6919c78ff8bb0
zb867152f1a1c94fd239b2291bdbac6ad0de0eb5700db904c0d27aee6c0f6cb5815a79e86f95835
z98aeb3c3edd71852daf0e579cb8fee186a9bea2f71b25c2c07b5b58475d565a886009149b30527
z904cb394a9707ede43d15ab81679f608dfc572ba28407e58daa21c845a34a2017336efa077d658
z60277f5f0af2c4878c535b464f8aa9489a938b8e39ac847f667ce0893ef79d4b428ad463aa25cd
z2a23a3eb225fc58da69cae683d93432180eedd2dcc0d893d51e0dcca5c533fbe9fb06e1514c238
zc4fc94e8582b8efe210a44571926f34f18b825c824d8a16c3c387342f2a399ec24893118a4637b
zcaf8836d99adb164ae1244e332a335e3b68cdfbb791acd796865925ca6ced02280018abd9fcd9b
z58c6540ef0bc102bd67b87acab9e14114a5050c3055338d575265979d1314d61a7dfc0beb8fe68
zc29b2614f0624b9259a60576f1ef209dc34a41c28fa2caf982d7de25b975f4c54954d8dfef86c8
zab01e9dfd97cadd7486d315d33cd40ac027f5aa84b0f4501f6e286b32f4fa682a23f63873fa634
z68e0bc011443aa4481932272a58b23388a0ccfc0a8c18c1ee87639c7056e11dd0992e9a47a3307
zcc2d3e8f555e66810be4da85d220e1dbe8184f2515c245886bd7b90d00d129ca51c37b05db0303
z51178e739850ac20815b7ef14eced9d6397f888155e5d8d56a48a4ac74ec31fb81e2ad1baa6d99
z6cf4f00c55831538c573fc997b07a17b5faf5d64389c60ce6728592b5c341ae9f1e6efcbfea78a
z19d3c11e9c1335c93e36e64947fea609fdd759af9b3dad12d097955c6d8112b8f9c3d89481fa91
z5c43679124dbfdaff33900812bfe18888b0f874ae84c9082473f0d0cf8fc0e642f9776edb7b349
z75c188f0ab34a2334645d0493bd1fba66ca59710c868920aa9f64816f4ecbc10d10be5b124b39b
ze7f8992e7438e801158da89b5f59715366c20bcc573e07f7200dfb512279c137cee42abac6c59a
z68fa7fc089cd5510093af086a8e714a8568c72cdd97d68f95cd312983da44d0db3bc457851b049
za3485c61d22bad9e59c5f69ce23cb7a627434b7baabc468d1b1ee4be3d9f05609132472d46bb4e
zfd3aa99ab43a7d8d65dd49a2f4467f3325fe9c5656ae2f4a4d373eebc9a427d14718dbadfd2380
zf2fe940ea74dacc023fe34c94b68ed94ea142774b4ec15716e5dae3f808e9ce54e1dcc69fdb499
zb7fa06ecedd9ec6e9917b86fa41f0ed1314b12679a14f57d4de93bf5bf7f7283830881f29b7685
zbf7e232278cee3db744d55e8395bd9006026f94125add9618c10f3a0d1c08ad54aa60e87fb1bad
zc4902a924f9a67157a24dffc25bf3667c0f745b493d0f985b351df83029583bff163560d883f3e
z667bddea4d8bb861ad2443239ee446b7aa8f3e100ddebcf1d9f410e2e05f269747b3a58a73a1ff
z3a8d94e588ab5d2a2b974d28a6350067d239d779d4d815ce71666774db9f28cd9c516fe93d84ee
zfa9d263a25f39d080a29642ad58419879e2b63ce1eded0bfbeb461817bc3bf4ff9bf256a25c7ea
z28ff9f2f6a830249f27c02b42ce010b6d9d0ab46677757e2e84b511c503a0d2f88b4666df24d38
za471b2594bd14b43841522bcc086d1bd769a160786ce0309f665cb86e5ce87930f505bc279f31f
zfcf97c7ebb1660116800d1cdb1d54d56beb96350378feaceed4791f8f65f18756c633c9b483d9f
z30747fea5440982aeb4d31b0ebee86b54f0f240890685497e7a6ccc1d968ab49810d56b4ceaf37
zd7a0d08437b7afeab9eaae0d97749b8bd05f2fdbec9f31cd1102c0c5174800f7e27937148a3d5f
z720f4edf1d164057b30db28d86452717dbfda1a42e935cc8b80fa4c9a7937340da26e820c85ab9
zd10dc92cf2d25bdfa00e8ef07194c635b6eb88ea8914c1a0d4e2b39df90776862b74ffee5a9cd5
zbf639be994c96e51ecd09229ea88c17c501a3973e086fea75a8b92e05b49906b9dc2fb811bb57a
zb76f84742b3424c7c087f69b6ce47d079eefa48cbcc2cec5346c4cd199d2481c1d54671da7a2b8
zbd92c01617eb5b29c6097560a04df4cb3895857428922d738ebaf137d9b79cf5a39d2842df196b
z0552cd690d8abbf290904e584c3381d7d21aee58a875b5b55c19fe3a13aed6482a7d60e7560ca7
za3249fe6cf9dc81fee89e760d3f523d1a91450048abf8c1f95d8d0e1e74cf02e665396d0857b94
zca60e1d75514769643ab80da6537830df63d759aa908490c6514312d12e4b6892d86b2fdb8128c
ze5890c02b9cd664ea1ecca289ae283d6edd17973e5956de8dca7ac25f1e1621086da3e613f24fa
z46775533fef3c6ef2d61c62dba80c349fdb5f296b4ec6f82cc2b0b7f15cb6aa6629dfca53b56af
zd0aab335b57d2ade08b137dbaf92516767837dc4eada053d766a359f34da4b20e3d57edb090f25
z66a7e9870bc233d03d7c66a76b7fe0b6b0df983f0351b1a6247733ca6ab702df100549d5d998c0
z367ac60d5a89f0e2893603f9dde6da859ce17ea9786bdee1bb5618ba981e764f4d0c9631fd2e74
zc41f5282b5455cd11a452728d296c4fe1f12ed28baa2f412378a412504d58e49a5bbf0f5baec09
zaaa1f004f8daafc2b63644003c0106edb7883bf10d61c513c4f5f2db6549946da940767bbf419d
z7ed025b36fb31a967226dc20959c7484aa6b3b73f40c9c19b9a61f58a6b2e6d05ef4a2f20e78ea
zaaac1efe0728abeb87ca6ebeb5ba38048fdb3cd01b5b1d4443cc06b98a74cfee0a0aa167182e78
z22d21045a26cae6a8a22ef12ad8a72ad7a37ba56d02b9591848f0cd6b72a9a0bcaf41f7023abe5
z1a478900f3b45b8e6c5f46d5523757cdae6dfc021626ae27154a2d94d9956e7df3c90f4c980611
z0a16e98e64b140106a25eb1d109ee7eeb4f5275ec15278aba2b86c8d0086796f14d98968800462
zdf438bcdbe142ad394e84a1d3b7231a99f211072d67fbdcc27d770587f72b5b74568f3de2574ab
z0497346ab93ae6560d7894ad084af1508804da2a88038deaae1569d0e845bef8dc7d68046fd50d
zdf0d7edc7deb6e58d94e1249aaf34ba9d340a9fc08aba935a2c9c6918a330e7e7f00d277af99a4
zbe19561eb1357552feda626139bd4d32301419ce5d5daa6a8493482955ae220cb311f964ab4abe
zd137c7d146d5a890fb7bd09b0ae17a0f8dd81dbacf5dfd982b38f55fdb475e8c5c037d11d4cd0a
ze1e7da6df1b978cc094436d37c46041075158540068d0f02d2b0ecb6034241d856e02bdc08960c
z9a19228e5bbe0b17892146b55b4919233075e3bd689084fca358d1512b35c65a4ff257b196e3c5
zc1397dfc80e171e28ab66c8d6412e378801dc84698144bce81c4087e95c8d67b4ba03f684c8a9c
z8f8b11c31c87760c747caf6029659847152cb021ff0917eb7208cfd509d68dbe385999817ae9a1
z045f6b36bf353653b31924d4dc9a4fba380d17e154d9222e3a8036b525da4082e4013ad21ab39d
zaabfb292ada6628a9b48cd49bee323d0c8c1d8e22783bf6ac8d670e8edde9e43b7479e3b8755f6
zdc9e1628802a67983294f6f1595f1c2ab89070b8291a851e429b2cf7a7b89eed6f43072190745e
zc842127a7b346fa3159099ad301465be30e6a837c0374cad3a4b49110a5392f0566fd3597672c4
ze427a4d4679eac6e02ce38d4042279a933aec8580f4b6063edae5f6c052cedcb96b38aebcaf8d3
zda6400b4de7862e7cb267b222e38e473271d9fafd820a1be3c42df2adaa67ba7ab01b3c10d7332
zb1313a1ccf7cc76613ed8ac018e4a39878d584f3c76edbaecf1f5a42df65c6e947ae3eff63ceb6
z04885f4ddfa6a3367f81bfd41906c22913dc279ef81a69631375c3a5331a1ba95e0920ed3b93ec
z927bd0700e3b18a98b3786b51a44cda239a819bffeab861c19415e53b40f66e7ef5e6eaa3b2470
z3e27a22c34ac5d62a8af54061647defa3a6507603838f440b4cca3b621ded002bd36ed22730530
ze3a278f5c22d0f5f803dd80276d446070b6d126577786f93712c5b5f37d349f4b9b6285b1601fe
z3e2c428199514e97eaae3fd7c89facb8936ba81548ff2156b2709e08b202f730eedf74f5d69ebc
z3f79f221f71aaa05e0e0d94523149d7972bcbb0c69448e1e6ee657ef716ac6d80c1635b148460d
z0f60403791bd289dcf358ab50550824febec6188f72c0502deba65e8ec5890b8891e0c1df1e177
z791c6d53a3e5421b4fbd071df5045518b2d73c67139ad8d01e6cca1c267aa723beddba40898255
z951c8d0e1298fea145c8fb0aad7f28d59110d8f98852e3a219f9b9ba290b0e32eedd079727dfe6
zdea0d2bf8fdd9a0fb152950b7683e8ef9ac2922bf5bfd633f6f1273e4f1de30f7e28246a8d2f28
z7d98679504a8abc9ad8fe5522a95d589e6aec525597e60db0a0451b947f46cb2d629cbb2b77ea5
z4765e51c33ff75a9297a59917f414a774e46d128dc44496cc5790b1fee3cb3de227c676420f2df
z98c6c73e63ca491b73f801fe7eac263880b72ae54652a35e7eeaa08d5e1eacbac876217ef6b9b8
z2bc1134c336c30aa3faea85c6c67094280ae31149373f97ed99f894dabb4c91f9eeb2b34886ce7
za3de15d2f3ab214b67b5f907c42966988da60534395ed3dad96b87e4320bf3786b1336d110787e
z133132b961977e322e3f750a666041b20423435bef0e791530e634f39e0b4300aa26030aeb6bb5
za04911151bc5cb16c92d149b8e8c0961ce9b529a8ac3b7ac81ccaefa9f13177a20526a9b07dd45
ze87d374aaf23ed700ed3e7ef1fbc153e197059046cc87a8c0bd37e9338079e310854b3d7d120ce
za034a08972df85a98dbfd17ea0124e3aef025ae728ef68074627428b4cfdb27a66d5e6740f7b19
zc600f6ebc38f67632200b917f2e3281663fd366e39f71868168f51db0a4f1597519dc7e658adc6
z1e1ee9fa259d2e3ca5c2fbfe82da1f1cfa4068ea1f615081b4cf9e9bda128bea8244b39ec70f6c
zbd72cde495163f60a44222bdd8fa4a4846091e8a93f34b81ade8082297672ecd948f88a64b5856
z00d8e512e69c1c196f5d816806227b9be40c0393bac4d005c1ebc82f0d67edd289ccf323737f4c
z8d9a136bda252d5bb73f78604d9eba08075139f8930f5d993374a8d8de7cd36e453c32f85dfb19
z3c83973469c8bd0178d6ac0d278ef6b0e662242adc7104dbf960e4f198ab8c9adde72f6ae04ad0
z185efeaf2fb81a6e60ee7ff1db899123621bfafc24607ba0e2517359c2d9467e5ccda8ccbf4fa1
z3f544d687b915878f326f3e0d618320bd42ec6de4d392f36cb6f312a5ea5651c282f33128a3a71
z8c9c461153a76497af0fb9908320a385b7110814ab5f57639b0c50bdf1bde557a99bd5c4fe9521
zef914496280c908cce1ed3597ddeaa0e362a5f2ed6c543fc9c57abe678c76c2ceaa25804f07443
z828b99856d1f7a1e5cdeb849886fb7d241eba86a3fbd28e6d9ff7a4ca3626c1f1f53bad2a9b4ba
z7cb69e8f1290f38a0a409e4ae0af992aa8db86332374a245a516c6f2848cd6bb2488f962f54519
z94626a02a72b40e76cbe4c8c61014ff7096da60fd24222481434f8d298916a053edd8066811635
z9cec673684d84c9151b469893ed9e1503944ea20050ddf25c9133e70297e7fe038d6c93e014cf6
zd5591e3561608b22a566be0351e4ec4070456cf4f4b82301953b034cb55e1aab6d1b0efe31a5dc
zb989715a60c05d8222a6b82f82864f6d4b713ad2a7d70dd2db512b1b63925ef1a9beaa5f6b791f
z573e1db606553f1ebae00e9b9c67735a88aafb182de43f4f08d0dc7e46fba650d69e113398b6d3
z591dd9f74d755b19c4dfb62f4c69063719f9d77c9aece625f0d77b598f927df78652283460c86f
zb0f52219e4e4265ca5b07fa16abf6bd5dea16e2d3eb37402ad5ab58f7fb61ab711ce0422d82a26
z9c66b5cab0cad24a1b4bdb451be8003955b0ba8de67c5949a42deea56adb510be753b5f1ca94d2
z627153db9719bef217d2b5de7d74c24bf25d18936853da31ffb7d8d39d4b3bda2d806d685c04df
z33baf71377e748d58dfb71e5b1a71c2aa81abe0596adf8827bd53485b7ba796d7a5840f644490b
z35242bc582e8151c8aad64a5523ac8c67a8c051ca3230000ae1d2fa681c9965fbcdae2bac1d689
z83aae6a88551dc17b85807b6e170699b3bc878718436e71f2040891f5815a40562a38020e43cb7
z347828cb2c6982b6a3d183065277301a2043727169731f3b9de70a1c2b27bb22b63ed3880fc671
za9183f3ef523d32164ca8bef874a57bac162fe5ef6dd153ee1069b14ebd6e407ee064aa9df0175
zd646c3a9861822c36a2e73213fe996e1bd29ce86356f151b940dfdb40d5cb718e1d9e2dc1a00aa
z6bb763ce20fbd1757e6921b66b4b73917995a037e914b9f8d71f02a481c8d1e1d7c731c9a07712
z29a8d9a5bde0b2093e43ca9b983bff39f0ee9b016899e774fc726a042cf2fabc54850c8facd1f4
zd37344d57c52b1823014dfa67ce873baf3cdadd7c447f94fadeb5cb5a2c70c6ff7ab420d3f8c5e
ze597d06ed2cf2dd1a19a41a89fd73133b1b9f7e08d8aeeac9d5b380d0f89886253670dde072369
z508fc013a2186e5e9d38e6548f37b02e3fd64b93f7a8354324589f44733c4a4b6875299a54f3fa
z7331128d95fc89cf2bbf355c3886cd1ae3086f9c06662b2972c733aa73d6373f3585d4690a8533
z22fbe2675f855b168e4c088eca601f1ff27e2f4c2d1e0d7cf00ded66aec6cf0cdf6eba312ddb7d
ze04088f5e4a5415aa2ed50c2c494f63acf60eb34dd13eaa32b1b4ea5b0bca2cf342dfecb3fe87b
z44dc928eda32a314152b63466beb87060bfe018e320d5ead3a6ae2ca92746f7da10217dd338eba
z25155d8bf68bde57715f5902c716f5dbd3f55c52876a6f45db6b9657a43b87d2f6df8e0c7715ec
z3387d39b683ab02ffdf6d2cbeb766ea4505a37f5359d98520066957d66d0e2c3f60616134d4cc9
zfde7180be117f8700cf096135fc3c2f1d592168b2233a020aa7e98c7ada56cefcc52411db0273e
zb9ec984cd26fd0cab68fb123525dd470546f01e699ab0b586ee2bb478a6e171d17345de100ce32
zdb4e2d9e56de571d7a489bc75e76ac4c12ec965a460eaf267968820883e65aea938db043596aa2
z69c558c7673b45e2d84b0baf364322b44c7cd9ac804fcb1d4ffaa07e651d14031df5347357eae4
z2da2d5dbd87e2dd7d06e5c94661b76b0794400a17ffa52efe0294fcab7af10dd5cc8f38e6f0baf
z8f0ac7f6918f875312cf4f22f39edc9458ab57da8f154eac5efdd8716dfbc83315b650f2e313a7
z1326376730130963f6058c7f36383b95078af6b93dda0798dd6ad5380a54ba7eff9cdde0be4fa8
z631acb8ca79e2f2a08b6133e945af091b3e60dbf6f6603b985386d351c1cc7d1096c2ad83d44d5
z5fa1a24f474f02cb5ed1cb630baca4a4a8773df7124123f148587ef3ac8753fa3c4c697735649b
zb7933e04fdc685668bd51d7acc933274aa1ea737f7a38c868324926e216ccd7dcf84564a75369a
zbb6e64c00dab867105d36c1935b6c66c14b136416f46b13768220b755a39d1be833903c8b8b055
zc2005dc0168652c44a4ba9a8b41ab7a39dd99b1f90e3e274374a09d6199461e4721595f9df5919
ze8651fb4c250baa85545821f858269417ff117043fc840e2a8bad0d5a32ff3df0f4d60a9a55c34
za59777017a689db0384a9aec05fdbae365dd21be8cab1aebdb0fb17011cb476806993345d0f388
z60c3303d0a64339512d5386d85369dbb7d7da513b79b5dfa25eddbcc20260946c59f9225b12385
zae99274e7a42370c7137543aeb3aa7ce4223fe5234a5c5d1bfc4b7bdb8b09696e88dcbfcaee733
z94e44afda486c982ee0d952ddfc8fede666e1946632e29e0a859453400b67c4fe007d387e6113c
z59362909af8dab91e763cd25c2584b4d27bd4acae8f480607382f7d450a0c682aa1aaa437f8e83
z25adc79b6f3aad2fc8ba63726a7967c3c24214f9d723a7269655ba467537a94f77eca226b006b5
z939de6e2e8b6a6e140af719c1eb1c171c4076cbc67324d14eea5b30662c32a68a19c0126f6eefa
z72abbbe5a9c5a23650f43d5fadf27b0576cd2c29c69f1ccdadf33453ef144f18cb60c7be305893
z8737da824208d28cc4db9cffeb54a68be827bcd312aad37ad116345ddc85bb4b050e0f70296c54
z615637657511e650fd1be3d35e917c0fc6a12d0a325664e4944cf4ac809a5234211bde97e657d7
z5c72d491d8b98343ffecd85c4e6c07425bd2331aaeb17684c23d217580da4c2707cac6d013bda4
z00d61825237e82ac3c867b7cc5b640a6706aec453d6d4526f0b1b8908316048d29664e78cf7346
zd0e90841df91fa9a3d893874382dd1f64d02193758710ce8aed30cd6849dbd90a4f23afc74f194
z6a0da1d593c4aca3523ac61172d679908b39d876506937685cda528a8ace8c122556f105d675d3
zbb27d1b04b125f473d5fe7e6e045c4664ba986886ebbe0f35d28f257b5a0d5b0c4314333930e34
z109e7ae13b6431139cb27cd64349d40e1504d6f16113e651384477cdde2a7f99158f23f270b044
z4e1f79dae42d750120b8dd66c7ca53e9018038434652f56391e47a4eaf27dbd4a22a045f5664aa
z8beb2adaa2bcf54fa1702debca86ad737fe5592bc300dab2cc2b6134beeec9bfca62b5dc0ee644
z2d5c81140b2eef23515f3bc64997bfd4db0ac34ce2f2e03ea918103c0a224d2ced02ad33c9b851
ze36a30c278bb70f9bc156dc9e7d0ec322968d5bb507edccc4d715dfc5eed6dd58b98ca6535f8f8
ze9d0223069807b094d6841b86fbe9874f7c1361dbef5232c6e50dede3fb0c012824ecab1a560cd
zc0aeb75780f7a5c52c81100dd69a25951311f097faf21c2d5852a86ac2c7349b0e3902bcd951d0
z7f0018f40bbfb2394b89b63868b3188bc1104fd360277152eac8ca7977ebbbe6b8416fec269068
z88a7ed8c021ecaab5686c10e29997724e4d652e8f7f3c40ae7d08bf5cf037eb18e79feda2c9d5a
z2198ed4ef72d73bcc4483738fa7c6a7fcfd42192b0c4c292939025b31eddb5d11a263f5b5b105b
zf13957b11cef3d2b42358c567503790c9d28a0c52e604298e81ba76031fddd7b0d274c07e5920d
z140ec8cc67ecb511b29a4caec32f6111034b668184ee5e15f949f5acb5278e8a79cd46f8b9c777
z13ea0e4aa626cc83f0260129c3793361ce5aca615bff74fc7ca2fbfc39c693e8d7d79bea050004
z66f795eb509e6711e239216f2e7068b4435324219321b19b85a9916ec94ee439a813517edc2c90
ze54348899b293b20f1d467139b3da4bfefd40d20c14d52a93e21d4b3d348c034212377811175ac
z6941374d657e82b6f595c30090a60f06c7762ee0300a256a6ba62101b8b3b07e36c1f4e7455222
z7107463268afea7a7c7e5d9cbe8668e5d9bd48a7fbdfea8d2f2ae57993d69e60f4e5a30de15efd
z61a8ebfaef9db4250cfea166e0fcb01a0bff51e55449466afe4731fd504ed97198e955d92cf67e
zc623b6b76ec7091713b7c7b067cc567df433128c2e15e28e081cddfccaa326f1939c61524642e4
zd9415e646554f624c44ccced946ab2cef0db80d75ad9560b0bcb82a76ef525aaaa02e67b872762
z2da51e4ee2f28825a49e2dcb5731fb075cbd3b7546ea74660be54922612bb5f0a2e03068689d98
z8e66e2cee04ebe415bae9b7b30be1f3040776c42abbd8977f906ac6dd281d660453b127887dbdb
z452c7eeee79a8230ad44f379455e39171786ff7c7720d3ea1654549a1d4df14e49e67107388f2c
z6c13ec61f4a00b91590ae3b1c6531a4bc834f3fe06f049b5d8e7c93f8c2b2746b6cca3ff200f43
za4cc2cf6f749f3b45c66f66621e94f715a87e380e095058bcb308e2817c37bd13309bb061324c9
z0e3477a1ccd04064a1e98aa240cb1c6f2a377cc621ebbce40b09f309aae88091346405546c3e80
zfaaf317963703bb10619288a27ef3ea3c613cbe962e652fd9414742ece714c004dbfdc7234f1be
z4ef0cd9ce66417d653a73887368d03e7286569563384467dde0f527638422e968f78ea444231af
zf01e5ee2f6560a81b9fba41d0a919e60470a8148bd7e202f6afb4ef30a95d1a9fabf3346f6b5e4
z7bfdbd59a49419d1342d5ea6d43ecb760eb6612148b4b55607fdd187ba95b59f5cd6651771d2ee
zb6b472f03d209aefe3bbf59e25eef86d2b78ba10d6bd3b901bff586992ca676cb16f9621f1773e
z84ae3e9842794d33307835362e60285c46c7f64f73e04777aa552a3d6ab6454aa8a1debe450cce
za405bd7d1585bae0fa1de0fb39625e7e8716b22bfd2530b5567fed6c8ee83d5589656d37384d8c
z32280082956457a4381c9b033a7917e07b14b8dbfd1539d5220e5cf7549aee8506e7aa8e776e60
zbb69ee1296fba2759b544d39e0ebb36514b5a3ff93e6381a7dcfed9c333314e1f96cabed71b77d
z7f3f9fa2056d5b0627c64381ed0d386f17cdf58a66f19ad09d0a8bff86bbc2f95232da8415e021
z5e9f74a7cb7fc6e65874c111a6dbf9969a49dd34942730b8d8f08c5c185bcf4e0721dda7333a69
z9aaa8702b5735781da9c3f1ace681ff79344598acb2dcbed87d32cd33c186379b95e4c28dc7812
z725fc2cf87c371eaafb3ce1cd2acb1fa665456cdeb9546edc4b64e1593150ea2538cb93dd762b1
z2ec19c6874f087f84bd5af89704e619a777e5dc90d9a71e2c814c62131e99027f56e9a6a0bb2a1
zd6e333af3a34f142b675b2dfc4165c4ec604ef5c10c12cb50c33a6d5c666fcbba4b4255ae342fd
z6ac969f0e943c5e2aa2ef9b3d38af5105532f0088e4e8bef5ec7560aa84b4a4440e11cc4bd2178
zede86771ba2b13b58c682f93c26b6582f3af993cff51b0bbf472196ddcce81c93d1661982bcd23
ze4e2ca4b6b0157dedcfb3bdf24d3b05537da423ad0e493cd27d9830256ce3da676d18b2c7332d5
z9b63e4bd7ca0bb7042fbda89699d1b59b9f887ad6e62fba4423e264ccbae056e7ea2722b255961
z5059d307881992b0dc2edf0588fb1eaa2eefa16b988dcadd414573a3a6758eaf363054d268f9f5
z57544e1a1a50195a9ce4fe22ace454139d38f3e5ad114b6c9ada9dc90451bb7748b67fe7703152
z397c359b5c670da9d8288a043d23a7bdf50440042daf1f0f7205df3a12804c301cf22634fc5fb3
zb6deb9add55b003fbefed70e1ccb05b20c07704dd1979a15f8b560ff3178a682427d8f0cbffb07
z2b18adede15099a710c070ad6960b483c4a2d9f65fc4cb0484705b2a393ed24c598bb02fadc5e0
z0da7602d4704e6cdbd5d3dbea5a5239a49bf7a15bfd732412b390065e64b6828c4a6e783f62619
zd641b212c739e419354b56e19984f79f764d028a4c139cd5a55e9ee723033e1874bc08a9411f9b
zf8b7fad88e8030749ca4ec84c8d8ddc5f15f20e77eace0e8dc8029cac9c8a729832c4ce121df88
z0e8ac3c23764ad43f008fc27f22dd581daac07e91a36600d92137eb343fe96325e3de152e93460
zd0cb5af48035d2a47a15445c7599307251d4e03f9cfb8cae4820f4f6e004a4504a67ea5699452e
z34fe771a67de13fa90d0e47078257177b2b679a602b6f540f954f598deca8fbcd3cac4b5d454d6
zfa8f643338930602853b9ce4504e3f56264d6def6ec8f34ce17f85328f74dfe2014b82f9fc53b5
z8393faa373f062935ed74dad648e7591449ac3cf4a6c62d3223b224ae930f1778089f74ea6203d
zf77cdd18eb348afd11b4beee251721b832405620aa37cf0fca92ab0b0aa1f232ae0419c4adde80
zf8e7e1fca3171a160b4798003e84a9f992e3065ef48fd55d3dd6d9dcd73f05011a43720ca8d97c
z000b107cc9b1564d94aa9ba4a59b014de047938ba22f9da035ddedd59953b3b2c0820b123099d8
z02f6e92f1a890a07305e74f09c108325848805307e5e0225f935c1fb6f592a8cae8896ca950f36
ze5b3ecfec24753d58323cc9fabea54375a3b68ff994bf2270e5541bf148021f527455307977cf5
zefb95d3049ad088c8c8cb298a8cc50ff133d1fe008a13d490af088b5852da04e331121a920176c
zf71a0057f08f06645bb2e8ecdeee6e95dc3115929c21ac8ed67a15ce246588171d4dc35b9843ad
za44a683a38ae1eea0527a446068bd001a6452c1f53bae34d6357461c9707e6a4b3c48d50a18629
z5c1cbf9c5338c219ed3e424d170918fefff1f1acbdaaf4c15d0f93638d6f3d0d16694318720f8d
zfbc8768cfc55af5bcfc46653e09b9da61690ed983938f2434d393e754e1c92ef62893458fb33ef
zb23e659319072daa22bb73b4c64c4bc6edfe3bd648ef73c7a933798c4a875b414db1eff42fd282
zf1f540a6854abc1a60202e4b1a9b89d4be79061d48aa2f348ccf3954e54f06a00c944f9e0989fe
zece2142ceabacf387b774f4d70f6e969a5d6d8ea18c4f49520b55e3b4ec0f3d753acecd92ed5fd
z49c4d2287c07415f19647b12196f652a1706999677e9f2a00b15f3fce52e29af7c4d1f72155d5f
zed486d91dfa0a44c56cd8dd9d838f2391306e7103b51525d7719932b37ecad949a205070160bff
z36b72d81d93466f4c6788a30c6b196d3b0157f6e9dd26531db62a6bbbd6d1e165aae56c401a5ca
z086da563c89aeeef0ed90402adaadaa2c55a07e82ad8d6ff591a7ceffac8bb2571c232a475df44
z499a4bd76d4c24cbe4498f0035e9e6aec78f23c8646295c129abccefcb3692715744375276e05b
zfee44f61a573ca11ae0e45cb8f76d0d9eafebc3fa3d4548e2c92b1bd41012e1f0ec56967567a1d
z0aa395f2a1274999fa10569ebd78e649c87dc13edf2c8b7a3d5f6e6c6ecb8372ae826314db1a62
zc7d1857df44861304e42646c018c71d9a3b2bd4db2626aa9fd03e80cce290920938f5600cd0e88
z35dfe316aab564da6ab8a9d5d98a47114ca20fb708ad2f0b6e7beb7edf1661b9368eaca8d3c778
z9b2d879eed5a55f00d8f29e5caee509d265e03724b3e19d1c90ebf06cd6f3b3ed987eda4f9208e
z49d634d42fd436629c5928d896d330330e7bec49dd49a2f9fa890b4020ffb59fa839206d6cbbbe
z592e20799cd37b720a12577f1dad0d538906f9c6e01b750be12581a2eb1a73e1ff80cd30fca964
z8657a71adc039834c98653aef87c4e0afa56f500bcf3e30c2d13f4a7171eb1152c2d91c89114bb
zdaadd9d85e2f5322473c4fd439697596b73520fe0a6c41ada82218596cd9494eee7f920ab07809
z86ee4ea6e916ddbce7919d50bee2f6f57a3ff98bf7301993486b16c458c801daa573fed924f8dd
z7ad9448bff033a027c13712728c2a6436eec1df9f71c071e096721eb82aeb667765cd4a36594b9
zfc558397001592ada81fe7dd739a9e5d61b87b9a8e2000f5c4044c4638fddafa11aa85334ab8c4
z619760225d4e61e18eb2a8441d6316c6b8f660493f850ee96d8273b8b97587e35afe0a266ae9e8
z7d68f3d55fabd4334835e12ca8f8e52e0d9156c06d6aa4a210bcfcf2ff8f93708926612d76f753
zba009264b2aaf89d0aeaf5f7f9e31f8943b06f122ca59d07fdc327a485883bdd4c98decd600281
zede323cfb9f29014d7f1bea16854e349c722ecf3686c7a26c89c4c7d0dc3446725ee01de7d2c0d
z5a72eacbd52fd44d31998c83373472b42828f03c7fce6466aca9f3fdd772eeca2cfa8b27c6373f
ze9574ee1e824d92a562d9ec852f271cbeaf0b958503d94d60f54d75b2f9273c02de3cb65351584
zfc1b121978f349ddf01d342fa3927e9dfbbde3324806b23d8e81b677a657f8644406ede8130fa0
zdcfa2d90b31e15dd560ed1e3ee68eb8d90bf959fa24736606b5335d039a37d0a99dbe3cd9f9268
z9243952e478017a47ddb1ee3d0445f2adeca44d5d9c4c80b6d2bce6147aa9f76810063382550a9
zf40287019eff0037905d5d572716a679614d488f52883d59f83a69c706a076b4fc7b67dd1b4431
zc715cc7de7c36c0b0ebe5f02abe7973be3c5839a9aaf8ad787f0c04a1713ca54329d7d2b682281
ze4d485682e14a70c421b76eb77ea9d317a84a5f5d4f24cb6e7fc1a5e7dc478fb2013c7cfae748d
zd27d0c143bd1bc20fe0f6707fe061f9348d5ec6906321a5710760e3ac2511e2ff54dc08a72b63f
zd877596975f0363e7f0b86d4c64de3a999bc6079e32a69188d5690910fcec831992c3ac404bde7
z51960fa5ea8de1d9d53f5a62c52b5e28026850697eae749f16b944d40714ed83be7acceb1e378a
z304b6b374b992b7598f84e6d91c07c3a69190d2e6e9741dd04ffab7beed96a4885f911a60927d3
z92aa451540d70834628223eb09b585134f4b7b716b1ea8be619bb4de56bebfb270fc54fdd40b38
z87e1b87adb0f672b16a78c4060b65c1682331daccbafdee988520e3c75bbd1860d5e1cbf9bc0c8
z166dab21689adfbf0137554fd2518382d3427a10749ecb6065b4a353ab14937bccbe754de28940
ze691edee63459b2f12243946223d9e8c2fcd57aa373e9ecaecd7c84eef6150dcabb6a94ab21936
ze93e32be018e1ef5a41a43f5bb8cc685e974580f5fd653a0c38382815bfd4adb91c16729225ea8
z865945b3d71d283e41e8fa783d61df43f64c15e0c53aa67fc6a783f5d4cae072ffae3476e7ebce
zf76862fa020c033e27ab6b29d6804d9844f64098b89131668b3c569da72b0f5349c1812225316a
z3cc05147adbe02ce1183822e32553dc9b1187546ce0e825cbac1430620f0e5456fbefa482b6369
zec364326ea47de032bba8625c6fd25cfc95a35a0f3a13b6c068c2952aaf6f95c8d27458a36e42d
z6f7511a63efda86f6f9e0dbb07b30a394c8b83c732d7dc95b20c4e7efef11280d6208d6e9cbba5
zcd2a8674a9d4e49648734654a9a0df9698a9a502a60cc3dd520f1d67abadf98cbcb649511e7943
z3317c654af39f28bd81017930dee8ae06ac70b521f1cebadb7a6c58aca8582aac4e3971ea25399
zd13a20c0cc52e93760e8758eb9887233443c23d75212b540d809a50a8ecc96b41160675251902b
zd546ec8c4abee663f10959c4518bb93137e377e2135cd0d70752f411601d08276cd1bd7f542b46
z20cae5985f94ce286c043dfbc6c097852b8db9c1248654d09d999efea7a616dc8478c068f9b487
z3a1b919a3f6343035dd5ed803b68112f150f582e0d6b7229cc810495a0e30bb93a0f1ec693d164
zb597ea17553f579ec44479f16ba6ab04fc1d5e322b9781c4df33044173dbf636a4619482f156dc
z26121338744a520488af1244d42b93ed846ab3772e1284f833f87c880a2b00b29ab9ef37704acd
zeb2c9b814ba82b1940daf5328158890c8de8f555b28204fa0c226f806406a6308cac04672048f2
zb8f34ef83feb92ec269761ebe81f3e4634f2fe8673e0262d322c968a7ede59827e86dfb5492669
z7e52fb7a201a0fe95105936bc68d56a35dd0fa5c9628c0ce43785948603463db2ccc7437633fee
za43b8274942b138564bcb82b05cfacefcbaaebb2555fcf1f32a71b8289bc0e8482ced3c2f75a77
z84f0343464c18b23f357cb74678dac08505bc6093e580272cd9e4239ab16ab8d92a11b04171c29
z62e246616e5ec5e6ce27758c826185dbe1c3178c6323b5c3e16b6046c1f0eb501a356f1d0ae89d
zb8909ff894e697920fa601f5a631e14775ddedc532fbc2560be8a78ad80df3f027bd3d20a9a5d3
z957446304f6afd39499ce4a2d5b6866f67d83ca361182b11eab2b1175eb75837c25feff9138529
z6ba1db27e953e90e012bc2508b0770d17234d6cdc65a35b1ec60b2ac678ba5f58244ca34d52bfa
z6fdbe8aa9e2e57d0b83d701771155d0dd8ea9c19a36fed74770b9f71c0c8dcc282cf611d8424b6
za0c6b19e7cebb78c3d1e86b41d84e5126f4443532f4c032175b9a0befec09c469a892332583c9e
z4e7b6d03932e70c4f4187025d53f0bd86fb2228cb7d2d28916103206edc51569a15c989a0cfff6
zc251657a3b29e7d78ce18e1defb3e3da3684e195b810c85a335b96193152e38748cfcf2d40a683
z2bf24e2620f2d41b41045b27fd17e594eb4f88049c356f72d6926e71d8a9b2015a34cea062cf80
za97e77c426638812db8faa7585389411efc6801ec9fe0be7ac8ebb8d2b1c2fff3467fc77fdb6aa
ze4b81512b1038c8d42a8695d5bd348bcb079ff36b9f7c2fee1649c817888cb47f6e77778985b29
z2fa93a1718b735feec60a3da36d95a287c6127ae2498dc3ca80aa09d45c7695d2c7255bc64ca3e
z794678859909def19ed8ef57a97537e839614e9800b5571b145a3629b2e22baaba6c13a46907d2
z901426c6115352a6a51e8b3b881346a91c6451f2de00ad83441b957cbf88a09b00fb84f51b7dc4
z9b2881cec44549ee0a06b02de3241d32ed0426cacc3c897c1810cd07eca262ba123c772177d5b5
z1c5317bb7d45d7c93cd048096e01a09dfa0ed3e368c626bea9abbe24d7298e03412b46b601521f
zbb05fa4365492948dd13bd71355ee3a85ec52e8d5d2fa1d571df3e23c298924efbb1041d61478c
ze8f23709706e0db662d6710385f915c5d456fad3c824643e337e559f32a096a3ffe6332402c0ed
z9c2e69e9dfe226812a145110cd937103e32c8609ebddde700e2f1d6330c34d90264af2e686a87b
ze84817fe485652b4681596dcc95a3663a39c094a6da4dec668436fa0d601b1f52a6fc90e7039fb
z68f7960c5865c01836cdd6ab8f03b5b8aa493b4695e3c4a1064ed83d04a1b97454afa7baa947c5
z0c1d27268c4066f6e7bfbe90cad0a5ef5d31dc82f37c859f2ee2c77769b0342bb40fb753aa54d8
zf81cd8989d3e6d840b83232ef4b998d18e88429ffea393864787da0322ff612a0198621662a02e
z17be99c8117c2bb29a519d80686d57a6a017074a1ce1647ac3fd0937dcfaa9378c57f7dc7c8c05
ze656fa9208b78ed1bca04587455adedf9c47174b7e4a8f8da7d1c3a9436ba239bbbec9a5e790e8
z20703bd1bddcca9f69b7c79f951b73a80828d714b2c12f5d93d752fc5d342b2403e6bd16bd006a
z2818973945ecba4defd9fef2926871475e6a96a7f38ab55c07957c132feb1a5f71463d83877519
z93f93786c313d5baa182ca6701828407e1fe1ac5376b548cd37d52e7974d07de4bf87fbe90e2d8
z0e3455b7cf823f07070ccd96d576c7df7f0986b52338d859d2fead4f0893ee3d75047053c4ff6e
zbbf739f568642a70e83d52bce8e7dfb0093907cdc7806651c28848cfd39a3b8d3ba303758bfc73
za7d2005f3bc60ed16af25a65169fc1b263d47ee43afd7612aa0cc790e2619d98fab910ad572d22
z98652a8f60e7979e983a176037c80d88bd5ccf890aaee2dec757786dac2ad2d3a361241d864071
zd3a14259799795952e74f7fc64188de392336ce2c4e326f1f947cc72eeb442ea234fcc767e3e8e
zc583b79e51dcc68c28030c11c4a4fe619e609126fd50f9fc0ff7617795d52ed0f734d755de9416
z8ff34e51289157daf4fe84a7acf2cffee158e8b7341e2e2de612caede40686de0ae765fa8e25be
z65a1fdbe5358280beae0b39a8ee7e387ab0c5267a53cfc390ece9fa8272315280f89bc734341bc
z05f8d619d89ef90161a34ef7b161a455a75f2e3a3dbce47e0b97749f1839626f474e0af9456abe
z7f4a1d6922ca4e25fd422f8fd289e6fd3beef42732a839faef30a0b6c2f48fedf5d21f7492e84f
zc019581fbc3c06762147302bc9b9e81f2767793b7fff175e38f1131fbf2373f18e5759c7354f36
zd5559c207da3c619ec57d2574e277d09171af97b4a4f2b9ee61233bc9cdb5d6358beda9f16fdbc
z35e2c968998b2d28e06c5f354c027e6150147a960be745e3d857647d9e629f76640c26593f3d73
z9b10028297b7b451db0a18738a9d7c1530baf5af1c1f9cb6e3b3f88234fc69118265f0f3cc3631
z2074580a2a4d8847ba1dfc9654c8209b64be71cd12fc4b92effea3814380d35fff77ad68920828
z9868dabe135db5c9cc89e36ef6de24b0c48a074d839c2c4356c5150d4f2df76687d40a46c3891e
zd8ecc8eac9f83dd39662f67a1ef3e842abaef53943eb00fd20ce696dadb3d769f5f9b80f82132b
z091e5b08405a5bc560680c897a424995f595cc0b7328ac3918790512b51f430d0066d4af91b625
ze0d4f8af7ce5baa9c2a490663d3b010c6f2f4a15a55de3719abc2ce79970e206dc2470e0321b75
zbf6e40b1b04759ac9af6f1948f242f25fbc8929b8fe50c4050a5e1949e4722d2d0ce3cb3c540ff
z4b1eb2025f39679cc8128a3ed52a56bb5e00ee8d23e5c6b6e7aa04b63580987fe484809235b550
za6d005d1dd376ffbcac5d7b73d5793ec93ff5dacf9f095fc96db24e34ce47f4b5c65126c716140
zbedaee6ad1ab8b0c6e1954f2240b07ad006e30b4633acf3a9bc555f0ea8acd7a3ef4438d43e795
z3c2f310c8c7c6652974b222efbb89ab10976cf2073815e37bf6bca1477f1374fd17af9de19cd02
z6fce4ed78896538564ed09d39ff6d310cbff51eb92fc12be94f3b1bd2504e7f1a4e45dea0c4c29
z5e9ec41b1b779eb3783b0c06aa7e9fb897e3f0119b7a4daa52b87455e1287736a6a36121005b79
z128e41496debce6a188e9c10744c6f70e1648f82321d597ab4cfec1d9626544c94a16380cd0857
z0b2efa12b7c093449f3286e82026bb1c1c040a79ab2f2209de52d63b39ef24211effc0781d3fcc
z2fbb906cce3191cd298cc7bb47d049b44b304a17715d30e75a752b2fd18cdcbf12c641084cf2c2
z883e356efea73335e0cfe8c380f9b6a460bfd4cbe44900364b15e52350364861085737f7ecd6a1
z156489bea1a0edf5a034a402fbf7bc903efecb7035b3b68731bb453a5fec849e51c9028a487f77
zf56f88c0814efeccee5f0f36a2a618b3df444a72a6fa7295ddba63f87d0e4c14b521db894f7cee
z289b995832db28ea1ced298bd265a08e19cd19c1f384d0dbd0f5664967ff6c470c6a0419b04928
zda294c6be2c32b020a5c9323c99c9dfc664e42a5431e0377071a3b3256f866fe79e0b2bb722b59
z08420b49cc6214abb0a894e2285b09b39514144294b0e807e7efeec65a7ac3b171dabb16809eb3
z5893d699a03a6c5b5c83e646095249fafe8cb438e053a6d3946b7f54fc5620fbad45c91d0cc8a3
z4cfc9edb993ba6d3a5049cc596ddf6a3bac6507e0d6d10eba33b1f25c72c5cd533b251c618ed65
zdf2d067d6e8ca86c8f7194213be37b21d3ec4e5d28003b5bbe632ae211b0c218f5a8808929bd8a
z6bb18c33b91f4297b653a2e30d3d0c72540a29f4a9f1464ee9fcd4f0441b4374688a82212aa847
z10e1ee8e33803940f66a6b0b29c056942313843e69ede936a5dfc20ad2f20be0ee637087dc5b9d
z287d7108c8baf99adbe11b03a30b478ca4e6d755e46be3f86d1cf30a1e36560e546654d1e2e04c
z57661b5a288ddbbd1a1fd4b4a6513568943c35a84949b0c01f9e462e26065ec508e82df2a2d40b
z820c11a9fdaaa920ccb748cd7a2fdcc4272df2b560a3d345640d6e120903b86fab9387cd501b1c
zab2edb5e958e510f1398b3b3566b59ca489ce3b3e1f1ba3ad9628dd85b5a5c4194df58b93f3376
z956b50368183869ca66151494abc7221d7d62329a5217b663f29e3f6705f173d222582e266b611
z0c517c78f9364a95af814bcc9885b9522975b47cdb6057354face109327b583e2da7e70886f051
z84b20c9956550592166f1bfcef93c50bf36ff4c7e547bdff7f204f0377b4edea6f3a328012aa9c
z11ec30f7e9458bf43157fba01eb438ca01b546594fab5a95c695ea1bb917125bdaa01f9a9ffc95
z1e4add75e8c0624cf558b730db6355885e21221631bc563b85871b67419eaf9f5fc312930d5e41
zfbb1644af649cb48645df72ed67a7b4daf8f1a35f9e97c610523c1f3cc2c518a5df0193d67ade0
z4669147e450000c70e71219f518d7a27c9bf9052a4bf99b5f3e71128e2c3f5bdcfbf47008c545e
zf8c1f72c726098f2a92833a252a7cceed44aff085248b50e7cbc3cbd1d3af3eb0dacd620495316
zdd08e6c3cd960c56a4c493d62d3da148306a815c42fd43c6104f99515216c368ecde6b80db9a7e
z1eaccc70dab6fb5a46f6aee657dc650fcc1176632e748e68452534104bd6d848e930a3d4378038
z812a113ae500fb8f8fee54bc7a9c357948c564cf36e6d018d827b5c7a47c44394ae36ac7214b09
z05cbcf6c0a3e987e21f4dc971c223672988fd69b7b5385f7d1068220f6afc9a79791a63cedc632
z783d9aa2c14bdfc1d2b84635f3d2c51d94c27edfe4cb8d6914dfad9acad90818dcb971ec090ab8
z257901e79cb8328d1afee1431b5a29bdff361d4041ba0fc16dace08ae4fae35b0dd90a2908a9f9
z031b8fb0da585a3531885105756bcacc43aa19cc47e76032a4a6da241492f2695968c37d6c1653
z09cfae89484270f9c6d737f91a5d6014378c6f09075aa1be2fe98dfba81b1fd070084cdf7b6dde
z559ee032568da60af099aab4bddd123940172bc6a27ac8c599eadd3d59a40d7225946477375edd
z88d9c9fe5c98ec29b87c1d072e002fa55033b7946f41ef1a56446cff5504bc87145b2b4c253916
z52e852f501aa21de7c5da0fa31fe89127e31d29761904afd2c0cf87d42052e0c0bf1904856c522
za346523863f2ed3e4853ef828cd5624524e100928a71a24a9449dcd4a45ddb33b0b4009d6769a9
z7a8d0cc0b73243c0fb8408d06ed58103b1951fc79462db0f74177e52346b3606cb10b96717f32f
ze6139af917cf7e812231f0ebfcdcc15a7cfcf64c7d5cbe917d693ceebb2f2e20d8134d6914c8f4
z6d220d2b52043c3eb6e961e0af5ff1938a649066b2f256a6407355562de2809ffd801b6b7844b3
z648be68287d2668270fd4259a44823049ed9a2e6d2c4068c727c50d6893a3968b2b0b8187914a1
z97802bdfad6174a12b62aa6f276b9ebd6c8f07ff6f547614d5fc5d38ceb9491b3385aa36cf4f99
zc4fe1e0b832893d3c515a6a6c5b75e9a0f7471f859bc526b3335e4f70a44397e6c4b5cd8d0c07f
z64b2e37a45cea661e5fd74f2b06d7ee4bea829f81ffd09dbeee870a26ed2d827b14bb14ace4e09
za2e40997c1522036bc22ec73e18a43e9a2e38d5517e43c343dea0a74c2675957f141ebdbaa6d7e
z9e561864fdc49acdd096f8b95c7d40e7c65be471cf2f11a12db59d56985b1e0ec9c635cb578d94
zba6d342cda82da8bcf54cc185b64abd43cace0b845c3721baa0716b70bf561a23945278b417780
ze4241d9a04f59d38da913a3015bf445c6a74bab1f2bd75e3fab66def74855bd653523b1eac07d0
z74c3ee9f011e59f41be2df9b29ba7fa012c12165c487920a2e54465ef1152d04f95bd787590b8d
z30a85d79a51270f5f9f22df2e5782df9880c52405b87365984d519d36b66bead267858f25ff176
z3a2864ff7985ffafe02f8ffc6ae4b2aee13a77a5271d5b32efa129055bf1a7c52ba8043dc5b261
z6aa181a01f193ad616d4d6fc5806527e9727b3766b6b7794b46250b38c2ea47746237358538bfd
z8eadb48d47247895ede488dfa855f90460567c8edb51cf087fb9daa4ee25d2236047b683fa5bcf
ze5098957f8de1a8b3814c1b7a4cc225d91ead8ba93990ec8a13b4a54b34b769faa64b8d3bd31ec
zc74d931e8b7839eab09ef14c35daa2eb5a5d1c69cc452b96b5756c9f3d6bb807f8d91bd99ad6bc
z29be5353dd783e38aac73e72138cbec6c78e142648ee53b3e6d3edae2ba6578042e701a0ff3a19
zc29f5c224734d6fe28069a3f945adb4d0f755137cc239df058a320d1f6c006edfaf8615a5dcc33
z0a7cdaa570929ab280660e723b95cb8553f6c263d91604394fa71e9e9f2690c79ed0fdaa632f98
z858a7ec724e6fe786bd7797368fdb641b7b24360a74e5a589b4351f73b30a39e2e945b1ab2eec7
zb3d20ecb8e5ec899b0db6f0657e2f1c628b7980f537fd40bbfde78daac5ac73dbd2a0edf7a0d64
z6bae404d6b40ae37ad6c8005628545b250f0ee15af461df44bd643b0e22c25cfb8ea3aff133030
zfe4599b71fa645fea140e82aa0f3331747a966b16e30a5308939415a74892ff71b58dd285882b0
z28834fa5b360c1ac276358cf763f67f487655784746f10c4284fa3619ac88a21f8eab6e47d350f
z0edd043a78cbd9a1eb973ee0db8b7fe0a3b5fc2e485f94c3ce76674b4e339af2ea0b4e8872e12b
z040a2e16e52579d7e70e398ed3d7081cb1a87cbd4fc81e5bdf5927212184035443e65b0159ad17
z3ee37953683e60c7e4b4ea2e4a0aebcdec9ca685753191fcde43a0c8e3b0f1ee774bd3ca1cf3cf
z3d99f5c309599f07c4b4553657d9d7bc170b8383fd16fa8e8ffdb6d55a2f8bb3c1d108547f48cb
ze9b5e2ecd6c4e3d562f2e6dcd38028a67238deb1093e860fae97dee5efd64b4f24473b49904342
z2df79ccbed6cc675253ccdd05ec8e83875b59b22c46ee0c86f119847914992ce9a6eae96af20d0
zdd50437590458586e98c9a3146f42e51b538377f7b29e72d42832e388da3639a835e1290f3da63
ze0796e578102477e68fc5db53db160175105254bffc6d686e6520bba785ef3d4b257eb22aac123
z33e7e4876555e8cfe7832cf0a33c2fae36862128cc97926e8c53d96cee7ba9d53a46493d68a6d9
zc94df10616487145ac0e9db686387f6d00d5c21a066f686f714e8e9fb6d8e4e69498e7b2ea43f5
z1a52c6e5ffe0cc3f8ee4804235ddf7c3201862f948a0b7551a19b6b7d4bfa203d11a27525962fb
zd52578406ebaca9a160df5cf33514d45693bb9ec4949519d259afdf1dc1c2318b03345611d88af
z439c9d1ed88feb5ba719ff9d33bdc969e8ff34f22798e6a6ad84ddeeaf312230cfcce3ad8a85ad
zfa69fc087033d3651e0c81c5490f74a70ee64b65b99de8dc685fdb52a34fc3298122a5eed4a971
z459b5f172add99bd702f37db901e37900be4daaae39bb8a44960c12052f590bc7715e13badde68
za29267e76d9d3a3122976766044e02d6447e89c4bb009027dce51e1e99062b260e7aa6ac406ead
zcb17391107166ebaf6845618783e71270a0daaec44340add295fcb96634c9fe9ef54e6e7170beb
zbc527829d2d403ca9a5ed64d4f34f0341dcfbe62c9e760ac7de3bab31625bb9069eafeeada1082
z884b381c96590a465b6b05f7ca262ad09e144f6e6ee420f028a8f698af26360870611f7338cebc
z061ccf9d389a0a282861295193911df9149c78a71158bdc51e1f4366e871d4f117b68b00a9bd69
ze8c27f3b32a2a0b920b45dfb14fe30cc1e5a1295ceebaa7d73c8f2b6b1bb8f795f9037c702ea2f
zed437471954243af6cfa549ff6ced09a163e0560ebf73db35e8d99cd12c83bc9dde356379d14d6
z27afdb8fae8b8504bd37a7162441149cd3b7ac1ae33b052052f808b47621f3c8630fbdb295ef81
z09bd4ca6677e40ff8aeb8a67b1f8e0b38c829b72828668a98a46d3c74cde2539502816dfcbbc07
z7e1812f3e25facc308774c2ba99053663cb18caf5746d0b742ba119b1a5c497739a1740752fa61
z7e2824f5b1a1bc2f136a0e36316f637cb527487c7a4f01c698990958f1bb019a8fddf911cb56ad
zbf3d468e5a45d1a30cdb8d09585733681476c7c2e77df4bef87a10ff01fe6eb2de58ab7f3c723f
z31d3e5aaf7e8d7e4883699da3200444e3b27b20d83597aeaf75809fb6b29672e356dd7c38bf4e8
z9d6cbb99f9e49faeb21efd271cfcf0f3efd7762f64ed700714331e61acb2713ee8035c00b45412
z4919d99911a0bc75b06a6fa016eb40a0eff141deab492ed0f98d66808c41290b02abffe52f1085
z4914c0625e567c057157a95607e306d142662d3cf9de692d884e352f4b6631031b2405bb98a08f
zd7a898c09086394722038dfd238f12668cb6fd6d4c09aac6c3d0095787d66d65ff32f604eb3ca3
z519e89194c2cff0e02ed47d4958a9adc2ddf03e69c2c59af143420061741d5e2aed80b296a2182
z87069fa856ca4fd86e2750cddf6a941b8727e4a6409a240b911f75d2415570f5e9ca8f282044ee
z00020926fd06881ac219485414c0c262143753daad80e354b8c78fe961c2001f54f27f6a086ba4
z98fc34027cdcac3ec1ee9cde056a339610ba92ffecde8abea9164ce6d970d0ea5e24dbcdf2cd8a
z385346888170c1bdaeb3e93462101ef740252fbf1d5735a19be2ceb23ef7cf48b9604635f2377c
z5bd5c4ac7ddb981382297e4e9c0232a3cfd239708aaa58d5ee96a1268ac237fc740e84d0f24e21
z11f7de7b5473faa4859a564733240ee4597828d4035968713d4e5600f7c3bd25bdd8def7241084
z906770b4bee0ddabdb49ca4f4f57984422e7a7a194ecf15e8a05105bbc6b6b815fd20cbeebd1df
za54562aec29f9768517f4bae509e3fa9b09ae62f40cb17a1bc72cb9cfabe9cbec98060add8dd43
ze6789d66c4d802109c1a6028150c1bf87f6fd90f94e5aef040c810a1abffbe1287933aaa49305c
zf7a49ad8cc394dbc5db6bd86146842b9991c325a9ef678c0b3a2a9eba207c06b7d21cada4b4ff0
z08130fe5a4a0731a7d463dfdc79a4988fec8ff3cae655387ce8dad6bc9c87d57a83269c2f6b012
z58d7f1a5d2badbb92828e23d5aa1fa1fb198e239dc36542668a95da0811a8d6e3393ac86fabc10
z595b723d7d9dc386c56607b45641179f87d9ea7272aca78df1a20a0f8fd597c8fc12c9a8b9dac8
z46b67503754a7ea391f40f311fb5b861c07133c1b76d207d7cb7bd4584b2fc45d72afd51968eb6
zdda2abeceb0bb39ca31d6ac995a6fdc7d773bb7797f92a033d6b7951a13898050db10d19029ba1
zeddc54b711e93574dd7bf73dbce7036ada13d35d4a1f9b410421a2de5d8095567457cccb065f44
z01a5e7fe2cdcb1bec3b0c7d655d2ef46ec4b120e41e3de39721649134e1c00736d0ffa82c43b4a
zc40dd662ce904195654ee15161607e9232be2f9f3457c152f5c66c57dde50a18976a913eded7f8
z44853c666ca394cd941e910ccc0b6a1c3ea049c5e3985b550af8d79e724061c80a0c9f7533bf1b
z54e7f50c1cab215aa869beb60e101daa2225d53ca445b37112425e1be5ccc7eca4ba155f19ab35
z4275c01c14989e96434ac0e6545c67f51adaf0c858b287c83ec231c8a8365f0ce5e9e6b946b766
z5b4ac4f6a8c91c75ea59ceff1ce3db18b06bbc731304a984ead536abcdc39af6e02d4cd4d33757
z577935c15fe6d20d1cf33c273cfb89d46e30dc19ee3e65b216604b56cb0860c41ca06d22b438b4
z0421f364a919ab5fad8f08728a307c97ec19abb7fed3a540d20407ff73bfde594197ae29e4b774
z1181b287ed8d41af870bf78fafc5dde6c558913e7c42be69fa3b0dfd17ea59109eea62ad15e610
z46b177df701bccb5293bcdbd890a6d9252f2ac36f757d2d2ea79ce60a31d383c20d099b7f1991d
ze5edc4ce79f442ad6957ed246b571f29b398bd80230e6b6525e0317b0e45a1832be495b71f5fd4
zd06df23bdfdd42a07e0a07b27c5513ce246c8ee72ca4d2203a252d0ad247d9f5481841ce28ad4b
zaf45c88733ddd45c9cccedd785402ec3db81882fb39bdf2de2125033b042e8e6f3c78ce8deda4a
zc4deabbecf61c141e34ccd9aab385828d16ecdd1a14ef787fad3463023678f03efb4cff6a0eac2
zf4b8efc4f97b5cb161b077827a1fe8a2f9b6653e76a7c2cf6f85f1a94cf6f05cac7a9f10df3fd0
z0a56e044127f0848ae42eccd73567c366ab2da7166b14d4488806d65146211b52179505649b855
z6840a7cdff86d9b1041eecda9dbb07d9f1001fa91a81ade94142e46057e60c7e8ad4f4752615ed
zd762595014983bbdf85728ef38de04da7c360eee3fa9fa1c8632ab6fd718da69e6537814ef1671
z38c9786e99916885e3d65523ddd7ecf33fcbbec975820367398fe8bab8268a42b25d086989d842
ze17cbf3906a6d5229b8607090bc97c9117de8cb2cc8bc283dc861ce31e3cdc02ff9265e8989f03
zf9aeddbc14f0f23593ac08b405ac7af5f54edf8730f4a923c28a7218958756f3edb891ded5d62c
z9ef62f0233b77bf8568df6d4f32255bca7e2a96fdd992cae5d65a55f8064697d406f244b43045d
z471aa0288be3c16162fda747045d4dafe7f4c1070e23708a94a42130777041a9a5c51c33b85979
zc699e734f0f827d592677d7b5bad7d084ac0cff823269d15c78c0090b70714afd9e3888f6a313a
z08491bda514d5b731c423da3e93f7af25e9d76f9b1fca6b8f310f4bd983fc94e9044c2396e1cc4
z80c24ba48a257d1e16c221350827f0fb613cbb020091e5ece30860881eafda28b32b0deef0049f
z000d02fe19047222d47337bf2690b2bcb4b81a0a13cc72aad87522c7890185692875a1929e60de
z4e0ee4a7d452bda2f34c0ec775798e3b1373adf9d3bdc050e74ddf4674c79c2d0ccb625d1d546e
zdb7ce1ec318f08a6612fd8417f86ba8d7e86e06c7f25e13629ae4916f2c593d7dffb8aadc7fb37
zf73080d94844faa13469d164da66c2932e1679fe3db300dbfde1b3dcdee361e82147dd1f13f078
za0e4a8958856e9e38fde9da0369f6f08eb7926071d5f5c3320f777ed77918f8aaa8af7992ea6df
zaa06c1e92c9818c71f6d30ef474e73d1904a6bafc17655d5951db52a039fbe7adba0962a6c5c0b
z81db35492f151b2f94959aa5f2d207e73fea15e0d11f59aad2e8a61811b5f19dcf607f7a8f99a7
z7bbca60d8f22d735a8c0f50ae81931bf72c0a64ecfcd4c8238d5701edab57eebbe839e99d72aed
zc58972ee90bf48f35adbcb110bda213899b0e8e98b8aae6589a8c867ca8a60a98599c78eafec72
z82925d0f3a937e52c70e5f1da9cd4a9e6534687d24bf31241858a86b38de55c7a8d68e0c0e8513
z9eb6786e6821bb84c11ad0b45146ae076f65ce62a50dadffec827ac2f107525951f2258a598490
z2fd88048f2382a248437eea439b9dddceaf18dd06598e48aa93810a67be993ec4995d297a24d6f
zc30dea50e747abe1d40e7284d522fc2a78fac6cddc31d4cfcf10acc4e5dd29ce91d32303daa454
z3dfc3c30d1ef3c1326deaf28133ec2f4a98ca4507272d5233c923dc3dd8def0c3c0918f84702cf
z1218837e91ea68c501f9767865872d99aef97a08c2e0e50dd4d2ea17605af03d1051ce506dbb1c
zcf15338c2988c0a25b72f5253bcf022129c5c705f49f9fcae242f60e2f2cb53c675dda31416068
zb75c6a1e594176aa12a32e08f2175b2270e6ffb5e73dbfb19d8677be1860a22fd41143f4feb2ee
z9103a6ba00d64422c3646cdeafa1177c3083a487b4b76f88ccd7ece54b1d5f1c070d93b8d2eaa4
z0b6d303ab3eeef7c62d87d9a8c1d1212760f6d82b308ae516f044faa6b950f799814eb770703e6
z7f4cde53642948405a144c5bf33ed637cae195e4333fa165af585695a8f202a0f1dc397b53cea9
z7edf55446d85d0c7ca4710417902596bc09549407ef9dd122bd321100d0c6b55813848db03b702
zc6f218762d0ea251d7fab0f5f4d9e3c1bf470a537beb876c5ef5fc1d550fcb294f89b470e108cb
z385caffaa350f24607ceb89b988a2380a30699d0a67b6642645addb904a0e07d20b5b7be0fb1bf
zee776e1758a503e6a9ed104dd6a3ee65c7ccf3e0cdac6905b981e38ffb178f1e11fdb5124bcad9
z040195141b008b650e1c18c6a8fc01051a09f1517639c42d45ff01095671d3fa7a8fe3b19b8260
z5a5a3a6e62f17ef7311f89f673d6e754cb1d2d777d96742e3501832b7dc7b04ecb196f07eabee2
z45c2d2db85a6b03d1b6764c287a4bb29dcb3b8659abad5820e0603532790b534f22b2ca34d788a
zc3878f508769a10abf594ce491598dd5206b7c7aaf76881bfa154ccf62e07b94aee6a20e31eb7b
zde744ae4336979a7b8fe2f0c5ae9a27026f5c16b0e9fb662af5d27345978e38274979d630215c0
z5a9f6dc2596aa3d13a1b35e05743f617ce14bf428f607270cfcb443a495fcd7e5ad1147009e2e0
z244b178526cae5577e68cd26fa4e22cf427204ba2fcbb7e6f236e91b7d42439e26859769b1fc8c
zad194a96b4c57ad43359ef64e272ad94518ff53f26d3dfe52a0f6b3afd646f6de4dbe2a9b9fb6e
z550f0c886c8b92171c474cd61a354a46285e8070502fb0622278dda4508ca1c3ecc69086178269
zbde59eea74b62b101fdaa5a574e024c5b1028b6589b4124aa781790a9b30542b6807a1afae188a
zfff73e087d75fc6053dd7bc88cf5f23e469a96c1dd4bd0b7c3ae46bb9b498f6639634e3ca2ec92
z88f3f57cf160f830bf3c278bf4158902aaed4104e723d95fbc277c8701794a5c1541285dc908e5
zed58d7e2dabeec24aed95097cd502ddbedc9a6444d22b48df79e6d090e2273ee7101acbf1cd901
z91dabbc0ccac08f27ff4c728ee9a35673c1a696786bcd290f5a4c557d9142b33199d00822561ad
z04a91153f0b53ac425cc3ef646ea907d1fab3d4e604cd471d5f939cd680490d7328ecb51bc3c22
z962754c6218068d2a62f56013e31a1aabcd27abc5c7e1b5d987cb76b6d73479a4109eaadc9d40a
z7a06e7fa7f77af5b1915d401026995fb96ae34bd2133ff9e61bc942052b5a64d051fd8c4aba531
z5f45a5c1888b6fd573c450bcedffe1917d3cc4a357e3031cd10615e6c248f6ef01be524bf6f225
z076d349550bef643598835cf8cbb0930550945274e772e51e31f9c5711880ab3fe7e806b3dcb44
zabab4fbbce55c164db1fcddda588076ce28fccea786720f5f3686494d4852b3d4e936a6a78ccb5
z047957a1436ce6a6c2d23c7bbc4a6c05aaa90b02f82424dbc7078adbaeabd4af37d53e21136036
z1f68837ea79833e68406cd469a0398bdc10e0258605083cb18ca2d112e32dd79a00072a72c2391
ze1baefe513301b13e544243428022ffb0c71f61edd3ab62bfc3bc53d14397a72d9820e8297916c
z3425a7dcde113c5dd9f572e8421d0a9dee05a84160eb3512f287b601b5b5ec6ebbaa4a6e8476ed
zf4bc69c751eeadc7951d1a36b1d79143edf88740d85533bbeaf4f1048e52ac5f1ccfe69c859c0f
z35a58154ccc6719cf04e1e6423894737f2748adbc3f1508efa05e5a9a00a4b1fc19edced76c238
z82a823ffaf4b29952d6de7954197ffaf9e3e3d366d8ddf3baac4a429ceeb41b2e0b05cab607f13
z477bd4de7fdd878e01d1601667f5f1fe0d470ca24a2c6d872800f040dd4e69402bf7d432082edf
z3d9f1fd270938122c5b2084c8a7e1b7093f6577192609b474c92566038d68fb8a963f58cbba694
zceb709bbe65981732ec9d7449509653fb4088285a86efca0424b9738a7f5cc1d892c8f2f3673c1
za123897953cc99c757a9b019ac21e784a29bcf4c6c43afe005269f33d1fbad5acddde58405d71c
z7fbf1de9ee157a49f6eb0c0e36d57be05a029a093c08b540bf693d8ea4dc39f4aadeb7f3e5f62e
z4de71dd7fabeca7e2b525949b351d7cfcc7e672932ed58b2ffd1d1a15ba3b392e0297d53eb840c
za430182e5d424c8adbe07a0c83b21cf34de4344c8c0e1a2d590321fea6af45f18c14a1b345c98e
za543806157f94eafa39aa53141ac3ec556b322e0dea5e39a3d2009375f6a19bed5da3175c859cc
zf6e90af98d045a5dd87ee74cabb37167cf9ae0878ebc102584bd98edcebe011b9d7ee2ff4a1c94
z67262b9251fe86e65e9a059070bf10b39848fba662890d08236349ccd6d145d2c3ac51a1c93d56
zaa69fe2a77545842fc5e6affbb1f9ece431793a098fad40e171cd02c4cd6a10679e98a625d80f4
zc8b5ac8f13661d5e643830b9c45f1fb90d843c722fe5997d978a047b31d73485db1a779c617a8f
z0705876312d7d291fa107e2f6388edeb4a7edca81ae8b84492d1aae7de92bd0a9b2fbf82c0640e
z0f4dcbfca777c49b576dc7c99ec0e2751ebd08255691147fc9c31d24bd8968ed6fecece93ed7b1
zde79845e59b5e5d5858c147f6cf0d99804610933727e2908119f6d1b3931ba9dff824c541ea50c
z1a06df293c17696a927ee10fefb8c1f76c5e78d313780f935f3b5ed9b5523efd37bace76e266f9
z8590c08b29ee280f088010a28435f8bd6fc3a4f16cd51f2455399a6212a3da9ad1b79902ee18f5
za85b990c0760d33359bc8836bd0f23533ce4dad40dd41b68e2df0aec8115e81fc611d2cebaefbb
z28eeebaa9ab41afebb6702400a50c4979074373229d13efe72be1a3cd006a1be690ec87bbf5738
zd5f083c2de0724a837922593c8842c4dcc6c265d99032ae21b898ffc6ab84aeb196fe0b9e14f30
z9e192216bea0be7d0f98fbba0891407a86d87fb448fa950aab6c3d4dd33d5a018d3e31a94fcfb6
z2ea600bc48126098102ec300fdc42e1f359ecc35eed4324676b3c4ff5b82512468b6b89b9b7243
z7856ad1c5214f5bcc5649174265b58e1041a182f9770fc792e55684a05108dbb6b1c75162ebd35
za1d42fe0930ad8640ccc2713f17bba0a0f8d999a48fcca1b7f6e8a952af814f669a839e3e8380a
z53a98a4e012c49eb5984c3e404ca81f164f21f8c0883f92a6195f4e26ccb2ceb6b49be44ee699e
zea2400e4209f0469a578802a65c5a2944a9e6cd14a634b55984596449bd675ae9c1c66748fa1c2
ze149dc28056bb0f7c7b37227a2543c53c9b0587b57e59ec3650161f21a6617b995838a2ec2e684
z1dfbf8822f02486de29384f5119373f81754dfd40c8f598767a3a051919c4f307234adef310c80
zf972bc66848ad203a44ae7752d579efa299e442f7456fa5d3124a1263d84a1549387375d7558c2
z23fa1681a3e929edbb6867acbdd67efeec65f16cb97fd98bfc821ad654bf5223b112674bce951f
za15095ee5fdb8a54d32327626fdf95e8522ffa7f802080173958be00349d265c2b132a08adbe88
z9e23b97140aa68dbe93fdde2901645aa4b579c273b31d6c8d15952b2fef9f7316f5090177915ab
zfae1f986f3badc6cb3fd433cdc08223e7a6bb72f2a9e074149a304689ed1fa0ad3c8313f46e89a
zeead90148045a77b52fb8dbca5b15b372cfff11aacd872a507f10446bf81ec7e17df708b5fa2ce
zff834ce228d68494d44296c9aaa5e2db45a72510f4efd052a41086ed94625ef863ef146705c37a
z5116a39c17cb55269eee996d66d6efad03d27bb2857c393dd74c191047ee16380dbbfeb5032ce3
z716b9b0599f96d8c3fb9916b1b238c321fb1e9bd1d70a376a78b2d3f903e9803920778c628f249
zcd56dd9075658ce798e8c774d6b302773b5ec7ecb2a882fa687621811c3471dcfa726628b806bd
zdd7fe7d9b3a220f242de32c95ea4157183eb4229c847e667a486a08885a15731867ca23dbcd92a
zfcb1596ae6964f8cfd6c647217b05eace3123397b925f6dd9f6e5a257c807ab09ebcf1824733f3
z908a75267aec00e3d48d7ad730de1a38c6c4fdc154bd6a982da233830d516a4dbd815488afd501
z006fa63a4b730d9a6a48633e5a148ffa6dc24a71d0fc2b84d22bcb1681c225adef664b21ff2609
z716b803cea31f8dff8871e8976999b46c54e20a887ba8da65878a5680ce9d3890862109539832b
zc4a9ce2343df47eb824079c0a47943fc2f90b43ea33cb6f09f42cb50672087153e8fafabd0fcfb
ze4f7b1f4d82b0aa9b1e398f5ce48e0847ed5627e8ff9a971f7ef0e58afcbaeb81cb79dc62e5552
z9a0b8c1027eccea934adc5631ecf14cd852b0c5226183190575ce332b3e3853cb832d1d9c84ff2
za8b3217563daaf04a166687182847082564c1f450dc9ec349ca4ccf09da9f5496211a5e678bf8a
z07dd071e089abc0a53c42d2ba0e0c6d50dc08b82597080ec80c600a5655b44bb8eb5709938b0ed
z8611fd097db53df375114d97d95abaf72a06a3067bcf98b5ef50e18c606ff43e539dab1adb18d7
z7533da3d37a60c6e0158730a8343dc747c27ea6add6234d59a47f654b331d96876568627f29eb1
z46871e066fd9adfd845a45b2f76b2d24d292d6a646f96f818c2d52671fac596a53131c912d3bd3
z58983fddb58db30943dd6fc3aa034855b15e4f3ec468200ffc2c12bb3060007c5da5f91ed29811
zcf68e995538a61a595811551e635f529add85ad44d1c11dec7ee4a86cfc0228c61259efa21bbbc
zcff764a3e9094d47d671828c0ee6b44914425e38d254f4b6353fb3fb0ee3f52d52f07fdc08cc20
zf5e54da2ce50875a5914d46457051b0623df1d2835e7ddbb3aaa8e4230d25ec144e686da7c3f0b
z127097307e017e3cb63b69fab583f8b835df115a82262efff0a0fb1d9daab6e1906b5d5e8800e2
zf386f01b5eb50182f8301794e29c816644205ff29631416fec74ebb46cce88012bf9168dfdcc23
z16680da08122f05db4d7576d218f5f605f26175d07bd4c3ad888adcd2d217075eb25275e5eea1f
z38e3ccba489d533df613e7b6c313655cc642ed349c6c49ef1f847b7f7ed453a6aa95e983832ff7
z6d9ac982049c25988d7cf77022aae8cc96c9086c80037e4d4905462a84fc2dd9705f1c8617a296
z8a19cd7424ebd79f083e32423e857bdea06778b043b2515ba1bab19a10a23f3190c15e2ea193cb
z7ac606f62da8d0246bc088c0230a7f37cf84cfcd89973c4c32bd6b83c6f1830702af9350794871
zdb4c3a58b1710fdf2c0502c06886b3ce5ad5757c583cf117b71f3bfe7064132bcdca46af39b37f
zd3a699b3fe2e990c9295bc376ac6a45da8c7af46c40d36b456691587161daf0a803442c024661b
zdea0df3b04caf02b317fc559f499a916596d967bac35556659bc2b70645635586ed5e719f3f3bc
zc72d211c0742723de9cb6789d1e82221158f482d72b19f5264c03f85cd2ef236b8635d687d74e5
z5b5e3f584e40421f892c75c9621a0d778458725e287f8cdcb1a8a385560fe8230c7b543d8587cd
z9c9c77adde2d075fe0725f44833c5e89f174a3f4cb2401a014c92688df013971a895b9e49ce88a
z3da14ac628a20e523d4db850615ae0e50b708468e49dc3a1adf776b3bfafe2836d42593f9b9571
z7757b484f37eee61810946340bb62106901791341271113f01a46a63631ed3ab98c43dd4a19534
z89653492009a0cb6ecab77cac1a5a6c7e74baa687a5cf8cb44aea38d02c36915f341ac5088c67e
z6952500065cd78755dde2af038f2ee818421f414b4853e98a758d7d0ccd506e685818f1f013c7a
z0c53021f5220b87244d36ce4a0404869411e182f89069b1ae24e54fed79a53377e25787575df7d
z480597c51cc9ae021d9590b645dfa7d3eeae044c3f93a95b61c22343a322f04b0c05593e6d8f35
zeda479f9b285c06158da01f202857b3672ed7f7f510a75b182981c8c6811d4009d37975c4179da
z6f188c36d7ba577694bd9f51dc1f0da06c6334d6abde0ca309ebfa0f613ba742fc7ab0a9a6de4c
zfe8a7a09f84eb615f7ffd265d1b8a515776bd9084ee7e7b4160220aa2c6d4c71cc35caa2fafd4b
z50edba866575728fc7e3976ce39de7fb737aad82587c6ab4b01e7ec781eb1c1dff51013b0636c4
z1cd8d6b83c4595cfcc3f92c8c8afbe4345d13e2581a2f726fb48710e98770ae16f4667eb806f5d
zb57cce7218f3d3505d6111018d92ea11eb310fc11161cb0dc8a42d9efce77bce5e496d7e0afe16
zbf880295dfe2ea36b3b06368f37be0efa9b1665f044c340bbe9338b1a601198ff831f7fb9bc80d
z0dea0dc7b8aa6d54ba2ee5294f7be0371f50228a4bb2348709355237404a909cd0a9a7223a6e78
zc561acf19b1c25495649ac28e9b9f6796f10acbf97995a310e85c6487392a04e43e4f698dfc43a
z49303241946cda09a8f9f322dc888e3f7ede3b5ef03d4abd061febc070ea444badab749f745302
z570e475a9a05875e40d1a746c9874796919db15f1b3f678e81fdd5cc82dac729095c1e90a321c2
ze5e85c93b84a4985a016987197821687ef1cce64f0bc23acfd0bd0297205a634854cac59b6dbda
z01b126446f7a4cbbfab38ec96d7e37ec9fbfe4e3f9cf06c46ca8da9f604a0327c5f7771e7953b1
ze4cfc6031ba57f3d2efe63721351e379437543c78410670ed31ffe7174ce473dc38cf5d11f5488
za5473fc706b0f6fce46bb9e704baaabf5afc6171d6adee865e3819b0927771d2c094cf754e52bb
zd441a4da70ed52e30faca95d58d26d9a5616ad5fd16d022afc362f0f9b105839a95b117a22da39
z26eecc165660d87da37bc487a79d8f068ba6b2b84edf589d5e2e1ecc3fe6636ed8188486511383
zc3702695ab68227b378d517ddd2df75a3d697d2510ca0748fcfa5cb7cd94c493b8a15f033480b2
zad7336e8ea37b9ef705ea5eddb362593fa9438833f0b14a23bc795b560cbbd84b502fa62f64c87
z932749bcde7797b98568b22e13eaeac02cecfa928bc509d6cf8105952156479300ed9f27854554
zcf9cd6ea9fe4576fcb92cdcc262622ac61cde2f2eeb6f16e107def83f1c58394a9b5015eefcc8b
zc6440b882fe85cefccd367c6d0e46803df004c268af08d09bb2df27e94484ff07a454221b5e06e
zc47cde491e696a7ab5bd5468ea78671c43ea53e7e0fbfcad30084e002d4917a0ecc21e58194029
z01d84009c0f2c5ec85c5595cd47ffbc051e26a0d1cc785f90dd003c25075915655d978819e3cf8
z35b0e3c82f512217e19481a9afd47a73fea07f423fcbbadf3c617bdf3a9104797e7d4835620a31
z293ebab641c426a0d7484188b0e5cb5536e7a3a66d768aeb0ee7a18810243b5709580c7200aa47
z8fbcd53bd777d7044445436c4c24bc7be11e29d4060d5469b2b8a604bfd8cbac0d21193680294c
ze638a411ac2ded769694dbd05f1c0c4ef8ccc44e2e4eb5d328f547a60eea01dd31dca5af7ab47d
zbd5abf5eabc7d35333c0845ec6708b4ecf76fc20c639616eb8b30c2649f6c4f01ed2a8f801eaad
zf3bceae935194bcfa9bc5f98530724afc550af40c2a3beefa24a0d244f0ee79ccecc2607d57314
za930e78573beb56e8ff301b6bff9154351e7e18da6946a7da462575a93da42caa2c3e82f08f7f6
z327e4d7112cf7f5805b1c9d0f416070fb40c7791856f999b430f7b213c8cb8fed9a45a792179ab
z5bedfae3836e57f7a16c29553eb80c8a63a3af82dbafea6831a00bd9ac08d344b604bbb812d55a
z0d9b32c7bc617148303f08c1adbd1fc397e8f181cd1efe1dd462c265c7954837d551cd08d8a237
z0cd6e6dec546dafe366c2bc77190227632f0938794f73a1b7c3c01325cb409471963b0f40f84f7
z78133eefbdad6044b2417a91c4243b3752fb35f2b3b615dfe8e928cfea7fc2bfc08d46d9e54e15
z80a91d4d2689d9c5e62a5dbe8d90e06b391b15cc684259f48c3ca37581dff6c63a97a167b445e3
zf5141496c638a926c7e20c9d912bf8db6ce468696031e6af37522e5e8075820375c965d0aabc6f
z7e23b01993bcb42bb9212e0d4341a1a04a7be12cec46b7952a9ac6be18d93df39d3f0fd940e269
ze0b5333e181f868bbd9f7373c0da44bd57378f16334c02710b5ca4a948ef94a39665861c093a29
z714472c3731ecf2675ad619da911aabf471603e6aded5c3209290b34721ef3a1ea1995137ca1ab
z1b85fc28c2c9bf88bafc59f178ef0a5332a1bba18820ec81c81206dec847ce6c9fb50bb4a8cef1
zbe6af10dfa893943aebdf5950d5dbd0eb964084e95d7c057fb3ca933dd0a4cc937e8de278d27c7
zb0b7a07b94aad4bc16e0498f514f4ba5802d13da77259bd2089d2e4c7926848133f5745932b97a
zedabc1ad674bcf3370f116d7d52159d378b1ba9c8015f0452178da7ed1d647f8a2ff0a8b748998
za6f6cd14739b08adb1d7a8ad1c1a6c4eeddeb23a845c3ce977790ead898babeb82b744da762dfa
za4f35567b953683b980a026c017d14c981cd754c0e5924e00b3415190d344458ea48f04b307eae
zdf15e8cf3bcd69e29a5f9c5ce1f1ead4a4194f9b96d9c997a7d32d4051b6703167a2d83b4c84f5
z82b728437c79f0c69639745171cf05480083376b27deda8caa4d7d527ae73f30e2033b2def151a
z1bb6a1a9f0ef7928e956903522f39d0c4618bfb87ae717828fd2673925c360e18d8974c0f66cef
z7dfff52f65a67ea7cabc043849df4baf2e0fdd4a35a603e0f4a25e505415b914e086aa3357a7e9
z6f1a19c684e471916e5bb50f66836ebd8168fb6323f415cc6976e938463a4fb228b95e4fe9d6d9
z069867517ab2674a45cdd88317496b3b59506633507f06330be70ded4a600be7fffd3aabfba8a2
zbca5a4cb34bf7f8eeaabd3456c16e6fb6c682a9aa4b391e09c8f77fdacbf22e21c74c422f6abd9
z39d2014982e5c416145ecfaf83611ed442855c37bc605a622dcbf658021e2aeeb7ddb18132b121
z01e836c014285dcb2492fb16f2e0a05f5d3503d2bfc6913c16d44b09e8b7cdd7bc5b394f20ffc7
z50aa2b77262183e2122f6f15c090f24177e72ffedd36ee27136c8a3c64d60c87c179cb8b1c143f
z8c0204196eb99ac1a2d59df61ca546d814ae7ba99e878400567ee994ee38d79929b55f1cd0f104
zd8f9b2c35f13e2bc78b77e2327e8b94bb58d629d1802c9eba996df8c5b00babae950fe16cb3a45
z10b2e03f4a28e9bb90e7cd661bc28fc348f58dab72c0eafebc1da35cb4351362f5e71162a02bc6
ze9a352686d95f5345263b6e6fdd1079c3b301c2766bbe3a94ab21bb6eb47ca1b7fb344f90879f3
z0061d394876766e6c360d1b0110361ba91306dcdd418aae451cc6ce8464c350e4020140b550e34
z9d5bb6fd6c5b03fefe61037766aa37d0e7accf1bd7c314a552479faad37ab4121e3fcdcbfb4239
z704a31f30b55d81f86c2a79fd65941a6ce36cd86c07a927d9b1cd6961b8b2dbd499aedd84e7b25
zd8327e0cce87ee67816df3d67498deafbe0c0647ac67d3917035c3ac9c4935bd8c6f076ed72136
z10d4e2e76e6ed50e61827f9a98fa1518f75c67c7fa06d368979873495ba5684daa95ebc7b61535
ze9ba48ba03017d2c666a64df1d23a11637a90b3377040373443d735a1a5dd7ab258e9ca926e68d
z06fe36397f2a1716cfd5e60ad56eed28466ef03d580343ba082168f62c46cab085e64e64f98804
zab0fe86db23efc76a8f22c704aa7617f9ebe960d54dc1e8031862134d085242ddb9c47f57bf1a0
zb1ffdef9b4282893040d3ae7ac52e75af12b9b680e21da409ada862897faba1da8874a2f25b1d2
zbe1f731100b84a408780d8c2b9ea0e17f4ac0f0b19a26a6d465f4fc7d5f0d82953e27c79cf18a0
zc0cdca8b0fbeac1f8c58f3833869c113b8f264d43c1f8ce1d3a42b9fbcdcd02374280e7d0c8a24
zaeb2d0977461daf175e126631012c3d6b8478013a2d47ab2450d98af3a4b0b0d2246319cfbba6a
z22dc289c2e4ead373733e974f04aacd299d9691b27c3dbd69c2317fe50eb9882b5c8de6adfcbbe
zf9c3b944ad7f91d328046890bd79a0e10a367fc63be1c4bd314d89cbf1246a9dddfc9e791b5d8b
z09896d256bdbbeeb6539f46265e6e6c644d439b8cd036d689f84ab248980884c1a0883f1bb7c62
z79baea49fec8f209b57f58ec0494583f8728858319d4aa90cf09d76da2c59b905d25d0c68717ad
z7c5c901fc8b3e8a6c889564ba1c899c042c05b4f84205cb81eb26888ace741444ac013e8e71b6a
zb514c5d7b73d61739306409f7c3adc63109c799cc9340f9d9101e73c341a3eadf8f9deb2845663
zd3c64ffb6660fe2d3a182433fb27c714962ba30242f4871543c435ff663be17af810166427d2b9
z0176a3af1e1dd378bbaa87fa04a70f0113114d5190112ade087905492598c2e7b1d6fd74754ae2
za278e62a8263d9a757e02fca729282d2d9165f1280b9e21aca929b9a86a9971ccb89e8893c06f8
z1050ccaecac77ab142c2555febcfcc01b5afc6b52c0ae2620502fba5a288d43a39169bf6b9dede
ze54d32fe202450a93884116e5fddbf29b02aaa6b189c308dcb9a76acec3b92e99cd3f2ef9dfa5c
zf9f771fda9989b3a9fefc9c8eb09abfdf7c9b38fc140bb16563b7722ec8582869a211df54bc3db
z877cc1b02c77cb2b5de0f4801c7ead91c5b9f3ed6ef53643c362166e6f257a541aeb5b94e17d82
z3c2b5dcebf5e7c46e9e81ed7f78c8377daece4fdc5c42322f67d5b04415b42927c847707fabb2a
zab3d1c264c900e8eb9e92a962fda3b2bf2b50cb4c1b880508774c78289e2e32f69869d3dbf897c
z87b999a188c2772305711164c4f06bca94b1164dc689365beb3135f5cf29a6d710d9ef46ec5ce0
zb0325ff14c990a2a4d85df7c94d10c97dc2fcc56a26b4cdc4a18a68af64669e62cb09b93318287
z510fa7bced778c5636fd9c3c90bcf0f250a503183e8fd2e14ddb0e0d85ef07c114e18e7967a9cd
zc1e7125b828aa69dcad47b6f11df1dd7e77193ddf9f0551dd232bdd1c6275b3d29396253b957d0
z41acb6fe6cf66fe82bb13665a1f30c1692f1481417b8967ea44218bfa0c4fdd41fd97efd7d34f8
zd169b505b999b28b843a88cb03edcd95ffbba0afc3481b3062ac6ca2fff8ecb61331c5ad2738d6
z4f38b010d8cdd1c7abd8040c34bbbbaf530be2c13b1782d691709c907e0c8785f7c5e5f1b3fe7a
z9d3c669d51ab05342d1391452718bb9ef6123e2df43d59e99bf9293880f54e413df0080a3eae0f
zd28aeb52cae2c1aa4bf18e2e4dc2abfc228f7d49863106be3fc2c830f0ba7dd0a39a0eb7c98863
zde81b46e3a22cce313f92875a7555f33eee770a978695b2e5957213cf2b1f44f45d4406591d571
z774a265e1b3d75cb466be7f2fddebd5d85fac6a8a025f5f50bdc6d09a7d25ed1d8cb4f61743f66
z8526e3082cb18723046070d7653b4d05fd6a73513f25b5a23d40f44f6e92d926836fd1ee1fa72e
z32aaf8b5066d5b8c0b85d153cac0c09b987053c67685e6617fcb725376dec86ac72e57833cbb97
z7844199fdc6d52c8bac88f2dc1f81e983f14428bb71b81d2bdeee6abd70a4e29970c4592b1f1f7
z001ea4c87b8c741cf5911979f20f42120f0266e07addaf1138c95ff47fdcab47099f2ed9e6c9e3
zee14de8516974312dd74fec33507d57a8b81e194f2548864a772d0d6f19af118405d4d1e6221a5
zf77c68aa63c32ac00c2430cee317a4c342389585e3c6a1985ac4c76b6846ba0e5dfed86afe6ba7
z565511f905e31c8d8509e6b9759b3006e3ba8b13acc3fe259e01b2dd6260d372b2079fed22a696
z8197550f03ff628df9dd2661a259d7add7f2ee363f4179f01cbbf43c227ea72da43e5b09903752
zf4751c38e4e28d689e903af6f79649eaeb4872854515f569fdaec8fea26706fcf20dc173a6fc72
z600b6aa3212d64357b4ad3e6769fede1e0119ea31f053f8c24b380d38ed53eb5629f9b8ade22fb
zded0702e52884060eea0c02e2a7840ef73deb3fe4aba764b758a1798d6464978005eb4707b49de
zff54f4bb5a868eb92eb37ee989aa2a74fdb906c61a00bcaeeebc1e56eac6e5d22e9c1d64a8d047
z79373daafdab1f6cbfe80970494d67eac100d1610a0cc52176fc10e3df75ba78056038ff1ec8c4
za7546f887e510a0d42b78936a3263a6239d8f92f0c55d192119618fefacc3c6e3d8aa04216ff78
z9c434bbf1c668df59c997beeb677394a11730088e5b130a3a7f99c1d287d660937e2c1b1a78a9e
z57e6bd05218c33f42dc6e526f44144ab917e52a13dec3d258d56cd25ad9af037398c65f50e59fa
z8ddb85820ae09912d23e23126b37dc81cceb59f45c6b69cb8d24c82f3f1c934252ca01d8784e49
ze6290ab4d1dbea3f608c4a7d249b9696d838044922cd887e6ac00a59fed22000c008b934aaa29e
zaef673cf4b35242eae5b875ae3ed6729985a4050ec0a65129c7ed155042451e811b5c92377b4ce
zc96a2ee1a82f193ec7cc525c4d23b2279ff92e64fcc1fc8382c56905e9654b9cdeb7ff410f35bd
ze142d085cbefc2cccef74d2081847d7d6e698b60ab8718b24a777dbbb9ad97f5845dc0f7aebed5
z038926c3fd973a0ea98d3df0dca326264ea85e4e86bbfd90f2c50507d03d93ffdef087085c12ee
z5908e998ffa812ee5f317c2093a989bd73922d5f037194a759db62cab6558be7f696524ef5da29
z5a40b5783f0f7ef78b9681ad7264cb6f4c3844f1fae47e614392c71fb7b55ffda745b365f5c706
z088dac389eeab33b7e7c8ddfe922ab3f9c9fadb874eb61b1ca1e7b7e459848d9b366b27a35306a
z8e8413873b2c9761e732964450ac123cd36b68fb7932d8b00a368cfbd68af9b3eaa98445214832
zecdf9b07ed5fae18c851074f252fc9d0d8ba20e8e766def0cf0bf79af727f1fa8a50889b7481a4
zba15f56c52b078637a2ca7d7d1322081c3b0d6871a56fcfa91275bbebcd81d74587bea0060e5e8
z26ee43f646f96930ddd7f381dac651c155ea78ea0460f7a9795d1ba4c8f3c95451d11703ccc2b1
zc0307a82e8f750ba367600e42f2b78529a1431a24baa5647cd87d34e431d04f0e95b8a325b3ea2
zdf593f2f6101627403e19139149663c525830ad662ddb5810f6c8e2bbf1491e97079619ebaf86d
z259e9250b5cc74f9f9b127de15070023f20235846b2925675b2ffd74cf50a07d14d4e041862c21
z95470aa12dc36b38004419b5109bbf37363b0b2077001e9cb579b18ea5e7427e4cc9c23e9d80af
za169373ceb2763ad66d07e3f4f5af2fd598d1b40e819d6821138f02fc442b2e804703c8c5350cd
ze97c088b996783b85973ac993244e85acc0dd134fe5f1eb059ac9822bbcc280cffb6f6a8da2ec0
z971df5aa6a56912bf0d32e6622a1b413947ad5d4330cb541394830fe0fda3ebda084a21d5e59e8
z766940acf61e33576115e21f36e739cd2920b1b0c56c799a5e130c41821009082a098f606a0eca
z4acec8fe5bc0f819548792e2056e4b0c0c633957140429cab1eafa97b9ad172eb19eb08654760e
z0a88724d88f11e13feb24058a5d6a20b0c8bae75f060619695425a881272f3ad2d298f40df66c6
zd5e1117adba56b240704ac53a65ea0bb362fa4388e96c2ac0c7d540d6afd3d2a7679fde0843b1e
z3b42cb9fdb4a00d08a8b6348488bba2856024ef8f5241994f5f9bcd5ffa895496a8ad7c035f066
z376207bc610805f9efe7f637f12c0857e2bbc23c386adfba978549674a213216e7df2fb6170b89
zbdf06bde1c7542a6bc3c6296f8cbbee61c96ea64a758d0b0d67b62e88d479319e832f710a64636
z9a5400bf896a365bc3440df0a0c406eeae99b987e8044a465fc92d14fa0d2a3af149c8ffb23955
za2906b7bdea6d03f446497d045882ba32230ddb84d2e3c902b20cefff1e9a0daa38a3c0405a9e3
zf6dfb15c94829c24acdd703c4268a563059aec11e6ab29d15d404affdd425d0ed5596669c977ca
zab3ca840f6bb370ecb1b7f3f5c5da2f3bb2726d9bae56833f0c52cdc9f18795d0427bc22db2394
z3f0f75c416e0f022f26472a880958b6ef050a89440fef36493bf07a7e18b2929af330c54247bfd
ze2e182ef2e0adff3a3ec26daa95304a2d18c23d77630504408f31dc219556d66bb2176afd9818f
ze6284c6869277299400ed444169be2f6c03f88594fbb1a8ec40b208d79e900cebc97fc12e09462
zdb603551b23fc6a96c7988e9c573f70e392e2d3297df9a0531bebb598df2e84534946d6af7989c
zd0cb286b90581cc6f1aa7d57eea7a882441208b6870d4715a63ea8c784cfd9b868ec2ccebce3bb
z4ae0946de896f8c23d2ae2a85671bbbad55e630e7634f0f37d3acb7b55ba5f83272e6d7cd8fe65
z5d48db8c1b1c969c984ea40e0d4dd35f475b9d6400324ad376b8b2ab025544ee1695670f6226f7
zc7a765b088202bc90ed4dc6e19ff304b138d310aec0370b22e415cf63579ba630334fc6e41e579
z387af4d4b7236473b0d0c55d9237aa8c99cbbe58214a1870a465985996aaeb8179dd5beeafbb6f
zf3f5f6dca8fd68cd9c2cd07cb6a2b7cd37cb3de493700da5266e0c869ee816790beb12c50c0620
zf4a2a432adaa0d58bbaebad66446eb3fc1daac792a540759cba30449127dc9443e677a3e328d17
z0fe9f4e0a0efa6ba45418eb2982beb98601c67347f6d138294f1a1cb2bbe2f8a30d243bd07401b
z3b4f3eeb7fa9e16476fea9f00cfc4b3e4518bc1da155b3a2e2c76a31199adb60b4da8f5bd6c732
z76da12c2f3a4ccccc06ab43c6a521cbe6546f46cc45d14d137ee9de0349d3f8358f4827f94ca12
ze3944c909b962efe00d824fb8d06b42d8faeee95925ed3c623b78255d90146aa2f0635aa1f21d1
z1bbace6979bc09824f34593587b1fcbd10e017b8e02715800946722dd0c9e6950ddf8ca0e31ec5
z4e50b4f8f863d13507471389fd8b65a6f9902f73dd435539f10d504997d640da4cd446bbd6d86b
z78d314630fae368bda9d1d42a60da1aaef776b3dbe07fb1b88b59aac12908368ec94b020d6a25c
z78ef5de8ae34d87d94f422e60aa762a9d23c83b489dab2b932c1dde357d82e6e04ca16401a7cdc
zb55efc3d0082d3f9a828c7191ebc0c27f2a78799b7d905b8f26f8df28d9718b4eec4bccb492c9b
zcbb58cd3141070c5b983de7ff97c662fb076c6ddf20d2f874316506a292dd022bd5edcad683ad1
zba57de4805f3a1f752fd202344a1e17975468565a541bf036f4434213a8bef83a4e9b845c39a46
z9f905d36713f9401de66e937c43f0e7d0a558280d8d443d0e5c37d8e54992e64cf4abe560f0dac
z55ef42e9ad7bcca65c8a23e475864fec7f0ccc28c9721ffc608f6cd8640095669542c10bca0f1b
zc648b1e956a0f39aaff05f816a65214ec7a43bfb7c65e95e4eef19d6e27bc00980c0e3ea1230be
z369feef46a41b5a73a69ad45d0e2af9a7b3a00a2e12dce6b0d31e231f26bd8004a0d009e1bfbaa
z1b94a34096be4405e1831c2ab3425070c6f0124807a335de47905275e4c8943f6e5cadd238f9d5
zba28112401aa4b2fba9650e3c0d6ffd37b6e88eca6340102856055db066b23e7e3aab283d3458e
z306466fcb84da9e4d5f2418458f3912ceb8a948d3cec460f06ed1d640063264e41f018e47cbfdc
z1fa881be5d4adb9de2eb9dd938f25f316eb452100657df763286ef69febb51a50f781448915514
z1f4c5d6b5b90852bd3694d932a8a385ba11cab0c051b8fd90d9e8234e7ffdb3811949ad855222e
z55944aca9d5ae33a0dd706e347f940040b2e92d67fa8cfa1636ee5df90abcf5da42f37ccc5b61f
z077bb2557fee0456d2b07c8b3820b623b732a41cf62485742af30ec8bf5cec590492891f11be7b
zad3019a83e915f52a63e4d2f800f2eb654358f54ab6d8c654685c1b255683e5c5bcf762d336166
z7529984268ed1253c2edfc32c96872452d1c771634ab20c282d7c59e2b09c7c2b419408a0abd53
z2361e58641ae816d7abab95917f8e381bf28325d14068f8d37f7b14be25b194ea8fe3e9ec69db0
z83c58381a3ae53c98910103dc31dd890912ae04bded7bfce4da6000de18822b0ee5b8bbe5a548a
ze7c1a624dea904fd89c1eb1d25d7b19caf8371bb47678fa5cd5f5bfb80cd78e5ac95ab219708e6
zf8a3ba3c3b45dacde60b75f144b6d6f7720b417a22047d1de19ba8551dd0377eb044ad044abb81
za4650086883a3f5b7726d2352ea1c1b85e3d165a5bb4d3915e22811c010a4d7fd2ff0ee00ffa26
za7b0ec23ebef9a6a5a9d08533e0dfd8aa4c06581f8039221b8888864940b5cbe99453893a4e3a4
ze8733861f11a6f9a3800d105aff2b79dd9123d2f5293d53c5f296fcf49ffcd14b828f6e8f35f5f
z3ce72339198b21eb220c84970403396b007790d8035242351d11fba4af59962222a9528867aac2
zc764a66f1664e3a17222b79de2705a74febb4d38f6c8a9d021267f3512e10aee495ab6ce2d1c58
z902d572cbd38bcdb603709481ea6e347de35eba0f7599bfae91ab3c490e31ad1dd8fda08adff69
z80ef2348c026b76d05738f410eb8a0a17a88e4d208c228c7f08e475d94e7172e17fada1ce39249
zbcdc66714c23831f310229a31ad76d6f0bc6113bae56347ef1350b464763cdd880908471ace1ed
z773c86fd7f497ed1e79dd52eb06e470a355f43500c3425947a5c0ed5c9e5e562fc8b550b20f9df
z35d460e2074cf5b1622cd4ac2fbab1984ab81ec6234b447be8d9c8f76a00ff10048540dc55f16d
zd72982b7e44f8188555cca1aeae792c2da569039c41a85be909dfe252b1100727a376b0477c419
z4e516c8c5a56330270a57e2fd2eca2a04d6052c92b948edd54b8243e021edf2a116575fe8ab451
zdd05a3cfb987e7db932e2ffa0c11c8148aeeeffaf66c8f48545ea49978fb8b104b8c69e69ba2e8
z64949e534c6897b93bb370dad995b485507f8e9e1695da9af980d16cfe8f792fed457c1bb69798
z723f1822d98b02b159db49727cda752f43255d290cc8382cf9c2765ea06e041cbbe899c05dc5e1
z7ea43252091120bd82bbef49558b016e279038fec8c738cd8ac149c2e64414d8e9f599e9283a96
zb679083ddab5c5c645b84684f76215278d5ec1139dc9ee8442aa8c00a9470bda5699f9f5d37906
za9fda72b62e4518c50d533d3e6a6b3dccfc133a9884ffc17a464091e2ffab817ed042acb9504b0
zc192d125633aad79c6129c8b8116ee272e5cdb8773b5cf7881a8fd548c5ee1ef3894b1940b2c61
za3c297562ebf497661cef59b4d009ba029879f5b6c7bbd41123f29ff2ecd334ce698b41f357140
z6b70d7c9fd86eeeaf905472ff1363c9e9f014dcfe2fd6e4de7662fa91b4baac1a1dff1f31fb54f
zf4c74e13fb13ec5087b19dc77e900676c98a52c91b6c44b28eadbaaa4266d140f0a25a165ddb83
z72a00f07c4383b28b0c24497e784a4b8096f02ae6229c681d478d161675c3616355a3e4af29bc4
zee8733086ae035f61270e83da0056d05259a10eba259a9a87251016ca939a38d31808be4c54c7f
z45424a709b01e373e3d5060aac36e4b2caac9463c0cf88e1e52179ac785466e50d0c204c051683
z6979938001f34dd46d1db58eeb7f37e3128ed38744420fac98dfe6b75c85dac342287ffd4f4397
z7f1bebd234ccddca5af70c8d35ac88d7c91bdec1d04af7e75177e842a7b3c2a8847eac2377ea66
z09c637893a486c999bc7ff24151d77da56d92ccaa321a8ea7e2f8ba2f07aca55e1b949e89acc26
zf0bb622e36bd1b9f2711f8837949e4432fc8126f8344d29eb1497f91ee8b47a3cea6ad27f9b0b4
zd5ba6ed7c6171fc90ab2f925cf9955ddef8a73c43fb47a5b85911220b1428fde168c3ca7e57af2
zce7ecd5714acf79b85cd292163531794d556989b5b5fa284e02ddb666cf0a7665a23d89dcf63d3
z8724a1dedd7dbcd9950ba620064563a84e0f15658070e773ce468dfcd2a2a25f7539999221a078
z75c5c24657a872facdb29661828d1f857402ba57a743579ce23492d55afb068ac7f7156e6c19fa
zb7e2c83aa50a8ec65c5d55e2f2c00ad6847e4dffd53e1b08dd6eea2a53af89859fefb3423c5f49
z15663c5dfaed212d4369fe25829ce9cb2befd1d4867a75984324b9520b4151fc07be1effb4392c
z64a5fcb18a2e5d082c9023e66abe16a8f94bb5c80e94e9bdece6d1bb99886f2a3017b958576d6c
zf411de3a0adda4b7f3dc2e6e4b2a74a212867f7ba61f226002bd46afbb97988c06c2754ef61207
z4082eb3f386b0bda61b282bda5a96bb9e249efbc4cab386295bacbd18a16aa0d1eae8747ffa302
z60ed48c2f84ed0d9c5c1e691f500dc158935cc8fe1627d69155a389ee97e577f500f7c2f9bdf8d
zee3fbd9a59bc54b312ec753ee0d53f30c6497110055ada4782a20ecde3cf290ca722310c63f5bd
z8eb0e05b747395089ca5770d9f23ae741e6ec0986d13772be84c3d4c44c9b6e0550f397536fd17
z1c3b12907eed02caa4601d39812c1efc106d692f21822b0ae2940ff7e7896b032df62db15731ba
z854809f0bbcbd0de9671682ac96fc7e0aa636cba2ac9b68e892e02defd57158e60c392a74c74d6
z12fecb268641e6691afeb8f860774afe1a1de35ce5f7c2ec3beef8f9e5cb81b260dddf2d7af6ff
z135ffc54d2a27f20b3736856d6501368c88d329670054fe6f5a70a46d474d8bc4c6ae903e199cf
zcf998beeff63b4bdbd3f264a5e7e52a3e882de7a666a1131221b2b37eefecbcc4831a60a0feba3
zafb0a41a0a283461256692b7b18f84f079c9101238e477532953f1ff300bce9282da3e30bf8442
z6407b26700bc826b75a2848f96639cd0df33d544ca918445ff32d1f765c0a9a6104319f3cb16ce
z21852b490f6e2baf9393a1d1078a00cdb71357c0fc0fb8810d992205ddeb802033a148a98b549c
zaa93270b8af6196b25a9615354abd051aae668803caf34e765345007f1269ec577bf9eb5f734c3
z2997b0c74b5ff0c03633014b553dc5ddf81d52d5191a1fe38cd1a5cb9cc6453f1e5d5318b58768
z038b0ded12fdd9c7ff36b54fc12e5398b3a2956314f78b9c5a920882059a79db2243e65315c722
z88da958b249c7ebe1f8b4df80f13752bfee1a814a8e625be47a475f27434f9a2a4bae651ab04a0
z5812bb0c12909d2d136fc82a597c8ab31c92699de0ea5be49c5c72fbd1c77851200d01d24b43ed
z4c30131b736521944a0ec71f33dc1ab989073e252e071a393343fd8785490cd27f94b504839e84
zaed010b68f68f36b5b5204c2ff50dc879a789d173c83b9bc30c2b83ed6577c19edf60e82c9766f
z9944beb7390d4a14eaa48abbce5f7e21a44cf8d07b71f77d0563657cecc36025c25e0fdede9362
z4e25788a69665c0ccfc1a89ac10ef40fb90b9105712eec9c934d007886892197d7c2ae5a9c8caa
z83c1ccf5611ad54b07f867e1658d7a3ccef7fed4829b0d2dba6912971203e4c9c7b292c112387c
z1f75f94083ec587994d5c3ffbaef6e842e2173297baaf4fb64125036b834e88725ed8bc8bd43e6
za2de0935eddeeb49d71384e25a5566d978f77610a701c4ca3dfe71220dc1d2e0983c57593a2904
zb287f4c44eb5d4d7ddab3971f15c309326eb7c28c1ef6d32d8d1fb2198ddadf6ab1730c3abe5d5
ze105804721c3ecb3db6afc23248266a63c0563e83bd65660bb862ad345f62cda59ba4abca1cfff
z50525a8b589aa48655e30618be650d4aee422dd5bf1ce36e9f9ad2e574285c2f502556151ab461
zbc2fbd0df06cbfc2e1a1258a2086f0153c6dc99345a9c0881fccd4ec9214f03632377469b3606e
zf8b3737644b2e82d232fb77930b9430e77ee9905d9c584ca348c0a2f86b77f0d99d3e29437f8ec
z1d75382183e4ecfc62422f79f33da0e1553a13dbb3ee48e2ca63f3a01a8a55d8fdcd74d4c44f5c
z7a9d8a583546766955d22ece31707ea6c2cc6f60703b481e951eabf3cf6608a859735b668cf943
za520b0fa3206bbf7fac8ff573559c9685af59764f728f23f3093f176e73a6f339850927415288b
ze2c1a151202b205018c579a98982449af6ece4a4d3099a8f27d8b85e21e82fa766750e0fb78cd8
z5ae60e66649fec741fc7f7f3260462b8478e6b82bfe97735ab4b7dced5005965d378d732658cbb
z3614b9ce32f6025ad4304aa96f54bde37d5999491debd5c08722634d11f9067a82ae9df2848946
z542af4e1cf76ba5ca014a02f60858a5b3f16f515476f3fc3d184de40df77b92e3cd949594c5d47
zdf9d17a9be39714358c45089dcb832ca9e99e7a083f2e8c523dac5f075e0a2ed6c8e1e1a9d4993
z1f79ba55d8e7f8f81448d87f534fc74a7d9f5fd9d65cda8094c7e066617ff8dda03f49c20f2580
z1a06e8580b5f0266e874dc9a150d35aaa50b6adab3728b3a8daf70a9593a63f8798cd5ceda37c0
z156ea333c0b3ed178065be689b4b20b016aaf441e9df31abec024552165366cb3c6aeb864c1217
z3ad8bdac47bf735b9330ca85b2ba1d7dd34ce55d63c496591d6a7ee6be9cb51035e6c793c23213
z6aa89571bba51ae78557cf062ab24d785f65db6d5446c2d2175e096434dcce9bf7e48ddb77f681
ze9852176363c203445988e48d966f3e437fa00c1c966c6cd606a23cfda20d7936201bee1bde16b
z14b8939686d2ab16e7e5a9865e8a01e14e95363135fcbc9696a7650264b5d552f474c22fea52b2
zd2445ff98b5aa4e9fa1e1bc9c39953af785efea93398dc60a172ff255bc5d472ef0940d9bde1ad
za41a90fe42715bef97915030dab8cf3734e618ee190907ef14be6630287630fffaac7d087073b9
z3863d011f5623d87fcf0cc89f34148ee6ceafd1eb9847ef4c0a8c2fcd97acf64e4817768db0263
z7dc755e65f43a42fad90d3ec4324429d0a7b74c0bb51045044552b4588d229357661c75216c5f8
zdadc80405b711537778aeb2cd4c90bc5acbe97a0da2e66babc32af9ffc1b9dc1912241ef230d97
z8b3075cd219f87e48a4710d64e157b98cc5e929173e939bad59fd21f784e45e9e781ae39ab2689
zc4dc6e15d5d61a8d317d8e3a9408b8eb18cd94639724c2e132e4db1a5f05ffffec7ee5f9d57b16
z8fb644d534c64740274ff0d98fb035ed122739b31e0e27ebfdd3fbff130181ecc6e298a614a6db
z059958b18ad43da1e2b2a65a1ab8b24e9cb30dc43801587615aad262c12b31ef74b1ff50b5fb95
z55174404bb8592dc7a58b0d26fdf0650fa029009d714f43a0ef4f03a79f9a029885d143385659d
z5da7274bdd364f2c1d34fad9cf2bd2e1c83c746216596f22b38f6b6d17d13d2eedc0f10fadba40
z53a11ec04c6861770202241dd9d1b2bd3e52616c592bf43c3bc48464b981bbe9d91912eb18f1b6
zbc0c52d8e016dd0c5d2ac651ba8e0311c3ad9eb450e5cd85f5a7109c7ac9935446d0df814933de
z559e6f157dcd800ef85114404aad8cbafd2e525a9eab818b5812a5f5351e1712f42d3822297157
z5da4a91a10cf7240bfc293a04a054f231bc962492577ac48949d9be079dda3652f36bef61d5597
z3a349bc10511605ddf6fae9b2373e5b71ebb78d7ced7e6401b8e782475b776ee15e1ad1fe63d7d
z3ef12ac85700a479b4d28584487e747292c203325a6aff8312ac506c0cbc70ed73fe36a6966213
z8e786c9a5752554982f1fc78ca4bd25287e4fcf0021b5d5a539d10f757b4100f6055dff8494b62
z1f5d0869a7cd03d7203b75a69de65696f648688e024e02ed59ff5116465a5b07e117c093614946
za697fbe670199c3d0cd9b8842175fe87856a2b769c784d4912cef75cf17a2a185b0fc8a8d07e82
z8e512fc2498509c3006aea9099e96d6ce32172efe5a416c715a090aa849a28f5e21df5a557b52e
zc18e9c6c971273e3f85efa42bf32a67aa8c0705c841b3995382ac9c286b95022becbde614d9e6d
zce039c120d1a06c9f49c98d4648d7cf79fe685986f015291aaca980badf96fe7d8ca8ae5ef6c27
ze03e1ad30d7d476c32059501436a68c253d345a828ee65d9848d40c0f9903be9aa676be17f917b
zc22b0ddfa7f8e55da99bb5cb3f8ecd36469affa90417d98e44caab34d2238538ed303d45bc5b57
z643b28e083a6ce470707f6ace7e6c58a90729699fb0aab07c2febcac785df6334875462556f10f
zb3122981217987ea0090d1f28272d7e3cad0270c2bd3145a903c0f9f0f09d1bd508ac5f0da8ae0
zc144cc39e9da16159d931007d436467943afe945b8646c68da915ae10b80d46217531c8a2fb3dd
z9d20f29a5c2f1c129c4552411f811122d53557dc456960a1e0a59237ac92f7f01dd84274415087
zb1170991c345ad2c870c6d309169b82d8b02e03d8ebe4ab70dc0432e96bbc0db7208dd47fe471e
z112cae51857f3d9793ff1a2cf899b001a2567bb442b611a0e3f98319e1b2a9442253c773502514
zb8cbfb714a0d2210f7e510f96653a91848eabafa5fa6088e6866dc0d50985529b3857ce459cd01
z617ee7509f6f2d0db0c6ec82c6857f47d677e23f77a54b3b76829e9615c638241112fa76c15b58
z41847a1f6df30320abd18465cc9a7ed03fa82ab57d4416c0d7deee2391f12da8983ab339f7ef02
z676df788b0b503a525e974686a43c9da5db65c2146094069566c8524cb55ee0238ca38d02e2a22
z0caf43ed37afbbcfe8e6fb36a273f3b8da402e3a4970c18106e3a9de4fea5e2cb63e0b6f64ce3b
zb19a05abf13965fda80465ce542aa85fdb0192ea37bab12ee38985c84ad37a179b695a0f392f25
z7e0d77a31296c459c8cee0e76469050c57f47e901d29f97191c0c27672e1b0156b34956061aac1
z1d077e535f1cb0810f91ea9dd35d7fa1c45499ac156a69e4c6bdcad382c0b937d9488ea227cefb
z5357f181a6d65ab09ae3965a67aeee7c886875f49a7a851a59a14f3eca2d2c97d03b522dd45fe4
z2bd70fdfe88086ba9781ef3f1dba28dec93099c8735a7456b1ed54b28a99c711f7d844d78c62fe
zb5c9bbdc54af7467964fe393e1f089069fcd1832114b86d812c17912a504200111bdae80362a27
zf90dfec999b28656e89bc23ee7b63d7549debf308b70bd07326d55874ef7e167028b3918927723
z16bcdbe73b51516b2013888f2f1fd916a47a638d2091957832377e2e7b0cc7da0fdbcfce053376
z89c005a16ee946c387df5bd15ce5d412f85e658d6bede82f8627796372c02570e292734947f571
z7744d2527ea7c888f92010cd6ee55a8e8b872e8cff3bf6e0c3d8745454978fcc4c62c0931024dd
z0f69065d02c564566c5467a6bc924214ad94dcc69b3e95a420fad672cceb6aece46895d750bfa3
z97046d2bfa6a76230d9bffd3219e7651534b0b96f0283b3d09b98e007f4fe1f1443db9ff9cc63a
za1311f6e12908ee3fb5c01287ee64292625dbb8978d10b2c1d2af693a8302f124062931b04c875
z6b5f4c353fd831f13487fc2bb08e08fc9c891a89d6bb8781dff239b0718aa190ce5492a3efa8e5
za3e12cbfc2bd7eab28d3883dfdde0c7230952f7af966fd390fbbc7495829cbb8da5f6765c679c2
z6bc2c2f0cc7ad0dc27dbecbb73a0a8db7edd330b97f6402047df8b9ef0c32b54d45f2a1cbdfd6a
z9335f6643e619c671e3ca838984922ec69abcf644523cc93485399e926ba960e5ee62c754a65f9
ze12c0ff843d738eb1b031fa713503770e7b144c22cf96b87495ec7721ea1937df41e28ee070109
z6e146ecbb1a552ea38c8a1ceb1a5da7a7ae9ddd84bb9f05a3b06f88ed5aced77a8c7364b83866b
z919f4840a6ad3b1add065642b52d5e7a3bd31854d194dc85e26823bd8bf9601438778c7a9af48a
z0b2c82074cdb95f1ce11d56afd134ecfb12edac045ecfe87c86628c450c6e3d17d08e642f9ef41
z3739ad07b4a0fcc3bf5b23298c6e465f09340f8010bf1ace178a3d48412633528085e361628fa7
z9b9a2812b72e5c95b2bda3c9c05dc0c6a0296105d5af2ee1158fb8d1bae991dc1c1c89eb3b9f99
zf086c2e752db0d59168a0d6f7aa35cdcea5ef738a81ae3970792e022fbb15e84051b4fa944d086
zda4b3d1aca962c67a40026648e521bf14fa7ec73e1d518b8d1caeb5b4037243e3bb5693c49e64f
z737e7adf14c643b340ef4a9b29be57b6e90931e72f5181e09ca7451ec2ee29931217f6995207c3
z6e225f1cb99dff19e88f62833fc576e9065a40dff6b79d90743e065d5ffc1dae5e27972357a692
z3ecbd165f31527136c0a5b90c9369e0f2388f2ead1c49dd09652c64dbf795b7451f4895bd20ee4
z3d77926cfe512d9f173495cb7e0fb91aa06de543cfcea06621b50f638736a74f74c6267efe3ab8
zdc5f3f434c640d65ea6c365423bb980cb288474315b4be5c3c140d583d6cb9287b7d680ca0b175
z1d40f809f229d283f78e05b2dc8062b5f8621b158cf74d7cdfa676de531afe7681d37a4c427db6
z83029298cd288762b112a5974fe4fdd1224b653ad9bb86bd168db4adad2e31f8933419ef74c509
z78ae8765cb8748da1e5b65f87fcea05a96488c33d52127ff0c235e6679f60489ba89166d567a57
ze768cd22a3781ac04742792e7adb25d8d3206c84955c28e1f091588919d153430719d19ae9086f
zadf906c6d972993ab876acf7330b5f6dc7d36b6b120c5d2ced78f4fbc434e63084658e206b5632
z251dbcd821342e07e519d0645961d5d38ff127426f60186bbe531e83b388bea55d9c82b0184553
z55b020f0aa0f8c8b533adfac0a0f15897bee66b7db0ce09b4163fd744e68f84e67c2594d1e6660
za0d1956c55f96749981ba29f51912a8096110b05201be687beea86c8ad41f1763949bf3b83c3bd
z4d52d8ac02b03c9a54e1fb59fb1c82492cb644948c845d69836292bb012a1844fd15f9bf6ae3f0
z6e6db5480a8fc44bd1704c6de91a263c4ece6169a7625116bf11418c4978149de994fa762f73dc
z4256b9d62eb271c342432125da67eb8d26ab46f398baaec112432e6b33663b678cd55989e7fc60
zaf936d8958cc5a54ef7d1c1ff399b73ce8661feeac9e32f3bf86fdb3b713b319940a87301b4ba0
z68985883b3ab50b4346ac1de0c1dfe4560e5760c060070f208b2982f0c2f4c1855812328b54f0d
z9ab495a00c51d5fffe3cb18798af4c519a9299741e61c80ec79c8ece36b792ab3e7c5cc23ecd00
z89393c0db063f0fe9a3a2c2c140d7bf50ccf686ec311388edf25152295c96bf1ee56284f004a24
z1ffcd0c218f1426e6ec92755640965591151b1058c36bf61794f050084204a82c81966b6cd3ee3
za525c02ee63e22077afcf04ee75ba6ec12bda630a2c3839b4885ea6cedd1994a54f9b23572ce64
z8adfddd61f9866758a0b5a3cdc88ae33fab9e6dcc73a5f294a48a64b421877418594a21c637b2f
z3359f05fd43cc9c9adbdde5e3daa981ba40b28771e0b3f27fc69fa5b182499a89273e5db620451
zd29f17b0f1245964cbc0b9b02354cf99b08e877407c5d862c8ee3178032157464359388803ebe3
z8a06af9371aa84b576f3fd4d16f18855a90e1e9cdc8714e79bf376b2ab00994b1e9d1e5e2a3ed5
z85a10c7b47e82bdadac240b1286106c8089479def1b7e90fc7a20876c262f87c804487551b4f16
z41c62627d09aadbe03e73b9fe53466e7e8a02f740e23de492b121af99772ece4aef24e86531f11
z59ef9799e72749b5ef8fe7f60ccacf331632cd50ef81057891d453c22099d30c9caab50d86db7c
za1dd01a0e0b17e486c6e56f7c95d5427ae51ce8ef70c3b35e0e94e0b92b81350b07483facf02cd
z35f84af665a326c0b63f8ecc7974c25ad7d6a64fcafc35a3e8a8d93ecdd31988ae4b08eb22b2a9
z3c171ec4737d687e5fa6ca1456f35e11b6dc71367646a78f668500e3ab67bfdc6335c43ec11ae5
z4dffeb29843e4a1fcf937e457b793da57c85bd0caa595762920d38e61326abfb102954fb188409
zff88bc361fe83c94bdaf75507080fcbbcfe92435fba449d05e371b50aac3563f3ca1ea3e34c0b6
z5216617c077eed5b717a3d33909bbe74f91e5abc90e13cc68f912d16549b0631a61509b9804ced
z080520490c20bbff917f4fd56273b458107c11df1278167464f79e8d4bc2dac79ffe921048cff2
ze0729d1d9fa67a1ac4395443a274c59d1dc9886a4e3a1ab59e01aa0c781aba62d57ce4f207cf31
z92fc81907314bd14f14bce5bc967330d0dc5f659d76cc0f694b069b067739e3b2458c8108c77eb
zb2857b7b7a67c87b7fc901c21a7b462a90d73c5154a0639e88b7c729f1a4fc89669b9493edebf1
z1751b2851f485dc6dcd6176bb9767636e1f65a52e9c47fc9518b4454f8e493084d357227f47a79
zd9379cfebb58efb4d0587b474f56e12fd177efe908235968fc7bcb68f3404f6ac31e6ec63ea9d9
zd2390edbdc7b32fb8c1d4db62252f6f312ef4acf0fffca9df241403af88ae1552b2fbeab62c865
z5ae0e7327612021fe813ebbf3a1162bf12b2cd17ea1f95644d5878d2aa00832aa8b813aac0567e
z33e3bfd0ace2ed9538c3782a6c790d03225af876e49919a679e2029be99df03cabfbbd8471ed7b
zb20b5a07f8eeaa46e1eeba3d04e139022dc2ad3056c216cdb1e7007daafbbbb9f5ab0a6d9faf93
zbad33078ac06e3b521b9bdfc1811a38aca4047e0b865abc03c84229b77483688cebbfa32a5372f
z3b52fca0d0b4fe3cd54c36067678c6ba2f22c65d5cf51e3d2551a062e8a40d1062090dc8826868
zc56d2c7134d80c43af66d0729a4cd191ec3bec865f9c9df0f59d40589d1c963b7df03701ea2338
zf48762262bd1ce70efbe6da33c01a73ba320df5a7d38dbd880c067df625fa74ccdd9d8895b9026
z87f82c7e07d93f71257e0099e38393e0d71337a841311767fa417159342e89f90394f18bfafa08
z691bb04e94a17ac58ecba68fadb62e33721b49972f5877d4eddb9fbe29538127207e7f745fcfe7
z48319f11323762655984fc11fd96df745aaec84eb3ccdbe6065334f8035f535239b573cc637405
z5c7548f0326a5d12716f5c0d5bae79b7a20958626a9f7a74a9b395e59577fd1748a4c37af12cfc
z3461506c219f94b81a5ad09eda645e0f45b54d7184beea17d631e38306a25c4b8b45a454515810
zfe5f85c9ee864f542d480d3784e72dc2664f95a786bfcd182c62246ee2207383023504f97e6995
z22d580a9fb30b6f9a29fcfdc01e90d327ef925c0b3354d49b8cc3488fe2528d017bee99b09ad3e
zda46461bdeea2065a57c8982974eeff4cfa400cbe5f4786ec9dd44f595eeb727ee19d2460af844
zf896841c9881c7fd8f7dde8afc46bfed47a8c5020ea6ccb37371c1fc3f69c93393bed45a64613b
z7a62cba2c890cfe415d7b05912611f3f375a1bafc0f3d282b34c6b0474aaf08569d7a6186b06c0
z3301051435401a09a069ce5396b6cb0f3ae630be8146c1999e1324917856d7d5edd2fc826ed077
zd232da1211bdf6017e8ff9420c1cca382ea6bacb00a23454b51288f27375aa3950ebb8aa508ba4
zdcf24421fd66cd7a07d11db7746823e07bb04d69b7935e19327d76ec253a6cc8b466feece98b21
z4e598dc4a42b1863113a2cdfc3d7cd3e6c5fb42115c79ee6be23f53256c77919be62dfafe152dc
z814d83922a51e0d7ac8f4b506d39bc8e2d0a857a6f8af21284ef84f9f070b45a4f8f54680889d6
zb0ab0ed6e6672fc4b05474d7b29069061ff91db9fe96f8a7678ada821f801731e73bd639374204
zf9d2eb43644338329eb9ce31b91a6d36917e624ad7627b1381aa768b3f080fa1e3be57d200a920
z6f20462671d398de330d1be5a2351ef6075511dc18af5784d9530cc1113daa86fca0fa0c6c74dc
z37ab13aa626fc8dc02ae06e1719491b1bb4ee833f83e08b98ec9de1650a8e0d11015aa7389d733
zd67acc4f58f715cffe736c7899a1a91a7d96051fc2ae284d4855b093ed3159ae0f951872740940
z2fa4d49fdbe5477529993bb1bd0e65fe45e0fce0120f2de4527b55216fa86f2597fab42cf2c81a
z0961cea003b23f77204c10d3ba21ddf5fbcb98f7bc4903834207a5a690f696aa8ea87f2e7b4b5e
z484b19a24504b52a050db009a348de8b68036ee7860bca22f4307d8b44ddcb31f798fc9255db36
z239d742a28c81b53f345f19762d7aa9d2ed618dcf8ed42822d305156b99be1057b2048a31ab92a
zff21342cd08a106821c7dc73cb01d6c27c4adcf133257a85ecfbeeaf360509075064d8d2d0791b
z98ed8b55907e129a3fcfd17d63644929541ae853e6a5c5890774d5017c227b522fc5b98c325dbb
zffb9121a8cadd158f351849e558cf9d721f9b6bddc82c8f32a2e5f1571f584e038f5a510ddfcdb
z5f17de75f4e5d0bd83b2b812a7f9d78fccfd9fb5ae7a47becf7317019c8f2e752ae89d44c496fd
z6d1257759778301f9f63635c3e6c954a0aa6f9675db6dbf13a7ed19bd9b89ac11ccbd5758268ff
z13743eaabc233eadc55be974f48b77dbe0f319b6b0d7d4d4a9a6ac3d1ef3995b0fed30a54026d0
z3598c5ffebf1f58f41c9964405906a2f29dcd2fc17d93ea00e578cd6331a467910a919f5108128
z5123158d90d82a9504997f2ebd80355da5ce25b29c09bd0ba1c1d5ba3c3268463343f12a66cbd8
z87e9a1ea98f7df2619a6c79face7244d77119fee27847ab87fe8d9a6c2ae6c793fb3abfa2274cb
zc5a67dabf44e3def06b7b50c3916585d6af7c9cbb4755701bdacf67cd7579dec15f3b9422886b3
z222f92ef637efb60f9ee9e6a128397bd3e3ea4305a97395da38cbdfaddbee1756070bb44c6c41f
ze8bf01a86608df2a04b45d7fba858428e8a16fb45570e0549f2e3fbeb9599272673ecf34b85dea
zb1689756019fb8a44bd045f4f224f98515370c33cfab3d79042bddee3dfd4290cdf43651b0287b
ze99d86a32d3cab88a495f0f2d148935e43c3a35bd8620c6c8b8a98f850bbe0da22cfff2cabe80f
z598fcac5652d8d726486a50dcf2e000391c571ced4dc6fcd56b40e90e4edc93cc070bfee1f83ed
za902f4bfce9730df35762acd08ee17b8b66152f10fa2b9d06cc3b13b1dd0df861bbf46164e5bbe
z97a966b7e85206c465cfecb1a134393c04e8315a6d3dbcc6a63c78ff559497d13e38b323357c02
zb2d58e7778ee35c5b0bf63f84b96a688dbf4549d98f6daa3bca3b36c0dfe43a12ed5a753c52f5c
z1e5a805372fe6d4580a5ec8f4f0a7fbf2fb4b5fd33c1347b986b9507b678394925451150809431
zf7128176f43b01abe1c0ff9471838c926966276ef8b6bba1aba96f7310d3f244b1a298961a086b
z3ab607746f75ece12fa115574b8e8d55e8bcbaa09dce78c63eb01f6da8820170f0f9c0a2fad8f6
zf6f4f0f7ab34dafcf6cdaa98ee2bb3fab91a63607a9a2e736e43d342d87ebab2ec2fffe34a0c67
z6c00a7158b56e4ce27a3c7a593e5f0b47c749e333de57aa350054ba6c4f1decaae741700033e79
zf7f5957c8b8c1d6d5e261df27b1577eae7147b047551dc75e49699b11945c31f77759c93435bea
z5177ff8f6289c7e835f3e9eaa4d05b46ac6c6b371a2be6d39eb7faaa305c5e3d56a7161a5afda7
zd9a7da9be1aa7c11de7584a37007b3da8153bf8d5db1e956186c021872118574bd405bda74e6cb
zefe684e5f398ffd87ec4097fae961682cc1cfef57ebf0ba79535ebc8e82c618491b9b5d134ffed
zc324f47ff4585e53734e9f387ad69e47f9a60830b63981b49dcbf41ceb07926326c8f04c9e10f4
zab50bc86ca8c2aeacf1372a4fd940af2a411946f9013a620e4f383cc5d9a2db695eb3bae5156ae
zb16759b57eb8f2cb3efa30ecbc23c8bae282812dd1c713becb1aa53a9d1ae3c58b4aa1421a124a
zcddf251eaa196268c234762c0fd897fea758a514a3806540745b8718ac2994452aa2db765b5726
z8be6c2a298b022c00e642eb6b3d366ef16f20f5c093afab8224ca1e28395deb8a3b6773e7be887
z2061b5fb07346e167bf1571db38508ddc1e61dd7e0e08a2a4e2a22293bb5a304afdfc4edd8156f
zb2f99c98281feea2c36499e5ee30abd7bc9c1565563c49cd9688025c7b199768cf82247877f6ed
z5bfcbb889912251c1146a2665501d4fa351b5b565dd715ac784bb4b61035238a80beb88978e945
z0ae5197f0f306f1969580978fa95704ec3d375941a34f83dda00af6820cf096daf2061faecd504
zb973d1e6d62c5687cf516c5f7b1baabf4267f93ef83838a08e505afbbcaceec269bba6af031e29
z4487e5b8d75b16ce7514b74832b2b7ac5297679671c6acd88589fa9e1500f1ff3bdc611448cc4c
z300b84b849a3a5f67ed8e2f2d53ae30d5cd1a61f864ec926f73142da1c74dccd87f6ccf83c969a
z7a86cd42b7a4dc0cdc7064547532e0984cb09c1a33ff8480fb0ec2517a02c31e0ae4e2bbca8097
zf46f13aa14f1098e407ad4e74736f15fddbf12124c3f52e7c90af0162d7af64fa78bd1a55b2a91
zf49ebdf754f8fcf12e039f8a54eed9173e8231a85f8f7e6477c1e3be623c3a5553cd4a142a5932
z0aff86dc4692b0ffe8b390380596d690c11a46c2a5220677b275144c500f6997cb71223ab43c7f
z64540e1e8c7b848bd839903bf3fb2b8df12fe9d32e3ac44ffc2418fa47d74c44dab9f2f3765473
zd6feba5ef5d32311dbef3a3aa9ce022faede0e7eef3802542b7af9dcc0ed73a4cbc82921950f83
z922f5fd5c15c5d6be7783daf35f88d95430da2f2b35f82d853d3359dcc8f5c1315d7bc7bd159a1
zd377193aa2b616af0194f20746a202f66df9855f74918d49ec203b1a2865dd77538055a1ea4bd9
z3c202c0de4a42cbc7aecec5e78589f348afc0c4634f8a1b89fccb03f31a0730b042e7540d8d82d
z3b6b76246350327f0a7a5caa6b2e7cd08d7e3574bfe7de684f3ad0b7007630b13d0b32c63b93d5
z9f099cf0461cce116bfb17ffcfbabe94f6684847f9f74b92b757a636b7b3f27ce2276bace1853c
zd4284466ced3ec87659cc9cd4ec8489aa86410dd959fb2068b68c7ed776d606a52fab38f86f773
zca5737ab32b084265bd0c97b396556f8dd03d5a7ba01de8d44e7ba8c6dfc48e590d78577c73f1e
zc14c864d625dc0c10e4e4ba18d6e1f413bc728a6a13a1bce2b6b7d3a492af94d882fc1a3e92dec
zf35d6be95ac32bb8c039b2638b945ff05e36ec28276d774555f3a6411eca72b9fe4b4d6f0c363e
z67b63e4e23f7d8c693f0ab126b77814aea410297ea6f5788cd7e0c4b3983764bdcc4ca78004600
zcd6ac26795f74cad74631aa2126ea200da382818030bcaf8f82229b3c6389e4f618bc4553f34ea
zd786da489269876f8374f3ebe017718d5ee2e441cc952a0a6864e7ee8b5c83abc785a728bdd9e6
zed9fbe19c80099c35e1a701d48dc84032f4489d7bd12616a90b95bce0a00702f4f780f61474ecc
zccecfe9923d7b3c19c7533c3cabe926bd5f6d85f4b5a1b8bf1af56790b1a4b90f97bad6014d571
z7f4b68280e36b7d23ed63b18899e1917a46fd77f325ab8bf17521852e1feef003c85983b67314e
zb37c06691ad3afaff323af0f78acf4ebd6fb615d97658dae57a1e885609783d6c61653857f468c
zb7ccf6171b41fe2f44db789738efbeefa4d8e81d10a1b411c3596ecc4db97b06cb9a5c271c4f28
z4dcc1e410b3c0ff812586ea809a9d48ff890663a44c5393d1f7e876d21bac65379d850e55a84b9
z838ea3d8592b856dd4d15983332bd1fe152911cdc2fda39146aa71ff8ecc073dd4e36d5610a131
zbe4036aad3e3a92f884cfe567855c55bffee90d4b4986fd3e523955361e60876ccb2e78ead9cd9
z5b47f93f223e49091a9a7bab761c2bcce531eb9d64f846b2eb0205c00377f3741acc8b1347145e
z72be0140d39d2d2a884e3f5bcaf4bcbf5ac0724ac8e437f774d1b5c19641497eaad386ac134ae8
z4e22c9fd4db74cbb1f59c00f58413a8f049845b91605295f46c6b67261deeb3ea2a5b2f87b14cc
zef0d52c9c18fb1507cf84f28d7cffa6c9b8bd2266a0f86e3c486d1d7b777056d7cfbeb5619d780
zecd04e35232e8fccaf703aecaf3d593e5af58d40bbe102ef0c395a07f94de0d98567aa7ccd3cf8
z8263482fd6a351b88f127c975510ed9d3b86230a67e5c78d5e6ad964ece5b217fb3bfb32a58254
z6ddc986e5570a9c0c8dd2a216000c9d574d746a22ac3f6cacb92c73785406d7bbd74a6414e6367
z4e9cf3067a01d4a843a4e5b6a5c629efb983df36fb07c529eb7b3fb9a403fa7adeb72754e2a5c3
z71417a558d25823c7af3e830d48138874c8f07fa1201891bd0c5634e56c8414fc33135716bca8e
z57441ca2e460f9c60da70cb6e6ce28a44c51eea4f40dfa6a65064566ebd953ab520775298af69a
z3a90f96b73c04f3130134e9155c56410ed4e34729fb8675630ecd6bdb78995ecc37c221d63f6b2
z0cff16d073d174f92148fd37d73c92e1f50d28593018a9198e8aeb9c3ff65bc3b33348c14b178b
z93e4dc40cb44509d97e908adb6d338a582c859e3a01612c7684d157b597d634600105705bd8b88
z7856c25193dc29c3367465baf033796493c2fa0d963378f9c5ae413b0064f058da7165d60fc07c
ze0493f6a3370c5954fb0e5361c6c84e6af9e6af5d81201bb697b0e83b4552e8727103364c1f540
z6b30dea7f0d36023a64fd507275d5af9e84623e814f407184ebc8c7941317480fb53a9d4d1ea78
z450e45819804239bf1aa56bc12ebfc04cfaf27b268f7e3cadafdea34df4d43e5fd0f0c2ab61cfd
z98c4e5ffbf8fcb4e985f71ee8ff2bb173d3f214a47df3963a739fc1df81e6494a8a3bea4ff3d65
z6aff02a8bc4625a48d62389b80f1c2715eceead567debf610d37911e1c07fd8ffa8d06061f7155
z99c91176e3c1fa61e03945a3396e621e59a715599d94df40730ddeb0a270f8ce8acbc358467e32
z50d9f495745243b6cf0ff5aacda4909417ab8356f1de61e836ab760c6a109a8c2fc0fdc1a8dce4
za3f236a01383e3f37ea1b6b0f88e010ffc60977d0a9bc1de9f67ae7704e8ed07b8735bc92fc87a
z83f680d4af71079aa660492eabc4f56146504109df711da061292ee12ced27bb2af496ba28310c
zaf8ed962d142a48a354f144d47e7de517dcc683cdb677c660bbdc23feeb6698f165ccad7bfb972
zdef500a16714b97b0f546ce81699d5337eef02c596ea523e7ead188e1b816f96d339159e5b964b
z78085e51e46db0846118b9a7f6b6e1a81d902c9e782987298eab4e98748430bc3fc268d0240aa8
zbfb219954d6468d49862a211cf96e4f17389db281b7cae00628ae1307e95c7b9d32b24137e9321
z2c4a0b73eada65178a75dfc3a17efb3591bc53e1cc3af283e950d4ee19ca756cb16f2e279132d1
zcf496a8661c31b860b3e2288616e50809dab208d7244fa690bbb82792bab9e2c33d1fe27aa304b
z6ab67f07b8ec71bdba8f5603b296c7d78613abf3cd82b65fa0fee53a18f9cb671b902a3582f05e
ze56057be43f54da846bb6f123020016620f96410e5af594733f69d43f22b0c204be6e150337c3b
za73312fed7dfc202367895a65f216207fe74f4c41baad96aae7537c8e2e3922764a6fb6f2f2621
ze3365920e5df71e63a15606b73ca05ac8344d002f75770d4b2a28a5e8ccd33c9a1bc39e4eee954
z8ee7bb1fa8524b41bca1ac5af53726f55fb0360efbda5c38fb183709377aa9bab50bdae8f05b24
zf1fee79965cebfac61875f0ce82fddffa7e711656eaf19812d8f2f1de07477b0d29ef006692ed7
z2749304000fc20b34db87e8e4a90ea123614f556483ff8e94966a6b7928309f2e69649776d9d7a
z5fe37730439bb7c7c68fb781f2a68d8d8eb4a0a5a7adcc1d4ed714214e14d32170d795492fad42
z769e8a3a12e55b31e32b10db4284957996049baf507e8d2e82458bb400927ac18d74f59c75098b
z5de1fbe2b92b37df4568fc03a012d4c0011419d083d9cc973ad469ae0049476d1ac0443c2b056b
z2ca7c5c2fca70fffbbec3a55e60782423b229890b432a86b77e558af716f02d8951cc8118ce4a9
za4344d64cb138af421eacc076dde4cb709194aa3281114dd6797661aca37a4bfc42049b56d6efc
zb3d541d564276c012bde8026134cc02c72012f8d78388c868b18ca95f1e4e8db815cbcd8576f27
z0b604ffaee0da0dcf444bdebc6fdb1a1ea6ec781c19219d578a5df48a4bbb8e6d4c98a4692b555
zc9133fb0c4466fb63dc23a0e1ff33d975edc20ff1b185383067a421d19b46c4217d42e789839b8
z16bcfcf3b7d0a4d35bfc0749eea73fbc9e7ca634fc3caa6439af9ae29e0f0a2d7bb43e61ee25f5
z5dca09cfa3908463e84f5f3fb15cfd1052fb5856a5fe3cd1b618d648878b0975d3851bb3736a27
z4f9fcec1a392b250e58406b5f8e1f1e271787d322db73d3003af0694bc4b1f7c2c542064fb4d98
z171e8539097954777fbd09c01124e35e563064e301f727672f2b87ed54acda133a0af5e81819d9
zc06fa8d4ed48108bfe42e655e8398683c455231349a558711805ee8642baa0c9e558a5597d97bf
z67044501ea0216b6cbbaaf14da02cc61f2789abae4f7b5d463db4f1b49886c206376c72fe03286
z213474fd79aa0f41a4fd46ad96684b608ea82016a8fb24355ccb705f033ff6301970042b000316
zec291ca098e39918fbafdbd06fa0b804c9b121aa56a1d00ef83cdcf09c9adacac83c0a26b5e181
zef8fdf7fa2681b3a22abeb09412775518a69168960a2ebf4759f96809b9d63a67dca933b58d662
z728e2f910468a31679f50670c601cb12e52566f86362bfb767b0ddcf9acbd247a8dc90aacafd82
zea0b49f09fd2f9a782c654d491dc644cfcabfb9aa5782e227bff47a91c654ad96c6250014914a8
z4167079b6792cd9a4538ae305974faed3d8c731481003ba4f19581cf3f1e9b2c60c8a8dc28d9e8
z5257d7f5236e7942113dc1dfb4f92f1e407900e37143a35a487825b5e2efbc7c8e8e70e7324b33
z2719a8d1bf8077b8991a6a00f42db204439ee6678c07d883a1baa08b04e80aa0c89c0d76497030
zc6d0585db6ff07530a684dea57bc21b3c29b97147501a10f6c6461771e95d58d78c95d2d0bc68e
zddd13f3cda06aee6017efdff9128ecfad80b9d20c94ef6784a94264955581fd84ddedc30ac11c8
z06784c862899160f201a6ca57a7057b11d94d54f83c9e36add22db830e3e9679c675142bd19b02
zdfe4017c2dbe3540e743724872cdf09419a9216e116b278b01124a05a5821566258e319c829de9
z1f630e58c9ad2c10907c7238f4e8fab05a9f6084978786ee5efe52ca68e308a59b5a2301f00a5a
za7a69514ba6a7468929be88f85e7482fc7689e41395028282e9c03447afc62292c6b3bf7b551d5
z8ac13def48071a359e81c20bd5b452ff08689ecf6f96d9da84adba192cdd54308b6ccce6797f75
z40e1c418e83780f2d88964a6a60df8509810c0f35b0e4e9a9126cd5ac1f2e17f8d2f2aaf444c88
z5ccb7350ad7c0837dcd76af063894a5386d547677968d80fbaa7c69994c886b818e202d5095ff5
zc013314db8ea949703ba3709f48f6c0c71c17d9a500b77ef31c3baef8c7e4983e46ea9e6d577b5
z5e053d754e2ef92da2df3b8d265650ad5a8b1ff1530f6052bbaae08d978f02ee406dd643660875
z39024661531255fe56d268ebed3a0d20515a8633b0e4c39f57339977a1a399bb38c6548cdc76cc
zd03370d05cd96b0c456904210dc12b99850d61b4a789bcd8ffe3c686690e0c77217c5ff965094a
z2dc7e1a24f26caa57ab194744c96653348777ba702ba373b1a8b2a03061591f9e92b9409564285
z1c05c45ddca3b981fbad4e1e890313167272ebd1ce79a6eb3fe086a4e5c6876024c31ad953c2c4
z7f1d2c5fda1ae87c805e28d3f3c2f2a0b0aad61034bf5e3aa7569a0108aa6f1a0ed56bbbffdb40
z923f83935b5c61763e713f19f4e13e5d9ec3427409e8827d4bf14867e7dc8cc1ea1af6cdb1e1f0
ze27e5ab81e0d4a700f03411d24e1c9e4f722350e34ec2bd02df06450cc905d6ef20ba42a40204a
zefdfa50efdcdb0901c50b2439eeca331fd0f48cb4a7f9a3964e4fb2e592e6816798a0812784778
z8a92a7e0746a6c5fb9827e36e33e3907d3cd4a0568179dbb06eeecf68baf37c0025fd99a0721ba
z7c217fa7a1e9234551a1721c6115615e98b07745fba3dbde02e2f6909c9128cc84de2471c69971
z388b61d2b72da58d3492e17c2fb26352fe0f95a9180b7ee1a84b94d6b1072a88467bded6669c27
z4e1645fb51fc5223b3664701b14492410f06cb96eb6fc72b942873338861954e42ac869ff6092a
zfe6dea17059e6211733c76c5c555a2835aef42467ecc9187eec255bd1864f13c6ef1cca7cdb349
z1682326e9c77da2a7c1663ebae438a2be8c446bd4410f5ec5f304ed4cbe531bef673da74f435ca
z338e36ff47ca7fe1f83495d8c73445139ea68de07608beb19b7b5c479737cf0f1719f5ee849534
z7da71bbc8afd796b6f547c2227c9b937a472f267a99fc325b0d8287136bc2df3a33e405bb654e7
z7f7c29a4e1748425aecf645f61bfaccf85fcefb37c3791f37ca92e1fb761521ba21b5d57c2d8bc
zb22c091edfb109af753723bc948f26a240ffe8e8ec58b0bbbe384224dd82f24c1b5eb4ee9b511e
z934b123a24cc8760ca8920c87432ccb9337b51e9dc853d44684880a38c7b141b7cdcf9c126a0e4
z4786cc7a1d36debe9f4fc1f7e1a71d14bc7a833ca10e931d5edebfec09589a682918611798da5a
z3655fb46ade7c3e8b89ee85cfa5b59c60e6a62393cbacf55abdc1fe6a160300cab36a2c730d9df
za52a09b8be2ab13167c896f58124f7e72cf8f4cacf4505e4f3274cdd8e9e3a5b8bfbaea04622a9
zd32a0116c7a326b2fd623b43ceb3f36a6ca9ccaa0f0cf42f5e01d54a276cc6519d729a4039e151
z73a1e6a9434f46c45cbf899c9e1dcefcf91ead7f06d5f7922a051f409b944f7ceb5de344da6f9b
z0ba4bdefd5db30395ff42267319fdf3ab0a6acfbbc762398041785e741b44732375ac78b669351
ze641e57d59c67d2bb1767fb2d7d000f89a96fce24030542db602ca3c939ec21ac8bdee31c3f1bf
zd84fa4d11c18967a39e34f030de0f4ea2e26e3664fec7c94287868528df8f8890e406319d7d6f5
z173d7b4f1eac18dab03d6f651cce1dbaa4c76022e07a791f62d0530e6e145859ec05ceac8f86d4
z01626651784d95cf4e4dc55d234e05af41d34cdf0ee7905562642bb7ac2dcacf7c7f6674cf673a
za01e1f8f21f627831a1e05bbb2c14a837ac51fc7fdfe114a768c0fef6e853dd85e852d73489b83
z417f694e486eea17032527785b10976625755c544c7a1522cf619bdb410fe4ff2017cf2c8a2644
z0aa8cb5d27dc464771e248b88d821239077e6f46f40e66f9b5feee3b8128ad2da0ba9f4e7fb073
z766d70e5ea41e25ce63db7644949667888cfd4c6562e6b8bbe4da8e639d7f3752d80ce3a2924b1
z32186188d894a9578533e9b8affc09a8b378f475d1ac32d790a1b0392c564df974c313b8a557f7
z66209c885a9639eeee902b83525ee9724939644c3b48a9422d15d8d97b6f2eee0294f370c50b72
za2fda8f68ce89b006f9d67577f5557d11348e58aed514eb30d1ff8a4c88d579d3dc75868a8b8cf
z54ffe797c3b7cd580deee52e703ddb661ec97101dd4cc778dffcc0b86abf2939c6d9cfb588255a
z3e8477c4650a7b309c79e55ba8bc02cc0581886bfa8573cea46a4eb3badd83b022e7a24f2c5174
z61c88c4bd7e385f46418178f165aa3753cd6d507fa2d4c4d0c4ae34f05d3b43f0da4cd172b022a
zf66d3f86368711c1fc1176dc833fda5abf7f6481a6407f0f50fb181bcf6a8ff3e8c629efe5ca80
zafb17cf440f20e2242c795fc45958ba7fb6200cd7fd132d13e6ecac64c94e92fe5635af5ac65bd
z8037f54c58b0e28ad78009202bac9f75e4db392c0a27a3af7ff5d91f07b18fe8462396fdddc692
z8c8f92a4ac36a901d2810dabccf393e219025514771ed384e5364c045d28f90c7fd6aa7a64686e
z227413618d4cf2da1fc3842cc9cce945f15bc383a9b9e9be783e47a3dde3d2f397ead391410751
z61094aed4dc1ff9490fbc0bb5ab7373e8107b5e3c7c58550e422d3d0187546665413bde7d7f833
zd4f9bbedd9f650dc22e13774fed78c22ed0cf405493ec014cd7d75e649f75d8752d5947d2ef82d
z1d706393446dc457bab52cbdae22cae476b09530d7a5d3ddb5987f27ca7fbc89b61b5568062bdc
zfc3042dfd19c03e60e899b3bab6822b3a860bd87e208dcc5f26f5cbd3bd2737aef9a9bf53ce69c
z946fc6405e70444c1000d5fcdc73c78caf93498984781df557fbad82b14c4f94814c7c20609e03
zed4a69d0d5b46ecaa7f400fee0c99e021d8178079ff1b5a50ad40e8f82a46be53a43209f094d12
zcd0178ac2a785d64e34d0fddf8e680f15cbba75a2da382b177ebc9df83827629c63f885d328464
zd80c0a0656cd534aead617d07196207f9d4b2a96edbeaba1ec5273dacd26b937ce78f5f2e59799
z25b813bcb17c4365a28c28c1f06ece8f2da83a64dd7138f80dbbbb19b5a39363e22cb9acaeca57
z41aed70941e6c5f4756c2a5c364972676f906f7afde6ffad3caad10b6612ef497d02dc93554d85
zc0fffc974223a86f3bd4bf89cc800c99705d2271f3015c00600b73bcfc4bc3853bd2ffd7438504
z6c64c71cc5010e1606af67cc021cc5ec5dad13f5a6ee8c5989f79855a624c53b8aac2efabe3161
z0623f8566d6d8fe30472c5c5279f548fcaf6484958c1dac7e85f5a1132f48ad67dc4afe7b24626
z33932b38e5f689cd62863d84a7d6b3fa6dec0599b67875e424d98b1746437264823b48133865b3
zc2af1e6ecd37e2cb8d24ca53e3f3254a2262f2988f0e7ddba43b9665409fb79966fd1c27272239
z5918bf2b081dc3887b1ea232c8d53436d0ef6fc4f1cfca851b7ebccf5b781e440019b3ac6fab6d
zb1b7d8a0272db3576fffbf5e14a7b9739abed0fc838419ecfca65f0599096cc6201f2ca5ea843a
z2fa560665af53d585fe9022767afa149481414b10c293f57da839e010ce40f554aa5bce9f1a3c3
zcbe8f566eaa0d2d1162c3f3e8b669eba1e6575499c6510aa22b4aab25a5544d33a975d31c43889
z1819f839e38624ca6fec5519e3a39b32b3615adf00962a48d30d1f8f95cf45d8dfdac775d1dd8e
z54a65b5b79452348e57d5fc26b8793866977e77b33b8f24f93d6a8d819e334e93e9f95ddc4d9ac
z10d3e47284b7b5b09c6ebd9ecd2c579d18d2b0279ef067680e001eee5a451a84c8737d2569e4cf
z5c7a8fcaa28486e59ded76af5fcc38463d4f0a8b68ff7209a284763a01d2fe8e6a6857c5302cf4
zce1d2eaeb538fad362871ba42e80052241ea2aa28e9458b12c6a7ab0cf7c86db61acf92fa54a13
zbb9646639e81563716b51e680a68313685086236b9d79ae740482e67b3e58b9d40861572be5df6
zc3068645c332c1a1007f02393373d11b3ed6d57e8447e1482c07cf296d48c031273b4d9d605e0f
z52a736588e48d74a27921169d01f8002eddea85e31097ab71f6ba051fed4a5f1cff71401bae5d2
zc42875f0d2a4f84d894859160cac641ebb099e4987252d2e1d83bde714f81a54e55eb2e69a05f6
z3d39850edf6f816df0b98ff87c9ff58d4f2cbf55bef19ca3f49c5ee07723e17b44d134d76a00e6
za3d5ae098541d87c4e432565aae95afd4c8242ef2cca5f1a17a7747e4a68e9776ffa9f62f2f651
ze14055d86575861f27452acbec94676dd324dc1630e2b4320cc346f20bec07bfd136be3bc9138d
z7d034d6d4b685d2833c70f9fa891f37839e92a73a4a3f04888c1731eeadf06077415cfd346c61d
zcebf27379972b99783b65b93335086f83e67d2ef91965e4cd308d7cd595478eead82381203882f
zfa24d9292c29cc853ab24699b3420ce9c112d020ceebde15bfcd032a6798980347a8a6dbf0b241
zbda5b8ef133dcb9ba68ddb707006f8a34ffc3b2be4a1ad2a06fed3a92740862be2341d4511e386
z2b2f5c5168a0bc9f36a60c66fbd91035bde71a4fe989eb213e75995c5a8f6abccdaf2c49358bc5
zcd6a2c15c08b3358aaec9bfb8c6324d4c22beb9225294c10c4eb2fe5fbb3e29eed7217b0bffbaf
z464c805666da0563ae30de0b69360c49f3cc3d4fcd705c81898699400a78f8138f701547fd8b92
z20af173a79682c19a79b13454b031dbc6086eba899277275d983e9c2c28867e4889c0cfe56f39d
z7cb6e3ae79ff755bdc9dee3d766ae26496e528c2a6d5cc2d1da44ab45b91741e34c22a06f496b2
z09c21b129b1ade60f9fbf13527dc4423470f0a1dc37b8882ce6d566a548efc445109f256a0ac67
z7c2c917668d3d11f3a01b66ce5b69f6a6650c3e763ed5944f63ffacf1b3170b6eb96444c026217
z95c165798c012a299c8b30cee6362a1a3087295cf7010d4f9fd0abcb9cbfb5def4d548f5e5eaaa
z0ca8c3cc05bc76b354bdbdd0b2575154b0d27701712b1b9e7c26bae0d5d3c587aeb3748a91c148
zb68d50761406c921ef5b1d5c0ab8ebfb48790574c147c2b93590dc093fa8f57cac77838f5a7c25
zde6a1aa02be38bb9e65b7ba6536c98306239c6d6590775ebce6f6bec24c981c2452be6daa47de8
zfd98db10ddd52108ebe241b0635ec5d5bffe8e2bceb2df55ce4f11d85bac5ae6daa999a1dbb96b
z7614e5fff4e52fc205c8cb1e80ee4dc2e30be9f9f20e0b083ea54f40afc8b6ecccdd3d3cbc90c7
z1174e3f475ebfef6f3a82d567acd948056ce7dd85adfd3a618c864ef03ecf4a7db0d067e422c3b
z8412406cdbf8c4d169b907cd8ac0b83e88d87edc8666b0314174c2645d8721d82aec45384ab802
z6c0b7c9c54a31cb009ab90ec288b1bb3addaf13eb9493c92e8d4adfa8c84dd81fad203dfeedd4e
zddcb65ad333d72b3d51dddd5ee07bce09ec50e72286d05140ff859812b809de706e3571f5d2be1
ze999ead2b4dc4675cbfae84d1a5a87c69b8bf334bed99807b6dd52c90d1df7908fd7d21e3f5968
z693aa11a5af286be28078bcbe56321cd582bbb58a03bd6e0a7e92004bfb35e552a82b0ffe2600f
zd9fc703d806066cca4f83e17b341b8aa0d02f0591342fe41a5cb9136fd5f438e0c57fcb107cfb0
z8afde6499a4de96c81b502fa29f542b8be3c09c1af818dc24361cec0c5d3d3a1b0cb23bd12af37
z1b08d5f61839ba617bf6039a04ea9c52ffa5f9c774fef43fc63abd525f07dfdf3c156a12aba0b4
z8e4b5ed24ce0132d6bfc980599b24240957adcaea533be9e2c9f58721bb1b6aa81ac85393e90f1
z936d40f860689b15f0b549bf73e7bf29589529af150c20b680c3b11c216de6deaf378199d9bb33
z4434de058bde53da5d9bc8f9fa0c9435d655af5db038e707740bf4d28cd3b079a2075081990674
z985af7033d0a02eefad2cda77798d331727b6565fd6ceaabd0d8630b11f0cb1af442715de1d6bf
ze0f9baee7f1937352f4d1a5cc1731d3acfdab4c84426daf51757ce4a08395771bac5aa30f36274
z59138701236bf473c37631895957080f87b19237da34c44077647e895df15955ab294da3e6b388
z2652421576f8e93a7b0d2559542d78bcb3cb23d8639740d65e22a9a3e0ef59d6fb61f07ecd53b3
zb5bd24275b02364ae48f62417dcf2becc3322a9d92ee8d8786d69f1e446c31468f3b5332774bed
z6dbbed06cb9ec82a59f305b225349b22e7300affab8d8c7680cfe795f83dcf9b2b71a9b2889dd1
z7bcaf674440bd93740ec4e972637881fa50584e106ca22d6fc40e92bce05e17aac4cd035b0c063
zad797cf259b264b5a9017fe08b5c85aaf7a61703cb94869d4a59c33d5ffb3fb0a9f92334eeafda
z8d191b017886191072843c9b7d5d8af35f771f8229a2b5845295c91174c5c641aebd47032bbbc1
z3023f28d4517011d4d1defb29cbd08db80df601e8cdc2e062f1bc6628de44bd767e36dab226fa2
zc2bb38bd91557a3672e65c9abcd9567309b5e642c5f49284cddac71b8f7ba905aa143b9126a3eb
z15f1ac7c8fb83f955057c2a795a05828a50c9961368d6441a6fa865cd47228807a996f7782a1bf
z1b09d1f1e72b14e9bf10c8d27ab28caf85c9b7eabefa41738f07a0460f23c82ad385afae148f94
z40e3e016234e4256231ea2fefbac1b23ee9386006638c659bc333eba8c9dbe60157a48b1940846
z737f2ff07cf880a9c8cf027725be1701fce7beb73bdec5bfb85915ab4154ef5ad0820aeec50986
ze6d9097c1826dc7f5bf1fe80f6a9d6c1f05cc9de70b4611261107b557d4255daa8f54af95f189a
z6004cab0f2e41c60ef441041df7b2382a9dbe87f6d1e67e17e676c6feb45f704a6ecf8929f6c4d
za1fef1f75a1de39ab1b841a215b923e1b59e631b409a5472181cca7ccd4fea62fef846271cdc34
zba6f54cc051834e700eff0e2ddbaebae522c89114f09888a1db46dd43aed70cf42ef03d5c904a0
z9ac7e4ae7ec5340f13f5d880cd385fb80cf68e86a407b9729be16af3b74140078ecafa73303d00
ze218374f740b621eb1c1dff61c2c83a6671e02ac49aebe708ef084afe64ffb11b160da15123340
z24dd9c9a5f73bc4ec97dec303029b27de4dd80f69824d8f9a1aa06fde0660a340b2c9d2c81c047
z9ed61574d42dcdb9d4240dd491d4f9c87a8cf8d465631ba21be0bee9ba06ff56ff3cad1a65d546
z2aa7704f6f0babe2f948a9ae3a75cd9d8a7f3cead5dd22d94d6efe1f3e9bd6ea1ea3a7053da67f
z205d035a1a057645b822174bbbf780cb6c69ffa42451a0eda496ed97f18311afea6e5b7e838a8a
z755faac5f341049161d33e4434bd474c9993b1c7a6ea4e63e3119798da107d084357f70f5f4ee4
zecf55a73a1ab522b3073c294b570a706cefee69a24d611734c17b54922b457a1bd5beda4bff896
zfa9933ee17bea8744fe5ce5f47e8e4a76358a2bffa4fd602dd426e179f5b27bdea7ff5118fec23
z167d143d3c6be2498caca5ac618861ccf9446f5242835229ceaf4a61e14984980652fcd87fcce9
z7e1602378a7de9a2b29a334e94421f6114d48fb925c4f3f41095fccf32a5c716906d5df0548991
z96d7553629b8298cc0172092753c49df06cd5a0cdf19fef120ff0bc4516df3efe5c7c19e850fe3
za40d5f3c472f5bdf60ee0eae8cdf5f237e443fbcd8b994b12615a159b1dc3a923178479d32043d
z142f7958361ed09ce43b9c81217cb9c0cb9b476b2028daa8da8135fb15eb599c1bf20d8b17535f
z2e43e92c0a13633de81e514d411c4a379e9718c9f3b3156ff12538f6e5d821eefb90136c3e7e88
z7437b10942ad3684af2c829cf6ee010aa6c3decd1b3bb4d914cc2e0a9ab60c81b8f4c7f87f6d97
z245c4f80b50e8faf4e5fab7e9deac8edcb3b85017474c83edb1da90a978684f98629581c305485
zddc91d9eea8d34c14a9c775c0a31fe85dc6a1ec0c1c4be3919c75a7e68464878269111298b817c
zfb446930b962449a8a67915d5e65bf4e5ee0cfdc9c5772ebda45631e74ad8c33d60f7e9f7da374
z12adf3e59ebc2a524ad7abb8525e8686a184c091e8045fedcb1d1b1b62c93cd7a883602d55518a
z79092c800eee4899dc100bee2aa4ae74258663acd33d690890e27a51c272b6148d71302743fb6f
zefac4b95367b531e44848156d830a44bd0f435acbd4e030c34e413ffe7208326651b2ab2248d97
z481c5b005804a0939af1ee340521afa746d5e51893f79ac1a68618993162376ee1f49cd1ffba8c
z2f61df18bc79cd674a0c94255394e74d9255e19b44344cb207cf49c0ca59d379e3a2d6d56901b8
z48034d21b77add73d55963471178376f566ce3f6d9f35fb04b4e3c9938cbf09f966d239d6c7412
z76e7fa8d78ef3dd0717c88b038fead95c451e60c73392a27f6bf3d8be43a54d1043498c3652d4f
z422b3189488367102934250a46870880f45f4b5d3d7b671bcae0aa9cefd15c5ea954fd07ef7cf6
z39db3de51e08fb93d371ee8c44097163fd26af13d8f0c6c898d3bdbe56f04c7ac88addfcc5d64e
zbb0d83bb2ad6b700928daf805d914714351c8bf7053e72a89d792472b4e33b4ce7ec6d36a3fefd
z3396e558e8da47ce1541cd61cc07f2597c0e15a07e6a32b438f0b3da4f2be3081cb0e73e4017a6
zcf3fed94880d063c61ee33b8191d19efce7838263e617324ce2f1e10ace1283521256a1f97fe54
zfa1354f34746543b1e2a88ebf0ec837f5958c6d33b032c3dd7265d884305b0f7aff25a78e4ea62
z7d30deb2725cae95717c4b3bc76ecd73b4d919aade53701198461e1ad926f75394cc01e63fc615
z5c709abe95a006d9c62ad04a2ec3311eb486cda83f44e6094e597e3ad0ba1926f2e2bb8c128396
z94cb4410687884cde9bd302cec9c7860c56c3a70143b0dc41f4f181459a54f9b2aa22fc60a1c45
z29883afe7d95c8ba97d31770d34ef5187311ce7b20a113f1abe08ffeb5932f1c9ea87b68c6af86
z15a0894ab0780c8b0be192d398580ecf97cec6d3201ee6852df2c431f89dd95105c4bfc2d442e1
z80497425640297e61a188aee2f827956852d13342cdaec76cf6f10ef8e58ea43385bdbfbfce19d
z939b208b7236040e178fcffcf4ace07c0da13f55ad4e8b1091808f1172f6c2176d688032d26044
z188abbb8ca6801f10dec9d8050639820db9b13df0770ccb96d771a7399169d96f9120f9ca734d8
z731b2e351b833d45d151957e6d0c7ced097c667ba32f73f441072ce022b24f6ae22dd467c3c44f
zaf51ddc1a50514bf57f59057f2e861b994552a72d4aa0217f07ea26acf3bc2ee25cfc44d65fdab
zf0c23c88fa0bc559332d239809614633811622c5b372bcfeed6ced45d1ea430b61dffdd9d48a8e
zb70aceefc9eafdbd82038d349e62bc2283907d23e3219f12b46c0e1b83ad187be9f1f7df7f50a8
z2832ac8028dceef9b57c5a31dc6bce23cbeebaef63e4d0c938a700f271a673b46a79353aa740eb
z5ea509d40fc9db0ff8b328fc671837cee6c681f94b79ac0f9721f3d7004254a54643275717644c
zbb1d8e4242d6c5d3cbeee2899150c233249195ae36cf29bc4484775f744dcb9cd0b5a231340864
zd62d91195b76f5cfc1b148d8682d9150afed3f840c2c4d4a67721702b1a79d50cd9bd32be190e1
z2099abdf9ab59bc9f637bbe89c94a75b08a2b473f06a87b072f390e6e4a85e04601ac2db2ae8ce
zae5f9d171868f866889234aac18d9c5e54542c95d595b2c62391269a1c22e307754d8e5c4ef499
zc95236592f965dcf144bc3f79ea29f90ef5da92471db5d43dada8bfc8f757d6c48ba9bbe74c6fc
zaa6640747dcf35379e31231b19bd611e7ccc6957842665987e7e6c48c8894510efd9eab33e06ee
zd8c4b8e3dee3a486d45181145d8c0f8aa951a7afd7ffc18bfdbb0701305034229165cf33c1dba3
z3f96f0bb87501e2b60f66bf073ea6dd10497102bbb81b7d264b98817b47f2ca2b626db0c05c92c
z3870efc43a13597c5948e0ebe811970d9514a5116b4ce1385e5f5f1c392fd730e150836c9a988a
z0bc6d40c9d0f8e6dad22c6c95ba6adad90f7011e8ecff65b03d1ed8e50fd766944d1b5edab7615
z321711b9f86c11b7fe306e71938b88e9297e786ff886e8452b56eda164f0aa59554b2d21724245
z14033e0d29ce40b21af2b353e165da93bfcadd459d04cc2463175050c065cd715493f3f72f9519
z36985949485a04b8bd0d06c9539dbb5e99cd308772144cd0d2c376226a48714f3399e89294a2d9
zc73851907826dccb9c8433648889260647629fe471252cfeae9b2ba0354a3bc01e1a89cc19e3ac
zca66fe5345cbd646d36ed9f8497afb9e76b43814fd3ae80f9310790ff684d8c7190bc68a5f7f82
z704475fdb43feede686a0916a073d208dcb681374d042db8ef7ddd70c9772920180601f097fc4f
z4e3d58585a101cff891f5b940ba5c0dcca12893ba51d835ba6540fb0a5508ee32d5003da76014f
zf87cfb870d3aaeef8765209e0022b8f022c36a6c12eb97735cc2ab94dbfe2c36060b5c51d1c13a
z47980d4ce2b3e96cda38242ffe1bc5313ad3662a1c76b2b964fd786fed6a0785e674c3471819a5
z601467f37836fb06c8b6c4ebb2b3b533796383a06b72bb62da377d60f5416cffc7aaabdb48240d
z644156c57c2cce60a634c187835fc1aadf25a58fcd4dad95853415792777016d4bbf547b386348
zf3ae48c38d33a811612e40964e5a707615ac6fd7e6a5f9bd7a8473cdd2e22d1ed761d9ebc732b9
zb22d9d6e3c7af4b5940d557598c47379cae508a0a6f73a52fabf236c99c53a22fb091c44676e34
zeabe24b573ba0144058128ba10a94c78acf1e85afd6722592256d8bb1be0744d68d93184fefb8c
zdd901c824eff0849a6b74d6475b2a0722ed9bce7cdd5196d2cbcf00fa49f271619e9f2b209080f
z75ec31fabf2b1096f7fef379e4574775a553a3e6c5b47364742940a3ac2bec8e09ec7e681817ac
zcbf87d0ef0fcacd11acb37774b83586405ec878a9164777b88a5a5547244bb2cc7d5496714d646
zc02a3e23cc1af0165acc482b99ad20ae75e917fbe07cbe78d9f6e8264ead1c9ec1122b951a91fd
zc90a1439e91ce372e1179bac79011514cf81a3173566c5e3badf513c3f581fb5cee15b32cf9f22
zd5190f2aa6b3e2d9dbf46ca34272130263ea938aa89d04e422b33b001e858e9cf62931ab3c5414
z536c62e8f5caf320b248aeb757ffc71d9ce0e5e2be62bec3719e5197000a89bcbe2c753a74ba7c
z54a5022231a60c2d0c29bc23c7aa4343deed99c500b98032daf89eeb00ebb3a1e667f4c6b7fd83
zb5d8674581cbb17b6b594b81aef881a4e005eeb32590cbd0fdc29cb1730a5b47e14f00c91c0a9f
z3c48b68a9b3d5b20b38cb7af11975a8f921551f4f44fb165b43683b5a00b37d24650c089b94ae9
z00aa23da381d88eb9af4b62f8c7743d93c5f6c4e0c9dab5c0cf64a355ed9301f9e721770ed3510
zd5144e6d2fd63b2c3050aa989cab690d6d543cc92cbea3340bb41d8fcd8d396a8af899e737e93a
z59dfbfff0a8ce2bb18dcbea0b12ec73a08e3aa2c9e94a358df3181f03018692eb6e5979341aba2
z570aa001469c91926942de168b94385db22726be25873afda23b6064abcb8e9fc9aaf2ad1f554e
zc2476920eab971c2dd4f9b180bbf0b265ed6320f041efd106c6fdcda9410a165ae6456654ee7ba
za627b71233f28f796e4f8dccccae0aa8ffbe0f5aa41cc74d07a777542d2805b5dd0de92dfe064a
z29dd65b133ee81ccae8052a4218a7a41f4e55337dd99f169b0ee4a0b624e00628886d94f578648
zbb0785594971b0df8266ec40294d18c4a93417b2be98c5333c9489562480e72c1c9f1e6defea45
zb4621071556052ebfd51182c584350815629a8e70c59bdb9f3f23cfa8ac2c41fc5a5882de71a1d
zacae5e4edffd4edf1e985adc553529f9c0e2e82cfc6b5c036b5fa3789b2d33b92533c5d430c86f
za66f8fc2bcb72723b52cb5edddf4906708a424a48305740b093f7d04c43b1f4f89826c8946cc75
zc1662c044a6268465981402bf0cd7b03664ddc6d1ef42bb389155b93c1f4577fa8a025d115251f
z942ed153aceb7eecb2963e270b8902806decf973e1af29d96d9d98ec3f8be7277abbd15ee8aabf
zb5e9e3dc608db829dde5a3d13771f6dbb386b0d81008235b0804786a312904c3921f9d592cdbf7
z946b0410a57397b9b0d1fc0b8c956fa27dbda39b0dc56040b351815feaf0c8eb8de6ef5a057f5e
z39826b11804c4463c5f7431bd39c68eb93c2ef4edefe1acde527e698e783aed7e7d926b8a13010
zc411009bbbcd3602c8c14ec1e6b0657e89cc39abe7e909f3862f33ee191db03f943199a26e991b
zaf8f9845864161eaf340bd4e72dc2e04d8619bb03432ef8d47450a6aa82f9034760fbac21c277e
zbd96dc6775e137f6762f5ca3a81f0f39f4a6d7879a556e50d5604578a026d9fc08643d7bf6df2f
z41b2e541bab4330f9d8a3f2ab0178e33cd474acbd51641b56be8182690c810e25d9ab52c5d92f7
zd94d40c8e02966ac0f1d0bd29ef6eea64303a740bae266bcf5b88532a179866ce6d4477cd89371
zd0d7d0d07b53ecf997fa0538eb3a8c4cf182ee1a9803b9ee1682c9a9118617bdcd56097e0853d2
z5821af65d01308f250fd0d15a8196e263c070eb94a91bac76cb632bf8c0dbde7e5cb4766450b6e
z8519c3e9ae2caab72376f97221e2b1cee7cfd0e2e9370fcd163de03b129dde2ca2ba9a5fe058bb
z20622dbda415c135b8e896e58bbf1aefd8a2ed262fee156bf28671744a313b287914055d4a0f03
z7b8ef7c1c7d13b5d7ab2c7857367444d8ef85b25e358171930d9c8f29ed847ecead6d6d03b7073
z879bb325eec71a974477d93a1f35402b401357817cd90231db59e054be8cee379dbbd3741b3a5b
ze0637ec366632acf694a6f887f63c9b867bb95f23a975ee380b28ae324a6bc6424f75110fefab9
zc79c2e91bbbeed4ad5fa1a3ec861be9818c4a1b03d78a29fe1412ee6159a5194dcfb5fb47f1fde
z839819f41b8847ee1519fc8fa63142073440fca3aed13b42e115ff753dbd649e6b0acba74c4fdc
zeadfee305e03474b2af8d5707f1a42d61f6cca1e9d3ba4242a9c13c54202cd504f648df55f6e59
zc5f33e285a2c38c3726d44ed7743f4d98f191fdbc7be9b9d14333b252be7694fcbb1a5b0c1c9e0
z7259e3cc24e1e749dd2a9e4fc2d759031f5ae8a4f6712f8e4588f41cd8b14d391cea97bb2dbfc9
z76195852f9b79f65188bf5366ec090360f4774a923e5ea2b549d41fb67c29d541848421ac10196
ze80c3b3de919ab7c836be81c90a648230d7840da034159d5208ffa7d0bd8239973fb2bad15210d
z72b4733329d70e2f1531869fd94558ae526ab5f091b34bfd51052b56a19e673254fb32d887835c
z178ca809f49d4e2b2acf54f07ff5d8825cb2572825b8f600e2cb224ffd57ba5365d3b498901355
z729aacd1a0732159c7f63bcc983b2007a05b274a88cbd234d2cfc5455e44b560228a349fe827d1
zf51fc537e13b9a96fd4c9a2b4fa61d04c114a860163d721eada4a0dbffce0a62d62ea0e00a81a4
zfb060025e3136f3f29fc77a59feadfb8afbf314b60aa36ad00de598a0ac1325e57ea8cd547f6fc
z50224ac5400d4a1b09ff642ead7958eec81c8256ba11740bcbe3059c4f40dbcbdd663ef7322730
z0d27741c6085a5e37f57e117b7f6f13cbf848f15635a079d77da8faebee49922934c21abe691e4
z0182c47bf9a2dce22796ecbd8bff485778059d6f4c7ce6993702e1c4ae0a54b7d76bb4b3ba7172
z0239ecee3207310066f3f52c8d4541be8bf3cb75844bf4b11ef7ba9969d945c8608a8c23d984a7
z8720593f065fd9d68bcee72b64fa688c8ddb462bf5479064ad464d04391d86e4418d1808d6f177
z24359686aea77f582f6e39c267681403ccc6694fac865b17d1a2f7f13a4d1b34dc823e3a93d46c
z7c2bc3bc0a1a04d41d80e50b91f1ee0be003f657a004cb0af148fd40fcde042ad7ebaf373d9a6e
zae0ed123a05c7a27272d2cb0c024dec51b7a8a27bc9fb3e86d744caed952ab47ce3dcf424f656c
z0920b744e7aad85cba062acfca411357ac20ea1c7f503c2250c261629ce07780dc39e29b101a2e
zec03935d744ccd7e3b2a9faa6b69a40f8fcdfbe8bba32ef61d82f3fda99ad3bd48ba66e600d4df
z0174f8465e054dc85e3739844ecf6c240f9e1c2b9e89dd7dc7cd91890be86fb508c5a5d9dd0a26
z4d5bdbedfed0892f0a6e88f5ba04a69194f8539e4f66b92de508d1655a0e3977186e77dd02dc93
zd55fd60517fecf5cfdf2428716ccfe5f32ef7aff35e945a91cc2d3f7dad485e64dd794b794ec7f
zdbb82cb2eac5f7fccbee6b5d22a490707d33af13be7c54d11fe138b903105975acccb951e9b929
z9c5afb13241d1d90c52a19debcee5df5d1c19fa97d1f23f333b760742048024d36dc03cff52148
zf0029fed536329c252c723ee630b7da9a02a3b6f64fe82cf47d6fed0d8d510ff1c63a9d0c35a26
z2425d361f2bec8d46aec839d6526a011e2ba941f91563034a9c59a05639468a0a8920dd471cc16
zdf1e2a2b0de019fc992db4df0ba5d09e2dd6d531331e155bf717e4d9a642a4328589673da212a2
z53766ad8ba2e95eafe469b65fe42f70f2c09b9f1efff95b1f22adc49fe9c84ae9b7b9e3a7bbc62
z09dcfc78939800d4a554012671e75769ee7d30a0767a45334e2c3d23d02d2b1108301a2cea30be
z4852224ae20b76aa321cce36c46011185ef3aaeb8bea35b429da4ef252777a23f63ccb6e537ac3
z33a29c63de28735f66fd7244585dfacf99b4b20296a12501b2834951c7407cb4df3209b0a0832d
za3a4df27ceb7d406a80d38dae2fec929706c23ae8d42b1ea9abbf5a8500570f36ce280d0db308d
zac3a1ce65bc52ef462863166a835e1c771c326e68f6871b50865b366e831ee64d91a346e8cb257
zcc45c5cb23f58319ae3b94f99747ea94c77e552c49ba179ba40b4313f538694c0517468b9fb1b2
z0a4d47637c56af0564d242e432a9faeff6632f2fd38ba6f5249ed47da36750fcb9d3b98144a097
z5d73c2ddb5f92649d3e9c434122a6d1ac3732a1f62c09d2c4f6109a5d680f7634dce348a73d934
ze7fd260830456ae3b36719f7562a53f49d16ee4de02223e6144b7a777de79a4cea8fd3245515ab
z9fc052ed2971d990d5878d0f38e59652f1b7a0c8af301044d50ebc43f6f57142fd2c587a029c2f
zb2a247f42ffc9000042b8e59cd16e4d7db5141a1f851d4b5e3a9ee5a96973a06e08f718b392910
z28f4482d4f8636193b3bf05eb6086c966b05cb8d8f72682df7b0e3d7629233091788401815ead7
z4af1dd26eb6694d6c7d4f482885349c53ce06b26d4fddf66111b0e080b594c30de786f35ff048e
zdc17d37e112e93ac4d0fb0077192c5855eb036187f0452e2767968cca244a77b6f0fd27babc9a3
zc20c8aea37a7c957469a0ec756e8028bbb7b3541e52b5d682196e9b5a8bd69a14f726a8ab9d349
z02058ce853e7d5f560584d504eb7a12bc53065887b14cbe0b34642b1192f98e6333f87257736f7
z885b739ba96753cedf713b50473e220476196a15cd1b2101e4f36609288de53a953f106e975844
z6de5a0372f076ecf66be52aa9b7bc80fe666409b7c7c8b1b724c1411b573e8752fb4572452969f
zae6fa3a2e457338ea48ffff589a1b3a70912b276819559170874e9682bd2227c76cfac781fe047
ze3e452148899e309f7a9b63f8fca7f6f9ba5f390eff72fc2b9e430f167de350d03d94c9ccf9e74
z03428fdf23aa985e7fb58e5c3757f6509799af0bfaf463cfc5f006452f0c193e9a0aa4cd263a1b
z68745cff13e7bc004d082381dbb1188587ced05d930cbe0aac02a33b4492fff802f6550c179490
z5f4e24a6aa2422bdcdc607080d598168dadff09b61fb7501a581ec6ce46f66a149dbd619b8e095
z2883d28740bd408abb8c9a7dfe3974813862226380f4de1d0910a9299e24bffff85122e316eb0d
zc704bbc5801f6eabe20ef50edbe1c98ddbb39b688af5544039592d724f241f4aefa04a341a6177
z912d328c768551bcc74dd78a797f4a540ce3040934c241afcecf15f8c9da9fffeda63328bb7ac5
z283a648f16dac501c38fcb3deaeacdf18ba7a9ed5a22b441fab39d7a2987355bcbe45f984ca68a
z54c1275398d40e51f32f07bf0c026110036a6c42156494d65cee2aba68d15d56c02267c7511b97
za7046790bc74cb7d33f3d32350966ee368e852096dbbc85bbdca9dfd42d0425890f073faed0e25
z043bc36b2c15617f21f0f0af653d2b90aa93cccd52aac47e8b1e94170dc76fb8e03a4d655f6d5d
zab21608b0f9b7bb6e62a8beaa70d8ad5aec0025187e35f9b3861dcfda7a26643904535c827d3e3
z781123ea2336e4afa5a6703534737061bcbf3f4f7241911709f77ecfc19897a81ddd8131024ec2
z4ea824716104ab5a5c63926f679cb7f4b45f9098cf4259f9b0620364fbef4e172f26cc1bf089f5
z41b7c852fed21efc9b41452aee01b3e16c9c53bb5b8bab0f292050f5902251f63ceccfc3017305
zf383fc2e50a147bca58756cdf67650b5e8ea2cde38b9a85c06af795e66b33fc841770bfcbfb7ba
z2187f2bf7fba2280682d8029b0a10c61ab7510e9bbf39abce93ef32de2472eba4ac4c3fdc26bd6
z9011bf390de3d33073c04c3c731a2fe6a5f987cabb4ab17e67bd89ae908192b4d9de6537e3f19d
zb807f3698040c125a7cbd94a040517c2e3acfad500d36ab9df0ae768e3d1aa7b5d5671d6ad4bf6
zd3b7a695c181b7466d55ea14c716275a73236bb080adc6e669d10a15515812e98dd9f85d06d47a
zc8b743ab5e707333a3e1e0aeda29d5dafa236ad9e45e67052930f5214651767b457d5e2bc8bfbc
z715974b6d7a0c98d4dd6d35d11320860ef3e62072783585f701e611ae40fdb07cddbca5e02d127
z900542a941fe7e341fcc0a0bc68e0da1607771ab95e82bfb240f62a5ac57c5e0a5ea364fa5207c
zb4f01a1e134828c3221c40205e1bf4674c0a998aa06bf20f44b98c795c67a78faeb307bd798438
z6dec94ab0d4da5f9744991bcc232379966c6a691ab24968b4e7285fa5889b5c80d6c5d49f8093b
za3349434eeaca2c163406707648a9ab9738b620c527f2d4b12f6aa2c51cadd6db070f0acf4d368
z7641e9e60fcd9201d801abe0920fbd9e620b8c110bd1356c3b4aaade3427f7ed276db7e4cda49a
z51e41c3ae18a57c44e0642abaf366bd3f5470195ae69a725a5fbd0b59f79d21cafde31491db2b4
z83fa4d11f53b6e660d45c3d47e2f5102bdcd69b880e2b76f684f8c2e10d8be1775a6246ad3a599
z49fa5341d8de66ad66887dd783b7785c1d68ca0a39bb9c7dd47b3905e5274fdad1f296bd109f9d
z963971992b6b730bcbba9b0195c75d0cb0433ca85c10123401792fb0c8de0b761ac4c7c248a2e5
zb45734ea45304928b9144076690e59ebf944da7e3cae4083859630071140ec6dcc9ae56d054e6d
ze772c2a1e650f7e79be661c913114f9d557414018c92b6fc504ffe16a69857a7d2bd2b16c57bd8
z0dd96ccb9fa294347fb094d57ae8fc94427ffddcce5bf6670bdbc07e5378d8b5f0af7243147f4a
z1d4f9bd7c3fe3435c834509792ef83d78e4ec88e69002d66e968618f014f080ffcafee6801b211
zeaad90700168ba944f77638d60715970a8000b8cc3f79e9daa6cc0e3804205018165ede01db050
zedd460238b31c9e91b94da1b476a4e27ceb26815cd15444a4c3a8f559a6912e474d259f261fc30
zfc668ac60aa04207176339cb6eb3cc56a08b6ef87fe781abc166b2c303f31d43041f79641a25b9
z6e8515fbe75a8ed6c1d66605445e5022fcd20abac6ed3ebd5796fb8b623789e719d420332503c5
z99da50ad642d13021c54799a16f6574d0ad8e54e0831c7523027b763bee211ebbc3ce04d905fce
ze1a6aa467e48af8ac9510e58e48bcf1b14ce132f10df7a4cfa1c436684415612df72aaec281119
zf53d36a91e4578a9cc5b0867f2d0f13b696813d58e43a6e5d39f21d8e02c121d5ec75d7163f985
zde367dca9baf14caea28a8417f9886b0a9a5551b6073e562e08316ec6dcf9ac5deb35059108a27
zaa7541284ab9002fb2fc99b03f5a84ef56691c1ee5789f7344f573bfe61d57b3dc160712edcd26
z6aaa79a4a6bbe86dd867c4648819eaeafed5a5f2df295754f5e89eeed5e54409f16cffa00f2c72
z76e2de64a49945906fc8a21963aaebd91fd0e185bf3783883c8a58d6afbb883c0fab8f3df15b1a
zb41155ed77066e5196ca02e9c3ca69135a3a76aec743acaa3a84d3c8226f2351e41f1614c58669
z3ccb1aa3eb9681920ee6a78e3f846dea0f0733bc08e7b3e0b662065b3a36ff44eec5c8344d06e7
za384bbe1daafa7979ec53c662df8de793433c304795be9a0c86a5da1b3ac5d2bdb020f9c1fbb1c
z000171dd15efced8536cce9652be6560dd0794e389623baae7f24adffe0afc42923d450b0c5d2d
zf3cf3157f051f0278561306fe3d0c71529cbef5cc9469afe5e63dfbaf0a30082b6448cd5301118
zf4a10ccba4f1d91d2a0367b99d291bcb81e89773e09aa59b6210db75992467ac06305bd7b231b6
z4f9df295e4419874628f62f98900ebdb3b3be5109ea6a9bba996e1df8efc29945e73ac81b495d7
zb45f0b9c07da50ac075039530fdc64c89e10ae866aac4eaddfc6d12e0755fc5d960250b1863e7d
zc5b3517c89bccac42f5d3c391d49271e29dd2cdf1770e7782954407c6ca5391a4d1995f8062e48
z243ebc8ab5784daab5bf2894f3b7d56f8328e7d289a9603382716ac1e3149e2a81a4bf9a11a314
z456b2bd1aff9fe5f245c2f7adcc00f245a80870eadd48a10e68971b7f568b0b0325d967ecdb7a9
z3a17fad7a713bc9a248dff95166fd9446552e08ee11e5d25ce21fc54165f99414c6ef309ffddd2
za9042b90a212f574d4a15f7bb339bbb94fbf037921420faef96fed1a7fc9f30fd259e6ed0c16b7
z33e2741b2eb2406aea7efbec58a5b1c2722286b3a2862c050d4dd229efdedba32aba3d322a27fd
z3510827e57b6188b3aa5e949cc3c9e70ce83fe35181409ce804ba792361f880d60696ca2f4b447
z43a6f8a29019dfe864c8f5713c0f98fda6f957a7b0f3390faf0fc1b01e12b5d67f4fde56bd86b0
zba605e55c207cbe7ed1e716547f3894b9e243b377abe0808836f50ed378c38b798974a1a30b8e9
z6bc23911f2dfe2a86c1fa72a8356d7ab3849a7e64b0a1b1527d65027be182d8527df7b6e80f3a5
zb4544ff7469752671ca8dacbc907c3dba90806b29a1442db9742ded6fd1d58753635c3ccb85901
za9b37de451ad8003c7de25fab5a56370c5aff43cdabf9096154da9856d033d0ab7f043b61bad36
z4b5367341f39d32e7f4f675e5a4cdb474524792be4b6f8a5a3998e22e0bacf890e933733bbbc2b
zbe740d1529fbfc3adad0b83a767d1646872c9fe2fe85ed54da697a60b1d57931e52b5cb4a5f942
z876aa69e14280e66ead01a85264d138207dc9c3e712a1a396c77ef2637ff6270cfdd1ea307f121
z3aef677585a54796c94a82b06c24d1bac78f164888de5f11b481d3c85b8b9cde93222f7b810aa0
z667ea9da7ce2123d31bc629eb8f64bac70400e70453b7cacf80716eba12510efed7fa86d47e5fd
z60a5af51094c388be21ba9a2c83722f5c3ae60083001bf655e25d344eb4b1f89de21fbe7c0a8f0
z2c04ec464f6f7af58654e8b46d992c81f78e4d35314741d76c9d8f15942de7df806160e155a39a
zfd9f976b106e4a28acbdd72805ac182d5a4209e8fef7e41374874c9ebd5f46eb2aab10f0a6b2df
z836b7a8261711282b23852ec03ce4f86ae167369d629aeee1d8fba0bb2a994131e93c1f3b2ea45
z3cb7af7f71f29d3c735a81ad3adc88168c631bf31d06c90b5a52ae3f3959b3777f138244b82a40
zc18b4d6e2bf25a610f8427f5212bf290a0ade5d1e236d9959ca63137909871d7df8a49cc85612b
z807b96e71af07675f598f7f8b76cf190dc9f98ccd9e2143c8d7b73edb7fb0c1cf034c6c59203e1
z04f1c365f0f9fd7acdd63569d12b0721e4ca287841e4076992b85732936ed5a8715306c34fd1cc
zf2cecf4273115e8ea0707e22b742b9c3745031ca4e74f643716bce7de071eea39bb48db8c91004
z496af02858e1759822e1f4f78459e80cf68f650c188b97481aaf11bceaac95ce2ddaced7405212
z902592c423926318c725535ab2174bd2c24ec8000001582e44ff1e7859a67716f4d3d06d9be4f4
zdcd6334285247ec3f0968623f584c9fdeca965f8fcfc5c566c1ef13338f2d2e5fb7e590f1231b6
z41e3a20d9bb1296bb108ca356b78602563a0c69820cb1b5a52e85452586921eb8fb52eed365910
z22580eda219c7c3fd253ea470cdbb2c131312b9b5d5077b8d3b81bacd056ede1dc90df330a2c79
zc99155e8392b09575d1f09f8c0dbe6a845a7bd6764f3d60c035e49c5885c356e628fcef3e0b834
z708e2459f0914853d11c02cda87d7f78eef9cbc9da76ad7724cba40cabcb9619d601112b9cf944
zca76046fbaa4bcc7dc9216df0cef4746c591bbb233d4390d3a2eceb369da0de0a885989cf927e0
z1dd907b2109a41e1aadee57fa40f2365c9f37ef04d73a830ad1979b9d0c3d26fd7c31901625417
zb0eb1d3a5beb974923a128865548dda02e93cef7be2fe184e02aa1e5a3a1a4dafec46950ac6457
z823e6fda2faaff15396bcfeaa4cead213ba011fc1cde16a8b3c41a96e7b77eb0e1fc1a37173150
z912be85cda2150658f493cf9cb00dcf6731a8294d2b91dfefccbcb95abdeba9f8906b52f8769d4
z3b0b2eace108a0f44af696633722f2df943d085b939e6fce1b2396f94f0b12fd28becd31a3f30b
z5403ced41b572487dfddb3007ddb30c7f41e64a5467de98a9f51698bc5d4e91cf65875b69e7797
z5af2a4f45deaab1722a03b57347b84bf6807d62d49cd6ac3b9648e0c8334a027888fd3f97f459c
ze8478b42de08536e3dbc8c372e8bba246454d92a0c5dad0dd96c5780f111015ff85dca8fbee483
z1153d3322d772a85f2dc65a12abb9054c9a782632f6f6af59f83256420086e205b874c432ad8fe
za709917d839b3cb4522c34d4b589a66ce15758418fe348f1ebbe13da51103a36f3a39059f8b0df
z1a5e1dda3aebe31aaa2e6fdf0a0888f51cb3670318cb000136148631f31f14cc9b590612bf90c1
z2998a02e2646cc839ff82db293539024bafb62b0e37a016fda0631427779761cd9f02b76b4d1a9
zf8a05c8054a41c37e4242f87d5f35d03247d7baede06b9535e4b0b104275de0c808b43159976b3
zd7940ecd3aa9ca6705948327b4a6c1faec69f6205a158efb61d65627c19ba524da9769a7a77aa2
z4eb922945947492b687f596a85baf9cc63d03a49a0af44d94f214d182f62139e95ba47cfb69944
z10eb13fba24f293fb34139e6b0df7b557399b51e36cac0c507d25470997f435219363ed4a298e4
z14e6d69e13bfbf75016cc79853c4faa435428c626aa9bdb69dbb5d1c13a4bc518235ff056f37fe
z17d681809980ff11db83a6536f69004cf04680453601e1838509c18520d7022bb0f71919f1ad51
z1f0750385c0cddde8e7a6227da86d43eaa2bf57a556aafd58c94d0ef45977fa7519f9c991ccbc9
z441995829bb3d7535569297db411eda52bd3a09e2b9492939490ed7f5e49521af08ff167236a4e
zb18bec50a4edb888c2e8182cdac2243fbdea36025f8ef36e0f21f7f1265304f7f5f0e6eeaf887d
zc443990ba3d82f88db4841212067c6e1083feee15046782fa6a6f1e6268af2e5133ba808e05ec3
z037ae76bf30f259cdb71f0f484ab3c6825cb4b9f832e9f59eda71be9e8f8c265b3022cb41a51d8
z3829c47d9115dac7120bdab819e562bfb09348e0b992f5a94514e865fc68aa25f1a61403433d60
z6a77ae737b9f86bdc1cd7b48ab59ab239fbae68201d8d9f5733b3dc2dce6fe13904e30a288490b
ze1388694e88fb217dd004ba9da4abac572edbba06850a1ad261731a2c859b716f71dd0c6775b15
z51a9dd86b3717e8b5dd2f6ea305c3a5822fb158832b93e50a8316cc0964f8ca96f307d740c327a
zf9415f639c39bc64a592b86d36a011d5132aa14154f36890cebfc50536452bb00ddbdf00d94c67
zaa18f4185de8a548703bb004c36aafbfb90600c9f8f1c5eef4ff2da35888a1b9ce11806d75de88
zcbdd4515c1e40f835ce07efe88aa685044e0a38f50dd2d1ef6a516e9f624075a6267f1f55b1d01
z9ab469ec871b4e9d5690de2dd74a7446809e13396ed720b9bab7771a82778652ef93e6efc0f3e6
za471b15c5ee33212ab7a7d55c2c061659993c61f41d2e6d8b235509e13d33e82272f54690d7055
zc2c0a99621669cd81a85957418eaaac7ba030516f4672988a3394b62bb8183408e74dc3c4caf3a
z6dd9fbb31dca2d80d56a49c99c369bff5a9a498f57553c03763e7100e695fc43b4ed2282bde570
z2766f8cd4fffbae7e331f1e10d2288582790e770d80e86f0b7e5aed1b98115baaa0660893b22e5
ze84ad09a5fe920831cace7893d351c9ea05800598483d26b1054da9c2e0e4ca5cbc87bf9d6473c
zda9d6c4e3fd2925c79b90f5b926227a5845eb81815bf836a5b223af4df0782471db4074202f823
z17174ef37bee3ff87648aaf55ca13a6a2f754d41dbd705243c14a28ba53de87a8100b917488f44
z1ecadebcad5756966064ac1fda2a2d599161e1f2dfce105625fc0899679c419436a908179c7eaf
z9a94892795ee575150e99f72ba04fcbd290aa51105b77fc190023f89079b47eac37ab315a53124
z3641f9be37d0892edbfc27189906e7252c4dce3b4b3d02f08f83d21901261322fe1e6f2ad5309b
z442c3721a05398f9a131ab9dc5fa9f50f928999797a19732514352eade1264054ad47a852f6278
ze041bdf4d4971cd8ec60d51f1e8be023fe1293ad0fe2b07b6fbd4e949018c65b59ae185cf705b8
za1ef7e38cb755a3e8b9581b7e34037d90de0355b4d3c662e559b2525a738bbc9aa5502d7ec2024
z28e95965cfa878595e7238714c58906dc5b433ad4c2b5703708aebd57d8176d450d79beceb3525
z1020d1193b70420fd9ab232b3bf9249220eb066bcb270e0819f1e1188ec978da4359c56df84e3a
z68c0a8e6d583e0cdc060a70365fa9aa8d63d70e785ec84affd4fc9b2c065385017da141a8b77b2
z2f1887962a71f7265e874b7bb5a71996207df836f72515a85f5be6cf62cf0ae1838173dad66285
z6f47d809910ec0c89381839b122bbe58cb7b1b9428bb01e2069a0f77812078ebdb54aa3cfde7e7
zd55f63eba16686aaa4160c483ff14fbde7626020ac4592d14a129947d3888f51874f6604a9aa36
z79d10afff597e539cc269afb416bf1271a58677142208f2e9827d555c343d115ab051fe0fd14c5
z26647c9712b9e5ce7d76d35fd49b56df744ec8db5f395a3ae748ea87f914b092e6d18bbe773ec6
zd5c7fddaa31e7a31a979076a93c5ae539d3b1ce6907ac6ba040df1400f4a40abb10730b24dbb38
zbc3a04de88cbe2c6568e33f44bf47585781cea4d2ba23d7bbc97bce0e1bb27e18e32673233a206
z95661e84d4d2892c9de1c3d816488f1924ae76c036a2107481b3b6c4e85cbc7c42b0d766565eb1
zbc93df90d5a2d25b98baac495ed197081a442d7c35f15e542465fc9442339dadf3bd25dee6bb98
z3373ddde768ec4679124a594f7f2a421934159a91c86d4bb260f4b7a855ef6ddc1d52c13d1ccff
z0c8f66e1feef9096d54f0c3acfcd5396138e747993b10159595c8634b354719b7be3efc0b62077
zf1fd6ff2b6de342b43bcb70a31b96629dc426176fd2478e55de8faecb90fb42e33aa42fb0dae9f
zaf71c0f9998bd538e5a54f87d4b7cbff7d61e7d594deba5932eddfaab9d11f54dbd0f7cb6f09b0
z63ef18f54276f4ea752dad0f0453c8fa5f908f558a11da83de71168a36f83424a00ed370f1a177
z1c32f7f1bda08fc21817a945b5e3143df34acf21c752a01221085b31375943917cec9e271bedc7
zb42a630deb6902cc355073660ec72ee6efeb3cd19b285816ecd6c762152a20f2ceefb7697a14b6
ze500848a9a9f9abf7ae32c57670337d86b857317c48f332ef7715e39d312e513b8137efcd1f837
z7ef15f6ff4f5b16f8a36ef2eeb1b530c266fe367a04205dca29dda5c9c6609ab9d3b097c190526
z5451dc3770ded7ffa2128dec22c225f291263c727e3ae055644768432ab97c833c164d8eebb197
z70825bd05b63ff80801a546fa8ef9dd9d4cba1d21ab943cc2f9b371bcc38a7d3513eae2a145ad4
zaba94f5be937bde74c3b93345292b740790f56378eea550f6c75d664316c2d1429c3973ec2fd5b
z2bdee6c918678e2d2472eee8fc580e74011c6393e58e845cff16330843d7c0c0999744ff507604
z69047d173df24a383976312fe10982559f524caee799cdd83aff00052472b8ac71f669ca94dc01
z6f079d301afd97060931d44bf5ca720d850d8148849981234561fcd42b27b0df30bc57338da9e6
zcf733f656b78f8e3c0da90e9d7467d0db69ff4a834fa6f8bafe77ef83d08c3021ad7e3b3bdb527
zed20a5a5af970a60e775466e0858c8ae797c0d016b8de136120f0a1138b048ba3496797f9999f0
z54b08c649534a70085e012a1e3f137ad1fe55d1b48855a54aade62ba09fae0c324ac315eed37db
z96775b32ed4914e04495a87901ced45964bafce9c4c5bec01d5faf78be427f07e8c16466937781
z4b733fa0cdae3cb9e2c8de0f6c0312ddc77f0e9231f18f603e44751c7e62047913e9943e96ba70
zbcf22bd6985af867eb299d0465077020108ab2ffdb8c111727cc40ac212e2ec7bb045c197eb780
z4b73dbcc4f8ce4f95a0c8c18d9ebdac88fb132a6b1d6126f3eee981bfcf35d0caf7568cc043943
ze8a42c8aa97fc4d46278f0541d09df19b106e928b3a3f86daa1e5b941903dfc807d35e4c934819
zfe511ffc9a809b256e3054395f66e6ab00c69c417f26ecfc66b84e08b62df6c611ca2e0acea441
z07db88c7733603d2a7b5dbd2517d08c864af7346b6b06a3721229853f316d2f0a4f16451d4fdea
z08b63d2f1b0fe060bc9151faf803e712d69e49a3bcbd456f5c3b0d564c6422bab6f6269674a0ad
z69c5da7dcba4f4f784141412175caa202aab523e805d4d2d394199b341cadaf196cfdf7a490fcb
zfc453f0ce2b071c7a5621b9d680732b2c525dd97d540f1955b598b92880ce42e015445909e176d
z8b87cba0e748318ca91f88e4469385f549fb7ef7b7cd0706c085e98f0c9e2f07d9d86a5c95203e
zc6b6c810b242e75c5f83e3e040f5c24e31b6e84192b2b87c5fa6f8281ac38c9b69ab41db3a4844
z8124f84663ef234820552f2f2a631351e6ea32c9a333dac5c4c607651867c35432e23b7283a5d7
zefb9ed8fb3b411daf05ad72d3349282dd40f84f36a65abfdd3dba4fa8c00b51a3c83680ab481e4
zcbca4308b135598a62304d3adf603405aa703a5391aad7926f9324e158ccac945479c61e5d64e5
z619d00036aced2e54b8821007bc9cdcabc98bc0b5a101fd2689abfb7987996cdc5e1906a550b0e
z093562db955773699c4aee0c1468ff7fafa0fcd576626e3e0fd39d9d923abee89caf1832a59795
zcafb336ad2b37cbb7b2434b4c7a031140a9139de748bc3ef6ff0646f96c4d8c6f2cf84746d9cda
zaffa15525dc0139797a6381fee3f615ec4f8e227f05dc6eeed4da78a797a72cbb916ffb216e541
z23bfe626a345b03e55f321a443c2acfb0b26465c1cbfe3b29b001812f1b559eaeff7189dbd5afe
z57760b107a57bd35a35c6135f8cb95d2de10134e2c0e544f03c60ec8c4f717ea84f694e1ba267b
ze6867041382f54f111dd523211890f2a0b63510af4497ab4d53be8030f47d25a4b005d50774fee
zc65f7e972e22b54b12de6d5d297c265ea3f31c258f6074ef4f72af813d61bc33d66da6eb82d86d
z61cf4f89d962fca1a72dd77b5dcdd04f88f8a20f2117c5647d5b9989e197ac2d32eb3248123764
z4528da8d30dc3070f96606ab15d7da80e44ea43be0f6976be7892d1ef0fdd160947d23041361be
z76b68322f53b76ee20f330a5efb784a084835b73d981f770e7e426042d3eb5b9e346d9e6ef048e
z745ff4f0e62e33d7f17381130423cece55f75f156638f2ba0f2c79c51405c46ac085743d040283
z1a2b4af38fcb9423d956a4938c4a67c630bb6d4c0f59ea15fd5e2fb02b7526dec44cfbabec6dbc
z49b2e000b56931db1061deaac1546c1151ee31dfe9962c665f85e25d5e1dc6ead0042ce867913e
zf664cb037207c68b85d426ada3e36d01cc73c37f2cf482bb5c2b34ae0f93a2c3c742c141f5b152
z16fc1215d291ae5d2777540fdaf04d92966f30e2e764193e76e88f5b6d3bbbb76199a38208ce6e
zf97a6a2873bbeeacc235562e4978cdec296b54b507a8ec6bba996fec7af3e3552fd93e02abbd0f
zc1eba183ce5d83b626803e9362777c3cbba2e8774cad7ff01270c4f0d2f0566b485dd44dcb5fc6
z47fbb78d62c17a17934edd860e70a4ce61cb87977e8df77c3274619211e68fbb8d542127cd9157
z01e30c7a4f305ca79edbdfcf400ff56a4ee93a646d29a3a793465932874f1b9bd5b08e426e2a69
z73c3c1a833d004850b91e2e80d935f11c5d3a0769f4bbd406111a4879ec67a8a097c83737ab0d5
z7557be73dbb003775f43705d496cae8a5bb6050535af87bb0c11930410ccbbcf6eb0df27a7dfb4
z8207dee3201d803faf5ed30056c1e3b4054704ee10e67f12c5c2ec1e830967f90ee1c2c71cf709
zab6b30f8b0571a47edf6a4eb0620e4f555a14cdd21169dd442c6be278554b260a0255da0de1e2f
z45c5db56338fc404959d4fd1b885daa6c8267366e4b42893e611891c1b207c25ecb7a7e41b229d
z10abc5b9ddf6e1d508a6dd442fd8381270fa34df6960838199dd55a3ff168f2e9c0f3889488547
zb70563cb993283463db210e56ad67ea665fb739f3bf40628da656553ea6ef8074def3a45bd19c2
z44cc3c77f47553f8a137bb4d583dca7421e460827932a11ddf14aa2c5ba734839367426b3ea265
z8dedd100978fb8d52657921b9e43b7420ae5dc160eb0725a046f5c197bbe0eb5041e08e8af607d
z57f85f11721be43e09d05f933e728bfaf5fe4521a7a6dbdf1b0ded78856b9c3ea53c3b09efd759
z79f43b0c9399adf38565313f6d61e81af25ccf901d7d066bf8bb62e895bd50610ce62cf475a859
za9dfc22f1194beb53f00264d1939c932fbd89ed933b0819fc01a6d78fc19fe21247f49ded58c11
za6afacc48ef8982c651be625aa229bded689c8c7188cacfb17a5974c9253c8829eb5ed0c65a52b
z03daebca0f94a439882b9c6518db22fef217ea9a9f4ef5744b59f751deeb019bcfa2e5851a8a39
z7ae2e6106f6522d9ab7b6190f004f0d2f333932f1a65ccfc5db7d71b12f764335ab8974787e2f6
z608aea0d463e40b44e07319e11f5be464894fbb9e5d5c0e108a0aa85f3279474a5cd11e99e228a
z532635356d4a0e0130a30b1d8cff8eae0f5b328adb3a2362d61a274f2b78e893d10f43149e3e3d
z57202d78b1266e4a7fc09ddfae64a0b07ef4f059363a5b5a725af9f3cdaaba89ac6248c0e437d8
z7f15e4dc7e894359b461dde9bd14aff389ac410c952b2e016ea6c0c7c1584c03c8d93c564201b6
z7ba03908a84b72c32200811db449778bd29b9b0b083c0663952c6911dbac45596cfb094972e2d3
zf72b522c4086346ffa86020231261508b6184821612395d99473b65f2b556d99e7fbb95fe69374
z00d6f27e0ccc3fc0b859bf3bd9eee38dd127d4a77ab0144dc1ec8a05cac7ae7b8cb8108a29b57b
z4d1ca7d61aa34428827e36b66ab3da6514ade5306867267035ad7f534c355adf61aa59308e097d
z8aec143f65e14fca276335862118643eaf56d1404fb3dcbe95bdcd116b0a84ac81370d2cb561af
zf5daa15d12f5ffe6e6d9ab22da6f84c719c3365d7ecc879a2e22170b0099df979d311717d04da2
za4f965d96388a27a569d9a65423494cf4ae27df4334bb70ebe74af393fdf32fe5cc6e3036baabc
zbe89a8f8cb49e5261baeee139f4e98cbaceead064692ac32c88a86519af9b3c31632dc7ae1393f
zbae1e8d9937a73d08295e647cb745cc39052c11319e74a0ee226839350aea2d4d6a4650c80ec13
z42e033e871532cfeec03b3b456259d37baeed51e553558311019db00017e0990707c0ce394f025
zf0fc9c46926a5cd7aa8042c9510846d42288aefb004f6ff7d6489b8a0ac286e1b462870cf463a0
zcd6c10c3caede5bb53141cb94045f5e18413881898790b2ffb7f3c6621b9c87f863a5617067e1f
zb055ea5f8dc333859b7ae4ffa5d2663564147a2c893a117b36734350fbd3c7a7adce196813c4fe
z854793546819272b1010460f65480ca9d73ce8d8e1497eaa5a390d12f4f6f3c0d3f02038e1943c
z4b5af93801d050369011bcf6f4dcb200d2467d4835cc9e4a7561b496ff9d78d51251d37661d2be
z2f18f90bed573693df148cea8fded3ea33db03ba3e9dcb3b465c9f62a94e9bd0ac61e5b70ad691
z0168bbcb8bcbf63ccf63d26a896c984e2669312b17ade2a028b5052e330477679e3257a38b3e36
z1e6e6c376ff4e849ad466c0a02237671d62fe9f4c309713a56d8bb23c07a6f1d9d67028299210c
z929ff98d7e3f1dbfbb4a71e6af1e56417a66fdde103a6ab1db49b0107c5c396f120db38ec395cf
zd8b690c9ecb82f7903546c3f282c63cd3ce70bd5b73648ec29a870392b6b5eb07129732faeb9f6
zcd18ba481c6375441a3e63eee272ab04e750dadf8b8848712816b74f54042d303f773ba94bc62c
zb5b8e97cc1895158b3b65578b83cc5d4261015227a37e37ee6f24b2874290ae740fc857f8bf054
zf8be18088014272ad1f851b95a1eed8f7591a9768a4bf8c49f96d7ad8b06303b8136430db0c7d0
z070da504caf707e34b1e9697f33ca46095906906010c94e00b2cd3875f418bd425e3971be96ed4
zab10e8c83b8c76b3d622f78eb19ee620bf9be13348a1452108b1d0081c8df8a81e7e2dc8cfa37f
z297ba66ee2af414f93947f238bf2364aba4fe470a2138b6e1c52fdf226dc210fa0a3142ce23eae
z6be25ac189346e5c556acf0c61ec7fe0820014b7c8ab5f243380f6af67bf99921351f387783bb7
z91b8209f5f1618ff2cc11a57fa48ee3eabf43a2b8f939531a56266be6b6176d6bc5abcb4cb415f
zc3af4e3bd4ae07a69dfa93dabadfc861e2df76130ecc312ee40fe1693412b1912cb1460ef1352a
z74943f98930fda41074b54af8d05c769e1244f7b30d3616efd4f745b57a471b9192e10686ac8ee
z502c0b4a029d661e181770f949b292f036c92a5e4ec8502a2b4475c1a0081bca3b788ccec0fcb6
z5d7ac28fdb790cc16047b0d6247706622dab1e7bf9963e4d94db5da3484c5bc76b44b307c4d7b5
z890f5dcab233f2e1e890e3806635fb2fcb190b8ffcebed8148a610b923d3e014da8117a4d0ad83
z6a61f9add43aba6daeabcaa271744b73953838d96bf91d1d8c46c94f787f324bc59014cea7a39f
z392180c5936a0695a364aed755bbaa106505e6b78349342c39a134f8eb14b950ac5a381ed68934
za790b9916eab5febd49b63fa9d7881ed33e0483648b9ff97e9f304dd75fb3d179b80c6286f6472
zb048c34124c7c5e08e6f56f41c7004306278662e3f1a66be8f293db3f4ea738a13ea78e705bd68
z9b7474c716fa1eaa406d0502e733766e1702e833ee3234eda7bd1e59fa3847a7d4c975d54f8dc8
z670f21b50efbb800e0bd6085882bd652c23b26a3c553668db92dd9c409a47f9529a66121706717
z33e62ecfc2ba7abc34195f3dda1aea5eea60d594d90cfd0abc1bb6d6b10c09a5167a9298364e5d
z4d0ef542402229507ad0b074e879177432262cb7a3087f51415be301fb826e12e518025ac322af
zd8936f3a9f5b824841a495fb7f5c8d7f4d85f74604187ab610b05a94ee18d5ae8baa10495c478d
zc8367921efd89469e390eebe48af8819aba6fa6cb06364752644266464cae9f2a676f623124b99
z4997c3b29e02dd087427127217dff983bf8c65d72646bb81f3a7e57e4d9b8ece1dcc01a5bc3901
zc0810f198f3fa2d7c4465c616b09f89b834b27c25f269c3b5e82be327108161cdd921764ee9821
zd8e7de22692e4e293f801c3c573fe25783634b7be2018ff1bf19aa9f785be5a44718f560fed01c
zbb54b0da84ea9b61ebd3cc42144fa81f9714365ca2b555137ed2a48b08927743511ced08e07cb7
z47f99aaf37f0eb13c2b0d1b80c6c54ef314220cb3596117387792b28fa8659e6792922023e0816
z1beb0906adb0d0965fd7e746238b6a55c8159da2053b9baa017970dae8d51429740520b4fd60b3
z7eca88609d9ebf9f20d607d392fe1958a36bd7e49534f877a50d582ce54dc00016e2c94c153f79
z310cc98f8daf533a6474540af64c11e2a61e4aeab5d2ed17ad7f89adce6d95898c622df00e573d
z8567aefd380edaa549a769a7d19e639545e4b2ef9a1d3d1d9fbe1daad15d275842158ba0e69f34
z843835d1b857cca6d6d7d11835bdff7c66fa67249b65120ba5f7e2f54253d34dfc8482b76dd420
z13f950572ef1d455a920b2e3a066be5ceeb4edd05ed310ca840a12d24eee8006366b7d2eddeefc
z75b101d8926ce28a7797c7621d6d9b1667acdc4503e4a77c69897fd310e5504ed45ee36d879fe5
z1c38c090f532f8f7361f89b2d7579ee4e844410cd8447945893cc63bdea18323516445a68f7a9f
zb8ea4cda7b779929bd1e18fc3b9645998b2a295d185694977617c9fcdcb4e96cf5ef46b580f52b
z29b3fbb3d100e5e7617a29786e6d28c87297327838b5fde2bcc750c10865c3a4013b471a1ff562
z14728f1f7b20a33112af11ccaf5c58a124dad18bc3474af19549964d7955ae841af2221d6e3bfa
z3a101f57cc96cc80b34991460a7e87d5cf7ae6afe6069ba360b9ea94095a5958f5d79cf21773b0
zfcd601fec7d1d6c15afa6de3eb33b619f35c4c8a976bc22bc80c5ca380644eb658725244d351ed
zf7249020fb1b605c2206fa33bb636ec06223d38f26cd57a4de26afad6db662697a49d4256d0c5e
z1b45a7b07cfe05fae5e9bf129239a37c345f8ef76ee7da4a37a22d43745cfb99aba34e3752685a
z0f3d19f9965dcc7c6049d5f399737ea6b3a74a551280a966fb370d003568f98a1cd28c2f2f5d51
zf8c19071527bd46fd6ed8b4161109d30d06561aa46dd71b87ac0c92523448e25183899688cf5f3
z0e53e192ad4f1129c3595020603160bc453ddb96e0eb0fbde31b18266a63225e0f97e445017ee3
zb615dc92ef4654220b49c856d65280141a0b4e7c1828ec0df977f18e682db570c1a14a31ac72b1
zc270493ee144c7b783849f6a7c18cd6dcd324c28fc07daf060d936f4263fc3280087f700e9a5be
z9eb66ecf66b8e9bba25fa30990373bc0452be38a36369db4eee18aced8b6abb820ea1a58102baa
za06e9c554b6aa50ca7cfc4b57f66c22b0f5fc5352bed0e0842285827db0abd4485e3917c8f9025
z4eec86db199d1cb695eb75405fc0beb70bef98739427aee3c7a37fca0b30266af91b8f89b03336
z1fdbc1cab2ece33e17d8c9b0352567cd42f1ebc6c39ead35c2f3ee8b94b856d768722c1f6b4b9d
zbdc651ddf212247674b3e1f9dcd52bcf57ebfc50c9f9462108edc6abb9b60335ecc8e5b2b19dad
zdfda3c45e5dcf4b3cc5132117d1c8e753075c093df411ab3cedb099cd8cc5b7b193a089887055a
zecdd58f389fcadf062fa290fe3f3c2fe7e16bcd1098ddaecdee5acac4dc396ed609b2976467d09
z29d839b7a01730402748d8ecb90680fcae5c2be07418d6c6e76722a919e5a6017ec183eb42681c
zef0bad8d3f7d1506de7891791bdcaa13c3f136aef748791b8e7e1990085f1d5723a4618901d4f0
z127acd4758d699eba91a084d17c22db5aa5a88459afe1e18ffd178061b12b99adb3ddce43ff804
za21dc8b9205baf9b0e119648362cde4365dd153e358a21642e424ad5ab1e3bdb228a822b9a40c7
z6cf92b7a10902de48e458ee34b5aca4920b915efebb9b1acce215a41970cbc512e5a7771765cd8
zcb0dd5be5b19886b203641607b66609ab17cba2a22c585c916317306d94c87e033e452b671469d
z742cdbe899ed5044c6e1033ecb8535331fde30db69a682afa4fddcc6bf243672d8fd3b5f0f3d3e
zfafbc3b26151dfc2af50b2cb863bab1503444242e66146d18b4b05064ef8cffd7c89c43007a479
z347518d88b9eac82a4f63b13a9e4683f993dcfd252c9227857c5044710aeba9f9ed6dc0d5b36ef
z93e6973989e3bda4fd25b1534cd7449fe41452c5c52a2cc1fb31c7c431c8614b564a691fdbb0bd
z3938f757dcac87ce1287d4c13bca8d055c474f5feeae40b9261bf8ca6bf4db1d5c9a5a3f23c2e5
z6d798732a2ff45db33d4ec26082e0a63772d9d35dff785d64627cc9c13ad1b4338779ba1573ad0
z137cfea4c815bb6cc8a3ed4965293f40544d6e8a2577095499555c33325a3d4c2cd05758d47072
zc837b26e146190821115bd8ec291310f5ce5dee0f365961f516e58fafd60133155352250d4c8d0
z95e7f3798ddf6555c134ba5b48819e114c900189b43c769b871e2fccd4017c29830b8d66bda408
z629c172e6875b2f4a3a640c27bedb660ad53aa32030431885c2f2e18c7bb9020a6b962bfd102c1
z715e05b99af4b7889b529eda3e4ed2a70b98f4efeb1aebd72ac8a6a74cba5094a1ceadd0dc9c59
za3e640cdd040da16073b24f8e1723f83242ffa9abffab6046bad5919bf77a1ad1a75cda3e7cf0f
z37ba7d66f199684ebadee32fcee611c624bfae71e2b326fbb6da56d0694acb4af4cc6b4ed12b64
z4748fcb5ca9c80ea8e504de488f1eb131abde49b3b9a1ef71d05478225dd61f78781076c45101d
ze14c28b40977767bab32822985ee8d035c6be7799027f856dd9ecca4044036fde077be52e80d40
zea48ac92deca3e3f95626b7275ba061fd21dd4eaca30c9c5d355f9d766595d3d1dc5918c07da1d
zda0d2ed8158b3bcd32a6c4f148db3d0a908c3436941a278c99331e4ef6d4eeb73c6dfd86313b8a
zbcc67c5b7a942e484612dbe12ae6b629f05c784ba3f1e66fd3f65bb80621f559f2d42e7d98dc41
z2ca7f0fe9e7e489f6f181286f40262e9ec0b016831798aeeb4a051edcb57b2b4aa3d8f0d894be4
z2060c0cd65fac8cfa32ed0d3ea58761f4a73c4b11ef571d210f8a5151fafeaf7e4d535d5ea9e0d
ze6ddeffaeac6eed19e081b5f249055965158c7ed2eb6262fc05812d4235b99e2deeedce763bb7a
zcec83652e6fb577afa0246326be72c9501fa9cccc2a7b53c0ef4d6bc233ec0f601e451f894e4ed
zcc4ab7e472ef2cab7f9fbd296f23571909206258b90f276a888dda122355bc384dad95fa7c660d
zdd501508f0a278329c4f3f15fb50e8e0aa31093fa9a960b4dec6a36db6184fb8d6c1d5fcc0a933
z791f09f47fe39ff3eab4c54e1af7811d70a82882a69bf55de2473f2de7377ac6d5aa0bcb18b65b
z894a3161ac71963ace765f9230dc52ea98a8a29b33653c3570ece9ed64e298819ebab4ae693571
zce11c0d09551c433b5ff6f028b90b81b8f49eab13c4947ad76451629276b3e325a327988569a7f
z1ae6b5ee7a1c94e3a9572df3c80d3c9735d257cfb3b43c4b236f62d663de806b7c472d8ccb66a5
z16e8ece95c98d7647fb79a51659b0ad948d628d503d963ebba369a47b844b55054597d265828a7
z384306c35678516ff13b645b1b87ba83ac6237f17bf8dd07075c94ac6473846f163d8f1879ed1f
z82cd146c74fb1c4c60a8f524d0481414233852b14b6abab938d7b7211e07f32beb234c06cf8898
z48a9a58d17ba4069815a70159b11a95d39c9fe48da99270501b0ca80bfc5b779045e35d77f0fe4
z70295aee83da0ab4a01e265500d96724dd6e4b8d974cb53b5a6bd394b9d9fd5f7f9ee1e55f3e1c
ze36973c0c258439e322f1fb2fd0714bcf2f8d046aaac0fcbeca1005b79e2733bbb2f506ae1b78b
z8690165f7b5b0ab20bfe5adf24e5ca3ac6d520640d8e64ef8bbb528253d2cb1f6749581bb6084e
z4945c7e157a0685e906f9a8f14ef8cfed9d2aaf87996a23db553aa27ee06bb9b56e42ed575abba
zfb4bdd3ccd6b6428cd7facd77257263900b257e6379f85859a2154a78c1cd57fc93f71d0704448
zc324f55a37863d39e13cca01a2acbc18393f418dbd310f427ed305dfd99911b89695b480ddd670
z783ab91e7182b61c5e88a1d0728ebb5747d49fbcbe0175c3ec6da4a4a79bb6e4faf561ca36ef17
zf0679aac0e33dc0c7eb9aa3c0879d61270e79f1f95235691dbc3d0ce2960c542602c2a029d5bbc
zea7d47c9e11c6b8cdc25923f1c9678d17866525051fe8bc96232567de60a94703f22ea242c31f4
z21153bf5b36adbd452eb1e91530ded5ee4b3089282c8b86ba09a64e2050b164aee8368abf8adc9
zf5e1c07f561be7232fbb86e710b88f2e933d392dfc7851f466f4affd2fcc5bf2f6d8d8fe6362fe
z82ba0704e573e892a1279a653dfb0cbf9b5ec49a3ff304f0d5c33b32ba6c5053547c70dcd6e894
z646c2b9973a014b9653cf8d64b292668bd82f65053d2c3e1d95319a812903d2e5a2c81fa3c0e48
zcad76c0ed2d335c2e5cb68cfb2154495f50de15b568802d4de8b3ae75a2ff0f577279cc517be1b
z36e16b4c6c632e022be5ed2030962794ce3e4cefd88caa195ab8ebe2f42d278e2c973a7cd1cacb
zc7ddbe1d3dd6c6e92353ee569c10cd4ca52a98967bdbe25dd864b4be89d2e2f1f9b1fe24e68141
zd3f072b965d68d4d89b376a531e7e3aa5e3eae2ef5c5cabad6dc0d65b4b31e426751b74555bcc6
ze95627729f6eac12d9f5481e41aece48595bc602a9e509431671eec7e588a75985dbbcce96a6f2
z3f9ae0ea7076effe7b1355ad072108ae090fb770b86d068fdcfc1a553baefe64a127d82c057c75
ze7337d7a47c31fdb416ad75bc9ec66d570f6efdc1183ae67d98e1b4ae40efee1d0c984a247597c
ze5d9a9c9989a22e646afe144fa9f5d23e78b4c2c22bd48e37c93387eff19ef0d829357cc3a568d
zbd85da34f153f212a002a2a4fff308a3a91e20b7d171d11fa9a12735763c24888672dbde42b7b8
zda218556c37d772ba43e625609e666ce0736c77e2b6272c1bc3361cced907f2f53bdda4b9fbd4d
z421319a027a8434f8b65308536a56917736c7daec053b5bb71bce5cccc8da65071623555a5d303
z87fa6f159632d8c433b3c8f51b531ca5cef4fb081b8420066b67a485fb783925cbdafb1cc8de62
zbc8396d36fe9fd7144476d1bc9af6bac4b1bc4b54253c22808ba97377e32b798535dce59d77ee9
z1ea0ac466bf61eb6b8cade275466374589cda0f5b6d39ba408fb3625b7c07dbcbc886aff6d7b73
z0354cb07d449c959285485e6ccd5a09f7057564cf39c21a5d8f53fa6b4dd158a26c5917425ce69
zc4e425ce0666dd2a05e2ee7c3a79616c8b4076fc23fe34151688f5972ffc1dd77722b6d3b1f8aa
za24a04ed2e7307e893f2ee56a54b9f9898f4caeda7a6358ae6110bde13d2b4321a307b866eca6a
ze03c78d0cde449aac247635b2a38a6bf33f918fc6240bc08b25be8585c52d02150ba5c6ab38e9e
z42949369143c2f788bd18a0f6a9832db979dbb3f40d086ff70416d683174b87b4a772dfc99a761
z7eb22b819877310ebb46d46c1cbd48598848cc63ec8b43fe777d13c57c17bc655f70bc06540e68
zee0864d62fd1b771f631ae80ebe62a9759f6f8046367256187389979432b4ddc07ad53d1ea3ccf
z40251c49f07f0a61459328590fdbc30a68d6ab00c0ac88ce35de0783acbe695ed31b233975326e
z9ed46ef24126cac0083fb6e8383d5d641b0f5e74c945e92e2c4c6006680faac9fe81b0b4648f9f
z073749dfe95f93a1aea5092b94d896e3a3d19ac6eb26860db9a943cc30b5ae0466cea711a89439
z2757e1cb1833d924848f8ebbd56e1a62cc81ad27276cd018b16a6a9a1bbb22e047c3bec0ffb22b
zb2ba160dbf233b70abf1418fee8475945da70b80a841d0a02c0d7c7763cf567ab8d03274f2ef43
z04051b2fb85a0b48d68543d3211da723922511500638c0d13a722ac996336211fe1d69f6700fa0
zd35e181c340fa3a921f49d6a78a40d0101aed176b66f6fd7f9bf26643955aba77eafe892a28e16
z7fb1f9ee6b73f0f5bc454b3d406ae9516d6d71d43d0fa8c0d4bda09cdced979051dec553226355
ze747dc108a579d2bff05b0bc1e71fb2c6a794d23e76b22f26a7604878a2cc13dfe168cfcbee9b5
zcc9e25bdf1964deea3dd71769788a7a7468eb5a0455707f243552a1d6acfc5c7921d074ff17202
zd8704f9667bb0124e1245635f1f851c1ee422c060194a1c215a8373109a6bf850c313682d480a8
zb0097efeb4f99b9e8d8981703a82905d2234f0be803f14cd775de6623d53ccc1f27f9975e43cf7
z74a1a535a9eb7441ad89dccf39c91727ed5b2d052c99a9aa11a6f62f0859512576a101bd27f996
z85d84a5faaa21d9b3eba77f3d878daae956b7f8632263c37218b39e3b1a76702078fe0a8fd1c9f
z4a4bcdcc1067a6c23db246822c118b6f51dc1b7471db4feb82726416c36359a16f148c21e033a4
zfcd91350ab11aa9415afdd36998ee1687c52597028d05df72032306269680aef120cb4081cc9d8
z655d21a2052a7654f7fa26001a0faa62e88f84700768092784aa089a9484d08b890b55d7d0b81e
z7c90417b757bbb850acdfcf04d0ec5ed7ac7152111212cacbf1ff71e14cc081eae3fd665b005e9
zeb3e2d8626a32e5d55ba1f59723844e458b36419fc3e137bfa5fd063a55088a20263861ad81c1c
z4442625fd5d00a9555164b2e7287d446c2f0803c5c58dca433dc20867e18f1830a115da7c18f6b
z17a77b382eec15d0b2f55debdce8cf18ead05e56950941bdabc0e2aa2803495004ab30cf053ba7
z19f435a9d11f2d1574a21b8d750e53ada673d905e86085a4c1ab0c4d311387d2eb43a38beae6da
zb8ab1f91ad994157d151e22e8ca345993de7a364a6cd20bdf08688db7ed3528f6822e1e474f89e
z8cdde64afee59901d1c2b742c8857f95462f408fa6d6adcc3ccaf275e67582d9b6b004bb74fba0
z029257e67ae70901918ccddac0834fa1b12a86fa11323cffd3905273730ceca7107dfd623e047b
zc355d81f44aae2ba081daa6895fde3286b57205b98e6bfa3698d9cf20c814b359b329c743c322d
z3316b3b8d69415331668e24a099105b8ffebc6f731c2bc5e8045353d9aff366ac8654673cce3b2
z7c19a336c0fdd7e15f5f4e5ed7e72de833ff2704a498db87105ca276c3df8414ca4d5cf3196af7
z16fe195b41609cd3090503f2e5f5d103e7388c3efb4c3216aab7a139962e32e203e1ff46488deb
ze9087f2859c6a7995d79548d85ed9bdf66144aa0a69c58a38e0d0109627a8c10e242e44f5d7cf7
z370d171d60a01a29d0c38212952555746d6d9d28c81cb273411cc31f143d178b35425d5ee16399
z79fce12bb350efa3103d038fb39e67169ff29fbc282fda164ad5a88de290e70393466b91d8e6a1
z18563b8fb1141fe6c2d6ac8f5e07575b841b8a5641fc8d81c5414fa52c660177faddfc523f0116
zd175ca329a72b0a4eed9a33a265a6b675e62a759b36d180c2c3def268c2340ba023b319fd984e8
zc26ba3d5cc613a5a1796d699468b364f7f32e76232894f50938fe7278a96b278e30b91cdecddf9
zd34c2ae7bcc4a8088d1e4185b0f7dce2abc99903057f09c267083d584fd22c8748983596152915
z2b07787bca293ed4e67476cf1451b67987c0beeb7ccd38a9de0bace7c869d00cd6bd8652eb71c7
zda1e0740ad2ab29bf7679d333cbb4b3d1c0c7605af1f4171717f40ab06db13f1c00dfe2b1bc509
z146fda3740ae856faa71f58cc934e59dc295f29486fee1a615395580796586418430ab22899ca8
z5be03eed9870e8cc2beb76cf4b31022332f3c80a46878177f913d82197f0c4976d3416992ac74d
z7eac70b7865981db949007a8ab58470e75384622e807d776bd7e8fa8b17bb18b7737eff7ec5941
za227884b3a56d20a40f1ceb18ebe04f11db927dbb0b5edd5a06dd9e206a0cbe4b9c5bc33cc9a14
zf2d794cbacc7b6b36ea3868ff17fc15373a7877b810372ca7aeaac6ed04cc86e18f8601d647775
zf906d912413b7befbaf8fa682d8f467c160575bccf442f9ca9890c3d86dc8c0960cf55e0adba28
zbe95bce7d18a768cd0b76f9407b53974efdd102b742b49bb9649256620f09b34f1749f96acac63
zceb7079a0fdd36e3e2b546d183d2b455c651a26e0f2390f282e2e7b4d6f6c85470e94fa4c0db9a
z75d7e7b3baba21903014b865f9a52db61c4fa6cc50955cdd77f2cdafbd575626fc0cc88f368a31
zcb759a333da96dc4dc6ffa869e7c448a9a3d642c5b5ec47afa3188c0aaa19bc9cee321c0e38d33
zfcd339b62a105ea4045070fcb99ad4a50baebe7c865d8cbd72e04925ddd83ff4ead0481ac46c10
z134cf08fc1c63eefe9b75707bb1006ec60c081395f8b874d98dd7612672ea00ea4ee0a18acb6e3
z0fba7ba522195119ab257091873de95338ee4b3e8481f2ce8a944861434d82b93e9e25749ef362
zdc1f0b8f7c91a6e54328754b15bddcc1b77ab7e3fd9eb4c26b52d9111dbf81498e3fa9caf7daf5
z11ea091f3e0db9db87b1a9fa11dd649ae7d1ba946325ce47f3b6db3948ac2642f3e1f8f56aa442
zcf75d51ddd79f846a8d0b102574599fc8a576790ed9395d5f55e7f9b189fdcc4afd981be7a1b03
z7c6b99a9c57bb0a3279854ee07898419aa811aa0af3da5adf8a405605f07acb0d97e4dd42abe5d
zc81a0bf44b3af976d6b8b4c2d3ef3847c2c71be039188c35836afe6e75a4fe0dc59a331646f4b1
zd5ad0d9aa6d25b0d962119a0314de0b50d72c5346926f91ae15aafeb10aa1fcf4dd0293ad530ed
zbeacd97ea707151b22892a69cf21b009a53b3ec9e9c622f0e87aa398bd33af37a140c1f5ec9433
zb59856b0479f57cb08a2ef400d2721c6ca0f51f27c5126d8199006b4d378814473910eb4373774
z1c4cd640c7f0f2505bedda5d0e9bcc0fa32cf3fe9e55ee7307756978cae04a82a6da2c487c2f25
zd4c4565bff5aa797b4d23063b9d1460cc58af7c39194140beaa1b01e0cb8ee7ecf032b23ae371b
zf79ff1bbb39c1f150f45e3f5f01141d5cb4381530c676338043c5ec064a26ac9c81d9bc2c8ddcb
z252361bf361bbe3e3a5fbacd58f4f5a9acc4aedaf0a1c38ee4e6f1610b2e62ba93973c504bb7d2
zc5c1c0229ccd23e367dc940be8a84e587ca6c781fd94b0defb3cc701b3da6a7a7c25686ac1ef0d
za23bc7b0af1f92588e60d1b4f4a4e03805ee43334a2b4fa97ee0e336db5657be0c2fb3b8d4dd5b
zbe0f3ce2042aec201f396acb416c46aca80880c46acd08dee4c65877ae563f15e3dc6fcfbb90f2
zb964d4696db619ae0e3a585318df58287187772868dd1727a86782ec0e210f676bcd855d77a4d3
z0584881451f2cc2e72aca2a084144a76237d811448b484f3d436ee1b932be536e5b5981debeae2
ze546e37577f2682572f698c4ef42a9c3f44b4b7d711c22f58fe40423179b7287ec26501da6ef39
z90985da6337477237a25b3b5b5f71f46a011519c63cfc579d12dcc39cd28615e9350a636935d79
z772f77bcb7069d4b7fac44a294da568bd93b36510169e4a0138aa0a5c5c40741c4936c673393c7
z25a9eb02e264ed498afd8eb04d3e57f9c2bc02f57e4d229eeb13dab042b28a0148f207cbb1fb62
z995f65c2764e95b845f4ed9f8a72a160618865affadfe219266550eec2e52fe05cd239f232db4f
zbc638f31c8bf73dd6b2ccf215cedb22640b251c025ffe08731248189909d0577febf703dae2d36
zee27cf2ceb7920aed0720650fac7b6ad3a0ec27a7784779484a16a80be82ba234d27c65d0db9f2
zf6d77f52bd88e6872afdc6401e580196344d95545d79a140b0019e036a9fc787ed790d67fcd911
za0b70ac7408245754b405b98a782bae6f7958c34e2298559eda5a1d57e1817a4529a04d8b1476d
z552a60f1724185c930a490f27b7c32beeb27ee2ea4b146baa6389d91122359bfcc84747d0856e6
zeb2395961620b11528dc36919de74e1cebf8eb62ad74324156eb1fb46efb41a9502c5c1260519c
z6fb48e2ef47e80b19f98c1bba972ec84a94c656a35cb230b3fe91fe8f349235661b9bb53ed07ef
z76e7dc5e45ba61b873c80630a5efa368bb400a8e4a2fb0de3509a2ba8b5cf869b9df5531ea406b
z86133276af7f79879dda6fa7dbfdb402c450ff32aea0d788a3b2ee7706995be860a7c9d6b608d2
z560e437875c319a0ae443a5d10f06f545d258be7015dd0a41ee8aabbba6490b6fb8f03f753a2ea
zc602c6f6c9209a61b80e678f63599724fa31a5a9dd2dda5a437c4af384dd02b168247726fed68a
zbebc1ca21e797eb197955dd054b27c57719010626195f170ee85fc83a0df5970bc3c20c9a687ed
zfb30143ec851670ef37338523b975193294d4696a28c84f2b26069ee21345fcf1c7992ec1f1949
z7c9701e21209238285c93def5569dde4b69b27edfa9baccfbacb0ec701e3da41994a1e28ac449b
zf7788b140f6e3f41a00df82f087a256587630156a55f4b8162bbf896147279f0812b9267c52d34
zaab80e28ccc3addd8e2da38a3b2127ed66781cae5d3d33502fcd6c919a9c3ea2b10e6f09813ba7
z0bd7b799784835fc8ed856368dc1971647a919c8ac64a9e338c8804b11b12b69239e61e4758cf4
z7d2570941c7a78ff789e4b8c42be32d723f90a22232d130d6678055d8af1ee765bf798abd059f6
z7079fa7ae4d5902a8d784700fedb160c133e210876e6add0a9be8c88a436b7c0c8f35fcdf6310c
z8748d0b327951a3ffddf5acb300d85ba4b48337f7140a6324260f1b934fd6155b116577e624a8c
zf7e972665e95f0bd6e6907fd1b745a75a169582a26e86f6b96db54e02a81a74de00942c8fc5cce
z9866156ebbaf85dc679df8190120d53c916a26dfd151b864881f66be6d8e379024bc04cc50bf4e
z1527ac8c38dc340a55dd00562aeb6bab2bfd1dfa2c7534b37b2e85dfe76eff4a13a36d3dc3c3c6
z7fc8339f3e8f93bc335211b90d78c6fd3e7736e1f91551f47cf86f07cb113b1957e1722ef077fd
zc0b5c33bf6b0beab0b7cb3a9365693cfe703e1d852899ca215de3fc64f40910ee9da574563e5f0
z526e13f31229f25bbc210053e378f7732d2aa0b07da1ce515e6d3b3fc85b9326c9b74f2d059e5d
zb4132d974b4968186bb852d2d28ddf1069e1ab6d180b4874acc1c8b046a270dab67c4696d921e2
z1b93a60d83abeaebc2ee7750b89a338a8617cb53335b714bc486b96b604cd5bc35147bfd92e25e
zbfb462b0531a631e1991fda1034bb642932ebc94f78a9083af39ceb36af8b3f2c0dc0d60278f7d
z0cd81d70f0ce8f202337d5d3dfe8e6acb6a768896d2e07353e4f8f2c910b63aaefa0cd17088c9c
zb112b8cd18fd8c160e05e1926e91e2c0a2e4b33e204878aee76521c8bd69cc6d27bb493e2f23c8
z7a1b3b121231f4d6ac3fccbdd821fcbe53e711ee33d7ae1895813ec6581f40545a9ed6b4686801
z3ea022338543482e5389f016496671c3f21ba80eb8717bcd8b170d535fd59e415596e3fa201eb6
z8e208654a2a0506ef8587200b134359599fff3254eec52c975d8e25f1ccca533f5a93d8fcc5e1e
z65989cc48faa11ac8398009c7885fa846265eb246328bcee0a0e372128ba9b40d660affd9812e3
z1380b0536d7e92b89397e28011d7336039772ad7db1903a49404926523194522646b75e9ac069f
z74b3e0328afc558b163c5061496e8791a21c125ab5c40bf9eef511ea4a90e6ad9935885de6c809
z60c3dc8e1cbcb6442dd8528c64132130f6f4dada5a1456301c7a2dd50a43d4507c4e24a10aed82
zdb82e110391453de155eb0fa75d12728f91f5cdc369217ef2ff0045a6572fc93a9bf5780137492
z6e92e32852e23590a6faa3884ee5295f286051a1986627c6caf8cfe6b33286c7216c9767d16ecb
z62b328cc1e20b11e53df3cceb01cd96235bfaae261e09ae3e7bd80a75d929cfacaabf6146a374a
zcf329af2c4cec4b96640953e9dc9dbf155a0eef15ac71dfb56877f10240f8d3c27e9d0640a5359
zc5936e8a613a49f2807f5e9caffff7e5d8d0e10e14ee190e3d8853728241e779513386520b522f
ze972b4786d8bf4ba938123ab1d551864bddef254a5b70830649bc45cb8070065bae56e0e32c095
z42bd199fcbb4671b1830110c21e7b334be94a3a5135703fc3f34f2130c0bb094eb928ceea355d4
z59cd5514908cb51f5f7c0344ee43474366b162ca6b48b84c70b8f096cf5cd4b58968e9d6817eba
z7e9d67d3825d57fdddcc6fe2bfcbdb7a7c99d087bad36b8caafd754c64ca1c75a7ed2d42b1dc99
z56c549d29784e75b31f22cbfaa5a3ed19dca2af138fc5b09709cf666e492f40051b8af718a968a
zf056142387e624bbd3b76c0de22abc0aacabb957755b1b7f6394d07a7e4c9335fdcbb27f085cad
zf71bbb3cff36893efb77fe4f352615fadc668291e9be7786f072d02115c437661e03d0146b00bc
zb0fb3a52ade640b897b909338b22c9443da6a7c073fcaf635703f3c108a102cf4738587883ae24
z0173a2efd4ead5ce8d046b8b64fa0c72d6e1d03149b91cd8c5a50ff7977dfd8ee7a6b4b7cd278b
zb6ea35499709fcf82e4d06ee4f07c856d46f7d47034b7267622ab5292b732777808ac85ab54812
z91458cabfca28eeeb1863f6ce82166e97197ac2fa6c43192b2a904b30048d4368741257142224c
z4645021d1a8dc6d97e4e01886160b9d6d75d7604850256179c1d484d4066869ba69fba2dd49e2b
z035b405c406eb782ff7c47bdae61c7581cbd370758ea9fa7caf9b13925c302d8fd987ec7557f8d
zadca57bef9f00a1c93ea527012fda0fafe02647e1ed4c5746700fca67bbfab2a5b812ed1dfc82b
z2c48bb71307b67beda8cd94d443645ad150e6c979dbc40e0bf9ce6b7d61a8d4b6434ed5c680358
z9123c72e667ba181776ea90efff5edd93580146408fdc3f74445faf48f5ced8f7211f29fca5472
z2e6293157956f09462291dc95048ca2498f8e5187ef3cd031b410b0b55b838ad60c6103ec36340
z5bb0ff21eac3704d065dab7f1fb113042f43734067a71e0b365087660056e85ea0e3c790448387
zebcc5163c2e351f573d9ae7f30bd9ba1a7a77e598c76ce49f96b2c05934cd2f1c7dc0521426a11
zedfdd6fa49f00847e86e6a34cec30fa29ea47a7ab548293330e57857be0ad785b7aa1fe0722286
zb40272e7528024b8961ebe90a777ed919c417660920e18f9f0fd177b79b9ad2362fae54d9bf520
z3e7080938baacb585371ecd03e59dbb95d7ed20a4c0a14157316a4f8b22378abf9f4183189a902
z8c6550b424d34c7cdc4c5160cb03b7c5e1756274606ba660d901d70d0692d408dbd390e568fee5
z481a1b9f9c60426b5c62f7469851bda4f91208cb235f9cbc2e0e5bebd7774811d5f86bc7d40abb
z42d2915b216617f77574a6b68b553d4c62170cb657ed85d7214396e41fc534504d163e7faffc26
z2018c179fe8a969d492e7e3c36b3dd41a3df3672e1ab3b6d7e95c3d78a69625babadf3284141ce
zf5bfd30c790878b8335f4334905f5ed25bd6de508f53124215bb9eeb7f08a7b6efbd9abdbf16ee
ze24cfd5b49112e006a9f52729b9a8bbd99137e072b3dfb6789077bb8884c0a854415d5d6731948
z6cd84dc3e888cf4c25da835913246c7700446db0d75c7a2d07718032d70779e2a2cb33b3c66d44
z82661a32b4e73793ea62562e05aca2c510fcd13c98170e8f12bd61778d3a29c8a42d6a3a7d749d
z28921804d196f174ff09539558243736fce44567b2fdf00654fc4f0426617ad00ed71343917453
z0c2445866282b8575e097471601a26c2da04d01cea474334ae47a354121e63830b902e8b031eb9
zd096e0a3d6df0d4c83c1cc5206aee9b96e699a092fa0e8ebba7849ad0127fe5eae0a29e26a8934
za01d95b9e16d51b8daeabf37ccdfdba9c4e53736ee91b0e516a0a735a36e8a8956f0ea0b5817a7
z17dc2ac154f6391ce8eb2b5ee5d0bc519f67450af38404c4a061806664c69f778a1e3cbd2d8b80
z5f08c8282d1b4c29ef4c556b6ce416c188f92cc1c9f97df873419b04e36b051f0907f0280f59bf
z1fe33f419ee281e55ba7f7e95b204a517e71685ba23ad989b0989d2d0631fc87a5d66294113c3e
zb783b14bac7b60e395ce723a1649a4b700a1ab5fb186ecf6065738c07ecfcaf87a972277329b79
z0f105a7240a8c83ee0f5121ebe3b08184869e1d19c987c2792c4ee3095bdfbd2e7ddb99434cb21
z3286ba042ede3e7ea43a75b23cde1b64c65c87938800855dbb1522695ab203ba94f69a066b267c
zb6256ab2fd91056786a9226c2bebb5ce79daa781f74b1fb2cec69b7007a331d898bf142432db28
zb45851462aa5b1820d43f5b7cabf90d2a0818f3d5dd9b06d3e91621869c3a89138e84399c9aaaf
zf0e2ad52c1a6a49735d6ed38964ee74ad44d1430c03a19200ce54bfa6899c28fa0e66a03a0628f
z3e676eca3cb3e139f7822128b033a61375c3803c91daad073700e48bede6f426c068562dec5d6b
z7138cdf82fb6f0d928543fab59996dcff084032d01a2997eafc22bf7374d4ea10adf4bd8d0e473
zca107cd99fc71f46f377388d53c0f1e5879d9174c49e93674418456920177196afff6e48ba1770
z56755ffbadefefc0bfd3d247736f7593575be990dd9993e31220b30dea10372f82be5eb142fe22
zd4649226cf073d52d2e7f3b7341ac39a700e7431e8cee19ea4fbc681d60cb356c5073b2256e80a
z739796553b5078bb4ead35b5ba9d0de5994b484db214ef2f7a4c0c398cc33eb28ec6f94efbdd79
z2f33c85e4281b9997bb82502d9327acfbc3c88f7b76abbf8d7ecc96b744299e42dccf05275a5a1
zad06ef741998c528e10e9c8afb5e9bafd98c452cb7e8bc20ca99531b08c1bbb42c9b71f2b72dc1
z468e687fc6a3e21c63deed7a64f3d015354847bc3dc6e4679567462b2ebfcbc00ebb70f2232341
z593b082f029da1eafc2885e128f74b2b38a40bf26581e3e842971b5edb8aa4638c31b620072e18
z113c21911f56ef0152875e339be6adf3c56f32034893a74526e4100339ee766ecb284900ff9c01
z90f8417e13e5b4f3dfbbba0da8502693a25f314039a334793a4e9f2532f4eeb860f4ea3e5f9fd4
z02461f517c824ad355ce379d83707cb84de5cf7121d001727867ed2ed8789c7a2d08239756d046
zf9b22701bbd83c3c9265e98747bf91294b90f7f72b874afd56c2533654518972f751e06cfe88bf
z9b90b6e0b8a106d77b9091f15cc6904bf222f40a65dda1b4deeace247534b228dad282b7291b9a
ze2be3bcc991451b7885f310f3aa064021176c8a0e5d22025f108a9bfd37a05b0a8e19853bfe3de
zb985092d039b2d0eb075b914343f0ff219d9de2757fc7f09ef73ed221cb358a7d0627a738f2d37
z208c44d65c1778b2c52ef13aca9e4c063de3bc151eaf6da25dc392422cfd2fbdc4707ed7f1046b
z78734309495f279889b5bbdc11318f90b9c225eabc44eaf89abcb5bf7864ff488a1b20fa6621e2
zd738cba0cc3c1e5c1c684eeb6710720b5613a48c9fb43d0f446a361a974ab1a893f515f9749d63
zb61335a7b80b10a845fd096689dd312e36664489062751d522037c1bdfb214ceafffc49766e667
zce10bcd7321964b717d17cde94bdee28425f34075be77952d3351158ba3d87b624d4633a37d189
z38abd171489c974877ea26ea8c3a0bce1afa32a1279edb8c120a1957aaebb9652696c58ba21e77
z6f53d6221b182da4c297142af28349cc56fb64e6982698b9e15758c57f3f327fe27cb06ce936bf
z4361eb2359bace3625734659f1a41a2a4a23336aedf7415a003f337170922f64d19d32f65ed2c4
ze4558e4868865281aedd38113898c3c2162ab4450c1c964fd239750aa81fa09f221ab2ebff4c49
z927f5e8c414f02209bcad27680e7dbe6b210a2eb44cf144706172f48d6f1f30a712a2cfe292e31
z36421b849513fea1831365523eac56a14c1d0254e55a99b6440e02cfb10f79567832d19854224c
zcdceab158f8fbb8bcd8534f65b46e768bfbd7d228f29f4efa2afd7daf94909e6265d39908f0304
z7cb9d14da9859b035b20d667b731b24f916340c54949f251e120db020df23e7b772ba1ef7655e1
ze1466927a6e0ba08a09d0e54071b860278b136ae2842301249cfb03cb98d536fc33c2e28ae9cf2
zf0ff18a7f418c5fd47e2a19e933ca1bc4fdae808e364b1cd13b8e9e983532d55c2af7e1b7a6215
z24bc383d11c11c39f25a11da45cf641fdbcfec76345f7187b0dcf093d25748a3f729f1e7d96b5f
z64fcd8866a288a6e74d2717ee1f0c439048da48747fc03c7f28a3b23857e61419c4864d740d69b
za4ea943f0ce64952ce37a98329444cbf5002585f480534a9df0cb6c561cb6821e6362f0a766ee6
z0aabcb2ed3b01bb2286d6640f8f2d5f418e239fff5656754916eebc1b0f0bf7103264d106f5686
z9b5134e92c75a9188ab936f515f32b6783c6837873b5f309ae565b0ed062de9d6f3388e93e8fcc
zb593518a2bd77152ed0c276217dbd58d5ddbd23cb4901d29a1993b76d85f4e15a116f93e078b08
ze13f100829f199c65db03c3e09ff354096e4bd90a1ea1168e83f2bc8de27621b3ee3a834d60de9
z9736ec2b46e86a668acaa7ec0f2dec31bc3735b637e0acafc8baf6f77bf14994578068dda8595f
zc8a98ac304faa6608a1c2ec1375b4dae76f7990ca05d2fe667f39427aadf6dc612fff9e39c0fdf
z5a422aac4c7bc0b9a0f2789fea391e16a9d89661932bbcf1e1be6e378b3fba816cccdd47646534
z03b891ce837e7b9bc995084aa00ecbbe16b0067795057c807133f2a56c1b66d40d9e5a09decd13
za3e6740fff882f288e8eccca8be09e0b6ada0c33491d2b831ec685e3dde539536871011b20e6c5
z3245f0bd799c601d8180a5e631ae210fe53c05173eabb41322cb228cbf2eec7169f763a5f1ec6f
z10655cf2c2ee9ea75c50ccf2f3757665db904e70b5ed52722ba5b3bcb48cbfcb105259e97822bd
z48273ef0bfdf2f1989d098beab427e1023160a0e7faebade17d28e4a8e89c7e6dd43d553a18fca
z7d7216878883a2d654f7833096f6163d19b368ad32bd8e0fd6b27cd7374d560a5e17864cf08f2a
zc1317edaa4afa2b1a35f909c8a4fa99737a0bc344ac0b4914bb16b6ae56aebe3a95cd3eb120725
z98ac96a0c54c6c9f010e76fef3a2808dfde5e39364520a33982fe61defec73b67df835d0ea468e
z400d86a9252bc4aeb46970a791b9f39fccdb3911d95d0e6521f351225ac4fe22e3d19e0522d743
z8aea6079dac3ff5757a88320236c50c6f55d80fd8d628d18f94724829595b5b67a61a418b4e36b
z3895ef423869570589a0c2d6df4c0e984093d4864fe2c44b136e7575a788b08b318810096ed963
z4939ebd6676f99e06fc2a6d38e09f8c9c31102d42d7a08785a51d81f7ca0c94ea64a7f96dc0894
z6f06af4b28f37014a38672fd7ccc637d68ac0f26e100e6654ab14261d573e5ea0e250574523b19
ze7dd702f3c3aec796e17962bd47ed10794a4fba3cf4e29e0284e1b45c88d0feda34d526f39af84
zee0d9e8c73722c9ff906a9f3edce4b49b768743a4be84a74fba87494d8899274b9700e20c7df48
z453b747e7f4d7ef59491513bc1bbcdfd1c50277d07cfc58bee12abf19c407d00b0ccc151130659
z0d95477d050b14c223ba471bf83a02b29492cbbaf608db2510babf75bcde38504cfbbe7bf7dd83
z89ee866fc57fc9f01f9f3426e58cf39bf1bed1e260a093e3940c54af9727f8997b38ca1cd77b4f
z748006dbf61c2d04dc91e9c4eca56b2a2a7c083f0bdd7d894a2c5ae9153139e58197257c5143bf
z859e48550604cd18e41338c62a6ba73658b38d71a0aea7ee1d73da6051ce15008a49fde97690b2
za5c964f1bddaf861c27f1078f1f429b99ccff08f1b3b7b3f8707d8661731d37509a62486ecfe49
z06c09a47b666d3e757a3049cd1bb32ebf491a70dda1f2d20d5deceafa2123fb50456482782ad2d
zbe14812f82ca52b368a910ac5a918bcdeea236dbf7da3872154dcb04bb331058fe31bd90849b50
zd2cb59579e409d32098318c07d54fbf882e5fd8804e6e3702dee72310cbbf78cc53926af9d1ce8
zc84f66e892356efe78ceb23356387625fad916df2fea548e5ccf8cbdbca76aa2b3c45cf54ef459
z56c4df34497dc8fd0331ea4a664190ed835e9196c22203c40b2bda3dbd133c6a427282011a4027
z3bf72f02efe97854a3e17135d993a7de1e4613499a22504329aa85e329cb2b03c42fc6eda7b92a
z397ed1d9b38b0b11ea663acefb43363cc74d37df8a98da5debf4ed405534e07b1f40c7ef40995e
z5fe87284c43ebadc1bd2469b2297a5b8ae866453a4a47056e8e341fa3c33ba9a8edb8fad634c97
z8dd3b4fac56e6bc48c4cb66c54205be58adc418a0a4118ed2c10c9664ba9c6a3b50296c661eb9c
z96d89ee2fb9cb7b41b3bc35bcdae0cb68e9a6fe9db38df24f52bb8e5030455ef5ed705900fdc21
zb3c47c8acdda58f88021664ed6703fb890e2147d3ee882acf60545be7854ec3bdd2d05401e2959
z820a989b71fec3bcc77ddc0737bc27543973738ed54944040c38648691624786e69e04f7aa9ce7
z201ba4c96fab693ea71750a9c67e7b71973236e6ff6bbd5473ed096a5788a4e575fca119199273
z5bec4601dcd284becab1dc42128e3118981fab8b5e9aa98e1fa3272a70e9134568d620601962fa
z897c0a925bee8ec5d25adc922b013c9a86dbcbfddeed40bf57d94904ee8ad7c35b9630444b73c6
z401053bc0f23fbbfcfa0b7b64f27d630deef3f34f773247c96afef531967fc127c37964ae311e4
zd0ed079bcbc3a3fd5370eba3cff4b6065fd98becf9fde0ee77630afadc039e9fbe8f498081e7e3
z819928ae72ce647f0b919243fc452c3d367d8f30d604bc98f2140891ec50c2dbfced141d06e540
z5bb81b363d0b72c34a09d00a06061ce5011705559f6594d1d6bbbaeb8d48da9dc27cef6b5f2996
zd4fa7ad85bb70d6bf76838fc456ba8e4e6f917be85627e087ffa82a71c1303871037e7538f86dd
zcb9d8aa83207f6cf6c097f76dbf41b511ae1704818110f5680e8f9330bc2109275ec00b46a63d0
z713276fb8b4f2f7b251dbab29b1ffac9aaf1ad4fb1b93f1de7347d82f1d2f0e229dcedc5288ba3
zf52498fb430ef72002828e282687ec237a9c3e2fc5367f0894c3a8533973e5f41bc19ad0118280
z7fdeb17703ed345f80d26de812192729cb4e7203fdc2cd8d40c693044fc995a80ea2b285b9219d
z742f2c3d25785efc7e0370851445bc6477d90a1dea3d22e7286d406740811800133ce9dee960e0
zb1637ab18d7f3cdd9cde80a89d0a2c49f1781644f0affe3372b3bc973f3f1fa02150c8b5075a8a
z3fdb050065888d8c8eebf3616e2797ad377c7e03485f34fe3bc3835b302ef67f5e3dc927f53f97
z4e59bc8f068f6b6b9547de4e9a474cf8173e56baf38e6aeacae6cee2733e698f00e6f696573b3b
z28ada018ed0c5ed33738a746a5c0d1e88b682209d1edd1ff051c4e289adc954d86a305c2b86a6d
zce345b31f9d4f8e4754e285377be66af946adb55b30e2cbbaeb7f7552f7c1a269e7da0371fe55d
z49109d5b421b51f0c92fde5cd0e6f59d1fc13e5b88ffa1ef367cd2654490022d5f41ae2d8d981b
z40a977ee594a7f5d5cafdc979c48f6887637b780b57b034fb55780d73f5dc5855e4ea02ee1a272
z041cd82cadf8b352ffd56e8fec85edb43106874bcfc5778c3bbc0c1ade0609f4901c205c76b47d
za33d018d090b0fca6f2fbce458d765a0ee6bb30c7b0a5976553b99f5cef3a71cd69c12e3e841b3
z51ad9f401a238e0fb55a97bc4b47f94e5ed840b94d902933b1ad1d0fbd25f14c2a09cd7eacc4a5
z30c12bc6720f42d67bb6fb56e6a33467f9f9a1fe6b73e60a8ec31f9ea79f46949d4c563f2e9a5f
z4c23cde74bf2717873b94c698c77a9c76baddcab63115751ede8b12ece7140d2a34df2a298fc19
z77823617071d8084685247328a0a134c9c399d36dbc7edea736aa3a99112acaeb2f32eaa143a43
z988c9281f51b32a535318f1ae79ee8cf34423197e08c852e363d1c850265db7994571b315e6a4c
za00273999e859770d9449a8677d6902dfc5b67c17d558f7a378bf54e869a24041bf12088f43f7d
z066b6bbbdd54399b9bf3500c63afc3bcd3a0062366708665758a8164de3fd937607c1175c0dbdf
z3b026a8e2cf5b7797d0df265d47e4510ef838a67b3f966f198b6ade87456a29efd2bdb856c1638
z343ee1681fb74e9983d0fbfbe9adfa310465781d881d26c72768ca1395d5da8fba8572c43edea9
z775ff33e88684c2b504fe217f30ee2bb45bccff3724e5cfbc855f67cea890a799e67c735a36cce
z9e0ba6acec053507825c7953d1417eeb854e3cc7026795f4efbd7c72235377654baf5d83b3a6ec
zb62abea30c3118f3d86f8dd77edfc6b790c2c37ab6de395dfab096d3ba7eb83a13356ea528c6d5
z947b8575a9971d8e484d23648b2bcd1633238456148bb49fe1736851c07c2597eeec8286a06588
z9db1288931b82f56c6f2c7e03b6797c8888c338f7eed47339aae3dcf97e54fe861e17521a11d96
zd67bdee81e050066406b867cdb1e9940be7c2e527459137e5e93156d4a3a200eabab3ad55cd65d
zab75abc085169fb4b2289f9a70e204f0edbf4115661e8ec73edc3d8a507c0042284350a22ea141
z724419e8e9aff36c5778e22d7570222d934c3ffa2600d782a515ffc0fdb5cdb3f306f7489c25d3
z79563d28ce4c5958916c7617ae38ed165c63fbb7fba348b665b3783e99bff6ab36a25ce0d30d42
z5c414059da3f498b6556fc7cbd535a1472cbb848f47781a8081ac15d96869e26d1ee5ec4897ba0
z1bef5d367240f40f9779a6d6d63144b5df32ad6d23bd63a12e5555d15618cb44bbcc10eeb42ee6
z7f90bef6175781935efa810cf528a0dc4c4834e8770d87538a9b9ab4c377d12b2b18cc43888ad8
z8f6540aa8843d8a4de93e1b35feb1425f5e26e8e408c29704e3ccbe2c280552c62c067c86fe1d6
z2a5f05c1f8561e180ef83d1ab3c13e4744885455c676add288eaa88eda8b5987fac898667f3d39
zefedc896a34ebe83213f0de493c33a9084dc364ad9d6ea231f781e830e2b16d130d6e38d6e2535
z46e65aca44df6dbd223b890e94c3a24e7f3a0a4d27438ee4ec0a8f3fabe1ccc74632a51205bab3
za8b65d59a80cd644fe2f80673dd2210b072c4f12c7c58d52b09d02003f90cfca3fcf1b68525457
z3dee16e003692a655da00677e47abf3bb0b5a6a02258bd8f77143f994609d8c0fb1b0d391ccf3a
z29fc2237d63f2d095971274b3e1910b45ee0d66418bec5a67628a40687025022fbefe620a4c258
z4809433fec8ac30e8cdd81ecc81524810946e9a3a1fbc5a2b514b634c245f4b8e3ca2fd85e0e42
zbb4f4da3ec855ac32a79df30b27ec004b97f1c23559b95ac5d37f396488ca11a2bb0e4f737bf93
z0f32bae9e94e3fc5ce5dbeafd7b4aa263c3a69df63ee53495140a0784666d16a8bf8802d734a67
z77be377fa929ab62edcf316819039f8525c5189eec4952cabdcc97b487959fe5d451ad2999199b
zc1f8b37d22bdf4b03dbedada6f8a8c9894e0df96ca868232801e2a00d59e690c5d86897f96f4f5
zd91b841df119cf4b37ad6194420d8f4a0999563547ce3f50af4be5147882884dbae5d00a65d81d
z6eabd30b35d9b728743f294affc0f7d76cd473575a878398c950002fc4df9af353572b88b1c322
zfbaf16a6148aff7f9c6810193bb11b6c13186a38304edda9ca8ab9f5e992279790380c7132a806
ze2a39a0a14f91042e4d813447b14d0b9939b944d43781732ebb09cf6e80c6ecbed547e2070c87d
z10130c3efebb920c8cba5cbf00482e6c816d0cf572234f99360cbd6674b66ad45aeffe92bfe348
z5c47112ff584ffe647ef01a203df4bd61f08fac0bc4ade47de7e722b19028d0952fb15736f21be
z06626bc3cb14370fcaca163e256152afc713fc35c9422a8f20be5d20b0f9958f7232c0c25a8eb4
z2a2fca0e4b13a67605408c45cefc3bc897349f6be7e52bcbbdc912f1f18ecbb448c9e8264c700f
z9d1d1a5e6281e2f1eb80a485ff2b1d58361fd8b835fe5d04af3f8bb4fc8fd6f890528fa69dcf92
z7a42b33b938711291ace679be78e6b374374cff83b4999c69f55f7f085b98aa505752c3f82f012
z370802e6b4759ba30282d755f955121d6e24db4c11755c5523c32feef68cbe194acb52cd187c27
z446f2822b1901e9985eec50f1e1b30ed1c42d07b74c545365fe0289a5f3643d0c1d0a9028bf116
zd36ff127477f6ae4f7053996baa8b43a4987bdf0e0efd7dd5e9c27a195416d963cd07951c1a283
za561db045a32c7977046592d2d7f56d3bce6239ebae25319761871f98308ce73bbd895d142a9da
zd58c1af95b0f9337bf5708dcf86fa1863b6a96f947704a38676078572cd834fc2a07d61393853a
z65312c6deeb1aae54c8383fd48cdc03bdbcbd8a4c1c9c684af48a8cc23c85aaf6031274a3b4cd8
z103eed69bcd1334a8cc7c482d7cf8df6442f2d8eaf1927562566fe9f6c16e00cbd7d8602780b18
z0bfb0917e913468f8f51e4cd7c11f94d123abdfe76022487e5da1c7a501aa252e61170477d7124
z3635219ded5209549f93cd507e5dbe4c2b64ff5c2eac347b70b0535b693d3f77fffabfb16becfc
z831c35c7376c596a7bae697c27266f3cbe0b97ebe8f419707a0a21125e316ba3ed21a7acbb91ed
z095c68961f6a20dac9824a000b6a61c8e7f8c19ff37a24e0d7a64ebb7edaf7b33e6e2380fc00e0
z5120eb0a30372760e62fee3483262a2d3d5c1925b854254e906f261c6c14e701f6db60b4841bc7
z9807fd1a0c867a2c443d20e9c7c3a133877a3c4184393c7a5f4e149561e2151664b65ea2e1b14c
z9858f3605dce1b0730c26ca324add05acbc0ecc88fd13107c066611aa46c1e8e22c8894933c714
zc8247290ff4f8d33cd5d7c365e1bac917cbebcfc88a3742d83cf71f70042077d43b658840d40cc
z18fbbdf7a8771f0694e89ef98b3b738ff29c5b58bf9fecf2ad27c4538e1a32cc79d45fa0799e44
z57613c4eb44e05ae85491d575438b86e398611142718966cf43e28522bc556a8d7ed47f18ceda4
zcc30131b11c92137ad760ab7d29e0312feb80b1299931579cc2cdbe2a4f0c58981a5d3a1b6b116
z6f38402c308f1597aa23eb383b8cae435becc8680c8f26a3e9b8a850a539b667e63bb56080cc9b
z7f7c1c5449bf0f1ee11ac3753954396dbd2d10b7cd8dc916a5cdccfc81a6f4dfeb4c0e0e2a7b9f
z1ff595c233a587416212b23eb5bcaf5618846a4bd1312ee8f4a0e845c445ddd9d043199a0ea99d
z8124b763c509d272d60465878d57d3c4372284513ec50536c160643628d5595b943c4bb85b55b8
z6c3c21351531ceb5d26c01f285f1b9fda713b5e6b985c832f877adb4e70f8872fb8de95b3ae463
zf02fa46637a6df025db826ab78392de1b844e1153157f9726d09d4efe2a52b58cd2006341081be
zc604d09743a89ea7fa4dbb703f1b3eaa7eafb3e06eb2017a7f7325cd41a7ec6e6a64cb95d2b3e8
z862d84a1e2276b3ecac684c0a7eb0b4da5217e965c7a41617703868324fede0be3ba107deb9e94
z63a1cb2ef5745388869ac5331f0f5dbb4def63ddbe8a15a1c0ace8b50bd9452bda866f14636335
zdab7f0161c08ead8e1fa53ea72303e29189cec8522e1bad51dbc01d2a5828035e5158b149c600f
zf64a11672d5354d4fe2d094bf385c7d36c6c1a5d5bd4e6dcafba3f67624ce8c910e33d9520c933
zee1c2d0ae7ec4c07792433dea6b74045b9ee8334a68462dfa7cc97ea822b87e1be3011212f661a
zebc9bc688f8b7b67ae4aff1640ab4352f8086ecfbb8f444c9fc312b88402806c7874772211f2ff
z83fc34f12dafdec95a88f0b44aba644bb99f02e500f01c88f98a860191d30c9b25a6168fa958e0
z7838d2846409e48a9d07bf3ff9a906a98cc53e2b674f00d0f2d1ce5c1bfa083f4f2e1ff47e674b
z48c195fa703c74ebf16e6e80e4f01e816f80a060d4c0fda7c1e399211e64feb20b7b974fb75c02
z4aaeedc95ad5c14c879a8e7e61024aa5501f128000fcaba9240e1ff0d820d5bee521c27fe7e974
zdb80a77a62944e7158628ee43f47a0f1e74a7ba5054bd0c39026aa4b4268ceacb1ad9b89bacc25
z641a6dd9b952d881edd6e2284809325edb5d60a741aa3d091ecb5d0d5a9ac4b494cb14909bb029
zef912714da9848cfedae470f070ffc18208f60321c0f1e967b25234f946a3f784df39c8758e2f1
z3e999fac963ceea29e718b5e0d573a3b92537b7d25ec28b3b5081c94659dacaf871ff4df3f30e6
zc9b4700caa1b6db2d18e4b7899b9a1741e8275a123d1b25c644dffdb6a0d93f9f65594e5e1defe
zafd2e3d5af5bb2616df6201af9dba6f116e4ac30a14136a974874fc7afdafad40f8a14a124b10c
z6df62df660d43a9fb3a181f4f7f1a2b98b2f24a07773785d31be414806c6c781d4f5673d652134
zffe490480a1de75b0f92cf2564e70f05678aacef52f432b4095566fe0c54869ca49e3de9e96f3f
z14feae10d2c7cfe4b3cc288766d346ce09bd503e5acd6a41c09b377bfafa4d8998d2b74293db38
z1422750d0838fcfeb322b32dc3e05eabf466f154f372c10be138d64da388f6fedbb8c150c70b37
z7851a447d9724402096cf26b28e9da8f2a828fecd09e9ad58efb8b702b50701028c2e68bfe90e9
zb9500e5287be1d469013b48c6be9f74a7dfb61e83dd1ddd4224faa5ec05a22bfd144bb9916dbd0
zc5763c566df284fb4cf10db6d9b1f0f190d5fae7bd5746a044232db816acc515ae70a5e3ba3695
z7d7ce6d6f93a48ed6507d4c91aec8ab806c8e1148eb0eb7743f0c664a374209e6bdaa8f86f7ad1
zaf9a774805ca638d726b5420d6d997884717114bec664ecf5a1da6990efdb431f6687e10a8b86e
zeef2125715930fa5fbf765c4e984f6a81b8a5763c563d8229395d9ee1d571f2b2616e8f0ae4c94
ze0ef5c6e40e0f75584df59e904e8dd60fe0017cc9e3849eafcb39c9154a14ed3638c6e70b49bf8
z8d449dafabb73218431bf55596392ad70bd1bf4e39109cafb6660cd5ce54e8135d8b05d1871d4a
z8dc42c6bbfc9d74bd39b601b2c275026aa45a24fb79f3d66ba508d4d6a6f4481ce8a190dcc3448
z589c95950419e5816cced318ff2e77b1f1311aa2300380d509bc52c9b7ac2c4ffb58d4c97b8cc0
zdcbe3c317b7f631e34b579d75447de3b4bc5e8fdc68f152db7e766df4c856bf652509b62e9efeb
z8cb903bb669ea3dd1df500f26dae2271ddf602641d8feac30ac658a7e5855e6cd754b05098bb61
zf6d89990f9c35e58601e700e36546721a0bf0d8123e4c2223a84a2651a5acfac1f52cf14a83522
z57a1510dd063603950f33b48b879676bb9a2acf251489498d35c1ac660d62985510966f9bb62c9
z4406bf70ed3f2f66933e104810e050033434aa57dc4f745d2a8957433f97605c1075b08d192135
zcd527b4e69e378c4ff536dc023f9267fd7c48883048c530ef4e7df444ed82b49218a9241a9a502
z75c249b48ec6a57b67d0dda9f8e4806b0245e4cb320796623a9654ece94b749a91af6877c87d55
z3454d1db35a0d45909c0e7432ba5552fe8228ed2e611b311e741271d68fa7da20a6bf8f5023792
z17592b56376e6dbed4e60bf087fdd97702f27fe5fe2670bb0c61770f0007c1ac6ad90aab7b2bd3
z71c7fdb03442b9c816777c4099307df48b3e762b31320fdb77614fb65bc71a4597f80acc49a348
z4f4a38784353bfb7c1f82c2b4b3461d7108215844bd2daeeb473684e50fbef3eeeb7fe39901b87
zb396d1d6a4e5196fe71f362e830f0aeb52e50f563ec7e6195edaaad27abb5c52042606ce3fb9b7
z09b84aa7a4dad8e2ae5b05705f42fa2235ccfc7d6b8942b67e1f8f3e9cd0d4c1a549e7683c1e11
z80cadfb28225f830ba5eaf3d38a159afd6bbc72a57e86012fb04456d66ae22ce74b6fa3afb9839
zf9884b1ae4322890158e93823f1fee4d8557fdc79f757dcce8269822b34f064524132a3d26fb57
z083a30807b82619db88e6ea6ae55fb5876668d2eac70fa17dca47df9df386a5d1385913e3357d6
z4897a97d98a4cd923c5e86ce441c808ac3138ed2398695de5e6bf41c6ff195a7b7e3bfcb3cca36
z91b9813308cbccf6248cc9a2536fbd7c524e23c296ff61adabb4ae5545faa3c158a1b517b4cef7
z846bb6be6ac950d28870d0cca415328d957c4893a076d3f1f65f85a633ce496c94238b6f614eb2
z42293c8c4d812ba9d6392ef6578f686d4e924303110545c69ff2f294e9f8b36e1556f5db0dc38b
z994da60df248d90e7b79588c38003cdf3df3973f50f205dc2258d7ec903719f32d70826471500b
zdf4baf5e77859492f3270b0a3f5e0cdcc38cdee8240a38017ba0aa79a08e28e261e5f7c115d6bd
zfee4e9e10cdbb7c4d032b26ce3c57d1d073c7f2d02f75f59530dd3a86e54c9d023edcbca1aad19
zedf48f0968472cad61a811e83e13b177af7c46ee83908c5a0f763d5f70fda93f39ad976c4fcb88
za272c5450fb65f5622fe08baf1d702044ffcfd5e9a0ed77b00568a16ddb12f420099da2c2bdb87
z197ad7db83d24eb244a902a59b6983eb85ea67750c9a30983808a4424b231c1b339503f9dd866e
z46eb2f27bd4a9737c373d7fa39fcd4f028d70a3acef3960b2d4b14dce9decc1ab2320cdc119733
z736c473c0a6bb7eb9925188a1958d77d03b4bc69fa9490bce7d98b14c11b057fb7beb1c1e90fd8
zd8bf0b1a12eb25446fc63ae1e89c92140980a464442d4c7251d133c4239c4a8e23794214fb4842
z700020a467a7774d8f42e58a9591e10bb3ad0470c2eaec93fd29a763b421d113e6f9de2212c11e
zd0f33373fb50e940c77f79a078f2a451553de2d5059298b2486374d30211e3c09a4c5aeb5a3942
z6494c40fcf64dec650b8e6a10b739bd0d631c9617ebd0af0b63f9a69a32a83ce69fb350141d6e2
z488565dbd0d021e884811226a059eb861a3fe5fa438b17d547bcb79be66cfb40654f834b500480
z31a8b17ff9c11b81844342e8755f77f28ea978a8bf4cfebfe442b3d2c2cddabb4b40777dd87b71
z896cb1ed8cd0212e3a07d839e6895f4e2eac4f6150dc30ffe8f91ce4c2969048ef3e90702191d5
z01bbc5ba371e4b691ae5ed950a498a31877280f6fd12363e1642779a4589ae0f571b1374ce8e82
zf458abaa089d28c7ebfbdfcd48745da88ff04a8b454d291028e7424a84498a9bd0f2f52f2963d5
z9adfa8dbc830c0cef7179a6c3d460dabac1e60ccef9a93ef98ea925381b1305d351d5e18a94f17
zd0fa9e69c8a9bcbdaa219877495c94674d62bbbe005968d279cadb131ee971b15b930791b427ae
z0247fda5f6ee4385f7d93a025d279c0d320e1fe20de961e5f774711417c656d3299e9936c0aa50
z6d4d3eae45a8babc1428d21d8a5f47bef75a2a12311ca583d78874b36e46b6e436ff10bff61a50
za39375816fd703d23141f0ab40fe53d5dbe65f924a9529b475c996373db3734db58ce88b52e30a
zabdb9b9559ed6e41d0f2a8063859b11d23a207d05b9af653b5c10d40c1a6af4f84f2c284c00df0
z9ffbde9c397ec5dd0aeda1dd5e45de17610ce57d0d5d066518e856243c992f40e431cb391cd8aa
za72423173689cb02f77a4150baddf074468bc35abc18e57844aa05da623126ce142b4b21ba096f
zfb76eeb8af9826f3393863b898cf80a65f3c12a4ecbeb2fc18e75a53899e40ae5b1a41ec1a3047
zc5e96c265c76ea8ea9461ebe3a944533f1cb61605b132be7e28b8badbee8c66d3c388ba800aec3
zf7489573599ad3657f2fd400c990d20af040da665fe79b9c01c96f234ffb267a00c5761ccbcfa5
z311425385a97a67082130c9c5733c838b52c2b0a2db326ad7c08b212f37ed09f207e9a8675e2a2
zb593507ac3e92b93726e00deb390e61bf6a5a7249150a63b28bd63b1d4fcb4a6e8ffdf95e6c2d6
z177e5fe08b90d5436c1c454407ed95fa0a070f443d9ffc292d92edfaf7363a0c4382979c574de6
z4ed65b9b9441896bcd7e690f010532eac7b84b824d697e36d611109e719dea6d1ff8bf9a7003ed
z783749c3ef7096e22e398fad050f9cbc9fe9071b3a84f2a47f3989897003f788aba608859315a9
za88b7f447e3e4ee8339183d768ba287e3eeae8b6d83f3640352879148fddf10cbc08a846e85f0f
zc3ac34fd7323b8e9532c157d2edf8def5b5d58e1f1641d50b4bf5b121ddccbc68cab2f963f6011
z506a524dc513ce1debde8b2b827181265e1f99bb2a8a7a1bb27f4fb46be45cdb3b021c5beedf9d
z5887e1a11a1e5d7fcebb06b72cc86a0457f32c3e01b81ca68e1a7d0630f347dca90546a6331290
zd41e9ec1c80b1a924667e82b702b86b1c8a3c2c1ad3cd48aaf5c12476afd8937a28b337079b13e
z34b7e33d5b26b9865005bc769022ff8a2256ff1c5286f5a70a44d7a059981a5dfb43245b8c243c
zc19453a1c9f1ae1810bd07e6d4b86d7052aba3deb8807bb949cecae4630ad2a6fb77f52770d641
zc16dbcc1c3feeb9306225d185f82ac66958582404c773926e0023490f70d738132cf47ee2388e3
z350a64b35d9d14a5bb7aa95725507ab9be324ae5eeabc48c09a43dc77547debf9d31319646689b
zf2c49ab9aec42a1a8a746417be569a33162ea5098e52bbc67a52b4a046ce587d6a4c242d39aafa
z84795fd2dce26c55ec29076c4eb7c5d5b74019bc03ba2ffa8afcc85a2d9f0c13cbc2bca56570da
z74be86c8e5ba2cbcdde374ff6f055d337f8fa216e91b5ccb842be287d92b428a7e8a70de6c39f3
za2d819b6d5674357b84bdeb1e2e54eba38f0e0fb9d67d7f02510770a71d6d5df1d44352b6acc0a
z0b09e24ef9e7861ce80c3a45b03505be8adc7bee480d633769158da115bf94685cc08838b86980
zf1431d06e5e00bff0cc05342244ab41211bb5c36ca71a4afdef1332bf1123e8e1316a1b593879c
z96ca03b4317b33d13902cdabc1dbc7301259eaf8d5ea38ab7dc83df05ef6a1923b0f0aa923bb8d
z4d1ef18b2dfc09b9b54337e27dd4b3691331f2435fc536e7b3d70a1c043d0cb94bc5ab20a0a842
za0c2b0cb7cd613c2029e1e505223b3afeb15bfb6e61ee173c0e38c804502d6ebe2ae1ee0ff4d8b
za993996f21a375aefe6f311afa4a5d1525cedac15a7012e5feb3313f6a63003b5c4983e5959d42
z59c4323f95dcae4f957b18431b4971d3a8fc754d753bc724b348f32118ba695bc21d0207ef31e3
z9473a67645b62ca7ff95e1614b7b7c29b052e3bede231f4350790b53bce81435b234ae2b414cf3
z0a8268e5c08ef437831cecb02b6494b3bce7ccf8c2f974e8079a3a7e6e1296f1e71a67b842765f
z39399426915f0cffc8f97a8f63e30ae7d0361918d51431009339f1008dc3487502c067269bfc25
z831dc1c842a51044b86aea8830715e92b7559c811f614ad79848fc7f93bd5cfe0bafade2c3f8bf
zdf5a3f9f310c210ac689bb7c317a3be05e7a027cd13c06c47610f72bfb6e957659762abf87e50f
zaf151d9b4c6fc2f2d08256495da2103716b348dc1aa0977313f0503122809647211535578351b6
z05d071f57aed86fccfbbfeda64845732dc5f1eff5d65b4a8c3dcb12d095fd71cb93ed6aa6a3b5e
z6731d04e3f113d83784c438df2919b699d798ae841bafb30bc643c697246290d96feedf4799d0b
ze936f9c07ce051f3be680516c267128c8a8d7cbcb038b401ab59471d2fb1ace2f59514b6bc2fef
z5ff1e33bf2bf9973e576686f2c4ad758577deadfa7f0468d71c12abf0a27b9f3c24ee93c75e676
zcb5ed2194d1b9bf9ef254b5bce6739f3a3e6d5fa95704aac1d2022369eea53d61bc33aba9faf2b
z2024f9c3c878004b7d2d658bc4004d70573db3d133bdbfdda3b761bdce2d54bb2cb1ca3ac94a1a
z1cd6791a2f2e2c1fe2c97d06fea86eadbb7954cefbf7ae8f8ea145f007556b60158d197e275d35
z905ab65d2954352309bccc1e8c7ede4cbc4e5362e19d5f42abe89fc09ebb1d381e31b81305e987
z4f80f28e7d6dd466d0c912e8aaa60a76d1a02a7ab9d0c6e2dc087633059e564b4e297501af2b4d
z9bbf187d9a8bd36edb4f045831b089ccc9fa3e93e826620c54651bf227665506840cfb926c8961
z681dfd3cb929c291b81d7ab13eca2e2c6410d929c20818d10f8b329f8a10a958ae7b3f2acdcd6a
z2d6e5cfdecd74f34c1ce8f89af9ec33aa19b900a439d4aaf537a16986dae15e9adedae5f01edea
z40ea8b18c0561ca13c809b216f2c1109845914b0e32ce3deeed50c144a5d372b8c731d95877933
z3dd4b3f077f96d214f03a47428e31f8b994e402aafdb5dc661a3c9e4d5712031b9ee33addbda78
z4c2e3d0976c1f47f88910c44cf73e8f7f4e9e8d05c4d003e4250d2bf1b178ef9bfdbd83edb0a07
zfb2149becd82407c9673944e13624c88743e169c447b0d4d27b04d5e4e6a29edd7810949796fe7
ze5b6bbfee696ed25d412a773c80cf4b033259a0651e9081662aa1f78d008cd46570e60b309fe75
za229fa58eb47131fe07d3f3f2c43f6a739c462e04c98fbfc140d89150094b818b47ccc49464987
zc34f08c4586464c968acb3796a8967868136231bd98cc0a28788e990ceeaafb23c399be8f14e3c
z9626899687feefc435ce063fafadfcf261bb14773422e85312d7228a38c5c1f6fb6367061dded2
z9387f0d95c1484ab0bc07a209d658caa4d9237f22470dfdc052e4ceb103ba87f9c527023f6cc2d
zfe3ee91272fccae206c376d4001c5fb3148fcda634e5ed06da797c6442771e119f71e4338c7bb3
z983fc5e0421874498b0a526867cdee04cb1a2c0dc6769121b5460d06d88945bd08bc849009cc9a
z7bd0e5de253fa1f0c24e7e0c8f9e9923c759b26f88d067c7533c911580302a63e2a610afc4e235
zc22139149c33625156a576feeae8609623fae7f49bb4bb314a7a246bc9779c4a68e5d8d4911ccf
zd691289a2efe68f85c2221313fd8e81a51e493dc44acfd3200f7acd5d8152f05a7f4a9e47a4798
z3d54da71443b4aa3f8180b39cf3ff968ec6473366d0a5180a2369f3ed4c439df67a8060a927dbf
z165e0017f90de867c093cf3d9ce5058230a9731717efc5297f6802df45c34814125036f8cd9ed6
z7454ce6f5093b23474b73b5992c2056754072eefbf0d2709ed6dac71fac494abee2fe4609d8dc6
z8bc241d780bb87ade200c0d86a71f78cb786ab3857723d4d1889f2b46254f7acdaaa091e68225d
z04a1034e20f2aad45a40270e27273817769634e12554fac3bb13e4dda41d9b45d38919cb2f5af7
z5e0640b0430332d95dfa25286635de89f6b84a3a2361366aaddd46a3d85f91e1da956d976691e1
z37e8c46b15b156c317d5b87f9fe5a8d73148e1959044adc47a6ecc698ab4108a41ee4e1438c2d2
z663cdfb2c98ba03e383ea1466d6571c3f5837d546c344609e8795d1f98042bc00a9f16656d1dc5
z8257a32a28e7170d53b90f5d5045fbe73fb687af0d95dddf330e1b73962252a5cb4bfcac9f3392
z469a59b0c0b4b9efeba396957d18596d4b82d98afc27c51220618fdb1e4f70c1454aacb34037b6
z0da1c9b8810f03685b5080c4d9e1bbd54f7c6d5c806ea2ad198ce2d0207c460b9d474a7a3308a1
z429a83c64208e3d9a98754a5653abee062d38b2cd837d63429d21d5edccf2c48d8e0186ffecefa
z9608c41cef7f28f007e154a09cb215f979a148c37fff2e101eadb5dce83939028fb6017efc33fd
z53a84d7e0275ebcc0bd91916976bae406ea87b9636062f95c18b240c30cbaf63562da443a20829
z55989967891dc4860cb95812b184a902a786a5e2acac5602a1ef6b53c8cb21e9ebbbec4b9a14b6
z302599f771c779fb18d13f7b3d5c8f2b983a0d8eb7d83529b3baf53c7c2f29e0a27116be349d83
z9f19428d2db04321446cc382270c3bcdb000facd6fd87e87423bc95dd8572b54c88b2a8473b0a3
zf248ddef79e442e60052d3d44b544161c52238e07953ee8aed57af0e1b12743a8acd8be747ad66
z71cc090374cb36cba2afc162ab753b53f2bcd61f778f7544ccf12637317bc9f54f37aeb08e400b
zdd2ea145a2dcde85c22263b615c9ebbb6f2fa7bc6d88d93b85c3c37c4b280051f35c4afeca6686
z3e68f2f92b21b335c29135bb907f1144409335d99e22cffb89e09a6515e2bf2726d902f891728a
z37f6dbdc1dd0907a4e449350b2647d1446309aacc42b50720ef189ae36fe07a36905278f9f92f6
z47f62b8dc1508caf9682d57562ad93fa9dfaadca2c22ddd19f15d534a26d74f771bbe948258896
za525fe3dd3acb2c57507795c264957aeae5e861a233662676ad9a3abbbc2e56fb52716dddad912
zd363836dac05cc54aff5720a625f11857b11226942997dc8d40658dc01443fb090d0bc5260510b
ze705fafb0104fef5ef2f5c65431660747894f4201fa362085ca728954faaeb5c57cf81d5c58c0b
z4f4ae951603ab91d02ebea256feb553007a0193c1a66f49385cb5d91e18dc7d8dd5c38a2d74136
z06054d113b00e668d82357fdc3e61ca90d8a7af8d5cabdb74cd0fa33aab49da09b889c8019d46c
zb212becbfef4d00b84fc396cfd70a0fc2ffbc22a0f36db0253bf77efff3c0d7ee763a6bbf3b799
z0beeeb0582005a25283ab7762fe27d4cfe89eb52f2889f92538507cbfc4c649ef55d1c2b5ac11e
z250bd3a1ed0049c92a77e2d478025c06a0750b1e98930f2e11505f951d61e5ec1829125e23bd5e
z233f99c41ba153ecae5e9c1ffa4961b5cee5eda0a7dec32d53ad0311550a0a57141feaa8ac9f22
ze216eb705ff312157faba83ed49cc8fe19898f440982b75c5320a4e2a14dce8cdb8936a979fd69
z5085d16f2a53b27599d3f2587388358808abc36633865f77b7b0be5144aa5287b2d003324c0b33
zf1bb14c4defd984ab46ce0548f92d600825817afe8e74d52690ea1c81ab157daaabef2b683891d
zcf2c675afb4b09fb0cded049106cca0151738087a72b53be8c8a53c12459e59485ba0dd2b289f5
zf55618aaf3a8065da9226615139846dcd8117f2af7fd8aed94f3f1760df3833cbe812da48b87ea
z50f95bc56b15187e1510e304946428785c6dc722a96fa5efd264bf95635aee61ce498bb815e8a7
z9b21cc689cab69a895dace82b19d2e07aea448d645cff75ef4f14d32946a808c0e98eb7b7fd809
z2adc4c48f0cc3c81ac6f2a484a73cc94e93fd9bdd1b8360dcbe3e24f1c154fa2698000fbdb002f
zb3bbd06674c91dbfa07e85ef620aa875512d7b07c6166145c2bf9b5a822f125ac124977ed19052
zebe04e464ce0caf5cf780402f1aa1b430d84f39ea4fab730a7ea2d28e4435ecda1dfc6aad5ca3f
ze18e9c31ba825162b3d86d24ac6d0e95a20c1fde512e24a461fa24c2d282b30c139929de2ffd88
zc57aea5fab3878146829471a4f8c0a55b817538d0f1a9c81cd019514466a4e8f2151aae6f7ee3a
z343508a46a34b0ed7a97fb496586bd8cf8b6a21a0efd3c442f63bdc71b0f9b7d974e95902beee1
z45ce9ec44ef07d4f0146413242cc576a5d0ac3c849e6223c6868835fb1764707cd65eb70b61050
zd62a42949f99c71655e6e31691c3b9171215472c5be36b7be33eebecf91c5d78d696cd34fba047
z554cfc47d16af7da25f0ddac19f6f7d9c27d1c9062b1634733c943a47adb884811ddaa19a65fe5
z399cb8f513c8dc002c21fcd7d8c0cc8d2b90f4018cf4a681b98625efa4af6d69eee210f784053b
zeaf63fdd94da50dc84671189a013c77f34ea4ac7de016348f9cd1b9a223cd13bb22d5cca0b9950
z743fc353e5ffa317a217318b6dae6f7e9d3604fda6d337a5ba1e8dc025414dd24467e52b4de829
z99b45ed79d001d098794e0b86776ca9999295a454d893772f0d77d79899d16e89261600c7187e2
z09bf14d740b9c67b68c717a2687b92a06d2c9e3f74702a4dafdf09f96906b7cea81451908cce24
ze35db119d07a76260f55f691796c0c6980282bb48ab707bcea396b577b16590a74253c0403bcba
z26f49c0b080a1d7657e5a2ea14b0aa77fc4f392e561ccd2ede298128e824c18403f1bf1545add6
z28f6dc803221ee36e3d6dd17d3041bcf40a5d6f32b8d735474c618a592fae828c1ca5de1a00e96
ze9aaeff8cd8ebd191da0e752fd20a3d4e2adde3b66aa6834c028e44b3e06291fc716a65293072e
z94ea878d012d7097ac1fe3e0f22972b89e891a115a882a3f2e56090558e4be3d11b56ac5469684
z0affdf62321bb65d151341fc8695f101286de365e46c5c239535d6d3c83dbe3aa753d605220547
zeb7c0cf97cbe10b277e4e24ccaf06027a096efd792c23a5e6901c4058852604b5ba7135282fbc1
z0d2f79db3230cd87c3fc1351ea482df2279a1ab0ff6646df6816e9b3735fd0ee59f89ad82ed19f
z34e5933462f62af3863d4976c2555a00e051e43c2fda55283be2603dc51bd035760e4f03cfdd50
z6c87580086c73064197aa6b147eff87af8cfcb29bb3613b324ec42c2fcad8e98b9ec838140a14c
zd28e8a338e13aec4094ef82d671457a2d1cb06cc5512077461630879effa9c27b02584385d6090
z5836fd60c4cd06271f0139c05fa67e2de55c1715543e0853838e74b1ecdb358567b316a89721af
zafa268f6a3ef76bbbf410a1013907abdcc58710ef2691fd7c74f9c1a37c5c1900a7a045fb039ad
zd66d51777bb9fbd99b1cc274c9f9ebb8990b30ea7551a521e2df4947d9b376df5d6e10a4695e7c
z8cecc385e9327e191d0998b17986404f9e5d6fc28a7d5b0b353f980d9741182e29ccf7d698259a
z5a81adbb70e3e6b665772d03867bd648e08aa7e8ff3aa979112bc73d2db1e9e9b33049e56b7a02
zd54a9c87ebfd33d1db4918c3e3821dffbaa6c25dcdad31d781e9f0de683126d35fec964102ea4f
z1cc77e3b7a868291b0c48056ff229bf2b41ed83ae3d2331a8d0a9e9396c3dbcd4828ba01b63ec4
zbeb936ea23716bc01f83343a985ea7864b1d3ea80327ee526222e87626317cb75f2274aa731aba
zee3cf43eb69443cb9b91241d5e8296de05349dc7bebea6317240d934a04db3937d8a3a335c54d4
zd98827ff0143496929000e2efcb7e063d0439861b2057e5516701e7b8d727de867e34f9ff637ad
zc55e3993d1c45b4f3ad03cd82444e44e6912b371ef26a5d69220beaf278e117693e60ae28fd7b8
z5cade64b60f72cb23498264dae65d49151dc321b1b2794dfc4ad190e900a3aebbe746caaf885e2
z41c424cbd1bf6ebf6589b462c22a888145f49340b67b17d4df9da452b462b26997f935a0b3fa08
z658f2472f69892c4fee8f7e555c52e445578214c1fb66d84c6b3f934ceef5237ed83cfd96c5e8a
z6a71a4feadf56a50423e4b6746af1005a527052559773d7cd2211a73d730afacd2486dfa1cda7f
z50ab587d1454506426701275650be6783a82a7ea79222e8d7701f4852a4fc29caf82d22ad20956
z4cd36e95bda8109f0eac8c28670f3523fa90d9a8fb1b5904763cdd932d7d2df64666a97973fa2e
z3338edf1497df9d35f763668bb3beb7d08b7c1a4b4090b94c70ad65952ff5ecf4be19b45e4ac1b
zae96d17bea0a2791152627ea026abeeff685fc28e144f479275e0e7e7602debedb92006c6f405b
zdd6583bc802a2efe8e7ce7f326badcdada1b3f4f0336d300d8905dd7235753076c506c9616a55f
z4169ec4b32a3329f019082edc66aaba0637a3d8ece3a035862e46778fd01853aea0fb36daca0ed
zea4515a4d4f258d0b47dbcffad957bd30db02e3635e6d039ad1723d411c91a958f482478c2a64e
z3ffe3d8034a966e48a1ebb59e472a84026d2a7cc65444d69d951c9d6890e6ca5c8ab575b69cdac
z63d30c5381e8dc5e63e4d1f26cb34a2b4ef4ef5562b8728cf32e9bea56acd10f0fe6a2d0408b9b
z6c80ad50e036ca2405ce5b1f7d117fde8c9bdaf1348f5ec734e4c80f8f7743947ea24040c98308
zd95e16dffec55bbfaa3feb73d3cf5d2a2ada4cf95a2fa75cc6b371573c057c29a61006abb125bc
zf0a116b7ff2f81e37bae4a03916679c27bb3d020a76168a1c5b1c8d807746452ae1a8f03ba51d9
z6a0da549ab7d6fe237ba3671666bb63ec1f3954cf260bd545416ea88dc2b9edd384f11efd73ce9
z05ee90f679a6a014881af9ece3f2c4cf4fcd01e0a22c21aff9b6820b0ea5e97d4407ac2809828f
zd61153c42102ea5987d4d2382ac01ab1cdb605f7edb5ba2e6039c1c3f6e40595b89fadf9683285
z4e8b85430555e526f573e37119de80208b76f233e93ac30a6576551105be4485401d9e08d7b4c7
zb8e640df899a68da13083f88f3917c2a25b3ab11becfc6a6d032362bb9424b12869e0fe00803d4
z5dca9f830e9b4e0e2a276964097468ec3aa50751ff18d1673c6c3611fc3db60d957479c5f5ca5f
z9c70c5c999fcb38c43f5b1320cc1dafb14a253edc68c732e3d1dc9d1018668a50d5f284c7ee165
z223cc293c51b8768aa8d84ddcda7326b810ac130a21f02af5ccbac814178aa6bef3704c6668ab8
zb0f1e4e3f8471f7b17120b320aa6e339a33161a8e4b02faa791d5cbd03cd5e849b21e71e4fe7ff
z190440647f14d19b91eb0cad8e553c45c0243d8a7764c74ce1eebbc53d9cad412db04cd215af68
z62744b86dfcb66cd0bbdbab90c6e2de974fcce3770b56b6923b46bec117416f993a1142490e8ff
za81cf44a509f78202eb7e8c1224626562aba2de30d5554ee4845c20677b25a2c237163eee57413
zf7e8644e99de5aec01c2294ce49be8eee0cb1c17821ae6b73787916e98fb56a24e2e7e2f779c82
za6c5e619c927f2f258833fad95f0fc006c7cb68ebcc351f5db3d64b41f0db67a565fd97b191ebe
z06a5faa8da5b136433aaa8f3124babfa777a665416eb67a48f1d6cf5ba46799a53b3e9feb8b754
ze9e041ab50d8f3424ca8eaab23458c5b8dd43b00f389ecddcee5db4b002ca33752f66213520ccb
zf98604c318c05f3f3ec909bb7d41d33e2a9ddbf0c678d4e5953ff18845396f0bf4410b9852b794
z3e974f4f8a3d7323f05f04d6578e09eb8fadd73255e71e7736d8751628d9f60f90e63f65ac47fb
z868c71bcbec09630ed9bd2cd8d6e627e37da8d98d878e496e944a3023c1b3d241ae086e995e737
z7a8545f1f560e32dcb50b5d4191a254667ae722fc50a0231b0035b8255c91b82a00a6dbfe184e2
z8243b614996a92107983448e9b1f98cdf007cc8c39b3a5b7a3cbbbde5e423a08cd1f86361b8185
z4496b7bb1fbae5c0e1c2bbdfde77dc14ba4bd472c33d1d2ae7e53cdeb80641ace9fabd9495e70e
z96175a93868b5c9f4764bc1f7f545c67416dcfbbfa4870a14442830ca36a0e9163bc581375772f
z0e4b4ed0359cd2031d6634f43876add1fdf8eb3c7fe30b5e45e6d24a0ecb580033494ce9c0a95b
z72d538b6794bf24ca8a4b21bb0b6e0057572a2b70576247a95e1ed0661d77f4f7d498ba0559c8f
z9534b9990726317a53e4deb55178d795d852f394ec08f94be65511a04beb7fe0a1bf8dc5c032dc
zac3abc13eff0fb5aebcefb8c7c5eee64bb589f7a83c3fbbc6815a3b73e88e60f1a04b701b12f2a
z9cfe9a0982e6a249366cf1df9acfc04e6799c51c496ad30db99d86f9c39ab1989a8a6de93bdd6c
zd5f345766c316dafe8a31225e620f5796eeb50aafab261b9f08aa201a68c387ddcf67c23295641
zd3dc877132090b8c51bbe1c13f4741fa092ab732790d17d452ae97fcaee0a761e04ef85d8aa513
z95f60520e4af4545a2cc8ae6a75f50bb23adc9c043f342e31389b5aad6bceeea7a006ded531f09
z48ee282819c2e21d5d73c29c0decf86dbcd85cc5801f9438f1efa810eb75e0cc86aa0ee38fbb1c
zb4c07310152a42195e80a66aa6144a19eb9fd04106b409a104db5c4bd74012dbfc63284afa105e
z40a432e1629a4dd405cadb4c8775979633eab420ddef53b6d4c40a763927119b1b6492aa031c37
z21e519cf2855609b0c5ace6c4ccdb54421bb8028fd39d89f1c893383aa9395a149cfe149d97ace
zaa3adce803fc8eb6c9f1b43ea21fc3344207b344081d8a2080f196c6101a5f098721b76d8e66ad
z59c55f4e50f64ca4080fd6cd908804812878248b24ddd78e0a60449f0a58a261fa563155612b3f
zba5ca72514e9eb1d37fc1ae05566bfa6d033f039d492d047b0cd01c3db86a97ad8559815f4e930
z495d8211066b66e5083703354f705a23b011bbc1c5a3cf999153c1c5c5dfa9b8b64b0a647a65a4
z7850a7ea91dc756283ba8d6c7837f43dfa16ec1bdc9bd8505986bf88841578e03213049087c45b
zd1fc0f214cdf8687b0376503dd4019f80e87d12f8668d812b261013d902c7c18780aa8587b0a29
zb0cb499244e65cb03d1d594dd8fd64c64987bb004ef8b8b0a824bb2a0f208e9d97321bf3b7e11d
ze0ede225e87f1b98abde1090238d67f8e246ce84ec175ff9e256ed9b33ff5241d500846da8042e
zd82e6bf41998595318f331ac606dc6b78c59d5663b3c9c7ab78a0871bf92254ff723d9d11e7a47
z49c66347c090cc8a8a69f2c8388282b25040fda50f2927345c156e03e35eddd3273c539ccd2030
za5837f35736220828a9fc9df9cf5857e1ad4d0b65eaa722275c0e3dfde9bc3debea4c35a8c9f54
z030c9b43d8b3d83181391eecc9a17b605afe9d40858abb98e729612a7e352006871d8985955052
z8c990dd247e948dfcb9b7bf8e57e13df5656a67991f65b2e918f50d83333ba30bd2fa4ba3c4828
zc1b3e5b3520a35b8f833083a9998427e00e3c6aa2b7225ec4181ecf010bcae5573292ec3e42a3f
z0a365b08dfe97d363c77a4cc038e45a4868e4f133d7e1558b43abd7326b73a250e962881584aa3
z6c2b318e19957c94d3f086d8684f062476e8b0ffdfbffe4b310585f160994f63aa8a2840c5cd99
z3a464ef9f68d8ca5a3fa1bd7824f15ebab919a1ee764228746c1839a9fb65b189a1cb7d820e3fa
z393b0fa56ab1f7ea9689788f7bbf969cfeeda42cb9ab14f2a834af9cfc34917704d81d1f59ab16
ze675bfcab99039d01f7205ef4077f6c80910aa5f360369194f477ee0b77aee3cd3095ef3832614
z03bffe122d6b783dd72d7abb9e92247ecf589f70267b77e89ba648026aeefb84e74207ef2f7ac6
zb3de056be06f70b5c054736b50cf40db358524d332d5939f17d57e38beb5a48d10d62cb0ad49b7
zd5551818098d909da797ab91655ed2c217c5f22a2e09a274968898bafbd72962d9e6f67ab2932f
z44abacb0c6670c4eda0c5b77a22f2b916f798d5376f0545369055f12573922efd1de2c4ffcf69c
z59623199c4550fcb2ff9b029785d812253b42c38eaa30164b523c001b46a1798332f02fd4f7e68
z833e2fea16777b494e20a1d586d9d1bde88f322a4060c316898377c1b56f85311e164283671b32
z1734ecf2b422f375a71d47ed92cdf55d88a46180401aa1b97be954cfaa0f94f0c5e7d1c8145b07
z7b722ecbc52b083873fb0c400d42792d0ee7eb56444b4dc774fae9c3b6e6f4aabb7ac56b1700b2
ze969e7e33086130b0917c85e44e9d77a214551409197411a5d0e7dca2ad499e4feaa55213e8349
z5dd297cc04e9720b3ff385a14bdf2f205d134f682468650279f0814534d566263597f875e10c85
ze7fed9685ee64dda417675a7c46426e56c3d32d70e4f4f7557c6cc266d8e254b32840dbda1b0ba
zed219d3db444f98fec217758404fbec1a41908c1fa4429f4a69ef3b0cfc70ee5f9827a19617e99
z10b45d0bf33f904bfdb5e086392df4353baa6b1b348464c62be5d6c2a36b5213e1460ce9a3f99c
z90b9a7b6f0a09796df9284ad181c75937446d8345de60bbacf8dd42c3437c2ad03b07700ced8aa
zdb2b12e0dab9729f484adc47887452f0f2deb34d11d61f7dcdffa762a7a94339fad62a17878403
z1ca9e0b0e8c26447fafa62c23a72daa7885c5091d25a6211393ab4dfa5ecac479a4e8341a7920d
ze93aaa179c8b6d127f2f4dfd774fa5184bc1e6d4aa580b3e95296df6e64ba352f30bf095107a3b
z75e9881e9baa1dff59b2606fd7091a515414de44cab172324908a81881b528d4c4b007cd7cf07b
z92618e90c22363d891f3220201f7faba54a051e4294f4eff17b89da0efa372797caf25beda981c
z0481f8670589eb782acebddd9fe7bfab187d72529454b3183f6371ae198fdc39c82532b066ca15
z515dea1c5996d265075438226e04815671d73f431c07e25ef02fe52fae8e68d162786d10860cec
z69d787512740a43ac995eb3b5749787e85d0398e8ed7d17ed6ef19785fb9f92b0a609c0824e5ae
zf90cd695daa957ce02e9e94574033125875fe839e0a17701fca9bdf6ad325402c8d574fbac9000
z5b63b6667b1c60e5d19225ea1af6a349a1e888f49d37a7e119018711f6ab5fdda313729baf01f4
z100c024f75a2b1c6e0fcff355e3e082aa33649b214926354369d76ecae32b2e31f52be48431803
z3f28413733b5baeef5f5e68ecc8d8f2bfa475d1e878eeba49164a96a61a8542f101426239b5a5d
ze52a0a6c6d7971eca1a4411bd7e973d786a4393d3d6903a4568dba614289a045dc8e1947a61f56
z155691ae813e7802ee2a892c6433eed1d38c4f66629ed2fcec94a1a6916ac248c4abfbfb71e5a3
zdf0ed1b8e71ab62a404892f5c2e52c2ebb4c0b67d6aabfcec7e66e0759546f152f62a8d2806378
z65ef41b38fa16218666ccc2c0da0e066272e2f02d54e2189f8c30591dc8d64631374052f8d991d
zb60fbfe985262cb0541be6e8445d4c4b4204b7fbb6ec6a85c27182e855a3dab8ba509e0ec7edb4
z9cf65c4fbd16e19f799ba23185182fcf449814861603c5270fbc5d3f7d75179b5326a468ab749d
z265dcb0aaaf5d10679daaeeff41634b9cac92d1b602a2ad749a5987304769c928a28d3eb8924aa
zde1bfa1d2ac77b3c3e86cd422779d6b3d17092bda0cc6c31a1133b8c9ce52be23884eefb7ad120
z961eb885ba42a1535923b334cd3431b69a0b4677376f5cfd01efc5650054b7d7454ffd64980c61
z74637fb0ec17d441c854006f8914c670c4b0db1da9bbb207bafa0c6f181a4586fe2834638d1c8a
z83a0b6166a37f4969e2d736f001a7b329801725fb24b9e413e7b695e9cd5eeae1cd178a3240cbe
zaec9eff80f5f251a839261e0c0fbb07851fa522f14448e20e7eb0313c8e757dc9b4d7219675487
z28af75578c5d3f157a3d49cf62e6eca9115df5bb447edf19e497bcaa43a8fc23adecb7d2e8debe
z76e184b8410d17d5a85696263313a985a53e8542773bcd77102a97c18d3452c61ae96e04e0a548
z03e4e6025aeda53ed7ff083759a4c31982b1b87cb9794b141affd6191f227ad7aca71752f39093
z1464a8c47b27af4f2723f76caeef4fe9b9b64933728eca47e885cbc6769cdd7dce774baca4bcc9
z261411a2649ebee104bf09c19f5753d2e7c6cb7aec9f8888e524fba4510edd5567088d8db99fdc
zbf9fd1e9f740b589cc80a14d870b2e47b5bbd8d8ff7fd81219ad48fdaf6d5faa486659026a07ee
z68b0d3944e4ba999f28b8790cf824789dd572b6e9eb1878df4c391ca4927a17e1ddef2a9dc7ffe
z93f50c9068ef4614e3bc37e01144f60a75556c815f438adfddcdfb291d513d10254a01d1e24125
z7f7b62c20012bc9cb3fabfba47898436837234e3b0b2aca28ded960a9d13eca2453947ede7be6a
zbd574f2a43bf1382a1d1a1a9b22114f94d18acc83b8f8c65e4c73d9d32ead1b7979838ffb2cd87
zb962123c0af28b0db2094ad2438c5c2f4dbb007089b5c71285f3e18ad3631f83ba16ea44ebe29e
zf71781a1f6dc69f419bb3aa357eb9c3ea7d50d30bec681c907c37dcc42ffd7286cb5b8b4be2f37
zf0ad661879f9936610af8c5ea2f8d3823ed76259d6669fa008cf5f2bf5311f02f83cc43b13bb5b
zacb084edd8a7ffae1a7c15bf4fe704fff635256c2e0e5a4f5e35fa8ee1f55272983d965fe28424
z6b020902ebeeefe80b8d3dc4dcb0f88ca98096983b6f953763a86123b13accca68b6159bdefdb1
z76fe68276a97e269b216f2c49c14ba7202a348620aefd48a7dd66dfdb2f134262d8362ed986c4c
zbd04d6c79741e3693cec54900d757c28ea52c275105c82071039aeb3957810bd93348f24c1c34a
zd3d5862136575281c42b3568f53f4f8eb889c6e47f0f13f5f0bbca4f5970a7d23e32565e6a818e
z07e286a558f45cf04217698e7bfd3d8bf2fb8a335f8db33f6b2b78ce3c776257afdd398c3c1cbc
z1836eebb9ef9eb238d392a7abb236b55ed269ee0f2ce9d5929d6b52789b00ff4398f8cab06ab85
z2c0d67bf6b2f791f204ad9173d83ce82df7eb0ce04a812d9e83adc5c297f9bbf651018530d8d50
z2f7bf276b1ce8360116bf38dd669da707c6a83adcf515bb779240f36b6147edc9edba41fb0f6a5
z16115bb9f5e21ffedb0ce562b6694a3157d7fdc6926c37a7d2f073dae5afdbe4571dc8f3052de6
z9e46a5cbb092623f48297d9f19a292ad9ce5ac3c8c5e1f2469afa0fdf75ddaab5f0fea4e0f9241
z04f3e75285423c4bb43f1d08c97dd9e17d2b719a0b6ce4a0a50e8abeba7f0d69700f31a11054e9
z1073184c6dcd05d7eb9008792945e3da20d9af9b20deb81724571a4399c3ba03c2830c73199373
z0a2d7d80abd38bedf9032404ebb2b2566f3e7b4e885f099080ae0f765b4190cb1dc84c75acc162
zef5960231ce2cfe2fafa0bff04c9f232e2153256be0682dc465277f69134d3ae26f89509bbf24c
ze6f5d04a30b98387a428af8b73bf8557cbcfeb40219e933390a7e30fc21e3de141e44e0c14f66b
zd9d044545fa2e50412c3860a08634cc3e69223df6e4d3f65ebc8338d36d090d325347695a222e8
z0c9e5ac8f9d2aeb7a0d0796890dd56323b3965d791663207d19c3f97da0f5cf98ca56beea72f42
z1f3f818435eb3ffbc5b89989b7a83b9a40948790b083c3d66239892c64ebd3801a6f01e0f0b1d6
z31680246182710b16bbb0ca4002b814893a01a7ba2df85d49c7ebfab5ee2f814dbb3cd8a1045fe
zecb48bfb83e37534ea3ca90432938c57a20f6237f874d4a3620732359cb668f50a7b8fc3dbaf73
zab5c9b7f6ff7d2d347de04e3f4ef501ca3a5f54a04487e94ac9f3693ef7c30003e8bcc0e06cbb6
zc84843c93289664beb974f83eb8a90fff766e87fbac961c9451ddacdb4bf0508ef3813183d4d78
z763e124c4fd739eaf58afa301e134f0834288b012d36d3bbb921e39b5e641903aa368fac603261
z3134c169dc54d10f116102b9aaa9c43ac5b19dd1f684e04695ed271ed628019a72566ba9ac17aa
za1d42c22caf26f0ecd7d62b5c0c5c0df99d901f3dfb59f1efa9fac6a582ff2d374841d1c742b0d
z8c543ffc1bd520b107eaabac3dea32b6404faed7aaac43cdcc2d8c0259fff64458ac6b9570e121
z0f0461a1ac3e9dc4a4fd1a8a529892dbe422c2a8bae36eeec3fcad938ee95d5006c7a4ce43a8d3
z54224d9edcd44d71dff0f3f38702fcd9007b9bf2a70d26f45d91f4f9891a5907de4e59aa946439
zbedfafdc4f77eedbd20b88015a2405690c8201305ef87c71739555162abc7b8b6aca8ebd0a58b3
z7815ba04ffb6e3b2a52d7c26539301555a04236880ceef05457895c092767a18a501530c9648cf
zdc842125fe1e2772b30d9b4a0a44c0e15541fb7cd2936da6277b58c8a6e27ac471f6cbb9458465
z708e7a2220c706f517e2e97adc8c8215efe839e40f0e2b6be1a41c19cb92f18bde480cc0d95b38
z5f1b07cc71bac3f29cb4ec59ee127ce2a0d7cc739c18c93a2349942e44cdeae763f01b66b19f49
zd8c3dbebb57006c8a4ca3828b6489dbf8d5094e14c04edc8c7779d1302c1fb4ce95df51cc26dad
z73915762a39c8f58a60f72e11d06d0653c3b3a0bcc4390f96454f932c08c0e41d8f830bee1698b
zfeb61cb7788d9c2290631a89583b40ab2a8b5000ac04e0b44f4a089be9d1d77c2216b9c72aac8f
z4fa4dd87404849393b157d4c480b70e3a911c47fed88da27d090e6e00acf199781cb7a4a11d227
z3365dbc16f2aa67dc20c8b6c74e9784b97e3e7e602a5a191348aed58a8900172b1de573cbcda0a
z76d062510995add6dc3fa9b3142161b2e1276303be9b2d879f5de4e629444e4a0f9c1c4285139e
z83204f7c6ac40e54dcd5251ef137189bbf009dd28a465082b44cece695ab46ef43c40f61ed6116
z1241d91ce83c9a5ccdc14f439d92210c45bf6b454e785594609d24b0276e950c137f1e00afe941
z4720468cd4c689760ffd4af8bdc843b8f92e66a1462affd1d40f0eeb5424f572d9e8599889fd1e
za8cce5eb8f9693b2f40a8314c9169331ff2eb319798a17af06133667f9b55d08ca3cf53a93db77
z1e0b6d255268414bdd9c6b4d655e0d6408d526983a7114edc547599807814f178a9abd2579b607
z422a2e33d5ad2eebc60cd98eb883d3befc3020f6d3723f4093e7f9a54acba32c7358aebef1a3ea
z5dd53821451cba2f5d58b86b85ec62ec56e521caa2694968197cc78560ed29f2196fa55f086f54
z36d5e9c9399ff2e7677499506c332c230cddc18b7b5368e806852edb645f06055aa083488f351b
z4654300934c3f92f2abb069cd7a17de5651c1285f6d6858b4a0bff88151c8af70bd6ddfd7661b7
zdcc5ee13f5d21f57ee350f460a38fd65fb6f28017a76871d7c481215cee99ae5e1fad1926ca2ae
za5e23393723076463f5b3e4842a1463dc93855fe3420275f662b8bf6c770917f12217355415263
z1b43147c92898b0592b7b862bab82ced1fc2daff7acb09ebda7c67278d44cfcce95614d3c9c2fe
z3373f8fd4d085bb1aca8a9b456785e06d5e909919db0d2c6713cb8b48c08050c43a18183847b63
z0883f48ae5c5a17c5630143c32313a06f18495c52b373ee9373194f98e81f482f1b6d2b1615a0f
z34e315e3741586de765ccd8674dc4b0d0fcfbddf14ba42ea22d691af4219e81987e2df219611be
zfff87eb1e172b24ecef00abc232d34faddcb42e1ca0c9645cbb507f169e484660ed6d6dfe0cf08
zb0336c1cb338f7f733cd5a69380bff06dd696eec325cc76b23dcd21d35c7613357af4a18f94a54
z01ce349d42e8cf7cb945dc1ebb04647be4cda87bfe53e7d1f8fe6949adbc16db3e7aeb1da7f3ce
z648d917ff0609d1b68a4d99c33aef0385ef5e4aae985a1dbb648702bdde2fddddae67e48cee11b
z7bc93fbbe2f143501a01999bb5e2f4c0b66dff546510c0691af1dc5620716009ace55f411d351d
z4aded38c3271b27aa2aa747943274439d65ea68634e812fa8543942bbba1654d149206f2d0fddd
z8d2c5de526ba096122ffefaa6969410ebb996391c0f0c78006747035380cdd7916e9bf5221e419
z7288128a671c8de9afa5b5a52f61b792d58dce62794a824dddc9dffa6115426c40659dd28656c7
z205d4cded1cdc1ab37fdb128c7d733521c6c5b74f8cfcd4d48dbdbd46fef295eee9eee0ebd5b9c
z4f57e53e2a2b0c7f71d7d0588b30361be3b3eb3740bf2f9aa7e7fe10b5796eccda3260801b2658
z8ee14cf4dab55f728922bff23080e82be8dea3ce51d5eeff17f89e4e899dab2da2b8e84ebacabe
z2e54f0ddc71716c8abea858d6ef0359cb3b9f564ce828da62ea5ba7b01348c87ce633c0717e3b4
z90f15786565d019b6137d63399e47e6d31d9817d0ecb4a31573859a00fa66efd5b1b5240806650
z7ee7af584618d3b68dbc302ac0cf6c483d67020c9681b1a81b335d016cb770333c6be77822b293
z15aa01226dd58d215fc8fc009d0da0f6ac0eaf793eecdeb0b14561f200e1586e49ad929529d383
z33e39b90015459e14de0b2b094b6db45be299537e79ab39fe0f96efb397ba06787d89b32264550
zd1fb503e70aedf1b78a12b4eb476bf46c6d11d1b84d43bad23df7ed30e4c710058b006551ce84f
zed0b28443700d08333c82fd8f68e7801e99daa77c4a0757939a769ff733069e47cf97400053f9a
z99e4b15b05bf2e04ede7af1ea5fbeaaf7e12513a2890dbaaaf5d7ed194bfe60c057cea5a6c2f1a
zcb37ae96afa74c0f652282c72b5a4ef345732d511c4ca0d410459bbf2783a251be65ffb671f174
za3b6b06f28b7cee41a3be9d79db4987305b3619201bd5ef2437afe4097bd8106c6abcdc669b5a3
z37c0c2d58378b4a2349822fdaf26f70c8e8719181ba385590635f3686a0b5ea61f87c01fed6ab0
zf29165317d5e4ce4ddbd1b87825ffc3b73d8aee81f325c99d48e6e245f1d0ba175afc2a90551a7
z2b99674961083f1029bc4a9a4e76f0f6e82e7861f4280686c49bcb7f0c84dec3c589c54eec0af2
zcb5f384e49377f89a7abcf7aab14690c428d0e1be730fc481f94a8b73212a7c5d8192af47722c3
z7639a172377b9b79f3f5723931ff80e05136bbb3d56d7d08776f433b526528a81481ddf3af5f1a
z6d8761b5bf2f809360beb31fe568e69bba737032ae5813eb3a037f27c72eecadfd5d92e0a940a5
z1d0ff8e9ff08d64a24e249f8009f0b974950a40f8652b760d18b33fcd9a24f5e3b9956c9a8cf35
z27ba2220d8992375462d7de49049b0f50aaf6de9cc991edb7cf3529a11324b2b66d3813faa455c
z38d903102d1c07e6ddbcac3fbfb0a225e4991c32beac5d119523c903f34da6f2031872633e0065
z7287e44c5fd2e15dc51e5aedba80e8ea325d2d5b32a198582323eaa03e85c47cb5e35d8b3046e4
zf848fc61e461cb0e746662d01bf7eea50c2d0adbfdc07b298a6a9d7f2a6b4c4d225d82a7eabc20
z032bd0ac13ae012a41a6d7591a5a93eaf70fc1e1823276f22915a9b1250a3e017ace1e6859f9ee
zaf607bd9f358fa4a281ec0c2666160f9835f4bd94e2ebcc52c7fe3d9f5a69c1846cd89f6bdfd4e
z2da635a0a8b6db978ea69217d8803ceb05bf36bff8718642ec0264ad8d87b4fc1cd0dd2ea11515
zb365e930d905d16ec3754e1862fe194ef0cc7687b90b2f84f825ba2b21655c7de89fdebda227a0
z176d9aa49e12b91e512b0ee51e3bfa89ec08a50036c32d5886e03f161e6ae1c956a41e9e2e9e11
z0a802652ce3424407b3a4b989cfcdf1afce53a44195130c4daa7845ca088a64ca919dbcf6733c0
z9698ecdb5c4852cb75759f8155a3441a2533d54d2fa63139245a884004eed4bba86395a24197b9
z6f0c1cc34ea0706f9f7d38f8c4692946236d456fa8ca3884f4783d94c5183636c51c32ec643dcd
zad1c2cd8cb0f2793d7da893550f32d27bc6f1f6ee2317ae40ed32bcea5ef59490192238833c1fc
z052afdb7d8a5c1bc8d1ceb4bd827275c1b64c0d8aff16e32fff171624a3b1d45ba70a2bf6c5439
z1fa740ac3a0de3665f3953a18150d3cd4f37a7a90203582246899d883dfc36a30a1cc04d7fdbc6
z6aac54770cff27b8f4342f70e043c37ee810ba5333a4624921f0a564eaadf47f907e46f36ed594
zd2fcc50957ce68da05bc0efd29640c20ed7eaf9629298d2e07d8d33ebe54b83bd71c51c57e9722
z24a060b980f3988c14c3f121bb04d35947413cd0dced7b72f3efbb837bbd58b61cb66f90cb827c
z717a2933660dc0eaee09c9ba0abb6ce44821572b99a48d8b34e8f389887db7436b01df3f34adcd
zefaddd89c28628e8c8394fe13c639d410ddf7985ffd630b4003993e14450a9532e5ec9447124ff
z4e130baa2bb02ab27517b719e8429c5ac90e1036b7054e7312890ad71072b1d5f645b9f55c4945
z6484d3f06f70623688cdcf5a51843a9014557664724a7be72e8db8c4da4393864a3097590826a3
z472f33fddd5b3acb73b6451bda86a17fa96d052e8a2690b8b4ec1d66944d08221a0ab29495aea9
zbccd4f1df4ac003ef21679e13b1acbb359a1dbb93e6af912fdd346a99055c620e23333a128857d
z1c35f0b908adae77129a09a732ec8a5f0fa36c888c9e075a80b1995fce0d3a655888d4e0ab6074
zd51490c42d5df6032508996f90f532b0b62c376979585f1044bd8314e2c232273189811d3a7c1d
z97ee66f8aa350373fe1c77184d29d2d45c5124e325cdd2cb264cdd4fa81d52bb5178799909bc3c
zb511fdd580c6d813e04f31372bf815673df40d6968eb7456435c267bbcaf4bd95e8960a9937506
z2d1841bf1d85e381de52b5de17a0cd21f049308640079455368bd5e52bc863490079ee43f0d3e0
zc63ca883f6ca1914d2b95f680535c523f1e2766f5a84595ba8c373f8e0f1637b352132437d6aaa
z7c985c7b5a53a54fc5c12d1a8278a6c29556c7f3aa1b4ce9361f51482a3d262a256f0d1693d719
zc2f02cd9735e44203ce23564df1fdb64d0f1204e9e9a2754f7425e3397ec25dccedf0fe9cf35c5
z52750aca146bc8bd5626fd915f0718e9d345fc849979c9c4e27c1081a619fc2315256215f3eb15
z49b7cecde1d37432669d4c9ea00e7f8114dee1c6efcfe054cbdf908182885ea66c28e073950cbd
z32a9326a15463ae1e34f6925d82ba981e153438270b6782a33be7560dfd161a859ce5fa8634b70
zae3d1c06f3965ee5d0bbaf4fc79194c62b77f8bd9ce227002809e02f6a1f59930afa813e0adeb5
z27dc4b6e0f8d7a37b955f74c7afe16060006d338f708a49feacde1990d02eb77caf64e798462a8
zab3cfae18827ffdd09301be3ee7e8d64ced7e0a9649abafd4d1ebed69e780f5cb05f0115501ad2
ze51832b8e195b14898d01685a508a07284b0e019ea0f61be033460ca15dc96d32935b6aee44653
z0d184a226252d993c8c98c665b4a2b151f29f8eebd6bac5c0053cc55422ea657432729f02f3073
z87dacd1973851ece0b1f9e22e5da7231afec50d433f38ff60526ef7373c27ee5eadced639e1d12
z2c85c88e00b72e94ca9663ce4aefbd3e78ae1fdddba4373b5186d66ec499975f9e7256c3de13da
z4abb64b04b7d1e43151de910ca31cdf482ca17f0b4c29f0e8351f5ac5e56d129fafddc0ad5a698
zecf9782c73b804aa94f799a30fcc96110b28af918da6f346ba7e81623e1a2e50c40d550cf57e7d
z7cb21b9843ea0a3af6384f71ff8bde14497114d359254bf388f5c39017aa97fa1c34d1f95f4c5b
zdc16710fa97eedf5c49e5375b349442940769287af389e559a2c4045af8b7f121227307101d943
z2a18b5cfa752663d774a9c5d57f30c4bcc86857c382e805b88d04c8eb3f6e961bb794edc1ca057
zf6b52fed32f4e243cf152197040e47e4c8ccb79a2e673d88ca9a227d38ecd1d3282dd851f10092
z8d7bd3c2b978a84e9222f0028584bc4d820277ef04b9632f88b5364ef66f557c4cd7fd06e23df2
z3449fc055470e7ada0c8f0ab8a5ae1539058131fed5b13658eff08c24bc38fc384690e48241eec
z86d2e9d323c7fbed9a7bf1f129150bd1740088465e1547b9a244a33c08d7e789679466830a3702
zc440b3de1c4abbbcdc4e839901bb77d780934f69a0594a106065b29fa7826d68cb898d089f9085
z50f363cfcc048349ceb62553075775098b9307af9733eebb285511253eaf678933b629109cba6c
za8961dd28f13b8d21f785d748293c9a4ad972b4771dfac358e9845f7855c2bccb81ee876eb6612
z54d308a0c66dd32d842df5d541af76b5a1743ac5399cbf0140ce1e875f5b7b6d9e3a98d20c0fc6
z785d38229278c5ccc6aeaae2188211af92451845a031c1daa64fe1f893b44de6e2d38bb834deca
z1aedcfe633a1c9c8c50b590766d18b352cbc67bb72fe94e163b65dd4ff130544638c010bb14958
z1b578ea8df1cf7ffe1e20931a908c14cac955ae8dc33ca30016e55ce9ad4306ea06bcbf8f69e90
z6eec549658833236da0cf47bd7c8a0f144f7fbcd302624e3e8a6ce03324ac4796631c36ff84ceb
z437b6c86c83874681d52d00ca013b2437e9bc16a87a2e7f549825fad4770e39d6b96faf971daf1
z04beeab37e45ee778f792ff4f97626dcb1848915137ebb93492ce962bf6a0bd169dd115d7448db
ze2a5cf7c184b128c57ac7c88886c25d12513a859cac8eb21c18eaae1d3183192d368b64981b414
zb1829840be706f2a335f18afa92cd36dfc8b6e0ee61e84404be3edf3553c462ab02aff0e08eedb
z847c0029ee20e457f653bc5f509d39eda371f5bfca0217fc472568ac34ca2e0a2455fce263f7b0
zbdbc783a816082c81abefb42001adb8db52cda89bbb7f7304fb7a8a228cf1aaf107d2d1283553f
zdcb8ea6ea8ffb7b6cfa245a4db4f725adad200829d8d7b8cd4e257f8f63e42a6447d227ee6a019
z369e6336ddd4a67536d607d1bbdff31482655290250a691bec9cf3cd4734587a8aad072a437a11
z3f38fdf749abc26f7a6f6572a22b8741dafdc97a18cff955c322b8787c2b381298d6a67c94623f
z9a1338ac1fb50c0e245fa3f0d82cff777e76ad047360c056449558eb13be3bfcbd85783b2a0936
z529ce255f61da1a6f7d16720b66eb2dbc1f6f2976bbeb2d0d344ca6322eca6eb3abba678c488d7
zd46ba161e2564a953c700d05458b81fe5f248e2501e6805bcf5a0bd7136c24aee26aee5db5e8e0
z0f31143a76bda9646fb2305bf172e43fa73f8056e31501984241290a8f7e92dd37516ec1ca99b6
z392bfdcd9a5eb35057ebc8c165199fd0efbff9c97906d54577f7554886e14b588123598740003e
z8535d7cb6f7dc303f0ff27e6d3277e82951a0c5215774c53ac16de6f2d980e7a27b17126b85c33
z9fb8ed7ad65992d1cb3b43478af51cd6b1decf7e51b37bb2ab50a5e7e4f3eff4eb2f3b425d03d0
z97ee38571e77b07600bf68749b2cd4886e8bc02b34b91a1b7cfbcea113b936eaff2e0c3bbf2cce
z21defbf751eb2403b4e574e2dd87d85769e27a4b20a4d7c149d41d9f800b9f637bb3587e70043c
z0bd30d35a4572458fe6dcecaa2e71ea93ab3c5d6f4b2a971a1ec509340b2bd583d6a84692aa483
z96aa507a847788a576bfa5c9bcc300409c3805363833ff188c23ef9f1a873eab87134f82a63fa0
z6963523c622944130be799a78929ab64666f824ba81ea205675c9e10e3a4df2d73ef4dafb07bed
z198e0c1d7f75b8c4947c18e9ac90beffbf16fef2ae31203b728fa1823b2a6e0df2e3be0720666d
z4ef2af8e6f24e24e5c1fb7062e5d994fecbf84651be6834a9be5e8fef9787c6dc755c4de817e85
z94d2d2b83511f87536af02754190333e1f6b308aeacaea7d1af03dc95d9ca324fcc01b511f1cc7
z51b4ead3c7fcfe5781f2dffeaefe5c29df45f0647f42e378624a71d60dcc235db87e0441d88e8f
zfe3151fdaa867ef02c4f1a7abce31822ce0524faf75f082f3109dd4074f452bbe4069a7e138261
z71c837e7e3925097eb122eddd75dcb4e8443b2168662af22c5e5fd3fc43a9c9a0e75841f77e13a
ze1cc4174ac58dc430bc9f4ef13329bc81cf3b70d2e35ed55af53d15f8dcf0633e5f2412901ccf3
z4fe7fac2d3a7997bad355e70277d677317ac278604a8d711f64fb17e7231b3bd1c7ab36c5eb6e8
z11670585395e84c22d9e97c97fef2e4813dbe3e44da5850565912d700ddeff95a7d4d8bc8f4d38
z16e47d4f05693d242685658b28b38ca88ee0a14c64de5902977af424e7c36711fe30ddc45bf1f2
z580b46863e857c0599640deecccc51ceed1cc516ebf1c05e288ee3c7ec150cfce7057065ccbf74
z21b8aa97b5789b29747772d9fdd53345ccb1a71910a0185232c38ce29f5efe185f7ed776070603
z4c9d0f6d3a795c390ec206c0bc5a783b8b7978ae7f39d3fd8f74c9b73f1987871a4e25d7bb7a0c
zc622c14ce92fdf1d1263ab23628d8ea72d0d3f8d6f171b84256bbd5449b92bf90cbe02276ebfb6
z2e3f300a31b0b72baf06682a06a9bddf02168b5471e492017a1b62206423873d93388047094332
zdbcd1a39cc71ac5871efcf48c2fe8defd5a8fa5e02819e5fc9853af57c25a026d2f3424f3ce5b7
ze2ac1c6e5be149f32a08a316901f483b644586286987ec3ff9d41808125ff697aa0369e1a3eab2
z32045e779dcb0ed03b098dbc914112643c6f20cc936b97da5d9e1958b229ff6724a9bbc7d3d558
zb7aba07d3ffd7258024f2d7753ec393df6a205cb1d97111a1312c4bf92c4b8c9cd4944e994f693
zaeac37688cfda98749d75c255b6a7afc8ec9bd3ed38b709b99893894a3532bb4ab465a56443577
za95b8727db858e2e176970a3fb5a952b33c0523ee78207243e9d0208684d945af514d0017edc07
z76440248d5d0e620dbc3335a318685079941afad2b1073bbf2da5e0399c42774fc11665de59e78
z5f11e080f27c5191ef8fd859bc36c42c54a354102066d60afee3b938ecaa38f34466234beb4594
z95315a68e1aa91bb10d0f13cb76208eb1f1b1d326bdc49dd33ab8ce477181f958a09ce7efc5599
z62aef3fb45c9be5b18cf0272162c6f8d9fbeae30a10dd30cb8f7858ac5c429810553ea3071652a
zb1299f0dd9e5dc2b11beb9571c9a704b65ff5775012b6f5ad81767c3c00ebafc7f2278ec95c71c
z4f71db16b071132f5142b28b548270cc96d9931a9e29f9c304aba0dd79e97dadd21d064adc72ea
z96372c5369c2b040fd187a89395b8f702a6b947c866cf7e88c1801d4abbd30d8679c3d1cdb4329
zc9bbebf2cab3387153bb7d9aeac309c42c609e902b59c58c9952dd6e866f2db9bbac48e1c30cba
z6ba3d412fc94d78121c74ec82d7c1010d942fac31003f70226c06b284fd4dae7698a32dbee8e8c
zb38cc74162c5a633d0c2e262367fcc3d22e0258ed72aa810e59a6becab05886040a1ca0300f9d6
z54882c60cfa24d7a5a70961837d143ef9a05601bedde157c1e22b4d5bd0c6712961691152e7396
z9d62efbbc7675e0f41a91450eac6b4c5c68e49da42d38e2c8282a4e3fb0274d45b798d0eb2e54e
z3343151b759d38a58e17db7e3d847ed8334a7cb982b3eb448142ab887eef58196196efdf859426
za073c96c45efbee579003e45bb1c22e0a54543a7fc8831ebc1e04ecc1ad3d28136bf9458e1a7ed
zaed77e6dbcd29c1cce90f038019f1d29bfc2a205983ce1e880f3197ec18e3c700fbb108355c813
za3aa3ef9e87c1f26596c3382255246416b6aacd0cd4631c248728576b56b34fde2b559663e4f64
z16eaad0c32c52087eccf2ff2577dc8878b3c5847a880c67a387e274ed0084f215e87471b236fb4
z8047c6b3e2d1fc8b603e46060a5dfd4b2e9338aa7eda3a236613a71a001fd50a9ad206955dd7c8
z3fdfa02c5d79f098ba89fbf75b45fa4f3d8c5a78abc97eff6d6d4f4a5d6d5d4bc8fbc874bf0045
z524b75d67249900467f01ded289b3b437c0e406164cbab07c3cb47377a69d875cb772549aa5c1f
zee7503a8be20c0939331d900bf0b9149ec3699a937ed5d36be30056167f402ce4229b8b6bc9519
z3c34ccce99d7e88f579e065baac7dece7e1e8332c8fc541ac4ff3a24c91f232534515e86f7c9c9
z142d3f3453d6d3542a6049b466f0367fd4ffbfa7445c79392df3dd1f53ef32620f776246d88e4a
z43652cd4af3cd7147476f2d7e306fb7fa0fd4f4a6da3ea2d90a12d946a22eda7007dbfbb3c5bad
z5282e2e94f99773dee94e27ddf8cc43c0c7ab88ad626052437fa0c050b2f1aabb0d5edbc10472b
zf22cf6e663a946ce710ca1e6a6eb8160f95fca260609da67372437bbfc7b44d81591cf1413e67c
z7e2b348f90ef3f12d84bb43fbbececbec77da9f165b49331b2a80bdb8bfa840a0ca51877f57400
z92da23707a5d906d31c7bc86cc391b6532a6ddb97a49eac5a83b6cc2f341cf43d07483a274d3f3
z106fcde6c6b32c119d8285270275d8dba0f828d495290d236e31aefbccad3f5b2b5671d6141a6e
z2af768e543942ca961f890e77eb790c945b3ba728777b0570298164b47d7b4ae971b6061631543
z146dc9ad762e0280ad34e5680d0ee78bc8d693ff616ebcfe1b4f0925ddb187c6a807d011e06f7e
z956a14193e8cbf001ac7e75175dead083f6d060bceb6be34d096e02266a90453d64e882012cb8d
z69ac9f2c50abde8eb42e226a062d32cb4a10b0747b07bcd43ce166a2129449b47a26bdec1192d9
zcea6c2f68e59c260348624416f58c32c7ebbd6c10e630e01eb95fb1b12f052b88d136d9e1e550a
z1630d95ebc925d2ab02f5fc316c02ff74ebe0f149d03b687d830d64669521d1c4698aacefc8c38
z2f45cc88f1d7bbd7fe8fd1747802eb54ac10130c2fa2f0e05a806390cac509e2c972fad83ed624
zdf80bbdcef15ba4ca6450103c176857c40936e313ee74d49223b2dc179c9156effb188a1785c71
z81f81132c85de4d3f9061f910d1876d8a6b4f26fe5f969e3821c9ba622a4db5b7297db4c9106eb
zebec21694668adccfcc29384a0e7e6f66b1be1b5d2fe00e95faa4b60a0e3f60646d72dc65ff48b
z61cf0392cf4205eac4945c96c85e5ff1994838a1e3956730b9101ae3d26ca1b7f7874b900d3112
z3ea8b5047f4e6b13f5a1649ca68edc78c4fd46820b833d90cc3512b850efcbce547b2a33dac596
z1ade98d1d18f475a513d13c3948e0aed2a8bdf2ea4d85bf214be76bbacdc34fa9be6b341c4cba8
za76e8e108bdf1d0e0afe6e7ac15d0b7718907558053f702ad8538289e8f4e9e33643a11d88c98e
z5cf4a7a87060e5f6669030e3a991b1fcf705ea6c32d5e05230c04028bfd6e191102630765a1052
z3b826d903822e47cf0916e0960af024cf807a830df04afd20355821c154af6bb6e3df1e4274a7c
z3101995b7e7214a97f7b2cc146a88bcdcbbf94bf34dae08a84a064563a1f7fecfcdfb0319bc24e
z2743478e0640088782ed07585ac3df86d8f3487f9e63519a44e081e7ca3a3c1aa2e13f4da21484
z1aff687b50e4bf890334b7c5a8f5e86146f831c0b59eef5fff91c97cfe69638459557069d23efa
z215f0e83d3dbcacb0a59c2d665211fc50129f6b866fadc1897cf1c3b656d55d8bf08d0296bc7cf
zd23065153b1527bcfa0c13df335135bfdbfc7d3c8bb3c1f23f18cf9ebe2c2ee4d4e00c35e3e4dc
za8d441cffd1405d6db592270bcf6f3f7aee1eefe7a96f5caec59e23d819b8681e6abdb8230f2b3
z466681c7b39413ed109df45ab25a6725075c3c5ca4182fba66d327d31d3b81d84db0306001631f
zd0a7fc0d5568dca00bceeb837687124d37bd24273823265b34add570d80bb5eb68e06cd21e3d7d
z56aff4dc9cbf5dd8b652b0dea3f793f6cfd47fd1cda2d706ae2438a8da38f1e64e18ac4cdada9a
zd0be6f09f1ef33cb9477cedfecaafc592949de2c3c872385557c9c5bdc4081c589baa34c97fd10
z557947f0228b5726d6283ae3e4b36bdc1ec0ab2f98b00c5d9725fa97f1a07463e51e02e544464c
zda0dd2d45ae105c5c26e984e390e74407190e9257e75d5babaafdaa7640ba4c024ad62be416cb0
ze08dce91e03392b4438f8c6496884d08709427cf3be17a15d1465ae0e05b0996b0c467f773f9fe
z1dbffb1001783bf97d84ed5e3ac65eb085a57f30e18138cf4b9f1065b2e2f740d66740503dfb75
z8b43098a29415295a991341885572efc8262b622131bd0a25c44064ef05b6381ff89607d0d0f1b
z42fb803f0270beec0973f28ba22d91d41b79af5390baa8437458f359c6c32e6395da96cb05c6e7
zad6175c4fe634eca2fa3cb333be13b87ef1ad2f9255468bd7e1adde5c6f30b9eb9f2c2f1b46014
zdca7fd58142cc43305617f8c69301633e49c50118a929f41230585c5e2b2910e18cc3f420590b1
z842bdd4eabef1f66ef2e31c500d033aba92d108aeebd8ee2d8b6e2348cfbefec8fe95ae4c40824
zd1dd9731b1c71f3f1b41ca8cb6a99c31f98d20e107065ad9eed639745c0e5c54525d269e1c5a90
za2539ea8abb7cf182bd0ff86ccbee6a6a9d611d3308fd3d342ef629eef1a00d9a3ae35ce83bf4e
z27cfc051523830cbb730ccaffa3bded95df27c0e3b04177c00d8f03a5ac13b2be8ed784b439cb1
z39e18bfccdcbf49b356584684e3fd39483daaed2304ec691a0a278bd46874b5660ca735af24a9c
z2122b3abbaae74ea92b0f65c9a585d869186c67c80b348af4a3c000616d58d4357f75102048522
zdba1d9e9a70a1cd81c451c7f67f79cea2674256a13948179f6d8a8cbdcc7510ae50ffee3c4f9a4
z424bf7177e7b870053a2e560aa76e72840779d466d986a8a50a08a4cdbd83cbc69de7e05215428
z8e64b2207595ab062bf9602e055cc3c6d629b9e4606d04e0c7c71a8211e4c79200d2bde6bef50c
z7dab02607c3b12598c38da2f64c6844bd2b69834a6892f396c0e63248551918e9befdb8f4868f2
zde6bcdd4706e4b806a0577b69eeb604aa49286eea05e44674ff5f0afc68cb21b8fe83272498e7b
zf61ac57efd0aa0f7ef78cc4f43375ad62bda7e09c40a98a52ff602e1c3a717ee46603354d4b5a3
zc27a4f8584eb83103c8373ec9e70cedc8b8b132ddc216e378004ba579f3c5bee170167e3012663
z262eaca21e9905214e48c6f7f3a0b212bc9417294506e91d198750fb35b4e5b5fc4c1b5e4cd080
zc21bb972eec8f1dac26968f779e7ad4530cffea3d05bcf566aeaacea6828000b9313f13ccb7adc
z6ae61bcf7ef3f9fac46b485c6288b0d55d0d1b204bae8785eb0b424424d2f53b3462b40c726f5d
z1786f727ab713cd07ab32dd2f363a7e9392965b628c6c3bf14229d6ae478278bf0789925713d54
z1391408703d5f022f8796aa021543697ead55e277a0f6b20ca4f468078aad83ffe8699f6c47a9f
z89e61bece26f0f40a67bfe6c0eee6f68b45e6c7546772c92fa8ec6983afa7c6d97e87d33b9634b
z63e375de936df8e080c39d9efeb28da76b3374d1c7066a9b5b1cd348dce983a7176353e58e23a1
zf15d87c19fcd7dfffb090977d3f7c73b96a7627f8983d46493acdfaf8715d4716c6523021e7850
zc56eeaa06463bd050a49034cf52ed6e2938a708f8408be16e79c808485033db91b9b136c6f537d
z47c6264164a19dee84d88b2841669d20b53663a3b3e967afe1feb3b6dd4dd286a9d924a2bcda5c
z02f33e11818b07ba9b5fa1027d71f561cc10fef6a003c3e392c8c27219cc99a72739c9b86931f7
zd1d05e9e02c235ea9f4c20eeffa2d89a6cc54cdfba48391d140a744035923c56890b7f3ed270b0
z00ee09adc052614be70faef56687f6096e0dae431a076d06df19fbfee042a8cb9fda045f646d69
zeb0f12634ed0f17a289dcf128ee08f0efc1cb4b78c94b71802534634c47da4da9a9df6a1887ba1
ze7aaee8b9df11eb4fad6c8293b5ec942a01ae3b9e236678272fad5d11be50abe2f0a5bfc02fa38
zf42eceef815bc6abaf4765f975573ec050aa3737c1269648aa4fe838ac668479dd65b128debd3d
zc9d08b352b37c074a445cc0df92801a413822ef91594a4cb6fd79445527441aabd737e87acd18d
z563c4e05973f04aa73da8ed5904bf1cbbaf9bb25290dcf290d1567c23b87ff7d115e1bc31ff053
z51705f588ebc972953ba398eb349fc905ec7e83f67efdc27bfcd21a101e63a9656bf9793e0c40c
zac1ec4e7084c8d55824ea644b4a63ca7bd2ffd1f0ba67cacc220747a740ab16a598ecc3b0696c1
z3d2f96e80f908ed76896afe2ac4796b3e2176a3c9b927c16a33996e9060432a31db8ce99a1dc81
za1b325e48a96a1f0325e6af67c5e2feae117edcbc04d8b5d49c2e8db8f09fa012e3607a0fffd63
zde3be2417dcf78bdabcb3c6551ade8ad1ec5e8abd4a2aa36831b109f8b24cc5a4d56620f8960f4
zd5161a2bcff03ab6dd5c0791fc71d4b7804442da7af22de61ffbd7be98d2be0e9a5ed277533e73
za30ebac09cb210d84f0d834b247b75eda125da0bed3fc14de9571d1e75c2f7e1420dc5d6fe6551
z9d16f3fb23c93b88562f1b1c315f5303fe693d8d2d1321e6d8ce4c2aef55db2fcd4412761027e5
z2e02678618d13e671ebd2d8c5c0ec1b3026f57e79787dc65cb136ae62927b0e9eaae6bb344af90
zf275ea92560c3b4e2e3d1994ec3728811bf3bc8964a0303caf8953335cefed3dee5d1a5101b3f0
z71e75610a0a06afd63c990ab63c3409a8141c4fc18e0e0b10e743fdaeb3f5dccdbd1420b2d62ca
z3be7b32f1db7b5bfcf08d18099d49abb088014b5f07cfb331f5cbc01486ffe49ec0babda83f469
z5c16be08ec1e86dd89e04bcd6c8c7956392ba66fa71cc6dad4e9761dee46a9df0466ebcc9b5096
z227ce60ff330737a5383e12de2aa7a6531c074f54b20de6db8fbf6517e66751d947bb60d5e6333
za63860bbde767f833483ee12c27da7a851167f56f80ce369bfe51bc6fa9ae897f32a305ce584fb
zd8df3ee9c3884dd616931078468edd731e096d6731f249f3725419db68230eee1cd072f1f22a75
za042161e912200cbabdfdd42172ac5e62cce31d50c9e8630f02d18e962d45d997902b2f9ce82ed
z2a422fd32f3423e6319655e6e0208b13b9e8af5147285027f42166a0383147c8805543e659e0ba
z4d4386cd3529cfcfdba5474a6295e8f17bb293e3ecdb54408a99f3592c1f8c3683d83214b3cbb3
z70f2e72bf72453bb92bc36fb51d3c6d86ad64ac25e5a721784b6becccc531e8ce657bcd9071062
z425b69f934b4cdcc28508fbec38a64da103747d65289cab0094ad87e0085fcc6cf531957031252
zf7ba20ce59486df270fb959692bb9fc211f34846d9d113926f8f97bbb5a5e3f087d886414d0487
z79a7d6c89a6eb729ed4c60f3104c3d7dbc41726057e1c506410b9c63d8c8550312655331a7472f
zf4038183c70ac6392650da06eb49e51136c2fec9477fbb49dd0ea0999541cfb6c2c05662c5d078
z3cc130102dfd56eb68dfd194f8e1309f2cb00197605cb05da70b3ebaea9147c31672e4deee110a
za59affaadde85f7e1c81be95cb86997906e32205fc4aec13c09243b13f12f4482985013490501e
z9b77a2df715443c98c72a9a87c6e96d564ca0cc6345306ad4a9ca15caa4266451ecfcdec70a611
z30ffd3556f7face4bb9a69402e8f3b7f2a831d3df7e05a9d61ac4fc450c0eda512eb7d4dd7ec41
zf0da57d0f34c418de37d6b651d683ed39dcddb7c22139d477e2117f214d38c7ca167d291b30fd2
z04c94a9fb3b1284c42321e2439c749fdf514c24a64db1defda00bd350306f4428711c58393de4f
z09ac80c1067b7a001dc5d83aee2cd4c516491a03f767c6506b8ff26b24c19a3c25bfe8b279d771
zb1127fd2c9b3a82e1038ebaee01b59d456de3dfa104983397d6f44ea33a6914d26d9b654d81349
z15381bf5c0d4be684ac3c7c6c7ae5665b398b69afb0988faeac5cee64cf90189078e29c87db7e8
z9e27dc844dccce4e61622e12f25c6d531796add82126ce7c052b00884d3ff5192af45ca6c63290
zd1c79ab6fac96807b1da3ecafb9b3f9cece8ff46a5abd4064ca48ab3051a51bb3c351d380d4c9b
zb90757e9d3d41915529a55325ac0e2c7bb774926e5912be130e25c1a9f83cebf9396bd11815698
z1675ab5a192ee5382f559effea6539a34994aea034733d209140b5be8c6f354c915b63476c04d4
zc6ad6ed99024249af35172e81d46e1212f8255f2e6f11342a12703cad476fad26db1b01d100dc4
z4e4eb606a64446c5ab20d6bf196db7cada2f6d902370035bb4ddd4f351f9236dbffff74301ff56
z2bab7afd8fc7ab9a23b82b0da9eb9285366cf7da255b4f75daf74d5ece7e5bf6ba39695638443e
zdb2d2b4d1e2e12ee34849ef34f4c204e2b9b46f9f79ef89250e59b975dd1ef06a996c5e6f575a4
zb910f9e427df99c254d1347646e075c4874e7b3dcfa5462ab2f4155ac5151cacff8125eb8b6a07
zf3019b2d1e460e9f544b518224cec9f83769bec25c91652787c9a376b7104cdb7c1c204357cd4d
z50768c59179df351dd5c95c5ec94632d803f79e3bf84f8b52b1d83aa4e953481febe18a1e97754
z5e2a858a4cca51976dd1c1604a5bef6d7fa2216120f3306b030e40bea91a2bfe626c39b902de46
zc08ae87492d171b3a9652f328f5e9bd53540037922595b3257a34841eac19d94eaf7371c14b914
zc1fd5a53208fccb666ac18b85362b5dd9a0e89b20f116a8205e60abc82450e8722c0de2898d6b9
z5ffb6da7d4f4662c1d330535bb6305a4ba91d27af0d086ceb902a41db9e3672fc03d5e6341e66c
ze4753d13a89e7a29137c7571c2113351cc5c23ed137f3dcf32991fd4ea6653194b2f0cfde5ea8a
zd5af682f61af5a44fda53c938607ed69ebe6bb43a9cb21e3e8e5b959355a32498063bab7f1c601
z6c0640d1682442211328549a1f0d9719398b6272201f99335c528aaa5f95c9be80857e36153e0a
zfa6d2a15ed9f5f8f14d592a0f8c6c8ea36052aecd8bc2d9bcc66b457bf35cb4ce029e24dd3aad9
z319c0aa7d9b125cd2231be6c5394220344d64867bc1c24369a2cc135898edb26096e0c4a1e9439
ze0259311b425f30780af7c2428d02d120882e39524054ecc5284c92d8cede46bb7bac5173c95d8
z0ad9c98e67b42cec0da497cd9520d18519872e8aa6d1613628e20c0aba493c600afbaba0957aac
z2522f5df5250c228d9deb7d8b18eac74a5e93141f4f1648a55b3b1a053548db1b1df74ce02290b
zd2cae0484d5104777de4d0ad80b85d9ed381fb8adbb5a48cb93e51ef003fb0d7291e5309b4e0d0
z7de0eb5223379bb59bbd4bb2cd51e691d200b86058c2e4ef5b9c8e3bb545e1fdffe69c8ecade25
zd7736b4488e6319ce6f12e3102efc3192d48310535fbc4d6539b3358bbfb4e62b33569b3c9f25a
za9334ed32b9054208617e674311dc2940273c960fcfb8228728415bc91b96b204b3dd7d85ae548
zcd7d372e13fc89c06a2e0512fbfd2bd86701bef391b256d9079f28d83d1577b276c57a5b7dbe21
za69c9d7de3581d44addca040ff7efd6e957d55065f119287435f7b6e2d10e42cada1173741948c
z9c44bcc5172fa7da93522d8c3094eb232c3d539271da222ecc8a4db85c276845f9534f3c5cff2a
zeea3ba710d7474092a78b71a7e5c58b6f967d3de1665829326a111dc95ec3b86b764f63a1636b7
z2cc3e72aa5316a44882f20d3b43e18e334f97f9f97711d8602630225cab9999d941d7ef4a91009
ze11ca80648ea60f9eda120da77be12fb17c19f43a70d2ca385cd4b15404159bc23dcb0312b3bdf
z28cc1117f24ee149892727bb39669c2903f89b59137eda4bf7cb3ab414d9e0778094283c8cc009
za8cf8b611c07ec85c5397dd379fc1299757937c1458752f4aff0e67db663ead7297a26e258433e
z59e1e4a356631ac2479c7a50beb16bda6df0d661eba590ee311a20da6ff7a8d4db8f5f4262fc4f
z4b51aa442bc7208528ed889b8cd1f34e469d082590680bf8c726f83f9ae1bd92c6a0c9e60d6196
za7e4cb26f27a116daa4b36280e0fb8590043df9da1aed37d2696ba2f934aea6c096bd230d76237
zc1316d3451e2b4e30df041008ba9de9bf39296c947cc785da24574ed0ee170a4448056e3e74d75
za089905f54fdb527ea26a2bf4b958b84c9f7940ac7617d856484c62bb2132154571d25dd1af753
z833a5fda950788bd20f502e7654752e45aaa18fd8e528f804970d900d0d5b704c57accb13eb7f9
zaedc693fd6ddeda86b91d39e7aa30c1e9b6618a7331b5b4b78028c22986b8d6749cdbd7f903ff7
z956ac91191a7e531316df313f689aa7a0020336edbf9666b9dde4c2e32595b2e4c0ccfe72d92f6
z46303592488fd9478f8819013f70c4fba480f6f97db64f83a6423e1adc569372869838866f08da
z3f21048f3a2313fb787e6bbb70c24ceadd5005027b13068490fa5ce478c0c9629a0caffe070a59
zfcd4c801006cef6867ef039117b599348d8aa36ef4b032316254ddfe264875469ebe3d68544073
zef57f6545c95fd845d5762daac7fb1ba1e8441feb0dc9e8f0700ffb336322f7a49f14eae11ea26
z553c802a5a9234939a0b4b796767f1805e5449bcbeaf7cfb926cb45448354d51368c935d922b38
z8a4397f8ae41033bd7ef31675d8152678a8a460134ab7bbc4041892e9ed9e80e4908cacc304123
zc28d6b326da415625518efdf79c7bd6fb640ea42f6397279118b348b77003b15a1b5c8d62db6c0
zf679bd7a795a820f28997b075f606dc68af2f9ca2b6133cc0d104f6e73d13562552a62da79a20d
zd3dffa12d3c6232d87ee80933afb02cd580928ecaa13d4f36191517194b6c95ffba03cd6564b3a
z16b3a376bb71ee61b6cd03d3bab08c7083df3cf88638676508a749b10568e6c862cafdd2d4193a
zb81ed6e841bf30234d381afa065d542122eaf79571cde3bb5555ceee3daac781705793653f59d9
zd2d2ae100901d921f708ed776aa2548e9d97ad167f24cc9d4739be7a671e1d5f5b8cbec0630f98
zde13871e045b4189113cdabc254b3d270975372b201c11f27a20e8d54b45b1b39cfbda74b8fc54
zfd8a0baba22241dea8222f53b49aec6082f3b429d3e5fba8656d113d9bf6d31959009071e1f592
z2576766c9e1839ccba556db1f8be7cbc2f32b63ea1fd6805b6a7f48bf229bc07e53ad9d9c1678a
z2b893b76fff9d47b8bc72062d7e97094c6bef9ab64339bddb1bac5386c5c790e85769c9c472979
z71b9a27379f9d1b0ff1266a732e0cfa2cd8d5d6b3b046b1ea563d47c77dca9c6204b81e4a43161
zf7878644260a6c38a33079656434b2ec7c1b19b1f0bf2faded5c590cbb540063171d123ab38b2e
zf30e26da31e953e7b05f0432ef9d4acff1fd9276e37b17f1a9c1b29c607cd4cc3bff2ba0fc2809
z5007a0611cee4644dafdf2857a960d82b4344c0532299c91394cd2af4196dc244bd7a0370cbe6b
z3afc507a963955f0261a93ba8296c9b77279ffefee30efb255eee9764c4f493296d89012541b43
z120f3ce4630294cb4e0034b54242abb99f40a61a21764816e93f7dcdf54495836682e472ecce19
z468a165076abee1cde4fcdafa48819e1d872996eaa2574fdaa0bd686c5950e9079945655d30485
z67f6636cc700491d34abf6997849ea95a14c57b99ad5f70f09fa2c83bb431fabfcfb8b7d8b5812
zc55ac46023655481f4b01d36c4f9d8fdbb27302d5e1cbf7d5cd9a1c8edb6939d0e8e64edcc0e71
z16a3be76c1d44dde2072ed2bc902a3fd4b1d1792641d149eb4ae7d99f8737b033b508a97101671
zec890e69aa2feb3e4dbeb3356afae836d02e2c06e9a7a48a8c34502974a5fc405a86c883514bb7
z2d9d139a44befa08db79846894c31cd8a227b6b208c1458cc414ca3b558e7fcd63d73280b789a1
za43cf3e7352e461701c0b9766f02628c72f04167bdf30cb4401c15c3174851c32169a0ca699da5
z78e19e0e263957d777830b1b48e23527a861124d3493b8c17b8ceb905ad581d633a21ebaec8922
z85f34c8ba832482d0c70a60cd7b99b23a23dc71a9f87992924a53be77f544843eae40e057fabfd
z280409a47a07e6583aa0afbc429785730806f067e1a7a178301a58bec259c4b6e650131f287e30
z7c618a9c11a79a46128258e9c5b2e0b05b5af544f1a665fadb209d38ba7c454294c4adf19e8fbd
ze062c5515f1595d0b887077d83887cbbdff9b27e79e6995263f4bcb1709ce084f98eb7b16a358e
z2b71b3ec12028ad44af8c2c5864fef984fb065618c5af5b69f515493febd85c8ef1411381906a5
z8c00f000096aaef95861d9a5b0b90ef427eb64e45828c4f30bc381170f1784fdad4641fbb6e1a5
z985cec4fbdc2d7e00284c9e887133e5fc617f6c258e95e1d1d83d19e6dc1ebd341a580e1fedf67
z30182ac44ec7cb2934e00dd1f67fd90f8555460b156af4cbafb5ab418549547de2093cd4088941
z0fbec30e23b932b9921db59a5c2efef92eefdf26ce49ce7580b1d029c1758c025c5148c69403b4
z0e81de19dd2b7af7e692e937c7cd09a383aa344e3d87b2a7aa7b7f816c4370d63b7c705926b45f
zc2b85f080cd7c898695863811809e53e17b3791c97196512fc3c1cc6d1c41c6ed7f87eda523b9b
z6153ca3dea3714f20a923a389f61ffa408c5df3b56fd3ed32a0c42fed73f8351f59fdd4c0b8f3f
zedd78efe888b53b5bcb5396e9368cd934e7aa9c28e1f2a84d11f40f7891d3adfeb05cded2ce760
zeaa8c82230c8d7c1af2f225f72f18fdebcd001929f5dd7743482dfef5aaeb0fe4c96da584fc0d0
z43e3ef836b2648bd2e70cb9b19ad2c61985c31c2c5f5f869f5199854326f39593074d095f4d8ce
z9207d9ca0d9ef4441629fb2ae730ab0b807993d4946bd5ba62fcd4a5396b0771a8bbab57c06ad9
z6c572f005d0812ca722d4c0b39143c69a852822e16145ffba79c6101ddc6f598765d252f35c95c
zb34c0e74fb4723245a6eaee3e531e6fb1d99cbabd61270996a6e0c3fb9250e305b45a8957db14e
z6617a5a81f6702c49ddb06888f3983f79676318b67fe8e42468e16083fd4fe4e16bad509b65d70
z86da819de45bde07e45aff75cb6dc39dca7561b430f096a57fa3c679e9e4fbf10e444bcc959d13
zb9ec607ab4e1f2bc5e3035517d117b97a9f91785d1ffa80467e8e8988ff000011ecc821b7bc762
z5d6028265b297cb28bc1a684aa00f4c5918c79f0b7b49ea356b279f28e600f2ecd9c3516297b6e
zdcea51a43125b4161427537304b348e30e49a9f1c5488c2cb1da7edf8382ef7d75e4b3018683f3
z0aee937bb2e4ba626f7c79cb1afc593e5537468fa342b242bce2bc33aa198af83a6d8f20901245
z4638a773bb3e6441bedec0b14e9ca208fee9a92e6d0c796322ea54fb7c97bd0273c78d4abcd35a
z8188f5a060154f1e186c6c2a8673fffb20d5ab805221f1388d538984d2289ad85f02fafea1a4e1
z4c23dd2ca488558d1e59feadeef0746289963bb71c324d863a8308735c682b9cb7efcacbbae037
z703f6e578ebf59a623a2624d17763a258c8b477b3cd482d4481242f74271e1db286d5bfe6cd62d
zb52bfc2fbdd311adc225387fe2516ddba3ed7435ee34a71e8e89c279f1be06241a3dfb2979c44e
z3eaa2abcec408360a99275bd5007bf38a77c9ea8ffca6837c98e1094d2c20511ab18549fac9328
zfcb1b105117a4ffb70f5ba395a7d637d99c566c94f2cc5623b1c68b504293682895d2cad020b47
z263572c7568b9f76fadb2c7556faa7a6f6a36003141405c5dc50466137d3c98a397240fd7d44bf
z1b60a75ed98bd2aaae5f9a8e18d4326eacfd14216a8be7bd9266afc7c5a2e6d5763e2c7aac9bde
z1440d6f5c70581012ecffe81c470f300330302028aff4a5ee6ffacf91bcbd978b98e13bd618538
z6c48787eae5535bbb2095ea9db3dc0badd8458be18cb20354cfcd3212ddf4c0b09c5b9fe3ef824
z1a5603429a3e2253ac658d2b54a039b1d0a76ead91ce6e8390315ffe9a931ffce92a8fee861715
z7855985d8ed543c7e7a2120ba7b7a310d6e2241e05b82bbd9028635c83680e15b6e230125e20ab
z1765b44746a77f880ecc77e58d9e8b81d658c415bbbd8c8de19673ffa1d241ce9b7506f313c96e
zc1a3b8f913021ae65fafbb7cfb763255a38729d4f51a2aa44118f29795f8b9c459647926dbe446
z7f235c016520bb819ba3ac0314596cb5f4281d5c87832bf7c387f790550ad82a29a6795eb3c223
z2a3959005a79fd24935e1991053fbece75ac967302140d6dff6a537172fcc01ae98c407cbd4862
z04097a2140b4058ca7cbcc2a9ef122c3217193fb71e40161ec420c25392c1909ca3ee4f77fb6fc
z1bdc5e6efce8f823bd2ea4ec54b1f9422ba1c1e29fcbba181a74f786143792038e1423ca1b0dc3
zecf16fff588143f86605e6213d35251f775c3c594a306a2624347570854728b43af2a9c3cdbce5
zd75f5fe7415bbaea2ccfb55ff370f1a6e6ecaa0d9ac42837cfc44f141c75cdddf7386ff4fb6ce2
z16a635b870567d565c2b9541db3ae2ab3d014d4129951f5e7c3167ec5153a6fb5c1009ce44f859
zd8f97a1a20a983aa4fb437910844d0577fce330786a70b648b2d97bf87784b1eb3799599495062
zc30782ea0834ae5fc7b00a24f7be765f5ce560c1cfd4dccc73abd809d270c52d323a15fea15dd8
z1f93fe1be16debfe26eb9196d40fc27cad1c05e85e56aab646aa179c15fb5a6b701c11378ded36
zec1e37cfeded48cf534386e4bc172b9ffbaf4c3da83491c055a7bd330ec1545dfea876112f506d
z19cd23c1aad7d59928f2b70149d7f3231bf57e5d402cf8bdc7b61a42c7af891e7339b476b1740d
z301467e28b04a4dbdc998000a92475d670332c878a5be4bf0cd6802a60516d3934075511f1f403
z4405f27bd982f433a994ae45afe0a5a398d5b031d41fda7b9cd0278796df24dbd813b9cef77b77
zd0cca469fdb6b5dea28ba0cd056b41e6a73ef89f3cf260ffadbf77b73bc942b7cca0abe22f26e2
z134d1cf5b31887473dfc55276421dfa2b1b32bef20669db15106b7d3d199778357eae31eae92e9
z20da319ed2e51c8df3feac5dce6ec058cbc2253316a205d235f827bbd1dd2bf7f6a0723dfb2e87
z8d4257e892e219b254f097f2f2beb6797c3fb9cd426181b2a5648e84003022ecf18b1d179f25c6
z395f134a4e3ceb508c682c23749daf87ee3321f6135beb97824c150f024bb755ce508d832963fe
z393bffc1d38843461f98d668a37d9c65f50e568b3fb450918e390dd2dac0636d2750eb7e6a2206
z36d648a8d22889217bfda7adfa9d081a2e4e41332a4f77098cf4bb6cca1e3cf9455b4356c1737e
z8ef38d61f0d924b19e5097c5aa53f465d2861db121c8eea48726b72d463057b6020346d8434b7e
z6f659ef1abe61d8cb76fa0566e2b6e67ad54d8a9dfdf85cc71506c72806a0969fd5426a9d73c8b
z7fba52a0bc4e3cca7d18a55a2d45a21db275b17a54a0c3eac76e00b59beae71650628f2578e415
z536ef907b1add28936d452b20a54cf5b818ccc6177872d12fbf4a84ac842f234cc82b5f3e9d91e
zb2ce0d05e5482e95cd46a6ab86b53274934824995ab376aae0c6cc49031e58b250207bfc26d05a
zd39acce0d77459ca3e81c164f054aee1c359df8c063816f7b70f0b7f7f75f86b4994e7ad33876e
zd1f5ca39997a6cac6cdd192d11cf1d6f39df660c8b9ad47a6d91790d7b5e6cde177232f097a17c
zd93a96731503b670935dc67ddfe6f2194c1274aaf30a691c1a6d3b1468212e9ca7623a9ebd03f9
z2ce3bcd35d0eebbac2abdb42238aa1057c8a65379deee5d66e64c6dafbcc8e358943036ce1e59e
z960a70a097779a5996db8e86fafc79e8a5e3c9ed1deff228eb2d03ffa8d0a7217d429556d3e658
z15e2949b92e87096b68c2e61f2890df10d865bbd1aff3563e59ef098bdee007f8ffa7f35ae9f32
zc2dcfebe7d124df3fd3b078946b6d60d8cfb330561c8f786957331b480585f73be4c60bab5b55d
z046878100c324c33dba66da3d79390154f1e5033075d4a2476bf65cc71d174877565d4db2cce83
zb068199fb81f7778428194a39b012a141ec996289dcb7a8f45d71a0ec86d1c0aab6c3aa91c6ac9
zacfddc41d4f9041d9923e1055bbe73e5fbdb9f2e1554f353aae919d72a4737788f5c663dc13729
z444e262c795ba6b08534ceee0446866c346f8362d0733cf3869032bae68ff8f9fe148b9eae69af
z6ca431ef62ad8466c43df4944d77296842902e61d916ae6e156a68ac4b816d18c9f787facf7cb8
zc615e0ac06df334b3aa78f48815a29daead281dd90efc2bf538d42e9e5c752f5f387cbb9cf32a0
z6f2f22f9a98622b07d960311c07882d6d84c88e983a2c3c602bd33d97b80513da3520c83beb5c7
z9b131473d90c7a83875d403635144d5e7b7495a73e8816aff450b3667c6d929ad5ce24199d825b
z50aa0ed66fa97b0d7e3fc5437f9da6ef51c65170812827518b7fbad49f014cffce04783ff19684
z3828fb6cf28a8a548f0c9d1f4f23d3a51d044f75abd53231322f3e62d2b42f67cec32cd04e3101
zec0186e520809e339060eab9d29f0f981e54ff2f710160814b4152a0415e31b1aa5761cbfda70b
z449bb6f570277e490821c952c9f9365d0bfb050ca77a5f6a662a61a75de371d1371380f8d6d7ad
z1312f22b52a4c54aee990b331b7ce34c096dd7e85765c1d75f1b24449291191e3b85642b3d2528
zc8a0dbb28edb3ae7da36073779c6062bb002c5a7165daff6df3e90adfa626e8fb1f3188e449dc7
za6ec3b5ea9a3b2f0076305802271751126b2b2858f9d20673fbc9c2d9b8e530d4bac44fa3dc3cb
zf53ea0b5c2702d6ab4a26c75e088f74095aedfc9ff2740b45fedc3e30d22b0b59d22531b0e26a8
z207a6579eac340a23c7bbbe1ab32dda0ecbd12876c51164745265a37ed07ca1b2cd960ddbc5197
ze18393c63a2ba1d125546a6c564245710d7cdd05c8c5173dbebdde8ba51cbb2b6514ec446ea9a5
zc4a82f6990a4c94f882914c636e8edae34219d39a4f28a0fa5eff4f1b2c1d120eedb251eb654bb
za45b425fda1d602814bdaea6bcf37ac792ac403a17a995cdb4416cf8de1a44164adba7605bb398
z416202f246387b14ef39f125f9317cdf2ad9c80ec057763cf30babc072636be5b4eb80328f6cc0
z269a341991139758fdbf0a664590431bde3e8cc829c5d7ecfea91e62d206eca2b8a9041e4b1227
z4f2f7be37480dc41d2305116cb362be206b6018eb17985362bc2e841442f2649857374fd3434b4
z16dcd66c53307b3c332909c286a92c9799bb59efeb601ff271a063b5e7701c84a3568766d5e946
z9079019b4fc482d64246e32b977a9696b61d7210a6ad6b7e8e789494301ec250395f8f8117de4c
z77f39e8031ca1ad88c937558611eb04e5fa1ff302f6b319c251b41dd84e771c020fc0e860f8553
z792e4ac9d770ec0fe1a726b567787a128beebe0a88804d9d9efd730274e7e131d3b795538a9c27
z2927d7462a2345b5a4f098b6591bf5d1f34087050c79586292a9337a4819ed412acf831bb3fb05
z1a2c3d43495dc944c4aaa85caff6cb2b63db078935896d6b3a524f8422b7c3e78c6c75c8c90aad
za0a6b374129908430901ee0f796c0ee69241e5ac228b1faeb42a86c54a23876cfb2725bb07c098
z54c5ad9b0289b4722cbff5b3498d2b2584eef04bfd33b62a2c1a9f88343affdf5d7276463ccf15
z3b7e65e3acc4fd8a00e10fa957618ee32077537a7496da090d4a98143f03f08d8e6508d58cad54
z93139f2c547f6e4fa96c4cfd0642f89fade71367885b28e359770c15aef27b5bcf19c705b797e8
z55032e6d7f6677f3f5614e3983478ce841e3c620720a35c91355e079f86a96bba13983d01ed79d
zcac5d23c5856a47838f5bc2dd714cd8d3fe33ff2c1e7ca82fadb9478bf489b33a1a2f875431b06
z88d1f0bac490af2d99b22bbffe4299f1d460644e8afa945ec043228dc3fcbf09dd9a64ab65ebb3
zba8192724bb0dbd88fc002c087be2812d2c7b2a120e94fa3f1ea9e4f4b451031cf9f2db6d60b44
z74debb3d6e2f6d05706a253857a86cffa8dffb8f3696a672908f884993ec69f67ea7702d0ce248
z64272abf027decf0943d68c6494ecafa57dc7589fe3a5d4d77fc70d0d0d71ec2f125fb01c067a1
z82ff60b60eb9ee1af612c9b738860e7789c0c67996c3b78cb7ce42e389f90b1260907fe7728661
z2b9b718f64f8713c6d6514edac5d5abacea50775e56f2f57a4a6f476acd306c470374a96efef66
zd0186ecb5401e7e2995a425061e19b18b260299a13d7a6d120bf8ac0621c721c4e05df3ad6c3fc
z1e796b4afb8edd34252a664ce4f70afa718c831a596a3b49e13ab9133a79c0daf3b0d9c99039d8
zbef2737df75f5f99705205a7367a4664c1a40cef33a8feedd8e29302ffa34aaffda74a49c5ea8b
za49ca2c42a1de1a0be39cc1e78a61a92674cad5227454d2bf254008822c6a4bd5490c9f286bcb7
z7e3e6f688c39302f4211b8f726c8672fa350d9537b289e86ffa813bf4591d342c2d2dfadcf0c21
zf7e0972f7e61a9b1e0d889d4e287fb57891721719f39569ed5cea2f57fd5952a0cee1a2e15d2cd
z0427df04b0cf75c3b48148ffd4daf4172b61e73eb8e80f4927ca344e737a8d32de84ed92d042ef
za0938c218e452342ec8025187cce57b8a1d626e662539e2c15e16a2d245e46946dcd1a3f14b8c0
zb007d3a48a1a50ce4a7c4533d553f03d9acec7986b1ba6f0d00a13be8a410525977573f05c672a
zd67a18b8f72de994dc29a8f7c7dff607da5fde3cb8b0ae45d0edc567e894de9acb6f63f3d2d11f
zbcd0a15507fdafce7131416d26a42f4fa9c9698b5532376546d04689239fdacc6c1b780f73c41a
za822e2134e66be25b775bcaab47f5ffdce62245de1e06b141e090dbad1c6e867c7c53ae1e79915
zdee8b57e2fcb368b2d44f3b9f88d0277d6e2336a308e0ca0a111ece1a9de1cedf7e5d6d9e4839c
z7d56e825381f5d81bf11f57098a4f36f157438403d97216c2269f2558197a09a63fc28a6a84fc6
zba8fa4422dabdb2192176133a261f753bfbba119c71a0ef2c6f6aa6ceb74de2dacb1f8c7c5cf5a
z5675229bf226c0abef18e3fcb31f882955c03980cbaaaaac86a98b0064394c309b416ada50bf71
z22b0708f9d830916ce874bb488dc8cf9f8d038a0d3878dc06bef199eae7de049253e928dd7dcce
zab9331136b41cd0212afa2d8e3142bf7bd3d87e821fcc748bd7de6a3a86bfd8bd3e8a0cdca9e24
z2deefaad0c288cbbbdfaa4a839761468719d913e7b3d4bff28938f194ebeadc4664f5fc87d9c77
zb76c965778990f59fdccbe2a608a899abad245fe575955f4a8a809be70dd6e6e2d0f36aa0e94ab
zbec952298922a19a0757c99fe14154812c387b5d2c140593a3747fc7774305b23d8369d72aa57f
z1b9a4ff62b09cf13c604349b3af715a0beab332188f1195a725e1f9a6c1aa8b87d73548be93341
zf3824885552ca1ce6d3c95bf5267d7d0cef976a9ceb9132b9168b1b13e158ea075f72b27f1895e
zd2cd89250b35d284c9094d1d95649fa3f8e43bc300375ba153a60e9c8596d256f0a3e09e324eb0
z13aa81469a29ebfc7c281ceb3e4b392df6072b73dccfe62990aac6f83661e849fe2c0ec34f9c6d
ze7be8545255e3ca1d5a07f0eee7e7a0baa8a0ad1135bde22851c5a12cbf5d0a2212ea929e3a7ac
z875dcc172661ec094313b517a1f8a6ddead00ee34f89704257d4daf945e23d4f3bb1a25a27a42b
z08ed0cb7ecc68d4b2dd79a44c67f5518a09980bd584e16c114fb271dfccea43d54c00b23f7829c
z910b2e560ba3c75e7be213686f78e134720296cdec8513430686d509bbdbffc704cadeb7837df5
z3008e153b5f790f96158b5aeef08ed6804efce5728baafc9ea869b85a45d967ebfed92e55ef958
za6126e4ba45d743b65fb25f4ba2730c6138bf3121556e9bf4d4105f9110b1c1d5af3ce88ed1138
z8a24ef0908fa3c30df6af31ea6c9d2983fae4d0d01be4a13383cbe9f173ec837b46baea516e299
zdc082eab2e875c09cecb7c5eb2f6458e3d4a8b7aa170fceb6fc4a6b0a483d6203eed7193ed8af7
za8ecdcadffa0f9e365666d6ab27e50c29fa24d704c1ca6405d84ed7e1162f18512808ec98e29b3
ze4d98663801e291fdfd55c8b0125d0d752344c36141b47eab9c3731bc0c25a9c97efb3ddc88f3b
zaeb66b34f633008ee2321330f8efec0773308c4ee91277169dbfd1db5d68abd29c91d555e7f600
z3492e962adae0b102bac09e7603cf35258141b2c1cb326ca61bd89282de9573d3e5cf6f8c0c8d8
z4638b13f4e98cd1cff58e252523f799653248b3c1c5a1981ce4940ce9158f6a8b28437bbffa5b8
z8119eeaca5144a0ba7a560dbddaccf222ec4d25f35fb2a14bc694befbe0ffc088302f797b443ad
z7bb4f92a2250d1b2a37acb3b9ccf00d081935b5cd5922e7088e9a02dfa180822e5107d99cc4253
zfc647e5a4a48f6c22f786d94be2fddabd1e802347bac4ffe2217bf0ead81a40af61529e05f77bb
z766bca187fa6e158932e5aab33a3ec401e308a0e986b91ac06a7cc42a1cacedb0c5cac38a4bad3
z793b269efc13c61eb9ed06d91407c6677ca474861698ec5ba165a251d6f321fbe466ce84cf9632
z2d208cb9a6f4718fb96ca3fe31fadc4e3ed78414a2854d09a751fb02bd459a882a914e8f460dab
zd549224c56752b4dbc13d898ba5f15976ebd7a9820df6fc6e4ed4e986893d17707336baf53af74
z47117570f29faa27884081b51d95543cfb55a4c61bcdeaa6b941ae1217095f4bb0e41673886ef1
z8ed7bbab2fda6a2f796d270caaf7a863548a11265eff72c92aa17890a784a3834a56e403a74e0d
z44dccd90bf544d7a8856dd376eaca1232d54cd6d1b60d80485c47ad1f43207e0e778381627200a
z83352b424e3fe148c588f67b70dcaec711a0f4fccb67f828138fd7175f6ca079023f0ef4ab8133
za3135613df7f0eb8bd86a117f43bbbd6e9abb211faa594a4b3070a5d1fb6e3f38b398d961761c5
z8f56af073e6472060dafc9353969cef5cb95419c794de055d01c93351c9789f715d270707e4cd5
ze0d0777f826b733f3baa7291902a684d17c3e98a0541b13d651b1fe699400d3a4c994cef8690db
ze36fb505fa07102335a8eaed10f64e32c39939c6a7ff7e782399b51b558e3737f8556e0a953387
zed4680c28d57f8af070e44545b6a3fcfe35caa6916bec9334d40a56b6a85e88858373cee614238
z9316dc835874446bdafa5eea08ae4d21a12fb348684833a3657838fe3cc8ddf0621c59d44d3e25
z8b8127d6da46eb24fd38b995e8eba00ea580567e22049ebcab547c0d8edcc8ac61b2f4df3164d0
z0bdc84a92c4ff1ad222757c3a1dda0d6dce6e373b670fd63df8decdc53b1c68795aedc80e8b977
zdd736fe304475a5463ed6d1173322f34d07271cef748a1e794087cb4c3f1d1c29bd6053694bafa
z0a6bf7fe3b6f8b0a671582644dfd387e10e2fa3d276e361677c0c6709bd6b0df563d84926e0c4b
z3be6f6378959ff419bfae400c0637aa981547cd1f5bd3a2d0bd79ef78ec623f08f843e683b69ab
z30979052d58fe928255743013cea7a3f1db8e474781d8af15b5376d5fb457221ce92a2111e9226
zfa236037b6b91bd4007e29e0a76e225743d49cf6efbf61c32440280900c0d91c3782a0d9b63cd3
z415793acb71ccee1766b42d802feffa896d39e5bc00af4fc9b489a180c3dc99942244dbde1061f
z2142da22823cd1542640e0d6dee718132005357ae9b979ea8233e524c2e2c4c499d5d27fae39f1
z4059ed5f1fe9f0cb0eea058d6ac15ca4a252dedb6702ad1e7756e903ad31fe7079bcdb4cd80849
z19714c1f7271eaa92afd0d24aa083bff178673ca9473f789785ab464c4019f060f8439dc73e160
z66760e5f07cdde0ebb2ad6244abba4eee4580c9158fcf4c0ac270ae236f74c7c757e28ac580401
z1d2845969fd2cc9babd3aad3beff3caf5adb51542bae70fae28ab293bc7d8056d88019296a2f1c
z5262c9724943a39a3c807a57d77c43678fb38f03106bb249e596dbc26313e7cc631e0b2bf82080
z5191509ea16368d285076cf0a608a7f1c22a51dd0c0116856a2efe93315d42a326322f68d01107
z943e659106bd451d7374b75053c1dec8fc95251352f3412e8388e527889886e9ce8e25ffb690a6
z9c4637dc6da65befcf437dc846bc3df39d79b131e443820446effb9c6fa8f19112173e79442b57
za1632ddb9c510a2ddc0a1b0a9a2d8d6dde400b4d9584c3080340983260e1d3d50bdffff5984de8
z2e6d295d71ec7c09b392cbd1724fa222546090d0dee1c19ee38df5d290c7ce5bedf6b6091044ba
z26b0251c41832a16f342adc86345a6cb087ecf9417adfc44198960a6a27fa67c67c6e6afb8d078
z73357ab22e17c63083bf794413e3c02694dbf43f2b5c03f825c206293d2555b284028538e77d12
z0bcd6e79471b0536cac6654693d93e5aed35aca3eb575b4771096ef1516ae23ff96ceb5cd51112
z73d959e4e4e51f7449cbc32424c6b3cee586bfb411a97a4fd42a06d863e65ce7288bb45b3398b3
zaece20c5e308c5a8248cf79196ecbf8c2e4afa96a8284ec977b80a31962298747758ec7a78ea73
z377c181d5a61f83539c08f228011c517b32a0cdddac3ee3295ab56173f0e6a261d57a21930dd84
zdb51ffbee57fe6c0c33c672e5898a1b6ea52eb4737af62833c4066b6473dd1ab318d7643ad2b01
z653232406bf6c1ddc856495660013ead83b3af4b7c07b39b3fa2fed52ba5dc55e6549aca567bec
z08f486ffdcea924b4c39066faff1e2fb86db96b556125b67ef73718cc76919127e644580c78f12
z6a99b2dc180aadb71230e7a9880aaf1bf621bafb140adc6da627776fe561568961ffefa257068a
z98e6150a343c674f5116f0f09672c8f3a9d61f4cf4005a8b630e1fe1203fdf0ce70e1864f237fb
z793f01a34236e084907ed48cd4b54b70dc095a7bcc22263f7a6b1dd9f5b0c570e1fb0dcf5cec98
z7925beed072da716026ce05055ed8814ca4d5db43ded1d6c1f9fe6d3239683aa9dadb95a73f39f
z0b793bb849996e4bdd657c614092aa364f3f4d56e7cfe8f3e0a3844b76c61885b269e33bffd45d
z04d035c91a426f0c0896cb1eda67d39356ab35335fea555342010ae76a7b0c646d79129cf424ea
z20d67008385debb8a68165f16bd29f9fbf5c0431af8779ae7bd3e73918bae234c65a0fdd79f9bb
zcaf52ca74ba03d021b7f968fbe85028760815a44abec8729f77a30ec64dcfecb497b361d239fbe
zd035b3bb282dcf1396cd94e27e8a56943184fb6ffaaf8fb81722e7533b42e564e7186ee4429bc0
za386532aba2c7c3c57810c48b0aa18bb7efb6ea2a3aa496632dffa0543921b3a21669544960330
z861e52ff405579129b4418aac008a9fd287cc090af123fa33785e7b3aaf1633d972b410124bd98
z86299e5bf5af83a72592a1b97dc20d0ffb5a0fdfb7a32d8e47394345bf1b4459af5095f6e0ef76
z9df1a0533adbc53af1b3b16c0f914a011d3436c3015d76e0c2b492312b2a6271411249aa388459
z1f4c42654153dc371573bedf22154711ef5756434724d8bfc3b451e22c68697972de02bc93aa3d
ze85cde989889aeddb4cecb720f83375afd8066c63fcdf7b0dfcda6beb37e42fbe17a4f38957552
z129fda9696fa1c5d266c555cb6cd257d2ad459afd76edd3ee5e628c2e69571167ba6bed0c66cce
z7c89e84566115d7f4796898c36aa7f17215f59c5f67507b2e76923d1878a258a4838f49925d1c4
z66a064a16047bb70b171dcee11e5014970fcfb5a4f2611bbbfb07cebe5191aacc9219b8a63b8b2
zc82a094521e711abf29a335a774649629af2022663048a9446485ab27350ea323780a56102d474
za3cc6389d1bffbd1033b1f034513b1f99504b71e9bcadbc349729baf24d4ff899b8385126bc1cf
zf845c6cdaa18f5aa69d2d05192d012fe97aafdc0c13563f28c57f3367353402b4823840f400d6e
zdde6f07784d0e378234433e650479f6ed8e877a7f8b928e0bb8d6652367c7094926bdde56bf527
z46ee2cf12b4f0eeff1387c69ba7727dbd235e4473a98beff36ec4e69b9e87a15a0d67c1284e746
zd56cf8ff97d82a9935f54c6db9169223ea08c45cb6a94dcba39f94dc52c7bae79a1c7d3337a32d
zdb83cbcbe1d78d31e48f1d36c0cd0cc4a2946162af4db8fea921d1da514f75c1952d3f2cedea24
zb1734d2f0938968053d25e9a4efabf6982d4246833f0af541cf84e564530fe500c84ba4b4e89f7
z58e21bab18f186bc2674e3140ea795c86fd14f0f31c85bbc81ce4adff40876c277c1164c576a9e
z91a2b98e7a32492f65bb29c4db12f92e2ac4157509381a6f758e976953ae35d7bf413447dd7cd8
za65b30770e9f4f5f34a3f443b6286b014a8c28b9455eac4cc108638f716cc64762986c6e429e17
z2c066bc7f7f4fd657e889ca2104e9075ef101a4f806cc9d9c77415ed0dd3d4d0962d42e0e7f743
z84fcd4ec1da841110286d410f5363f9b0b9e128016b665888cba685bd55a06cdd8a8f451bf8ff3
z4e4109d0540ed69a0efec16be130029031c36d57b13efc09b4b760eb7af78f39a2314e5b185ddf
ze15f1a32e4644fca222a89435e6c81f0f9368c2e5a6004b78d76b2d42338739a64d4790e371d9c
zdf3fd97c594925c938f664a0b3b7cdd91fd6c3b90e24b7f79ef738fd84c4cda9db92f5c5c11b84
z1513e552219a9795a1f27701466a95557629f2082989e6c4afda45e258acf9d294feca92d906d8
z6dcfcec28bf96acd188c6d89ce0c710d5987ac3e733e836384350c2d16effd70559718bbe51ab4
z42a9b40e3795b4f7d8df1d3d438c65839d36cbac614b2e58cd351726d7687a6e83ab9d56537a9a
zd950f95c1f0bf68f23f46bd7f449e9550102b739be0d61f49a4d26201f0e7bb10dd0614be63579
z835942c195bd5801f9db1a3944e0e7fc4d1abcd8de6d2f110e26049d1a202988746e6ed0e8e264
za07b8f1fae84ed1611c963be8e9ecc26057e22afdbdba3d8e761d69f046e79ca7bdb9a9fb3967f
z9a655d3d029ebce64b067afe17a11c393f672e441217d9d07fe6080dc70057a2ffea7af8a4a95d
z37b5bc50c24989b4c0c3e58c1be6d76bf043cfd72a4eb126a70b5c191b9dc1a1d2c61c3c2ff194
z8ab934ba630c8c66e79509e7ba134de7199a3a58e2c8b19c8b5846f6fe04d94c90f862c34bb0aa
z768edf82582e1c1b5cfb9320c07372e6666972874926b52a8f1ad0d27da3fb3ab6cd78f863da37
z4c438454c93271cb892b2f10fe3828099f4640a4b59da429032590a85fa000004a4eac0a1ace59
z0fa7aba568a8b5d770dfd66fa3410bd9090468f14a817b7e7c1817067c11dcc55616a540c455dd
z05ffed37646a08663a9d4e6ba92426cd67f6109b9ec2169c10049e5931a49019a0e1a72a38ae1d
z3f992009e7516807af770ef35d944b66dfdd947a7ffef48f09419c930d628a2e4b40eaa171425f
zec820015265a3634823077671034d4af934f68dbfc7ca26c31cee48d407ec3d1b8354e43bf593f
zc3b71dd833ef207add9f297503db290c9049d19c4c1b943489b8b45e763550ae3215fc50e3af3e
z9dcb42cbdaf2ae1542895222dad8473cdc226180549b41de7a317a51ede32f21e564b6fc4568ea
zec1fde5bce3d257e497f91a81546e4eeca3081a14bf8742a7877423314fb748ed6ea8badc325ce
z4fa0e3f1ec8a03f688960bb4f69f0b2ff8a6e3bbdaa79f6e91a464f4605459c6df5ab7bac5b492
zef28939ca49ae8cf9ae1e08bfa04f254afba106d424fa00c7013d5208b9697f77ca1d0baa92d63
zb0ee8ff074640817f5961870b0d5ebb8860665bd5f0e92e48a85e76a1853b1a12bd7d9e6fe8678
zb5a65a8fac019374e531ca746f52f658c3c8e19f786bfa399af4a97c643123ad1f9e8582949663
z8ba99a720578f3ebb33c3be76a05179f9250e6526a8e2d824c10d3f8423360c06e63bc51fb9749
zda0c0fb8e7c297df705eaa450597ab870ff7a94ad17fec87574ba4a5e3fe50f10f8965580f6e4b
z23d1c4cce073235bb2709b09c895e28dd26db283e75b08b47df76209921a5ddc0c41e156de6e54
zbd2aa6917fe76caf8e5e74c2b8894e1c7c2e80d6634921060137cabf248395be85e91e81293fe7
z064c5277551e23e2f1f946dbaca345c2fdf70e46b3d95faefbe5908f14f30013e8447f25a73586
z2d3a5c433c68ab0341af0a8f20111023bcff1d4e2ecdadda8e991186698c769d1adcdb6d40d3ad
zcce54de7c7fb9bf0554cc1c33c4bf14fca219ce159330a1699ee595a9a0f8d6d8dc81a67989126
z1bdf1bfbb23acf29ebfda32f9f8e7e49b037a659815d7a752f081a8687a53f3b69f910d41b2afa
za2b9b3ae8bbe1725b9439b09e079857c4b4867b8b5f4a6e5003797f1a13feabe2322946b3b4bbe
z66fe40fcdb34f502f74eb01dc4dcfd5df8f349fcbc4b4269b8daa73d58d84a49ee77a3d7917165
zd324d44432b156ed6178cb8ff6f9155dcf931853751862e8d29df6b38896dd0f9babab41de384b
zfd42a24f42cdba07a6ca73bf1a8004ac2064860040d5c61dada7739b7839ea7b45ba3b3c4c52e8
z845d5795da2321d75fc0edd9316a5e5b78a055f8b3d04e8097b1a86a67c08898dcea5321e5baf2
z5fc6adb79e601c1e41d531c06cf10a2848e40983dc24fab114ab38fac11718dd2d5b37d08707ee
ze1c775f729294de9de2cb45017a76a14586d1827bb75b803e8bc4758c755553e5eb7b44622acb2
z28853cae19c931edef8545848588f7db4766790b629da3430e14fdccfc004caaf1cf5815dec8d2
z6c2638b45d096c58cecf232711efeff1579a1d558ee42cff54df2681923e404cbdf47dfaedef78
z60f8d2af7f6e98b365af55a86d01fc1639844b5ab4b7da08e65928d74a7ac7995b19b8bd1c5082
za900f433aaeea4b434189e6b54916f6a510c634e4d40fc337bf0485356bfc0a41de6ac7551385b
z2360af1167ca48369e672bd17e6dd30a6f8624a3f133e1bb81f5913d5d9008fc0ace02ccd6ad68
zacde598e7e0c4e1b15f950ab566cff3b60e7470e88d86644b6d4c38dc9b8fd72d631f9b179043a
zc73da9ccf6c3b9192c72787d1fff4b6217c24d4897f2e594c7d0b29f00437243291cae6ea5caa7
zb5a532844bc00e29671f9a80c0fde63696e6f4b81b2d2c539a5ea7966ed90838c4cb6c96dca07b
z4f2d77e9d8331481496a8bfecad63209d223ce7eea1f050c867c5eaa95bb92c935b3424ae67051
ze7a1ee88a1b27b99974436c11f1a41f3ecc4c68e1224a8672a046926d48b2e147426b0b425d9ef
zd38c0538d226992c44c7e147216e49fb9d9eb13629ecf4dc02a248d8b9fb0eec9a8887c2c3f8d0
z330c8b354765faffd688c55ec596bbd851f238317defd8dbd138ba9c98ae374c0c8ddd5869e4bf
z5d77633d7307f55d6ae7dce42f19350ecb3b21e53d1eabfd138735421bc5aba5395be2db5766ec
z1d903664319b27eddde60b78c79f17d5ab0704460eb975c671e041c7c86d5f6faf4828fd3a85a0
z2b10d97287ff3b9580c8e36885599ab4d021b91e62a82a18ead978a21fd25de2d74bce5fd1a98f
z7730dbdb4e6a38f8a049c7d0ed2ebea4e354488104f345b58d18cec3ef9c01ac27380470e47d0c
z0cf1695c1c724ab2eb6c155263902dfb926b41f393be2bf5958adcf1a4e52cf886175974c07e7f
zde4ead2c31c1c46b0f0b8d23b21243439815bbc9e8bec0ee5592d2f2d3aa5326048ba185735b2e
zded586a824752878e0df3e2e4ad2005138e5784feebf90ca99bb86b8fee648bc3f3f50dd07d69a
z75906441ab9e0f8017ce82955ba8e42a8ec2fd556f03810321fe614dceea08bd51e864810752e9
z66877367f543e6bd6b6cbbe10f2a865d30e7f8ec64e2927b5b23b5401aab354219cc931d307457
z3b19532e9f71afd0569a683c9c3c439e665d99545803aab5c992f50782f68cedb9b39ebef8f015
zb4c854afc6d567b4e407f3ae3358a58cf5f602a0ffdbb842e5d5a8c6efb0263b7c3a133a417e94
zfe2294c9b599eae1aa11a86fb18ecf6c305dfd1177dac5c6354a24eacdc231b1ca5d8e1c14d7c3
zc0b39d294cc53b91ed7daf8b976c0aed681b870889aecbc191d353fa87253a10edf06ba99040d6
z8b8e484da244d5098459c8af1e0189fc44ad66a539e8a0d72d5aa48ac838a48168ab4a9cdd5a3a
z05bb332a38a1d28bb387abca5f2b6b6267df5dd59d5661666513108645e36d54a33ae39b9a8d85
zd256c143c31bd16103edd8046be0e5b0342ff41e11165b6d0927d6b14b9913c19163e4c3e5b0ef
z9c8c87c0966f628a60d06aa43e85e245b9cb32c2b48a1674666459bb1fa81285a3afd36372fee7
zccae96ca0f31089e3c29abb7c8aa1e97893f0469193c12fb89331762f613015ac4db0ce2c2c393
z56402bdbd91a553c888d76ba705f7659b9964cb67b32e209786c619a8f619c11e0b5fd49bb353f
z25f9f9859374c12eee4a51e531f3bfd492203c61b54b7574fe058b7c60e6f1e11684de5e429aec
z2d535565d4bbeaea454370a331a5b11d5fc168f1782edd02b0a032cdbe6ea06672742710ed30f5
z040051ba50c0898fc4258b3db9e522a210feb16f41d18b72f88b4789725f65c7792f6af04e17e7
z31928179cbee59faa6c3c223e30f76754ad0a95f827732e9da2ba9b4ebbfd010bc27b5e5007532
z05e3e9b4838400a24ada7214baf0dff5ee4ff6439ca3f3e46bff6fbf51ee577653ba3f6e611884
zf3fea8c64e57cc0e1f882b580805984ba20bbd3858e5d742b0ea0ecad470f4c476cec64beeadbb
z0865459fd08ba973fca97fda0541d6fb97ef35c85829353490245aaeefe9645c96306028db5205
zc54d4e8dc3f7b00cd15746dab63511b6f886ff3a9f5ead76a6e82153df5f23b4fcd810b032e2e0
z13a970326ce67dbfeba6436a487998d2c41a392fe0db81d0857fdb9e1e7df6fe241cdf47a1294c
zb7088a1cbf57c7199f173dde3dc68fe64600ade3c583d73ff7b47b1779b157196a582696ce2418
z6f533637d3194e5cb85459d79a5b99d8f59b60f9a216b66079f45614929cf02528a22eb51b8d25
zac513d59944ef3fec9db08c4b31f8e842c883a199b3efe3ba1e396a11df31c39e3e279372868e2
z1173a3e618fb4d70a9fcbb782fea3ace6877b5f32fc0b93ef0c693f474d39327b927037582e5c7
z05c8b373e2567e297eb7a53019e1b9c58ce59e8fc19da943f984d4dfba42fe170baa73df5fe640
z2bf97a28e5b112180352eb498cbd98de0840776aedd11ec7682f51855628aec1733eee0734920d
z9727ff8280e6b9f0bbc8589edb962c7878c4e06f7b3e6929201afc5dd5bbf5225924057676d2ac
z7a4df9c875739c364f1d4e0f864f31f790918f6cf789a3908b92fc9e405e146b554281540e092c
z813084927a13c4f88e2a198f057006a73574e248d008c150f376c491482ef797b819233ec99692
zea39c2225d838390d8d2997e31674e9183fdf82283051fcd2155513f342478f861a98b6c1b76bd
z5cf1c4e1cf4b8b36120a2a9147b71a64a3d60611e8cc25e9688973191a2f47b22657e4bd66d981
z73dd9e448375391b71e4c7991e4e7da6fec2a9b71c7033ca67e47ef2cdeaef55d7ed3e5be8e83e
z8e01f7c2428bda111a3db231c9d1c46c19faa5dfcdc0aa98f1bbd1b9c981055ce2e42cb7567fca
zefcf14cac799618742632213b8583049f2f68ad511a1e406fbf8cd5f276dc140b4eef1d751837f
z0301f7bfaed8bd767dada1e17edc6fc444ff759d1decf62d965c4335cdbfd35b46eeb111bc1fcd
ze1974bc97b325f55e8426dd55c024352ff3a1d9e4c5cac1bfa74e3d119097fbf563203c70d28a2
zed2f49578a5bee4978d53257076af1223594b01debf87bc22b2b5083be4cc12ba21c4ee235aefd
z9af9d1dbb95b1a1da6f6c847969c5f3474359a5d8de0c55a7538887cc599c505328c5d339d92c9
z85792fa59027ed055a00cfc6bf7475523ec74142d4b90ab54d5ba15c20c410f895cfe9b4730011
zdb2633a00b98b65b244434f85281207e2e8a800cf5ed61b958d34653309476b636270c26b4a6b8
z9765da6faad0f91755ae4a8e663a8e436367bba3c18d5cbcfd8038f779c3d05fcd101b8f01fe76
za5b4ffdc66ddbb2094956d11431b090d140ecb49bf9c8cda6a79d838b35cbbe837db1f64561d69
zf2f841044b0f83bb424e21ad637bf00b70c0649ed59bd5605b9d691545a93f1d9731d71d8ce03e
z91523f866d91f3b0acd7b0baf8b464a8887de006bb086140af40e090cfcfde2f38fcb34ed73419
z8b9fab2f11c6683b03b977691ecaa5c6d1e6ebabf16038e6a72e8afdfaf3b44bfb3f52e0d12dfd
zd1121a500c926036a3e9a8a5664a2f90222fcfe92af935549d9534fc847059fa3a269a9fe28e84
zbe125043297ce3778d0c41bc6af2935f880abf1c7766434658d3bd1be0371c6e66748145753bc2
z07b23137d756fe890ff8400ad687e84e3b9339b5c0fc3b5c7f9b0258d0b7607e790780bbe5efd4
z6ce073eed09eb6e9a9cc25a87adab52ed70803fd4ad7fed06e2652bd6b3f3063a120ff27f89e11
z380db0ed1e277821cf7e1796a30abfaf86e976957b5416853fdd370a22abf1b79a05af4cf6328c
z37719d5627df3f832a750bc937cd119a604768631ebf8ffb3e2754b86991778c3655f663d955cf
z2f64e8b580373c8462520a1c3534d3aa11461d7d4a6cf0e7b470826142cb764f609573d9e77503
z623fa91c3442414271a7a5be12bd67024c04b92e3d2b1345c7a963f7f48d985ff449fa24c1d404
z55e6b29305971afb7b35d7fc5f0076cf0c55737138f24d1d58badb5e576d3d3cad3a95c902aace
z48ecf04f209b1d8fef78c295a7c808769a00e9d0233648908f1dba239bd59d1592065649a57319
z0bcde610beb64732d5996b6365c75f6bb5babf21a2f25afb53909f9aa04b55be61726198804287
zd64d7cbcf056faab97f0a53750c1eb9622488dec4a56301f64cf1b1cc10b14c2a657a34ed572cb
z2b06f50de73e2761ec293931078f62c918d5659ef07790aa90c221c1b4716da45eae0a6ac6b80c
zf1b020026ab8601d1bbf95bafaf70cd7def475599361870c1cec4dfabe7f200495399a871e851f
zf6c6997751d26aa8ebf4c8941f94068fa9c85878f17006fe0ece696ec52661e17a99c1eaf3aec0
zc39c7da4d27e2142840652159559c4019850ef72365a188fc0002e4bf8d144eb151de82bb726b3
z7956e79a5f3e45c274e54fded8949e6b6e4b4bf7226cfddf46ebcaf2b8e1914c3aee4a52c9adba
z1a646237abeefd1b3f7396a7a29282528cd6c951c6ffbd5a56f4c181199a501682e3ff443de0bd
z5a7e377f89e30e87873bcb51caa47e22747aafea5c7f95c5fdff8550a5260e6d7a29a15d2fe2ae
zcd0414dae302d6e4fe5900f7138072536412536b4d0047599b8edf91bc2bb129d44df352a50c0f
zdc4f7398fe92e3c586b22943bf2b57eea1089c0b8aca7552148512f5d0bff112dfde2ecbc8eab4
z13acc9b0f7bb230f6f9f8c5e3b38348090f547f3c27418fe77a77fd7a34ec7199bc44dd2ff8c08
zfefdde3832a4539054bcec1a20434e13a70e4cbb6ddfed1d68369531ac2cd6e91e3e38fa4ddd9f
za88baeb8a032ecd1a0d435b2f60345950290a196cfcd2c12d9a5bf3b61b3c48e39d32d0eb60c59
z74c9162f35685632d80a8d4657d74ef5081646c3c869652dd57fd4bef7f6faffcf83c5710f8ae6
z542e14296766d8157a737951e932f4b49ab50fee8c2db5bf0cc2b669ce0d3ad43ecf128aef6e3f
z2b39bd2b5a28211b8717734af204a66a4cc1aca898f424486c4baa8e94ada4a96bbb78a7ae931d
zaa7dadf58f5e5648f59796084210284d0e48a0c79af67b3a449f96be6b4c84c124b997e9be036b
zdef5d906ecfa601cae4fc79212262e0ba9f7acd6e87c97e117a404fbf0c332d30eb4978843e060
za5874f2d8932ee6e3a03c4906c687a393badc909f08a4cb1e386ad3e44312b1ef60b5601c5e41b
zae8af4a9aaf59274247f580f331f2cf3b54279f6b08621d6d45cf8354b94914168fb4951b851d5
zf356fa977f91c383cdb4af49fb97dafabd9f6a8057f40cea2686bdf20f7aa95e492fb020b99d72
z9157374f8bac55e263162bdbfe59bf71cb9091c7db5056bccc3ba9022221224bc7c8aa0c78a40a
z4a7ae05ac8768a3170632c272fb04386693d8b3bae1bf7b52759f3d02f45475a9d6a5101288c7b
zf75268072bbfe68086885ecff6eb54e886f02b9aee82991081851a9b86c0494d0d30e27de761a5
z0b9bc3a0e3c5c8558701453cadb6c20af2be458a99d54472a173bcd3483afa0930d69ea5d9caaa
zb5aaedf7ee0b03cfff497052d0c328d36f37bea5c8a577d8129f754401c951fe3a94ebcce9b396
z6c5e092469884965060956c68dbe44e34199772daea19526b762dfd160c277b43a030329ff784a
zda3a82faf8b58c385d240481e7d0a8929223881379b12e5a73cfd8183991caea3e7842db03c18d
zf382823bd8563b607686c11f35bc172492fd8b15fa0d3d91412d89f6a80aa1447084a7681dbeca
z8671cb54b30f5ceac7e5e62c1051844324f384ae9c5373c49bf9b4dc4a8f0ce2c255e89cff6e11
zca79066e31ad307ce916f3ac25d6c99713d4f429a303b65738f293d4c0e3c60c1a954afa93aaf5
z0c6348cc9ba4f24c5b6de037f7e2f2bf7ce4b374012a1368f0649dbf129fbc42f41a24a67151f6
zc8c28e3f7f875069099e5ed13562491741a5f2bb44c6132eb39a0d0c2e80d9ce668eabdd371b71
z73d427e1f2a43b89987b23e33128339917c4fe7076bf8a9a8e105785e96cd64b4190d08fef1f8c
zf9cafbc2441ea7e543f85fcd60fee4a228fffe7b364e966e0716eeaeffa0f4b0af2266faa4a028
z9c28184d8161904e0ab371126015474309abaf9966468e6654c8670665249f218e5a5d31e20ac3
zcaf1bb67d0fe7e6a495e86a12e0215977acb9252374b5942dfcd7b31d34afecf690623f4fbd352
z491d3d1481f18b463293b9cefa4eb3970abe29154dc6dfaa96243a2cde6b6503099857e57138e0
z0cc64c923fbb6898e2044a617f094f1c01a63522c2d6fc58204b7be22848d60df122d6b7be3e46
za9dbfa2a963b8df34eafab7570e706dc23c1c9dbcb6e3dbb9963d7ecab537ee7b429defd311327
zb3c7c630d2223f8ca6779eef5fe499063aa6bd5b71e5ce9e3cfc0d46cb8244ee992ec206231ef2
zccb1de358c758bd20c40545ea1bff4e4ec47895bb6385c9f7914c712cae7fe2e6747ed0be3f281
za160217f29f952450d4794948d87a32116f088399e984461f322d4b7cfb4fab1dd5933e925d3e7
zb1769a41748c7a32cf32e836d1e4d0e06b05a8a9411fcf4599bc5a0852d6298a3c0c8ce6dd57b1
z71a451c57399a7292927ca82d6dffdc17d395ca2a5d3d26e3959524f76638eaeb99fc8320d3178
z9c324d17f531cb2f56e3cb6740a80a41428c9feb59c33563189026849ff065617fcc3f8c865872
zba61d25c91599ce727c2cd24c8a724934aa1e7a9e14622b3e5ae8a4d46df3ca1e814b650e88549
z5b903be16e1d61a2a61c24fcfeadd6f8e1bb4f7f0306b23c5527bf0796db748addbfb9d06206fb
z8bed02bc0ac0fcbef5773a1829a0403ebbb7491ccbd2184ad837c0547ebf06e4da0456e8e4a0bb
z30e16faa6a58cd559466e759256c231f55d90964d6c9434c1bcbce612fb6da5259e70bc2caef5b
z578bf9106e370c0a4f540bea296d2e3cee08008142cd37115e26f89cbdbcca8bb531667679b190
z545dabd88a399d96400de7f19ce79e9ebcaf3b009fb9aa809b5901808cf3df1653ee48a1b18684
zd37d5fb8e4875143f4cb8b39dccbc59500c1c6681333afd9abe70b664d0264b4c12cf235bfb77b
zdc2a382af27976c77d5b83a5769315c2413b8ce1788a09556d98220499e9e045a3d025b33b9c0d
z9804472efc833bbcb4d9d0dac1ca86272a42cf6c0ba31131b63885e1c1817229d046e6c8913b44
zb8b3cb3239224e10cc5498c4cd69289a553673bdffebcde711b5c6014b3afd683518d12a6a0a12
z060d0d43e6f66bc7ad481722fa0be530ffb421a24e37449566167b4fc51a4ef76995cabc3321f3
z4e896c5d9146087ec8b0b7dcbdf889693805b0d43476b696bc2892116af391168c50a20694244c
z92364bd9c1deea46ece2509309b734c6d370d9da46c8e65ab65ffc94bf67c755f103c4244e60d4
z1f044cef6685b75941b8c3c03372d21a29a08a2eeccf59235fbff31fdb42e590b7d48c56fe7780
z13bdd0ab5e275d0fbcf8103417c0ac06ee34c7f836a6d2da531706d060a3ad48831be832eb7504
z2deac045b0e07f139682831bfe4906cc37ddc559c66e6ab059171f10fef8532c4e1879625f0517
z568347b24bbdcca676b0b0b9ee45f11c3e609e06ea052d979fea071339dc84066664e5537d530b
zf6200f6b4fce65b54ad90f1033d70252625d476c8ac733a4ca3329f065b0f9f78a9f1338d342d2
zb10c0c9895c74497a7652ded9033ef781a55d8f20e95de6041a7ac2926ece4655123c8ce58772e
zcd291b107ad72d561f470e06577e8aad7af7b7f2784eaf4be07fbc142dc128a9a11014c7ace7ae
zad7c7a8c421b7a23419d6ee2eef17a1709ba7d1c0ed456769bc0656efb1f708a2303cc5789d1e1
z22df11d89266843a93db696410586cb1e85ee9606369228a48f842bee5eb57e4c96edf6d002abb
z359f7742f514cb035c6280358de3564844d77bbb17b9b852c88b1d6fb49f69bbec34b8e5bbe11b
zc629141692b503be082bdc0691e2c3bc7f2b6225cca469685d2753c23854fcbf0a3054921828ae
z12558a86ab2e4603bbe6e3c60e88276cae7195b5ebe214495f73dd8640347fa5715cbf635db8e5
zc46d0ac49e955fdcdca0f24f9bf20a157765eb31d817ec13a5198876c64d2a47f676bf7c1c889c
zeeb668b185489c295aeb46f8230acfdc912f27b21f46b6c6e3f58a466d52cfa9bda939d2e54444
zd58850db752399a6d91ea688118a209f4cab411ea4355560b249a9531cfd5b1af191d1396a4cbb
za5734bb54b7f34d39636939038a742fc706e43aaa98ce3ceecc1d4bfecda2d1fb91e7eb53d36e3
zf21086558f9040d288c7afacca2547a8dba034741287dcb7003125657fa6482f66aea138a44f5b
z9bfd8892d2b88c597495878c3232d39f9dd848661aa4596242365181c23a4c0227bcb65a3308b3
zae1c9940b875fe0acca2b23640675d8c8b2e4d43f5766793f288ff48fb23cd5f6c60f3baacbc36
za848072a1def3c6b808f57061c9d50d4ea123bf9fa2261c8d0302046c8106c5e5fd1ce95e34a84
zc306e79f83e7c8fbdd6446d386201a8892d0d615cb97e97f70de06e9933b16995bab72aff96c2a
z229c18d42546f833bd252935dd2df1385f37b9dcee155a8c7c9d0f26a24f874bba03e132458f34
z9d12406c472113d499f18c0adedb17f0241dc1d32548c554bbc40cfa0342d037c81e2394950dad
z8edf1b8dad96ccc4807bcc330ba7fc49455af44fc5119b3671892f36869a3187b41a4ee080560a
z2e80beeb8f7b44303e57f962c26a96cae1749c753052c1eed8ce2ee5338eb25110ca05dd6fd649
z822b367de771361fe461f7cb6ef31204e9156aaf1ec5fb23d7c6dca89672da08c478c626823b73
zdac15323f857107cac0f61fb32971d4a3a45141e7da44702be01844197427629e344226f53fe7c
z769341810249420bdc669b470be8f5614aa049f254bdd97279faa6cda39f617ea1614f461346c3
zdaa2f4784ec8e394f7a793a385df718e2e89097e1edfd91daf26f0a02d73c1ee93fb4760d33ffb
z51ea7bfcb7874e2b187165963e5014736d947320fe0baec04913de0dabceee0d4e8cddeb55f6ee
z977f539d68f39db5bb21b88d6e9d24ca32341f6466bc30b9a03522bb547fcee3a8797600aecefb
z85af5c8907beaffcb5eb6e1bea8b3eee5105c8eba8acf15a8b74928fcad9cf404d36ecc2514cd2
ze40022f102e18b3fceb47c9771653444caf90314ff9218ff91c601d3ed8c5a84ef9f03ae66d27f
z7ce31c1760d6e16722f8d3abcb7adf021a8fa2034a8b6210c84e5cd4d31a409079c0a0d54b90f0
z9ae43b1285c5c0ad6628c563d04057f50550eb9a2fe68033d093f41c6b56f8d16c65fbe86e7c2d
z72776ba9d12d0801739074dee790f300bed84f0cb32e6a29bbcaae44291127b98e20bc7ca54052
z9851a152de5b6f19ea7708ceeaf5ef3f09e6c4dd3842cf6d48957988fbce640574f9f83029e562
z26fe12ff432b4ee6ca3e32179ffb5ab467149346ebec07e8741c9297e01ca4477536b0e4747f98
z552ff88e1f453cb88adf99f0d63f49689591c74911e834c9cb92e1acc06eaacad7fea2aeb47435
z0fb4e77b0b86c6534a8cea25a45641986dba6084fd466d18da044fa99c35fe88733c7694e26236
z366f15875b2ba95a7266e237ecfb44e5e59adc327dc6f30f699ff5b49fd46e4061bd1659bcf77b
z0e6052a28f44321647ff9927e97ba1603b8fa4a3fd35de99a6d43263932a8723323d9aa1ab2504
z7b88113b87474b036a946e87b0ec579251ddcf6ba213a7dd2dc3b4a4bb8a1bb490fe40d4ad5dfa
zfe328c75c9fda0ba776106afb623ccae4f632f449cac69902d869c54e7c0a8e8e24c0a6268c86f
z6f6a1ec6824281fd4ad7ab523c9c3961aa14e1bb598234a2ea4f366798db8f2be12f9081d216c7
ze6a0fc885f10111ef4c6cb64de82425a3da5b772f25f87ebd7b5ba93a6260099c6fa168b287640
z2128bf28e6ca25e38d2df4dcd37e073b1fac2c26c2fb934d291d008da3903c840ff6acbd1ad2d9
z801ac06300c0304841741fddd7a83b851b5fd57c7c3927187b191b2b07dbd4003da5e234cd143e
z3588dbea855f303541abc5f8c4edaa6006bdb13702714bd2177bff38043e64dd201b6a9c48ee3c
z2e175fa8901a01f74275320ea1190f8ebc58b6c2d915373740067cad756eec04a493414952bca5
z65989a728ce12e5b8efc01409ef24980e4e9ff7c968e90627d7c78ce67c748c1ef334d08514234
z17b09692735ce2f50067327ab9355a538a730e6bc5851bcf2f12ec5d7985cc918e1742906416cf
zff5d795fff98449583f891b97808c037f48c9527a95ea4eeb3082e0b3fff3724d6091a24e41634
z62b26daf5f73bf6829b5351db7910c197ef57b5b982e42300e129fa67d34ace092c7a9e49635a7
zb486617666852117bdacecb063efede13762cc7fdcfc15402eb43495e092542883114624583c56
z7d09316f03850294ba575288db3adafaa1af0c7153aa4553e2cd1709e0f96cf7e313b6a9eb7716
z610f045f4c891f6f64e3f245d2c66988fbfa7f98382d514bd25d451940bd5db87b2c8a3e1d8a19
zaf21b7d85a9fc095fcf46c1a7fab75046cde6d43ae70438f1c2031a570e7ae538e9249b050c0a9
z78a4b8bccedca1f2759f5f1e49d785dd47511390fe940f43811e97f03df086d346195d237dd533
zb8d23ef15f6e4de78efc00f11b5f3f7fd509a30505eabd3f71bffb2bac10de566d7dce8e29f5e5
z367aecf71049e173327e6b431f2e173fd3c47542aa0c29a9a131d0de91c90d222d4f2b65d10c05
z7edc3eb1957e2d287f8c7075b485838d251074f325259f63174a789757b95e2d21c25f296deec5
z66f63812f6206bc833919f912f8f7761e0256fbe0b1b0b4295e13510567495d672516681ca3424
z07f50e2f1692211335841501c72da1c9e649c8ba97c7ac11f7a80b6f062be63323ccc522a14501
z05663104ec5d2b5a7c2b378e87aa7279f6c883f33cb280f8eb94043602b25e67eacae8091bcf69
z111774ea0122c6d47876512bf635e4ceb6ceebe30f171ce177380f85586c3f44a3e63c4bcfb00b
zf672668db716af22a906850f8ce3adbe6249fbe43c1a32179b04becd09aed5cac3698d95932779
zee680940a88000b15270d43ccf9c33fb431fe1314d0adde6032ee324062738073e6049993aaf07
ze34fd7bfb6db7295dcc12b0d609110215138ac9bb75d55165bf1ba396dbc7931f8836503092a34
zd20c48af989cf2135ff0145016980ae1e0fd1bff44a2144ed9a5bee3cc09f095b8e3efa7b5cc83
z1148261ccf62493edd41c0dde9a2e0adb3332b2ea4e956032a452efccd337c2e802b44b5ef579d
zf3d5c122980a30051df32e456bbe761aef74976894d076c7e9fbc86253776a3c5aa4f27d31da9a
z2d82505ed68e0252ddaeabef62cfb2a89fb563d9a4997cbaee4b5f398e5fdd9710b860425fb52a
z83f2fd9563c4e64d04dc2bdb4efa7e934df50ac721c2c37b4628886c4eb120cb92470190588074
zc89afab24a4d5219e85694496275732c66233d1181ec082d2e6d2bbccadfea5315fe3627e34b84
z7ed0e47b0fbb7802c0f64fe6531d2274e73483fcab84cf48970c5d5a79d4062cca26813ebe4aee
zc9393be3bd857e3a47678b141095b13a13f2a02fab815f7445f4fc1badd4832cb383920533f2e9
ze72edf708c6acd25c2800ba2737c6b974ed31565419eb64972ac3d24a755d74ce17b5c7a13bc9e
z3f85244a3d4526404a4b591dcc5b15a78c413bbf14f741a9c307310b031c0c859a4f0e4a98cda9
z32a114ed26969d451177b238acc33b33aa74f638e88b1cfc6ec6936a8dd1566501653ac52bcb26
zd8013f571180542ba1fa4f726436fbc9b9829489032eeed2beccfa147135c42a46659b4d6590bd
z344c9a344fa29a4549306ced1b0336b77a50f0bf905e95074c87a968612242a594d7eeaacf7268
z074b82484af59c5bd5464a3c437c78a15dff8a6454c4c228abf69462dbaf7416070bbb973beca5
ze0e37f735af89b2ab86527fa873ddf714417a5a874cb6c8f3505fa2ad8dfe1670dff5a348ff800
z294baa052cf00ba0b426065887a79b806f77dadfc1188d46c5b7b2c4a31bd3f5906c2ddb2b36ec
z385c2516b3a785c7038d856ecbcc8e4cffd59f13d975694c53087c8c5ab7eabfb67040c650821d
ze02aa044b82b1c27670684c751a40cc984ff50e189f0471071007ca84a9a0d0aa3a45c33b46761
zc16ff600ed3a7d701bd0ea270789d86016bfe34d7de957ceec1ee897d66015183b905779ce6e63
z2026bcb22565ad714de1e1e7834b87e3038e3fbb6dd08740abbcc5e534e93ecbbe656c97572d41
z275efc821be4b67bb62c47980b5d5595e550878f80097f7f67a2f9bd5e2d0fee24fe71021cdf62
zab63ef0668d7625df9d8bfe09fd8ac8ab80d01f77c067b9b6d0fa620401be82a16fde11fca83a3
zfcfedb2eaac7001a42594eb2d55a845c37a585669bbd9fdd5fce170e1a248b3fda677d3fe2931e
z52a8021707549ee1fe20d8fe558faccb3c6271a533d0ff8ffd8513d57a92eabdf574c456a22513
ze5cd4545f70a4b8c070fae0391c627182accf774388be8e512668d4897792c7d5e18b3a892bd83
z5db4f0a3ba5e7a1e395ff0143f94df76b4c6063cbf302cde709a20fc482734c591617cdc3f83b9
zd5ca722e5d463168e999cff6e68553bca23863d5410da539c98c9bd65440c51352d0cb4b81752d
z07e38fab5707aa97977561864eb360fe64ff8c4f8c261a5c861171af1c446cff80c44f5fc1d83a
z62076c9347fce476afbb0f92137b037cfc5a6a5619ff1b976d3e106966b78fac83fcf8751b7322
z400d5d84f2f073bb4acb79ec9dd4af15af316750ffbd39697198e15c47a4482fe3fb3cd88e2a0d
z51285ef5a81e0d4bc0ec3b09de050568439b666a318ac107f56e4be8924b918c31c373eb82af0d
zb98249c4a07658773499265152ff3da95004da3ed80bdabb1a668166efb4efcdc91434a0b48f2e
z118eb5c20a07620dce95c4efafd17d63d50dd10d50816d185ebba72a807e4ea9c876b4aaaf0385
z2775377270d46b943b5e4b847b7d17568d3dcd7e624f247c620ee79d5fff1106e4985768f1b441
z16d3be0fd482727dbd1175f8ec0752ee182e020d5fc6fa2c226349eb8a9bccb6a3827a38256d38
zcf5b0409416507d07bce3ff4ec0f3c4104dee9696a1e58e2d2761a29d08cb6f0e9bcd2f015641c
z38438c027e8e813c502280da0fb2d4f1d64322e288f020c095e43ca7998e544e5a8916d4adb5c3
z2bd8f4bc43ee143f7b975570131cbaa4027a15595b7959fe7a07e72f142c5d0bcf42e057db2143
z9a639efebd766a5859faa1bf7339119200a7305ef49df16b844652224afb55e1d071d8837d0eca
z78655edaa5a663f24086eb4e6edb2b7fedc74d903583308d143f94d4d1ccebc0668ca94460c0c3
z8ba95a4eede786d437622cdb3a30f1414dee241e82762bce30ca2dc1a5b9507834e833c2c828b4
z9fb382a9458a492cf1e1ca7c8025d26a34f7dda4e28b9cacf5a9ddc8c4ac9dd6637bfa45bd5979
z79e44acc6c531d79de8e924954cd15ce0ff1d106585053b5dddb367601361ed48d3f0f6384be1e
zf07fe21f02dbd574ed1c5617ef148e0bfe7d4443dd685b326b54725c9329da1a7c604040bc32a8
zd345839005bdc0be37fd8983d4b1793a58a259d8521d355c0ab745b04679d9322c4c60f5c4b77e
ze200088c084386892945994631ca01ab3a5b45365994a3aa6f2e9a15226e6ef7a58790dba63349
zdd411baccf5ccbffa15af951618446bab1d0e93a16f1407aa9aec3188e8f4a1a45335e4622b6d7
zc22ad4fd2c56e172604574bb6cfb523bd39fd11bc9780c9d7f00a5e8ba88430806d202b1f77bec
z1317da9e9854fd6d1fa347b238e1a4f1b6fbff6227e302be3cc85571d80a74ba1dbdd4f23e02b6
zaebbb80329234227a9e3141476949cbc8748e3fb5bbc97c96e22b9cd15d63087f4a0386b032db6
z360dc5a1839f631cf416e92cf06d6f6cc794755c136647f637a6662270312f88118b638211c406
z33fd8f4425fe79489085f1ba9cf563b71e2d561e90a906add2f9eb368164a8b18a6b09f9c8489b
z20f9c28a97aff96df720064b0ba1a4dedaa8e05119713eb1a11238fa80c9546b04752a1f4612e5
zd925db3479e8b08cb777746d8cf31b2afcf61b1e1081b54472dee13721c923259d52a3a1fbc348
z533564d119af60075b6bf4ac48c289e6ccc8f1564c416e893fed36510ae7e24a709a6c7a20d8dc
z6bab8ca999d8e0849bc2f5268f8fb5caba569b0ff1fa7bdc8f4cbe50fd0987711da524d8599c5f
zb6ed2a5bd76320c96a7453c5826c31b0f8360ee5094156b3bb732ebeb73e84cb37c2d14535c854
z73fcff0cb6bc2e3cffdef3ecf41b54047c3b2946d9f0d98830da69da7dcdcce2a1534f905b93db
zf024b287155112ccbda092339d147339d80ef2a7924f3788449f28afdeb86841fd156287e5255f
z1406822b5e2ff5c8d050dde6eb603fcaf41705fa7921a5d35a5e3eb105c88aec07ad5f4d7788ff
z9a71e99eccf899ab549637e74d1b1d5189d5fb64c18264953c13fb6b3144d7928ea565b734743a
z8ae9088d623d3720bc5d6995bbf080010bea67e5a203ccebc8f3081253ae8902eb6df5fafeddda
z28d47d64952a6fbcfb313a5489dd3a7f44feea32a40772dddbbc9592eed53679d096451004528a
zcd6dd475d91c2d2b92bff0cdf6f74144586545802997b1273eb3ab46ea2705af1187804aca71b6
z01b6922413a3260c6de188c98b16b4b41b96a8bff2dfece8f7f29a03c5ffe64138dc7c5becf6d1
z157a062f32b397a62d8d92e565ad78f1400ac8b5f283c66ee6270442e96d349467285caf97649a
z36ff653de40b1f55af4e909db117c7baf555bbf44e10a819b43dae8f141862eb5b2119451d26e5
zf1deaedc2f4cf7fcb7806ee6817733c15740983074fe1c14bbf52f6470599809d21aa1fcec8ce4
zf52927e770a9113eb1ee5240274d200f2b3cd0c5e746e52307905018781e63b3106b2260ac988e
ze2838575a022295d1b73afbbb579ab628909d812ea95a6e202d6da44343b10150bafb21d17ffe2
z80f66f361ff961c57f26170932f4ee51ccf2ead8dd487d33f2262c58b561822aa6b097c0be2ca0
z763702d7ff289c5866258f9dcddf822be1393b5b17210a0470ce66f3deb00aed9be208aa8469d8
z6d18b971c5d1da800a09b0ce249b9ce7624d5a7253e74d7bf81c8bb9c9be4d00828805a2d7841d
z64ae00bd3bd82cd95b290cdd79fbd1b6ff6db3928d780d757bb4df8a467d7cab3b5156a2c87b40
z2a176288fb328f2a7fdc00b942b0212eb9d84108468b9bf49493d4753a7cca48c6f8d501897589
zfc62f7ac916d8453976f5e0f420608bb77648c5e6a471b2db28bf1d0e42c8decaf29d0f776df97
zacef3bc06f2ed96efb485e0edaf5969014aa2687693db2f9a1d3edf7ecdc149a34ae40531eff1f
z7f98af7a1e762360f2205e8fe35aee663aa1a27453dfeb99fae1301db0df552997c8f3372f7cfc
z58e87f3641c29fb23bcbf7c5352fa0abf233b372805cfa96f97ba5f8e3bbea7b19d64fc1fa6112
ze8e2f3b98d495befb51d84cb4f8d7414ceec378b6786ba5d7a0c5a5c19339b30fbf0a67f7aa2f2
zc8629d4004a10f8a310814756b1c2344e0a5d2b2cd59249f2f7c95ea016c01af98b1bfdda791b1
z78e7410c2b94f971afaf20ddeb0a65a412ba3c4f20cf14b72e2496e124aa2a2b7ba53e55951fc9
z649944b994579a164f73c0b1e5a537d3ee595e92eccb7fce0738ec5dda9cddd51987a162df08f0
z150e2972482527e800131fc7d66f0c48b4016d9a61b298531e5e98d218abd810a9cb378328791e
zec7c3a0085654bd4def5c8d8906d33593e95c38dc719d086f736b0a92bf76a890730c5c0ac11e4
z7f79f3bd83bec0f59414cd7b4de0544310f842b67afe58eacccbdb3045b95d356ad85d4fd9b1cf
z90fdbcf30809981e38decebff28d5c83bd29082a1898c1c455bc6837e1b8e472363a9828aea4e8
z9b4ae2f4c004bd24684afe82393bde2b6040138c52301fe372f06f7955cf524d9bf27e719e04c1
zaedf1c7abcb82961fa71adb2e0a95d6af9b963a3318edfb7c2850f29aa36e0faea6c6eda906e1c
zcf8978964826befb3676632f9bf1eadfd345e8ad5cc14972dbc472ca2376d91cd938c740db00d5
z73223c9f6b4e17ca08a4b3924740d9245b8a3a98924db5085db62d768a30424d107bba8e1df486
ze8002b3f022500586ed1396bff22cdc9ecd90e7d455fd8c53132a760f14180788675ddd5e612e1
z2cff53ab74608843a8d0e59e310c9bce5174c1aa0cc6711a8a078be9e86b29971fec240acacfb8
zf48062fbc2685b8af1400f1e37483d9221539b0bdaea7f6e4b185a241f2ee9af9cd121f21a4ba7
z2c3223792ee8e6ad77218991118852d5ce90ca74d9b7b57e630274eccbb9697f0f879bd68f2673
z02338b6519d35ece8a49d0bb3d326fcdd9351da3117e189dd068b105fb8d1b67d6f59bec73469b
zb53221722ce3490fa69e5b8743af689830127cf360519ea3bc0d1a5da7846d460bf640e65bbe25
zfe6f0b7362523aaa39c723ac026a9cddea9703060e0f4982cc2c61e8df7078abbbbcdb80feac3c
z007e2ef00e9493d2392d49676dc68dbdb79031c88ebcefc18eda9742e86364b802fae5148354a5
zc5304da4ad76f02ffad71f2666e48d365db797d16bbe2f1bd7d27f438de885baba161580a06773
zcdc0c961209354e41e72ce0ca45771c21244e139212aa32008e17959f84fd978c6d5b691ebf582
z91a1f5b1726674566691c9bfabc734ae45d25fb14e3d85ddbcdf9f217a3d04bbe17f30d8268601
za9e169cfa10597f0a2d266a9ace0eb5680c16662cb53880ea61a827177b091ed6b9acfcf384942
zee3082cefafd8d29f9a743874bd55aed378f02093662aa7098825119fdfb016a992a1cba36c97f
zec74bf5017ad6586cecffd3ccb1e4c835260a60f4096541b669d23fe2f30b88ce7b0467eafea1f
zd130a9d8b55603b00e1f0108e238dc308328ba6dd5632de59c32e3de73f21734a08961e5dfa32a
zec240fa4b89935a3e7d177f45abe55c22b77445e95840dd6cdfb3dde4906687a7dba6467bba074
za606eec36cc6b0ca4132e69320d2497901e1a2d804a11849fd9ca3d3ccd3fc600e5017426b4ad6
z740e480df047b5be348612b26255b8f3c9c4ed973f48917aa2a2f53514f194f1f54fcdd66fefb3
z3cba50aef56dbb2898483dd783f5238e5548f0d4af3178a4d96fc51e838efc4663e147caee7acd
z059971210c989eacbc818055de2c0dda476e7291da5f34cce3abfe7612ca063abe77fb11dd45a4
z2079fce992399dab01aed8b9a0e149f1a221c28ea12a0cb293fdebd2f16ae06cb2d97694512bc8
z7ab73291d3ac10828856988087d70d0a4b6fc70ddc094456786d02c2707585cc2fdb6a0f4c4357
z2a90e15f09259025e60ad6741154a652526dad27e6e9a833c9efcd3c74dbf3f86dcc51f6952e90
z69b1ba492d7b84ff060f6ed333c38e53bbe350ad3304c6ab0d4100d6c61bf1a698e08591a20444
z0365a2d3786275e3d26cd1113667d0cfedac38ec29a30e952be20bc42260c525d01c33e7764456
z20f92c692d8000555b8450d44a2b944da829b25a7e3dcf403c47600665b4adb00a4527105402c2
zcd7e59ffd1668bdc58008c9c182b99d4f0a76629de126ca3da2def308b6cd52068f023314412d5
zeff1387137da32b9b4ea80aefe27667718ea8281a176829b368eadbe6615a8e06c2366a67cffba
zd71fb678dfa1e8f607dc4fb5d9f20606d281055d33dc3fbff365b6e85a76d2d8c19286412acb5b
z07ba2368ccebacdc3f768743f7ff001a129b08f2a783ae7f5e6a12177d745aa687e69bac719972
z6cc65c6ac2468ad785f7e79e86a4fb2d4d59fb3a8c343d160e4d89628830ab6652ea09d9763d61
z7a525b44cfbe67f370dbd2988cab405c40ad329db2321f08e5bea0f66fbb54afab2715a7e1adac
zafe7658ff6a977513266b9cfee595de5990c1db3e3d4ae038f4914a6ad5c1cdb749a78f8e9ac3b
z33d98d68aa3ba3885f87252b392036645d780de7b466032a9f8a88b5381a472b1c33b2500be06b
ze54af957fe7038b1d68b9d67b4d6f566078844cc4b4fa7e2af8499f6483adea27e4de718727f6f
ze6d02d9bc2e23da4fcbd16f596d7f234d829180fb892b7952b828d31b1781f56e43243d1d6ffc5
z7b233ed8c32ffc947707a5ffe5a79bf26e80325b5e9d64ffd4ccc49689d1c01a17a39b54507de7
z190317c129a63b95d578ae42676d3e036a7cbf50cb70e4bc9ddde653214a04a691348e892fda41
zfb468c38227545de45c5c114b2fa97a768b4703229c1071d641ec33e1f2bfd68bcbe137b35dba3
z5a29132da88d204f82c6f586480bbb968bcd283b3a622ad7c315f286d34f1571ec5f94b06c403f
z3ce1fcdc550dc66106ea55fd2d284a2d2b6f78af3b4bf8e2fa276c49f05ba101f5cdec51c28bbe
z2fbb899270374c5815a1e6751bd2d7fe371f2e6a93dffee38319b451a1c222dac45e7eb82db947
zcf154cb3571754f44a5f6c6153c1f37a5e276c9dc93bc2c971692548e3c74a4179c7f39b5ad74f
zd22b9e04c38d7f27110872721e4e1f9e323f3ea1db85eee4b7c33d540f14554c2289a3c4d2e71c
zebeeef8ffc12e4a612dbf903c856d58899048306995543302f0e5487ab2bcad3cc4479d972234e
z59b9fba706de427b63e6b11403ed9f332652abcfad5c11bc0f4dd94ebc53b84d6d32835ec5d15d
zc8c9440cced9d17af2a7f943b6b54af7420af99687600050f0a822d74a0a225527941f64bc4fc9
z24d563119ba649423364784e5fd28522be1f1ae82819a59d0c96c7fe46a710fb7a711ac94bf0a9
z1d261821aa970851dcc9c11bb163c54ba7943ecd73f319b55efc7fca9c57c0e9e5254dcde32002
zcbb3f14a9685907dd8c97ee43df7fd73a3e53e456d519b1a677c9378fc34dd2b9898c92d966648
zf378526901b3d5128e17659d140e9c3583b82d276611c9914fa64889846eed991317c40a6b4bf2
z5279eb79b094a5f197cd14a4c686ff55285b00c8aeb2ca55cf04c1686fb993ace4117e279c2769
z02b26133e15a393ba31d17cbaa6e96cd2cf4f61b634ce9398698205eeb1172888d4b15a2f25f19
z78bce43b40c28ab7e2e5cc465f84d04af9529183f4638150bfbe006241ff94d7823ee1f11ef2b5
z7628110616bfe4d2824bf9f060ea576c7772f718170436103440e4e60284383854eb3f5bc5d97b
z8641ae6e0706f993a82998e8bf75ddcb14068a849563f11d19d6d128e6dd207d19c4907f63b14e
za88bfe1987442f47d34a7137f0b9125d1ec9aec3e3ac10f4110362b624b2f3790eb63afedf8ef5
z81d7cbbe9056be4d198da876fccdbd0a4e812530af6e2799e12d67444f05503b22ac0ae1e071f3
z52f0fada84365d5bdafdd663a5c5e2fa81a730e766e069414c7e18450d40920ee5b322dfa1e59e
z9d3e8fcc72480332b017a4c68c184e70352d2e4404ef581ac92d622f69c4799797352460e6a0b2
z3ddf1d4ea3a7511f766bd6bcdfe65e4b4fa9fe38938e1ce9c29247bcfd658935119f6ac1ed4fc7
z15954147b1fc3e9082949026efc5515eff626dd8b29460372e5cecdb67641cededb601cd24e9fc
z21f17de0db20c4834ca0730d139962b444f808cc2ade4f93bfea7933f979751cd17e4b88d4e4e8
z53c1d05f0675335f512e68abf265e983c59bd080ae3f42a2594c078ff53f77bce5d7c79fcbf258
z29650a8fcf4a2b8cadbae2011fb1c9f68684eb8246a8a42d581264866fb8999821ed303ad3f33e
z6fc2bc686f5bead80a7d73b99e8046d9c822c7a5976e04bdd73b1fa87b0aa8b1195bb4d4bd3418
z891138f224cc4cc17a3ee0930cf30cfd7285e8afcc243006575f75c794739a9f8c3779c3c74c20
z5c897f05a56ed1c71ac8b2324cbaaf6bebda73a171b3e7326d951b40f6ca6eba51478bc4905459
zc4bcd11190341d6eb1a0ed527be82675abc762560972bb5939cd387d5c399ad3cd60d0cf1b7eb6
z30366f86dce6e5148b0e71ec2cb784854967071b1a8a183223713dca6ffa99b28f2a5cd5ad8e31
z540eb64200e492cdd3f0a95c7f00d45f5a7b0c672e8262bf0be3eaa230998aa6841ae5d04bf591
z0de4b99a7f3cb73916066b500de97b16560e590d76c77250626ff4d4cc0e1f4f89bcbfe62dc687
z67509afa82c3f0b303084be72ead0fb45633c7fe08d0f44d637cb238d95619f51ef07c2e387d9c
z0c6e8f918ab0dad839327d492ebcdb3babbb034f87dfe89b693aae815243cf376d8e99d8e69df9
zac3cec25044c038486c72f83df15756a5e84c19002f33386d3502948a6d575b2d6772c5735ef7f
z5d74cadbac1518dd724c7416b80071487e14d5ef2abf7e801b572d6189cda06a0528f2075b456e
zc1006117bc828634732bb3b0560f2799a65cf0b33f330b610456b002f6f7d21cd36ed8aadc7756
zeb01814b2f35fa0d11cf6a04acba619125dde8bec942b452bee43762f6a68bf65256cc98ef2d34
z653e6f5731793361ec7a1ef9e7a08575effc9acc917d587a13bee3992e7e8eab0f87e3819f42dc
z0ced1226922c3803c5a64aab61a4b81a46e6723ea52be4684e1a127a91a6c0b22c79af75956855
z5ba70295139a1224a26d67f509bad03b04458896f752e21eceb5bbe21bc642d634ff38cbb872cb
z58749e0ea7894107a89e2b3ef8b9fdf150d7e3921a01fb619522ae1c4cd8d8dabb566e10c66433
z23c15a0199ac0d443b86ab853fc4a73dc34ab5945d23a6a4827864bf1597bba03446f22f36208a
z67870a749ced214c4230108424e8eb0bcec0b76aef07dd83495c2fbd710e5c8d165705b37c3617
z60c4f6d83ed9dc2fe2089950aca1aca266917c4929e7cd1249c3722dc9e91e82bdcdca7cc0bd53
z0323856b7cca1ab17c9ec294707493f6e403ef1b737e3c72c5411bb14a163ffab111906783372f
z32a5735df0b4c9f097a4941847c6ac63e8fc04f65ad204e2973d7b34eb3c4d4f492ca0428bcc20
z0c54e518624f1ff99cb251188514f56ba8f28e6650b1f9964c30dfe9565b05b24ea2b23cf07c12
z72e44fe5d19f4b2d25146c5c94166996bd8cfd70341ebf40bf957b0070703b107da29210d062fb
z6972607b5259684d041137c1ee06349711f9b102ca7602af14e0fb4cdaa0d6901da8240b7e60ec
zb9f2aac394c71c3a3d4962ee60ff3c4ee0c5f92ed5ed7a6c580213b2b8c716a9dc61fe3159bdc2
z20bf490782bac09652b23a1aafec06133e3fe8bc1a317bf57e2617dc711c3ec42b581163ca007d
z7817d0b8c8b150bac158d8c40b00f3def34828dff9a6f2a32fa0a5a371875642693e263ef6ccc4
z819a4c57d2c47105e5817895f4bd2bad2b5c01329ee381f843da1a5e9eb1be0b9fb7e920394284
z5051ba22e6bff38a750d6f45d3bdac40c82dab0baf7b9e7832fe5591ecd1ae2f7555479bf700d9
z048c894934d648e695d67e2627d0ec904e91aa5b903d982ce2b3a8f13c5de92fed16d042668e2d
z69419e044a8d4dd237b9805597085438700751fe9b8d898c8265b721474828524adfaf5d9836ab
z26e08d3fc0435e1e83381bf1eeb0806cac3ce583018a61429886dc8fb9892201f9fbb157ddabde
zac3588f492a204e075ea578b5487a58532e82051243daec276d8659f083c4691391e461ddd0599
zd739aa06641e79cf50130f49142c60d4659b1c96a5664a3376e6d345cebf96cfde59a281f90dce
zb3eab7bde2c1ebc6abe16e6f98d5b0e6ffccd75f3638efdc514d91ca6997ab6dcc5c7df8c402bb
zb0708ac750cdc14f20bbf5f730086f3f74592097858295de7bf96786909427e75b67d6193e5736
za6a51046b70ee700f4cb10ffc09eddffbec9ed083be43a68e2cc7129850b9121c7a2414e90cc5d
zb08b750a6eb236aeb243c52a8061fb3616ca23f36889674be87141eda2ed22be0ef877b95f86f5
z116403818651a5bfdb2db698eeca426f1ee383931c8c3e69278050db64f886c4bc08b2111f1e2c
z2e09645944f70a4d4f75118b231862394fc90e9040507198c8f90fc48e2d1fe8ce565fb95829a2
z399759b38c95d74b008dff0468ee8e488dbd5b719cda81f917d422a40db859828865a93a92ba7c
z170ee2665fefbd4852c55f49c4a3c781bcbf8250a78d83a859fb6b5b6a2ffa222e17ce6362b85d
z49d77ad95ad697deb3e4192de2499b73adf2650d5078a3c1af21d5213a84c5f96699bd4002e796
zd9f2ebdc911689fccf6971e1abbaaa618291eacd5b6357d7f3c93af81297a645fbf8a9eecb8616
z98c3d01864ac5fc8627858284ff0646ea7a586c904a62f557ee725a45094e1731332ca1f0cf87a
z81773dc5980a31a8d2f881dc2030e73795e655c0d1ca8f29482d1ec8a2d9c5f6c5237b083b94f1
z409e977899b04df37f2f044d1aa794eafbed215d00c4c05ef403767dd09750c0021985f8f9e4a1
z33881b4ee24ceeb60f818746c770eb3cdc8a3249477c7eaf0830a81d99ac8667f49d0eabc41377
z94e9041aef74b217dfb507e4b8c27d4fa39eb3addc49cb65932afaa674193ce39f737a52f161b7
z0757a877c948340ce3578a72fc2c3ef556dc685d7ab787a4c2d81f7e449375a7b61e7dd9f21a78
z049bb91430be52b454fab4773e149ec6d5947a73d8755984e7155b0191ed884cb86b2d9bff89a4
z37facd0ceb8e0cfee8f2c2db0575f0d3c12e8d6decd832ee5b2fa5e4f21660259211a677b92c0f
ze2d7ccd71595ec27cad5581143708aebd6c97b934acab0f0a038bb25d8eb4c55aba6aa23a2f0ad
zaea22b9da4a23a7cbc608491c31a4bb0956516d3016dbe19a8a11cca0c72635f2315a181382bb7
z5a556d1d1d3b8416dc38f3a934a8475c94e6258b55b668ddb363eb1808743331732f34df5fda66
zf915979606f0460a141903937b94820953d36b2e448922d0c6f3c724c1c74b08978edd97e0405e
z9ebca392980267d487c26d482d432db9a23f9215e2d5a04ee6696414c2a0da123026ce93fbfe43
z00d6d12cb94ead15104a8db3dbb9da9cc9330ae43569fbc9046c929b674dc8d19ea4b3e86837cb
z0aff8728b299e9b36e27425104e90049d6e77e484239966e98c72dfa80c799b2fcce34e8a72459
zc81fea0f69f7a20e36c7ab3d7f44f1f8745a395982ea0f53758d75ef0c0375f9aef434b346447a
zaa948e6607c523aa51bf73083a2a84f641b0fe4f9f5bcc1511c3a4ac275d4a7153d09bff095dbb
zb976beaa2f393802a3534352ce696285e544542d33f13c21c67ec46c4527749f33443e29cdac3e
z440f080ecaf382882698970a50ef3fa426229c0a70ba749631557b8e90cfc25f139b02e5316c0e
z1452727c7d65ed22c5ad194d934b355f134c40cdacf87abd4f2ffe3ec7c95abad5fc3e8e3a00e6
z8374ff69aee9a9baefb33f8e4d66849179ba9762d1e17132a2f2f462dc80b68af7c85d6f34e44a
z102e7f297f1632b7412e73f55c30eeb4307b85bfeb6c61197623f01714eef9dcaec6155c18fb6a
za01c653eb3730623d3d4009bafeb55776dc172a5eadf44e902973160dd427cd544e904b6fc83fc
zf58a3f20b01481af16edc0ac74a0a1acd97e811e05317cc7bc08c6e7724ed931845f31f3273d7a
zffd838d10b33e8bd69f621e941fd57e83ab53b53feb3409af9c01d94458e1e8f26fc013fd03c54
ze153f401a5727dc58142998810fb6411a638cb27f5f13b7a0dcee7dc6fa4237aa69ad99a72f150
z3faa438ba6824360a253f8fc4466d9e0b817043da9472d03986ab7b16c06d380c7ff7ab59f86f4
z9b971d3af58d42b64c9d98c2d0f651372bc785535a23dabab02cbf3869cf2fd9189f1e15dc252e
zfb1e568b9d3b84cb78666d62a830d550a16ba66903d694b640a190e63f26784d02fd7b70df8bac
z65088721fc004db48ac417e77256e0190591ea01f90ecc5ac6edcdaf515d242b635f600f5bd393
zbd23840303a4ca28357f2e5342529a7c62c9bacf699cb690897eed07ed4c1462aa7b7a074e8b84
z23421ed123a9e706e961e68425c25803be9014b84ccd7914a39c21da1da564f2332b296d3df620
z2a03cce483edcde2f27f53932db28602187e92a23b503b13862863dcd57335e584db853aedacdf
z5202e338d9c73ea0c858c1b96ba661abb5e83a7efb1f683172134ea9eacfc5eb9147593edfb022
zf16fb130e3b63ecad36b4492d655762b1501efde2e9bb91096160fb5c90e6a2831d39d2d38ad9a
zdd13614f0462166463ae7c27b5036a6e41ed571bed092ecfc622940e60bdab6ccad15833d6ca5f
z4e48c9f8406b8304b57e38efccb3751f571b1513ea8de240a3ccc9c3e59b4ba5b6e3b1f709af94
zac2a854e9bb4939f9d18fb38638047a2a6db6828529959862ab3298aac4caf75eb0e6debe31df5
za6c64db096c62c63f0cabdddabe1610406ea89db3c4d26e85382720041706558711e324c8c674b
za922beba0d9175c2130ac404d0fe60f82203bb971609ddaecb7bd0b9dcf40718604a5ce75aab4b
z62f67c0707d72232c08d32e244c56cea92f87f0312b373d4aae8af396ecd1c6fa9159d49466976
zbaffd67bb2e00845cfb702a0c7645996e3d165fedfe92d716224512e284aba28b7cf07cd6f9982
ze5865cad3deecfe680d78557d2cb3126e1975affb7e364deb87eeef4724c512a471fa8787f5d56
zd0ec14212df6a042fb7f3155a1027a703fbdbb634e736b037084b04f7def9a11a9bc7503d4586a
z39723fd0dc9d5fc1fc2b13cb07b0ebc4db802c8a583c697477baadc0c35d5cd4476e0619704603
z455d4756d29d063f37a075264eae73126c8c4846860523be851e067cf1eed2ea5b90ed6a66eab8
z27ada81a94ba8953571a0b003fb883133d0e27b7b4da5eca7c52a33e108599946324129cb5fb03
z4e63924c01a525208336685f2b800741dabc212489b7eb72e3d9ee9ea2daa8967e3f6a7efb3248
zf2bcdd0afc07e9d3d8956443f5c62d6fab9d16fb7dbaa88fba8a0289722d59f1f57a2c6e8eb82e
zbacc208263777dcb08bb5816d741b5a1b877af943c46f7a2e82d45b6125581545dd09c2003338b
z5930371e0f8b46aeb10f53095df3d7585a7c211362c6dd2e8f74b467b63ed10b677f29eaf47a6d
zd8b3c167990b8ad1ecf09667eb36aa7faf848c531b7a9c83b27dfc299faf1eb67a75d2414eed9f
zb57c9ee0f38192a84483990571bc4bd2dad77953c26afc8cdcbc4bd4dceae7cf5e76821012a52d
zafe1e42b8899cb0ebd2ab1d4bcdbbad6fe30f3858f0788162850b9eeb5ee1c05613d57011713df
z71d6331bdc025e50510c51ac5521aae786121ea7a5153731e69a62d2cc301c677a7e9638af6c46
z53e7fb546660a4d442a93df348269adf855e419a9249e726e837581bc0dfd21e19dea0ff5c93f8
zb54a9bc3c9f8cc559a5c19b30d23d16959516d23855cb5516cae04101f64c52d2f93491f5447da
z3aa0b02b9204954397119c7d33c963cd21df85197f50d2946c8296c0c5bd20e18e0722d7d4490e
zfc9b47835eac258348d25f97f39d0976b34d35b44bf9f224a3e96da7fff0d629d930610a1b7bcc
z7c0cdcdef5ba06a121b5262bb0f6cea09a702a0e22e3bc0d1fde83deec2ed3791e9a5bed4cfa15
z9f0a8883785278c2ebdf30783b8cc1b23302b2da16be3f1ca50eb10694634003bf4a52f2389645
zbbb04e3cc0f96f3ab6428e4d0e1b1ba99a28e3b694fb22ea3f1646b5044d896f468aa6df18950b
zcc019d5d803827fcce0f1bee840a7342f6bdb17f04b851b71bfcdff980f438bf41e604bd67138a
z8d398a97788647343c960a52e9007d1a9d775601430e68ef3fa56438ccf76083b5eef30a49abe8
z2c24ae850fe1bdbb22758b7e06dc79e6c806a5a34895ac47c73a66feb898b6fc37d99e92ea224b
z66dbb2e36ee11b80aa1589d001b29264aaffd4d0809e8e03ba5bf70ad1422cbef277f2b7a655d4
z3ae8a81dff857e232d103c2c0a5a5dd90333f5f4e00763f3270679e8170bb5158b2e0247025ec3
z624530a8f7fb9133b565faad0b9cd5409c5963107f879b7bb71b8bb404f33766347f81e000c6da
z9d2917d9f43216282b371962f91bfc0902a33ad30484bb831defbc4e03307476215ba2ed455a78
z54a4bcba2d94a455a4219bc593c49d50f4f5b440dfd0502445e2af89c35a8bb0ccedcca4260942
z58064caf418808aab20f623106d5135cad85b96c2c280b400418ff927d8dae2e553a6447cf36f7
zae1ca62c6de719defd8d26721b5d19f1941dde238ef3d8479fcb81bb7dae803d6e563d3392d5eb
z10b66191d5a8a5f270847d71e00e59803ca1769ddcf9820f3db65a0cfacf21da0aed8d6312c2be
zc3e5f46ae7dc1abdd27c69dc67a941b573a14d84300e68e59462cf0a30650042a4995d21cde6a8
z593bd224e4b6ade95cb6dc28a8fb8429988b7686493f277a4f573d6f8430738e4043db308d3c38
z7b89ae7f5f70f3e2bc2bfed869a4882ffdac00175a5bd92c004971be9b24ebb9e38f70f6a940d9
zfd2e926c75d6456029c4a493246dd1d5b9377bdb13131416c55b0f7627766f26c7b8468f47943e
zaa0de81dddb2b65443904513fefe2b39d72f40cc020d70bdf867e255b0128f303fbb7fb0413922
zb2395333048130caea99f75fd1697a77065ada468aba23394d69c2ac22eba8aed1ff77867f473f
zb1821f8782378c3b69364416e976687536a249df4bf26c86b896273596c95556dad55c88df1413
zb41d32905b772642437dd7d663adba734514da8cbaa5441f779886d7fba0e3b01e76bc46d185f9
z713c1da04851f86f96ed06dc1568e76f139288433436f93f2800ee643e3762103dd889e24b3211
z715862851e5ddd2c05abeea8f98f44330133074894e4e332946c14d9080617a448e3dce64ab10e
z595b1353e5407b2f23df651d6a810d0d7d257972e28cda0bfbe63f647b18e5dc65279e97b27e6f
za7c1f2ae49d59e00e0a436a16e05dbd40a4cb7d2c029076823e7d55ba91f814a862cbf36f4a5e7
z839e86c0eb84115ac13c3d812fb08079aaee70a880c2b9b1d765471068913242fcc73bed718648
zba30a9421ceee2edd519a8391299beadae9c0d7466bc1104bcd40c970351d5e1a365b2d7bdc09d
z8ff4c30ee9ad6ef717a5058acee7bf5dfd2e265651b00daff37d32891d62500cb23e7cfd3ca4a1
zc5abcb824704a866703535a1db55472c9595bfe84db3c1f4ec3d71df55f06f309df79201283f0b
z9cab18bf9fddf28ac857103e30f79ddf048240f38acff02aea8f7e8b44278fbb55f6b21082a394
ze409650b5b8678b95a9176af06009a68e56000d53cb26dd8150066a8f7dbeacd82da69fee30a50
zd5b96cb5d9d27149751445629e0712fd5b3980fde98bc2da8238a9ebb6d2a945c0dc00be09e520
z58630bfc436cdf8674d3f5d93933dac024a65cb5d002a9674183e3bab58b2b9da95c232aa33faa
zde2bd1c4910ec13428717843aa58003855d45566e2af78280ebc8441713ed6a2509ab990d3dbba
z3c4e4b66386385b540f6b4a1a2b3b3da1abfff1c566f42ab9e57034a89a226c08b5da4f0887753
z3fe277142fede300a109c62dbe28b2b14df9554a28d17f9c9989d2bf31f47631812545440455b3
z561bb1ca4597406fee893b54b2a7990b96747847334e37d73929dff406a926871fc9ee62f501e9
z015ab7bc3374f09461bf7a6daee2b3e260cbfe1451f4d794839a9060af807ebcce90b0c02cedd1
zc05996537f2afed81dfb916a0bab67dd83bcc9adde005fe1357f3fe4fe65a8c9906836bcf09e3f
ze630f45068b5bd150678a1d27aa03085ec5547301306926eaf666229571bc18093de0dfd4524aa
z279454e0369a6e611a6a70906047aa76118783c7921ab68d805debdf3430cf7a4696a8fcbcbf57
zabc335e33a2a3ac14749e99f6e5f1c752f0f0740b23cea2976384b599d7f50236ae3c3caefd441
zcc1467b1217e0f57c45bb63c2627e22f195bfc7288bff52a81fbda3e14968f3c7323a0b61539d0
zf017972135ec23fbc502e43266df151f37be24d9a99f73c7e45503af6f289a24013eaf850e2e67
zfc14247853fda837a221e371fa1aa2425e438826ffc5a5e25dd50c3355ca4a6978901139c34c3b
zece0de468cfcdf9c42aab6e0c7cff6d092ea977339807a671a3bf8d278f0b450d2c3117c4a8908
ze863d3bf3155574a78f83e061a270823d7a2de96270cab0f99dd2376d73e1fcffce095330e37ff
zd48a268862fa6147ec7371772e095591727c7d65714277b6fe9274e9b5952397b2fe20516e5855
z898dd86b028829382be920d160f4c1dd5e09696536e7bbf3287cc18c94effcfc8d67e5d93ed640
z5dd32715e74a9a1f488a07b0c23c0777a38f794bdfd056ca4df378f2d18f6786951f88b9e05f42
zec971f69f9d296a9145326a4ed881f6fff00597212b3283b761df4592db345d7555e4b54305a2f
zcac0a07c0d8a2678e208b0e67499d10a2ca0bbe5250fd68ce166e9bd60e48180868bd5220cee2d
z78fbc77b6f51bd9f7001648f724384e19a171b156c1532ba4adfe1a1ad80ed555985a42332fded
zec86ef257331f44854bdbb2338e6bdaf0ace0a6424fd4bf52a55559105b745a5192ed48fc2b50a
z3f7764ce188c4d36d0d59044a27d0603072ea7ce68809418f57cb05a8998d25b51ab29ecb95e97
z463dd1f7ae164e4d0b529a293fbcee51d4cd03a0fd91072acfc3b48bfa270da82e02cfaa3e3f5e
z3e24ec8e33dc73f2e9b1f68101e3151a14f2f8b83f4d5c8827b8e428d5ac5fefe1eca5389df866
zbf87fd581a558e1d349ae1e4fb0afe168bcae2c87e76fca3b86bad91e81708c77b9d322608c9df
zba4a1d51ad89bf9bf6bf88f28178db48f607aa4857ac9a30fe756195582cfd50fbaa7d9bab9e15
z924cd11e1d04608598b159c50bce5d2dc568ae89704acfe09aee7322dedeb744d359acd6cc9202
z6cfb9a8ebcbf1318ce1baa5573e53dcb42b30b8ee4e4db3afff4dc43a4f0f285e2ec0992027b57
zb5a6c9bcf26475b5f7801cb9dce4bee3a20ed136543cb4df537d11b33891007bafafe7b61f827d
z8c8b57ae1adeb99a204bf814b1b2dd53e1a453621b87b37d4f86e48a7a69a0d63aa3f916d9d802
z161a56165941b3d8472b3d8d39f22c89425ba81fa3c511d214af2df95e59e3c57905a02d946ef4
zdd995221817125651ece1ef482c704051b53ea1a94b377ee2af15715c20ff2848d55827268a203
zf0e240620574948b6f39447c1fd4ddccd811ca619c162c65b3895702468e50d65f266ddbbf5ff1
za5cdb4f1491c4fa2ce57f3d56859b6af65a1318c8d434176397c3549c0b5fd0c4265fc2b860c41
z97a9e40c5770c8b59dbca18d3e8506ed68e6ebe81a79b0e42355478022dcbb81554387d6126c98
zc45845fe160da9f4f1e9a795a9334cebcf4994016b648999fadcb478be97259f09582582ec55e9
z3a7d9ee033057786cbe3488baa412366d9f98b79a38e958c2f521fb1b614bd932b365e5a1d0e90
z778e986cc39ba84959a2a9f5b04e4c7194e3a0df3fa36d58311a652e3bbd17524c2761de083fd0
z89826998c1a9e836e88003cd0311bcd504babe18377ca93ea6edccc0ac9c55450a0b53f7cd3a23
zd7d8fd94988e40b51ba47ba659a64f05f54ded0c30358706b0ff8dfe8e764685a7574669d431c1
zb2c852dfc68c85b56622345858396310fe76e8f759c1e5feb3441549811c20d1e939476afb1515
z6ad1ca939a42b8daba66322eb30e1a7448625844a9c75261e5f86a6dfe09f42e1f31882ba62a23
zfcf264e8c72f6a9a519b6c6bb2d1f3f6f68f6c0f848e499f0a55708a2001731390b767c76ef70d
zf4103e7f9775f07775a9de0a2fc4a712081763b96b813fe87239c3420ac1028599012a5156296d
z2e3e42b2ff72e4095397a0a073fd068473ee58358bd7e766180596aa87e4c8a89c455ca9d158c3
z80c03a4d81c385d7ab3deb452377969b9f0d154d8da8874747d22218718c6178c1271e75d5b236
zc72e4e37964743091e505f3d058608968d0e69123ca88e21f384cab70e8ecce7f8a27354fd4359
zdf31c065fcbf930ec946ae70aa1b7e8a557823c215132e8582ca7cb3b84378d26ccd9bf0746eb3
z8e41f2697f0e56fde9e8273dc639e6e9e033cc41d697a019582516414d707b62a7d5c35d670c6f
z8c85adac4a426dd24e13878ef555d102b5ece3d6f1fc50b96117dcd67165405d07c293a6ae38e1
z331496669b7597b6a2eb88a816908d52d85ac465530e5db522ad60c9d8272fa8348458ba8eddba
z5d5dcd6045ccb582a0c9fb36f3404da46b82780fdfae5d4ea2ac3c07ff44f44b1cc09eceeec1c7
z687448d874cc456e5ec37b16045caec7c3c1bf64787c4a98a8ee3393bbae46eae6925fb8bc6c7c
z47253e99553f0da1ccf83a378af8daf568104a99990041f2935fa5fe7ee32c88e11ab09f4ac8d2
z40a10107169f203059b1d61527de3e860d559d7fd1b731442a1daf687b08e57bd4ecc05b4cd0c5
za18c3cf1a2ed9fa26573799c4407d6b72e6ccb1ef28266d372b4483bce64b4e4b9f3e58189744c
zb1038d11c4fad8166dba02a4725af6fdd124d0f60e2eb382548fce2f60dae0a7dd5283becccd19
zfeed2767cbfc7c955e67b7af68615b72ced5a298fef1c0c1c7a287e4fb2b4ba542d6f05effce3c
z7148c6f8ed629b979517adc9511a66aaa2b61fe37fc3facaaf09b3b5190ce7c397d7a063491615
z5c1d381f293ae886a7194042fd990488b799261dc3c53bde748422d694c9fc68551b3f1e2e2d2c
z5e593e8931ead9a4f2a634b2e706c87f62ffea97e30851ddd03a0a970e46cfb51564dc13dd5f97
z47ac5ec55ad9083174965967c0b2f96a42b81085003e2e6bf254d194f8252102738e92334d5c7d
zdf8e36ef84dc4913f40ebd24a41018433d9a7f686cdb75dfaa6bc3f0fd4656fab83a7fdee381de
z0fefd7c92a75d5571af5253a4dc3ce2b9405d7854789fc05efe7f16ba5c3b0f25393c09175591d
zc640b1962f38b7f86dc33f89fa0870cdc69f0b9aad310ad52980502f52d4f809429742da07e899
z566ff50767654fafb38ffb428d7ea870a9353fee26f84fee2064c6976b1ec8b91a5138faae6533
z63cfd6b2cc99fd0a53b906af415ccb74b82e9226eb533e765184ed571b5b44ea121b6fb8df42df
z5ae417d27dda07a503bacfa0a5c51d1f693c39c031b2aa9138b751190ed4e54350306e3ff0fb7c
z816d66080e2e92da528d0e8cbae1448679423b9ac8348e72457fbb68d9d344c20e42359390e0c9
z70b83c5db839ed9ae3672ab27852ff8299a1c325d24b8330d1223c3477f6fc07a9e3be51ea6bcf
z2af32d0e14fa2e3acbfe6fbc3dbd7d9f31314a917c40582e670a4a7c4dd0aa245e7123eef24520
zb59912d9f1e4d2d569917c046e233364571a3da3cdb369736b9661751e4c826399d4954f95cb67
z6c160d3e799dff8248d4075c3e3a0df8933ead49a9e5b52ed6fa12e49d715d70e63a26e2d7606f
z56ad8ce81f31aacfd75ea88aa2cc6e6657a45e8372802166b9c3f9e190123cd9cb2531ce53c603
z8842543974843bf5ff66917ac900e1f82026c6f891ffe31b42308d5b6af9e14813c6ce488b45c3
ze128e2a9c9253f32feeccddc44cca0c6d4161a46ddf1d0aec246e5940d122b1da054bf18b29fcc
z8cb1f607be8a2b69a88a2753ab8b29ee8f1aaf1d9e413a05dbf6353ccd9961e012df865a914630
z569b1fe381f4148b5fd3a60aa48bb0dac133db694e7f711876ab92174dcf822bf1130eb2d6fdaf
z545819f18d7f7b7e8229b512822ac26230342366e3246f39eb8da8390a38bc4019196dbc06481e
z3c449223b782effadd88c3a8e0606512c2d561047b04aa429d0a7ba27c79660dceee0e2d4ab222
zcca8b4721779b7df28a766541ba178d895a07bdc87217a152a18c16db70397a7d41984e5f644a7
z630fba56b774ea841d751b11e0c49cb659ea2d1a870373c3c93175f108704530a8b2da08c7079f
z2d2a63980e9f0c6189c2a7536295b5dacb8f6a159a7ea021766af4615e51ee4e2edd0594b496b3
zd56922911c261dc2bbfba4ed556c6ebc8706413949d74bc17022784058653a6972d7a0cc9f70dd
z80a4aa53a7f36a9b69ef73fada8457c0a449891cb942add3b61aafb364cf727b15a00ace9fbd0b
z71311e0c436ff624fe728e2564e68e2d354f92af8bb1e200c45b229b61377207476053a51c19a6
z9235b605faf979d502ce04767a1c4203152cb1c82c85f787e410f21d7a498b6e844cf9ae944670
z04f9afcd3b8f8c861167223196df77cf74e63abd456b8e7ed8e4da48ea89a874612ee3bc2bb345
zb8465678878d2b7becd4db8cc027117838eb137889c389b6a81c73a180eeddc042ece52b68e877
zd163503bb6b1cd44c28278f26a57e4ea749e916bd2bbfc54d9843a97bf34765be473d8bf09a1de
zf392e1f46ae43a8507ddbf608a407e546f758b8aad6df6e1abfa8710657ab32f0fad8d7d8a81e9
zf3ae3dde33f0965858eece197914f2b78d6d3d1fda0afbc4fc82be2c5cc3aa0c8977eacc5c5c6b
zf872d677e4cf44ff03f8506f2e9249aeda9732e1f4cc786df46b5111f5f967757a2c305761e2fa
z2f60938522d88b6d4cd82ac6ec8c5b01b3bda4b98df7d988348b25f4587c3b1fa9148282f94b20
zb00eda7618a62781615e0d8b92d75e90b33c5906f46c93d244b30e411f2830ab19ff48b119a0bf
z4f3b68fe382a63109b634b6d0abad4231229d8d41a2b7f27259f389f6b49f59dc061c464a9760e
z6295c10f421380b71b6f0405eab6c32dec3340f632262e9dfc8b45db1f6fbc96c7a12bb8b9d6e2
zf80c9c86a50577488da990e7f58bea6dcb63b9f41ab2d65245d8d6bd6691518df6f0d20da4a3d8
z13f1a8c13e0912d6945e845044b34f85018d7e4d1c264e1c8d4fee6d14ea473d9bee8df2e12ec3
z40caba6477c74b170f4e6cf473f2aa4be24b055978802de015bab064d9e883f84166faa3b0d1fb
zaa3a54a57cf5399365bc591e0a5e970d2912aa944fa420cc53f8ddbfd932e63caef44e3b7740a9
zc631cadfc698ca41849747bbf89b8cacb00a00e6650f9af46033c96c4dd6a96135e93ddcbd0811
z9e9c7b53bab4ea144c42bf0877874406aa70d8b214f7532fc0ee319c7b9656aac704e6c900c7ac
ze440995974e11f7db5f24d911f7c97714755f32a111d5b9b5ccb41984146dfb048dacc433354cf
z7dc98c553b2feb2967eac45509bf270e351839dfc6858d0e8b8bf575c008258e8b59f2bf143e92
z75fd0da719bfa63a1126421e50292b737cca654fb9beea3808b0f8e193465d12254ed6e643e430
z822a7492a98a0f28997f254bc95b6eae8c9801b16050d415ab3d41d32ab04cd0dbf93a216a09bf
z1a3fcf49fe5338564243b14ebfd5ce22e035572ea5e701982b85526def035a265e8188271cf4de
z2efa92ec91f149990ab9bc03c81842f5c8039fcd28f6ff3a909a4ca1a35858655e631623ff373e
z5db325cd845a7078cb3d2534bb8d6aa3131add6ebf10cc6c62b93747e6374d4f47afeac0f81094
zfbcbfb0b9e98f02ef0dac5056cc20672989cac1324d6c9610352183e414495cf419157c8cc8522
z748ec5d8f9e0b28459018ca09139f727d95c36e6a9724d36d1a738e56d694a285273c9686d1b76
ze3601334e426a22ad7a436fad0c23dee4d8dac5125fa38ec1a2e328f709807e1124e379c68ce43
z9800679fdc93ca7d0cd7646b2fd58b6a0c4159239ea7c347ac2285aa80642003018118f39eab09
za0c74e15492b1e2d7ff295313512524ffbd5db288f434397a1942c0f3f6b875c3922b5802945ab
zcd64e6e20d2926a232ddf26b5b93fd55b070bd352fd5ecd0af994599735477d274f91bc2fcf175
zb3d506d17df573fa439818982abc41574090d1ffca3c49c955331b8ec9a2c273abdef1ed283030
z1fd04b7dc9bbae9c083f70e56c9854a9c30ec6e65f45101c945292d019f96eddde00845c0ae69e
zf0eeca4e8d183830834cedc5529d4e5dd286f4e3f623e240e8162c9fb75c85f73f7d5a19bbf126
z724f09f3a25cbe458fb3c7825ad1b9ed7736c3b480faa3dcc16079cdd830c237fc0766434c17a5
z9dd54ac7242cdba7d4989860f65d314aee6b9ceb228913643ff290064f05f208a9b5114b530df9
z42f261d457b4a20a015335ef3969c9dfe45c5db16110aea1c291adf40e58f69eb2b6102df10e89
zd715dbf10425f64cd3bbd7eba639c22a5efb81582dd34df02a822f9d027b34ba6a2cd9c668393a
zf59b896f478ad8684bace12928f04c21ae32ccba853b2b4a36477f1136b311216225877c50f1dd
z80fb240967c1a710490d205b540fd16a5e0907708a7a26b9f1ebb6201cf4787ef8199353cf712c
za0fafe896ede90a6d22ac3005335d4a83f58f25ea08978d92dead8d656d1b74bfb46748072c605
zc2f8e7232cdee5d76488693c91125c7c9488da9b592c0637be80fab19f539e248537ec3b964df2
z720a986362e80ef9ed9fc910044eaffbb4890f1ab0fecf83aebae4c67dd46cc520b9d646dd687c
z50d82a8f5ad1e8587d81db82a2029e010755995952234f11927008648982f85feec5c6d6edd169
z186c01d1487814a074c220cf0dd0b82dfcd54fbd1bfa93de630ccd77e51acb0c20c1af9c29c34f
z9a2439fa3e64a8f3556b937ae37f27ab5c125ee00f78fe989268b16398358bccc8faa8a0f5eabe
zbedc139f7aecef6dc13e96aad03fad4d0d44deb690e9decaf188cc6b0943b0a39e63279cedca8d
z08fc7f09e66402328ed2b854ec8ab46fabb4715907c4e172c63d969a7448680708e89fcb6e4426
z3816a93ac2d2072a3b98afe583aa8055aa2ecf524bb5042262707c71e1b8bc27a9e357fe3af368
zda0ad992b74b21de4374ce41096c48c82657648a0fc2bce7d54cf6479f2c0494d9ef4f98ca8eea
z8b21dcaddeee12757d1b183cac79b1cbcce013163bb54b2b979e311e6da1ca4d598ec64e5ca027
ze2f82ef0ef149d21c915e80394f035c64b40dca2949bdbbb2261683e184ec1dbd59a5287cd6e92
z93caca19625f352e3508727213ecac9c4328205d810ac2798e0d09e472d28d5ecb58db59775b5a
zb605d2af7a91fb0750fcea413ec91661be7220f805274d1509d03e5e0c04d60e1e1e5486e4bdca
z35c6ac3200d5d5cfa038529f76e790c69a9a07db46facfee2744180f3d1637f84ed920753d31b8
zb086508bb0171096f9ca32829775aea853f34dfb0e0904599b1e5c52d89e5d5c7bd5ab50f18a49
zdbb899548d4550160f78f6b6c1e40f7db8acfba04e8ec1e5d9d0c70c6e119f1a6b97616e4239d8
z324ceb658546ddbbc1857d82270bc72dd367c8979ba457a948b7a6532d43d91fd81d8e25e18dec
z54b42b9ac5e6b02d2850fc2367206bfefdd11f325b733cb46c4053dfe3bd5b79278bc019a4619a
z54a18c94591185c33c3d80d07602903beb79d29a7686f3a83b4e3b66bb1a838b755524b2416d54
zdb7590c44d6056a313b2ad6e37f00d9e595f2f1916ae1fff256161e3655bef08e01a3739dc9555
z5c92fe26bb0cbf28ef9334b152f772f578fd1cd0a02a98dbabf76f3d7fc1e260d1d241a3644ef7
z664ece193bbb4bae527744a11c24483d7e524b8cc7fb4cff5a0d27d3f6925aaf29c720dee42191
z230742bcdccda11973fac73ebaabaa57c0dbe934723f0a45582f3c98fc99f7826185a697dd783c
za46d071ce8dfb223d2335ba337c0d06bcd1d6a240f7437575a47dd41df151c07d8fe91d8f34c80
z59ff274506494a3f720cd07686981d0ac3bfbea82a921aec58906c650d50d11cd7f95d7ae1e75b
z2b4079383ab56f57535c3a70f7c27109255fc07e27d8cefadc45f7a99ebea20c338b159de3b996
z59088dd212feb1361a5e88f8d76c44a873938873d3906d6227317b2d7de4897359d3b421fd3831
z990eaa003b809c67fe3908519d8a9ec95c7857e91a7806f1991d54631ee01aeebdd7ddc5165793
zaf7fafb4842bc4194253b397c9011472b10b2511af0149432fae962b3acf423f8905695daac7d8
zd2515d044bca9f1dbbed0c0002d57d88634c4391a0a2f821843c24b2700946eba95a7f8f4e68e2
zdef461219afffdde3a4b48d89f67eef2e95c898d8d877e7cfb3845e9b5c71f691d86379936f6f4
z0ad064ecc3c058ded2d42beb67914a0040a8416c46f552fdb9fba61559572d6b7e95c30df77aff
z90ee9cf8ab53fb53ea64cd4be0fc7af35052af78dcbdfa0d3b71e7a7aa8683b56260b385f5f734
zd7691eb95b940084294bef4adc44a78472f387cb8cdeca22d8e035bda532e21dad839e8c0b9093
z5cd15b87f919eb68de9e13f76c090d308efeb183af2d77582608dbac4879c8e3de5c0d1f52f646
z8e603a243312d19a0c00df41e39e9b5a03c3e522afce0023db47599ef2120374c9387cf3c98f8e
zeefc084118eb42e80dee217dce36830ba440abef66615a395e0b4f316dd3ae54233d91b08af0d0
z16179f1b90cd6a449cb3f6d633fa7c827a00e091257822b6c5595675ff19859665e6ba6b263e69
zedb54fd28ddb919b310ae1fd455882497abf3e416eacf2a6855eed7afda858cdd623ed38d42830
zfe00079f0da8f9bac7c1df4b50fb6a92f12451d46a31b93b4584db18a347690c61a34dfb2a450c
z7d92c516025334488c8346c5e0e4b94bf6f7159cbc9ed91d59d13e882452d1e801abd5852a5a56
z54a249fe617bde3e9d51f2e11bcb24069442ba8fca8c1067ecff226c993a3cca9fe674058a89fe
z91dccdffc34150c849998819bd45d4814b979171d78c7f475dd7f171716f8a2749766b8b41dff7
zce4593c70402d37fdb6deebbb07fdb9b86f65aac58ea6d023ec54f8b569f2052b6c2fc79ad6c7d
zc2d92257d30818454886b4a53d3eec2b013c56aaec52ab501622484bd8cb408c2f06e3652b58e2
z740c35dc61396a5a40a688bcd8614d6f38427cae750086a0967f766ecd66fc8a82439507cf152e
z47ad468afc399c858d9c19194387c185a6dc7f19b4b3fea1123f09df7654874c3ff6e5c847dfb8
z17d747586d5ef9d68010c06e709176c7bd824383646a3990d8b766ec401207ef89547e6c4ccfc5
z109d7832693b501a1040beb71acfd744745536c43328f99fc418c89120a4973233c1a282db22d8
z4175ab42ed9df65d9574ba71fd1d9a1bd72ff4462d3523ce69b6169318517c3b299d74cd777f72
zf09fc96c356e36179c9fd6c1f84c53ccd339b46ae5152199f132597f3b25dcf4245f626ed6f672
zf247e8dd8b651f0362c0d3da6466fd928bb8cb18d468098b1651e8e818392c3866650cae21b6fe
z49e3ff901ddb546a1cceba27f04c682959facf3c476b8fe1ffa58f6cd8e26ca898aecf96e5079a
z24346f4e92a118620c0179e95626f6544aefde073b9e790c8c20ee26288e7f2143dbb199ac974b
ze7c59913e1a215cf3db225dcb311afef89249bd2d2cc70e8f5f69496c1a26329d9b1545eb6e118
z26147048af86248be1712daf9bd57d2857e6bb120b76a7345699a31c68dc278f71aa8ecc3ac341
z7ca81f9de07d525160461077ab915439703251307ef021acd792e7a71b61c2b489ef4980d14315
z205e15ad3aaffbf1293396ca1c34f408f68fecc94ea32b34e7315d4ceeb2ef859db3f52faae6bc
z7002ab2a8d4ecbcb59bb629534c646fef10d8b0ef8580b031d58116d0937b8abe8606dfd128d4f
ze3172a8b173dce39395f88fb87f625cb67cd68ea37c72f3e39d37a169aa7e6087813b56ab0f31a
z453022e6adc2f04fed60ca4017493e73859968852a24a1ce506fde8ac8b99182bd1dd614f115f7
zce2e46d126bfc48d33a8eec72c229b19f94aa1e572d259932fd5679317fe84abb5b94c63af2308
z98235c5684325577a3c7fba878bdccf1e9e92d5ec7596128168433082aff50c67f97677ef42c90
ze90b9a64049882e9b107a7bf1975e49995a784d71d585f414ec0f89da2296e60d0d7f778c4af75
z166f508b1a59333eb81ede6c94f62b30b6ffe271cec75484beb314105d9222fc39ed2b9751f16e
zdf9ce0cf04062c0a0851f32f028038840c794a4a8aaabb936bf76b11766b93c0371b7126dbd7c3
z3096073c3c7f0bd9340ad3f384345e42263daae7b9085c0417c3735d969432b59993ffc05f65c9
z48cc354cbed798545a82fc1da6f95c4949adfc9e235ea4bd41b52c8164743b6c78694313461877
z415c1a9b7fe9949ba8551f1634193a257f4ab506500a81f6d38f6880be5f55bccdf0c0d756cb05
zdbccfdbacba1c30afdfe124eb138e179b21690c5d59fcd00caaa69c03096b63c6ddb5cc1da3067
za187ddced8039accf813405c6ce9fc0f0a8e64183f440e352bbfa2b2e0dd91632393043320e55a
z1f435c92012968232c063f2e40e0c906c7e97e70a93b1f1819c397de9a68bee63b704b3d51dfdb
zc996457c612f46979ee3395b8bc87d440d9347e218608290bc742d363f29e2b4e4f99411861f17
z3915d272171cf4987297788de7ccb9a515256efdfa364b348f2d9f935f36f12296128c6f51a7ae
z476df7ecd095fdba2dca50a6f58a22afc666dfc4fb291feaada8156584afff81cb27d9c2105a2d
z36515b290536094e29e01bcec7b249387574626f2da9e844129916179ea8dc2823c6a863fcae24
z101a60377f38278d430c03548cbae7b5406e4e6cbe51ada5d524f8e57cd66ec4ebca77ebd5e1ea
z5e0c05560e067bf880c8c41fc23fafb9151a7ad6d4eccff00363352dbbfa5eaa6d766024386fac
z529ddd9f051d910754277db77cea9428ffb151950b915f701980eecfb43fa8b4ed53b1400438f1
zf4ba70334c3ca3a0afc74fa69d83530dce6c9ac6751e5f8d971fbd9cd589db70c7d75455b54b93
zbd988cf353e00402511bb873bef4c0d1339951897acda69c8929cdfdfa6d4c4551efaf6ab009e0
z3b9edf49c27696dde782fefcc9e5fba0c0dff35307962b87444674021cd90d93431d5af186c817
z18ec7390725beae6cdc6f63507b100011bea4bf7ede78eb4ebab8066861186ee25bdd5dd0c3740
zedead5968f5ad91c89487bdd185ac9bb8bb7f6564a823454113b4c332504f142fd9c7c43dd44ba
zcdbd75784ad405570705f85e5eee2c2db7bef6149d868d32bc3f5ea9c6d1865841e2d6b269299a
z7bd2f92353b0cb5a96f7b5c3fcf07f755f0401f50ae420847609200b290744212004409e352027
zb800bfc38c251a7e8f7bb41cbf3b6601a573ec3787d9c8e9895a90bcbe8d819040299ce25ae161
z52000f6fafc937abef9603230a0f55ed55d87e522b2fcf654c1cf6a3b57e204d148f4e60612e84
z04d1bef4987f17956831d82b70fa820a01d63743c871d3cbde70362e93b7f7d1d5d2451b108435
z92f685195ed7b29d854c232096f1b9cfa0467a50a64573cb120d7064433fe76b526d85f69b7874
zfe3ffecfd99dc3d8539c07a209c138a151bf0ce17500da74d45982696e640d5a788786ac4ee81d
z20a1cbb2e34b63412b2cbc4504194c79037572236881fb79abbbedb08fe1762167af7361a2a41d
ze2b9b6204689677b8344572d3a24887fc6f88d22ea6deeea59f4f7a7d29a115b29e4cfdc31c230
ze4b990cad783fc4256bdbcf4155b0b37f91b0fee42315745d99ca57c5da114309bbe0bb05044c1
zfc5767701564ea19c9588914eccd5612cf31c32b934d7575a4c538eb7a84700629b4a35c73fe15
z0249da44b12790c9ca0242acd1bffb6407af12954307e20e6713f898a42fe5c32a772dac5d0f9e
z231eea8808f999cf075b85e4c727b2de6178dd1083c31033b6eb1f3bdccb8a00d1cc9215e448c1
zb024de5e1dd5abe60589fd68c1f900651991a7e329fa6905bc71c2fa1aca983ce455373435ae33
z071fbe9e7ebc832c178ef06133e2131c1cd562bbb88b37364f9fa1a9a36fda7c543a37aacdd0c2
zc6a5c481c1fac02e20b13af6e00d8fd732a20d192fc8fde9bc6b95fa5a74007f2bad3ebf3c6854
zef56f94147535d57c8af7a2b82971b69e4bc14e4d578d68360a53f6aea411597067cf5528e6182
z97584598f35fa22d53738e913dc794d77fcb53d7aa69de35e6f697e14a0572650c9db09ce18d48
z3df56f2ade09c3f79826100740da5b7745cf6cbf25c1c052873c1061cdc8aa49999c2233fce264
z36950210cb5ef60909870d65231e56e6241149abc7458ff3eb0a607dbc2707be60960aab79c31f
z34b3ec1d7d1d57a7a81a30d926f330595e8a9eabd0b7df985546f462125c9e226e0e71c2204414
z93961e8f2736268ed57e57c8c76a55c8d90b575400bc517d1ab5b1fd8c625f40fb4d7e15f457af
zf37a876cc83ee6191b74de1745cfa4be85e15c368034aee820d353e359ca82373eca3c5133c6ff
z73dc73c09321565fddf7c1ab199db28d7de7350d4b3ed6be183ade6efbad3041abc3bfbecb086a
z6e26aee8ee9480b34256e463a3b6e58b6a8c7d0a6fe9463017864276518b30c6425515ec4c7a6a
zaece07d3f282713e58d05c0d2c999d5a00f66be7f6c0ddaf9cb1993b0d3119abbcae26920b2703
zeee545c3bcd559a9364ab02e1f6d3595c56b0bbc8f9b5404b9b8d990f24379ecb0a57ed3285405
z13019d320d29c1363de37bc2ab2e19cabe57e82236b1db48fd3517b6e283927d435a6f52bb02b8
z5de790d71a99dca0235bdb0190e4f8fd15bddce2517d2f9bf8dc44e06f413f1300ff66c373cad8
zfdffb0bb6b14f05ace3b6db6e9e54c7985cf75db55207d1dbdb1d033615b76440e372c5876e74c
zfc147aad9b7298178ebbd6e52c128cb6890cba2420f7b7a98faae119f7d105aa4bca212eb16810
z13c122eece68b10280afe6ac81a6cc18c600471c9f2ef361df2118cd6f8f2dceef853a9c1f873a
zf557901fbf30d1ee6338ea4463c8fa108d13dfd2a94e2b7b25f09e6deedb78b385c619561ce9f7
z8915cd2ed325407bf64da0866bdc9efcbc04862ed958e0231f169856f901a69ebb0d3946aae434
z0d95ddd21c60de3fec4e01b2bced0e2f5ae9aca77760e7acfef55d61023b50b7091b46a603a0ba
z8dd6b9859b63ad0280b6274dedbebb3bc9bab7c90e21e2aea4afa42bcb4b90e2128e6e1af1bfcf
z11053e03da9376b265d93ff3049d63f9b75f774198e6cae6b318d673061ac4978edf289ad7f36e
zf5f61ca65bb81f68fe7be9331c9c5695daff3183d53ce665e0a29f0431055ef0f2017dec7eacf0
z4bada10cbaf4d16fde7980c96457dd29b67c9de05e998e117e05b5f2ae404e730cf87205476df0
z9b2b31b7ff64115edc08f33efe819e51ca483a4f3b3e0d2667ca7b08412c5d408b80b89af69735
za03f51a6aa4fcd1d0425d9b6067bb34b6bb9f37623f0c67e0b4729dd0a36782d86675f63c71bc3
z08b5bc72d4d5d5ad7217c367b3d82a129b379b9ddbe657e0ba73f6a3ed70768f952e9a42f4e6fb
zf9af268d2ca5a56a0bdc20e8baf6718b7c8ffa7f69191cc4ddd03a81544f41ab71c5918e1aa6e7
zbb702c0ed4655255d7ebcc769fd2d46340777e3ecd0e1a5f34e46031e08ed8197d5d6cb08aa872
z950ce152ab7843cf7046d9f854be2bd5f36954f41b183b81dfa0059cca8dd5b7966a01e45ec684
z931012c9f48dbf9d195f3cb3270affef62cb56e0201486012cafe75d68dc31d12cc410ffb7422b
z089df64ad1b60a4749aad41948699534e088a86645b0a729f70600ad2e0acf1b2069cf5c403857
zb78650b37d4fcafe75f95a1f3ba2f699b1d7a0241fc8a573da999fde58b0c94db3947f56fa6a53
z99a311cba8a25be143b4ccff2a98cb91ec2c0ff488574e52dc485590a243bfc3270ed490bb17ca
ze9eb95056e1b250931baf2eb46b2b2eb87a93bbb81971a5d6a4877d268cb8876c3543804428f04
z5b160282fe1f897cc67b8f5703a56d5ba70d138b1e58ad051259f87bb6af2edcfd2485370dfd85
zb9cb7e3d462e68cd1c729dde5385f475c1a7313db06bb5a626eb80cbf4354ec62d85945f4693ea
z06fc6d3e792a7935a74440b692e9dd6fdfe78070574ec005ea94b4381e677a274a5477609853ca
z123cdd100a00665ef79e56987e22663ac5ca3de01e5466a4919d30d3290a84bcf1cc4eb5a53a52
zbbe6c342caf91893f92efd3ad8c2a6513e9bac0ab25808b7ac64367345fcd0b41dd1a2f9c711e9
z94c2076990e32dc72cffcda798e1109a19814c7252372202b6dc3ddbb9029806e6171daaecb1e1
z042bd875717e849491ccae1145da33cd4474b5256db59c68215ed7741fbb2a3e8e17d1b8a7725c
zd6c3a9f3f23b363ea16bee1c52cb11786c7423574b219391e79adecfd9386c02b8aab668730f51
zebc579f4afd99c2b9b063e509d7412c72997e2967fe656368714a5f36fea6f4e97bca37767de5c
z99bb1d0a0410a2024e138be7c500394d5577ecf5e8d59fb88a1caf718d7ab80000af0293a2e4d1
z1b32128b6c92caca66d29dfa91315d9862f88b91217ee11b81bf60f2232dda06c0aebbcd318553
z9cf93793af5e86445400efd7050cdda815a29bfafc36eeb715381fdfa61687532290382b72e8b0
zd880a919e0d2468190a4005f084ade4030fbb680b4eddb87a2fbe11498ca35dcba97b73b2cecff
z19224ae7187bce945db623f0fac432c51f4f3f4b52b42e445bb35c6c99ad068d88831779f297d9
z1f5ad76afe3c8d8203bf5b5f4adf395e3aba7bbe0b69f7c905c24f07c0cf497445ac33bed08757
zb3f01f0315ad5ee0835bd7aa6dd8497f2adc17983744d764ab4f3f43ee4084a6d4e219bcec6869
z634d8e9075bdefdd55c41c3db0e242751f0b75b8af849482272a8b1d464615dd8bdbc544f8ecc2
z5d0c305b60d67555cdd64bc4d452d43ba8848de3fc096b6714069f1802d6f8a54090aa676dd9bd
z1b006cd77140a230cb6c26ef09a7e235dc41f754802b9b0158da13b35b3534b6225ec23e4a43e8
ze1308a290a6e57a259827e4799eff5d16f689a0394b37965df2ccad326821a0b31c418c148c0b7
zcb75a6a8ce27885e36a9a246ff17346719b3e7fe3c5ffe7fc07a2c9a2bf0400a3412efc2d5b7bf
z317630ae528c6daa8adf7b43e2aa80905370e0a23e79693c5b1d8e1d602db689d294a953650261
z28f8332633d026f6454e2be31c33e582875b7056075fdacf88d57fe0b2b67b775c42dd38bba14d
zcf991f9e6d7b13b888233a77f4408620fa5eb60a96c90cc2547c1f2e3018766489018570d16610
z42ea4f9eb2c942072ed77a54af2c2bfb73105a4d7ac4f4e2a898802410582c6d48a2ab23afe082
z5e12bb38d762a67a7ef1242cb423dea5b7d20b772d2928b11c07c137dde5c03546fda57b21c078
z1775b2f835547c59c8737af3ac8888fa6d3cf24eea335ada37a13fb2e286dc2ac3e013b2b061c1
z9ab80e1da6594337b82c26c9f14c858b4129329bf0b2fb5bb4f2f0556408c21680c0e37131bc3a
zb1f78edc27b198554d5a920122b34e9c77ce3e83e65eac7548df9cf638e1de27f3916befeff90e
zb07b962d0d98f36f8ba85cf601c0ce9a08c5fe9a78b2bb2664ec08e30ded2b37b9bb6c2ec72db6
zcad2f795509de6e143663db2a00cf3aeaec0c5719ff4cf2080be1cac7b540fb21f5e7d3b91a3d6
z55bf6485893a5824550b4975bdbe4f40b85e40bf12ea1b5f4a0c75bedc8b9ef45577b94e80aa82
z110c76b179c3b02b0df8d4b1aa2fde8e79d8f983906fbbb5b85474d77e640bae0f4a7566d806c7
z10f3b47ce58b77afb75549f2543b41f5311c8467e7831725fb7b89a5bf79a873d9ed58d4315fc5
zfce7f46607583ddc207649f8c186a9acb3c1c5b36caa4de64c6f5a6a1362f3dcffc9b36edc29cb
z0b547c9d5502500c19af84339578830567f4a57022443b86d6128617581c19eeb134c4f9067deb
z7158ad75fe15261d09b386b42092594a71300a10e33cb9c2dcc93af380b728775ed2bba8da2130
z31ab96caff3de5411e5620fb1a4d9557815991b5689a65041ec1b5c52444c861a2bc01c41631f8
z98f86bdf362da2202ecc19cc5c2f04cd7d47c557a95d55e70661802becdbc66aaf4db9bdbc6640
z0c12f0e2fa28b99bb41dff99e619128c1a520ecc9aaf2846bab50285c08c734e02e508f2a9ae08
z6d8779da6b629e20ad442171d8d0be8f0bc4b1e54ccd86a4521e53d504fc2846bae65c0c6ee257
zad1cb40c1091dcacb1afd933d5e6f7b2fe2215988b3084cc2a9391a0833642b90d0cd86423ec42
z9b0cc7324bb70d507b037dfc169f1a78549fc942f36fcfae64abe25e4866227e7eebf48e861f00
zca46e9608bbc6299af4e5218ac46606fb1eaf7ed1a3e10d0d1bf9b71a5bbfb6882b010426e04ee
z664fc2e2f47e0d9f92a869f687ba1eb4b744edec18747c72b43e7032f70a2dae9ec8ab11316362
zb2608cd94ca9398f6ceb1dd661cdb167f8142bffc47d945ccfa718461003dfc3602f54d610bc84
z0d49088eb573ae3e892e89d2e8ba8d507928807d768b7921988bfbceebcee753191deda7bfd321
z1421851c4a4ea943b33c228db944b683a940f5602518662fc7fe15923ce1f7b249d12aced5ae8d
z8bb44d2b7f11b86ca103b2851cb9cd5dbeffb304391f5de4e22e51c82203d101818335b75fea21
z80fa9a8da13457743c7a3ce29eac388dd7be493cf0a902dddab380d2ca00b74d46f31d784348d0
ze86875a72c7e3b0588cc44bed2964caf365c0c70dd4ba68a9aeb12c86e2a75f539258011db3a39
zac4b45fdd2ec58fc075240b9e03626d8c57e2b05e7a9bb281fb9ec95bbc7049400c51412794d6e
za2c497eea2d132d78ffbc9bbd2ecd2cbc9ce9ba4e44e179ac1fc191c9276598bc43d428999d559
z400cda7df10985f30817bd31126c7d88525e19ff319e2f66cee88ed150d629e05121bf5964e83d
z649031957b4e7009d82ab4a1131afd04ab4bdb3e3415aaf65f12693a74beecb8c1739e5df6e722
z076b225fbfaed2a47cca739919e01eb7e54a6ac8ec64ac53f9a9b19c9d2492e53344553101ecb8
zca34a156daf9718a931ed2061d823fd6ece74cc208a38b022c184d4cee71fac9eb199ee12a3d42
z9935cb1816a92a44dbc2deb0412a4d92ab7d21262e6291023d0192188e5ee5d1e204a7bf4b0571
zd57f680c666914587a64dc83bb76bdd535328b2ad60eb4e93d3c674eb8015bb2e3f012d5379bbd
z2ae6b29be1e85b15567ad678c51ae240650c3113b767412b8434d5ad706cfbd99cfcb66a5b7457
zcbed3dd38f78e1a178856497a99e98bfdb1674f72275922e4daddf305b582329f07feb36a4df67
za374e2dd5b19a3a54157c76632631cec2bad7081b7fb96057a55c733798402c481dc82c16e6c8f
zf94be07a65f789caca79cf08e231abc16bd2e5484942ba33e0ee65098593b8f2ceb31b71093a85
z0ad428484f2de88fd160035cbe4cd975666abfe1b5aa39cbdf9b7ec27aa00b808ef1e7c44b2db7
z9cc6e115ad0fee576a90e43f30674d2dc672aae7c92d35e055a3858cd0ff3e6a6e2791a36b6679
z8ced60ff507ffafe1e655c19c8a5f886f78cebb0894deb6919895e16f7fdd94833b5ff5dbd4bdc
z46234cfcd90b509779f08c0e527def5a5c1602b19a39f5a4217b058950515111744370e8197930
z1a4124b6e4cc64d04c3abc35b0dc39c5f708412072a725c9415eac7ed4a7cceab1f90da3348f8e
z2df00bc8bb94203f8543a3358b72365b85708a8dafbd570891a6c46ea1c6dd682609f95bb761b5
z3511649ad3068129fde1f0e666b8d4f6904e546bac9c6176636f93529d2bca7811fea2e3585ac3
z61592bc1ac026ae9c9a5626915092b46b125c61225972e5ebcd9ebd11f0dc504cc0b6d07484df1
zdf78294288ddbdbf0dd1ce95bd4cb2dfe6c7acd26854682b82cd593de649cfcd31daa4a0620808
zccf0b174fac8aa6f99b70c23c1e9a6eb4cca8d88a72ddd0cfd26efc627eef15f837efb9d9e0263
z4ec6562e06b8aff222bf89385de8afd6f34b24ee1976626726e02a72e1ef67854769de3c947017
z740ded282501f20e29e27da03ad8c2897c14e74351b2d6cc42f27bf946f2ee142475dbac99e9ec
ze3a632276b9b3bbc89c4bfba59e4152161870071213fb63f78dccb850ef946a247eb751d8fb92a
z47d4e0d003a94de58757652fc8daf0de861242c7922fea3eac65d1a0425af7d0c5302069ccc2c8
zb06c774b3af066d505545319c4655db8173a12100b89889b1ed87cef9e9b00d5bf23de0bebb50d
z74256c13846f99cbc5e8695f327442d211dba08b26710fbe8e4fd7e8fda6bfb4e6c1dff59747d5
z84a4448d80fdacabdcdb2fe6acd88b3998739eb52f903d6c5d739e862511e94ec1fca7a99a50d8
zddc25e4956e57dbedd1075dbb433b985ee3584f463a14dbf512b5d730e8c1325e0bf4a36cefd04
zcd1b262ce4e414051bb67827b831775395d0c4c5c6bdd111708f1ab61889c7cb3d0402bba385de
z97bdf6abf4c617492bee421975f7c2607bfdacf10daa55a093adafcd1fd7db98f8a4e0ccd9bc66
ze798c0396b418fdc2d20fde6160a123c6fda4b5d75ec7cdd3dfdce9138200319bdd4977db0b1cd
zb8205eac4285d81f5c9ba62cf2e5c082b66ae21d5dfe96b129c1a3e92f3078877ddc89fb222e13
z6a8dd5874399dd64ec74ff6ce2fd2b5bd2b2181cd6b4740540fce68e933b4a2f3eae3191055255
z869eee0cdd5920115241ee7ef1bbdc84d4568ac815c5841d424dc65b867d5d2bf8e6ce5e4ffa2f
z3ba4c0c2ecabbdee00824a9cc9e054b7689a7215b8a62ffe0259aa34190fe86d0af7d9e2a59a33
z3e350eab6bf14abea5ba687ad96de2c8cc6319ffda1ad267af99085a1eede182a281d05c5a48c2
ze8f8d5759ed2ca79009fe4c65f0d6be6bbfe187b91a3dc4c62dd86cc06133bbb5fa2fe30d4048b
zaa91882b4400083c940689eadb631ef965c7dc9a8f0fa3dbe84c50325e85d28cae959f5443c763
z6007c6b5feaa7d803d6d87cc82813633258304500c4f0f8343a7743bc111b15c41371bfd3c4ba5
z21073a284d736916872dccba778e7296ab88dbf9cf7ad08d5bea6ba40b764a45a845f8e07c3f82
zcf4d832ea2994b3ab42c8b0aa9cc80fe4643c8232365eebcde737178370e7731be5b7ff630c1a6
z2a249b2f26cf6d9c50f7f6eba2f5bd1386a7ca6881641e16897de70da7c92029041c7068694dc0
z7515ac0dfc130437e7f588661a17017fcb4745e9b898559822982f551a16c4f2cfa906a80b6dc3
z2a8965aeb9c894e3c709ba00733364e5ceb5c8677983111778de8248f91b36e656a58e60c2dea2
z3cd4f098c73d72dd8b75b33c38697d0f85c43aa59f0253549d279c309ce68376e4de66c77c2599
zf9dbb85615fbe54e6534f0a133e559ae8f37d6a06c310cbed5d1479072f0b5a97587515e9d316f
z1cf26d12bbc55d137e8d722bf475e6eb265be8900be806f70d1c9a63b930cd57d72a6667685c09
z4641e4af5f73571a9e35f76d594722ebc5829db22578af39d6114d34d7672cf7d4ed6b58b46777
z5c1aa5bd742aadf35fef3d023845b4b6881bb1aba255b04ab84adbe19aa1942c8dc19a3bfcf663
z55fabcf5c1b3cd0a4c8642c2899f1dd84d9d8a71c80119df4975b58ba453f0b5b6ef97a8bb98df
z7174cdd62d3b652244cbef439fc0b1c1ad8381c324598a7cc5c0dbce93b1113bf9120fa2191f18
z9f9cf7376ecf71613f03b35947c8d2a56dea3e650c2461b7a3d9cb4d6a786ea9b9eb1ecd51dbf8
z31c99f093186cf5dd4ee4de965c6f6392cd255bc8010447ce4c79bdb117be608612bc6b17d8a34
zf163b680585316387926154fbc081b826bb26775452e27d1383ad3525cd389ebf6e686717798bb
z3fdd0db8caf7f487cbe05cfacbfc673069f06ee8e06fc1a5e18e411ade2c0eaf54aa32737a875e
z49b85ed8cdcb36ec6349f0f6a256cfc6cfa53f741a26c0afbc6fd44c460cfff305e5a26c5ed274
z91177ba04dc306d51da5fe2a8f47fdb7e02766d95a0f06ed4f9889efdf153bd9785d47fe1c7dba
z7877df173f86dbabff8aef51aabd2e12a6959c7f1213de4893a4e10f0887617efdcf5d8ae31d0f
z13ba0c5fb0fe1c61274990d4578d135b53127afccfc0a8a336cc1b8976e82c1599d439cfb84c5f
z6c4da7160fde776ce63bef6fc9839feb0010ba470ad724cf70d46dcc50c77e4108c9c6405516f3
z5e761432b46164bfaceb14939d880120f6e2e9bf8ffbf4715b05db21ec6e2c5f62e15f2286d58c
ze9e721e7dea33fd7f3fed9dab19be016f38ce5d7de2215f3873714dba40b93fd9a163f58f387eb
z5a1d3b131b8dda5b51a09af4b4d26bd744c08560bfb8fe97aa9f9146e936b9c884458dd1eb3d93
z045d7b549782dd56d46db7232a3a1241bbc274ec97b09404a3962d0de3feb7618ac7f9edb23e0e
z3fab3f646f258b35048b53e7afb61427c187ca31a810c27e6acfd8ede973ee63af967f07c25cfb
z08922b11cb94650feda51e48fd4b51bf4e7066086a1fb6d8ebd246fa00daa7f83b1fa2e3c4b760
zbe3f2c183ed81d9a5b8df252d976be44d7128a6096f26244ac02aa2b56c8f505f5776350ae57aa
z09475e692ec779b56652a55249b747cc871db827aa589e323041ae07ae77c7cf908f4d9dade191
zfcc7517da9fd542c4b8bf18a5f803783466b6d48233e439c49a5d7eb895edeea94d6a7e465bcaa
zc596b8a7c82e2d387e344fda47eb27c45b261c45998c9ae3011ca7399961ade9d9e8b6c1252d29
z96f1c7c5e54e68051a9c63d5f4df2fc2f28c5eaae5aa2256eb55ee58737b5f12a1d5e0469d6ab5
ze26fe21c764b1f5892d0498dbd5c099af1d277dedd7791dd098785b7f93c180659bda318e55758
z54737c21713079ccb921930a8ffdf5bf5c97506f07ec3d2abe2f69796f86bff650f76040065d0c
z31de0563581a5240da37d1b95f06a664e8f3cdf46452d0e752163eeb990585da4077e60581abb1
zd1c5d476c8a765bd8e5b71ea56ac6ceece01f490abae2542bba62f67384116fa0203fe42067c64
zc7cdfd2071263463853eba87aa85733e3ca0adfe172f8a1d272e550a780f6b48692274dbe5d36d
ze8225fde7a99ea9a6971b0eb49329c84b05e1a5171be5cc354ee2a392dc5017c1925358a8f3a5a
zf3879c0e070e979ed96d1ef732b08749296fd2bc0f36c0875bf65db271a67da6dfbeeba214b9fb
z9647b33013a2fc37dde3c53cb0dc0eb174e47cecf7a25af0904492d73bdd542a143088f5da8850
z804beedb140a474791bf81f3b3a9b5b48a67c019f9366aa9f3e01a5cbb81038411db1adb
`end_protected_0in
`else
`ifdef MODEL_TECH
`include "qvl_spi4_2_tx_monitor.mti.svp"
`endif // MODEL_TECH
`endif // encrypted_0in
