`ifdef encrypted_0in
`protected_0in
ze74c34e226135848fe16db9ffd31815111b6d7fb642c521a3f628cf6da949865580b22efd062a7
ze90adae0e65e66a2c36a587d0a790699166942afea5fb71013544a379d857e146892234d38e3a5
z4d7ba7c62fa3a65f2f4d7424646d44b510488254a74265698a7d7061e59dbec7c6ba2d153ffa62
z9bbdb6b0d94277ca46d0799fbbbfd05e5840c76a44c76bb8827cc70fd94aeade2e109c923d1800
zfabc4556bdcc931c4d75a1f77e2bdb07e4b5791f120f631958203c05da9a77d6b8e1bf6b79359a
z3867a84688be35edcfca5755f9e68eb0fd78d231d23c41965723f0fc86a46cc0ff42cfa62494d1
z800bfbea9764ab39642a354d0afb1e579af2e5c001982f2b3e975e5ba318f3a2f581ed37f38a80
zc76af5372f18fb93935913bd7c8d9c9bf519a32f6bf92658356c3f478657d5584c5e80b7684085
z74f8f041a1934a4b483461bc98df97e0e67587f1df5140642299954a9ff9286bbaccca2303e1bd
zb9a41b701250f7c71a330e5c2348325991513a035d23151d5be51498c4bbb70c0bc659dec2f66f
zf3d0679b2478484e3adfe5c5920e8823d0f93906e4991d2aee2b266fb4594e543bcac71f972650
z3bc9b677abd4e007e7e5ef3e86b183228ecf4d23a9cb90650922949608a704f2673b1efb9e289b
ze60f10cd03a5d19536c0d3f2b78249e2d85c9b7edb06bbbf0a4bb72ea6af69e181bc534e3a7c96
z545c7a3faff1e5582096bf20684132d5406f906be4fbe2d602e885f14806003956053e4f7f4676
zef9cabe44cda41d12acbd88b04b83d78c1f7deac7f9eca38fd758de0e91c9e00a89324907288af
z3cc303d9f263462ce94dee2f7868ef7a9b381a8479a4216003071bde43eb349cd2a0fbb2ca5573
z0e622674fe8ef3fcd4b8ff4caa9c5c4899ab6d4d312c7c6228dfe09527494dcc4700a689e39ef2
z0dcb2b7fd7d11ed2d4e9ff0573f496f7633186513b4384d18a1dcfe0676276af02d4d4a72dfbe9
z2e2e96c0abd728fe9f5c1608f9d4cc4fb73d3816c8a993dd712ff89a3e20b1a150d78bb7494c0f
z5ef9ce037de29eb7015ba41202ae5a5b39482d3d57bf971c9ba76d8e13f47675de0b5d627ae081
zf600ac9e102a4555ed319b6db40d8ac8e24ce6b8aec170df073fc0f17baa1a1a5e5c99ec1f18d4
zbce916d33ad0878e5093151c5e60d2c4c96b0c788885bb27bdbe5283f11bfece5459c2c90f52a3
z6a13702ab29756f2ac44983baa649784121ffe9bda0f06d639cd581e05e9ddf60129543d06fbb1
za7179f51b201903a84df17ed41d8d7e8f1e789a7296267398fb6ee01313f528fd634fd235404b6
z847372bedf7d4261d4e9928dc44861df5b4177eb3912060a78d1781b3af825bc3a3d1a43e6f7a4
z6a8041f995b092ac4d2dd52575a4dee24ea026c4b56684ad55878ece68582fb12e5619e2a0739f
z4906e0a29e1cb6b7d7e3ea3aa94f6426a118ff60d44c8872fd2cb22be7b9fcb1d0de864f01ecd8
z84dab66e9374132ad09636d10edc707722f554310723e39b8f6a8664e4ff1a96fa3185648fd9f0
z6dbb33a703abda8c0bc6ea03a014d1a96237e2da44b476298413d90de2f70068ecc020ccc428a5
z076e8de09f8185de3d04a43d3dc1d5a5b13494b0dc838eb2950a5430cd5e68630d285f18e5e8e8
zff924c02d066a197a87d3147ce8350583757edf2edb7df512b223e26ffa784d00e4d6f1043c959
z691dede21fd3d2bc0b589b90773482ec5dd52a245f0d98ea3e9478f8fa3f9daa590ad79f1b1740
z74f5a1edf4f4fd9d537d309a4dfbd94685c97a93387173f4c9b0258c3254d9ff39c558773c96a5
zade6453975f20f3e81abdf076ea11137e765b26d6b8187ae97caa5cadbd710afb9836c0fc6d37f
zc709c87e88f9b0a2223baa4909e5e25b8078417fc8ba3beac34397d7bdb704be0e171071b2ffd8
zdb201c8c862a678b2282276d65671661f199fd5c264c191311d76dfdc4f2447a815e8051e11225
zfa1e5d6686f618be153a292261a1e1c5b1d7bc184354257ce29363d564d4dc466a688bec841161
z85db370a251c1074dbd91ee30202791676e8e7f6c7d1ae9adcb1b0ad1a16b78ac5ff832769290b
ze759df72732fd690a27c9baaeff0f275cab9a3a8b0a30cb832a3e642670d5bed28e9810d7a996d
z228876bae33d7bdd2d49e5f9cd8e699b0ed19030864a4df2ecd34f1c3cef2d1e367d1be1f8bd17
z9f52decdb85f612ccb2e70cee401df0789609bd2182998b55b38fb232cf1e306a994ad70e902b1
zf9936b9715ecd1ebf665fb3bd68ccec91bea6c6762fb4dea0f2e15dd42f71f9885c19a1d1ad716
z8d6c69c29256cad1174194b330c88db32828391e9360619ccaa51591cd3d2410047aca1978e688
z91af87e99258d9bebae51218f4b271dc0d9e4211f4ea78ca29c6d7c8a057b5a882dabd14d84621
z16d78938e929afc03de915bf6a43de6ced825a20d38271bf9921077fd2856940a89299aeb2c21c
zbba77ce124b8d559c58c65935fa31b17b40126045bb88e986b36b0bf14987226e08c07efccddfe
z1ae63c693816e2660ba5c0e69196c0b0c0ec10b6069eb0c142b2b9607949f3f20c0be2437e3b24
zf77e55f5f22583a4244a637bad623ac723f0e9175a76cdd6b2c37c5208e9539f5230eef886a954
z252413e8dbc25cdf6aacea445f4cae5d54bb799490e9c76e289c12cd8d3a262eb60bdba3fad717
z1f2b6b2982fbf97223fa21fae551878fca8d8cf9d00ba62645136084af544cf44983f7ad3c5b1e
z3028bd4aa9bd5e6ea8b08d313ab47ec2b277b37b00c99649d36522d0a8c7f5f0c471f361cebeb7
z307909808b8eba926ec7869f3530b3f7333e209643487a046a4a25dd0ff377c7a55ef9fd46fa08
z46848b302d694fbab04ca0a0aea823083700742e3c92c570ba7b56255bb72a1bbce7990437c2dc
z75269b5f7e5c99dbdb89961eb1ddf708d77a8e3c1029e4faf1a409ef4dac15c4acfd18185eca4a
z2506366ed93a34a7ddf6e80e6b6c63299f3cbe15449ad06699db657a2db05d749314d1325c38b8
z1d69b68208328d6fde09a7755510d69600f942129c1bfc0a43b533cf033ccf37957882ded52c51
zfb28f096a79a560c8e715867e9c2df7c005c593567ce96fbe3b13eec62acbb67723ecbfba07df6
zdc26169ed9e49d06293c6fdba94bc654e9da2ba5a8b0b2b4e8c6e5c69832288471eb115ddd89b1
z7c1db60a1d564b955d327bf34799bf4ca31f392b375c1449dd0e1fe41245e4d0465082d04ad888
z680f3f4f7d1c29c9c6d8ae472681462eac25d8ca45646b4f26e96908c539f04d09cae3401885ca
z6fa9b6e50b335dea8f955e80b70cb6f2811f6d92b6967d60684e848bd526de26d7a6a36838b594
z5e011fd4278d5888fc1a5c4f654599d77ba7e73281a027cc076ba12acbe7a9d47fc85e71d1d4b2
z72133a2b44cf2abc985347e33bfc180b9ee439908cb74808246b1c8cc91afffb2c8e9b44633b40
z8e0aab4a89de5253212511e19f18d48316ea78328146c2bbc9f56c6637d1bcb9683ff5a1e9f2d6
ze5eb7c5b0ab4ceae03da10cc55388cc0b82052631f0b852154bbc84c4bb9f784f73b251919ef32
z44c2eff0f97ad9fbe093b94dbb4864b8fbd4f3a8fc3590d49152003371337b8ddce4473c722938
ze8a8e798f2b02734e5f40c35185c92ec25e350c93d6688c782cdaeeb632b6a49fca6112b10bee4
ze61cf030c942b6696dcc3e99bbc274062eadd0bbebeec10a7f7095f43e3b3d42f8b79cbc5edba9
z3d1e7399b01777a67edb6b1213d111823188f8955a0094ef9cde928d244f8988a6f32a27e8a9e6
z3ca08c07536db8decd0c98fd5ddab50081eca909facc02103627b98d9cca9bafa17b2ca4b0835d
z96e8d4dab93cc8e88d0268fb2e4817f967fee506c813d6891214f81f7d802bf869f5adf308216f
z5deae32ac39035c89cb7eb12f1a384c6080f247e3b60e317c4988b4356d833fc69601637f63c11
zaeb81b6b7dab688a3e71036390b3665b82f55c6739514c6bb99b2ba0e56cb85046c3fef5eff812
z9a9a97467d34426ed45780fb95ed0f15d38e5845a1a9a958aca22b57e36e40c4cdaf66203bce05
z7bb78294598d93138fc5c341d7af39ec7a93f02fcf063887fd0334e6c30c51f88a2511604224f4
zd14503368958c5ba500ea9ec68d6bec1c348689a7682fe8430913c0b82f2857cedd454df3ae2b3
zbdbec8c22d9810a37c549aa64a0bf3d1e46ec2a90bea5d5f6aecf0b9b802f0097765bc9f8e0d6e
z1509888e9c827960e9cef2e4459ffb32f6dca78c7897b39ce618a9302100d91547dfbeffb87b3c
z5dffa6a7756a89d980355156846c59fced17726adf370e0f817419cd766c6967629f2c84432498
z291fe11bac7dbf86c704eed51c45e547804cbb210cb31943a1cfb9ce32de889e2d797f5568908b
zfe0e57d9c27315b51055bd3c2ed5e592145614186105273c68b8635035dfdfcbeacf3c6a126552
ze1546ba38294972dd8adaaec79ee381e0bd4ca526898082d6d677991fcc62e277a8d55824e3e39
zad35a0e76066cb425bacee955be96eaf7af656325bbf8da0b55c07740f6bc0642c5bde73cd7b21
zed6c8660bee65fb893ca1403bb958d1488e46dc0f3893c358b7c8e9927ec42904210ce32c004b3
z6d9c85b22f1972d53e32dacbdca76b23e786456839586c7126d1905aaa7b2a1967e7216780761f
z71759b9249d9de3fbe1efaa8d9634738bebe5961ebc560f24b59627b2e7ca58c73717d21c37a19
z580033a3a78f22fb589433c6d162c39022f42676bd453b8729242f4f94766f32b6f8677bc94fc2
z901d34d3bac10bf27e48f5da43c4b73e3535137fceaca7780f5ad32a53d6573b461d9cb504fca5
zb9eb9fe1d570151232e28bb2705d8051cd2aa16fe1b6c9fbb438197968c0b02f7457398a3c72e3
zd7f7a433cef58fc50b308c3c4bf782e4e609d3c0a63da1423072a49b5c7e338c5e4e3f69e778ec
z415336ef8de82d8d5fb60cd0b62d1a60865454b3686b0b54f4cc8a0e3dde8bb6008270c161170e
zb0e4ca3c671d8df01939af1a91a6df6f63889253972050d242dd457c912ae1e4a140d2f47779d1
z7af3c6add39f1e35e99fdc5d935002bf760f44b9b1cc79602c46cd680054798e69f08f2bbe738d
zdb19c3dee1c5421dcefc6550cf5ae84b2e56e6b7e82bb9ca7a2c10d7a5300a1957adc343c6db76
z9612bbf15265da6ef64f919bc617456ed37967904e5d9c25fcccc8bd8a2fce41dd9fea3cd39668
z98b42b8418bf06715860434dfe45e00c5c1b92247722ca77fac215fc4fb1db39e1b2728a3ce916
z483ab8e8cc035ef85c626185eca5c556d4fd513badf045c652797ddcbc5da9f323c276f1863d7c
z8594f887a177aa4cb86072cbc831dd0ee75d5ada9f19c48fbeaf398b226aea5fd90db5a81f315e
z76fd83f449787edc4a7d3ea5bd8db1ebd897dfc988f3312233182e3d10beb670fcd041865fc1fb
z7623e4f01e19bbb8b1c8d41b5b5e34f217775d766aea2446d907cba74278dc9b8a4b19d569b775
zfa2f9ec59556cd6a80d87e43bef60cdebb7bd5aa72983a88ab0f748a20eb9c9e6ba8c6fabd7de6
z4d04abf49a0a6c1c8d9f9fddf4847b757d42b1e3c0170404d000e60293ea92820c324ad269ca16
z250b92a29b6ce0fb380e635eac360d08c7339fcc0972d97b8b428d799a02ca0b6c1bbdc14fb774
z0c97982c8a202779d24901b372a48e57ce9f4fd53a3c354637a9fc9353cb5cededc1c6de4c6543
z65f3ed75c69b05d74c843effd9dbdef3f1c05300b87ebe35a1aec86775ecf03a0bc9f0c5e5a699
z7f48b56558cf21f862560c74d3345b35869e63e520110a1bc3e693860f76ac89d502a743be97a8
z7b8ecbdc9be2ec374885f25a57f3a92bbb2e9a7af20ae8bb5d7572201d9aa851fb753c20944d97
zee5027708631fab81e61b7083b5758790c889f0c8fcee695de310344bff75ca9cae7fc70eeff7a
zfd0d380dd81b76fd403950d677d83242251c4c44b09a4dd3324bd2d2c3a262b3f85a0939ed67d3
z7b8c5a52a86fba02084b01b7256a34a552def46e636872a853b40eecac5eacdf1aa2227d0fa0dc
z515f40a827d901be4cf650f430add111b459877e7c7ff8f86c234f710263f04ca8ff185f457491
ze5a33f18d065f76fffb2ad059caa0f96a5be965cfd7c763ccf139e0b20ecbf88ea08a94e3e8eae
z71a3d146461e15ae279b7b01fa0ec025a1319d4e547282baa30791c77d85caf40f0352d3c65d35
z5731c18e5ff9a194f6404d3b9436abbb8e353e77f6c9bd8b42fdc31d517f7dff25c13e761d9295
z5ed1c91e5bc446c3a57fd09c824abc90d4be02dadc117fc3565cd8f03bec9138108dee50bd4f3c
zde856ee989ba0ccfa7d08e8fd1f30af380014943b48623bf2fba16f14def101992e7a0019e4bee
z5959332799ee40444f76ac3ef5e186238ee89990b69cb5f401ad5d1429c3b340150615161ede9e
z04248cb1888b4c5bf0760395286df7ebaa7c09519eb2d743379a0098f7e31a49bc7cfe1226de94
z7ed0a67518b6eae09fe0dfbb08549ae2d9e9f67c482107fcdf68170a8bd640aa9b147a272d6ae9
z81417ad74e83f2dbf5b58e2981f5378081f059354e3e085cce91105fb13e2941cd50d9726739e8
z6a27a77549b964db0329375bc4fc73ed781a89369e254748304e92e8dff2dc542722562ffbaa65
zb9e7b383b4fd19c30f089a4c3011a56ab7a938f2bcdc834d2ac7557f3e4173da3b9ca35c0b1e4e
zb45456d2d72cced18362822ab397a0d8557a05f266803322f1ee749257c8851541b530ada1f384
zdb0a2cccc23ef38a023cf6f76071f77f1d99a65c9ef39fa8d5c6ba19856228791b5affff9c2c7e
zaadcf2009ea5424ed77f102ac9adb6082184aea4262837186b0212af7ea25551048a0766b7b51e
zf2436d412a715f6f8510a07d7a7d19b0231590836ee6b21c108745872f6a614eec66244a0ef77b
z5af2e81007d2fbd38ca2c4e43acc36a958364ced475d9fd35ff4127febf6e82810847402355dd2
zff545ab27f1c24552d40320fdb4b1bfd91a0ea20e7753b234c396cb93de236c6f286564220ea74
z9712eb7112ee9cf683a87fab1662db417643f5fc04640ca8bd01f85abede67388cfc7367bf46c5
z932b8be1602f6b84615d938c1c6e7fb41c0e495bcefcd48fe576a955c8def998157bba7b9d205f
zb61ae7cf2739ace03ad6f107825e84d9ca715a7b12164f94c6e8524d7bac696d87e536767e2703
z8eb841e278dc873c7fbcb8fbd8f5a43c610a0e134645eae08b6993338987072cc7fe4f42210aac
za2de0c8e3d54e69553ee201416a58c4c6ff62914356e805882b72334e1ba1d98d555e648620fc3
z397dded5dfd45c43577f2b1bc427696afd0b6b41f34e0ff6d28b5728884b5f12c8c7a4bdfd50cd
z8787002afd6f231a9711e21359cce648a29bab5b36219f54fdbd5dadf7db5ee63dfd801ffebc20
zf855fcf0655af777e9db6c88047d3d1dd2126324f833d6bd79ac6c1ebf436fe0e7c54642fdf7ec
zeff5911b28a14bc07b0a24ec093e524d9e9d9a5ce7d8fe1a53e0903a3cf66c706b82c04a77be2e
zb622b44d25884a40559fa649a8248b029b10c24c576779f2e83a56e12f7b71ac06c86fd8efb506
z7ddd2583f5d703e62085d49ebc272fe55596e56be5930dca466ad058e08a9b1cff0f93253d220b
z9b3f76dad8a31e3358236aa2035a807f785965bd0b653b87dcb7681b0ecfcdb33d7d0a3c641be1
zb0a11e829b707bbc8964589efe376245110609fcfff6adc548bfba0e126a0c2a09d6c8c97aa1a4
z92e29c3dce75240bf226e6f937b37f707994a72000bd9871da27803e338f40502d2958acbfa9c6
z0be85979ef21a8188dd876de3c6bb59539873e1d983aae7206983d09692a5c07985e885aead4bd
z6f9550c719c3a4ebb8278ffe15e606ee5bdc83d584113230f16c9b1681148d3a3630dd060d0b1c
z5f6999fa5c861c5e0043941105dff5dbcfb765f6b6e16a2b634f2b5ede859993bebbf72caba3f3
za2728478ccae23a11063ae7918d85b9de4d6747c4ee102dc2cfbdb08010d3aaff2341087dff320
za5909b2c122db909212ab6d56bde5de0401542ad9c55b5091e902be86f586b01887f6e0d3eb302
zc22f6966dd24d294e5d25caebd290476b1a50e36ba86a48dbba3ae154c70d954e622f15a473ee0
zc049414173087988cc25002c2976ae6154385b165aa4f7e1aa2d9f33208f7414c6b4ba435969c3
za8fe0fa6a67794e797a296eb1209eb076c7a2da9f11e229c52400bd30872e386d2763489908fc5
z0516071e665f7e38596f84349220893f20783ea4a85954e466e1f61d752fc921bf37e8d5d8d926
zb760ea6494b661c0d69b360275bf38c53a03575eac1f882b6371acc08942c191faba51e912e60f
z61cc37ca5072de1e0f2147d800c3f000c096461ad662de890e728096b680b7239da398597127cd
z4397f84ce26db2124c91db8913880b37f078e5dc77b4e98411a9fca035edc5438d5e3707b61e07
zabd7be14032c3f4de8c1ce9f90dfe226c48f65a06e6c292be92d8104a6eb4e405f82af6aa18f5f
z774cc695577c7037012731c022613f36a883c91a8ee13d50f82660032e66077a8196c0c25f5ac5
zac7d3fca82a8c44817abdf0a4d49496c00431a7e7ce4d2f9145f499612cdb0bb72fae242ca03b5
z11231f266125007af035c7483c4a08cfce84978af9fb0c3b2508d3b2fe178753e3024270237c6d
z45d619c9538bf6e1811fb5420bae5219699f128bd1e4bae14346057c62c1b29d8ece0848fabd88
z7bc9f0ad180c1e49799ff186578057967adb400243c75dbda2ae4156b0c45938a29b047474b4ce
z3f86313db03cd193cac682e1d3858f4519ceb155a5ab9c0855f7bb27b02bf1a241c9bd89f98ee7
z3a35030f105e83e304d0c8ae44e0f0b713406bf10575ea12cc3955a73ac9131915df3151dc35d6
z332c2d7609f85301e1cf5f3e11e878262e00677cb02769d45062e8c64521c8e3effd345b5ec018
ze2c624967f8ce355957e1cbcd6a5534c0c277b17f08be95747d78fed644c06135d26a90172fb1e
zbf996cb53e6854776600c5d8cd76f3780474ca30bbb67008debcf3b42322e6c2afccca4827d4f6
z39249a76fd0e88c633f6296d8bd19c878f1cd2e4634d30d33b5424c730604623e8ae4557482e89
z4eb77949ac4fc50f8e9eb499734a4dd5aeb5d45ca6282409d4b3c1594a2293b2926df59a61b714
z1e6552829f665d930332d2b0c59f5a68dd5df8925e6eb7f1af7a86a0affe29961560f02b300211
ze1496c2566a0798cfba536335cef84b8b94f0facba1b108e018a87f30d7c250ebb935cb3423ef9
zdd6f8adc95e8b31b91cf974b9f87b59d6d632282c1c2736508db41f2d7d619d4c93b88c430db4e
zd0233b15c7534441aa4c2974089d3818e907065e1014dc47c9bde571e2a36858f7ae8b92f0bf5c
z8c31e537373f70932217ecac31bfc2e26b362eafaaba0c1c3291e212b5a842fa813facac9aa853
z1413fd2aaed8ee4f4632a6168cce693a02d760d4c5ee6c667dbdd3a1ea1bf2d9183aa9045e2042
z0c2e470803cada2ae5572ee367dbb0a2cab945848a34a14c7a43e7611452ac903a97802698b079
zdf68b06452773dc9a69d20074f4dfb348c8fae884bfab660492d9ca4b80bad3b4952bad5e3ab29
z6583b11c22826edc14bf83e3c8e9f66ee1e0a152e453c71b5bc256767f7299cabfbe84dbe49818
z5d81d1b38188f1e09d1989fb90766e58e9627eef038c02ee3d37083f68e2406c39847db860d2b1
z102ba04b29605cf4ec2efa49aa231e6c1d01b81fdc86ed1596c83b585764de91e669493fa2d560
za39548f72d25a5a7c9f426e5056d7491b72b845e915b54c018490bc2c6fbb4652f9305232c41af
z572339c1ae2172d5da3acc6180cbabd4818d1129fffc350f44a91eff4b9d0bc549d831052d1c20
z41f7e22edb274cb6b890097db8d6688c9b1e85e75a99bfbab9ce61b9f8702d7987cd746e401280
zebe967c5b365980eee042dc6e48302883bbb56af9c49f69b1f1a8ad43afd7bab1898f770cf7030
ze3b95954c3b4da586d2b42aeee2859b7d57f0b3158a44020a81b1685639809fda6c0aef1bcc32c
z71403252704500c47d9009c2925454f9eb5a7c87d99161498c9ab403f2559368b3f66f348615d1
zf6fb47331640818437854c26c8e8fcf47b891afba0fc09138bd2b97c1bd9f65c5892c1aad32fea
z7303c3399330ceac4b0cf45bce07f009230e2f45bb51e94b73bfc90cfaebcd833c0bbb03898bbb
z18d6f4324d6f161ae1026e2db1b073ec9c636ff48f281efc075504458bbf6b63c9550099d1baeb
zfaa078bad2056abb8d77fb3181bf32a086cfcd14df4c795fcd68effecfab56de287a10d06ba57a
z495f517bc52ec6aa8e4ba8eabf02812ae6a0bd2d2b70ad41cbc7ba4f2c07e1e66f04e04ce72928
z39d1a0c5768a20736cd20a16b84e5cdb0b41e9efe81b2fcb70b83b6e75b0d2c46803343bdfdc15
z73281f80d27e1601a3c6e808d36a53ad0b1aa1f93f469e06ed560e29d21887edeb2eaa12cb1db6
z8606489f5edba17737ed39b4698159e3d3f426ecdb9eb6536f76af27d77933bb0278e2e87c3544
z50369f7cbc3f7f781bcd6112780f621f060e7c985563946dc734561e8aa1efd3e5ab6cd9a18983
z1419079f3b99102cb2f4ca1c84dcd6a8a67e96559261d3f3698fb3c89d7168a606fd9fd4639e1b
z36943aa69619be38613e427afcb2d15e0a482ef3e2fbbd184801073f549752bb96907f952eb295
zfc468485d5f8bcf87bc75324361bfde898d7dfc83eeab8d7b1e7eb573ed8b394715559b9be1c95
z11de1dfc67ee1c15aea2a949fdab849f4b7dd7451f75fc37b5e16ef2775215df0d2916f1338422
zbe68d8b945de459f56a2bab6d785952246615734db1b7327fff6921a9dd45234d8af3f2fa0160f
ze0e876764c4db44d881456888ac64303951ef41d0aa121395aed67a49fc11f75459ba137c3cb8e
zda08e6d6bb9dc5d6a122d6f93e40d643e3c1e318bdd2cd54dd6410944f37b47f8a0b9354feb2d6
za5caacee69c3a9824f58a1196c23818021be3025fb35b0c1f2b8fbc8db467d9acbba71a5517ae7
z1f2ddc31f1ae8bbf2bfc6ca2a572d9475e102fd8ef8c759058790fd82c40baaa4abf4f41a391e3
z0f04574d20f267417665421de982349e2baf997912bce190fbf9566a8af1efd155b5bc22c2d572
zcd62a528ba723bf4ffa0fe40ce0ad75dc557aabb47d354bcd4f149b1ee4904d04fe5d5946ce9d1
z617904e4ee492fde3374baa352668c8563d9517198fe03157f576a0d7138a1caf8847dcc306820
zc6014ea1185f18706b2391ab3caa1bf96d760a61ccd4e074fc7504c2858f97d808a31f3c225fc9
z05d40a1c9934b6d72a2ee723e56848d768e1e9fb59ccea408613cace1c9f44d0138e8a5b65cbf2
z92f91f3491a72f8af33b6a5bd606a5d912d7be71a5f909b1f93174e7de2e463867b82403dbcb74
z9c9987759f57fe1f22aec07213249baa931daf6a7105ea7aada3c884124d705ba361f496766e36
z7af3fa3f970283b4cd904ff2a99a65881dbe1115432fc90e42fd343eb0e21784c5ba450e137a81
z9de0c523eeb73be1d67a887ed5dbe489ed60c0643ea3e6d1d1c17279788379db7807f452896847
z308b9c053fcfe461c660fc485fef7ea40b8cd87f12e44cf595a5722103062e0d75e3454bca8d44
z2fcd571ad3ceb4cd2fff7614b47c58cb088e6227a2e3810087f97c389cc55fb224bdb19ad84f1f
z9f331fe65eca945df10dd6824d946e421d4ff84ea3ad9643f5a9ef3d306e0561873421b9a48aaa
z1acc586280f9299f58368c8dfdd7af86dd00d29950e9a602c06944684df371c2d728085e63d0d7
z9bd6ba3be483cfd76b068572681a01ab35d1642386d75aad10caef275c78d275f956bc458624b8
z4b4df7f6b947925adbe16762fbfd030f5f863b0d1c3041e9e2d93bf11f0d71ce469de0225822b3
z3f8a374fdb958fe05e508ce2b2544b0402a0d57c82f5fdfaa242ad0497928d9694ddf0764d636b
z34aee32aa1c2cf15dcc0a82892e849cbe2abcc03ae2d5c0c0f92cc5180cf85322994761795d5fb
zef00b14d33b3ebe66e8a0966bfda6d5c86cc9411b39e22ee95275a7a7322292eb16473d7cdcee4
zb17e082bf9fc7bfa40897aff49728d60c22ec89d9d5c31dc2bfc8ebf42b53f7d9e447f22276307
zf0941b38e15b893f6aa11909f9b97dfde7fae4f3676f02421397efe54a634c7cc99e6478203dbe
z902ff4cce292195b3f3f47c70d312be1a23b6bacdb31c86b783a7713301e976bae78fac3661c3a
zbc775418d5f47a74bc169156aa0cc5fac6e381789cc78ae6702251ab2eec27afd90eb484be0903
zaa901ed425285279be48a494836b23eff6f56dbda89c5d0f110cd86b0cb6fe54aaafcfc2dbc3a7
z0ceb6207cec3c918c158ea83aaace5e4fe2177ea58340e0ffadd28faca9d60121fbe9606acb929
zbfd489a0d60eaad334db3233b3378a475f44aa15685544564d5e3cb3ec3d9507fceebb97a48df6
z1b5b44585ced103f6b46720285dab2dea9a65b131b28d71dfc3860b38903788168db28d9d48a35
z8d9ea1cce0e2196cec91bc64fcce52a1f7a94f3c0cfe954e9e4b13faaeb0823f1bb4500b1ffcf7
zeb542e0ddb26a708cc3a429cbefcd9b24f8a930527389b6e677718864f0b9700a3900f852d07a9
z6e07941eccedb56cc32c0c19f8a90e64ea12b12be6602eb1d4a6a48ccb40ec2fec82772811c906
ze0655241cebb832f4c480b1ae30cc4144e1b033106f1b3654aac0afd12077228d53392d2600b2a
z54aa8105de1d8fadac403c245529aad0ac7d5270ea0e136442349ae92dd67e25139e1d7e55d145
zccbf6c2b8cae632229051d0acc20730ab286b9a153d9f026f123b72591197e9bc7709756794065
z8dbdd7b01607014da60f0333439aa40ee4f89039b474b7a133c870b0082cfb1c0d305a958293f9
z54748700b4797ecd0ffe383806a4c71b8d220de3b6ca24c07dc317ea873b01f68a143aa73d2a91
z1f89c6d9e41767f4aa2d86f4ed9fa2c2f320d4b5fc00902ceb5d074e623322084cd317a7bfc873
z463d4863f341f987e659c3af0dedc8ba2dd48f9bdedec6934e7dddc1e6dd7dbc63b75cfc55de6e
z6b4b71ea6d0fd9152a9c63a6dc21d3450826e22a2b9810726d6bf60f8792d9c5a8c44f4e499b7e
zfaac6b21cbf259850fe87e343109bf72b03c88b9330135adcf88bb1ac28cc877e28163ea71b8ce
z5e3320e80c20d071bdcf9212272b4ba834fe2862a7734a0e0b53f3b16bb9eba92798371772490d
zb04a1e3e878eebc38ec22b59420686354551c682e81e3c1995ff2b36ba96339c4a1a60f46e7bd3
zbf02dfe69585b6288d222d5fec5339e5082f23faf4c33adf745520045e46df088ac134bc027517
z0bc7268aee471e36d9448ed0d6f989ccfb94eb25ec70a24bfac78211f064b97f6f7fe271d76df8
zdd97b42e27e296556f64102aa24d739941fb2cc599b66aa13bbaffbf597d2d1ae9897144288fe8
z151c30e8a7ba03e9b99ce73537306fcc33bd1ec30bb5aa470495e2f73f7f170c16166a1b07a1bb
z6c5dbc55d578401fc5a205a3eb2c1b941be92c941adfe8f690751b5e2cceb457554232cd46ccbf
zbe123f011b7534167baf96b296c28e2f844c59999065dbb5890645bd0fc52c70893dcee46bc2b6
zc0aec9345fa0d2dd3a251462773e8f51c2f99481ac39186863b6254fb5d04d5c95aa62418f5554
zf67263610e8905286b8089287432d09dd271ff97bdd6fe0e256e81316b43931cfdeda309ef5b11
zecc126e0f81792eff1931d9b6ccf7ad782d2bab8d893477d9e46416606169b4558a0741aa02c31
zbecf20fc16b49e831c90d7358555f39f6e78b351186148975cad9576adb88a649108f1ba05d55c
z5cf9ea56adc07bfff392abac5663837e1d795e075c43c8d146198c7756a2f5aca3d1abc76fe57b
z06ca4d0d652c380d5d1439fa6edd9d15d42dce2f11beede0d1e712b61ce6101655a9cb3ec9cd9b
zaece8396de087f8993b85e77cce4cb63e1d1339b8d1f3283e832df0f25a0862c3451be5d8307e6
z397cbd840150b140e6c344fdc44679e79324276a1636a44fb4f6acf4eb86637b76041aa40e809f
zf18b6a26eb01527d9f5cf00599f3be0379f75f253a1637f2d90a28a8222dd17cf66f2c0c562756
z7361b0f8c74841e29e4a67d937ed117ab7bb67a537cc4d2d2fe37058dc2d14d81ce3954647333b
z6e6bb956ce813663ec41e949003e86c6c3bc846f823d497bde7309bd2cbc836fa74d61b6e83ef7
zac587268a2616c87e0ad9cce42b6641bfa389c267e2d54ba233392e1a1cab4f16143b807e991ec
z1c2bda6de9f1e3a13161aa99e8a024abf278456b084622874e8913f7c36da470e2d73c5c4eec49
z9cfae845f042af4ac404b7b0a428e56ea970f32b46814302099e38cb89332debb2cf08c9150f34
z6ba30493efe6b16b4d2858a067057fce6dccaee92539e3afc886c5fd07ededc00a39abac18b7c2
zb16259d635b5fc38caf331e9a06bd6e5800c0e69ff7ca5add6cbde49b87c93635a6db059c6edcc
z7bd7cd54894c29accc6b905215e0ec5c0883f49c10ae0e4a9b3338ed8d3ff00e271e6496fbc321
zcffafeb27c7a8bbf5f0d4a6956e2d0fec8333479f8ffaa6d4d11518b747ad114a5bcb43d6b269d
z2d71cec351c56cc652f277307810d346e07f01cd419380502c1953a74653207e6a8bd3e63517d2
z5536757658f148ad48663ed4e2c1ab7df2309d5155af60d5af059ae6dcfe6e4ba92df0318e3fd8
z3dae24b017b52e4e1db370e6d68c5e486fc5e07d5e663d65ca79b69ea782c84f35243ee1c509f1
z911c3b4ffb5fbf5e57e8d9717c1a8f445aff8eba3b6f550129b028c21cb2d0e907a1727f6354ea
z7eb5fc8a830f936bf1141811f00ce5de4dec64219570738acae8e5c9a269f4154e8e42a2c3e84b
z406659ad6df20e36f4d6298293b71dc83dd7904cbc82c61284627275593f51e21d78d464f3ed50
z41ea03893ebe652b195e2c4a96df9298b0aa773d019393543596dcb6a6f5d23b3329d3b00bf8eb
z1f163fb4f4f86acec17c816bb2b362682d65349e1cb5ea07323cf20dbe8e9846704b881c6823de
zea6f435d7c834f3f0c57d6bac886afec9e248e47cf693d8fa77111f1b55269fde835810f7d9840
ze1791f5972f86bd976878db8086aef9a31e1ad7fcfbc420928724b65d04be9e9f9c4627028b84e
z253f3f5f0e41e396a76f795e1548a2d61b2ea9c9c686cd493dcbd8d63356532a0728e5f4ebf13d
z8699f02864d0a44a7300b36ec06ddb002d52e17bd8cb30281b91b69dd272484b7f8e1543ec9b63
zad349df7a291b1d2dc060bf7fe9f7439b7c314275b2c71a802afc1222d9ae8bad2c8cc1ec84a7b
zb6a7cdffde42445fdbcbe210cbb0a66f344ed123c0ba8d81d25070fa3eb52d2382e2185d709517
zbeb7fc2c0868dac7192c22d1c3ab6d6394c16f2e3fd9a4cdeebc242808b378febe06342952ad33
z280f54f345afe9e847cba160dd8e5bba0c868d7bfd9430a59e5e87dc34f4e8de8bff00307d71c8
z9b4fd23e6968033f4113615fe32d91eebe497eb919e7704be04100a8e3e62a5bbb1f74f020b6bb
z364a219da1b0ba5ea7742ed6af83eb607d9bbe56000721cc8a844ecaa6726609ed3e02a2501273
zf41971e9d78b263df642417fc8d241019d5831bce2a3edf7de161b2ebe3da8bd6ffb1b96f48faa
z84950b867cc54a5af2ec95768dcb5442584cb632e078e56564e5a8260ed3d38d42303bdf50ffda
z4e77bb9b9fa8500bb2503ad09a07c6ae9abce344047364ed77fffb366631c79c6646e435a5bfe3
z3daa2b217831775840ce638140d4f9393f8a62d8164db19c1aaa460de124a722e9f89c4c837923
z24db09e07a5967b4c46748ebc2c890a8d971e6b8456a0a0ae4761186cc31ce284c4d8a8c84e0e8
z7fc241e5ffc227c6ee0433ceb4e8902dd463a9e6e94963cc401461fa2392b6741e2d1edf45150e
zfe6d7c2447f58c996dd60ae5f20b9164e7d5a21fed8e2ae342c426a426a5ed584c4c750f82a7f4
z714e3947b5ea0489024d0b7691bbdb2ff4d188def7dbb1c5f46e831dbc6be0f467083ac7d7bcc6
zf7fce4b34bb50a1fc70b66b1a6a281534e3ff8c715c8b766df4985911c6956d8aa645d6e684fc6
z99c51493cfdd59571f23679bab032af22b55b81cea12a729897dd6931031278950dd363a938c34
z09c895e73cfd94f01d404db0bb6b0576a4bb9dcff572c607370e16e140946989dc0eebe5bfd325
ze60022b5e15832f7b0835c18b159aa0cfacd2b4c8bb01cfdf6aca06fa5673f27256a80800b678d
ze7f8243c484dc0b8771feb2c7868b4576fe79fd95b6a30de8ba9b1f451d841e9e8e2e907de99c8
z734c06676a765987e62df036ef77e61d1856e99db20f40a3602f8b31e26719c9876b2d2915e260
zcea789ab1b9c32653b8dd698f80b406b8c41e28ff2d5125b7798ab408bd74b581849f88c2cb2f2
zef19bbe1cdd2e1ee487b069414051021448e30c0a335ee9b5f517eed9be9f83fc52af8c4bbe512
z15faa3052a62e7ff490751d8bd2d37c2a5f15d696c386ee104b44f2e026d7bb41ef1d68e1aec8e
z547504c9966dfb4afe1aba5120c2ef2c93d8b4c8c3cabd1e92991b128c243b021ffe45a6d55c23
za8f97faf276316000c64e0f0d4ff0bc08ef272a9c52eee3165e7757bbb188bb4e9e9487e9d0b2d
zd93f6b6fbbdc6c2c0b79d3dfdab012e295a3cc7584f02be5c02d34674696f5a968b546888f0ff1
z1c1f4e28442e7848742a2183abf0b45632f4585dde755b6dd01e951f8e84e1c5b38ec901be1ee4
za4b53111b4ee9ec0d817333717e9dade3557caa914ba69299557bed9cd90b71cb06e411dd3ecaa
z6d351d0220c11fcc3925ed26a15f17477f36c2fc3c188081b92c8ab6dcccae6a9654046e7f03a0
z35e2b4c03f3aa7f003b12184d5dc2d4eeb0b7e5b0dc183058dad9d95a892e499680ed4a6c5e8e3
zc8bf433b3a3c21b8e0a45865862cf4f89dccc4d23cec54862b5e4a048a060398a2e7517a874fe1
z11c4d84efc0d51589500095dbdf264bf2e2e8a4a66771651e651d6369ff30a8bd87d0d3558bf1a
z433489b53f9fa0a9d70191c6ee46e6ec30d1a1f56993de08830df99c3ffbf81545a332cd2d345c
zcbfaaec3aeb44538c07c961650db388623602c2fac4b14468e7c7f1b4a767bc644cacf0619794a
z514acd8dac4dafb4cb79eb628ae2ea3834c2e0f4e909f6641e4a3292d05c140d1d95e5c4ef33f4
z78541a0d1ade2dd71ee3f1e2cc107f5f21fb5e3cfd9452acae11b39baacc29339d59111e391a40
zad9fc5ffda7e4e313fd0bfc24dc2bd5a69afddc4f701e93bb10ccfe49eb4426a6f96751012e681
z58b664c7a68a5519dbfcbd911569c7106debbbb103409373a8000231de72e20ea8a6b631b47478
zbb5bc646cb03d844be3594a26c9d417f6b672eaf6767389cbb5cea70156d942072654ab4bda590
z7a025e84882cf627d35812c95e3a1f7891bc32a4cc069cbdd0b81229fd90b45039c0739f8eb899
zd407703b5f901ebdd2b50f79a52847dc740f20d3d9479dd687bd6bcb1bf55dfc471ec98ba00a11
zb5824158b9381316662a45bc88a03b34bf7e6eeffddd1e488fe811bd35f9145860badb0c8c5b2b
zeea79b396b69d213a45212636050f9d3477fe0bcb5fac4f7a4901d607f8455121cbadabfbb276c
zdc69a29020971fc95c479550dbbd0117d527fb6cf612960b9f92690a90be92c44ebc0f13a8fdd4
z93d9081129c18b6020af7284a934e816b582e13628f15759268a633d5f985b3229c418089024cb
z5fc3f54397da2a74d07fb35a563e1fe2a2331fbdae5ca7a431f0f0c26abf9cc3db8ce81528ef0a
zac1a156fff405c847daaee101bcdfd420849e93d2a5a761e1dc14e3d7a635b9ec458679d4c5ac5
zb85259a8e48beb962c864f672b4f778e9ae71e9194e9aa8a0d39fc59b375cce9e187e0bd2daa33
zbb7ddbd6e3a2bce0966a099ade63f78331d6ec83353714257f3285e157abd34060ab0dfeed56d0
z45f0956982550f9ca441f89dfdd07c5c8e613f802c04e6d1a9e3cdf7009b051910c9207d3fb078
z87a024b8558d034aa34733b09b4ed26093c937ca54ffd96de18fc13652231bfa8c242e81edfe86
z98d68c34d2b36fa056cb1220df87cd186a71a512da16df2da160673a115bdbe5fdba1df5507624
zcf10677a75e64f61bd7a3e658270b43d8003ef54550865f33a478b1d45654f1a5796dba3a2accd
z4676f55b562bca3fd823bb9092d47dfdab3e0f6179f7218f1ceebd255636664f19843250d6e49e
z12fef0a8867d0eeea430f070ebd39688075c30a7fec6546065c6caa770ac0843f99b0010294885
z15ce1e04dc17e45b01d25d313a9c191b6e56cef9f12fbb2b18b32791f992782b21b5b6f4e79cd2
z5373659b0ab306c4162ea02f11d29d53ad393c0b5feae90fe0fb45ca0f43938b8254c358d10725
z91c51977de4560df6f4bfa37f6821db7829755e005cebdf19b2085ade49f71b52f34994e7d1dfd
zf690345c694c94be20dfcfe75ab4566b1befa1e1530b13cec0860493e1de8c1fb59c868e330355
zd6caf6a9be33ae0402f5c6f998d0ce586355e4a4b46b244c65b3e7217f5096fc9b34402abfcb63
zacd1f905e1c1bf5dc22e9799b6904c85f1d17defc4088f1395b16ea98f41ae63f9d1fb81c3a4d8
zc53ce0a895cc09fd9e5079230ea401fc9a8a7b2ba4008bfc11a9c4dfff95c4b3b01317090e8ab3
z973e8b63bcf6fc0280aa396332dd3cdefa080c56bf7173e11bcf7edaa6f0a4508ec42ec1d3db44
z339c1e8fac02efebd3de5a5a8fcdf7b5b3ceef5a9f31b8ad6952237f5f2d27d4c7a33e3936b47d
z094cc29ec3a40403d2abef9b064cd2fe6238f96e9e4de50b34c98b37419b274b0afb01641bd986
z3497e0b2f11f7ec1ee980695204bad1729d03a9a08d6c8769121d3f06e49c9c4310b574dba6de3
zd8f7c36745785184a6f66c08803de773d4fffddba4546c959f3880e9a414d5c52f5b58a0522259
z49c7ec515b483caf1239301a017b36ba5f0decfbdc29bc798d0a0aebfbd915e2c06e3271e6124b
z34be24dcd2b332ff9282b8fd14932a06439eb4b3814e407aae38318ee21de7f11f9868bc6d7336
z5a1460d9179fe5e284581f98dcdf38140d51040666e4e6550e006e5e52c2d90083cac4227e4ce4
zbc9a493c9d643a0a6648346cdde82ed00ad3bcc747818c0cfd5fed590084582b1a7eb46fd2f048
zf038f2367f31bfd91da9763367310710554a156162c0f39187dcfbcd1eda7a8b4bd349c3142f20
z232f374931995722c96cb10cbea02f264675fc3b337dc4ac04cb0a43de63a13e5528252ed17911
zdeaeefeb9b7ed57054463c7214421a381171c5ec232e10a06e4ccea61b42e9908d6cab7c17a692
z003ea95dfdeff4510e58c0ef581d12019ad525182c8fcd32a095967f487707b3777878a461b3c6
z986226ba17719a893c9734e943f0cc0169f418e03e385aa56cb563a81fda8f84d562ef962befc6
z2fd4ccd66feac07fc546aac06af0ba5862899f31bd536461f522fae5cf79b64b5229c22ceb3b2a
z716bbdc9081729fdd8b5be8f93859f50dbc671833f6ad08fa4c4ce5269b5d39dc78d15f89e1b74
zb3b635682a1b3c665aa4c6ed760778c23e0cfea672bd6d6d5997baee42f1407fef7ed7fbb9621c
z559c2e471a6a762b39f1cbc691fd440fb0033136000918a9b6cc5cab8686577b89f0cc182b450e
z4331bfae762ba50ba00be341076f60e38c150876a9a0e89e2b53c0ab161a57014adfc4d294ced4
z355b44e518b81e7b0cf7634ef30d5f09e19c4b431bcdb3647d8e1db4447a4405e6a1f47e8b5dc0
z10fbb410f8e1b0fc2ca935c646bb1228081b8cdbb42ecdfb195dd19cd4c7be28db91c34832d77e
z75298b6d881da46913e514bd7dbafeb27083c3e8f94e8bce6ffa623b73ea68a7d20becab022579
z65d98404c32f9de7884df5ea3bde7237ac0930d8eb414b9fe62a4f114dbc3d8b38b3f97fea4df7
zc5b41c7b3e8ac84c1f5bba0064e964bd982bc012d202db1546f39e2e05923f2c575a89262b5b68
zd1c1a3b026218d93708e333fc7397981ec27031f7117124e4a2e4712c38d5d4d5c4fcbf7ee3b18
z7b74c7128d73f796e0b289b639817305f066de504279ae7649b01fb0a7c0d35a3c561f1620f3ad
z558fcab16feb5518c1f8ffd8a2356074327ecab5e0a908581ab8230464c65fc1a2e0c938775f0c
z30c5ba02dbd887f15525097b73296c5af69627a896ca81d506da3f4b04ba0a650cbbd559aa28a5
z83c88ee47b5338e9dc38fd95b1ff1c8aab93f790ecb18613ec955f5da8819e605958c49ea277ba
z24e251239e3867355f61bc2fc252027160737ddb90553d81aee12e3f74b77f1992ff49b02f43d2
z9704e2d5478f6d898fe8e72bf6e35a231df79b3caeb1a557ad690ce1b5dcf234b3c50d5538a5db
zaf74ca3498e1bdebd35015dfb3185f30c299e9e9988b1a32f10448b6d2cb46afef909d98f625ec
z27b943d9df3637fac0a1e75eafb89d0eb428fb9c78ac51173c0b9f6bd252d01a7d1f5f7736e1a6
z9edad341432793f9960fcb145810061fe8b5d9a07310c568ad0ab48b2b869608bbde642376feeb
z801131a4e77ececa1f51c846811c3d9a3de39e5faae8a72a896b88fe207021f7414cff5957f9ad
zdb6166223c99fdbbcf4d0de0ce91bc183a3ec5c249423fd0b6514bddeb2dc5c3263ea5cbf823c2
zf62a33df46e4048e95f2c8e74a68a3a9918373ff6979ccec1162274b607ad8a790677858b53a26
za2826db236fc0c9ef7781c5c56a44304842cdb1c930bd0a196106ea064ba22cbc1306b40768851
z676f0ee5b2a63215f52c9b8b07a8e1ff12d06dee0febb2a38939f1150f1489a501a0e359e9b358
z634e3c5deb7d9cc78476e3e6a13fe4c8a9afccdaedab21bddc000d9ce319b4618618e28f56761a
z4e007157cfba9fc56b3f8a8d330dfc181c83dbd3ef5bf5acdad68d830dde58de4592d0ae182d89
z853b6f3107911bfbd08981c2eff643b74bedf18d4f9fb0a2e205feff15ef9d227bb517e4e3d777
ze75dbb3ec4bedd309c4c1b777110f434bbd3f14b68c84f7f74c164eae764fd349df9ca87146099
ze0f29d4a895d2ae0460474aa8294618e2eca8beeda3527ac971f0b41e5ef9e9489b26c6a46612b
ze8646c2e5612796df78fee7b02e47996878d3555453288341a36bfc6dc564a877b84017c889b24
z2b9b2e1ea934e2214b19247804e15f7eabc62fd26641eca98e51a0f3ad90ed9b6cd2aae75f5995
zbc956a1f37ba1d88301d2809e67b19859f046d6689a112426a2f1dcd0f40648f30f5e34f136e46
zaf2df847d4e94aef8fa72956e8e9b52d4e2de1d949d113afff4178d3f8ad28c04d92c810219df7
zacea2f69d70d2984e361122b54dc74d6847c384d3653c6773e86426038b9bfbfb4d967e60f4743
z634a36259d2aad5f15d8f97e1ffb41cae6467bcf4a2caa95e9a52f3bbf8bd554f2b6c2e87782d6
zdfe302f2fc085706f0c61269a05d832c2b219878461f0e92c869091bb06484a7530100ce4f9579
z2d49dd3c288fd186eefad0b175631b0e1246c37d6c791a920c46b288db312885d77828c748e827
z4a4b27e6323030717537c8ef6e4fa5e061f8cefaac027520af8f6427ec8aa8b71c6f1f907a4d09
z26e8f6ef721f31728cff6a59be547140631adb5925397148b693d5e1c51b0fac61a31e35342def
ze78bcc7a8ad032226c59a6ff43bb4d55fbbe1c82e23a7c5268a2e597999420fa0dbcd65b0798b7
zeed67798a66f31a10a95f89c1f1894ce9762cf3bf5a2f63151d5cb5b6220a9101351263e6bcad7
z851f9470cebda5b4574824ff7013915aeb73a72c5b894f8ffad8d6ea1bc45d06b64afcd8c2f006
z628e5302399636c6ee43b118c202ddc8cd045db02d3ca0bc61b2918467b2361775f5537e5e47ff
z97683eb150f677f3e97d41a9bf5b21fbbe7c0d1f8e32b87fe43baed73dccbd19cb8115bee79fdb
z70d1afae6eb7722b43fb3e985d6cb3dd1dae37294fef84a559ea91d77b0014e3048d44ead91e3f
z5432dd74351708ac2d5ee4a79574026c23a65b54a24a458bdd19380832f6c326ec6a627afefd3f
z7d98759c175b9087c31928084b0523971074681f72c8248be44dcd4d5c366615fbfc46ca4f5740
zfb257f8b6853051abe3b1fb1d965ec86bc04f2633cec06861c95938fa394b1f239292c65be1010
z296f150a9755f9db2464637a21b7d82a286ec10e9edb6bf7cd5c651102f403e45a6535be206d6e
z698ff98b12eab538db9ae5edb15bf10b401cc0dc2a511d17dc85ff0cf7b63a6864857b887b0b47
zec348083f790bb5234b555c5ebbb167e50ef45a278f1684df5eddfdaa21cd81e914ad179c4fc73
zaa15f417c25389f18c58c2d4fb36554f42c1e156f87defe788883d8200a220915d73d45d308853
z7012c37fb069e9db168f83854d36f06b8ed3133aa357e8d1c06dfada6342fdd4ed67346aa73a07
z7def59f1572e1f82005d19be4ed5070e410315bfe2734f2f8486908e40ff2d0574aca932cb258b
z14a204d1c0a8e52cb4593bcf24f3e9b1ed4cd529adcb24697589132a774529dab6d74b4d7e152a
z5589bebd8ed2b58614d833023c907363b87a735b585cc90b1a8a3893c893fe9bd8c17ca8456e45
z3f36226106f7a258621a7b371b27d87abeb65fea86f0bbfee34efcf46f4cbefb2dd24c6abc6e8b
zaf5ff6119a14a14a8d151c163f4bd1d54fa86362a1767fc877c9721bdbdde68fd80ff6deaeb9a9
z1208184c63b408101d778db033d7dd186e39a0b904b3a50676a0bb849d009582c42db58b84b109
ze015434e6763b34ddf9404bdf3d98c05d9034ab8f9e462bfaf3a270c10afe540d2591bada4fab4
z14c82d617d326deed2bb942e5f0d58bfc33b288f3e18123e32f623971b0ba7a85974cb6fac7b14
zfe9d6a2b648f42011c8b4606ab17dbcd0b8d68d04cb04165c6dfdc9dc330dbe303c135ebb132a7
z4e2d72301247b335158d3d223d52fdc31c995a03b29afe6edd8454f1f05b6488a4e6f74c2dc72d
zb27762b236f92d35fa6c70805ae2634b852088475c876131ae37220e50108c76d7f6d122fedaf4
zf7337eef18c128082e876abed6327a42b186c6e2ed0be1add79fd043ef876e1f498e9ce4bea7a3
zb0ef0c06dfc412cf0f4f8f8bfeda255eab6a5fe67fa48aaa8d431f369aca280b8a517210e6f826
zc9f74afc47bac97b24d003dc92c3dccd8b1df59306c8bbc52571abf853e30ce5fb0e3598a35e90
z23a6b36bb6b6d27f81e1569bcac5e6aa7a60ca010a44e5756b42642b2ee5d6e79f4ac35275cd80
zb69199b95ce937a32f2c5750eb88b405a799310af2b3f917d99aa49ee182279d77cc2653ff6f0f
z9a0dd8a96b287eed18320edcdf25bf4169b878efcc85e383d59100cf54dd9bf18f0b3d847a921d
z78d204fae2154fc62d086833331980a9633fb4b3593e4790868229808fc6feaab854f5ed5f93d5
ze4cb16824e5b869d78123651c4ff0f2a849a6b34378a6efa5147f768ecda91c001e23cbb4c1367
z1ac98c7e34c1428feaf45dbde58ff08a2ff474e15b46b15c1b77e2186391bf71f7ddd537eba739
z7667efe5fcf8975a90c7d72f1da979492351a10c1dcb712251e39990645c6d65a6f828ab7f974c
ze8688daf7f2794368c024915914c95dc62cb71403117717b2c1240c0eeaccb112539decb3eedaa
z6cc2784028ec3406263f8b0f22dba727b20b34c679ecffad234a5eec88ecd28f512de80c3fe1cc
zce08852f18f99fefba9d6bc8b00a7f330ef97837564388bb94432b45161644a06bac2720601ee4
z745218849ae22ead679f28ee2ae514ae432048554cdab539f35db8e7c8db3c16f553c84500edf6
z9982e311402c870837be3a0b779ba365c0bf8fcb5f1dd829f80adcc85777e64e56c4c854e44136
z88244e8d119d954cc4dc0caf813c39716625ca18b9926ac50e5c0692a3fb6531437a65002d59e0
z838efdde5547bf3c7d708329ec229e49281a742ed32a2ee3b0ae9d55d0ea0efae338860c937ad6
z675d8b1dd9656ed7f395bd6aede8c382ebb6f666432d394b628e155ce82383b1ee6a03c2da2199
z5a3a4a4b987c51bd88320550b5b80be9bb65c0e69a9c8ba46bc105d7b52c400b3a2ae29d38e7f5
zc387b7994881acdbe043637a71fbccc3424cf29c39fc1817b008dcb2322d2ce6f43816b44ac2ed
zc4958a345d2a63de1e11d325ebe044ca59d02409b757035c1cb285cea7787a050e3523b488762f
z332e6b8ecfeafc17d77610e8acf289ba7e8c55cff1c1efbec95f00248a7138715ac3adab1e6da4
zf943497ca68f49b7cebae107c993e153cb253dca641174c81f072e9819dd92f73f89fd5084c8bc
z5e1b53596ef83e56ab2a790e1bbfd5cedc2f0dbe3d2bfb047e75c8da6407312019f8f545adfea7
z155d272fc132a80c3f5c54d5f1b953a24645dc411f7132df9960bdf038976feeacd140288be9d8
zfce12a30629456eb96a6baf2bb9015bedd22143bbb18eb8d047f162255923adf03c43328d0dc25
z68c9a6513286b3180e233d237267becdfc17346b94bd59d70576e851cbe9b6cb1e77f431f51ff5
z0ee63fa74bd506f0faa0939de13327f9bda0943b195d9a2c0f1d01b5c747d1684961f5a40ce62d
z57d69e54f01e95a318911abfd9d4705d89af3994b918ae3a9581871492dff7ccccd6a68e8aff09
zab4d75cdb6cc82a47ca55fe18c6883d26ee71a4e3e0cb1678d72679eadab3e17c4b6d10d59c9f2
z6458710c7e5152881f2393c542c2aef252b5a4ecc2be1824c39dbc8b37d9acf7758e1e083c0895
z8483e34b83a9d6d7ae124e6ada6f77d1c8dd89f5f24410cbf98c3199e91d19cca5fa6fcb670c2c
z82e01a40404d5b7215a6ca02e898205bafc85cd86c18511eb9c919604a229eaaa33e0a176d07e3
z553cac9a4677fd7e9c41a4d7dfe4de5546b5d836398597bca56aab9571078f208909fa13350deb
z1413eb6c178e625a1d14cab5e95d7a073b2a397159e7615d701c276db0c631c59014c93f3fa66c
z14d2ce5e28f2a6d0ad8e0ff90387eaff882f7d1616a1f087da475ee16b73f8a4c12c03c27033cc
zbb596a0be512bf26136dcd437b05af250e86e884dc79488f1268b7984cf6590dd39caeeb2d019b
z370fda704b011326ef3ce29918630732b935f652f4ee4699ca086aaf5879fa9f7ec7e2a7713b1c
z3199dd0917c621c5c9771e039cf9833d3edcc38870abfec5b1686ecb3fcbef98bf6196f402c2a6
za4eb85dbb26da40b4fc3c2e4b8797f46a2201069ac841eeebcaa6f142c6ea40c6336d519922ae2
z12f03e65cd370a3be02b654aa697415e2f3c58fb5f12b8599c5d329e8d70070e5dab8a391c494b
z667364eb7b357596e1d952e6c6b360774306916b47775ff177e32c19a91e281f83eeb857694a46
zeb2c5b74584b6aa4607eb31218cf382c835616a9abf4e81470b10b58a8733038ab6a399398066a
z12585c97a114596b7a7721c19e933d080a7ce35a3ab74138baaf3ff65966d3efa952df9e394bcf
z9c01450fd7ebf4db0a14db3b294c50ba4c51ebacd78b62ada49547281e38f9c059fb0d6a80513a
z9ffad9b8895ba5fe5221b73c0873745c3ba2a535042fa99a8c9a47499392fa27ca40843649b582
zf75629ed22eeeeee349f7b40d11e6ab577ed030f9488d38a9116aef688c0fe5662bb0f5c95fc41
z2d181ef8455e442374a087572fa6b1bf025f0a49a0f96a8377c6fc624e7d60ad1cfb907a181ff7
z85749d8970b62bfd6771b527c1a9a31284b549482926f2a5930ab1616ed0bd8db3bc5e714b8fbd
zaf4eff1028ba231e2658b56915921cb796a3c41ff43e99ff7dde85116c1cdd379acac25a9548e8
z541b2da70809dd9aedbe1b0846940170663cffbd1e1eb44bd7a9ec7f103c31fa0a95a767ba89e3
z8010ff79ffccf6424b958a86808ea9da341207645f5d47ff5c04bd2cb37eb7761bcbf76b0a6e4c
z9babf54ff6a1c075ed746e48a97d96a815af9c7febaca62ba7d9ef478ed1820446653b42f9cd20
ze96b3630691093b3ccaa239e03a36261f91d9fc360fbaaa01f5dd5e2b212c5ab072c8f93bad96f
z1cf4726065e6e16a421ed891f52f4fd4974f43a15ead358b20c571447e6351b59a682c3ca41974
z1908fead3a34cb6bd8f26f042ad6ff91e2be8c8d1d3b130e3956941a88737a85f5dd64e578c3e7
zc500068631151cd09a709981101d44b7a55ec0324b2cc6d36f82f3d74cae61c6b585948a725401
z965d32f88c15576ce170fbc00e0b9865e17a6868dd35630fbf3cb86a2c1769367b855d352a64c8
z494a0b80752545f2e01d8ca42d8347067f718de458c038148f365fc6a358b868587fa7a52aab39
zef8368f62efa3b705f49dc2d05bad22b57fbcb2960b9e1140f1dbd2afb4df75a37eb9b162ffe0e
ze6fe26fe8a8f79d41fc14790129cfaf091c61933d0aaebecec99e8a84afb2df734bf83447603c3
za514d06731789e5b73e6e00e8a496086a70e5bc12bfa3b291afd7f9b1c1aca694047b25643d33b
zb8ba565a7f7742ffedfc2aba22863c7dc7a941c564fb39522c32f054b6eed51761d77848c8ae00
z865b1d5011107f8758e65fc0bfd61041368d98edb2993822cabcf3b7af2b32edadb780fb6b125f
z68224c56f78a9e7f0721d34f1525d426b39348e3e54b133d80ed9f504b2e618067e03c44233c17
z707be567247cad9f22f0c695bbf52940407c29cfed8d868e2bc29aac796a3111f7e621d31523d6
z6316d23212f2500f44a41d9ba714a4e25f8afe231e6a5c3e0a1aa2b7b530bc407a4c5812c1b228
z10530fc9257ef72c4245c7ed12e8987bfccd86d10caaaae58efc2d4460090fbff0d9b8d485eb61
z40e3fff56749981861532368995d554209bde9415ca7f487e1752a03e0ea2532d393618e02642c
z7ff8edd78e029a5a51b90ff842a310929c1ac61c4fb68d111294b4eb35e4da1c0000d1617aa116
z895bcc906987158613c10e7cdcdda6ccf1043595c567f5040928ee17c11cf0eb7d04fc525e4a2e
z8a60bae424b0832e8a2619e1003d058959a62d155bc49d69b0ee94aed6831b2cbb7edcf20cf2b3
zc0e5fbe3002419f1ea898ea9aea44cd1b2b8fa16557733e5d27f71a882c93c6b03cd448ec79100
zf27034cd5559f3a69d5ce55b01c7c10787bc3b1d3f967176540b0ddff58521e20ca52c02c1047e
zc70a7e70d4033ade2934e852625e64d051155fb0c58e206d72b98503e8d7ad3b1254073768b112
zab355bba8fed099dce6a14724b25163d8d2be3f75c9970f2cc1ab4010ea979d3038943f1712216
ze7c8ed208052c5531a549169496cf82610fe6133674d7767a722b5f079935752e528ded4312bce
z57876941f9bb79295df61ea7d7630c223fc5ebf4ee280c5f5c823421371bfb1bfbf634e949b7f0
z0afd2832f4c8c98f922c5b118ea1a5b5c6fe5dd77ebacebc5d9b1ee4cb2d83af4dd01ae733ed3c
zd825572e800b8648ad4f8e7043df30abf248d67f802a317fb9bd2be65e7578f52f4e68b8b28f59
ze9dde05566cdb9536239dfff18059c766c88d0a11d9c95dc0782502c4acdfeecc623e7532b60d1
z6773b11a9e2822826337325a0d5030ff6ed7c505272b000e925a5ccbccbedd831dd1814fa624a6
z82b0c6b5fd3e3c66aa553b606415dbd176cb0440c49c286f6d4f893c84b3944160d5ca6d154730
z6f50ecf1367ea2d4724eaaf676936a9019be70c9436c6e55394a86014be1b01ccbda57ff76c058
z491ec1e60cb5fcd1709e04399b691177a34c8b134189ffe81b999489be87f75ebab57a89449d8f
zda49abb13d9749745a13738d2714a6ee4837efc8352e2d5e8032422fef899f1e3d25d407a3649c
zd2214d9cea3b8567732f7fa63832ead5d4387683c21eb7e4593e9605f52a7e921e56d9fd79696c
zbcbc64f5b48367d9c572f9450e94fdf128b5161d1871066505452b829c16f2c5878dc0e2c7a42d
z4e3bf47ed8fc20990ff1316146d409ee1c5d9913d3f7b448a255b2f2b5b8ab14e5b78140cf03f3
z83d67df708ed263433a76796af46046f06bc988f89294c512abaafd528ed3158f68f7c1dcb0a7a
z392014783a5c521cd8d8bc871b22dc25b14c540ea6dee2380f21bb64566057782940ea17e6ef9c
z0dfbf23c52b8274d65ff1c5cb053336f12b33794642a52ad7bac7b31df9d68fe7cdc4f53b21df7
z2dde538ff16b816f563dfbf4a794c4bf6c6813d71df4b6e3fa09943698ef34355a46918d52c9e3
z9cda1181cd9d60ff8f2ae73d72ae6aa6cfd64649d089e471d71adb681d85c1248d703d3a0af7db
z4342d9e30a5ae2404a1e86ed0afa1dc9eb480f9f1dc680bae568e5fd68aa3e39f486a2ea8ce020
ze39ebf01c7596308f24b84fa76edcf984d79e28e51db0b2492f757519a34419cd3c9553e7fee0c
zefe20450afb79ca78442f1005c78fb096b2a5f2d6afb6051efb0bea1a8ad76a7f11b8188af251b
z8a6b3499ab62f7ee8702030540324910aed4864a56080a5342079f8da06f6f006fab8b04aae38b
z0321aa6370329c49f9abe519b984cd35fa1187fa2a313494d97d9dad0fbcccb1b795cceaa846f8
z745f9a43a3e3dde17e735e8478e6bc601f14c59c538c90517b2646879bd2f9ec2056f7b5520cc2
zf8324b4310756662b6ced3d3f03bff0489735cec619edac9122a026f972438aee3336d9c5c5b74
z97647370d35bee5485aa065aced15700a85a19dd699f659efbf08481699436a138d94d0ffd7c58
z57ad1cc6151ef4b9bc6b4ed7d809141737704b24c11a55427f0f9be83ca4c7300e25356dd3c0c5
z863dfb7f46f136727c7702b4210bdd91c780770ac433e1791005ec803c5cd135020ad7af8f7b3c
zeab61e54167c37951ae421e5f634bce269dc8ba615d6a71efd76baba947ad3e05c26ed71142a8d
z6bf77a8979760093575894858af619ffbf56703cde661e5d377b26aa8ed1ebe7803950635b763c
z70bf62898ee967ae97111a7c9537ae30e3fc4cd2dcf1f00b51ce679e70084c50a3a412011f9364
z809e194da04a611c1aa9ea7ef2d5efb28927305bc318675c9677b2af7e24b34cafd1e68267cefc
zcd01b361795d6eb47a985b6488a875c3c36709884ba7005dc4cf1fe81f06edbb18e0462d1410b9
z7414163533a06b0cf792309069128353f61b5177a6c4d83b7a7c1b95c3a17a0adb57726da707d8
z02e1513729dba0b5439ecaa91e38fb375f73ec81fccae75df733603171b271f1e84c6db575d13c
zf1332e50daabc46b5b1feadac9662d136473c2cd50cd34551bf16cc7e4af2a089f9c8bf36a74fc
z75ae8ed7ecf6fd28619eb7906f783ac24ed50c863bf20e722c7c92ddcc1604337f97fc9e2c6fe7
z2d1b855ec92cf78976467f468a78b8d944791e199ba67aad1af00195b50971d383693aea607611
z7f252fb2d93aaa615a60cef5010817adc116e3f08b5a6b9c83a1bca345ae69650a9766094fd3de
z6b9937ac95c14969cc19ab161f15f1674b489013a6b973398837cc1512f39b165a1b2b07570c41
za6927a791586a3052d34dc95a57cbe9b6cd4819a130cf407006b4b5719a7428c601a2502cd46a9
z83732a6ae960d4ac4178b8aa2ffe6247e7ff2117d239e299d7217b93c171d174f3dfb0c048fad5
z56196ea4fcbba3b8c0be89fe5fa036e04b89b9bd88ad02b085aaee6d769684d2c6b83fa15bb7ae
z4b2180c8995a1d806f6e17252870c95a8eba309eb3cd761ebffc26335c3ceb2f6da1cf1f26c6d6
zad5fdac0ea5a889001abd187a1f0b0486754fbe99813e47b39ae73e9b8bf84f59a71ed42518965
z92c2ca1b28f9113010f3fed8a88b86d5bfb8098866de4201239a6ce32e6dd91b270f1f77e5e4c8
zb926e983c72a95cada1c39c739b38f34df3ed1fd533f75330f4f971e5410dd1ea5d2acc076f38e
zaf92bc83cb338faff6cef86abebc6a17d10e549d7345ba1dbc0edb3a0d5c7730da9d0a68539296
za94a403661fffb29b42833b39a94e26dd950f203eb97102174b4200472d8799d997dab4f677d54
zd2157315f6e1792ff0d3485fa979ea97706e009b30da31fa25498bdb7146ec8d290de7f7a7cfef
z0cc9f48c1d9f8a01b07a092fc12b03b4fc9bdb9e7a5f526412d812828fd3c660cad059e413c537
z4270299eeee8f62f815289a692fe7ba2cf5ee152d9cd860728faf93f296138e6c66bf1e19ea89e
z7e2ce4e4144c748f3e541ecaed3ac13ec548009423362fd01e03272cc954b235583dfde741b94e
zf94c16a68a0f47f5d151a1475e37a1d7aaf3c0f4a57a45110085ee04a2c6f5a7ed22d0bbfc7192
zd7ff1580731a9d33697136f22a1222a8b1e72dae627dad842a1fa87d1b0c7fff2a00f6ccff0e44
z2a45183b49bb35bb7ebb34e2aaeed4d0918a75ee4b95f3eafbee1b99e24fd6db8ec769c79d2bf9
zd2601ad9c63981bd3e6fbb8484bf124e352d3539571b9e248dd6add551215663487c9aafaf833a
z51e187143a2f26bfb9d3193c6b1974f5c833d0f49fa6b2b3ff7b40f04b691494c4eed76a015bc3
zf555c9eaa6f83220bc66ac42203b60289103cb4003e0147a93
`end_protected_0in
`else
`ifdef MODEL_TECH
`include "qvl_gigabit_ethernet_rgmii_logic.mti.svp"
`endif // MODEL_TECH
`endif // encrypted_0in
