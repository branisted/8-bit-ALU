// Accellera Standard V2.2 Open Verification Library (OVL).
// Accellera Copyright (c) 2005-2008. All rights reserved.

`include "std_ovl_defines.h"

`module ovl_fifo_index (clock, reset, enable, push, pop, fire);

  parameter severity_level        = `OVL_SEVERITY_DEFAULT;
  parameter depth                 = 1;
  parameter push_width            = 1;
  parameter pop_width             = 1;
  parameter simultaneous_push_pop = 1; // Note: different position than in assert_fifo_index
  parameter property_type         = `OVL_PROPERTY_DEFAULT;
  parameter msg                   = `OVL_MSG_DEFAULT;
  parameter coverage_level        = `OVL_COVER_DEFAULT;

  parameter clock_edge     = `OVL_CLOCK_EDGE_DEFAULT;
  parameter reset_polarity = `OVL_RESET_POLARITY_DEFAULT;
  parameter gating_type    = `OVL_GATING_TYPE_DEFAULT;

  input                          clock, reset, enable;
  input  [push_width-1:0]        push;
  input  [pop_width-1:0]         pop;
  output [`OVL_FIRE_WIDTH-1:0]   fire;

  // Parameters that should not be edited
  parameter assert_name = "OVL_FIFO_INDEX";

  `include "std_ovl_reset.h"
  `include "std_ovl_clock.h"
  `include "std_ovl_cover.h"
  `include "std_ovl_task.h"
  `include "std_ovl_init.h"

`ifdef OVL_SYNTHESIS
`else
  // Sanity Checks
  initial begin
    if (depth==0) begin
      ovl_error_t(`OVL_FIRE_2STATE,"Illegal value for parameter depth which must be set to value greater than 0");
    end
  end
`endif

`ifdef OVL_VERILOG
  `include "./vlog95/assert_fifo_index_logic.v"
  assign fire = {`OVL_FIRE_WIDTH{1'b0}}; // Tied low in V2.2
`endif

`ifdef OVL_SVA
  `include "./sva05/assert_fifo_index_logic.sv"
  assign fire = {`OVL_FIRE_WIDTH{1'b0}}; // Tied low in V2.2
`endif

`ifdef OVL_PSL
  assign fire = {`OVL_FIRE_WIDTH{1'b0}}; // Tied low in V2.2
  `include "./psl05/assert_fifo_index_psl_logic.v"
`else
  `endmodule // ovl_fifo_index
`endif
