`ifdef encrypted_0in
`protected_0in
ze74c34e226135848fe16db9ffd31815111b6d7fb642c521a3f628cf6da949865580b22efd062a7
ze90adae0e65e66a2c36a587d0a790699161455169ed55a01f2084f11770a774ec4c588039b380f
z6de9c5084882a40b79a175f5c2114b2b6d78b070cb806e1c0aa9258297f4687ab308bc470f0040
zb0b1de382961eeeaf2e279e1462520fc31c119af8f2b214846f56c2b3cd2eadbe4099496abff18
z15cec83ec4a77b868344aa20ba7360908f5c0de2a79abf8b3534b883bb12180f68b5d4beb444cf
z3fba8f13afb0abfe8fcc4294810f75afe452434d2d0f1166236c82f76edf1e12979f04bc35693e
z32ae028996dd85737a8f5adc1ebb94f39c940246e887647b64782cd7ab429b0544c173176cede7
z01dfb26b1f73408344a52b7e1f117f12bb9c8077b34876c2e6fdc085981637012dc9754765e1a9
zc512ce062e0b8fb16a214591f5c81e1353b900a611fe1f4886b57940b41b7f2ce99a7b84b04b90
z916f717e73bd10589c81e207ed77ec660a8cbed5b487fa50acde1b055c8870bd8676023f21ddcf
z9c98cc47cfa2d654ff1365d1f45035a045a66c5dfa82790502623b57a3af03bf0f0c0d35b51558
zb8b5f2d29acf03737a9ca2a053b7a8f06800d50b465c41b30eb585f62f3d0c2c5a43bc89607e51
z10be237a925b8ba7abe6c5c8b9c4aaa6ea797a95e6129eaf34f520a1dcf43d3b93588d5095b277
z416b10c78989a3e94defdb00bf6a8d2ab27e566b83eb0a9e145a0b185e90ef6debb8bf7d5f63cf
zc053ab961159cb0153a3fbcf83b5bc2fde04eecbcd6d4e656171e795bcdbbfa79735b8e3d5f8e0
zc89a1d964182f58494420f17cf6fecb06715113df7c956e09363fa7fdd2c717c5c1994d8cf51e4
zbd03ca46472b66d9b8dff7da0dce58263dca8bc89ddc3e75f8b70372d9c33778a887a530853aa0
z5459c50439a82d1c6258c9892675bd78fbea967104a0a4a60d1e91372ef44338068110ab5bbc1a
z81d051deb1fef87153f1ba99d5fdaec70548bb11568218224a1088126e5add641e8a5916254566
zb0475e2b853b1ba91b2375a93a1fcdc393467ba36233851458736dc8fd538b9052e109b1e8299c
zd5638a76d33356de1862cf8b7f54619a655846fdda90d5c8434b81f6571a02960eae0727b52746
z7aef979275530bc48128089fccc6a74d17a225445f150a952979fa313d56f9be93ec351b8b34ad
zc36606a68acf2bf9661ead2f571d8645f3bee0338a125d080d8dfcbf350ad3aa29fc1ad18dc496
z3141e4f44a83b2f1f41d7318a26d7c26157ce69ccf2a71f95bda758d96d8a949c535d1ff64a135
za4f3bf4c78c30d28fb354db294c123db5069dfd386eb05e28f57e4d817ab6d467ec7ac692b0fb2
z4f2fbaac689742612a86cc96b8fd296626cd0a46a93fc1b2eac0577afa164c516677ec7aa70b15
z69b73da52a01a9f21ddd66c37c40fa0dd00e0694fe5f9245e25df6d997d7535135f668050d258e
zc22bd308524299f0e83ac307b83e2a4dc3edfe5c61bbe997d0d63d056c5e90bcc1096e5261bd35
zb8bc27a573a052e4e028d0f1fa97bbfbc60e6e1e07f6e542ee6bedc466ab5f676912e31a6825f7
z4e91f3d966a1dd21fcaca4ac5392dcf5d5f9ef171488d6433ed1a634964b06fa8cbc1b49b68eb4
zf9b813cdd1841a35f7bc05c7318ef1737296cfd55244a0d6cea290f71c0c55f32690d622a09156
z40da63fc79693aa4512fb2bdbecaa82ca26f772f39ff534666514a0fcf5659e53ba25aef19faac
z74b92e8fc4aa17cd6dc9eb8cb967055fdf18ac4642481910ff5934e63a32d4a25873b039490d53
z388e33cad47386c27f18c4ace7ee9eea829aa205fae8ea8e7d18962aa543372168270d00296813
zf01bc2a942451b9e4e3bc35a16e80aee134d481b64c2f145157880c9aed3e06c616cf559e8589f
zfffab9d8ba8c521f79304fda9350a5f628dacd79e62c8405f86253cb0e7d824c1f51378cf6d8db
zee8383ed7eb05385dbcd0aff1ec64c10a2d906eb42494fccd091cd6176a273a567e7962b33ab4f
z2b22a2c1789da1b993dcb0ad9242b0d624697b968b0915d6ec04450d4a2c8d60c75edaae762a1e
zcbf2138daefc71bc8f44e29df3a2c384cf1b0a0b5152e2756cef673242450a98c14d0f6693f7fc
z6ca98ba89084d86679346abf39ccfda57372fd1221797ab0b4510ab17c103c006eee7c013ad8a7
zae4c6e1407e605f2162fb300825741d70958aed31b6fb49ebdf8fe01b86381b451410c92ba7be8
z4c6518f7257c1ee4783fc1d415e08c9e4c3b3173e27bda72c8754ed895bab4b812f0f7cf276d69
zd1a3db0e310d0240210f1d51444b7afff92d9de78f596dd88d42d006c80cffb13c2443b69d7c2f
zacf017b1a90b7959664df9a9f3bba073ea2ef8ce1af5afe7e00cd91ba8ec1a6acb9985532391f9
z81f3843c4aeb4d3d02386ab7033d4beff1f0c2f28411092842817a0ef45293ab1890d1abad944e
z3460073af173becde4792e56c528480eced4d34dc221c06d9be9e8d5b7470109282b3754c5b42e
ze82b024bf4c2a4a0600d398a6d2226eba46b1c18e831ea169208e505073b0a351f9a607d9c977e
zdc057ad46884328e80b1f6bb9eca88715c7e0dca8bed6459ea7be6398d16a8002383b67f513f31
zf40cf68635ec6e8e1c4da3c47e4f520ad589bd41ccc30f3ae879f0ffd3611321a626648f328f0f
z8869f6e21e58b05c4099c11cddfe4fde427161aa1071670a8c8a57c7a17feda34b8cbde3e537f9
zdb3727fa09988bfc7ae80e688b1006252550be3de676e8ae38e740b07a03f10d86571ac15bf320
z4e75ca2236600875f449aae256d76b9fbfb5a0d2e1e2fa6af8a487097da3b540402a98d7517af3
zccf26ea29fc76d236eabd14744a8ae61b06a9fe3528a22d5e8e5cb2e04e1017c478baf0fe08761
z529fc4be04f3024781a2bb6763488955b83ef16cef4770f4360a4f48b8b3ffdee4dad805b283a0
z17ba8824fb9f862a10be8d9a1489de10b50f175d265ad10ec37a7ad02467a6694ce63339ce6cb0
z55eb7366ab26114aca7d07a1f44d96a1239d6c1348b09c68e6d8d5d641b944d8a4b691b79f9e64
z40e0096be2ed9cdede07d6a63ac6aaf5068f210e66bba90bdb9ae904161f3a8e67cc562d63426a
zb60f6ea4042c847453b409734595d457d605ab1e007141c655a8bcd3fa306777d5bffb9d31b485
z97d25144c5618b03cae5a9a057a2a0bdd48f11766786773e8c0309d6a2e0607aa3c3f417809b43
z691cde44ac5d76cdc52a4a58cc70a955e2533268ce7ee41c55d4d704f0f0379d01ce831fad1b83
zbb76c31216c8bee6b9f6c0e2b879f724e97822453c89fb3ce0be8104c40af16c12a230195782f6
z9e1c52f23469d3c56899a2a741b218b16c1477c499c20b68559763c8303fbbdadba930d14952d3
z4a5bbff095a8834750127a3b12d9bd52462d9b7d0aab396ac16f3ddb648792b6115a3e96816210
zdbccbd9425c1f89ce2845a92a911e627ae35c2668ba9d84a51765be8971250dbf653d52f285e97
za72c9e32f119fdc6a2c01abc365888e94378dbd4a76cb29c4e31b633d4f63cbcf5e3250dd9be50
zfa4d8a7e40a4c7f431bf1080f4661b60b343d88b4c5e56c451d32d04f7f87cb185929441dba7b6
z68970e813d181e4c7b7685faa554b3d75bd69657d10a614402259a1787866d3e69461d08fc580f
z8f3900dc18dd40ccda78663560da187f9b4344ddc3d1c60c55b0bf17a40e75315193e724e00337
zcc3bdd9146b33890e9c568b7c5a78fe5ad2cad89c02cda613764394a1f6ccdc568ac505f4668ef
z55d97588724cac2bbfa4b1a1a3fa408c4250e62bc00e2c0d89bdd02bec0a0314512ec1e621f1ee
z17be65c80eacb5c7143adb4be4835810b26ab3ae8ca6381bb4daff723d8bbe89b6a1e68f37a49c
ze4bb60d340caa1872a6acee43e177a85c2f132ca5ef9200f77f799ab841caed4dd93575453da33
z2171cec231a7d0b32e3a54caf7aa4ef2c2bb6bf0952c3acceac225a684e342c4231e45a571cd99
z3cdc8687e20344d1ec9ec7b3418fc57baa2ddf5efc20777972842ff7f2fb958931fccc6caae59a
ze3c06d9cc4f0906f05af6319dcecf86dd2562bbf054a6e8891ebe03affb7e331f50cf44b6e7a80
z9611f9653da9a2e0e34b0e6208b7b000b8185bbdf7abf0a849cdbb06116777e55bde02d96ed1f1
z23e8011b96a58a3398ba5bf290e1c9f3f7e6ec47e7eb4127336802c0d1b1f0fe4e6540c89667ab
z356b66e0f0295165851236e366ac49a5a44aba12d1169f605ef2e55b6fab85a193a23e9a3cb98f
z9446c031a727861e667419df9306ebf0978de4f90c4efc61efb07e3f3b11fb595ffe32fc5ca092
z187374077748f12fd47713b3c5ca2c0dd5201a5f26537e2bbed44a56a5fdb7e05ef66cca265a1e
z4eeb1728fe54e05a1169ae0db6d4303294e0037c8737397af4827e527d0ecdb189a3ff324bc0a2
z593d97eb3f868182836729b9d7e4f30d449ca22a5b24d641a21b8577842d167b7ab6d3e1253133
z8fb3e0bceb9bceceac37eeda5713bb0a99e9e1551e2dc083344b6e4e849cb920532d40f437187c
z7972d998f1fa71fdb290328732cb2dcbf8ecab961d588e84f706fa583c290e999bb9bce53029d7
z4811dd09ce22debaa9982146ad79344cee5543bbaf0b62f538ef6e19b441d095985a76f09d3b8f
zbbd5cb05520ac44d3eaaa645f16f77bceed6e6fb970213354f7ef66e0cdde6a15a4e0b7e66216e
z40e3caaead2aaa7526c8f1260ccc00db7793cd834f28eb998a002d53f0797442cf3c887727ba68
z8f7e0bfbe81c98d24589a9e9e161b1d0d6ee11cccdc682eb51341409bd808b67ced576a085a821
z99e40753e7a9bbf104a77e4fe36176437370f30e2eb3c28fa7915cc8b47a202fdb514fcdad3544
z07cb902aa65831fc7f6a3f1cb3205285e07d903c758d3bb94d85c65bdc76bff887374781707e5b
zbb8e0a9742a6fd917b6305c779cf7fbc469eb057fe1fd9407320399d617184d615554e394b9a07
z6bc681b714fd6b3dc7e386d17e7557f580878d871679295c94897191e9f71e0b42bfe34b858f71
z836d0c8f4b4ea56214ffe7771c38e059dbc42be7c79ac66a3efcdb5cfd88ee2971f1eece98d327
zb33b79eff7821f0de1deb05355d6e049c62208d26c8878038dad87da5561e481d12b5ff05bd1cb
za03ddf4b4bb653b6d7c50f9ceda3196a37269ebe4b1adc26df549e8b3484b3854811111ac186b6
z8d43a01a85857a8ab25240e489fbf3d197fb0d22b4f7f820ab967fe1f53a09298ea8da12ffa11a
ze6080f5b970cd8075a5c9cc9ec397cde77109e80295ddec64dbb10aa6fd05851baaf4ad90ad149
z8f7dfe7f7fb9c1601f9077025b85e4691c40c37fc2c8ec3ed642debb9bdad409a7f383bedbd891
z96b8dc08dc3e85e293c5bcc9b8197f2c0a8bde182a28fffda8736226d8f91b059b117b9b2f5d24
z9118b3eeae118fe39d00d9c9070c6f6a87d1741b132586ed975d039941d3cb2bee7fd35580994c
z6bee09315c4b9ada23ff8f8db8405ec8e518b9ac5368091fcdabd87e784cd11e2c95fe4936cc73
z736432139f9e86bd573158d4bdcaf12791b96e34c0bc478b80baa848a7c43487a1d837dd44bc3a
z7f885d20ff0c1d825cf1cc79ba2ab56940c928f1ce2a941b63ae441f66fbafc42a1577e48220e0
zc125df4510c063745ec25074ad3c976100b710aba160c064aa6a72aa31ef913bc591e0e03c678a
z20169bb198aeaaca212a456e0cffb2fd3820244d6f267811fe6c44118484ef3822f086b1373b21
zbbe5e09bc8ab9b20b77213e2ef8fdc367507d9dc68659fef5045fba54809f480b87201564bfc8c
z0190588ac288a92b79fdb0403540e2da4c9cd8785d471953ff1f7850cf804f936ed7227279a8b5
z1b7078f8e855f06e22d3659a2b523209986c89f8d1c73a04f0ed0f51e0765965be15d58003230b
z061323f41d9b28a7aba846e72ba96dad79136933aa079f9822565820444eec387d206bbf281172
zd935d555321ede4364091f71e2a347ba16c9907bf43961568c331541c9bebee7a1849c4964dcc8
zf1ad97b4783cce15c6c57119ce05fcf05fe37fa88bd2418d9d61af2e51ef09c96f32e5a8b7fd1f
zd85fafa7cdcfa4be66e2190bebb2581b98397b594505156bc8ba5444bdfa8967aa2272d991b48b
zbfd61411edb8a9ffecca4a2b8f6ce2ed0b3ef6783b20d3415d7a8fd0fb9eb41863ea81ef12a862
za3aaafa74ca0cbbc2cc5a1b8088f57e0dda8edcde4fc8848ed53f8faa16737933a0569648121bc
z1ea7b0749077849a10f96d839c1c6b7a9b9cfb0f3fef91a7ed151256b1cf1281b6587b626823be
zff8a957973cf65e1339e5a97f59c5d065d98f70a460d4746dd3370a01f1ff81c9a1b3d661a3cd3
z52ef3e827cd2a4b85ad1f8b6e95f975bfa7a1cd546982653e5b15e4b49c5c5e24973d8818c46c0
z9585ae4d30e5d1658039c0d0a1e639778b18bcf1c4eaad9394b1bf082506fe922d989f4b11dbe4
za9a1db1232ea7e0f5586403e125e5f3817e5a346aa27039ab540ff6fbf4ed2a3cbd658dee36894
zeb3cf4588f18d32c820717d4f08adb23a782ca87b7c4d7cf6fea5f3bd4ff9ec9f0f76f3503eecd
z2739e66235ee68617747d69df63d91e675ad6dc02818985903e3d68f1a2091c93bbdbbce24b1be
z719ac48f50a9677575cbbd63af1bf048ced8a4d1ffafb0608f7b355ffc47fd74246d7e2ffd3e5a
z020290a10529303f61fb314b8a1a9e79e69d7e5ef039cc9c81065ca79aa03c2dc806a8616ae0a8
z4005a600740d6ef9f0937ae4f2cc4073a1fb07c27e8aba592c6cfe33ccfa7f2ed2ed77ee7821c3
z05ad080c959ff38068be684580302216f998ac78733f2831cc0433ca1c0008972ed3e784516d0c
z2896b34df3d320d267363000a91403e4f3d74d3d24c14c26f803365b271b45c175a103f33dcef2
zdf59e2e160d355664c9359d4639d85382ff1b52adf1e0b320cd90c17e342c714bbdf327e2c64a2
z23b6084d77f92fba4a119d9cce330190237b162538672c608c051347bb7c13654e01d628307bd1
z87a89d5f7ae8c51bf44087d9b38d124810758907c61f6d0fed49b693575b06e4d94a7ea1aeb652
zc26ce6e88ab24762d6076c05f26f88469bdf10b2a7ed738dcdcdcff10415836a9af6a835a11a0b
z3709035234eee31bcb2da034e9836b634470a195a38097b81c24564b982457f35107aad4db82e5
zffcdf4187e5da0714a17bf816acf09ca59040f3b7f5cff9861f4ec50b9b7d66145b59724232f88
zd3ae74aea8842490581539eafbec9d178369aa48169506d7d858a067910cb846c0707ccb1ad250
zc7b8d9bf482e71e05522aa0af95edde41af740130a8b30735dde9169138db08a0d2303c48a564d
z7f1bf6dd64ce4331210986a6140249805a26aef6a01a3c7bf66e239fb2816e5c397bc3302e798f
z2a11794d32a38eadc90956344374ccd5072e1e0ed311261c0747c69d073ed3a807988c4246e4cf
zf5bca0dc78b9f8ad315630328c044f25ebc7f569dbea99c3a3d9b656418ff6479929567b646d76
z8f538bb619054690b2c829d066e39811bf342846040fdee3b5fb1be2de13cb8bb1102c848fd774
z9ea38a4403eb0b1b5ae8b687c9e765acc526ff92517ee91f4e418d66c5022180d70e4fc501a615
z72c28071622dd6e4dd7c8f2f51662d8672858f867774363b5b1fed65a70b807ac9d7ab9da4060e
z2cfdabdacc89ba2c11273de7f84ec0ffb17c6074118436f791ae3c60dce22cf7463e904792ebc0
zafec8220cbbfee6b40ed2c39db01f97ff8ed98ad6574f4d65c7f1293cacab478906af3a498228a
zbb2f9138a5b7f464fc4ffbb2508457a39cfa7c6f33068792fe5677a8622ac2219f83ce9d5996a3
z6b0840c0a8c8ac74e59f66ff09b1bb24aceb21cc8ee30db3ad220737e17a2655df8e0b51dfe161
zb06cb1d11e1e8a56589dde6c93b285dbb856d98b3d41b5de99127330f2d4e2bb2d40fb50b070db
z12ea0ff404f0fdcb8a83784e86453320885a819c83282c9a2e47aa265342b235828a531bf0d85d
zdb58e89bda0f5cf52e2adb4a9e1e37f02c3a9306897290bc893c9ebf0874128610129a814b932a
z3cf524775a865a73ebf78e08acf4c7c91baf1aa6b81ba7f295f4c2b5afc0f79ad436468c6e1787
z9d99cc73e0b1b53f6f180203d3d30f31de9cd23d6236808dc35b36deef65e37f4e5567f1ec09e9
za9ff27dd30b309aec5fbc05e358f83cb74e85119fa50b074fb750636c17440a450c55ec48944e3
zf806ae52a7eaac5243600ea2646368e18c64a9f4e7aefabb6d8876958d7d5e27b1c2b4304d5c5a
za8ee3c2a2c0bccffa060c2995d45a0c53c2bdf553b03d894260d612f00abbb9eb75cce6c5ae8a9
zc0991758ff977a541d8f0e0e01cfab51d769ef2afe247c2af3470cb436b99879de51e95e97807d
z626b08390a0cabf2a4ac33d52272870cffc6faebdd34838688cf76e74d45706643ef62036adf2e
z53458508a5a22283c0e4a2fcfd0b63285feb5c6755baea7b9e961c4d5b9431af8c8a38c5971e4e
z7732838ef30d65ce00e4a6f52766611800418af8688737ee1d5e49f98e21b50e57d9926957bc37
za456bec741bd925867a4075d7a6b04aa3287dd0011b12326a4702b1aa152e2db4312ec0e06b2a8
z3ad5e0dcdf1dc6504666cfd0a3f6bbd1ab1f57bebca397fd5a55171716a5485d07bd0348f6b224
za8e093d74c6690048de8a083aa34eab315c8f50edf703ff70be17739810a6668d3686d1ae7d540
zf5e206ccf58212b0355aaca3194bc1717ddb20c8038e9c6278b47e2c76ebbf386f59e573a25987
z6f546756907a11e7e4c3712f2fe4a102b1570d82980619dfd86ee58eddcadef4949e29d6ddb9af
z2283ff46af455816819e776d6cb5a68584193192a5c082e83bf11d8008376561b55ef96278779d
za7375498096bacbf21d46c64ae16d3938b114cde3cd07a8c48b1e62ce937b0de9b87387c170a17
zb82ab132dfac2b7a782d9ab2eb82c2085184086070604ebf39638565cf75fedaf5e4a1f538c473
z466c3aa214ff7862f5b2175bc3da192f0d6eca61492f25fa6be4b6bbcb632af68ad492f3f6eccb
z5ab55f27fc51f4481352b742e4c6e16e1905958d4974a703e3f2f2fafded83cc4d9aa7618ebb87
zb67382738302522c9482951c55d80386386fbbe30f02fad0b1048554d15a6e90ca91ab855dd5a4
z6ffe49fed45491baafac53c8ea0dfe7c2ddcfa03a78167ef8cc41ffa42887386e2a1966b8e1174
zaf89e3d9d29631daccfa1d1b3b0ba38d6cf950ac327ae4d6bdaaec5dac7a56f8bee6262694f439
z849ad6696e6126e3cf2d1b62f8b8a00924546478163831fd93f306e5ee2f1e5b31e1b0312b5be6
z48bd55201467256a0db1ca7d2eee92691c51c9f6879b22f233ba1c46456f3d72796682bfd96700
zee8d57ba26489e496683e549bd3b1ccc4f59acb6130b325d030bd3431184a6ecb118be24526dec
zb0545b09fcb3da8a48ae80dfa019d96f55248732ae063b0159139548516d6654bf6c719f3e390f
z8b70edfd9d33a9ea39606fb123c654769f834bd13945686a2ec988b05795b492246ea0f3f1bc67
zd02ca1bbd06abf8191e45f8633187ddc87d5b4fce6d7d4b929f0ef1eb66300952ce3cadaada7e9
z6dd77764624e81915eeb0288a4c2e68e4ed71a3c2bf37123c39e7460cf53e0bc99e23e738057ef
z243d2e7aac71ca44b4f6436d69bf9d636e1296974c0ffd1641b8ad872f260f392785738eeddd6a
z0fa825e049e427f9b6e953c37f88664da66484dca32a6b5c55fdcfe9d215dabb4dd5b82b52855c
z516b296389b98b4e748a78182ca5886b9aee509f20398202550544d7ef2a2b1db34f05dfa1e0eb
z9312f4e4ede635c1533f44c427d97b8ce5b8667850217682b6d0200620979a7fc23b28b8a10dc4
z4baa6d3a15e0c20fd1a36c3b420639bb8594f9d83c584add02b826a5d3254c2f8881e8a59ec2ae
z4ceb3fb0c6f142f31ee35d39e9abf53f46c06a49621fc6a4bc32b3da1edfa12f9c21bed1803e3c
zbf282b4ecdee399708c4e543042fae30ed65516a7fb60235710a9f4ef0049f857144fca04256c6
z50df1c85e4013a17090197db4834eba92ce6e55179ad2bbbd3ca42e35e11b64e132872a9280a33
z023f8293617814c93933db2a29d2c48bdea91875f9adb8f44b8c3cbf98bf02e681007c872d2871
z6c1a2803460e20c3ffacbc619b9816b4f3b7640edc4695306818ed66107f310808230b745d58f2
z675a3bd9462ef76a98fc355ed24ec30fe7d2c383b89c0467e94d2e1b383caddbb1bae535a13ff5
za720f3ed126fa624555abd6a8806e4a325622391c5d4adbcee5d9f08603c94a05e9b0d5edbf9d5
zb025dac7b859efe4dc5c7c7aa0812e9319f87a8210a3eea7d423da786e60d31da63a8e89273f21
z2f5a259bc3602d6e02a47aefd59637011aa64632108652598dc3c8e6a186b3353366218eb85c67
zfae1b5557c05ca004cea0e26dd86c74087d1cada9401ee802d2720c56ae2aee4691fd6f76d8a63
z8dbd1b96ac537c0d974ed3470001d70fb640f53cec9ee13f9a0c29c8e0efbb5356393be4077b10
za3c2ddecba2ae25c0d4be1bf92077960d1eacbfc5924d9ad305f95ec0002ba53e979f7641c5634
z9dc41f694898e506c4eec9ad8616140d71356716e7595b56a7f6662312b6291918170cdad0d248
zf105e312fd48ef55ed23841b5641429170e4e1e14c50affb0242d9886592e972ddbd7a0e4353cf
z894993010af785599c77737eb5e9e851311d3bf93f909cccf33ef374821d950887b225bd5d6a04
zbb136b46e98e0c3ce535bbbafd5c463ad617327d6b3b27c64adcada20f203ee562743104eb0220
zf260283f0633bd7f8d8477024ee97446e07231ab31ef489394e9bb63a8cfa90d55b40033403a0c
z6a193ab684f6eb1ebb29375cd4b3768450503b151c548bd75ddfef520acf3fbdadd7c1c257ea59
z24fd7f22aa8719ce33269267a5bf6c4bc3f575d346f6feae51293208dc447527b6f925ac7ac3a1
z3292c6d14db36abf2f43852ef34a08520a1056a2ef1aad6096c96cb09df0c584801bce17d72ce0
z341e5ff2913a5ac0bf85e9a17f7638b97f59d17d885bb6727b3398d15ad5479283e75e61fcff1d
z97695927882708fed55bccb1784cd533f651c36deba15c1caa20fb9881cee3ef5e87d315d49022
ze8406014c320b5f2f0a8b6ec73e9a2ed7b67387142083e235805597df0b36539eae2f89ba22a38
zc64c57cb0ad773efb23663aeaa34fa485c6d5fbd398228c3bd617913af3a04f197635cd2b5f8a0
zf657ed511b417fb29b941c1640c67ab4ebd0bf46a0ddc80393cbb73014bf776ad438ea3a2387dd
zeb804cb9efceaffd41c1cd17ea1555bf43e2c515eb333e718f885982146f9c09a18dcc411a8dc9
z88c9f962f9aaac99664fc39bba4eff741f8b4846e94f52ce678739e72e2f3d6c41b7bd58b3a6ac
z94bc8d9cabba494689fb9e5aef9ddc2df44eeeea2b0d54281fa6dbf1a7c9d814f58f49496e3b3a
z33c333ccf6f1c440545fae3857e926188247a238c86e3395c44a288eb2eb1273f6b1ebcf322578
z443e3f4736dc14c063595c5734862a1f75b73566a16fb49d2cb322e4ebbc1a523f92b5990a8358
z0ebc5ab45cab8809c995c9a39455973e729c20f990cc48f067035a6b79e00b4ecb17f4f732caed
z5b8a2bfa5c9ed1bca9ca8ddda75974c6c9dbc6917ea6aaa8847af6b3521234abf7b1ded1e3d238
zf85917bda493cc43f8a23b6c3d774c03fc045bd88618e1118f84544dddd607ffa06755fcb8630f
z5df1e35a70cd7c886721de7f27f40bd5ddb3150b3db379a4d797b71f1f3d17c9c35409521bfe40
z8061a308df41573a7b8953ddafb8c9f1b96ca5aa41f46a3ef671b9d64bd405f9f890fb0ad890c9
z2514b9f5300ed4eeda28e300bc7d2694dda0922caa80f0863acd3008edc1fde96aad617b6584e5
z522313b5fb05232d853e64179032179fc10b98d1cb6d3de92b322656fa1f4dcc85cba4de7cb44d
z53750563836ed1b09d684e0f315b41a7e13fa6a11c4b52e4ee38c4b45e0863d5cd4cb77e4c41e0
z5cf4a39db9f7e31794b96e9ad2754272ae01283b66e3b087879674da28fd5761de05c56917f3a6
z111da49fa934f5c8ec651d8fb1a48d59f15f64bd64656cdaf105532fd6949fe7eb47c799b04fa2
z3c4278f93fc98d5d725c7a249297abeaca8697d46f341707a196eee3709e10a14895089841892e
za65dd089f05c8ba0f44864cbda501d48074044eba3791a8c8170f7d614b210e7e2a35e0620a6a8
z589890b2608d7bcba804e3733169d7a76937ad74bc7c408efddcc406ba3d6a3e8267762e184475
z3d7e8810b57650f0395c23b6012162dfaa5cee914fe0604f724724706879f512597fff57968a53
ze244c71a39879b7fdc7a35d7811df0653e3c5598b39abb6e8b2e991e9225adb20bfb3968a4ddbb
zb4084db6b30b18aea7b48d3cbd930a82a307bd15c24a67ac9f2cbb082359895e00ce7e71eaf957
z5185f5be5660222d5680d2519a4f437cdc41af89079ff83abf49057784a53271a07c5b14c34fec
z09ba5b8376f1005d7ce99ad7f46a001f6a587a914cdef37d3f7dc8c245dda014f743e52ac6cce0
z183784cf519b54085b9282a00bb5c2850ed6b7cec6cb99bf64917634f3af85f1b4b7262ce29b57
zcea496f3a8f27c09432983c8cdb99c9527a8b4a35845206e217096ac5df2c3c50dda2261bae47c
zb3ddef514fef3c992835d859848419b7e644477adc334ede035cdcd29565de5a958a83e3358b6e
z9af54be23d25bfdb13d9831cfbac8701bee2a6060e77a0b2984028b663420c75632334b34ae97c
z24d18ab8e8cad4be7ff1749659b3c0379fe6ef59876b83bc98ace1783b143662ad0ee2b489e869
z6ec79c9cfdff1fa3c4089168d3d82c5158c8406ae0cb5449c91b52842e1ef12c1089787e706429
z15927562ecdc8923f668ce5b75ec90de11f1658a79bdfb30cd4e10ebc78c38dbd2af27599b2eae
za3879b26995acb16f4e6bf9c9c5a372fe51ad96eab830e7ea6a638bcefe70bc6aca11de6579b73
zf23e9357c82af05d3b7e5d1bf2a38649a5add12091bbeb34b801f278c2345442d905c072a12549
ze90af2e3aeb754b5fd99ecbbd136a922374a0c9d5480c2fd5c9185c01272f82ed26cea491fdc96
z21b77613050ef5e01cdeab0f4df317a321fa4bea8bb30167293c2b0b2eaba47f279d0f2e6912fa
zaa840ec8d2a1bfde6e3d019eeba02085e752d2359f951879e0ca4e4278b05c5878114b50c83a56
z444864a2f362b026e75616e33a0a7230a2a368f52b6c3e11bd5bc2abc46f192c2bc98b01df2e86
ze38d098982e09a6c862700a31f845105468b0767e9c6af7bd83d5e362918506cbe27e0e85b5720
z0ee0915cdb3636bad50bb08f7611a394a370dcadbf6241b3658a5ecdc8d2268d5bfda68caed9a9
z69a5af33b5fb52fb4397eb9cbcfcc2e493b9a1a71b82e70e96646898b98e9ba50a8d69c5690c0b
z432ee2239a689a7b1886d8df774831c8ad7751544a3eb7e947741335db88eb42d3ed06e5d9cbfd
z6845e4d363adab39e497d6bac9f935a3bf15527a8d5a701c7ebc8e89b28adeca1f9b66de9fcca3
z9711558ccfdce618ff2ddd35b8664fa3d9fc8c78634df9c94bed15736ffd2db2cfc1cad52675b2
z4ef7fde1fc32acbd11b729619862eef3ccf27e3e16c6040331c0d905867512661e5a88cd2bd57b
z1d1a1ea638a9c9e966daa1f72ba4af07ef3b0d4afa704d4c5f86f125f0a12092733e40558584e0
zc985279f0004e3d0b905ac9d50f2f6f4d1ce03f3b56ee25edf01f8e82b51aae10fb07331afad1e
zb5391757bd3e3a0216b55dd53de68d991fab5a4abd9ff2b1a17c10058e5598f0b833073971a581
z7ee3563058576bc1ba7931fb7ad2974637ff347633709c5aa848dcf446c0e7df82ca559f46168e
z7c0d29e5ba35a607337c1a34ff292f152efe39f2c70730a7b44d2b08599e3da6665592b5a5a238
zf60deb148f99d193ff4caf3b67f0efb891b616303d9617bb3282b49d2f34b98128d727818685b5
zb86cc1054d7565ca3f2d26bab9748de0f928f278dfde5f34bb74957a71fb8e8c5d747b5ed7fbc9
z149407b6833e410e518c6cdea4703192bacbb6e0ff9bf534ec8a602a54acacd5a9eb204cf518a4
z5a88c9a54474ee61479163665ae356a617e4fd73d54d8d3ff17b290e75dde18454384dbec23aa2
zb53ddc578e61546d5c5d6b181507c0dc17f0d0e46c3b544110663e0c7713baea69a18cb529ad7c
z409dccdffee44635bee77eda1b79d467be0e98f0c130157a9d2ede8f21241e7bc70caae02883e6
za40b4836d2e945b95d67bba0ee159bbd7016115de51496131cdb8065b100f3c1cc865c5cf12b60
z0488aa32012da34354fcc46547093f8209c694e4ab2ce5ab0a90d259d702103334d17fb7dae75d
z0ed23b9bf3cbef92f01408e925017fdc18254c2a473f4a016607e1add49506a5658994b02a014f
zfb6db140c43f4f0a66c4efef00e0608870f03f8a090c738a2c3da4e5b9a05c7eed9daee906c015
z8bc490ec3013af954e2a4addd8ba743c759735d19681f199a399d713251adc513cb80292f7a7a6
z59cefd722c76442581658bd0d9f1b0da9dcd1b63125b5d5dcff7492e1721f24f20722eca55f0d1
zf8ec2988bc80c55baf561c7bf02f77c52d6b7fbe96725587f0afb139de92ac465180046a738e52
z44f176c896b779c51d3f4b82df4c06926f0a39b1ef3065468ac4d3da74c22e5cee85b84a4b06f9
z84f5687a8ea85b91cc3ee5b4dc96ee83372452ac7df22f13e667c4e5a0d32817d5d713e3176b30
zf1568f1f2f37fb702f72f46373888e4864e656a8e916f489bb999fb7a71e1482d59f1daca1c012
z424d1156402e5bb014256111bd9df5797bbc05ade2d9eea0d181a8aa67afdb420420cdd1cc3f76
zb9afa870c84e16745ceae7a649d11efec20948b37efa454c8bdb82748e917136079149ced05b71
zabdb939bc9f96880d78766851655500142b558d0e3e6bcc8ae5e5f502f40b38122db5b61c01aff
z41a074b9105b27937766ded356304e44ba1cacd9f5fa33ad1d68347418ba7214f92773730644ca
zc150f77816cabd990ed0e162155613c725f5fb49c6eac77f4231b73a54774659526c0c7f672b68
z61466596db04e358ff6e577455aa4a2c343dc8d5547c31fbbbe837885bc1768a06003395d46233
z5081957d5044d63feffd5768370b435f420f054421d5f8b6518809e8758f9649f3b157d998e031
z7a5062d58390e3f36798ff2b08a24675f6d5b9cfe060b26a7bc665a68c8e6b5db617b81ab3c6a3
z560179e66d60730d13c57eba9ec9ecd98b5b1b5bdc1048c532ba1416b745a637da0edbbda13b37
zf87d0391aa307af7f574a573395c80799cb696d9ec8d5af65995710079d98236799cd94e23bfca
z3731064579ccb8bba8b9737802716ad770bd21f5c6d7c146d7bb872a76763da17b4d2151817acf
z1ea8697478489e6fdc5249810ee08d58c84f9493a3229841a9e24644e24887ca659dd56bac2fc9
z79f7684173fd58374fa43d7e92176722e182cae02ccd57d3c58c7c9a5179e1de5058434ec9645d
zfba7767d8049d833f84ac4e168adad0e37666d16a3c0f362e0772809279090c6887d131e6f1a68
z4f38e4e6269daba2566d16f9ba2dff87a160214b8969d7c9915bc349bec6a0fe59e8bb104f598d
zd870b991e1a2bde43f06959400a8f9e4cc709c099cafe8a2bbb93f135a5dc344dd3f0c3553c986
zc0c51a34ed4865e3b8a097b69b30337d8aa0f9b5a277763eb87a43b6766534b158ebb847ea0bfe
z1cfb78019a64654a4b6f26ccf09ce1923f702757c4499f9a0a9e9bb507fd3eb8a1ff5abdb4cba3
z8f1d5497eb3a2ce5b1befa382efb8f4866f7e21516b2ea1785041908a7278ae325fe646d6a3fe0
z2f990d20f58c2b9eaea2afdbd885acbd9ecd351300975b680ca9b28087018945f9ec9c37774bd7
z9bf3596ba0071e5e1900fb0ef1b001699c2ad4cf9092fdb4784be1f06a1ce06673464082982cd0
za9a9ef44ea803b0c5133a7f2b1fd3a547ff89fb4e93e56ede02c7b619bb0cc49b21aaefff3237b
zc1fe1ed524392276725f1bd62cb5c04d20255c06abf2017859774db55e8bf53dda1c3512f4e007
z5c98a7fb0922de9aaa92e5dfa3968af413cf6c194d3371eb82760f5eaa6fb56db3c1beb83de083
za38bf2dfeffb47015bb0429390319c2459612779e5e4daf5a02b2282ef8f875ec3fae8532a1c87
z41753687180d276091870012a5db31e3049278a5743174d4726ebe515c3b32520ee1693f95c1d7
z26c82390ee426ed6b1e0c9310f8373c553f3dc474b6de5291eb4d3a1a019fec39f920d20f0f09c
zbbb84326f5ca736e0c6279e63a741c9319cd66fd2592246cfe17682f91f7bd5856404420d8f52e
z4a86c2c568988d4d9243b5a464313f6bfc42ab0b128165f3798ff187176a13ca5afda428c88b9b
zf4aace3d2fb151f4a7ac1697bfc35ca403db82241f45e5479e6c42da08f08ee0139d528cd35afe
z267af82f595921047ff130aaa967ad3eb9e470102b43067a0f4464002bbbf903ad61fd9e682440
zd93ff76c6f4ca4ef91314db16bbe81b8a85616a5824fa3aa708405ba2462d27e0faa245d327140
z537b67c9e8618d1467aebd6af4c80fd8beec084945630f2fdf0941c9797429e727e9b1782e044b
z8a21a126102ad718a054abbba9e7693b8b8dfeeb482b4559f839cd439e8a80797f4cbb52ac48e5
zcd24a1b45ce552fcecdd9b18f85891e2d470cfa06f86f3653b8838c1812f615661773b8a433d18
ze70445706c84b361583150dd5cf34c07d3bc4592daef4d3f21835961ecf20aa0c6d5b0bc5f42d6
zc2fb3afd7840a9435a07e54531a7954460728f80e5f84d3acc4d4d43b6b2a967819a1770636abc
z2e98a6bb5b2df64ced12e69f3e0a61bc32fca5fe40b5f7ba9985d1136eae88f962eafbff916140
z20fafe16be2a579f132367f292273c1cc86fbbf7478591b10023c4ed40ff51c8d650fd66b99b09
z65bbcb84365ee23cb88e80419644ab9ea905895746f1e3aff9a9371bebdbf6a772521fb11457a6
z9dda6fba950497d837e3b18b26d27218d99a9ea8456ea5b44e21868dad4b4480246cee4dee7405
z73d1a7204704afe7dc49d2d9f11e850fd39c4fb964c94bbac6c190df9f559e26c66031a0a11d6a
z5d464588938a54a1e2362572e12e4dfe157e9e782773beb9a347d8e3b76993c923887a7319a39a
zf5692da1391a6247763dd271a3cfb918a6830e48b226ced5145236547788210f7e7c31d6f29a68
z384990ccdd45b2efa5200eca66ad014ed745f3104660efd2823c3e6ce84bc6095ce4a9cd7a9653
zc49250518b90e310d6f11c34cd8443e0602c218f5e2e4d58b3c8b437d5fe591fb39a07f7825266
z252b69992a3ace2ed2cb126c5da6de603e507ac6b49eca02a32c86397e54b442cb4791eb3351d8
z0f737e6a4228748d2045651eeb414f9d1e540eb79e160f51bae77acb0e792f329a87b9f3de188f
zb1c6733cdb46f2f1b609925bd08a735eeb2b1038f1af6d3f297f2a18138919556b7c7f7d8dbc71
z64d291caa3ec8b080d20ce985e92283eb1c31b15d3e7abd4dab0c2fb783a8800ebf27de1489b7d
zd710b5a504e5f67cb2442bf84d01e4988790b8eee620fe4ec7f7e88fedb6df771bda45648de2f3
ze7ddb7b2be11b6a1d5123d65ae4c85734a16784f28b9687c7b86ba090fd2869f1007e338969420
zf35fd26c8a56b41512ee367ab4d3704cab1711fb084527d792c8ded8d7ef966232a1714bf8dc79
z4c4c1e695eea4992a3e3c0cbf1e2ae484edeef333545a5243d57ed521529154ab01207221891c4
z080206ddfd38f08fc9939e723c411a0a290dc4360ac1d7d39c596068c8aab6f5b964d7a322bd6e
z0a7c2d527c4745c78ffdf85e1540a5a2640d05f1b04871c9e0da168f1a0e420260a19a62ae2beb
z34049a74bff717ade896038ae8fabe49f5e7e11d1c19c4971ac7ee296f772575cd647af6339d98
z57e5df86519996b96ebfe374afe71fa0120c4e710d5c22bf88921f6740b539e8b18136a1fe0a55
zb3ce159e79d9e1597ad442fdb2e5c864fe7397d396de16fdef61f587f355451c5b6b74201dafd4
zf493d19fd6fc747cc4caa065431d32d11fe61ededbd065da702858e211ea34aa1b219f2c1b6323
z6b76074f88a450f7cf0b65669c6b9a7dce449cf1a5066709da30b23564fcc6367384cd588f9fe9
z7e05d00408c9ef972337c93874019e9af20b9392816c7b786a47a9cdaf32dbd1ba2a847d375536
z0adef450d7f31a36ffe83c4cf52100d375a6fd9284e49bf6c0e1a5ee29a42a451dbbe047b11fb2
ze05906eb9ae5c34fc6b8b139f0d1f71b72f60c7227342fb82dee69bc0c72e9635bb16eea5f11ae
z3ca98a8526bddc8a39fc238b43f1094dd27c9766656b1ab44df93a36815e01d16c1b5eccd56275
z6201eb0598fd454b72d423c65609c092b3bc1abadb50a8ddd149cda67d5140367296beaa3062ea
z14cbf04550f157faaaf37ea32a40417370eff1059bf132f323d25cfeccaf8e5d704845cd611b9a
z6c3ef9622fc781570589d9098d033ea537c5d2958afc1251af23de082122b9903754f77d931afa
z8e2b0b43ea05e224073d4a699c500bbb5bc6b675e519922d1063c8c55a4562af00cbfe9a82a739
z397bbbd456a3654a15650dfb030d0c036d3a76270348f71b490b6887fc15c560b7db1e79fe4881
zde91af210f447715639a0be53152d95f81af93654a1a1639a238f098773aa29864a7d467b8e448
z4233a4aef526f8b542ef52ceb989e2504f29514119f2a5a09b9ef3ddc9109694bb2d070fbca97f
z41530928d33aa44b66f8372f778fa07731164278647d7690331260717ed64c68232bef30a71f33
z5ab6e2ad7ee32d3b9fe68fa9e816ce6660c482416825919c8d97e4d2285d794aa9324707f2efd7
za221d9189e0a653551dbd6eeb9a954cac9cd3c580e28c794dd715cd7ee92f3de4705c608a7563d
z0b637bd250acd6d826133df8f791b52c94ae906b1b2ecad5706183ba79593a21f6dbe10214f4c8
z53356f9a9e53f11b10ac08ec62b076e498d3c71a8ac8988e5fa534e95862f72c6e10e73aef8745
z1c4a0398d24d618a256ec0b3f75f8aa48143941c918b87a902acceadab3d8fcdefd6c30f34fd0d
z6b30b798af4d0df03fdcba4d84bd2cf7fa3e905bd515b039efe7e1725a08c706c66a009d66d81e
z6a2ee9c5225c4e9e0392f9ff3e023b5977fb8e9906ca70d63f6882b6825ca0b008be1aa0e1398f
zaef47f1d18902fdd91ecff60c1a9150f8c0eb8767a9bdb059099882a7f998c2743b7180e4ce304
z96e223fe3b8147c74a7d6144da4b58d8ec6334aef82d5331174164ebce6fb53f6a27f0c4cc7bed
zbb39daf133a2863ee7683b3a6539b6cdc323d6724739f9319f4930ea56699ea269457107032d21
z5b1b534f05cb67f340dca587b7d0d9b5678a0c0eb8b16a0c77989953366eec4b37fa39d439d179
z55e940164a285702d0987748ae63d4b47b3a2c5579506af61df4304c7f2b54e1720aa2213d50bd
z20c37b833090be891f5a79e1aef75678b2ded62ecbfbc804717d1bc949e01acb07188c60428d4b
z28ffb845984682e32fd6e24ca8fa1aed44324b6f8c2cc14780b46164334abbe50ade7952254b48
za71d2bfba53c7335755596d0d830565387a2e8847680b8813530696b5556801221ebfd76f11ba0
z98cc8fc45e92a42e9b730dcc58c58fa302d44bfd55c50b4bd4b2a19255d05ce0d406fbef28ccc5
zb2dce3e6a9c17dcbf6d1bdbbeff044f8949b843f8ee01fc29da3c3cdaa5be86c44eb325c00b9ec
zb2bbebd236358cfa5a82d985ef3bafff9d09a5dd8b0397786eef3e358728f3b885e26150bb7467
z7e52606eead8b8a6bceb61834ce4fe454f3d4755161a7d88fc0116a462ebef2fd3d1484fc711be
zdf6ca0c173a30151bbedeaed71a6c65277eb7c191a4e7d10965974688387881dec46467aa70fe7
zb1368d9ea1c4d27de201691a67c16a5a75ae80a1f1f78048d6f70bf910adf533579d80d6bb20ee
z3618d1dff05dc15caf006af61c7311de04dd544595c4202a2ee67067f784748573e12e89f6bb0b
ze160eb4371f56b34603b17f5a2ebba9aad5c403898a74fe0efe1eac61c135342cdf5abf411c629
zffd19d819728307acfc753c513f3b30da58abf7b0b77c252d790251368654b41a26c02cd8ac315
z57ba496481083049a8e4c2e7657dcbb0c203934e5ca27d0fdc953c0a603f8a6a3868a28551676d
zee39cebaaef86ef13a3307058ecbe672c5c764df8e592dd097013b420d1131d739bb233d8f0dfd
z0bb8ff076261a00719148de71cbf8c35a71872c0e86c1d2840015a0e53bd9aca86e1bd0d5a622c
zfcb9ed59795808e8e5a06aa817c67ddf0c30c102a71f2f19d7bd18ef3da338e627cf4012b737b7
z2d96577ea0346c19a1ba84ce925bab46c4c316200161ba9d5ce832369ba247dda5c9f237c6ad93
z5eea9681fbb88609d0fbc5306055968816499713faada5c2cb991bb3cd6be73c042856e4be4a71
zb7879b9e9d951b17fed9f05522751f877ed2ece29ff657510b81bb2c9b08fcf3ee85a51695fea1
zbee314a261ca30483f260df9089da858be4ef79f643207aeb8ae3646752daf1355b715f3f56d8f
z37247ddaf0a0f626fb9395d753f3f920000113f1c876e045ecc101c20578e728382ee22d974b4f
z169ce73ec3f6d445186f32234f4a8610613ad2c3999c93747cef829d439bf63e49bb1d4e29f057
zc1e7655e24284dfb00e7c5c644dbc417be23a243864bd61618382003d44872f655fd018c08c91b
ze38be7926177985d9cd6dda27d9dd027733f6978587dfe9929c3f618f90126a5d172f27535706a
z9d10aa3dd55f248b387f2844efb42a0537f159c0f108f5ef5ac1ee50141938c5133e18f83d8815
z808a0b9e1ed97519a7cb322d8a8b6e6a427ae0b9d189b04ea504dfe0c225b34c4d9d38accd1472
zfbcd6374360ba6a09e7cbdd0904bf6793053e795945857642b7f7ef0932b719f90175a3525bc61
ze019a02bc4c242c9c473a81c3cfd4cf381077cce732407646fa39cc6e62510a016272418f4e291
z54cd5b821e822ee1927a8b44da8e4909a979b17fb6ef4bf75d416a6ad612e1c004102860b48666
zd73456fbcc5ab7c574e2bf2dc47ac0fd575cf4ef737de68b102468660ff4c3b4c92996042d7df2
z742155d159c61a4b765507ec2b21ab0519579d5ebbd04f4b88e9610593d43736ce82cc594bfb28
ze701298abadfc3fcde44c257baf5a5394128fe38161913dff2655e647d9b8d6d573ed11ce634b2
ze53d203bb797bf94b0e7d75efc3009f4c4e0404930fb25535eb215e97070c80b812c50914f0935
z2e89f4f0605e95ca6b88e066f047eaa430e6784bd8e74b541d74b75f448a7d84d16eedcfd8c0fc
z38bc3baced480fc2bee4963a1b370ba7f001cc6c2de0f54bcf9869a230d5ff34a702ad90a6db01
zb6fe2264cd1665dabfd8080bcf0e3c3f48eb2551f4558a91950f478236ede24b534622587c3bf3
z5f2e03a9ac7744e61a64eec4288b5101901ec2239d915a50998a66d80233bd575f8acbc9a24720
z14d8e78f9d3508767e9a2023ae98a441cdf82cefa103dac814829cdd46126aac251993df9610f6
za9a4e2088c27908a308ca2580967493d406247cfa6a90ec2927c974a6c26ff57adf53df8567461
zdcaa7c774fb6b6100f57ab0431f74e6996ac450f6265c0336fa8eed62affa12baf789dd7d510db
zc714a4a369aac428ea64d29e89fabc59c637784669f3a34da33a8fe230df0f7cf7b38e495677c6
za477ee00c22b3ab890129cfe3f22a857b76c62cb34fbc6b49112ed61be47525c248cd09004d785
z16017ce69ab787acaf513cdbbcceea7263df74764c1fb2c1cf118737d1d55ae9d7badee53c8d8f
zd727f6d9f51c88d9a36efda04fe133e8a7fa215c86ceab380e87e64cf2a537209b6f8d5a6ac56a
z97e287cc0dc2c39d92532ed4cc7d17c22d045f6d172f09ac771996a7ca121e578c6187f3ecd908
zcc1aed53130c2731795c677bbdcab12fb82041a806930ba0ead61764cbe1a563a158a7d70f3733
z818e39042374425dd047e817d53d5cedf7314313a1cbd6f646ff476945f47807d616318ac929b3
z202312401d6c0bfde9623cdfa66fa53e9002e2c2d0cc4ba8b285c91ac1d369f2fbd02521f4b72e
zd5554cb641a0d7a58c117d9165d578e82151fec8f16473d4d6324f8e24a29af1c0bdcf25385f53
zfb4f109aa899e2fb5c13c648e67cf8081775a04add6a5ff58ec453944017db4263a16f0bf23bca
z97632d3ab3f22416d217f1dea28ac660bcb1033d6d3fa9a163bd93c4a2c646c5978eb179c84064
zfb1d1e64ab9cc0b25e11b51b510fefa59afe656e15b153cd6c698f1f56e1923ebe69cd51baf58c
z63d8a2ee637d3fc7e26447f1fea6e6727327a48e96313ebee78d80d4d2d5ebf95ed7ce3e126545
z9aabe2c3067a3d311bc0dfbb2ec4f6f21dbdabba31cfbd50f6b0a322bd57736d81e8d251afce5f
z81b46adc686adb2c7f1148c971d3fa74b053756885e3c7b98de3beef2929265c0bd05e8a9bdb29
z8fdd2e84db9b74e4e5504c0b5a0c0f1cb48c6818422fb2a5f24529e86f12083f22ab2670a80bc4
z86affd90880dadbdeab13af67063e1c8aca2ffa9ca5729533e198f2289a596489ba4b5696e76ea
ze5459edc66a723075f603f4db868b15f32fe807c5688e446ea34ce9892ad3bb5cffc3ac978c316
z96d33f49438ecd20ccbe5989da5c737d088e6af329aa1b5789779700ff0d0f375817c86b2043fc
z0033a29f131acd415d9324c59b08d684c6b153a48037fa28a85efe4798ff6f1bfa68dd1494b807
ze6b471756327c3207f4316810c26ce5e4506663b76082f245242fa6c7c8c64864c5904ffedf57a
z20e7191f4953b4012fb1ebdde49f8043f5410d7db065bdfd1d68558c7a816e8dc16e33354346ad
zf7299ce6b39cb5afc0ed45dbe6961b9491ffe90ba188d7e64f17217bc8b68e6e670426a320628d
zb91860be82fc48cc834fa2d3fef63e5db1f3bba41fdfa0623d15247089e108014aaf678b47a47d
z17f044837275219e89fb3c268918d293e59f997958321113ebd50a8c61ecde9e5faccc93b9768f
z286ecca99c32e4e349ecef393eff4603ec5cb4581d218ae2fc28010cbb8e5ad49ff58099e66ae8
zcfd0ebb0cdea8f314bd337b0cbdbae2ca69e728995933a6b5fae335a34c5db98379b4b0ccc7ac9
z7c9567168fef5d07332d54d6783468cdd00d2a9248db161de703a729c4e85eb9fea04909f25802
z9d2f137e588e3606ae32d8dc5a739ccde3a3e397a9177aedbd0c1e9144b14918ece3a9dd996101
z0bad9bb08b8a44f575d2894a780963aefc922a7a7636f05a1786ae7833f758d041ff048daf5407
z00d0fc7e035d8db81345acfbca35359add535a100b863aead325a8857cc2c8230119c98627934c
z614efb7257d3335b7d234541ecc2b1aef6b180a99a1c5a55377b8b4a012f252d05c98a13771729
zf1aca56ab8a7f2b038184b444b735ae33b147e1ce07aff9f114f588fbde8ec25ac212cd75b6abf
za1a5d65e65b2123fd8ff8319c0e303cdf95fd2a09b885f6ae7ec33f08a79ac99ba2d0c7e29b761
z2c5fc23477e5867bc8b6b79c42989d8f70c19d57265e5b73f00d07a2f378a0e967540b3e0c3b04
z9f9516343f1b80e2e9548c92b23f8068beae785316220a0dabbfa8cceaa5f73e89e1d044bc5b20
zc91932142dc325ab42f886637b21a0b9f7206b2abad9f853397f554bb5a2b7389ecc348980db40
za0289479db09a1ac25085cf8dd7e2279a64192bc6563974fce2c1cb7de6e29e194d1aec189d959
z18b2964d2483fdd64c888daba5d4b01d95a7be46d7c5943917090bf7084216b68abff5bae2001f
z7b0da14dfd62dd0f94a665de97a67b013386bb04bf01f716133dced2437a5e9f1a61a4f13def26
z4700537febf7bf4a942aff1ca14987fe469c35406cb98d4e93d524773fbf5e031014d1ede2658f
zd56f355eb964afb964957045b5a18a8972be727cfce4b7bfa5898d829fb97aa5303024b8bf34ec
z733a6772051d289574db805d66a7d1a2a224e55d581d8f7c11efb04055953e5ac855e5e44794f5
zae6f9efe346b10fe001ddad481fca863c863a3327372e3d8bec375d6d6e5087995c3c59225a51b
z8f12b30a624b49bc1c0588069fd8da86ca488e50d05b0578a696d4f9ab4d418bc449984074b210
z78a4e4196eb198c145407920a3b80b8c61e2aa06c016eff153a48e6cd826b99b60f0ee3fa86cab
z807148657f1c39883313730f03becac7a134bdf90cff09b85d758347a25a1354be1ab948947f77
z9978c7e96aed8499fb990f277e7f14c1b56cc8f17d511d5104788ae7fd5c1e87792f6f688ef924
zf3005dbf5bebd45c5cfce607550fd60e07fffc8d80ef7857800c3e1eab620da037f679c0e84caf
z1aadee8e9ae385ec16797227fe32035e39d61c5e2ddc53d16d32f2207aafbd5736b5655bce7118
z0173fe3f00f943f3f63b769141e69de565ef0dad4c2b9e6cdd68e48a4364847578b0a8dc3e3631
zc9470f05d1c30da02cceb59171b544cfa635584b9f0dda446a08e47f4c0486e0fc8c7dddcd356e
z394c2a6d47e2a808b876458f9c6c0abe41836b4f2ad15b29e40785da1e32357115802878cf152e
z316937e692897476ac259a75ee6363e1ddfadf1700af44202e6b62b316b9ee31ca4df2d060eb8f
z01c0ab54bcd95b45c31fde09c113f249d775620061af34dc727274616c55399a902b9aa5fe429d
z60553c72eada116c3e614b68f315feb708daff6bb9d6ffd5a128389d6b90e85fc46cf6db68b34e
z2fdf590f4d54fd1a602a1bdfad8ff3cdcf0f166e0a4cdb4e4bf2a81765c0a863aaf3eca2c5f2e1
z5dcbeffcf854d7c84628a2b06207cdd3cbb1c68f23884953809138d1787b5b0034aa766a6af58c
z0fced48bbd8b605b63586c9711ff59bfecc484b68bab993e86fa6248aee4c5cba6ead15b88df5e
zc81b1cafd1c34f1d9007f008f1bae7236178dcb52fcf29541ef77c899bd3ec88e7c9e3717d44af
zd4c8285d43e710437fb315435ea7fe76dad420376a3c963a7a3a82e8963a50ad79da8a00d7af8d
z8bf46fd1ea4ed0188cdc2b8450e79eb3f2f84516775226b4b0d372e41319017c42b19172a8917e
z5d2e18040443f9284b22d4edd2715d17e74e6712cea2cdd547cbda5474fda582c7a0ece957c8a1
z27c7115285b26c3964ed42fcc83751b9ca06c342f5456c98d82f992bb0336a92448322c1d81c5d
z93aa645b1ae47651acd2dd13307fac82cfd8c30498a69ffe30272b153e146f66b9c6bd1e31b922
z6be3e0823d77c4733b2dc3433d8022a1f39e6689eed834222c9bd45fb41adced3a6525406ee110
z578fa898ceca4b59be7c96051bf96addd8a7b58b478417d1f1f7cd983b37eaf334950af332835d
z7cffa93a1c4ec126f36097dbc855ab00653a64feca0a47aa262d21feced83525d6a57c4c0f71de
z28999c2d511d6cd8611ba3eac7ff635bac20c9349776ef1683b3896bbdc1a962d335ad635f42b8
z4eab633a41c0c4455f90722ff6e794ff0078d5076596fc1e5d2a990a903fd76e0113d886c11a93
z053f421c8cad48af3cd27e9feaabd4f17ac38572e158f5da6335242d0a190c45a89111803f784c
zc6f6720438f2e2ca1af5edc6e96e3bb6583c80724408e0f37b3f12ec3bddde621c4f598f17184f
z3caa04e58d45b4963934b36801575f3226b3ffa2db2094258319e54cc0456c686d482e5b59c2d1
z08024f72634f3de6389a56f9c96fa41aab073481262235d20d5ed62305acc27d02203a4bd81ed8
z05372e7007127304740f301f4dd96bb669da3713d644ca10b87ef9e32bde4e50d5de3ca7dea04f
ze7dbed6591748886113452955ca5d204a85eaa43c79432bd05518c559a54f9a3bca7af85e0e850
z5f693606bbf48f84b59be6fd7b395df2c0ec6095eee12f132f91211bf322c69efeb1de2235f6c5
z7101ec29e511fca207648b0639e5b4df1e9a71b71a551de35595772d45f7507cfbf5bf1509eb62
z0447e3baa4956a3b3b830735ee23be08f2d667bcd543a63d8371dbc4e88daeb06c0ef315502cbb
zae07dc1357a81738ceed0eb8127aa3aec6c4eb875dd799b01632e75153f708a30112501d2d392b
z342c76035e3b4543e0aae45c136450fa62f8c53c104064c897f0a5a163ebf34f5f0af0eb5bf4ab
z35f5318309f32782ed473b3c4d870311ab20c5c7017ed74c9e5c291dffeb0b48ffa28d163d766b
zbe2cb879528c4609f34315e00a731e951c06d7bb6a1d2bbe6713df67e4206613c9f912e95ed5b3
z44ece55aadd7e3155a41fc0b2654ea00060a77cc30c43674589d6994314495503dbfa0a9937383
za2071903ca98252d50a949b77f1c576e3d7a80681950cd6a8a646b321d060a25d8b0eb72956a0d
z8ca9706df85d2b8a1e76d7f7b1c05477e1d1c49d429588d4faac24dfabb861572ca7ca1f6473c1
z381ca09c81350a7a1d0253af940253d5173c358f8a8e647cf604ca6baf64ae8e6067e5ede901d4
z45cb942408623ed56d9154049e7754c5861555a6ad97670c627bca23d49100c5c4c364ad5cd666
za1a1d72392ce33edf3d301e8cfd5328d375e780e551b0d1b8288cde71ce17387cd4acd74e55028
z3cd155ac986a044f0756d3204c1267099c96e32221dfb3c13ad07b325f515139972f13de958357
zefe67c45ace32bc24341c19dae162aeb15b29e3427e51d73f4cff84600c36354928cbd1861573f
z4517c6e864be9fca674b782242dfbaa088294fb0c6e192a76f803d264a775bcbbb1660a4985bb3
z8770359d6ba4e16151a02e4c61d17d44e6d095f66e3c1275adc266efae4d44bdd955b803bb9059
z5f852972f61dffd545cc252e480739dcf7c4655aaf8e944fa022ad738a4e1f990914eb22f7cbcd
z849b4457c9566e0a266525bf9e4eb6e70978c25745283fcb56498385f72e70451d372d186554b4
z1c41871d680c2a55be9697a9d5adfd85d12bf4643e3b80fb43ef97ad86e46a681f7268adab75e0
z75b05aa2c375b37ad953de4331b48660d3046f8360aac7f2912e3572dee36083f8b8e252790be2
ze6ff0c6a4d98c7bd1736e024eb9abf5729066b9a6903f4907dfcda3ba3ac6b79c86993a25f071b
zaecf081bcd1562d915c60ab9b6a6f2f0f385280e1796f71e9626956e6391cfdfa485af9d62b4be
z0010ea7d3188fd6af89ae10ad0ba566a1db23e46cc8de35e23c8d97c0d66bd53f1b6d79c28515b
zdf5c74319618f375fbce3eb8d337615e78c8d3b5b22a7603f6d2047c67b23b9621d07b8af99706
z797a62d171cb06a4aff554c14fc1efcaf485446f193fc93f97b4ab69a48e7b588f80548ef78ec9
zdec39d9e86989011057774f4e7c700caa833f72843c9f087019b162d2f934778d355be95009d43
zb5c98b95fdcbd54b2619980367f15203d0424a93c0f4a0586226cec1ec8489080af2f09724e78e
z9c0db078a4a9fb81d239a4c3bef6d7776e00853fff61982c7a57208815a935b332ddb87e784cee
z42545962b89c97ef3ef9150f79cc834f095e95fe452ce25ef09373df97ba2aad8b765260ee0e69
z3a52e3d75f8d6a169c9074c993c98485cf6d820742b05681248a383f185ea62d45dd00d017dde6
z681a1c35a7f5948bc90468cb6098ecf788f97299f11602b121c2cd56b5e4eb1592742a208696c5
zda762e7c79aa3bd2d6e4008a3f1f4d09114dcec3e6bc86d2b9596696a5159b9be52b55ac9b7974
z2730bb3d0c371f8644fa81698107f480d9b3b2fc1b430733ebc7eefceb306a19bfdd948d82419d
za212aeb30b209b891d25f317bc7f4a93525106c3abd50587f0302034124823df3b440c5a566b8d
zc75ea490e6de241f931b4b7bd8540ab7c8ce4f3ab052f5a9491843320ba1ca0bb673d9a83c47e8
zfd60d5bb4655acd6343ecdf41fd7184a1945276de044cf617dfb19cc7f3a081118892c89a366fb
z9e3ed522efa18852695126dddc1ca5acf92778c209bf37a78fb452000ad40bdf5173395a37a5df
z30ca27fd830094434bd3a1a3064d39997efd680fbad6aca719736ae838b2b14cd77d69b7070f9c
z9789a21c6372b9a3d86c6721448233e3f46ffac43bbc3073f37a15f755470e974135e1e46ab339
z8a973c5773cff0a69c724c990c6cb6aee8a0e6ca918744d0caaedf7998b08905a50e5e806a5157
z32ee3553845dfb2896db00d4bbb4d7c8ddaae825fe77ac54cc0e2e29fbbd2e54f0c8e40e23c1d5
z0ff48b290e5bb77431e00228e6211b3111872d0099c9379b3fca6d4756be493f8145a5997dad53
zc60dfee61d2d497e2e93dfac30e7afbd13a6e19e1a598502908963cbee0afbfa731378669dc013
zab7777f10201308d6ce1b1c52f2c0d4d46f65f20c7527702dd0c3fdea51c33c272c6fb39678c81
z48a2fd48c359ccd2d2154ce69bd8c2b458430d820d0d818f2b2ce5a2f229e952c540b333c0601e
z42e7a465412e3e0023a4b1759a313b215e7877aa50ef0375474c0785657a950d535b831ab5a2ab
zb966bb136fb576ab24cb26dba733f6c233df7445ba2126971a39ec8ab940642637528594a77620
z3994bb9bdaf145d969fa2c0df0aaae1d43ca054dca47093bc77c5ff4fd3292b7b95f7d06668711
z4a5ac71e5546e1189401931f2b15c4e6923912124eecb509baf1478477ff4493c45209a988c285
z222e71ff9e9472cb6093fd1995510dd8e67cb52926d7a35b271669bcba08c53ba0b1d70241cea9
z8e3440ccef23193bcc3f075a1905cb743f883ec7756bc15b420adc781ff9d2055668a5e80a6690
z2871cd0dddf42203164dc3c244b61aafbb350343aae597ea19b47fd9dc54b5d6f24a43f864c13e
zb4c2e98393a20c9bb4f3dfbe1bd579d53c0d754c910483f93c92acd9b6de7234e07d4f2170ab92
z3375e495b4dfb12f5137cb29973d61cfdc1d705b85cad1cd2012edb8b309ffa9fb90f1e833b11d
zaad085816457bc5adfef4929f074efc20922b66292bfe3edfd1801ed446c5a07947c81d7951f40
z110a60e266f49279854525eea546e0d46ed482d802271d6a17650f7eb3d19ed63e6765ea77b450
z102c4d84577133b30d53dbfee796ba42f86998014ca53a18a4f6c11fba4b1495d267ed9af8567a
zab4895da2fbb3558cc28944a9271d9184be9cb685ecf1edad058c85c70dd3c029ec97691737710
zbdea3a6fbc44ea81134979f5396eb0de9e3754db9246d39dc52caac0a1d56d209c1645259cae8a
z815059d7ae81242e20c1bc6b57a1a9dbb01d3b0d4e8eda10e7a0417c42634f4b2e202c0ab4a6e1
z2023edeb4731c56aeacc715e6dc4490dd8a915ce0c875e3333c5b46c93385a92660cae4909869f
z7ffa48e52dc1d8999ac21e3b16500e85dbfc6050b817b69f55e89aca4caf57c731dff4f87a4871
z40957503b66b34d7f68a27e0bb620f4cd1cf61f9065feb38179133c31f7ecbef2fb685705e4ab2
zb8597446d9acf0ffc4c7fe788ae8a7e304b7e8b707e15f1be0a2818eef6022765c316d4315e179
z3a9fa18555316b5bca742279de7a4c11f690fca4b1484a97d0ac7c9c5f8d2899b73b068978888d
za1f8ec8c06b8fd8b66b88a9f8a97f7b582ebc8f879e4c4f0fa600d1cf5cdde73942fd484fe62c3
zcf6d2d4a002fe5ba2244f8e3bc01a6077d71fc4690c86d147f3d020d11d8c2008af40ce8ef39fc
zbf94a1a32fbfa4b80b4a208ecf1ab1a27fafc684c2252ab7a0514dc7ae23d2d96988e518f533ab
z0ed9a0b3f1667425d12588e7b2f18e49f7d6e8aa10576227885c919e5240350085034557d9e917
za79b15484ecd6217fab4cadd23d6f2c5c2f3adb134f64b69af4a578031c195603c93dc8999a5f4
z5f73da03f9e36ccff0639f4f034a12fd5e0cbdc1724952a150b3fb9b8d018532645ba72782c5a7
zb0d3dc1d3233ec5967f0342e4c4c6795a51129e9ade81e42cc5b67265915f710fd3f6dffe56b82
z11aa925dac5dba6574117db482715be98bcb5f941cfd435f23506accf6c82cf9548fedcec1d138
z2ec1a89d2a5d27d6d75c30cd71c75c8b3832ddcf3ede9517dd2dca1a01d6a5b6222348ebe676f6
z38e383b02571bef2366ddd6cec0707866f9150b7157cc6b6d0320df4207376d0950b5e29f8f0f8
zdb9cc67927dad1695808ed46a4dfae789e7437501411fa51604b3f905bec4f81b91c75dc5ab39a
zbef74973475414cdf076b64abade853902f2a854839b1b67afb2653a87ab16810b19044a1c3749
z32494d440792fee2f6439903da511497ed45e2599160db38de3910c1106b408055994d4a59e50d
z5c3e6cf75baa62d42ac0173da7536448a98febdb54bcf4cff9fecd259cb5ec040b854bbebf4172
za00e42353e55cf3fbc5ff10d7d7172da112424d4a80531cd3038ce547b7ca7c4f350cc4c16798a
z2282a2b90ed3b5a0197a9bdfaa2a01b13041092033f2f10af1958e4fc8f7c6de2ff719975ac946
z777ffa2ed3ca90b953512ed43f1b16082c9f9a1db7607cbd32d19c957c2cae9b191e51ecbc34ed
z5b55b4c7db2d38db0d802d8be2faff7acf81f6c00a94fea7ce9a622b2209bf87e40c4c2fc76cba
z458eba2dd3e025be6cdecf88fc84429d122a8b979ff7aedb513af79e2d76672e5a5e73d05f7959
z6d91fc8466c73f349e1204538ee9260619b8af2befc80f1b2b5bd7c15a07c241aaa34b590c4223
z2da2d27935cc674fa5695a37087e22e5079f31f4467666a766de77f690025b605dea12658fb2e1
z7b9a6856f45486fa1ef83497f2afa56ef9a9cdfec775dd83ce9386608f76ccd6e2bcec069110db
z7a4cacb57905df6de87c52ffd69b72ba0e641fdc5654e5c6646003fa54e4f72a63c72ae6165dc1
z0bc4d66b61c55003c26bf64be6e7b53b3f479467620b4c98c3597c0ec24da4151234c5e5893d91
zb66386a13fcc4626bb62cd30aafe23b6f2772460e47a8a8172599879636c535d5ccbc8ed87c284
z8a04ac9b6adda8caee5d1992237c9e291b7fbde2cb1bef163c28efddd32aec2b9cc643691e50d8
z03fab5d457e5649dabd00dc24421400e7eed920c97c9288d6d2b9b86c298bce5bd11744316c850
zed2c4b0a70961e28be41c5dcfff240197c34533ef46cc75713ae8fc41977d0a8c8fbe14ac4fb1a
zc8ca4552d6f8d4d9f1fb965841752707f4c50dff6c5e70bfcc2d7d4c9c3447533f8b3423faa0a7
z14656815db9a75cbbc50fc6fd33e96474c1679ca1a926717e783a068e07d21a848765f5d2d651b
zb783b679b674dfdbe28e3476d92b66707ad7355bb54f704bf9e0bfeb2a56939735aba485b1df49
za78c4a6b6864db531bd5e0b811708858b8c5d8d34722143aa91006e283dfb0beb0820e66aeace9
z3f2758b9ea18877ba8b0dc6f74ba94638013b711d640253b997c28ede4bb72b8b4c4f7253a8fe6
z068752001e657a7adbf04a92a91243322f84c6a8a7416003ee09d88bf132c2eb55783f03f52cbc
zf291e955822f3b9a57b19cde048f5dd30eba4e94ae1cea449758171f4c9a764518c9ed2d3f2e29
z19c3aed64c57fb79094e8f85622b698a97e9b810b2cf8b591d658860d15959ce3e051d814bd969
za6e66714930aac14e9f4c15b64bd8be42df060892f399cba50cca1173a18539fe945d5a910dcf3
z0d1e2cc84adf0ca94f771587811cdb2d300b59c37e6045438177938175b545576e8112ab0247dc
z58c20876ce294c08ceac92f1386510687609fa81737ae97dde5e5c8269d73d114fb85e2ad0c157
z34a835021a357356aff3facfcc34643530eda0bd7e5979bfa40c11866f74eb9582bf6f5cd715b7
zd00f3a2d1d8d0eeb7c6ea76fbb48975d9412b101fa4b2530b8cbdfef7491bf7855eefdd1d26eb3
zc155189dbcd9b1426cc3381adc314825f1d0c12e11510b5b1bda16e9019ee8c6bbb1087d3c5a57
zc010c98ba3a8cdc61b90eac560f7c0f615f281ff794883fe8e3e3e26994122677efd092f66006e
z6c5f29534bcb1b310d2d76ecf261f27054bd5db54b92b5db2b970b355a284b55eab6bbdefdc54d
ze71417f4d6667a4dc9e42ab580e7aea7635fc4babe7ffc4e068fd20e4facb8a816346de6fa4c99
zfab49b8f7fd6a3e3e577e6b553c6b425926785df45f3626ed2adfaaf0c55585bcf6a77eaecd99a
z168b243d7a52ddc8dec95a3730737447067edb28a77f3fd2d952c55a3f0f0d91f9c2706b41fe98
z3170ec2265b17a877d9312cb2bcff97e891a6710a7f74d4b95552956ec7433c435f9b7fb9ed0af
z98fd85fabcef1c9c4e7db04f7a5a00894383c36e8f2825efc6f49fb5b940c4edf752fdd1ebc2cb
z99e3f0eec78906b48353cb177a1499bb03a6a8ee406dc72c177132d4c657ef8c4fe6fd93f5906a
zfd97313c7f0cf3b69afea1604d043193208215555c77012ec1e99e68cf5404188bc24291f2f750
zf898dad9cfd3b5a27987f4c0ca0066665afeb05603dc58b51ccf1e5dd7bd8fb052f210fd6ff73f
zd9ce55cb902e52d2f5715c9b3d2b6d8bb3fc96db89d39c28d1ba7955cda7fc88ca41cf7c00a87b
z3e2c0a7f98471ad9d4005c8b4e208ed7263ff9c8db150f030f7f84c193e970528ffe8293cfb37b
zd0b9496b83c8c10c28b5aa051de65606fdcd058b7927e023acc3b62921c4e0461992eeafc56ae9
zac1c371468b3e4fc8a0b8614adb2e907c975796394cb76838c8f126f42316ec262d62aff24d47e
z94e30b1a7e34afad5215ea06090e75992e6ca2c3e1ee20abfa2543d0f9d78bf578b77f3dde3b87
zabb42097898d4e75c35916c608458626774561e3cd58f72a7935051c41a4e8b489bc9826dce710
z5ee0933dd1567c4a36cfe7d0cab3a82c0e862d00c6b10ec47eb398feb4e0cae6865833990beebd
zc2bd4592c748d5caf0e0805cdc788ea0d72e5cb898c8991bc86d5b28bc6a7464e046f2125143e8
za0b5ea7af7e4fd8c5f5b0415371229af44e2ad12ad1aa0bbd2d99b94b83494cda6de163521cb66
z55dcf9f9be8e118c8687ee007b12da5c7916b616a45ed7d94706d877aa6d1bca82f5f8ed3e9b3b
z1cef56d08a9ffc5c8ccf3e5ca022e1e668aecf0b8b93c69dd30c4eda6e81265a1b81f1eadae681
z16710c93e191714b20e84232b1fd0e7bdea42d52d3c17c8389a5749ea44286cf7dde2438ec3c16
z2ee385976490b23ab825d20b58eddfb25bbf8a6160140404cfe9b8a6cdb6b7b67a16d618f54478
z34825b67aea2ef8c8a0cbfce38f0fdec52d84d8543ad7ac8ab7a50926be3450e5d9d050c653b87
zdf90247650fcf650d85f9641581b9a2b6a60084a79d11f0e6748e57c2dabbe378c6586fbb72bd4
zc6246073316b68e4c875f957beb7599e51f5108d762a5ee4ff2a77ca4edf8133a3a7bdd71123b1
zbf4b34ae759fc76711777846287b1bd66993335ce5d8c794e752efd76171f86e64867179453d27
zb2469e57c408ff8958519ac79d03952602ca6fb34bc4b80ab699f6e73133aa5d662a78cc10ff79
zfb00a2fb534960900eea4512308957fcc3ae7ba1f8eb639e068e982cdd006502daec9c15f2f0dc
zca99a1df19140dc28cde25d9da0dc74d248e56dfa3420f3e0afcfdd1bf4bdec958885292e26c74
za279c3e57830c6cb7c2af70648b4512744d1f5e68e7493d24e417234e8befb1e5e72276fa85a2c
z81ec496d63e641592a6cd1276b983ae852edc2288e68c69b7017611304ee50864822dbfba1a8a7
z6fdd17848f145341a9626aaa1f0fea12983c6419eb3f5d8c11f6f646583358229317053142123c
zc04b15e27512e22b1ac169eb534599d92934a5290dc4f1c35ff1075a9237c8d5b7c5cc18ed43b4
z8f7e9fb6d17dfb0193fccadcf1ec0057df6eaa249711c4d5e5f18bad11969fd691e2d9fcebe237
z4577ba7e2672cd1eb7d6ba7a2a8d8fe0edc37efcc1285556b5aca7886fe774efd570ff894b49da
z1ec8718e231064241044128cc802f8f690b0b323a2e8f81b0d810056f32505e4836763857ae42d
zdf835e64d79dc7ae1a0208c62982828ee097637826b9cf66db36b1bc151b44f0a09d97db373f4b
z95acbd71c6cbbb01614be888a724acaf639a0b148ca8a34d749ffe6c920fde0700bf4f0dcb7c7b
zd85f054aa12d5e87a18bdfa4836e5717e8e9ce21577ee27d4f885b5dbdd6f130695ceaa1bc8224
z10009e0782110d268023cd3bcc6b49ee4a5f4ab9427da58fe3dae6eea6fa753df33b18eccb6e6b
zd3eef8e1b67810ca52802b90f6801de7b22f508c4b3158b4de69d3667fb53d9c5ac1f265fb40be
z4669e1ebd4ff895f410912ca610d5b84926a8a329315c0fd34ff9d01509a889fb783950ddd0afe
z4c44cb48b003cace60e751e42d5a29324bc216bc933909fb886117d742a4423006221ad6ed21ca
z6f294b301402cb2405fd177b248f7e4109be5c9fed4fc34c9d9b0b67e61d038c762bcde6abe6dd
z95f76eec5bd7ff7686f529f777de595ccce61c4293c1fe198690e64843030155f3afeb598f2fc0
z5f16ee94789fabf0b120ac75c5b0a5a0085c0f2b615a2523ab5a3896da46270177f1c7eca5cd48
z4bc1a354392f10832f29c6d5f465a35264be42e991636d19e3cd5f83bd6d68c249b3a59fd0fd9d
z9088cf4e066839edef8723e3c78bed15519d27d1f551c628da17035cded5d7e326aaf2c21f261b
z9ffc4058b660e14ef0e372aebbd24084c428f168c1623dcb37a31af96ef84c1d54f61256cea30d
z2a86566fb2b8642991687c4af42514451ba7912fe9416cad53945c0d75fdb032e6948472f21710
z4b8895273d66cef6a2f16318106b1d8638237627cae4779fbd56e494f6df826cc747b6b4a929f7
zc95f02dc776012259a40b3ead201600c77b22e287672118ab75b9cb2d36c038b1c9515148113f6
z8831b20b167839acaead995a1d48c4ed44acb24bb0bbaabf467e73638dc00fc41b37a717c3b4d4
za48083ac1287288486083deab03358de8a16f7dce635ab0772cced2c173bb33e7e8f08a40652fc
z33ef72e0fc79c839d6b5e1c8ca4d9c1d6687e1e485a2b6401bdcfe3233ca36dacb2b4e1f808e0f
ze3ff19b09e433bf6d2231940ecb4dd0bf3f620f6a9b46855c225f8f362addc82a45a1c6307e184
zdecdc109750454180eccf931a99830e61580ccc06f697acc57c4c1ee627cbf6898ecd7a326669b
zb7e016a973e7a219d5cfbbb0b196a1dfde88ca3fe86ca67e90ce090119489b84943355aeb27378
z0d1c8d60e9081dbcbbbee50cb5735fadba5e2a9be35f77534fa8189992807e2961dabfe8efc763
zebd75eca93a3c432e21ec67e8c55f9536ae9cd7a0283e7b83eb5f69aa5cb1c9f6c89b9f63ec941
z9bde17e34b4261d0ca711c4f69109e868bd9fc2b8a94044bb13e0c8a3d8dac2825433a7643dfa5
z9fc85c469beeec7504fd6392707244263a3bbb70cf5f6b8416c1db38f14832cefd9153cf0574ed
ze0b804bf2119c852039ab4670320bcebf1e366005e8070f540b263bbcc7834372149707782a57d
z4ee17ef55582ab7b31538ce44a69de641ac438e0cc513e665776f7a48877507a8d46ebdd39a746
z5b265ac187f1495f611acd5e32f51272f1db95d72eba40709c269c0f5135353e7cf5244a9009c0
z6c553a20cf332701d3c5be978c40f70e45e9b53d7fb1d065ed091916eb042c9f9e5b2c8d83adc1
zadc5650dd62c9878727c8a7058af7ca3597cc2337c2a82197949d6b6667230f1d130b261060025
z2d6a976323ed77f2e0a0b7e3d5df2b972e6232f27ab4ef62a14e3e40bcb358d5a1e636684cff42
z08ab16fc68026c3b8ec0288a3cd7c2c21bdb254da2a95c2db27332f39bc28b4aa246fde2caefe1
z3952af177bc745ae55a422c7a4c13375efab13a53673919e650c142771af7ae20b1a1ee18bfa6d
z1f79b8369f7e9ab5ee5fd53d20d587a5196c7ff617c5c022728597c778d475e4c95809252d7991
zeeaec2852df9cb5c66acfeec306d597b9fb1ac8bf30cb49b5c74020367f92309d7b9650fc21f8e
ze95e3a508280ed24a4d8ec5492664ecd37da2c17e869adcc25c0396bd2f490f2ca34c5ee625573
z28918253182b853d051bc3776c27d56cb0ba53171b46f379af13618acbe3e1f3af91ce81135ac6
zeed08ad154f8a5f2cddd4e3d657cfcc7f480f480a54036594606fa0ac03439b1dd835bd5bbd0f7
z52ce0c5821272454ef2eebd82eef01323c73d7f434f7073c1c84a43a14045d5012eead84d0d874
z44283ca36ed11969580dcf74de0f029baed339de7e6b8681d8eb19fa2eef4295de92881f4f4510
z9cf2c65066970e278e885ddcfa6690d09c048182134b33dabb067ec4dfb49cc6d291a8941ab57d
z9e23abb5a0574a87d371c60aeb2e2f77873a09d61af523494438d1e90e9c3b2f72c196ce126774
z3820f39cf273379dffa3a8f89ae6e40fde6287bcbf555c23ebaf3ad70427bb6d319898608ec832
z4d14b92e646c41bf1b568b9be74805caed53b463857dbd96a558104e8b90cfc1b106d3faa2b5c0
z55a3ffbd1315295efa1b705db551dcfbdbc1dfcd9f4923602573555a7f25ae4a20495b345ddaf9
z5f784db79c828d8a14cefafd94360a022e81858e7dd517227fee33e35e78a59c8258961bb4dfc0
za70afb74871159359117a718c71f49c0cf60748331921b210b1ef530653654169065474741a070
z0e89eddc64015c63d6263c755a052177c68704a08b3c539707773046c322a588408b9f3e2789a9
z3b38f050d1612b560068df5a2773c2217b4330871a6b1ba5369fd5b9c5b91430e8e7e9ce234fc3
z552810165eea6e8acda37c652cd587f4decc70eca9bdea2af31295e4dfb7fab8e8af9096751e74
z01f7b0ee1bd7bec3224b5356362469fa1907590ec3078e382f1f4a9fcbb3a5735de1c504b61383
z598803f112662d554c17487571698c6f0e2b5a66dbaeb725d425fcf58b9abfc848bc86d7a26925
z1d67aa484eecc43530156b1ab9faccd54cc3e8a7b034a267f6ab49fbfa210e9b721784865dfc3e
zd5211d07ec1dcf69165e6209c8f26f555de48e81f11857d6a8462046f7a81f9c93c8fb4ed40357
zab4899b33055a6f7513fef32586a8941d423d7f916713651855256716ac9dd0911d5ae7b556f6a
zb4631473338bc64ec26521b54def836898aea051f0f0133d3c37cf6963ad818f021dc98bea01bd
z9aa20bfc38d58786267be6789c269e785f07b2388a6b3b6677fc646aefdc6d48776b52d4a28f01
zcd4d7c4fbb684541e197df9e5972e2c84d4ab176322991294803d3fd5a788fc1b3dad7be6d3a75
zc1b0c295db4eb83eb212bb3268eaf6d37ef457b141c4aaa01baeed7a73be18def0493586905551
zfada8302abf3e7e653d285308587809628744abe6f0e118881a72d15be012261301120607fd15e
z151c98768d3a1c096256683b33fcd46c6baa8da5d7ee1169b0942d108fb3ae17d8aa9fab1b124c
z899bdc7c3b4afef071654ec42c9c5f776df1d7bfafaa54b080de5d124c43df7bb27a9ded444391
z6e0e86f9c6b2e22c83292e669739dd0f8411f8bfbe5274cee324d1bde1a4b412297433ffb3c77e
zd796ab1622613edb16c1312d1b43e077820934c82297dd4a02201f43dcd4cd8774d584a05ea98b
z72f0b8e2b0c6b43466393fa6039c7cc891ed8a66bc8be228f2924d1363766520e3a8025fce006e
z9f36fa9a6305499ba39b5859f0df107be92a6d952355a96db2a8892c63f0c2d2a4a69c13e1b12a
zcbb51bd4ff5cf9733c19d49c74639015720001fbb8dc9fb6e69553878d94b7745f6d5fc091b885
z4791f24d050ea1eb69780af986767f4da738161822a7660a54c32224d51a8d1bbad146da70026e
z7f57860798eca45efef6218270438d1121863e43e7c34f7460d02a1fc0aef49d1b955cc18b9995
z6b97e78716a18945a09b14c1a0e200c279d18b93af5f2cc73240a63482b1fecc56d2e841fc8f7f
z2e61d3718d3d2bba096744ad3562531474a917a54209972f3c578d2cf03f55565cb87d7bc4fd47
z4fddfe749cfc76ef1b3330a6d562e94221f004ca4dc393dabd1eeccd521a1350a9e9c24ad700cc
zf24ff62bd3c4a59a1234fba001c9b16980613ae008cbfc34e7f233d9e562466a5994b87fa3edc0
zf6a602e62b1860e91699e2cfe2fa8d8687fc5ae7b64bd5a0615f2a82417d8cd38de858f8c21b5a
z56d6db65beb8d0a6bf99b9aba89c98b452ceff2bc31a2b60d514df998bffba5d54ae4d84d58aa1
z43868f31ddb7dc1b6281308bf10da19e60a9d2133c7980959648c13fb656bccfb910d6e9d83a4d
za029ca14ee8aad50fc67d9a53ef56d1f9c1cc690c5c1a9d7bd1763c26ab960ae88446b87476f19
z8363e77f15ae324341e22b2280afa6bc201d75a208d7abb14a4711d09c1ac4fc6b6ce13c812c01
z94f2a250c5381d4fea93b8f5122b7537899cab59cbe23876cabcb277af75ddc058d973ad41c2a7
zbf7428a4abc24d308763bd8aab9d984b945c4c23d63fda4d9f073516a75e188480c17607ddb120
z7a58d8e6c2833d85b3819040f2dd4897ef99b87c72a683c2a2b290e212a6868add8adcc576d540
z7a1ad90102f26664728031cc68d2dbd19fad063607740c7e2037f2bfa44ce01a6c3bd63db4302b
zf7a5b4c97d1169c02dfc60b38c8a31088e19fe38850d1d3d2acd710cc40d009f38d5817b11e44f
z2d449e62e183fc37cf3b5834d38b1da0d22bfac43bb0acb6b35cbf91ab45d4ba41398c201fc626
z824c22227e14c2f83fed7cf4970404f497ed0f8d33f22446896cfa57717d64bcb0f8a00d9a0c36
z226088b6933b2fc979f42b22eb6388c93b845e9688545ec490ec8de48a496f8d52c9512fcb9120
z60400f5f8fcc199f4d0b7d6e30e366e3bfe5de480a2abd3e72b0b60f71a6fa3a011c680fe78233
z2a1ac9ed6172044c053b9051a52b97219fc3aaf57285c2009f3667b8abc5c9c405968b48030de3
z43918c17b70d945f917b44d09bb23f2543b30a7d55060bbf1facc5e58d8fc35d149c3f1c1887c0
zd7317bd3f7afad2d2fd3b52b5181bac454e02e0b128f67ed611ce2261be66fe78d81db6bb9955d
z06b4a5d1d9f01d135352b90507f81a2f0bd52819814d62f1cb50d15b6ef9126dd81b49a0c90814
zfe321c79a9360c7b84adb8d5e523d4e829db8317ec82b0e44f316ee959e010f6ceffde7626d430
za1c4dc0d05feabbdf5da8356a721360e7c44355a18cad5967206d8008ff271864fdf6385129dad
zd3222adafd8f449042c976e0e38a783d474fd29469b01c3ff8a4c2a54b8c8a4153932fb88cce3d
zbb69afc362ba813761c6767db7f52cd735d5400771a5d38d1b051e713ba5881c87829d0c9f5c1b
zd29e5bf2319b359883174e65b885412ab93305f1d47216b6be206953bd71c96f47267e8c1d86bc
z5114981fa9c6342cceed44e56bdbd7b286c212b9f6963e7850a8a33b301662619d1fb626bc8f4d
z6ed89df255fcf110700563540cec5ad5e8c3818d38a0155d544390d53e7a5669aeb38c17f97db0
zdd86437bafefd32c41087b2e9e164de0cd1d1ed8a76d7edf2d63c718d81ae951bbf6df473f863b
zcf1702101307f69bf25407afebafb9f859e03726109fe9d773eae5234853faba76bc170017a1e3
z76d26be549ff63ebcc3902e0bbb4bf1c35e607c7da23cf4c7d677b47522ed03bfc6b3769903345
zf3dde397331018731d93120db86b3763232f8402b50ff73c3cb70768b851bc3fcdbfc9dbe36a73
z2eb49c40a3ed2b730c6353b36c3b1493ee62495eac61ec7bd54d2394466f380efa81507c564802
z5572912ae5db77376abda970b733b973c1d1b16034b2bae6ac78cb457eebf2740860a231b4510f
z1df7e76b7952dd668937d5b34382c35c613c818a1100e58e900ded21d364d39bc01f6cfb6bb1a5
z35ee6f4e82a0a27095346c825e10c8f4217faba3a248f9d8d0ca11d14233b452244d9305362fd4
z340331a5c3ac78eaddd1f59aafae052725e13c56fac3ce5a3e29a6ccc96d6c45a7550ebe12cbd5
ze76e47d335ecc4c5522d0619bd66b903ba1f7712bb94c49d0c873954d5a3edb7fd50978c0e81e1
z06b6b4b13695d3ac00486581572389c986f94581fdf8913291a0b526382398dfdd190b9e712773
z1e8ceafec571cb4132fc79a9d9fb2da41eeeab02b928c293a548787db7b32e406df6b1d20160b2
z2fd90859b9ca72d8d7a359c3aaaf8b3a044df079ff0b8cd76f84d127972813c943b4398cd06bfb
z9f2c7e33ae556a064393c1a805bf16d47d9993a1f3238ff67222678899a9322a5644f00e94df56
z5a3fd30ad6c0e983aab8a7bf3733fc4d640d955bf56838f5b61ba397b744e4bb2e4d6386b6b783
z3093838ba13cf3348fe91828e3c208c215c7178e15ff5c4437530f3f3963f355558f6258a56886
z37be5f39951dd374c13649911c900a005da37367ad2defeafda72ccb503e75ba5d0fa6cfe07303
z1d0b201b493a7175c9edf8bd770d88d1a76c3f76eae2f133d30fc8d0a0d73ed8cc6dae8436097b
zc0ff5de17bef043b3c2a68a5ca4ab7eaf4ea0de2825733027df6709f02f9d3ed37115c7d7be00b
z09a57a8723bd90abdc8dbbae943b58481b486d14886783a51590ee8327e232e90927e54667d89f
z0c45fa1ec09c4addbe95e3bddf0d6335d6af6c80792ce025009b2f71bdedea36595f10c93bb060
z60b080201a8bc7c62f2284173dda8f85c108abc67b243af7575f80d315ab5566241538bdbf3122
zdcc28c2560f7e72ab979b97ad62555978e539d7f026e56a7a18de4d3ccf450ec4647578ff5cbf6
ze3595a8a1354a300795f0200bc6465cb6b9a299d747599864c5c12b05e80f4e6e23403efaa327a
zfc738bbb7f895ff227bbbc8ecde045e2355f4a38bdd977a8323749b6c12bb993409e1f7976ce73
z7254285c4d17d3387b91ae8f60891396acee209362c52a8edbc56831ea6367a3880c4b4e93cf10
zf223a342d5bdafa2d37893a7d06f91336d9d722f124dccf593bdb17dd0508d0db462d2a4958388
zf6b79774cb5def445476513660014439c52cdaedeb9812a84b00b184ab1ba1cfd723dbb2b9f3f3
z48020a661214410f3c177ceab750f1e135784cffdbf6281f9e3a44b5fe34398fd61cb2b110c483
z2d63551b55275c15860ab6ebf4910fc56b791b1ae120545bc5bcbea12d2a8a27aeba0fa8608431
zaa9890fe7ce1c64208abbd232ed2c50bfbe47000547ebe978496fb1a14f11aa200e4ed17568802
z33f893b0833ee25a680fb246a6144d53adf940247bbbdf12021f6510a3948cbd2a9ce0ec0d2ba5
zf28f9a52a6a91d9b892a6286385f43aa91d9547eef738933b2a64ce96b0c42e39d7d7452e9c124
z415e6b9cb80c857a277b2f5f9a6016909018422b5d71e9b33372369d4766476586ea6ef766cded
z4eb9203b4cdc52b9befa2e7aeccf63ff5f9cf5b7d4ed8c08961f5f39b4bdfbc471dc6a919d097b
zf75a86bff07b9c95e3d74e8149b611459a99f27e1b5a7ff90009b34a27a839fb1007ff5af15533
z205dbe5e7cca47b0e4aa10d65e1ac713375dd863d6fccc2304b4c2891e33d0ab3c6cf912182d3d
z0eb04e464af01230684b2ee82b0e0894a5304a7ac0277d86fa0a0dad38052b7468dcefde400c07
z8783fadb16ff92adb0bb0138c33863707fec53b88dc1f14a5564c9e995109e024b98fc63c8e3fe
zd611262c77927241657acf2da2a2a22d167badd542c08085e04d0da2915389f5390f6faf36f1a5
zf5532b0c716d69e94b5ed3eb2e345c3d15708fdbd2c437d56e4478769d0fefee038d3d4ee2ed17
zfdb905f558745b371bd02b471b5372626c6ae785c02d05160599560f294619e07e94fcdc93e528
z1faa667476bbc7852b17f052f2871c89b0ee5adfa21bddcfd605111b52e5d05adc3abb82f61ebc
z8dfb231fbcafce24608ebb10cb71d1b39f25e396a3b12923f37b416f44db3eb968736e238fb7fd
ze367860412ef5a621da9eb98e4bc85707e87af27bf9cfb5f15c42c2b1459737ab98f7a4f9c9acc
z33a59d8a578ec0cf80c3d38be5df62a9b18cd3362db0c5015f5db6bc85fa7db83c966e2cedd4af
z96ecfe6a826fe8a4810cb2bf97648b5cdb7067a208cff34155a23da9799acb78470f519a5278bf
zbf2ac3f44084f38e1f51682c62fbb8095d77e68afa72e83f72081584188216c98e79141ee814d1
zcf523147438f0ce7b8fe762532e1806bd92202b8d2f44a0b1bc81e4efdde835b9de648e1a0132b
z7355f82c915ccc966f94b5d1cfcd945947719ee5e43607ad469c805cf223ba622844b311b8a0b6
z50e9439b67d8128271c209141e825bc58a1acff16d2c953334858fba60bcc54cbf26395f0f68d0
z4dbbb35609236f235df87f7d7020649d27df506946bcf70ff228115008af80ea4f3d3dd74cfc91
z3927db378df6526d80dd22b6b78d489f68389695eead6baf0261bdc7d8fc8c466545dac06b273e
zb88a149d095883d4d24a1fb60be0a829fd4e17defdbe63ecdfc8c45d106e43e3e9c06be3b0a3db
z856d7fb1387f26cd4d25202fdd3574463d05782122a32d45c7c7851a572a60712188d4939403d3
zc538b458ef6bad51ea77ecb296f2a5ed6bd5b6929f297bddc48f33f36de63bd193863ae6c62f66
z28970780ac4d37e499e83027f0501a382c799cfcb1f13f761ee588bdd10dc3e35faccb15a53e34
zb6df10baa11ac8c4275e54cd6f9b979caabbc082007eea93a19c9fcefc10160c79879fc9995e29
zcab058166ed1f9b81d989f5e0058ccb4c32faac7b13231b87d2d5d1013633623048bdb3d851ceb
z065ca58b8b0416ee85ff2b16b870f80e2f30098dd095efaaa14cb8ce99fca8df6b130187199c51
za4e6cb3829b016bbf22db881bebcf595a438e17547b2f7676e1f62deb515f2859a4b5795006647
z3156578e978efc37cc73ac42f1a1d145e0b307787500c20feca16f4df4cc92154b262ba6b442cb
zb63d3e1c19825d89f6d2a87978e1d02fd88785d5b20c6fb29a2e8178e5c843ccbdb9e7f3a2104c
z84de959d6fcce9137cce0ece191ee7eccbeca8300c90993f2c3cd61d844940973b62f279869fa6
zfefb377043ff6e1b5b157b230ec426e5152e8d084c51f413c30c385eb1e7b6c27980275ba54120
zb693bef91cefd6e5476b7222dc21258808eef29ff628eff922cacda0de9fda3299fea5420a4b58
zd26a7f8aefff7b72cfae3430e78b11118f55bd306a6c5d4c03c4929ebcccd3df0d2473ff76e761
za7038dce0290f17d433cfcda72d3b9625a83dac32ee92fa648533db3e7bff2b4e3e4413afb43e3
z0f6c43b71b16c0c73e1d9b47dfbc1e6bf1f4b6df13d5c95b3068b539a93c7ec7ccf7cd563e71f7
z64b7aabf674ec8d08c3ebe1ee7529ab773c8dd8793e0caeb3c751f7fff554a44bddf9d84d15910
z80052c0a91d6c4508be51bf4f41203dcf0d58743434299845f08f1fde407facdc4289a9049c567
z7eea7a4dd947929e4632bbaac7c9a960942017f2b4b5152d1138b5c2d02244f17210d79b979a3d
z4592b5aefef749e7f014885edfc52ac5b73cd5f98d56d29484a822c4aa44ded71e78b13d728cf9
z305dd9c88c684e99ae141f93dac5e83d2373c5cf38863619653772ee25aadf453e5d28f7a63579
zb9b576bb41a6860f14be7fdb1fc48b10daa2f8f4c5d862d9c702fec1b4f76e065494e42475317c
zc53590f1328bb45cd7d745debd9190ad566241be93d0ea924aa858d5175ddfdad3b29dc30ed59a
zdf4d2efaf045eaed819673765250bc6d53a84e11501d4a7845aea926479d429084b9cfbfbde8f1
zd0e8a1fb490b163fd947fc3e9ae6b8966f02daa77a71fdc9d63d215927b9180c419f9957197153
zc63d56da7fbfea914095c2c641caf1101985687b170b29f611098beb16f889396eb46541747682
z30c8991df38f4b1ffa8bc6ffbcd85047668fac54a73297d9c6b0201743b285a56e84030690e759
z7f308e0996d1f0d08480db6c264ecad347be2f0829ca2a1021ad9aa9ae6f69cf9b4e94e6183766
z1450c8ee8880aec2497cd2af129b15a9f37a74e4b46b4342b84f193e3a66bfaf076882403e3bf4
z0f3dc8de3aad61097c00da30a154d2ad8c07e48bc0b6517959e72d75acaf673a5c4b0202f9e6bf
zd31b96e57da198936a7b468a6ecabfa15e41206e032854c6e811fd1c307c00f9dd2c43ad61e2a5
z73ba21400a1ae9f149e8d8cf1958056f3b792f437e666b1f21bf4f58c7a9bb25b3dc20b8bcba7f
z38dec4621603fcdd23fba64806b8f162834e3887fe3b39be69b59c761d32fe989ed72be2c58d6b
z06b4ac3e6b99d5f607899701991d82850c53b40f7acd9d64683092f08460e6253b937af20e08c3
z83bf46f2986805c72ad143f5fea48501c688b63af0e194d7410562b27fa74252a6bc79ba235c0e
zb8fa4c7eb85d0d6914e4a30a7d9293f4cb6cabf0797b8453e8bebc38e3ca4e1574765414b6cbe3
z3473bb08ea031207af5cb9bd8c244140d5affedf2528310cb67230a589f9b387eb91bcc79b2d7b
za3d7a56fa9e4fc24d661664aeba4a9034f020deda5622d7b24d75ce45495529558313c44e07aac
z8c16979a358b829ba6394523de03a540b4155d63809354f88350bd8297a406d9f79949a398b8b6
zf2f4f718a9b64831ccc0d50d98aacf3a8f4d80b1f0eb3e88bc5e6f7ef16b296120deaf94a841e4
zb4e1326668db6878207a4fb1c6a716fe206e1fb2e4dbd0cfb9d591e6491b01e19f826f5cac6e42
zd48d413a69cdf1dd2d50a090874da72433f6aa38f1cd29c7eaa60d9b9e34f055640879c744644c
z78c67077114872dab0f5fdc249e778f5f8fce7e3ca5baf045ac8b5612c5d42f287bb9230bff737
z84773d5008f1867f43455fac2047f9d5dd95caec64a7e99e1c4f30eb295cde451fc0ea785553e7
zd8b06ece45b65863c15524bce7059e1ec6b9981f9a6629dbdba0fdc90f1e5d78560fcb7620aa0f
z9a99b4436be8398230af511ce2bcd791aee07661a43b70208265d8f0569f971a752b1c75c04e88
z51364dd7ada3cb0cc5824b8d38da21b074cd33a0c773cd1a64445a3b94056f1440d766891a6963
z899cd8147cb6d9cb95bc5472c2eaf43e53edad9b12c55dd23b6852f882c23a42480cf91dd82b43
z3151565d01a92ac2e7de95a69a6e1fca1b4842a7804d1ce7b13f5855e7c837fe4f9f4c9277dfa9
z3b4a08cbc671b5ac45861aaf76906abd1bb1fa890a204d200cff4cd04865d7c8549bc1ca3016af
ze1a16f6c0030cb543fbda08d0bae9010d0ff6710fab83ac63084b0de51201098fc0972f8b1944c
zac2b9397140aa6f2d1d07ca213bb1a590164eea7fb89e268bfc18efd578a2db3a82ecadb175f0c
zd24bc25b454b77229145d8e3b9bf19a1e946471e6cedc89d1b33120da38e0404ad0cf2fb32d296
zffe61554b35ef3c6b29abcebdbbf8964880dafd073dfc3797d50da91290ef4c886b14104f87eb9
zb1e05a0bb47de989d822649adcce9a3f1b4b337d44f1df83d81d4e154c94fa0ad81095ffa2a749
zf160f6f53581cf6d1b05514036c7784501b896308e2f05edaa317dcd597822ad7dfb197f05728f
zef638a7ce5dea5bd6d92691b569bca7be196e6b00cef7d07bba025a4197c88ce1c0ddf6033a2ee
z2a085a7c3e0ff458bc67421ea034d12b222a15a3fc8748536e6a3e36ddfb30b13fb2979a0a7a28
zd65ae16d54d2ab4983dfaa1f41ea57eed123258f471a21a249e490793c618faa02090be7445626
z918f87a28053bf0d1425daacb9da02316cd0bfae4aa7cf27c2b88b92660e81e3fde32f5a3b1314
zd4b9a0b330de8e03fb5f3dd1bbf7931dcd4425feed92bcb763f6e425bbeab75bae0b2a97396b2f
z73126e7c34764f44c66d77b02f2de779f19c7a667e60339a2e71155384762abcfdf32e92dce4b8
zc2604bb680dee37869c8b2393027c53f88e27ad6bf2879d0467af4e78dcac0b0928531e45d219c
zac582f600715cbb1ee2b1829d79dfd8daa5d0a69838cb121f6af4eb93aeabe1094173e6a4508db
z0a5fc07b949c2312b800f7ee8a0cff0e9072bf4cb2edf8f244f0ae3902ccc9f57bcb1089ce2d9f
z37e8bdb7b154d442073bcba49300b333f3daf8bfff79f7b36b3e795f855bbebccc88be4db7084d
za61863249d729a264eca21b1eb7d73da59b8fe1a6aa132e95f6f9f03a2a58ad406a696970753d4
zaaa691edf20827c8bf9ca45ece586788f14ba4c1765104aa6a29bde8c1744a9e77d24199de1ecf
za9aa5123b14d141f93cc0ea05f15374e0a9866962b9558e45ce7def111e5c1e7e2fd4c6ae932ea
z24b647b14b9a6241652da9d6e7b4fa3832c10d463809ef09b0d9cde2d18def3a5e2d2375bb3513
z1454c36ed7e04bfdcec241ab1b9a2ab9e0f5d3d95f0d91052c8061a85ff95cf4d8f6d11116e9ae
z76d67ed247303da7f2ff548386043b9688c59aeb7ca63a2ef0122221cacaf1484ab2a4d2cbacb6
zf89862c8b9673f11230cceac51654f332e537d700d78ea5023338f111b952604694204339ef6a5
z60fb021878653a835b0f65032c790bd1d55c354cab83a0034ab1c66509511686fdb8758d234abc
zfe6a6c3ba3a40a73de86d9f642a222e46fab214e6de86455cf579347c4b8d89b0a6ef91da3bdef
z4efd862e005c7240e33c1a6fc0c77834b67c767ca8f14c5eab02827588630fae63c0242584ead2
z44029c1c78cde9abf83378aa38bc83075b380c77315251fec3db03f57a8e896064a10501e700d0
zc9e253253288c6d060a206ca82930a78984dc7b4d04d3265dff35eeb083dd62f3dbd82011886c8
zf1cf6eb03595af45130ce8413a2c3fececc4f8e9774bd7ed27af35e7da7472033335151387bd16
z73e6bc623c336f3bb284ffd8a49c5ab9e0ccf7e51663fa1583d98dd573633edbf05fb1cf7e907c
zf2747a882525299ad40309976c8aac45f698541ada0dead48ccca11841b6d830fcdbefe8a91ead
z082160d904349b3e7ce4376e6ba895a00c607bd41fc0d80a93c7ab4f0da974be85900d1e9cc17d
ze794e96b1a6a0a6498c3c3f9e85a21abeec3e66642b80f99eb8f0fcb57ea40fe64543cb55bbd8c
z303d065764d29e99b948dc2d059ccda3edc25162c4ccf2f9796163c00e555439278bc240e62c06
zd5ed3753d0c94500c9b694b71f86b87b9e4ae83c96e3c46cb9f3592e02e2a8d2099487c34b05ab
z23fe43edebb899769af0781e8cabba343ea16cf07ebb1bee8436f841ff21303d279b020e5ce9e4
z14862493478cc8394bbed36bbd5df1e54ee8b88768c86cdcde6e97c0a6fdbfa5e8da6a4aff717b
zfdcc01f2dcd2b128ddcf2bc40a6abaa9481236568af2af095836ac9fdcc8049f15e0137352a129
zfd30ed6249bf59d534bb871ada1e9b92fb5e7ca13229bff15f0ed3a185690aac2531f3c92aba9d
z5726b611cf82fb382afaaa987bd7459dad1b50d9fff60c6c3f0f2bbd8e9b55161810f608b44ac4
z2627646725985403ed654b3cb72b333c7995b1decbac4e1134487cb475a434c8029689a6b73a67
za2cdf2716c9034adffbb515d1b342c3abe7e4ead9aa792156c785d6e854baacf122cdce49e3a41
zbc4fa9cbf08ee34953b1b04ba89da5f21408db24eca0b5b89c560c21e919343f8afdaff2285382
z37a818c4eb1806bea533902af432480a34d59664a2daf8d743f832d53c1c6e10db5ab6f1a29e90
z2826e1aba8827dd45499542052816d52be56d1340f76d8dc16f814c4bec3f598e72a0996bfa6a2
z09eaaf496106fbdc25ccebe1747286c7dfbf566e5783c585ed3b0ea4ffe0ee83939290458b88dd
z15b78a79b169ca2c910ce9b7bd0611152584527a4d322bf4fa21a0fa00225b09e36d8b5d584ec5
zc8ef8b8fa83c9dc805fcc271a266410e351bc7021d4b7cb2b0fcd1f1098de89cd13463cb7643c9
z2deef30240c818696dfbfb25e5e45c98410a5482d8883b1105c6d66fd6370f725dc736ed70e1d4
z6fefbd270214bcdca6a124858c1d9c065423b791d5dd1612b11294e1ee4b9e49581fb2ae4f4636
ze366c8ac0e878a1c8c6434f7e2975a98909b26abde04a7ec9e44554afd01e65112597a0fd95994
z8eab69027bf134612f2c5592d3451aeb16575f06e03b86f6705b913b0f5091f13eb32ee984c077
z34e22076c19f5ee46ef34e463346c1322c6e6ea2e9b4a5462f457003778e13ac07b57c00ac4dfd
zf1dae3892cf825d8f3627ac80eed162a498fb2b4cdf40e769f5906d7214092815a790237375391
z810cdb897b12f0d9a4aed45d444378e221097dae69bccc47833f552e89a1ba86ba6e1315c60e90
zb97664b7979d3028a4df1fa016d143891395a4511fed5bd0b0d16bf0b5b56fe88eac52869da485
zfb46c1a54e41e35639ed291a05ff6379fadfb9c7bf2cda3f1d4d11ddaf4cba0f96d776661d41bd
z5854f8b33efb73989f20161378d0581aff2bded1058626fe50aaceee42740bc4ce072e12519272
zb8c76308
`end_protected_0in
`else
`ifdef MODEL_TECH
`include "qvl_assert_follower_assertions.mti.svp"
`endif // MODEL_TECH
`endif // encrypted_0in
