`ifdef encrypted_0in
`protected_0in
ze74c34e226135848fe16db9ffd31815111b6d7fb642c521a3f628cf6da949865580b22efd062a7
ze90adae0e65e66a2c36a587d0a790699161455169ed55a01f2084f11770a774ec4c588039b380f
z6de9c5084882a40b79a175f5c2114b2b6d78b070cb806e1c0aa9258297f4687ab308bc470f0040
zb0b1de382961eeeaf2e279e1462520fc31c119af8f2b214846f56c2b3cd2eadbe4099496abff18
z15cec83ec4a77b868344aa20ba7360908f5c0de2a79abf8b3534b883bb12180f68b5d4beb444cf
z3fba8f13afb0abfe8fcc4294810f75afe452434d2d0f1166236c82f76edf1e12979f04bc35693e
z32ae028996dd85737a8f5adc1ebb94f39c940246e887647b64782cd7ab429b0544c173176cede7
z01dfb26b1f73408344a52b7e1f117f12bb9c8077b34876c2e6fdc085981637012dc9754765e1a9
zc512ce062e0b8fb16a214591f5c81e1353b900a611fe1f4886b57940b41b7f2ce99a7b84b04b90
z916f717e73bd10589c81e207ed77ec660a8cbed5b487fa50acde1b055c8870bd8676023f21ddcf
z9c98cc47cfa2d654ff1365d1f45035a045a66c5dfa82790502623b57a3af03bf0f0c0d35b51558
zb8b5f2d29acf03737a9ca2a053b7a8f06800d50b465c41b30eb585f62f3d0c2c5a43bc34362c5a
z3d9608385c2cbacd43304ea39a46e6842c8b74b88b67156934f45ddb292f1ee039f2ff7a9cfc0d
z77b96ed0ac12387c4e43b77e8a0278354e7a44c4c7e932861ff899137d875679c86ef4ede12628
z15152fbf2a4c1d4d7d20b6e7da6bab21f71e4f9e84daed7f565d0b628dda769ae6285062e2a074
z03242216b4a69691418638e818e19bfe1dcdda02ade8a09fc9419cc1273e6336ebc2f67a388931
z8ee5938102a059bc1c59720ad454a7b6cd53e056bda4e2144029d73127ace5899cca54864aec4c
z0c8e0188fd13ab7e2598d3741d8013e8b6dea6a56fc5db254dac430b7fd7d3019132366aed6aed
ze2cbc46a76e5f898d056d2f540b074815f6c27ac94f4ed3e019c54e7acd7fb9297361d303531a9
zd81c574d9def5582de0d599235439e651821f737a14a8abf464b55bf3582ecc00204e0c1ecc8cc
z6890dccce9cb76ad20188f8cc3f47301ec21903b09269bb229b82c30c783ea976701cb8c0cff52
zdbb2636209478d71eef84626fe986a746372978a8857d5508abc1f10b02a5ade00e3bccfef60d8
zef5ffd5508078d39c7f336020b513882bc732d662a1851f27c5e94694c09872089543932387077
z0ae8d6db5a98f74f37a574bed943f2fad0f97d84d00eb53b0b241a27699f274e8a4f2cdccc8058
z291cd48d8876f6936679cd4ccce98798a1fe3e3f036d18ef2d92fe41cc63517a90c1fd17593335
zdf7ecb4daab3a77fe02519d88623111787dc659a9007ad9de2b6bf555432dec1e7982c8b455338
zb84f26ea5bc1258d256c9591ccadae18b42283bba0cdc48baa509d38dff0f16aa9cfb3a5aa1161
z4781fd6a48af63cd1f6a8d1d3c6354da9a524ff76d69739b050faa62eca38ca223264c2b496c0b
ze38444883e2f7fcff61f57fc70942717835c332064a46a481222210db1d36e41376f16d44ff26a
z9c16a78d608327607f4901c986016b1fe582895303aac165799809df3318868e0c9b120eba29a6
z8be754ff9a9dae0c101947ee36e0c8ba27d1ef050a788b029476ffa327a2638393a9e4da3be33e
ze863ebed68df07f8fdbf8487fb297b70f6ad6fb6aff9d43e35d9adc64d88feed36dca54b128fd6
z41a3feedf03033c20e135bae2f621095e87ddfb0864e2b56de425bada9aea9a4d3357950a360ae
z0ea46ede3977c7b63b36967551ff61a3f314d25205ef60042555310b3bb940258c63301112e92a
zf75a9e08eddd6572289ee3503298f762c4e5ea75e920ec6bdbbf49d76ab02a63ed858e5d131c89
zdf0bbfff4fe35d36bec8325106b98d8297bfc233085bb1a3c192537d538518682a9f34311837dd
z9640d217f1dc13b3f53298270f11aa1c00214c146501f07c0212d95282c815c74ace872c5cfd44
z66e8ca77139d9bbab46217266d096a6c6c68247d72492476d63f16e2467e703ebccf69c352de3c
z1fcd144da0c45a4b645c27cd6ebbb7b8349fefee07714c7f4b6b7c36ee1f68cd883ed49ad80985
zf55ffa506ee1dac8ca6842376e7eb02459e8674cc004849d14679474083c855d0163987959b1e5
z048aff5e6f346b5704e2fa30f633c90d4cd51d05f3b94ad5447662ad94ac406a5b01ea71a260d7
z0287014154b15f2e7a09807111a5a49d788e7d4919d5543f14ee1519fdd197242512da7c1abdb3
z02abd3bcb6f123eb326c56d49a08b94b74e389e77f26c6e3280f1790f125e9a4139750c62200a8
zb252cfd040aabafe1452d6c3763b8d1b2682d24a57fac5cb0f3bb4140d78f00f3883afcc25802d
z288e1a5a4df63929578b854b4efe684d64ed19dd739ad538f489a59c120b5427d914b3115be3bf
z1600d8e42d0608f407c2f98cdc3503189f5b1e1c6db2739f6fbb777b176c7e8ab12d6d79622df8
z08b70bd5fd46bfa364c6ad63d121215b705c0be2603572f6b0c23c54bf950fd0f7f8cbf8b788d0
z55e1969f770101464672f731b7aea28311fb027daa4f11a681d6ef4abe821b3840f78c318c7a3a
zd238fac14ba9c4209ee1693808a3db8fa26ac3857112f1ec354f51cb542d4f90b60e0d75110409
z461038be390a5bc401e21ece4f041f0bae97e99dfffe76debc0f7904174794251cdb4abea9ce12
z821388c2852f952619553147c46978db631f3f09e7a5d5ea4a6848721472a5530ea54fc7cbc81c
ze7a54b2bde313279fa41e44cd668f44a065dc18e59493e14df8dc45b7c2378128084441d590407
z2f495422f5577e140f06607f140ec53bda6ec911a323a8eda581cb5947f52f6d4d8fc2b97b3256
z3bcf5dbb4b83139dd5faef9a82eb2055088b91d396c5d99dc701b6d3623d1200dfd89269587b52
zc11dce8566c4db1499e9415f2e74d71238e8bcb20e8311727906fa4fe6c5bedd271639c24c2250
zb67853c6cb50addebe47defe8f8ad616e10c01cd883fbc804a1817c0fb06a49a808cc0b145bd69
z7dcc751e379e32c5e2e5c964fe472afb41136f08dcc29d515634ec7cc642343df9cd12518f0136
z3add75e741b0105fcaf360ed5493e4e251fbfb67960dc41b9ed434e7918dcc9d8e943b28635ee5
zd608a9fcc2e94f3a2074971bddfe21e1cc1a50082852f63867ff036bb06b435b955a2f6f1de382
z3bb0a32e76068193535dd955be470447512ba16c867e1b546d27c330520855402f9e87fe57c70a
z5faf075f06a28e05bdaebf8c4068109416e73d37b3e2a70c470430252bd83a05a5272e74b684af
z0edb00664c275780c5abf3a00a04cfca1838325b8beadf62cd6f4e6d40da56c42b580b5b3d2902
zb2feb925795fee0b2e5eb4a14b596700aa28379f061a2f218cd9cde5430dd9eec947fb38524b5a
z032c5a63d42aa71f9be54e723987a299a0d2e358c6086062a7f10633950fc3d1c4f92217dd6628
z94d9f76a06b08086b2d6987af96b92f84e02bc32e299e3ef1f04b5d18fb456ac988ead141eec30
ze6f5aff4e1d945289ba364331da14452e7bf8ba6d39c124e11a81c48326bdb52157c6fc1d41d9a
z367850c1341df486ea880d55c33b58464d4ce4cd68a212a894a29db8689335fa40a66761419b81
zb003ad5fc99d635f27fcdbce3f1f2fe062668056ad9b7e5da47f980790a523668536d2624ce4d2
z12f80dfe807657f239b521d1aa1d38adad47cf1483da72f643d4ae98c9f23d4d8480d5f0ee5929
zd171e28d108c4a9c0420b3caa1fb226b90d44135f147485b82354f70bd6a799c79f1f6e9a7ccfe
z2e3a6d34c4845459f3f94d6c242fb71500f0447cbf052f31d23b1168318dd0e967567f3af235f3
zff9f9ad019dc1fe20e00081aa20e847316e414def9d18dbd1f14c1a8f1b57f777718e6bf82dc22
z13a3e5419c1e76985e446b654f81982f934a850cfc384e3a4244b6247318fc4f06c19f94089621
zcee7b10c02525b053e6cbc1b5c4683dd07fc379b2261ade6d90a227e9ba7952652b099a6f2c283
z50eed812aa71e59bb979e087c55652edf5bd5b7a7f26cae43eea433d03c5daaa128e8321164ef4
za2e4457d97492bee286a230c1e281efaa0c543beff0cb02c8e16e01e834b0d43d77137edf6cf51
zaae5e7438a995eda2a5ec8361aa4f306ca0d3595f637c7752c2c018b300cce3c66137e84bf9084
zf835de1bf8901dad60a63a389c2c219c1e14a807d22e6351ba2071d85f0e03ca3018cabc06edfc
z004ea058d5dafd88c8269cc0d726249ca285e7bdc3d52c3266bfa0ae871393fbd4d44723121a18
z6076e9115ba8f48eab2dd9af92af3958514adedf5574d1c69029de13e2dd41354e20651e3b2e07
z1f4176f8cde77e1e6f8dfe2b87e2fb5c48f73f849de0f5349218e3d7b4cb7ccb4f5da927c060d2
z8083a1cf3bb009595c2c3bd02dba63d25231f75ca6694d43c738fbcf5c4e8ba75a5216b0702de4
z35e8bd7c43c1e0153d71672264e3f534bbc62e4db009c50b719fc9ecb1bc1968db6a574da2764d
zf673eb914e5da34806b819ae34c56c023c065ffe889671eb51bb254f4b657501476f24a2290c31
zf35cd0330ba60c5df167a5dc25b96630a70f27dc8698e5eae9de87a5a9820e1460b1fb7f29c62a
z47e525e54cba5bbc99dcc5b447d3ba5b9580aceacc44eaee7873cb5e45b68d3aca1418291d388b
zed0fba6e56e8239baed6fde759354a52d6a75b8d0c0836d716993ad4bbd1e68dc3de17215b98c0
z2e5092409e0ded694d75d33f51f8ea0dd0aa9d3218ba3c9131c98143e49e9600346be74ef406e3
z42ce947fa6718f478a76a17ff8749d966de2eff8c33eee9a704a910c41a86db63a9ec2e02bd46d
z5a3d701392434624f8541eb27d0f05a01b38fb27226452d680fa608a278b0acca1b7935c3d1fa5
za993fea34d2a15d1b7d2199afe288df5efa703c5222910d0c9cf04138869f69ea8a8cba6323809
z65d4d49f04091a60cea045a830c2c442819d0df147ac6723a17aac127c9855f5af5ce015f14830
z9debfb636502b3928c2b6229f7ff207663e724ac622cee5647e271b2571c94e036c8664be01d6d
ze17b27a5939937aa7690a1833f3690a6a9e16c8e4650a1b6d279a702d7dc4b31ed7ae2069cc254
z190767026a2d50f76bee42929941ccd34e48937139f6c90cde0a46087278d4bcb432b224c60f5e
zb2c370de4bb4cc08c99b5c02ba32bfbf96f6c7e6a8a6ad8a00010d94f3e7005eee66389ecadddd
zdc52a40e1ca23a2c8906b44f2fc1615b12e56c19468619c3823a72b70499949638b7ada5347676
zfd0529c23ea891b4762be5e7a7cb683eb86d55a6df0cdf65e48cc235a61bfbe427f5a0ff963db5
z14d9b1b9b78b068f734c0ad7460c159eb272f2be87afc607339215a2e4a0a02bdbef481fce6404
z63fa0dfc26be0921a0b8d394b337fa83a4c664cb0c1d3c02997f99bb06950e4b43e88afa9a5ea8
z292a1954c0ad0939269b61f23de3f5f7d669c9d268a4ee837d5921e37c8f91e456f2a0b752a9ed
zffb5d48e24414c7176d0ccc4ff6c64662b37436cd0b21c71fdbddac5800a7bc2604755891d66d1
zea4a1cc9bc8e09d84b1878dd193d15fe13a58a4feb2b73df0be51954aef2994769c83d99c5984a
zd09b032a7dc69a1bcf83c14228d276ec2d44dc9c84e36964b7238449694f7cec2c274274ec40c7
z34a1d027b2b322045e9df2eaeef101d374877c7680d8bc315a75e41da186b4abdf379dfb961ba9
zf049d19ddafed6bce84f5adf7834df5dd936d2457097114967bfba9ef9f8a7428dbc0d66557fb4
z15d6dd598fe2917040532ac641e4856b12129463ad6c85a5c30b231dc18a8f302b51627d001f25
z4dd4461bca232b079b958b4e3c6d802caef1e004c70d1e90fc226bc68e6f4f1c60c1cc2de7bd36
zaf9136ceb2dcacc8683e05b7f636c10d76d840ea8658c4ccaa5a41486f8dc87764051515d58baa
zc3ed735efb33a2fe4bc99672a7ab5d00bf61c2c28f7b288acc6cbc7f1d77b16a237d699a2ba7c5
zee9f04187725364f6628ee36ef49defa480bad7e6c761514a34f079945737be2a8366c7f52d6c4
z1ee22856592c2d04f995038348ea75a6f656f57c47512dddbca4c83d9bc9b35c54a4594c386889
ze5bb2b917cf9d757dc6c6a43e11a83d4f642818ecefe8fcd9de84c18ecfd5392d9e30922e23f33
z257bc004e22d3ce27c87e45703c5e21787386da9bc72454f0172e704bc5ce26124d5f7189b853a
zcdff72ae2fe88351f0da2f055a816b34e4ac9f616aebb3954d8ba0ccdbdc83b15bae7fe6f5c2be
zed09cf45d3ea697af421d1fec1b1971b3994270d5ecba081102ecdccf3a36a807accb56886593d
zc180eb09f8d1fc6bd5c295f9dbecec6058c35f3e043e7976d68b261fc83f7212a9d3433460520d
z740b5036dcfeb727c2641f6a73548a0bb6e566a5d93a00b521dc910fdd939756bf1576d642667a
z75b5ebfe5e0feedf46fe78a7c3b2b34fd3486ce3a7c1cd130c1aeb1e6af9851be180efac7225da
z5be19cbe20cca47a11eaf1ccde6c4589d15803df7d2d817b8b21d7ddab1ad16435a45ae967228d
za91aeb0e0f588ce8398a2c8f9bffaa446d546b0d5b6ba45c838b8149e4b8b3da5d4403fa8eb939
zeb5713565b398f9eb9b0880628c19ab4e79373e77ca0d2ee13cd1dbdc62536eee30cdbcfa5c57c
zf2728346f9492f7ad95e838e666f63f645a17aa1fc9331e370e1d065e0d7a70e618152425707bb
z95d4bb2d560ea0ac51f97994e4c1b2504cf0219088d11285acf0990651903e9d7755227aeac4a5
z849fe60bba4a7b6de752e06aa3239f511b4ce1b8789f28c909c8918a858376b50b2b1cc1cbe2e4
z2ab059f55a30f41578006508dda6e42730583c2bab328553418e409fdca9c16acc9d84811722f5
zb6b2ef69a25379141ea6fd2a5755c20151ff2e190575d3c55bc2fd4cb38144e2a8e316b79caf7c
z138afe55913cc882dd6dfc100681bfaf1dcd0ec26e100d2278cad3c7f1749fed34ea17762cc199
z965ed041f6d86a11a093edc1c2fdfb36f8604543164f087ec234013887dc07571bd91dd73a4101
zac69ab378a6c6a82ae81a436527724107696e0b19851e557f89cd7a436357a88ff6001a990ff4f
z1142143bf499ecfc3c14df6e5f86bb6bbcc6586a0fdb117515e60ecc4a2d820fcb33d2a0b53b9f
z9fdfe1d60cc8140ec165762743595310c9d20151a62a0b6106b0668bfe0a4d9c2101bc51bf1006
z24888acd6ae1d9263b59c7dff4d618c0bed22d9582299c59097577b846cc60752c13a7685b8761
z8f79dcc652edc17fb053fdbf14ed5edc55501801be9a339b89e13d3da1af24c63ac47715117811
zb24fbf214a26deee30edc76cd7c689ff3b24e9f077ff4d896207fc100ca7f8c04342071cafc8ce
z20566f31a391cce6f6b5b814cff0c219599217e7f43b5e06cacd3ef9dc64b4408ef711cbb28024
z88d80e8ebec04ec33390d60f48b4f7bc946fa7960febe6ff9544ecc8dadaafd2e16bd34ddd1fcc
zd5d34c01d4fb3e9963328c0be78a277898b972424e2577524a5e3fb7adf276138b66547acbcdb9
z8c3284a6b6cd248a81f7d8686b38cd55c4978e8e4af8e7fb3b6fa98868d8ac8b270772d3b8f521
z09215b043569733ef1908617d10cec76ea6b5fac7e7d93571984e62befe462282fe35ff88e137b
zc68ef6d6b3f4230c1bdb3592170571abea13ad42331f0c409455e6859da897d5fbb90c6ed9a0eb
zcd43a0c5eeb7c4fe7db935fe49f944dbd53ed307a9f182450446c72c14861050714674e7de3dea
z8dff1c95625b18596bcdcb3e4ae8215db5bf654ff25205097a34de990e6a8d5c184d4997dddcf5
zb8a06ab3631ad45b886fe79faec021e454a310f2083fa1ae0721c7f852024559d832b795ca0e1c
z71b6285613207e4b3e7ce272b71860a1f8effaa5e287c809d1da11bc26d89339e8bed799cad7d6
zfdffe235272b236ba788601478079c9227e9ed5f90538cf67b8fa8190d83fcce80b9db503c7160
zc48c380bd6ff5b9f18b6d2f2d3064c6407fc906bffff65631d46ab19a1c5e4e27d0bee05f39c40
z85726a7325280fb47dd97d52b42c36c9880559f7ded5c20385a474ee16988737d7ac8110a0d81e
z25ab87d49a404dc7dae87d1a14cb4f8580551445d4f1993bc8c5bdba0cdfb537866a672f5aa279
zdc764b630091daf3d14c6a968219f9a5014690e9e324717145c367f7d19b232ae1023825a57965
z85582477c2f2ed8e03745e7808d496d7345d9c403d08983fc176b657a7e3f738f502a8632fface
z9c54568279b4465c3e91f0d231bdb5e44a75e50a1979d2dcbdf3e3533df73f00f8cd696787f7c8
za54c8756315ffc5d619a12a68328e7b0e805797de1be6ec1112709cc4c2c447c101ce803c08772
z3d3920a870eeca79c11284b4aa804cfdb4f53778376fe3aca399d316777be39e7a3918d3ae89b3
z78c4a19ba446ee07dd2dae1b2e908a145b16b7e4f59bd5169dc75965bfd6ab63733450828e7eb9
z4a26ce41875a4b01528182d61caed3aa3239c6c12b02554d5c39b985ad317d0c2c81208a63e7ad
za4f4c3147b0d15015e1780e770fddb6b8b1cfdd5b4e545912aa128a8b1104539fe18049af5bb05
z22c42e178381e957b9f7897696196b73dd741348841564e5d769e636a72bb08dc5c37d0bbcb8f4
zf861776d61a04e82499214116f4223d108fc27193fbe90857cc05c9c603d2579f35a90b09d9a71
z93a3330fc70c49805cf59ef728dabe6af36ca06452f928dc508192867f5c1c8f9f2f84318cb3b5
z38ea8c52462d8f99a3c63598f21ae2f98a5e47fb27921de10c9355f26ce6c394f643554e140ca1
z74459b2bea6b2305173f8c7502b6b3156892d689c8276bd16c7a0cdaa69f2ff9ef0ea4c74f4e41
z817b3b63899d27f2a7db9354ae559ca08f4c1511bc2c44a8110039ef89ba73597425e0c422f542
z59de2fefd2ce230db954d2ca80dbf1e76d3f9437fd9350c77db41c5cc02c860e83fffcabec01fa
zc7c46fa2b0fa5ddbf8f2616ba9c64b0fc00be57043d579c657c99cc0c5ab41d94f246f6aa240e4
z4848bc3944c9131d4500b1361640354d90b47cdeaa84c0d1230fd8c500788588bed40d8bb21158
z4a13c42589cbd7822cae0e2a36338ef6fb856352815ecedf6571f7aeba969abee0d2da4917d672
z078f644e46b7f96c837b3f27deca23f8a791c848b3b23d15c4a810027ff7b1ef3e6f1caf652f09
z860e5117bb4da424eb8a6a859a8a5122a1fae7e01f3855065407cb64f73ccd95763cb4961e456d
z697650be115a0c1b084747a94f839e29812b24a6b89e0bafa55e33f23a7fa30c0759f919e16c1a
z82a50d04a9df243bb098d922aac991a2fd84adc61116322116dbdbc659c6c76eb6c87d49e3feb6
zb5e74d33201b751f7db9bbe17a4c19467e68a17114ae98b4ff1c127f3cd2ec9ea59f77d2e8cf78
zcb839e8995d7951495bd35bf3ec26f5c52ca48ca86148467f92358d2d1e147aadcc93abd30706a
zd8186db3492e86f18bebd4860fd642de5b7454a81cab3f69e5f331969bc8bf7cbd80203a222183
z693709c53f1c8e1996b8e504b6cbc238a718a4138ebc90591f85e70dc3a8d22bee1d76d4787348
z9901bbcce37ddc2b236cf46823bf5ca91bc04879ee2a405599955f8c32ebd644008a0bfd2dafa3
z9c2184a8e1a1f253b7bd0feb9091e2710c09355009290eb7f55175f2e8a04eaeef9d729dc9160e
ze4a3df1f3de59311bd59044ecf3c71b19b75e891da65b136b78d3a8dc947485d1fba23a0830c1d
z5f0264baf41b66a6b01f1af14f0c4fc9c2787cceb8cc3d6c54a353e7c308937fbcabbb91c7827a
z34b4642b3c3c14aeaade7369daec6e5e6a6b0257f5b284f45f19d7926e7d2b3e790e9c3549bf28
zb7a35804af51edae4ddb9067968e342b7cda4e1fe77b1881d02e5c604473b129efc047426de552
zd79db0573d08eae0c7a005110d89e47742a3564b6ad813b443e1e27f4c0400ceb1a7b92796c5cd
z8fb78264b745e463ae56c492258c340d036ac072f6187f5d24d28fee322f8809240f0e1087a450
z87bd5dbbe3ffc5ca8463a13938c6f02ef26d6a199e65e4709ab687f7c2dc3176120f27223fd4e0
z751926a4fc68ec74cc2871be9f7e98a1f63e0ccaa2b384fa77c4dcd609fc03666386cc06509b1e
z2fa114f488591d2dbba140494f450d7c3437ea5b3004f6a8b1bcb41de30087eda81fd37698f958
zb82d15e1904c9ffefad0a880358c23930389c3cdf00d29a023096fe4df6988d5577f3e12f21935
z9afa837570c22d5e901539a09f4104336cfa3e661a396fb1f0c6791f2856e2bb425c96ed0e5ab0
z272a573e8fee779fd50d51eb841f0d5ed1ed6e953de73e8fe1dd6b027e306bd5175410926049fd
z54f5fe0889c4481c3bfa813bfc00bd4c4b90db404262adef570738b8868845f4355f0afc140b0d
z70b8fbac8a6f294362ae99665f7e5570795f1b21ca72bb7f6c06bf4c53aa46d2d51fe795acedfb
z371bdd0bf33bd79067a7eefb68343a0d8cd8d51bfc920d08e464ead85072bf31d498217087d87d
z18b16eb46daad718280ff84cf775a837d3b2eb7ff7af898c86d08d65d2f7ab2756c266d307060e
z9484f08d13831201d8bddc40bb75a0f020f5e54f0e2f7177451dccc636c9f71274bfe1ef3e7221
z4051327474ae4b465ca9d55f87127a1fba974bcbc5369bf1489aaa40b16c28ee4c572579081e23
z3a212c92176e9142fa2d0c7c0e6d57a8049966978fef0bba9d8db8a8698f9afb4bc10747cc9e77
zce1adae949d07afe03959f424e3bf7b215d913871a8f7974dee45615e98f3ee92b3aeba10a16e6
z0b5a4697ccd44850cdeee319c9bdba851c8b6994f9f836c5f3e440084e97313534130bb602f459
z5c139a4875ed6f8b477d408efa55e57e7c03f036486d9a41a9f9cd9bceedcc0bc7268ac29f9d0e
z7cef126f647b989da109bef30305c78c01b977e072da8917e7259cdd2ed8bedd6d1c2b638dc06f
z94aa7c60e74c6936ac369f83bbc829c3f28aa23ef5e38ee1065df4a86427154cbd5f0adea9a59f
z533f5a8b02b173f3ed890b14f3ee8a99346b33dd4f55aa74a182c4b6ee833068be106ecdeb6a35
zcbbb42ec6827cd14c77f858440e7564869065fd94f38cf4154455a7b04beed4b4fee06e9ffa755
z2873e2b119d579922f3e7101cfd70b2791107d3e7f5c4ffdb280c7f62e035693819774d2df6d35
z2a71046ef6cd943d2a30e3dc3021f84e33cbb662286a315c253d97fc8b130d36dcca31630e0ce5
z3cbe202cc2c61c24ef07857cae83491374cf8916122b0f066b34fe3db5604739345880bb8fae92
z7d08d1efa85bf04d696fabf0f700558c2063345fe5a38b322b086a73efda936b3525f2e84451e5
z48f29fd4f4e8e723ef3f364415c289fedb80f514dbc4ed4f1e7b3b2e261cf5e7825f797ecc632a
z609351ff6924f8e64ec8d90697f5983c41de97a25001961f6dd96abe6cb269ad625e2e121e2570
zadea2b400336b9541ee0d6e7b5a2ff8c408bf3b3d9bb2c2ee9e56f397f0bb51e1539ee6cf1b2cb
z7ee954125415be22ac9790a61e1f86b39d3768ac8301a78427df58a29f184c0f1ef4b42487d451
ze3d32bb1e211c918128e25b6cd0a8737204caf0e9d1942b11ac58f3a4f0570cf6af4e2474be6f8
z58843f475ee6af4f84796d4614aebc190929f8e4769981004bf0dadb2dec0ed4636b6c3b0d7f18
zd531823a589aa284ceec99f778cc23d9762b3d7b7847b619bb4f218b1a32f8b97a84d3fa01493b
z96a6324b9983755e16f1ac57d7d37d87d67b694e1c1709ee105e6fce6321c25902ac7e39d922a1
zce0a4281c521d12aef5355fb76497db89a846c384c166f1d344d9913cef6d50e34c0434b1d780e
z9f98455e21a1ef4b3724dd607450795981c3c35eaa38d0031cd37a36081597b852c00aa92454b8
z1ddd98d9495f6942910f0045f780c7546a8c0b0ad30ef23a1116d6b4b3fb01ed3f74e4dcc09482
z9f8e2edfe5df23d4dad9f7ba9a6d96f57014d10e1dc604e20232ce8833194270dd6c73999211cd
z0ee78cb5d50d4eccf0806e5942b97dc65799783b4bbc54e82dc85a633a85491813e173ebd0dc16
z0736908363b00c7f5ab9e442119249c070c4a2ea56abf3ca4ef146ee1cbb987ac95e1d8993bd10
z27814ecb541273dcd9ed966c1de94bc152309e49bc30bad2ee3a49b67a27f741d08cfda8a97ead
zdb4f5a36a01039e79529a264a1a85ff11e0949e3eea95124379a8d1c267cabe311e780d952abb5
zf0762cea9811c2a5f4dde62e6be6aa251fd364f96249fc70df66dc78c53ff444c6083bb18b3eeb
z5c9666b2d17e154f8a6cab0461ddf4a8ce491dde42f69e4244cf5ae776e591b9e942f6fd4203f9
zbeb358957fa462b69a2e90818e79134861db22a77c5f07ebf220bb21db374073ecf6c1a68722c8
z50fec032e0eb17342b26657cc7122a07ab04241eec02dab3ecdf5a6d9bc39f6796d89f011bb9a5
z0882b8ab5355fb7d4e9ab7da6598e92415f262d821fac940b14f9d1b24c7d746a5a91d1a450c90
za3795d2c166dc662aba299d50593abe207ea344ad17ed6c4d0ee39a6ebc189dd70892b6092ee6f
z7e78aa51caca075dd8e8670051eab094df5d6814602614652251580ca24a8c7fbcf853b16f232d
zeeea2984a48de451aedbbc0511bf13e272f1d0f58f225bf14ab5fbb06bb9757e9d47836d5695cb
z582a778ed72ad989b3ee12085967b921ad7e349b7d4d8b65e821178170f06253d35d3b5cfdfbbd
za084732f77a3aa23db7948bd8398d67c6a7d3a38213a5518638216225d15e85c65078dc28a800b
z27248ad04a8fa68f7dd058c80b8b8a42620b0c57c648b7ecb158d86233fc147b87e8d8937fbad9
za5bf6cf0e50267406b693ee7c1c5bcccad3764fb8e3ce75d79634ae6f6180d6e67da5a0ea8bac3
ze051a52b44877f4a8ee75cfaa66be55a3fe66a81408984c106bdb38638c0db5646d0b88d46fcae
z168aaace40209aeee61b3c954e5405640ebf65178ae94b560b695470bf43116d88674852731e5d
z354f1364190e938f8542e53c851aa324f1e6b14292092d95f9f7bfe000d1869f6898cf073d5dc9
zc95d597f45596254c37fee876920d545cd20693d81bcda44243bdde28fffdd236d2538d4e3f9ea
z6fef848839112b53aacd6d8213828b4098800f60274c57c282e6a17f2c5c53fdb1f908b052b1b8
zc39634e845280cbb853243cc3d9ef6b28a45997f4b4dd08a1ccedd297882322f6ba947e810856a
z0bcca2f809cddc69c277ea9bbea03d945e83c0b9035ab93682d6d41d049b345b8280fe235bbf79
zca972a2922a51670a16c96cc74535141b639d348b816f6676b137321a91cfcf06d416352a7d4cc
z943ef15dc34a9fc1933e0b7d1e51afb10b407b9f54249a6368c7188ace5c5e21e0f0b5449f31fa
z53ef2a89f475e2a5c3e529c0d5e51334e4c7d4b3a54ff9f0a2ff93da7fe6b9b2a647b4dd59f3f0
zc08efe9ecf6aa9e5b95fa4f7debb09cfe931d0f3e4df25fb6ce6b4c1ee259b6a4680aeb46f51a2
ze9aa3b7355283017f5f3bad4864319e73fae9bd1908652e1ca77e0a4c9ac59eef3b03acf26d67a
ze9babacd80f221fa43948f0900aea876372b33f75cfa67a53a805825f439387bea33997c692929
z9a80ad888192c89ef18206ea07e0070b77ab17eb55c71235ad4e561b7eac6dac8b8b2b2f1f702e
z38181fbffc3f0587eaf7cad4cd51d9f40626574a3506eb921c97c7804061ac03343c03ef8f00d1
z6345bd398aeeba74bb6920c4345582d4f71825ac75856dfa8f9c748d0b836786abdeaf32bf5ca7
zbc0baba5f9a334933082a6e3b14c04ab24da746c3476a8ed344e6b7becccd20e4f8569d297dae2
z8985e17ee920d11975752ab9096e81cdc5e4ba6a82773f73bb5788c73204275730d1d8b210e84c
z4d9ca63104881c64d9c262f4225fd1ade2cc50f39a01c2de60e3023a0299c8f42440bac081979d
z4b090c6ae287ce77d014c05c19b7493edd32c0ef5415363b3c792783554952b2e3640686fb6b3a
zdd9e2b464cdc0df0dfc4774cf056d0643d94b4bf8e3b7d05e47c1daaa8a10969c987a723869db1
z47373eacb5a2aa0cbcd5914673efb01f2cbe40f52f9d41e8d25dc3269045f486e936cb0c83fe3a
zbfe0f29967a273152609cbd35a3ef1778753d385e6f26e24bcaa95a8d90e2a72478ff0c27645cd
zd4e644ed1de164ccb8755d5446c756a9fc18577995ed34f489ce9c9b26a337188d00f90ec6c885
z892f76bafaa1be85d452a1605b9c3db483d22a667c958249088604e5bc1f0580e71c117c0c0d90
zc99044cef5d6dfde74b8702f87b8cf1891625e9445e8b82fedbe1ed6e097d860b6f2dfeb9a366f
z6317e4942775e5353eb3aaf190fcbc199aba8136d48b4fd0976e56718666a27f7a85dbb54b8f7e
z5208523ff1abf900161d9de7e8bb762bfbe37991d2cdd9dd90e30d3dca5e04d7455a0bb53c5892
zacdab93c9f3914e41963cf3ad419ead34ffda72f55a4966a9008fccdd2cd0b017c431542a9a4ae
z84ec3d00c4702bc20a16e0824c4154ab72e3383d29faa46054c94b19940aaae15fb1a1006a10fd
zce5bfb74fd175d3590c702640d7754acfbcacd0125b3d6c804c9c9b616faf8385f8dac50935570
ze9bd57645cd1925264d9dd6b2ebfdb936933e6a9eccdbb210fac524e82fe15186a1a1ea83f90fc
zea5eba96e133b6d90dc59b5c763328b922702b79a672fe160d4ad73f5a1b5a144ab7d0c2e4f1d6
z4d7ce0fda4f2dfb622612e20c253403e1e58ba610e3c00ce416b7a6ca822fc261d7626124a5a22
z28ba018040a854e91c92599d9d3a748e99fb396c65229dea9a1789f6c4f30c836d36f35d171266
z6f97af2bf740e61d64388a993d61496b7d8a1829cb10e6bc31e32a235b1ccaaa751219279490b4
z771ef3b2dfeebdc255c70ef98c202ba4d83b9d1faf291711dd8aba42ee48d1b2f9c90fafa5a184
z8b33ac16b6314d803e377cf33cc6c7de39d6975f831a56d286f3931e0c65df738bb3ff836825f5
zd42d4a53320e6ba00bc3373e2aff790042287f4bc3154915891cfeb04b74221c5d33f4cabbfa4d
zff5b4818b02275f08b2f4c8d299b053fb1667d8de345b7997f619c064e3ff63eb6888041a97810
z2f027093db9241b821725a5df67c9dd557779562a1263ec78ecbe62e9ab4846d12cc11a4ac16ba
z094acb237ca4ae077b156ef11b19fe86165bae54bfe7c813e71008c2cf66784a22ff909bee464f
z878d24814a53dcde36230458083d3daee8682126af07e4f40b6dbfb228ac15bd28f987e1a8d3fd
z883194b3b7aed6ebf24fc35f363358eadaa2a73b2666248a3dd7218acb51b7dc07c0d6d8875296
z8da71591e5d29bfd496c9776392509aa797214b521fceee7dc67168595ff8d573bc62b86f2b24f
z4a61ba6350af59a340586a0943ab023fd52531ef137117faaac663d5ac5c0ed883bf87a8296604
z7d7cac0ed9931b5d813c8d14dd65bcaba660dcf70e0795aeaadd84b288b50655c6f52fd47c511a
zaa6700980493dfd151713ab426ec06bfdd6a0d9c2415ae9b0557d89d237c5897da7fd4dec0ef99
zcb4b27d2865afa17f435dff426ebde629ed7183165b76d5ff52f5906f113ad79291819a7d0cc7f
z69f319e7040c523e549ac65dd8b130312130a2815a15dab1181c021ab4b75e1a0f3d1201f07660
zc79a87712a251bda29b42d9a191f54d5202ae0065786fd7e076d66d0cecb6ff8ad306768648849
zbddfef3ac80ebaeb7e452263e44b5c83c386107a3d099b013bf4d9cd82d5c37ff4177252230e94
za3081d26116fdd4939424d6b6c112e61dba5053ed0bc0c70048dccb61252d7e6b1134272bbe375
z5e215c8de0a8ef62c4450490732b4a019739ba5a95530fe64b3785d97746f59d24d56169186234
z91bc164a9f310bcc1ac9c5977e161adcf9d9e4190127fe35b68193e841e7ceccdc066414e9bcad
z6ef9edfb2994bf2c1cd13723c6bbf8f5c332765a90d1104ac7f8a9cff2ce4f06662b81f4e52ef9
z4e463647577aa549011d1e9c803b5da3d9e8ed1aebc97afa841629d342c5a67a39556dd6b1ba99
z1ce804d73b10766b7787ddbe0b163881f1510db0b9380afcee8d40e248718319f9e0532ae7f3d2
za23a7fb16d4d77d1d21ac556208ce41bb416ac6a42126b62ec19b63224c960b39b31c2304a3388
zcd025b22aa1aab39b34a291a81abb0c44d30863f3e568dde2bef460eefd90639863dd00d5701bc
z70f2547297c0fccc9686cbfefdd4a03381040d7b62d1f79f0d229e984ff11b58ac3037235c9c4a
z321d3d9156efcb38ffa1d13344bc206eafa29cdf30fa05b19b35f11a216a5ad04262f6a1a7dbac
z919ddd7320ce89e3271c11111156236924661c2edac35d765f9113a9c42885ad00e36beb73b3c9
zb0a9c1a0ac47861860d35188b32f3279a497a2f17798692627ab768d797a68fb06e4089cf8ee0d
zbad2d53cb7e08d6398b39e0b7bbf5a0522e19bd0d6fe9bb81463c121cb5dc952f50fdf2656a89e
zf1d5f83db9669d718670c98ab8a87da05c2c1e32f87456ae662307ea636e7886f66952b6ec3207
za2d0b4a6e96b6f91b9a8d20cd4f6d0f68d0339201917700857cd30e727b0bce2288f3fe76529f8
zfb2c8f8070015d66bfa40ff849b629f374a5d042aef4a0e3f53f0cecc92aad129c46dfd5963dd9
z86261d1f7ea640e81f5440d6f85fb08ffb7213213679f89db79bd0c71449dcfc6577265469f147
z4896d03ff637160cc6f902c5841e5da0b5d4394cab5ec94d0686b5fcf8b06004f14823c7398de1
z41240cb5da7765fbe1ef43cfba93149e533684cd385a083452f30b8324339d4266c6cf23677c07
zc652e5e9aecffebf0f5ca5d72cf8cad0773ad888c42a7760bd943a95f3087096784190b2c14f6d
z33caf7cf5d840c4c956f4294b9b7caa12c9a3e2cda76e1282dd0ab149d170802bb4da973c57ea6
z034bdb639d3a75f1517e50e41a078cbc4fc9acbce01bcb4163cc714551ff1501b12c6aad3589c8
z7c8e9aae2009e5be76d83cc51a6f2d29ef3e283248688787994af48765e093ad2ebef60e4ff026
z530b1c70ca619497a0943b2840a73b661ffb695542c7806f766ea860a11b2df8226a9b277c45c8
zf989f1614bf06bacdea8372cfd558e5f0ea54f5120386da002e7fed1a908bb117dfa6bed9f046d
z580f6213969cc9f0a42450861ea4e5ac9d3fffe0eebabfd7b0a9e7c7be15e4e65e119e7555a8d2
z4986597a30500282f50c968a9f54dc6386f405d0fb2065a3700ef72ed05aa02522e35630f6b0a0
z5eeeef1ac76355de148c976509bd1bcf1ede6ff32eba08878ff31495092e907f30c963d70c6a0d
zd88eb8076cd956a1618a69adcf557d03ad15c28e400bf097b2cc74656ce3612960a8a993721506
zd84533c967720876c9640f7efe006c423f4f55df97190b41ea510889a28172dd5765ca346fd4dc
z54494ab0496e780eb6bae1d0ffd6966264f48c09ef5ed8706365e9c21d1700af3578a446f50e0a
z31102d8fe422fc56a25e902551b991c3bb5e763e23c21988e592ab22cde5f6170c60a4999b1834
z49e2fb3b7f20dd3029b52ece01503d42f9d5f9cc9d572ea3e7fa5387fbfad40d8fe3069d10476a
z0169d516a83b82d7bb683c77d1e9b641afe14c5366861966f587a85197913a996ed602aa686808
zfba86bcad0ae3fdbd4e37a3763e6202f9457fe9467aabcc90bbd2c2be266afc0e1947084f5589a
z969c8b40faa08a0bb853db66590eff34bd6bee24565e4a1ff63befa022aeb5474d1e8bf13eaeb9
z54d896b7b1abb1b6e4be983bb612de8d70db356db3bd6220acca0c3c2cbd11342d2ce02bbc3fd0
z56fa0e7b98b7939bbd2dea6647f71a8748042a15fd805190d0388545d9af2f32fb51b17ce28dbf
zd0503c9c899ee10e479c056de32d46bb14bc776cea5380a2732f34bc4e8416c5b8b3c2cf30b7c8
z8be92503f0d26521859f4b394d25108c33b430ecbc88108e8ba0ac14436fcc99171a55558a0543
z75c0a98b8a7abcd8c8c2e7ffea7c9992c9ffaac2ea013d2bee3718c61436e1cc5ad32a30e8f130
zcaceb3fe0b3a2420bc135ab5077e43b0e10f20bbfd7720799c578a8340ce8c14398b338e97edde
z44e0807ce829b711fa4aff35ddab21490f51ac6c096212ecc44c90a30e480852819edd9cb6e563
z827a6eb07965ac0a0cb3f1316b3a8494fced1e600372e73b62301254cf38f112bfffc078846f93
z72adc83493bb3469f78076ae7156c2a4c4c83edd3c64df3d35c366b99b97298f704dc08b7a4189
z6f6404f4cd5faf8bccb5e65b5192cc68c1cd7a43eb621928e28c33a503ac32ac66fcee4a0be48a
ze2eb00836b027e0e7dcce58d35dd1138f7521961701d9e73844f3a7ad35b6ac9dd93eb24791741
z83655b8173dda1faef9b683635b2eda089134de70c1e31baa1598cf9b7f60979118eb4819950d1
ze5f79a7d2a6b9982fbad86ec3170489d9185936ac8105a0f777ae9532d10620d29c298593b5b55
z40931c9151d35916c076ded147458921a8bdedbf2905f6eaeea898b3dd1edfea31fffc6ad56e1e
zd5212546928784cb741addaae31116c00d3edeba2fa1441a3c2aa46b53306a34b7385bb9f75493
z39443197ca0825f7d25fbd272d71dec6e6459f981424294a9eceeb913b46721e4443d1177bf2a8
z3be1c9d114f51a13dfeab0cbf15d8782504e26005fabbad72c290cb026073d7b431bb971a0bf7d
z165c76fe8de516a7854e5848a06aeec8cb07a5190f3b44480ecfb90a4b27505c0b7c0d5cef98bb
z7e8aede9a36f9f2dc54dff5002b12c75049256bcde1d30eb696a6d6d0bef7d6df6f5def0c3283e
zb159ef5d6350685158aef458002b2ec982028fc54fc43f528e77ced448a79b8bfedb2d60ea68c0
zeb9787547ba11cb0f6ce0ed7f2e2ecd3728956067acdc8f30c00db281178a192272433e1cfc7b8
z9b4fde81611fe038cce8b538ff1a66e1c1bdccbc2b7e35b361e093a7d51ad41e74054f101b0900
z6df227a9b39a6a59b42818e2b0d5ab816eff710d5f801cd31c5a2ed9fb30510abd5405b28001b0
z226128fde42dc6821b268142a1584ee18218397021399b794010d7359cfe3704c3b359ccb34961
z334df290e813baf809cbbb122278e7e2e6824bc9f5e7ec2b2590603741b9b1dd80620b0bdf993c
z2da3757bfd5a2205f608ab76383bff184fbe0a2cbb9eb8ce496b4a95ef203b0ff6c61b74307e86
z3d66858b5fd9363214522b44c44271d1d9f176e0bc35c6b8e1920a1903bb774cca13b0cbbf0640
ze9c7eef793af85741fc4d283679a315ae3ef9d131a6a1af7970cbdaf0c5ced3ea2a865b3c6b09e
z8dbb003bb3c384a768b97df8a77578430e5bae7b6c42eab1d87ca728dd17ea0d5d835796963388
z9f748f011dfd0c9968323605ca3d0ed51f8e179a5785e79520d1b8e7813dd57129f0316fd396db
za306177f6d9fba65be255608a66268f4ca6f3af5ba6c3f245771990e464ec761c391a9699f17c4
zf4402c1994b2a0ed906b12f287284a60c6c92c450d9f87d60d7291ffd731427ce952af7dd0bbcf
zd6f7f7d0d70b534cbcf476b2bb311fe4245018010f3d89451c1678b284e4be62a0e6803ef18bc5
zf33c82c1f50d3cd3e2e9c654f9faab5b1b06f16a3ab1eb69d6f8ab1d74a89e50144b9113650709
z385300b75a8926faec0acbab72ef8ca60573cd288d5bae181dadd4fe6a1534785d4e99d8dd8d2e
z50a3638d3ae55d5ae5b4b44731c1ea1063bd6123b16f4ea5da4f33c0707a1d12a81c0ee5ed2b13
z1f1ef2ff9b88a7d9e2214a2efc02ca04c719feb72a93dd7a51dc3a9a0be3f1252cef3181ebeb84
z758516a09f40c8803f5c9193504502d7db06ec85d902e523b6e64e5db169cf19dad081ac0e51dc
z08f9bba885794948a0da41e0b3b3022fb1f2147f8c591807bc96939cd108f5fef32771680d2bf0
z627f9941f880c445f548f4acb0430e03bc707fc003c46eb45b612a6d4a23c6973786c5217bad65
z89d8f848a508fa4df7ad92fb68bdff37b3a846ed09586321283aa9a25d0964bd619578cba709a1
z3e8f8ab518d8123aa54c8fa85bb9bcb6400bc16620edc7ce402002be351c8d5926ada455bb962b
z16bd791c5c351ce1d80da50a8f85fc2903b501a0dba83638dcf06d45a43c678a11568cf1edaec6
zfcb136c18a2d4d575c2fa71534bf72e1ec847aa7727d448d11fb8ded49b0d81102829cc35a37f2
z95599f9e428e25dfb4f67147ff7897c0f521a2144ce308ed7562c15e3e02c833569fded1ea9416
za164bf76228a167aa806e2df467c6bd16d4f53059491a8163c4b5ef252406bcc7518594043457c
zd82dce80977e4f59a662ae0623179173fcbafc8adc52911f343e7c72b8bd9443ce4db853fbdaa2
z8fd2aadf802a7a88e91c6f0dad9e810230a696e4e93924096439612d47f716f4379b0beedd33f9
za44e53dfa21248bea433e45bb4945fb2a44970b9cd72bd538d463ccf11156d09f47e5607d0862c
z51e69b93595c63976dbb657e5fd065a34daaf3bf476280b4c15f05b8172e3259bc01abae3c09c7
zfa9dcd194ee198848e2931c32d8030ab3b220fe3a6f32107cc0cbdf93146e03b8d60dfd4487114
zee688b7969edf92978d554e19e0a0ad09e19615bb4410a408675be3750ca4a563f90391dc7b2e3
z82c7c27be03a3802a34c0737d7b7e3f7f2e653072cccc40642f1a8c380635e023c80d23ba87234
zb3b8187063e4dde15c6aa387a5da4df0717edc7da57bc48f9072af783517c69ac19cbf93ac170c
zbd71c07e89ea3d1ff800966cb323182d6d86e150205e84ba7572e8a2fd709f368afdbb21994e8d
z5e511fcd22990a873e16ab6b8a312ba3c4e2ad0794e7510fa4f67586d5ee39a0495857c7ccfaa9
z230d1ee12b32af875e0df00cf5d896f1d64bbdfdb93fa9d1b90e0a376856ac990d027b990cbda1
z218e8dee82c16410e5d98035a82f36eee1af8d239353f07b6172673d4e79ce62222dad73fc7cd7
zed73bc81bfb1ec77f8b9f6484fcc0ff1b94750d4b238e80ea738ea89bc3d629c6c8467c44f5ce7
z01c1229e8f1aae9083adc2f910d2083cccfaa36be6c7450b7e57cda45ad015e3a4dcdcbe794840
zc51aec0d4697aa7a0fb898e800070aac906b344d368ac340c05b3e53689d4b0ab914574d3837d9
zc3971dd3a1b9ff854b795c39ed55b5b9fd2622711cc3f54bcd77694e104748836537de284983ff
z89d6c04d339b107a2293f8e691612f7ade76c4c0e3da67392cf6300746d04f106c2ff7ce665e0d
z96f4c402441ef72cfd21ba614f0b92fc3f7bd53cd7d27faf24d50eed8239ef5b3cc3b4338980d5
zbf92d086178e9119b5c140c9e679b0a787b20492a34920676b2e975b868dfde967f0de96e9c964
z83b2ad26f38396ef0fe490317b8768dd6b6ca992d884dda75232f471fe17fc9d8ab0e6e50f135e
zda1a4a02ef4ef4318c654f680de5d1d270cef86761db6464b69fd179981c5cd90a2a1b613a7095
zfefbcfe14da059a89814d796753000a16ce4bad0e2e5a020d9df86ae8186a5165f1be6933f095c
ze655b0e6e6878a7157c80664b59c4a54e1f7e236b75a5a1eba26bcbc8b27af8a80b70463a59016
z0320e670ed96e215216a36ec1651cebcd71e32723ffe84fb8bbda332ec5b5cebd18387cc015ffb
z3ecfb549145962318136f3cab50da866ac696ceb2a810ec322b63cd9382fc0f735d3988e32c691
z0f1074aac73f329bcdc2531d39c3bbc3b822bc8703d1a97de31d63348aaa7ffbbab20612c001e9
zfb95b01a9620be1e4b42ed260f56f7050b8cf6db4f986c5f922f59e359831ac2e569968dab8109
z7fa9c7c4da662ce28339c54a06055e785cd5e998fc625392c712e8b2a403e8209040f1d4e0ea2b
z3e849b44ff991e085305f1da7e8500c5d1ad6c96ceb66cea46999c92f560ffe6621fe10542a2a3
z74dceab5972c8796936932457cc74bc88e5ce5837c12d85e852cd6187142a6f97bf73719d19652
z89366fabd8dd2548bbf5d685207378fb023e3b8a3d2126bb285cd629c78b12f9c4b854046eeff5
ze31f268d526729d99af812b329cf3bd52b71df9a3531008a0f870200719f505b2e29f23100c825
z5dcd052593f2439b7b84ad4f58e95992f968d7ea7f0750e574ab9f1e9866b07cc283b9949c9d98
z445025f5c5990d87eccaa85804981cc45bf776f6042372f7e932b920a6912464621307248da18c
za642b9eb76ea8e9801d250a414a52c7a635ef3a8cc237c636b580a32f9f0efabcfb2d6a62015df
z13aec2ba6309f326a97cff0646d7d02a7303f8c4805b2026428f5331cc5df2365ee6b9024d2674
z226e010fc359acafaea77c1ec06dee118e55af2d6227200d53cdf4679979717dc01beafb42b01d
zf22a4dc27d392acc41c560b67a2e101a700e805fd1857a6fc49a55a26fe56f48eea961ab838d0c
z2a2f130ac35d34c48f524aaab7305255af31ecffc3f05ce30e5255ff3a72702acbab4bde9999d7
z4a1cd69b00a6b04dbe59db26a67b113eb86ebe5bb7df4cf49d01b6ca96f88d6cfeb88afcde8696
z8e11eaec522a644144f27ddc7fb53aa22b4ab3f39618433288e2041fc24f26f74dd8555228c1d0
z2ecd9d610236e697fa6cfe399f5ee3efe60d9df4b0de54a14c020063780bda25643afb070a18de
z326112a97ce806dba057ae6351f02c3d2a9c575d089a6373264082a074c51541e74e76253c280c
zb41cae046699e4c304f416f5d5224d0bcc7e9f370bda404f9529a2996f252126a29690521d8025
zfaeb2f61b37a9c36afa365a2a9e6cfbb46b5faeda12064c03c8a48f857b7ff8fb43249c31c00a6
z76e696a8e34b75e971b1c04f7412f12ba8fb332e6e54dde9c213ea009e9951fb37df71dde6f2f6
z8b73df60a51e8bbafa78da1e941e3fe9633a642ad86e16d2632e5750c4672622ac2ca39d351e67
zda5ced9c59144f07c946c09668e06414fb7ca4b1ba6b655a6cee9f73abd74cc61473b3b1abe5ec
zaebf440e3283a93f9c4f5c4569f2db89e1827d05577105066c829738560554032c0e16e79f8fe0
z02fda9a7f7c80c7b720d87bf183a73c2d68a0737b58d2baa5032965c71691f76cc33a924879c75
z5aa029afb9c676f191a8fc2055f14b4d37993c68b2f2f3063c90627112bd212b851ff4a5d8f267
z9e7832951544b049edd7ec4d2934aa02cf1db4743cf6e8dbca6016d9c16d9901cad4c93f635bba
z7c7c0358d9204143a6ccc1eb89e8dd2e80902395e8d45dd0bafaef54a96b0d50f01d56cb460611
z082c4f23566ac34a46245c77a239c0803b02919e91ba5886715ebf1eca54bfc35737051502bd65
z205823d6683d96f452833be16119d56a293c56080ff25bb964f9292b452503bb224a0fc8bb6c5d
z084e07542973054604970186fba0b7493fdd6f89784513001f24cc4a27e4ec4c1e812ac624508a
z204d4af3ea77c27784d4ec469122b25f7da0f829e4feb198473a3de7aca78ac11869550da26fd7
z9f4fa366d11b6be78f27f1436d21f6407e068f2563ff54bd6d8a3cdfbf78b6fbfdddfa5d60449d
zdcdb605e87c245fad0521c4ce18aa533b911e7c87ae5b053048a8f5907d0cbd4269593330881a2
z6a6ac086db18fe0ffadd9832497601c7c86530d1fe55f3d13408f7e443a2d97b901c57432861cf
z8bfd064368b4428db4bdf35554e46b5bc9bbd49cf9903ae1815cd33627b6bb62f930da5ad4c7d9
z3e30715a9187ab750b332e0fbe7dcf7e738ee350cbdf5d8a6ff8808641df376403a0f5979c8ef5
z22042765a264183cf90280568116caacf1c8a9c6625ab0085a4f4d1870cd457e93754ef8d65741
zb7edcc5e1ede01b729a3a75c2232758e56cb9b97eb053af8731ecd1387cac5e5672480300f0b51
zca0111d733c711fc4be2ad54c0464b5bcffdb8fdaecf07e1979b7ae8af8f0946c411aa973b3804
z39ca53630875e4708e1c32916fb1b3c47b774b08ad2a30a442220bc1bba772d453dbd25e1e5168
zbede25fa819ceb74d94731e677c57b09628584a2509b742ce7efa5d6b65751b2aea4c55df60f0f
z4be813399f5b1281ebb31a32e6edf277ac3d3427f68db019cf757e5d7b02cc4d029eb140b5330f
z10f521a5abf3501c9dcbd4bff2f3c658964c9cce8c8240b5f8d18b8649468efd8206f4b4cfb41e
z2b38fb4ef27db655309a181138930b69803582900adc7062d55af5c76e3b4cdfd8cc230551816f
z2fc3f7be02ef191f3a4e4b4bf3f09a7d979b0d18180ef837717ed6cf24a3f5873f44d27a0f9382
zba6a339a1e9dbc8ed34ede28dae65fa838e07ff217c531298c07f5a70d16f8c972016f11198c3c
za21d5bba6c8ca73b0f64673d9f27be58e28a3f2032403e351db955b6ccf6d1dc440f3bdf1a233d
zdc6547226f9ddd8badd711c4f2bbc9c2b743aba294e7facb1d3fde886a172f2f54fb86c0dcc98f
z134462118a2f29a2871ef2ffd0936f812a70f037d0db59d1e8d9cad1d3b6718e416b680882ef1c
zfdae64ec904111a64efe559b414fac4429eb429a4d18608c3d8a34b88e86c952d2271c7109a70c
z5c79f79276562433ba81573e814e57262a3568689a37ab0f24fd123536d14b52a32ae8791c5777
z093c8cdec6a211742b902e6417c523cd79ce0d7ebb5e6018aad5da20c101e3dd63aeb7dd6b8f37
za26817fae75d65a465da60e245bdd63f8d8717dfc90c175a7b0c12eaa7b2274bd8e80c6f3511ad
zb5a66c14ee397aa553d9369bd62479417fe7e01b53de9b4029ce5c71b80b4f0e0bc7ee2c1b5c7e
z9b5f277705ba082bdf81aa8dbe7a26759e04e8059dbe3b7ba6a41b0a92cead9c308f4261004b23
z69c110d12fc4f0bd1f6795605b445d1b16d19ae2ae404bfc1c4ec360b1a0d4876c37c03365dcee
zeb62936075f5ff8478d0f1b55c5ee8d8505a0eddf76f1d480be4e3197524e5ecf766ab8418389b
z225c838ef8c19be147ee59b66c1fbccaea6c0df25575c38233d13441075851b8d54dd81ed84a73
z79e1483414df0bfadc6dca49ebb65ef55d0f54acd2a3a59e34bcfc36f0bcb488cc1e5ef2b95607
z17b1800b4210266227365b70fe651c411b7ce0086e29d06ef416fa262944d55d12afbd70c3cce3
z8b4e91f715269ee1012e03d9c438f849dd863f1b6800c81734122b877b949800174d92dc4e5260
zcef01203811914f19bcde1801675e7bf7c1172745e01bf091af843632ac76881b6b62e8e8b3798
z4b8d16f65322d4f12451658b0f5506d474e680747d3486da8aeca5aa43a1b9b6dfe5559473a804
z596bc127b61df58891b33d7590f6478247250d0ec578fbc3579f923b9d6b5219d68fb5dd240f5f
ze1becab3956fb4f9ac30a9cea51b760fd07c5df4e73a02ee0d2338ce45b639405871f36ba1d563
zb59c95320736bf91d70b58150f9f697ba20af7df43546ab1f38ef891a0ac61cc896efbc5a180c7
z7c6adead44fb54289a551a4d25221c7398cea7aa3f8df87bf503790d347c8fd74614edb4f36f18
z94a7472fb6ba473979c24b1a43a190d05c877e0b075d6dbc2eae6c7c6bf837af1bcdfa4fcabea5
zaed0c39c4922bd5435c80c441b4c83005328f0fcc15e38131a7c73ef837645736637c4bdec63e2
zb9ef3d2f525fb1056864f0fc22d0a228d128ab3bef3bcc186d81841b0159743784d7eda52152dd
z570ea2db3491582fa4efd56ba4116115a0c2cfa4325b7959d9992e1333ca5c33282492c16d974a
zb1c7205bf34b2da620e6f04da766b2ec291e5add9966b4d0abebb2f801e43c06d258c0805eae05
zb1089e350d38a452402e03198e44570af2ce703fc4fedd7ad79f05439e3af47e6a160947758d5d
z552a39594177101264eba64a9cdf6c8132db400e6615b2acb2529d618d9dfe897e4cb50e79885b
z46dd88ef3ec7139af4244d9ab1fafd20de0dc2229efe77bb9beb0cae92a25e715a90d74bcd3c57
z810456dc81f62d3c4c65f9eeaf23d89383b37da280aaa73d25d8ccc84ff08c445762e1e72e4082
z9924042d35382dd9270ef364f68092d45afff1a50cc198b09d1fbfc09089283726798285c31346
zd3f3381126b62188f531de2b56d585f6671b68aa6cc6db8e49ab65e74382923d55b349f539b937
z83ebea73bb64c38d2edcef302766e4e0f85e7ed18e71f8f9d6a8a5c200cfdd90eb4ccf9a333713
z3ac66a70b172de2c98efdca3e876f0d4e5b6e82c9fc589cf31ff549675d1b471d0a20b4897222b
z723f231947d5eb922240222e70bdc4028c794eacc268a61e50e2bccd8f3853936a06d5b4c63fc9
z62e4359d68aaba1ba74c219dc55bcafc6992b969e79b607b75b3245a3b47766570cfc5e75fa1b7
z600a441e0f515eb35650fe97dfb5cb216b1f9e0fb5ac04f1f22c01b646e6d3b2e95df336f108d0
z93c1108152be9da00f5bcae3eb6a4d036cde81a00e09b7c841deb8f571ba7af71594ff9140e4c1
z3cf0337346d635e35932ac6b48980afe0c6c008438a2e16b0d15e1f6671ea6a6d9d14f23b3b5ed
zdc3ec7728e8302c60a93fd3ae8843eb829924aafcb4852a7fbdbbc631a94c642334c7c49ec9b7b
zc5576cf4716f34a410722e94420198fefe1988b31f7cabdfa4a7f0693a968c994b3432376d2a1c
z1c1e7461cce9d3c2487013a8569d01122a43a5349b49330dc8c4cff12a55bfc62ed4584b066631
z753519af9db1dbe4e73f53b587c55d77a4bf2da49f09b7be31fff84172af551967594fddde985f
z907b15b310ad125153ad192ee9651a7f0a3156288140fe3390ba527e733b20d4b8dade6a3b15b3
z3b4e97b026370aaec4abc0cefe1fd514976b80194091941ceb148213bc740d819a04b535d6d998
zf59bc7d146b9e949975f82fd46aa18ae3a760a768ef9c2ae10f2a6e6394639c684a55966c60a2a
z9cce1b4792044e8054d53664db1da7a1d7d4f8905ffc3796f4bde73a186f7c6d41bb05b884618a
z4e4de3caeaccae40cd9fbdfb471d2b613becafab5b59738c4811234a5a2f2582f0720b35551cbb
ze3f197ac900130d35ce963ade01f66db0bc89ed05d33babf48faf51daa5b9c25dec0f371395aa2
zaa4455fcf7fd10fa72d2c8e151e44bd1b99024ae4545fc58dd348ba52f06d1e7416c02b3d2dcc4
z7b97c1ca6ad8ebdad9aaae891272f1d1c7740f06aeb4b212918713524a391fd0b695a2ead9f294
z3222bf313a415e34ba862e62e218feecaa055d8950d421468e4bf7065e8a52d36670a82c37d745
ze293ec14c613feba8f5658e4a9043a70975284e93e1bd55197f330e7fadb366abfa7d924d44cb5
z47f0e8b1fcc6975c85c930c529c51ae0d2b065e84935318fe268d40e2f04b9e6ba806b21143773
z35baea03c5e901fb80f11c191e42c6c6b8876c83fa2cad9c6c8466b498504aad9e420e10f6e62a
z2e12179cf899383d0346705f4cb127e8cdcd94ab609710c7e6e82f478fd661f8bfc95255018977
z3aae5e7836a5086d18e349fc30537d6e4ed0eaf06c11c7c43ae98556780243b81666e31e78a76c
z08533e83265c24cab739173d92db1b9e8978efdb6d9d30d5781078e8cf96d60d2a76bc148388ff
zc9bc1daa6f27fa1a1e0f00a6e2078a618f66d85791c68c330fb31fbb88785092046f763d1e1ccc
zdeee30f59698e64457171d0847b18926c73e81c4e49a689742b100904e84b90175650cb95afd54
zd269647cc5b3c292904abe2cdf09dccc55c090ca2a392264182730f00985d1a995a273e57b287a
z1fb37795384fa011329c698c0f0e137519c3c83c87462448074e320c980efd5a0cc396bd13be53
z4577b8076feced41a1a0c54460b283cd2ef75d658bd60bd712f5a0e3907a26d8eaf0e8a75c8c09
zb380eaaea1a19c08366a40f4a741e31658eb4be0054829a8a0fa1dc40bf9bf34ad313361591b80
z6c56bb798af38bfc8a70ba203ee962a20924ed1d4cafb0f2c136794ea704a79fcc550bcf593269
z75f9166e95615693e4878e16ca27eb22edd4b03a822f6cf7c2f0a047eff19effa6be62c0e7615c
z0e18573fc5622d03e7bf45ea89aabfbc6037a12e56a8fcea72b267d7faa43cae00d69050d26933
zc35367ad214b8600235cec12b50ef7bd47c39fa23afa38322284def21a214683ee7a05fbccdff5
z25ae57ba84f160c3072a85fcc3a6fece817b1713b39c691b970d89f0675e8cc90e4edbf5d3b4a3
z044b345d3897810ef0635aa50762b6ad4f8a8d91d9f8ce006a3b7e22c1229dc9fb9f78dc066a24
z0d156fc47e90dec6c670531415330e53a9b9481dceffb62bcb296b4ca72de98b3858f05e5f9be1
zffa8b33fd8b122fddd733810db5888d91580daeb30ec7a68e99f1800505de73d37c3802d2c5fdc
z621085247a94136f97288ff01197e478d22332b93f5ceee0fbd0ef976e37aac5d3d772c99798e5
z12a0873933504d0aaeba42071f23e3eced2d67867ec3bacfa482d596583ed076a79841eeb4d6c2
zb5406910f4eb79074bc9a61a5f0a24b1bb3405bf1a4c6be41e4160f639828cc3cb4fb9a70aa429
z7c3a6624fba4efcd3b0df8f0996c5ca882f2227bc12017f6e9cac6881f30da80a510214449136c
zbc72bd8fac0b5d8654825c6abea977a31ca2c5ee386e6421d78176951e07f3eb66d68cc2bdffd7
z1dfcf6c62c3a1c064a894b053a295086fc9215f55ea47c70b9288e37c2692bc80dfff4338d67a3
z0fb86dd9ac81f6398d44ea92030993f9f5c44cbdb46a80f61771c24cd741a1ecef9d8d69629384
z961575adfcf65cc503b92e51c378d75fa0b0158371c1515e1606ff4e99b55c32f938ef5f9b8b32
z3e58f19c8529faafc29eb438b9f301c9550a31a3af8f8f7de488be26c571c87bb6d1ba8ab5643a
z03af93f94e6732af5bbfe49adc2771a23326e644ce83d3972e29580a34775c5098e26836643c04
z2af15ea25c51b04ec6de12b2e35dce103283a46a0be346c3185e50a48cf623fa57a624757dec7a
z75fed4c0e9aadcac9bb59037a959b4ef1078e7cf09ef5ded47fa2187e80204fc885d01e6c54681
z84a4b55e510d18a8fc0a488bc511ca3477b698ab59aaea943f3253bb24897c342a15eccec02a00
z5c5b6a4ae98ca236defa25911adb0b35da60eaa4bbc035f2a04a90e6d38e84bfc2031c810f8ea1
zbe279948999152c40f3f8a5028547abb51768e4f5e999480934a3cd97a3814b8dd9278b71ed03f
z89adfb3806209aea0bea205a9a15258489f0c40966b33e1423fc9a4f31a840cd5ecc6f9b3f392c
z267df05cc137b8ec1976938878f05343531517aaa2b2fa038b74f3122458c30ddbaa7c7e4f2f21
z82764526a7868e6edbb5bacf669df4caa0b6b45ce491f56f7631bd19febca953d1505eb199d7e5
zd63d8ec1cf44c1d641a051f4f9f673821acc0b53ab6302cb1b938dc843c90cfcb5b2abef36c575
zf3fccc4944da02b38a9b34d08075c15853a0cf4e191c563fc2bb84abd8556de141b6a29b07e549
z65ff8845322e076ad01b05ca4face2f0f56ed1e06c4d9281bd8da84c985ffb446da946d15b9786
zbfd79937d2a8349afa606bf60e1b7e7e305fca8ddb2d4ab3b259ab23058f9e163aa789a0c4acfc
z52044a7b41c550144597ef9caec624494da613d2864b4cac81110526355495748176abc181c5ed
z723260627e371489b35c2bd20423f9005d4f58cc25ee00666ac0e82d7a2138d59733fb0dedf64d
zc49ab93963aa62df61a1974b7c0228272b3ee08e5c660f80a92f9716deb108eefb4ec4b495ac73
z74318b9a0313700dcd31cf935418686488822818570409b4acfdb6a80e94e4dbf50321b11fee42
z4e022834b64f6e161ceb9b44515702e58d123409f9d385b3d3ba15820bf14376dbc8f449c82dcf
z1954e8ff1fae32c5b6a343e3241b5a477aaa89e060daf4d85712888eb05ad24f6b0b7dfb21c389
z6768d88a80ba393144c7ea5b581695f6da29f2eea9c9360a69f122d4ccc77b2e41c1acb2fe897a
z417a31e442f3d4db41353cae52c761d37b06d286812c4000aa97a792ec182bbcaa41171be3f98b
z04aef6ded30e0bff4ed7ad4dc1110249deb7edb643835d798731437e2fc2e9b6173d2866c4d1a6
zd45918e2ad23f5ae6490e30b6d315d2a5f464199d7ab7400e4736c5bb8d9a09841856ffe952219
z2f561d0f1a4f695485979b4162d656acc2b39c6cc3da311e6355c38ad4c06d3d87b767b916396a
z8119cfe69aa0a54fbfb38ba52815683bbd7aacdeb268f4338219d15205ce749517ec54993c9e6f
zd2d2f7fabca7e74ef12cdc2609327a9ffd85f11026899d8534a1790cea76c65d79e11487186d41
z32cdcdf7d92e25ccf3992f483e83d8c078927ef461f303a6bef227a77241a04c957747d833467c
za7239eb6bba4f69bc75c12c3cc1ed9ae02b56d1bf879fddc3a3ece416af9ded6b97475719e8606
ze336e2c58a916641e2ef14457b9ca410fa63876471a69070a450a9008eff2fb320a27712ffa79d
z170aedeb0ece8947dcd0f6743adf3baa9c17dc1eee1c9e8beb1752042babd2099b2c42ce899458
z858b7c9705047882003b4ca4b484c150807546e5b3bdcea269f1e55756f20faf2368f3f6c1e0d2
zb8039a8d63e92b42b7e4f3c7662673eb644c908128659628140bc453f876169b192a79204239f9
z7a1de089b18883b3f91a9f32dcfbc18d4a98f03329351878629d091650c52ec95e85839edabf79
z346efad569dfad4c642d99dba10b1e55766a1377b5b9cdd6739a1cc840e82dcf99144c5dbf0821
z45a6c5f86c66a4ed01de2e2b31a0329794a1865f6f5fcce32b9a0290c5b561443b46c35641de62
za9900a5c13318c5b3b59ff2fccaba1562c1e9f301ace7fa317a5de296432128d4b3204466cfa09
z1010bc00c1dbc25e7ef758b3ca864b1d646274524419e7d5e388d313ac58fdc5d12be4795ffb77
z803129e6750b10c5a99aaca91a46ecdbe97ba5ad7ecc7018a00b58fa6e899cc3253c11ed5fab02
z38465bf830fd8521646d691efabebd000f33284a01cf13e7417f2161cd02a8675e34ccb81f7c96
zf6026de476ccd9d034e568e0842de8eec05165e7517df7201e0a23b18597032b1a34f60218ff21
z7119dc1451eaf6bac2e55ae0f874eefe1f56ec84d2668a9aaa7a44ea20048abc54b12ba0dda38e
ze1f881b769019ac785f78bd42fdfa3c337d6684984784e999018329cdaee50fb2c9ebb39477104
z225e869c34279f6c65b0966aac433c9e8c777c4367a5be89e53df2ef0432b66f271556bc4399d6
z51d5aba0e324967ad2caa5188a37cf4e0164b49cb26d348eeca52419dc1ab169a9376c2b9c5616
zd17251a1da66f218c401b463ce526dcac91a6413a3b7f67da052e9ef7c9d410a60e5c069d4682c
zb0bf36a68167a0cf448c7608857e762ef64a3e19bf06678ab68030a3423949aaafcd9854fde9af
z4856c7551504e540c862265d963c681ba6e939f3677fbb0769985d7965d3b6ebf1d214491c820a
zae364f4623c54694ceca62ce235c78469b82b18537a24ab4884629ab2a981f237696e3386342e2
z8fd4ecfbb1e46617929223bd70ff61526545578cae5781db3f18f3575bb862b74abaad70feb926
zb15eca7a5158f5d6c325746e5740ef99070536dde63b9de396fe492a9e1264753a4389d6a8b1da
z96a9ef6da4c2b0b8e7d23b7590b222aa61b91b559500794b66f0d46ccf3fe04b4a5475e8fcd391
z8fe0602eba76dcf670257ce3e38430dc825f10bb2216c38899869cdc69a447d3726f8440807822
z7e12a6c68869a99a29971967b06f2dedd384bf81ef1ac424fbaec7761a509d1d3777d550b91865
z9c76269a2b0dc94d90a89f91ee672d96a75fd95b673a73bf7b729c0bb5fce6a6eb2fad0bc47e0d
z16f7a57f6b437ee69c58f0cf39e0992c91fa7e87c74468a7aa3a1944c95598231e965a8d9d0196
z2fc7fcede57528461d22b9149eca2024f3fb60455ef1bd6a44617644a378a44714d7dc36a1eb76
zd76d351fb3f54b4c31e8f417a11ad140325c4ccd69ce350130544c331428de0e36eb2d6a5aaa8a
zc226a8124891412b3e10b89cbb5b54ccc152fc7fff27ddcd737d03364a831d027b813f42669af0
z0cba0f2c959f00b40866b4cea83ffb205fe4e2f6ab1384cfb7ea96740d8b21a85e8a7e62215f41
ze1b7165b238f624389b705b56987882717fce0e700851beaffb13ba2f57c8599d81a3fd49a414e
zb08754cf307866c837c5578d1b8bdae198ab6ae5499038000518e08f7262c81f7fc62c93c6f525
z0456c9ad9e557144d95f402d1b49878bd11c17479d558e940d232976570d55014a0e2c71134315
zf9c987cae3579206addf40a21bac446b0f51db2dbfd821860228057cb82e1f974f57207dbd7165
zd06e03a1b5153a6253d047008462e999d76c1986e52f9d1b14503bf967d516b9812e9ab1dbddf8
z9c31b613bfa503d57dac93e535959a64a524986aed67c78b0bfd74663f7a803f8f914aa7247cf6
z190410af7c9b0946f6be267eb88f151d7c7f595211bf1d2df8fa703db8efdc4c8400519a54d3cf
zb8bb649b2978f632074b55f6e1123ee6ff1c098b1833f042d151214dd6faaed8f6de1d13d055f0
z415857201fd7c695de84e496b07445f75e82316a85072c68fdb698b146cf947d240d357ebe884a
zc0599db094b7d3fcd600f5d3a6fd43798c6c7248715773257d057f40cdf2df5b51cf48a05c9f40
z790737b8c83975b674fa24aba12854c1e8dcd41836e6f8f3e363257820e8e111a7be27d4dcb132
zfa24ca1a7328927c8e1b84e771f06f8dbc409c6ba39312acb00e5fabfb0cf3ee541ca609ab0fa4
z4e37cfbe50ba6a0d371a34cc4e36776db01913d5a74407405e62b3fee49b6a6cc9696b8625de2c
zfc0f2b5d99eec65160c8a0aab16bb406efd9d105a37ce0a9e54b5bd1c2e080d5f5fe3ca9f17311
z6a0e3137f63c7a8b4fc109c13da54f899eeb69f6f3a2370cec5994b795dc3bb576d263a5f00ed2
z174235fb8ec29ac401be599386a72a9ec8ecc5e8439de098ef77f96ae09dafad4d4939bf28bec4
z43e5b7b17349b42f5f00f5ae1514c9f249ee2687506e386de4ffce60105e3eb930131cbd90a924
z50f01be48c1f0be99503eea0b2f59bed7c08866647db3bce308ab7cabbb155b2ab718647efb896
z86a7fa269ed5b99beb4c18a5f808d055d710fcf4c6904b4c0e58ecf84fea2012fc13612a7fa0f4
zddebdfa4c8b43c96452878dd68fb3cb5a56467389c1a6234b14d07920938f7f3f9e90d969f4e38
zbe4bb981ad0f00dca178b58c1267577a8f18c89759907b9b65cef3aa969fbdf2ab8127fd2a731d
ze46073b6644685710f919589fc01ce69e8db133544aabc2630afe2b474efe8e79a2e4deed04729
zb1500e16207ee44ae565aa229ada238faee75bee88a8b4d37e8b855e4b683c324153aa3c83d959
z262a636cb48fd39eeee8ddedc318efcc0964e359f0478f94ecd9edd9daeb24edf1dd022b70fb3e
z987e8c88f6295b4c69fbc9e15a168d4150f865a2bcc1ac95b4de6099cab2e2a9e780875f601ef5
zd3943b0591c68b07781ffe5112d7d98c9e095d949d5991c9004f0bedd7c3d6c507fc34cd26f9d9
z7979f781e90f6bdf88e92838d609a3f165760d46c427fb9523e1599da36bc92925ed197fad4b35
z46e4f21e01cb9971e10032b2d016499378f25f3c2ab03612318ad64f4702e3bc175944513e708f
z8edb1770988be21e1e20a44a0864d3f541f3269a4ac7dfb07c1503814c6cb5c987d224d3e4e91a
zaf2dc063413bcd7fce4247ec41b6adeab74481703392879b2fceac3cdedd2a1fe707a92ed4510f
z677a779dc46b5992797bf35b98460bac41c6a27ab6c00c349619744a2bbd20ee7c046695638dfe
z5081d69603d37f5e82669d6f46f15d39bbee1b66d708694e8d2910713cf7c58122dc529789efd9
z03dacb0e05192f6c84afad3bc2acf8f3f9e5af00e8886484bcb68541139baf08e2e0d1d7039511
zd3ddb1ba38978091ba82781e05864dc11ef00ddb96ab8ce76058a9eff345ac71938c42b5d68467
z19a4df870a976af5230543de898c7b634290eb87b0a9710ca6916c3601bbdb31a96c5530096ee9
z271a323a6fcddf9a9f98beb22fc586de06558801d51007b18918ad18b38e8b3dea7614dd07a428
z0af7f11feff33ad0c2c88c8b831b8aec490d4b65257f798652ed5ee3bde86930977b951b23f857
zc737cfa18f620994ba902d7837597648461577f415a52d1f3f015b42b5ae4fba222f73184b8bed
z89071cf866c7ddff1b628780983d3ea3e3796d828ff9a22caba9e5ec92cb29396c49bb075fb740
z8ec7dc626a40bb31ede570111a396cf7fe3e60dba76d449b0dcdf728d5e7ae9564c69d3bd4a13f
z824cfce2515217b23ea752a02bfa01860a1ddcde5d454fcd6f18088a7c8b59d2229e35436a9173
zfd6762501d2599d21d10586bc637864017c6b04b54ef2711e1ad0adb92d687b879563dc2c8ff6f
ze3839b7da3b896071e7754995e2b09ef8562ba635d0d8a6ec331b5242af31cddf39676a840fcec
z285c5a2ad29a3bbe299eb470984365025c8503569c09b1c5a8240fecb201bdc8ec511b18e9322f
zc46ca816daa8976ebdfce26aecd264bf2e2dbfda5e6092df93b25706b283c8c9134b64a3861552
ze5339f431512ffaafca5ab2cf428a455e1f172c5a8529db371aa064afd3aa63d448419ef93bdb1
z62106901a5e15f11665f08cf7571076eac639b65ef0dee83c2fc2b04957cd1087a806c57c943e0
z0704dd86337340281ff6b53ae7b278ba0a5d95983303a62e1092e9d5d956cbfa3a15c01338aa40
z9bc416aca0423d94f5e97f3c5a3933bd689e8b2a5d941650a20c63d99563c3151d233fc41d95b2
z6b394c81776e5ccc77ba52bfb39ab84e7b11c648d6a841d052687c5834bc6156642aa9fd80db79
zb7a700cbdc477fc973f1862f512d5c79a3eee625bdb7c770eb9f639b9ed972bba3b2c3a6cabdbe
z50914a4530a8f1f328478eba4aa251ab5938be343f330515b02161524f096ecb2e96a83a3479ea
z864d76da5e318131da857b62a3b804726721141a69b6e144a405b0d9eb297154af2a9817bc9ec7
zbaeb367490a9e25e72c85f77b8c8296be056150302551298e8ed4ceb07083e760ce3e24588119a
z769f6edb2a88d5a8dfc0509e6d6861e27bed33adc4d382c0c0652073dc894d79b8ad7038000b56
zec69fe121395eb968f85c9338b272baacdfb71b53207cdb227a12e22b3f06315e05a77e202d518
z262aefedf38a9faee8d0ec45e6a5d004127d469d3630c04fc8291d479bd05c818a79111b48b2c7
z8c2bddd1c4584128eb511bcc7371d0fcea90c08608296f7ef765d81add121a0991b6b20ec893f3
z52e39a31c4e982dd0d58d991582a64d3108b42bdf8d555edd9ef5925c3b82a8bd72a9d37cbccd2
zd115464b24e48232e4cd8123f6e108ea41f004d561cc027cd7120fc49a0ee6741b791e463c5a74
zc859ad375070eabb976fc4d843af70bb2d8c64893af927dcafd6bc8b0cd537e8cd6b56e5763ed7
z0aa230c4220e62d28642c59a0b1e1bd875ea1f2b773d2df40164ed3917de14720dfa19615ab2d1
z624efedb4da3f08f00c16729380d181bef3352598e3b6862664a43283fd71766051056a6a09b55
z347a6973d958bae294ef3df397ca7a1087f6a75d66f944110b063e68c638b5e76325de91181ef7
z393269250a90ea97f740355379b18ed107d3276569588ff7f01e1dd1eaa0d41924889a13eb1d0d
z68e7b2a4a97b936bb140685cf99889152be37be7bfeda09368fac2c57f1c06930de5acbe3ad9b2
za39dcf8e285cd320bdf2a9856745fcf4406314b259b43916d890bd5d5f1cb9a39cc9d5a097ceef
z7895877f5043a27eb525cf238c61c88c20eabfe9597cfc5aa433feac14b363298c49d841415ce4
z1ecf2073a39bb6496925c884e9b27937b9d8059ecd44865c428d44e59eb3984da3d256f2a804ca
z9f52d1738071bab5d8250beef286c2101e4335edff8a061736e0be4c5f06fd000844f1be55b61b
z429171fe6f8574a75a46dab67a667a8d885cf8b87e23ad0f3847b61262ba81c3f6ce2c1fc2a195
zbc50a547ace22368e08944800d3f5d52597bfa8bef6410a34d3b254cfc78f25cf91366055e511e
zae5e2483b8cd26b0189a65e70084b3a9cae24884148dc17e59e366e40ada42c8b017f0e12a5380
ze7eafb20d3f029815dc2afe69cc123f7872500839032a7033172e4ffe4656209a841a90dbc85e5
zc729e4eef6448534dd4b82b975f845b943872ae684121bc042492086ae20491e27222bdd34f638
z1cce7c9f95f955776fc40394638fc8b46319f6d324c889dd57f0949527c7925bdf62f95b71ae56
z8d70d778181573840b94a2ed1cea219d7849e859039cf5dd80a4bb1ac0dc68d1ff0ec121346fcc
za8d20d8ee87d33194cbea058d73454b684f0f8e56f31d60f87edfbf0e76e434b5f53f7dafca8ce
z8cc526c0558d7943054206af88272538fa3268a62e6be9cdd4a0b1cde86412b0269ffe181d25b3
ze223fd091734e116d37cb335bc05f59c746a873e710fe42da09de8ae848f0c95e447d9ad7ea6a8
za7af58286dfa0cdf0e5ca3398741e21aa71ef3adf4dd6c7b1a5b63b1bd3f891bddb5e5f954c683
z228f0b81a5d0ded510e5b264684963969645d209977809908c9b5bf6e67d26d57140d344ee266a
zcfeebac4b4bc70971599ddf81cd4ca31e87f9b558994b34083672e27178d2288a4d2c1f404f824
ze93c8e880329c9ff313c0046431abf7970321e032292e8a7f760d4b419fbebe1051bfd427796dc
ze5344878479c588a40918bc7bcccba7b505786e1d74f5bbaee6c7ccc61b78b90dede79d710ea7c
zd94bf07113761a7e1a54ddc18e9d47a36334f87f6f5b20a62a9fcbf0afae234c7ca6eb55d8feb5
zdf6dd62abd661e44d90007a5a8b08282e765164fa514443a129edd6424a6a5486d2bf14bf5c61c
zd8f4a11dd28806752fa8d61d0b4fc32d527486d0380c57dc567b8b67338176743f963f2fbed414
zd5e740f88de12409c770309c46079fb8d56a7705d9d21c39d7b9ce6b0a09eaefd909f95ca5f2f3
z489465e2bfc2a48247dc8ba5770acebf9acbf8485ab2671eca596c5aa1bec3f1fa3821b92f5ac0
zec4d9a9300d94b1e6508c2dece6f03b288158e7648d5c92fcaea3bc7550eb295c04d7d97ffa239
z38f82fd57a2390f7b6ca3b22403e086f1f3ee9cee4af3ce752e1e590a0258d8fd330356bfc0af8
z4a45fd69216cc182a0965906f35c6ee67fc027877c57d63c76bc6e9257d3097fe88a7b0579796e
z3957acd813168376f9a28179057aae2070959bccfaad6cb52c6b5d67ed0e572895c120c84c690b
zbb653e210edb14cd34b4da2335bd574e5923db013d3b0877fbb9d74fd73b46e03324cf63edb6b9
z3d8696ef1c6b58347ada8cf661e197fa96635ddd1df185984353169be7a496585860dc9a94d3c3
zadba952c36d2ac30e9fb0098226a70a6cab205d57e0858b4d97bcb11b4f9028fa494310f6e8364
z5470bfb8dffe9205a93bb16f412883600da9b2832e78e7797e70da54bfea6baeaea6b5634633bf
z782de1bbce73bd9e62d31f7e1d99eefa0a62b5b8d5d44e7e1491547b8f7558cff109d69bf5915b
z4c64b49f7ca46332e8917bd54f55d725d325c52093d788fdcdf8924d129ba95c9f6200b2beb572
z7bd1c6520a37b20c8ec300420d2faf5f37c2c09171f6b4a16d0d491954ab9b00d962d39a187f2a
z99fec8cfd4e29aa379f9ce13ea893eabefb76eba5db6b41b0e3c06c9e7af711a7758e088d3535e
z9e1d6d57d1b46b995c8d557f63fc4269da4fa6b43aca87f889fbea08f8b8ae4fce730d3f7d91de
z3f4f799283ca76caf4a3eb71e669f9ba12317dc61c9519b1230fb21f66d122b789dd85ec895ed2
zf890957f972e2f2d8a66577a07c3f8e17e653017aab8ad53aab7b2cd631f7ee4e20ac66bcfb9f5
zf801c16a468da352cc526f1dd7d74e01e7a7f582c9de930dc44d4c4de3d0716586449fedbcd6ac
z0b831c7a6b5b384827d9241fa5cabeb97289cc92de39a380b8c714e2bdb39cdfa3768300df4a5a
zda225102819e078ab12fc9a85fae6d1c54ce0c4b157f21f01893bc14c5bb9c935d02eb19aea37a
z373c3a6ce7901354ea22d7763a0f5ce4ea9ea4711d086148d5709bc07dc437e1fbffa57e3f9a97
z4946d984f1c8f1328375d1357b72b62c55cc11b7619cd45d3fc347b42836ba6b897a67812c0737
zf438db713dc010e0ad0851476a227ef510483f138e21064c87379d4cca126116ad5acf18467182
zbb25ab62fe04fd2f6af9b296cff950371b3e9812a875b9b5c3404e471dea8faaf7ed440fbd40f8
z8c1f37bef3b80e9412bb3fef0ce4a7887dfcb604e4bf41b8f6dc8051922719285236ca1c6dbf90
z4705d50318f6b6f2162e8ea428a09b75550082be0e3403c5ebb087613f0a7fe03da13b3bfa7b6d
z314041ab22fd05a50718ec550be89ce6e9dcbd4551a6a612a02fc98882e9e4203a0628b7d80758
zab2b5d03e8916bd651223f279c6e65cc862a6b3d9af9d68ca15ca352dbb9557aedfedbcb204390
z1a7aee985ff4c0222e225ff33b0f1358eee7c486d4f840cb6e8251ccde22bc74b8b99611982b8a
z457172af841c66cc3275b6e0c07c5f3bcf61b3b997f0350a715189cb33066e52af8a3b0cf64242
zfa8c08ed041be951218d6d99de47ec0525e075ea21dc56fe199423d2e167cfe0f81352f99701f5
z2f2e37204e593960f3da1857a2c1e3e41c6ad1588bace60cb9afd339bd1d0bd0cfefe88c1d7ce7
z9d1599639e144a617ddd284473cec780de08523040adb1c839fde3598a44a629f26ae9755e9c2b
z9e636ab5d8fd0342628b195b00152f69192fcf8c6d3344289240ba1a127dc64a323eb2827a07c1
z1249669d7eaa0066a5be88ed4eca9a6cac74aa51a43ef7ab97950d822ece1dfe2ee78d75542cda
z3f614e6a2f91b2ad398d9f0ec44c4c7edf479761af3731586188516c26d96de4697697e63259ad
zd5a6dec7d9a9eefc290fbee3556fac0064bf15a6040e13dc258201fa89799cb1726ea630dac83c
z078f4e79aec3a9ec55307df64f9a0005b62f6365bbdb49a3a26fe6d9c38dafb2eea2f1e8ec3247
zeab3862d94c1d17a8e2631b11a8eb08c60646953f9119862efac2aa405964e818ce66e7796e154
z65c97d435e1cb46d5b9e5508046d0218d2fe9dd10e17fdda1cef05f8bb554da9c06fa6d908579d
zdd66aa7bb20c665f60c3a5a0d418495ef95511ac1dff66e1f2dd6c19298e6d0e0e97daf2cb0f9b
z24e45fe85a2e66bceb3079983fdf064a8314e99092aca18faf7b6f605062bf1387ba766fcd3345
z52808507951148008f4c4c764c9a4a44365236c374278e24d7f303bdb057badd3a29187561b805
z2b52af3287ed954374e2e8e033e20c8a08453ce09b00df04ebf4904a3d486e12105c240a20f342
z353802ce4e526cfd0c9f61307495eb720ef2320554e306f66e160335945ef5d1136612fee00fd5
z436029dbb2df5f0c8569dd3fdb6e0939f6a663d22c1dba4a62db3284f1488bacecd23fc040dd0e
z96cb732d1da449b62ad09be89b2f176a9ca5e33c6c01a0e22e0cbcd8b7faa43627089c2de551fe
ze4ab553230323fb411d6f6d3f1ea774f872d94bacd131ba0e996c80720f9280f5191088bfc75b7
zc3c587cd4fe15652b6f905995a5c49a63567bbff55fb75c935c6f116dc27eaec67710e4cb64df1
zc3eb87823724f7f187e4bd7891392d882a31d878f31ecbdf1a7c469028253e7f108e4ee9fe578a
z08d632c629cd5af20ed6da59f8e6914b7932b448a3d7b40d8546031e041ef8dcb8c24a6b526a94
ze0088d42ea4066e6874199d00a21b6d4758d0df8780d0c2212bb1cc14ee1dda0e59b987bf66309
z319fc3f9d233819409ff738751ccbe6d8c01aebdcf491ac84efd890677ebb46cac88cd969c401d
z0d85148ad6cab742236971ffed9f04a67ce35257f21daba86149eccfacb4b61630f67d2bab88ae
z69e63c1b9be9fe61cb47b6e187cb2a38a7cca43833d0a9b9855d50f69d52498d2b273366f14fc7
z0379bfa18a102d3b3b0c80b6616a4dc109bd88dc93b4749b19db0e45340c4d94dd92f36d40d0e9
zcf9ee941e8bc2876f1c349ebae94e9f046d4f96a9d64a3a66f90d864903d02dd6ac11475cc50d2
z118dec6ab9ffc058baee918fd08e42a202e9f434f8fdb43f79d5bed895f0041ffaebaf27b406d9
z9378770820ac9a633f0376d60c75edac53dd60392b07167cc50090fbf89d528cc6df4ae170788e
z992763af8d80532565edd1c7d25351a459d41ca00f56a9de17f5b1d1117dff6be1a19ea879253f
z46ca21a77063058c95b2dea0b60c03a37b90886337fee1a2a4df3cb8a19bd4f65164ad6594dcb9
z672e2b4764165a1eae3f23d4501055af615c3f51038926581a0a33ced052d38eb2dca9681e009c
z517d20c8b47914b6f609c768d21ea74794efdcc8661305170a214423f4e8b6ea25560c1a7d3e73
z9abf9556ac79dc6f00278e8bb36a3679c2e1b319806039be100c6293bcf5fb673ed280acf4eeb3
z827ccea0363f47c75ed95c0f37baf9edbdcfecde615ee3aec5edd1c4f2fadb9b32b57526db82e2
z4dbc5062f4580be3c3ff6831390c50cf298bab38e7865ec0876bc55e91ea3664801e2a69dcffd5
ze711545e76c82a2aba2106d7ff3443952e032d8375ca857704ae17c349ac7bbc5db7ff81541dbe
z9b98c95953226b0bedc70c49246324d57424dc8cf9dbc81effd362b9b54c6cf9b29e2547da3cd3
zb439f1fb613e0d16086241490870c14ac46d290ea1212869dc45190ca3b2d64f3c3b6ee735c727
zed7e869b6e3e52b5be38adbc86ba289f1c845f8bd4919846d7f03b0cd7de3c700fd3a010e44306
zfa2b331463dc89c371c0377fb211ef726a7e488e55a5e4fb5d62abe344ab1adc0a9fc7096cb86e
zaadd988f7fb0737f65941a678547885374840913f597e1c59751f3ef1d1d306332dcb938a41b44
z89a8ebb6a0b5315af3ca9b072c44f4416d02cc17a7fff0961daa8e30b0acfe877586c5be769011
zbaacf8c8c49613b8eb822618198595cbcd9557f4d797421997a33273f9fbceab80193f4f75ee00
za94ab45891630fb0b753b9dce6deb268014736a3bac4c0938964e134a378bce0f6f22b6d2c0284
z1eee4cc06fc9803e836ae69056f2eed5b1a059921a99ca739635edd9a224a1d442e02669290713
z626c8510321479e75fde92ab8134cb0046f5907b9ab02bfcdf1310793c98630cadc1fe7bc11c20
zf6afd2757fbb367672e85b6d42df0605e355964cfaee75447bb69acd7ab5dca6581b8f16e06e67
z6c8e485f37f69787f1318c3993587a6bcbab73d0ba6fcfdba62168600c55b228bb8534975766d5
zea8429c0c1a7144436dba8070e0bd1aa2642011b6f9018c8805ff821c7a5b827eee73fa755d37a
zc2e07135c7eaaaa1f4413a62442a55bc18363a7c34b4c0914a2a1440347e74e57f06bb6596d599
z50dd71967e65624561677b9443177ce4115ca16aab88a8616457db7210ac4141c4d433485cfba4
z70d00aceb228f7f061e2aa5f870a973ecfa9ff91e4113d0c7bac39c356e278f0f9d753eccc6262
zfc759bde565e79247f03f129f1c1ae2a65c9e01d7866a395ccad0dfb5b41ab34263673e0114c2d
zb04d4098190a0e1c755811daca133caa981e9fa1915dfa58cc00390a0ae37758be8da672212f68
z51137a4388061c428955e0bcad4a6c01981ef1664d70bed9f0ee0aa963fc577163628b822445c5
zb4da9f9319e4fc565696cc299c6e4eb54f1dc693e5ed4fcec5b97e53f7a0984b725fc45e5c30de
z0443758d8b2fa178b8da1ffaebb8cb44b2e22efac45092ac985f99a9dbf1b8186c96b69a661b0e
zddef1d4385f6e29759f57fc21d249c01abdd82c2ffaf2e3da3a3bb0c979acaf1ac5bdb549189c8
z6dbc145cc9ccad35eb6fa9145cb537f659487ccfc70a789d75b3615c00b534a6176507568ca315
z188254cf5629af2fb3a4186912d76ea93a73c447a0dc2f9d87ec4fbc50c380473411653327e241
zd8a24b3371ec055ab96033e2160210237ac3e2b6cd77bd4b187120edc165f8b524f0d721406730
z97ab2b9ad11242c5e77e3b76bbc59b3a96124beac9eed370338f0ef2e7e3bfc4ebae59a0da9a88
zd1b5a444609239a6ff2fbb190891c3d560493a8103ed0bbf56618cc80b11e258cf74ec56f73cf6
z6d230f016aabeea240c4840234e66890366c868154239b2927c357c5876ea00470b236c7a06aa4
zf08f457aa0075ec3828599836e004609d3f4d37a7db75eefdc43de2e61b8005fda56d693d279d9
z9d4d7d08ecc2c63a1c9949907716cf999d7393e0d405e3e60042eaa9fe0906630b05e7074171bd
z0eec294c7703c909e7f55c3e0cd7c478aa7adc4569f59f85108da118d6618bea142c430a3c9bc9
z1305ecacc9c5f684ac7e91334e0737e1df828608d968541bed8013f582df890004d6ea92b97437
z3e37d4e58503a3a43dae441c4fcbd58417fc22d2c61b90507d2f705b6a0d23f3d9df5070794761
z254a8528a9e6c91af2d70b27b3bb524a8534d2dffd6a3d9cdf437fca88b454d9028409b2821078
z63dcd0dd7af669dffca6dd42e33d3a0845c035d61578ca48c165dd7feb65f23d838ecd2e3bb663
zaff9a0071995643ff8f7050e41f4b6ca8fc4208c7c71e486dab2cebcac9575bd7d8b27ab53a68a
zd5411b2f2b9c6c429e94628cab0fcf2246b3e8506bae683b71e4d97cb3615ed8cdc95f3fd2d6c2
zc091bafccd839b17751ae27545e279730388dfaebc2913f11b74f606df3d8945ba71ac66a4183d
z87cae4e0282106695e7fcd9285987e8372792b365894764b0cc18288b8c9e388926042547e4f96
zc61c8542c1cc38549306041439da262b0868816e10dbdd84005eb7fa2389deee92d1cfda76ceac
z7f7ace8e14bfad54c0219e8a65ff6892bdfbf8b1529950e81fc6d2932f607367e6e035b7efb922
zc9601b0f26aeb407dbb354589806865c4ca80f8c46277237081498c38e12c8476ae046ebe0c5c5
ze274d01ae7af1513f51c7a99aa0d5a45b09a6c11a7da2088e1a1624efdb2201cb06ad296a3f2c3
zf76fee42e8a3b78b6e727149f9fe76aa95bf03846041dba7d92106c7b1e5c8b4f8567b69520adf
zb2231c5868b36ed25d66095bc69194df2e227bbd54a7e2f2246f43ffb4d5e405927f495c8c519c
zad2c53992e10aba40df7e2798c79aaf9abb041b596094ada18380ac4b81639f87d164cb5936d96
zde47ac22c3bbdcbda2724249954cf2a871c042b0ad2c01c65cb99bcbf90bec7e18765ca3f46ba0
zf0d815ce6417673c0d0868fa0bf59ba1576b5e001ebc1dce5e4d42255e98d2f23eee9ce1729e85
z559698327de908438f09923d522cbbaca17e79354c7d06bd3bb37f853f22dd5972457b99b52477
zda6c04d7e07748e221acb39fd8f32f0832facc9767138133c4e65ac652724c533a368ef5a9fb96
z73998d5e782fdfc272dc7d7d577fe2204211e10af5730ad63ba082634f03666b83085a7af96156
z0d0a958c2c3be7f8e8af6b566c9b4cc74cf87bc8a74ef4727cff8539f0f57be64a36d98f44c370
z9942c461e583c71057ccf01ea70eeb59939400021e2a54be45de99157d5fd0af24ed38890e10fe
z8ff1caef3bec9419811bb42b269f529c3da53fd8fcdee1a9eb457302c55a5460a7dfc7bbfe249a
z21e5b79055becc2b862a5526760bdf0f0a02e5638e0c859af63e8f341dd5cb52be80fc8d4cb3e2
za3df2a81d6767f7fca403c83935f9421599cc1e75a57a8bbb296aa492bdc57769b99c296dd3087
z2aca54cbbe86f41c10f996c28fdf1a0bd811c86618d91f428cc4b9bc1f460c69702ab71d790899
z45f2a7e4ff5cda861c35277f2f955fdb7ef62254f92c050c9bd6bc7c22ecaaeda8f011604b5d80
ze23e88d57083c50768e72dfddaa3abcf60c421a4d9c9340827349deabadd1df39e226f5200a293
z1faf01d08f99ebe1560d3fa9c61bf5791c7755d567e11655feb8019503b3087d4f758bbcedd1fa
z1f430982abe4fbc35325258a613b4ac0608547880b9e11e6a538cd9c469219e2b4b16edc145bdc
z771423c490a32d92698f5c403cae43abff4e9864e4114a29a5989c62869fe3eab511eff7fe9856
z203b3340bb7e2797baf5fdc2ffa608798d186271d3dc316d03cfa2fd7c7b6bf8613463f494599e
zab909fd6fc98bd040ae7dddcda91968e53742da976f46e6b300ebf7acc4de03f90ffcdc3cad7de
z363e8a8e134e17fdf74dedcd417e22fe9be455369454ad0eec8995b49ab448529becfeecf3c5dd
zafcdfbc3a5bd247126ebf247ccf4d627444624b7ce20c618e677096e36e71367a572f6a1ff482f
zeef8083f61c934da9605470ae018eb099d20d32a18db6bd4d5410268986b60aed99c5a414bbf6c
z293f65851bd60bf2487fd0c8a3e3277fa4d7013520734d3a83dd2bd3c0109aba81bb9364b83218
z35ae6b8c180853b63b14ca9485dc4c4734a34a60d15013dcccb2fc62fbf6072f2fb95eb761c002
z078eee9cc5875c0fac9e5bfa8fa6b7cc988f9ae78a98907522ad99a1d845930c5a0309502af8cc
ze9f01160e804429cd5f0d3f3e408a5f08f639a4ebbd1ef2ccd83968b962248e2053e984b1d4294
z9b4099a61a3bd2e472caa7f20158e7ff5dfd2e1958556d17cebca7d044c7160312d2f186828319
z198ec188546127a062d544ffb585298fe8bb060d14793a8f4adabd20d97018a1f544fd3c3cfca8
z3228ae9047f214c11d936c6a409ed19c45c64f1d27605bf44630b77297b5fdbaf175f0427e31a8
zdef9e8f7ef6997d05c30541e23a79f4675f9e21dcdd373afa215bc0225cf6b97cae1c6358e4b1a
zf97636197774a3cde5e1160d49b3ca7b38c4534347863ce1a23dec1966f6daa0eb7b429cbb3a37
zd04d1afd1f68c1a0ebd589213c4279cc8417203422a77e3f36ceb246fd929b95567842c970e69a
zfc5218855b8b5528fd4888a3aa62703134db969d9daa439114d1154fb599deb747007b5ce9e151
z6adde8f44fd5d996b89e3bcfeabb412e4759dab093313ba33c1bdb4fcd8e0fd55fb2c751b168f0
z01262160f159887ef38ada0bf138667f5996b380b093b09792b514c29be2bbebb205a83ba255bd
z409f2fad5fe3296e7010f37a5a981ad96ae0164aec823e55a310947b442fb07308f8422f33a6fc
zff9a7d423d9daee3c5ad83badb5e92d8f31f31d05bd01992cf35c68a8a238813222f7decd639a9
zda889aee92531deb48a9e3662d66f8cdd3112d52becb32e32c228794e4a233b372b98c7a0341c8
z8490c48ba237a82acd917ac1d20bb0e7210bf40a3954fafca2dc8625d0a4a69c8cf43164c560c6
z5f56d7322d92db1514fba1df530ca3e654e09db7689ddeb277939fae41719e08989f74c5f3764a
za754245d8226845785e72d23342960b9e8b8384d9b06bc96a5a8b3f40999355c8af30dd66452ed
zb70174749578ad2d4028e3c68f868d065996ad2c4e3a08e3725495b9512f7b8018527e3e354735
z464e5a786c1b5a39f23df350e852f661813d659551e11c17f0a899614cfefb26fe1f2fc04d6dfe
z31cfde627d881a7fac54d36222394f549fd9e3bfce727cbd3eee47f7d327cbd6540069cdc81953
zd704d6db16cd21e0936c755840d04879bd585d31bc55c63a95255f36bd3ca9c3eb07095201ed43
zbf042882827d45c425c8732a723e725b4d4cc930bb0d59e82df26c230b8fbb87beb1b9a6de7555
zd82c1e3d5ab76ea23f26e0807896bd73f73e1917ca8f7b91cad6a6f32255efb91bf39c0b51ce20
z7eee30e020aa282b62ba9f1079abe80cd1a64fdb5dd239bcff876bde21b956125e11bdc10a0534
zf9d6c06ef71fcb52ecc4a128b309e1430010a3c7c85ca0927b6a0460b04f248227d520dd14242c
zd568d65f93b425727fc0a33f8e2e443829578db6174b5febba11c3c6dd35fe515bc97cbe8e6954
zc311e86d20a537d5885824b41b269297594e8b61142dd7e7c4ac768f49e163a488e0ed29a1e279
z0ae4806feb77a8d1c7a8714b653d2155e1a8d7c14bc687ca2d2daaf49f2b8c6649ecc7764fe588
zecf26bad50dd91dd5be10e7d0a993bd99cca71e0ce199626b1c1e271a60d5f1cc4a18244acf8e1
ze6e4bff8f06b263d61c07c7087c54c06113539b41ac7f36aea12dfa0ceec20d7b275b4834c6f77
zace43cc6f3c4953bccc914d44d3eb8647df8b7b0fcfc4d5cfc5ed274d837e4c8bbb62b92e4b9b0
za47e30f48926877084ac71fd587e974ca10225a3c5058cc79b0b2062795e6ec96a5651cc30c79f
z7f48d29fe565c51c4a3fcde596a8a5296f796e12b30a678c936730fef8306f9a1cc0d2ed44a14d
z01f39f3ad9a40c66f012b815814149449808e439adfe36c1838fce125dc90ba90ccdbc03797b52
z4c57345f19d0ed7d69360e21a638e58cdcf6e5af3c60031482db5939b766c9ccaababbbb16be48
zc9f2229f49acfa1052060c087ba5e709c33d521f0586d53c6e2bcf555862f45c7e03ab5a0e388b
z7ee3d4a4f3369f82532d6baa6c4b93d5c0039f33a9c1965122f0225674e6ec4e2cc867b6db1fb3
zb56281f1031ecb1c1dc8a8a21cdcbef888a16af5e2354e1e8733a6599816d9335bcbfbd0356032
z75c990262202c40a30bcb52b428bb49e67c64caf5af43838dbc99ea3cf977dfa96c8782da03b58
z3ff372eda8d1983fcf442052bae8ec5a1dca3ddcedc242f8c19ea84795da309dcf4bffdb32a2cf
z3ed22881bfdf8f94f4e4350f4bb6d4a1293aeb424b352e78602155b30bdd89c5de8c632a0916cf
zaaf32753a7db4fc6335f7de826d627e99fa4cabfe2e4966aa97e2ded8bf2b3309513c8bb5fa9db
z5f461e56ab407fecf1ea7419f5a12cd64ac0c4620f481d3ea9fe427a0aab51edb91452fdfca1ed
z401d0f73e2da42664889cacf1878d888a051b7b2b5ff43ab96a8987f2e5506d0901ba56f6f6cca
zb3326f4dea90637acae3b997cc280f27444ff7c2f1902208f3854202f55df3fabfa7b216bfba2c
zfa1449792fbf4aac0a670480361471c58562db34960cfb71640d0f75eecdcb2b796ce849404877
z10edef2a7bc5e951c0403114f9370ca7a11386c19d6056482d2f3cb8b05560c2e8aa1dd010984c
z52577cb1110ba7b62f50a63afd5268cf40122b1695f89b52a1448e5c8c300bacc735340bc13541
z839d6ee81804d202cfbd1752569300bdccb47a07fa0ecc48eada5ce5aab56eaf127fb6d6548695
z8b6bf434f117a0e41fa0bd478e07a60909108907af5bb49c978b159a10558a3fe945a031abf4fb
z754ad739bd5270fdfca1d64c2abe3e880f4931c8f500c21dc5b2d1cf2e6e10484a07d4581c1cc0
z543e00243ff90b70239c5cfebdd0b19ba095adf3a5b8fc4588dc4106b72e4ca7aacc56296ec9c4
zba52e07c08f37afaf8822bd457986e1468d811f1f0b4590a8a9f3f319aff761673a47a4a23e9f0
z5696a0860c71a972f9ef7339c5b8111ee3c4345082a47156684f6a6977190492ce39d9cfb6e3ec
zf42607e0a1561c5bd6a529e20cbefd4b47096cdb1ba4409f6d9c058421d9985e6d56be93ff9219
z6f4e0880755b4b99135f67eb05288ee89882fafbf04827fef5d3b8ef2ced7ea30bdd70521f17b2
z501f93cbabcbd2cf99ac390cc8c536671feb097f84be1c26e235da195ebe0578302e4664d5d80b
z18241e1e0bf83fecb0398ec393210b5ca41360b48aa02618b6f593cb325c4b09ab7cf97e65e610
z0a3adfeb311f0e711a3b79424d23dc56ab519653dd982ff1ae7cb28fb4bf03030cb46e929aadcd
z9b8312886c90db0d9261df8d336688e355cb30f63684977b775a3842979208c77ee55536ed4d35
z22a8c4256d1cfaea51755d89605f27663e910ad5b742d3b3cbb6f384dfeb0d8aa2804dfb25a277
zd8c0d0921e9e154b920f58a18fb0bd22df60b1182bdc2ea43218936e3c9af0d7ee29cc44cd5169
z85626951b07fe1fe90b6239a6c78d8bff880555343f09ad11fd7327238b7dcede7e1a14d4fd4c3
z8f86ccfda708eb3bec349da5c1f2c224230e068f5237520c9987262594aa6ebda71b5fa57e1fad
z69acc5b52dee4653ff75f8241fe59f6c237003badf4da7204982c94513127e172587e7ea2cb253
zeb8abcea22327cbeceb410afd22c0e9770a25e8f044dcded42284f0efdf6420a29fcaec48a5318
zbab722b1757b0497bbf0bf0fdf87e770453c229f30f244ffb0b1b9f616e2ce63c3e565331eb459
z6bcd8546d08e3c3b705a1981a6a99de2a2f598d701eef2c8ca6daf9a8897edcf86e1fff27f410f
z378afa049a45b27b7626e44e604b83f45f2db7fec3fa9244a836592f31db7f48d2e53b3ad4f2c8
z9952e9f00ffcf6ea82427eb56a2aa375309402f57463520f4fce6faf5d8aaa994634d35a37390b
z26ea9791b22ee554540586fc3261db091ec415602eb4488f17b8cbab8b28c153461ad392bc9fd9
zad5b467d0fe0a56e494b1cc8ffc6a61725a3d99af2b42d09491f37bd50d387bd3a5b936ba44b21
zb99b6e66fe6ba35be565bb936e61d28d7ce2b9f326a1d83db207f37558a0967c1fefe22928b780
z8afc69a18781e7cce375ffc3c7c5da4ca28e95d5c4605cbae63d469f28deb6344d4e71f72956fc
z1144e946a71f494ae62affc661479d416f73870336ee28a206dcf7e2a3a490b2be42d8cc61244d
z2a1637c76b6ffc84ed84a117ed7eb5643b6c31e0882e41ef28674439d40ae0b6391aa9cb0ed959
zaedfa6afd646c46e2e5d01370a0a543cd4ed59eb43e3de43155c875499e8563fa5924e12ec4d72
z64d051fc83ac11057d506713b4c624d2f663c42f27495e5546a8a598f704962e246a766eec7cb6
z17471267968ee429c894fe7c42ad00c8addcc42dcddb8e672f1e7cfe5d6b3daa56831898420115
z886db406d0576a22ad4e7c70a74040b99b5e9c1489951713a7da4880026081582ef3375c605d53
ze42e35e78bc8ffe63a4a6927ba5181f77167180b32e4fccaf3b65ed7ee11b2126ea34a31314ad2
z8c99b9fe9d733a16e051a0579f9122fb817c767f6ade9f8e21464a159efcf745649e5435c90359
z31049be3a0e5a5176121969dd9c900aab0e47ab6506fa509a7aee7f049c3fb3bd1e2564ddc87bb
z14273782386e683c5aaef53cb32524601da4da7d5583c51cf7d6e2b688dc12d76b1968db98f315
z88b5ac804700c6124689a60988c9a7dd1892466c130656159435e374e9dfa74e936cddae4a9b63
za3a1fb919ca4b22f69540cc90e05414fd60849bb8c01e1cd22b06e57445ed45072d38b0d4a5fe6
zb9fad3f0e90818dec50be8d047f40ea735a42e1aa56fa4fb9811ca9efcf7c08346b9d64feacbc6
z62bc02043a3ea273bfe94bd1d6146e04ad3fe4b3349af61b893245f7c150392ffe120934bd039f
z34b1099847dcf2d4d64144179cc2fbcf44ece65473acd2ee300abe50b306ab39289890efd89128
zfc32e33066e2d85fe6138c06c69e13cb4fb0d20268141d3d2a0621d0edff7c42d6ffc0ffb1a58f
z0369ec6c754f4da8d94001dfa97a496bc189ec8d1c0de7bfe1967b20662db8fe4fabbca18e19dd
z0d685b6524717ab2810951e18c468afc171e416ecd6011382caea466e62db895fc9fa5dbff09b9
z672ca22eb7f623ed959245615d9b8a9b56b0a083138da1abce8b78481ff5fdd99d3ce2b9425a83
z8f780c4cf52a339f1aa68c5d45a434ed6b2cb50d6655a44700a6a26e17dbacaa5fe9c506a40f94
z3fe796343089ce5f50ae97cbd5a199ec5f0dda03861ca5709b1571b87d8aa076425671145229b1
z63af7b5cb11975d559371945d0bba7d5d7ae3896289ddfedad0aa4c638db7c85b7e15f5c5716ec
zbf8ce94e0efdcbbfd2cd9a15fb160c9d8dd3bd45c42bae75f126cc67a9ca424bb412c343ff8aab
z913fc0a5916a7eaa887d033a28aba0f086e70766750397124f23371c639f03986ec4f8a0332808
z7da57aef7856b8f135c1c6757327d61edeab6aebd9b15baf45a406d89a951bc1f6b92b53f2ee9a
zc97e5191caf77feee043c66ed55c5bb9cdce05acb319fa375a58bc67b85b58cbb0bed260885b2e
zd717bb74ecfd91de8abdbe1ea9e50f699963011cd9eba36d001e0f9ff047860fac2f6d0ead3b56
z21bbcd4aa9c9b202df850b5df03e720b12bd043c451c908e033ffa765136fe264f99775ebd3701
zaf094250cf78867b4d194921b4ac732d17398a3e773bb78d1c3ac4a1871c53876e2897b33fc336
z9aa1736504036dd69299ef468e6bb5b9a45e7575e7dfebc1fa31f549567af92c3f273f9feb2915
z3ac87ff1cdf6250fff75604bfb28a492150b8ee40041451326e180b39c4c82a77e14407e10e765
zb0cba5299b90ebc24d0ccc5a973ca5ebfc1f5107ef8c6c7fa7a0f8d1542c6b910d95a3bf033ddb
z7fb2b9c96109234c98c8a447b6b18daf0c0630390cd9ebdbecf95a6395be519dd4c55c295897bf
zb815f3b2eba95c1c386816e98fd78b8910bfaf64e6a819dc093247289577e581a25b06b0222bc4
z6bc7c6572178ce56927f55eef397e4a0a0dc7cac047fb37c6489417ed630f2fbda44e459a0b98a
zdb8a81ba01ed7be166e2bdee17d7d98cfd22ae20b8a9ab4259ce2c60033a381717d402e67dc17d
z4b926d69dcdb413332edb8a1685de8c4ba1861c6938b7b292ea8165a913393f3f89cd4785ac4da
z201d7ec0145174e6d6d46578fcf8a8f09b384e868db81cee2622e8dfd230cbacafbb8df92d8f2e
zf9b1563f3bb78829173deaa65d1598b15cf7756ec1fcef82003f8f13dc5c9623f23ef2e2602456
za061d5f1096626e94bbdffbb637f535e29b5cea5cfb706d75dcdafd6bcb0084fb4443cb3ad14d8
z868d98b84b25a20e0a9adeb0aa352ec3a147387ac99a11dd2b3580e621618ce7aaf761e7f28c6b
z97d172bda97884bb8a318faf42305a2f25406c7bc9944d4df42b422cdd77ace0a41db4646d2c28
z6e03aa4423c2c0851ffe4204631a1aec6c5aec2d3741aff9a0bd7efc4a6703bf5f89c0852d0fa6
z10665be6759e215f3540fcb6a13d241fc9b38d245af2cf03500bd4cbb2ce3923c70724da92ca06
zfcd998a2c4df138150408672f7bdb1c4f6133d3a807c744452720b0372213accda57c55671395f
zb58bbbfebc3b7205c2f908661a74ccfccc2fc1f730887daa3c9b640a51c2eda444d7bd3abb35dd
z9de3e6477474e9eed2482411a34b937dadf31a4121316a9424129e5f14f08563ab211e9ad025b2
z5a7242ba952fbc5d767189222723b8a7f02329d5e5494b2f9a1b3e98b8a0d05158780e9f6c8c8a
zf146b5959041e04a57b187e411cb7debc151cec70fea23477faa6eaebedc819d69bab3b2a34a52
z63199bf5a37de121b3cc7e69edb31a74b2640a518e827f5d80eb4521c38af0dabf3ecec079706e
z09048d84edd500e37626cf2297e2ea073a2452f5c1d38e83a33875d8b74eb904a79803ec9d35d6
z14fa7e5fb79dea85ad0ab76a2cca74d08ab7a8cb1741518f4b04cd2adf5f0fabce074a7cd597bc
zaef02fea92f54ba78f8522bdb2627619a801453f1268af7a25d73142bb1148cbf0cfe74425b0cb
z767be8df0d662cee2fbda90bcfd754f3eb3c5b9a168f93e34feb41bc7af4ba402e917d74b09aa7
za6a2fadd35fd35bce5f3ebc1ea4935e82ddf144cd86e76b6112e317f4ab07e54e3a96c9ab48b9f
ze5dfa1e9c51bc151e1abf2b317b3335b9c42b63f44948f84c0d503328dfb24a81cd108ce885cd6
z9ff9115b26d3969fc315aac65aa7713060e22449f5964afad1f1bba864d360ba50ffbf87df7e53
zab33b252d8e7546211a52adf3044edf547d54d19727806c7ee773c31bd09a4412c06341b5a602e
z6d26f6db36aa39f4bb2c2a38b1013e30fb3c3a1b95808e4b444939265a9355502932dc8040217b
zd2a6934b15b3f7c9e4be6bfc2240c9bf72a23293fd1796518f5a190920bb11652f908e8b1ab90c
z0137ac65de3741630d9252904f5d8a2b80cabb6048f3c16d64ee161bd3668432a5227cdbd1bc75
z8bfc43e9316bb873ae02a5700e06708865b5a66ab6f4889d1f17f59da88a6eee8e2df2b1222ea6
z3a8b427ad9ba08c58d8ab70661d180a09dd197a87f8344ce99233b0546c874d532a28da67854e2
z319cee7d87eed441b60bd8ea108ace0b072807bff1c14222249bf1c127413e5f342c2e9e9f27eb
z5d01bb87a99a15d15ec130ae661c4357364942cb4bc6bc25339a0709e55c89ca6712b52e3cdf69
z1f45ff6651350c339b0f4f486339fc8f972162628d54d641ac247c5361472e869593db766951d0
zffd5f51ac126250c1f965a0ed253a4549dd3194c0e7ef8dfe2e5513750f38916491ee814087edb
z70444bee23f5df0f39e8c957cea1816da457cfe7abee21cd46f76a2185add7fa269c777ec24053
z965ca9ebac6caa1c769e03d3c9d9f9f922a8f99265e4b5904924a43e3fbcfdac47bd7b22b4b522
z759f47c19e2fa66a986d87c7d6fd40ea1d19acffe6ab640be02edd6d589f3076f624842ab507f6
z458285d545122e0e73b28b89fc4a279b497e7780e71cfe653c7a999b108e584cff8be1d085ea84
z85f379db8aaa2fa3100f55238f18cd5dcb12481b83fb5c64fd5082511f298f071164b973173bb1
z7aacc45b3f6e47b9a75bc1a3c31e5fb461deed81b15def750481d369025fbd67055be1b9186fb8
zf7f06b235e19bbaaba7e4984d2b2e128d9bfff901302e6a173cb124ae9447df9742dc6a381249c
zd8e1715a6881eb430468041434f78d3b4ba041453798bd02f3702b23136762ab4af17ec3a5c744
za2449a507b295bb53c2b84da412a12252802d143c55ecd746c25b442a8cd7c910ca0939e6a0777
z5b6df0d6aeb082c59e0cfb60079316b7b4cc4e9df055d056f59cf54a9220035bb15f7602805820
z9e5ed48fa0fdfee0cb4c24b3d5fe96e1a361456ecb338551d66708fe98f0afb1bb2c62d4602dc1
zdf75a8c69e24b8172cc37dff0d858ffad86183e3ce8275321f1578087ec4686db0a32634f0a1c5
zbab420d5af56da32a7101fd0116943f55577336856543ad1771b97d17a6aa2a20376edb3a1055e
z239f53d1269df70d48d8bfd6ea25153f9594a57d2cb83bacef7bf4025abdb18302d12f14f29c85
zba0b7edfd0243ee92ed211ab5d36ce8e355b07112995f118a1b424c577af7a42032ddc4287129f
z1705edf1eba7b1959a4196a28a038b246766a07f6f464108cbcb85140ff23bb417c2c47e6ab578
zec7aaf6a7cdfb71454d31a8e1181cbc880a5290ff179b008cab5373ee05d303f08a7c44eabb13c
zfafc57daa934217f40bbb4dd3420e797f0dd1ab769c26bdcdc2e802c97d74b4396ca5578a35716
z112a2ab8aef954c9bd5c49f670751b2234fc7d7549f7190f73ea94cb0de10d608af7540bc5c8ef
z675b83b52a5309921ed8e8b1b97060f397c174a468aef758e76958faea3c58eb995920b22f47cc
zed88eaf6784bcb79bf60c66f6bdff656de6003f1479b9a109b424dfffd53a41c4064586fb375bf
z9e33b9ac3d5c10d35694a9fa6a99f21a62b3f94627c6fb586a9c784b6539de076e100ca9b3f7f4
z1995765ac8f2362cac8e05388c080d7a0ccefbfc1a04ab6f3861287c84482034010ed0ab7579c5
z89279881b1525c96f63ac422b06518eb3e6bd479fca0f9a5f9f5d0aaa01f1cbeace62cde713448
zfca18d3b9d37fa4099ba6e30729717e54946643003ee6cee261cd96ee9a8dd38aa770aa2395f79
z68f7a4dc49c60b1a1130e5731c503140cfd38cdf643c76e47f054b498455941be318f88892e2a0
z364908fba10c56fd347798168daf900bf776643decd0bcca2b0797422a505f81d20fd554e5b3f1
z7f9b40debfa01cdd42a22af4f800c7c41c49c752cb37547302ef42ce33c490776faacce78916ac
ze450a33fc9a8d522b3d4d6737376d2f2b0199ae45fbfc03dfc261194e6f2d5a1792c9f0983ba33
ze97ea8110dbaf1a1e8866d0b57d88462421b1941aec3495de14078855d72ae87372479457c50e9
zc08d610b8cf4a56ae7cc53c4f87ac7ce26d110983cda7e1bc81084e0c5ddb7991fc14b10160b0f
zd241df970c5e12432b9f48cffba71721f77ce6880a82bad1120972c62c569af774841a23fd1caa
z65612e37767880c7c9ec503919fe9d84a2e42a14ed6b4d59905b859836fa9d239367a4bf4a07e7
ze221bbdd6ef173784f29f14592fd376ddd75f17c296e991db8ea518eac4047e4ff5624db26e87d
zd01c13cca57a47611579d5d018ded110d2bd8580385d5c8f67da32aebef0d0e4dd61ad4b508baa
z37d8a9eebbc157b2fb0921684e9a72d610e526c8a553544f00f8a691ecf9314ae886ab3ac91ee5
ze8185a8485e56b852756b494275f4b1ed54fe384ae17ec18586de5ea0c9b81e2e8c764b5603063
zdeea4d848eb20c8cc42db17c4e6bfdc9b1d472c9a5515c9ad40eb666dc7d51d57f3e606497a110
zf6e7615439112aa7c8e0b2864086c3d16a187cae1b7ed87035e021f30c12d98b25680565b07cbf
za64dc96f8db55c2648ce41e629af24909e92b31a18bb981763a9b40b0e5aa4b4bd130e8db199a8
zf1bd65118967bfe545b6d32bfb695bf49f5c83dab8148094eaf05b9d406d43f3e84a21ec978c10
z81ccaf9cec0bf4b65f35d6377f72776e422c2a80b946fa37290def69fe041743a6c5aa1ae5b56d
z185619c5491ce1b0a2ecc80b417287241d14045beeb25b9b442cb08f3eb7e49e2377c54317732a
zba3312c84195b57bf1b2d55443db6108a54cf2bc0a951b0c4906dc0bec9dd1e3b5594f89bf9fce
ze782e7ba6be2879de20fdc5114732a2b90a517670c53874c6955ad86c541a3c5ae356490b79de8
zd8f4d4685244e8afa9724f693e38843e12eefdf6be13084f612a33a5b7ea5507031d5e9ce0040c
ze8c7fa83cbfc40ce8668553d6190eaddd292cbed24126c1a4daccbce36aff6e3c6a767e6bf72bb
z5e46602a4224b249d8884da09f1231cbfb2d39c41c5f76950c8b58e902d96034e10734afb4614d
zb1414284849686bb1c21d86f2e5d522f10fad3043df5f547c95dcb6a37bd8117917ed2e8f2a02b
ze6eb4ed58d101874296055b43c5aa2b1c0fa1edd03604ef824eb68440dec25ac57ab13c479c794
z15313c5ad00441133d8ab45fd6cf91e856f7cec9a645a526bcec64ab80d4bea9f8b4e54141c112
z9afb62eac934bdecee8f1ed1f3b5362457ad222fcb95c431389e4bb6b8b19c440a0e92c2ba3be7
z60c168b3d7bd57fb5af88b5a2d90e3593a4086439841ceca19d3f971bd8aa9605d43e0d91783da
z3157682d15d03a752f10bfe4f228a4dea7409cf08ad8559d95cde278a6e2f7deac61b4d07d1f1c
z9fc4a83be661555de639cf4be50d555f2cf61b1b6c76255752d2dad0d3f1df7b6b435d10785327
z4ff07f2f3e0e63a7968a44880f17f7e010563f4dbdc73858ba2751e0d1c179c79005b865abf551
zaa71a9bf9044e23d2a407cbed3155c754fbe25d2cdd5776ae16f43d1e4585fc38ae206f47a0acb
z26f74bbd5bf629f465aacb9fdcc1269908d9224b8660ccc6e78c150c5e6da1d265443059afb725
z4b7ab9a21ad1b36b123404c3fe96e0025b7614406dd07d411ba0a97e99d9be001ce7ba559694f7
z2c0679131a27955c3d74482c02f8e3cd811b43d55789e0b18b37b15eb8c316ccc2e6fcc140613b
z6b34222a5d387426060eef70f11b724eaabf060bd0a1a4d2dcb2070bf51a3863fb35ce89ec82eb
z82f61bc5b07a4c88ee39440ab483d78045319b860378ad1be011a3359ad6d031c3763186c7a337
za2a9d7d0503375021737c72f6d1271943154701f06d86d3089646893b2650a54b8971ef79bbced
zf5215dae7a66fda60aae0f2038f7638476c1672193642f25dcebc9a48cdf3bd50d5bcefdb8ba49
z570682fd58007bb5198c52c80ca0398823f8cf0ed43dc084d79e137d1cd389181eda525ee43c53
z0cdde28a14fa7e3c6353bac618f3d87e9dbf9cfcc81434d6528b28ca4f4dc4f210ebeb2c422feb
z804f19296bb83427ac652218bae10d38711dae8e6e9760cb48a83cd500e111769aed868eacda52
z7565b4277c18e545e66940529d8342aabcf78cf63396d3472969fd06adb6fb0ed3d9d73fd15a24
zcaf1b776360c54a77757dc62b8a28f8f9418718cecfc70ef9bcd24a5ab848563f039660d8da6bb
z10c3f318bd997d2ceb5a7b8db8aedf4028c3babb3db2103c500ee994130256b7d6fa356bb68e6f
za76492fde24d90118f49b498c779257b742983435e9fb161c71139187599e6b83b26cd9f3dac6b
z380bb5c1dbb82bdb36de23883f09046a4f2e67bf87520de21101c19cafe89df6f95fc4a026f431
z7e50bc45dfcf5ad24d3a3f8267c48bef91ad9b8bdb8ec3ee237d91c0385793d04bd14acdd0fcc8
z163e4939b3dd4a5f9caa05b20d8acefbe18f0b785775072eb0cecdece7bd0c5fd0fd9f65e2d707
zb73cdb11e52751d1a4d6502cffc3c603f7c719543d020f34416af1041ef0da6a7380788b703f5e
z4499dbd9b09533e7849ee4d0941ec13f87735619036b4c354117328ac56d9a0f832cb0141217fe
zd8ccada315bd83f58af718c74db370a74fc39fb920ee9b13fa4c8fa738ddd9604042742e539e95
z1d75a2cba1795993e166ff32415d887ac64386e21d58812f79eeb80b4ec086028c655bbb35c95d
z1bf9534a8a611a94b1fdcaf2c7abee66961481bc7ee09f37049759a240048af86fcaf7ee71fee0
z5a9cf4dd045e32c31470b7649cc8f7267ceaaaa390a30104eb9edcb545ca1febdaea279cf35573
zb5b520f73a8c887bea3031086ee962f4bb22e890a846d19ac5c8b8bf40a1268fe43962196ce1c1
z3f74fae4d833323d4bc6bc2c77460bdf8b5c9e3f2fdcf38470a61a0c35a23e5ac54ac40e1dcb4f
zeff8a7f49a56dcc46201bd5ae18fb8bfca6cad9f94ec9c1bcdac0ec70ace07bdd41df50f35d4d0
z45d0a8f7b5e6d31c92670901f1062cf5d97e3fa9bee086b04febcc5867834fa4c124ac647fbbf2
zc4a497ed59103418203e84681f00dc0a2cb91759511c8fcb929b6787a2493a5388ed11dcdc21f0
z8e74c7819399442e6a911b3fa50a07bf163804e9c872f375e361447b7182b6bb9b7a3a098abb67
z0fccadbe311360737069910ebb1eba2267fc7c70a80eb01d3561c8c6ea8cf4ca1699b5b6a6f215
z88
`end_protected_0in
`else
`ifdef MODEL_TECH
`include "qvl_encoder_8b10b_assertions.mti.svp"
`endif // MODEL_TECH
`endif // encrypted_0in
