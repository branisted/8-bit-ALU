`ifdef encrypted_0in
`protected_0in
ze74c34e226135848fe16db9ffd31815111b6d7fb642c521a3f628cf6da949865580b22efd062a7
ze90adae0e65e66a2c36a587d0a790699161455169ed55a01f2084f11770a774ec4c588039b380f
z6de9c5084882a40b79a175f5c2114b2b6d78b070cb806e1c0aa9258297f4687ab308bc470f0040
zb0b1de382961eeeaf2e279e1462520fc31c119af8f2b214846f56c2b3cd2eadbe4099496abff18
z15cec83ec4a77b868344aa20ba7360908f5c0de2a79abf8b3534b883bb12180f68b5d4beb444cf
z3fba8f13afb0abfe8fcc4294810f75afe452434d2d0f1166236c82f76edf1e12979f04bc35693e
z32ae028996dd85737a8f5adc1ebb94f39c940246e887647b64782cd7ab429b0544c173176cede7
z01dfb26b1f73408344a52b7e1f117f12bb9c8077b34876c2e6fdc085981637012dc9754765e1a9
zc512ce062e0b8fb16a214591f5c81e1353b900a611fe1f4886b57940b41b7f2ce99a7b84b04b90
z916f717e73bd10589c81e207ed77ec660a8cbed5b487fa50acde1b055c8870bd8676023f21ddcf
z9c98cc47cfa2d654ff1365d1f45035a045a66c5dfa8279050262529d2cac9e64fd27d9c7de62a7
z731bc808811ded9016570962244887f98fe5440167bd0088f2f049df882af501358497c3b28776
zcdc5426c7f52a851c35106bb93e16fff984784052d47316d4a026d12324c22b69566cabefdbc15
zf430a9b815bcd65d9af292f33fded2fe9486202d62f3b4af3be6628570b1cc01d7745db441817b
z9a5c0d54605e3e1f48d27cb7f957d398a87a10a5fcb6ae1dbbb1e84dc2d3c3bb2eb89d3a77fe31
zdddd0cb5808fae1724cc6827c574daaf656da92984db0908d95b40f1a66bcac6f983fd2ce7f5c5
z465f22326a80490f6d92695edcdb1ac875da5d3d6956a02e89b2f7f0b78f3d1e4b127766b73755
z0935532e7302fe5965c7dbaf32bd89ecf08e00087f5c2250fe97aff057ccd0d1eaa623060741fa
zc9a2ed26eae81594c34d6a4660fa212b9f2aa7088298c592a5e6421a42f37ae97f3ae7e0e10e10
z75ea705015da71dbed49c8638109b3fb14607106367fc1dc0216ed06b10ee149d1aaae56727c1e
z916c84a8de9861cc1d73bb54bb2b8278b109486512291095c0714e9b37789f492e8a84ed9649d4
z03c5c08eda1eb680dd1f73fb499f2dbefad405e9e37b1493f6686f610a136e7c3ff4eb94240a62
z6a26dc85111ed40f9c95bbbf5108459523c5e5a70a7b6d8b239a073d46758ba7b0a920563012cd
z3225c6a9792adbc90b1b567b26855ecbad460d4c3e74ab68e63500040fa520e83efcdec3b751eb
z39a4438d26e2a9cd0178e8a2a594ccc92142b6969942032646d9f48d955d6398c2b846f2ff1d86
z7728be8a2d3208129cca5776e8f67731ee12f5312862b7a9032a892c1dbf624c66827c0780caf3
zb0e2076da57ed8d207d55f5537534585743a4fe2df50a6441dcb09eefe3b93b8da2acd5f1a7b39
z270486063b973fd41523885f281393169b796670abeff51a6047fe7b9da58130a45e3f54726089
z285711129be413d340f0cf4f3f2c2812861f4f7c7111f3130d13c2d1ba16f500d2bd8ee7836c82
z37907d4560b5dc662b6923c4e7262c39ee25ee05060c309a7672222db5685eecaf53fd4b8f891c
z7bf0b4765fe0429f9f007281ff2b2ef9f299c622e870b12181aadc697dce065fb317dc7f340f3a
z29a0b258a7f30c281dd86068b7566d0d1ef9f833b92399b14d7b99372ef9b36c2112761f654f6e
zaba903ccd4c2949ee3421804eaf2f4a34fe0f6417c2b465e3ff7616533981f24f24c168bc9d6f8
zb32ec23755992ff59bf5b981d75eecf1bc402127d3016c02a536fd575de556c45bc055184305d0
z1f09e081c270ad60d5a31f127e415d903ef453a7ba4b84d6a4bd589621f8c4b08692c764306ba2
z16700158f46771529cbdf78af20d775a8aab8feadc404967b1ca04978744d3bdd8cebda8df9425
z9809585809fe147dcda030819ad21f8dd00035a799da6dfd59c97c8082182c084811f340e56a68
z22734c91b5bf62a2a50769536640120829fa9b621d4719275a0f8d7b99bb18c3920fe077cd9a39
zd92ef9115f01963c96c4be91fe5bb67df084aab526a8ed6ac8e8ca00f1cf47ac5d4f791d303c52
zb8364877ec0866f0e8701eca44642bec7b51e7c8cc24346fa61d945770c94e1b3a459c4039b66f
z89f0e545b486ac979f910fff3e3dd4d9d414c495b6c9e6ee82854195bbf32a86394de5d8abf96b
zd95f89a1e21adff81dbcd36138ed687e0a904062380dd11a00603d2061dc7f1f58c08ad85c67a9
zb12256eaeff07f238e84875323b655b6173d797ca3cb0745001f0650ac83a459882acc017b740e
z3e8c285fa878c31be03ad0df6fc686f2b02990f4756747284b7a68a1ce91adce13406d7fb64928
z675b006c0ce9d3d06fd548cbeb372107e60f13c5757d19a1503fc9069484899730d3d3f9a73f5f
z63e8edadd77aa3d8ad8c3c078f8899fbf42f81c3707382d60911314cfaa8d45ba7cc94a5cebd3b
z895419ad616fac9d747b7a6e5676f6fb63381ed2f78e77ba8b179533acac54270c8b78bf2f0d5f
z2ad09af04b19b2b5e040b6e1fd0a487a427e13444bdcd26d98eaa95bee75239d8c7e0e7fc4d31b
zb8ee8e643536db9979a9bf91e335ccd6b64abd523e88e914f83588df5a5155ff170fbc339af4de
z4e502310c850d658d7a9748056e14b54eef37a6d2fabc9e9cb9257681472e73bd062aa5add53f5
z02c1c3a3ab714f6f46c63e7dd9f0731987442c383b8a0e6b295c4723c57e754cd5aaef5f4568f3
ze35aada04ba917647a525cf6944b3a74f383c8c16ab182cfd18ffb36f0cb7cf8c41026e9cf9575
z3b7959f071456713deff41efe7982817253b6025820bc21efa6ed179ec2bb77f1ab6bf9df02cc7
za5300ff8ac970098669d8314cee3e1cc59a465f70a19ec526d31da6b5ff56b78753f1acabb0e0e
z13b199719e29d50b87b329cc690033adff016304675173a40589a4ee796ea7d07269fdddcd09cb
z389154aa3ed44febba665a03ea870b9d65fcad44a1b7327659b3cf30baa30e40c94ad35188595e
z2a3ee5fca3550d686d258c0255b79ba0a7ce4adb7582c20e541534826503ee7ebadca71856ffe3
z4151adcc6d6ba6c6abd0f086370c33279c2bed0ae9416a1623d77cb4e4449097a0faec6b169d7c
z3e6b1d8c7f6960c45c7e826a4ec5dfebcddf27b0a42dbf7ba211476e39ec7e509e31a47c0a8227
z463010dfbd8d3fc76b24fbd56795d92ab26f6f9a289056934d1bf6099e9a710b390877fe6b6bfb
zf22cb370dafa2f20864b2ae0b7e4168cd588f7ccadb75c37e46e692fa116d7158408ca73779e1b
z50a0ff5d7805bb1613644ea9aad0ee24f5882d7fe2cfe130438e6ebfd3bbe6c94b27c0a814ffe9
z0eef8bdc9911eac610ddf9398f9174da588a11cfb6a2fedac67367e9a54d34478e7560ad2af780
z655ebdf436e0c60cdb88d19f2aa5125e528fd8463e84cbc6ef62002891f4659574562c4b21a378
z3af5c16bc52e96d89abfcd6e02dc54042d7f912084d7d3cb96d314075757cd3720e779151d37b1
z530d73ec49e39c625f22e52546ee00515bf89141c90fdc6d710cc1f05a0eb4d474ad65b5f1dde3
zd491fe47ec9fc66ab377b2e835dcd97120a02d06b4d04488ea8e318a2fa8bd5d6dbc4c61df0086
zea1e7c14145ea42d7231b28a7956f4c041a8ac43b0f769bdeabf9fbc7ee9d7811a333c47d8ee96
za0f20ee0496c3b8faf10ea85895b44add69f429acee5acefe288d326b29413b37970bf550792c4
z2afedc5868034b5cab9cc9c1271b18e2979983d533e791449176ef387fce1cd59cf0864e596105
z9e8e0e476ea436d7c70f000811dd4e482610f160b90322b4ffb8e3562b3636fff00a1d9afbd2b7
z70d19969fdf96a34a0a59ca0254edb6e8936a242d09ca956b45d7b613eb44474ad150396d04691
z69d4c18ec0df7728541d8ca0bc0713e46a3be9d39e2ced35809cff3923e1daeae74c6735848bab
z4cb3455b94306832a68ca96de83071f3f5c37fa6339598d9c318bbf0c2e5c672d8b5c68757f4a1
z095396d634ded67c717a2a723eb7d7ed56d06c87b97c0487601f5c3cf8afdec25d3d01b26e7a2f
z77bd389b1588f35779c6a4d1ace85643a4c87fbba54951b372fdc879022cab033968112954d8cf
z76711360cedd7614b99c9b0d906f4abfbf7d85a54fde39371ef852a104867422959f3ed88c7ee3
z1a43b0d53c53c79944884988c279b0fdaf6116913985934a5220929c7fc9212e132472d9e3ecaa
ze421526b55e52d6e15135355b55a412daf4bf902413347b18c4d68d27a7b0f0c1ff49e7918b90b
za63caebc1598df8890e7a1b3db09b6694afafd790066fab8fbf34a8aff7b3d397fa85a1440f14c
z53c3606ffc1e8a84a14d06dcfcf6994998ec50d18f83580177c28612c8c9e2665cb42cd4dfa2ec
za76fcf94cad6a3d608e0f34e236d7ebe08e871ad7d925c65aabe906cd19c2cfd0ced2a50e819c4
z62444c3a23a972a183ec304aadbd847bfe2ac1aace77c8321090ea8c0f35f7e046353f439f40b0
z629f16a06df1de0ad96652c8b69c848813102ceb19a6e3cf2df3a8536898b334fd591ff96bb6dc
z0c4f8ed9565d16ea30fbb557a69e003b5737b8554a7a671289dfd6bdd1433d6d3145490a5f9e35
zd2b4dbd73af3323a3741ede2da3d2ee04a8cb3519714a27820120192a11640c5bbbc67320eea79
zaeb5051ec7080014864af45a7778d6d7c92f87270704ae297974f508316e98112ad75a80d0141a
z490137962f0757c8b6dbeffec34c53f57c344fb62a29f008185a940fc25148e09652eb9a27b731
zeeb48a34ce3051bf57a94c0828c0aeee3a181053a2b08e44fbeaf8532e4d7b066b9e6ed71b3777
z0a70fb0860aa872e4103f5eca3c5db0fc6339ce3362387f33ce13f6a977c9b992c58069c34721e
z2635204c9301e496adfeea06b0eecc12c0047454da3172f8f461547cd65ff7e745d332181fa54f
zd8b46873017b098078b6874d3a6064dd80dad2e879a78ad0e9feb50577e076e9a0a26048cbe1e4
z4f1044f4d7fbd28659ae2e0ecc0be78d54411b220425bda866dfc4a501e55adf14a931e61485d9
z0467de45eef6fbf504e28acc99b22e4b9bcdb3eaddd752950b3977bc6f7130beb65cf2cc0f20bc
z41a923bad525e1da1e7b447a1d3ec3724074d7eeb8f60da71f5ea9ec81a3f4f548daff62eb6930
z5beb56cd5278194e95872931ca295f3637f6912d04b1974b1991fe8ba9c6b382a459d23ccca0d7
z16076ed160b80be5e59cdac3381c2ee64b029a2bda1b3f5f0eb61b8e0a95460b76e3eda1e61afc
z6e7a483667e78f05dd7d8348b98035475274878071162cbbd865687d619bd1fd32a30fc121ceab
z431c3eae4697310531553f97ea05d89b634b936b502cc432cf7ae5a17260536f0836d17fe52540
z416e4c6ee61c80d65033a74aa3a581c0a5954ebfa5919dd6ca45aee93417d4c1d34a26498b638e
z306414239145e93b5803744bed848002c8a4d53c7843c97d3373b1d946254afcca12d25a6d2702
z1cb8310a589a863733e0d12b69c8c55c1a20f4f509bef37e5c046ae5852fdac90282372f81ffe6
z0516fa79c724251805db80d9ee25b5dc671c83abd0ccb2b8102643401eac40b6e1385d0fbe4940
z85812dcb4f8a8662eac5c214bc009d13954ebe5b96645f47c4c0e436108e5bb5083ede58eeeb5c
za6653396582a0a5bc57e98f11b54cad719d8b3af9e9524c89762fdd805dafee2a13ef2322edd51
z6750b6f001501b0f3552bbc210c63071908f193dab8ff90152634190d25ff57f0637dcfec5806e
z916a0ee98d2428e4106b04d5a137ce52271dc25c8352dd6c5b51cea85a94269c60102496ae06c2
z2c539c7c5a8772878a781f4848e02afb36811837811a28f2678c0deab18da088cba7326385b717
z2d324a177cbb1ff10d1e03e6fc5cbfd0d0dab89f8898adf1e308795595b4444093b11044c8d833
ze40d36a3eb2e7e179b3429306768e256953f01d1ced9efec45e1c11e9caba9c85f38fab12b4c0f
z066b3de8193d08d687f0d3d7688c737413035f0aed9206dddc1a26787b2117bae98204a2aa01d1
zedf19648dd676841e5926804a26f4633a6c8c19c74909ca4561686a8e47f9bd8ad8f5e3990257c
z66e30313ecd21cb005ed8d5eebe834996f13dd4ec9e2cd4093532a94cf98991a80f5336f586083
z5cd32ac426e1cd8d4323a7bac7c36aae0f6a239f0937d8191233705df111992759de6e5d8953d6
z4e0f9e194744db890f5ac35b5cf7770c6f8bcf804f4f86c84ad7bb03c25e76636f17e58e57cd56
zd909e8b1e83af889d683aff40c975f3839d170ae8f0bce4b1d32b912b1b9f7662c765ff6d2e6dd
z6554ceee969ec69a6d657d96a2f94d5551c946ed79cfa9259947d783539f0e483eb97dd368cd96
z93c4c6bdbbff64655dfba05f5f095753f711ce9ee22e0bbef6820289cdde1f8a9171cd537db3c1
z9ba4c090b2fd2828e19ac9508575959d04eb8449ea5700bbb9594005a428dce37b95f094a1eea2
zd960596bd8ab05efdef048664b107c66dfed9538c10341c6bd16dc11ebb48bd102586c2cefe41d
z0ddf76ad9547077f33ebbed50f196f2d18c66109d8c4b5aa7fd651162b4d1b59ca40c85e8a11bb
z62cc628d4f6095fe29158d0a80c10c83570afb18beeb5501add9846a8700e81efd8e3daa584367
z814e59d0e3ce714ea3a53f525a6ecddc3684005397aff929044fad2a72942e667d5d61eb1505e0
za1f63c7f0363430eede03619266a8fe7e1232a0caa9cf9784d2af70ecc85d124964d7918cd98c0
zd78f0be030f45af30fa5dfa48f9dd263d607fac2389a369be5b2f9e8ea45c74b600a17d2e982a5
z030c638326d512ced6dedfc48a9fd21b2bfccde09d714fb4d5270c0d260dbb312958af7a4aa617
z1410c26f2a0ce570f963cfa03e5292ff4f5273aaba2625c963200c9f491cc68db00632bd6ea888
z196a8a80cc5b244eb8d33f354d922a899716db98ab083b56c3fc6aa379b6d55e15c691f7b60c40
zeb8bafd4e060b99f9710c90af9164ae28b622a79ac2a89b230ad2b046afc51385330d3ebbc5d78
z24746565f09c4b382e34e1281228b076cc8b029b1a6a140ecff40e1a65c87b847080f0998e6095
z1adbcd80051c3575dc5f35b84983d76ea7bf0b728f03ea01536845b147df3156bcd42b4d9c4e2c
z53f1fd027556dcb6ec7b231fe4e80722d4c360af3099bf8db276c3ff005d0fc8cb3a46c18b2bf8
z19acbc35ff8a78824868f8e16fd7453cfa9bd0ec45f435dac9e661d5e86771e12492d89b5d6dda
zb69f84b155f3675ae88935590352a8cb4694a5394a0a2fd55f3f6726acba2c970dc6c6cb200761
z91126010c4c7c23556b3e701078dd650f65607883c5ca57e5427f3c7711185a7fdab846dd32b51
zc39f0c0973ab20ba5049aa54122dae10e71bcbbead7b6b68797946b93766565a7d23a04ad37ca5
zf2a39988dd8328c3d80078308d94354da845bd51d402af9444e8874e6a2492f9de012d6873d0ad
zf00002af209056eac7bf00941f8058ae8f53a978ad9b7bae8bffe3fcd011f77aa25e8c00f7aefd
zc3404a2a0283b54209eec97fe1c0c8f2c71549d7b014c8205676d1e684cd664c0fad30c8e5ee55
z195e78c5305b05e041a16a38396fb4f8885dd0c39073ca4641c46622a562abc392b5e99cc739d9
z85cbec02fef7d6f669a482fa8dafc71a5bbe8939aa2b37f62d5a3cbd94da69da5fe18eaa9125de
z307150d9ffa8e77ea3e7f56cfa1459aa1d82a031589701eb3bad73cb893a415e166224f4bb512b
z14d8f9ecb3fcff9c063e373bb07a737232f2f2af3e6702e1af90a1774f327a741b2567c776aeda
z0b36ca39a1e269dc7fe14e795bbddd308d92cfea1833edcd2de0ba80950ab34ffe18c8f145650d
z52e6218833ea73d944c7965d19644b571fb541d4d22872153a724ec9e84a3fc5593d505676fb3e
zd41673bc4ce0abcbec7458eb9ec599e4cd100a16456562666bf17baf93babf9b9a4369adde4589
z8a943ed65fdc8d9c01e158608931619137c231424ba319b088abda073beea7ea9705d723c06592
z731d1224d7ddff33003dbd8ebc47336bb18b4e5a3b7b22235b88b8e6904e99dae6e2459e30c479
z340152b2898acd2d1668225a7a7ece0239e96b83331a7b3ef8c39de383e7daad26db327953ad08
z200916be2116ad594e73a6a419ec15350805a95afff7aec844458b399400b45280dcf0a73e8dcc
z16721c02daebd8304fc418a802e9ae514a2bfe0300802b3767694fa05ffe2c9acf8f3ec5a73e3c
zd4ce890ebc6875f34c53966153a69bcd15621880bf68686e4dfff4b6ec86acdfffd5e9d2e45348
z59cbcedefa51e8f3d0c1d51bd476d0b865a23ba6b9fd27150644447b021b39cc9c193b14d6183d
z5b082d887e2594e6e72dfbf774f2ad5d998f7dd5af4f28dada81d194aeccc6d9bbb0f61710121e
zf4fdc546f5946e25a8225199b3ebf0b0433716a6bc4e1d59ba8b4d23fac2ccdd22d4b96790ad45
z744191eeff50b48eeaad5d7cac9f5906ef5008afe17165de7d139369c24617743407e7c8dd952d
z59e6d55eb417f25d129837acb8e094632e27e126c9b57eb26715aef22a3a07b5b81a3b75689a82
z4d240c72c6cd9c34190c75e08fc9ea788e95bb6275f84a4d94b9e3d97a3286ae187074e3975166
z5cec2a4393dd9781d443902b3a78c80b454f711e811c27dd64de3b4f4c59be92491eb3caef6ad6
ze87b0a46b126cf3eda2c670c890e60fa4c2f59f94acea2d071a9d2386329c7f07f24ce2ddf8fed
z52408de2a0f080e6057ae30b898b2da7309545b5ef5b67b98ac23c205935d43bd71b3d014c7660
zb928096cd94afa3562a8678ad6eff3a7b5491422cb09e3ec69757a152561999bb5b4dc7a10f938
z79b184be1f530dd12db6623b3a15967b658592027ac906194d6e79ee5e627f4eadb3d619f912ab
zd753249b3295a6391825e908a14e32c535481cad693b7875fdfd6fecd1e8e5c550309e71b18ff5
z11cc271c7ce33c485295d5fdba7e5dd37b04bb9ded1cb2fbed908e8f8296495530713eaf36381b
zfecd94ecd5e30da9a9fc5d48447bb2615d2e77bb7c137816a528cfc4a71d25d6ede82bc25c6199
z3ad56c7eb0b3d682293dfbdd1e45fdcfe8ecf3631a5b9e49ebc6a526544f917336f4b99096d373
zf207a2d4ac34ad3fb56d2aefeacd762264fa80ff89faaa3ce7f5bfaaa20baf0b4652b116e5cc9e
zdf756f371ad1cb134627fbac9050dd3091a274af1c56aa61448dbbf92987ddb160217ac94d9c80
zdc77ca95d2d82ed6bb50af16123ee05c25f9db1abdf3ae7dfc5be385e605d0cada3dedba930e73
z5ea4c03c6c8868e11e5d639f0e7fbf8c6e33ff8c8ac39c4cd3be0101de5111510b18d233c89c79
z9e1f094652a03881be9d69eea023fcd9161fb9a4466062b6ee42ca1c00ffdb11a08922897be076
ze4fc127bad5dd79b45a4e9331e15d35c6b8de9f6523e5b1c776a2e0b0e2763f5adfe9caa7fe67a
z1c16f9463cba7fe990926d1f5ea1fc5808dabeef4aa17eab7b9952a4f75fd9e26264a691714b61
z38133f980615600ed3faa0e8cbace7b37710b76d8a8ea90e3092c2d3fffed224c4ac7589f0d76a
zde021bbf019688a9ed99c48768b89aadfdc867a3e372fc99e58c3df5d87940fc30fd777e315e2c
z1f2c7d8ad967e559f9de103f9492d677c1fd012891247d5901859fe8e723e7144877a02df66269
z41c5d66ac41e0997f76eb5f67aac7b996d6374ebf1233755bae62244be68005a71eb0b28e6f227
z57a6549c2c72a219a90a790c6c358989de9487364c1ac34c505df9f0de056ab612bd445f5e37c4
zaf630647e6d5b9c1629d5f0aaddd58fcb82086d02e1213ecb9ec170c8b3eefd07ea96e733961f9
zf910f9b463bbbdec12b85071fd494ba568188ccaccda82b64c61dc0d4cd5b2f2db4a07abfef09b
z6259d3d656def4ad8a1427785b563d7d35899a99b733a36bcbf575826037b068194bc63ae8d996
ze20f5423e30e4b025415c6a582db41e70185ca2c974efa339dbb27bc8292f68129e26a40194dd8
zb1602e7f39b47579d89d9716c69282840af0031ae17d000ca6b7903a513f71a349e867668ba11d
z604f9f034605a5896d133de77a9a1bd0e5b13044cb8eb365a1516b56a6199fdcaa9f4bd8b4ab69
za4d59ae1f621931a77d712f29953007a3b205de93d1f43b0c04dbaa4ab2615935748f09ea0cc02
z9d1dca1aeb3b668bdc364a8471350bcd4c4db6547a7727ed771c5d665f62ea7eaa1ddc98bc4ff5
za143809183fc8ed9198bfd9aaa8c3f7a3d4b50046916d4ce6cb387623ff2453af14f727500b556
z63f44efe455d9728351e75150657b7f42011dc1f1b6f51da1b578a1a9603a651e91314267540b5
z28031ab987f69f600a676a8701976268b342e3a169ca0e4f3cf0a7eb2ee694c0d2a4ee799c57ca
zbd24e9dab478434d64b5b1a78ef7b72297a4a0129447121dc573d2bdb161e1da4bc7016d411f3a
zba4796f43a6e4b696d8d3e871bccb1b188140d443678a671608b9420073ce59bad54ea27c94661
z6d83de870e1191e24272b07f2dc7c1a7cefa282482079816d0d560e072d6f831f99b663b1055dd
zca53e920ee36ae34b037a20056532f1420699953e61e56fe525118c7f38ad685ec6dc6a9719eae
z4fb6d4bfbb88a7f65379433a3758fbc4e21459c146d53e663c20a6f70f3a9a1759c31222a391f8
ze3a8c1aec515bb2562d0877a3bdc1da7b08cf6c222835a2994d5e5778f5727566b7558fd8a1d8e
z1c8eda28235e6a5ce2ee7d007e178f10934081b35c3ff3402353f7fe853d7a2814f7579740cae4
z8f7a838c450bdd4291b13ac7b5be21c188b64233e804b7f90e833d99b2f442ad5c5eef65c05b56
zc159a9d64211e54cfd3adb34ec9b80da54a13da14c77254652e71c59a7bd2483ab9b9e90219e8a
zaba6dfcf560f76214b819d956c55c47e154a2be73d80ae2f80f32be7127e8e669f49408ef50f56
zdbdf7407e5c367517f716a08535c52d6db6bff60879f12828b72c98336c3950d27e01d591cc5bf
z63f934d9c025eafc66ebe800f280dd3376dd2fec5b50b3f074f9c612f7b6267a2ec96fa5449dd9
z30a834449aa11f177540ce8e74cfaf5dc7bbfc9df490f279c461901b76196cb735738a588bb038
z62f981f1a5c6b13ad76d3dc9e6b5dc6991f6c3060d8c0940fc9f661f63e91ebe1dab039531c4ad
zde2441ff6f148fae89372f2874c1d5967d8fe100441a92b4fb7cd610fab30b63762f3799533810
z3cfa3183c369a1d47dbbc5690080ddae15ee7c1830888a6eec12ee6f96429b2bc1c46c26e7e64c
z6b842c110e68690880736cdf20ec646b010a5dd414720f99ca09f8cac7652438cbd21e33f2c3e4
z746fc8615fa126b9040ee60b2e4a19b2a52c989df54ceaa0775acb0b72c6d2e1626842e88d4a0d
zdfa5885d43c2ef7448a835825ba910ba107486d70f5b78b52d49998f1235333231276088563767
z31ab251508ff87047209eae26b91b511a566dd2e59198749b9efcacba064da2e94846a74019510
z5c7adddd8a6c7cd29958be391056e65e88ab9262093d7f3e7eaa796b5d962ca62db31da4896b5b
z0950ce8ab98e3487613d9a05abd541bcab4b28d0320c81c0222e5490b5de8901a1c9fa5aeaaaf1
zbe9fbb8dbf99b04cbdeedaa5fe92c7787a597d900a77bd96b20b5898337eaa5797e54f271ef5a2
z835cb698e82d79ebc25bf951f1b93e7ad70b7a38a13c6a9d26464a65b25d19533a7c5f7c134a74
zb3857591f4b6ab17f021450bb8ea912e46d08eb0a4c560a4ef9e8fa36d7ea4d2ee29c2ac904d36
z7d322b4711eaa26788e7d48653bf226ff77635e63b2467b3298ef147618973fef397162012c6f0
z828556adb169d898d1e21d4ab7e1d1672533e93e3aebeb2da06037f4a4c56475a3e9a1135f409b
z91e25e74cb2bd3c8d48f437bf30e52c9f4a3eeeb7af2e107386e01cf88c31ff0cab9b264a40154
z4974a2209e295c02f90cc42832c8b5fc190b65f15a55fd8022c523aa82082f0410eba8815ad719
z6d929a8399862f781f3391426384772fb58dbd554d5a355207897333fec51a0fbe55898ff7d0a9
zb4fe3d23bef5530b3995c235b03c7d9a24befd6a34a8ef4559ff54f439aa46d6116de8cbbc2f5d
zaeb89206e100d6a0121b3971ddafe61e146a420223fffcd485be38a1a8cc918b9adbbc4d88fa34
za7e3749073878ef2a62fc3244b444b9570d07e09526aca2f33682509fc4faba4b4f9231191c249
z9364b8a5e4e68e889fdd29550d8f27a196841b1d7f7a172a73280d806ed064459fa86d33b03a0d
zd8dcd04377382e9c283071d8bfec02465ad84625b83ed96925993352bb204caa61b9a08b1f9cdf
z9f9103dcdd39584af03558a7385aaa29231c18a5afd099b5005a7b9556312d64ca0c1be8a20129
z3e10f7444389d41a6ff1caf5c3f025871497d0c951d78d60f3848ae46639daea10c38738f80343
zc025b42905d92e106451b97a2fddfe92b9da346e50f9847902fdca1a9428f4835c6aacc25176bb
zdaf0159eb6f6f226f4016048904af9fcb2597a60dc66853d5515d7d5438f19139649798549fde0
z3634c2e4549a82793708ae88a4953b0dc065912e06ec6033b9dd123e87453a9bc432309da0161e
z1d9dc7831666fa8ad8ff9423dd19a46589ae63ca9b7d792ea77cfb8b1ff66d1bd8325d8b692c86
zfe24009373b9b3df22360928605bcc98425be8f8b1863ab5391a501500bf04db425405046ba75b
z35efc1ef1cb4b39fd809750368a44258661b6baf63684d8fcf3e73fc8d0fef5be8a66d238651ac
z8a775bbc6369187ab626e8e6f0d04c7058db1aeeb4370a721af3b5eccaa8e8c6eb9bed2f7b4180
z689e1c7606d4c56647f66d0169538145a83ce5b1bf16111d9ae236dc8d54464625d9d5510f85b5
zbe094e2a847ec3ab66c9c9460aad163d4038750dc89caf3d3a938d0cfcb1b1def94f4794bdd028
z472067b241f13474eac315d14bb9022f488a9a48104e5e8e38170c7cf6d5469c1409432167b362
z6246fbd1c6a5365eb4250ece08473cedfa9df95372b94e3d5b6ac92648246144693a35b7de0040
z5f1b9847492424620b06847230d6b55ac11758812ea359b5d5d00b0781f68c3ab879a4beb07dd6
z572eb050c4b8fd3fc3e9c5a92781631509f9ba7df3acb4bfc2c12f7b785b59a7c0c05f77bb0b01
z92dd70ba4d4d4006eeb6630b042ebc2e5433d0ee7f580ede51c86baa07621665eaa3977bfd55cd
ze942ee506416bcbc98eb450162d099443c68618c03a5b4127cf53b75f946e6d24d04e32dbe6434
z4cc703cfe91d5ddb34c7523bcbdd8796f74df1ac6aee12fd41b5812c9e994f3fb555275abbaddd
z0d2740d666b2e2cc6e33733f1efbaaea4b2845198c0ac9942b881f721b7b19e9db74d892d43ea3
z3f77f991cf8342369d6115e310d542fd91e1ccd3cc050c9e23bd761fcdee749abe44ba8d8c80a5
z698941c7a139ec18c14fd9808502c6d805abf703f9d098199ebd24e3c2b207739244102f329d6f
z604f972cccf97989ad805780b4d44df1b1720001b228d7991866e5d62cf0b8cb9b8dc72dec42f1
z12d3daac34aab272275adee2c3860925efaeb5136159679522b55f3a79bab2838c26e34492c439
zeeb1485793077e6925992bd516f35fe501ecc6fad97ca2395da57c70abc0c3f23e7aba5a6ea8fe
zb68a0ee98bc1677dc49e317b0f5f96cf3cd4356372224f82f3730228c7919cd069e14d237160ff
z83502cc33f25905b049689585b58eb2dd28aeabb0c102c0f102c713de7aefe43caf6958562b511
zb558246335c46384c85301a49e38c2d48dd0dc3fda3d164d303de718a8e54f462d14efaa1a242d
za3397ecf10926c26394580f7a92b0d193025b73f93394e5acfbf6d2b448fee1838843ce4f06f0c
zf92e0d66896dc3fa9778785eb4d9502324245f7275ccabcab4b849b5cac6b057ef046b961e81fe
z103785ba7d804888c2ece348298cea2e961a2f1bb2c1ad6eeb804167de48b26c9311c3c1e8a585
zfa6c0df45a106c1e95950cbdcdbf70a92def3129df3c2511dd191010f0929605fcb4bc90dbbf43
zebb8c45a1bfb603ab72c6248458bcf5f5998fd79e622c22b7a97395aebf2806885e84d597ddb19
z81bb8b65b99c9439b6829bd6d5a3cd183ed6cfdc2e97e907cda309cbe3b33c46bb42f9928a34dc
z98cafff8f53d4d603dad7019d979fe819253406485093f804880279fbca73bf2ac38e6efa755cc
z96d089db35e1fcd3e52ecf363edeb56f75bdf9f94dfdabd53c8a77cfee78bd89aa5c9af39c1bb8
zeef66cbc6d1109e588ce7356f3e4dfdcb575a7b6608963740d3ce52d53ab166355135b180c7394
za21f0bb324ad9aee7ec041799c1b2bd3887b06e86894b5d8564900dd3f6f21e95d35191faad4c6
zfdc63316eab9388fe082254781a669af5bd1910f386bef8f584fbe132ffea529b3cafc305bf376
z848d97de23d5afeb463de23fc62f755a607aeac49b890710b87b2bbfa7ebeb4cb954cc83a07753
zc2c1e93bb8525ab1b723f8d554b415d2c193b137da1d4475fbc960d1182da84aa938df52e0e10b
zbd255db0fded1fbe96b583f35d2369ebd4e6544469f6a757ad45b95f1ced650ff61c0f9d787b91
ze48aa14017a975c128fe00137ea98efff36b5e5afdafb68c889262bc8445c1dd683341fc279b37
zce790e3916aef6e6bd90280ab88217c957db4cafdf7d5c636b60e2d28a53c6d090314c5ef553da
zec4be9208804b269a9caa579a31103b853ffea8f21bb479ab040c5e7d2a434ef89ab3db4e3d526
zda55fc8c78787b0fb31d9bcca93543e209eb9c07cf42a843ef5b812d1969fa13fdba17d34b4138
z6f65b028eac2d13fc5ebb7e758d97b00cc7cc6ce3487b13be2125219298fbdbec075793d58ca6b
z874b7c0d9bc9b8b1da471cf7009b1faee14bc4d736d5bfa1883eb91126108d0d4197c3668aabb6
za20e58aabfb2996adfaeab976c836d066d33cd0bb679ef0154e08929a95d87dfca393779eaadc5
zc585395c5d9403a5940dd1a5fbc03428533ebc13aa6c60b8ade8f9b46c35389fe917fc12449d51
zc2f8460f0116d8597f7e70041ed641b30ccde3fba2ac4111b52e6784fd4dfcf4571f588140d57c
z4b72c072e252292659bbdbe2623b82c22075cc49bc1943ae7cbe53cb00cbd494d36e7ec2c8f4b8
zc4c03a0237ae69e3f275cd53af112451073243b0fea2fd0747843ab3aac7b842767a5ef512906b
z6581b2834e70137c404b5df73139e1dcec2741ef1991ffa2dbef9640937b2f4fce55d8a27a3b87
zba16802fe64cd63946d1dcb88c140b73d740d69b49296e1feaae1535ed991127c1f3b9718c4fd4
za5431a927b436c1af5356cd58bc79dd579815ad3a0d5afcda0f8f279f397b869fb7c42777614d0
z996aeb072d11f86b7da711dc4dcc3971153d488d45aa56f2cd1d0caedf25fafcee9e955460a62b
zf142b22dc3b2634f6480d3bd22795a431d687ce10fc2ee9a15afb7ad36690ac3d92142ee895341
zf1fe0bf8c32b1aee090d866931d80e62fb7f3febdc34c3d8d6653a2ca234ecdaabff787116b7e7
zc4c5feed760f5020c8865bb76613e5c9d4a3cc76013691e74019b93177e2747587429100490bb1
ze4ac2da2c578541218bdf2eb4d1616f601a1f56a980b37983ff1dd7faa702827e018b74402f2a6
zefdb869ef60fea6a50d1cbdef2a8969deb1cf37d756f2c33883a29fa85e37ecce3417ac723c2ef
zb2594ae051c6d37f169a7ad2c57360fd7f7ad9c48b048d7e06582663b2b9b4a951af211866ea92
zac506064e15c62439c19ccdf7a6526655c45f82466190f31ca6ea27263643dad3497f69fc5fd57
z03f0ce53e805de01cce1b5dac3d6fc4e56e4e1ecf70c74e4ffcf84318673a5e9a38bd7855c63d3
z0307373050142d13ae2a2e26a9abc16e7641af9628bfa892b346303b1e39e862a19067917d6861
z193bab79aa1c29c5da8cf54944b8116db2e8c320fa8f526f6031b5b810cd25830b4ddfeb0cfffc
zeb4b2e6e9ee908b5d2d2378955c00c8b801c9f5098eb72377c424c6e2586fd66a2468ec21ad27e
z144c07b5385606fe2a96ceec04b551fc161aef47004f9e71a54e92965db05d646992a34557c4d2
z4080328b085e992f13a9c35cfdd8d50e7d30a9bded444a81ff3c050ad1c5a53241d0445bd93550
z167108dba5f2ae5a3a6e757b332b9b9339f6ed56724fbd727450f6325d5201a507ed447c59d9c4
z3bf04a224300949dd8d7142783a371e44896a5236107142e31b44448f61e9a7fcdf4f6b448b116
zc1901b9b6fd7e606575b20f747ea254eea321fba0504cd1141a517336db5f52ceb571638123754
z77e9f22e2d76135135bf9b58e3235a53f5d3d194ed5bb8cc6025768b81d323688e9847f955c2ca
z9682ad685fda0e65d7e13117de48515e1aa910ceb9e93310a19d365083a2c89968498e1d92ac91
z92bfe306c7475ee06e2d06f99e3f95a3d30adcb5b3eb2e5b3a2e4659af6a2cb5908fb098db8aff
zd265bf3f11725086ffbd53a93b5b3b76653fb3a29aa4fbe39e6a0d21eec9adfdaf7d590a8db62f
z5ae0309f8e046768a3325d3f33ef9dfcd881af9c02ac627bcc3de4ae14c041d10a4e216f27b70b
zdf5baee8dba195996e1a5125d08887b73424776ae95dcddbcce41e95266c4de25656a5cdf14541
zd2c74541ff06608c487623544a205bb56835d9780554da6cb32f003fcfca5c344785eefbede112
za564fcc5b4f3bc68096e83c8c08c7fc508f40035322bb6bbdd612fd7d0303e7e0961430c5edc6c
z63ae532805c0c0364434f44e5797c05471da0803701fc13c42a5e1084b0b3b331179c6393ec69d
z2faa66cf2e2b8bc58d4e2da507be347d8aa1f906501a3e9629e26a7e0b04c4ad7f373be3498d00
zf69748cdbdf1fc948afa1a1e7bef9a72dfd4a65693ad7f82bd422673a68556c3be8938d64a3cbe
z779b2cebd0b385e248fb0919f3b8e3e9454c581c0c661d06b4a3723ec2a06efd6b062a7a848128
z4edac30b91985281bb8321695ef35c24bd023ce30c31a7df6c0d2416fcad481c4b58cf636cbcb4
zea8fdb2c44c0dbfafac23e057ff3069d421f8fd7f0c6a99d0976be787aceb83a78956f2c02e545
z3baacbd5fcec7f1a74b37a2ded8103f612f8a49af8ac0d9c41301da59842de976d6f691b1a692b
z4a7752390000e6b70a150dba8ff77c914eb1fd89868c3c258a2b4d39ba11bc9dc74f88a0776e73
zcc61a7efc7ff9e80e5fc2544ff3235d137f28886ef616b3265c382c328688339162ecc1cec6f7d
ze4aeb9c73b040fac28559eab3fefed677ce6b741d8bebfaea55479e753a6d75c3a58690c4924c6
z80949e3cf6fa8b43f145d7b83266953098ba070317d3f48ae6254aa9d694e36210d2b7c5fe8f77
zcf264a9db7c77ad0bfed3cbaeb1c11cc582bc44950b324928347ad30f4826e4c3dfe793e692537
z3682c68380df32a068cfe350180f27bfeb5b1251da412880c30c2c28b985da6de6141d0e2bc174
za458ac4d1921708841ac5c013969b399f5b4ab8b4d491da117e16e58bcd6586ea52de40ca46e2c
z0684e8f9a51ab30dedd740887d86516b4625ead7c0ef207ebeec870d8d1a26d02901d249c146a9
z7da4150f9535b862289e9c8b19348b5e2a79b8b58ffc76fd51d9f521a411bc0a2282de0b138d42
z817c5f1f9b6721f115ead088d5c157518a9589e539b0e45683f29d49ae24ac808c1494ee6307c9
zc13f6c6a6c130f6301c447ad554b90fc6f214a9a7dbf0745014f8d1c9fbc10133917089a5806d9
z5bbb68ccf81d909ad35481356ab9ad62f0f6036be77b6df34fc0dcebc1d3b4cc43bbb8ca766f1b
z6ee90d0e754163c0132e113e87e262a5bbd7801e33f524af3a14ad32441d667a4804a144d8453b
zd983c7023ae069dbc1dfc479904ccdd57583bf09d37ebf9a0f499b6a0f8ff1b5441f5476582950
z289f1407166ce98bd8efb0f291ad0d93c082bfd557c36d32f42d2d2499b400e467da83d865bee0
z045ef593156d15afae7de12f50829edddb3cfd84bef9bedb7b62ae9f37197f9a2cefee157532db
z4700e1604c5fbfbeb4eba69fa8c34d9ebcf3905c539a1fd731259b2bdcf3dc2525579aac70c65e
zb73e0708c354b935308315057a4f34b1d75e6e9778ac731c4cc6757bd38e6bc6cb6b969f5ef839
ze4cf41c520edaa48db0ebbbe1452439060e58778034e1e1d4988004cda7e1dcfc650559cd6b507
zc4f043ffc7ecb34ef50ea53e2ea0809a3ff5308e03c41b85e69a0c947a4da968ff0c80964a691c
z4342cd00c4608bec75ba61229269e72085d2fb7efa83284ca1595fa0b688d0724b96b76018431e
zda246b37754905d4ae8e37d846704cd4a2e7cec7dcf8b8d3c190a3e43106b29da57e8bd3070d85
z88f2358925b134ffba759e424113d9e19857cfa98ac845c15b93963e1352abe8732513c7b88205
za6eb1443073c30953fea519c5c48eb90b0da8d14a0dce95df2a27cf62a5c87c89a0361a8eda631
zb3f0c170fabc2ebbb72ac0d1855ca8e94f301cf186ce2d53e56cd8444dcd7cf58121cd7109110a
zab114fa367b1f75d1550cbbd0876683f58ff32912ecf6a4664b9a6f21ff26af90ad0c2138ee4f7
z0ce38b04e12dcb100f7bbe003528643ebb80a2052dcdf1864843a5c94488eef33d2ad4d1cdaf95
z381a24fdbe56f28a634fd75e7fa96a68aa0b01c77f6374758967639ccfff05fc6fbe831eb7243b
z07fd5754b7f87b6a550193f376399f75147f9cc3239474224ab3b4bbb836b8641042bb334e0841
zf19c5a92a46fe7b119cdc33978f16652c83e9ca1b4a5b15a029c5afd6c353fc0d89edeff1eb8ba
z90e985354cb861268e7369ec110636b53f3dc46815b9b8a2f669217c8b8d2a2140849e53f3c759
z3219025b635e02e7b6a616bab78071bdde946fe7023963df718ebfc7f08802bb6e10c9035fcec8
z1219366ca2a25d2dd469cad75a9191f29cdd4f96b7d07b945edc8ad7d96fd29a18d615a9863727
z20e6a03a3422f104247b8d1ca200d2d288952d879d0618a1548ee44712f00ce84bb6738657df52
zdf582eab3dd63b3f7d4c8eec3cb8526e75a6394bcf66c0a91de28d821b56fbe038358f774de412
z0c20e0e9a80bd667e9218f21b8a4e539ea599f555607c4930d4c81134d48d2f3ee587d82352a5d
ze9290a027610bb4965b66cd9c5345a53b9e1defbdeca84c8d1cfc840e6c1b78e808ea7e8388994
zd0f8f0a6a2a1cbe269bd5d5e36407221c41dae5893dff5c7dc76ae0becc425d1bccc9054c226a0
zbc4cf6eac019d652ff9a5f4fe55fa52f518ca6cedaf583afb485828b17d317d7afb45a92c43764
zc0fe014cd44374d9ce64d3f771744d51d9350a1c40c46ea11309c59dad0549d8a0e7739a6a536e
z4414ab3edeab7da3a8518baa7d543c99aa69e32bda252ea39ff2bd516f5e57605d02d195a36764
za18b98b2066b25339a45663172a9b24933a40e4bce41b1fb6d4c309fff50372312db902b802c31
z0ca70e0765a3f3702496f9d4ac877bbb5830497ca8739547dd6180bf8b5efe75dd22b9d19fbc17
z56450fd156ce803150f0cb9632bea01686910670f49bfe8e0f1d1b4ce69cae0904b7e522bc3539
z46fd26ac9c23242923023d58a6fd1deaf9c093e8c0e1c6efd9f017e208ca5bb2f0c81521a3fcec
zf22222361082cfac34c959258fe5e382bf627c551588c2f8edd305f1fc261e3b21b0d57555a70d
ze6567cf29b28c6a5a1cbe7e49aa162c151a179439b4827809b1f37122de38e49a9e77450afc031
z88ed78b1c0a0c0b28549b2a6fbb333ceabf75a522a51dca713dccd0bdce5dd2c81cb17252909c8
zbc0fb4a60cfba63cacfe9100bbf2d629a59766d76e553ed3be52c230a9e185b47bffbbca361e4f
zd986b22cabc4d365e05af1d55b0a9ce969c3b02636b8aa15a295a39bc9a42df56676f215ddf2ce
z47717082133498ec49d5503c89b67a20da4deb7081ad53d10662f69434e0fb816187450669161b
z769a1786291f13dc620b8df72168c4a6b253db7cc174f5e134dd729ed140dca3a5ad572aa3b6bc
zbb45107f1789c64c84641117ceb470a8a07d77d0485e784608994c908531760a7653a2ff06ce27
z393684ea52197cab1ca19bf4d073a31c90676795d68e589612eef6a8bbb28410a4f41ffd5a709e
z96a539a83afd07d3e553134cf31ef746d13c51294fe04c14762b71d35bb64464f399251c426477
z6d7cafa25866b80f5054a2a5cd2d75953b7da6099affb0e389bf8673a82beebc61bfba0a7fb83e
zf1b63ff575bad74ba82dbd76ca6bcdacf41c83917a7a5ee30e36d04c9c14b758845e7f498e8d0d
zda9c880f4d27a20d52d9a5c6a35e391a9d8456eb4f9a562a9b78dd264c54956e8e4a4cad92d3f8
zf56c5578731bee14d6ae440d08eb324860adc11cc39ad432e60a3d0aaa5692df9bbc97999e5a22
z6ff77e568be667c995276547c68f767f0a5c90383bd58728254fe73273b5899218c94fc8214baa
z70e185242f0570685314b071c0818bf7b17b187231813eabebcd03c511e661b9d7b85a97a9e332
zb583820aadbfb5dd5196b60675ae670b6ff85f5140f84bf1cb78f571826efccbf759c1a9618fa4
z007de98f603b420a19134ed3f15e41777fe3222778fbf63d36b42eb3cc412acd39afd53b442b38
z7f1ba0a939c29056f692718983bba509b059edaa30192df1e696d7811622ba417b566db0ebae4b
zfef15a6e3109ea95181e6efeaf32a74583231b6d4695575c032e94040dbe9761b67b6cf9c25dc4
z168abf06e6240f8e7f82a2c50f6f6e8c204c72223f885f7597489f8457d5e51ddd605f45eb39e8
zcb16397ec3e7cee01327f983dedc98de79b3aee05e9de1ff575a9f0119830eb4213062cadd88e8
zc329681d2985f88f888e92dac6955db5809c988443290903fde9b75ebed116a572c1fcc97afd4c
zf8345e2a6fa62de4697db1115f5e3033135c1b99189fddeede0a194b10b6f2801aca1fdd4aa675
z548f612ccee2354be83363459230b6006a6913a624c2931c846cb736de6d05f3b207bf7ace3562
zece33bdb44f7d222995a7bf0597679898ac48fb1269377a7cb5414cc3faeb290e52bd114ec775b
z2cd6084f6f56551183d6fe4eae72fb56adc25d8fce0f96f8265a660487faccab04a0d5c6b12915
za76a793455a8acdecd8cad929311ce4ade1b5afd22c6e1b791ef7ff2fcd7efd292623fd4d9b651
z8e083203714652c20ee036f1722f4ae7701928b25d62293af69ecfca29c728285c79520d2ef708
zebda0d5a839bd0bc6c4ba697e348d339324fa120b794894cb8a8496afcda3baef611f5bbc598d8
z2e94c39eb406b2076667e977ac5f2b2f5f2eb3e19d9c54cd9c38b497015fac75aca087308ddfe9
z6a09384baf8f414c310d919dd5b4bd1f531af1a4de8f2568500b04711cf8f510c3310d7dda9275
z394f9ba595df7c19cc5fd5ac74a4dbdbade0f51b823062f2dcdc145c589ff09d3320b8db49507b
z5bd4fd0aa7706fa092b670311a225b8cc72257b924688a010888676be15ab65b61a65cbaa0c921
z6bec64d7a855165f331f222ac0d0d3d62304f30924cefedbda1ce6b7a775ff4f954472d627c106
z86c112e5c1adc909cd22b4028c0ae4cf7002381e0baa306e10c05f2746e1e02464132afebd63e8
z6fec089428a4a2ededaa7c1c816fe7a9632a9f0a1dc1ce0aebd0bc6f832956a947d8b287941758
z80f59721d9755302d325cde3ce6d670a638abddb624ffca291ea6a1c20610f54e4e6ce2226a6a8
z9d90195493a85a89e36dbff865fb1311320dba9db7744cd47dc0e98c0d7f910db4ad6bf6ed0b55
z593fde92d8a5ec00837c7a766b2c18158551558854a8cf98233d1489a04f8e5877424c1c6f772c
z808b09cb4bcb6916055f46fde148135f89c5d18ef8e6afb9f1742df5732d859cfb8da5fd41aef4
z6c742cbfe65ff76d2856fbcf113ace6385eb0233906d53d26a9948a5da3c6295dbf4db46f5d9dd
z17aab6de01c20e368cbe37d08091ccd68ede168ed7d1b3a92eab42520a4333fe5bc5e2a6d6a487
z5d182923284f20362d185b632d19a580f2067b6c108fab890c02e8c69e34793508c54892613210
z55eb97982f6b450a3ff045e1d2b9ad9187fc8d2fe46df1dbfa88c782f22c62ff187ded70e171f2
ze07db5d457c8951a50485edf8a170778e94e6de5fe05cfb55e7b01838656598901854e4e7b6245
z1bad3ff43529bee1edf859dafed1bc1d3cddfbfcdd7b6a10c5c9aa2cfe730016517eb890884ce9
zd2f9f0b8ece623f8d408ebf355e57f743a156e49a633b0a710bc5260a914e35a7402ea887e9c8b
z4793a2461669be0f87b8626d4c4f0fc86bf629df4f46e9e3a3d2c9f0ba524e55d3d9c2ced11e51
zcfedacda8dbe884331db971ae653b077ab86de0dcb867cc539e4de35c8b262841c37c2c9c2eb23
z25ee41fa39ad4d950d4c155348ce00882291d13470d1d177514ee53d34e1c39a3b1c68f6a7a121
zaf49e2a6bfbd8a0a0ade41d36cff93225dc93d67ddea7b09e515ab0ed32df310516c5b60e611cc
zb7b93379c9da51d7a5b8c928c17ec0d0062af8340b5d897aa46036605d675d2c34fac7467594b7
z41e654ccdefd171251104c88172ed7f79001abdd56aba5387552c4defaf2334178cb7ab2b8e655
zd1e60e9abcb9e0b5119b16eb520d4b717f6c8f06ba565a7d2594b84c8e27f2cff283c7b407e149
z3f1085f1a9dd6e86824b0f4061a346cf9a31f1e96a806f0188f5009f28be2e6b7c7311c625f05c
zb3ed97462729c34e0d2370899a268ae01ebba4ab9234e6f7f855eca8555cee475c7804ba707937
zbab4d0a91bb17a6db3fe9c4155d76d3f440adcb2cde540992a94ed3a594d958af44f8592a2f751
zcd105108a2f59bad486fc51bc4e509ea58df0abc93979e23e5b3f88f4a1cedf3855d45d10ddabd
z582f3dcef57441eba8ec4a0f93855fbbd44e3ab7ab07023709a27dd1150461a284051406a48f45
z68ce76001735c667552a941fc99b1df804e2b60e280d066244aac84439f61321416d3230f06c38
z70a75f144bb12c50a38b41d06d28bca46b00c0e31153cdb813d5d1de524dc0566e2bb4b43bb45d
z0b7b716f5ee1529a952adc90c7a2ad8a9a9226909199cf1bce42c022dd7ac2848283477884f0b5
z62fef55a0d2f04e88490c745f98e8796554714f2a2a369194c428a9773649bb39417ddb14c5a9e
zc9ff9f57835bce649f4950a625a29027725586e8137de64a025180cc21053f2a0d3fbc1a3628b5
zeed795eec25742106f55d436d54e59c9cb828cdaa377febeec09295151c15106b6e48f4b002aef
ze2cdb56a4c5f543a2d715a3e35cc7c5e00aca720966358fbe16a9d048332a6a176e9f270449bca
zfba718d6558091d07bf8c50a309f467e5f98095be739937c8bc809fe7891951f20dd7435102390
z2efa401799888f925c57d65c2c00765396ca16f08dee1a518e78f1bb41e625bea175ac6ea85f95
za15e9fc05dedb8033411b4f089c642c8666e3cac5ceda74d69a2bd91b5eb999bad28de392133f0
z4e5a40ad83327431e7bfb2ac01610d05c97129f635c39a21aba256cc3b5f6ff7ad600f4a9e5242
z77b58163db3ef7f990e35d1c609d1501474921253b2a4b7aa7271eb5c8737aeff3847079805cda
zcde5a79736ca0431c5662a7f33fe080b9dbcfe54d67eba4e70cf759f860176ee9b5d9e20a18042
zb6e41de5594ebf3453eaa5f14d38a3ccf507525275ed2ff4f2c283d2cbc02055923c412c017b33
zb54d67cf781300fede33151c031933cbf7eb43185f5f5947bebc76c9a44c3d7788b5bd332afae1
zc67502f378b7383a6ba8e2901955867db98a5cd5da5f654a020c88fee36118605df8f8594f578f
z219ec654ae37ddb74f7e5dc71b0aa598bad19777f783a66cf61e578316c4ce69f228f9766f160a
z5fb347d016ec564f195d830175b14fecd6d0ec2cea34ef0d1941b04284457501e7ab6ef2bdc6e3
zba0ebbcf3241c9da0111863e10dae58f22461c292d9ab9c310d4f86ea6b427614f639016573101
zc716abb4bd2f8858b52e2425109d71575b029d586dc2f221f6e5e8b90384cc82eb0f1bf7d6e5c3
ze7148d8dbf44c3de80bafa03d16f8201b86ab851d189e872e5db5f187e8ad013a75de402dde2b8
z7e5be3d4fda4012a3281a0fd8588cb388729a3a9d3c927648c2acff40006c2ea22921b1f290a7e
zbe10da907a61527365b80c2b796c5d866d9d91c326d821939ab7b13832e8a7be84c16cffde9a08
za5d2b5c094dbe3a30d00bf1944e66bc73d8f65989ad73092be09a9a627ce17e03eb7633a62757d
z4b38601cd8fd71ce13e10263f46ea7b4c2fdaaf2b6c858ea61dfa0904eb84a1d868105c49bf568
z306a589dfd2e7c1ff9eeb6f3c405fcef110a8b8a1ddafc864b47e9bc3e6b9ce1a2dc60d3cda82e
zcaf35f2ce18cf3a6b36458c9b62b54db1b90adaf1005f10e0d3b1938da17e83d11f1828ec8eb7d
z948138c67da5ba239f662f9787e398738a64a178ebb854d4c6d1e38adce0911187f0b48e07af35
zad89e172175f1565de1abca1a8041c2c192f928f9ae0f84e25ab741631e8be0271bab2320661c5
zba4bb02aa87f02a6ca94026b6216dd0c905120a0025264b4e8bf9972cf3fe77fa792b2ffe7f9b6
ze333cdf6b610b929d40b08afcdafe24e678608046861d2d1a0aaff9eb547403468d92bb66012c2
z1c2f5bb7028d6304ea2bf3b98fec639afe5e6157d6552ee767a350c311f4c88a24ba30f49fd106
zbb278eb00e85fff05ba0bfcd8b63a5fd2204592345ac890f032ebb9594a7315eb82ecc958d51fe
zb89e4022900bac014847dd8b8a15abe5a04cc917d9691f12a9fc9dc05b537e6eb1d52642226bf4
z6cecfc6c69409ce26e96a89627117bef46a5db6fa4e93da98ce9aff86257677a48a3a8797f579f
z0cafa77381f46c9c17487b6293814e4b4a2c0a62a5d72df6f3363edbc29136c4b5d58d5d452fb9
z1550eaecaecaf12c927923bd725cbae39b3405abc485132a2932a42dee1e2ca0483e26d404b9fa
z288ce4bfea3d06981be77e504757a69373ff08228b7b96dc73cb5543a0c32294173241e8b45f30
z5a11f41b1ff37a336a72c438eb2d1acf9da74555cdf0b883d36b1ea9acb0bb890a94e14df1c280
z86fa494842e5c3a0deb564ca0a4758e92d6d68e780b6ebe7fc973d44f5c1e896e6ade85f74462d
z41d0987a8361f4ce7d0bb737d4f03ba33a94e279be81edf8d1e8a563d05cd2cb76383dab1292ab
z93a6a20a679d3480da62d7b4f675dc267a9c904e814e61e3f93207e4497c33664ec15b95feac52
za82a53e0494dc7b10b1d892c4a1290d135ee814e24f0b3c3f496ba42fec00e1203390ef6cca905
z1278a3e9817c8933a73a3cb444a44bef28a0823ee5d737f86b49be0abfb9aca8b8dfad2995a5b1
z33992b18ad43b8b4739466e1df0d3b9cb98f6b7508db5deb71c09d9d9fb2112f99e30a7b6b3c18
zca8bf80ff8b89c923f89b8d9b2dec8609918dc9ee0dd571cd2d1e944496d9e3a9ddfff57cfd983
z7162b941ff04cadcf3cb92823ab2c00b4e09df07414af465376d7f63eb2231f820df35c81e1698
z9c2f924be76efd468563897d0afdebe21006e3b71949f31f9c1f6fe08065101627c6d2dba3771c
z0efd5c453732b146b8e94f36008e87132a86915b34179c5d5c9f5accf67628b7b0fb531a803885
ze954a1b2e011fceb3c4bce2aadee991a11b51f3a7eabfacdddaff63eec38693b250d619c829bc4
zec8eda81f084f6fd707012748fcd2f4eb7858c07cade7f9f12e03abf616bef6a941b11d2fa8791
z03bab697682786a7b8b91b37e9dd711b6367043c6c53818105b3c8099feef5e6eaabf0e3ffe059
zefc7fc3f5c176ae953c27df4c53e63c275c2be31b9d363b600cbacb107eb5c7ec85758b5337fcc
ze7dbb1f776642ce8fa86786830cba93387c193b17ac7982062d27f7270b6ff13b6d72183427fc9
za6eb8715e1a2227529005df27ef262cfb285216f7ceed83b5cbe54c86d64bd3d558682b39c0700
zbe523124275de45a04e4f63aa8ff91f77f66ea2ca6e88668476e2eee89faeadf3fe6b5072dd15a
ze6f71c5a703cfe2fc5216b591bc7fa007f01689bab9b46e61f186850338116da1bca11a575ead5
z3eecdb016d6425793eb2800ac5e04179973312d88ef6d74ebfeea088b358f51ba69ed42534e3d4
z5dfd3da1a97c2f601b4ab4c457abca68a1f143eaeb0ef9339a61d88f03037af4709f88c3fbac8b
z1b571adf8f880db38faa7c8a9b30032d804e5c2cc149c488aa12b27f20cad41cf4928965d5bc27
z8ef41bc9ab3fbe00eaf6e651a041379fa187ca3c8230138d041ff0100dc6bbb8ff4ee0ca003c27
z6799bb21f72c8e08a4b2a8d375a133278240ae04f0c93a40313f70e420a8d1471080a6da34ce15
ze6e1303fdcdc7f5934d9b871df011110eaf8fa8dbf71b3ed44733df07adb099089f5e92f09e6a4
zf43b5c338ef78764fa425778213fe2b575363a94ea06b27e5800fa3c4a035cda19f42d79b909d1
zb5772dca334749d162ae9c0fb288cacc856dcb2a805d6b1fe41329941cc4295eb83e79742d43cf
z5a79758e9c0a4765589261ab49e247297316d0c1dd5d727078b0cd8b4da0e2cb3faf079499bf34
zd9514408f8d30c207b98317b227cb6081b368eedf01f99f4881624853f1421c4c22a2812fc5204
z273a3ac30cc06ab11dc325bac0b32bc8f10c94a5f060680a0dee831cee0a09eacbe787e0f5475c
zd1ccdd3ce73fd2c0be57dae481b1cf13f70e2d735e2c94f608270b6df61d6b3d22697dbcff9faa
zebde279dc0292edade06bc9e9cd8d457eaf7f5830452edc9b2eff9b4c3815571f10b3f9650c49b
z1a377fc7c111c14d2bc7444c70fad78636176e9451228049f8fee27f7471a9fac8d8069c7feffe
zbc8d89bd819a73fcd80f2e836b2aa9891a3962cfd974af749b61335f19445f445fed11d4ffb519
z07a4a5857b5764e641c378de671fae9bef34ac2e701323fedb1f8162b8ffbb12bb350d82aaf50a
z0ea1955184e1210e882a84de8c5ad0ff21d18e359a1749b6fab630d90df445c1a91456f921512f
z6b83200accc1a3d971f8fa89793a797b3eb4e24c6b590b78ea363266ab39ece13677aa9f9327fa
zb365324cc674effb2d76051d8d5c5909b7ab8819cab199af280147e07462e9c5108a35d0eae071
ze09275464e8922071162f8b621cfa44c27d56d2aff2a507e61c607c60e3f30e0552f8d44c1e188
z5613c5b4f9a68b9fc19ebdfc01fc7b61f93c82c90ddce5a22747954b0a118469216a1a9b1d1694
z28e2c6b092979a052db7d6cedfe0f5beea01434c930a300934ff7398367e93168fd53c878340d6
z2ab4b6d442e8d8c49992fe56fc889d0930f8090590bc881d0d3b03c677c9946a40ae28fdd07b3b
z868d288fc8de64c276b341878d12765d3fddb0a26cc86338d060379256d5c062e937de9d0e3c75
z189e2e896952fcbae461c93fa135e84a9fd170f5517db546d3e1cf6dbeee11ce33fe36aa120bd8
z4150a93df0210353f0059e9ad5747ec87e94b3d15a6d26141ab6b274eef6b42513955fcd46b1ea
z2d47b5ede92c625a7a29835690db62cad70d6527e9758cca2d1eb07ae0f1d5ac2d793aaeb2b559
zb3629e628eaba4832af596a7875fda324b3e5bf2d1c062c0d2314fb532ded69e84a7cd77f06bb9
zdec021b406b7f394a52810f7e3d1f0ccc8164dc01b71d5e6e9a5fcc94e580888688fe6ba37aaa0
z9e1a5a2152c09345c9953edfaf53287289f0510680a88c1ff04d14a4c318bd064e90dfb962e1ce
zcfb632b2aed2cf84ca2456b5c1ef29726defb18cc007939707fbc6e243f6bdc25def19b3661852
z40af86fe7c02699264fe4bdfe12e13e3e464d3ceeef5bb1a5a5d54fc3498dcd882e4cd44a27d03
z41e6625a815c440e2cc0729baad733b5d721eed79a264fe5ccb83f37140e05f402dfce02b8267c
z94df7f6125ad7aa473df77fd613ae48c1a7b634d8fcdf3f1ea6dce2dbd35314312b45b9d0ca5fc
zdb6783f3f67a2e966205e0007e05dc8599c08aa74ccdbbdbd62cf51bc2c8e3f0affe04c49dd0b1
zef27ec7766d0406e481fe08145543ff0196021008ea88d9aa0e38b9df4f1796e79a7bf82c81de0
z7c1b423d1fbd3f8c5f459d045210e82d601c2d00e617f702b6b0271cd1db5c28bc77d86d1d066d
zcc9e67e2eb8f4af7f4d7db78c0906978d311c9d42c42258275582b4b2fd554b5b0d38db75ec87b
zc32e996d4db548e9c19632dcf7f18b7e141c395b7f2a2777524ea27a6711c24461c6ed64a3a0a7
zb99437b30dc9d3ae742672104623f9e9b609a714bad20e874b13c2e6170f68ee002cb5d317d085
ze843873ec726c71d74929db51bf6ebf3027d1d8e878e5f6ee88b14be9e00049097499e0a2801c5
zad18cc9632b63b1acd2d1f776fc3ef7bfd8f86660ab063d8b380c454fdb7cb3033df77b07c28b8
z541ba6af41991b612efcd5f25d17dd6238196a36d1ed5c0c92debac63ccccce8b03487b255c16d
zc210336b025898f5097cbfdc091fca7dda3336e85a891ca8965fc137e4e5185301090901278974
z2435afca7048d9a853e8d1b89b51bea7169277a30523a5e850b49d22469f6d2c9cbaf4cb39af96
ze4a5feda3ee72b6cef74c53c78d1c041a8506a4860045b5c76571b480c24ce22dfe1d3750f2326
z8957bc371571494ae23a96d00e3d6b9d325650e26ee4e40f58cc427629e22af665119e24aa7609
z565de47ce56e863cf0c58abffdd4717119442809668c9c307d244b48b99b7353f146effa154ac0
z35f2f22fbb8bb1e1426ba9143cf50b0afd7baae5584ee64b1db2e31f2b74ee3c169d50b8a39e79
zf4369fe53358ae647fa358f68533d5834b0640bb48e3d20597b7c1f531716fd2b5364253a10bae
z5ed30dee71461c5ac53e712fb338b3195d3e3e9f61e1e5dce8c89b4547a395fac6574d576c00b2
z4e8e31dfbef2fb825088bc997063a471aa169ba437a7535fb19831aaf05958057bc1ed7593ea83
zb0c5206961ce3eb019b71e13f87ac48c5e4ce139c38b5103e7e34c5a0323365642bcb505257283
z2fabd3033c03586b9414e23efea341894a6566ed2f21377457d937aa1ae654a3dc5fc5c0eb1a5a
za2e1269ab8625fe56879590b51ce6f14675d65b54f3d7d6a367c87579d4eab253e8f2e82111498
z1cf2ab9372dc66c72ce8615ec333994651bb2af4bc5a68e98839666059fa1d69d1dc9c95fb44c1
z5115c5ff80c7419a2085fccdeedb2c22c4c9309cdd1f4774dc832e5e9008127fabca26b40526d4
z9b104c0e6dfa572fef4e7ccb2b858ce18ca6f0b38cdf58819fe9754941f470444061f638db3083
z0b9ae8c3dea46e1d23861d0881e9e0cb476f1e3eaa5659b48a9c9344d6deab897b414ee8b7498f
zde4597c91d954227801d3b3afd63e39456d9008d91e9d1c03f94cdf7900f984f6d779172514cfa
z3dc6bc8ad3333a500aa63c8cc48e9186b909350308ee7ef488a34dd7613e2fecb558dee9b46dcc
zbc2d49660dbf610dc7cfaca5e87c1cf3082fc689c4420ad7dee70175d2962c8800482bc524afa1
z8d9c2d71691accb7ba760eb07e0099103a49b5aafd2211cae44f984a391bb3e4aa72b82620454c
z3424223bd0bc00d04293195518ea40f59604842ac5243d81f8d3f6def3ae2f8b7ea876fa0ea9bc
zc09e09a393c546f452bc2d5e0d47b753a2a28a22c6cf7995b1661d5672a302b49343943421f3ad
za7110c5e1aa67c15ca854d6c9d116568dabd06b45fb5a119b25f1ca87a1d2b236317ba529da60c
zdd0c6d3ff6f9e7cc6fb95c37553b3163acfb7dd4c0ab8eb1240a8be0117cfc81b29d0727926010
z5df67e2c3ee84c28813baebce475f40bad316642b543b4fb3b2a525ffdb98a2e8297c2b5af93c0
z93c5f8f97dea144f159a92737f8d58de81cfc5f0dc002a986c91e7ffb1b08287e5632c8b953d0f
z64f54bb12562a7520290040c7e35a791f829b433583528f33f9dad7d8cfe251b5f36f0c16c3052
zabecbb41cd12f78d24f95d91b5043e10a29dfb462544692fa283dd6535ad513fc2aa5073fbcc5d
z8055fe6b6b7ae6bca9267120a372dedb7ba52a4d5406420f6e1c2c4d77bbfdc062a78643715032
z57dc16648acd52dd2da459d1789eaa496edfd5f299102329019227ea9be8f37a348200436faf9e
z2631ec146b8e63fafbbd3b47c3975c4f4d43a0c7598e0f8ac71f9dd066dd3475be43c8c3e8ba95
z8613567d1db02aa636ed925e860513cc0ae0b7306db9093451778c8d0e81a8dab13b2eeef19161
z7081b1e5964992aaf6412d581678b5c008c228d6e631504f23f783e2ca5744b5a7372a7f136b38
zf0b50caaa16b938b5ec283d3f990bdb0c525903ebe85849c9562dc9315dd00914dd9f703d25629
z18868c7333f7f802b1d61ebbafdeb26d51c78a54037350f1fdfb148782e50a3c93f9618e0ff317
z7883229ee29f94c807a320d27e39d8cc194379dcad6b26ca9ade0f81f0bead5fa0a699706ccdd7
z5e4e66e5022ed19354024319c0309f49bb2daea51924186578033f59dc7a7e1c1ddbb0dc63644c
z9c8132bd2e8ee2b3388620afdd4b626d852665c903f9e290b3c4ec0e34a4490cda4da301ccc440
z11866f23347b2fe7038e3557eacfeff91340f59b40eb78685d4d5a6303d8345b5f3682fe7d8583
z0d60511ca8cb3257fbdb7506797e8d59435c3bde5fe7a352b32e1dae1ca734a2104af7a7959c27
z34edf2ce60594bc36fd8cc09a02b00ac51f76eee8122233afc0df938d086377bb74bb11a76a3df
z86dab9e814f33488ae5db069c1bfedbe161ad9a2c774734e494e9c1df025c36551ff46c388beab
zd8853c89c67acdfcfb291033174c1ecbde72136321b1359acb5b91534943a35622d7191dbd73f8
z922eac9837bdc28f0cc017ca086c09d453230702c2a22c0b49e54b0bd4c9451733e990360e9e97
z2e70bd3d3a1d30d4edf625db96b7ba88a4dadabacceea612cbe89cafbc357e1f234cf598ff98e5
z5e65502aeb52bda0f24e5f7209b567c1ecbad73b7d397e9ed0495205271c2304d1eb0cc75163c1
z570862f5866ce8cc7e595d9a955e60cb41fb39ab0235e694fc005930964e80fe283b6e21e8c372
zbdc8198a3f28212bbec3f5ac11d1166d7944b4d99e3753543c2a731fafec4735309e44c52b7f6b
zb3966cf896d21fdc2beb9fdbccfc0f929d0f6c0d34eee511f69fbe2cf830b7b0b139f0e032bb4a
zf6dc5cb883bcce423232dc6b89572a7f5412580e0377ff255ac3342a87db4b241f02887d253076
za3a83b4eed2221ce03cd25978291b06e96c288527ebd118d89ec2867ecb20732ad6a0a62a69dd9
zb8cb1f9cc3e922723c2a6fad37aa9156033c8ab9ce41ae9130b52f63dd619d917f639f47ebf0ea
z8f2128c160b1db69545f37955a0a264e473d4f5b83f3997bc3fed1dbff6dfada07e0911b87f726
z3cbacc3cc85764752011b78822f642510f17db99d1bdd6d5246338d00d3c3fcfcc3cf73c67f706
zc8b03c3c7e3be106dd5cb03503e5c93afbde925a949f46f5102e522cfdb69a1a567106a5f8606f
za51b4b38da71337ac6cceefe51f555b25d4006abf0379019f0e12bd40ed406ee61acf3c8101342
z79f3f9bdcc5e43502ac179a85ef9aaf5fce8d8ba5a3ddcb4dc7926e65adc104dab56225e78ba1d
ze54e01ab888f439c8e9875a365522107fa0967ada30bc1c94d76e3783dab37c4ba56eb7c566aba
zfd595191fdb42064ecffdecac01c9756ee7f0da48d615018b02fd2244c01bf0827f290d7b1138e
ze1a61b93b33aebcb32c9f8749ea2f0002b97a4a1ffe3d0db086b0003284849dacd5efc1c7c9f9f
z71b63136e431a0708c39c06cc1fd858ea0f914aa12ada475417bedf3e02349149e675ac9b534a1
z2e44eafecba22c0ca3243f204eef19a002d9396c44b6c164076d6f75ebc6b1a1aab2d2685f1d56
z876ed82a51a71ccdf011f569230d6ae02202ad1fd60abf1c3cf2e6cb8e0d2711b32f83f0ef62fb
z63d668d064c3468b258e3696ce50fc191a4acfb1d3f1cf70a247b3c51221de60ab480760a5f5b4
z1ccfded7d359ba8d970428ba7237e353a4e52073455383f300d0904be3f59a07c5e56d694ffc89
z16870feb6c5245567a629ea6acbbd623bea1bc28951c97c9e1133ef610ecdb6202a2715636259b
z1a42e2f9c557b735223d0b3fd846f13357cbab0bdf604cc6bd0af14434c0f53d878aeb300be87a
z00ad2215dcc8987db03d4dbfcf814739d99072e7b79d7df9807a2308a70f3f535f27e1fcb8178d
zd66ccc0fb248b04aca38645b5b1c3a198372fd80b73cfc7d3264271540571ce7401ffec70dc176
z2b7e3b7a2168d875e3506e79f2c586cbb4ea1c68d889a7ca3781f85ea53c737a18815f9ceede32
z8e2d14f538e63a53c6ee3751f87ca2d97fffc91eb93f56d917b8421191f8e1747076b5d775a6c4
z1d6678388d52d2d42484488456058776a309ce00ef5900943673608a62ba047eeff1490c18f68d
z5b08a1a50ada19ad57b14b733830e3549c4ccfffc75d43da02dfe16969da31d94c5fdcc784f642
zfe6e04554014523567197a250263fe97ec5e617833e3f807749a235106fe6d4b2d980bea3029c0
z8fc10fa4eda833d1967a15ba27626a3362c7e3c3095352bc862df5db81bd6134258e9143a434f1
z53b3ee96d795b3d0808feeae633f2ff00119362a15ded6a8fdf977720a1b92cd22b51877b84fd5
z09acede6100f1e9e762ac5266017a115b6bde49842ad7a3ab3ff783555a6d45e35e757eea585ae
zfa02b5a43f7f172bd9ac309303f986403de5443926c19555e0cbcb83e485a48fee104f4e0a2a5f
z85ca1e5344cfea6cc78a9d18805889a174f3539d2bed8fd1f27c0b87a1b41377aba591106c856f
zed222a8860c9b6f5f2be0a00e24ab2561e367cbf9db39e2d80a56023790dd2a4a64c8d9d9d6fca
ze62e2bc0107949f5782f78d05fb78deb478fb13b2efbfa14b6450dd9333faa882008d7b76ae46f
z2ddb8b58129a9feddccf2b35e62c6775ad3e7d8e306c821c7ef23115f0dd36ca9419cd7dc643d0
zfcc7e0a7a86b0b495e6472139b398c25f2ff2fc37a20c6437c537897c4f742eb51e0abe5979982
za33eacff4694077ea456c8f6a9464b86c02bb0fbdaffbaed6dff275e88be4af74527f6f481ef41
z05c2639521b0d9f6ba43ed3132f44fcf9d67b79edc505372a7bd1e961aad39df4dfd626f5bb89a
za101cf5c38baa9b422aa4849e342c5da2b68daf8b3dba0be78d6ec189711327f5741fa399d293a
z266de5be19628308b837312593087907b4eb2a20d27e976477c1d43ea94c5d5fc3b7c316caa0ac
z48570fdd652f31fe6d7c60b9c860372476000539505aacbdaafd4a86d2377e7b3932efbe240d84
ze4a4ddcb8d09c3572dbea5ba05e3f042795d1fd5873b8ca008028d1ade1b502391095bf32ec8e3
zed609146d96dbbe64505e72cbfc1df51c08ad541c3d7a75377000f54bb826d3ff3c3c5d24dc4e6
zc046659e4a2c729cc9f77e43eb54c612ace737b6451b582adde90d3957c31abf775cf59eeab846
z9eab2c61b605d47b1b9c302353677cb0e28e1ebcd91320d8b20415dd9ef6a93ef15509450c6427
z14d49f4c34b8399cfe504a76173b91af8fd54f44ae11cb71c7202aa73109315663bfa89561b96c
z3bd41a9c0ffe598ff9a1a1edf7acd75026f1f61f6926b22ff88584325ccc263d49219996585bdb
z8100fe0860d7ddc739c3a376a0e437d00a218f5c04c48c3288079f966976ac35658cff9b83dc72
z20d31de696e5c49b26626f86ad4b36a725eb9d39a834b21fd6abf16fc95a538eb940eabbc86020
zcbf727ea190b1324ddb9242797e0d4de5312249e17d5c8905ea4002595da02f83a554064010e94
zb0f5648779f547ca7757602e42debba26e34db12829b7a894c0ba2bc5fae7ad66de7f4b847e83e
z121ee7d8c16ec33b3acbaf3a1d8d5072944b671390d4a0038e07f28962a9313d266bc465d84213
ze1c5b9ff97c1a9b9fbf06056a331a94253a764070e7278b5b9e8c709af6b759ad439460986d0d7
z54f9e564c76b6eaf1b8588ddff391e3618744df72cf3ecbde0e04cc45804dc536e66fbfb9d21b7
zf06512534d9e330dd129f8fb4083eaf1f61974eafe005335e548a0380d76c52cb3eb3d082dd673
z6fca95c4c432e75235ed075f8b1ae012d20068bc7465e01897b151582a2febd35eab94bd088ea3
z8ea9ff62e15d0eb85da3893d71d21626cd41143137321e306d0df43f5cac2ccbf4aea4181e64de
zed90d61ff77442a56c90671e5f2751f228608ea02a6fb8017b0aa4ebeee84cbadf887930f0ac22
z0c8fb26291b37cfb1d5db1d4114e9164be0312f3e030927fc951cff68a5c95e5ce481082bb0faf
zd67b83185aa48839a7af5da78ec16fba5f98921612bae390fdbd3af4d420c2c4d59875ef75a887
z557f7fee5b51b7dece346b2972b5eeb817726ba3193ab1588b50120f143adf91490a56eafcfbfc
zef85a4256460e76524e21ba240b53ac85851aa0a2112be38c3d7941b7465460f08935ff4f9bfd6
zd218811f732a470c421d3c5fdf109b1caf8072739cbf96bcd617926eba0dbbba0873ff5f10c732
zba73d773ed0266e5f1c76ed8cc95ff5034f9b085c5e045cc0bf42e2568710e1c52cce2348a3f7e
zd6719ed39ecd05152f0b5cd628f86ee7b20232bea9f6f0de14faa8ec2f7c24afa87dac48d59910
z80c06ffa555108cdcf2413956f1b58206b04efc547685ed95e23d97159b51e4fcb4ca185a7bdf1
z726594689d284922dba3ec0cae54b913e3b3b1c5b5633f877434ef21e9e7ac371495d9ad283722
z1c59564f25ceaa0cfd18bb9c991e054d90e1079796ac9b893ba2a2e8eb2112276613581eb0e24e
za20b04ea26e0ae2fc0dc9367e32a3d279533a6eeb8e4ac30cc5f8e26371b17a43782afc27e281e
z3a6c80d3ba1fd7b9254072762423f17dc41193cf6e451994b6de1e561f591f3809c77a242798f8
zf3f9084d0a9388cccb817acc9011f6dd4d3c42c36a6bb8cc6edd4d358f41c6b1d5aea4f489a87c
z1a79a4b60a220e1d061b271e26a37c9c54b10576ccedf02734fc429a5f1bc3d74a2efff329a0f6
zc67868316fd19c96ffab333fe9b7565d2157899f3112799977d6e5b15cb5678bb7da0300190e65
ze5bf7385858d6bac05563f6ea27efd923a78d65875e50ba34edc00080c1eb5c02cab0b4cd64fa3
za333332c7c58c67f9e213664002d726bba6c9cdadf559fdfd5a85b4e02ac269e1f713116996476
z33906a0b10f4992e582a725f8d568a24bd6818db20248f80c6b7fd2a6c5af27c86316ed2f26493
zde469c47ac0663102468fd515949a99968dfc301dd83ca437c38e62ee7a319ea9f4b5107ee0ccc
z1fee3fe8391c0d9076e4413d348e1ae4c745ed68225790a133870d8f5ce8870f0b779fe40fe5e6
z72047c4cade1472c008cf0fcce4ec9d199e783e5f533c50805f187e1cbc7f6f80d65c864b5cdba
z58e0829664366451c94f38b81d15ecdc75835d2486b8d2081cb3d71728aa7319968662666b7ce6
zdc788fc95c4df55efe08ba4c4eb277045dce3322845aaf78cd9e4a9991410261e75c76857a7196
z7c74e4adc9d4419c28e38035e902824132fa4628bb78c18fa10085a039b8824344e1f3c400187b
z05ec72028cc63401513c3824fe23732df47c80118d0c4d77a11a595464fb5ce14893fa3ac1846c
zbabed0a6a6237ee90c86d5ad3d70312b628179b360874e09a35fc401bc6aab14a927d9c584615e
zf653d79ad7a939b02278db87b7bfde5d55abaeffdda3eb89699ed54078825b4f8f4e774708a746
z7ed18cd0dc49e43770f14a55b6489ba5fe2fd6ec04bfc4bb9923797fe486142b9521919d4cd5ce
zce6c4ed5262533afccebd38be2af885fcf484d4a6f2a271838d35ba62eecd925300c40ba6219a7
z1eeac54af777214e7bfeb831a861ac03350aeba35c5ed94acd855d5cf1d6865a49935d41e1a6b4
z22dce76c30b4858e1d8f4633949ba9cd6837195d3a6d309738ae77c9f9061000617b9673e69dc8
zfc3e8070209a5acf79dd81aed07a1eaf7cf31d0acc65719c12d6e5d2ba71001c2a2dcf86378d93
z696c0715cd2a1af50c7ce1053f849d0f2cd127e38c8cf87032d0709067ad12a891976551652d7c
z9e3b5a35252b7f2209378e59440952277eac4f8b90cb16c84fb93fa0b7193e02ab53e7de383fef
z958c3829c0792882212ce6e6f28bf68604cb1b65ca9f04f3c8344e3f01f4e42f01499b1f938701
z62550d0b60b4bcba5d4d2c392caf9f60f902bd6e622c127d0c99e1e3f8162e3f5e72694777a91d
zfb6bb556baa4d48bac186bfe6f4865cb0beff2836d41aa34fee6b79d18f12a5e4b20e8f7b58a9b
z3278be6be3d2f3276cec6d58ab49a7a4de01d95156ab620cf85b1cc8c5edb5d7c72865dead0457
z90039870303257612a07434eb64af393db724010bd00085b01e144e49045ece9855ce8499c3fc1
z4a3abc1b341e25c1243138accd93c935f02f3632abf7826ef401c0b4144a4070e42596fb8d3575
z1cb8e2ab412d15a378ed9eb59c70e076c50966e6f61b217a2a4f41019bf1c752c9934d0c05cf4c
zc8c95d53b430510003e0f57e26aa3c452ef77a9ba96b8d0c1eee86e4fabd3294601b28cade92f9
zbdcd45544ecc6a4511a5f92fc3465c7c9d382d6c4034d7ed8c10ad8b7e68be22705df79a097729
zd617279924a0e77076ef319a8974deab914eab821140d56d46e409092311f13a8e8ca458dce59c
z7049ffc70f3803cac51c124c02f912d1a723261307925e0a675d2881228bfbaf1b75fc91681984
zaf17e93f179ea781859dd59a1e1ad476d1562baae39f97b0a041c27aaa6e7ab55f2554d1c85bb2
z26040e553db9ba81ff8d2b228b563eca6e219f9a86ec9a09f6343f9c7407765635a2b98b70acaf
zd4cc648f6a862250b9c54e2ab9833c638449ece966097fea47597741bf058af4bd73f585b8bae9
zb0f03c31af3664b4b0318489591d162e936ed3350276feafeff2f6dc2b61c723f4f139457fd3cc
zfbb7240fa2c7c6609ddd7413b8165e760147c5b2846c85ba9e842d515f0788faf2363db58bda99
zc7738234c0300e42b2f36865da7df839453dcb40393bbfc3a621b2f9cf9d1f694d4a89d32630c9
za0e899a5ab8e364767bc743f19f8d410309ae20732666d972411adce3ed0d164910863fc44c297
ze84e40232f31a95a6f233c82d0093d6af0c9f29c29c9d0827977fb860ed0ac05b6a6399f71e3ed
z39e19304b140e946474870a8af3b0d866a1832a1f9f5404898fa4d9d47bbd2d1cb71e438b4630e
z7843a8d4ec23a19922bd34179b927253eb4fa45715b039308899bbddce20dacd94bbb1789342be
z85cc728f6d3465ff25f59b1e5d926be30a3d48a7eceda23efcdc5740fbd5856cbc14933e26b224
z902487aaa2c33918f5d2a4f95eb34cdb43cd6008d12ed284af6297c39c71ccf78ba04405d0c7d3
z5f07ae09d9de2e1fbb1c10f8b4997f51c710824a90e93ea537d5db1eaec7df8da95b5b8c438caa
z8a5b0df66812fa472ae50b8238c9b108469316c01208399df34cb6ed883b3b6e0a218a6a911aa3
zee393470c13f683ce029e636170cd837e43bb872654a9e357b9a5f20a9c4262926db8b85e34b36
z835072a1fb02cdabea100bdb0702d54ce8c15a091c44363b7f2d22ca4cf365f4754ef84d88fae2
zef22592e668bf10c4d5bdda79ae5f7411bf2cd882d80180a9ee12c25f7452195212ae3a10d48e6
zc078b6723bb432712a368f1daa6f1c01d946856c7dab079b4bdea2ac296497b851b682a6261827
zcfbbeb01ed4ac2d5ce2e98bd13408d159b5fb1c540d3122a8634aefec156eab46c89b5b165a7db
zbb096537a8db9d8ed7a8c62854a32ffda9e59e4ac8e2fb88bcf7f4e6f6ed8b3a0caa89a8a5ae8b
z52d38c2b3cf4593804b028c7e3c70fff612ac5db1ec81f4b4768ac4977ba451f0584543257be05
z8389e97602e7b949de4241202b70c76c242b52600c485be1c0ec1ce583cbc4b128238f9aec50e6
z4b9cd3523658ca4ebe907a0d4caef3211a932f26b2da872a16344e95328f3faada1d4050d16e8d
zc03264ee5d95c402d740b4ea391a6d342c2d891503a3cfaa9d3f731a075895ef915c5c830c1ca1
zd0b3b16aed666322d80c9d7c26a3f6d086a66a6bf8b77bf81b6952e734afefc49d32eed68769a8
zc64e79214175834343e4b3602dff1a782ce23b9db8e131e5867b37ac7c1a194036e7c45629bdc6
z238dd21eaeaf889ace75fc7b554e766add69dc9b7372599ee386ee4f54d2d09463cbe45c5dbe8b
z4488d2549e74f4f2de097189b500af9c7b1bafa32284365e0a444ea3adafe3e936192c0d7a918a
z22fde55271c789fbb4dfab3c010b779bc8d228154465a8262c16581044390692ca308d1b26d48e
zf9e0638d1db2f2d82e3a788280a2c3db9a20eb6e01ac8d43d3d81bbe21a293b9b0a17c66116ae0
zb40404dc443e8c657a345b50900675b337443ce28af818ea1fcfa9264d8cf96b44cff3d1655765
z79f5e89fa2ea7ba5425bf25999afb5c12ed3351097fccfd89da240aec6d478391a38384aa36797
zf9bbf44bc77918c41315bae9ef9cba945219d0b4b2aec5b9a1ceefa3d4b26b53b54df3d924df11
z3fce36770f12c3f36130a2be80877ad3624ca5b14fe2e25d7d928c1d6dcf89a2fd76eeea75380f
z8e19c50c5f44d896ee0837d25807cd9fa243140871acd875991fe8d8d17cf6424790969f82a8f5
za87dcc0601fa4c6740836493a8affebfebd3cc8dffd6956e093f22664e7421747fb2e02e6784c0
zda4726fc7da6e20e338d22db32d3555725ccb3a232a78dfc51e8d3ab124ea85d9f249f6c9cf003
ze7adf505998a84ac3e5397fafb2b458db0afed5e55db00c399957b7a5d8c34c5a2e062d407c07a
z7964b30d9100bcacfacfdae64ac8bd3673c0c2aca7d85947e3f6eeaad99306eaa817f4b9ba1890
z7b634bf9ea006e971ad07f0a901c78b99b6eab6e620789a9df4ebf2ea839aa0afedc402c00d581
z73b172db843dc64b818ab7f3e5b8070c3862f53d191bf98124fe76f5ba0331fe69a72ccebb4bbf
z544aa2e67c9141e7af8f7ad1b63c2e9a8d5b54ca67d35d7412bf3d346c87cc34b38a1d632fcad2
z9fb715209f30867bf8677a8b37d5cb34e7a0dcbacfe6df36008984e9603da57a686e33ca6f4bad
z8c207d141fd040028561b1bf7acb0561af5a5be5c69b58ebe730932131bc584e7a2527caa34661
ze63620a005bb338fd68e6c78a1a0235f03d54739f98c7f52c843794dd7f9872740df096864567d
zbb46f186b82fcaca49f1e8a36a117ecea313ae50adbc85c6174bcd835697e8eac606bd3230e9c2
z4c51afd8848c73e365fdfcafab9e9a15e3077d9504641f07485bf0e71662a46cc45316b70170c7
z0b10d5a71d90632db3af64bc146952b3f20d4725bed7e64bef9f5a9a6fe78140503125583122ff
z99cd4e89fa1ddc661a166598f5b2fe0f72f34f7105f25108fdaed992d02174031d601968657b5e
z3dac9e79c0f9c94c4f2610422d72aa50c07f079d08046b6bfb528f423c140af2ee5dce0ea04978
za6ff2d10b0415500dd51d41f59fd8743fe6e004dbdec8c38ab02de9393fb57e9a5fc130aead942
zf6ead8a51e44dea8978b1187eb7abeb011b849f258e559ed3e417b9fbe849e0eb01234bc9c4854
z3f840ebb246f847b2450d5fb451a784cdcc031cf2160fb4e5368e9d34cc2739c135470bb127fe4
zf798e291d0b67cd8dfd52d62f2b5b7ed90a5ced8cb7927471bda9fbe929bbe6e92a7038ece7e1e
z98b934987256cf535b044939bc7cc870ac7bc543ebd02a7d26a20c1bb0543524264e49e4928ce1
za24f6c9843268b45ec361d966c76bf156db1b6bbb81b8ebd2603f6c5e240ef479ffa4ef630f597
z20864dd7fc48909a20a8fbd1acd2a51ba92d0a57ada398df96524c734e6cf1680ad64a3ba0df89
z73abf7122bbd7fa1e9ad010fb3ed3115e4a3c7e93792d7ecba0f791e1a761e6e0e794dfb168176
z6df9163ba96012b9a7dd660045a50edeb796394b93922897b063a940359f862cebe0ebea53feac
zc957604d04d6b639b04dafb1a208cacaa48e7359879ab7a583bc6fa1b7fd758de0f50f94a66799
z49dc3a9835e23fccde44bb01ee624a76923ad88e1724e77a54d2ccab7b67661e026458bafdb5f2
z32e3708b07a6524958083c2ef1ef78b3c185fc07ed3ea84b768c6d787710cfc0e1ed7f9d9eb3ff
z32f3587a371986695de02a48db1b07cb199e6946fe5c307a228667cd4c1f2842119f11b3169e80
z90f6b7da27e788970d0426594ae0d321454ebd0eddf3b6d2a0fa91e635f372194c9f2e13e9eb43
z9312325b206d7156723ceb569fdf581d14cdbf6cfae6072c0e2c5dfdbe9d31c287b28615a3a291
zaa96065d21ce2b17a70e95f84f281ab48ad3888ef839ba5b9fff921237b64dab6c4ef6bcf065c0
zd2c61806653c7c8071c48ec87924ce1eac10f768742d8e82e3fbd02e7a41a6b2bd05ae2a9761fe
z5f12fc4ae85a1af9df3f2ff36dde7c8c6f169d91c5741455ec35f4c1530d116a97c31ea4ff2304
zfd729638478fc0d070130eab44e5aaaeb7d5615099255cc016583219e70261ecac1125277fa95d
z4bc8455258a1ac5c363e7d54ded9b78e5457ec32d18c226603491086aee92a7619b3531f0aa063
zcdb67f0fbde26c6336202c94ca13cea841b502709a86c46b8c61487d3e1567264bb506b4130856
zc5735c00588d472b4c1d34204785ea180653725699afe5b8e997d4ef117a0b6ede0ab12615a46c
z854a3670e6b4122e287bcb08c575bd718e6a1e8adae506382a1bf4f6d7c6b16ec877cc14009905
zf5dcde0461251acaed98714576ac785cb61e403283bc3b62487b7e56746f722c2f59c78d5bf9a0
z034c2f5f3665ccc3b6a6fc73a8916e8b0c21c011c7dba9d8b8e1f0b9495f1ed791da4455a5a3ef
zb2b792d9f50cc1dd4434d5b2632a222667220ae9d40b213676bfb16e87a0edcab35d7bef506da9
z1860bec62ddfe67b01cf31c922010ea691baf347247256a1f9ad977de148a3703f2cfd30fa57f0
zee0856f0572b6b5210070e10741697d0e3855e0371b39403e47f4dbe96921f9af6293b098eb3a0
z623e690764b3a62ca09907b1427940479fcec14e6ad6391be7eb6e684623c092e2dfb1be2572f5
zc09fd4b64c9e26d7bf7160da456a06563f43b02d51e77e75e3a86598d88f61dd15c1ea193f4f47
z81f31d7368bb9c113f5ae2023489ba9b18b36a780cf4b5692284162f14ee6051322b3b47e3aa89
z7036dcefb67ac081eef16c63ae013dda17ef376b34719d170515ded2183de1be1e1cab0b98b451
z16b56c24e155726ec26ffd8e457d6cc778736a1f2224d9907c84e8814a611f1e186cdb782b2afd
z2bd10bcf2fee8deec7d84347fccf27b4a1059b7686373db6f1b2f848eaff05fc94c40e22ce8215
zc7c5865487fee1453ad0e1f7360b18d7464768c404662f7775648ae64a9f67f813ad37b9aabe5b
z7517c2759d730560ea3a36a9ba5cf3c0adbc084ccbf734cd4b6a02de4ac37eaccd951cb53261bc
zf7d63a569d27ff7c648c8d1431d5b4cb481ce74a5b77d49e5a4ec6325c87868895485c2a0ae774
z9f1911f00322de8d6a3cdd0a1d36b353ac35273371cf01f10fc8014ced7357c5f8a61a84429bf2
z4d1b492dabbc272cd8774de915e066ad4ace58865d4d9916523033f19b3ab33af41ecef19d25ed
zdfc10b76e737ef9d3794a1c820956b850712ad8ec30a0324767fe6100fd7b89fe50fbf68dd6410
zded9b7bb58095606eb3abc9783fdf57e8e08d7a37d1725978ad6d0bd0d13b61b83dd663ddd8d9e
z5d9f3aa25dfcc47ea9bc50a54603f4f36a3ea038989c47e5ab4569840832dcd6d404e31a0234b8
z2829d953e48c64b280db1fcf811c598d74614aa7b1c1d5a2fee89b6745b00ac97caa025d0a7ca4
z9af6cebe5d2ea89d46f6f4ec2cbebcd511b50c8c9f6e65dfa897cc3ecf222c4e52a073b93ac281
z0f6ec6eb5614963e374d07508a539c935145394df65b4575f84eac071d87df647e4386cfc238ff
z2e11975cfceece67fcb624566ddbcfd70cfd3d39a5afb62f9bac610a1cf690fa2e60a7e9b3c17a
zb559de04cd7669dcc2277413be16691e2c55b14aa64798f93a16464420d3798ec7161716e73b96
z4f7bcabd04e08a743207191b4fd1d0ae05291ebf98f92d5de5d4bfc24423926c33c0e6d7debcb4
z12bd3feeeb2c0d296e11a2e5748004bb9048bdfef8d02032525d84764bdca13a8b80b3b8b5011d
zedcaba740eed09afd763d3f6f89330b9ca25814b50368b5cc53de877bf6a57f67557a3a76e0928
z1fbb0135e1a649b3d53d1ca9235e4fe996542610af5bb6098b19aef0b87e52914804550a542c44
zf28181b4dbbcc6d28651f1af52f8827647ed66fedfa401ec99f62452d61cd1dd2c83ea4846e676
za9188d249b9a38c5f8c554f37ca0013e943ddb6427ee58c39a38cea75a5d3ea7906a5095dc83a3
za11ab3a378a9141bc1f17a478bab33aa531b6b770e05aa594be4b2f77bf0e65734d55c71a16604
z2079ceff06d0134ceb9ec1045e65113181b919953b9d8a864a8c3ccb686704d9a12e113b73c19e
zd8a49314e6994400e67f6ea92e3989bb959f5df53b52fa4506ebe0fbcdb0f03d19f905b494d9e7
z8f7e625e6b3bc2e4a5d30aeb456328d84c7e4973fcdc4514c56620585c90661da452acb58eb7d0
z852abc6da396bf6da3439e97d451da13808314faa805ee12ff62c93fd8a227f08495fb4e704def
za4750ec704ea989522fb6a15bc5c0401c067d8a34d0f30780c658644c3ab8ccc6fc17cc51ab602
z3e5d0b10ede1576137e822a7a17301f7df8b19809f7e3dcae79d277cedd8b5cc9cb8bedd0df7c3
z18910d4941e7e8885d0591fc7d21950efb96ece4ca5578e11e6fc1da312a630b45fa0209272c81
zcd76c7294a38a3a430dbaf594650eaaadf9dc53fd731130198bc7145c3a06826066222a1599f24
z57c9e93874b3d5c4222de03ee1304ed221fc0e2f843684d4e4d6dda5ef36824b2421a76d6a12f7
zb23376bd304587f79e9e7310aa55cd5bc280c8d06846bdc25aef57c08148bf9437a38d7474f0be
z79c2b67698d4d38bc5f8c3a3bf28c58049539e2ba91a378aa955487be3e714921a5a4d6d29c9cd
z979f898a297e7d141ab89a980dc4b85ac3b5c2be7a22f3f060260fc40f9126e69cb83054469742
z1a37fb9eeddeb4b56e83f359ac23fe6cb9c79a16c964a5c8fdeb6cbf819fd7ed947f0d8d3ffab1
z64a0f3e8239d2d151ee6431dd4a7dc85c93e7456f25ecf6d5603e61da8a92ef0c4dfd1ff7f3550
z595ba2d4cf6a8b935bc066242fcc536d3c9f5d9ae872026b4380cee68b469ea1a6a7661b1c343d
zabd9c665862279704d5fdc99654ad26b4c3af0edd2a2e240b106084d2ee4bba6ab2e0980ac395b
zebbf8e44258f071d8e224bd152215fd72fbe543325ad3b7c91a74fda746848680757ef3a10ba6f
zef48c0fa5d9940acf4bf597ab0564d63b0d1f8bd7354041032b354b8e026fa46e67b23bb51d846
z3a1edb2bd50f761bfc8a3207910ad87c7db41dc347e16a3c8ad750035c72040664b2e8cdecb728
z3aaeca3eb609d2e5188667e754a83c8d3a08f57dd6f5e49bfbd265003df3565ba3bb4664ae275c
zaa59f8f2328128c3e06451a4b60be267067884165eb2600da17c6ac7544d4bba8ea74e8d06635f
z5c8ab19a0c3e0460039650e63d16667518ff9840ef4437ed0a5b2f95478c3769cd045c9183a9ca
zf44fcab84e6713f143a777f8001038496c0a010b3cadcd64745aee4f959c65f9c9172b82f95eb4
zba3c9f94dddce4e30f5f87406ff8bb694ac6f5b653880fbc3458a15d8fea602998dbcbb58dbc5e
zcf643f5ebbcd51a4dff765c77c7685c2d0db0659a40bf07c717350798bb8582c74b630477c0d0e
z4adad3064f0a111b7f0565d76b04fb75b7d24e2a34614fc432e6d40839b428741e2433955d94dc
z3a8c4be37be9aa8a8b5e70b8e08be0818114866c53963087b794137645ef671da007f560aae05e
z60550df1aef8b7494a1c1c75fc9b31d347f6ed7143db661e5c9d15524241cd0938739528cc2812
z18dcbe6a07cb7d7a948631d9c203d0a53253dd151da0af164b38e055cf28900bf9062b1b5be7f7
z65909a062b83d65a3137b9d4cdd181f64fa0e8f90c05635599f44ed2d3c9f4b428f48655318d10
z6a3c99c873f9c8111efccd32206fdaf385fe8e4d24df6a0477dc4fb2a64ad632b6188702eee170
z06d7f70c1e60d0c89c550bc35046303d2d3c8bf34bb8bf45cefdf0bf1e1eaaa7d737c465f8413a
z40faa1a2f617a10d68273a8e5bc6648057b75a349794ec0cfff2d87450a8e2f1dbaf7222bdfb33
zc2d58922e363512d3885173c2414682fe1c0610a027d8ad70380bf20a91d9f9a2226b08b32fe57
z54d5fb97738bded90188706ec6a047463534a9d466e9549607c33f2ab61b18b1c922fd3a701b55
z613dadf55ee083830e692c3977f040b79d3f941d2fa5c227ddc7e43fc9563a2d1c62e8ee30d24c
z22d9b1acf3f8c9b96eec7fd2bec1bb181f2db6a3761e601e9f399d83ad598e3e3fc5595260433a
z0bc6b554058fcecf6976460b00a203a8351ec30f462f47e6cc4ab771dea5fdba3b082ddb6a89f0
zcef07b1fd36c1e5273defd7d15dd369f32d1257363afadbacb454890c0a19979110a376b387ff0
z14694a72c427d15bf0cd27e8279a30fbc41e2592316d1db89b07f32ecc0945f247c12085a4c338
zdf60f9dd4894752283cfa5c746a6e42dbd8d698b55f0595dbeb135214025972a5ba57e086dad14
z85966ebf5248365447d5636947b90e394e66db542ddca3de7ec37758029f502c41f5e2a539720c
z181663d0face40a11bfd46b74f7c594992201001f795150b8eacbf1c477ae2f5157215a76d2e01
zdb94630295c3ea44cc1f78df122c12983358a448cca9910d4e55bb871242f23f4f29cc4f74c260
z14fcfd7a019f240ea3227513e4dd4403899747b8fe250c9f0f480dbabfd53b8482ec811e942094
z2e83a9cb9ee5ad709ccf181e26ec30cd43e2df806181cdc3574964756c4cee827db83853ea0bc2
zbf1f126e6aecac41f4ac7a0737055c8621af44a17a568b87a4a313004cefe0cfc947822a7187be
z38d7c6be281640a36065399656d7390e6483b05f6d32be47213dc5641428206006a3de84b1d4f4
zbbfabcc2e043a65cfbf4e90c95d76c26eccbc14ffa6b14d4f1ff5fef6784f9a11f60bca57f13f4
z8554968ab223481c7e3161a89fae3a6def76c61bc9d48895e25c49404a9f1617ca1bbeb10bb704
zbfd2b35dd8314fba6b33b67506242d5ee2ec1a2a1a1dadb8a9090ace3a85034928e08794b3c035
zddf5f0d5537b2839279f236b371b2e9380b28c4bd3f2fc000f6f7d4bf9e71db9af217f9388c16a
z164535b10659141693e7b103cb0489a7f992682358bc6398a3075c79368f0ff23122d8c702e940
z9ef3aca31aa0d1c3b45ef2966e273561ba37ede99a6826471f44b27c97f180cf5c26e33701a5a5
zdcf77107999c72dc67837e5828f02f8bdab6f9a424ea0d65793e914352fd5952408e4739494d59
z8590767e151fd8266c35759c7fca9753f972fb9783cb5e987e10f9fcf3e75de89d35e162c1df78
zf20a123b58453dfea27ab252926d2f2de34c1e355e55e167fc59c9099388d9cfef7d6ba59e9eae
z18423c7d483a6416c69cba4a4683c2ba62d2765ff5177b06caca42711f298688ba7b4d157048c0
z1d62af58e659fa11e99fe163f1417c2173dcf1d701302781c29011eb8c37127f4e79bb7171cdfc
z68ae06f57fa2e35f3193ccbad39b8f8c44e2e57daa85cb408714b9efd8d7224a026f99e9d2a757
zb66198293f7836d6205b1247250a5cfdd329fccb061cba0ffdad01e4fe05f9804c3798324f9b3d
zbe10961e7ad38222d354c916e8070e17f73131ab5d3cada926e2467b462fc59760fc96a05ebbad
z87c54af0e9f82624797ce8565d9f34b77796c8dec2f916e6a5d4dbc62e3fe32125c0697e066168
z180ab1809a6b9077ea671dcfd5bc0714e9c184fea109bc0ea01a76fad196fa121320d84860edea
zd9db8dec75d8b8347ea3f2ab2e5bbb243f4bd8bca02392860d448ce52726694167788a71c55b00
zdadb679d8b5f981edd801ef383aeba50756d1aa532bde2cb21f54c0aa40f6df05a5e45818c59cb
za3750d48041ed0e6c4d613e139f87e5b89a73884cba3f89407e0d5418f972dc05acdd287d8ced7
z090544112d37dc87c3a71be124fb9fd0b5e38d039b54c39ff0cae7c6ff4e2e2f81004ab9ff6710
zfd75de767c119af47a7ec111d95d2bd634f92aabdfdbd5f5a2f0bec2de26af1b050974870e9fa0
z8264de211f8766aeeb991c9190c960e1bf4dfa38dece54f7334598826ab6e4fce2727717dee6c6
z50ccd6e301dce2f25092071fe770ce6ddcae1f0411a3d1ce2a11fccc0c096a792322715081f1dc
zdf780acece8d6c5e1403d61da765d7a2a6fa08964030d573d7b2ef31102f5af847615d8f82b387
z009b728164fb6a915e3bf66e0763d04b69f11188e069b4510c8fac10ccfc99c176001e1e7005b7
zdefd976561e668bc910fff9a2977deb0a9f9be011b12550e609f5e6d0cf9e29931a85c7dbc9df1
z1c9bf8e831c61c9b80c943caf93bf8691392384c513fd7d1e199e96659704cd98d4bccee861c0a
zd6c4cbba960995aeab8d22a277cd404439f91af74f5bd9a24b5ba01d8c50623f3da45e489a7c4c
z1e9aea7d03c575ce7bd3bc1e1318e40da978483854096bb507672d90916340cc13f5334e4d54f6
zd0ed68a51bd1dacc329270e81b91e84775eeac263185c7108c7b292e3f090a77cfbbed8cf072cf
zeb6dcf7f37d646ff61fd603c740d389fb392db0b0fe8a4fd699fbcab8acbc2c817ed312b1fc13c
z8329bbee71402bc59b9577ce2afeae6d07c3b2a85ec49581ed4564e6896c0e47d259c1e7a2cfb3
z051dbdc901a8d035ad6d514f9da08ac7157ca1151486f7f38724fb0e07852e993e45bc77cfc1be
z543249ea7650163ff6f2051941c389a4a753e6d50070c5183a5348c36fecc652c9b086e0f02088
z48ad992560d9f14bdaf05e161dabd4a90deeb4441e4eec9c92f45c44406ec6e6b2a3f562b61634
z0c25e0076be7094af53f207c21852bc5d1c8cfa0570b06f35a39e30cc8ec10d77230d6f38f1455
zfbdd8992f19841c5a131f9e326f097e984a0498c03672105e8aa05bb7908cf9c770cbdc918e341
zae282adddedc1f23cae7c30b3e3aaa5913aa139b02dae93bf5085d3d35228d892597233bea3c18
z2d514fe0c920efca9ed9960c7978c60cb94262244257a89fb4b5fc7c0d00b4d8954868c3a87897
zf64606ab44008cfc790060f85dc59dc9ad3a4c0e055c59d2a1666926b93d937afd3b4a5625d87e
zffdc22a373717fd4b54933e0ab83aa307b0b3b324f8ef35a83a7a2e162718561d853b523a43c27
z8b28beb2a51a872829e8ec2c2cce6357b52f7751b79aaee1a1b1720fac414fa8514c038eb9d75e
z86d1e2ae97b155ebfa6d4af61b89120d36311ee6f71a55f43f77c6f1167b15fe39f9f73c96c656
z4489c4792951278a147d19d537ab4294839f098116e51f188d81701f46e1f206dd2c10358e8bcf
zb3e1756178348335475838248e2ef54f7b8ecfdc3b744454296b74466f338b530f7b1edfccdc04
z00cd41ddd6b7984d32d0a607f6011131c8aa921cd29b39fd3c96da07e37612b2b9e3f3ba66f940
z6be373e27ac3028dacf87961bc039eee270180e8c2df6457c829f152964f96eeb535b1e3228381
z0f58bfbe1ab33c8b2517ed4c72728a195388c1b4f1177506b1f84aaab3e27f88fd1781d9d92543
z5168d0065642481bbbff29791892a1d2f24251cf4b2cfc767aa207a735408945a61d6506d22c89
z87608137e1554a190fc58c0968518ba91267b496ae54c68de394eab46aece85eb3076545c0d606
z756177c49ba0df2645d866ada1d7852ac70019735c5d753900ba0ef3679bdbeb442eb36859334a
z409d9099879ae1be26b4fef418a21f7be424feffb5fbf8d92534039d9aea63afbf0cc551821bc1
zf98d766bab89ec64d3d47e700b4a4ec8566a66aff7732b5d1902bdac1834209d47e42c38113330
z0c57b80ef17e7fd0b1101d8395416585ae99a5ab9aa895f79dfbd7890f08d80563309267e68b63
zf9d6a86e53db7c3fd7b430c2922589a2349a417b069700b652cebcd1683baea1adb8f9cef8a087
z0596d36fb2e41b1c039473beb3b1f6a00ccb9ac97418464121b3f44d4fcc3ff05750e06b48226e
z3cb706e77407cc3d51c05b8420c0736ba10ca50f82dd0eab358c5f79e5c86385356d7a7e4465c1
z789658de5e818121e2be115d3e5d23c0d4837fcf401b1bbb969d245167c41f517422a3852574f8
z415a5b086b52e749b45289efd5a366e2f09e83cb714a806be7c19856a8c5132f135ba8a9bb2770
z8d0c31e6853a3a274a9dea72261a9c3e44811c60677ff93e60028c2dacafea252efd49f68da58d
z29e5c788ae32d24ecae43ed0f9d3a3ab0225e932b403322fe7a2a94abcda4c4c4d170631792462
z89a05572cbb12c22193dcf6dee98ab477549129d84097622386aee5479b8a3d2c440ffae153f3b
z3b872082802f2a8bdfc2292feb192748b28f5dbb56802d237292b8c87527765b677200a688d2b4
za51316237eb3b9fa741ef6084f3c467ef9f69a678442082e208935a72c3eaf3951881e898dc3ec
ze3f3b342d43e5aac9f6ee206e9939f9c838c6e838687492b13c89e3862768f1092ef2f0fcd5701
z2b225e9e673bcae5c98a037955ea29325ee426170769b9781a1642df609bb949f717eba32ccfdb
zbeb8778059a67990e579982045cf4359dc62bff5b25811db1bdfc6443aa6ab7b1ae345918c7a37
zac7b3ea2eb15a9c209fbf9d316729db72e37e357e5cc454d1fa6a249da7556a3997405ed129f69
z8e700a41a0592b3d0017aadd35be5ce0b10a0d09b272299fd0927a4c35efffaca7bfc68963410d
z407b3b1ef254414fe0c893db5be1c9d9a5d6d02b568b07d230ece4fb7debd2be867f6e22512bcc
z20e3436635cc9ede1e16a1ca15287276933823f8c6f3a3fa74258ad04abe96e1e54803508d0283
z53691c8ac2c8ef72d707e2ae7e07b895ed303a9c56217a8c8d3c8f79cf8de8f9bf8fe89ceeedb0
z4dc0dac67b13e821335e35a38f7b25eceacf2028e0c5491ff97ef5e5e5765ddade4b3222ad289a
zc87c2bf9ad90ba93d9a36b9305e50b2ffecbc6b470447263559f7d0a1de75230ddc7f96510283a
z6852c54e12100db659e55dfd7ebb1eafa1b154bec92ee91332a456fc7976170d8756357b839781
ze3e7ec3f12677fe4d795234556ec308691cda01a6c903380d127857ecc3518b0b97fc55e75c0d7
za9f208f40e044bf13278bc31dc403501ec1daa310129ad779bb4dc1f0471f3794bf8ab620194b5
z180286d608160c757371abcba53273cf20bbe6ea3fdce955bf037b8f0a9994552096a043bbaf17
zbd478f2fae0d2587eede662a121400c06a2512ccaa14c073e1f5f34699433839cee704cab2a921
z72ea1866b366fd665b96b018a628786605ba5f023a21bd0da3caaf69e7fa346717bfa3defff8ca
z4b5451c55b8f4c66711e4cf5ba20cfa24bfdce7d826dbb31fc0433b747233003d18f831e2d557a
z3a736c67ce13687bebd90b9bf62cf17a1ed0f90c52b03ed3565014736e34ce7a9d7ba14a982e51
zdd995b8f57c9c1aca3cc6ccd6bd454de3ccf78b89c841ee4e32cd054181eca23386d083afb6fd8
z82d2cd6c0b2e6b52f6ad9500e71046bf548c1344d3a7a9595c523624049560f09f1d37ac983b40
z6601e763b732450cb1ee24e1c38bd6c5dda3fde67c1ae13c1180c813d7705b2cd9aca9253c4517
z07cfc1fb6e063b5e0dbccdc93e4e8999c034adde9a641a2ebce970163027f04a1c282b503ad075
z5bc985ecc8db8d1cccdc6f57b20d990b1438d6047e959b48ba796fdd093b2a0026d4168325f528
z62b2c194c577c4c5f212e376323081b0507f05af0c8d3be59b322276180320d44d6e600d0b26da
z5f581460f40bf9076a08e4ad23f2f5a265f9dc9f192924ac8858b535550e9df54ae74223e93bf2
z6f1bb9a5d431c6f757848ff0cd8203905afcdb3e3076fbf73ebb3ed94b01e828a777225163ecc2
zfbb36b2f00217fa50b54842333eebe3d9ed56d881353d8e73b4e2a63d3bac161ab328484b41b66
zb471c5a226d9b64f4b955f1e4c4402def7fa6c3708313b8b034b3ca53a319c9304eb73a09c9898
z57a91f63e5e2dd2db0242ca5c1603f739ed06341b0e1df4d6fc3a4b53978987b0317f5280b00f6
z754efd8e9f650c0e89a6952ed313c0d163e7be154084b1696130fb7c1e02a3780993d8c9b95566
z88848054e30279d9a544d626846e20f7a10aed5ffccee5baf49427c978c8701e5acd883956dae2
z1e3c103e01cf723b97c2eaa16d111d95364d477df7b45ba6cc96edfbae1904473ac7d3f3208106
za16d7d684828e077b2fcb809601352083869023a30178dab32d63423a0d25ad343d94b5b81b125
zefc92456beb1347b92990ff3423aafb4c12347491b6125610b90a0ea941e902b56b5725cfef0c3
z91d530ef7634ce9d19f493364c970b203a50d3b664d351f4da67349120d2b236ab69b7989c377c
z4dba95eeacfd26f72c8b478b6bee22ba58adb3ab9fcf2ed5da90bd9815904eaf8fd4a261225735
z28a99abef3555ee389f1304890802e2bc78441eacca702e77bd898bd6bc4b2d8c1cd9a4adce487
za3debdf587e1ffbdf1d9c3ec38d8e39563e202ad67f81f024ee186f6f55067b3d1507b9ebe4c1b
zc8455cb0aa0725f38af594b410fd182574fad225575afaac135ade63ba67fcc4cdd16b79b96549
zcc1a2611bd13e5f97e51a8e8862e2247a9578e1b562d613847452cae7ffdd77d8163b9cfd59ef8
zbb1f2c7331835e3654665f410b7eb5c281fe61d5775a0433b388f4c8504beeac1abedf6fc2af79
z84667434aa2165a0cce9f43a8deac4a967c36d833c783c71a5ea678bf44269dcc7032257091c71
z56a9d6ae3819bac2c70f2a2def745dab0df1ee201d4367c83214bc184327e921d9f8fe28315032
z73fb3f0264e24a3afac2cac1dd72d4e37a3841fdc5ad5dee460561701de01d302a1074578d46b2
z3f059571b62d6f2e9ae1fe2dabdc4010c40c1f6d9ad5f2cfce5349858bf0b05eea61a558004662
za8917cb883980f4095a37ff515999a0a951eed607caf9e155d1d2c388d55bdb8e05a4b4cd520e6
z2cd59bf862100a7d9ceb706158498b2c5e4222cafebf26863b315e4f0965b67d9850f7a6bb7f26
ze3534da3a1a0856b28ab045ebd979bdfedaa888bc1963839b5a54c36de7a2c67aeed84fcadd055
z76c4caba9b4a2f8fe9d09dc9ef598f63a4adf8f97e27631f3a311dc86e735dc911bbcebc1301c8
z4a241eca3916fad482179de48e395882ec844a7bf4dd578cea11bea785a7afe87eab030b89e007
z1307b5c3a6744018e96a1619451c20d2e96ae56b1f9e2e9f53b0ab40c32cc71e1b402dfec1d41e
z7cb5d10ab14f02a4dacc1e13a195a76e9d3baf63c63347ccb2debb96ea041a79f65c8a5604e6a1
z47783af62e7d3892816492e5974bbdb56ea3502f31aaf9e577b66cfdc6453def241fc9cf6e7d9a
z28b46ada886eebbed9ec59da2fff8cca5dbeb0f3c578ac80811be7f6160ed3fd84b79e286359b0
za11e6e7b11a47c119e0e22e028cac5ceded805ceb39d4ecc838df41f2f446ddac280a9e0e68f09
z2965a2ce94c1d5d352a74e12ccfb4ef21053fe6d85e84cd2b6f3749a7ba16a5547e4b2c54a0642
z68c318b84cd681d42fb2202c88aa52455fb6fdf33da237483ddb636377c065daf7ec5e7b570487
z180e9e7400c6385252731a6643489c4cf8c757e094f3ff344d00615efb94877c2ff68e28f85877
z2a64e16400a09eca2971df8b15328d282023d773e67c866b8e4a739ac02cdddbddc2c543975205
z55d905fe33b33401b9861d1673b4a1201f2e9ba4e90be6dc00b0e56901ce808604c91fb1cac899
z27dcf7ab084f426453bdbb02cda6ca473166f46e5c002143e26d5fcd76c5bcda838ceca8a37217
z67c4572e87109cc14a50b01aa0b962ee3532434c35bda5da1e92dd6d5ea4e7fe6493ce2d6bf29f
z3390e58b811ee8abea523e6c33d1e89156bdc61a4d202db2d7ec8aa0ea71521a9dd69fca695301
z78737ad0ec8dd3d4167e8ca3e6be9ea06d0bb3c2869d5bc43ab5a941bdc1f422159484fbedac53
z982b0497d5ae3d2021daac9fb2b3b409730adf06fb2b03f17abc49c35f2ad510571f2372bfc989
zc5e19247b898eb262689523a5006ebdf8c389033fe6a3399974826108c26ba464777e8e9237534
z00e63811618747d7b1de8cc57b58fee79545f80a6e5c0b4b4636f1d4a5e765c6eaa82076c3b67f
zc1ebacfc5e30666b67c890b8b33ff71660373d1b9641281165aba2c80ecaa3523833ea436bb4bd
z60148d13be5c802f1b5c52e37928d585c1f795db4ea893982ebe3010b8ef961e53dd85d206b423
zf6355d538c9a738420b72ffb4d785fa6a443bcc01ddc2df9a5a095f6a438cd95e4d9a51278b554
z0a2334f6940e4d0a912366208a343261bd8ea1d08fb0753b049a85b7e8fb2423038675f841e650
z4d16c112be00c775c2fcee66231ea87844bd2aa6513924794d36f81bc457dba5829f7a2302a34a
zd93ff4dd40dab80d4f5e91d9f3442b600d091feb03a687c83d074e7502786614a6b28120987fa2
z756ba762b693b0b8c5d09947bbfb3d409be03e0043c653f1589dd983f270a5eb06ff6c1dfad52f
zdd48c14cfb83d758cc15b6523c42cc08d22e6fe00203f94899a6c931552f9e1268fc7e3e12d2c0
z0e64f6b49a9a070b880fed01789396b799bc8d5c9f6d4a026b053e1202d7a585bffaca2be602f0
z517cbd6bb2e71cf9c5412dcac5ae503538a3c6b300b8126afc861c9f347bec393efacaaf0acb06
z9122b6319d14158c290051b2cf32665366869fbf1aca1ace44478fa70546fac5a109cec606a4e7
zaf95a24a2948b96224e08aa81978eae6dd38c6bab017b84c4a2c16c1ddf132d298729e2cd020a8
z068e238c70a3664918f74dbc44fe012d022502254526f20efcb35ad9cd092003f1e0f3f815074f
zaf552751f92bae8e78b509789a870987b59d96aea1aff432f740b5c3d501176c17df6432c06440
z14b45ab7b5256fce5412d8ff2ed64378cc8d227d69bd5677e17bac3dd5db0c16d81e8e5fb01bf2
z647373011167eb0f2ca8334070e2d37b7725ab6995398e02b6e43e03890317a7aabb48de356e46
z792cb018d6a11e4f3b0d85f8dde60ecc5073161caf2e938732386e7e2493f14ada6c3370fc5d87
z9acd5318bf03734e0855b6b8997a4fee7e709bc9039cf01f0a412485f51484777a4c24477e997d
z90e0eadd6f522c3bcbc4e24716c775a3690e08b8450a80600093281f5133d11fbee776c4681743
zcea1453cffd5bf592f303fe0a69d4febd4f563729a95fc8fe4efd4590cffcba0b497dfb1698a95
z8025bfa1f1cc9e15b7f6e0b9cc384837aa74393a1e99049233a8ccfd43e5ca0e84d302b752b49a
z9799a176d51d8d8a54e9c3c10811ec8ef9b94c569acf9ae491d604b4af8f71b0b5ce39cfaa3230
z658131b921f713d660da90f1218c140999a00a2a52ce477959e9ea7b5050c155feaabdac9e22b8
z7f5d3aba9646d4731595c8c484788658d44e918e2bbb6f1e439862c663c6d05e1e54c7dd0368de
zeb79f22f1c2e0d5d73ce68a9804c72ce0700675d6fd974244b484ad74103d53269a0edfeeafa00
z52bd8f13ff3a361ee8a8a2e7f9456186b25a2857ef816597f381e127288a5e9d0acb2697597d7d
z79f124901a294466f20c895ccc958c93a46821d961eefb1281cfaba64a28609d2fba6c6d5c201b
zb5110c37e8022a8d8beba6e7bed55cd884806c938d807675efc3b96c23aa8771c70930f23c960d
z40af5882ba56371bfde05d56d1db0c31724981fc8944c21c06653fe81afdc7b8ebaec042afb785
zff92df5a2353dd9dfaa51a52eb41835a4d6412661ae0e3dc7449bf72172d3363c35214bb117641
za46861dded5398b2ab69afb82c24dbdd2afc354ac8261b57641e9d0f4e4685437f7c75e7164aed
z18560194b64c998ccd8c731ed493cc3b205491dec0d1407fdb8df6abbff87ca2aa000a6dd77f34
zd04e40de44f4ac66be7f39a3aea49d6e29b8f7c44e4a546927941c8ca5d02bf211e9e239bc1a9d
z904fa6070efc2616bb810ca11cb37a59de2f5621882deb5d40ae51aa16f7a3c5f8b5ba4918fca9
zdb9d3509b39e541386a56c151039d7fbcd4f653f8070af87af8299bb0df08f58d93a094288350e
z466667fec515766d0bda5ac5b3ae3bd12d8e2cf6c9b491d7c1fbed430589127eb9871a470b1781
zcb8bd8f301f4cb57b0895b1f00044ebf6a9f39dfa818a8fb14ba167d112bf2bc745f3253651a6d
z847a462559bcad65c1146ca87521d20c7f4da16a14807de6878b9757b11fb292beb89676e7064c
z462a9cfb01f3d57c2defe490906eb3a9471ee6a0c5be8d980950c03583df6ae48323a640c01af6
zb76e13c8aff72856ca8d3c5a41ad18d278725c9c1804afb2e06ddb53ce384180b7f31471bb7b52
zf2c0cb0bd2b35eb838a15ceb5cccbe5e32f2c9e57b41b1c073f62d18a09e859f19cfe430f6fc42
z928f246a76bb881c2059b7eb26804f85156add041e4e10b38260d65b3c1bbf9fa81e5b2e3b5823
z5883e09ffacf0d4c846ff8a02900bae4bcccd3091840814b63c4daeb7faa29888f2e600b887017
zd86c2d2b681cc8c20391585d500954b96fed0cdb6cbed522db5ce945be6c63434148f6edbc4605
z0369f21dbd06fd63d8eb997aa54b4de4dedeba6f11f3efff7f6cd4c4780f5e69b4d6d26464967e
z797db5aca7ebffd44c21fa42058562c4ccc070a187dcbd4daa4e132fb293efdf4e07d2ac63b352
z8da926a61850146d04867e9c10519c2b6d60fed0c714397dce941c9f5393a9fafc4d71ec09945f
zb3a8bcc5b4616b074030749592229ab2740f847d821cf21b92b4f2ee1d2a7c517568eaabca2224
z789b873339156d28848e90c37b5cbd2d3fcf67f1c49aaf836035e0d79b007fd2e9d5c990edc53d
z5c9a35883f92476e0750ba59993c1b76e6dccf729dcadc2528de2f720de514229cd3ea3da5fd25
zb1253e793c68e1cda4b9daa7402d62727939bc01bcfa18fc174cb5daff1388aa79e6d85b76e2b6
zf5769ddfefa30361e2de4b7100120fcfa227e674cb680a0b4e86b8d28a835a998edb9062eddecb
zf5ea9d58e0a928a9e48230d0fca01650fc486b21a8d1d628a1af392d68d9dfc9aa1e7454094cbe
z0110de7fd871b3ec34e290763dc6c44c291816f478e5aaf1602dd79147a4af8a032675d0a947c5
z5136ea506755e384d69bfe275b1f10452112b71dfe487331d2f29734e46b4f30ab43a5229fe0ea
zb00a4423958ff19be591a01d71431afcb89f59f03dc093d5b5722c724db272e9f2c6f4d20ba541
z21fe5c9cc6e6627da64fe7f4810bae80663425743f9b9ac2462c94fbd76d347d119832972a6596
zd592517dd3953d736a6137acc620eac128cdae9ee4367d2ef31ce58bb533a32a53e5d794382e7e
z7390966abee3ed97c5a159c5730055007dc587ff6cb2f599a02b809a2866b1ac44d560185e1568
zfd78f48daf1e1baeddbc6a26a7d707c5023ae8609e41f9bc6d452474099172a1a42a5720fce889
z0beaa24ee6893d96131d541d65d67275ffc3b35388bfe18471d31b415369d9ee8925c40590b290
zf8600b0e22c55794e97b581fd7537daf64c45ffc1f0ee7fe8ec1943384fc1d487ef49735fd955d
z340439f4ad000bc3597ec6072ad5c18a367111e560874bcc7c89f0ca4b6b50a234fc9c4b438761
z81124eb99fc5a39fd0d1d7a9a3a74a72335dabb20855dce7302901ed78a7e74707a6e0a0e43acd
z712c00eb8a7304475f91f242280c1c04bb0db5a2eb391edc7cd6dceb6504f355af37a3743bc657
z4b1c66ec5dc837741b40c9175a1bf948eb625a19d336bd5b27a13913a6e198ba53dd908d62a9d1
zfbd4079d51e590529ef544bee4c4aa58e9045d79149ebd823d8a8487094e16a75179c762b14682
z162c34867ca2fd81557ce55353175c519de34e91feb91bc764b674ce8b06216dd8136d3349b9e7
ze014f5c3f9e89fa13753c42720571c45e12ef2c125715452fd8d84d61704935446b8cf9abbdb29
za38f41744c0c03eeed535f0dc35ea04fc9c9ee0d227fffb8676a81cbea09f49bc01c0bad9c7f4b
z2c6810cf4d5364f3dcd80b6fbb613626f97474c0cdd67a20dd09e293cad5b15f3d61c51a87920b
z01cc2a6ec0445cf4954d9372d93ee3cdac4f0632aa061e5035e4770b786a8e3c451d3a7aa53095
z8bd7357f8a0a0e420e542a79ec0cfb10c628e599410891fdb7f8a674a2b7cede7df63b145eef3c
zc358062d00d1840e77c7baf0a65dccad86d169b00d4655442067289d67bde63f001001dea651c5
z436a3ec4ee6ccb5c426486011b699bf0302fad426d143a4e142ae55c10abd3f7bff1d0b9967132
z377dff030239046e0179e169db87ec7f15b8d5ce263b6dead123517481bd3b2ba953e65f22a6b2
z909e4e645419ded53695013beee16ffcb2c07d75e8451f3aed5162e9ae72c202495fea7b2fd9bd
z78bc4326baec2458a58139284033fc040957e23779d4fab54d8787812d7dee815ad19b8c2b5150
zf370f2b867c35181a630bd28d05fbc0a48ddb902d11f9bea2282c926cbda0a825e4698836ae51f
zf81a65cf43588fb1c8879e0736ad37cedbc782bdfc0b6d42c47787b07af69ad8dafef93e9f48a7
z4e5c03dc4563c91d1a384109ff07d0f7890c8b8f2c6655ce60bb93a91c53bc58eeea205a3926e7
z2366d4dfe8ce591076004c41db5c7619d2fea40ee8ea3df15433e42f30d297c13ec17976fd8cdb
z68e143f2be8985e93b84a1ad503f8e26092c660b14a47bb6c454859a2dd08443a3854f14d5ea31
zc5bc9afc1654b02c159f9c7e5f8639cb53b75bf9dd079d9406fbf90589a7ba48942edf485b2099
z78e038e044eb98ae16e84cd3e6541bb690271c2fd017e5bd07a21a94d574ef7ff596add472c391
zd504060a4c96eec31190032ed02739cc167dfc72f85d335c4ad9c110d2e3cd2d7960f72a67c9d8
zb8d7347c4e18b4573b7257441e2a471a3e58b3f50d4a387d00cb685b1a9b6027e4ea4a3efa1836
zd112216f74b58be28ef2d0bee3f49eedeaa881c07e57d56edfa5165e0ce35fd5687eddc6c59687
zeb09d771c062e5da7e517dd0e272d7bcfc029e5eb56f1b7ada3164596fe150076a0e387a9c1b70
zd586a2c0e6a28d41a14dfaabaabcfa18685d96f895c0b6132560611041136caa876243a5ff7d47
zf012fcb0ebf1940b8df028d651d1de303773d1a1491c2c89736da95dee8434144b835cea882f20
zfaf61a574c2b210b8be9044c8170d49b2568d8a7335715ca94f5524f52cd1ea8a76c5cb4485e1c
z0089fffc7a278aa13abce7ea3d875bd0ba18a14da7cf01167fa699804ba9a138da648e45e88cea
zf8abe7235beef8502ec2eb5a14b02db58bcd49d3464ebd227d78cc2330af72d21484ba11c42a54
z31e71644255dbc825b356e81fd32ccc0d56624bfca792f4eba84ef612edc7b915f7a4d744d3eca
z357b9f194afc6a794f00e73f15617cb6def4cd8d8365009a922594209cdbf96a7d27cf536ba5e0
z92cf5d72a2911d3d10ae0e4921e8661d16b494cedf63ad44e905084d7d2169df39c629a78bc424
z1026bf151139267d68958a51642953f89e1839e0037f68d64b03dcd344e7d76e6dae9866351742
z8ae269767c7dd429561fb1ed3fbf3d0e3cb28b2150476064536012db6ac0c5482e403f8a025dda
zff3a5141fd615ee0d0dc1a6309af905d6dc4e706ca4343123308e91a56c5798d18f312e074e131
z7a524afd0e0ec7f35276995b9ce9585474b04824d2d7188199a0bd31d9a11401434092cb771b1d
zf9256ae038ec72f6b715d0a7f20accbbce35eb9bea5b74b4276a1717e675e141af83d22e0636a1
z1c0ca8fbfead9ab1877ad7910818b0a25f719bf970dafc40ab9fb5411587c6d3810fb1f116043a
z5d242f5159dd10857fee3555df19abcec739afa1520ba2c600b065dc2a6cd3ab5a15ee0875a921
z005860d0450bbe5f01297f77942531b730303c0b4a645b70b25871c5b8731741b1fb824c98266e
z363155c69f74907d50baee2643a7a9063f4db8803167e18faed9cc39111ca16071ef952c6ffb08
z15038be88584df19ed8f0bdfda2de9e0f222f76ec19dfcb8da47bf1cdecee41e179aae9395179d
z1eb6de3ccadb84513193ad5c8976db534cf9855df0a6ce34e838b7130bfb420d005d1e7378a1fb
z0d090b8607e58afb51b6da58612a2bfa4d6bfa130cbd2fd84a789a0753534083889d26e1b8f942
z723f2ce8f95737f29a3c28ba238d195cb7f06ffe3eea596a3fbd6718e11ef1e9d08b6ad897856e
zc0082f691682ebfb554fedcd7541164110b7c0b9e33f5cb16d228b2a8e0208889b13c71b5fe948
zc2e314449c4a2b21fa8faf66216beb28bfdffa0ed8fb86663e5a97f788490992de79a87edd4ad8
ze41840c880950999d8fff61b8bffd75c9bd10c0ef225b6f105d477ee10a18f77fb1415e1326a52
z11112da744560da097b4c56130071459b8de7c060b1ca5f5eff12b640cf57dc638266e58ba217a
z2adab27a838b148a542fbce0443b311d69af1d4aa147088fcfbc3f7a587af85fdb36f4f5a422c9
z28e0e97ffcae233ca08b364939e8c155ad89c64643c989fea8ef0857c79b6b079b9804ccadb799
z2c123a5586525f5158b85fb998d27b81b4b7ea31eeb1063ad770856f75b951b5ff781ce8b98106
z662fb3d0be4053744984cc96d9dc4e73fc73f0c2458bc976c5dd2bc5b54b3ce4905fe3aa5c4a59
z47102e13e958cf50cf1daaf5dc7f5d4c3d119b21a6d75ab475026c07945c957e91e89b1631cc4e
z99d0628c2d096cfeb8bd7696b9e1b9571ac02a460486f81c7bbac020354db0a214a9fb07da8228
z3a382a796aa298043ad52f5a16e14655b738b33fb6f9a850e7c7fb75e8eaccb4be1f9b15504e3f
zf3661ee752ee657add60ad2d5a31935b920265088cee3beb2cb696ce447cb68e8fe239122aea5e
z2bb671c43a44a6b09534fd36291b7ffe667241b6866ef5b5ac811083e59d61a75828dcb32a390c
zcbc5f734711b229ae74fb37331b87e256a81c709ed068398a57f95364790e5bd7e52304ca3de83
z5e827a22acb11b70037e4fb4509a7d9462fdf35ae76ac7e1652a9aa727aaba4701f653e2f8c86e
zb42504f815063a38c5db09a39a183000332d67d62b692460102e6ee7be4b8e4a8f2acfd8e2dc8c
zb0bda53379beb534a5db4505e0a30f2674fe608bb1c9438116656da38ea9b774d5aa2e6855547b
zb6e155c733ec88141b9dca33df098308b67959f6948cd7147acf01ffd791e075fb3a93d84971f5
z19430aebb75cde00398bc482d272d71175cbd7c1d7c5310bb65f145a933c37eb2e0aa16acfe774
z010a8973760e00b52d00aa9ee74daa28cb27dd88242849270a0af6a9462b9bf9d6a219a850e6fe
z0e7b4d70e6c4a62abb49ec81a4ae2ffcf5d073f3c7575b150b43bbbb1f17ebea36ef6ffcaf629a
z8684d3b3cf796dcdb2003ea669d1a4821ebad13fe7ab0bc0664f8a769df3414ad743f31927b20d
z3caf4794dbb82de50b0c6bc19bd7b4e63450978d26d31362034e6989db92a1a586c0893f960bb6
z3836e88757ab52aa8c5b31d9640a89c56dfeb162ec13b57138c791977f8de430997e03f41dff42
zd32dc77e4d8a45c7c49529e00e09418f17a975a1aff182014e8faaf5df41a6ee31747de20c180e
z784b785f9de28a534ac4dbb0195fac84755926adba06c307742c842a34a07cbad15f12668a9ae9
z600c4624907bafe491601fd8e4681ad0f7ec1e3c85ac9793abb5fa529c6d5fe3d92127c0eb9b6b
za8e2d5ebed9309cf7af5f5eefad37349537ffea9b4eb363041c4580a55d061e956f9c0e07d5727
z5390dd6f2aae7b5964a152940403b8233a02d745e701f914d9d53140c07791dcb981f37d25572a
z7a3d5f09b8a212039d585a65bf2464f9e2623e709a7aed22de686018a0f42c447cb037e25b846a
z4f405ac515c492706ea71322f3f8bfbc0c18c8b3de84f0d7147dc92f4a2b77a54a37f58dd41d76
z679d5b7e10ec8bf2257b2d89e7c02dfdb23c2898f7459082701b682d37435804484bf4fc214d9d
zfd7b8d318122c9900988feb3c5d9a615856c5373276b1f1ce8999642bbdd4f3b12807faa911148
z5b925d0d7659a587c71e367acf7db253ad4ec17c6861d8e55c7529538817de9ed52326d6f2747c
zfac555d8b4b9d426efb59b91d527e71255fb7a7402d519682721a1723dc3d0b912ac43571d8c7e
z3c03a59ccbc9ace56a26f1ef619fd536c1ef3cf9fe0d8ace7e62d9d90ec487c5019b7f943caa09
z81f54e5a3dc8a850310b1e2085388fe6c8723d1e9a40d6dda6c98aeb943498dc1921ce1ce8d50d
za3ebc444860dc8c71df7ca29e943691e672958ab539b79620735f47cea5f20223e550c84cd189b
za9a1da9976cdab2fad0a4634a878211110100f36872347ddd8d202749ce67dbc4ed664890dc7b0
z350833c5ee68431862d7e917ea9bdd2b76e4c750185b75348e9b49b2bb19235089b89311c868b9
z80a0c554c63c8d03cedae188726ba349454b1d39be0fe5e3117366320d36cf5bcb96382f0e2469
z540ffe265591a819149f54f6f56bda844101da1db9eb1401277e464f9a4bacfa02647275ac3ae7
z9143c52049961ab58a12cb7cff630537345cea7a06cc8179450e1e35e1b082de27419cc0f9c052
z9370a4305ba72727bac8c57c3d6c9ebd98d111736e5a080119a32d251b5ac7ee6e648c9f3efd68
zdd4b8dcedc2a1b811b6e5c7e9ffd4b1286fb9a5bf9e6c886c41df22c6eac5d2aef1ca041d9c598
ze68788f52b521826397a42be57ba53afbd74ad16a0d6f9ac4f08578658e78747f1b869e0db80eb
zb74c507d189323c669771a3e90ba02cabc0e952865348aa6c1ebfe338abe8beef3490fe4b56424
z93b43b85a9fd4ded9d71722dc267404610179a1a12f9a2370517929d407f00d2a2a90045f33bbb
z5cc5bd049ae3df496b468b7522d5693f612c215da344282e3ae0680dac60ab2767404c7f03b3be
zf379f694839369885747489b4dcb0bfa0687eb5ce148e2380c3232d5e7a220fbe7e446f1a057df
zf7901a004db63c9de99ab6c6790b8f44fef0b05bdf2478e262ef04652c98b016df4bfedc187ac6
zfc03f4984e735987f2b35bf8fc3e434ff2d6b9e3eeef9d3631821ff0f12f8ce076e764c93ce5e2
z1645b5f90ea2d0e04bbae691b9d3240ef7e6b6ce2b7a3999e83497c0620c056ac04459bebc5268
z66814c2cd9ffcf1f5cb331643d28e4df77222084d8e95bd2424e52193a4f4fb4d924fe9c967fc5
zb9645aba04d6fba877c04e51c850e0ec48e41062f1ca9b44957c79fe9a89733fdd8374b4864c9c
z2623672eb6e72a455cd4053ca37dc0b6c7fb9e594d7dfeabc736acd18ec526e00e6be5984985dd
z6a0d466a9c87f46aec4c5fe2f29924e0f4ee16483cc5acb3a42054dde08df322369804950330e5
z906a9de15fe2307e7434d82906f7d40193e261a88c7829956c8f701088d4a6a817f648a79f101e
z7a5e0b67eb5e0592a59feb3adc764380e7ac950b8cd8959dced1445529575f2501110b0e5a101b
zdef4d34bc69bc756bcdfecefe6e0dab0a485d9df1a736bbf008bcddf3de7b925c7e2ea53fcbcfd
zda910e2d8eeecd9688bd813a68c69def8a9ea500cb611b227f6c6cc82db6a870f7bfbe440a94de
z1f0e3c7502f981276c009503d9c10c1705c21a89b9ad56dc3d3d9b94505cb1cc5acf0fbb72f7bb
z1db555c17e7d987fa4b2faf5f802e983d1ba1f852eaf3eb8bc13e0f45325a12ca6d55b09f007d4
z8418cbe731f98c446f89dcd8962fc744ea12c5db90467138c319da85d8c153cb8b39880b6d18d5
zb90c3eeef12612798c60bbc15540df5d1aaf7b62efa302d490334b3a3588d3e8e0efbd4c9b84f7
z5d22373b0be66b596d99bee7c970f404f15dada880de8fb78f78ff3f4ff9bee568c3518ffb56c5
z3f70ff0b765d7d772730c8a7fc17b46f9679772798a8aa5d18ddbd15535bcfb668463c5df69bb7
z1ee0a1fb4cc5dca69f3d44f7d88eabfa45ee75883afc0d197e00d3e0850193649d59f50a03dc70
z8a58c1410202b287c02a9ddfa445fd0f6252a37a9540e5b0380848d662fcf396071e9e4e2f4a33
z187ee446f9fb427ff03cd66ea0b0b0c6c7d5f07466437b8ec48debef3934a2cee159a2a7fe8a5c
z037b568fa3297a85b83f4782a932c37268aa9e44db6b8dbb0b3bd1fa1439ca97471ebdae23f864
zd4ee439d45703047eb42d4df540b35f322a6cc228f02af6e490bc9e393079d14e20f908ce7edb0
zcde4553a9fc8bfa38a7ce15cacae496dfd95ffd5e343bc93c0b7a34a75e302c4c1cb6ff887b1c7
zaa1b15797619a77acb4a55b950afc645c4e36f0437de6867bf0bf603da5ade44f19fc8feba45f2
zc6db189c4bb0689cf34c279f2501f9c81c7baa6e6d743f42abb2bee0159ce37077969d44dcf9ed
zef8efbd8cd6d5b1d38de8f465b99046ba75db575ea22227841eb1685c34857b4e9cdc4e7c52f7d
z9db430b6ff6b13948342cdc9a49896ab0eeec7c49c8a20b49af50c8574d104844519c930915e58
z513b61af4f7b066950c03533d1e8dc9b600ed9ebbd4f5d71879ccb3b475b14e924f3f1f27c22bb
zc62c1b8818de50bdd5c6e2571f8d1af2c186805e24d671b2c8fb773d1f7b896b85e87b9352e26e
zf430b24cb6c88944935ee1805e1af1e5cc3078010748e1b42416c4bbaa346c3ab6f7d4ed516d0d
z15a6f84dabe5cfd8a6540b0db832507b975e27d4de517b8bf23ccd4d52db75a0d59bb964da1ae6
z3c445d579d7d457584752ad8de3b18653a6c5de2353961a2b80926b7d9b8e71dec303f4c15ac1d
zfc0cc1d1223079c06866c8ee5edb7036a5dc8bbc4df2249a1ec57d8eb6d364af11a981096c9848
z3eaebed82f6e40adece3dd47bd5c023772982063357f6888bcbc74d19114459595ba884ba0b653
z40b9ed0420664679efd728e6d066b51a583802e49d43a1890bace25d644f6d541ba7c5ab722fc3
z2af4d86990268cecf9ccb6cc645eecbefd841ad2b763c52b3308798d2ccd101695ee1b60408379
z7965793af8c9e27bbbfe5a77d451a7207e8bf1879a0830ba5852cbe097ece78c2c8d4838fee63b
z3e46232c3f8e8792d4622e41fca87cd3239fb758de46503c0d518ac95f82c40563fb323ba2e138
z1a2d55c5c6d5146669d0ae3995903ff6dffd2ac29ec1675df27243a8bf26ea71d9d30bff2218fc
z1b015988b3a85daa97a6695325830d5f394a8cf6af6e7f41a424ea497ab2b1a977b143532f73cd
z8b44a4a12e15826d7c64fb4e51cf00c9bc7f8da99a483e99270d4e582d1cd82ed6048db0f255a7
z8727811f3ae095affe6bf78517fabd69ae225424df5aaf35bf7d693cd0b737e355e8ed26a32bb8
zfe37f7c74c9ff7e4b146000d49c2f6713e5df8769e96e10d94ceebc6a6aed782316f4c0efa4820
z1d59feb1f2b3d6039e0e0b10036d32a9afcf1ec04c64bd6b507a7b8b0293ef7f656a4fabcd5fdf
z207637020f60b46423cc431631378ecb7a63e59149636479c2cad84b7379f5fcf629f243fffa9d
ze7f84d7fcefe3cde9887e60558c0ea3d73882d14f734bd2b81aa8355949f46e3b52b66a8ccb0f1
z122909de0913b2455744fbc7425056257e4f17721c1fd3d96f7a06d5076b963d80f428740257ed
zd2fac6cdd202c63c747005376ad19a350ef9bf0ac19e1e5316fad728c996975ab2d3cf6317b850
z715855dede2ecb426cdca562db40cb347e3d6b544c01914ec8a686505397931327da0d652e50ce
zcfe06229441cbd1a312fcb21838aef3f4b5a9d671ecd20c21c2a2a5e6a6c56ca756f417e1cf629
zbd72b8417776f889a6076c38b7c603e935bbbb4d8804d16e729388621cd129df551b72e2655ea0
zc7ac378f5131dc56b9ca128de8f1465195b5aac68530db6f497120d389d8951de2fb67ef79396f
zb4e85b71c2f465005c6b68d5dadae3a2d674efc8af7a73cd256e3f4c7beedf59df8f262e7e6d5b
zdf3da7c87408774ad8e88626281f43db6fffea0687db7fa9fb1631727aae34baef5146492031ff
za46d10b13216f07983a8796dcc97a3845e6d13bfb3aea5a9cbf8dca6d7d21500ad39b36aff4674
z09103d6a13425e0aa90d406b9d307a6b561bc86add85deb6a2452aa8fb3e65b1a595347d66685d
zdf2eda26614f97e567c011714c9ed1bb9fd1c263ede7cdd23772b4ac698016fde996ac3fada92d
z5e72ac74b834cf4895c62aa0708f5fbab835d97cb89ea310e63472e4371e84c7bc4080a1011ff1
z836391650a33406225dfad4002d26412da1733174489463dbd90ca6c5192fde94fe60add3c5584
za094d0b9dfd4263d89533edd660b596143b8fb49649357794f8791d351114cbcecde29468a7aa8
zfe56dc3245b325a7e02695d786e60e48c89eccef0ec03894acf1e9f149c55211bb9643bcf6eaa4
z2cee1fb902f49941c3bd2787f81cf7d96f1b21261ce841dada5dc5ffc807f08e1c96739451be38
z8694f50172ed27c0573f7b80791832d983aaf83bb5dba674b94aeedfdc8e419bfae36632664452
z781cc0fca49b81f824664b420c6f09644692f845b1f8e1c5c2827b67b3633dd2e2fb07ad371d1e
z92b86ac9dcea5835ffd99568e9e5de00a707b1ea42643a5a1550c1d69cd5b30e64f571885bacc1
zc635abb7c9e883b2cdf3f479a480c570a8c7a023dd5da313c0ab57368075f3496cde8b07604902
zed498c3fca7db52310405603b0bc8c7f028be978a3051adc3a69c994a1ab2542f84242a8dc5934
z089de339cbd69c6239879ad62b22558326c3dfc5203ef93740887f11bdca1c5b330eaad06ed4b7
z1e85c79809a91035ad79dbadab6ba3543b3a05d37f4f1b3c703c2863bd50140fd5f7189a7b39ff
z7ee97770943c5a575b0484c6d7954b1d37c74c6f7f3f87db887c1fc61537644b52f41041328baa
zf799d14db44e18a86731238a767250d4536afcc040224c7afcf5f98c0355e0696918f023642789
z9c56ccf20643fa6378124fd08d98b90d5c27dad2e2ba2750323e6578a696abc46bfe29586b866b
z1baba015d66253ea88ebed6227f7f9811cdde08b0b0c5b86491ab6228b160406934a6d86b1eabe
z13d02c27f93cd1e3d0d7eb91881fc22dfa7d39a5517f9af1c09462a5bb7ddbfc497b0b92720604
zec42fb357d9f9a1c088119308db86c1347bf549d4569babd27487a55444132b873482be0cc691b
z9e405c086d8240b4830d99ff9d90c7dd96ce93f8b8ed7a2e47a25055d1d78f840c76b3b6cd50cd
zc97e75466bc377ee74e9811a2182b5f91d6bb4190a43acab91207b772b802cd62506bf98119e78
zbcada9067d6176ce724c8c96aad86c3ea5c516a1eca2b72d9d1a24189cec2d62d631d4b909e610
z462a0948f953b052d0a31db9d19e1decf89ed79d6b23242e7c9358e47fcc8ed999dc966658ee4e
z075d82297651c768b1010793f2d1f73534088f651f288689962444882360958382df14d6a836ee
z0b4e08ad30d29b9ebfe7b01182720d304ee12f312c2eb63181b8134d9780567e88f042d7ed048a
z3c7dc9f1661ed1fddd6432b0611e3cea31ffa67973f186d8e9d4334c9db3353e2c17877cf06039
zd45d977cc5a7811493db5cc562b214da17de2d2157c86fd1c5328374d014e248477b9b7fd71ae8
z6b43da15f23df9ca21e39a089d7bf125a7c466cca02272ab4b99d02eb6ab68157143d55238c6f3
z8d87ffdac3dd45cdbaa24050dc7f6ad013ef96c9620541eb0f65d9c320d5a1e97de3297d7806c4
z7c3ff6e8a1f1b89bcacd2845cfe45ce9956c6b5c41cc7bbceb27dd7d69508ae6258f5918f78ca5
z5dd009efe667e0ed8c6511a3b97497e476b46576c77f1ab7e0b828c70c6ed1b00950d24cde2725
zdac1ae958e152c6b1ca508b1e71719ff9f0824f727cecf28862255945b93bc3fe4399523651038
z4115e4fc81a283d0162dae1070df9b48c687e614b220393651df190e566fe93d1f2f95eb2ff845
za84bcbbbd76d639cde2fa29f8b24babe8a1bf22e2db84e233f7b2d9c562402c76f34fc3b3363e7
zee63ed5ad93fe84f89fdd3c4a56863e0db3eadf4e7c1c082b5b48856d5255ca10fec08d64de696
z1403d5a9bb35367923d7163b64f5d307f6b02a3170e331cb66365d53a20bafc33db6d0af53f201
z8e19ec49822096872145f1c4185671022e13fd76824b145260d89d77e51b50c93fccbc9856c19e
z6ac0e0f23c1c1e77af6dd3cfbf4d54aa187f5fa40f8fe9eba79fc29034089742416ffb344048f9
zd69d63f72cdcad8cc785acd559e5a1d7a0c688e3ee01b3f799b809c6914c9dda5d64cbddc413d4
zbad1f11d03a8eb26de37110b444056cc213848f4b71ecbb76ace31a1ab2dfdf5eea5ae63e9d9d0
zf29482db62b8b7a35d7945c5960dde76388f830c41285c5c3b26811de31e1fafb2deb71a562d24
z569e52bb76a3b294fa474b63d51370e862b8d3e4972c903b261c086dcbfe67bff5ea6b8e46b4dc
zec7cb319f1bda55da0a19e45e4ecbc6d2dfba63f461329204f78a447f717373a91a120f31febc9
z6b6f446b9655763f86d750396005d32f370edb08c0a49dcc67150c56e5dfedd9755df2f2ba9f20
ze81573f954670b50955f1d6f62e9007833f88a4eaab523383c872c6cf0c69fc977b5784049acee
z2bff1fe21c7cf054ab7c87f60858bad16b14ceba688cd68d3d2effd170abe247df1909efa8cf55
zd5f6b575c4c43c1428fcebbc6715eea3730f8dacdabde5143cacfda79049f5ad2da7236bb602c7
zdf7f822612329ec2d573a6c39d2360cbdb32bf7b308c66d05363f54620cc13933121aebc8df2db
z80ef2f666a194ed4c0f3e41b5f959a8de3065c0d67bd7ba94fbeeb46be7397ca2cc9693aebca0e
zd0014c3ddbf84f0a28198fc0a9c00639853545ad1fd87142e642a1fe3a31fdd248cf7ee8b94a9d
zf4fa89f4a2b162bd6217f80897cd1110f156510917f76b72e10043c35821f2faf2ce74584cab7e
z976ed8d9a58143cfafa87274ba0bbc5895f2d0062bb2b84382347b9b6587596f32576cae956fd4
zef7b261a276be8e6470c888323c4a3db30c8451ac75315e4b721475e713a427b0929f48ec11593
zdd4cfc62b14d958cbfe54ba721db8144aaea2071f3ef4a6fe6b491486e6d5f825ee52640a56aa6
zb0d61757ceebe22ca08ad41bb8acb32b82fb098758108a9f4f003506351550b515debca261a845
zf54e15635ea62f09af0c669a96e5f47df2d060e234519b3320974f1f5c031b1b95f8ec69de6bff
z563e356881cde9060ac64142f488f554ab363b2d1c01abfe45e1c8a503a682abf08c8d77bcd651
z8c7774d8f9409584a1ea29fccb3fc7f9d06ca6330a01a0e58c3725c476d7d636523197061ebdd1
z10769d7bc2ddfd59c87673bb3fb8e076e0324ff8917d5971cc17df72daf8be65b10e103a4b30c3
z1fa301b6248572acdb3a7b3b65a033f44d5381aa045149aab38c8773189e5e66308320bb31cc93
z8a0837a1648fcd996b09c3cd25c0e811e985b2585e8de7499904e8ed6ccfb1070bce4e59985267
zecbba49929ab9f741a97df42b06af7530a688764dbfab345e8368159e8384537522fc14390534c
z14313df31263662039487d2bb7051410f51ca951ba0ccb9819ba2386094fe0140ac6fbdb54b743
z30eec1592bee2da2d36ceb83249e508310a95aa4ff29df6e280c94d47fff2388255ef826fb3d00
z12f9192beea166e50e514a86a6acc615a5779604a1f4166ee887ee43a61953cea6228057be3ca8
z16162dde4e18e13343f52725d48d5db5587505e4b7f66dc14309788ffc8d4dbb53e2de0c58bde8
z76125eeecb9009a8836721447cb46975a1c535ac76f8555fd31aa89c4a0deda68cf1d8e0a1fcb1
z21327645008cfd7e61eae8232a3130e8d2f6e0e1963af2a8fefe26cd49a99c648627e9383f1cb7
z2d5716c27f2d7b3fe761e6bb37ae5e1df33ec44a3fcc83b5893b43a5475ec901ea13aabf5fa5b0
zf1ec0660aba0772e06f972114a416f0d31c6d8f5afbe206187f1746c9db45bc36f9d4ae02d9877
zd8ee7dc9b4177f18ed73cb158c48de62cffa6354a06e341cc40d492fa5b96290d284f3eb9069d4
z54de869119196e2e5cdaac24583f98272845b8a9a86f23115f086af575256b0497d5f9d0718d37
z71a77dfa42cb3ba08a8e1e59a7033b61c8161892475a468ccae945411df0d8c9d242746ec25c8e
z1320cb746cdeef9652408612e63ff9bfdfc92ad25f66ab0c6c2edbca180c61ba9466320ebc70ad
zae201baed0acb31f609a8f77a47ef58bf2b8cbe6f0b3c3105f14c7a7e20e8db3f594afee504600
zd038e1506a480e2277962471e6153a0af9ee65358c48603db0ca53d49fdcb3e0a323ad2f53f3df
z88792797637d5ce858c7fa78ddde2718a32d7349e4d765e0847b5fb8af2a039be1e12f3b162c8a
z8196f97a0ca2d74cf7406f0cd585e876dfe3acd82cd14690387c7130c9e0fa15c671f1eb48a149
z4a19bce1940bf8acec4caa11b7b792a926456c3e3f4e7de9d4371896862da0f9850bc459065920
z7f46630eadbb9cea25ecbc1443af6659f8491acf3fea72862ae289dce75273bed3242b38c37044
z57b2f0e0fb04300dda69b157dcc224bdd086351d018d6b2ad1531f7d60a2139891ad61dcf46da7
z964298142bbd142cf2685e363620d41ab2c7a3e7ad1d0a5d07795759ede5461c15bb335aaa3925
zd9a3c60e98cdd0684d5a2562d1781b71db80c7ab240dfbaf8d9cf7ed12372b0fd01770b0836d1b
ze93739806eccc3fb9400f8cbebcf3fb5438b55569f07b63c00fc043d4889115936e1ff183872a4
z88e71ce850f6ab2a248bfc1e9717052fc71bd7a520d342d1962a4a76501e5e6f873ee96bc690c2
zeb1c498b74f4a3a31fe05f5be3a6bf12e85f57e31c25b31e769e5eb075964bf7cbdfce29e0669f
z0ff9ac9c5a05d87fff8931d9abcda1581ce678828c9d29a24a6af54dc344ee31d0c51239b1db06
z39d6406198fad73e0604bd8742da326da7526e4103c71fee966cbc2bc13deccb36ac54a7dc102e
zd38bc4b4db5df79676b7503afca64fe64273938ccd3fff94ecc215ef4fb4bfcec03899fcd420b6
z9575fdf6f7f24eceb66ee793f242a2521962e1b854268dd956e301a1cf666c356aeb48c982d234
z1dc05165f8fe0de20aefe21c0c251b017ee0253aa8cf381d6eeff2f3d9a86f05039b77670b9f9b
z3bc30bdf849ea2e68943049894a14a3b083a252ea990290b2aa1df6832552b4ac6f46051bff46c
zea31da668f90b535efff000990812e9f151ee83008a27afaf48c5ecc4231e2d36e61801750bc1f
z6952dffee13acf8b2961e1d60041a20ebe3230c8b61588dbdeb4e5de286f05507b5d9c3b087109
z495a8e39539973cfeb95b08c3dfeb194a290313d7d0922422c0b3482a8a472c0185284c352a816
z5b0cd8504a4b8df84db24451276099fd988c5df047330bb73a65dab4e3c816f2449e31ff0e22e3
zf6baebaa068cb72e40a77c54a6b0456e70634b20f026a6e9612293bfb22d2d5cb930775a828cdb
z294be2b2bbe918a42f76a061f7a295619f74e148e017c411cc06a0ed671408101301d284ea7bbb
zbd9880abd4c32a8d0ff17fe3ecc98512c555365b4084eae6a6c14cb597a714b52584e1a030f2f8
zd508272cbe735ebd49dd50691fc1f82c8bd673c4e56e3873a7c68e8120e9996030a918e0c482ab
za5e3a6c83d396fb8968e50076d9ab6c07d81104083a19e3431a66f3522a989fc0c42778b30f339
z5a5cc8edf5fc4f971691ae3ca89a339f9ef3373ddd1de2989dfea8a5be79a4c60ad7f896e498bd
zd1b80f2c7c24883187d67f711372e57ed22cda991deee71934854f6ddeef5690ccb7be82e0d944
zc309003e569e30dbb3d0b6b1e14d858ff71e5598b3fa96394ce2df58d41c2891f66507dae02a44
zd7fcdfeb6df1ab785a2a3cdd17661598f0777dfb79ce1dadc7a7038738b4bb3234ee2c22170ec2
zc48c979d880a7996840d4b6042583fbe50cdfbf80f5202cb472b859e9a3d79ab04913ec0a498e5
z030f275ce132be14ff5aa5619714cb399d76d0ee76950ddf6020a514ff2da509a8effcfa051b58
zeaa84ab58fc5e741490adb28f095a028b3c99c322be6bbdaf63862e56e1c4937a331f193c7ff83
zf22346c231f41d83b7c4eeccc454bb03f6a7b2ac62fd11d15fb42dbb1f7ab5356acf6f52dec50a
z245bf68dc9ee78e9a9c2cac2ceb7cc291dcd602c7e6a4bd0c40150d420c2161fe122340861cd62
z7727b08594ee51cd7761c3a04a603d64e7136c344ce20054d08bc4cdd424ba4ccc8be936723e5d
z584b0c5516b2a89f89b4e0c936b16b391589a5cc55f0d93255cdb7f9f4af7beb121302121283a7
z2ddc6c06375b327d3a3df9837ca2687d21e0328321af99d4208ee8e16ab791fc102e256d7287c7
zd1e7548342305588882ef85c4218c5df65ae799e105def9cc0df8d8c0bea3018dfabd6e6f9c62a
z1d9e207df54008c6d8699ccac7e99381bc48a305e7dea65f07a336014d348f2cc4bf79916ad08e
zb3bac51d43be920caebb55e6229a30023ae58174a0237d4bb4a977a71857c2357b7c5758b0e991
zd1d446d4f7af1cab5817862f83a08507105daa6a40e16bb9f7055238789b84ccfd9581f38046a5
zf00131a86dce4212e78040d5ee958b5c99235ef64574559de2d5dd7092ee72bef68341e51e98f8
z780656f4d9ac9b8ced896be11fa85fdfb5bab31677ac3aa96c3feb313cc309c48cfbf7ded1ece6
zfceed47f8e2adf7d1ff584a614b8ab919b852de251cc69b3ed12008b6ea5645d260e2029681c77
z04690efcd9a380be42171efa1f4136a7bbc59401729376b9e5e5640a343f849bc66030fcae6aed
z1d0130ba80537841e50364e4bfe949da194d129af9bfa83b3251b77df69374bcb3331b0d4ed286
z3ad1512ddaef8d89db138c586e48f9d9b913eae299f2fcfe4bde6ca8bb474112280fe4e9e72fd1
z1453d678780723e46f2e9619e07fb38a47f6da1a88f5e654d8d1aead881040910625c616b0d6aa
z2554ae9496cfe57b2cdb8e86c949c557cb6948f4d7d84e1a7b79879facecfd6a6a986f4b2a5294
z31cdb3d0051bce2be4d60562a27b90ea1e76d65a3c19b7ce23705eb36706c6c42509edfea97fb8
z74c756df54ef830bced5c0f1c97eef87775702a490fceb7a226a73f5268ca506f677a0c144f41c
z9cda3fa42fd1e2c8a95c284c881ddb53528702295019d39c48f8cd250039d0fe1fbf295b01b61f
z48c65d9edb2a403d6a0f967a9454c142d61229f6ac58c5035d09d22c69bb2389c34385f86c72bc
zfa6ccd08627820ac1fe6cd7d2fc56bc7fc1d300de4e7885ad975ebc47dc9931afec952279e3804
za060716b0b08557dacbea735ff48d4c31ad10f4f568b6b57d362f75138451611f9671aa6794cc4
z10b7c2c3662a4613f43e0f1332764924dd415232f7bbd9583464987f02a17aabc42267eb34c976
zc93ed2a5e512f501f9e14311e94f5c5697234bacf059fc179c77bbb6fd1e4c1a17d8899ed8842e
z4055b5c236d1bdac7e2ea54fdf83469d4114d999a3361febbf0787396d0cbeb6d6cdce76b943a9
z67897a9f4072ea19ba50e24df78f9374422af568bb95ce85aea53fe070bb290da2719493046b0a
z703f26908c8ce3144fa3cc1d2958bb077f1a43cbaedba4286d229b695d419647860d84a26921c8
zd49d3573832097fb2be51ad41a12e969ae21832c4ea3da3aee7818d4154811911360b4c364e798
zd6f099e0a5acb4a27ec60df26bb47a4da477e7ad6cb35d27e293472a69e0afb34521ca4ca4f8a0
zb925f1ab58e431ab72c4ac5e03ad7412da5012740f131b8121fa559c329ebb364e31ff65ca95e1
zf0183a00bf568568c37d6c5e309195ce23b23aaaa0735fde1027163b5d98ab3500c0b900bc7329
z85d7385e00c426fa0374c7c2382f2998a95545932f01c0d839f36bbf71341c9022f40c4961f156
z17956995ba3fca15f4a6c7748969e74053f8ba4753389f396e7ac9bfc90122a60674fceebc3645
zccb563266e7a322dcdc910116715d1a30f21196f1bb6acab74088327edd464c3d1eeebb477ae27
z5bb752e1d3aadbd3773043d2595f018d796088bb4220dda9de41c4a6ff2efb487a4e56b6664c88
z543dc9a84f40d7a9d28926abd34418640e6f3ad53dea4332116dda2cd3e84b3edd1bb4ae382d23
zd936ee074f5106d107a22bce912563bd83abd89d9f304884b2df43513b16737cc665767129e92b
z135e1fd425455259b1923ccd4183c2de1e0666b400d9596c44128b260b4e23966536dd4bbb7ace
z527075242ef58b314b38bb53ca37f3e0d6130f359439ce7da3c3d9bd6624ec19591f45641ed9c8
z6d5c394e630755449722c6dd03d5a7e6ad7544e9875f0e3f63de41f8e89235176f7244f37fa345
z931dcbd833c1938228fe4e00704669a8649f64f97930e5ea0ec2d91bc932279b9f31224b5cad52
z24c9d1aa743bb6a1b5c24c5e656ba80cd43012efc49947ee19f555e34c43b1600fb6cd752d8297
z3176ca1ba9ce633bbf74de9164dcf108f991419b06c33a0fc33ab515725506eaaffea1a5cee322
z29a2508c68681389f53553eed67a5774a3af09f327df1ac734f489973d593f1d7c3892f9feddd9
z31b903d7a6f087dfcdeaa5a4c381a5c77550f5c275a1ee3832286d62e94178758337c9da68e3b4
zff1d4321e9934aaec5c753cd664ef7f0d37d449062574632f649f932ba0e2cc73f3a22986f66fd
ze3edb282268b589f8c499398fdd16a27988994102a39b158e5fc05748ec66a016420910d7b6a08
z2c818e83b438e958767e02cc1ae5da70e9fb091fc5d2bcd7860bf4d4df07115c67c4c75fa243cc
z892fd134ad496205c4e5f874f8dd01ce3d72ef5128da2c9d8e5b3f675216a5325707543f8567df
z3d299bbf073cb164413644f99c56a2b12e13f7f69cdf41a71f5c571f169e374e5d55529eb84bdb
zc9aae0120469d99aec56df63eda51c02e228778a314b9e2c52a508723513ea6a7a2a05ba2c3f3f
z2f3b8aecac9818824e4930313168950a78c0ddf8f7796d51cc09efd433aa7c2dd37c189df504d6
zf764a34969359e0f361212df2b4f4f9cae75bf6e3afbe094df489464f0f78d57399dc2cc900579
zef3bc4f556963a41f5811d898bc4cf427b942c00460dd2354d3801b9a849a19a1c39c7c358e973
z4ee70334fc5daf1df394c9c460031833d72f4e40984f9a9b7ec393457b646c6257ea075f90fa2f
z317eeefee7ae293565267cfcc48ad4358da5bd2f7ce5030bee339537c52557461faeb7be704742
z929aff38a03968f758417cecf39ca94ee321b22de89fbfc5f5535ce57e5fd0e87169a7c8088c15
z5211571c30441e53125fe6ddb0b9bb470810c8520e052384b4d6444313b764668aecff5185d73c
za98a7a25d404150a9c3a7b7fce819dcaf7a77c2526e5bb98bb3e42f37385d583f4fb6f5fa382a9
zc8a0f6ad666b081c081210d84d1400fc48108ed010d646b9c10f0984f81ab01dbbe7907f8bf810
zded91fbdddb7d1c98162594f16946ed613de42b1bdfdce5bc75ad85aa0fc7bac2024041c9a6cad
z5984afd15ee7d51f43595ba6d00ab47df4d19a0c82cc0b54dd3ed6836c3dd9525a5dde0a34fda9
z1c362ca41addea5427d31b328fec7000cfdbe4f4fd160bbb78084d959cccb9759999bf13629f20
z716d3e09283a8d303617f2f909cdf79dbaa33ad4655bc07e718be33bc99593629ce2bdb2062f64
z8984050fdfc77c030c7a4f54100109af92549e69f46943102c9859a5dec464ec061a3ebb7703de
z3ac1c1220a511bf984e9c5ce8c48069c34446d6be258d2f6c356763d9e444c4cd04bf40a509eaa
z460673955a99e75390665b57fca3f624c087a40748d50be06c971ad46e363f654e2c0b84b89dfb
z06b2c702a8b97b8741d7bdc0801437668b63d680220ebb6e167f79cbb2f80db820b34ed629df4e
z18ce1b02e89269f26ce0f6dfc2cddc0d31466e8900c7f7ee65fd89f601fc76a2760a9be577549b
zbb5e43d1f50bcfe7fbf87b8b6d8569adde44961008dbd4aae7b26f3d6796860b3c99c69c1d243d
z5b7f62bd4436edfc20aeedf213e4291a28647cd48e4614a863e67881a33e644f45baa2652df995
z15d444c3a4baddbb55dcc8852806b909f15d8a6f536450de092f5cdf6be87d11b4172e3a63a48a
z51a301c096b9c93e6cef381f014447f470c5b423b99754795c14dec96a34e348a618c4ccd97ac1
z4c15f83b39312d2337df815e142455856ba6872e42ab0df844a9b1957bd3d2b20e305dcc253ae4
zfdfe50a2661a6ff7c24ebd98dfa47d6bab4c6ded7cd333290d6ca885975054c24dba2c87c63afa
zb961109ed289785c890865012a101f09f6a37c3fcccbe055a95e79c8dc89153abae10071e79372
zfd9fb6ebaba16156ea530e4a2ea3ec60d0746a7e57972cd6bc747061101f6156f6f5056d51e693
z42f6612534b6c9f96f863c9e738c8011eeb1738492d7d6aacbbca4d1bebd6da39ce1cf84c83137
z2daadbc6352be12197f7ddb67890d60c1f24ad4d5fdab5cb7ec90f53173384685fb1b99933ef7f
zf3321f47ab7478f1739963db4e5e6d1ae030fe8fd57f27d46209d42fb7e3e22ab034bd973c086b
z4a9ce1604236b1c2d9db02bf1cccd008a0a626992e56dfe29fd23a5e23a0b177923fd0419b8eac
z194b40b650d49582178e39b90a393ae4d8ad3580e8f337300c453ba11b386593fa35307e30b414
z03702047bbff85045774864698d2d3924869f79d8d0199b2621df752820b2593654a930ef7ba8d
za854ce3d89b033e347a09d173b2930835b09e1f20b89a968523390cd9851400d7e14509a178c3c
z2a699c531a2ee7021adedb48b72db285677c35907e229c9707e5af4c42576f1ba31192c859a2bf
z525d1f90aee7d986f0c0dac8af54cdab4298aaca2e0c91d4be4aed860227e9a9476f49bc306d13
z2b293bf567dc91087c9e9d86c165abefe6e481f1287a2d0568aa9cc7848ad16c71d4ba99cdd06b
z36873cca06167034531f423b1c1383938490edda8a11125801d2268030fa3f82e54fbf561f3a2d
ze04cbde6fd601a735c9499d6fa61a2b44fb95535f7263e910cb2422281aa95fa0de5cc77728f50
zb49de5d6f0abb870ff2971277ba2c7e5eb1ca0e5c5ced72530fdbcecead1d7788c674ec29e04e4
z022cb02d4baececf14649efcfccda06c77d883971204591d44ffa47e7ee20be47643df7b8827a0
zc5a773c8da65a3cc233a4edbc9633d1f317de66082fc336ce5b9ddd21d74ff897ab45fb3f02905
z58fa37fb76073776f8997fdc037893760e192f0c52018be82c86a9be6582ad4a46a91c595da0ad
z8a2434fe6f910a24ce61698d0b3d5c9469f5b93ec153f38a850b154d208f6c43871da1a72bc7d0
zf0eff575c8267cac38bb2fc8526daae2d12cee05b911acb31d6a1cda3f4c44708ad0852489ce4b
z24c4976e5ae08e40d06b966cbed59180e6bc2cb420db7e35d5f2e7fe4814d3e945bbacb6506962
z42c6aa0541a1849f1c3c65ff0a5661e58a5788585ac76e28ebb45ca42374e3dc963b63cfb9edfc
za54c557f077eddc4cd2ed387a0a10516b477474b3810424ad25dc3b3d6152c8335af6bbdab312e
zb127c0b5d50a373aff0972c14f08d4b4183a441afd9e88256e1ae55d8ba24d42b87e17dab43393
z17b4b8a6615304fbc134ae9a153779b7c3e09c11408fd6f304c5725641d0c1bca9983a572e5e62
zd45840583e98721a3f4ed3277355975418106369aabf6211e9e9fb8b6bc05fc7c66d296fb8aba3
ze7a276ae279688f0fcbac69dd9b842dc294b4098f10c912b6dd08bed2d0b09aadc16d9aef24629
z6cd600f678f8020715a185c7d788117457aa6ab046fe89dc19fe74ae8e6bbcdc2c811e48aa23de
z8dbfbd022e381b806ac5f1f4f5d5e4d70df5765f9f32bad815a099501fae64c971d68657b4fc7a
zf3b026acdaf737c5f4607456bc303b8c557601eb716f68fcf6cee0650561d06ce63a25c42c9c03
z8a37af68926ee72711847cba9d3f4f73716a116859160ca83cba6288d873f4959535d87a0a456f
zd4b6c3c509034302e26f73b2d96dbb8eb6c569a79fcf917349769c73a467a64991af308efd71e1
zc9c072fb185684231b7d8590955db4aaeba6048255f32340ba6ddd3d427c5610a36d0317f88d65
z39f8a60325fe3b6beeacb6af2dd831305615fe9251f76f88366f9d6b170fbc95f1157f23dbb7b1
zde41ce7d5b4a44c24e3fbbcb318eb29fa484fc30321f88a9eadb0e564287c9c0182475d3a28ff0
zc565e462d4578071c051396863e7e28b8cac3812279924ebdbb5524110801ca91cc1de81e7414a
z8c38c67a2ffc6ccd9b08c1579790c0b16eb663507f030f0fbb39ea0fc64a5142adb3c06d764856
z6e1a9057aa6219325f346e52ce851b549351815e97e726f2266e79fd5d445c10b9339d200c472a
zd9d0a7ff0e5356fd03f7e8ff1a5ad12930b5ae82c84f8198fda96552b7246484e3bbcfdbfff1f3
zf160c6614d35e3c58435dc98dfa7fe3456c1eb98db25270fff6fc2873ccaebc182767c57c9bd36
z03ec720407d9c7abe5b1117309c3ca697c631512873926cdfeaa5ea8a3ea5bfe829a62e1e0c756
z005d2a678570d3d54353cf7b8ef0400be75fbf64d39162280bee13e5b73cddc252f4b2ca43b879
z88c1d2993fc1f9787a8f21c102f62c5df100ee139bbe53c20f5432e062f789ff8d78e540199614
z50c7f11c4cb129a34525365a03c60c9f9c511d105e24e9aa5a4bff650c84c61689f2a1e7180263
zf2fb0e01a6119e4437316b4bc231da83a88196ccaf86b42bf53a68b1c771a3346592034a1162dd
ze9d7bca2e851b8e62bb5bd479877a8513f113604b8c5cc3b33a5d2ed730f40c0a447a03eb8773a
zc813f1e126b18dc35bf4a86bc0f698eee0659267f1fd1294efad2796afd527d4f876a7863c89a4
ze28fed7a7ec5796bbed1965ab4a46b448dde9eefe3aa48429a9a83e6462e49100940dcb9634609
zb3255bcf6daa3230b816ad3075d89abb3b756d59bb31ba9aac3b9dedab6b88e4d1ee9dce95c2a8
ze0487c077355d1fc5d4da76eb9bf27e5c88185e3934fac7c041e106d1194790bd7a1a08b8251df
zdb20e252dc598ca4993b9195f47d6dd22b2f3287f02aeaefed961e23bbafc52adf302eda7fce49
z21e00428eeff46bddae3995ac4d2ed5e9b1bf35cbf78ddae348ff9e95b26ae01fdbcafa9c37f32
z1526ee9f2fab22de0d324e1cb771250d0fbd4a69973fda899b7695600eec694fab5d57286d4b3a
zca961ef910c6052ce6c5ac1eaf59ebc6bf4aea4d3da78232da3f7df54179e60aefe86572a3474a
z454c95c3592004818b34b3b026912d2009c8a49f399d1b67fc83f1163d10ebace2567491809c72
z8528cba9f2c6475995bb4e02e8b3fb2e7b93e82af0eb789e75b188aa32f539534bc4469207515e
z40d4092147b0ee08c974db7dfb4e65bf43f72a673467439c412db798ed93402f7991d34a8a336a
z5942eedc7953743daa444138395d933e16e0c34f7fdd57cbfadaf0d8e444cc8b0fe5ff9f5b5e95
z9cf5936dc813b42ac30155b85f6fe6c30f4ff7cc48d3c1e03eecd8ed9984a47133119073da4ee4
z1471d7d39874e5902f4bb57b0bff68a7640b49874e55a5e91a236fecbe20b4393380f7f08b0fe5
z635751e12aea3d07307c66181b4a5e2f44e202ecdf150fbb805b485828d6caf474f6b5bf0a7b10
z4b35a709f75e57f01b4d0749013fbd8fee8c4598303967c10fb0450df1a5646652a6f32aa90cc9
z240489b6425fbdbf90cd0353080635fa93e82f45436d2ef326b510a719a839607ccc09790cf7da
ze756a593ac9e6a87f1a0f72683f025f6a9cd9fcc349ea89599c268acbe801d72799c3e6961441b
z8b0ea81dc14d77f4b111ce8f10b31ae1f2f549a99fa37d24d381aa4a170579b78b9c6de0088567
zee9bdd6632ee436eca9f5d90f35f5f705263bc70d5a069d85f53393033ddfcd612025d2604747b
z403cb792c43603f6fe4998679e377c6f621bb3115b4a3d0d5c28a9f1d130787f3b3800102d90e4
zbb9be8c8b8d1f001a6b1740a65680c5481b9e3d0cd2b6c0bdf49817d26a5b46fd3d6cb10564eb9
z6a5a0a4409594151184556d43933fceace2cc8cf96ed4f0ca71c4b5f20b4e8fdd11f6bb891bc11
z412d5ec5f71b22d2fe192226ec8fa59a5468b55e5bdfb6009643591bd5a5c99a0ce7c2212fda60
z034c31876248129135bf53636cbe38a4b2680178e46e2b80a6a85c237eea4ff497789c8c304bc2
z24eecdf9f24f815ee241cf001b9f59a20cf6071add466b9d403be84df4aeb81059ea4201c98c44
za4d417591f2a41de519ed4451f25d0eaf3a91b9e9871c0422083d12e10403af8162f7154826711
zea1a07b637028f4bc4fed23d9224b2b54cbcfd05df6f24d2e58fb16cabc7ce0dcec12a0cf45195
z166c1dd8204cc0484d1c6cdf55f1f8cb8a2e158773ad8f6c3e6a49d13a3ddbd11a7b6ddd1ababa
zbda1c5af8adaaf25d8d5c8fc41c8cc8720618981754744e4edde31ab4db1280e06d201f4a1b13e
z1c62ea4832589e82147f1c934a0ba738cc66446628362e1b8a26b0adf76d1e4aca084ca910820a
z496c0856f659616e30f405df971f453f6a05f496bc0dfb694d7be1083becedbdd3411e9a9aabf3
z5add2a1a92c6d420fbd2c103827a49a0bcf10a8b8818da081626822adbd92ce01d6ff1916bd54e
zd1cb1976da4c52e381759e9642b0e686981cc676a2d79a8751038ae9c283f01807b77d20a2d628
zd9f8a04ba424819428ae9a074ee86fc6c90179ce7c42c4dd179f8a0100110cbc8ce11b17d6d6f8
zcef7ccdd314a6a0e543b2b156a1ca52d64b7d6691b2e114d1da8f612ee584e00f4c4b04ae1a23f
z9945e7840796b50d8200c39ca2a70d6854a3c63de6a5a528b81f85dbf6d6b5cccfe0006125d86e
ze5986267de222d5fcfd7675df75a0870670aaf606a90b4505d5799a5dcf8c54f0eec7638060e4d
za26ebfb3a83dd480a0a0b8dfc6ad09719327f410f14891f3651dda2ea6328d8ae58bd52e7d85e5
z54ce7cf6d13c8bc2ee146ebbcc954c19ddcaef8be680a1b4b4475c3e224cfd88a05b0fa5da40b7
z20bbf6f1b9e402b3c967d84c8f4ead514748613a168c0de8dd84e7aa3f241f6e566d972280d078
z2020ca9599c35ab06ba57f354ed3fdb64652d6fc77c63bb313661e3261982db6265afc2cf86ba9
zea1e2e832295ea613c1c6e6f54e222f1903e645279da1a2db5ec89030eb0baf08d51a8abd241f7
z7c8ce4069f873112b7039ae826557a87d17e87979c9e5e5cbc72c38601f0d1621e8afe8f0cbfbe
z63c8330315296f6fc373222241a5c26bb1d60de14966ad17e7c9191e7f76a068aa6061b2571993
zba0a666170317181d3e8eaa6185948bfcd2133d971651f7f6edeeb4ff0d27d1ca54a3c5e321f75
zf8c07f9960742eaf290151d60bb74275089a183394c21430e2033e9c1b31e5bb54f4f8078100f3
z8029b40578d0281e6dfb39f6bd9d5f3901e99acd3f6e0523af929a7c096d8d21959665b2062a46
zc43867b9e473271da5123b5c89b98101f3e652d672527ead2e650dba1ae0819e678f3d280d6ce6
zdfbe251139013b9f4cc2d219786bd36a6300e58232652d89e17abf70474eb765c800be67471321
zd8b5f1cdd666e1469b78fcbd62ddbc5d09b84a7fb4f53da7e011c6cadfd1b30adf3bab3c07bb99
z81961c0d2e814bf804a51fc9505e4e9f4675cc69a4692e0a0759e0f37681282ee7bae833a91016
z519fa22dd55aae5203e499504f3c83f19c64f3f12996bf9fcb424694edd4568ff72f8e16601cf3
z4328a9ba9aafc9168fc0ca174b6cd7f0626c038d0cc4c88ecb7519238f2bdbbbbc7a14fb145f0d
z0ca8a1b69434e01146a47ed9678712965f3683b8a95745b4cce38c89d7e2325249eaafe3a8b218
z9359957aa1dcb21d5ee0d7aa46a51943c21c659524c5c9d553b7a607372a0468cbc023fea76d24
za0979d12f2b436908ee108cc16e3c335529971749ca31ebb67301908ea35e5ae02d3463d3f9942
z6c605644a3801c6b11e884feab308eee5b8c8edd5d10aa37424f669fc3ea47eba833c600b0666c
z96800eb6d79f696cd8eb2e34ba4663585e404952540411a817ccf9f25476b473c817bc2fb53319
zd23fdc133af3974c9c56184078124863ec320250e6660ea6634ff71820b619f38eaef44a27290b
zab9814ca8b6735182a78c91c7284bc9d374f561a59501ae128b6c7df5e773090ba5356a8636fc6
z2b86b71207e28a8f0fea7f7a02cc242579fee67b0d2bab12071b2a7e49222b6f4d61cfa42df0f9
z0688f4a59f418b8cb3c3f653c2ff1b9844ad6a52e3f2cd2202e1c4850270bf3038b3735b640df5
zb9ba2455b19a2a861cb76779ec8cdc0b64783cb2578a7725ed6566078143ab79a0c54567683b96
ze1f17b1812380f47c6aafc50310ecb48d505f978d2e4013facaa59778d7104e20b6b74e3c8dbba
ze635f6546b4d66cbbb4b9d2db80bb11e847f06b487b8d3576a18bcbe73046c05e10225912b03e8
zd72f66c79d059890e03e38fecd172455d5b6eb44e536f74ee492d4c4eb13ead3d82d7026b9f9bb
zd64c813c8605c867bc15a4ab0f3eb5e3ec4260af7af3aca6b1e7f04d9f49a7be9c3d5337b03fe3
z8d4821001002490425fcfa2c5a93d5816b02498d57f80b484693cd90241a2c3774d19c9c268741
z92d9ae695931b14e2b215b7f4ee9f3778795165ad0c29f220b4f2a43625d65d3b455158119e422
ze1d480b16a687b7c84d07bb7b3e6e31b1aa2db7fc547da9756a3bc824497a157194b6688468a59
z0b82bd7aa8175d94d22ff13ca89311663efac484735d66acfce19d635b0a17a6f7a5fdb83f416a
z26387a5267aa19802a61d527c3b7d6f0fe741b9bbac8747cd28125dfcdc4b5e6a663763826f4ea
zcddcbac2fe26892f53c198a348b1f4ac85660f3c42ef6ece73e0cf51dc27bc674dbacdb80ec8fe
z647ea3f2caa9040fdf8dc7199ffbca620ca1607b95182fed80bbfb5a52afa8066024bf676c8345
z95c98c18a8d11b20c68987e5d640c414621ad9d41f1ebe2715156f5e9302e22bc29d3c7fbe80f1
z3d1a1cadac8f864e81875ab29d6b39208d0f9219a35cee137aab1b0ff833d6b32839dbddd3cddd
za7737ea9f8addb85f2b6e2bb2e0c01615b617adf300f7e4c815f3f0f418a86621b2069d49c1ff4
z413fd795539154f3b9bd0c21de5ff3de6b382f3cf6257744d0ce3d8da1be197e13323af46c8114
z9baa3ab5e05d13f009eeaf54ea992b4efdb06f4e6d7a9ba09cb894910cf5492b635aa52cde800a
z2a2ccee37b5f9e9b2eda193123436bb24c5943c54861a8f7c97f888e82e1ad0661d682066c92f8
z247548bef46f48a6ffbbf7cabe844fdafce2466c0fd2038fcf671a1d78e10d4a27ef632c656a32
z62df3b743ebc6f1a8ced77461cd83ecc07d511002c816c37ea29eea4aa74479a0a51fb0e0301da
zcba7530d34a83fe8baf5a75483d7ab6dae69f3a99d8bb0aabe601ea95c4c5160ca809c380ec4c1
zfd33c1fa2f421b605df8c1dc1e5af76fc908ca78baf6503c99756389f46511bcf78f022db9dba7
z2649d27dc00901ea0f0b5d0007a38514c4aad2cd913a6dfeed37ea361643924a8f3c6c6253d8be
z66962d972a242ec4f75dbe0d9af7132a52dadeacc35f7378aedf6901d50bb9d3cb8a3802e94e74
z37ac40e291a494c9d2445199e2d1012082382fe3fc017f6f0c18210058fc8b8258c4fbdc80b117
z658a0cac388561e87b38f890979a693887b438010f0baf2974fca80608cf074638276382c518b4
zfcbf91d84e537686d2810baa05591d43479ffd7ba7d75ba3ae1cf1ec3c53be22b18f1ce95ce6df
ze7f5cf5dbaf9b91becc43863c2f6087cde14eeba3dab52dc9ae175c1732394422a948dbc17f72b
zdde7fe8ce5f83190160c9f515b79fb1c3a0088762304d6d8f0fde3f77c79f76339178bce577821
ze3ce680954019072c7a89edbc17fe397a246577f358396a0e6984fa5227dcfa8d43b845bcfbe90
z6567a77e76e7c5a78e53af1110090e1bd953e37127a6302aa62ecd3cce18bfff2decec9146799d
zee272ccebe2cbf0dadb1e22a154e44e099c362ff8f5cfad233abc57c8784478e7a6f99879edf14
z10ac5f9eb396c92390479af5ee1b079404019d3b101abaa13b976ec5c7d780c036351af81be566
z1243049f621c22d21975b7ee5440251a442a9322d3504b014b7cce1bbcfe6e4afab7434d7944cf
z1fc94541f921c4e4dea99f79a937e8361ee88359c233e67911102a0bd80700fa0a94ae6719f53f
z86a0e49b3740526158d90808116826551aed673db729c019d58d9ae0dc241c4f873343f5c50d78
z99e1fd5be5d51802119e5c60afc92c226422753ad7c1b5b257522186453e3d7d8077a1d8d8a2c8
z203f20c3eb624dda75422b04c5ae582f477e9341347a129bda93a86d0d39cc538d8781748f0ac8
z5007f547067f9e8555d820f9308e3a517f878c1dfde2b15f12ed0593379545967bdfd1619e733a
zda002d95f113ac4d19a30d95839c423749e343f80b0de6fe0e552946fceb4074a205fc448cfe65
zfe80f245ce7772135dd4a7f8058a237e9f094767bda8bec18dd1d5bee1ecbc63ffaf1c057a3903
z8cf0868435e4a841a7f80fa2991348434cb6d41cd2a65367a2c4a2ebe7c55ac6cf242f1d94af63
z5d076c584e74a53ff8ad13ed99d32ea118d0030752c4a41fbe871d19198fc202314f4ee3545780
zaee76ffba5224e204899acab3ad6fc6197729e124b9d4b4506f78df42b382fbe0626ff8f3da10c
z783e132f06c08c45054001a09c0dd1d657b1e03ff8ba99e1d4f079c960bd25ab7e497f8a91a2d4
ze5d68af0365c73d6e42988400a389749d7400653efb6d3c07bd5172df9f132af2aab1ba4a6f2a6
zca3aa5206b7278234b0a368735de0a61c01df1f21e0eb1ca43ed0b48d9696154e5f1e0e2551af1
z39128de5a85bb2d22a6f9f43c3c44b0cdad5c916b375b15c9935e54444e028a56cabc1b2db3896
z7caac6132a99ee0846c5b6e398640a3ad6c8c07bbba782340fc13c484c45d4c8ab1bef071fcf36
z1b2b0b37904f8dcd6aac2505cb3f322e0f93892fc165afed823bb1ce7c8d7ab5597cbd0ca30353
zccbb2d1f3472c72cf63f64d883ffc785fac053676e7a504fc98df04f6033a16c57d77c8494e98a
zd553c193e16293cd4ef30c01730130ea6513d044888f8504c19500b03942d5fc89cef5336e28fc
z241bb56f20247e344497a02c2559f283c76e5fc85f8d344fe6b3a26a48e63d7ef50f5a3e5ce734
zc476cf52a4510c0a84419a91061f267827bfea123624f8da4804af06af7cf09070095e40824a55
zff1927b98208ebadd4ab33de05c1ea20a8be6dda403912ce7d92d1498e95907077610411c3d21d
z72aaacb86bfc8d93ea93e90358d0d3a7dd1a272123cca42b8bb496b536d25a8c7e43b6acaec066
zfb87b99dd4e9251260fa124cb8dbe6f3f35f1b24b37c29fb0d3c52e4f4aa40ec545ebe97e370dd
zab2d6ef1d90bb7567d85c19f476cef92be8f723667b2573e7038285068772d1a34c86bf67bc9df
z62b8b4d49b6a1d13a2bf5558f044a81fe14d88e490ad5f8dbef17af0c8e0fb8d45d5b5464fe207
z427b7a7fb96b01c98a866ecca632f9ce5fea866929ec520a7acbba7d48abc6a73b4dfe6cde5bca
z3840ac4e1de3f56de3cfd9dedd6a67f18f4c918872e26a63681e561696e2e8635e59415eb0c9c6
zabf20d81d52f7039a713e45e76dc18d03afdeb0aae87c59e30ced9cca606d1f391e119c80affd6
z7d1bda08e1ec0d6f5d9b9388eeb38c091c5ada235307f0666a8312da5112521bc08871d6941315
zb122632292c961af478d2e12289ecfb84b60e5c6a83b4481d2a5104b79425759b3822d6184f494
za00fb5b565c29db8d350e55004bdba8b27888aac606d6b5fd08e09b6f56072318aa7dbde09c706
zc5fb51ae594212a982688976d2534492d694b52a2eb31c7d6c5833dfafb70281619498a2d92c33
z9c9e5fb6f4a947da334e6030681240aee4c83413bb1a72fa61dbc90976e17c90d9f4476f44afee
zdd2858f9ea62f9bc812b82587dca1c341c64654b569f2eaa273458dc78b29ae9ec01a08299e66c
zd8a949f8510845941bb2a44b62316a994035c732b459a5f2763a9613972b5d168f52f7a868b3f3
zad80a9e86a6d08c8e2f6413134eb3bfc0bd9eeb4c93bcb5c6478b5e1d2765fb7affa2dbbfeca87
ze7e044e4772be6dea6e536da842bc01e87bd1553f0ca87cfa3c9d0275b4926f6b19acb9c0838ad
z263181b47450f4ae92be62f62f3501cbd91584607ee1df8f2c79030887a9dae71750844b1f664f
z8b307ce0f3a060db71148b490feef3259d157d10ab855e815cb1bbf879adb2eba2896603eb251f
z81dbe29ac6f9d484dfee29fb22cd5bf498a4c37bbcbd8d00d6196ec03a796a2eb90e200b37d1d8
zdd4fc43c0a7b81445ea296ff56b796ee8b7aa9e0235216e6e8df7456bfe17722ebf82f653364e9
z0ffe87a357d73404354ae71056fcc86d453224d270ee937f7476daa219b56583b7a5faae2e7aad
z1f7594363fc25e2938f970a4f8c7b147f2e8e9379a5bafe2f35c654e6b23fdad401f77d7c2093f
z46edaa67f4f31240f10cedd03d288d0af87d3470914bf414f1924362eb321e3f73d47eea1a4ca3
z56b0cb9b5e298224d812b588a53e24c211c1428aa46e532372a870bf3ded45d79952a5566b8efe
zf182ead8eb3c914a5f7e6cb6eddf071dc93a2ad3d98eb43b964f0940ea8f47b55ff41365860b77
zed5c7a7c2c62667cca3557afbeb408b09e188f0a50cf1b3d6cd6bf67677cbc4f13c0550f0b2d93
z09c30787df7c8642ecfd41b43119d8366c62fdd76d66211f3d0714742a2f62b8f730418047bb7d
za187425a3add1fe4ec6d1813002ea7563f338b4c3b588a14fa512b5d4d6dc39ba2a3681a1039b3
z8275eb1a3feb24433be4996fa31f24e57f8de1c3e3d45c9ccbf791c30078a495c7e75a0e42d727
z28ccb181e70cc639dac530be71413f01a97d9357b210a4d2ce7b951a0fc9baf4c02792e09ec7ce
z406899bfb9dc9c5d1fbcdbe3a716bd72bbbe19858646a55c5879947b5186be4be9fba21548f2f0
za2dc343d78f1e1e9febe0229b4c7c3f62defa4914478303201dfd1a7dbbb782e6fd42d661816a2
z1c8631e0ad7d151d0356985032b001efd508b5e49054baa5387aa9cb7d3ff5ef5c785b8bbc9b60
z4f90a14dd278c12f85584b74e0384711bb24132590cf3c6d188ab6902eb9dbba3632968d585d3d
z0f15f51887b6bae45e3651d17b528692f340ff14061d272af9e1bf444f5ebd6f62c1e920d5dbf4
za58569cee198ba9d27753f7ab43bca4d01ffcd788799c2294cc2a75a5da74dfff0441812838831
z22b81c17f56b63d9802b745279662bada2c259e6b5e6fd967be6b19132102441e90b136df47368
z4f031195623dcf48ee825c320076a9accfc341fb0a4abed0ea109ef73ecd2efdc1eb310a89aa09
zbc6ba24570e0afb4292e53b3a65219d61816a87f138f9559d6f3044c7a677b0a6acd7f022b8430
z935f5de0cd4054a2b1757d6d271871180476c3c07a3b028677bc1ec05eb363849f10b0af3b1676
z46c510c528562571c87dac1edb4465682f7b0a03fb60f301adbda624c68333dc2e8a194f4ee08c
zb97be628b21b54514204cf020ff6cee5b16077875a3b00c68c636141f65c9ecddea39c1c363399
z35292d428d91fc4a28acbd35a8d61285601f4532540449d5b07d923ea35f9619a054cc0b569692
z776af83027ac4f5d5748d3bb67d3a0430e5c14d688ac3e060631dbce24678ba6517e041cc2ae55
z26a33cc5190ea2dcd5d6592327a81e493f506d820901ed4e44eaa1c22237fe4753048fc90c6aee
z9208dcaa100cc35a05190088f244380208d5a271b2fea098959886204db57219d33724c58bf7c4
zbbe740ea9077ef028ecd71f77c171f13d56d897b1b074d7479c13fb1635ad53ab3a939792ab91d
zbec72aa06d78cff9316a9f5630fa460774372361ac4d2d7f955261200ac16416525613dcb6ec81
z9e790a73a9e107b49c556685037a4bc1b5751786248a452c0619dc228c0ba1012c787f7f02e227
zbd30c07404c11f4eec44154307f8f51269c15dbc35917e0d8b87d8e280c3a2c2a90af9524fe397
z12dfdf56cc0d50a9870b1e6828161ffeec2a2e5b51efc12174dc90bf337c57458b3ca8f8cfbb66
z319371f5735a3decf6c965eee1f14766183ae4ae2fa7bccb49f0c26fa3c36a804023b8f625502c
zc6f0643284bd8a77714c7ad8f87c236e39b4c62832a1c51e327a40cd0b0a0b82af8e2a253db251
z664a6fd5e8449b5ae65bbc53853ba5bd32104251bb8d14b2815dbd6f8b404b377b57ec9619b1c2
z971ca55dd8b563600e7719871073be78b9a135da0f71389116b5d19d3142324a86975c188da9ab
z1b88a5e1da35d2f58460838aa9bed093122fa010cf85cd1ecc8953d3621afdd6416e68ae10a2d4
zb8f770a1be6a92f063ae7d7ea9983f9832af9ba92516ef8f85af2cc7879abbd75159c2c878cb46
za47fd7608bea17cc946a925c32967bfdabc2ebc95c8436cf8af532bf4d392e806ca070b97c6d10
zc273ee3a999e4720ce2a7214370946ea2d9832c26b4df764f48d54b56a1cbc1851e9098bb4ea89
z81511c5e41f8e4cbca0ae1154dcab6645efa5eb0b8a3ed431e38cfe63897b12ef564995a20ac10
z24c2873da51b5b2fcc7f25019db45c59f599f7f73faef77f21890b374cdd004e5c6aeccd4ef8c9
zf03aafccf9400de1ce3046dd4fd11ce52260ae9a3a6503e7feea029ba1d78eed1a7e39818690e9
z3cce96b476eb2303bd4c72caf03b60b5daa9dad343f45597650e6652677f74f54291dbe5139805
zb2e080aa3ce98e0756c747fe9e6a521e2134c52ef1d325cbbfe13b02ae3ff4566bc44fd8dca0bc
zea0a33f3cfa7d03a56e6a8d2eb5dec50b9548b983b8f56586741fe160b39579182ba5103f9d944
z57345e9e2b67620ae896b0ccc48ce40a08bc1a87729530e4ce2a1c5c5a0e6f5408f5106dda1126
z0355321c951976077b31c323a7f954d0bd0510e4da05f01413aef121112b9e927b1a03c1f49ae4
z9613dd6ae8fb73377861475ad71e9e3e426d1f196aa73cb0ddf3c54a83f43d2f825416420c26f5
z86831511d67577dd21bc4f83a9c34c3cf122de8c1319cc57f52297a38ea5bbc51d34fc7a0c86da
zd7a383a2a6a593d3b15e043d45707194ccd0cd6a2ab307fc4bd2ffe9f331c6f9521e73d93c0c6b
zbe98f0d2435849f454cce639e49b5616a9d7a8b464c9427a692bfdda497e912a0e77557cb52352
z6936c2105ff8aa9b4ed3a50e23d0577b7dd42e552dc539c621f65bf200e2c91b6a842a4cb22f52
z3a45ece013172de7637561eb282eb865cfa82cb514549ee7b328399fc3c323171fc9a149d2e42b
z497dc924bc777aba2315d6730b99a9fe65d8c0805d49f59abb5f3efb11f43de6128f0f9337c056
ze7d921bff69efdcffe77000cd8210e8e38509f5ba375bc67f21b31786be1b109b53201079081ba
zb07afb404b5874d3fe57d85b859fbd8573c1f11ad579d3e0ffc8d1ad74f528d994dfa9339c608b
z395cbc1d58d3370e2da6b96340ace89b6cf18a5c6b43cab4bd3f0ab56f4b54cb38e99bf1f829cb
z0b866c1da5c56c2a74578ad2c6ae3110a1a244ded14d42424c4c62a2d08aa9b34057dc3f393b89
z20ba5934d66b000e6a1a5549c95f87ee88a532def1e0a1769641955ea4bc98280b27818a75a3b5
z18d56522d032e576ce91ea835677c5b662aed2f821f48d30f683d970173a22110a77b8a7e42426
z5b0d32992e1ed81a6b2d02bbfc9ac97de4ce1bd31c3c0bb897a96a0eb11ac7dcc954d71491efd5
z3f121af452578fd7b1d7c73bcc17c2851fef318d11e142530b420d4a86dd93658db2bc7cf4ca70
z0f62f2f94bc43e320710faf77e85e1398b19a66db78f46b6e956e338c04b0be3bf9dbc163f182c
zd75d7dd6cd9ef2f0838f78548e2ccbf51ecca5d33d75308dafe7b844d172f5bda8d249bba836b4
zd3e90335fdf93d0189ff3906f1f6834f6a7bf80f42f5a53db01bf8431205ef3101cca8ff799db3
zc9f9bdb94849dcc843093547fc26e112cc6909206cf565927bff72cc97d327d46e14343a98b94f
z44d4fab53eda4a31bfe450ca57b096097d5a1ddb51be44c79f79804b2921c62413a7c0261cbb3e
za6e0ae374792e8063e1a913c7710fd2324f8442ddf62c1e3518b61d3a61024e354402d4f6cceb1
z70c7570877853efdad494b7677355cf67b05612f087877c83011777e5a3b94a02dd77f08e3aac4
zf45bf83ca72b60193242fea68f81c14b66f2f3c0a8da5de85019ff199da3b249a7d2405757dbc8
zb5db35c12da81118ce9c0ec11c971f49f16c7a4e07324942d759922c74bef420e487acfbb91440
z3f161b93c0ecd72400fb5675db1aa7205a047ff3bfbcc72a1e71a25b2e416c39f2622941721e7f
z5b3bfa092f742d27e9508ce06f098a1340eccd2c8a88689818d403311531b9189155152b265349
z3cf817c4583707bc60ce543ee1c48f3eef0d020e996fcb8c5bd8bc6f7ec5d0012f71048edb952d
zbc9d04056f0652cad9ebc4d1a856cbb31ba4dbda926cf7f42d66044d4957c11f75c71211e12754
z0fc3643f25b8e407206597c6f56c935ef63b195e34e7cc9a811543b637b4cf3be835f0b7fd6173
z055794afeb2bacb30a66d4393a1801c684b0aa64411e75dafbc6636d5e035b8c95cbcfbe5ede2b
z02cf9d77d16eb3c76f2fcc1c8102989d3abc6631f747f7993e940a2865bc3f889401ad7d3cb88b
zb33adef975c477365e52d6c20fe78aef3428127757a2d1c59ed20f484280e7ffd1123b6e6f6f55
z121fbf683a94e4383e03d3e8ab7e14e3afb9a2aede1c0b273a98ec172478888ae7c70cf8a9f72e
z4e8b59fbd27c1683f00f128e46250be67ebe4ed686998a055ac8a9f7c885eef36d6fce0540dce0
z5fe1beb870817da1c10af6a22503d6a6fbb7ef2d5d227acaa13e7a6905b26464e76756f8392b0f
z961837292aacd12ccc7fa9eb68d5bff34ee6fda51ed83792964b4afb167775f971cc7546fdb67a
ze71d2f7efd89c170f5dfa85b184698b8e7c1a06cc625de0c78c1ecb493cb44063d5c6b6af62bb2
zab051250bff9d2963eeb256262c9bba0c1715a7d3164c095b3532831338163a833df1a8d6e9b60
z6abf31dfc9986c63803c9a51670aa10c592ec26b5eb1787e1545950a6d7883abff0d68a75739bb
z52400c55a0b9156c1d8228dedb1e3823d219bd31aa72f43fc683076782423cccfd3eb3a9c9fa23
z8b974524b7740478fc081a748441882dc20c575db5ddabbe9778a256d4911391a42b81d075ecd1
zbbdd28b316670090d59e01ec9f3db15a0a5bad51369e2602337bc7645f09a8a7e778967509efe0
zc81681cb3e9e8ddc2068a7404a9063b17420c1a5e1fdb39686fa0cd167af39be128d1b3fa0f366
z2bb35c48b914bb0e2f2ae51eb4b84eaa2b9c6afe5fa682e0e5331300f575252b936784b45f03f9
z98def39ae446c6c766844d8234b5a3ca1d272e80eaf70207d68a2cdcff1ab6cf630c359eacdf3a
zf5d744b6f64632facd7686fe352275d76c912befe1e46c8242520150342c613d2324547cf59941
z7e0f30474354b2de0f2f3031b37e5c80dd235704985c79fee7a23d98c82593199b1a62dc0c46c8
z862ce3458e77dae29f8d1ef6a7c53cd65521262af2eaa2b9093f8839d0c7312de7eb2132c1e97c
zf774228749cd8f8584e92630293acbc696a3fa58f8b97a59abab8b17eee68e8720a335f419c19e
zd8fd167bda9ed05a5979784153ff334d89ed4d90dd5988db9752b2e1385c4d17dae51a27b65f75
z5f2b4ada58b3881a1ac0e349c5b7b64646f843e1787aad2f5523c9e294cfc22f7ab54c571eddd2
z65eece5eb233522ada36cec413c3aace084b3d4f4832dba6292db7dc654ce1c9e92b8f2469c654
zbb8d0c6977331123d9ebb906cf492e7eebd225bb3324210f382fd4ad66f606c6877b14da9fcf5f
z9b1fa39d8dcccc3eb85dd81fa8e4add16e0268c66e33e19e647c8d1a15587c54217694f3838341
za5edcab147543b210f08e99164f55a14b18e3c6b1078572290fd8758a74c1cc4c564a9b0eba8ac
za75763d1de4dfe2e161d74f918e5e3eea34b23435d8feaff2637415fd3a85167b262119e63a578
z20299338d71d9bed936acb5807338fd191f5203243a5c827cf619a81923d8c084b0c25a6ff5f02
z1592fcc827272b0b55a69fe0a61186af9c05fdc10e3847c6be5abc322ad9b317b7228304895ab9
z3994bb5ce19180ebaf0de3b36bd2ea7a52a87bee7bcd5165235b76d16592fdc8da8e3b281178a2
z1401d8544c26dc653a03a6c406a8427fd605b7e43500b26520dde23f32793cf719ffd34377b87b
ze83923af52de8e446d785faad57c21cfb0940df5e4ac51c3874d1c64e3cb6adde4e9917d5a6460
z91986d25ccc5fc36149db880e52a439fe454a6a6dca6990d74f5039c8a8ed4edb8fb6e11926767
zdc6104e95f0655e5d2976c17eb77aef39c7f2ea05dbeb97b5b183b24b6e0710724a19deab66658
z3c84c41adf3012590ae98484f52a35be1fe0a0df7c92b8dd7b7cd233c528a42260c4da6e07f186
z0f41f33cfc7d771a03a82965d655a525a50845f00590c52a6c6caf98bf0724d1af2237fd50e054
zf22b2824ac83af9930e9cfa4296d1fe22eff370388a9115205f4a51d1eab592ba76c2745fd0614
zb810bec2674d7fe5cf44a00ad3ca0d15fb1e6678c9367d94ef6d4bcf7b0815b1b3c59d978e6def
z5d12bc9aff079bf0e8719931ae6cd54c612a06c93e70747358a146959a1d964b1caa169fff0fc8
zdafc478938a665dda09f5f333733d8991a7393f9a5a9ae823c41d92a4a051b5265f06ac597dcde
zc3a2b7beac496ea1a72da0f6c0397f55f6a6b03feb3e3b7c03fda22864b188292ae613b2b1cadc
ze2b35a2e7aa818b18f72b85414b01d6633491acb42311fc6e0612927e7720eb54e849410239620
z2907e34b861f7d4e4020a6d06b79c040d10bde04853ed58f2e072aaf7d4868d8d2eccf9edd00ba
z3a750615b1294312cecf97f1f7ad0e7fc07e06682302a93809c2589bb84b5f2e8d941210db163f
z5c6344fad6962520158c91f5ccd9e3e5df75bd7d075598e24af4fe36cc918ff3e7985c1eeb399a
z7359e558bbdce6516fccc445d5d064bcf4718602658a3b9dcd08358351b44bbb81f56faf145208
z70991c53a83829cc33abb264bf933dcfee23774ec3b6d6d94d12f919acbd2b5ad903f9f447e6a0
z6ce68c3c422d18daea59e6de3008cf3ed26f83071caa957c313850ce458bb508e4767dda4b8565
z0a39766a7dbe4589f4b81a5989f558929a7b2186f41caa31904946feb05b4ea2e708faca0cc28f
ze151974dca8ed07eec42cc19d7fe3299f4036875e31ffb9617f2d9fa7568ca0ab11aaaa338f8c2
zf700243bfc98f589ca69d0965ba84e0b16e40d2777b81b22977a2fda7643906d2a9af23a91a7c7
zd995dcf0903cf5f85e799a72741dbde64458546ce65a9911568ecfce24662868c2900baaadd4cb
z63fa9b7cb675bce773e92e06ae30643d678cc6f407809efa220e49fe6d9bd496081cc84aaca343
z2851470e2d63ff8bdfa9dc34fd3767bf16397edcf5ed19fac4a26323d25c9c0eca5acd28a616e3
zb0845fb459c3ba8e0fb84f635094808f485ec37f02a58be443b5ce494f09de07988390605e8d9d
z107ad2f8581b0ded02b95b4cabd90e8f8f0eac19c1a9e082fcbb1fed7f1b22e91b022220acaf37
z85483b09183eddd373df72e6dda88095482671eab0697a3886a4cdfb8b7316b77cd0fefdb527a5
z1c9f24aa967260d6b5e9d8f8374594c2e92ec7f7c15885915ca41465d479964d96e0a32946761f
z996ebac95fd14f0e8875f17c6d7b63b2198596af418829aeeda2a05ec64e13ffd5dcd046ca3aa0
zd923bf9389b09284d71b3ce38b113510ce20d1f71e856f46d1c415e6da86b1929ddefe0128e078
zd1468f1727ff51fc1e858187936bf1ceac8d06a7d4c4f9a80065e15b14caf826a9f917b87ed694
z1ae0d2113b571238dd39485cb863d49e5b7dc4f5795fb61dbcad3a702639dfb9a30693fa8f188a
z2c4547612108999cdb0b922a241873b0492ad75a8c949769564e673197a225736dd5856fec2f2c
z485e870b4f556d0023fb075177102e91833418bba51193c21abc6f045f3f7db4002e18682bb424
z9a3e7e638974e30637538247679011c0e8033eea2d1c82312506c6b98251ff105a535198d81a7d
z5f8ffc897a216b142729557fa98a1245c2fd6db8932a0a807f93c1c1121f64c2926cc6f6e7846f
zc9dfa43654b90e46eacb814a90b2849c2e85d6a431cd347a2167162755a1a76e8b30df13faf032
za6b8bf174b7e6d2bd5166d96812f32a9ff7786b865360be0251e5b1924f9faaa737241549dfdfd
z2c9fb83c1daa453ecea9d90f2f97e72ef4731c9d44f90bf3d708677f6f91dc339c86c65ae8161e
z858bc9ed7ed8ca6aa68126bba24c566c2a70a705c6a799f16859408291f5d662c21bd1b5672906
z9493f4219d615c9e42d79322a4534c4c03e5d2b9c80e02705426db7d615d4842976d580ca72d77
z1b9b0c729cb95ea65a0b3aca715a93cd88e250b62ba1593170f4782ef08a7ebd3940c835416d18
zdc283d4e8cd8516dcd2f89434ae4c80ea8354a3a64e491f5854eb2bda3939132218b1296510fde
z782a4a104c2146332d634566fce8ef0c0575328fab525ffcf8afacdcaab0aa91481ec74f2230e9
z444ecd6e787064d6230e5be35ecd676590b1708f8aa220b07f515cee041d4e24db1ca0de89cbfb
z62c12ccbc577912b865ba4908a87ca9f7e7db5532a82c9b6e1e76c3787475edd7ee63271256b15
zc00bc4796c73a4683f368c2f2e3f5af5b707efa33ae2c4f872d5d6dfcf209c9f57621b654d289a
z67046bf43524a4d25f3ea7f32980c41d1a3d8971888b166cc6436b00620b12c8a237994cbb0139
z41d1e0831691e5b113057e686bc111e2815bed6a5383ec4c4a4ccf8d5055100c1edc3d055c1e98
z62371779dc1987b9fdf26dd5ba41760419863dfe877537b8e288aa8a680eb28819ee58753a16b0
ze26ef74bb3cf13657656589df4d8a1942def120f7ed27c4bd3a04e64559f61eff30c67c3ec08e4
zf32675e94e6311cf87dc8f5f55c32d647209df00699219d768104ea2afd2d7bae17ae1a91f9b8d
z4d77f1a763084c233e35cd2f35609fa4715f2a781f61c2f12ef9890d9c70b16518251dbd496b5a
z236132b7925526b68295edc0c3c40275692c0c0037a6e5c3e2559adc0bf5d266972c995539886e
zfc84e3ccef927e9ff444b01b246ab0ef4df73f67cde37c74cfb482ecfd3914597dcde59e6fcea6
z465ffa2d4665617b907f7106ef5bae18d7dec8cd18d220bfd12ad277eefcb4b818f10a8d8278bd
zd8ce27fb74a20d14ef1dbf729fc5ca7ea44af43fed3b44d4fd9df5d0fb8b71fb3a16825912cbd5
z787001accc303b40c8dc32cdfc5f25536e673ced12333bf73a8945c036e98733c3116c08d87fa9
zcdf22955e7eff89b1de835cf3879aa5d81b82a6a83d87300cceb796beb595ab9c665962960a38f
zf064f8ff5d060fde3321d5b718df8ad8afe57cf9390521add87d7b1e722c4fea8901ec5ba6636c
zafd6cfadf18f068c6173b5b16738d1b18441157f2d1da7432484584019df6e2f0a642d7934086e
z64d1271badadb7bb3ea856c5480cdb04b767383cf7cc929940d34b2c629d6c5874673202c707b0
z3a870171029b42421d3e8bfe2dbbc78ab0988c9f0eae98d56d49d81104b7148d4c0650f9370b8f
z6d1ecab8a14860e0dd775f6eab9530fd25e349d2219a4164a2cd35f2113e02c61b2387efed344f
z8c699c2919288ce165d0e9661531d3e3eefc9fee88f94f442411d76717195dd534be9d56ba2318
zf215e3e27258c18c9426d32ad1cb8231b9fd4c9c11fdd793f99e5bd6fa7637a7aed57f8a78593c
zbcc38f3af81d905ccd7995c5b62760766693523bf92947abe301c8fd42f3902237b1a1cd44a2ec
z4be915c97f19815841cf1ed56cd84219b7807874310518cfc1c7891c52f7b091e2fd29606b378c
z6a583cff499fd0ca5fd27151439fa4c6b5ed5e876d6cac7e83a6123bebffed91cb5c74f54961d3
z65cbce306e27bf827731aef7255e3b7c87c563ddb35e2a6901a1dbfa21720e9e566e3efacfb63c
z58760ce21289bc83a43f9aed37ba5caabe2e1d9dec0d130a15ff33d29644a815d1d0324ed3ba14
z991f465adf4f5d31ab349d3e5bbb168c69057fda1665f33c790619cd68beb5f5c1c023e3ae8d53
z0faf0652cbcc019ea7dcf159d8d319fc0c592ece7dd882ab84d798525b79d08b6944bb4a425e6e
z3e2314dc191cce9ea33dc374985d9846f87a83ea8ac643421c287db59c58f2e56176109a33a98d
ze0d054b2146e9f35a6a71dda2c9ea3a196e72eea5e4441d7cb43b4a485dca2f177cd3c2e6239bb
z6f545abb584e7899e26b071139425c2dd89bb5523e230130ab3312dde5390995dbbe8ff53c9a69
z153f6e1da1003dbefe69e30d55327861e2b635039f97151d33fe62bb20f023f888edcf1d49e8fa
z541c850bb6439787113e4f548aedba0c82c4aefa6c05a5411060e71456f78c4bd836789fb0bd0d
z9ca1cc389b79228ffcac43751f4496cb11c7434c750d3ef50db59cf23d223b0367c91411f3b79a
z189b410b3fcdd8d1fd8773504157bdbadbf0aa7ec7ad759db5b037a25cb30f7a0ad47cc2f4a0aa
za24a0a6b7536800b8ba77dfba6155a7d55f116a36e1cbd0e2bd5a1da3e431cf14d3e9ac63da0c9
z3b6c1c7d3d258287123543485c3345ad529fc21b1004104e62c2cb3ee4744961bf9f7e3c83530d
zde35fbfa0bec5258e22010bc3a93db42187b3b5d404eb3460275007370963c97c662765d48a678
zde207bd431afe6517a6aa2b8496cefcd36acbb2940c6e5022fe4b87303cc9d4389f412cba4ccc7
z010731e830e1fd813c7ec85b9de8664b60f4b1b999f3dc3d8f97e82901dfccdc6af93678f39c81
z3159ad4bc0e96c3de49a680c19a865407107b2687ccb09b301f0086917196aa60a5f7e4cc11d1d
z7d3378811b7efc8dbe41f85128cad43a6aaf1662461ce6fabe8d7cfbba4d69b941e8a5b894aec9
z156ab752f662f6e899311d33df2dba4e94b0d3b6fe49e26ec55ff9fac2cd99ccfd9ea6e46fdfb8
za3a6e6686d3bfebe36424d547756be47246dfe64c535eb2d855836a888683673edc01418dba73b
z9b071cb1546db5a484eea0c5e31821950f630552e3dd7d1db6898d1cdaebe11db82b26e8716ff2
z9b43791fca457ad0e094f372b19f4dea8088e6de8f34a44128db3ec79ab9cdf1ba42ac678d7daf
ze68e1aeb7632e2137e4f90743e0193d1994d2d6f3099f729481531359e348699f7d49fc356abbd
z074714ca493cfdbff0a3ab7de9a4aaa6c1f16344f4dd71afeccd6458c4306ce188f3720c69dc5f
z780d83faad8874b9ea76cb73da02d5d4443d5570a04efeb845ef5f49fac0b359ef1de56c5eeb66
ze5b2c6054842f3543348b041ec2b47f6eb0264d10793f5b6f41ca341dc6dc9bc108c436ce934a6
z740b2f1853e64e42853a811167c10dfeff1324ac4ae718e5b6023a2fb22fb21af8fc93b7bafd2f
z41d54baf21d568dc053b7a20f16ed459c3c173e0fa6e7b5133f062732f76b8da89fe47932897ea
z518031718eac4402504bf4733b7f2e8a00393e7eae192b6fe5ecde5752215620152708532ff70a
z3f481df3010c651ad514f60a9edf8fe832e60574186bfe30984fbc3bc5f50bbc9d8218c860ace6
z0647ba79a04e0a7f69d658823b9beac91aec5410beb5e63f287f721c0397df1938c189bd3bc59c
z0e0b88f88e9a172cecbe717a7fd75325a95cc8bdc328f6989f7de0775add5c1a3ac48d5a4dac7a
z88d1b30446aa01059dd414accb4a461ef0aee6a8d0f08fd9a52498bc9b8ef7ff020d520fe6898d
z8405f64e81531ffe6f0c099d847d846c9015fcd8bed2896b7eb088962ad63515ca5685425a6d6e
z28661277848aa805e8506782b12778cd0f43b027077cc2b9c3e250b4002056237995be9a8e58a6
z88fc30e1ca45d1cc4507ab548cb8b31b8f61f55e9e26b1e6b82ce59fa0dd572cfecdb3c2e2a702
z00700d106ec3fb1a1dffdf3def249a6dc49fbba67300845cd246a19eb8beb057848ae5bf085bc8
z66b0f954c1cdedb2b166d0b347a454ca6963cdbf71bf1e018aa05aae5d98af5f8d86cde831caf2
z9634be468de266e6a4305f91d093e521fdeac77eda06dd5e5f21bd106e69766998c9e9b4eec8ff
z51b72fa7d302574d6b8bca93c49cad49bd22c1dd28a13f82004d0f746e91a36a8b2f1f9564565e
ze132ff759184045e7eb8b49342eab4935bd371e1b40d97db20e56249be0b98f13810b7f33dec6e
z28f1f76432c0efb5fa16e3517e2e827c827781374a08517c6e772b9875177818d28f855f5f69a5
z1635c99b4763db0ce401a4d5b39f093e6a7ec6395e53117869b7dd96d6af5882ba4576729d5a1e
z48b82ba58f567a264b3b9f90a2f4fc1f29dd932f8d03937fd2711ffdafbd39fa4a364161952683
z733efcc3419e6175fd37d45dd18767bc4b0d3a7d3a26fd1b956f568d50345e077f983c066391c8
z55ca69a54226b37c9c4adf8656448d37ae6760fe8561b4a1f114c0492fde00381cd929ffd495f1
zb64d2fe1c1c7011f397a7a626ce11f6b99ab8086395d0b86d310997778a85d35d2ace86902a947
zfd548edaf3b967d5a09a784b13a8bc1bd6829bbe49bc6934bce34583b463b61b7b7fb601aae818
z5853efd90ec8a97a0272447a11b80cba47ec575dc920fc7d078c9e421c7df656fdea934a3acc10
z9c75193fd0e31d8f3a7bd451b8ce967c2ebf060b5354de524473579463c151cbda81b358ecf5b1
z0d9c47fdfeeb871060c65af3863f02c594b8305e1565a52d55a7c4fa092d6726ddbbc026f96017
ze5f36e07ba6289f741a897b27defaf20b6604ac1f397b2a9f856195bdd524a8b845d24a7088b4f
z9a1fde89b7a13bf823af01c3382f19e92cc71e77a9927c40848712e881939fc6a7c3b7f4b5d26d
z5dd63973ee5692decd331f595d6a3271bc5f4720c074a61272d63be101e5007aef4f6ba30e20aa
z4b808f0a80dad79cd94b3d9ceef3ac042e3d7ada6ccc68fcbdb5736aed47f789d81780dabee3ff
za79b63b9ab7f6e608e6e5f08121f1d429f864079c5e815b54375fd7b935f2237490f2f226076c8
zd93645d181f9a7fac8b8021f4659dcf3f9d759bf7a7753b6baccaf9956ef7fb2d7c35a02daeca7
za6082bb15c418440fce829d7a07cfb889c29b86d8bd665ff4ccc7c468c586d6e7be39ec77011b7
zd3d6d260dd72d8d7818c33da3ac9dd1d7a3f4a1130d161f2d6a72fa4b6257e34333a1ed0c7a257
zce0cd90679e1c4a1e7b054e3843f20325633b20fcf95a850eead5accd5adccda39a04b94285906
z5ad9465d741918b41d24810966288b2d808aeb9779e27f025a99dfe1f14ffa3ac419bbc926efc4
zd8d42b80f684efc2705514b3213e9eb1db5c440754f31c42eb453984c05277ba063a5ad4fc65e2
z23f09aae8b0d54d54f3657d93a7ed1dd0cc1101dabc7e6f19de42704ea36bbe5916cb700de12bd
z2e08cb1b012d2a87015b2ee6c73b6554a8c796adf1bb432f8e7363dcefebe4e08eac37689717d5
zd449e0dae0331c83e470b5968e831397c67c3fb79273b44b0602e8442964d2499075e0b4ba780f
z5aa19cd6d49bac79737b7a21abe01a8cce96cab70621561bdbe93d3240ef10ac21a2a91b509c7f
zf9ad7d973afb2763b3e3eadf96422e040e4cd63669178613e2c06e3ddb01524380bcc8e4fd8b89
z680efb765d5cc44848a240e616e3b9d5d05068061235f979ce548428739cf46af7c95319a40c62
zf2aef46bc307964dde58a68ca7e893fc50c6e1fa6b687ce30269335a0aad9b10a11a4a34be69cd
z3685e4eeda5e11c3f475f9f62ae5f993b19e2a149bd8b0ecf271af079adc6471e0889b4c2c12da
za073e44d2670156002a3382035d0609f393d59fe2caacce7c03dc41d75ace3ea3077264686558c
z73f8780e433fe65265c8cede88dd8c42988c58903abbce16673631e30b07074e9b42e2ff88da4c
z80f9fe41a8cdd1b688bf535f5a5c2dea74ac2b08533f0bc913c6b961083e051395663e1839c0a1
z8f33a71291a01173185bbf7117cb419680bf07af20362be08579364a195b12b4e3c80db41d5f33
zb7a6c9c9ee3895024179c9df5faabea4f652e16ac7233421f6fc02da467be5c5da59f6c0212867
z5abd9bd040347c0197bb3fc2368669dbce851cb44f33ac34c9c446fbd3f6f27367eb823ad9d6dc
z4e3206268082cac4588e89b20bfb518ff49176b97151365fd0e58def188fa76a41ffc2e6586e8b
z0e2196b8cc111ed6ebb7c810be19ebe8e82cafe59cab4c33e6fc2834ed072a0a11b388f695db4e
zaf93cc55f75719df1b5ed6570703fd859feaf04660931b994953ba37782f1f668e6626cf8733f4
z0c7b85c8fb4b6ce353ad17e9c38e936067cc334b3cf850e581dab89a8b4333246534efc0d87d6f
z77302c2857de2b81a7c554667c3be126bfa9fccfbf120a00a390a89c16146a351c970fa2c8a818
z36ea214e21579e763c6d307e4219c79a3c783951740a71bdc6212f11b7de8b20906f6ebdd22eb7
z38d3176e004d99c29691b1612e7c108fe3abd14a6c40fb570cc28f7fca4821a5ed8bc654513c2c
z447538ff7e59c60eddfaf8f7b2a40128981412f2ee0a3699aa090a3d213956eebe281d05f9edef
z1a2c4bed38b38e0e14419fe92c859e0693949d6a0142e0e8ee6598a57ee57375b289a7558a5127
z6a34b866aba3a64b8b716a578c2db13a1b5ab5be1c4c87ed8bab56a52858f3933b15b18d07e6a2
z303c17c33e2430a943f602caff101fb5c1d39527ed8432f373610c8e79576c77f1ad9130de32f9
z82cd6ad2f4b61f10710908c6f7ffe5779058498d03f34fa753524715d2c198de31b6b24b271c8b
zb055b24a4c7c56e37cdc62faf0ce504b39300bd1af703bac196ac06d08a138509f2376222486ba
zfe8ed37f5318f3418baefe71054557f34259157011cc36734838da9472516219c0cc76a0999150
z7ce315f284fb95433717cd6b07f769a516d336a316343e8859856649d0fec51182669bab5634d2
zf55d2be048481b29271bc6a8454b948f6def5ae5e6b4a7196895387d20c59b1f33a53ef94032de
zaa06f5ef095840ac99669c28ba2287a4bf134193c74201e01490a0fb531a3cf1096026d327b0ac
z7ba8c15bba178e74113d52711ebf4381870cd7d53801ed319d9b79af245bef6996636fac8b720a
zb2d1bff6684b2473c73abd1d8efbb3b3d83c40a40c1311f1566435dbc6677cc26516c8c5c7e4a2
zc63a45bc524505aed6f0ebc0ba49b7d01d1fbce7154d86ed4bb26e8dc56ccfdfd491b4f5e2f602
z2d570f7d6d69840bf35e8a6295ffb96993d4ef63d4edf5488c2b93150735b1cac27b7dcc4b646e
z35c698c654b9e1ea5b6a2bab6b123b598fe8cb96325a7b28754e31c303e0f17fa48d9f6b9d0922
zf17f0def7e586beb5d8f34c97c57eb283adc0f5c9321d61c3e8de140e91baba0293e4d5b68dd15
ze69dd63b32a9f1e013ce2947fd77ec9169110c26a53a739db3b8df0ac806c5d670a61a1b82af02
zeceb3ee2fea6087857fc4db053044591a14a4e483685d7e6b6906a900e4f63a4629b4ad45487bc
zb279520c3efc975c99d2326ddb3b2070f9fb4d39dbcbb14474164aac4f273a19db0813baaffd7c
zae2fd72e1a105fe83c545806cfa76c289ce4efeced0ce305727851e869aab64e9e0a10fc8952cb
z82f43f9ab10fdae239aebf57abbdd0bb39162d917756a89348e40961981cf675066bd0eec15c0a
zc13df63b39c4a0d8f67e71f80def7dd1808b5fe72266d44acdccebb7b1905b55d6b28f07b9b76a
zf5b00aa70bff2788e4602bee93632c77e2e7932baed97529a6f4de366e223e6e8bb9d236b8a793
z3a84025b7ac3dc1bf3bf145a80f346b18a39beb8297655a1d3a68044324ea4bb3e34da7b8514bd
zbbb71b9776d7ff98d60ab0d64fd9955c4f23640e580e9c48eebd500cc7e91055befdc9d27cbd03
zee8da5d80b3744d688dfbb9fcccd7f915bace32fb8b3164e074fa15c117b45bced48750ae0d28e
zd4f2e67043dbf6c502bc9e2ac7e60b085d3c9be6c696bd98365d5e4457f42fa061b819ae37b47e
za5da9d6d035925276636c9eb2e98ae149f57af7c25b8aa9636646bf473d824c7e10c51077ef21b
z21c5da955771f72e041cd88c03defc4a3b06af4e34037d5551bbbe55fa98d13f736b9d0b3a02df
za1478a077709b723863db148b9ae74d6881c446dfc9d304ddbda080fc3a32d81a1a87f2a39df7f
zf5e43e772ffbd6e26904a74f0f02994b87d2a1e4687344e3867ffb137d3d4d691f2ea113c2bc9d
z0e2baf0fac11c02404bc52613804992b915b8df147e01e4ab5d568186ae77807890698972c5285
z5750817553ddf0d3b0e42b25f5c834d4680f7af14ac0fdf4c9969c12d91616aceb98edf251b978
zb8257aca058446d630dae2bc32781ae55118261dd8039599e6960b0b5782c0b50e24087b3686c6
zb6f9d7e7f1ae5718487d65d72c8d9dd3b99acec2d7147524b2d820d8487624b9434f0d20aef879
z02e0927ab174d1363e413865cf98a58bdafc9b9c75bbca640c28db0173c04d1b5a143bf6fe32ae
z9dbe9eab5d7edcd94547b4fb6386f0d5df14904bd323f0bcf250647f1fe2e6eba542cc20e84a15
z9cc9caf7214a7ec0a132750ee3e963f9330e20767a1210e5d0c28299bf97ce35ac3c8b0a8249eb
z84cbba8289bb34d9cbccdfee3574f0110a0f88b9b48ec84660398be0726c5ffc1fc6dc2ba895d5
z3a0808fbc6ba9363cf8b72c2078ab64999fd531c5e950a2550577a7a413e70f994e2888bff868a
zdac1088b170cb74de3517549b464347512e8ee51b1a4df9056159071385551e9d14f057b57cc1b
zf7e182a6e0236e1f412daba0386e09619c9cf54d65011db37f8d0429c47e7a2f4eee0b75fdc2d8
z903b8dfb9773e19c700eb2e004d20aa210261ba8eaecc7425eb565dae0a51bb73e0e07e16f594d
z7017ab835af8cb117d10eb86ed829be0b206f74b75dfe859c8eefdd60fcf25649077a295b37e35
z20d7671ad98e056991a19d306c886eea4d91310b97b569190e75f9fc9cc2bd4b3821cdc63d6ed2
z6e9993a94a1fdaf7e9db74372480b733f1d6ff3a0525ca15dd23118688c03288b9892310b53123
z075eed976c0918ecea590e6a8592b86d408d8dd827743d971842ff314ceeee294d0c25892325ca
z9b164667c10cca9f4d2edd62316a4beadfaefdc32dd07d33decaa494a28b5ad3a9e8f960a95847
z7a959da76119d3460f59f202513892a758d29b14e419d83e9a2ab17e7ece0ca39e868749488192
z7db9447943e2d9fb635bba398bd7738adb2200c04e9124e0864d3d918d6cd023c111884e8baa11
z133b5c2f1e5f3fbd3755bda6ca8eccd73bc5132eeb98d369b17a23173b1b4b3fa7f5bda4f13df9
z6d342a035c698d0cd29f1780ce26e8b16b6e7d8fbcca90fa83393e596ca90174c5fed7bc8b34c0
zc6b8c0e0588964844a72ec0ac08f7232a15b86cf48903a81864eba3e770253ed6a179c06dad275
z06e25e8135101b4165f2259bfb947a37a8fecb2e8e1c7f483676c71c1ee45b312fa74e445cdd0d
za7a3609a82e818386fe392c9a4a4893db5313a625b0495de03e32a80ce6a41ffb1969a14814f55
z7cf7548313791848703ecf35e580178538623387da18ccc389edafb4b0fb9299398de991c6d968
z2dabd5ab9bea077fbf89cab60ccd9f8805677f6a77c2c8e8418aab58e9174adb259c0dfea56f60
zdc3043054fecd62786b85ee6472bceda8bb28498733de5e016fe981483944d73285a1c4754d570
z843aeaf515955d51491bbb9564fedd94991c9d2880cc5c38945b618ba8ed34b2069e29d66cddae
z51d7ebb96e90f35159aa28e498a52922b379e7b6a30e6599e1b5eecfcb1545848a19fd602e707e
z2bd7dfdf217de2e93a22749c812a4e6fbbc839bda6db2cf44ab0e0e10056fdef895678b77d2aca
z8f8816f8407e486230edbd1429331e2e1b57aee453c1570d9696d41b3e9e596d481aa9267d262f
zfc98d9c8fa3b47effb437312c1b812381b7de0a7b2e1bd94a8bc3940a68f1054660b62b18b1496
zc9f3d42ce804bce2be616a2bea51c4a9ff3c2c890e4291d94f04a177abd2f94a4dcd940715ed66
z3a1ab26702622f70584522bef45b8df7f636b5f7ba62ad882b8735cf215377d1b2f1da2eac6d5f
zd746213831ab84f99440445778e182a7eb7abd99115e040fbb08dee547b0a982857e32f54528c7
zfc77082c387c686a4018219cc3f685e7b9a609080349b2e8305e9dbf5d20ef28913f5d3bc61904
za743521ffd019ff109f7b1c8590dbca6ba2b031011eaecad48afbfcb547b84a68bae98d372d951
zd3be8936da842b5782515bd2be105148fa80e55f6db96c7309518f8b99e3ee930f9b890fe374c1
zc3176ceb96005670f7279a3151640c494eb8c80f7415ce06745782fd9d9eeab3c0fc40df5c4d86
zd9f999ce70a301a51cda3b34ae2d3912d27cd9bc5a86e2ca54cc286f06b121a425f1b435fae94d
z25a0a2962a84e2ad719cbefab68a5b4f9a1ef51d1d98610d4c89494a1900ba466c03bd499a5422
zf6a863a758df6b0fec3288cbd19a0a1475bb70a486b11f9e25f506d3387b20931288c393c3b72f
z1a514f33bee27adcce601e22c4f348f4cb036fc4517f8b059f6c39d3157052ae46fe23dad6857e
zc809f7834aaa02ff84fd484478cdfc37de3d66c6f284cb84038716ad66f1edd4c14530335f8de4
z0c42a7a062e2a68602670df863e49dfa426cc198d3b9b3074a738df7d01e553b3e2e4f9ac880ea
z2507d57080a4cd70d574e1f27a0cbbf38d014b8654d06e72fc78ed65c0801146e6c711b413726c
z4d532eefc24f895e7b4440da97435ee102f8a19a6779ff99dbb7344c2273479898ff8573582c52
ze5b1038f3daed0a36f4642463fbad17d49153024c14a31fb975a8ed76d8d1b74ae52084b5a2244
z83c09da3df18e4b01c9786f7d945f3eac197c2e4e5ee5aa45eca291a5d0a92766a38195bc702f7
zaa4fdba66372527d8cbed8140650563b006fe391b7126c61cb3e6611358904b520e8689e95d8b7
zcfcf88d9f85b87342ec86481c7b9a5129854c79f710bcc1610509ac582b37874ca480c8f22a775
z33a83383b967a571c0eda2f13281d6ffaa9b0ec417594ebe449d9926a5eacc253c7df604c2d3e4
z66376236cc4699d3539f8b3b3a6f88e7ae907266cc9db5ee8d35f9e1d04fc2099b6b66f5a7ce7d
zcd226f0edd5fd106c012f3f7d32e4934123f95017cd5fc6f50598710117b128ff26a046ceb2af3
z10ca392a1b8726b5632f264aa62e6985b50d47b361341298a2b75172a0f06ef46902fa6655f3f1
za67191f048f091422f619704d15c0c2efe1060c1133ee59c074ae86282870dacf80550d4ac3778
z33bfb3859c6bb5090c1e8413380d3beecf4f8c61d3764488c02dac5a2b7418521b52c3c14b849c
z905d6a2c348247f6003d0212188ea7a65e0550c193e2e61b8c41e17d891eb2ae51031ba7e95dae
zdf1af08131b69cb3ce518cad0bf5d7782d8ec9772b0efc2f3499c9ea38d616126590504ee83b76
zeb9cf7ffd04c2d2dcbcc08f37d657afacf264e714171d1b6b688ec6fc228be3d57d5cb3f7fb4fa
z3585899a9f0b6496cd650fb803fa409b4b27c75a881bb96b58cb6200d0bd46a7486ec4389a1c1d
z34c314496d0facda8431f8ebad62c275edb6e53b7187d01a78d4ba5cc2f43d021bdfa75a3ff54a
za4f63f1212efcd7f125230d98a6dcfba872113ff0d6207990bd8d4adb8a8f459f17005132279d0
zb67178c883bbec047e048f3104dc16295e39c6f16ec2cee2bc8581d4beff94e9c51b5aa229fac1
z7a82a58482be2e9bfb7317beb9996eaaf4cfc75082b8941935cbed51568d5291b07afb122b1d7a
z2c3d30aaad03b82f9763d1bbbba135938c586fc81f63aa1c37d442f2348a4776c130066bd4db0a
zae73163b1ac5f2848e9572b82085c27d76ce0f2c33817d85a4ce0ce4731d394f427757b7097119
zb4e715c04fa95eec114254158c158f9a796cef4b951de1c8a2e5b2cabf57a84a79ea80cbc85153
z5345e3ada2eaf70f547779c73b1c0b56cc34e013c5f6124d727d4e4c1e9726659da1f66f0414fd
zaf7b6c52e05cc0923c7c2d9dcd36e19fb8bfe7a6e1d0049c56911af05acf799780d82e2f47f5b9
z0bfa967cfb13fe73640c4247111a4c20dc50c66dd7a5b7233a1b6ea381243d959372aef5df1710
z421dcfca3e5f84b3f0d201619ade0f77df480099aa9560d1cca4183584890e46f73764a6f1d096
ze674311b8de2d5bcd7f356192d6d3b32f9fa77de6da25cf45e62748b938069403b07f0f56e5d83
z1b291e205f4c508079a5c08deada2c6de9a2229c09ce0c51a9e628edc93d9acd8735a91d53dd8b
z4b20a0b23eab6a3b23fa003fa1a0d15a30b4772e5d0bb72aaf53ba603a3aa0397eb919c134fb60
z842c6a8b18904c3257e7af1fb8b7a899b3b6e3fba39880ae3cdc0e75268c471ac0efafaaca572f
z2ee0cfd9ad2c33de81e621e67a6d4d11efb9e24677bcdac87444b51677ee726ce217a540376f0a
zefd39f3d799af3493ce152676180a3f996b28891b37331e264e5fbde48b7dd90e80a3de3dbc26b
zc3374e97771838bef042522b1871ce4c0441aeca01be1f1c52128bf298599124101c380dce7810
zfcc7b13ef03420bc47e803fd8e3082b33ed1d24f2daa29aa27ac571821b9685fd389474a824767
z4f1e4e2003c337b0b60494861ab8346301b6590496a17b17ecd8464cb2ca890e3296d59c0f6877
zcb4f9c7b2ac25636b5387e6a43e1441a936663e6e90db80d9bbeae12e5f8d2cdb308f41a042c60
zd74822737ed0ff2dd693db1b31c8aa5989ed70d08d77ad0721e0a5947b5f76013f43cd21b27e8a
z4c88fb6858555efe9444329892aa61bdadf0ab2c751d14157b3f74bb232311ce715aa2b453b835
z91c809bc4e876b9f0f20b302e8b5a4fe9288cd5f8c7c55e7c94cfe10b1a6360cb2e3741f556869
z59fda1e52ab349f72b81e0ede6b632c9ac6d0d25f984fd7ad99fac3b8d388296f7991afee24ff0
z2b747feb33266691564ca006df395123f38c056f949a91a9badf54b427da00bed165df3326fa18
za074ec4c01450ae87efb390bcac81ec22bb9c0c06fcb055ebdd59956e334dfd73010d85813cda9
za69788d35829d94ae3f7d7bf29ded4aab69661479aff7053208902a40961f9046d2e624175255b
z0e85fc389fa82d91cbf31fe75c9780ac9e5dc0f63cf90e733cd827c4352a173f0d16263af79fc3
ze215ce782874b1ab5e2beecd390899bf3080a129210b02131d6224e92340e6d5f1333716fabd69
za3b891d07eb1edd951a7f3e2ac6b917a0ca101bf372c0924358981b4bf07b085a6bba973125a13
zf6e70e7569b1031f94514e16800082496c60450e4f55289c73120508ef2c5dcb478d131af76559
z24a15dbaf013a5fecef5c0004dd011d99f492757755eb4fe9c95c19684815c38c2bd639fe59115
zce44f40971afa97d9bf926e7515590452913240b0fb5ad71851dff8dac11e0f4cad0a7518cea11
z52f41a744a5a69647bdaf9e448c8b1c4262d25f5d994266aca664580921cbde8f0da41ba6232d7
z994101f1fb4efa0ede51ea4387e5ab5fa4736843a1e04c2d1f0a14320400dc757606f7f1b0730b
z473f17c9c4e86b3f1647bf6de274a1f949c9f3ec1fd9c9a9ea13e0cda5674a98a684be0df39bff
z8e9d1d177d11374d3c5c23e64fc6cc5c83e304581a32213accfd980c12f2031375914e6f5c19c1
zaf53615501eb0208f3638b4ff0452c6328b6fb81e822d161f8a1fe36417eb56d683d1ab5414b3f
z644a4c1439e48a74f526034325504273a2fbbb47744dabf3dfcc735455250a88b5c3bd6064becf
z49398836e808f194f86e2fb18f956c5a70a5466185b432e2e96d62d66d67944135d86f46e8ffed
zd0800c1be1cc6692334b7be158d921c7388b84886fb37e8352a4653f4af9cc917cce1f5b61159c
zeb5a62129dfbb03910f63cc5062307834e134e248de7a96d18480e30761de7aaa93f5c94b4d9f5
zaa60a0932ec01b3dd7a5db47f4a2eaad099ba2dd158f75c14c643d2d8a85426eaf5fa23a96e57d
z106046d9de4e08ea73e957ac34d5c780736cd3e9d5c36487c1fb3f712b5bd63d528a1ad52c3992
zb6e1e75e6f728bdffb08ee24540d618f63b8447886a35fddfaa3e80b5cdbdfb1c999ccf9ad6288
z136628e4af17f74b5cd222975b2f676529ecf19efc122469e00feb48233b8375a597a305ee2daf
zfe12f58972aadb09a548ccd6a045168fbea2a99aefb37a708987d5fa42d756ec52c67a9ec79253
zdcde3a3130912fa2fcff5d399c5e8d967c7f8ee95c92295f992e471ff92c4c3ac744d81180c76e
zb81274d0851f9d6eae77c7af35d437f347620d5e025420236c8977b23c5d7cc249143efe132017
zcd73b4ef4ded664015d2bf53bab9b26592c630d0a6a2e6eddb667a1ba96ab5ca33a6ee45a1b0fe
zb711c5a33f1628009401ca4f0769dcd22efedccea1d54d8d564c6d9f8a63508df964cffced0a21
ze563fa17c58bf4cf1d3ce1c4222486f6baa1504999a3b2503751f1e31868e2d8eae7db37f27ef7
z7bb95866487fdcf7f208166533777f3f7c565db328da7fd089ffcb77ba7721b4c2f897343afa7e
z1f11005418c1a21987d51e5fa2b8bbf7e97e5f5f526718b08e846c0d411175b1bf7b3b963d5555
z3aa609e378cb866d0e3d26fdcbe65992f2f483d8b25315a78890efb6307bb78a62859230ba9b4b
zfcc342a67fd8d5e7d3008df6e2b959c7da47e75473d0b76754c566d40a8645a4969ab430607846
z24123de61b42e5aa1cc981628148081dc8828a55e69f70e5458287cc0c97697dc45db21a8c7353
z510f73c2f81daaace2a75aa03c0d8b2b90826034009096d41a0fb17f90b7ef8d5cd891f0cc2c28
z535dae2c39659cf23a3d50bd18d32dda2becb5d2fb52971eff787523f1dcabd5d05bddb6e29641
z7232135c2912b9933a2e520a272688736e79128dcb34eee6dd7935c521cd086c48936c48cbedbb
z2bb38e17e3535032f3b08ce3f29c2b14a174b6cd3c91cdbfb28f4c1d05614dd00617ad2f15d972
z4d2cae3fd27738f7d27decd3e976b9c653f5a88765f746175f0aa938b5eea5a34dda0005854eb8
z85f0d153192aa9df4827834ab47a5a44aaf1f6172ff7076dbd472bdcd3e60a69097ba133b64bba
z9f99ccb072c19ef80319f78f4c5d134742abaa4796c256f07366c253db3567f9250ec974962f30
zd8be913f5badc2506bce8c46f9866085ede449cbda095a028dc465fa18980c4cd24b8a41945ac7
z68a1df6bfca497ec75a713085b31f37fd1bc232fd04e3f0a5a13b0a3e95f62c71685942ceac995
za86e7ed78139ed695ab202a573fda089fab594469ba4f09a920208e37274f90a69f782f4860107
z4f2853d71b7778f8ddfceab9285c2ce1bd5b68c056395ea3919d40caba52288fdd5557e2d205df
zce6fb2a550d3e7b1592f01cbe3b9e024c4f16290de4ba5a7a421b21afca9986ddce26e7375e0c4
z5d4b18c4319b7b7cb0d1f2b06b123625346d9cd77cd3a413e6df457fa0b01d0a32991fcc2e4a9e
z326e9733d60221723fb211db7ef10cf1a36f166aa28338a269e1c3cd11aa02862a8a2d72b722df
zd966ba149d25836cd65f33a2d1a4d466541f4758bd9c5f95925645f8feff2ca879d4cf28713abc
z8e962886ff2f20a384052b1690de296189cdf44344af7a6714563dee9b0a4daa2e02df0de6037b
zc805eea2f35c19a730d68a02eca57c6c8d96ed445e5d9de0719ccceee44cbc3490692fe70fd72e
z9bd656c3c73c8dfc2c5b28988cc045c4acdcca91e7260a993b4b13646d7ad66b5a00877e4efb79
z344ed6d4687de9b53f3c71e2997309f35cae1dc3683f286efaaf880006a13e47276499e80e6e8c
z058728ca5f240013f77751a138aad898e77cc0c4228fad5926b71c74188beb6a8de90df38e178e
z347ffc9b5fc7a1bfd300fe2a3a742d148db1f03bf4c6732b4899f700176c90c3eac1f459fef1f0
z7018fa20217f89288165d6d6266502f8a846754a156d421de178b01dbda30af3cf1b171704ef98
zf1f04db2821a7a218c663f241af5cd976062439661005ae0241dae00d822e7f7b6abf36201ea48
z75052713189ed80ef57157b670efe27bd6a96beb0efce1d5637d964927f1f0c486d1773b1afab3
z570fc1fdb343c1eef6e07ed9d6c2a7c4d0f83588e5439694307ce2aa2903825a769856305e57f6
z7b6ce24433ee9e31d9aee016cab976639e0358c9996f1b6b9fc08992bb31d9b5297fec8e9ab53c
z6cb44fb42c8b062dc01ab4f480b7e0585d44692d7f1793de8b8170ebc0200746c80703e3b74be3
z4989a561fdb988f93a934e45ad625159caa50788b7dcb177cb769054079338aff3752173e34e0e
z4dd0c58b7702b07709e1004192ec1dee9a9c118dc9c6f966e78e457720c727b57082f7545da801
z632361d58211da5bc88266ac46453be819d3e102a0049ae834123eb871c9a506859607b8445d0a
z5b4b14c45384cf66ca2915472252f218b0a94eea7427e482890b8108cd749d4f7e1c7bbd3d5a44
z3a09961ba02a2d47b4ef87e272f995b2be42609b46565bc25301eedc2d204e7b83e1dddd39877a
zc86c7a949a8505df3c8f72a272718709a813a6e31b214a65dc2edfa0e87fd8ec2700d1a976c8bb
z431a1e21523f6f96e953934fce6d6b4a485b382a77945297ebeee252cc1890ee8c76394604d299
zf1e0e3fa6ad77e7d418f4135a295eaf44945784a15de041427499dad05722c840b368d3294ab8b
ze2364e935a496b463792a87c4b177448c66311d31f17902d7419c1651be58a5461fb19d8b77582
z9207e1096d6dfd310204b66f5fb84be11544ea03647f265f6015c47688f8424186f5febf9dde75
z36513a1bd748da4cbc785c5731a0b96b835cdedfe1b45c1cd578c12e0d6ccba87333b120deb229
za9ee149126dd2411bf4e6962905342bec4febe0d635eb60eeeee1206881f2a2f94802579fc34dc
z7e78efeb3d8ba9d643a87cd62d35b4f2a149267f26d697c2d9a90304240e45bac27f97e916b70e
z2a0e0dd14723d88e431a709f9237aa23615f5516d7bc5d17e7c0663c1fc0a6f57c18c1983d3543
z7d54de1ddb8c6f1c9a18b6c78b2ccf3a514194dce508531760a536e5fcb5cb7d280e9d20b43979
z889a172a6cb069cc60c8548cee84c41b9be8fa2b89b651c64f1d220f8a4be987fdfd969fbc92be
z5ccb3491ccb9c91683c8dc0b7555023655dd22963e17495d28d3b87813c5bd49a05e7d408a0dca
zbe2d937dc326d5e0bd6093eea5f363bdecd2e5a6f878b416533d7ec0cec4fab3454abd76df3c0c
z5b017a5cb6fdc300a32dc117e3bdd75699f53bfd13e4d3ff33bb3375c8a89972d6459a090c105d
z8356625cf6f1d833481069e38ca3aac86d63c7d58c740f2dd53799982d0f043abe819f5dbb42eb
zebc112164baec0b9641da27744b15fb22957c744affb90f5d2788a0985281e5436e66650f0fa7a
zcba655f0a50b217de2b8feec023917e705eb76cf394845aafce583576b0c56c27a19e08c003b14
zcafd63ec13440668a181b7dfd9f1d1b6a3bbe233a58ad8176ddadd172d9d111d07b7b161319ef4
zaa982be2fa90bfb9f24d0ff21eee15c83a3564e9b8a9111201adb2425f9c0b8b49086e72419000
ze4e60aabfcaa286cff1dbc31e8dd316fa52ca469fe5cd154ec530f3e3d3132903b6435566ba18b
z8c75475639e07d0fe7c00c7df62e203ad4c8d43e23a5939790523da9b121ee4d202ace93535fd5
zbd070476b16b10a25040100ddd35c994eba1b30859d514a1454049d6e7a8aea28da30a0a449fb5
z9c118e71290d1b818fbdeaa6d61392a7fbe2f81a8ff0696b8a519fdcca7f084e16b7f4c0dcbcdf
zea4d402e67a15f30476a95c5bb46ea0b2d015b29af1e8bba2d1ca5867f6c3d9530c6fa1b3cabaa
zc20eadfde6adf3a3b97fbfd7aa6c87aec20d87d70e300977f033d50148e60424169a5a46883669
z3abe31b8ed379d35a38f50a63f74ac2fd710166fe89e2ece72abdf76fd7234b212dfad420bd26e
z98b8bcf0f19dc31e84781209a62a41fb6979cbd96cf8eaf95910fc78f3547ca7287393784e6174
z9498e429942e244cd9e338a7d36e2ff52c702dc7b312c9c978542fd56318b3dbb4de13d07d53b5
z43c724fe0ed3da12772259f2f6f7f51407abec5f58ba36165484442008996518ae6f69de4cb848
z37d15df3557d4a5867eebf3c5a8b1a7c779edfd514f8ca3937b0e601299a969992c94a6f067393
z7aacc5a338b77d7257ceb4937ef6a151dcc771d517870ab860c772796b2fbc50a05b25f8cdfa80
z94ebdca94be3a3c585f3c73ecae2278738a24a9ee332e72b9c7d5acdcc894944de7beb18c63a0a
z9e809e022ace52866704c7192931bac5eede129348c79aa8d1dc3ff2a31db6d89299ea81e0a8fc
zac0dbcc2444201450f48ae3d00965d7e15329a344cca0542a899647f20c030efa98b3c3d344692
z9f143c8638f246265a65f9411fc72d48d2193fe0a582fae9c69ee776320f25d58ed621b9da4dc0
z0b73152c19313774acbb079b72d6b6629ed0dcf0f3b3a740daa53b97966b4476e98ed5f7e69283
z226247dedd8bcf8c8aed034fd27d15dcade5cc15de76e0180b654c6de69b7ad32fce3deff2d8e0
zce8df0d79ed7d1cdb28bf3ddc53a2f03d5aa27c70e729c24436a071b797a9449e46cda7c95428a
zc9d79610f00afedd74615a080cf617e58d8ec3c0e4c09128e037ca5a71c3cbd2effb69156f3bbf
z66fe611c6ef9c91e0549ea66d228f903ce813de04f993249ceaf7bb1892bac481552339c7c58c4
zda0f7c262515c5a2aa9a49de663e720f09c753061cd6782c0c0b148856f766fecc8e9d4310914a
z1d5d79ab161a24dba8427f57450cf65a4a2c60ad7b3a91eed0e6dd6dd734e400acc1203906d646
z64e52996ea2caa686678c0ca092a2462494f3e5caaddd89febba7616345d79ea876a44d172242f
z5ccd2a44d3b94f406972e735affaa1728e61fb4a6ea4c8a64e8508ae17a640fc925f99241e545e
ze1341d621e0badbbaa2681a894d4fe965ebe00d3e6362ce8f237526b19ec6c7ea3c56bfb7b0fe0
z8fbc4fc261ce8c248f7fbaab8729d2c3588e6a64c8259c47334f2efe1269e816af310bdf103d1b
z9313359989a9c720d820feaf69513dacca2d6271dd8ca706b0edd2f08ac89f4489dfe7a80859cd
z569ec42002f40305d6b2cbf43dca110c58d7f714c43faa349021bdf3b788352d1678c7d4c39342
zd67af86349ad975fa70d88b4f6ee0f470905dd306ecbbac899981f01b57f13a4a36754bcf86bcb
z35ea8a47aa539448104e33f36677bf427613992f4cb8933659caac49617d9a693a3a7d15e564a2
ze54aead10f9768ee10b4bb7812479b09505290bf15b84c3ff318274ece94939688851bdfb39a1f
z0e71e7b431470cfd105865ad4d16470ffbdf2639c8a6614e386d0ee05ccc3cd786fd84022ec054
z677a505f6373e7371df22f868f05acde782bdf58e3426efb46b5bce4e337624dce9c9c0219f80f
z2c9f2a8eaacb66dca7cd756e435bb5d070ed5aaf7c2359dbccb3f86b6a7eea85045697b42fd7ba
zd5e71c19b8d2e1237955ec6b6aed67bd0975b87f66ac71aeecab8de4ae05a89340d878ffe8c828
z8cc2439e7862dc7795664136a0a0f0bee2a019c2fdc88527a5e00b01bd323abc6692c2f205b937
z6d52787c7274522e7cbdfc9cd212174df1b7970b5ad2c401d6ffb1c1d41ec54dc3001167117dd9
z1553ca087b243a849d8cef6efad7e35799f24a52c381f4e1c6e0be743c7b5a13c52c8789153abb
z97858ab5096f8db599710cc47656c9ebf6026055d01e4a5c6a2a4038cc7dad7f3ae0464db2a8ae
zb21f221e0049b51a9c267e457913f8198cae2184380015f4a63e9e677df1fbb240f3f47751b66d
z0232bf6f1509d0a0a9d903702d01db59d3e8f13e3ea7b90e18a02659b8e992699a334b0623e639
z36ebd5e291e86c5de1f5a1a92deff1d8f867f7fa49bb1594b440d93e67711d15edbf57e8d0df6d
z9fc54fcfe8a58405c3e854603f98b44c030e6d3cdd384eec5411bd31fae6c99545ed1d97ce77c7
z28272ddf6842149f51b736d3accd7334f57e4900a5610f4d3f75e067e29bf6463c1b9cd9827e19
z42f1fca02f7a814417166fd22f66dd7168e2638208967ef1b3ae8b02ef9ad7831ccfc72a24a3c1
z80c79a4fc7832133bd87ed4807db6dad370445f84e624b08d6fae23a8a6fe04fb6174d4693dfff
z4335a55307bfbf5031789a20bb79bd571362b550ab292343cfadb43cb375c0c903fac8e32ae372
z8e9b36b2a613600cecaee1a1e7f9cba5a08276e15a3972e88faea770e6bb0a7014015a8bdf16b1
z986694a00ea2e935aa6439e09ffd61cce4cce711ed702c9b0b2816697706a2210cc01bf1715349
zba561e6f8b038321d8095ae6f9af9a2e60e7acddcbbd2a1f107050bc7e782577940c522f3a698c
z0e4a239bb8c4b53f4f4d954187890688060207587fc5e97cf3f27ff74aa63e1cfacc09e1cd2406
z0f0277b9d77b7a7e61acda5d936db9a14c12ebdcc2688b6b08322adc4fb5684031e121d4db568e
za7a44fc2ce50a9d683d7d567ba78315d0f445b655b350fcababbc0b65f4eab22de94c0d01b2197
zc05161da7c42abe4a47da9cf0dbbc64c61be4d80eb70b4612a71394c29a41b925af8d8831638c1
ze067ddf52cb1ea5e3d7bacbbe10b41dd7ebcba3e8dd16712554c66e7103b1591bb52099b5e85f6
z2fd07d55de47e5f628a33510492dca56955f0d6cc5c879783b310a3cf9eb56b4b6fd5314b6b3f2
zc8293dbc8bc7c0223405742384dbb41ebd7fb67921af4c260e307371089c709ac23493d06c03fa
zc99b9522c37024c00d6c4a1008dc88f23dae5a5adde1247ae1d32a6ef2ff50797cc3d97e001e94
za4ea2fcc0e0302d6dc1a0e7eb29fd037db622a3c23a8e1cb136a5b8e68e5e7ab4e93aeb7a8b05b
z9481c740a5f8031fa43f797989cf1c51098355d14dbf77acf880adcb82878aab32fc50408418b1
z9e81ff42ebe5a20fa1d9215630298edec1b6762b57fb64f49f593c8ecd0e11f97852dee9fabdfd
z8b5e405f0bd6db472c7769ff19ebae1c2b3bd06dc1c8a1a7540035f63d3b801061c32f5e2318cb
z6c5316876405a6c5cfcca278242378d50d94ed605f867dc07eddcfcc46d877327ea0e89d18b66e
z236e370c9866ceaae0b1770cd6c27251768765efa47c8bc51566cd8c1f12824c47a2258096b288
z02d612624a2eb66301fafb892ffc38fff5581bb790d6defb53ccef20d16a16131a69c72626bb8a
ze4a3ec9c51309d51eb91ce553eb43ef2c4a4ad625b0147e476c74c503860d84fbb7aefdaf58d15
zeff31160364f299e6fab13850f8ad2ce5563653e6099e70290963abaa8a8a61adbbfa8e7257a51
zda662aa081f21c5fa0da0701c645caddd91162adb3528db2c1f20f1a28f5ac09785bacc4da0030
z3945e2fb816e6542faacfe529a830ad28aca42c047d5cd9aed1fc713dcf3af156829ba55686f29
z6a3b90f33381f38587d98527dc47992362bd9bb239ff6cbf1eb3476eb44647b49800e1a030f707
zba1bbc977542ad3f17dc42cc39ad0c8c468295d7fa55bda5e85b1e7709da8d4a1f96fd16299e4f
z14c15f7f3c05460b307ef59ba813965d9abf6eb28d0cd0bf8135561659a07e3630b5d0b373615a
zf15838d24e4ee5f8ee1105892ef462deae590510fec480136efd06de4f3a2418d805f84ca3517a
zc5661e960eb1e524b7905aef6219349549ebd8b7817d262c5b561e40058bf2636329d30a0984fe
z7966c812d519fea8512ef0ba60819a9266421d184edb41162687e1fefdc82f4e11a0e360f95105
z3448aa25a5f0631d0bfd345d44075d534186a75e8eb81b3f871e59225068ee5a46dc017a450ae2
z4f91b16a0142aaf1eea299142b60efba885eb3c71a6a791fd38ef5c00e800575849a0e7984fa77
za355a8c310e176b4d68852b91f3a55660a960900986580ca2f4e4ca2d9544af56ee430c60008a8
zf9cdbf89336e017414366453e30d6760bf3f86dbb52591860806f5f1e93987bfe2734bc42d7823
ze47cb5a81b23c69cdc2cd6e10fb748cc836fa16667f651a1d102449e7d4ac083766f9d01a2f52d
z51591b5a4baee4309d1af5774733ed1fa5d0085e2476913adfd45e00395e5173f850f19d2f039f
z8a8fb5fdba2950cb64a75aae369d97b0c4f8cd8bcbcc1e299484ff0da6865e800365bd6f31f7ca
z06019ab1cfe205c65924f6101d5d7784a00255769bc454ceeb0896587bcaf6fd2e76eed3a22fe2
z733b2d8d13e3880e76173bc6440f37339687ab1e1fb2bc8b96a595dfa10d57c33873a4f728ab7d
zbd81fc805cd1b441d6cf121b76e45a0584b04f2c1142692306fb0ebf28cceadd4af43d395da70f
z029cd2fae46dd0e6899427cb4bb83c9bdb7e130780e350392071317a288370d95880ae995a99ce
z0007205e548e95bdba0a1a4f92415ed7c0ddb89d2a61532ea344e61f5d83dd05c27d58c8fc5651
z9e5517abefcdd37e5dd70b4cb142a8411c1693d4f1259cb4f17b6836a93e47fb33cab386cc058c
z9915b2f77a21a23532b8c80292d6be70ed0d7debcca6db6d965c128efd6207625fdac5889a2be8
z56914ea58864a0d93edddf8519122310cdcd91875ab885687e4d57fbc077085c420bd113c2c9ba
zd04c5bc1c2178216f0979745947bbf338296e3864583295eb84665f86ee986d0d6a71c91bb3239
z4dd93d97624e186b6745f6cd211267be6e7bd9820e7fd053414f2bb0c18dd0cb46ee7a52083492
zb4c5f67e050a65891bb5a8f3149b042d851239825e591911b95a9f510fb3cbf4c7a82ad3e4f645
z2fcbe8aec7fef6ade27a1da88002d27e933e29ad6fdb14e3e9736d03557f6e8f028f7fa4a598d7
z83c1ca1221e50ee8b77cd55b7c1f0531b273392ce17decd9c6e1affbe650563b65ced7610d2deb
z2417302b2cdecd2a3a4ce6e52e64c6d63baf90c6a8eb201150b6c89dd7ca9cd7af154de88317a5
z91c1df8b038bbf432d6d0f37bafd861b9ad4c137a53f56d60b06ad3623c4b20c2cd717f0549e87
z4a54bee691cafdca1f4d643d0a8d72bb95b6f38e8b157357069031e77a7160a461a0234df174ff
z0e160ef267d9f5fde5ced950672f28218706cddfcca6bbe1848e7c7eecefe93de1430af9177a74
z0af246690b0b077d3e74992af6158677ed13e98a9c326a33a2406c5c54ec8adedb8b8ca45a565b
zeda1a70360d1baf68a79ab9883ee131812e7466ac44eaafb5f4b6d6bfe9162b7f9cc0a7120f40f
zf9308b423044fbbc8a1e9f436afbc092f23a9b06f2b76d1927919e53761ba5e269d56a8082238d
z5c13e865bc3c26e2be51fdcbc3e763e4ef6f947dcfc61d1fc85c5560ae9d49d3c4a8e302d96d6b
z22070d0c6f0ebdc82479e407bbd259d46c557b16b4fe05f9c012fb9f9c42fbe171d93b0c61b8fd
z46205aa7a07a11c5501a6dc24f5098a385b02cc38e917b3bad3c999bf6c27b502bf14a695c8963
zab8db116f11f2f115ebe23d479c606157ccc15c7c2de52fe122eb2fef51b1b43f399a9f6baad77
ze1ea4273a110ed6d90003aacc2732155ee19b54cd82f822b414c1e4e5bc37028796f057568f185
z92283717440a530f7b93a4c0ed22f03d562415f8eedcb57988ee2bd5fa6e27642e4027e177e95b
z7af6723f706892c8eb05476daace2736e139a7f99c6a1a37f46b5256eb923d2e017745c43c7a96
zb0716e5664b0006c1f239cb266260fdafb5062c67f04ee7c081e43eb45144ebd1ee4f28c225478
zb6857f61fc3b9093184b0e3b616e674628f29a41e125e012bea8b7d00777eecc7bcb0841883f44
z7f98e74b2b35fb415add114dd0656cfd39560d1ef26529ba2198f2ad61769047333bf49b9d7e6e
z3ffc353f6947e9b13258a1a836f76f89d0d00f5cb7d4c81732c7b644db6f2f006c457b2f8ac0aa
zfca78162955e291eeb1eeae2f52f6144e3ab83d6a627b007eb956885e0cf4ea584f2924d5437e5
zd4c622bb6b8bd331b84930a290751237ad632b44010195c69b99c6611bc60731a9351483e0a048
ze4febee6f4d31de421d502c154466c889803e686570409b085227779586e58fcb89701a9f8b8b1
zdf47c2c8069f080d430fa19c09cfdea75665783544906938229be2b35519603b1773f2619d54c3
za2c38c34833213eb04e4cc26d9e21829476a415626c6b76560264dc4423b69f6e106d21aec9d19
z9a78febb6e818148caa809f7f504104c70b42e6b732c465f6c0b6b6101af5496e34efcd096fbaf
z3086e6ee745d1b9811d5f61d11c66de2eef8eb8d304e9cd532ac675899092e71b90ad876212782
z30674ba50dd069249629f9f7b8d6bae5cc14ba60f42ca0e23ffa32c4a9f18b751875a4580855d5
z9e3ac16c2e1a1fc9737bafb6836cfc2e0a3b3625a72f42cbfe99efd4b07911c2a036b991fa10d6
zbd5f2e3a82e92c546c7b93bdcfee7ea1e1059188fc93e59b7a981285d9a88cdef15e767caa4987
zffa71af88d3950c25c300c28905648074e405f079b2549654fd9845acbecd0f8ce6c4e08d20b9a
z4ac44b280d32be9bcdf568c2f64f03a3e836eecbf6a23f52726c822db899e0c5a45af02b3ff925
zd1864372824671a1e7ccb1efc8119d09d787701f96a6ca466d9e1da2294d1bf8979377a66c1ed6
z4a9254f5fcfc79618eaa3b2af98c62d8cca151521097a18c8b210bbd4c88ca4fff92c25c2ccb45
za8c47d22b430234de744805414369947844c97e0867aa9b09978e8a4f0b27aeb97abadee575e06
z5e49fc1e3d64843a896c91e380d16c85795924e7888ff57377bf995a18e0c634bd46699d950662
zbf941e571d9a1b802f2c314a15683a853263b2d598f1c69fec0d4852ccf1d13828cc5270af7a29
z58f5b773b5a58dbccb9586d089e1027b9508b162b9a3e3d35de576db4bfcc92369eaf5578e86e3
z181b8adf936f8afeb254c8da701760ed19bbf96efadf52ba2f2b48719f99aced474fdabe0215ee
z2bb98f6a8787b090b57e922a045030bb1950d38b4804e841d0d922e05f1761b14a9d6ff4e2d96f
zff0283272aa7099fd8004960c0c5d926227f07b816e43bbe527b35f0f056f997b4298f519cc0cd
zf5f60534a613a377b857b477f8f3d3bed699e55335dd59f01fe8647b8bac2e31a096e13ee84d26
z8a06615cbee8dd1d218829768a1b57ac818e64969c0ba524d5d92838d7b7a84a1ebfd4a21234cd
z57e2559746c6c8f499bd22cb93777a92aacab2215b0e8ff6e9c40b8c5ccbeaad693dbff519653b
z8c700a6a2600a95909fcb5f17cf42548ae2143c20ff2271084973ae92b4d9525b5065b99478fed
zb3c621de6adc3de9a1e74e11b5867f80ff8c6903d8e200706de2cd1634dd4604fb02c827f797ee
z0e339fb5c606ed8398fb132eaf7f1a59ef219319fa649bfae4fb5610bc1fb81998d988280c5d05
zcb7aa15456124b6ab3809e52485d887bfc0656cd43667728b6c75148357801e1bd4388290a95fe
zefa99a572ec4e5470f55972c560d5f96833e0b862190ef188300aafaa9d88357934ad76de08f5e
z378699eb94d83ea5b192a644c06f1ffcdf9a99c28ec70bf741c74b75c2b311223b5f5ef048ac4d
zfe26f690ec955bbadf698d55c05b6325a58e77ac1a10e87d57367ca94506088ffb987be1a3e9fc
zb3e67b12a4517f6c978762ba7e561c46638c315328cf73c1fa38f905f7f268073f7f2e20c91a3c
zf2280282fea6d74025ed59aa3f2ec42e75f80cd8fdda2cb0f67030b4ae14680c5c507bfa4f2ab7
z071b1f9bef23279500438de3f897cdb5fc3beb0674c4fad2651a985087af5252d3b213fc9d07cf
zf629c502f622b3337740f1d79c04735e7ea2a141cc8a881f39be8f3ccc7a9c549cdf4df6059ff3
z8e1512670e2841cbbc9627dd13c38ec35e47d0cc91ae58e69fdd09a8945b4c480a8e2a2fe2d05a
ze6ead46ca8f6e2e5689de0dab0eea1d47009c5d3e7bd4910a93c75dffbc7dc8208cf417b089083
z7a28e775a5d89e0eb1527e0c8b1b3b1243a650c6eea6720948691e42992671538b096e36a3fcb9
zfc34c8020b45c08d1b251910ef38e8a3798780888f8363cf3bc03f52ceb9f1e99350ea96dfdd53
z93a272310b3ba6d914ad070c67b1f34118445c07f167506499987ac3fb057bfd7b7d1f88906300
z9c3663c61879ee943492c53821f5e347b37cda90558bfeae4823ff78045c1b36c760818a313e1c
z4a6f2b327f862d9e2fc40b02c68e6a6502dbba07bff23f6737d66997769ee7fdceaa4b25424764
z31bcdf3ccdba6447ef8d5b6d5ec3eb1873635fbd83057b62b6cfcdacd664d8d6a3f377b0e9069d
ze15a51e06db076d19a1b2088bfb61002e99ed3a8733dfaf36ae114c703cb331588131c80da3a93
z3fd915e014d99ee946fe57fc9b39de9177c98ea1a2616749dd5b31051ee975a6aba01567d36d8b
zd9e486811cc508eb9062b8c4435b43995029d41ff312149e834d1f85949baae80a5ec77ec1075b
z407c16a5ef0971f9c3b2a5ef0a300a3782d3584cc7d5535f3a2a29fa150bdc1fe06c8beded4b97
z8b49fe8b0394cb84ee482ba9c69b53241a1846120966d24c37ffac984893ef7c40b9745deeb371
z48666b87b72073460795ba73da460ddfa0ff1fa0304f8d395f2b7575191acf746ee30b9046c81d
ze9ce08064aa249d3a2fd2effa7574f7d75a4c13976aa7449ae116c85b3ad612411cc5f5aaf64c3
zf72f3b1b36e1381594acca836c7629ff947c265d364bf4657f61504bd459493b89f164eb82a85e
z74d49dbc6a0c3b84713aa714e856740c58305be175ae759db937717a6bf6298f3809659cb23bb9
z683ec64bbaff6b4614678d58816b6a8b84b6cef8b0f611c807892b82f3ff1b2102e824e66ca25c
z21a98d7d340aabe5ac9b8c3b934ffd75419f4df5c30fbded1772a41d793668d9cd499d5bea5bee
z78a8648767ca9bf83e79688ed074e6c51a39a026f2539dde495b26137ad5c92c7ab84dd7ce21ed
z508dbf27e02c82a54e320641e94c1210d6b2b2c7c5bcdef1b7cc34537eb59fdae9ca080d00779b
z3fe5ff10bf0b1838aabab520c7292e538fdc27f8a20036affb7fb16ef7e2dc288c884aa9094fd5
z68a480505fa75a8f627108d697d8c9891c80d354fb6173fb2b04c54801dbc0b2b077c043e20755
z5995bf09a2b3f8ecafd9d8a77a721f7cd8a91518cc28363f5fff455ff4b2b67f4c4770661bcf16
z5b26639c0db1e74b75e149818072c09a11afab04e45ce565f5f60ecf65e2d2507c3173613c3c9e
z4decddc8a1498f9cac62ffb6444e7edb843d8fcbb60f0c2049d795ecd6f18c11acde023943a2a7
z3deaa966fb8287e40a2989533f044608e6ce53b744b9021b96f4ec253c0e9b0096fa83509013b2
zeedde73bec062ec83e8f953a02fe8f9d8c66391636adc5a0f27c42cf2c74d425266f0bca9a8b08
zde297f73539cd6f5279b8c6a911f77272f66bfadd5cdd5e49d1a8ccabf6e120dd6745b4f89a525
za3d6bec57a2c9437f8b9bda0c3cae080f7792c37777b2b325ba7f88432cda4250e84064992f41f
zb799155324ea8b4b31a093472a82887366ff1ddaeea24cb700e0106762eb8cff01aa18ef531574
zf151b74408a81e3eebc81248a8f99bcf0a7c639466533734f07792ad3b5bcf8b3597cc3eeabadf
z5df54e8d86d6e113a1ad861436b0fb904c5caec548ef7d69f023ab21c49022aa38fa2eb6bce470
z44cb3a82310edc649c6080a57f5e91149fb89e9f49f10da55a73528ebefab6e928530f998cd2a5
z600a47ac5fcd45627663bc0c2d0f363edd4b26186a2cb408f6152f197ab23245888cf02ed9d196
z6ce0c442b6beecc5590d1a5a6a695a4cbb0e2a2a48547910bf4c3d85fa4e14d83af8a75bc836ae
z1851bb19947c467c5603d3bfd1e33db3b4e836b546183ce0b964140a76cbbdc12e8664e8f7d2f0
zb21f88be365859a5285d091d407b43bd71bd39af749d8c5e9270a98776f57d1ac455d886b18873
z25444b1720c922b210e7b2d44e678e0d9f413474a667812569c97c380c85ebb09b27e1cafbe1dd
z4993dd5db133662a68ca19f7334abb8efd3ef52f76b2dafe92753c01dcf7198da61e5e502145c3
z833e8719106e5b9d69f3c8103c3055929eb0617313b3c71b223c54e1861a169a1c0e0f084c8d30
zc4ef8b1341ff39195c1e655daad8c7304bba805c5fb4f1470ea5e6a5f87a4c7213f3e4d1c33f9b
z5f644e0741163b68a5d86edfcdefebe8b042b27e5e0e4b51b14187ad8c7baed5d6ac37f2645270
z42a84ec298e788f569fa0ec3507eb28842e7e173f27c8a1cd1225233b0985824f7b3770c083d4c
z5134de10d03a82a399da7bc8e9d488573aa07383886208af8c4891d35e35c836eed382dff69711
z68e891275eb7367168d90ff7ab8d868c8e01352e132c8d7500ea7b26fc7f4f75da1d13203f5857
z17c1cdc99bcb2e1cce28158d63356e5889e2684aec40f1896a72d69b6a50855a75a497e0037194
z2655c6969f404e220dd6f58d2230ae5ecc2c571b49be841e5a2c1cd0eb15cc3cac74e92f011850
zb401c306c01bcf906513b6c35c8bb90146e371d107b0c7a028fcb24fd287d2654bf71b33aed901
z675148f99fdc32893ff0e317ccfd010ae979cd64054e0c58cf4eec25cb51660bc333cc21b94236
z1c4a07bb0e96bbb8c2d49b99f38eaaddeb03a5a805aeee9b17d79fc40173c4d42fbb0bd6d341eb
z21da956dcc31e59bf8f0d2612fd9d83ab435d6679bc2aaa1d6878cee255e29adf589722180ec28
z291b949d26cccf8b5cf38899bb6e36ccdf33c234ab5a5c4ccd1db387e13617e4a9c6500a2108b1
ze044ba7a49a4f180d390d265071526188c4cf4167855a7e1ebe1251ed733b1a0e2e2b89e29616d
za29f4ef5fdecb01b33e76503dc18ed8dc818e9aeda048315ec384c3f1c1af3516f107de418ebee
ze6007170997c5d5bda22578300b3dd07f77980c83248fb72e1671f8ddc1e9675311ce59dbed441
zca4ea44028bfe72434c50d2bb58afa6f7f340c7789f41123b676ee74d259a772e77e2fe2aa3360
z56cc0f172ec47fed6cd8ca0026e157633d283612f018158355bc3d303073ed5011f9737d50c32c
z303913da8f284567cffaa079f311a06d80342d1b128a737275c175871319e80dfb4fd4cb894815
z5475fd6310b070afb39e1d390279a591909cf4c75d97a90b0079f8ac3ee9c2a70801daf8b4f66b
zb65615fb30391d30bc7c8a634fd6586ba3b2ace61d9562f3cb5dc032107b3d7fbb938c41930bfa
z39f07ed5bbc391f516bf4da215716a0fe3438af8ae72ce07a993085c26ad30051860282f33de95
z5406c6eaf4737b6ba295c3aaf1dabffba2198e412d7a71b52be053b676ffd0b7a6a74ac163e233
zb3729b707933831a33f6d3d1163d0d27804d8e0ffe4636f0319c32280bc030876993df5233ce40
zef5ae2a08adf3e04ae0fb1bd8a319a69eda14a96036eb6fefdcd445c96b25875e61f10452cc8d6
z5f8904b42dfbe411291415a39a7a0f9cfb82a8c38680f86832ef76c6afee0f0475bf81254ee5d8
zb99ec35ad71a4f406375d25df06b8664b2757975dcbd016708de9abefab64658986df0453dd370
z17453ba55aa668678c80b056666c3c09e40687ff6f80023d5253c956cf7d56c63d5721c82d2bf3
z2974f0e1675220f2058cce53bbb34a6d72e14d5486ec756103380427a33b9667e73ae715da506c
zef14e2cb5d3c088916227430eea15a2dc1ae347478c32e5f0d26a8d37d9cd4730f32ed17e70e54
zcdd3256357fc8624e8e7a2ef7cede60a3752715c5be722e8daba8022d6b5488596b2857a0593a5
zcf5cf49bb73e9c6f912d6c3b23a5edd6a410aef06844a37512a0e96ca44be24792a752e07a59c3
z9fef6e672e1e6e3816dd1693f907ff7dca444cf7f7b4696ff7d6a58f764ca7b16ef21c1220bcb8
z8c776c7e73d7e322fce22ea86198c51dcd346d5abffdb7da72615b7fb855486e927615342f18b5
zd62ba76efb9cd1cb9aab1d7f3e56a48492d396d825c9d68214c5f944f7c94e6b05f771d5aa9cec
z7efa526bc2edb2be4778e56ae4cd9b62740ba74ead3df546f77d53e018f98a3cdfef8da8f4abb0
z77ae14f15ea8a712927089195586721da80dcb357a8e00ab6ba825cdd18b6a286bfe5776f7b7c8
zd1c8020fb30a5ac2e310281d1c374216044be2eb1b461bd97a35e1c8aebd3a4f93d16602713e5c
z48d811c5933beeb34530a2c8d3f87b5904780b51fb2d7498dfeb374932b3da0a13620be1b645f8
z3ad6d43fbf8d6d92b3560aa4b8d69be41fbfb5102751054df43aa638498b6f960c791c7394c01d
zfb91235275840637fe73fd3dd36988da25557a5c6cfa05fb08ae49a674bf5d6209b79c37c9140e
z0856b6474c2e1d92c0e0123cf85027ca0518478fb72f067e3b6acea1e78c8d00bf5a853e8ca5ad
zb9cf5df9ad8e42062b4fb2c16f1756cae0047b4855bf2587e78f9ddf974c3cd8c1c3ccdaf44edb
z4565e56162316686bf7d793270d2bdf78ed5b4c5250d6382a9c1bb09040e6e8f0a1035e4f69720
za1689f6f8ca60d7c0e493cf7dfc8caac25e0bda891f73c22d09a7fa74eccc7e4bbe73c18d040c1
z2a1805a0950eefcef89667d7442efec80b23c6b0e85d883c0383d885f7905882189b06ba94cc46
z9f1da2da0f3db9cbeec0b1abd80bd562222e047bfb66babea7f837546a7d766b1513f9ed5d5cf2
z3a08f644cb413411678f3075056daef4f96d5c77c1270bc18e09dccb29a7cc1820de9b7c94b060
zd8ade42fa8327157a48bbfcfbc82e6e01608b4a583797ccd0103f41e14445b58f9e937b70b9bee
za9bb4fd58ca038d031ca20c1339adf57429c1264459d2c80c6807359a484ce25c917d8bcd6b457
zfddd1ddccdb43251dc4418f68774d75399af5bab9a00072f01605d4f2de69a903af0c8b5e411a1
z4700aa87e8f8e79e4c7044174171e6355c8876e2f8d13ee1a504d2ba920000ef0aeed93d3ee2ae
zb02955c8aaf2632b2bfba150c3390405cf34b40c9f8e036ecd3333b5d6eed9f1ad678beb7dd289
z5764917e7fdeed99132d773c4728a3f0f0297d3e837998c936f0e654a0162d309ad9f559eec316
zd5d06e4052d75aa504d51e1e3231b4b293103f93d4ade1c7201d9375ff6b668af2e1c7f0f58fa1
z154b659f1e30899d940e615f3aedb28f949b0c3a158cce54d78e975b57325a17776d2cca8b575e
zcd8d9922024f2df35595acd661796daf1101e714618c7b9839ec81b047214015d2674942097518
zb2c919bf803a0b062c2711f75ac48aa0f61fdefbbab015897a444092b08b48bea817e6c5e893fc
zea4b595c89e854e3f6116d2779d4df1cea1bf61a5cae1307e405df4356e0f0e3c6e32d290ad28b
z4f5dc0f4212f7a2a8e187714025f0669cb5dfcb973b9bbbae9e05e3ed1f265147abf743f3f024c
zbe5f5ddd2e8193472ab37b5a063ace0e426b2064de174283498d6c6e092a88b08e9c3623737338
za3ed2e690a637a6e1b2e664a8d84f2252ede52943c35f22754e8be519bbb1920e94474968cd933
za59dba8aa31d2a0abd96b81023b71919498338a1900d3cadb0ead915c96e4f1dd4982153035683
ze5b8a5293ed1cbb1801828ecf9549d84d81437bb2342ebb8e72db195be0326ee13232ba8044ff7
z3674d3b2bf85c081ca2c94977771e5ea114de8747c9314d1333cfce020248772289f513f4252c4
z87a063221ecdc232ce6b1c9b899072155b03008cc7d3d021f55b2818675db4ea070c3485a2aea7
z7829c8a8d2a486653c598495115cdd3a18d37f6a6d3b913b204fe047f9263edf4d728d58c47457
z4d5a28822b7de233d9e3f18b8ef528ddff3fdd05b53a740e70efc80d13d8a710eee3afdd5d093f
z3bfa2c3f7d6a4c9b31b3e289596d01d90bc81b8d4564ee9165a93c4391a2e6bee38acd40443f58
zb5e80b451cce9c3d53655ff0d2f8a01c66b0399bc161ef6135320a175a9e5e52367130acea8fcb
z12a2e05f175fa94523a9b7d9eb27517ee30f5d4bd2341455587b84053736314e178346cea71d12
z06e920f5472d7831ca04b02a8cafaf5756c0e8972db3017cca908235f09138beba6750962fbd61
z188e508dff691f640c0d2f4bc414683801227e1b13e2f4e3701ae4daef45988502fbb8b76773bb
zdf6808242663d580adc3cb4b1dfacc38fcfd1226e956612e8cb2fa1738780ea185b10846feb3a2
zb78cdd0ea5aba93b9437b8c0347364dc90ac0fb8c2d1d9a02d6b8e3800f7b04a268ebe4051dde6
zf9cf7809b5c163046f47655362f2a9c615d39d352ff6404d24ded68fc78d13b8e0e473fb23e292
z106be2f161032fb1dedb0e259ceb7b3b97e0466a5aea437b1dd64afec6996ec011ede2b19a2fea
z9e720b666fba1fadd2539b1d3f111358b944b499f7b79da1f0acd7095d5960cc79af79daf98e2c
zfc04e0219e1990ba88eb99ab6d3a467711aa847bbc011532bf8bdb2af810d3e1024ba7d0ebc88e
z605a69f4c582cb1a7bd081bef3a0097452e477187b20c9b31b8b85c678e19830e950492968d036
z909f899ccd8869b8fca76b7ddba8509e191796acb8040e7c45f82b640574077170f7310dde7789
z874afa3705c3359c22a665446ab09726aa849566d94779c4f1d692907467e884ed4868697f8b9b
z2d5cd2d66c3b16f633b157655fef5a0744447c1acf74da0beae6e8dcdf7274edacdb6cf8384c38
z9ecaa1c83ea7c9b4f1b247aba5b9889eaadf383e064c5b37c7f3b474b221d3218daa1314996de6
z0788338fd38f8e41df47f80d1f041089ee616d09410b180ed5db234cfecb873265267c6115c540
z8e73136c95cd43371e43c972c262d43404160b853a1a925186549022ad1bfdcb43faf9ec1b4f70
zb3d1e433e80385451fabcc6f837692c5d6f2ad4dc3e2a1e46cca8a61c9560ac4b4324f37d708e8
z84f9356987d28d3858f2b5a6717b5889e4494c3e5e3bf1493639abf62f9b12384aba2b57482ff3
ze89879fc20bf65f331dd27ded55a5ffa6e0aa67cc90fb307f22fd2a44f97fa5fb6be7d96c5bea5
ze67faea9a38e71aba46506b93df943c3855aff8410cf71864b5b3fc66d7334d167f8ae8d67931f
z4f15e588985c4048d0af5c9f2c7e7a06e3e80a9b91e49fcb64584985d06b12a23b5c30c9c610aa
z936546bf6fb50a8da71581b00629ed69c1b205a7370c55141bc88613a7b6136e9aa139819452ad
z49df83459eb57d5310ad74f47ac209412debe01a9eb81a0ab6430084d277c6cd7ee50f6084b733
z12b00f8565ebc770189033b437e82d433d0278e1842f147e54e70953ceb5490975af7ed1d67878
zc07517970f36d5da09cc23d28d5a704634542e548a03a1bb9db8d24fed852169d5870cfc1c9e8b
zb319578ddfe678790e6e2c381cee391983bf92896f59dc0a4dfa5f002007a058bab3b943d0d8b6
z6f2c7e40abbcbceec2b3275a46ec14e6f31c299d48d0f7141ae4f2f0b5cb4acf8b2e117bcf3a9d
z94c8d564747848eed2e719850ba5fa755e75b5fae7c50d39d465f3b6df2bd4c8a847a89ad6c037
z0ab4bec6861703f8961590bff1fcca6f3f935d5c5e70b3f1fea74a6c3588a553dca2b062f99ceb
z949da81210eb5562dfbc95916deb75b9f313aedbe617cfbbc38660667eff10c2c444282a038129
z72d7033396c8cd7e7a567b16e9a149fe062bc296f884cd8f0bdf9ab977afdae6287ce41808cb31
z55285aa0f58f04baf280a4739553232b97b7e0398c392da9d3c0dc8b1908acda08c6c793a92af2
z1c15009d7a891a57e50756e781f299d1e8c6f171cb239d17542cb6c91188921408f56fe44ec439
z1cbe74684ea6c805cbeb6a1ec280122bbb4e4c45f166b8115477b82277bf5de665d702d60494aa
z26eacb23b8023a8207dc055f7b42d7f48f97bab75fd5622c35b2125c76c30afb8881a609a6e3c6
z9a82c3c95195bc573b4cf73c703b33e20188a9b616199ea17db1c0359aac5d8cde32322037ddba
z8dafef909ef9ac7bd541bbf6d0b9f69b2d7b939ca8722548dec25807dd6adac9ed161133e5a997
z3a7cfa4890a467c2b1c45287bf607e1d4bcb39f520931055f55f190bd7cd24ceb46b0c1630cfe3
z692f036fee42824a6b6aedc4038fbe6a78354ad0530b445a40a1ce5881d908aecb38278307f3da
zdb546c9cd403acd674e7e4c616b05e0c75235fb4a5d0d1c478165494c2649358670f49ff778580
z84ace8675218c048c0f68a7e7728785d50673ebfa1db46f668f07ffbb33cc289c70c95cb39c762
zf36e06154ae3b51722203164f63fd70e20ad4b510da94c446a11aa9ea060be6824ea537eed2ed6
z42fb2abb925f506aa1ba6b87ff7c4b2bdb094f55e42492fd892e71d008903b8c6c275a7d4b7990
z551ec55d1bf1d03b42beb455000e230074ac1dcb0887d3ec6093e40442a4e308f4b143268b5fb4
zb63bf0f37c54942e2eb0305b242c4e8680fd49a153c909e7e87d71d4364b79e77ac8a03663c970
z31682f6cea414b3b40e864f3935a895a153c15f86d27dc487873d1d8c0bc91ec2eef0bbd28e59f
zb9457cb165c900d4bff6ff5eca2bdd26107c26a60e609da5420908d5c44c9c20f8b5c4a4204209
zb634553402090ed30ec5a168477f92f00a3d233de479b85d938f928b3534ca61243ff19dce7c9a
z466b2e8cac8b1553701a64914d1ca7f4f991bbe3b0d1864cb2c4f929fd5d8e6fccd3758f68ba34
ze0a4ba12706e6d965339e6a979c34f28fb880a03da04da873c715b48b21390e72bba70492cbed5
z359618adf34cd3a8f21a40ca52a8640c6f67d2688d04da1f492727f8f0513a6f5b3880e676e725
z928059c33780ad1bb013255c7e1cfe6d6f2e48d091722e9e08f6e14a928b1560658d29ff2aed9e
z69692124f1cb1fe053cbd321355070cf8ef985b95370b05563242069d738e48f9ff84f8eec74be
zf12945f7668788ef6c7bf53f4162303d5ae1744ba6bd44b192db31aa374cb84155cd15411f116b
z4b95f78f5e6a6ba1a1dd65cf0f33f9fc37eca1ebb44b15118bd506c88a159803dcc60979aa91eb
zb21ec3a4d30a154a5c8362bfef1f9dbfe7a8b2947a432303ca94482ba635f8eabc4b9000e9bb21
z3e4123162c3d4b0e5b1f130eb4ef7fdcb57f7b23bc235bdd9c0b8b26779747c0235c0de0655fa2
z300b8e4ce73c13df244d82e81e874f29b056b8ff78117e6c523ddd11e428d106c16ba4835150ec
z0f4fb988b776400f9ef5843d836636e4cf4e40cf8112b2011eb2849b2b6bb2fe3972eee5af8df5
zcfa544988af074b5e76afff1873df8692a582bb6870aab8ed1722a638def649df5b4c78caae2b6
zcda91fc8e8b6234d31861bb7b461f7fa2ebf4033e082aeed4528a0127d093b2dd9ba0dc2644479
z5fc0a70b87e0a09ef28f172f0af210c6c4f6bd57ad88441a622c9fe3ae3fb7ebcec475e41268c4
z2c6effb211cdf918cbe28a62c780330f657534fcd79fca4d22403dd6d5b5bec03ab98b9e578402
z8a2f2e1edb1657dc0843d6cc8939175e0d907bb8c76d4bf0ad5e7d19d9773835e92661573e70a2
z3498c597df74f486ad5473b9884a740a6b2463b8c9d699ce4ee57e18fe56949e0ea74c047c67c2
z970dd0d69f198b1bc45526c289330de2dc284857c3a26bb21ed316c3a89d446a90db8750f92fd0
z19f1feee4ed75ceb0a50a03de5e1e65c782faf3f9b2c7155bf1da4245477716ffc4a6d26914d93
z1971928999750adfb14a9db51537c129e071b13a0f433368047de623fec82aedeefcdd99be04c0
z668f862404d82ff841b60af65b5db0ec5c87ac7eebb117f421496fa7a77646d4d87792fbbc39f8
z7a465ae5d4ddfb9bab937718c73c500d23e74702b87385d4a66c2082f424fa1f437e3a9319ec79
zf393e9aebefcbeaaa7c541118c4609b4fc51069ed877004b8970465021337cd08715a42dcb66b9
z63dca5eb14763deb225bc4d8c6ae7807eaddf1157ef1b89e9e0ce78ef36fe3583d248c658b9297
ze340b45725f56d49d54c23cf1d549cbe5689bf8e6ad5569bfc0a8797aecf8391931a8885d3710a
z55b50e6db7ab4401c806fe8aa437f47c694146ec6ed7e58b50cd17c8d2541464fba82bae3dc19b
z7fef393a66e57fc55c7ee046d5a4f56d6f42a57d2d9f956471441889c689ac182bb0a03670792c
zd0a3a94a12434a3ed3ec0784c7a6b4552142f48f173a3b82248fa2a89f6255d0925ff8c8339be4
z000061c244e7d98309461cea32fd1490db22bb8d8723593d9a45fa655763a90b30893c9acb322f
zb6364f4f0b3d5cd7a083df69eca7e7e7c09d94ede52987c85844df26da7cb1870cd23b7146f25f
z94a24a9e91b191c74c60e6999e40a381e9beae82574d132162949db486e5f4d4fdcaa1ffa2a3d5
zafa4aaf0620716f0b50f69c56f0b0307194082700e683c15b5388238677a664bada3382d014908
z7eb50187da692c8ecea23807961f64e5191379f30c509cafd386df7d8e9b0a8637035774b45d17
z0a561d41c0d1d9d3d7b1f2281e516f7760aa64b92c45d364faba27caec1a78a7319b1c5f4b5925
zc5c6d9ee99a6d5333c5641e765c9a5f671105beddb1d4fdd170e6c7256bfe79f33afa275fc6f3f
za8664a878e09ea7d55f6322180c56e0bdaec14f3de4dd5c5019292350c5f968ef895c37b6ada40
z99bbcdb6f865dea7feedbf73ee06ae319f60218e68eb0bcd89e40f9ab4c07eb48eb34f7943225f
z6ad32210fb8e06654cda3f8a38a3637ede0bd70401ba988c468a1b2b12cee129c52168933f97dc
z17f3e4c81896ec348db039907a621a94e4fc7c21a56391d7cd4ce64e37a0a083c1d3876dd45240
z4bee473e10f92908b930c638acd0fcec0e065acf28f400ee7b338f5f6c969fcb50c424614be3e3
z292aa713c321faa10ac2f4fe6a222fd566b0a8021e6707e44f3157d5b963708e89b4a8cc6a92c1
z0545d66a01eb956ab640d5c3a243b0aa4d03e446be6edce9b378f13b56ee4f6486fab122aa9802
zb099c6dd9b1fae08562ada98dca566f05a2dbe7f939ffc324b2d3dc65a06d3d2d53593c6deab65
z711f1ff7fa5ae19f6098b614287db5a853c38386b405877e5df49deba2da17999a72903a74ddb6
zf1f093fa93bc4932c8ef0042d5f3cd5605227d8d50777ab45241f948f9cb420943bcb94178949e
zd4f7856c672c3e1d6701ab45def50538a823cc52b583f06832dfa5f93b06bd5fe8986219f202ea
z2a7e3c04ee65f21407fce5756d0c4b6caa7b03795c11b0190841bbd372122c01e39a8765ef68ab
z39e76473f4a4daef0c808367f395f4877661629752c12088b46e39dccee802c7c27ced9d87056c
zb684a3d21bf5b40d3a8e57c39521b8ffd5e1c8f8f3a84e722e74850740746ed0fac71a361b17e7
z119774ca42e2ad325dcadcabc67cc2c6f86344fb4c6b1e32225874f26b9a904fc20d9ff6c1e11a
ze8673bed54ebc8b48041a7e0d9f7e9bce4919bbfa6882303c6fb8a5e03bf1e982d88df0d26b859
zf47f7fb4378e57ad2b75eef8f884f1a8247a1bdad2ff8c8e5688207e3844e1399fe42f7119de32
zba1a8b3ed874fbdaa4a0f93b6c97873b2c991deca105f5c15a8c9f3578f35e599ffa88f9dacf35
z7d6c7ab99b8af73409aea8252ecf30ffc50305ef6332ce018057c3125aaa474f0a7dde9cd0af1a
ze533936528657a1916ef9c7eb654617b4d0fab5b7c269f05780a51311cc1ed2978afcc38980bdd
z8b130e6589da09c0a791b8613856aa40b996585a5903fbea7d53a1685004b0b241b3dbb63af8a0
z5751cbb425277f2c94ace7493006abb0bb14ad7af15335fa7581c7114b8945c743e4db409cbdb7
z09239f9bee25dbe7b1af8b108168bfbf42fa7e4977294a621b95b4f154f54e4b8b7cd0102a7cf8
z0168596f9e43ed07d637f38a7b3473121078fe7481a354128c9229bc5c3cee24021f25f1dcfc56
z88218404aad6d7902a4c9efd3fb4341eb3a588a7615bbc4eaf5e7ebd84f7364067371f9f1a0040
z08f536b49272218539cbd28c394e3b6310d8f947acb6ced5345f9a511b1745d9c012b5f17ea2ec
z917a09df6697359e6b38aff569d141431eb88ce3c4203604a5767ff1f8c8a2893558d816afacee
zc0254592c2e4468151691742f5bb64a639435c67993a7a2c0ebb976ccfed87aae5ba0590605887
z8a08a30f8bc059da8cd706481b259926b70f968579e67fae3378912ce112814942a497e09613a2
z0928abdf20ac8c6430a57dff90c85b16e2158c6b28233af7bb8ef4503bebef1c70f419fb27ae01
z3fbee1bc7f98390f3c49abb099461163ac376ca3da26d325613b5a0a73d78c399db8d72a25c0f2
zc9812d049377923499de346c2d1ee34c8fd2e8c41c7fd4fc70528f7dc64896d134c707b7be987a
z744c4243e45b259a9b15cb36df2e064ca02b08b349c14353099f7947b7d649fca09ef2f99bcedb
ze7ee95b8974f6a5ba35eb5f40a7fa62c8f94bd45750bcb456d706421fd8982fbfbe91061999c82
za81143cea05b8ef4a9eca1e35fa15cb039d174ebbe8ca8793e5bea3924326e9e2a9d1e09ecf135
z9dce8c1de4f119471d92cd735b0c9620e2de38e8682b76e0974dc818ad01047e0904c6a3365bb5
z8c6c441b17db6b894de2218f812e6f4c5c7966f39e061af03ca3c7606b9860a1338d43a877811a
z18281b1c17ae4df1ffddd0c63da8bedab48838fb8e70fc4a0749cc420b66a68baf414a6eb949df
z7681402de2344f699b95a4e6f5084e26eb187fe67a6c837ebca09d421a41d20f3a77d2b7615740
z06bcd003f5b53940bb85cec964d0e541741cb5e982ff49ac7f34956eb53c3745e2b526859fd8e2
z029a0abe7afe4b80888284eee454ad9772a472e44d9d0dc10f558f442384b2edd4489c7a02e7e9
z7dc8ec73289d2a5bb022e8d6e96054636937d6d04ce9dec21c238cb52a219bb94432363b13ad8e
zcee4a209013d81dec59781f3e0615be5ec10ad40a77507afd09e421af9003cb6c192a937779f4d
zabcb047ef6e0219c275459c62d1f60840c73d350e825876233c30b4c9e9d59d5e98d95ed5ea6d3
zb126e4195cfd50ccdff0a32d76898a026b35e6ebe7f9b5cd3ddab2d63e6bd1ae0897f2776643f1
z161aad48c4b95af52a931dc605e9fcbba45ecc529cefc85361babbae6fa1db393ecf770ad77bdd
z2d687b03a63bcba09ac468e8ee084c6890201bbbde53f79bedb740ea98f661e0c908145ec9ba3a
z271c338f25bd7f8cf004d63392b23e8b1d4ba150aae0dfd2050fcbf24218b0fe40e16cd84b1d3f
z5a13cca06965fdcf472de95bd820bd6699dfe3cb87dedd0f6693c9f9d78a4ec7b47cf44795a6a9
z0e8278226b2c56ee19a70f5d6645c8f0d04688bc7d33d5419c3e0a521c2a661fc9649f9a771ffa
zd9988a36918d24223aff805e98977739e266132dea05d37d1e0cefa83b283c3835b69c508029b0
zf1b6de907ab1befb0b34bf9f3fbe201b8de4c2aea285e2a00422f874d19a2481eb6b9e89a91f90
za3840ace9a4a239124203edd14ee112ce192631a3abc0489c3169b724c79dfb45b57d266849745
z5a9134e0b982f752f60ea2bd37121f19796efe53301c1ff8bc3aab1c4942e310873d86f4bf72d9
z5997c9d50d6741b2eef48664fb8d77ed6e074ab84f4aa1eb63d8c6096da11de449ddd974ae8c5d
ze181dbe96bd2560d5fee4825a78468689a9da992755d3e0907e922a172da4d5892f07f3cc706bc
z50d6ff2a12f5136c0a7f5bc2660049e685651eecc99b371a1295496124421995d72d157581e03a
z41623eb3c3c63a2e53cf9250a969f78a2fb55f3007b4685e3833835cdfdfbc7e5d84ff01d31401
z30029804e21c1f2c4d1663a01fcac9bf139ca22eaf87a3542113358fd91ae4e47fc8e6a7396273
z7033dd95699d5afd35006bc5923a7d28ab564ac9c8b8200b90c3b39bb93f28852e3546970aa29e
z20e24f6e7908f8f7fcea54c7bbeff6f0c2da418856e747186528a87114790f22b29964cd5a018f
zdd63fae9e54f715c6fc0018a719ffc510455903be95ec1d30751f2fbbb3e8e3339c78527132ba1
zf96beb0138447d5bd73f7db5e48ffa25a3993192bb0ea1ddffdbcca571d144f79c22b27771ccc8
z870f103cd4cfb44013bc4a59068467e5ef1704068360b08de9f4a059998f8c30a71a8e535f6bfb
z9ddcf14c48cc36e355bdd2d753c9225cd14e1df2dcda718f45147f9e4217ef3f5ac2bc9c8265dc
z7fa338324378ef96884d84d9535137af6e0a09e14b5b618b707468d300319fde13e5df3e53e093
z39b84fb6c885b4d55ab43050c6d0e763a3f7101ecd0cd4680af6c4a5a90bca9906692ec6e06ace
z458e9f48be3706fa7ca299daa7870fd59e839cfc91618c4a296d0ddbf851b94bcfb86fe4735858
z19acf74d2bb328340d8239e4e16aaee66123cf427eb06e6d528485ceadd956a2644498df0065c5
z886b047cd734e0ae0413109941065bedf252e0f63d35a9727e96e321bc2f273263f44918b2e8d0
z14942682863f677f7ecf1aa2e5f03fb04b93e7b2dfca6845f7a01a94239b104088a9fa07b08c1a
zb253138925b0cee81a8a0a097a3fa9b9d99474a0f993344044cdde6cc55b40b681ec7af16617b6
zbdf94882b75e6f434a39cd871c6beef12adc9faad23fb93f66aec604a02161d24f8ece395ea372
z4bd7223adcfebc8ad6f200ced3a395735f6b79f44e05d27e88d857afcadea5adcb728b61e577be
z981d57485333531b7bb184bdbb7da76407bcdc125d0aeef02c387457f522d5e591c5e426e5246d
z70af2cef03173870f6201cd90b31295532453223cabac9f550cb4c20748dd9bc905e4a07480d86
z3047594b98e251a4f8587b4a1a77ae38732d9158c16dd4798eaa8cb0c9014b9049e7c1cd0124f5
zf5dbdc2c22cc311c146fee48746e4ad669ce6365f6c9e7525ee3bc7e5bd23049023cf402512b06
z2fd298f45f679972be673dc1f037592ab7565d0f01ac75f4b52de26d1081182bfe88441a9bf114
z74122985a6d4e75317c031fa83b006098ecebd671b648278dc6122e36ac0fe76ebf36b4543931d
ze5a216e8527aefce5ada08ec8079a7c3906ab8303cd7df36dbb4f3847abf8df564ac64a5a311be
z851b3c75a427c7e238504cc15c1f991c731613dd024e0bdbd0abee59ce28fbd6246cfed3427ef7
zebb638150f2708c40ca4102a523f433053994fbe54ad7de6e46e62559eb1407a517a68ec4ec88c
z2ffb662dd9c3af57558a0e7a3aaa5ca754c3eec95e4c81e349d0c8c74b2adff303c8dcc57b7106
zd3fd33864e371bea5aeae6e54f01199ec77104e43e96518161c6623430d4cb64f2ced1b26f83c8
zb255f2e8485346d88d02f648eeb4e9c420a1ef83d949710e89f9c6a80e9a48e50f884b129b3103
z3d7aa58475ff69428b3c12224304724b467e9d0807c6445f1c4591f9d17371edfb42b579266efa
z8dda059fd8a55a398d9cbebe06d3cfc6946b223795c40ef153ec10d8ec3c1d69fbd725d32fbbeb
zb827ca6dd457b8e88ce6f6146318e01734655b4e8bd2b75bcffe6435c1f42c88b52c07e778c127
z31bc35c79fce966d311e2440baf0863a4c507d94dd0a0d79cc7d76df77a6fddf8b04d8f4d032bc
zaa52863183647b1122e88419808007e5280477d377cb7352a071a13a26c6708baae287acba15ae
z7244c830420bac31847130d25329c6fdcc3c889dbf99aff258d9ed58edbf6ec15e9dc8bb33cfa1
z2855526efa484f82372dd7d8d2ce3629b7072da64953535f0240991380bbc2c6bc9d235e0e1ab3
z3d18c9aeb2daf559ecc76f44dc6e5c16abfaee1569c6ecd302d6ee42093c5b82645a8d45cfce94
zdccf5e2d100bb774c18a951286bae7849df18fd56a79464fb98d4d743e7365b2a7975428240f0a
zbede68465de1de70b1098327cb93913385b589187833782984c87037185331052f979fae8e9124
z2c8185d8c551b50aea130578d3acb15edd0bc9999ae50e303768c84b5e5411fdf722e422cb5050
z8abee601a8c709d34b7a367865693d19a05c9dfd37861c995ac8df3a067128eb4a18ceb97fe82d
zf8ba07aab0881a7a066af2f88b758fadad0ce76b69cac47b0d6b69d6042c30b3f7a2704b9f2294
z6cc0a7c3e2043f0cca7aecac0f064634883d95abed3a019e9bd412780e9fb97db6a4896aa2779e
zb7ee3e91d3ed03c76fa380d0c5f275dfaa410ec8b6a14f7e4bc7fde9b6fc01967bb726a9037c4e
zdaebcd5c87f21cfdcc0d7c757189375f807c25bd937f2411da83ea3e8cf2a2795fb5b9927acd57
za882c5e886702cdaed9bd56121de09ebb2ca801930c685f1f1014ce30f671d1136571cb34c27a2
z34df93e54230ce1835e3d8ec825e467bab5dd465aa95e656d89532e5ab61fe40f4f5186ba737af
z9803fc7a821561b4b0e80a49b343c01dec7d6f8b0456f7d5d02cb62eb501d157a3f8dfd77ad5ec
z973d2a009aeeee4d225f54989d6c4d6bb61beeaeb76c0bb9ff5a841e826a92914ba1bfb4a12036
z63c30502f051cc4760c328e515c744595e01f568424ae5ddf5fabf3b089748b41f9bffb658fd1f
za4dc9290cc9d0be67d28c3c287b1e27d64bfb2848687e1ce655d6845aa2960971c9fc4d9655027
zc4e4f60589598c511554eea27cf6887ee669cb531f536f20c3c9dba420dab9f91d484408659b9d
zd995ba775768dd2fae23eb95bcccae777ed8c8c75f15a370a37e96fcdbf854ce9c1b3817affd20
z64b4bb08cbc4cacbd99a585a8c1ee742f1b9237ba3e92c93c0baf0a02f90d0dc974ae17f862c03
zecf7be68df677979b8d88ce865c86981c6c268028f2333756c7c2a077b3035f6463bf1f1a4dd22
z137fcfcf546373cce9e0efca2227755a584367abcda24e94b98e953b8ab61abed50e1c1c5b2b8b
z3cd0796598490d9dde7ac3e38032db1d84417515da935be07f7941ab53a0c6f9be130c18806d82
z2ddfb9a83b54f2852a948fe9680dfec6e5340e34adb1f6b00b3abf73bf8a96d35830d708da697e
zffdbae47b58084f8cabe9adfca3826c0a9e315a7be699ae0c4425df4d319c0d17853597ed0789f
z02d4fecfb2768fda5266d575eeff312526be96d19e27af313aac9db7e8c18af7bc6441fad33f86
z6cdc22cce374fcc1bc3f0b8ab7ff0561f207e6a61bdbc203c8ffafa6897ac54760a286484fc861
z11f736c075503ef661e588826e3779d6ce1452bb45d9c181d98b1089f92bd2b8675a848064691f
zdbc1fd2ba9186152a4398d02dbaba432f27a0b7c9c2fd96c8b1c2b320f1e5762f00d1796129c65
z44aa2e5c738821d46401a408604dc5d0aeecf8addb50951cfd5dd913bfbfd42593c4147b54ad7e
z378adff189cfb592a0eaff0855d5cfc9a159b90aa7d3065fbf039fad8f49261f1f1707ac50b04b
z25abacf5e06f7004ed1f6a71a474de08eba7503f2ff3f6b2cc73428bf946df8cc62bdddc51d805
zdb43c1ac80ea9ae765bf8b0a8a373a530f1a2b593527d6709183f485610fde88bb8f74e4bfde1b
za3b3617958679479e622a461a1b1da4e9f6d9e7ef6eab6a7fd98a3b0b0145672f753501e436b26
z1f0d699250ee4e05de7faf1f9eae098ba0f8d25f2a69e05322be00f335f3003d673fd565efbaf8
z2cd77c9853b572e38cb6e79ff71ab022e14513e2a63ce4fc3e5696288af549db25886ccac8a1c3
ze28be2e0dc460f7faecab3b6fedc8605c1a1234b5428f9948ce374d32e72454819150ea649831f
z418e1f461c41c926574378fbdcbb63a9e4144d0c0ae735de38232393b6b7ffb830a3b4abb460b6
z03adeb5b4e1099f99bd79cfbf0d26a32688877e31ad58ba11a1a439269758cdfbcbac6f73b5c07
z167f4e7f6c03ebf3df28131d98d65b7254886608445c08045374e77dac22686cd8e8764ea4a096
z96c44ea4d5a2cbdd26f032ac6709133a3d737e0055d4a654588b7d257d5bb77f75033215e08d73
z7cd233ad82e6d04d9bbfaabacc55886d962dbcf19b5a5b04b84210437c21e4b403e419a89a4337
z1e48ef89c92dcfa92c90eeb4b5bb6f61d2a1f72dc2f7d9e6c7aa14235bd5807733216fd7e8bff3
ze4b8b3a4373b260eb965e6ccd16db7fcf608e4e55759817fe15b86557b5f69eb29e97d5210e6c0
z76156aa3cbf71a8f6ebb987fda0715bf877cb034680d74eb8aa46b248cafe15278f8bb1cb3f815
zde075212f2827b8678154c11fe6614dd09f0d421d8c24af41109fca22c041d9ba4b76175ea197b
z68d466d5a398e5cfded4fc694a9a1371ba0ca93654dabe9384be2193abceaa421fefbe7bc33883
z139675996846333cf26a7c1f4706d22458e1c4feda774a10d4e04b8494f85285a87904b727318a
za397f574c23d6160cb6f64887ac4eb43d38da4babb41aec1e55e6e0c7bd040ed2f693d93209200
zce9d7b6c383c958d4f4ac14bc9c6c957090fe3ce43a274647f35df4f43d16e02325c685b63fb1d
z5eb9d72ef69a28a6148df979a212d63809da019043c16455532df127a783dcc13ed241d76b1cb3
z0c780a71db8c1d8b864d57ef4a4ff81dc83a578d2a5c85d10b49bdda8317897e4f433c27c7afc4
zb44883f386e13d20b71af67017836c14fe1efa80fca6d5767ebea4787822878c89a60e855a8859
zb944ae42087642d2ab6767f0261ce129ac70955acac6f8e6870f5bee312e7e1ddd0baf0615a321
z53d4399d622edaf61045c029418a532a812c834b053de5d258e29cbcb174b82c4619719e6166bc
z0c0d142297bd53c7ba423e8d2524394e649d7eb23233a60e5c15b0b7f5e727d196e6c56834909c
z420efcab2b02e95973fe2e68d80757bf444393e9516ec482e4951d2418610e117e08baecbb6734
z52e6af9f7205d83785ba73834fcf33ee54e748d99b1d758a01d7c4dd632dff81602e4038b19667
zb858eb8589f64c09a8ada03f6bb0b94d58436f9dc70765471a08db6c3be83cdbd3326ec2e32688
z4d2d9a135a043c1494250bfe24c0f582c0f5195212bd896a0396b3b00ff73d365f0ad1768e92c0
z5db30d12bccc1c22190ed3ec53e389734260bb4620fdf0e8ddb872d1de3ffe58aa9ab2e3e17c4a
z0cf04d20afdda7e1c44296eb73be1795de4acd36770133fc4f5ff61a1409b31bb112d6eb83acc6
z30bcf97d3f653964114081837ac0e95156366a933dbffdefe222bc6f109ea4cf8e086bf6e6ac4d
z7f6030886e96d188639c9287de4e17da0601b800525d2652005694efd39094e15e9765522bedef
zd47e94cbf921dc343c309f621e1968406e0585dc7f8c8e8fb673ff67c1b597baf391a38a6672af
z048b7a05083113f22886b2f2fa3358ab609e405bcb18fe9aa095b48aab772225371ecad7e357a9
zd1166e8b44936c5d9899a465b0298c6e583ef691cd389f8fd8ef6e12e15c924884abddc29d762b
zf310213c1080c9cc62028e44ef319b451d02a2036c3d67cd7ef633f365809b223a7ce8e1d4d2d7
z495bea3a8b9d11991bfd2e27d754ec466119b338d92a427372b4f45689c870b813e9273d8d0b6a
zcc708c123268f8755564ab3c342288c68cd659f1b90a4827f6a46319881649ec90e5a2de6d5540
z24ded822a2b5ffe9f78d8543b34f6138a900015d930566ac640aae7634f7a061934fbb5d392acb
z1ae170fc50b1a9fb2eb0b8cf9473d6b9cb6e23e7788a7e68def9bcdfcf139aaa63fc84bc09db56
z724fc6db2ebdf272df8f6b5302076f7570158de765bc58229734b48cc9339f16f9598f8458000e
zb6b1b6d2ee2ebe2301426fa51df60ff2ad7867c4ece1d8efc7a63d3fda8b59c9aafb5724706f61
z9b6d35d865c6b7ec8b36e0310c9e0e39467d53937e3b84d5267290d6426b6d68cb2ae61906eb77
zeac65155ef38a3ec771f3519ebd0165421a82e26d6c9a0f295d3d08e797bde78a0ad18e9b44f6b
z32857df7e8f75b796d23d96eb9e211c16877cffd8daa281fa1bb2c033bc06502e74852dd4fde85
zb2978c87ac6b51e70107749957026dd803f93070c155fab070946f8dcc83aa52c707a7875b86ac
z2f035201c313443efd501ca7ee535250befcbcceeedfea81bae27716cfe1e495699328be0305c2
z63a5832ec6667de3b274dddc28bc08d195071fd41dcd9dd43fb165def95db5a140f2f48831a285
zb24a121b700d81a58f98588104ddf9a83b9306cb92facadce01399c96fc37c1eae56a6c39d2333
z42a05d63eef87c3c95b486e0a99c42e85f7b44c5f06d6059866a0caf7ac8a079a51fae720f2680
zfa11d53b89d546f550c51312cadd7f46966a3f32f12769ca752dffd4c3026068f0052b6e836476
z59e221e2e6a948c35a7f63d833de2cd48106c10bf53f4a0ee5d92971c8f9f5469104ccb235d32d
z352a5919b468ea100d5a2e05fe3b6d481ce6acce9cbea069c6b8f2328eec780b766a8c1bf8b87f
z6bfa5f2526d2979b641d632ae7c089703fe6a061a2495590b64620c25e49e4060707b444219dd9
z842241e12fc0f0a887f3556da7eb81625782bd2411575ed81dfb8755b96553567b817495362045
zd66a72614b9c87eb86e3eb6b62d07149b8d198eb06e489aaae2f7e932bbfc0274ec6e8f2341700
z9edaf6142d9d549ba53ed172653494506765de207a0b7d742102229ed3875625df02b6d499d53b
z885e29bfefc60a1b97ed8c30ff684487645ec463183074f204e901962b0ae04a5a476e5bae77ac
z653d501330d7632f1fe38fcd9eb6ca014b5750bfeb8e25be795a2dffbefa8f7a72d0c319db5bc5
z012f94df4ca0c8bc69e189c4995add9b8befab3abb6a183f664490355d219b35f6ff71015112ca
z0b407a4a147205f289975d90e09694e13f8910718a88512bb115cb713e2ab7c8069408d4300402
z3a368ca107d2d3b81bb74df1bb4263c0026605418f83205c018dffbd68f43f7af9c695a02ef825
zbc42e2fa47dd82218cbca99763986e8e911df72462013acc44bf68990dfc1f28720555ecefeeca
z546d282aee2fd52fa27fb54f3564a20027b19e541aed6cc927247b458d3ad714bc977859b4a8dc
z9e2dc4f20365a2c981f326478dd61553b22d918bf82e6edcb20cd32d2b5156202ba3cd8bf03a60
z741e9db2abcf7aaf61a87286268a3b3f56218be10662351d637e43f24baff1cdd9a7e7a43260f1
za68ad3985148cc96531e24dec55091fec313abff8e4bdb6112baad7bfb74e3ee6ec6c6956dc3f2
zae2d19663d324650d0a39a432f0f1fc0d8268901c23348f882d2cdc84ea129b8cfceaffe7d98b8
z13e7a76d01b6489889932127d1fed197459fae2265e65e31425424e53196e584c087d8b3aa85a3
z3982f966b2437fe253fd5d109fd6d38a3801d5e989435be77e40527af81d65d5af4ce25c0d0631
za480db06fb4d2870aa42a481b39f3feccb62039607517a27ef7d97409dc7dac907bdae8d8d71c4
z6556bbc483089b17902b1ed76f2dffdb344bdc304c0766ec402b67ece92ceee0f261f850e60fea
z0591ce80c6d948e9d74d6a3f9100f87ed07a979d988c3d84537d5387f7e45bb4a12f6006e492c9
z557cfae524fe01a27d2ac383c4226a667a2bb27c3a1b47280c30838717ba22468a5522800d2514
z7ff0056a1e0bc9f48d235a55857beee97d18b8387a8d91d9ee916e5520e47633b5089b0312f597
z0177012894170e09df0f479170d0c3ee481ec873ceba0d58fab00df13f3b683d26a3fd3ea331d9
zd4683c33556aaaec33194a5e3a087e494cc06c17c92b3314e1b44c164b01bccdf8407423c16f61
zee136622584f8862e1bd05076178ab59db9ebc0ed7e9497f76d6bf79c5f565aeff68fab667524d
z0af2bff8d37ef07dcbc88c37bb6413ec673df4617f22431dd14d94a668503f63b1cd4039bf890f
z1e97c1c8a981ea8cdd6783c926fc325118a6d857931dd77d1a7897736cf67919c37f9323d41a00
z9a5779b26efe9044437036665d9444af5c7bb7c473f46e19f7db15d3c5aa90cb9f9bead3cb6864
z7852ec08c9d6bce4d284e534111f9c5ce7a06c160bf6e2707a5a5637056f0dea2909c54e74a751
z8b97690f47074fec3ad29e99263a16ee570b6efca44243e4cb1b8d72d0e97c618b628a03d88794
z5129182eb8fb0b97a9fa8cd51eb9c69a91ce3c62eef85ffb05ab987f2f5c1812789333d34e61c3
z1b1f9b4e88a459052928738b9870df2183d411bd40ad0bb70cbb9efe11c7fd71860f6d48d7ebc0
z600170f60798a888e95fedbb29d4cc032d92807a08d1424ee57de2cf28d81b4fed817fbb4956a5
ze0e6add24579bce64f1d4dafd88de95ac2fdff78dcf8e69eb0c570633f0c65dd6ee406f3f1553d
z5ea3a7e31a0bcc951cbbef62fc397865f1200f1e7a0ff4e927c68491977fc46cac27deadf91807
zd08be61ca7228f2d4443f562b9c5f1d11a62311ae30f33902d63f3eb498d13f09c1d0a2c0f0b5b
z6ce8b82dba7908c12005f1bd1b46865e9bec2f09f90393271fabbaa6ea5cdad68a6e9aeb92c771
z6f28a0bdde3ac910d6bf2c1bed5b3549cf5d3b25ce0d72ff98d41080c790cdd716580a743184b0
zcc503d9e22db62d7dc23e0d22c1d5d10b9ec48aefd235f544330a63ecb77e0bf09b6584643069a
zd699d42730260d8d640667125f0cd2d668b985f14b4aadc6b2ed091d7f08adbf116ae663384fe4
z67d6fba7e3040ad63fd7cf469a16595c26380b8efe168c02931dafcdf22ecd393d7dd1839aa5de
ze96c3566796ad0125fd51e0c7822bce65bc87001aa41ca95a11e3389973230c775113773e603d7
z6d2f51725b79828b27695805261c95120753b27f876dfcda21fae8876c0112fd16f7a9f276a984
zc75fdb9e092e2445ad753988d0fcf0bd2cb176aacb1c28c68e2d855658c1c59a894890eb230296
z714afcb4abb1c2abcd5b15a3988e45d775d6fb9f2f23f291f9a721b707f0dd6bbfe80a7db41f80
z2851003b36562c4f1b554578f7ac5c8d48a2d0492117724935d4dc553e53aa64ede2b7ade9195d
z263c44202220a227195e304f7978dee5138f169a6d3ddd76e8e07ae83a7a22a8e7e8a1c371bc6f
ze7d90f36e398bbf5d208d71cf0a8137fffb71a7b2a49603fea982d17d4a2b6abff27e15dd89e81
z22dee254ca080c6a51e5199689144f4f014d2362302e1384e7ad486563b5a25eeb033817e55c82
z73df9df2d02cd1faaa79380f94058449466c1358dbb4a951c922494950090d8dc2a7ef0e21390f
z549e05e61d8ab861701688c2695cf91c4b107287627de6aa6e27de39c1e63eea9aee1f250e48ee
zc074dbf30182e22b87f75d78756fd8360f863cc345ee8b6588ae05e1a10c4c6097d0f9f32accce
zf5cb298e1a9d1c53af3212d1f35d82ea307f7e6c20afffa05cdccbdab409684a8fb01f406e3029
zc65616b1a44458531b8358d084db2fad06a182a66689b9b6827f31f2ac06176800ef6110f4fcd0
z1590cec2cadfeab603e5a5f903423958fd5ce9fcc1289faad47a136d6de9d989b3841661b289fb
z7a5dd5a6f6b61797b1f3c52e33253ccc2101bb75f3ebab871e01b763f40740e81e5ed23d61c98d
z76101a064602f100ab4097bdcb17fe68f1ec2a6e117eb8901cdab9de587c97656d14a4dfb7949d
zd03b0d4171fdff891fb9e19fa586bdb0bafb794f2c3e2017373bca6c44596fc17e5500cecabca9
z3f35cd5474f3e78283617fde7f66d067aca0ee439e9c83373e9e6fa1c0846d990be1a6c94f5642
z516a718dd838e27708624ceaadd56c7870e629f703649716dcda33a9ef7bd5aadbf756a22fe03f
zd9c4989c1b992f4ddcbea53bcdeffdd6d8cba0797d19e65f3b7edca59b978bac0d4459f7c59b88
z3c861d9e7bff7dd9537305b562be9235a11c21b626f280fb07d601afafaedaeddd6cfbeb2efd73
zf2b959807bb778870c27d30bcf037e75598a1892bff0d6aa0be28fa099baa1f1a1b71c7c239fa9
zdb14973811401dbb1878ea99efff4f5223969c9144e5698a5a80d4cfe4164b869b202d488bce0f
z67bd6bdbe28bd28c423e2eaf48d53bc44b459714915c136425c3012a11c32dc40c9a2d5c4b32e3
z0d89ff6bad77e612dd9b2054f5f838cc5940b93171770c8c6e1dc070366d10d280ce8ba9c58d2a
z34b5ad411af35ed7417f9db5501142a0e939d61e571ae945784dcfa954139a0d16ae88f1c6e4ea
z9a39deb6bc215d72b6e6f13ccf33a3b8117b4652fa05e249213386af86f89f9fb7f73367f1234f
zd9b5d196e53b969141660af28a754811c53ff35b204d8e581bffd998052a27f5eeaa27bd10ec71
z29256394297b5033c53fcfabf2dc2359b4861d1289c1139c78dae37e102b5aea93e0b6e0104e89
z8fb89d8adaf8cb001416d5ee498c24e93981d93a991d0d0dfc735b5be7d9af694acf7c52a4cb94
z914e31ef642bbed48188401190de9587c4f169d6d2e45de189f472fa1c255e00d4609361e94940
zef91dc373463ce80d41fb488f3c80108065e5520798f4904332321a19779a78a01929ebc88dc8e
z6d994e4176a46cef13146e2379ea4bfb8659c9a0133783752034a39bb5a07907a5068f3f115dac
z6a38535fd426a993f078ec476d299d388d49b45b2b36d76f3d659d59b646ac4fed2865bd0d92fa
z586a152c16211d9dec0db2b4f2f46053d7b59aa65afad80b04f3bbf46bbb516d4b8513e655e8f4
z5a0349aec3e6bd72cb265ad66575708884f2b3d19d3b2a7ae82f39b5acf4d9d3cd6e71d2b072d9
zf5ad36622f24252465825e56ad1c536bd420753be79b1bde30668bdcfc0cac71ca12634b4d2999
z7558133bc0032cf366c8f69f97eb6464f720e5fcb6f78e7d9092671a4d531fa87fa4b3df20dc7d
zc92e7d4096fb22c166b6193bd8b780bd6197639caeba0c1912a29a7b76758c0749871b32c20912
z19b3dd40aae34c62602c61af4fddcc785c17fda47a6b512846494a3666854772cf0bdbee7c6ccb
zeccf6a9d2d7355261f6da849ad7851802c428fec9167d42c54e1acbf1d8ee6b7e2947189e77a99
z3e6be38362896855d0e70350b5a353a705bd972782ea82700dac369ced43ad935ad7990799ff38
zad65f082bcd68e01ee160d4693ae562106558428465e370bfcc46cf1578dc8cb667b3d06709f0f
z71ec61ecbb829a86d9be2580c88145b2c9601328704ab8f3efd43ca306e867d78e8ee8b6cb1196
z95c33686ae4d24897f16605374847d1ef18f5e374b53ab803cfce051eda926dedebe3eed452107
z1bb603607f56f5b29c314c07bc999aad63353168461fb1fd29b4aa4f93a77c202a1a5f92d1ed36
zdf0a6883619d0f70423ee2a9ec546d08ac0f7c29cf53ee931b20ca5b83550db1389d2588d235df
z454524de09ce624c52238f870bb1e602b5ae231d64871d8b94e315b76848ed829568ec081f4358
zce1e11067c7b52a7e297227de24c10bb407efb7501a969f5b0d385e820b332be3ebd5382414d8e
zf0979945674e377f100b902506a3ff6ab38c88f4b6ae9620e28647bd9ac12cafc30053402c5adf
z28f75311d1d71001d4ce2f7848d018db2eb52c7177329745fb5842095b0e5755997f85744f6959
zb6c55e69932f139e7ed901b8daab6b3e3f0e7b072270ec716323eafbcb91a9f15d9ee201a969f1
z3c224e3f5bd41e7926e3c0755a95861e23639e14e654471884352fb91e3f77b47e930f14a6d90a
z90d07140d3f01b9e63c2e1970fa034f71ce3f1a55a31a30127dc6f8627f38f99016c1bac422308
z6715750ffd5aaf2526268355a94fdb88e40337c2eb5412ed744b317b43f386b6b23aea81048b7d
zc77647b21844d8f863c7b6a98ca7f0f0cd008635fcfabae0b4dbd66024927bdefbf617025de865
z96df0bf9b6b2caf44ada05b23598ab34ccbdb4b956c5b12abe30a8658b41127054197a11741e17
zf688bcbe05ef6493b3614a59bfcabe151c2f4b4de8ca779bf789fd836537a573f298cea1bae9dc
z28725d663a2fb07cb989e53816929adcf794ba19266f2f8b5cde0b40a74b919bdf5a8c5b435eec
z68a0b8ac631be7acc1a475b3c9abfa426e4b4f408e309bd8fc75a56229234e8c5c7d3fe27cbcf4
zc3fafb9d9e17011bc7d093479a05103f5ff48b63ac097ddb941c0cac474c3044055a3d1598fdfb
z2843c8c9ffe44ea20688d8ebfa70d232e854e16dff9a1d33f10be491e7e3eb3b47f1c57b330780
z8b998a0cfec06f104f1902e8b38298cd8b933cf7cf5bcfebef27c8bbae0b316432b592f9379b88
zd347ff53ec29b668f9b4471a1c4ab84fad132f6fd6fff9dd569e2c27fce419d3148a6dbf3c4fc6
z1865817b36c55380d4d93d8eed0de26c3678ac5649820f0c90f1d12338b3184d73b3d300fd243d
z554ed2b0504c936ab3f29d10e87cca721dfbcb91569b7f31a6027ee616ed602bf292d3520f63fe
z7ee07f45fdaf3a875f097848fd2a021e4b0ae53e5021df328d4b52d837036a746e6af4d0c92d2d
z37e75f6fcbe292ada945c195c8a93abb982afa55ada933b7f2511ffe95604694aec33db8bb4fc8
z2fd6414ceacf1eb2e6a7f1eb060a68f7fe3a1d39b5da8c4950c609e8549a9a09adab1e96e8e1d7
za3b55104ad54a44f54533b443082ff412c923599e59347d30da8246b9ad0aa767094ca29b4aec8
z846c3b2b8780bc966dc5a0d14053b7988f40e3d92e4c6b6d0fb48cdd2817e9d4ff0833dc11f2b8
zdd60943b59259f680a42d9c7d34e432d60816e514b7ef86f55b45e12258c82220782869a6429ea
z1880297edef492c10a412625fc6c43560f6f9308267141daf0ede3a9cc086a478058124e19dcd3
z456603d324b25083f12d29fc8966e2d0e07c876d3fb0f3501e3f97a9fb1c7fc35307eb3eade63e
z245f9d844fbbb3a5b0921136f3b8da7b1f71f2071a282e2b2a0230ffa5a846feeea59517818922
z95a28e3f9e72ad0381e4974a6df6cc62a43e66da6739583cb00897179a9f02f625bf91a8d0fef6
z7a89edb28f20e85a114c52f4a8ca210bad33ba707355093bf1bdd13ce67bffc8e8e938fc9e1cd5
z4379c78d8fca6076c61361db35b811199ee84403e87c9a17d4d0357db14a528e0d18449d402bfb
zaaddb762607d8d000e79a87183aff2483b25fac5d19fa6de77684e3e460fdbcd788c7681692b2e
z6a561d619a995a3d466ea9daf9e1db76f44fa129df25cf063853a2ffe4ae508afeca99e593ea33
z847505e6f9dbd14bba1974a6f31a787fc5deb2d0fcee5b7b9a6491a138523a1542ae6986070d92
z72b261fb38e25be696442d862749758cb181486a45dc64af1758e1150973e084c156ea770915e4
zf7707d0e97e0478fdbf48e482987ca5a02ecc8a7981f214225131e59ffbe66d1bca0645c0ed774
z918054ee1bdd8bdc1c18f62ad7b7b601692517804fda239acdc888daeed6325a95e61d97adbb20
z131784219064574730f6583f599b1d8219af804e299db0b4b301dec86cd21e06a89451f821010b
zd5db97c08753a55cdad557f00bad1e2b328d749b3e603a04570a12e49b7313b91e89d9d52ecd39
z54114d91d9418f715a754da02ea8e8fa2e45f6c204becc4f4486bfdf0c7164d431a707dbf25156
za07c0e968a867144071ea4f01243f4537e47a7bb628b3599fcc4698473ff8da5c4f24d7de484d0
z2e9c4fca654e7a69a13b17778769e2494281a3d54fde790c13b2a208d601f65d17485507ad41a2
z1c5998f40c76b0addb81fd68ade4b95f9470a08cb4fe94829e28449ed159dae92a636029cfdc36
zbe66aed5f81e53c35ce677db5d3f4e06138acb468cedb82ef1dceff5945b241d5fbb8b06f9838f
z8838cf9a409c03c9133d5d56fb893235914e5054f1a64c8ffcfd05d2963d46f5117e68348c4d25
z5f2f62937df69daa25dc766cd5dca9c2b78b7ce08009105a5d0c675f62cf1154707d4f9a85714b
z3d34bda49ebc2460c750d1effcfd3861351c98085abb826b47060a0a92547d3ad516cb581bc9e2
zd9d0cefdb26b474844ff36901f0a08dfd6d324cb0402c7a4c9076a287bd4a6d7a3556840f396ef
ze6268a1c4fdb1e7a2544d9a30d49fb280b61f340b9b700376e5b2c3cb8b03f1551a26ca908ccee
zf68d90288b7282e3a2a9e23b6cb58124c8c7f961d629bfdbe3159bb1d61290537ff4b3f7c932ee
zffec54b3a38c2a79f9a339a343fcab2c6ba2eae238d76f6c3cd03894454e71d5f9dfc0ce19974d
z2b20c531ca5465a8698c4be774c5a042bd17f103c054a073a6b86ee33fca4c8f43e8778e88c067
zd3c6a0ca27c8ab6928e149319ab608820784d10f74f294f2224f2f5d7170c50e3ee9acb9fb2e42
zb43647dcb4ae4518c359198e32b5b2c092ba7fd508fe50c7a3ad15d5f77b58b5722d308d25e4c9
zecb617178e6fc0ef13f13e0ff7939143ba3073336a95787ab5873091d7269681428ed4e5aa5a7f
z770168bcf6abe0af517d9a7f881649e090923147a043f06c0b426be44716a3ff01ebf65e92eb96
zcc0c83d1e1c8ac4f1ee4ee67ab85320b289390d052e33c0dcdfdc9ac97e050def5ec2c67b032dd
zf8efce474bea2ac52246978b635a0206a302fde693174eecb28c2c5def9cfbce96d92697af3ccd
z8bee51f592b6eb844faa74914485889f965c6ea89fc8351483f8cc231400b0d8d9b7f381e52140
z92d87205e40d9c55d4a94c5cd28743a85ee14cf8dcf62cd4f21133d2a863414ec9ec672b4879ac
z5dfc38e9134937d234d821b1904308faedc132703913f03b1018041ffcfca9effc69d2b0ca8a56
zddad277e2ab199fc751a81f2814a82f42522ce5892b29ebb9bc6e4ac3340fc21e894b2c5bf6acc
zb3cae6e24c938b6cbc865a80aab020e561592abf26859fa23fa4277feede5a6fdc4237762240aa
zc2cb6fe13a73ec912b456fde61d005156878200c4c31a52cd02a6bcfc57a0268ac765b4f349caf
z2ba7fc4a03156e8b6302506e1561ec05f1e5bbde85623f620b49a9dfaeb0e248b215aaa9b08dc8
ze16d2dfca52576bc459a75486c8f3b9607cfa9f8b9e92cac187c263761a40745dbad0f354a0622
zc3c40aaf5637b1141bf554dd5858d3f06253d1d30c9051604b972895d42c48966cc516bea8814d
z468d107c396c7374219d3adacc8351e27c5338b133d6314407643b9bef56c74554fbae7d6ad835
z72110a66d31f04fe52ff789f8d056796342704be2c5d737fdeabf45d6e42459836899fc25d9ed9
z12a61f422ed71d78eec8894a901cc417d9fee2bcf204c9273d48d19953dcabf6735e33d82a9f28
zbcfad520c56791ed6a53e42a4d76177ed34dff0b861cb4b97e017013285f9934ece3b30af95e1d
z958394569357a454585cb0a13226ebf15c2d975938b315e9d27c960aca64d9592559813faa9b57
z6e2dc060113477ed1571025cadc2ecb5dd7fe566886b0c7a3683589f4913f0f40fb4209a8c886c
z35934a4793c3bb732652db7761f118eec8592151aba5980e41735d8940bcd4493020299cb75c96
z018f0d1232e4dc146c090812353175d7a6bcae056677d808cc9aae6fc23b012999eed5b5220275
ze73c1d2e61a27f3e8dab7f69b202d392c7f85540d4e39f4977de160527ef8d6f4cb81ddb18b9e6
z0464641ce261ee878b4e6a7ba174bbce19be1a369754783c2e9c25e970f2b28a61585738aac4e9
zd55f38e4a139dee87cfa5b1f68761e0d7970a9cd8d9a218a761ef3a3641b859235ace27b40be81
zd41b2c146706fb294ed213979af6eb27267680149504432192d5e98f92ee4f1d0ba3b46ca44252
z7b84033ed967b554a8097677b68052214a758cfbec5e55395dc1398d3034c2098aa63669d1acf5
z1607419ca7a869a0e8d88028a81f455059c62da115a8eeda34399cf9ef429cb9a9933587e88988
zf8a2eee78370a854f78d951b3a7cf397a68e4c254f21605bbc55e4abe33cd363a4ce9b4d951440
z74e9a51d231f18b7ccb6322ed2172f0b56fa486169cb7e8a47f2385f84a129f792ccb172c6ffce
z0d21fc39f27ac213ced3acea1842a9ad7d9a387e5264267eb6db57d191e421c38917b49ca9cbc5
zaf2b4ac7d7ec0c983a364c36769c12d0f02f6c2b4038fc4ae4688ad8201c03dc1be7c020cee132
za3f66c68ebc82cb3e6be2b9360f645797683ebcaa7e8cb18ca394b645b0181c933f14b8a91c96e
z11334784ca749b956d5c41d55be94080dcdceafcd68aeb160398d529f9c7ae1a24ff504f940584
z850f1748c85668b32fbc9c8dbe06bcd79fda35fd43a52f621811f4bdd31f5e7d928fa0a3973ff7
zec702e4b23abd73006dab2940e71287e160d48015a0718c444cf9caceb7876982a469d98781f22
z11dbe447c51d141371dad7923a9d75b42274c32fa4aea91b1a82d66499cd047b1a9a48b9428203
z8f2e9298612bd2857646f3ad7ea2bca1424746ad20ba0c75e9dce4c7c6fd942c03c21fe40fda09
z40dd73dbc240d24d90dfa698f422a7968d355f947fce15dc96ea4322edc96681ce5fd315333034
z5a4bd76cb74121c6fee0b3022ceab192e4532ab0d6aad822969de03663413195524405a6640d4d
zd5e5fd4b89d9fc69c52c20f214057197736f4b5cacd725e6b2465fae6445340c8b7e5e88277b4e
z6e18869a539093f281fdaa9e5eb22a87335575adbfb934eab49b3bd009c88ee0e93e2f61a72d0b
z569003c0d6453767db293ac24cee190628a59c79396cb6731df6d950ecd2ee2d0ceb4bb0c057ef
za6455fdd78d81991e4c15491db9d5246dcdf7b601b094553d2e433ef4dd96a6922486426a83f03
zb541c5fa3a2003ff540874957e55afa04968fc13088c4e22d57d9fc57ffd8672f7c035c5dbb344
z1c666892437ae50411b1f097b3adba6cc18adbe5d84e4aa2d65b4b411db44d132862b8e83f7d00
z9dbe1a56b0677afce61981e220f8f013e59f30eb1225d5fc0b3a925b99e1ff71cfcd3dc4de9fb1
z747f5416e1f1447cd5e06d70ea65e08a492d0c7c6f27c13eacd383769b151e22e4fc325f9e93f9
z852325b47e8b668a29129b0d4dae2e2f784871e9bc948bd55dea43d0c8125fdb2dadba762f39c2
ze0025f82301010e35f5139a24daf8ba1f36d9b0b4e7f42f2264e7cafdf83fd478cd54f1463800d
zf7fbe2184467f667c13d338e204c3be926aba263bde6309a7651cc24e141da7095ec063591c478
z7b35c3f2b3814461035ebaed477525a60ddf3ad610f4a910120671a53c55f1f255a19fcac7bf2e
z45ab9a6cbd44ff573ff037e8cea0a20b907668a7d878469401fd3158d62744ffcb832d26eb7053
zb9759019a9b6f718251a89fe683edbde21e97b84a6cb9c41aa3a4340dec875dc176b276790abfd
zfee0d30c2aabe26a88469768dcee0e9810f9fededb9dfd19e6380d194646a032a16aba9edcf810
za77cc03200eb53d4ad950131edde5d621f6eff324457e04b3cd3c76642f26495bd462179dc003c
zd8bb5eeaf108dfce6eb96197b53eece6f78e29bbd9d108f71a243d70c0fa31d064a73b8db69be8
z3a042a8ce32857a731184e28951ffbd15950ef3d5a913b77ba3e146746edaf2bf4a1a01c14e8e0
z6226f1f4c1f13ce309480b9ff13a23a9b55d37e9bd67f775855017158d7835000c42777f2d0e9a
zd15e8c2ab1013409a40517e28a758dd870454cb8f9b76124f2eb219f73d4a2c59716ee2a4422e3
z0e15a601e8c5f3f0fdf765d09c482a576d0b2451c9c0778725251d0908cb8f58165f5b640cd026
z5770b44c655f53d7e2cbf744642e2e739dcac10d60b9bded1b6e42497d2bb967cd64024267de99
z75cb1762c1613e6c87b93c9eddab42776f226ef010d91073f7ea689b63501fa092682cbe700eb5
z5fe3d4b615b490916ce3e91da4e08afc4337a299ba1a68bb65ef88032ebda0ef6a73e75567cadc
z5e27cfe4221e332f93012960ddee51eae43f5898283c9be5da94269d6b901a0552417afe34c550
z36e1c6884a1aabdfc4b6bb293ea2814832ba92e37d2a3a9f1c49eb7c7598072e3ea3ed048fe0d9
zdd10e5932fb48c91dffc697daa2b4c0dcf2adc8301101b96a9e29f3fc16af6a9ad07770be9026e
zc23502730b20e283d34f8e4b43aa0b430538d64137fe7ca81a18d353f2f0a374d1e752e268b5fc
z146b72ea154ce4ed1f4f14e5f27afb4306e3105d246dfe44a9829417245dfc3df316c6084a7c6f
z70192a352fbce7963d73e68bb071db212f1a7f3dd977e1ab994c6006dc5bff1450a633189a56df
zac33af012e70c225e7663027b9e2380f610e6184222070c7453e804ea0043aa502fe06eeb03b17
z00cd2b4c222b5b5bf05acc750bcdeae65c1657760ffea9889155fc172ced5a74d99c378757bb09
zb8150fe493086fb1f43f4af40973865815e2fb6de5bce98ef2707c5f72d80f0aaeeddae54239c1
z71dc2cf5a741f2bc91906aa2f28626883ad27f89c7540b5f91a0ddae9a2dddf9ddef7a3c3c92b8
z55a074ad6e640a87965f0f7880d33743cda18dfebeb9549af025342efda4a763d6434e90e7cee4
z94b30f38ecc1a01c5d861acad27ff26adde965155796f1a5e6b92da045e4ba170300b61038a912
z9938193619604bf75be9d6ce19f35afce24dc0037516c164e4703f518bd07009ff64adbc4e63bc
z22961e31e74d19bb121a8d1ac0d5591a93e89989cbac64290d966c60b7d9837b70ab3253974a5d
za8940d3c90366b3f2ac3a35819d722582a2571f51fb274df5c630fbaf0b44d34cf94d4fbc3c5c0
z2643891e37be6321d021324893d32d946db334e4dee30b71d4a5069a6a12b2011afe4c161191f0
zcbe4db3d756e1cb432a7061717840b665a46a85f31a2fa740900323d20bb378ebf9e7f042df17d
ze7f591f030182d8e541958a83e84814cfd170296332a5472c93e6b59db251cf44cb5bde355bd3d
z46dae2e0fd99926c33344219c99ec99c8130cb70c3bf5065f7dbf993d2e5444d89f667ec371083
z70ff68e1ecfce09c380b84ce4b8a8965223913588109e62382c292d87c6aa13efdc29eb11192f3
z68215673e97156ab861efb3f41419def35b23c261c87af8779e8381ee60f4f28f3e6db70c88d97
z1a8984cc10a64a598465c3ac827c02630e28014015ccdcf4b9f9c418da6df9f52185b6517b0cb6
z75f70b2e25e0435ada70561faaa03a0d5859fe6a8b0444d0232570e14a0be67d100584eb3e5291
z2c721866932cb3cd29523e658789455797ee6e789f83472313483784aa7ce85a92153d3a3e6c2f
z1722f3afc625c8abc4f83eb60696963fbf5b0774c6aeb1f72f3880e4623889338b9d87a5f1e240
ze96309227b72da3c58dd4a26b9678295a85de283d271568a7f73d5e3e0fb1b54c8e330afc4fbb6
z352971af97b999b7d0e1cdc02a2d8d1a58e2bf77abe3c26bb8c48f1e346e11e11a411ed4bea72b
z6486bfa7b95d458dab6357bf71565b19ae1112ccb870618c5d1520a1a54ed1e3423309af0dd553
z93da546e6519cc0530eacebef3a116d669839380f6d3a3fdca7fc4ca496de52d01a6a085813823
z7a00f3bc3087e417e0ca0eb1d7997fa92015730d3b18476fbbf2a56164593fe9d418e71f00740d
z9a81bfecb37cee45de2e62939435c61d72e76ec41967ca87d8c1ae0382c130082160c42605d355
za82fa5e84df0cfe90470334236b4312641c858aba748a892b90e78159199243611753c79bee680
ze01f0303131a6f76d35f4b52c9f4575f580551d5616d761217c02d637df37f6d521d9e069eb915
z47a7d40c949ece80db617c64d5019427063e47f5b9d88d8d6ffe2196686239db97e17db9e09acb
z9288d1fa2f27eda03c3886608e33a3fe275dd5242badba5779d06c25e9332e64d76f6dc4466135
z63486823c4b727de4f517c9f73f157803b64f2d11c7df1af0776372a4d6a5c50da726b488104f1
z6bc72b1e31811d4f1e59d9f489fab9a77f79b933da192ab4d0d3d581715046cf8ef91fe911def2
zd71e02dc50cbac395ceb07216fb2e15d3421a6635cc6ab198b6cede9a2d4026556be5b283246a0
zf6ea16cd6a847780845ccb7dca10e7b11082dfffffe57115ab45cc406ae9c1f1affe23a965c0f0
z5979625035c758dd4ef5cdaee26cc53cbd1f101a85573dd8e7ff23cacc8e8b96410edab27aca04
z2337e4a227ccd6fbb8f644197f11b84ec6a3e2549ac0a147a56420f4006cd267e1abd57e9f206e
zc2c29fb8835d3de20c2eff3325b89078817b01ed1dee1fc4c3a8c4728e6d537af4a2cc3b21b654
zf3b5fbbfb1991b41b5ad916fea50f3aa593218f37c043646e39115b654232cf1342ec378dbd7ea
zbf3b935e2ae672289440ea9baa454d39c3e452db38c429802315bee88d3204b0934d551cfa2f5b
z93bb67860c614e19c28c4526bacaae052598b3fd8f005070fd941b5f2c0c338770d49a45db595b
zeaa9f45a471d3c6c01cdd8ac23f39472c851618bd8417a16c0b7ee84e76753ec47a02ba35e1760
z515ff3d219c19dd920eaee496aca81368c98190424587f23473dc6948639db11fe97572c641659
z027cb3f54c6a34ce15f8b80d7a63a2140174e57e694e82cb0b8f73b3338e35d0bdb48cad7dcb35
z4f95a1a25ebc182a5970a09160a996965941e7b7f8ac251a7c20ddb0ebf92c9fa36475d05c3a10
z1daf4d0dfd154337b6766e6fedd7b259123d10013b8621ac0e169c220c84cdd6423ebfc814109d
z0e5a7f6b1064efe6fcbd8f21e9b9f5c2a51bebe426a005c5616d5e027581dc64b36b693fb1c325
z4e018924ea3f3b89ae36b609b0a0fa27a4091c157889d615c5aed4e3084a54a8a72f63432d9e35
z7c72b649ac8d4b931fc9e1b378f277d0b4fd2ef77b024a5a09a7f5f421e5f21f8828f62c7b13c6
z29b391a9bc7a3b8d268f1f2848c83c44d9064ea1494703fd5e4d1c32fd661f17dbf93e3f4dc8a2
zbfe53530d725c3da33325a54362efe3ebd5104bb9cb3aa1604bc3d30313c9fee25c06e0f6c320f
zc390659f24aebc96c819b5000987819f39c0b98af129fdf035e773a6c2f84deadcbd0806407ace
z04a0f78e5a088848d3b4ae23a138dfcdcddcbcc94a928b7311bf59b91ffce50a0d9d200f27e8f4
z038d9dc80c55671ed9190efd6b22ddcc6ca7b77916e7108f97b12c287877ddb3bb8ef5d4fe5971
z84e57ef772b04d6e7b2bfb31185d9403222a72c1fc95e95dac4a3776042667c4f6638544329c55
z31d76474c1844db8380dbd6547a530745f9b24bde7fef172110cd18d3a182d9565d3713ead718d
zf1d72a6e0e6e832b408dbb36b2a45729cea86cec1757e6b52be28358f636934006afcf7f3ad0f6
zf6af705636695fb3b63eacd98843342c2336288f63c029c24f27cef8b3e671cf8f7d31be1aa980
z17c2f7fec7fffb221879dbb627b0a02e73896dd3950f44ffb9b85a9370c78a62616c83b0b105e8
z221842e993988638faa82159a26449b781b8a42b2ad5741209fb79e9589052dc6ce498458b3277
z1142eb9ce85b864339a96f96c613a8f831e3793719d9b7288b81a49afacfd890137a878de756f6
zbebde19327eb09f3ab055c4197a6c43149c2e75f9de4ca545d67e0cc70df42ca50637d46e0ccdc
z0bf2f99e3a814f28f13d56e979c5c8690a4298df969c36d796996a71efd02fcc455d6954916fd3
zc72edcf30f112f73a2f812d83cf600642d4b8324d8ad71c7235b9ec9987121589f59f44d6524f6
z71ecb070b662028ea36fbe4f195f67fbd8e4fa5dd772b96c8b7e98a6191fb76e57f2cace6c3f6b
z3ab67fa6ca138e780c66211348147462b540e8279320d3b79d6f137cba80ccddda134e2955421a
z0b94b6cd4adb8b4aa7141390d64da9747297c6f4d9e76e200857aecfe64676a6ffd753e0952e0c
z1e7c09c33feb376926f2406d9d0d5535011be052b5d0a1d3aef32518f340d5e90c751026bceaed
ze240f8b249cdf589a4b214dc528b36699587d4ae6825dda9cb1ce09ab41a9ba8d636df146c42c2
z1b503bf40ef74f84737238ea11de253ca426c955c6c6489dd6935d3c6473f2ce200f83deae005e
z3cd9cbe96481d3b49804b971203ce33e78d609ba6b85ed8df3b932c142e9d95b3d7b6a5634b3d1
z0eda27eb2c29800925b7d31b0a8092f39fd6b02ae3353e742f0ad249d30bfd651d4d19ae730294
zfae88c3003f41a44d034188114fc1150c8ca9c9f7112b4ac20a335ecab168009cb70c1cd888e05
z6fdf55cf67f179ed728c661568ee0638134cd95da46b3b0ef2d2a52492c1920e0d1a3bc9f11e71
z4f6cb6a7b78c666917cb497def9a60fe1855e9c0b2874a29b3dca1872e085a84e4802cab167073
z64c526bc0ae4070d76a36eec13f03eb69413e8b0ece5abd35570bac22c84a5fda785bf41b38966
z75dac767c03f4bff2388408e2c81f6cbc0d9055e3e1be46d1e92159a04d1d86ba09ad0ac262bd9
zac7cb8dc3a0120557fd8d367c1f97175de6b969c3ba36b1b413f29ff845e94e20668b2686dcd7a
zc925dcb18f01366a5efcc603e6a864d53fd0d3a197efa7cf10eb4a097abb0cf0329f723500dff5
z27f0e5b9c0c99c903b9478f41d06cfb7c1bc27262641ae89a98a51960d35ff68ee4b3811189939
z4a8a59ba2e1109256a7717bcf3c99fda297e4ae3dd6a7b2318ce86bd5652af023088776784f67c
z42acd2c23bb6f373407409b98a9d4af8a8b5785a22b0a52af888362d651cdb22cdfa60eb9f2877
z4c98abf423703424fa7beda3d10e7427df98b4653795ac210359dc9e33b3edd7b42737d8f38340
zb68025450bb5cf95da31ab157f527f26cd4c3d0882ab68544034c5ebc4c31bb61ba3d9c51828ff
zc4e1912adb2857d2760057f9bd33cdff212bb6c899fab4bc4b07823e54e025b8fe87ce799d2382
z8c3ca73f68816148e4b8207c4a5b061f01bb5d2bc348095f012be917eb5ddb06d5298f7c482db1
z918a6b49a153e6b049759794c5037c2dfbfa85a708cb0d2e12569f23e02ca126a375250f14b232
z4c2098c5c087466e54d5d948ba2df65d11e66febf486670a9257e92e386a6cb03100c57412ce74
z8a5940d76fc77c6be4ab2c6d8b3e3936dac53b912dd38e9eb1e38ebb62c4e13a0901af21ee4785
zc666019d495816d0b12ffba4781eeb835ed68d2063f1b03e8d6d99dfe8b89f4d40e4bd651a7b97
z15098e75bc5a3f2fd7ff72d5368f4931d031612a12cc66182d36206376829607d86145cef29e4c
z983859d9243821191f83f8116c78c648a620f075a741033dbd61d9d477964deb8e72664feb5050
z31951c52ca53535bc95870cd197bdc9b64e5abab66472acd85adbc30c13345ec949aa5bf5a1ed4
z840ac4be098f5babeb1f6995e1b218f5b43db77d978ed4f6a49db436226fca969af352bdb4822a
z62dbaf88638d301c663badba4b8f3a953d773f350cf9b73e50ad794063acce8e08d65214987952
ze31961ec4c64550be71f391873eca5b0dd36b25e44d59f903b53571f45ede09eb98808dea96f2e
z2642cb5194776aaf7396a6d9cdaccb219a2dff56c38b82f7342887cbceb64b648f0cb28249db47
zdee253e1697f3a17e16d87de9fc873ef4fa8e7e05c870d265c4b6f3a6ada47f3acc3a43787f4a2
z075f30dd5ef516b97975b4cc58c5df7f998ed946168b5ce546222351ff896873a9a16f56e6dc65
zf72e5df08df66bab4c240e10daeb25f672a99899c67725931b3120ae6893f54831e38b91b5fe7c
z6d5ffc4a2efac5b5981f84ce8386ff9efdd703e0544eaf290307c307396e181ee7a2d9b00b1f9e
z59e312e6209416c16d6b68d8e418b24f9dd635131668dca18159e26c35ea50477b1475394b3672
z73e3563895790847b9a71c5318dc9d295f95fc758fb02e50a891cece38e2a422d1ca0b4a7acdb2
zc2aca1906af5667ab4e3cf3a3e86cbdf2b2a222f968e4dcf8297da777fadf6b56b41b897487ccc
z06443de40e782fcc394cb3d320651a51fb9073da03f03aa56406dcb58324185cbf1994621e0d6d
ze67928e6e377e1759575448603bc882abe773b8c9dd786299684ff50fcd6e9cd6a864023fb5a6b
z7884ac063d6296217ef7a6cb2bd64cdf69ff5484029f5e766097057ac20d249295d2584ca3fb79
z2a41151544d5282eb98463b51bdc45b486825c9775707bcfa7a80aadc4c839de3f3a92fbf72782
za0cbd737dcbb88964151ad17dbdd8229465d0767da3940a210f9a197ec86d924ddfd4661a812a3
zb4e3a2ec096bc655b7293ab8db2ad5e2bdaa4c1e0f2181f64b8ddcf2ebf44b932294c1d9bd6e0e
z4a120b755ef51420f8d0376e212208d6da60cff8beeddcfbeda5ca19eb2dca273a404f0cb6b986
z995b91292884a8f1f93b50f0a6357a0be1bcbb51e11f9aa0e907b13c4be6454d5838e72df98a00
zcc554722e8dc03365f37e2f4e8e91eea72bdee7e436dec8b412bc4cc6615d52046e6d9304d4cee
zf2bc90cf3738ac3746ed3410af8712e24bfd16b29db5f1a287dcb839becb206d9b2f5fa56f79c4
zc50ad2317568c7ab183e0f518087e011daf0f0aece50bf6739cc1b9cb9000da13261b0e1e14322
za31378a59438aaddcb96ff2ee1161e60f37104f81f7245e74092dbd222cfb1c01f7cc9027ebf66
z70538e7ccd78271f323a161719779dfecb3789dc4a0e1e46035691cb8c20388ad5e8093e675a10
z875ead7a2626a04144947610078ecbc4976d405d6438ac84726f1896c1b233b99ddb409b20a533
zd40faf0bc469b13f576f6c3698fe48ca5f1601379060dcbfe59ff33facc66e18f58fc5142610ea
z47f90c523b4885f2d3379926c37948eb77a8770b41c641c1126c078c299f92729f3519256160cc
z75de4f8630532e47ddb74c81409dfb5bed20ea71dc8c8284a990d9ffa9be8aae231347c5aabeeb
z9d481c9b2c391e37225d0e72fafcbc14f2da53229a486c745b9a0298355f61481fbbca5d09f529
z5684268b622b8e3581e17cebe25b4ce78f94012174b6af433f3b217fd8d6bcb280db45712fb79c
zab03893d8d456af284d1347501de713bcfbdd61d80f05286878e42d8359c7154cfcbfbbe3fc129
z5873af406948905d82dd17c9961fede94461a11db7f6319febe39cc5c270d8577fbec363cf6968
zb471d9af6208040fb14615445bc06291f6e77e831c44395bccd1981e09a0ce386eb1382b60ca3a
zf7f5c1ecaa22dc2891691e6d46eed24df29a3b66c0551fca17a194a0bc320d0a8ac42c9597f7b7
z7c350f66c69b1f0c56dd3fbe306e1a1eaabfe6059846d7e9f1c77183058127ef50e5c2ed2dc17d
z0235ae13237dc8e4c67ca7a89a0603a6f3669b60db58d8ffffda4b90bb9e0396bac124bd1c566a
z37d06f3543917893914d537eaaa87692443d3178d462d011f8c588ed6da9cf2c16bc9606a5e1f6
z234318721ba6b86a7f0f098e3fda6267c043437f5cf7b293a188d8a3f032f3e24bbfd7236548ae
z70199a6e7aaeabcc4332723434e6ca2cd45b96852f284b2d5bf192699ffc2acfcc1f99b731c17a
z2967a9081fefc3e5fdcdb39f2fd5d37a845d8f068879dca11c2416e3b767d47490e8bc2f0bb3f5
ze680474a6515dca9faaee39850583cbdfa0eb90c1b70defe6e545609ab0b4b0d2962053cb5a08c
z886e68b4b8144f8f2ae7f24594a4bef3adc97bf820d32c426aaaf3cf74dd9b8992c8d1864b039b
zbae245fabb814a47d2d92463569eca452dffa6924690f58b735b60f58e94fee8e5830185431815
z84b2411ff143745c2458e0364dff53227ea5f64a60d4464bfbcf4fc85244cdc60dbd7f8fa5498f
z1214261090ded5bbb285e64f3a68b8e4f73a149895299769287efd82282d352f01a96febe9d931
zc3dae7973c8eb212bcea05a33d94743d4039f896b4424d77b86ed4241acdd0beb227f022764db3
z7fc37efc5c4f04386d2334240b74a6959f4d5e27c129fc9e8f120ad78850650612cb0a7fbac095
za4455103918b01f037c9eaba588dc0a959a48be4c209137733e6941eb485df84b2b8331a31a74d
z12384f16b92353f72745d970c9d81c51e2ad0589bd7330145fdf72ec8528e5a87503a63772394e
z2ec41c3dbfb5d43cbc698360ead76e441936c6f029f52d23e471def9aea4d5a7ab7adbddb5cb3b
zd0f7916fe64d8f42cefe3a81428bafa2338f4695fac5a890026d4e3efa5f69857873ef1bdf931e
z07a81a912d874c2664c732fd784222b65e9dd3051dbd0a7a3e0a4b27f843e8f7666c003de6e690
z49c0eecf568d1a0711853a65c296637dac6e09bbd876803a6019408d6e2ef7208f6c61576a244a
z5e4433b597c0c663b58683f815fa9f84b9ea88ccce8d266c9692a72a7ce4eefcfec2fdcd289fa7
z16b1ecd1cb2be9ba9afd720f75987bee5036bca57e3d59a371e37f112e952cdf4a6f7a4795cbf5
z690b511ba04fd0833b43578f116ebb2f7860e8ab198d6d0e9d18d461fda6b7452d60bf41b151e7
z1f73a175f2029ea2680ef20c49e9c3c6deba03e49f32c9b93e0256c27620f2865f52598be8f42b
z5fe8b4f1f64b98701daa2fdf39cc289244d6e96eb092c1540e2e586d8dac6df2c08719d5c6401d
zee4fa276ffb2e5c7e9b7428c04d7edbade8301dae4224329e646805e73c2777259fe8ebc1a9519
z9fccea7a146f53a4a7d131a72397a9c6029916fbb42f32b6895c3316572e4af6e91241059390db
zda1694f32c6cf376aa0f4e27b76f39930dd59e5c17d2b0aa97138db7b1623dbb57b78202da7658
ze35f95c297eb43525df646e4ee0908441e437ab2a3be7c16272db707bfd7a64fcd38c79776efe9
z31504e97641c576737879d537072d102c0ebf17288b8e0aeabaf3dc1d498044e40069405633df4
z10957a1495c54776bdfc1497ec8f0ef410d54e0b8326300fbcdfdf01f17ab6eb8618e460ff4f45
za452d2f6fa033223663eec131cfed0dc7e6430da02d6c42e7befa50c76c4000b62cc1ca0dada6c
z33efab74c1034ece344302a16095039d850d69cef276dcc523ef4d476317057e3d805c8659a787
zacd4ce9f9ee871066f0035404d4c91e37cac7b12cf08d340a2dad46fc3360eb5eea689ab5ddd42
z231fb91fe02df38db014083abecfea90b7f5e74d8c43d6d2706f04ba3520a93afedacc8b025717
z9ae0ffc1efa96a9e5378316f688e67f79279923730663814e84cd61c774cb18601f82b386554a2
z57806cc1ac7202bb27ce859d660f73a05bcabfdcdbc534b3113864d90b08aad77afb495456d643
za2192aed05e974c8002805e714e1fc1eaf47865fc96c2a366d8bdccc34e983e5a36ceff6219333
zf05ef5f384527c79cd564c0056869e0ec458812009e78ecf725eddb7a82c9f78cfdba0eadd7143
z5d665d41bce0b30541c9b25e3a0830c3fd514ef8598a5b8cd22af663387adb1e23dac2550f479e
z7c75eb174482586395a7c56e11ca9db614a37bef6ae0f560d860ecdae95e134b5b6ced514c5096
zc90063b98d5e2783e6e93e96df335d84c5ea18e06f42abaf3f4d23c63db29fc038805b55b7b5eb
z6652ed965ac3b5145224bb309e042e7ca595c3db5854a86b082c4cd677fa0a8aa939c2760248aa
za7b04aee4c6c552d614df94d633d561cdc8e86ee477d21c0d5de95a300b6dd877626bedee3e423
zeed673681e542db76ee637e5b6ea27dcaf30865755b1917f6054010120c2796afd520de9acde13
ze57203920ab780ac8a8f1b1a2b52c9eacd479255d8b1b7b1cb039596d16f1b1431da4cf72e4fdd
z949bca2ea4ee2c5c93836254bad659a0252c66fca87d5a12c1f84c75039063c1d517ed6a4532cd
zb6a60e7f0e8280259caa1cb705c3691f6919491e2996377be8cbb73a7603d640c8185ca2b7a32b
z9a257c9d3425fe4cb494bc64c742309e0bf5ec65038e2203d5f6e74ca9f573b20248540b8653c9
zff144db386387950304d71d9503240f1e66bb7a31d32ebc7f79c2d25ba5158202ded10991c007a
z514998bc32d945def381e497c9659385a93a91659f022028c4595589e2a8941a9bc4954b1757e9
zed140888e2e96a3114d6c12d500611a6ff0a989534eb5d406f3d2a4089fbe6301d0f296917ddae
z74582e03bdfc007b207b3e27b93df6dbdc34ee3819a292e501f864afb0e1657c7e319a75589956
zed17f5d26764e42f0e937f87a1b6f973c741784dee579ed002de9ee0694b35b064142c7f5c3bd8
z7750721538ef05406ec576f736bc726cbdc47a5c7ac452e29656b1534b8b3b3c6f4c387413c248
z5d3d822cddd9e15276882da453fcc49e011cba98dc9a50bda38a9eded6ba4e9be676202c14a80c
z63f95cebe64b3c1951c7411648c56dfa9348f9359b6a97b6ec13048ab05db1f856b8643c22fd31
z0f8e5354d61d37025c9e9253df0466358b2e8968bcfa44f56f2ded74a5b4cf537d40c015b3ae05
z2bdf52c3f62de3342333f4fe0003166ba2f3ceda9c0739886cb313358cdf6ab32dc1178dd7b97e
z3f415a2173ba0c3644358ea8a4bc18429b0a6fa57bf3b77e3fb98f33bda46851bdfda51c4378fc
za50b2abde51624a52cc8f76afc07e2e401ab253e1870d999c5cb3fd0345e3e141213ecaa452e58
z9c2de71fcd8150230d9c7262c667d6973ca00421d71dd26cefbae76445933eb76c85aceffa81a9
z203ccb6ae0c5c597d46900cd455550cfa17c6da0bcbf1569c5d88e70b1f688e23f399d76686359
z9c5a7b1f9bef1fc405d07118e9ade04b1d49e72aeb2ba0be6e97932f9fb23d318131115af8550a
z57b189f93e059528560983a3ae57b364d7e0eeabad333b26da1851e6484b69e3dc29e15d4f5588
z45667a7e8e818035a0603e5d2a893188b9391858124541e7331ff0f40c5edb8e2215b9ba421049
z5c7c41e41545c45368726e4720f065b161e41379edc68d94945cd6268fdf2f21d6b67f060d5b93
zd428b5844330190ee6a7eeb6a789fcacb52bb8135127180f7fb71218fec3e2d18b9ebb6cfdc86b
z3841f2d128300a40a30c2a2439101a59ef95651b2baf6805f268bb6c8b8c83f63853c5bb67d4d0
zd78577809209c9ca72c9ef947578486079414020f6dba5884666045d6c66d8c2a7a7a618811fd5
z39b213d947012be6c9d71eec3b9de586b1b248e9d5a736d989c843cd067d236befe6d9b100e557
z0d8fcefa9fc8ed7806f480550d2d6d9cb32633b6564396dc0e22b01258c4ba0e21b41dbdd17f4e
z958b8545f61fbd765fef021f94d778a93af7b892dd10ec0910bef62bffc9696c295dc258028a3a
zbac5a9acd7e02ae96291d5fda3961b2408780afac423befc64a9d521bf8ecae9f065c73322a1ed
z3a83fcbe0ff184bbc6b0335238ce2fcea19a7cac130be9b65bdf7f0e7d2ff3e3c357cdd6419d42
z2e45fcf156fe6ad8821d0b6ea97cf19b9f53b394e4fe8a729aedc8778f1ec610509221551fc1eb
z32dfad4910e39be011254ed0c95d64e5c1eb6f12d058dde4ab1972949b3f8d677366fd61529318
zfcc90787bd2fa4f756e40f5e7bdd30e2b7b888a6d4adb40b2e49124f6b571fa710b876d7e2ea0a
zf4e8671d35ff8f828f195f47ca8ad956fd27bb805a594fb7da6e16a3ef588dcf2feda4ef3d5aa5
zb81a56ec3629da11907a86294c60ac1d44af89211e935ed8fbb888afc1f252b2872c5473e21c7d
z54a7b2e0584c30fd048ec974c75698924571c03ea9a852352e6f2e317b5d073c1f9fbe0f62d0a1
z8e442889b64827ace114a889efb16373ffd78a29be0c319e68e398f8b5c1e324d1fc392e80491f
zf311792116d2f4c89090ff0e749ed5b447a4c190b84603a591953e4e23f693ca8fe9caf5371104
z1dcf7298684a5f747e1f68511fe4d02282ddec32a84fe3d2ca24524c37d23a54db7ed6116d7ce2
z28a50d27607192dbf2351d1e500e676bee224a9f37290db6486e5df4d98df4f12d65bdb38752bb
z2f623488686cc08ec359e189018c13146b590d2c3dc12bc86f771d4baf1dfc8a38d66a48f96fd1
zc0c2168d61f32b80dafdc49164a1eac30513ea019e0caeb451e44e72f24071fc358397e84e0384
z8ab2f6ab5b84f5153386a7f8dc873718db52434eca4bc3d340afce6f622b24c2e713556d83b1fb
z6564ac1102383711ba6fa34bd9e4891ed06ff637f105d9867faffcae344218291eb3406b94925f
zf635d6a8a0e1cf88010523ada4a16f2950da29243dbf8f53750eb2f7bf7d68ed642321229c96bf
z51a1ee702497407426cdc6e10836baee2416687954f16142cf3a636cd4b84c3ccc8c2fed586903
z671fbaeb1e2515c3cdecd643f088597d83b6babd64aff976b641ea900adef39098659141066cd3
z932d84f05fb3711d13454430b4aed7012af5bf7e183f6c179b23e7301e51432097b53c755bcb6a
zd33b8be8dc5d34d69b390a7e2f70f5bc110e069cd9827f507ba1a93ab582cd92cc29c5e3a22b00
z2a57fea2de38379e4fb3d96178a0375368e6e1e25b941162ca11f3b098f9a969f403851adf61fb
z3bc04b6d2cc427f23881cc207bda6df4cb45410f70f80d8a066e2ce23d461a6e8d2bbf17c1bc01
z8d59f89565183dd3fed2891644a7f423726e1abddd0839e496ec700d2e997a044bf45df91e3ad6
z05f668767dc57deef233e0dc7ccedf15a13f1bbcf9075ba756268e13ad3ab3a7462f82499d77a3
z04c227ca61b2559210fc0adfb68ec6e8a70fadbf0120b8f6b5624a70c40a06272c1661fce4064b
z3b79d90b2d5f8e245475d92c0bcac3588c9939646e0011c29ae3106b6b779215aa3ff2a569415b
zb91bc4cf3f2fa3c62bf092c2b8ac5ba80726d276ac9b4a76daeb285b65eb4796f3f940dedcb21c
zc68c1b154442319007bcdb6cf442cf5fdfdbb769574a894d00efaa4c3b5865e7b80780f3889193
zdb39dc56ed340629d24a1ae65effe81f5da8187d7c18069e86d7c7be82cbaf8dfacb1b486b3d48
z290a276b6e1f41e08c34bca644df93925ac8ff894b530832d89e20fa519fbcdc255b50291f4db3
z9fb7517a59dea8be90bc4825ff996c94e7a171d07fc76b8757f32a50427c06ab55b7d653ca2fa2
z11af5d79b15654a1a4f069243084e2b922887aa966a8d4a478222c0dd94f1d9b3bc06cd75b79ac
z4459e284ec6562362b73e7d3970f1b9703cb48ec9d6b013ac12bf156fb16ebe4bf6f9ba77d4afe
zefba881e55f8ed69081eb0c824a7025dbba2314fc8ba73cec45e84d9c76e1c11a7b82f4b6620b7
z17b761ca8f2c670b6fed97fec5bc0be4351ff3d980af5b8845c831518eacd62b1044e2411cd96a
z5b93361c4a7a9647e06180532db88740d46ef12557dc4ec624ef3bd1031bd18227ab85cf959761
z351fb4b3d5bc1f8f18763b88e9486edc6ff0d9d463163c32e12a5eee02c1a75ff954ad08e120e8
z449d08442d7d98ff366f7153ecbccb25759d804bff565717b80b8bcbb690a25b38b0747040e9c3
z02284246f923a8787ea1f9595d790a6aa1a7bd04c8b4f79718de57fd8f3766ab066265bdc6311d
z939363cf110a8cef38b7a999b51f9fc840d282634e0ae1efeef9bd624fa0e69e79c7cb6b1d79f6
ze5a7f1e392e4f6cddb313a55bd386e0df4ca4e2cfffa22eee1156212706515d3c9377a248fed99
ze6d064c6658668f7a272ba2ce61f2e2cfd85c2ffa3801b1ee341ece2aee538bc03c3f545d1a75f
z971f18f6023f4154dc520d5e75a542db972cc816dd54116af79551dbcad5067ad18742a4a02fc5
za1e4407df68ddcfaa178d046fd8b5da761106b5efd443c5a6c8a374dd4379fa10a9cdd6e1ed061
zc4ad953d130c8c5ac95a872c414f2bd817f77f6b0c5e35216138483f7341b98e6b17102a4b5b2a
z30957c60d23fcde4ab3f36f1b024c93c77565f082feaa3246248b84c2a8be9e4e4ca538d4da91d
ze9bf9e3a5ffc2b4d770c7e3e0c02c83df316851e2cd42a019e51ee21160c90ed65f4574a3d35bf
z5da63ef809892c80844ba1a8d09f312ac9ca1e47ad942cddc763d794f984365bd6c84f2f2ff7da
zf94282fb598764fb4ee1c61159e2426a9687bba77666ab7718400bcedee4162b85ccd08f75b91a
z2965b3c989dfe02752962f05a07f76323a5c516177345f42fe54387e185d188ef1bb25897f8fdb
z502c49ad396fba246a85eb3fdb1a49e972b11f74d9d55d09131f1d139b9a551286dec31b167ccd
ze34bd2c0687d331d6fbff0402cc8fdc3be286cf8377155bf96893ae8a4e284173feb26f0d13450
zb30abc1715bba6f9267dc74c72aa1123d3a396301b63e5a4c9b6544a17a6f77c6b994d0ad0539e
zee17db4adc028214ab15a2e514efb1a912a04c1bff89d158ac14381a4078e40f76c509606120df
z5a55b705068285a19d9e4916a0d6b869ebb00f19a6ccf1d4897a9dbf4486797294d9ca3c2c66b6
z84c30492e935e9899598976f8320e2cbd98fbb3a9b6dfd186ec62ed317a7fa1408982856841dc6
z9acf473a205528a5943aedd4df6956353855f29ab5a8aca86504c7b798d12b309caa11fe04d0bd
z03029b2d43498e8c973ffaaf9c6a6693924c1f910021cd06c8d6a2fab1106b908dc5a568528a8c
zfb2896a14b8919813bc1f46cb7d64f8adbf2d3bd90b001bd826de1ddc183eda0bb8bd6b5cd1e54
z2dceeee9cc5d508afa0f5d0dc4e710c8e3cebeed8e08d4b18591d609f5742f110eba00e3b18266
zf1e485e47f4dc0c0153f4d4c6c087c6da03b81d4d96aa64698b8b101fd33c9b18a57566646fe66
z2211d21f441c046c5864e4f41f5013c47440c74f5eddff7d4c3990f20277f262c7bf40939e08dd
z31cfd667e3099089998de0a07f0ab93f12a811ea59c401b604998b6a2d831f7b8b228f6f6e0fcb
zc458e8a7c8e4676ea6972da37d787da2e5e242800d28cd1613a2a6edbe26e72d57d9519342415c
z034fbf724549598fd0c08b31c9e870fdf805089c2bf94f1719d5b5ff0e9d063ebcf3fd8a355d62
z18215c4693511ba5c13450b7b58a2c5371c0460ca54757dde81ae0533f01a43325b5ff8d0c14f8
zb68caef8b94d53c6e650c7110b98eb1439cfa8ce81c2d654e074ebb030c0d0bbe8a59a095008b4
z1524f714c372be05623583593f7b2f0544135f43928d609cdbee62a383216ca4b79bc2100b65b3
z61d51b24a2865708225dd53f7cc298a6cfec2b49528f0500e6ae7166002be4d963955dd8ec094d
z0cbb0a90bfb421af68288ee6e9207d9cff446df6d305b7f0eff6f41142dc2602eae698ca2e23b1
z57f7902bdc87b528c4e54b8c815642c7ba899f13138d31c533c25d8de3b9a790d825c9befdcdf9
za616513aa9a44b99985e3d0ecb5a5d18f48385dad8e6ebfb15f0fcb16764fc5f5d6e32d261779e
z4e89a9d664cdf5a58463dbc6bdd4bcb270001fb25a2a280aa904ce1a56026dae0edda0fca25dbc
zee67b8239f26a42809c9f5723fc24a90cd01943fcb5f42f48dd2bd203ea1ad924759abad215539
z958e49b8180f10ad84da3e83b05fda106ad65177ce770c829d02610b6e5296e322a8c8cc5b4ac9
z7d5c3e37b59a255415de07f39b13a0fa05bcae5c043d272b5e08324c1be41b96afb2b7798625aa
zc191a63cbe6c5fa143118b506e49e8d7aa336cd1bfc5a1159726814f73af880471f3127b023269
z58c207a66cf78b80128576a36aff201d0327e2e2f948ec870f0582bcfb1c7d203172348b1e025a
z6cda5bc50a27b738865bd158d63f234f380ed5c1fc3c59966439e43a8a035f4e9462437bab1b42
zf9e0ddcca5d2c977433603464457c69b1380e004fa9e975a1c3d008758f57d4c0b35d796cc76bb
z16eabb3f5f54d8536e22e2f2f3975986d9592a754cca6dc6091b30639057b29b5a197a32ded837
za836e7c11bf42a3f5982b27b9a5975181b22abd1464f2ac63cd9e2d3bc6506aa338fec665e3baa
z0392f3d62026484f9b73d1074804798f10159673b44a61833c7dcb0c280dbbaa4d619a05b3f2a7
z90e0d2f85495c5bbb0cafafe7ccee759c27574517e9beb5fe2222ccafb93e1ac54b6403404b05d
z609dfdb1aa117fe4449b86a0938e3e2564f1a8fa14dcae3a6424ec0e06ab642044ebe6b2962bd1
z1eeaa2a0e1988e0e089817ea77c402b0bd1f370ee73332663801b907749192d8c1e3b378a65c3f
zea72d55f8b45ea19cc3c3d6240571baab1a330bdc00ef901bd504dfc58988e59ea198c435434d2
zda3e75c30ddf4363d076060c8c443f7d1adddfa1f755d0ea1cf3d2c20bee017d9dcdc3505f80b6
zd2606427a008a84442eae0d733c37db58a9ca79021f5ed69c21b158b134a14d209fb263731bd92
zaf61b04e67b7b6e47779e6729018528ddc9ed5dc6ee87527d293a5156f31e9fe4fe550e71257ac
zdf2287157754e22184479f16f17143139a85cb6ee92c3d0f23b2b8a4825fd1b82e235e8e97469a
z9466aecf0f7cb027ee0a1c5c37e4e36d01a5d5188ffadcf0ebcdc39d84aed5116c89c6f02a5ba0
z59df788b9e6afba97ba53e78949d29465ef514fc13a4ca8d836fce8cf647e9d9aa61c924f970d7
z7873f9dfe037e7bd8dabac7f7524f27c8d157b5738eb970fbc00893e88f8ab26fbb7c14a92f4f4
z9d2eac143b0f4768f824fe0de59ef6ac0b7ee5dfa00c0928784f247ef64abf2941a6ff1e0353e3
za28513d55053a1a72dec4041ca8a2a7de0efef3711095acefd049788b2efc7f29e716edbb4825a
z1f0987dbfeca0435ae0ee0a31c170bb112bf95f4e96bcc078e96522bc43de3ae253747647e1a8f
z25b80ee28428d037910b15c11f24e9527cb928befe717b14409ad70afef84fb409d79114f97f71
zeb51b8feee90d7a907263e049e3ee06e56710cd7714f4a697930a979f0bbb1a748865da4cd7b3f
z7df6f59605884d1a761e3d721e5df373b3029afbd7d051ffb017327c1688c7228bcecb07820a82
z496c377279e2507468604e56675a83f3ab5cbb048d2a719a74b6e280d91cc2f66417dce3332ec6
ze22f9b1146fdc730733156e0f72f680e2ff98f5849dcb0f18929b8f3013ef6f6857da55c8f5f65
z98a3dcf021bc35bdeaae7153f8913b3ceb24e888b924daa41bb667eda6f8e349318a69171075e9
za576c05158a15b6ca6dc3823dc1710f673eb5b191d30d4713d46cf7c2c9fcd501a65c317bdb2d4
z3eb59b9bec16e0310282f0abb9ea05e1ab99e2d3482e9fce6b8e8497e220e2b18af6683d7fe789
za0b011e191b0fc21554505421d9b29939b68fc881cf6a225f08ecd52a4451cc8079e3e7a115d47
z682eb95de4cfda03112c00009058d509e449c28505958733bb3c20089fcf5e68d2bb6e02a3710b
z8520609d2fd2b2954b0fb6727573ceb567f895bcdbfdd18296ea110c25411f93dfc3b9cce3cbfd
zc72b9b04665672cc0d933a6ec41085caa4c31bd96ce42477b08fca88cd7e0ea1d45ce9e710b296
z2a58c6bca626302d89ff0a8f409b7b9688a047c84d3c4373e2df5c7e09e610818a078e04df703c
z71f78e715937a65562d33c6d5733c7d33ae19fb9f141e33dc1d98280a579d3d36ba573c274002a
z2f2c0c323343c8c8c1a4d9c3ad76f4aa04c78a8842740df5e1c1897a2a22c9e11cf1941412bdb6
z953696fc8cf5d7127a2febc0deffe73242c349ba0532e2aa615cc1e4b09639b6d399df5c174cc4
zb18353857fcb0a6b7b94b96d85084dfd3526b5dfc186bea52ad82c5b6df99cb489e6422f925b95
z1b37d647002722c8ced1b30487769fa6d0a47e8687ba71a31ed2b10dcd1deb6626d91294026c8a
z3ed8ab20af027bc51f77b178cc415b33969cb4be6f5a6981cd2c63a280024382171d49c46f2549
z67edc868df7a528abe3f904347c4049629f36611a6b516752e1219465b14daab6981ae35920ce4
zaba1f812a2c342895f1bf3b37d4bf4ab5bdabb83e1d93ee776139f8823ef836ea77591ea23c569
z830e543b581c3d00dfe67fbe06fe1698d2b57fd7a401565d2deb9394d826a727256082f80c4585
z66de44b776bb100424a5109135c1e64a3ffbae039c449be455709e79815fea72a83020e2208011
z734cf790f2edb63a91616a567f776f0e756052543bdaa6622d80e6cece175b05a294bdb2d650f8
zdef77c8ccc6f5eca81e34adc909cb0f5675511f8faca7289c21157381bd21207fc68e3992006ca
ze1eebc23798ef6a9db757223dcfc49381950001361c262a95ca721b3968853dd138bcb56250fd4
z18482578f44acc9a0beb3a7490d8b94f1754c5523a5b6b8c98dfb5ba7bb9d4faefc84e2d2109fa
z7448a711a59375ed11ff4b2608658208eb5ed4600923f837bf31b28826ac1bec69a98b3beb2749
z77eb6ec6e9b407a84bb2db9b239fbb961cbeacc668e49ff2317a9f06c67eb4edb76df9a7576b89
z350d302510201fc597e39edb1f85880506b01f81c85cd447eff2485ae4d0d3ecf631cb2ff76d79
z0a291fe98cbcf66e4118b94e7dbb2cc496031296167f826af6317fbbf4403342bbd456d96cfbe7
z2d0a35fb2ac697e73c7598aea0e372d46a6bf4c175d7f36e8ea2d2ed20da72046affb2b848b386
za0c634512a811cb4bf63216ed677bb7dcffcb6068e54d50b386980e46b63f647f3df218f2f3d18
z8df8c11a2cf538deeb44d5a4f6f03eefc7fa902a3a98fd4b9e3528e6405f590862b794ccc7873c
z3c2974fa00551a55b58e3576eae22bebe0473df5e527b7bd005e37c0336aab409341ca47537e83
z20b66659689a30e5467dc7dacd2fbfb03df981843a88a7ccf0a1508889dd96cf182c1bca2e41ae
zcd9bf0f2ba6a8fb0c4706aaca02f477cc2206e99d4350ed3ab78c61b9323be0b9859d4b7db023e
zd62e7e723e0feb52346f5d490bc154972d4d6cbae81aad274889df77673e46d238d89a9a897591
z7ed3fa6fcb077e77ac7261ce6a5489a8abff47542a5020044ec1735343e135768007971d215ec9
zff903d782dcc34e9a80a80d2541378474fd19ebab6d1734105c746607a46c0132d6f7cb7ec6101
z4b82609495aa74543f806be3fd54017c08e96aa92a9d5fcbdf07b80bd2762c101e573a31739340
z85f55aee178c35a0ea81d03d0e03597a8ad716a438c6433ba2f40be2eb8a03ce1eda2791606196
z57c53b2cbc64e0ceb419aba1d916d949c9fd275683831b684ed1e8850b088b1cc6becf59c35d85
zab1996b6cece0a4eb07761905fab6b7fe03751c0a4294fc6f069d990ad6df7feac5a2a895ee351
z05faee81a5be801f7b2de2c4ab802db597843493654ee697710e8957dfeaeefa99c849aeda88ca
z245848df121033c2979c7206306d79c93048b79b9f94066b2e185428ad5c7a112f1774783adf23
z9fd2f47f02dcc72a23c8458f02a54c9c6c5f7378c279654b0cdb7492cc1c877ab262cda14409ea
zedc52f36ab53f53c36c64de668343d589b505e41f30f2c4439e8cbe34fe9d76f5deae0cbe14bf2
z89a4d55481e68ffa29f9376baf8214421ac4bc12eb51029a4257e3307881afd586f3dbd9c7feff
z5319e0f5bfd052c45f3102d3509b47f72e33c400a8bbef477a5aab9173efddce33fd9c8a38e74d
z1e8ebe8a8a136bab2c283b5a7e3dd13a823ee7e5ef1c45ba77af859d582f3968690dbe52641768
zaa2d4e809db355be6217e4758cfaccd7abd7eb53189bc3cfe487ae7edaf56c9c12f7ffda818e47
z0cccbc77da2cceffeacd50a162cd6023fcbc29114777d443436624b79a72f07e71b5dd30090fa9
zcf9b7167546c7aa7a63acecb3bfdc3b44c812c0cd2cd14229e350b48f35236f7396d8ce1ea0c8d
z202f4d8f20b5541a3e15f196051cddca7dce695f03ae2014f7efb6bde6d1e2d2269bf8f9703e70
z8c10459a938e750713f03cb5e239f8089707a924adf1ea1714701ef6737ee4e0a248c94c4aef61
zbafcb4d6eefc3f755ebf7f1a9751fd1a57a4018495999064454c7a6d25f8987abedb9dc44d17b4
zb71d890eefde2ec4dff7d5d2e5a2255ee0e087e840f4df320cc2559693ca54550d691a6a1f31e0
z7964c8f16f90ae7be7aaea1704da8a15fd0c477aef9d93778d88b34c5b42c396a180f5ddfe3e71
z1e6d32fd25b3a7ad97a15bc4eba07e13ec09fb1f263290337f016a4bf7a135ce1eabfc256ab86d
z6c6c2125b3dd6d29c4c54eef48b6c41094d5ff0bdcd0b30e13e1398c1102ca38a15d79685a07d9
z97fdb6fa183ab8fae221d4486aacbaa68fe9752237ef96edf83876c444d6948479ddc2c9e925ca
z695975f0196e947e21657c0313a627966ee447f1d4a6fcaa7fce292f9d4c51f4b673d66450a55d
z9e1bc43c3003abb24fcae2ce67c2b425613157d49c5683efc7e070442a540d2355c185fba6e02a
z8b915fc8b903cfa6ef5504dafaa7431c9d2256b65190e5c5d7f230730709dd3b3ae0e8b792685e
zf8d5c2fb6aa69e817890746d313e20712105ade095f55874871e613c38c7b493cbe5fbc41e0789
z45850e4d15f25d3edeaf0eb6db50bd2082f354ac2d171453b7b0f0f6dd8a669774ca7159447de0
ze445266fb7d88c12fd8c1287fe2e5ac51e54775b7e4da864b7a0e326c4f430af5ea04d2937a211
za92e375d55e2cde578cd6708a1d2ebe90b9957b5807dbcb1b7343948ff182a33670cc395a6d031
z2d4cdcc0127bc7a145c58e9932aa8c1849e7bb7620872275018a6b9f6f9253410bec51dc259d68
zdc6349c2899e0401ca8f86e5e4793be25a875dde0b45144ea3e98d6c319280e01bd23d48ac05be
zdcb287efbca8217561a8703018833a04d14ea909e095ccb4613060ecf2eb4b91c21a222c952b4d
z2437950ccefc6d474c5ded666e9807d156b6a08a2136084e53827d2537376955b31aec2fd5222b
z163ebef25ab8c67b1b2f9e6a0a99393c049140714c984a7d2562548a0261a37abeac0c890cbce0
z783ea0b13fef30a3043db1477dd96104a88e6d3e1fa47650dc6d058dff43de402ff5bb451d7466
z3b702df89bcbb48906a0fc9728310607eba1146684c1ba6b74f3b96723fffc63f876500045accc
z0e0473d583545ff92387ef8821126db1b2cf3ec3da54aeb318d3767e126cce1be4207fed4755c0
z5d0a1e65e123f79ecf3b5a311288de509a2180c05ab82d03dca76b4f43a37f113c6c799ebb26c5
zeb4a2c7b48f336807aa9df9bde9960ddc037f4d385db4f00cf5d499feba01aec06a9c6b0d101a3
zc2a9fbcddd99a11cde2f075fb6e12f75449389f6044b6f608ea3e1a1297e3026c2aa3cc32d51e2
z2442cd0f0a2be9b9f46bef81acab3f36cfa79a62f1d5cb3064d3dbea964689696c5599ad369fdc
zc514e549882261cf347d92f9364502c2bf513b8448f4730fc5c36fbb7f53ee826ea1a845bf95ae
ze868edc732a522706b9814d43d9f6e1c9e6a093f3891120b851f5437e1979c2d631d519ec76def
zfb68562129b89b527a12d2e293aebfd34abe5b37d163db254c5020770af7ce12eea4af2bb098fb
z317891c6d23517ec81da9cbffcd2e815bdb50e52e3a911632074332511bfb3771673c8b349cf3c
z5762c8e3f0d62f466f426e8669abd485b3c6aae79e010e810bdea6db604720906e4238fba82b57
z0f8ab298429c778d6db9233b4d6a331f020542cd44e3feb39129c2286889b78b54fab165dfb5f4
z02a0e1cbbabdf68a8f6c655145e44b35b657ccd5dae3e7dadddc8f4c7d5d5d2e3af0fb10410d74
z93f85c6dddf01b1673c70d72341fdd1d2ff51ca0176190af6ffef83e2a3cf1a92ac0e093e38e84
z2c099028b6dc9016c94be1046a49c27ebf0c3daf49f20abaa19576d0b62725fb2f0cdd508fb887
zb3f1345584c3ee55de59a82d9d50e5b066dc2cf361ebd7eb3a77419772945d0d010e67b864b8bf
z33d27dcde0249c7e15b383ce00d4d52c4c8e89d08de05fa24f73bb5fdf7a5eb1e5eaeece76b700
z37661b2709957bbad74ab1a4c1c7312e1d4316cb7c8ffe705a980902cd00b2e1e2312f24608b01
z12ebf49613b6152861eb2d2fa951468bafffdc9d991808c4f3cc613b57512f20a2e3cb6a7f9c72
zb4496ad89e48f92673a4bcf942b48979700b52b2e3a3d359706d344d5da7e61471f00182b2b84d
z65d68a55b0335fbf37c550e679d8ccd4eebfdfa4403888e481910c192ecbf5a90df9588f96e99f
z9ae17b111b9f7c0da5c902f62573096f8a735239e562ceb080829dca301d1aee4fdb8a8dc67fe6
z0830766b41150f4edeaedc7cfb1ea1be747b327894b8c56fd606cb3370107520d332c89686b0ea
zea886db89f8ceb175f8a177d3b72f6751eb7a7d3f18c5e23f2ad9728e2aab3286f2a5991ce7aac
z99a6dbe2b6bcc11a09af6dce4c951acc26fe79a0fdfb9bf8db7c1bf643e1c2a018ff354ef17c03
z3b5d7c9a1040710f3957538802dcd6d0266efd152e45a6421f7f6f56e714c115faf4b926f7470d
z969489240df68955ceb146a399816e5af2240a310357b9f3ed8612ecabf34f481422a4ef14b952
z594b680d03334d1bc3df95fa199beea91de6ae4ac7d3565aaafd6e77d9ff9d6e086d86e4c000d4
zed7d72801123e70d28f1a8f3305cf00aa0ce5168e5d39e243c3b479928344e2dadfe46f0d7257f
z08619a625941b149b6979df558b98191e91ca4b710859dad62fa996a248ac68dadca3cd8fe1ca6
z3a22346d5055dccfdb6f0de8214df87a1447d4a29c506d99d2bfe38c6abaaadcdf9cfa8ef68b96
zed69f78472963d9ab0d5efcca13b2ba0cbda00c7dd9c22df7689aed1b4586e22345fe866c2e12c
za059c2a3602a0bd052b75a9bd40370dd0168b383254c7640872097ca0ad7738ce9ad55758b1460
ze7571ddcad73fa61cb0825364b29ace811b82934e18f4bc2ce751ba7850ad6b623b69cedcdd504
z20f1daa7a593f318b92607b81d3c7ce13f3ccca75ef6bfb6484c49191a38910887f84f04fdbd47
z1929b7fb090ac6d43e7d81a5c053a654248fa2f661f0b31aeca664166f984fef4345f27d11e006
z7cec14f4bc8f19cbb6ddd24be9a3e55ba2ed68bd2d439030f348dbb12b02378d7c8c7c390d0565
z341274127b0baa5ad0ba19e8176186e0cb57cc36ad5c44296add907d9f8dd8285b09280c43848f
z573b8d3497201714be1bef6f749e6b7e5500c97344fc2332910a8163e4adfcfe2f2a3ec4b21416
z84507ca0e0d822206a02c0bdd297641d5281db58d42bf92a3a92ebac573357975fb84267d45c29
zd6da7599e6460bddcb2545a74e96948654bad8ebc38f83eb3fd85285bdd16850c7204b1f7c281b
z9b663ca94e698eee2590c3d564df42c90b115ab060f42e544523e03bba54dc11d15f8cbd4d1625
zbe2be15176dff0804f8c46e76056490039d97035dd15b9fd7d4698798f74583c2bfe0bcb52547c
zb66f3a4fc17f5d05c1cb4e91e53f08a43aa421a887f0ad978d79cd9c3a73d60fa7bc0a381f11d4
z1e082bf20354350713b5b4bb81d96230ed8e4252e32d014d2e82dfa4b55ce589eb1e8515688388
zb8766cf0fedd81ab648ed0763b05fb0caad508c0f2b2328c3576aa08a817c0e06c8ae3d4f0e9d0
z6e3243fc0e2252bf4ec058da5f65e08cdf3158e6de6bb6f642b14733be6de2226c7a20994c50ca
z9f4afc5fa1eb924a58101aa9dc1e3f3ac760784b69f477466f8d52b922d999349b9e82e9c1be75
z370222e78289b322b2259ff642ddb61413024319b5df57f92412d37f87f4849b8612ab05e805a5
zc196357e7af364d14abd095f2d3ada09a1fc53a6fe338996dad6eb9927c22b39e5f1dcd5f5be8f
zfb8cf7309919f7ac3222a662a3809f5d8f31d1d24500e4df685b0e9ae067a25fd6a91f94af469c
z654e70e585ef65459f833480de9bd7786c72a1381ba2e0dfb1e008b7fbbdbd446105586528d3e3
zc667ba06222ef577fb85005277e69d9e7582440c48bc99fd2c14baa365b7c9e661dda5acc8b814
z6e2e71cdf1e4b60ed11aa21d0f938dab821d04392afcef0422db121e565437a7eea1701ae8c12a
z39dc82e0a1ad8648de13cca009829ad781784832a5f2eedb4c863d822a067384b65b213431284e
z214c1ab409660e9d477b5343028ec4bdd9d00d119c889c69905378fd44d482228df983523b794e
z704e1af90eb8844ca8bbbcb8481d4c1b6170af50edbf1fd8ece4c19973c04d1faac7d67772fe4a
z83474267a4b84a80332ae3637b24e0e79e96c4da961adc426fb0c8dd2c7feda7aa5211219ca172
zc3063e5513a452350cf9fcd412c60836bd9635c5a7c8b635edf60e7ef6bc5a3a133ad0aaf2d563
za51a5cc53964477352a7a34fead01ddee4008021417db1523ad6972f76728f5d0270c77dba89ea
zffa65c0f8585cff04c88caca2a0e3b121642359c41290f3ccb779bf7eae777bdd6702a389ae9f9
z8f23587225de2fac287ed111d0de4aafd78d82fb283d0b619c1ac93f9c05c23f48e7138773d2af
z4d567d578b68ce4ee3d6517262165d3abf56f7c80490e0cc5db5d9bf0ea8f78af957b0b4a145f9
z310da5198d5a1e67fdfc5fb4ff4fb21ded08ffea938bfee1d0b01b87a803ed58d830b380799f4d
z5910b6bfa45af33f964f35537c8d3c8469b59664c0cbb0a7b867e5adf38db7208cb992de2176f2
z48dee4b389a512ed65859242bc97012e9535ec4601264a836fedf3caf57ac80a1cd46103ef1cf1
z545df8c14bdbe3e401e0abbd66327edcf9cba18ffe12a7ff58dd7de71047fd358e845991fca151
z0a2eb227667a8c1b142ab5710566cccc9889fe801500c03f675532cfb96baca521a3992c6ca511
z1102565d3870758401248ab51f3fd640ded9ab6694ed3302ecdf4a0577a7fc7794e1640a71f556
z353930c5cce5066b9e4e92dbab19b526ed8c3e90350b544ee502b0688ba373918d411722b13ca2
ze4c68a47f06f80cc9a89962b773d42ccdb2f155aca1fcfc61d6ffe5a41db7a5d5c80fe428b0283
z5aeb980f6f68c51dbf00feb6f557dc07ab58937844df23ef9ccb1e1d85dc52fec728e42b6d6d6e
z10db115ea1512dd38bed00a2f39f7ad6e3eeba7249041c1eae51eceee97d1324618e54775e9d57
z6d611a394c622da1a21eb251ed7b6b39e4ddf6bbada05a59ad5ebdefcebc6fac95d02da3a0173f
z3add9041a8ce76c05ebf5fc04cd7612b3c6b5854fbf914d9484d5bb3f14ac14b19a338b94fbc26
z322720d381c61b2271496b7222736beda4ae62cb9612d5a5d4d4513b9e23455208d02efb8bbdfd
z23cb85809a1a81a2ccc0a514cd119a43134201d7211ab155338ad187744a897650294dfeaa1916
zd5916c4617f7358bf9915de6e53347e97b99b2304ad28a0fa56170baee4782322025a33549eca1
z8ede7a578fb3afc573c474f2249a907fdbfaaf15198dc5f0c0aa610f64f4fd46c79d83cf5151c1
ze334e995b054b30b418cf708db05876706a1e8d812449ffcce826e6e47ea99bc47b511c76ecac3
zdcaa63d77120c68d312c17b0a15f1fb367d496aef53176a36d232ad54962e0286b62154f4340bf
zc1dfd4069b58edc7e4e389bc517a07472b68cdc7e208e761043e5c4096e4aed1177a61734f320c
za3a0668208fbddc6314755def195ff09133928edd80cafa2fd98bb56139381fdd4954e64b7dd0e
z4a6345475399f3346a9b148d6216672f9b15f846afbccb0bbe0a261ea07b9b739fd8bc9cfda631
zb0440306ab81cb2b4cbba5c833a105826fdd2a51d95b3ace90ad1ff4fdd0667cf3948a4633d9af
z0e47591c98a071416b18e40ecf9f901c7777878e31cf3a1d2ef4fc1d78c90d45b1e68376bf7ea6
z82257638e44b4669beb856baef8c33ae290221c64c4cdb437dcbb7984befd0d5076a80766d55a4
zfb39e3f5c424143bd6b998daf236c247890471059450347edc9178c2001ff6cb1d005880e3dd94
zd73253a754c24e92881d1f8056db919141408fe1dde5f0abd1728b5307b81f5d853047f6148edb
z1a7f0c59d862c0036ca174a538744061530f0c3a81b913f587792352d6e353045b2d791e8f6853
z08ad8ab36f8ed81f4f34b6a7099e5a6d7587c7dd24a88221cf1cbc1325c9063fe02b0becde8e84
z752c4402aed28a1f82043ebfd770a5e3a286f9d050ef5ef8646360c473e6899be51b64b927cc01
z7f96db302c7cf255cd47cb878cb84d44ab555c06f6ec64c585364251f744c33dd58d91299e6ac9
zb72fa4b8df8ec2ed2e25bd9479c88c814be7b203706ae50e51e7d31865f6ac8c6dc2ae61e85377
ze6959c97fae11d016880b29e5a8fd2dde75250231a6599e463f7d8330c81ed23d734e5c2aea90d
z368b0b64b072933f525d18fe6e41fd909a99007307d8e516ccd19d92f9d602aa670a192278a498
z82716faca854ee566c192cff4a90c92c38ea5ef8729fda962c224cdc40589ea3f46d218678af93
z8dc8c4df22ef43f917b80e08d2dc18092cfb4a11ed21fcd86fe83c01daf68f4f7c3d00e5a059ee
z164908f5e3bf37a0f8a3ee53617d12139618d38a8da8181e7456ac2d561823d881bbf0d9eb1f51
za603b017f76fe82da571e734c4bf7934e8f448c8d32228f00ed32ef0d81c6feb05544030702764
ze05812213938b4750271c8b132cdced220cc67f51072ddd4d35bf10163bfd0a98d2729698db8f2
z9d920cbba8f496e3d6afe79cfdb5be8069733933e0dc339c3516b610eda0d826518ec67a302bbd
z6a2d29e57aa4982d744ddff682a2737f8cf5fd049e20830fdf4b942560bf8a71472678f6758e67
zfc7a8e37dd5dcf6f9f0897fd30aa8c289e9e906ac6a107c6eaf5966af4de41413c3279fb08ff98
zdbe2d5708b7eedea269937a4dae1d6be600580189da44ccc2a8e594ddcbd67bb9ce3a843105dc2
zf0316fc6bfeb3aefc49142e8c81d8a838c4e92b0598a122236a017efdc420b68cbcfe661e08847
ze1917157a4603bfd474509defeb520e56350e048ebed5af18d65aa418a4adcecf6118ad8c955aa
zc2dbc51ec6eb84549aaa3455ea1f900db109e47bd64077503b0dc79a70d1058a0834f7ba36afa0
zd9d8816eb703931df6041b08cf36b9a5ca58c0f6bde98cc90cda67773fc97fa8ce5452fdab3f30
z529d6cb64e8788f60706bd6bda20eb95ef73a3b9371a5c0d925d73ef6f1c789b58b8d811fe37da
z6a4dd2843252855f9dc64f42477ced557abe95ef5fc8c810d4130589140375e704a3ed60e6815c
zb6a7f9186a9fe0480c37e128578c0cece200ced4cab6465ccdbdd0edbada531fbc0bf4640df040
z6fc6fa33c370eb3a90c9feaf82c59f28b5808ad3fb4cc5878d87cc6fe8dc2a3af3fea9048bdddf
z5daf37ab345d15ac2d406dc274b7058482dc4c579952567b291821b4fd1645506d5576742ff4a1
za87c6f8f628b89b14c828f17bf6e41327ac728a6d0361a11f628ccc9b74aaa752ec9779f2eea00
zbde582f879a77ae35a33545fba9599407dcf4bfeaa82b4bb2d2221394eab31272ac6eec9a5c9a8
z9e8a598c5bfa5adf62bbd8af54db9fdab914a3159dc5ef35886a1fe7eab39a8df629586e5b88d8
z3d38e95de56f298adf009336fc9810f49cd1bd578fb3ebbbf440d9a30a987cb4434879bf18a57b
za3a4d2e0389dce482b54652d6d49c355f21de8b14680d60b7857b96b4ac5eb0b6ba8965a1f3617
z2dd8300aa57ce8b88d5ee7aa349bc62b0bd503f84984cb551e1e6cf95c816652f18fa70e849459
z715acf4f76cba8a6c04b1479fcf015a38203cdcc6b50c5f81e6a69449c3277c9b1d5138c77f95a
zb44643813930b28559b6710c7ab72fb46aafd7f0ed309011e4208b395c3d33c5aec6b77a77b15c
z88f4fab8b1c9598e36a608d4791d2318cf0cddd7485cd43a47d7e54ea92eef2722b5dd37145c1c
z939ad2c0a3c3046b5f5dd5de3ae1ba56c49950ff27d3cce37ccbff852ec78c6509d1b13b07f7fc
zb844a5da15811a9624b22c49d79364f8c49ff16bbba3607718fbe50c9f2a922d820e24722a0a87
z7adc4881a06755aebb9a6c2b71ac39b79e78533d1f7c34132a91fce4370e1f6e9d0d872af59f06
z5ed5a4e112f2738c968817e51d201bd7a76ea454c2a0347d7a919e84a5db9126420c8b8d0ba3ee
z6752ceba039cfcfa297cf8709c91a7f38a2807d6cecc68f633f6c242a211a6f8b587bde54b9bb2
zae16c5b8fb6d25c860c4dc30fddda23b806a92ea8bb9542a5dab027978d97def7d96cac65a8939
z5191d0df4ab9930287f8b596ed87db85e5b9e1e278b2c60c2ffde51fa53a3f94359f24ca2e7c01
zd5d15d0aab8994df44068ce65e6ed44f4aee6c8f9be94eb122dbfb1fb6899d4e64b389bb97298c
z3d91026b04825dc3bcc3423d8a1f219650b1ec3ed03c2b0c8513dba33b1016aaa1156c48cefc2f
zad97882c54d3f3dc9bbefe9e80c3fac7d84d5e2995ed38634a07a53bf210260aa205b0cd192178
z25fdc921a3e7c938e63e641c45de1603519756c02b2a59fb81658946a9af97378b1a6b80e9c4c2
zb5a009d43d61e68d73a01c6b87e3fabb3cf126c33a676c48e83f5b4d15fb3d3706d535637d9285
zc32927f2a628ea45b55c8be5206f8332bfc2b3898a84087a5a043071aeac08553d904ebe0251ba
z82b90e4124e970dc7f4c5b2b82de7286b8660a388f81df3c3c94b2643c1ca15161b1d54fe70011
zb3886275eb8248f93b93677f4a7306852d1ec87ab5711852b43710f6dde53b0d9421b425a15563
z43cbcb8e6b8f11e35cfb1b07f44cf2291899341ff9f4a992f92e7d074d53e201938c99aa93d27a
zf350c26ca0d5b6edea6af7932cdee7a048a26e2f988c9aea3aedbb17c63da6e2431baaab4aa71b
zb65dd769797ea799e85be0eb8b17700aec19597e5851d0b7f4003ed1db4375c75a25811ea14ef2
z837cf69c0e426144c39f860f34f4d565c0c700c860c0ded1439c33933e7ed26ec12ff088ada632
ze26e655c725184a59e9a0e098dc42b007ba11dddcdfa5fcb2c1d5f575486de789b0108d9c7f89b
z52b5d80be7e953d6999cbc3399f2e47272ec19c8cff6b9e7a7a2ce01a62483a45f6942f31f1e1a
z92efb383187433916f72935336c6affce1386fe8653f72e86448ced3d5a692c9e1007834e54fa2
z67ec1538aa39b8cb772d90458a763acb7866e1d6c32321bcf74fbf3f18883dbd296336846cc541
z91f2d2464d0a892c7ae8933c27451f775cec2611843e9dba492e21663dc9b0144c18fb26bb3713
zc207f13f57a68c50b0e167630ef649b8325e008e0e52e78480cb9daa09a5cd1bb0d666b9afc297
z706bff796303962d970f9cfd6de09566a611deb50c0a058a6c8cad24f5fb6c94790953c06bb002
zca6913d2903b67e784dbe7401259ea6dc17eb3afe7e3d79ba79370f983abcc49e72325ca963841
z967dc622f84b4959f53e2004d70740234213cb4b48526d7a9f3c2a144d6d5c5e36724aec7a09fa
z1a355a9cb05ccfaab7f9289086e08beb17a680957f529bfe9c32f47ba3272e858d6d28e9714322
z79d4887af0894243ddacc9e8363b4446175c10ae9498297a04c022466b91b74fe2c81a79cd69ad
z057bbe9796b8fd6f6b9a1626264ff7bc77953098603b7260f4d79b2f12812eec6ca4eb94c241d1
z17ef3e2dd65de415193e8ffc8c750cf1ecedfd42a3724871fcee785c9d724d5bdb3ec1995c9b64
z9da339f0b4203a4f38a0a7d61053a385a991bd9a4479140a747a14c1a3379e08c53d30cd12517b
zac229e31251efdc6da6c10a36a98e6daa943bd605962d4a36cac7b7526a53796d8608878355a2a
z2375120fae447975df4e3e39d0f1aa189495579c8ecd0b311ec6324baa732d9544de49a2d83b72
zf2b8dff5a3910f5ebfa6315e74c791a21049c71d1b4d29b41ee8ec59ee6a546f5b13c386ae4cf9
z657972847c2703dd0f659ae974c802c56ac276aecd4e6a20884690089316261fca5f2177800f85
z835b0c6664bd7e863c82ebcbad5171609a9d13ff99f98a17e34eef452d01a0e7b92aab0f54961f
za269d17911cf035fccfec68d7155d659f705aa87085284adbb90417af7878baab648584a835d79
z0fd1ccf509317303304f089c52c92bf3718eb2e6af120ac5c15b12a6efaae67c18b9095f8a1543
z10783f446f0028b3c95e4219123ced37140807dde4f43f75426670ab7780eaaf2562e56734c8e0
z08fcb9569894ce8471afe79dcc0da26d2555c6760d716d901eeab5ae8ec94b70f3fbd5ff061cca
zfd5cc06692fa86867aaed053407d3a87ff776e89358fdfd51583744efced7284f7e8edd88a1d73
z9919e50de2ab0165a1170cca2da3c29c46b9ae709c972cec3433b70641cfed675a88b7225a4353
z620e005082e4245046542b9c2e15d2a8d36c790b430d16b908223941ce809dece6fc8da75cbce0
zfa7a8759886f5f07086556c738ba0c2940032f2021dc4042fcedcdcf608f877cae809703e6dd8a
zd28c3fb5e2c8639146ef5a8cfab129bd1b6a50b8020f606fb7ba27912ab4b4301427fcd20a13fe
zce777da2d2fc82c32a0d94f4f23da409c3c5a2e091da874fae749419fa09407387db82fc6e73d2
z4a9852247c85838aae83e6b08bba85c13ba5be226846e4da3509c89103bc4db505daef570f4221
z2b29a8bdc67a70764d2d654f38a699cd5d3ec7691187afab91137012515c53aba6caf92dfb4025
z181413d2c7eb2edfe4b159f48a6345a0375ed1419ce086e81c2df7e72dff1aa7ffd72f8752e452
z1dd86ca356e0b29c9b798d11478f4dc55b9bfea7d8aa7214412dbc5f62d6fb6843debb1c942b1a
z7d47cd06dadeed93d1840671a70525668940c300aca02db016e018c1e809e6f1116185a5ec29a8
zde52063403231df9328c54a369817a880e63cbcb5f4306877944569ee348ceb1d1b0e17492f693
zbd3f10c5bb504cd0dfaa9448faae2acb1998e2883dcdd176bed5faebc2789355ce30e36603b47d
z0bd2a399869234d5d6d5d46eb5720a634e548b5cc9c550abb5c2459c41e634cd8dcc0578f78840
zff3c33a7510ca5b42b304c9f33efc3f60b8c99b71ab7213b961d87efd8f70caff6cfaff015a3b1
zc5336b4ca7b0e847200c17f7139974aae52decf911a14a3a9cc39eccc7cf4b14ff1cb6b4ec66fa
z11719ca2ae6349f08613494eddfd4787507c1f63ae4d85e41372c3fd2ea6c5d0b229a32991da25
zbe0c3ab4d098c4a97c58b09bbb22c15aba202c4839aa4e88aa5a88c5e0789ba00f4e88554949b0
z336135158ecf48377938506275e481db644f4946b581deb104f54b1c88ced8631afa960791b34a
zb675193066a93f50fb6d2ce5f062f70279e1cfef4340f4c89851dc82a75be8857faef89532d885
z0259a308d35648fe5d92a60dd5876cdade74feae6bc6a881bb4b68768840b8df57d15b83090cc9
z92c439e9abf68e81f05c0897e6f458571a4327e597fdf40be3ad5b2f30da40db2b5774e9e46c77
z3c4971a066d258817143facbf35e917e47be2adf534febaf094a219b8014f7e24ef7353cd70e93
zbfe29ffec746795bdedbe520323d9a88f39c6f28f1e4469b2cc4de784cbc2acd1aa40039973165
zf5b99745d67c058a83c5b24e18f51ae7b86ffae3ecaf2c91ad8ce1ac9676d18c86603cfe50e9dc
z113b3adff6e1377bdf72c95948d715978fdeec2a691db3650e85072d01b06cc5ae55e2e4c12b78
z6c5ecb511cb43c88b90aa443e06b8ca8ca07e020a46af3baca32ecbd6ca053eebc9564f0f42c3a
zb51d6bb45c7098cb1e0df71c3865029b97f785ef63b180a7473232c5b2e52b3811f50d5cf22439
za3c4a1d0fc204c84a508f06af90da5002e7fe763c0d89b7f6977d040d747db6fbc434f13bbd9fd
zee6c08a2e3a719e7e93f2cc9e748cadca541e9ebcfb7cf5d2b567f9d2135f433355a00a1d5cc9f
z0bd1e19dd5cc0f9ec6a0cdb091da60b1562f33c6d1eba39cf13df9fdd9210b72a15e37dc5c4ab3
z70f677929bf017c64e0921330e3001545bf17e6cdf73fdc11d86534cec17470f300bc24cc5b7cb
z39d926e97d264e003c8f282e87480e4833b60a15b19a0ca06b87656977ee490246f560ec8b8492
zd5cad700162c9dbb40192e7cf319e9950fab2f7bd10bb0d7139767c25515ff343bd04edf3789dc
zddb64ffec18bcc6247329673b67666ac03b155433bba070d7bf50fec472f1cddc3028220723047
zd999438011428e7ddf70ecc17c0d0d5e49cb5517d96b05782d91af9d248e6f98f1121452e2f955
zf5fea7156fb835668d96449a641ed8a549a8efaf2ecf34405be5e8f14b4a072136a94429add29b
z48c7817dba69edec486678cfd98b9980271ebbff4e292b80358ecfc32e8cf2a9918b6ffa6565d1
zc3f7afc274f99cc2472d6c36963f3567acdb025456a1e5404792c903e6bf2e891fb3abaad084a4
zbc16d4cb78e829516a3cb42b5c6c1bad4d4b8ecc2e4859341ee7e2f9f748fe7c2e36dea9edaf4f
z3366ab92cc5d49cd325f9622fc39184f00c64f5dc6514e8d25471ccc381837a28fd46a7ea33b26
z62d80867874f6ab9a2b3487353b4e7dce86da609de6d18af4643fe13188e9194fcc216f82d6f7e
zdf1c639409d4a0d60695605b1912f7036328169194c0f8942a713b6d46a5339c0df5b346b7ce1b
zca46cc616f60b28298758cf7ca1ef897e27d003a84b49eb0911a752d4e7538d1e8a36df7f9500c
z7600c73cc8a440752bfdfd8f07d98f4e20a4b37e13ad5c0c04d476f3784dcf78e70a24da0298a2
z1255d7e768bac6031e6061792a4cae18d9e73c4869a0bc1dc6f374282d301d3305eac4b460c3ae
z4fd548017cbae35477299637d4aa4c0668732428a7c5f1055649e1f7da222ff533aaaba0927f98
z910bd6972aad107ef4c747ba8fb91557155a97ce8936a09a777c83f791d3c33f06f4f5d1db4757
z5d6fded0a0dac8575ffaee2bc7c35ea1991a541ac64d6d8e603101a91088dd47cbbb789be584cf
z9a1d12ea3d115cdf56848e00770f7fa96788f80d6dd6888ed3ba2faf2bec8b4eb76ce895387d7a
z6380c9ae33445918c084462cc0c79c0b845ada42eaf06a372411b6b849bc2d41155677e82f4dd5
z26dfae18e01ff99686e990774360318a9554f0be2d3bce7c197a1309b08503f6c9e0220247096b
zfbf2af214a66efdd83062c6e67d6c0e097e2c47d9d8f1e4c8f684302af62edf4a746730f5229ef
z7562046e3645191cd7d93a70598ba3772d02fb6d42b1d0f52c5f35f221f5345bd1da521bb52608
zdd15537e991d85df6bfe6952435e2e1eaef14623533210c38100f56a4f9ed16846a65186bb454b
zeb6bb4a7c23fbe503447d95f232d84a890efc924c4f8a0dad6c1ee4aae4fe7a8253598ffdb21d2
zf62ce94592ae324fa6ce11756f9146fc90042a406af32096e2f62f38c600e05ad00a0ca2b3748c
zbc7f434471fe21ded1cf300c7f3b8255214cf7cb543f2e79e245c09bd087ff17c6decc66ae04a0
zad43642b5423e6902431f8ab0de69a66d25824975a3279d27cb13245123f7d3b9a46bce09004a5
z8d286dac2b64ffb6d8758ac0904854872e78180ba007116d3fa9104f224fac38673dabe8243d32
zce0ada192ecb47aa274cfa355ff3b49eb6b9dafccc1e6a3a5946fc41d167c9c685c75207bf6ec2
z9b031ce81182b050dc61a12bb9254d8890c38f6d4aae72b07f431907a586dbac9f6ef83c4918c0
zab180aa255d64083e20c5c57a6605fe62489fbf80efa467ac346e9a421ec004187e448a5586bdd
z83b8d080aceae04db8705c832c099629d54c7c9b7cbbb0ba7ae39e061af5f191a8787f52f63af9
z405bddf6d761a5d2ca0ff788d1a229eff885d7672660d882af9fd1490fba868ccab03072ca0139
zae435851181c05c46d49d8d52aa57795f6d07b132a0d4cc783800a6ccb98d93814ec29237ab7b1
z55291e8f43dfce3b41dbe38ab65f4f6267c9758b9e6440c9cbf685235ba7ec0e89f591a43a217f
zb49722266ff5ea4698319802c6ed23c13ee6ee9fbddc16010b92e0db846e1acae573e4f4378f48
z0e552ddbdec51cb09d68056436f8832134b22bd041adab25f3ca3e7c2f52506ec40ef909c590cc
z7b9dba01b79112265647ab312377ef2f02c650067d55444dee59e8265049b100d43a51b9e1911d
z0036d93abde504500081af0d9590bd3884a3fed823534d3ce30464fd905dfe1d29b86820b1a4fc
zda504f201f7eeaa5ca2d1347aa3a0d1709f2c6312aef992a905518f55f2970a46161603f98f70e
zaa1649685d068bd95dc2349d6328d1aa54dc08987c0c6130e39c5303137cead01bfa770286d85b
z5488def9141f625212bddeecf0f7d30443724b43f7c22a93fedf9df4048044fc08445c4536d5fd
z15609b45b93b0031ef3a611f8b485ffd725a61ae7b7f1c040c63de6b00a6bc5300b6a4ea9394bb
z990c8fec9bc38127a796fcc9aa49d8dc47b8c87b15de04cd363e7a1c8b682bd9e663adba2be8c9
z88348bb2d5910e900235f8eb9f8ea3f216dc26977464eeab362ecd3526e77c736df40cab1bca89
z2a8fba044c438c53f06fab25efabc8bceb7370281df62812c027c15de2b2d2d742efe52b5ab6c2
zbf5bee8df8d500b076ec41cbf6b5a8c084832776e4bf6fe09ccaffb84db034d3bfbab17f24bb3a
z1f6edf32202a2c8faeb1a8517e3a6a8e4e9cbfcaf4d1f56dc42dbebc623a609c26a8dcfade98ee
za979b92a045f5fcb69617b79cf507a69af78ca1ddaef3260d8a37d02ec5ad41cdecbda029c0f32
za138a239f50679d3cdf685e0d25b059167426af277e8f843e052977077d4db95b35f9c24c6ba44
z115b55e47bf1ce892122d5c44738bf889d1bd77671fe454a109ca34d06b25f14a493c3267574ec
z3a59a1c8c78c0c02d428b1817ee87fac3f5f31a88de4cdc37160aae88859954e2d31038ce5321c
z29183840607262fe44b6fad7e41181a8a2e7a78d3598b7b859984f49a50909a55b8ddac41078c8
zced659ea26a96951565e6a1a76436cd766f21c9967b24ea051d4bd0609b8cf1c8a18d72d49b32f
z16899b8590170e1366c32aa737436e39d0911465eb961f352236c0322008c2915e51281aa0d71f
z45f82c21abaa2119da655c9de2079af24daa7ac9054e17270068af527b5f7aa83544439b28ce74
z1af36b2d46881af46ab4c9b4c62b8737bf184bff71e07342acb9cd4bf165f5f15d3da3c4ccf9ad
z7a97811efb1ba7ca6bd0a55a5d205e94dd18be9aea32d4fe9c3556258a12b4ac72edb0855c0e4d
zc80227cf77ee377b9ad8ee169174a81616e17ff579cf8e75f357be572396b9243c3583f32735f8
z4463f03a160ec7496092e40f9b28f17f79faabc46d92440c49040f94fad9ffe97db40a0805027d
z080f695a2155a49f9f637d10adaea5aa2b1985dfd01551f7b3f0bcf7e5c02065a3a5546e9373d2
z0046b17abd9344a1c3ca5b3058e2e48869c5cf00e27e265640838909d16471b0e9da3760738bda
z02acc4b6e8678ed3929fd6ac4573776e0edc5b6f9a50c6f4a1ac99280f82cbd2f1d5d73753ccd2
z505cef05080e035c0ae1b7306148140efb457d3f93b801f6a23004ed307550ba1230a9af2cc27e
z599973a9c37bbd24fecccafc3ed0cecac83b8fca310d759a53c4002ff854714dbdb9aeefb8844f
z9e7f2bf2c47ecb3f70547bf5098c9453adaea35322f3e9f57a991dfe1b032530996e789cd65ee0
z106f9c6adea4918db0478149ad42df2476ddca6094d19a3211e05f35af0b25744972c203d57b08
z2385fe8c94920ddaad863b137190235f2afc2d7b54dac0f124a5c0ba1c1b442f121319e35f0052
z0da6a419b42dce80bdcaa33dd038f925369b42f1f4e8d16ec3558ba81e85aab1428d36104bdff1
z6ade5a50f6b105934a3222a8e55f271f07664155c417c3b82377428b8130727bfc7cd2e77d927f
za7c3e373b98c1268b7d038551e7bedba4a5a7ef6e83330d3acc0c9469f6afbb756d07b90bcc83f
zea6f2ede8df0ed5238bff77e85f2c00164da474ed2ac661cf17c3eeb04b4e6d0d9676182cd40bd
zcf3ef015a595f599fa6b6208a6d0a8fa0ec899288c12bddef0a35634a993a51a0b410d24e56783
z7bce682b98abc064bfa607a4f08a36c7753f265689cbe8463ed02f48ad11aa1b7a989b24e743ca
za03b0583d311acb4d8ff8465ad8447963f9786b6825366f7712731b6525064e97b42313355caec
za0ce61c75d3cb6fef3f7508eb380e8d297c918032f9ada8968059cfa145471dbaee777e58d0954
z53543fe5f519420827d79e830f8ee8cdd74222d6f5ab4e43b8e0c50631bfe4ed6abb995611ee41
zf0a5e4d0cc96ad12c535ce913942da2d2cf1be917313de3faa16efcb00b0c2d520b629dddeec5a
z52ff66a5ad79ac963d618d524fcff42015184875c918e5977d2475f9f19ad022152d0e634968a4
z637b090cbbe5b7019ad5440f759c2f9e817554dfee83014991e89628a0e0ed7620397ef0c0ab0c
z2bd7e6cdf4b9c8b1f883a4cfcaa644ac829f1dfd25fdeec68db114e57269c1823864336dfe2985
zc3a4aa17ebf76a8b31166363add87087df876e365054319117fe668e045219e1ae7f1baa5b2a7e
zccb92c7da0971ed79a1e80ee0f70cfae037631b8667487c77c623474aee0f8a9f18e68fb235db6
z1b363dfb47021dd4a00cca0fbbae81c62b3782d0a48e79b2f754813a33d592a5b1d8e36cba383d
zbd923f432ff7a4bbdc652fc4931c45939ca91e0b8d137284091a2770f19422367b8b67d4af33bf
zbeb823761d0489a3e8aca65c6a78ff4bf6de5cc153f7c3515ddd94d880567521e1211dc34ced0f
z6ab6a635e6c66850c974a9743da550503e0ccc3a5be952a31562f02cefbbe0541ca798cf34dc57
z650de2bc94477fc183eea59d68226cfc88d5fe43fc8c89a75d266e0f392bee64501df897119dfb
z8b0e865aa00727a4fa545290220b263caf80112158b5a60311707f58d8fcaa1a3a0278eac37350
zcd1fd451d16bce0af7b838b5ef5bfc695746b59256a79ae6cca0ce3277b66875db0a0391631086
zee295142e90067709ad748e3a4433d4af7613fad544014994453d1b803259816011c508c397efe
zbc569619a527125079935933bbe1fe4f71f90701064248c88ba0214f694f9247512dbb5129dd96
z2908ab048a9e5dbee4bc843cb436768961d6a03743d0326b8a65592e88b99993d7de9287a016d6
zfe18ba3836200fbd7ee80cd67c2d9518915d66597d6ed9a114a36c58e7a7e13f3826915c3e0bb8
z7d293fed59a8fc51ae1ee07c2d54a6896adc280dc79153a833a7900147954caef623a12be249c4
za133a071c857103009726d33e1cf46f89505dee554698fe4d06533ff2010d9171d25feb99003f4
z755627581b820d5d8c25b6c6bab1baeb4090d12dff1aecba125227386167ad7f53b0ea32aaf729
z1b56673f8fb025899752af5a7e1f6f2345543ab191f91fc6b2a9ed965dfaa09423ef16610a007f
ze2c840b4d3a673e64724e53abe245b58cd42c406fa4973e884339566751ec48c51c89ff4aeb9e4
z7c71e45e39ae5f57eeaa5680aa883b50ac6c5557efe6e90322ab34220aee28c180dd58fcee19ae
ze09b2451bd263368cf561dd250ace66240b23af4f04ec4b5fd18966cbc45415ab10254a7f36262
z66d89feaa726157286f2bf0d4dd2d6b1aa487da53833c7bbbaa136b928cc251021757f0ff5d93b
z13c0eddd06acfb509c9559e0a125e77b185f79cfcd6a21d962ff5d1b6389ad42e6689485d67f1e
z3ddf76c642c97bcef2c13f2b0a11e475d9e5e876276cd4ef8faeb42ab3e82198bb6ae6244d55a8
zebbe51433cd642b75e1b91c282631128c3118d38be67d5e99d3ac85e1eaf39971a2d14b942f660
z5c7ef1424c0888249f546c8204f4bec9bb32fae47d57615eeb56f0af356955c0a4c8fa64d7d62f
z18959d78e35a1ac973535154bd4248824e8f834c317bc17cad6f3217f11a5530f2ec25c58372f4
za65d9acdd73119a3c4f6b6428ea9bfb4129e905606c42f4326de5df5d2ba56713db6c2e915a0da
z4c0776b1f1405d26513e4bf8d771894f9bb8e47dbc93d45241f8c6e1ac582e375baa524f5f85b7
z9eb388b626d83d4c79c4ff0578fd3fcdf036cc136670652c04034c6f7519e458ed45c615554ebb
z704f771edbcb83327b14055450029eeee849fda3961f7f2a4bedccb14422c510683d389e86ea40
z7bc8aaec28e85d8fe8cb76eaeb04de6b3c4d07f339c3d12deaf1859ce454db40e362207e1e1093
z88d733d51b7524b85f4d5f8252462558dd3f036d5e90f38a7e529f90619a03874c854968f436d3
z353e72db2a86a07a21d3b38f64c150628b41e4cb2ada355720face4e098d762d3e523741176ed1
z9362c12640111c3cd43f25441a0b497684585c8326e0e8c12ddeb77b015625b9c423f8d50ec3e3
zbc1b37caf9772d6e4741ef7b31367d684b6626b695b804337e911fd22672ca1bebbdaa6cff9403
zf741573f0137f94c3d947bef12272a2d3310e5a77c507d04d4e6d5308d5bd8c8652fcf6a9db058
zacb9490cb15e7bf2b3fef40f16d28efd5adf8d38bf45f9e5b70b5609f05a593fcb4481c422be6e
z1c25959d4dcbd651d95ad3925ef828161066114e94b88823546e5f83e7a37ed7ffef8b7173612a
zaf4440017c89958b15bfca9701548ab45c3d8a8976e62f89950194a56121f93f04313dfb0ff694
z39f0f03ab117849d1bc746f864688fb1016da3a469663fc8e9ac871516bd3e6e14bb5813b59018
zfdaa2e0db7f6b002969929b3e27b088f0702efe7920c9b76a3ea73d1f0026bb5c24af1aa6283e3
ze5d75b3ae3ba8d8e1812ddb7c00b9c458e75b39a74df15480321c8fd62bad9422cbff210e1a3e8
z54267940b65ba76ce2ff167c602233075c31957e3c0a9a3d13db17ad96be4ea3f428b36d7a25cd
z7159901626dfed8570d207163964a03a2bca91b48dc551f27aafe8572a434a879a972b406ad9d7
z9a19c2acaa0fdcbae600ae603cd1c19ce1006b9a8d8b2a7f8bb29234ecb350f9216cd3507c979a
z3d7982c92dc3735000e7de1605dd720b2e4658efef7d14ef3335894bbebad5e896054b92bc418e
z6998c12bdb3552d226040703dc7f5dc191c8dde4563a10550d3aa3ffda0c7b30fbad68d43a632d
z1f0edaf756b3d357842fe9a63dbb17c49563419872f688b6c4ad157c1330ab1f57cf8a3d1eb91c
z76f560d48118dcd7d1cae51310a4fc19f52ecff9638d233e9b967883327734fccc26db65c1b82f
z032f4ce7557659b05eaff45c57364f7f325266f9cea8dd701bd2d11e6665c379e37c751f5c743c
z7e6704efcd68962ca2d81fc3dcb956aedae61ba078e78783e0f800b6a31f359012b0eb1b9bc65c
z212b4b74be3e56204e38ac57ec662e578bc23c08a7daa1604041e26f80fdcbbb6792b5eabd38c3
za510c1b205e3f6aabee4935b0241cf0617fe9e47f5d92c03ea7eb19a6a7099db405cc33898e001
zec89699133c71228f175ab75083d08ccf2e28803e3274f5a8d5a400d17876b2194c488bf1bdbcf
z389bfd7ae164cb9c779c21cfa5b34b41d63577cb0b87cbb9b95643056fe06c4073ff6def88d005
z258479f525fbdac21889c3f97354814a57822865445fd0f6b19b38c5ee9582e752ea2ac6595f13
z96e205605b2b0de1d24e7c0b6d9af3502e80978a11df7528ce97236e29dfc3bf9524e518c64b16
ze677882329b27a5985c300e467a6a484c7c0f6c47be58b955feb05a6c848a39cd0a3f522184a3b
z5d8bd7e5d6881ab45ad7ae79a87476405fa0ed14701d036779aaf13e3fd51e5949629c0a1427ce
z8084c168189ca7e743c56d0ebc520c827b5ba2f7961dd03db472ea191c9d0d983882b4209449d2
zb428e6ae18a3a1e7d40328cbe881e124014eb5fc4019df5bbe46fcff3c303352f6a42b5661198f
z3778d76685a592356967811fde3310c1f5e91b2814105894c4f2f9ece290e7c484d835bcd5c58e
z2ca3c78ef982c132ed71e803908e5355ed28dfe0b83875d2b8db562c536ae59eebe6dae26f7bfb
z7311045e032463bf03fe42baaa7c2646d42b4b5054cbb92e65d72e8314a99c76bc86a412297fd5
z7a34c087f896bcebc53b357f7be0c3a8cd14ec7565c78133328a6bdc635552c82a7112748c19a6
z7f9c651438efab681d7a0e6ff2621399f481e7389abf16458731161a1f4c7f35024ffaf918ed57
z7dd1b1a86052ee645e1ae6c01c82ca77cf1d5539ed599adbdda15d563b95b90b75ccbf9a698153
zf5a9239053361f1273d41109a80e15a47193208c4a651ee8a0aa35423bc72ed88e396033317f94
z35df06ccee2cc190ed2f23ae5afa1b8dbe2f39445abaeb49d5f5d1c239514befaf9d066ae456bb
z8c033d08e1fde98f34b7a87d5c509b6842516e557cdf2cca0845076999ae2fba4f28f81ffef580
zf1dcaad0da921c759af9d3e04349fd083f2c29d6f20af9e2273f6360fbd61c57f517f29e9ca598
z90c2e0fb28329bf9a4433215c9486d0bfddaa80daaee65eb0924e2a166d9fe71f186a2e9e2c30e
z83959de64d38ac9d99db2e0ed3966cad372ca3067f21dde73206a04a7f7a2353592ac22b19fa8d
z0b240939e717d05dd6f30714e518cffec6c8ae80f86ffad6cf90ee455d67ac8c8d7af53df27047
z0eec83668610604c57f5be0a7c9d62fdf4790f3944747544a654f28b7bc22e0d895ae1cab6832a
z432c69c679cd5dad0227a82c4f571c26c0300417ac1f8e10be99cb5339429d6b06b10f2d8da39d
zcde3b6d66edd7e6e7073ae0360f4e35e107394171c2c8a114ce93bf34d25828b80d7784e9bbf55
zc76a1f5ded5a0325b18546f1d8d9261e8d77b098b7bf95b80005dcbe5f5ef352b3da265dc6ec47
z78c88211e655a578571ded34ee06dbfe36de6dc98df3636478e44cb5da39dd384b9b4fbd57b153
zd268b687a6b958d021ce1c62a9f2e7761b85e0674dea0fcd1f10d938e46d58c031ad437fa495d2
z5dd582452b634a21158080755692c323e1e390f32ce5b2c6ac63627973a14c7c2c0c5ceee30bf5
z80182ad3849b980d77236d77b32dc8f9c4b46a298b33f7e26b5f3c853362b0bc4de468b6678502
z5101841bcd599e2d7d9f5bf7a2a64f0c959b64247f5dc30fe2cd3ae89f706e74d293de214da947
z9b8748cd2a77e0f0c0d174e47f3fdfa7718a5b8ba6631f4f3370558b7b7ba1e430ee66ca6708f5
z04b73a59895b9e901414a5844b30b18752e0b9685f555d5ba97a039fb260a18827d3529b98c3bb
z648be62276fdb9e157bf0e49d93f5f3a0b047867b2f041d2e47bae795526e6d00b15c0d5f47cee
z561c5d626f7f6d4a57ccf8f5e2c8559a80bd4f939b81865f2d9df06283135007eed468a46a8f0d
z010499b741440decf80f0d92e850d2dab8af5204c5e520679a9c44771b5b8b5e4dec5756c8ca96
z6b34e7b9972fc27013d3683c036e84e1faac8dd3f8c9022e983a4766cef9f6511502d4ae88982c
zeefb6fda001379010143e51c9abf3141d8201827f5a1331dab4f351c06f05c7012261b3cfa408c
zc42c2ea6a0ed8269dc3c1ef8c24f29bba770f4e128a89122747187c721d88f951c342d605d79ed
z31e8b4cc71c81bdc7d964b21c1511822affc24f874558d3c06f4f3948ff0eab60085a63c1dfc34
z27c57912d3169f88308bf8e5bac6c34d0c1016c5ba4dc158872ab0c00668384efafc3754055fe8
z24d7a27445cd5484a81bac4c570d21e0d0c535024efbece9fbfa39868c93ed63ad791cf0959ce9
z55271be2ee1d934bdadb5adfd841b490fad96de082158ba115ba4e53c0b09e23b3f84f0b84ac33
z8e8879ba9bc17e5ea0f6853866a64d6f1562cbfba51632b9d83e0e1bd08381a20e1ad5b64b48d3
z0a6679176c01e4ba6594c99dfab9d161815584f488ff9aff8a9ce438fee5d6d3d7fb5d546c6ddc
zf7617ba12f2d3513c5a50b9af67d3c40ea3ab0a65d226b3bf6cc88cf6a59f86b65b429ebc3654b
zd5bbe06f4955ef9b9c2aad24f54192778c991b57f34172cfe61117d89eb196b8a9b69b98fbcc9e
zb0a03dffb32dc50b307622f918515f32a36c97fbbe5c8a86632271aaa9cc8adf0ced252c32b53c
z5124a56098aab9d09c204d16c17f4fb491fb5017a13aa992eed93e4a6021e0e942d32904f66b01
z8ca577f7f9f021251c8d254e2e532a027eb81f3c52518d0e9b6b3956e6d3fac12d3a9899089a18
zccb34cfe5b5c53eebc3f64226c990417fdf39421328d70b3f2fdecfebb1f8eed9da0b8d225ba79
z9e4d346937128b7b869093555dc37a3a6a08d78b4c7c162f1719d164046e583e0fd205d1465983
z3cad3a50670a8c7e510551d427ed081ff9b0086c4729165073656cc00d3fc5ac9545d84b68fa46
zf2f3b3324d84815458aec643dfd0ab3c940348acab46972bcc3f18d350e91a4008e2a00640b819
z117bb48fdfb7f1dd33a3a949e2827c840dd2cebf8f7eefafffceccc52e74b10085bec66dd32472
z2584b55139074758161a033e1fd87454a63ce751cd04e768d48dc7c15c6174410eec0fe915f682
zccfd177901f20730bb3f8b518c1c84fde8ebcbf35c757e3c80b0c31390733828d3b712d747d50b
zf0ae2bab495121cb3f678911a33d6008fbaa41f8c91b0dae9d276aca2db24ef65e8e981d5828ef
z9ec4e8ad80048fc809db503470f85e75e1d4147e190946e9ccbb58cb9145c869cdd47860fe2641
z9a8ec58ddb8f0b8bd022eed8c5a0f03fb162f756fde071fd2a9519bb7f21f3ab776576c0a6186c
zbbc860209ddce7e1e6042ba5c3e0db6e739922775a9e3748cfb4c61fda2118076d47dca9c58588
za4b032ef936aa293bf366c873eff53105b8f4c6db0db5f0396088c266428d970942f08613183ac
z1e32a80abddcec7cb166a73ff881b3e935a21d723a119effc811f17e061515ba6bc0987d13509a
z49e4a1c13864d27210e1a34b3898d90146fbca9546c217b93ffb379bc71c4e3178e8ee65ddd66a
z71a5dbe78ab284d2e41f2c0168b4114f7a63fe291efecfc6715e10c1a5d8c25e565ea43442b586
zd45aa2581e18ddae848a84a96497f9dab0203bd51a2d6ac474d71a2a982b6b0a5eae6baefd67cd
z5a31f08e115806b655b86366d7a0e9037d556e54dd0513c19bed571fc6c3740ce39660769909b2
z66cb7137111adbc021d2229383e2cbc46af5cd35ad3196587c16b5cba3fcf9a2ca03369fd19798
z44c03bbe44803eca0d0b6576b56bbc3eac21b51391f6d128be0ca783995138c7410a0f8ee61c45
z64f54cb3c7f1880561b409ccc3253188659ab03c76e6ad7b70fe8dbce60748eafa9bb45c8017eb
zb25b819fa1321ab5a3ccfb999bb47b9a03af9c2bb1d5380f033fe28a3cb1e5cfe8a0b2c67808bf
zea5ffe703e407de0b7af0d4d48137ccd979577e64605ad317b8c0366570c2a7f4817dc004451cb
zabd50fa66879de8922b56445efb8b81aae3d874c28ecaab25edb3e7cc2f39c19bcaa902d67e132
z97d25c8fb36326f09885d47ab7c8d90d07ccea4e7719ae956cae33d1f32bd31f65c0d5b0121cd1
z9b514ba209470d3f1acb70c8be9666c4e919239505aee22eb21b8f29840a941b9a63622474efd2
zce0193ce52df80e837d3c0a2e892e53ef9588725201848778b83e9c89d773da75942a3b0dbe03d
zb8e29c1c0b1feb407c9c42b44bbb99d7d0486784ba6bf818b9ba43406b3b0abb13ba4b37aa162d
zb97bf0d375a38ed072ebdc6e349de1c35480f6950f7422769c40fd78b1d57eded7c51e17626b21
zac7ec1ccbcc28470e54a98eecdbe23b8df50d17c973f51ccf31771b16778ce2155ece574d32bba
z977fec1d20d7dcf826b8a768d4f9c64f76f00919e157051d35da5bca9a52b665e628222e049f1d
ze274bc0419cb197fa2f1f5d27adf7dc2b12b4dbe195b368ddf73a86183adc898f34dd3eaf1ae96
z42f9c362e71c6ba56224d3d07ef8dcdbfc1e367c058c14c3c4200dd5059f01104379819e9eb1cf
zd33a199b7d918f3a34338a6a1a35de760a88e90fe4c53c0bd83fc946ac8527f18ded22308b4e4d
z89458cd9e8db04831ab84cf380316cfa8f1dfb300149b1a9ea74c5e13fe26448a73e37e21ce4f0
z99d9e4dd04cd700665cdfc534d4a40d1aa6521bc85cad8a31c385c16c77b987e42d659302850e5
z5b94050aecd24b36465da41d3aed69a1324839e8cdd21b3dce78cc983851525f0167077e614e64
za84fe2b5b6c790141b8b3d859216c9b1838e5b8c520e384094d483eb4e3953a0377d1f9f0da2d7
z996d48f6efab19d6543825d6ee231328dd591dc7e55c58f8e0bf0140a8f676d5f6d955459efb1e
z85fdee59cb444418a522b96b47207dfc6d2338c1e96c87a4bb384264750d0b6b4491c9c48f4a9a
z8e0511e08bd31537faefa3b80b17e6fe5dde0796ea455ec4084eeac6a8c5b9286856d571277aa2
z0f54639c27f49ccc1f7e098faf3a4ab0d48ab35cde5be91d4f9a13a3f03efb683c420ba991ba4c
z274ed5b55e61f1a1ca1dbd1a735ea610d4430c2b75651c826d6fc6a31cb291c88d0405f26b9c5c
z77e92acc656ddcac8ed8c34a30227a8bd100fa7bf3ea1890cc210fe20b4094df77a212868641dc
z2bdf0646f0fb9b28dfb7fde7ea542053f1ca0bc7cb29aad5d40027e19376e8649b605a1959361b
z677bba0101bd800af79c84deb641202a80b0cece64df78d1fd7a9b461b5609979528f1431b4cb7
za1b60368d4145f12fe147a4283f27e4eb49ad97a473caca360ac31c58ce26acd2257bedd3d4972
z8a746cef476d6e29f58b04bf52724af2de05bbefa6ef4db7cbbd96662bf6df1a75ad3ee072e1d8
z3d97c4d403799a1e0b4fdb987629a5f2fc187d3d8bf7086cb2c6156ff5201a6a9184ee10a2ff69
z4039076d5d205679353e6897a00e26dff472ef913297884baf7c866f8a255754b183725a148931
za04be72bb6b27a353bd0b082e199e49690052dff5cb805f3fa8918bb63215018b6d6f9d7909f0a
za94ce8fe6acf1ebba80a09ee6cbaebb13cce38bb5a42fdca9c75aaa64fff0d6c2fadb7dbbf5f7e
zbabccb83781580d047f1e948e8bec293b5be8250df64b54ce58c32e75fa79b7a20b1058ebc2f88
z15c16986b37f92d43db15160ee7faf0ec1a3c4626f5ffe35fe4bf844383353c4e2f1d509b28aef
z3cbb6c125031dc7e9cf5495c48434f4dfa4058aa131453b096eea496a0c7ef1885e0cd4ab339b7
ze975ef1d4dfa99fd937e84cbfaf5de1e082e625dbc2101b05639e6d82df30a7bccf01edf342ae3
zae70c391962633ba90fdee289913f72caf06fa0e121cc668622bde7d13e646bd218950e87d74a1
z47d6036f73e292be22dbd062cf4015fe5cfedc2896ea66a435ff9e9033e86664376178e050b2b0
z65bf58037d025148bc8f8f6649e28bbf9912e329420ee3f1d6201c8ba0f27eec275edcfc42adc3
zb5c498683357522b55c34aac455d3d41e7d84c2fbd49695430a7c8fde6d379dfb3a5bc025d345e
z1a950576d2898eb1349a3047547aacb5a0e8e64569df27e50ef5da7e0e93d7e9c18fd596b22da3
zf0d45a44eb58ecd35aebf23e0b05778732a1a1a6ec6f781835545905cee0f1bab518eb67ca82f8
z2239051675b23d030e7d2f5f9214f5f37b6fe74b85b8f76586aa451dd8e02088d562620b3385b6
zd5a068075ddcd0531e1d5fababc6c6d47c2ebcbc17f3ee8925773c5c468157b556687af31261aa
z2e485f0b20bf8798dcd5897fb1142180a4710db4bfd8ad4a311c72acce69861f8bf68638e0102e
zacdcdf39c9015e0c7ceb0bb1fb4140abfd1485b1f8c93be972b6f96f64977f849ce038fc6b4220
z18f2fdaf62253275a5f06d521adcf0ca4331368bdf4a8b301396e4acf2a6c5a154e272d3968ad6
z24fa3ffa1960e89b31eb591ac2d7c4092b3bd1fca509aad738e024bec4625c0587be57a66cdcab
z44644e27e95944ec8d3bc392c75321a6035e70edec724c0a46dd5280044668e9d5368ec8326a9f
z6b2197cf4b48be5b6b91d2bb0398cca52f6f046c4bc782d5f331f07374da2d610e68a8bd6df006
z1e51f977af3add9ee042a035bda735b7a6bb43b3eef6c76abd0a302425c7400f9fe5223df5f5c4
z96d8c22cc7e64c4b71be41083c3422df1925757aaaf73167ed85a57906aa890957fb476f886609
z53e2e9a4448c2902581e21c7c18d2d8bd9f23346715a12c370ba70a2b51b2eaf9a78364aee5809
z3ac5f1cde5a92c1b955763eea6ce5d987f5e4c8ebb9fac3974c6d2aa2a07912eb2bf9063b83e85
z90cd880c09231eb0ef012859a922bddc3e807ebcd6a8aa00ebb755a3dc13c1a571c42e5e4050df
z88c0093f9ea64cba88c33a27a12be98c09202d19818878d02d4a79fe9590594f49825575b8f494
ze8839e3925f03208994fbcf866140ff9af020e10161e2370002846ed7898dc032f53cdae2a24c4
z688ab757a124df8db7935f3a463edff16b31b2e0db3cb084faf1e96c6cbaefc0b60f45d8512e80
z9d6c5394df7014c7dc5c74eac5c0ec0b0829c183dead5bd08b97bafaec7a02727e4a78e94bd70d
zf5808bdc4e05b4605aad77a99ac0aaee4eec682eca1a086974292fd2e08fe3e7998783a8ebbf15
zb4f6334d7ded9f5a696074f511220df5f42b8fc844726b65956e4f3bb437e9dbe5bc6cc024f7f4
z640083cc97c522e3e2bca551b79bf5d325c2f1a1dd8e1f57026c3f92da5a02143d252f93e5926d
z13b3432cc2799decae3a8b7b148decaaf849b6705e561fd9e51a6a1a2d97a5c1a579ae5ee5f2b6
za147c59df08b903d04347c17fd63a08753fcf898f34172499522d41418c8133775c81c50f04307
z85d724b67bde79f9987a7ed5dcaac890ec3b3162c03ac2468674a9f1465ac32af9c3d93dd8f0b6
z596063fba3c862de6e52b3f143872d004212be934b51955661314a04035d834c96284bf52a767c
z57159c4d2a7673f7cf57a59aba636453f469090ef7004a3e66eb59c9c0b225931d73d7ad029c2e
z883c2f0925db67441e83bb12bb2325abc89c94345a5f012ab0c1409b848859db4e314170de4639
ze65debec54892f35163243051ebaf98fd3833ca684a4493688eadaf1655dfaa32ddedb51ef1ecf
z470d5f09772af0243d22b384554892d09ca003c4ceaf14f077d96bfa9b132971ee62108f3ac59d
z1996bf3630ed3d5cbb587dd2a311e03d91013bb1e3845cc36dac8605829bc1e475b24cd4a304b7
z5738573c59292f6c00e76b623de887144491b53ffeff7901f8ef5d53739cc18413726a8a3cf911
zfafcb092f0ed0e4716150909a328164cbb4b4772f6c17acdc3bd76133219c3929f9c5b4b0fa9dd
z47eb84f52106253ff78f552b0d49735d962458d7f04a2c2e4089814ea5a4d2fb497209698301c2
zc0ad523abea09749c1e915ba03ef2da6ac82b77094b92646fe5c55fa2013056370484a3a679817
zeb767c0f77763741e70400a2b4410ddf059ad4357db13f8e06b4667cf18e386e5a64958cdbecc2
z466869da2ff09d75dbaaca4cb37650050ea281d7f3398f1019c98a0e6a5ad185e05230a3c025ef
ze5c9f1b50bff02b9f2020bdb35d5434a5cd5e973e7f08cdbaee87fe3aeac4fe37bcb0851c33f74
z70d81971cc005d881c814656ff2ad5fd06ddeca8725a0d0ca2608f6ec9dcb54e3a78c1a6e16dc2
zf82d449768153e48c93fb121deac4454ab602f204802b4b444563a84afecab298337e5f8310820
z5ab71869839a776ccda22925f55fc7896615bbc4fd5c4fead6fc3865219c82fbc13a353203ce0e
z74923a23b9bb0b90c2c586202203137cf883dfa2cea60b8052b61e3b716276ab41761cde2a0255
z11dd73006ae80ccf61978d92fa282d5c907fb0fc802ff7cd0c78cbf9768f3f5eaf4fa3742a8ad2
zebae0be9fccfdd2e07dad22f8a355e7ac8a4b1f5df9d1ee0a761a39f6a5f4af6b2d5f8337ac000
z09db534202b6884b91ed3e1985c027bc789f2e43252337bad7783735d9470409cb5a5fd7d5384e
zd8d0f945108e03485865370f6ec7d490bbadb377d56cd315e368409facfb9785ea308a237faac9
z9be856d6907a6f878abe1c226439d409693de8ed1cda0e4713d9e0d508790702bdd8ac04bb440b
z8e8506d6d915b5c4dd9f3bd3d9b9cda6489c115643b0d20e2fe0a8c92eb388b2150a7ace425dd0
zbe60186c97d99a85148fc782ebd74b732f71a986fe30a94c821fdd7ec581c45202984f122facf2
zea4ea17139d175c6849e11bfc3e24738a7bbfde09d93f9c7bceb78e469b1d8b44f608ac5c01efd
z906d88fc472f0784ecff0d237aff59803cb7af32a27c7d06dbb3fe89879e0f6e6d0013298350e6
z30f7b1479395fbdbacd28d7e2bdad11e1bfc6d2873027c6be230f87d58a661692240449959a3e3
zb183a7b9a9e14e481b5223f795a32ffd693fcd80c78a1ef8c302d232450240e0ab3f1c4afac44d
z2a5bfb58b50bb675f7191cdd51ea9851bd3355ad7c4c00821121564ac4f5910fa64f9e4c25e70b
zc96636d636315de474312a67fc2e941de98a4df22e65db7ad1905ab9dfb44d1ae7f35a2b955160
z73f9b4ff8f884f4ca03a2ff5ad91e421b0c503f52cfe604fa2a1a7909fed5a389554b9fe70fdd7
zb36aadd0e35dc5ccafce667c2b626e9abec82754f173f4c86328f53a307d28e0af8fbfa53bfdc4
z27b66f8fe4bc2446cf49e332003a0c4f7269843a27f009bc3370434deea95440e25b16184afc9e
z4ddbee7079346c5ab6e12c62be1bbad9f71bb3d39241f2cc69a8680120150283df0d3b938348e5
z2669417c71042c294efe250a14e4368f69d2cb1e3d5b778489ce338c963ac2902809ff20c0c864
zfdac47609fddf40b1b6b33d734ef451da5a563b396192a047996deda2bc36f346d903ff6b11537
z76189151571c0478ae1499aa0b07f7cb041c415e15109e7405f0ad8e283efb9fdbcd52b7521ad3
ze509d47201cbfc5113ede8188fb843c5114973a551fa74cde04d779f8eaac5afa12a70ba824452
zf973b3599669876cc46bc5b23aedca973de5ab0a97c138e9a5349907ae4f184088d5819c367e0c
z8ceec5e9938000af51b8939b690a35e4be47cadd88242958d3a4ab2c20e71d3059f319c5bffac9
z88e0f4165e1aa34bf8a935625cabd8f15aa6b5888912af1797cef1928b90b023369b6acdd98f37
zd5b871fd62de7d789b0d4495a09ba6673a17aa5a13fcdbe7c3eab1284e116e2b7c167425d5aa80
zf86e353e0a5f22007636c243c29c4c448bcd9e7692ed662b819f11869eaae02392ff8e708769a3
z296e4dcff74a352b7bd077b988eb1a6c49a538ab3a76901a156711771f7395dceee67e183c7416
z156ff60f7f888e53ebb350fbcd345b56f4f31ab1eab9a3ae4d3fb752e24b409b94c9ca1fd239b8
z6523109d6e4f755eb6574e1face11917ae553311f237c73b80d3de80f8945b6e88c1928a21fc27
zc823ca7d50ba1595692911ff86468704b7fed87f16ad5ac17148ff44df63938e8c5f12b841697a
zc2f55442e380ca02484b747a38a7cf32cf093c19e8903d1bbc0d27f613fb8838ddb1eaeb054fc7
zb94a7ba645f846bcc239d73ecefd54307f42e4a7716cfac1fbf2ef88d5fb09fd94b8a7bec3a285
z6cbb66c715b6305492c480f358f9db85f0e43215d5e51a0814dd4c911487364acaf5bd531f3774
ze47b2a55db1d85221c60c77f5c029a25d46d866ab89074921a4a068fa88972d1130ac5d0105a3d
z457876852b41a9565c105dccaf3e0c0c2924139d14d05f858e945decdff08700e57d1d5644b973
z8d3e839be9e51240a352fe65af8dba3ab1eda69da95a430ee4f6a7ef562ef82153e5be765b90e8
ze5e3ff4ec10846c66e75a6dde088b8a8c63b69977dd748ca65317051546a0f021e9efbe265863c
z23fa4ff434be11b72c1aa72737f0627130e80a6fb533b9c629b6f88d56b1d6f3fef31c8cbb4b4f
z8caefb986b72fda43a7ce9dcc37ba222f4e9d938baf0e1743f65a0c75217957d01ecc80ce3edf0
zf09570c6c9fc6a7639974f4cf9a4ecf7e60e7dfe8ac669cf081e7125932ac5c724999afee79ea0
z27c336067c915e1e402b3b5ce6197c997fc7db55adefa1ec08d30f54d830d207d7ce7d7c13283f
z2749394d6736ef648a07fc2b567f7535fbacdb1b0c873697331d7812fd12b94960ee7f0534f8de
z57105fd8b85ace37cd10447ba2f26598acde344f1c512eaa1c1a60c02049958eb48f4e8d818fc1
zc25f8b71340c5dc9e58cdd42338a39971df45006beef346b7eec4e6b7f0f3d8ef64cd9123cbcd7
zfd455e586e01a8ab27fd1bf21d494d871a0f12b3259768da986bb5624bd11816a00803367a7053
z20e0032a74d4cff9b3df55c72e06d0746c17a51712cb69a1d6a5d89e3a99f51b9a0be5d70dd833
zbaf9af0f442169a9dff685fc5b971afa6194ff04a9db3bf34d41930db1f83f413432ebe8ffef4a
ze49659894ecad6bfef49a1dab3fe30120d8f782ceb08a42b0526106bbf8a4eb26f7023b2ef5b7b
za96e337641906f92685d88fb13096d2bf195a79bee7a625bf50b1b4d53d7a647e1a15e6ecce02f
zeaa284303ce3edbd32b243e83ced3cfcd86166cca7e810f79d0f621a1b40d3293d3d4ea78774a7
zb2c6c135baf9d83de4ed655e57ac2daafd8ffb648e539ed2af51463154360c3de82dfb80006af4
zc09b32552c21920552431a1220de0794a11164b5207be15072c5d2d4f1cc74c8b520d3c4d3a04c
z7db74661baaf1f808a9b75646091fce65dc79ee9d1a04ece14a65e2599bf0a8100da1276261dd6
z23db7d5e2536564666f531d8b5a9e2a3cf2ae9a64c34cbb8340bd852f12c804e9ac884eeb20984
z454a0f6c6922a564d98403ba6d042aec58ebd330c84a2a84c5d2b95ad24be1f3a64357eaf14818
z9ec348ecfecad584910336ad462a9e5a9fe089ea056cec67fbefe997af7a38599187f219167971
z3424871db831adcb96e9909d1be649101c5e3e262bf1a1819242622347d3618937358ee6d24fdf
z3c054533a73d3c12af5f3c4c1d9a97bf540397b20c894798ad9178786814b5a1d41bc17e9f0152
zfbc3bbfb373548aed1e52ec8c14f5437a19755b03d4f30a9bd7946874bf7c22b194d94218de43d
z8721bc856085eb4ec5c491c35ab5de78cfc9bb890124357af3a3705a440ac368840f01c9a29359
z5ec8a551659baa925b7f51667bb42919c8136c3b03efb42c69478152617289e8a9ddc4d796dca7
z2982232f8b33d973cfcffebf5e6301494c510414e9a9fa8ce62ac154b611596c14451473d6a539
z6b1507303b930061b81e117de67a0e67f81fa2f552c6f76e133c660277c8d440531e7de894d36d
za86c8873b79b9d21d955732cb166beaf7c7523fe1af1af00ca3089fded4549adc4abab9f9535a8
z89d76ad9cb2980dee0d7dc777e6ac744c815f2e2e85d1f338eb2d289cc5ba584ccd051c42ac383
z5b938debb69f286cc2f7b1b9985a4ba8cf0c1f79c1afbcdf5b0cbd155f6c839cceb1155d7232bd
zddb65b72af7faf0fa089952162d5e5344249d7ed7904d2d6394b2a1f03a25c1d29b3b1012f176a
z87622a2fc118e7fbc2476538a46013d78354449e7a548c34278458e2b809f72ac37fbb84396e1c
z54f66d9b4f3b4a1a64bf06413c9f78b65eca96a04968b09766997cb38c669fc18b3360d4999ab1
zfdab8b5c6b211d352a9a7d6e9c1112189b937d33db84d5380247ce9ff68e31f3ff98854fa78380
z6e55490d74dec33aeb8349abdb6bec1474f8fee3dd8f4a931269c60eeec8082add6d29931e764c
zd1237704a2e0f1a1d3acbabfadd9abfec5f8e8d441d221d595460c6ae41cc055cfaf32d7342995
z0722406815db2d2af51b403278c6b1b5f265783fe7bf61cc76a09322c532891a24679d7d043de0
zf3048a18fd491cf14cfbc32cd86d2f7fe0931bd3cee29e568f3c0d2168694e58a2be3d0abc9286
z39c71c0075e2fc7117dba3ac8af4a362cc6c5257b74f0798057a8c18e440c9ac9802c35ac937a9
z0ca6622fa492cc74aa2dd3e3186e5f3eeb4eb7e8eff00ba19081888dca3647fee17f9dcaac8420
zd9198d01df22f2019dde79f82e37cd15cde530675c6fd9c8bc542b9191fde4fd799a8f49eaf6ce
z90d8520fc109487163930871206741fad2bcc5f71aeada98e93c4bd95a14011ef32bc19da4f8f8
zbced68ede92aeb7224020c6f2184642e41c6fa3f15ceab32d866da5404fb0db6eca3de2cac4ac8
z1396f57efd0618999b8fc30be5308afa566f316e87d3500d559029a5f3ab9b68cf42a3eed7ee34
zb311c329b40c699b76aa4b44eaf7c71709443e7c101bb71255effb5982403998c742f96c149ed6
zf1ce0e0d63f796ae189d6b3a68fb93216fc3511d8053878a4d3e9f8e65d7f1f8b21ab782853243
z8d11046de53fd4913f6f2423a26a7fc917bd765365a2f41390592b86689f5c1985b3ef40960e13
z339cfff8caeea57c7b0a39264e89124327b95d6f13e1f826e98430a0aa92376fb1ddb2124bec3f
z3baf1dc8775705c92ee05fbebf42dba2b2f42402e0c5ad7f321f68d2f34d2431e176cc4cbb48eb
z6f2ecbd003889cce1d095aceb6c19a1652bc4aeef81b2f72befeaa444760b2e3e32e7d1e57736f
z9b5a5c96b09765ea92420562ef7823ef081933f9cd6731a5ad5b2f7ae195b0817d565c0c040f6e
zf2c410d7fb7285157754fb113dbe609df26dd5175ca6be092dd8c81e83a51f3bb2592158a2fd3f
z18d7b82de65af97c785edbce6b7037960aeeee4b46e82e24f5fdcc9e9a0b7b7c2e33c6a30a705f
z105c2801887f45bd3bfe66ca7ed119b081ef643bce09a6e124d6aa79a3bcfe70b2798ba236d80e
zc4240e2f9fe98befe316331c7212b67ce22a4f2403a5c2ae47343cfbfb349cb273cb11b53384d2
z9cae7c385feab6c002821d3c939b6941f1d34251f9e114633622ad22b0b311043d02830629dea6
zc905bc71b9e6c97748f3770b7ea52923e20f310ab3da9f7cb4eb38b861d505ccfc00b352e105bb
z200a5f453efd44c30a1beaf2cb39f77eff1df1951c4a9bad7ca9bc710a3493ff6e7439d26a1d1f
ze23f0349a54568a8cb02af34d4201bfb0abf30edc0b7f3cf412092139d0300698982d184e7d1bc
z6dbfbbf6736d59f96040c33db40ea75daffdbcc832a6bf6d1dd3566018ff60ebdcaafbbc007c8a
z811b05a88b16dd0a2691710f8765c19aaf826b0371ee5a864a813d87256adaf602e48e8aea019e
z9730b6664b21cb57a9d6a5397b128a155770e5e4eab3dc0e312b169f5454270a8b2253dfe1272a
z2bb741857ebdc93a77dcfdebef42de52ef0d113e11a311158bfa4c56dbc80a5a306fe7fa0c63c1
zff1a034285b1408640ac18d19a5aa14479b6875bab003722303963d3c69f142dc96ce86b7f7baa
z4015b6620e60cb7d9a35ccd175207f20b70b5685af92bbbd0480bd669e4a23535f91c068b6e1f4
zc8264617833081ff54f57b5ceced87f55c3e13a23349aa9d9b16963b939b6428885644bf544626
z538754ae746572da508cefc85afab55f0d98fde81c68e61588ce3f70b8fea7de8bd7084a945887
zbbe67e84051b093b5cb099ff6fd9d6a7fa36195d0e93e7a95836dd36cb1d1645c9c622813d36ce
zee0412f4b060f8f3a55a293eb20aea1c4bef6982a7a427084cf96159023f396d94653472f8939b
z4486671b0497a8ed10b050e52f8560b024e9d5394328413c7c55078691b487428978530baf531c
zc9b3ed1d5d6878dfb16ae19f2e17d5298914b6c899bfd1cf4ee559b9a1dad39c83ddcccacd74ef
zcd7f081d00e9985b6c0c95d8735c7fbebdaeb3d1c2d0d4ebf0176c9283f8d39efffabc4face15e
zda4f72d9432a94419bb10c596f0e050e8214bfd7c4e83c429fb6940839b9783e1aa9398c6934cb
z80d4288d6c3995a259450a50937f125e88ccbcff5910add5bf899b68301dee401edad35dfd519c
z70b92a89d3bf1ed0030ff06556b24eb8b2052f0d01c4503ea22a39f6d7faf5b80ba5ae4162953a
ze5aa9c116474e011e4ad877300c7df1989f108f8a4533a2e94de21903fb5565b9c8194864c6e4c
zc1ff036edac468e499c33b28dd3e9f6be6c7a54c7a74b1a92bfc0b69ad36db656ecc1d1ed88a56
z94266c7cc3ebbfe0418d475d5e3c06243deb2f8653a88269cd65b0ddbff9bc3373a27e08a9d892
zd967c4b56e18fb37610f3a7176c264ea10ca0e35c6d29c358606072cd8b9966fb4c28b33f131c6
z47fccf525a98583d3e334306eee26cc3325112b05760304cbbd0e381f595b5d53f097d9bc35c07
z15c6db329b15a4a344ebc77def88a6bc2717d568557452f07b65089b8233e481f8d1c3081627be
zf31c16da3fe91daa16095166a8f4991cbcdecfccbd635e5fbd67f37dbe1002ba554aa1ef1d8f03
z022b7700d71e2d22f7f1b7c512d4c44ac2787f44592c1dd8e92a5abe30adc2c7ec633400722e73
z41294b386618f9ad8a25f350709e1c0b37c8c00622729dfd0e59b9955ea72c990a1fbce1cd26bb
zdfa8e28376b6be7687f02cc11c9b734ada98b0145e9c18e0dc823d3cac20991ab09b6858a9f873
za5cdee7545ea2626638bf80753c81c360ca30416265cd2aae13d7f5f2165c86042af340346baf8
zd4211153f329a75b87ef2283824ef3d4401c210f232f33dbe0ab825c85208e5941b8847b82373c
ze6f71c5fa020f8c4db133f3117ae6c4e1826bba70bdfbe9e251bded859c66537b0d7d2dd022151
zb65778be952fb614bb40f1b026a0e34df263923d4d7fbd5661a99cdaca8091ab55ee2e4ca404d4
z8db94d0c21a1b75f083093dde66b0f0bc15442310eba8c12adac004382f2fc2bf86b20fdbc239a
z9e895ef1cb843edcd780a3b5cbebbdabc62cea76ce856971bf009868a29a8934aed02f68c3fbac
z66ee6f2e1b9b376feaf6a5463ebddb47f8a7e5e92f243ea676c8c4b5f7dc3e91a5495ffd1a95a4
z5d009d2570fae6a0f529825f167e2d3fa9f254f0e38a7c21f7ca80d467a1bf5e9eff97fd6a5294
zefa883048867a2715397e9fae95ba4a38b9f8d7a622469ef366b772693bc7ed79527a4fffb4bcf
z4c79a1c3eda96639916a7d94e99678fd63a0c2bb0f3b3c7955f4e34380415240eef36de5594cb7
z999bacbc5b418ab1fd869ac95fb9449a0f3fb9c1abbc8e9be0e08f075c9726b686f1032b03430e
zd18595e191b810969717d4f1f309ffb01cf1955e862c309acc8afc7e8d7cfee870da571f1e7ed9
z72c33141434f700286a44508ab6b442a841a53e87c80a113e52d33371a13243f9f84bcd4a4d3a1
z3abe823877de0459e29cf90036ff42a11aec8a7a84ea5839f29999ee900c1543c8ea20669aa67e
z4f97433ca4ceb8c887bb3227c4b832779db80d5c2d167c298c0000ca236e528188420f68712dea
zf1349032ab30e0549563c09afd8b021b3852b708558302d3a065e32befa3b0479eb461d36648ea
z9e648ad847a3a39989ead16bee65b8075381b8e634de5061b98236fd0bc5f815cc7c91145aee50
zf9a096fa5a59abd015d3689705da8545f45e7913f1fecc98007f8f8ee5896abe2fdaba615de56d
z8d2075ba9711c92fae6645ef732990571ec14d53a518b5cdf3891b884a54d62f97751c82223aea
zf39acbf59e2cab78b1434def907ee5c3e8cfab94417d715eda8a92299ce158be763cec1d633b9f
zbaae81954cc80c602c5afdbb6bc4976e5d3a1951a724a6460ac8ef205dca287cff35c3366f6482
z128d61b345a43b4055346fc6a2c20d27ed08897ecaab1c689383eb526c0077c862345e264d693d
z112657c548956210752d1d0bf841ebc7d8301be195bc7230b5623b3ed2f0ff1a9939b9f972df8f
z5146f2d0c23df766d2fd1ecfd791ba34986936b812c00a94af7e22d656f17e1a485580ff8c9e1d
zaad5dd9842a3bc0dc75d916d7120d80a7528a8e7295be3ca7649b07f418e531f20352edd31e07b
z15982f315a0d521bc5600bdd7f7eae8cc8be969505ac50f7c417d265664530b18fd66a032b2f61
z4e5fc966a95f98ea9afcba39be256e30a3795a6f220e642093659fe2abfc39ce80961ebb292141
z223a2b668b4d37066d4ad3868dc934b5569a58f26b7e3b2778a25d6ad8c6031a7a7c007c382f2b
ze2aa9dbaf4688335095e100214334261868d995bb6ca255ca986d69beee799a5d26de652428248
zf7eeb9c5bf00e1f74e60bc40455fb00a52b33ccaa21638299744a864948891b0316e1d32951ee2
zca1c8ef22e60d4176571d5dc745f2292779055151251033c93547f1e443d72dfee71557973ebae
z12e5d7b1d3cfe4f4171e1127a3315be307e5db7564285c56810043756035f48d3f8bc47a3aa667
zb3891581e7e7566bddb2bec5e6c11bbc05d3258988dbb096cc04766f23c18a43f684fa2f18bfff
z925a0c047abb1d63149d99903514c0be7affa9c7d7508edc027b07d5ec4d619972cfbb2791946e
z3065184fe6a3cc0befbe14916c6534c01923a7fcf76003afd070954e788f3049268fa209144092
z977075d08c63b6dcce70103318412ab8789a95a0c7141feab7358a09b7d75c21b7c47f9a131ab4
zf7164512f9cde7dcb98d5d92de4d6ca67ddfbacb8cd844a6972ac6bd9b5d617f3f7d9bea37ab72
za6f46b5b4f79bb8d1571f48c43651f445246869845121f99057a6090eedf8f1b1d803b402408eb
zd86d6a252cf7a3263f07ddd38658f53400288c4f4b9e193e7c02e44c77cc4739cf715b7421271e
z09d763eeb64fbdaeb781cdaff189b167cc082c8a67e5103f66012e6c45dd897c117b44e3ca8e4e
zc4bc032ffb32dcc76327a684d5d97a80c96ebcfc8d2395588fb8b7afff2951c53fdc277b7b88fe
z8a9a6498db282fb6cc7f021b6633aba03c203d1fcaf80613356d6c582e55008be1e69c44b7b180
z1bddff6eb46bf05dc4c3dcfd45e8eba63e88e129a81621dc085486c5e24b29b2d0de9782657b8f
zffd813200176f3963bf8b5988876b63e161ca0464f345a887bf3e6ff99013e25c7dd0648b34e96
zc4a2840635ced6e14ae352d50efbe6bc34103defbb82de3da0ef39956046bc9c9b17b2ba0881b2
z63e78c537c847d73057bf7a4b8800997cd30c0f58fb1853bff6699fb8b2e47a2a79cee2818a3ed
zbaff685adc90ce71ad323295c611f1f248f1a681bc5747650bb643d0ce16f99be2ee9cfa3d4a05
z1d789c1c218b5c04c4c951eb1aa20cd0c9d8e22557fa735bdad324d44be6c92ef0f363a9da0a94
zc7005dd6c42d8b9762c5ee703e9991e2de7112d662c3ed033372acdcdfc46ece6a21c7141c2cfb
z7c19cef0722365c8e32624a11f012874ad4500bd676722718678e2436919c650b08b3c82fc0a88
z985c4beb9b159ff06c40f7a926032f4d10ab3854213ef61850a03e6c0d114ae5c792e190ba5f65
za93df3ce9c08a4dc582da238013798836267714778e9e172d9c51558351f6cb76bbb165c85fb03
z5914b523d85b5b7d69cd2f5dfdc251d094d6ffa7493e4c07e80cce414dcaae6e6244391e4f1908
z578a4ce0026b867b3087489785f3f5d10c0f5ad1058cf6df4b885682872210d9dcbef41e16b1b2
z597aef5bd556c9956148dce67fd9805f7c22e9d8cdbe31b4b3bde35d4e07f04c680bea85542cca
z0f1fa215e7d2542fe976d1d7d5e2d0a9c67ab0d42e66a92ff8348fd5b8ed7add3cc5d15d4f2a69
z71db2e984966c508bac6493bc837e2e825d828ec16a8316d195bc0a16015a15f7bd0329d903af3
z1ffa836d4dc01ceb3894ef91a61bca4bb8279af9013d30b29f00ab276040507631771a992f7a48
z077dba37fbaaad2cc661bcfa3c2527a258c7f1d7c7830a42714d05bda761ae4381d120d9cdfeac
z3fcbfe45382241e98705426e31e1fef0aaffd820b59d3fe1717ab7a1634922ece625779b4a7eaf
z65b7b5814f18df2c3055d81fc889d0d42bf4e2ce74f37e7eafca92a0ab551ea39b831468409f69
zfe564854e3c92c097d07d08e64588f8bd0a08b1012ed996e26c95de4a1397942f814a0a0dfa38a
ze086882f806ef72aa61a7f487820006b3316b661cb6d42800c98f712afbdfeff0965d407516713
zaefc24fed00175a664680091002ccf98bf49e57a444eea69b015a22b4995359a3544dd7d29a417
z7950d44cfa94964718824abdc021ceb4befbbe77e4dba419e0d61fabc7001a5737ca0e3cfaff3a
zadb5ced88752233915e35912a654219ef32293d2ee89143072102ebea9b078e8cd423cd1ce718f
z7351bfb317bc44bc2ebbc6fafa818de273f1ad880414df43c868ae6fcbc482200f51d8b4d28efb
z33ddbde112bbfc4d6435349916f2f91d2bcfe6b6df567c50e71e4aa8df3e9e97291c33010d01df
z948e5eb52c1c4166d569a50e9313011436319392ee134dbf53b8af7371ed1319ef6e69926b370e
zd75ce8daf4ab4554d4d1389064ecf46cdb94111dc844a01d917aa66489629e5fe50b201dbcd1ac
z830e8a07cf094937f1d48fc975ce4f61d882632e29c763abb254f309cd14799d8e11af9e2af993
z406ae75dda23a447886cbc81deb2621ceae118380974b8fdaa28687baa9e776ad770cefe191c1b
z619f4ce920d07b858c6e14f6c6377e3831c48a1939221673e6c771882a0b18458713bf50351d6f
zb763a10bb9b6ecd2cb9652ea096837bf7e58f6e5fe87e0523cdd273d409b23350c095b797759e3
z7cf3934ef889ea6083bc2bbce56f86ac38a221146999baa268373c8a1263f0d74c40bba34f2f25
z4cb5347e84c289ebf4738d38716bb48a928148e238289515ce358f86c75a722a5b8bbb753fd413
ze9d57fa51f1fe194521de5d5bc38ef3038c95fbccb15358df373b1190cad27b0fe7033dd82b8ed
ze8b3e0db11a166a868f686df59eed3e5bebeab6f958d30822199c231094435678a1da2c8f36481
z78327d7d738b0e2d38e0fbc783f1fd7984aa62fe6f7088b9690966f2e7bc3278993d6a32441a1f
z4fd78355828bf5fcbaddf5b3774f5fda341bf35e2e73a1cf08eb51c227d66983d27cab57d47a71
z62ec43b2259dfae0747d4609d042fbc7ea93201062407c19dad19f2487d2d90684a2fc481f6c75
z544595930e7c4bdcf3df200863f2ac1e74ab212fffbd26f192052800ee1222deb81db6c83b3cb2
za5118e51616300f44a88d1dce414b72a2a50634da4cdd901068c139de7c46f1644d1a1bc98b76f
ze19af7b026841b6d89566e25c20663d08753644fbff66133d167117e7d1e9d96c434874dc62a55
zac3de5ad5f4e36aed281e803fbccdd7bbc755a804674fc22cc23d1652da518adef8c480f4cc113
z74e3868723abea17b725d195054e49dd8c848d127f796c4f673e1783b3ccefdb15c2847effda9f
z44c44a419220675985df822d1c3c1a2f7e06d9cb7cc727349cbc9245d60f5f4acf3ca06d3445af
z242c3260977daa84352e8ac40b708b4fb2c28bd5a7e01de9197ceec24558770c912e62da223391
z1f1d04a9b44af7bf3131a36366660c225c18ab2569381c50ccf1f704fbb33e45f99b5352677788
z83e1de1f07cb7b96d7a15efc5ba3870787bab165ec99d77cb0d1899ce1e9c5ce59ccbb700a24c3
z43b1743e5a8c2bef75741309fcb0fcfaab70bb7952b6414fbe44b44ab49bd5eef942478eaf1704
z9586ef91eadb66c9704008253b327497b11b9260bb67cfc9dd5c05699b76eb3bfe220feb606a76
z53bf76acc851425400c469fcae8e2c0b126e73ab3d678366074bdc13aadf4f97151d97159dd923
zc7baddaf5ac4ebf0cd07fb5bab75edfe05a012ea9da8e17758907bc3cec1ed6b84fe954f701bfd
z6f958e8b33531cdaa8529693e7ce0087621dd9d55dce09fcf76adadc4b52fdd2e802bcd88b6475
zff9c8ea8f0d45e88ff5fe0728876e81c0000218874b1f8626cee53f9a04a813ca22626c61af884
z70f73d56424abb15b373a56a2afad12070ab8a773d07828eb8a70e91933184adbd9d88bb5f3045
zf4f63c8ea8cd68c7df570c8f8e99850bdb45d02857c5ab918341965989310434765a9e58679a1e
z8ef6e0ea11765e2a79110e762c1670b60b4c285fa18e2ecdba6726c247677a7ffddc1ea5019b2e
z400872ee7d29a26c007253747e1c47cd1125cd1f80918643a5e0864ae0d233d3f82087ef2b917b
zedbeccab41dc8974872534bef76c784896a36723adc2c410a642105c982329f2a0ac730a940274
z699753ccf32e8bdf0fd1e13ac0fcd92e88a79cf32b6504aa3a3f42dde505ea47a9c36a2443f296
zf2aaf9c45c0a6c0a9eda0770d4d0417a8a87a9044a1453b5051193f14ebf0f7e68bae1c912dd95
z38c7ac8cf4218b87dd54c9401cc19ff32a9cc148e9844fc1f63657b4d47aa546de75f9c8a61b4a
za2ac1566bf97cc237cb2ec8729c5b57d5b35902e4ab09b3655d935fa44d23eddc20e550656ce67
z85e984985616dd43308764f08a010942f5c730e87f6a040c287cccee18006ea5311fff7d42fb7b
za2adb112808cadb12c2dab7dd43e003bfa3b6c4dc3006abd3647ed5053e8e95854508a9d485627
z0678edc3f50e5a78eba99f7e104424cdf8d58771eeb61913cb2fd0693d308c1e35851d628103d2
z7ba82fa46ce4285cb94391494d48354db077640a8a0e364bbaf30f70c80fb9fa3927fb9064516f
zc2f75b1c6199ed24d022c3fa975dac01c5cbe6579cbc2376d4f668756397777e20df86f948a5c2
zfe12303d85fcd7e98631574083f5bbcb1896cb44f982966bf4d1c9934bbfdd5b5df4fd295b79de
z4c0c6765c97cf100a1c8fb3146bba45023784534ea57ef372a222c11d913ca036eed7f2616ce1d
zbd4357dcc04727413e45870c2497c845b74f510be5d97373395682b910412c8177d3f5de7e0dea
z44d0eb1986ba725bb011e590a902bca4745fe82b51eed8ef710f68d6174da19edb7947a0e82217
z5179695a80293fbd298d46c7125c80de38b9dc5a90a59e99b8b230c2fdd1caa7d8bab51364d249
z607052f85551a2a31d24d45533be956a0dc22976d0657c38e25b065d5ab011152823db13eef157
zd204b389791cce9dcc8b9a327d49536189698c5541ca41daab381bcc2a6c1e97d0bafb1b558752
z679b2f389176afc6105ef339b94049072e628c6d9f862f6843f38e97c70bba5eac23540544dd1f
z1046829b5739764e71a26a1d2a9b5796d22d0914ac1ea47869e3e9c1b940e0b077302a15a9f9c0
za770b79444d2d62bbf9d9ee85dae7e55758c0cfc0dba7e7cb1ed1dfd16ed4782729553d7ff2a46
zf9ebede523088f4ea730e2acec904a6f4a005823c7d0bfa05b908ef11742d739a21b97c836e810
zb53804323a1d2f8cb45e6107194615eb13b634cb5a97e216561ab522080dbb10c727b5e126e4da
za412df53ff7716737872a1fdca4995f0972b24f5dc1ae166445f89c2be2b826b89edd142ee7a5c
za9fb7277255d575ae50a9f2197dccae243a04b115a980aa5c2ec607559b4e9e1155f7cc0b5828c
z19f5cdd8228b247a4c7bad85b42f41054737bb5be892d9faa4719eee1a8b5f67e8d04b9e9a5a69
zf33bb97ec7ff2014fca2bf4d70ce7e0aed40f23de4df038b9699482cdee1a0b12990934f903a8d
z32e5da9ab710526b4b6108334de220d6e3e77c4d925ffe65b4db0434f137070bf56e7ff2c2396e
ze97d1db72ab1d4189e765b9fc82267f0ebdfa8515202428c4143bd51535898bd0f9a20f49e626e
zfd54aaf322cda5bf7fdbfa9446d0de8a0cbe825deff7d95791a87026323af044335fbf1422e5cb
zd815bb6865826400f787ac46267feb26b844055f1a3e7fe7764a13f9e4251d0a3115664fb3e704
z5aa463dacd36c9aea6a46dd1bfb672388b567bef6b733bd1232d204cf0a26b56a6eb35dbb03798
z3cfb97c8bf9f543a0fc3bc52b3eb29483525b574427f98a12088ee01d1ab3b9a3904392c7b6376
zc0397a66d193e6aca605e2a7e0923327ac7e713c68bbd130a51c5fe759698c74e67045c85d3afb
za90a068252539944ae4cdace6724f47726b524665b68b836ba45c89faf762b3f5699354d46f2b3
z9e02ab1e63b6189a853ef89c98ad3112382299fecd682c0a2eab210a1a58266a13bd76a4c4ad38
zf4c6c83000e4d5383c07afe73eb25a53904885577b4e5cca332ed13653d56349391021ff08609d
z0eb601b2f9fe2623291004c55e32e6b6d0c502956463b925c7ac9d41a98850318cba9ac23312e2
z7df13142d1c22837d0096d9c0924a19bb8cece360921765ce5eac5d8fc11da40b5ba6b42e8d0c5
z0ed8d8f63e0a1a3600208e1a274893a21d6341c4cce08c92034be78a3f9b5336eaa3d0443849ed
ze3dff3415a1f7b5d69fa8dfbe842355b1eb0d1eebce0c3f2f07f9a59bb2bab1095cc71434f599c
z0db463d586d0340621cd569636a45cc41ede47f27e9284c08995f381128203bf42ceb6a033ad3d
zb79bcc05991fa2e6b91daf58aa63285a09efbe3f998ba67f8533659bd06efe87c8a9acf8e5e26a
zc47596d264cf7da809300849ed9da2b67a6afe5fc4812fce9f1c16da897b40653749e3c533cb5d
z364bf22124a4a43446ef72dd6d62e2e0491ef996f419b39ce44535c71f4ae7d18f2198e15e26b0
z4776815609940f95a21fa3a43aea648021ab0c760b1996f34745207b000d7bf981a5bedf7aff7e
z78d0679bcfbfbd67af51e0d6bb89dc5c961375b8d93480274d82d3beaee6f20b526c3851bf5ede
z949b5b3e1e14c5d81474178b1efb11a6b88d6e8a7cc5653deb4f9685fc77450a089ac01c65f3c2
za6830a22d25198de22b5a775a0327281e23e6f6f391b8f131052d25f3b7a7bc1cd83fe1386a07e
z8ef125646c81fcc087fa90d8906371c9658c1d41dff8975662727172cce789580a8c5d2e4b0324
z6cb14f6445d5dd3bbe3ec2073440b248406f71003671ce62ae11ccc50cd5e113e4088adbe76ab0
z0e128b4ef82d16ccf59cfd4c979d1b0f41e334a17c38881622dd3f816dde7f3690570245216102
z1a201471082477406ed69e23998ee7775d241c0c6cce28b0c34f46f41d6e40b7dabb065599b7c2
z26c64989f45e42f11bd5c3fc6acda99a0514569d42d5a376adcadadb48beb403cb391978818fd8
z125b70f0ae3cb295b58c4c6ec678f1fc16e04e3289bdda3465ebf34bab8c558834e42b4e85a117
z90a533d96128cbd76c67dbf7c2d0e8dcc4d99d61d3cb7d788023a5231893dbb3d14aa5972cb3ce
zcab2d46f033d96b1db3a46d92b56a1beeda350cd8df43460e706169c3c7080404877a0d50574c0
z905bb3989291e1184b689e12f3b12cb332c95b2f65c066d687b588b826baff882315abbd68a319
z6d443fcb2f74b813cc41786ba47aa1061dfc134c3eadccbbd5ccdc121b3156491bc8592bd26629
zf292fb8a7cf99d44034a614b2e9953e73eed89b4e1a982d3edaef89a7f53c89d43d4fef206401a
zea3896dccc9db943e47f9d9d60082779540574e3b560f99eef686f7cbbaae456b71d8813d64a08
z1e653451d5e5ae69c376d54abf9269e743d2e8dab5495c1b9e889a3139adf8b68f0f7fbab0a4ab
z33a92d1a6ab37d97425bf32cdd13789cc6ed97eeb56f2e92da7ed34e348fbc92286986bd50431b
zf91408e8875f41818b816d72b1cd0be3bd3a381e94ff3a8cbf5d983a900ed1e4d4e28ff735e485
z076573a741b92752751e3e3f2dd1f2fae79ba65d83bfb2a8ac00f1da4a49d44125b93d517d9e7e
z75a2336e1a6a5396f13a59c447bd19f0d9aa865acda38108703abe6b75e805386b903c66bec7a3
zd1611b550bea538f9b2db8c7478e8d810145328fb25ba8eabdf955ef2f0557e264f029b0529e64
z00b161b1206a66b9815f40875801ea112e2e7b05a9666af9953518f27ccc1094c0d5a0486a7736
z3923d7c187fbf2f293010ffae7c1381f8bd603fd77bc46958126e70b94e81f1b68a68f672a1fcd
z253c114a6c10f7a36da93a0d1c281cde81675fdc9d1c990b1d1d3aeb460bc77cc4233124c23283
zf12e21be5c0bf69af29b584165e6539287e0b3800b6b1efd97d09f5a6d3f1a0bfa5a11381f720a
zbd86911233fdb8ac86fd5b855b80a955663f692b943dbc14fc5e47339f4862738a4e2af56efd48
z4185554ba48d3bfc35827bb11428ca2122bd16f5e7f669de706d8b7f8f3e92035abd0803a88bf7
zdeda07322d6f41e93771dcb6e19d6582600cf85694c0f6e19b2b2b09e357dc2093e960c7da5971
z987c8c195e34772b8dbc0548e9cb7bd15a0195ce7b5d9560f2656ab36fa20a7d27b66a937fb216
z01b6759d6bdc05441c2800429454c2ddb16777248e446dac1e102736d6dfc936bee545b6350f50
zf47f809335af292175c96c1d1d4fd65b1602fcb85e8bb09c52fff67873ab9452a860fce6a29905
ze6c095bcb1f376f42e40cfa6e8fc6072278a789bf4df563343f1eda173f37bc56a108912e14701
zf140e8993102930806503f7a19165fcb91fdd06ea3ebd9b9f0272c5eab276abfd2225319e28b0e
z237e180b77897a87ebd8a6c826333d09fd22e362c0e251c93dd53dd6bfd0880ed2f8b7cecdfe86
z596acb2817bd9bc242771c703413561a02fd060387c0a770166d623b9d1f6eb178b48a6121254f
za48710f6b1740836d46795aa964e4f578d449f35748215fecbb65334a11c1ec11ce9f21ba8b705
z8289f61d5a8b1276da2eec37dc477a392a437e930719dfbbf8e973fa22d86b8adfa593c24e1c8a
z33210edb3bdb0bb027a565fbd39f5ce6375b0d7002169cbede38b49036c20e30fbc78b2ec96e15
z43194a0b682ced88c2d7ff560bc8a175d2198176d1ad78c732e81e4f56286db26f3c2ac9eb60ef
z456f95c6201639d457341a47b5dfc3a83392ee18025371c890f9d16437e3ee4318ee7a97b4aa70
z4a9db238de6b796b08bbb17d6bcc86e07772d2bd295b8cefcac14cb392676d9f0633810c68badc
zc9495ce7fb68458f639835755dcd2bf6038a4a7d2db7ad2d5cf970ae77efbb412df193fb02ad02
zfb1bb4e02ca1f8d89a4d658aec9530a9a2cb165f43dadcb6af8a2cc67b9e2c935a0a18dfe4a902
z02c8fb65d9bcd1941b2cbc9dd6d56d75c69bfd80b901ca9a3be5e11d1ca87c20a4bb226fc51a08
zeed43937102f77767e5782dac311156c9eae98e4490ffe2cef6ca68d99003e4258845002e3ac39
z87095c8d0004e33498fc13ccda4b1fd8e856af1d7ed62fae7c523df6437c39540767967ffd6fa5
z2737ea0e2f64c456811bd04f9d7a30b2b9e5bd6f4ed6bd756fb9da4cdfca8770cb8ff535cc1287
z99536331c17e09566731b1b841a73c9270b8cbde5b3e3a9d16f5da9ad1fa917e9aacb860653e0a
z769c7542de9ebc96e051cef4917360477aa7b9c1e5339d1cf0f1055bff7e6b9296d578b292ff32
zf7dd08944d6aec89d54f07e2a2d1574672db59745ab38e289f420de0767a6a9c56548120ea2bac
z46a33fda1ef49f28b11249a583ee528fe1f347b9f84f0fa09f5d7a1d73b3850a4c6d754bb79b05
zeabac73981455826aff3a0332c5dfeb72c33d3914d7a936cbb69967369fa426c817e99313ad5bf
zf9a1c793861e73cacac1366a6d329e3060ec457e031a99cf383d60188cfe1d12a5b052447027a2
z33e59b84403bff0f17682aad873b9919bb01af77b0dc8d0d3ce1441df1fac3be83baac11dca4a4
z942ff2cf53a392a4fdc878bc21d7ad3437bd308756e5c46bf0ad8ff1476e4fcfda4f163ffe755b
z6286609555a45b54b7003763995c724e76c43588ec016e0bc4801821e4616a7652c6658a9a8d9a
zdcaa53ac37179fd379eca92af7acedf570522f2b4ed996305789b5ae712d7dd9bcdeab9d617952
z12f8a4369fc7dfe8ddcaec86f4809e5a1b90f7eeb9f83a9796cf322ab44e5d891d1be83f38ccc1
zc782807f3580032c96e80298a9fcfb52bd6343b8b27ec9832d2117d99867ffb7513dce52ea4bce
z70c566199143621bd007494eb9580e9bae73db83912812c49a3df7fe8a29c0f46c57d51b138b6f
z4fbe67cd79b552fa08de15d5990174c4417b72cff5a4e910a9bc78d158a8cf5452a953a690fce2
zf156fecf82e484812955336e7e01f69e3b44e23f9947188022c97c88992fb28051c066abe7cadd
zd8b3f25d601086d284036043eb4d6b219f56ea096ef8b8bb7def4b1337b7ba1668689e645b153f
zbac00d9e742e58a36cbf2004af6c1a9a1b71a63c3ae6b7ac4df7589f54b4ee38865ae3d80313d7
z3083f6f7aefc64b0aa7721648a8b46ec083d93b27ec0cccc850f1b1613bacf13a8dd37812287bd
z6e6990eb7a26de09700040dc2354aef46b3384ade7d7ccde923b2803511fbb01af8e0826e7869a
z3030f732708c98167de4972d94a4750ace290a03e26d514e571b754ea4b7f23a5ee20e346ca3b9
zbfae006566f1fa28c0732144cd8616dcddb0e6b9b46117ef97ce04acb08e973b734276b2af5627
zeda67f15c15f0ec9eac003890a988b50e9ec28338531ae4550d6afd162a136fb4ba797e1528abf
zbd9aa5b89df9dd4745444d052fc8c55665ff2b996fdf7575423f4a949255388db43f87ff0b7e39
z8f8cfd6342c6983d99d2ee984e3a2c7a97e14fc92e574a290be8d4589e6611670c8cbbfe623a08
za5302c74cccfa867211736da4308e48fb360052f0ca0c4b0e01158b2c979546a7de09783799128
zf0f34a0e997da6f374c506dc7397484bf9690b6adb0be3522d0a89bdf4a88497a53ff672bdfb9c
z2403da4f597fbfd368ab063c59920798e4e8c9672dedba33258bcb9d8a517baed89b03ea31333f
z91917bc2ed481f65ee8d3b773b21dd1db3c561e21edfe9f075a93717aec36f613ad58c7c276521
zf4846081557ec9ce674f22c8cc6708a1c71e0ab4762a72fc5f90a094127cc1753bf5aa0acebbe3
z18c87c496340a28da88489f1fe5994d62d59ef988d13f69730ceb9b3b8c1c1e7faee78be41da7d
zecaae37956a7bd7485f1427efb6ddb6a64df97cd8bc3027ff4a3acd5e45785c5f92065b11b335c
za064d42f5ccf5cf82654a66ccb78fb008040f0ff468bec2de9b82372e17e2c6823263704fcdc40
z25dbe15d7980b645de0aa9093a6b9097fa4d24164db578c15fc9794c770d7fc8c61115fe39d23e
z7e12333377b8add7548f6f05bc07ae27df1bcac901acdc1ad5eec23af040cbf80d60e20f4218c9
z128bb2e3746d1e98d5d9b6239b74962e110242e99f387ba0b558c4738ffbfc8b0d1e13cc797acd
z69ce4fab16b69fb3de91a27435dc60c5a25211b64c577d18438802f212047a774b1f0ce828e0fb
ze7fbca9c634c786542eafead1822dd63af07d354c3a61552f88525c7a3ed56e8455a650c76a240
zf6f8be3f0604601ebd060b108b7cfeb7e971bc83f760bdd228839c7218501838bbb3d68aac277f
z8564549f0d165ed6c7b5fc85c3308539444457415eed30e19bde7e32ac274b3c602429df7606d7
z0f31ed016964908d4a077dc3b057fd8b25e479e018c4d8ff8f8ca1e6d59b582fd8a9a19ee626d7
zab05d53cc88d61458dc1e607dea7015cd724fc5ed0154854a26cfb9e92a05225707f917ea5a899
zc654d83b3ddf4f0197acacceb86c9f15389a6fb059c06903a4fb3bc523295c81666ea042fd2331
z64923583dde7f4f3ae54c8de3068768d0215c7fb637a1872e6a521c892340fa522b1fa301381b1
z439b631cdc0625c89ab2b8a576dd9bf776eca8a79d6012b04df44a4100ebeb73514eaac79f874f
z36df263fe566a971d24cc2b12c11847a618b91d72751a17b8bc02389f4920f247e9a1aab30d4e1
z0fdd010d8f99964c8c41f5da055113d361aa2eb06c0efcc6b4edb30d2542e566710b08c6b618cd
zb45516beeba6fbc4e2062d6d3827c39b0d9e9c24a4197cfe9621ceb70de3468874ef379e345a2e
zf5b053b1828a9815b3928ee046f765a52ec8518dd8f3bdf58f5248268894263fa43f7ad88efd32
zfb565640a206a849ba40d5d864a85dad1c47533ba3540c6bb0395eabb02fc4a2e0562cacd4534d
z6fdf263190688681a3f7fb1e61f2e4629c0b473aedab43449b66c927f142b6a57d26377a501b3e
z4973e523cfdca7e2c2ce7bd96e7bdde730f695182ae24a229cc415e7760dc5c7959f153fa20656
zdaeec18de1000615fbbf170c420d4dc50ea7a2710a45dabdcf4b4e60ef726e617dfa8d30d1852f
z5c9bc20d89fc2d9addfb389e2eb7e04c377769e894fdb3ddc5eca6647206b873f690bcd335fd06
z9579a2833a1db83af0d0dedfdfcdd0342ccbd12acd145f3b229d482caba939180fc135c00b02c0
zdb9e66d7758cd5c926fc6dc4cae344fbacb39d3f0a2e4a0903708f779edc09e207be2fc47e62ae
z89e9edb4d6ae91aed0a7eadf8a8ea5bf4a2472710b6231e63632ddda1da3e120113e5c6c1b46e4
z168cb249c36b722555921fefe219f75ecb436d011e7a74875e245233a4fd34128294423e5efdc4
zd5b4fd6f8cc0df1ddc521866f6bb631e0ce372082cabd0b96ec9d7ce88ef5bed35db33304e8a7d
za70dfcdb120b70bb452c14a9d73b43c6184e3d9b0cc569fd0448844e8188e3bc95fc8ef4c8b630
z067f1808612b1ec54ad37da045e8579a1b953c8d329c4b617f4fe0dc77af2989f734e1d1379b00
z9da9bafa108c8321be99b746bf4a29bb270a0f16cd525e305849fda9c4ee4e7ad6e96a6da9393f
z3147dd724ce71875ca193d183abda460d66d1c3a9322a007168a7ff6abfd878fbccc577bc8ce10
zbb37cec7cd238b8157b71c27dd0888595a172f3bdf6d29e9804d59d65cc81970ecf84236ca2867
za43b23cb02b5b9472169ea877aead76d6522dcac950bd588a880cc80e7b283fd1df99c7ce7c005
z00eb2531ed8f1c5c1a0fcccb76433a7c76a26ebe0ca2eb11a5a3dbe05c91ce62e74dfb7a9f1da4
ze5814579f3c3ba4ae0404b2271c642f2756352d164c366a2f891fa3761220d1d67eabd64632c86
z06a2aa8a1061890717eceb9ab60b316e1eb58d4f6d8a38fd910e0979f482b2a27b148d3377fb01
zc9b568dc591412153c3e25eef112171d4f4fe4689005e09418a099b93f0aa19475dde9d1ae530f
ze8f8210b39daa622facd52a943505c2254a165ec0a316f3bcfcf47d0bc7da34fb55fe1dfdf4914
z85fb59acd33a1942bb8b8b19deba5b6a52daf79f62f705a26ac00dc23b7a7502d265f4f2caf48b
zc41c8fa40bc8513e6b4dad8b0fff55b9fe67e9f0e9c02a721d35c34c4bf15ae70c8cd2d4364019
z1f2f7a7f8d1393eaa61c842a14f20a1abb2dd1fb08c888053be282eb2d220c24249137705fa60d
zed99e37fc824b536d2c9c0487ea319ab69e084fc81634092dcdb8e724f4bd878ef4585324315a3
zed8620094b070001f9b4b6feb3de5853d780d8c61e8c7f6f15702deb374f8de23c6d8a1f1cc942
zc0754a668e51b0acb35f866cee085d07ece67f1e8cdec3b62fae71e378c0da936bfc6d6acfeb95
z0e09437ef1facb366d221a581727a7cfe60b99fc8b87fd267fb1de7ec70e4bb245093d26a848e0
za457e5b2d17cdf633ba5700309ad8beda8ada5b7b2fde8580a757ae42bb35bca1d7c754d741712
z8dc167f6b7371dd1414ccb41057208ba34eb7ae76b228e247e597933a2fc4377264c7d2638252e
z432b06a3078ad5878a0bf044be99e811e5330ab69492b23a0a4c9fec2c992f5eb5bbb969cea7c5
ze5326f945eeafc81295aad2b4fdf605cd28ba2752ccac9a24947fda353ba87c97711d4950881b2
zd7ed5f98603747b977d32747b8cf75750bc7ef5b067559c4dbeb7dcca81c19895fa2517388920c
z080d5a8a86c619cfb39484cd5ab769fc1151d3527d9bef3832de93702e3923ddb684caee7561df
za6de8aa292281f64e01bd1558bbadc18390f54f1a78106ee7e48b63d66010772f9d68776552927
z4027ea4e84ae0425bc5454c423f8a43155dbef88e3711c365f05ae6fb618dc79ee5b6fbdb43359
z566ae5e330c94153a6d646c2a5e4e81debf8e8facf65e116a7d4a74d56fcfc4a3c2af7b836e904
z88dab74fb583bb1211bc8e2768e5a2f306053416cb255ba85cc45294bebdd50adee00d431e1f47
z4bdc06cf8bdc3dabe1eeba8e2ef3bd9388b0bcab2497ef5d47c43308f7593a30034a77cd548004
z56e1f6cb9e9a1b3c63f02b9a3372bacfba4b880df87954198efb80045bb7c5dd21595f84715d74
za2674773af9b5a651c630dd3727da14b17f14e6bd41912408e071c45a603a18bc681d24ea62f38
zbcb19970067f066ad9f09ebeaf6021f1b7a2d3118368bce53111dd2c9b175c00e3b57ee9071e30
z21337faa05695ea0d64b43bea7548b6044895d735b8b816d5d055e706672699d5eabd7144b0159
z2e345f4b3a84b06f85fbec2950a3623e8cb130295f6fde732b287cdbad1c4e07ee340329959467
zcc3ee14c361e041801616197ab1b008bde8ce215295d2a32e807862fe9da7a430ec7f9a632685d
zb9b9aebe07a28ecc0b76ee5b382d56905685666e930414e589edb65d906630d20dfac387879312
z47a7775358e285d3e720b1cad37a8123ff56070d0091042a8d6c5911ba02bacb34397aa6104b93
z2443657233878aa14fb23d2a9eb6cf4fd5da0d92974722a6f542729992c3d1a44e30632c529fa0
z1f71a9e3bbc01dc9cf2cdb9dd42e7dcfa11f1e50eda8e7a57a41bd87bafb586a89e19af42b55cc
z0d2712bea072edc954dc9189e039af9aec93a87fd3a2723e696a01cdb17a558270bdd0c2da41a1
z8b84de3d401e32978a1bb9fee17985a2e1121ae05a088122a8c80831b49e0679e74f81a2e18540
z7eeef89f58178f152b74bbac97f4c7a3c9050898dd05ec6e6ccab4f6b73b6c52706b0be1ccc189
zed94fed26c118c68f9ec8693eab231f15cb2b027db896b1cf37653cf71c403bd2abe917d8b738e
zf4cf5116cdb80546ea3f530e61052b2054e6646dbf8b0e1bbb131f300aaa2ac272936af9ba03d7
z0b083b912d5d8e1ad30e417c5c70c9da5728f76373570ffb0b5192d6febf35cb1c2ac610156e81
za1cc041e86e965bda2d6eb84c84d501ed08df8ab2b9b88e067f9f56c0c92b2228d4b971cd49acb
zc1760a57407a0e0847e2cfe3e672831d41668ceb6251f2fdf55a5164bc7632132c9396c8d8310f
zda83c15013ab07dd903af726df6474ce0e46a6248e0ea9bb7772e2816592ff63ab276830cd5200
z2fa059108930ef21ebcbd39015ae5b067e04ab0f5723268f542b53bb480e83fe546fe38d283799
z56a0ae96da6fb4dd6e0f2fccbc402eef9a6b9338a0f3fc6d4ce3407b3b355d3aacb1a35a69194b
z5bc88cc183301feeb4a7cf02184690c00e0a0a0184f97376f5ee2f2575d9e63a739df8a3505d56
zc41aa435778383a005b2aa1848ef33b552b3c01aabe3f6433579c1bb4da1c95446f563f1fb723f
z840496e646e354c2b44f1759d295fcaee5ecdc875c357cc73474ae94e9c4d582aa1a6cc039cfde
z5fc881dab919443c919636a234a5ff4f170682e76f8c28fa21d6b55ba63a02f57573854b2e0845
z7dae40ef1ecff3d74c5c61ca667c32e80446fbb5333bd5780e80e11809b17a3af6d378c5da6151
zfa9c65acd91d3795421803e0c7d6c296d7d68501f1969addc4bd9d19152e9d8a42dd5e73134120
z6f0707b5da519a4a762b22090032aef937e36d3651770a65efa822e198c029ea6a6509017c1541
za6aafb44563dd27c90f86f61e0fdaf164da0c7c071d20d9f719d8d483feaef1123f4b41f50f868
zb964ce5d49bcff0e7a83159e72f8fcfed424fd463b9621fd121c5ee2d77e0204ad02a5530dab20
z9b7ef6c0fdc4d5fbb0f627e5572879371aa231bf2b880b768e553301874433c8d88fe3f923ab51
zd3dd1d423ffadd0f769a7d6c8fd8114e21534c70ab3aaffa489558b5d7a14baf861a1a1a32495d
z04e75189dc1493ce4dddb465665b47a78b6d44bfc03711e139d080f558995ce101d09d1e93bd92
z3157447d18ee114b000342c9a7f9d0ac79323bcb5a83f4d8d17318eda0ee632c11cfb2fd0ee5b1
z3abba98dc411b5b5215bf778f642ddc6130548b4fdc2ca025caf197c1b11523b9ac44227186a7a
z956f4c27cda53e9942511dc714b1fe1a1cfa8eca2ab2cb2a617d091911ca72ddf2c91ec5a8ac90
z27460fd54335e438911d52b8eb90df208848033298959421e89eace3a746f498230225e0987bf5
za914db92199e24c581f5296b8cb6d7336ea996d53d310e04572530da4bda31f277d5c754d35180
zb4ebc82ba8ea304837e71d7f94411cd8263fc313e027f0081475bab8dc98d1020f9cff152b8b5a
zdd9e5c6839097e6c857199733d9d5f4fc3d9042bdae07151e94f4d64746a5d288f14af242e137a
z0d84219ec260be5a73974e9c959655e99ea7a759112767d752e893ed674c88ad58eda3da749856
z6b4a34aaba47beb64372bcd1ae538055080e86a4e7e8c40978b0e30816680973fda521668d8e5a
z3b8b868943423377e483f1e0b7bcb99c3d00dcc6eab8140b26b969394574f70970208785c749ff
ze9a00c0a090a31b14af049bd6e04d520795ab9bd9d8e4642ddea0054e4c55ad73b43f848b8d4d3
z44a75b4e9d3d56eb86a2e0f44ebdf80fd9dcefe2a16a256a714c136f1cdd026dff2535290fe6c8
ze410a8842264a07a97fc4046c5f82685f81a8c1b35e91cb31c5612fbb27d8c4ac87e7cbf5039f3
z40f763111905b05a0a32c9c35a05c59204edc0e144cb3cc86791d43aabd3883c56049d88829b59
zebcae33ab305f5eebe569b8fd02256108de5568522c613e03a7726c8b449e6f1fba01d1fc132a9
z03d82c97cfe548762cd191c723e29188eae53d42806d4b1e2c278d39c15cc55dcbcd59a44db73e
z73ecafbf0af6c5694dd77b5b7823247bafb4955c92ff35ba25b55573e76b99b845f983fa2112c7
z252b2a24316923ce2eb54761d34f4989f0ced1617d0d6fa24ce7c3e776fce7251c4148226eaab2
zfdcc7bddc2462d31d7bfa02c3bb1e5191a8c4b8ce95e4daa36ca6d0a5494fb066f424b165f86cf
z0e354eac9fbcc9e27caab42b58b9dfcca9506aecdb63afda31927e5b91d7646027c831607ce378
z96d2c8b99cae4e83e6a2bd9c53afb06bb628e4df75d57afcfe7aa3b9cca9c354ee85300d882397
zff0d97e0f1a7ce2e33cf0f872fd6ed4539f3521e8d9cbedc85130493b44bb01867898425fc6a89
z7f506e0d5fa53e95d953546b7eaa9e49688c7da858db7ff79e2068c9b54d7d31f6a835f0a6a19f
z77ca46e674e2b00dc6e9bcb409a9c4a34ae62844ba4298047edf68394189aeec0c9fb47e406884
ze7e983b3d4bb34f2f0e282dc448f8f686bb1faeb13a15762d049f0efcd7a9414f3c521e926e683
z5dd6280138abd80fb1c4b5156a9e181a2de95ba7491ab32d63d0b3a92e9c1fb16f4a474a86d99d
z646c7ac1561bbe0261ae3937f866e755b60ff59da6809d3040c8ce34dc5cfc9b6f0c3758fb3de7
z106d12674e252aa28e29c26b7d17e9fae9cc8f1c906fd260621555f7d6df4ca42f870f842c63a5
zfd0b9b3a6031461dc5755c0d36a40368b5bdd5a30a6d898ebf48bc1ba8481c04284b5eb83c6a0a
zdc926f4faeaa9ed67ddabf0806adae7af2d011491afe000114e43f9dc17e90c02aec5854d4bdf5
z995a160374ebeedea5fd90203009c0c860bbb45cf8d49e6fa42f6aa2923359e95d63e3fe480e1c
zaa0531523b4335b2a4b83fbe8b623c64f60b049178f5ddcc469f3ffe861913cab8d527c2b8ce4d
z34f3265ea99b2eedfdfb96a6429e838d40fa15f0792b4c3a88106611ae63d697d09aad6b0334e6
z7be55a004389d7544d2de467374991d338060248d7c560999d623ff4417f6f95bad2666412d66b
z55c1e49040e5721afc9a5696d9eef1f8cd9f4d17e8514c758764053619fce19bba81bea2e6b4c5
za7869d536a46ec37a2ffeeb213f0ea2617c92ccb7090142b656b8a7684ef61f0dce1972d6af5f2
ze82db25e4eae7edbc68abd3d618f384f4f29ee4b54d38ee488d2576b779b18da4b37b841f3d9b7
z1bd95eb774a9634c15511f3518c07356ce34531eae36ad99083bf766295264681f98f9bddad1cc
zeb3dbd11b57e4493d7324d2f99127e7f68be8f5863b01166287dbab54e58438af7ecf6afeef4e7
zac1b620733a777f5b87ed1441b1a532db9096557ccd67dca931b406afaed50b83b962d5c658005
z78798a1afacae5ffacaeba25d9e5a6e84de4d16d2e7f35c68fe0019dcadffb06df1b4bf7a6ecde
z95b4257158d429837e3f773cad71de24184729c8c788a0d5db6fb42a6fac85a12013cd4e1f0d0c
zba483c2f50dd25ef9832eabefa330b845e7d225ecb5feef5e0ef94704ae5d02ed38fb29a0c9d1b
za25da68497bdf6953b06b9b10d76acf4626ef4240554e2e3fda78a03b733d966e63d92ee6e6be3
z01f64b7c4b1ab1958b6c154f7b257745b35eacd4c32b76e5bb4458b985bf1cd1d88ff967f4d54d
z1f1e44956aa86cb1d373c058a00bd0513d10faa7a87f574abd2c37bba67aef4803885aed9aa318
zef5e8651617e1dc2cb2dc08825989ec1a38827ae20d111669867e9be2043403b8dce64671e49d2
z1bf888348b046d29e8775dc2badf85c638ca773ad134136d2f248710f74a135176817d00f1d45c
z413c866098306ba332547bf9d8f2aa1ef8885f1258e622a80f00b6c84a80754bc41f64b68b2c9b
z9ae8b6d8088b1c4e524fdad08983e00206cb7ef73ba1d9958e376ac28672916c21b37283aebed3
z4f79b28d744cc5a58ec3715147fa7e66f666b83f39d17da7c999cd230eda5f8cc355bb3d669a4c
z898a53d460bae30929a8be40a2575c949efec183580759b5df67c0714a284805b6c4ec0d98d1b7
z50c29a86399db4b54418908192938285afb3e918f4ce57f12eb8aa8d42b912eb5b7c39f03e99fb
z216d4dffc066e5054d6493c65b6e2770618a0499a16692eba897a6ea0eed568fd05786faace549
ze377863521bf5f0d45b6639d7da431df8c20408613b49cf3d933893a4b38e8df9f2107f34a791c
z6cbe449e02ca33ee11257c9cde5c547dff20d3d1489eac9bb9cd01da2c76fa6aea1789fc3c5286
zdc9070c59c9f19f527ae6edb7d9e144251be5adac17d856d8d9d80c71572368fc165b37d730a57
z8bd91f43da55605971150a1f8d0de2ede74345d401baaf889c793ed6161beb322ae13ebae77d63
z029febe5b9ae6187d7b46357e52614dcf657a39d085a5a845323f5932e1603f6b0c377c0d86e14
z2e2788580f686597c09add689f540c685c1bcac212059e5836898c91ed718bfcf05cd40d2e84f4
z3f1522d01a1cfbf7f400bbe16ef4b7544a24a28e2e1c3c0bc26f46d84a2f28da5c2a624642354e
zcc4b0ff08762c0e3a05b1f0815c07bab1c479367c4f2349bb3c4ac1455b441a8e0da02fd2e5af5
z816b215c6518c2984866a5f1f10c6b2ba307412d47c1c05a335377af051dcf9036ab14aa847191
z4a9987843be938fc9175c5079669ef337c437347af5f71c5c0f8c425753217bf52bac826a9cb41
z19516fef305c486cc24a22f1e9ce500ed641e4a7d75b0e613c4057f460140a413dc07a1d971a54
z07437a92db231627655d740b165ceab319c94350d3d0099d84a09ca6a93e995d3c9550bfc0329a
zabf4bcd5201c4074a2295484a48f51aad61647944c2fb19a03c006028cb539aa49a211edb45477
z830d5a659518e6c86d049ce9e3165167d99005dc9fb242b065fdfdd7dcfe0d50bf7bdf8cd9d9ed
zb7b890fc0071789ce1fc3f9dd74f81eb923d06b8038780f706ad8fb88069f80f09219759ecedd5
z945019777cc57f92c47a9e2c2060385c5d3cbbe8a5f68316ee5d4177fc77b6141273723ca8eb02
z50f0f0bcfdd5a69a065146c3367114e3f89e0a0a56ae80d453402c438f55e3e8e6a3822164cd98
zabc9e5ab77fe3bf2dc72c62d8b9097ed7a994afb4768ede49f07f8d64ad58f484a61b2bcbecfce
z7c13ebc3bc68eebe92d3b0c57e7ec9d5a61c86bcf4a41b81a06fa7479f8b5badc686d99a547916
z84fbd629f66eab6c0271e6ce9d9897773b9e25aa50496555b62d1b9ec57f19d312a41d2fac13e9
zfde3ca2f9c103e441b1625aeca7f81d30be1281c98a0634171af9867e14990c174ebab5864c676
z0cfa9a697203321611cc142a880dc95448b0990fb83cc8b433dae608027c40a3f03bc95b802ef6
z482eb934eb267c15555ec3b3c922c3afa51ebeb66c4aa81144201a2e53979333b8decf66d04d5b
z2c5960c074560fefbcbd91aae7c080a4b6bd91215f7440b1ee6b8b77d14340b31322cab0119570
z777a298227bdc3c4362136e58ce0f9f4fe0229bb398a1ea28aee8f514d338c4d833f0ff2aa1d41
zfce7e329694074f2df4b8b58955e99b1ebdb4c98c97d69e82102250846c4d0a4871a415496f293
zbe4e6264e078f1e5577a7ad7fd54c151858006351fa102b602cdc063f3671d6a13e7d2b9a427bc
zbe8b71e22202b3ca7873af38db289a70c05188ed6d315747ae44e412bee82a7ae997fe53b222b4
z5c5a8b7349d2a06d52383a9cb48f3b88bb56025aaf104ede367bc15c7d5a119dc6d47bb6defb82
zecd75914b394138c8143d5d09536f008979f04db479abbe07cc13ecf651b2c125b22760d5bce5a
ze7b895be11b5610f9e24c0c9ba46f99cd0cdf891e6d56b69459fe0550e6bd629c2e51c4477f2d0
z5f9ca52a347cafe979fddecdb4f6c7b2d3eac92395832827297f59217008813b7fb536eef6c472
z8bc7b35df58823cc4b195aeaa81a6df9a48f93af84c940f4a71f82ff5939362038370b18cf8d41
zaf0bc25390bdfe5f742cf9c848b86c3d21809ae45315bda760617f702b233d4a90e9bf42ad123c
z08c997fe01e2aaf697e413c4306711b9644223330d9505ca035e8943afdd53ef72b02282f65ddf
z250b905e409d60cf05d8c00be6852224914b68900e9e93eff210edd1c8e54924244597988d7980
z0a398fbc84f966c57331f0e43c67a4c6f91a84f61dc231536fa44cbd6ca39f007b430816a2c685
zb814edd7f887fc76c8926800770c136ab40b36a6b218452c1a2735f9e7683357b65ae4cdc424a6
z3bc8b0e1a3a775adaf2d92d036ba8200425ab72b00a65e4f1ae4864d32ae3a13022f4b5c73d3b6
z43197f8fbb27e7c730652e0a5b993c55c7108efb457154c91498055bcfa53cb8588d3567547121
z867a49780d26ed1fb9ba37b94d19fccb5472ae9dc19bc21ce208545ba1bf76ada9bb3e8ed003a3
z11a03c8ea093648b4906e9514649c41dedc826a9e3ad12e37f2b11948e9727a4b60f30ec3bfda5
z85455ab769fb3c220c3969c278b1d3858b36ca143e08d18a42e7d9205cfd619f6e74c1804557e1
z5f9f299da6885c6ac19c34ca8c9ef0253f412f2b86e4d539b97c2c0367ff2a3dfded9b54047e34
zadd40e5ab0520645f5b7ce9b0bb28626e78584f4917a35a11edb210384342aad4ad2bd79010e6e
zb3c7b724380ab06ab23cf34cd02d3c3e6b44a9f35fecc1b77ea42a3ddf21acb2002078e7c90984
z8b9ef952958a2056fd3b1bd38b5bab8acfc921468b49e2117731f4500c0b096f241917d1459661
z1be6d505c4c0d84e2cea5cc1f847cdc61ef718b5d89fd105e6f0c657062a24859bb8275714bc73
z5a0d273409712d103f933b613e7938a81cb18b91b71de628a1ce60b56532e10405ff125dc8ed2a
zc8a657156d01734af8e0bcd23c9e6319b03f2c6fa10fbc3f09439230044add3efb0eda894d2a94
z6ffa444a6b85f53947c3e3745a5efe0ded59562c1db48f8c609c999fba1265f0d61865abb67efb
za77bafee195f2e5fae452dd087a820d64c140911451b2ba6f7808ef45d306ebdd591d5c02c45b2
z306c8672ca8988814ca56f4656fc3b83346ced6394aa640e2bb579e0159f8bd552ae919429910c
z4e56f33474916f628b0ffd8f4744d1b57994e31de1420818af378f770c0d8443be0de40a2088f4
z380f5186779e72e41bf0b9d67e6c80a776837d90530a7d9e24d5982f27b3fd96c3f612916bfcd7
z28bc4f43d978314cc9cdb9c254fc7b4c88bda83ddd207358eb456cbac9640d44a9e7a39e5e4043
z410ae32430c49cf8d9bc7adaffd320557688e272a5d07301daee6ae0d11fa92a5f8057fc48a2a5
z8c28701e45a6479ab7aee76f550669ec8390656293f6327882931d7007c7d9b3b7a6f84aaffc3a
z90939054330da75cedd68a027c9192f63e180532f2fd6e7989aabe93268ca9b1aceac57601433f
z0a887d31d0ac9853cd00e4f1502756d5547af852cef11c3c255b3e0065fcfcf874d8445b302755
z21984ddeef70777c115db4345d86d9eda4800c0ce41d5ce30cad7850fdd7e4b6084ecea374bbee
z3562b733eb6b1bec7d9266c2bec823e31a0f4db27586c3a3a7c402c9ec6fe3e44258e0fa4d40b2
zaa8ecf4570d97e92fde21a58adb6b6fbce23ff8cb7e0034342be7d9d1fb8181ba4290378e75207
z59e3bd1b1ef18c635fc3df6d0afc73bc235e40dacb7a0c530e173470c9f6543d3c97411a76b0d8
z22b22a49eae43f6b76f58d8f46096c4ef560834c53d9071f0ec2c7fbad233c4d5dd1efaa65a8b7
z9a06f4eebba9c7ee8f320c561c9d36ec3e9b84fbf7f1798b89355dd352455db5fa176f8a9bd227
z13fb2be132ce4cc1e0be535051e8061024ced2f4e14b5a3f51ebd4e397267a47c5a7b5ad0cb232
z0b8681fcbadfea4e27089ffb409a5c53f1608be32b2d6f6b9649ecc957f0e9de0e455a80da6553
zd5bbff7108bb66a63f1cd16465b50da705dd72809c38c895b9e144d7583b35932d6c6f045ff92d
z46bbea6035e1b60543570f9a48b2ec2598a3b764c839bdc316eadcb60fc47da30264c690ff2f4f
z57c21d6f6e8944b25cd30db5f8c88a9509cc1461f3d3ad760d6827ae43c39f4d69021ba2f65434
z312ae8279fe15ff9c580bd4793cc0ff597e218a1b1f4d33cc2a1826ed53c41a1b9e79d30a7d7b4
z6974d758a7f8d951c2669724e3515dbd63813aa30e7d102d5b707397a1c661ea430c90faa4dc6a
z7fe00e7ba82ce210ce24ece727b1c5556bd8b4edcf89efdf64dfcbb906cd48d200d19691e23184
zfbe02bd6a713863ddd0215892a1f692ea5bcaa9bbab3b08f855cb96d306a6b86fabb67909f6d7a
z5bbd03c9245014ec181d886208482fa04a54ca051c1267db7f48a8a9439deec523774b133d0844
zecda5d19b162e8793346f245f7808928ae4983a27b77653df05108f9dd0b40e1fe84250bb72163
z9f70de3d04ad8ebc61348af801446e795163e0be5a37aa8eba3968f4dd6fd79fbc4b2625200180
zed13b50fdbb604b204db45588e41eaca5f54c2009aea5316b5911bb62cd1d845f50e8179456d18
zd7bd64341e9d2291fe8392d9ab8448b5f3b4ca6877bd7766a919735f353bc73f8cedfce258d8ad
z99230c597e3a4b14310852c07ce1ba90192fcb15049cfa7a57d36d7e40910d58258e417ebabfd4
zf1c14df86b3f8e03dc55365f0950973fbeb5914f28471001c8df3fcbe5c964cfc10a04d0498bbf
z11a7a3085f5c7e40749297ddb9e377e3a8c7685cb8cc14d3fd0e88b8744c70756ddcca01274372
z918b818c2b4709ba8e261774a8beefb70fe56ac5b2bbe36860b75edba3242437e88b6de4684aa5
z4f8aa8585b43cfdbf4405d1b069e72b1938e9ce6af4b89be1a918795f417c7448dd90ae580a8e0
zff628aaf05b4ca575f25620c2c25c35e02a836536946cdf45128edab486ea7122ba0a648a8ee91
z7eb9d7687c2274ebf93a2f026b00b7f3808ad2fe2a462fdb89a9a0332738f144d38f5dfc419185
z28f49d3eb1bc4a6bd0012ef2d38118752bf25340241434c8d90eb32d5443916a33c71a2c70e562
zee132b506de357bbbde8bdc9e5b78c2ec1daaf5387c4f99098262836bfce7795fc72a835f0e4ac
z2f9cdc865eb788fa004afba7b1a42368ebb4eb808347ff5829d73e268a3dfe3773abbe9a364469
zad7d725a8396cbc2b96f33da3b00b26170e13b418fd8633025b46e60126246c18b9cefc2178ded
z6190caea71d8f8e3e159757855168474e426e4e8a7218d38794d833cdcb5c8c221ef9714d91ccb
z5fa6c8309b658882d3e3c71cfe3b19406d92ee1736f6423c079ebccfd35d83c30763ba54fbbd2b
z718ea83da42dd9c47e15c6d381e87618719f0038b4390984024788425cd7a48cb33cddd73644dc
zb773988419d021a1bbe7bef865334b953f3437ab93ea76ed12ce65c0ac1b9b393b9ac8c66850ed
z40af468db6b548942bb359c7755fee7d20b19e2a4e82dc4a7273619c94b49be532e10f6a37be06
za7657e84d392e7eb2d58091a6f1e7433580d116c8940ec68bbde672577cef60e6210f397ff13a7
z0d8fa8cb0ebf61a5b3556fef328ae6b2a386f780069a08d808ae72f762ac78cbebb02db9308789
z488ff0d7682fd89888d69044ca8c832ee1c8bcbd7959961d0cba0107552065137d8a6ef9957d55
z3a88b91ed25015b59bb4a17f8e609aaa5e8389ad1a88d3a7e2550837ef6c9270c58f88a030e6fb
z7bd86b7826e36b317b412b6735ac20350b495b70220464e056b244a51259873e21d161da9fa75c
z29d640087ca4ead8a4187592616aac8c4b792ec56851d7468b56f330848eca88f93e08ff737404
zad09e80bd6a11ec43c2cff07c2357522932a59c51d3267b641a9e8746387c1975e8b2cf079117e
z901b8509b540f532e709c8bf668c0503227d6f13ba24af3bddfaa1e563756f4d04158b12bb15ab
z592932a7e70604cdd99b2dbb6a3d957ae0c1af90ea78b447238333e2780f16c71ed4d4de27b403
z55e5fae391bba5575ee71fdba67cdd47d87db8bfeced98765540709e3cf7eeeed83c24a3e3b3a8
z1a5ca9bd3e26ff6ce9a4bf5e3dc997e65f29950b51683c3c6c1529a5818b7dea05745962e89927
z72ffbb303d961170f2e6a53ed608f9f9dfe25a4c0d9df205cda46a6caf81c7038ac08b7f9635fc
z4239070463b2b7e2f70e8fe9149625e9e7a9e4b1858247e6ccf267652029748fc6ef4f7036a84b
z66a3d5472f2815d7d74b9127caf36aa4ba28b71a4d40ce26c1e5ff9e218787b7640c8f26543fe1
z1df3a1956af17a568e3295f92e3dac9b9b7efa7324e04efe7c2bac7313a6ea688d46653b4b7d47
z62f62e4e9c4adcd628df6c4ad9c95f65cd835a847b4f8d5d6747841a683474fb3923a59f560915
z563f54de62bb3a9cacdaa706148b4389bf0c919b7e02eb77b0624fc7bcd06d564ab07651fcc11c
z3a95b1fe52aa2ec221d5ea17ba8c4b9327c354c8768abc965b0eb3b5002201f04a56d94b0b6448
z523f934293ea34c92d82b59cf92513dca0087506caff898a4e197e75515aabb1d1066b041d601e
zf04eeb48e3da25779eed09eb26ea98d6c56b6bc8bb79f1d7ae843b57ee2458f34d4798c4b1ee51
z97645a259e0be013377077f5a2bbd3d4bd0a064d4d1cd931e0882184fb7a8822f6ace37a0c1a16
z136f354ec09ea16f57a613d03ba07c2df795a8e24946697a268769831b1fe040cd0f702ec0dc36
z684721a105071fb7c4b5144dc1debc647abe5c9be8bffaca14faf9089b44a2cfae2571da577c9d
z7818e0645f90b99d5f3de1d60cd78e09a59dbcfe9a148553e153d0f2ebe1d9be4e4d8b1bc47bcb
z8a786b303f09a48b4459378a5d2fb1c323263ec6331412eb20eeb45e2a5e552369c9bf9d64cb33
zab9c77424d19c6ea7e3ad62d2dc1a2efa60a8324895178c16f68035a2689c438b9e0a1af55de8a
zb9682ba16f0a903f42d94f81d699ac2544b0f99176eadd85bc7f31180c606c4e8bb2fe99c82023
z80fe7c132e2dc7745936c4c8f762c9687939368ed1c8c6aff361749aba5e6dab0daec80f440874
z648c3cb0a5ba5642f563dc369e35de4c11403b89545187c928093abe4b420a6706a522a62f4139
z5b2cd374e97033d8238c9bd78c93873f8e1c238e1192ead5e2a87b04b1abb4b79acda2d211250b
z0566b3fc1175d212270628292771b4d17d015da1e44a902be08bd8ff316448ad498526b0295c22
z747b15a916c52ef3ceec9e882a32ae69c4e7d662e373c87ac14231747e807e4f22684bd29f55f5
z6f569357bcf8792bbc66559e40fa86692b147b364a742dea35fc6423bb14745dd713c948fcc188
z28fb891b1f24044715316cfde24b0610be5d0fa7c0bf8fa056ffebbf1e487127265e81777adebb
z923269ead1e0a17fc1cbcb9b4b2333680fb54ccb0d938eb93500a066208b27d083bd93d7d9d1e7
z9237f446ee144976575ff33546a7bcb116058e6c86d092247a886329b2050952e8fc4a710fc9bf
zb8c56dcc81eb22e0b85ed8fbd142368c0941a4ccf1210d816d8f1be39dcafb642bdf7a4f0724d9
zf5cb148f18911159da03a62ad9cf439ee39120bf70806edd31bdded70257f53d0017a016a44174
z8ebf4d8d282882b7442a6d12e984f4c8e21a88223fb23f9e549bb88715c4f75a461c7a935d89fb
z2928252101a5ffcece11bc464a9265af2d21ebd388e02b320527ce02f4dfa98e560e39206be4c3
z0b4da26335006674aaee89754672d42b1510e4a9b7418dcf1e3f77834cded615782687c0d33487
zb1b5cb8199307d6a45bee6f1b67c50c6d9b074ca4ec80cbf3bf7abc9fad99bfc03b94ad2007b10
z8aa3b00ee22ce09e78eb29382b8cd6b226d91fe02e877ba05418fbc4b7998b37847cb10d803c94
z41c03972a82e472d37a76c800ba8cd954ee30c98a554d2c509ae500978f2d6326823b54dbf1631
z5a896b30d0b5a22f4e74e8bd2fb4f1b73d48724c0b750cc2848b1bac6c459befa99b20351d8d9e
z11cdb86278c976709a5248bb6b72e9b16b0f2d4046c0e5189bd1817c1bdb3ea87ef7ff05c325f3
za8465fc47587be8f3eb5249bf308a642d06aff7c321d0aab3beb9a4ef6f8eabfd33d1dc4acce7f
z0c412f0d53747225d8ebc978405137a298ff76300e75a8402a17ac7a6f5de3b386fd32be2aff3d
za4a586a23a9d57d1f46b7b0483061e1d0de1fc639213a5d1b6860a26cf3615c159170414bd7904
z4ece36b1fc79589ab0b97ea44bf3aafa71fdb91da207dae863f1eff5533f53cc98aa4988b743c1
z55194a993f1b5792c251793af87ed3c9597c8a4dc21fd45a9d83e9016c0d1418e3e1e34900f48c
z63ff7291630a05562e80b41192f656ab5418f0fd1a9ea3a54af2b44c1bcaac2fb5d05cee265dbf
zb17dad4ba00529d7e7cbb11e8bc23f6a4a912bf7effe367fdb107e80e64ff5ba565bb7357454d3
z0f4ce17d642e45e1c811a6baf0375fe854da07f8a080c4a75769169eae6f7f184327bac147987f
z36d1bdf83b9b49b36456a7c388de87b36c4c4da0d794accbc55d3aa400dc54642a64c26370badc
z03c8a4678f3c4c4def7de5c68ee5a4b95b69fdc756885cf58e7872481e7c0a8c3eef8f7db3bea1
z3313d8257490a58edaceee130610d223ddde0d1e011c3c8f82da1ff32f11dfd10dc23cb4811c9c
zb2cf888c4d0968e65e929b37955f82765f185ce04e4626cb552412019e01d8371ee3d55f1cd74c
z262a2726433b9931609efef544a9b1f9e811322c6cb8417ecffecb4b0ee2d8b0d3e733025e17c3
z8240a13374448bf7a459cb4c07a6b97632497d198f9b26db360239e94fa4c58831f1256b93f1aa
z2a4993d3abf78ed625e7b71e55ac2e0e7a33e38b822df5c4e186af13f7ff3441f4af7645c26a6c
z9f7f7373510b3f53c5cb4034382403d8272727c2c51ff0958d5f59b4ff7d8cae0d16b7b0801232
z5fcad77da11563e65fa30da2b0a81ca041b72640dd7e99bd18019f051aae5ccd69f37f5abc1f38
z70341ebac820465fcab641a6dd92da4e6a58bce40cbc24830a58170c444cb38773cbeeab4e620f
z219ee72a12beaa03745d43cc89f160f7ae1a3e4bbd78384c84a10afbb601aac54ec8a527b4bd4c
ze1c0e8543c6d256782d467e71be6b30882bda68f616ba2e4fa9a12931e4d285575cfa5d1170b53
za9fa325e8cc8f5eb6a73c9c719d9c6c92a2822896cd297741ba284aa84f66a140e30f8acb51451
z167d242b1967ab554677ae2ba8fb798107b7a25c79a257337293e54f262435026b84c8cc309562
za8397c0fa3f25c577ddb059c30b859980f3e35d2d28d0d2a2422e014e4fcfd345392c6038dfded
z4e21393d859de9dfb7eec673003e08f5d39765c308e92e2ec09b533f2e6b2bfc2659499e8851af
z815581fd3c7e9f1cb85037f3a71db2047bd56aa5de4b2842a240bb611d5f7fa0e82c98889b926b
za7faa45b14da98b677060338c6b86d2cf6335632afc1df1e344c6559bf1c367f04c340ac8a246d
zee9e043b8d0e3ab24a04e00884ce8991a500e1dfa6cc08d1ebeb78002dbb24a0f48f03d6c74ddb
z44d23c0fe8088c58b40b57dea70fae9f36fb9ed0d5b6522badd1e518f3582672867a22a05acdf5
z4da8a0308465eeb2633667ebb267065f3635971516cad21fd14f75c8ddf2c4942c819e7d2e656f
ze8f8f91eff36a16c4877e1ebbb32f1f1ddf0954aaf38021e5c8486b117a0861c486d6b529cf99f
zf3a3353e0f8b08f606f5be5a7a726b8f3fd2de4a4dcf265eb65c58f812954778af8fe3058eef6b
zfa0d2b8891acc194f53c4c13eb8a414107003645ca4aeec5de385d2fbf41657640ce3cadad1205
za3e1e07618f7b96b43ff7fd5ee63b78770ddb0dc6f25fd26f8d1e47c5f417d93118b19d497510d
ze8e879cd51d55d713253f61943414f695ce84cff349ad969d31b25c120ec95c042dc815d48265b
z4091784491ca00477c4b78d0560d185f9c734869a9922113b57afb7d3745da4d0623dca7a3d1e3
z9fe23dbe3d48a7b53ff6361a2dc53d39f799fff177044925993bfb1cb44d20a952c9f15f2f77ed
z9d5addea1479f62a88d33d9c8f6229e4587ba92f5171c36241b354c341986b4bdcf3ce11d8ceaa
z43e0e302634531b1027c7995b82ecd0773e7df3dc0202c9f100076fd213eb72647dd5c1f1a1fe8
z37efd092f36158b316867167daceb73de7499f199ec6549f4d652d965366360ae065f2e49a977e
z532d26475e415a60ee33dc34db1609fd32de55ed59a2b30ec379cf44b46e35adba155c4a2b742f
ze8e63663549693ec1b52563570ec4517867e21b6ebf75b900f0499ce4c44ca316b03a577282d75
z1aee9b997eb8a2dabac79a65ad8555295bde34122006399bb6704483a54efc1f4a2b5c085fecd5
zaa0c36fc61e48acf7e8123e5b930b7a4389846d78340e8b9e6d5efdadfcf729d5b40054f844590
zbf497d33a6fef50a8e5d03b17777d9ebdd0cfacfdc5f27fd6540da9f9fddf73e7ae622eabdd920
z20ce42a0eaa8ed5e8cbabebbc38c1898e0f6bf3f65bdee8a8151efefbf4019b516e6f5cd182c38
zee0319089a9e79e168aaeada7866dcba6c6ad7e649f139ce401e534d90ad2164709ca1041022dd
z3c8ea44df5f98dff07faea3d03f891b7e6f7ced957a3639eeeddd2daebda88b234b65943c71b09
zaf2c5748284c5fac01a67cdf2934ad942617d81fcf53d722c1a73eeac76c47e95b84f8db080ffc
z47d32783008e553f1f0295d0eede2f9459b4eaa66291bf291a5d88f6d8b78f8cea23e11c8b08cd
z2420b53fb12a55bb8d5484cd6f0dbde56c45f4e2c9ee9f4fa73c66b3db90c207b84424a4081d91
zd8037e6587cc5d87aa161e0f72ea7a2f68451b5414d0a9932277aeb585f00a3a1e738141893852
z7e126cc7c8ac0ceaf79ef7adf61378388faceea06a1f7737720851f58e02a401e4c1ae56b3e0d8
z3ea803ee5c392d41cccad20cc133a62685c437bfe376277b37b08f99472c33f52863fb7a70280b
ze9378aad6748c35b0f21cfaa329b7340fd5aeb725126725e8493fcb10f56711a7f0b8bb723cee2
z3fb85ec362b5d6670c88322cb89839aa0c2deff6b5249b9b544eb84d16747d0edfb64ddfda657f
z09d62b27e1ddb69c1f6b88d608fad5519015b2cd24b158355b625a7afa38be632529a705f14d8f
z20f8c7b9b470b8be8f45edbf3bf6b6b4d0f1dcf5fd8074a0a6d04693d6b3bc466f78996f2fe828
z586c776acedb4c67fd84898e93800780896da724ca9c581d7de3e560cc7efd2e9711c9a0d68df2
zd4b62fc796f20e2bfbc3794cff7e1a8f0105e7231d054073f7a68a504b460a0492d1d51bc1d201
z33d0d6de9645afc66d38414cf902486c5f17efbf5ddb3b66a32e930c9563da46697a3e41822527
z9a52d471978622b06e73624dedce04cdb7aa7cba643a2e357031e0476328c340a08f6ec38f84d8
za5c6fa455faee509571692dce569a02c60c7fd331133b6ed9727dbc4416d3b59b4c7cbef3ccea8
z4ad61eae9ec740a1dc7612949173598e2e85526c924f4648e8bb13441cc00b8c332a881d7d2496
z90f48ce72517d86911eb5fc362e3dd7fe187aca9f80cc93da8d68710554e3dafec6136a9015ff6
z869dd769627b2fe68f966abb4b9f7e41fc2b3172a72e61f070c17d1b883f9754389ace5eac5ce9
z9eb0c356d686fc14bf1894f7b6ad19bed5d2f1e9f73559811add2bc9e8e3bce26784bcb53ddb8e
z329b27351cdbac3a6992f6a779b0fffac50defd5c362c01c2ada808818ed12c05e875c37dcdd1f
z0be68a2062ecc8d3efaacff220e2344d7ee5c7b39997bf829093b057ce9f4b5d7817239810f570
zb1fbf64b69e8dc2f34b0b43e7cd9451701f950e6eab137a25cf1280b595ce6d232b57009757ff5
z521bd77508c18b55926801e1ea414ad5cc95e30319f43c37dac53a5ee632a5fa3f0390937c20da
zc18becf0a83c83d3730ebe7d789661856f8ba5ed7b28fdab8eb2c235aabf5d70ffde0d0faf7e08
z0217fa153cca9ececb8251149aea9e7f38c4c20e526b6e7947accaa30fcdc4aeeba3d80ee94e6c
zc29b693fe757048460f7959ffcaced14344e3f3bee4e4ce4bf1e50bbb7fd05928e80acb8eb857a
za3b3c2dd835790d7a76b10a599e2cd88b9622627a48ff482bf5b4d58ef0f1bf17789e2e5ce139f
z85c93bc686131ef2d343585b271d7a729c2871f9ac023da7b1dde3a40f4e1ca6e3108ed6177aef
z2d16188665e02b112ce3b20f87898044da688451586960308d34ae2719b8c9e98d7e6814c5af75
z716e2cf72fd514bae0adf7d06b41ac3c038b50a964682b64db1b40520f4bc6892f9dd1390c8424
zc75ea5686b02c7b2b60af897f9b9cd5843e6972ce39a6bceddaada197e283c1f16ef93a115b094
za30e59ffaa9577e5c03d3d1830dadaf4a5927a25ad2a7894a3ed57bce2002640e43bde3a96a4f3
zfcd2ee05cda10907f9275721bddafed808d700d6cd9cdd019392fd3d2804ebdd6ecd0fa4028a21
z3f067b177e0f4e5b7edd894dfcac8226df43e421aa85f50ce1dc2f3aa4acd318ffbb7aeb7d787c
z799cd96724d859de9c4cc402de7163b66a7612550467266c2dc9b835ac071a094524ee87d3859f
z1243cfc3b4d3380043f056b46eff47c5fe721d43de1a7725986b844ac40bcc90ebed6a6d5049f2
z8f06adadab8f3d6ea37b12487132e42596dbad3bb27fd9140015d57a49f5825dbcc6e09d610f05
z8124e2de90a829acd8d0bf4cd4cd709aa812394298e3a3bea9cda571c774edde55a25616a919a3
zb4da857895432414fbd05f2041bda62b32fb7e117f9ba4dc66db50665f632684a493d7e1949c6a
zff6a5a7f41cf1b27019a73b729161196afe170da0b471c6792e9da51b336e0639b452192d334bc
z1f5939f8c54b1a1ec9aeff2e2df7ae827dde49a0c36249656ee07b43523ecc6aa908755b68d004
zc112a8f606283e3705787cd24b8aba63c03e92915eecc90a8c8dd86bf38d03137849a65606b9f7
z2c67f31977cbebd07e420d6befdca42017ebe9c853b5a0c3c19b40c9ae954bb95332777b3c86b6
z8bc02cfbd43fd37919839dad2fa27695e261057c1e07744d6d42056a62ad5601f1fefe84febac6
zc3f09ae8152a00a1898443c3ac3854ccc35d20bc9aa034d46d86b83d35a82b2672d78eb2ada005
z2a21a3da9606e6e30d578f04eefc76ea71f3c4125086e76ee5626cdfcc946043fde9ae77d6b1a6
zb843194ec3746dfe7bf82b1fa91ccc4925effa0d729d78548ea93cb7e17106122755db413c771e
zbfe19f5abcab2f868e6856e1bc333d3695c67fee9f196b65594ae47e50b37729a7c5950750ad13
z8402e3275e24b532181651112b1053cce59082f9b245ea10eeca2ef0d61c730ec953afb9f67bb0
zf2b225d8739619f60114722254b6848ac7f1fae24c385a36a36911e57bc424c7fe21b124dae4d9
z03f14b986b8dd7c00db5278201b8e454815f34a2fbd0c22c6ac8bd074850eb64e8e391c3709944
zcd53a0c99ac4f86c8a6ee1671d42de6c15e18aac682d6bdd80cd2fd02b118a8e89c477d5ab660e
zc2f152de403a7944c90603a4f97881de78c0cdecaec11456e739b30d30fb9d31a78b226ad593c6
za1f9889a58abdd9de41df5175ae608fbf8f62c1fb9f2323bbfd3d35d631f381015f4751c0dc992
ze25db36f970ad5d9feccdac322bece55879a5a657c88e30c3af266ee203daf8b8d07c40f76a2db
z76d4df9fc3427bd424d6b00e7795e2e37e1760b6cfb906f1f1768f83100519240f4fc8e0f30ca4
zd335409ce5ea111fe8a84c1e6aba6300d2c42d5a885b3120e19ab1225bc4787237d59b23557482
zacc9d9656c74e322b3a566b31b8d7d1d047269c9e9067c4d10d2c8bf2dff959545782ae668b4dc
z5f757cd565b389e8b0fd3531ec8ac8cd76df1aa0a5ffb261bd85649a94ebe2ce30c4a1f8c60920
z8b61afc61066c693d550ca0d874ddcde1e496fb9dbfe9d582898740ed4e082bbc430a1a9553170
zc8bcd6000da280a4d8920359eece2cf427fbce5266e9664b2fd14eda61defa29a6c116bbb60db9
zae12f383f029b132de9063e5f6d37fe90d42100d331cf92d9af67872d4668f7c4e0f44eb000a4f
zedcfefb603b6394f3d743be84cc5d0264132d8f5dc34e2463b19a6fccdc7b045a39c0064d7b848
z2e18a3a11841b1557afc12b1df74bca156d04cbffa3a9684338c619d84775d9ee1c896f178c435
z8c49975e7eec32346706bc1dfbbf2da4471463ce13c3534b0c7b614b69ec0f509c8c954886f200
zc5366fbb9b2152d0892b22c399abd359ec286125f74699429ed3bbbdcde608141f9663c7e5a502
z7a3ff31fd6e321d6fdee525b77c58735cc3d20109ef54991cc0fe5b6a86c19643ec339774d3ed5
zc89c733b20604adf7f7e8997006975d2f40aa0cb9fd0903ee4bbbad7f58c4923d545f9a0260163
z8b30d25f71d4a4af382fa4c5f4d72c891fefa3740590f5349b74d892d68682044edae9e60e5bf1
zd106d44b76a7b39bf089f9bb2ab44455561216cbbdd85f3c9c8953d2da1ba7e17ccc471f75c97b
zc93f6f0320ab67b05464c4f61e14d1e5a66ebbc5b714c9205f7bf24fbae1f1c214c80c942853e0
z658867b169aea3967fa17a49e60a1cf357b995c2c1803da75bcfd6db88dea6c5b67aa86b732c31
z22f5850b685ac97023732aed20b9c56d2740a49b40f430fe95ee9cb99a0dfbba73b6d965219bb7
z20bfb13801a369c71a7335c26d728ae394fff68e234cf66ae032a16c7e42b224c955210ffe590e
z02b68e3ccaa07ecd0aadf94f5eb9d1fcb419040877ba224cb0d18ef4b378f6def9da0efc4e10d3
z480b45095bd28536aaf80acedf49bb383e36bbe1d8864d357a5cbbe7d1641dd1aa418e54b8bcdc
z95f9ab0ebe79cdef4961b69ef6f06c2bbe6b52d60795b80a4eb0d5efaa699587fa35c1b68c4043
zcc4b16f5b1af4a9d6c80407c5406e8c39baf02e543d2a9f030d114d0f4697d6029e6207b8315f1
z4e7f6e50183a4a7341ab9ef93a063df4d3c441806edd4032d16e430be0586094f55b4746d816d8
z55e55466b8c0a6d677654f68b6ddd615513dea8d7d305c62208a4b6c777261960c9896083d7699
z74f21ff8dedfbb1643725431d37e922fd68074ece5aca4d74be386a4e886a08e1cd55cd952d6b9
zda8fb39eea9782691ad6e1c370129dc4c30782788dfcae2041f00abd6fb59ad77315678153acb7
za339c55c1c180d9bdeb2d0693f4221ba4d219e2f9e064afd3046379f46adc916d6c0dd51d4c173
z8c7eec2c3d0d069cccc69a524df53bef955d0cf22a25e520b9c8509da0b918ced194708bf4928b
z00e3cb6ddc423e16f5d46f27cf55b4606f0fde3eda2d917085b6720c4504c69d71843931a57d6c
zbe5618c35af6c0c1cbc9f38a453cab112b6139cbad00ec185b356e2159c66d60f6f1c2c9142d2e
z427b77acea7f7400be2c82ee3d987a6cb015fffe5f23bc0741c91def7018fab98cda0cd01f4ddc
z256a47a671369545aa78add23270627cc596e66070371ce7a76270f32285c3be15f98704ef6692
zafcb979fd77c98b188a5fc9fed03d4a3458c774d940868e6ca6c7037d99273e5ea86a3b6fcba3e
z3a393b1c03747ac15b0218ded298b4c34ba4508f93e573fa84047ef3da33d37a367af84a7605d7
z71ba28093263b2aa58eb5adf05e737eaebb28cfb1f23b162b0e1573667ff295eab8054f74ef861
z4d2ef618be02e995dd32f7493ebe0914ddbd7358e3f2b29f1e7a36006816032b39ec9f854179f5
z3028772159301761e1c052d13ac22be0a5d51e4f41270c2b97adffacdb4338f2a6916baee94bec
zb768a06a45bd27adf304207a11c707a31278a79364f674420c7b30b84d2a132cdce74e094f953c
zf147c61aa86f6da844d678bfc32297aa3b8da431575dc0147abbaed9820cd7e081a4742411a371
z73f1ada4b5a65e649aac25cf7f7051e9f26f30c1bcebdc5df3d202a9b930935bd71487cf6c1387
z91fa9b5db4961ea787403e70796c916bc54518b67192b4c807a69091f27f9f7fab20fb9ff9f2ac
z98200135c9eeaaa7e0ad61483f9c10e81e8c77e6fc3fbe76170f290c23a93b8efbe29a2bed1248
z6ed7cc32d1e33d7761ee7dbfdd0e7a2551728426538cac55a790a1a21603efda86c1c12fcbb505
zea00df80049ed62d33d29115e3ea3c92ab4dba41fdc07053fcb6fc2f880baec7dd8e2d6e1f7af5
z8376baa0a7a44af4878a1b8847f8e44c5dc96d423943a720920ceb16f36bc9e12d5ec54e1ffb44
zdc87fda47e9baf6b14ad6cedc309fad97f96e1a4e69bb4e7d33459a07907b4b773cf9e7ff97162
z9094e5925234c7963e28d3b3459f718969f7a32c7e90829181c0ca51a04b0893e0980ed69853c3
z9334d7716950b705c22c4b5a8bcd67390654c111e6fa37be1871b0fedaf427674607b9f4873e33
z1eed4f0a976eb3299d8df2e5aaffbaa940593b2f7ab032fabc4bd3c346a9e54daae7a25da8323a
z8c91b7798633813aab7f0a2523ef0d982d36f52e6df8c205186f0291bc12c9fb5c78fb59579010
z86a9c9d06530e88366e994eba8026fb9a1c148b71ae2719a4cd032c1567eee9617e766260f7a77
z4a107970e430a9e124ce47ed1e76e1415df0245efff40fc47897eb7ac2988503ceb799d7f2b78a
z0be36b675bce0ddb3374b524a1a4053cc2d0e00a3b194fb91d69f465d136c76eb24391fe7d956f
z065949dfe7294ae222b9911ff1c325d650c9722be85a0f82ff5dc216079091af7ffcc3a6f1431d
z6d31a70ef91b3fd86637b9a73f2931df1b2b2f6ba2057e146b4d01d9a0fe68861499670954c38b
z622404ac95c79bd6f29ca5d6be016fd0b092b8867db8413120bcd19411fc87ee27138cd2fcedd4
zcf20dcd1955cf5e734c97f9afb4858f1b7a7890dd8c2b73d9d514d8e3284bab2083db8fe4c6244
zfc54125db00eeca6a620efe7b1555145c2019d3a41feddbcca121545d2d6e9ccd74120c9d46161
z730cc14fce7fb0544a039b23d3fa14b4bad43c8572fc5e3103bfc8ac22b8ff4fa92e819e17596f
z5af74b6b6f9dee8b5d1bda99bbf99405bbf6224b3eaafa49131f40bcad2f0e6c98e55c67680431
z8bdd7ad0a2c72572dc97e80f767ac555becf52dbdddf82f46661864def64a18c8c21135987a3ff
z29547051e5d9dbdfa2bfcec146687b607a054275f2452bc15fdbd926071037d7c2a8add66c936d
z1f4931a28dbc4405d153c913760651c7405f8106e55e1643a0cb8db8c20e5f08371f432a89c183
zc6437648bd734132d205c607776a653bdf44d5f0ca6751d0cc221e0b00b6f527a1edbb0e79164f
z5313eb8638c514f9aef5dde5c4553cc5a024b4bac540e97689269f32320440e2c21849a2ceb9c2
zdc7372987066ba29e40c89e8044166a1e577d68db5852eeb8318a348c924111b88630ae32d2e73
z3c7ed83f0856ebb8034cbecaa53b9bd70efca4d5ca21353184516305eaad8c9266c35458f0f962
zcf64848e6ea2fe1944a50f23342ce31d3f3ab3548b424890d1d74d168d7fba7e7ffa9596eef8d5
z8365b5c3b674efc22abf97935abf9855c2cefd873f01c6f194add94bcbca5157f5180627d42e16
zb25be758e4a51cbe1a059c33cfc5bd02d1ab1ebf86ac33cd5224dc79f6c138cbb057a6706724a0
z5b1074b04646c45faa7fe074dcffbcb69bcb30bdd0d873741f414951da702c4338b49ea8dd086d
z72cf186a8c40822eaecc9924e7d98204194be79d5814e42a9d4c8de862e32202e48e2659748342
zf508908f420c142ad87704acd2955172aa7351f342594c64f4ecaa4557b3e946f745488e8bfd75
z5983ae6e50c542a2bb6deb96631e56e787f24ec445c25d71838c4b89b9418284b4ea87b8d5fd5a
z864a2e8e0a516782826fa52cedc1e77f6be0519ed82d59cd9930628cffbe1f3c4c135f2f756158
z28dd93aa5cccff540d19926dcca5991ab068c9fe0875d50babf0cc7ead02313e87920541abe4e8
z903467617db38aba4a736da97d19c909933d2d964883857d3b78b18009430d34ebcc737d081c0c
z13f06a51ea034f54062c61f11f81e5ebf5327efef84068d446cdcc3d4b7ce87e5d6781971c2793
zc1d2bba3043b2c2d992f618b4d1336d7a78f9ab289cee79b6317d93886dd50ae63417ca1fb70c5
zf78c26920c6cc53660f38765a3d13c741573a18978b47b3e78d5707d0c52af3f3057236ac42ea7
z2146a1810c39377f4a0169814666f0fe8401b5368c2f76fd66dbc326a21dbfd0a463b6384ef7d9
z0bc224f245477ff78686d56b23018752045e5150a989a1b870bf2688241131107104e59ea567ca
z367e5a99d2e07771eba586c6d64c39776b960e3002489dc4524c0a1c686f38365283a2d0fc7f82
zc2bc4cd4d0484bf134cfc01e394bc134c3d5fb26b2c509734118217cb0202646c85c76b6ac7a36
z1079b991fa950fc0af9608679a823b3a05dc31b75d2f8590d412d0238f3ce2901bca4b72a9779f
zb11310a8b83741aefcb1d1175c08a916018a735b73fde625b677dcce5aea8512acbde3035d55b6
zcec50b9006a0ccd2ad2cba77cf3dec83a2feb9f54528195b23125bb4f6c000f57207f221af6b19
z25627487c3ff5e39a6a8e0edd6907104e6499dfc06f1742c5d2b0ad89eee8261929aaf97a5c315
zc3e4cc93f6fc9cb63956dcc5be2b8f95f29c593101c618395d8a156e9ad25343b87677db2d99e9
z911aa7676057fea4e25ab76176bf064d849de180a260d6553df720bc3d2c133de84fc279727635
z7975a8269475d292bc995f0d48ab9666c838a2645cf8ab81691dfe8fc26735d66669927e8bcfc6
z68c04928c884aa35a1682af07d0a2267cf309a620439c9d47f76b3d4e0d55bc074f0e7f4627810
z2e1da08cdc5b26c7fc3d2d469ca54c805d8ee5921d9e0075c7aa4ba5d006200cc159b49e0038cf
z119a54c8911de191a17d2ebf6abc97e5571ee240f4d9dd09330b0e991ac1c77d0ad1dc6408092a
zf00b16e0764f4af85d4721962b5e5b44f4e9abbda6d48474110aab9c0cf4787378b5b6600259d2
z17fd5c6772ed78e956cdcbfabf0fc681cbe254c3620ec9ace9649742c843427281fffc8be7ab5e
zdbe87ca4e1878c49b2ed09ecafcb0434579c0ddaf62fa27454e40eddaf6bbfb55721e9b5763b28
z48cf46fc7b5a73f860731ed9cbd3751612c5f8e03c27d32bbe8b94cb027b4ea3744b47c6dee7e4
z48db9ba1260e5b2cb96bdc7277e6f16f0152b1ea6962ee448d6b645cf77f27d304897828c00f1d
z005255c6f9b66acfaf29bb2924d557d2b0ec2665f69fedf9a9ab5b8b410796d4cf218fd4918e31
z1fa4953cae066bb584e3cdbd0d8bbd08e6e160ecf91e50a1d67c64d10c828d2543d82f2a77abf9
zf9e4d682664d7def4852bf29c9c0c3480c74090715b614bec75a27bf47397fa00d5872266eade0
zd566898489aa7272a09cd0b4ae8a5fdb10e6bfacf9e806acb0cb5f9f093c9e4274d9bf396a08a3
z9204822b4dabde124dda7c37c4a37f5ad7069be82f0bfcf908549886606b6808d00577ff520edf
z7dd55db2f4f9fbfd0dc0b6a0936c75c05d535bd53f951e576096e5df93e4fd86f5055a011a4b13
z2f22bf0fdeed6e20d7275fc965cde1e1be086334bdcfb86962ec8954f2d71591497c89dbed022e
z9b3f59a76f4af11712e0ed9ee90878a509f35cbdf861861ab3812feef9402d38bba569e829d6b7
zd602aa892d8fca7d3636eef64a3f8180ff6da2d8e60a553ac62589f0d537a1ebfd0eeba4c2ff4d
z93b12fe95342d5c363d8608c8100f40f5f12b375b4acf9cd3fab2da7e8917aa37866277ce00373
zf49b00a782138fda2397023c79ec5b2a703bc8cbc50a69f0ba98bef35b985a9cfac9175b83824a
z84344c4aba720f5aaed696068864bbb7ca83e83346253013dacef4d64c36b03163c76bc2a7594f
zc22ca2f99361559cdfb6a4c5a193b14d9003a23fdb662144dc4cbdaa45a6ec72fa91f77058b554
z602248d9efa662644971ddecf1cb82b79349b246a16df04a0237d01581ed4ad2edfbdb23e35082
z84478bac1ac5719b6c1119d7345450d7f70329216a0ccd79539cddfc636af6c64b7029458de780
ze6c38d3b85c2f4ecfbbf06e1b7f2bca0452b4b5269727f11dab7341477b5cd6119c85ef16dcc3a
z8d90a3c9509289842dbd82782708a743526fec40a2d09d9e6c4cdd291378c9d30718212f131706
za4efd877de2fbc00809c62d6905bf1a5338de519636524a330b32443a3d5ee6f430c5e5e67203a
z6645601c45f1a946971e25ca05c7061ba5aaae74750122c545a535b12bb352ca537fe401722b4f
z54425d795982bd004d4f78e49cac16b4c6d02c198b09b6ca567b62058a5178c26c4443ee559589
z54932b004a1dd17eaaddb81ad73e41b19f9f13d1babe2a909c3f14bff7af2f023483089c751cda
z1788f8a3cc536d76779d1889c03aff86e12ebf55b2cbf3013fd966e49f39b081bef7e2bac2a1de
zd1d1dab5a0efd931c25a55d34d7fcff6e62e391ca704dec988b7bf5acc461eed207d10eb75dfde
z9ddc883fe660c78a1a29366b7249c93deaab1349562fe623926394788f33ac741868e9d707549c
z858c2c390e57ff489f66f473498df6f33656394f052ee83015afa3088f3d4c5d78dc340f9a4521
z3d3f160cb5854fce56fa3af8b93391a2b3f963bd778026fcc2385c8a83171b4bc7b079bbe27eff
z5c862e9f1da8b7caa3f2859ce29d77c85b84b44581cf6a153b7d3e80cba547ddca465c46187baa
z13c2e6e7a6333a76a741d27bb7e8a0a515970130cfb3686a89f499daadc6311c2b160e5b2cc52b
z7d9fd2af9b7af90646478b7fd9eb8f58c8fd45128e2608a7ef5fa0b0c0c159432a67ee099ec5b6
zd0c4094a60ae448de6f8490b17770f851eb40d19cd3c889244827334c5c081baa7d3a28575e1d2
z2541931350af003da0c05a6bde54293f0f5cfa4735a68937cd9c7f9e889076e129a4ada62068e9
z7fdaabe2acc3be7458864832c039eb8091485933d05c03b151e72ebcd3a1248a8d7d2b591a9d2e
z8965c249af8f5ceb244156cfaf3ded883ac8b9b02eb932777b33865304311bc32e42de342fca77
z0dedaf1ee66af0432d5fa2dc14d78a271002419e199c3742c616159daf2a7722f7fea83aae05c7
zc6601cd14e427150c3f87da6a177cbe85e145381f32c7a9fe9fec237a128ed4545a3765f267cf9
zb46490cb6e01d6f13ac876209bc2b11d890324a53ede897b5c3ff7dd883839e117d32cc1d69765
z30875b51bbe514abaa6c25d08630db4cbbcca26bdcaea8ee0bb54f1c05f3804f65f3019499bfab
z84ff02347fbf26542ee67f900ff3e9864247ef4532da6005738c7f62d87df4673b228fb1d7724a
zd71eb2a29460e4604583a4c1ca339b2b5a0a6bb3d9e1204af64ff3e589cd5e5446b84d3726d86f
z43e4e241aa72e1ddb361f1911e85506e29a16bbc5130d501dcef0b2a831753f6fbb8a77927f81e
z59443ac731c08712ac74f82b045d8a35d2f56014d9ce4f08a95d3e627c148f67abea9f0330c952
zad5a40002934dad595f569825c64cb4f06b83c3eb4b73ea16cec5dd6202b29c69155be67ca94ac
z3c7f5f19f3b9694e54b98a3b2981f0fde790c7af718df15bebb1b62f84cecfee278f9ebbb8841a
zdd3e5c86934bdfeea00f3af3bec60706af599971bfbc89c4fa3f7fc5ac70a512c511a9d1c4b16b
zf807b04e0644438827ec6dbc76568d9c006a11ac8fdca4341b97f28612782cdf7f5195f5468763
z6fcb18afb376fdec34b9a9c20a6c6855e27961501f583b9da769a094285867d0d9886be56f094c
zd977bd58e3f4b99f12b53cc835471930637c10796bf7f5120299496bdc9368100830ec6f02cf1f
zdd2bfe17920d9cf7e9efc0abff48aea44e2af4a56c6b4d22b5c070a07b1b7908891d4435f3956e
z7a332ff84ec5fef0bb1fd0ed1f58352d5ec587ffc9bace9d7efc1def9c665cb48549002e2f6318
z20d2679f92125bd96955fe6a128aa759c78db9746ae87cc195b56b7e3e0b26a179d16061816ed0
zb324f6de75236f2c512836e2706608c02b4f125fa0a1dc8f95a7d42c8d78c68ee3a4971671261b
zca6a87fbf067d0db2c4ec828b772960e651628780fbfde20a49b3770d162762d31051343ae8c2d
zfe31f1eb8fa817b8da44f2670b44bb2c75eb88c2e67880e8766e94f4479535cfc3c6fcdf94b3cf
z8863bcd1e49539156ea7f2e31953dbf9675ab7debdcb53fbb35f87edb62b219797e6d13b2efe3b
z67b9bf438e1f7e9892a2a78dd1892b80f6a0d2f19dbb66075096f9212a15a9966ced3fbd2a34fd
z9ce16b6a32983c30351f026d1ec4cf199ba5ea1534adced0f2ac2071ea78e248f37e5029b38180
z9160e1a91c9434e9c31e86cd38df7f7c3ddcf86bd02e415f5ab1290a1c7f745aba381e683ffa88
zc548d5feb1426b2d653772faeafa63398da6d619f5f3b8859f1cd77015ee5a35131a2c3312daee
zc77812f88a9b42db49cea32c9f08140724a8002e522379f52a611a8f202ccb645818739d61dcce
z51b968814e436a08fa8fdb41b5f5b214655525b8460d8051502bda22d42195264604b9108f419f
ze5b316517e983c4f782463c6751a4335ca52700f8f03122e05e88d4963973e4ebe88ec4258f322
z9a2ccbbaebdc65130756de0d2f9ee113a7dc2911bd301c3ecf369560df5558f1bccf03e13b43cc
z5d80c07b3946dbc20275d5cfbcc39557e44a6796ae109e2128bdda4747acd0b9fca41fd9157756
z0f48e7531d436510cebbb11d4022022d475c5643ae067237423cacb698b877d8e3a342a9cb25c5
zf81aba833645812026458a9e7f3ae1ddadb6cf9c353e4a6ad6cf1b785a108c6f4aead3dddba099
z31db55d341fec1686330fb87a7a0b7cf469fde3fdf072beb04168fca7353b599d53135f1813063
zdb5907d6a663e06d34cc65e29f48e2a227587a00045f4802f0341c5dc6ee98632a4e3a7823ef0d
z8ad5975a2e562d2fc14f3109d66f7fe925b73590992c1472920f036c2a8221adecaeafb1099cfb
ze9f7e12ba282df6b51cb692ef9d3f193f6b0754e2e772fd552090e6297f00dd7d1f40afb967aa2
zab02c1561d0826caf2fd4c90aec8ed1147529f459d7f77cb0400b757a6957346aa56fa26ae9235
zaf340d54489bf601b87b19e6f2bfbc51c4d6b982cfbbc766f1cbfeb651dd5063653f02e8aee1f2
zb39fdb293f3c57539cfcf72a7b3385b3ccd87b4e3b4f587748f0cb0c81ef663bf64fff6c3f71cb
z1961c686bf0cb8fc388edc60ee3b80d2782e628a85609bac05904b72501d6a57362879647c189d
zd219223faf3f1815c43c0fd281f4c5f5e135ec1d21da14d09cfcd9f1eacad603413f9dd0d725fe
zfaf19cd4a47b67570e548f6e4993b20aabea0820d2f6a6f4f88bb836432e7e18e75b48305f3119
zd7952634e74bf540603b1d4d094d82094e2d2e1fd6e04e4e1d16cd4f06317dc40cea90a0cfdf2c
zc7737071e119e04f52ed47a2a1c9af64e3448f18d4170375c609c6cd18dc5636fa774ddf153815
z31d224bb42e4703d596503fc2c5ae84e01a2c3ec0e984c0b4e9480707988a977b5b5c57eff19f2
z5b975f63ba179e402d6d665a1c24aeacefd33d6c266b2d0856298fb2f7dee4550521a794350016
zc9e94c3824403a87e74cc73d5fa711b109e694e959f18f4ce78da099ce7c8186df91cdee02c7d8
z2c00351786dfe7006036f70b24307bfaea063d4797c3202bf4178b0038ea86c4212a0e247bd624
z78015c0102e2b5b33e3bc533e7f8f4d96ebbbc1f5631ef9e33caf138c107e884aa05833862298f
z8f5a1c724c7b558f12dbd30bd77606ffa604e40c42aec73fd2277bd19ae33cbb2c0acc1a868f6d
z8d652a2cd54109b4677aff6925a50462665cb2f0bab55948b1cf65d874c7ec44a2f3ee07247dc8
z839df94a384207e99c49d4d6172de94f6a2d08a6e1b67caee548fea89c098e33cf9c1fac698164
zc0a0786692a3d31bc509f346177190afd617d6425a930cc349d10c8857bc7e1fadfb6d0a9d66a8
z39b2a9217d9bee18fbad4512f62d84caac54e33552422dbcf2d79568336a045720cff110f798e0
z9b61ec19e181c8955ea84389f7523387c7aeefc63ac162f37a82d2c9a51c20da5fa7a1b4aecc21
zd8940e2480cc75fb5075958384f89bef3d78c3539736c2c1d0f69db9664cef66aefbaef79f5ce2
z02464dfe79813aa84ccc296be316f94b3a26e87e8ab9e836e8edb270a1895dfea7ac8731fe24ac
zd1516cf94d28b721af0898d649c9b8660ec6ed98436f7aa0fcc1647bc00e378d0f30e3fd27ec70
z7310e3b88ba722596433e1079a2068c4cab6dfbcdd49180b5e5e3012d8fd8f00846d785c4d706f
z4676f5b3c2753badbdac07f4b4b7e72ab5b088819ac83a1cb6c2f75538bc364d232e2f51c71a34
z08c8eed463b52d24397ed0e3ae601eaad243246ae5e56aca99d1744a810fd3e4e9d1faf6fdc13a
z51afafed53f16a96cf3f18e29e14f38d191e9e6dd7f53098a68fcd1b9c993c6bf373a67ee76ab6
z3cf02d19a40a10cd35dd86dbd26a669a9846f9f7d4aa4937c4c10f2708fa2c434a778a793ea611
zfd5d434467edd915a645263f664c7b00c0b0576942695ad6538a10feb83bf3dde0777b8562b996
zd95d7a1a4241e62bbb27fbe4f40aec8e165d741af3d9d77e7be3075ccd14d0216a33f5ca369be0
zbb979c307f3502c0db77137f6f4b7fdabe7ef5690f20d5cb570c28fbdd1afba62d300b13eb7bfd
zd9339d683a1f316bddd6faf454b45bec8ac97a4ae8d3156595dcf1fd1c13a33a95639453385365
zfbb34f8aae27f611f362e1466689d551d1cfd72c517c58b6e14fd2c63e188de3865799b4709a9b
z9c7800116592f8769b1c426fc7a2f0411ae05221d1673e2e112cb88939fe19de00b335e02ffb4e
z5f746b7d42cf45da68492940bb4083419a29a4de6f7c935bf195743f9acfacd2dc0cc2ab033a14
z7cd0601ba77083c256f246ef6b2e600f66fd6864ce9b894ca8e15780685f597b2de544060edef9
z990de7c28297478a76f25477558a48778a32e278a46ea28c8f17b548833cd35f2ba95b9cecdff4
zf2de6d5ac97bb49e2b36d8d7c8b51ab2bd0c0027a415a94d023c3dfb224ab2ec7a829d743c0c0d
z6b04c84c6c0cf4235d79d93666bc5ebc4b6ea2352d335d2e9f7fb74d5b9440adf2fb87ae90a76e
z5a1dcfaa2313ba132d60a13c93bfe8673a7730df67ca234542b8c851539ca5fdfbe5cc5573754d
z6b81be2e8fdefb61b07ef0d8a294afc72f20d632ab3baa3bf9ee8df919d9145b7c5d88f905f269
zaf11dedafd7cd947fe0c21153aecf1179b1b1c1e71bdca0cb143b52cacfe3ef9800b3a1f565288
z275aa2f428d54eb6d0a6a0decadb67189394aa6dcfd337e0e25d435fb023ee5f940fe9e90b175c
z67d85e675ae63d0ee75cdee39fb9aafa779187c5f73a850f425a80c0cca18d484705cf3bd093d5
z9a161e7b7f9dc096fb9d3089d4823fe61593da0983629ed13f84d290eed00c4103f8672ac9287d
z47a62ae7922df544f531924591101e54496ab568823743babf4d77f508f26be8a80a2b869acd1c
z52755d7924e2d154a059a43c3c339ccc45ba2d0f1ce6ed26068b941eabbc16eeffda189eb48e38
z66c67640ba2845c765cbc69e4ed47da6f16367689147e73f65bde9d5196508522ecde1f8c7c949
ze66c36bcfc138eb30e312048d07d034c618677849f1ae29ed92ac21d0aa3635ed5c044e602442f
z4c5cbcc297f791c4012a880f0015b62b62ce42af9f7bede0889d35faaa54a40edc31c42ee3a7ad
z3e498dbd2e93fe44372eafbd29826367295e87e79bdd927ff37f83fd17d75b728d3dd6a1ac6a22
z3ef5bda4ecc6b187c93812fec0fa42e3492438ea5ab3806fc28e397e90dc496b072f2f0f3b03db
z5180587d44feca9116dc5dc9060ed1f456c4c00e15a8afc2ffbce6474d094b68daa5f69c04b1a4
z815b4f95839861e92061d753de9fcd9b347801fe44c4b9dec0503b0215d1b623a1e6271acad4b0
z458e2045cf30e7e10f4fbffd65931f8fcc5cb3d10f01ab5a70fa0fa3dd935017b8d1e6e6dd3d2e
z5a5e8262501fe37e8b277ed2db6e13675fd6634ace8bd4abd10459e2ae1d3dacb440dcf1d7879a
zf5c4efe6a00817317eeb0359a58c8e321d3dffeae392759c41a2addd3b5b3d96f47fe482f23021
zf3844ef7e977c3d33da344175f331adddd4043ab69b908d546137ca751fa118cb41211073cb689
za3ff028b72428372d1473eb042d8ada507855e67a96255ff71c75873f05b718e4d96817b62e417
zb0e0e4a06091ad35e81af3677f3320b44bc6a0b98c25e43ef06863b70ce4827434d313b46c99db
z3575d9260173f98495732515880917ea3e980613c674d58805820cf5a92a61173df2d53ac52c7a
z4895904693527f638e8721acb6f3693248c467bca66e6a60ea29e79f94b849872e1237c2a48e48
zf19f27800ff90965a8224e01033ae0152b7df825603bbb0e7997e4c507a8741d922ad058d8575e
z793f35074851bd4b9a936364f0202392885d74d85678192c70529d8872d4461c1e3c0f99224805
z2f701a0ebad416b9429d317669816ba13c43412ae57303c2ff38870089cbc0af7bbcc89f0e87f7
z59525bceee61751b1bc624d875d42d880ce64a046509aa31f7dffea9680615ee6f4e8d47e9ebd4
z95cc7ad734fb43dd2c9926c46bd0bbe2456cc8b338fb210f4629a8dde53ad76073262ffda7f8e8
z6833e41cbdd9275738041aa7695f14463324367def5824838a0b35359faa0b05cb2ff6fdfeed38
z5bf4f6c8a28b85313b723eb7e4171ce73361650fb33ab5debdaa322cdb8acef5f48118c3dcc678
z758fa68ca838ae9e5958a452a94856caa8eab0c55900134c9b191791006fe7de1c129434303906
z1c67a12820bc5083f99ff7b1858fe4e45652c63ab2ebc8a4df220b8f1d3e207416bd76cad26bcd
ze4a68f328ac5833d5e2dd15eec9d2ce1c149cb74ce3bd715d571c3394161cb2df9e25db221deaf
zb437bc72028923cff3f6273e2be3b466724b491d178ac256a3bbdf7ed16fb8e4369ed920bb57e9
z3b84c51d939ff11e2aa7aa07ca465f42b942113ba05350598eb40d5833384ebcfa4c0bc6be9dcc
z717e1c52c776ec7c50fffd8be5ab06cec7f209a604a0e6327f3282da7f8bb3006b3ecb729cd848
z3b89abbd00ea1285d21dc22cf7c0c87555e1294bfb12be0cb8d4b2074b594a560d76594edeefe6
zce51d2afbc379ca27de046a8afea31d47910b13c84216c6c1b591139566d9ddc24f6ed1bb1154a
z8dc4ac552339f5347471e13e765702019044ff53ab26ed03a97aeaba4745f329f5d26a2c7e7a04
z6806d0e981393737cce34afd62608f574059f1a89e8eec232a582acd7d5554788a9ca8f0b67227
zed7c1cc95245e88ef1365c9481537819b213352240aad6f8f4f438a4fbacfcd08878f470ea1d78
zde1ea40b6229beb0ae10fc13d59a5c798c887344356f3540cf745e21fe4bf1de85092a6a2b59ba
z638172013b0e6d21265147d98d59fdb1801a23e335681edda75f8f9b18a4b60c43744f3e7278e0
z508c7c2af7926eeb18e47145583f7be950e93843bd6cd29e1703b0efc4af86a08cfe5b1d86f560
z8a96d197b91ad324f55fa2f8b3a29d76c6f369acc14a5b5ab4f86bc0613b10a7044132812e7a9f
z2ed76a4192995dffe6d7902a3d03dd0281166e6f525c3ebe989e786250cc2cbe0bad31cd0f2fa8
zf2374e3ce30084d65f61754b6c094ed8acd285e83341b694ff31bc4b83be3615547fb256285aab
zb4ce46b1b0aace6ca46fbf9e36c5427f558caec90ab227e6f362d07f33604b31eddad9a280faca
zda65afe886f1fed15ffd7fc22b6c7e3032114734fa3a80280816eb8cd831d22a00aaabb8042961
zf3edbf392f946e7707db502fbdb0ec2f99f7e1605bd8c3b4470b783c53e15a4a3e7cea9cf3815b
z5d9e482624fda2051b7ec5e16d02ef22f4dd731635c590262a6d754c1304df10b9a90d1cc13e46
zf4f7f7e72e4db4fd1661ef94cc64f5581bd7eafa72c9b61c5c247915731f48b9f22fbfe8d03d94
z32e3ecc898287f0a4b9134be851c09ba878fda1c64ff83a8c7ca22e926fb10e0ffdaf76b738f93
z1f338f6274c2243cd0031b183f64999384c1d111b110f5616267cb92df5082473a9cfb19a3e4ab
z9bf38a90879c1caec7a8736698b8f5f61a90626591226fe775f4951923a7469fe9f2e41c5e5564
zefbcc189339052901c61bc192b399aba838467c8eecea74853a3027675fcd3fbfe7719104353c7
z3300a1d62d2ffcc2fce24cbe7fb7af21a7bda96910df6b2e3668c5f3bff6b424d464d2b64625d8
z65c3595d21ee1789aa6884d8fd530eb740df25efdc6e3cfb6e3decfcdbe3f16a69abaa07614655
za2184da9512b54dd850e56ecd2a4630b9656af7a9bf7b89ba371df4c9520612248dbb23d08ca7d
z16719cb399a0fca9004956712e3cd362a150af3419b32b3779fd6a0e0581a14f7eef9649aeb3b6
z2ca7d1162aca9adc15619a3e6980eab1d9cb5f98cd5301eee094a2f28b335cbc711d1223cadb94
zf3b7eed76d5c46ea3ac85bb5e075eabe3e1ae3551fba4dcd298dbee9d6b3c9c5b6ec4a427a6073
z9fe35d90599c7421804f1aaa7444a83755852381c150f5cfe84d98de74cc4e2fb2f3447a32be4e
z27f548ab19dc1757eed3d8221e90343ae5f3220edf5f40f398314de2cccc3c8fcd4918e4615bf2
za8665d550a064380686c2d3c6d360e701a7ee01199da9b638dae6fea72642ceb2abeb191e9c087
zcc091ccc737946954698c56b220a3d96b5008826c30473bd5e84d12ac1fbfe5e80f00b06c5c463
zdeae3abb20e2e99bc53bf48e19d2d9b2bd2c3a74ac9064b91004656440f024b4dd3b043e6dab11
z28dfd0ceb6fab34e8bd31f2962050605cb9493a5083ed342a9d442b22e82a59cdd1d5fc3ed5324
z504865f1b2d3dfd5de425566857bbf70f187a4a350e95735cb0f76e2c3ab75f345e8b2c8ee198d
zbc6929c2f46fe80cbdfddbfef347f5c02f42e2b3669bf16d0a596c69bd339d85042046e84553a9
zdade6fff994b49a8cec131e355477c46376aaee07bf048c4180128a81a4ff442880daf7699ffbb
zff9140bda6c40d13a741ec499531bbde9809cb858b8600e6773a8de60db951aeaaf7d5bc6c21a4
z885e61ffc5b7b8a08ffc16019abeb69e68036b859fa1f12691d65866993120d4c4951717c31dbf
zdc2e0c65d8f1d6725bf72495b47c5ac84349cf2f7064e91c4eaeb0c6e5338715c22361ff4ea09d
za24a64b21a1fc346e1ee99496eaab515b1ca7cd6461bcfa95e852d0ee18f8b97641bc53237977e
za74bf716ca6e89c367e74983648d9e01e192c8f89aea5a05a185ff2d27bbf1a89abc733cb9e483
zf80f17f03f63ec06170c027f97661574c25bb0454020bbcf0fd276edb3e3918adf35b8d617f697
za50b86790147ae34bea5295588ca5d060f22013e850bde2dab7d442d2419330a654875daee5f65
z3bf6fe5117159ddd23342315222586f21fddcc42f8c873009e0bf039c9f7866be3b0c85a2a7a82
z4844437cc4ba88d6a2b2d3b0b9aeb900e6efc8b6c907cc99bc5bd2d5d4e4d022042d818927a12d
z01025df026d8ec20615057f32154f9ea3abcbf818d28e816326d0bcf9a7c2a0f1af434fee577a7
z7a5b502672b54418d8bd0ea499f69b95e9dc5f20ebfb71c8855c0236734de403cc9c76ea576e5e
z9e6715ce7006a36c5f47452b2f1a549927e7d7f9bd9445ed9a0ce0901b5c87a93f209d34fe9edf
z433c85dda1b2d6b846476d92b74cf4e9b6c3f605fcdb8ad1bd59b5a29817726abe8a7973f5f2f8
z9de7ad4d9de577fd4f69dbd750b7d4093255da128a62938f2507dd0823830cc687cd22cd4b05d1
z2b3997306d7869415537ed3b9a86c5c66713f19877a114bf0ad3565424c9341ddc878211e794bb
z145e5ee78f700d5295427d6a2a23fbbe8fcc1527885f0edcce6ab94dce578c247fa3a56a57c5cf
zdc37cfd0be7b33f0dc8f2772321a97a9749f9e0293020b570695773238c54d340c3e191d8fa611
ze1b4270b629527feb02166409cf3c45bf8ee15ab66d68f0b683b52dd1237657accd55af51e92ed
zfb60eac99f8187533653f535c76264faf1940b17c9a61a14ff2aecb70da543868502a2d337791e
z0026701f1057056b1d2add9f73239a06b8caf84806f14bac1c2c6970e195225a107d33b3b667e8
zaddd7cba500ebb80d77358484fd878e72ca736f11de3148e731540bc9ddef447e8477df0d3db93
z9ee79f5cfd1165d688a7cde3b32bcaa27e7471238a2c6dc69b2d128c185254bab3f6e8362605c5
za1d04ba97d572556a9916fe2d4ad108a0ea458a4daf84e26f027afcc86ca7b1f69a3848f71ef50
z708a39331775722317de70bfe16ff23b5f2a9fcc0392dae3b0d5916b78c7a9e5ac767f5863ac36
zfb5e017082543d35276813d944f13a4cbef9f813e7e37bbe58ed7b6e6cdf6dfdfda95f7be60b33
z4f4b8ab347b5b8c998582fb2fdee37494de8a5c6d9223a4e0d47c0a24f25117010dc55ac58cbbb
zdc8350cc4ca783b1dc40079ad0f3b74f6b83358f68f2cf729abae96fdb7ed1886bf45e9966f2ac
z80e2ee888e7989b936a4e69c8d595cd0bcb47fcfa7dc81a3fa7e3aff12ed0658c6783bf43c55f9
zb37e03afa05ea9d390d9c9d31aeb2f5422a6c125dc7fe55b958718f4ef2ce106f51d0df02fc5ed
z94ccaabdd25f5f0f407d80e5bf88eaeb5731cecf70f2240e751291a6918488e987bea7812be947
z88899fdab5f13d2911fde6498736bafe8a3678d6166c837dff580d3e3744d75cb306e63155a133
zb6c2ea17c82b21661a73c533cfd1a673c96e3c1062021db7aed4e76becab623506c5f86143edda
z870f4bfdc9f17db8ec48ce321b68f1aa8702365318e578434075d6c1be2ba4235ae005f4df04cf
z74b35652e3127dd0bdb7eb1a4f13759c1534587966cb77d0d45d3be9adb3162330ef1a8a5a82be
ze0d39320bda180bb48ac956787410694382477bd73b300e804be00b8e3a4bbd866ad47139b92e1
zcdb1f65f2d89f257d1fb175897f191292f219fa64a1c34d4e8e867e44221a84dc7e989741a6ee0
zeaca97ed477653e8f8fc2c65fb993dc4091af45693e71492b335b1f73b3a347fed6738de443cfc
z520f5f75eb65294826ceb2a653a56767ce1f98c8f921b1beccfac07b94b1b42046913d7d87d372
z418e1fb4762cb10859ac7390daa4d2a69959ae146f9d6509c6b755aff6c541dabc83c2cb2f1222
z9a0a9699c28f5c6a0f4a700afa844915a07b6099a20dcbbd38a5493635535d72e0e13eb8276d30
zd57ead3e60dea1f25dc5a7dd64cfcba287f1a098e6bdea67b2071ec1a4f05b09ccaae7aa46caa1
z49713d0ad44216a757715bc3444d036417613a006e57974a02dc1792cd4f9af19246b5368ee498
z222649a0c9c32c731fe124e402c9173d0f0ddf0e92db06c3594f99579aabd17c01f03f2bd20740
zd0a9e532ad18d82fdf7cc9fa48faf0995f578c66c12c14ea6a685331a3ef00c98f3b525e58b4b9
z93949110a832bc6a5a7dc866cf5ae1154e400fc9aa98fa544639e7422922c9544c000aaf53e396
z0873dffc106154c318c9922acfc87ddc7be7edd5bb52a0835fabfd7f3e9e48668dc7a9e3696501
z457ee4154b035095873bcf7a40da352709c3f0f9590d8943b48e299c43e458b27e68024ecd3ef4
z162aa3b7197301be3bbbda3d2d16b3130400f6ca9bf807342b80e897f2321a16951911a200ff97
zc0878a5f888bdb45ba47ce128d5ac17906add3890b331657d2c5938e77f372dea023ea865b9edf
z4fcf0222fedba6e02ee86dabe3797db3e9e36037495c44a7c7b920b95f95bad081c0f26b2764fc
z24b89481c37dc322bfbf99bad7679fe6b0faae00dc8caef956f1925e3ae9f44c357fc0363b3bdd
zf7c7e47acb2aa499262e60ed1d2e5b132dd1b1f21226f0d615c88ba27f3e8e109bd7974b8ba3ea
z414f0635d6dfd412b941627d9caf6eeee35cd2da1774f164ff03d46cae168cff7f5607d70ad252
z3624b239dd9ca7ddad8d5269fe3d3e554e21b38b880be6b9d0275afac4fd4b1e9217dfc46f5ec7
z2a4ae0e9d312924bad4849546a9a162dd10b9bd8a1c14c55df7748ad51410e5385056d77e9f976
zf41b0648af4d64c4bb1746bc44927ca070f4b6cb57b85d34319ea33bec2f70994e298f889b99b2
z8eb0bf955bcaaf91ff911f12d589e2afddb61426bda29c2f908d4b7b71359502a2f08a64fa8e7a
zaf3d61e2fa6cb5b4cfe5a895dd7af8a7f8dfd734dbbceef9362ce554fab58cba1d59871b5512f3
zd94527386b718cded9ade97b4e4f06f48ee221ba152b337119776e3362e23bd8f5b941e4b12714
z062b37ba87bae4160b4b2a3cb10394397737f818fea015987ffe5b0febc840d58da5ecad987a3e
z661d2ad3718405c280b680690c3e22cccc0da4b541cb630ea33ed2e64b836f0c922b3ee57e988f
zecb3daebcdb9ca6b9c84487abddce434cc848054f1642e30f51b4c1649827878700b6b05a10164
zf6b74d2c04f6d6a5d151a2109d70610551a24d89f53bdb0fb071b89dc83590e8c92c6479cd5a45
z203c1a32363666a3e14285766119cd78ac745244ed3cdeb4f8504ae1bbd7c966722ef4ebb09613
z889546d8f1498a4eb475ef8dc9c50c8e068b5859e9005777d2f59803a92e5a70f0744c9b03c799
zb778925ddaef9644695fcb289703e6180b41cc0c43bb0ced363bf3090f2aee010f694e9b1a899c
z4cff10e3347f2469e4fc4f06b76fa4a3783232aab8b388b95392dc4a3803ed652afa7ab18c5b28
za7298daff035ff5532beda982d2116155e6031e64263e08f98ad14ccfbd8a62a22fa7a373b043e
z68f71ecda2d89425708cfe07fe9cb2240f6a8e7602d0914ca307d4c2637503533f20003cbc8715
zccce035d6913df654c5803f4200b9fe3354ee9256641f23b2f5da1a055237bf871e3ebb51e8a37
zd773569a0e42d921155806881d9c93d9854b990d82f2b4d3f8e24034e50e910b95fd4456a1526e
z6ced7e262082ed2179f2f21645b44eebf0fa3cba3f6255e55582206291476d86e5164e8e61dafb
zef6ab381e81a20e9afb381c6af3fdee9020849a9221a18e236e51904ff39f7ec5d647c7989e102
z7cf9d420415a9efc5e32199f5053268717a1c835822dab74e7c3e0cbf0bc789c7cfb64f1441221
zf51740ae4a331fee0ca6a86b81a3a080e7323fbd4b66b57a1ac1c5f0615cc621f2de117198b295
z501152908747bc9daf51e95c3ee77e95faad6b92b9f6a24ea586b90c5cc4a037ff059249e662e8
zc1bb14664ba25f62c38859922aa69410cd11cf57b02fee2104617596637212f6ca9c20e666f823
zcfb2a69eb0d5ea63f46d68f6d49b3f4aa88b75013cab4d68e39b2795bc22ea51c8ca0397dcf964
zee88d88c7a45bcd64c5401fc8bda3ba3969922771ba3adb8ac05717e0a491211cfe188aff7f0b5
z994270bd95fb2c65759e97a6ff3074d2a2a20ad5532d06489f4329bc8eba90653e79b234e06dba
z822240071807a7f39e4ea951ac6cecfaf76ac8a753b743afdea9216b104569fa4280dcb75526a6
z983b8f26477386f13dba5581bb7037185e1fb233b88c08d3c267d314d9536e8121727251f5a98a
z242cd1cb0048be3281fca652128316d61153ddee175b4dc79fc0dec7378b6445a675554ef069c9
z20ae61fdfaa429ebd1c2eeaa23eda5da96d0be43fb2000f02a656f1a90bb3fad3172fdee1bd0ff
zeedf1e48cd60ff53f4b0ab67682dc8d3d3f068948abc1e7e12e6f445da39df1a644a3bd52ce103
z383cd7a8c096e1ff6e8a7f8fe156e2442cea83da5c8c5af11cc361f7e8a43072929feb3d2a07c1
z106f2a03c6b5452e30fd93c9f79467f135df2a857d0facd2ba490f4939d14cc0dcda94ffa83dbc
z08ddbf87750c549235da4860e11f817ba16b95d07517b1ed5312e6a0b37086f8936c71dd12110d
z885f1769b354fa6ce1ded34a44190a6db8abf076367436e3db24748fcdc71e82af60f156b8a829
z8b966ee3ff23021c0a340183b79814709a795a96f92565cd4ac473edb50adc5f5ae9c975f7358a
z5eadf43ef4590fc08dfa54b193a8865d2e71164c718f187faf96bb07d2f545c6b07f6b2114de74
zaa8f55de1484b8cd876c50e5bb4f05d360e308bbb274baa6900310afcc8643a95a33f6aa3c147d
z67986c0f0afecad1e687b6ba671dc0244621063404650ae19a39ede6cde3ddfeb9f497f9f31bd0
z75621c2f32b668d387b1821798b1c69ad573bf104b1a644adaccad1d378eae9d6a55443a030fef
z0bf3efc98f3044a6a40b24c3e33e1be7c887e6b4058f5498edb9507f367bc64d0ea44f717a9416
z9d7ea2e7718f233de5fdedc1feb4d4a86209f038170b3c9ce17e23161bd0eb7042f878cdf63455
z6fc309385fe1073f51e2ac24456082107f61ddad1f9af97a5558a166caf61cf0fb7403628dcb69
z450dadef9f2b47189c891c065c0a946501297698b3eb42aeaa0241f399554260493000bafb736b
z536dabbfa2d5027877600b58cbbde0d96205844a4a9311189527545063a8bdcf465fac8279ca4a
z3fa8de7a62f278bc87f497a1266d82df99987995594e7e834fa73fb25d806584ab60ea77789aef
zfb0539cf20d573ad401750071388679403b47d292dc0e129fa32f9d42dcc5e61d5ba501bfb164a
z4396b7ecf4656117f6ea96c3be1ff930fc066780f349569593b754b6a682f570070e453356124f
z396b35595e2b8b0ecca90b2353282fd2afc10809d77d22b6c5bd4eb9c876ee76612356c8978322
z934463f6c042c0a307e53dd48caba13bab330100e0e3295659bd85240015bae9e989257d3e589e
z4488f21cf75336b493ff27887880aa39a2ca85544674de08d78cfb92b55ea51bd1647c9a59da5c
z25e4c812a772aba6baf09f33c5045bacef44c1e59faf8411ae0018c935604dddcb9733fd6009de
z5a35a55efc6e5188ae4a744a109e6c3262d3a0c4d3c049e72da4b5ed35a2d23a428208b6ec0630
z8478b950e59f3a31983f297bb53e2e71edb55e9dd6a3bc66087fc00f75a0e24e7893c952e5360f
z6a5d70f4592dc9495ae9366382a2849b27be00afb2ff7756584a89b747fc5f67c1d465e01c1204
z382b0530d5e369b4dc23b2a517b3d29b8efbfa6a10bde6d094c55abd2f9e7da9a223257fc11201
z3a330fa064f67b8c4f32f819b53499eba3ad55e16a34956ee08fd2b5e4cb265323fb8703b86bd3
z0aa3dcbb05b1e492d9cd0ee75cef2a82293a9b6ccfe004209a1fe9ce0c7562fcc92083f5940b13
z856b0664b563171f6119efadacb0fcaba069671dce6d587f08df48c6945e1c865eeca8dc1b5468
z5adf6b62915bacec9018112e1997a679270f87f7f2ef5fb2b37eaa67c071ce22720caecf21d559
z3fff6d0921b7a9a9401acba98ecd445a2f7be2d1c52a184d562d3c8d518c4db42c46488bedf293
za2ce09ba7211834cc98aa4f9f4329d2c452fc08b847246bfc46cce2a7b2ad49ad0f16a250a386a
ze141d136cfe192b34d9620a5dd17ce79da59adbaa4b747bcc25d91f977264f51bf876cbb67e886
z49ec96e0d1f5dc92ea7e543d40a1d6465b18221741f7348b05fb8eb4041d2150cd6405b422842c
zf4bb73811c0587c75e4cfb0aa98a64af2b2e5413ab34ee43a09e9212f439557678228ec7be0a70
z0c0bf8c836df3bc583d4412f6e3fb9999832640ad15a9f19923784d79d74bc311abe612c51b0cc
za02717a538583abddb56f99cf86197adf22bb9d1785210944566bd2c778f30e3f7c8ec1c3dc2a5
za24979b98b28b27699dd8b3dc687de48f58e3382b076c95e492a1aa7d0e26890be8d3641d15c68
z284201d1a10ff55c05f331d5e803e6f13eacd7c707013997b5f628f11046b5d8d5f605719e203a
z282bf1a75962c29aaa5977985746611b6457112b2e556aba4e9d6b20b3818fba5f21da1912b073
z400a3420a4e6767a5e83272e3ddafe0b1bb534b0e2da718babe3d96988ef9745e5a772d83236c5
z3cbd6a2e1521d1469391ecf3f51586ebc8adf29158c4c0b7cd2a8c33878132a95ad8db699d03f2
z120696a98d175f1f823a71e6852866fb6728ce6c72a8afa8c0a0c2c6a9ce9677b6ee5545f6e2ed
zfe605020fe6545808113c77ea6841443aa2823dabc2bf91dd90354fe0209cebc49d3671405d487
z08b8d936dde8b8d1542b63ec4dedd300f36048921fc12ccbd3292328dc16b69c8eef3cd3da19a4
z3da78c1f9d5b36825607f6251867c8ab07e096d1e580664b337ba971dab2841b9135c66a1cd7e0
zfd9e11411b615cdbff88b86c76920ea08f0b9c5b84c428601222f56582a2729f23e0931da9f7a9
zb838191a8e77b40d287e83b061a8f8583d3baf5b92b086dd20ce022f1aeb9f454f4e9dd622cd8f
z1144352c316fa2ead11fad07a4125a08abf0e785467327c7bd952341274858a7a82e6e20e3ae33
z5a9d22bea4a643fefca218357afe76a5abd8276764ee19230774e5bf88e67578ab85d2c7ccdefe
ze5c6182ba40bb1cfc0d38bc53dbfcdd29b42163bb4aa6277b76329f0f7a690cd0e5b035011a88d
za463e7f0050aa44675450ce821e6284f0b039715227ab860d0b595a338edad6b2f0f57660d79f7
zd6b0c7f937197b699b8299a386b71c98aacc1ac81c502b9492f49c52a42fe49c86857033cff189
z4c75ec491cbdc2493d757e51cd4b22b81c991a29700ffc96512406083c6659638d870131b31341
zff15f7f0670140f35ff160398b87971c33366e514f48399b3701efbdc6123176991202ca7f32b4
zb40b74c81f582b9ef738c020c4d0ba65f50be451b62a2e57d7397ba78bf9bffe62d77e151f63cc
z78bd6934bc704e8669debc7b3b2984ce2d570fafb17b671c596263a0711d84170922e891e536b2
z36926da1cde86c68cdb7ba3602ab9d8c7da9a26a28679af675471141e8d199d492e272f2a250f0
zc55502528acf8b8096201df3fece6358fa1eac85e7255e15059d85ebb551196025b3637ac0f00a
z107159a2377e055ffb284ae6184233c79bce37e686c1adca606cb794f280404dc58abcad9ce353
z1425a8a8d7d95ccea3f47768224ed136161a24a25449683ee09b315c1c33b2282d1cd520a9d162
zf994abc69756b1216a8ffc97edd401d66b54f5fe1332f770fc836c5f4748e26df959ab90eeaf3b
z8eec0dff5084b4e2f0f870683a7a48c5f89cf31f4482cef1cf3361dfe21a8e052dbfebcf7dca01
za377d8b3d18928ef011cdc69cd79cafdac1e74f6b605d1a25c29bf8efb4f36fa30db8db21ff937
ze2585fd29ef48fb7ee2e9b8c90df4fdb3dbbf6723de2ae781f0cafaee2824e2a6e4443f6fac42b
z7d4a61efcafcb9ae0ad88b21ba58806b0a9752a90b243a4c53227a64ab8a714780be864079c3d7
z1d9f964478afa908a2a0b735be0d2b67dfea95bf97a321b05fd0e1642b0af7fc76341cac538bb5
zb296703bdc5b15e95a98424764d3a48e443db53fdf8d2e5f031ee6c93c91885febd5d6d5c32e2d
z7abfd43bd348ad1fc907f57df3c2687f11277f7ae6dba5baaa1b4f29285b6fb5cdb9f94724a250
z095a4afdb799aaa45ae217843e3a644a4604be374c767948032fc0affd95069901bc46cf9a5a89
z9845e36feff1e2e4fd1ddff52af6b123bb223a02283b13def89c2a19f3521c69b4abca11e95402
z10cb51019cccfdf4540f2bb440cb6e89885cb029b6fe53c7e97ff1a87cd69670ca31aec18555a5
z6958e9cbb937e6241e745c3adff3139235783a08f8e9b2a6faa1cdf5d54deb84685892e7f534fa
zca2a9bf4649c1f6bfe1f297e366626c6e2c58b3d586e87f533e366fccd66d0e1ba3c2e093f1530
z1d96977cb1d2117795372852dc755c469abe9f48a0bfa34253be55918d193483c6ea42d1716c88
z29233d48b20bb43b021bb4547c2631630b4fc0ea27aa3ee24b13493995fb89c38844b6424ff096
z3c8f2f9c89c866c3b2222b29ea0df725651c06386d1e8a2493fbab8a846722c90c2927d37714a1
z69b49f6ccd7c78552aae1cfbc06d916d36c43d13d4bece1c2d801b3142fc2c5127604fa18641dc
zd519d410b0b5ebc4c0eb5c353cc8f0b0b7fcd6536554c743584ca311243d5998bf3f223bf4d036
z91dfa7c675d2649f37028419e686daa5bbc4c26733fef4729c9415657f116e0d6d3180bd902c90
z9aa199a08ab2b102bccaf0cb88c51f8f3b983575f0431671a163e8562c5bda1b8f1a5ad4560994
zc313d83fc119378421eab567b68ec12553adc002bb626b916476e8c94045edbd57221bf10b78e8
zccc0f05770d2b165a0cc6448c4bc5551b4c02ceb87d22eccd8a75a20a6b596ccb75f127be961df
z9abb119de6000ea24d6bafc050c24fff0e56593995d20945eead5aa37ea8d7b182668fda44717b
zd2d26042b3e9cc49d541b10da4a0e07bd2c11ab577605511a43438b0370968aade6bc1f86e6275
z47cc2e038dd5f0f92918c1623b5600f421ec283ec93cdf6732e1f8874ec06d857395ce390c69d7
zae0417ba5bd5df0c57a7ea6e4d1dd2f256ec9c9a28186733af66a4c1506f64781836dcbbbb84a6
zd8c8114441e004332f5c1380e59d5228785b5f6c0234bab4fad615462e3b5381605eff21f6954f
z5c97dcf3f6ce2cc3d5be195ea0aada0efcb85e532afef68bc7fc22be546d1d6e42018462198a8f
z1c50a7ab27c13635eaf95a20b78e1fdd32d769650ff6cb64451421d0f8f5a015b07bc42eea7078
zb4f6a4b8289e2ab103dde7f14ca975bb1795ef2228cba3f7c1f545195c60e33e8370384402846e
z089cb5cc3e5d069787977f54d33e6b8bdc69425ab553166e3913fdd355187a7b28944414ea18f6
z834546153e48dc5b0a5fc9654810ad5acffb581f3dd06852f2fd4d86c80922b3613b64c96d9414
z338c230c735ee2d83cd184a8eb574cad968efb19682e021892fe360b539349010ddee6377a24d0
z2385f2b0cddc0d06d9e43088198da2192d2405d929cf94d15ebe1f5a5fe940610d8ee5ac0a84b9
ze0ebacd6ef4df24b1a1d939bfe3dd92e7b9efa044f8fa9440932123c38d4863315c2857347fb7d
z55b9ea9d484dcd615df09b78cb7c68d463947cb3f79865137a05b983c9711492b0a76e8190c8f9
zf8b7b1641e5b62553e63c07f59d8299d1c03b87703531838746099816dfec2818577da14e277ea
za8e9c6569698f27eed2bb50571e24ddeef5a92dc632b3a6daa6f4a5a8a797e4c98a115a3ebef52
zaf87b6b5f0fa5b4f1e9d150b32f6c7a2e99a07f0f4281ab7da958e6e0abea9252dceefd1219d94
z70efe5d16ddc8ab6a85612147de16291d702fd62c071f38455f419286683c411b46be3d7e9848a
z18b84e1b70b50db6e101160c085351f3b17fc16c0c6fa241d5ccfca5a37ef05bca4549a67a5d90
z673a14b984662e52e92ff51e59668c42ee87bae2ccb04548a21e0902e6dd5442cd5b705c64c636
za03430f15ab2dd58c444cb28b6fb4f6f746c1099b277eac3d911445862bb3c939f5e6b14361d48
z0b2a6988a7551448be921c74d99503aa901b0ddea200b7869f713a604060d4176fce501622cdc7
zca3a5120496dc4e15ee7772be16ebebb4ce48cb87637c13f8ffc529c031720d8ab2e385a79543f
zd4aaeba1c1ab7d3c577b36bd5aca923abca59bf47ede4023a52e2a366d63c0466b7c05340c7266
z718bc589c13e5d797d1222b7d228f727a96070d4303a9e678191b0665d94a10da07efb480e0a2b
zdd513e323c18e5a88898d40dd38a3192d86dcce9478f38d91ae98a8405a6380a5c655bda61b26c
ze56f709092747376f45426fb4c7bfd011743774461b3b15dca90ea5d604e53ec614e8245fddfce
z26ab1ec828025fc1e6ae86ce1d8ebf6f73f8259d9aa123dc8313f730d669d7da32a7fd8c0ac12d
z4052f70d9cbc41faf83cf9b42765430bd00909857a193ccc31495039535c1b225978d8793da108
zba5e64a76985b3466c1ef4aa42cd8aadade0e00fec302f40089a061fcabc507ee05895175ac2c4
z9d997d74b2fbc980fe85dd2c0eaf032c83d07e6860180f08ed544097cc4b511d00f5d8bd5e6a73
zfce9f6111cd62107b12749de2884752375f922ea0f4306eaee7b70cbc781c148db1d140e0eba59
ze67f54e4c27339c623b465416b17d6e6fd3f95e05e475b6da13bd024e3594f56dbe296263cff55
zac57d134e47afcfe70d8b65b4e613bb273334ccd1c71aa23bb663ad7b58a0426b4d998112140da
z2b933d5cdcd617d1cbfedc40f351122762106e1ac898fe667e4df04bcaedcd24a2f53d75ab5d75
z75f253475ba4c64dbed1086c47132dfc6daff7998e8460bb4713f81d16f0437f1775aab15c2c9c
z5172fdaa82a7072ace281ab7494c902c05bd868e2e4a257d1a0f8cc3bc916820d81149dbdf7e65
z20a6d3cf2c72a11e6a433c14a76d6c34e8cbfc02129874f9870f7871017f7a94091b05c61e5dba
z2fb409748c29220b5031a41c461e59b1c538b6e7d764d0e6fc6bb8f70ef607672bc54bd404406c
z35734a01bb5b8e112fa4a3c5305241cdce393bb054b47072c3627d699ca97142bfa48b3dfb80bb
z0fc2fe4370002a7d20155e8b4d6907c801264813af0babfc96baa5f64e912160ea345e66450fd7
za49ba70de5ed63b515d111ea6234eff737b54b661bf0a6b136fd5ed39766740cf270c3792c1aa1
z5d23428d428ee3e91b7196b106a9ba0d7ecce95379382aa7768a455e7756cd27e076e02c0f1f74
z550efe5541344fc2e6643e80694537489d930ce7c1d0eea17d988735119a7d1a74d5d658572c40
zb9319b3e2451a2d6841dd48e2ec07f017001093c5c11befcd1c6123db8a7636409bba2e1f21b27
z58b42bec83166a042aa91da273803edd13649445839277431d14013e9b6641f5f067c2dee51d60
zfc6fa564acb50ea654cce64785f8ddeb664af9e4e1070c5f5567c3790efc9154ec6f736033110a
ze6ebe8111d02c2373ff90e0b2e3291b0220fedc861c8c7d24e01991aa9ed67fa1a32f92a639437
z5675fab5581fb52b6f89f9f1d908aff42e59a7966b93c5fb1e42188662134c2df700f78a0d0ba6
zd369324f9c4d2a0691cc15dcec1c5e212c2629296073e9fdec69c1c9766d979c185c206bd011f1
zf4cf7f779fcba5fa2c711911622bc474c0136b53b3a9171f7c911b815a0861f79cf4c5b47988cf
z6bd0767af01ee7ffab1bcd97439a9ae879045809972ebd9e5e79039b0839b727ecda4488167c5e
z6828ef3be7a534a200779a068c23344e0933c1e693b9d21b1c716d14ddf8dfbc9d45ad8cf6033c
zb71437fb2051c8c9bc8ca71cf28c688d98cc3c55660d48a07c60c9469f857d6894fb934dae90d3
z282862e87d180072f38001319aba592e11e9083ad61e113fada17f7f86624e136a46172cb17266
zaf47e6369159f7914f5193a4f62d200d193c73f0421c5a43e8bc6607bfd326bb651f3135ac502d
zd4cf56c04c42c58ee5830706596e3d37546ad72ddc0e84dc8b3f7acc046f79ee8e197650d0e859
z0bfda991ceb6b7ea9cc8ddca2942de47f286c28be5cb4fdf54d6d0330c464c585bb4f3a759e008
z165485a814c5e401e6eb25aa1c3744b9791f938059bd65f8fb061c089a8847e83553f4d06d90eb
zeb2ba82b8dc079979834999f306f323fb990d7170950994cb150c86d84b468a28b62261b194332
z27b2472d3d06b127642425cf2b5e042f525d5e22a61d1665c5167abef6e539e9fe2bb0d3775660
z0d60df9506ba15798959c95e2733e3b705b01439c5be4e29d088ebcd47304e459db8bb33d09f75
z33cffe256887dde50dfb64c419d859272619ecc91fa49d55dd6d33c15f9e7df8618c3a6c8ee008
ze435ac472e741f580612e10e77e463271f902abee05773c183b38f4e44079d965327ef3fcbc53f
z078ca5042910a21ba15a1a0ce3e3c96a48335278e68319721232ad830e8b3670dfae48473ab72c
z55bd9b0806108120b3a2b4c58dd03775ce08baaab04bc3ac9b7df1f21ddd290a6e6072b3cfc688
z96386dc4cba316548bfb2500cca3470e0c98ccf2e1101f884d305a37c147116b8e6a299a55887e
zafd6fdd2f7940944aa9ca17e93145d707c66dd5b36a9018d252a61306d4228ef35a30cc531e38d
za5fd7cec5a07143a45031194c0c03ca42974297944ffb11fb3f0d407eb1921c9c652e0bf1ac96a
za14858f7b8a8d290e835807be677d2f8cdd3cd6c0223c488957be1ce35c62f593d301c031e7733
z37d31bb2483157bb842535bddc2bd51bb940b73e2970b1e2ef34a4e167f348946929fc945b0f13
zb1e5e297735bae84b7afe5773d56fd8cca509c60bafe78ac693845c7fe3f471d02a95c55064ed5
z997cd5dc48cf669259d1d61c5d4f3821a6541e624f29e20b248623a540024484aa1fab8ff2d3a1
z0543e1a4371aa1f1607675c1a4486ffe88a314856b21d91648b91e26c54c171647d37c0b19c3fd
z8e9c64f0869da94cfa9ee4eb342585e7073a82e6c8d649443430986fa8a13269d8ab91b5a28eb1
ze8ae2ac431318a38aca259472d410b4ab84ac3b9762ffb6a9702613d90dd4b2f7f3792e60cdbf5
zff9a3dd02e1fa7184cddeec12e1813f14115d05228fe2de22df2fdf3264965283e149f60cda784
z0c057d1422ba88370f6ce7ba0113e77d259b6abbd8df201a794bb498096a17e98ee5d4e4b400a4
ze961500f51c5d4c436d8e73689bf267528e8d2d16339940855c3fb359b69d511b9bfc6a7ba521e
z6f55a57f946330b14d4c837f4984227b8ab7c17e9e2599d44299841dcb2da35dd03251ca6a8710
zf9648536a91cb1385bf3eef7dc77aaf8ee01f31b245af201adcaa303e387484c5b8797698b17b8
z74114a4929c1d55a5eda6bdc875d548f6c183735ebdcedf5b7f636ce58840a11b451975f3920a1
zfcf97d38c516b7082784856950b27ee253e8f45b5c155f0f3de2a4af33ecf4935035ba1336dd6c
zf743e6a3961dbd2349b4ae8b600c40c86e2233b15876c0c365c8ba62174c0dacaf2081d44ea43e
za8f371ed53a098638f3453f0173d58b85b8d089b611fe2fe5ade6e71c6af0ea286d2d727d9d785
zbb634dc09973fb8e359c2b54381d92f2e07fa75e6b29bd284cdaea989bb23a2723acd627a54e83
z71e276f8addd3813d46a7f42287e6251c02af463ea249b25981bed7c25d8518572acedfd4f9440
zfa2aa91af2ff08ae0f5bac543c2edf0f3f0b80cc7016459e88fcfbc24e6d57641b7adb6529c06b
z896110694befb642491b795f441ffad5b994938049cffc87097f52c484f3eab04abf117f931e80
ze09b61dcc647645d4170951bb6e43ade09c9ae50cf972f6f14980158e705b4c24ffe1e4dcd42da
z9928a58a94a52866844d729fa7266f7a8c83ac3b42a09b97648d507d61b12e4ee1a53001515aa5
zc99fde1b93d27a4f5f1e55982ad59f5a66e37ad4654b43c37efbd902b06f6010d9ca99248c54fe
z886dee7b4d62e0082542cb07fcc4289b2ab71ea5b0893c03919cc08200e344ca39e8d9e8d717e3
z24d201210eab7e3242a23ea10cc1b3cf8fc3e8e8ce3e1731475d97d57afd09ce350937a4539630
zeabf35ab4ad8da753fb7722293432c277ead06aa34285bd21b2f4f0eff29a06c20871217f3a688
z3d149cfdc91a006cc6ca6f91e20cfcfe4a9b8822cf05bc4af08366a87616c2c1c164dfeeddb01c
z38efdebd8f4080de6f26225170f6e05aba1c3879874115b5cfd288dbaa25c166fa480ee6143bd7
zdd68d5bd5a4fcfa69e42755e7a9266b26a5c5c700c8e4104cff0ab8a7d2e6fd3f899e31d0d929d
z6aacc3a716b417671b3265a28ffacee1c70a36d2c324cad3cc9f5a3a095208325848aaee98d3e0
z54eafbf1e6696135ba112d5cdcb7672571fc50f8669676c9e07044b8dbcbcfe1f20536cec5a829
zc92c24b43624f6f2afb51d393763dff97109813219d3a5951529402aec4f16b5a10b3ee09e0ef0
z68b8e1c0b1585956e4cdc4911789d91d1dd8f37626efffce8f2201a7fb6ed148927934b4146f71
z94203ecb872d3c946980c0d4bfeefc407aca7d7854df92560e43527f93dfcccee852781226fbb3
z5892fe042ddcd4753e3e261e89ad2fea17ead210a6ffff7db9e614a8db7fe620ec1dc5966d178e
z0d07ca13413355c636f4d2dd93336903eb76c6736ee8f78006b997d77ca07118daf3093afb71e8
z2a728b225dae7ab531e8fad97b024015b0d9d3ba61324c77896ae7d49f829696c10054561e02d8
zae3293899fa15eb8f327c6f95812e5858faf74b5daa8a8ae31adb5e46ed38feb715811ada18fc0
z0125a51b540396ed9a17081de6398e8449a3693e43ae147eaab36a921aec41686a82e2debf66f4
ze66f27b9eaf8a773d01df0a9afd1f2e88c6c53c68412b1c3f220da68ba51850d989819c47f6257
zf7f6adcaaa2c7c773ac3ce83c8eb39eb86ce8e26d9ab2af005650f40818e3cdbc0387d09bdc4cd
z8f46fd5bae4cfded88bc0a0a8c97245ce9d8abccb440e038a118c2df3144ea0cfb4069296f1aa0
z4822856e62d1d4fc80b8333ebe726b0c85e9df619f94b83ec033d5808b0e24995b0d6449a2aab1
zb2d8f5445a6c99f3a362795c6d79f64247d2a2363361687f52bbae117fbf336250dadf17a4240b
z8658b5c7ba56242fbf8b396514cb07dac8aacaccbc59acfc896af75f772da51b9e1b9988aaba8d
z70383e499ac09f56ce515dc8453d1e4844c8086d26d804b59a51b467a139283fdee7ea556e7a0b
z01e3a0cf97d93c4536decac0ba797f7dd1922ab350b8d70629c45d25597e09e6fa978423448db1
zb11921a5b2caf84d157e13e9a7cceb9bde177b7c3f0cb1aa64c4b9df1d43c851b0777e2990b66c
z4f5a897e7ac6acafa57404519a53d4cbe931babd172c600729e2dfbf4b86784dbaeb3300faa4e0
zb4371d4f703c0d7eb2ffe28a6293115b61cf7a6d2e1e08a1410a8c2986dc45849c800b44fff5f5
zbc01ca255517da0ac9609e9f27edb84899ca0c0f5be8c85daa1159279eacfdc3cfc078ce799cb5
z655bb4eac1e680cef8b2d36efc9028e693c7d6de7453e4583942e5431279c0f10bcce3951019e0
z7bd56198d24df63b16f986c670b1f38c9aa134adc8de41bbb7fa6f61df9d3ea94920b5b8763ad4
zd73191869b410251a2ff42f3316776c474ca60ca2f02656f1b374add8f71c8be1df89a0b102b4e
zf8c6b528bc713b208be031012bb9ec6e16ec9246f4fd5a7de49752b288831b4645781c8c6ec9f3
z14323f2cfe33334bec7b36822d3aa1e1b004d618d9e6df1d4f114e621722d36fd34b6be19ce7d2
zaf28c2a74464d20e8eac9200a4e14b0957fbc65c4e1791408b61fc71bf1744e28b730f10383dc1
z6a848f3d10625db4ba3499daaf8d45dbfe9c78ad4bb46f4984ac134212a152731822f0583c250a
z09c3588d0718b4bea37a03ed38a3e85ff918798692618fcb3873d109c1b2a56d24a2d6dc086f8f
z7a7d99bfde01f8233d3f74a41499d8a683572c4cee644c8993fba908a2bcf2e859156ba872f9b3
z4acc978bce897e18331aebf9d0585b013fd66e8e1cb85790efe9c776b12475d106859eba538deb
z1728c58591fc2e2a2e2d4e0b4a8604f1d197b10d8b1c0aeb1e7df7465c2165d041992a973a3177
z6a45fb9eea26db47547a5f2aa2712e5965a8383a7026c6fb1d3da6d87f2a931c34e8b365305d34
z93288a7e92ae585c933d53aa95a4f831ba0426d611d377886a19c4e9e1fcbb2a09117783f6684d
zeb3d3cc5195cebd745d95a667961f3d6d8444da18cb17bd6e36478c9ef609f5d1d647c25c62135
z3bad49acb7239e1735c0296b7335498a3a7865fcdf60c18723711e856310d7d36201b32b6fe489
zf7f112decbac0f2dca9ad3869fa34b163a8e8205f40212f101caff695dde204d0e7cdac56dc277
z703058b6fedabfa3c1bc07fd3b8cdb6294a87290e8d390599a29e2355a87651b50a341f56b813c
z1d9860bc3bf629540aaef41d95e234e2e54fc7d51873e15f60baf7b14b25ffa28892586d7dcfa3
z0e77d6145be6c032f8dae085fa3436b3e31d7729c50607cda31784bc01c634598d3cc94e813e14
z162c434ee0298d0e5d9ba94e2ee3f47e35aed07551d5339576ef46e3ae8d7a009b4f69e88910bf
z0fb5b3ce1d631bc0e7dfffceb2d109450f97cd6beb77b5d6ac6542c007379bf88d3f2fba1c8d38
zeadf6b8d62e80d8866a300e73530e77a7254a764ed2fa0e53cf41ed08bdf0db19bb9b4a03d3174
z87696181c795a10c7473ab32c6e705b94d4a770fc21cc4ede5bbc9e04cebc2fd6d0cf8bce15f92
z1c782427bda462920d68063de5db8fcaa5f09ac137dc9653eb845fc2f9a2c5bb668ec2f5effc1a
z5def4862e542d9a9de2c23a466beb8a6ccb12b119f5231890aa257e6afbc4aa280d11675b59c94
zb487b208f3e79f4f00b1ec15746b14b0a828f9ca9a503d9e82caeb82741240d7f2ebe624519910
z9e7a3092b4bf0c61467576b957b755e52f37592e4850875aad0ee0147cc338be83a6dc5b2910c3
za9819c417c0c903fa2b360a8df6e9cd1d2365edf83931edc6cbd3a80d91886e1e62c0a9f122707
z484125607cbbbf02437e85d48cd1087c41481cb4b6b471dde5994bae8e0ce46f8a0abfdf06e15a
zf23e934efb954428aeb4fa3ba55e091568512025092d59521acbc06c01bf8a60e2e563b3684a96
z7451384e300a37229979f28a97805e6246f8c9898de3f13706d1edf8754d7ce762b3beb7842300
zb64e5c29764a921a5a61628992724b134071555f2c225f7d622f4d14a61e474bb96069cc3a6b05
z6eeeb76786506f213750c9969f43ed429ae74aa4a8361b123f9fa04e75b52a3b8d9d61eae8cefa
z659633d5900ff1a6a090bee9a85bbc58a08c4145d1dc925e6d621f80c00cc29df2340eac00e471
z0646ae43fd92ea61649d8f3ba8f54e275d7985eec7f354f7ba7c254a9402bcd81d0a841f86b839
zb5995650c1e53e6903cbe7d98d04febf22bf603a3f7d5271dc0f0e721db3f70cda1d57952d05e7
zdac6be304ffd75bba6c0cd61df589565123c1efc3fcfd31e8d340b1deea8ba880fa265a2b09df6
z2608270040e88642eeb3b507d867863229513517acd56e108b3d63bb5abd8391ced555e9f27e9a
z56e0caf5817ba50e41d2948f3fa0c1805c21cadb8f3b15e461188468b4cb517bb188e1d01d8525
z19713ac565a2847164fb845921e86edcfcc30c6c4ae8857feca05d1ed2ac60bc681b58be884456
za4b5092f05024ad678c32e79e87cd68c84fb638af3fd76caba9e7c7166a6c727ddf08aae3da25f
z36841f73e3a8132e354e75882788db33ebc6b5c4d8a8c56a15f84c5a97ffdc5d0fdb5476a3c888
z02d42a80c14a4ae44526c1e0db341c358eda614107bca62b695f4a58cd463a1308d6f41e15e10d
za8e4c2004d0fc291d256db2ccb4857e96e4678c6e26cdaa6e1ea267795cd07910b75c0e6b94d42
zf211b0460b2acbdc04a66b3d1133ebb4de75670be36b915926ed7bb1f4b2e8080eaf916d639716
z00cc28c22e8f69e3dabd78dd0da7a6a9e89a0506d3a834db67f1f85ac174d0b58dcf4212dfb8b2
z567b732f72e69c0929496026f7035cb7348bcc358bdae5f7b5704be0bf836e7b6d4ce76a1728cd
ze20d4fb43a707a1f4886b4621d6aa79ea530785a7092dcf6b8229fcbb1478953aa9915333f4a4e
z5938cd772cf6c3141db25eefb345235e1632c678089d993267272963f4c695c85d1253ea1ed914
z22aeb5dd4e63a2e88834d7b823f0658c6d3b69059977b46512f973a9548c7c76f53035b749cd22
z6608f629e7dc6768647e8f677cbad5cd9f33012a020739d6e5d2ddcad4e7ec3e558dc5d193e0cf
zc0d916fa2d1d2f92ee6d30e5b97333f910c6be73bad90b1ce3695d8e38da67a246ddd7d652d0d3
z28462a1d89f274dcb6f9e040d3172e0173e6a96976e317f0eebc0cff940e529cdd3a775ea7f5cb
z18b652524f666f8790575f83b7d090c2834fbd6bccf4e71f2abdc66b36e1e237d6e4b76e8c5cdc
z397721cc2af303fb96742e56d4fdd2d905474a2e3d771c9ebe2745edf59bc650b73b64a56562b9
z78c3d3331ee82b8126b9ca5169f3931d16a1ce8df0a6350412c501a9579014bdfb520915eb0fbd
z1578ceb4cd8fd5ebfcd43ce1297009d3ec5bf86f722559755b39da2437cf60dc333fe1f7044346
zc63847be0b7847268ce0c8382a8c6c0211787c35b2c66f2dac1cfb98fcda0f2b5e128309201752
z9d300cdd481687c52a75ca25c84e5eb984cc8b269eb1b431780b87da62fdbe406a3a66298b8814
z1731f3954e25c7a12ac76752c102fbf6f66eaf959d57d3f1d5546727dae564fa21f7bd6f0d7e12
z82119198c77a2474e01e3888fc9611a0a39d3f6a60c3d23f659a5c9ecf087cb136dfdce337538c
z1fa35a4deb41410794093be3988752d7e3c79b6fe89e2c279622282afb64e0d223a1b5a794d22d
z38b7225b7ce3f2f578ad85b5244391d87363a925dcee5949c2329d3bc02bb3830e623b53b1aa80
zdaada2ac4eef1012fd40786e642e3e497e33b327e719162b632fb45e84c2d1a6a79b8fe777a3f3
z561d6620ef3f125771def0a027642bf7fa9604ee9a82f4ee4d870cdd6da14dcac1faa30a733583
zd77ce28391f631bcd3a40c6cf5e58389ee11401869f82ecb8a5f452637376412fa103258909621
z516305c40d0b6df0b9611b6757a1694aa4faea45a93a3019be0c947c2c53a5e59ca856e200048c
z9e55b95a3d90ec321960e3f11d9b40def64cc529a397696a249ee33e88a74dd49171c0885f39a3
z2558044c500c7d7ff2f18abfab69ff5b7f1f6794ed5be3ff7613184cc67d778e200a28ccbc709b
z6007ec2dc5dc26dcb3359905928f3128ca0205e4d4270eae3a5d7ba8ddd4508211e1477af3f77b
zcd89d531aedc5a14286542654a05c044832c28188ad65ca858b389058fce2ba5c7e5dcc2659455
z5c411ae9bba1a264e0557523e4ded3edb3e68db83ea661461467d5e386124afcc9d963265de4f9
zef03ea5a4d498359ac0570abc56b1fb3649030908d7bfabac4b981bb8ef255bbae2d928fcce60f
z9f2a8948c6088297d2b18be6618ed529ecaf517f805c839e3b27fa7fbfc4a05b00b19539c25052
za8ea4272b720046bcb9999caf360c984902adef72f422748cd13f835afe2d6df5ff68e793c42b4
zff935673e101b3ffe3d5f2c68d491dd5864bf69e5e14f4b71b43f47126b2752b62260dcd4225bb
z62aea96f374e77ff7d34494117dc04096bd7b079dd9974cc5417bcd1437ce854f0d4d5787b81a6
z0f64d4aaac897b2b61d8ae68b651bd4f86f77b859f5997a56dec7cb84da0b919631956e5c61ae7
z2e3327ed464b11feb6aa7ba4362e858c620cd6ace49d248fa43fa3b1b19eab851d1e2ddb0d6d96
zc867568aa91e9f22afff564d74435599b89cc80ff6abf325c83f39785fa14246f496acf14185c1
z1895294511496010c4eefc2489762002e13aa18a6a158a82580cfc3253c77dce45fb6a02d0b9f3
z02736e6a2fce500da21a981012efa304c7e8c6a68bf03cb31d5e3e54b478a7a9c17f727461cda9
z50e1f4a14df3eeeb87027c580b96370edb237f5a398e83e6e49cdf8434a4b0a004779bd8d0e46c
z0587f46d482479c8c9a81c6ab8f5b83a2bf2bd078f6febbc58f2d3ad3adf492bfdfe000e74e167
z24a4cee551cf5cc9aeddbd4804d2bb5b398fdffbf35e034ab1bf15581fcb72aaab71ac19fc9a42
z7473bf2d4da2f941347e5857c4522f936c2141fcd4de0cab52f0f9b92b4fceb75dd24b67895648
zcc23f0e035f1072c83744ac72a90a145a3553e7575f72d8da5cda5a8372c59aba3a8d88f39490b
z058686751c0269f744e32b9280fd8e6aa3a2712fdad34c08fd589c55b698e46130b8b03cb5ed55
za18a8dadc9cfceeb158d98b1ded4803c0a518c303465189b02a131fbe1024797e5a25c35ad5acb
z036f152a564c7ef266a6503d4a50ef2b13675e79bff8dc7953b45bd8d70d7eaa01b449bf07af9c
z51893a1b51b6d0abc4f9f3596e133f04ab5bfc3bdac6215544a7d580ad56abfc57bca74ba6796b
zc7f87c80168070877f581b7f056d33a68e0113fe2f9689ab41b58dfdef0a4e05faa91323e4591f
ze85029db5f556f78f1d1eaa05f21d056dc5ba0a4f313cd9bbcd89af3def5c91d9fea9134c2e344
zf096435d30cbaa480c61da995ff68ac8475a1e4bad10efbde87e16b8eeeb070b3da29d664a36ef
zf8ad8809e6e989f9b0c8e88fee9e31cfa36dff7d392d79f270e7a0fe364d265a45e0fbc6a3d604
za13f3bec2fc6f9cbb3f7d1e7902aa95e766919d4ed42ce4e5ed621c8a7940e4c489f72a0bc9a9e
zb51835149b0270492a1401d92faacb44b486aa838e9bd0f5d538dfcd18140edf8a14482f167757
z132351ec490106432e5901bc9a0899d9470fdf2d8f59cc68a23c0354e0b7fbb41817748c440a55
zbf3daf5d926e5c3cbd92ec97e311ece0d90362256304c1ccd589c4195c3bf620caf69bee6758fd
z3d74b201347e185ea5453016f905e7b5bdb4dee41b76707261e6377967e358cf15b63cad75718f
zc622628efc6d71b670804a1c0b047838757b045e2cdaf82097e7017fd5b58b3ee7e8f83158f0b8
z9d2d8a97783c8b5f5b56bde3433559489932f57c8cb8ba61ad2076700c8fec7f76e97a38c085a5
za9bf23a706a20ae0d3e597cfd1941a5d4acdc7d78728fc0aaa8563653f36f910c7a8e681cc8e1a
z870650c3a81f2c1db42c631106cf052384cd75844697c0985df0362cafeb6130bf29a01b4e4fa0
z162c729342296a8c5d5611552cd0edffd7bd34793d469221a00eaa4c113fa648c142dd3ac5573d
z5b1e176dbcd9ee2d8196f1eb58252a155cbabce6e394a690e61f4611ffd3dc729538ead093985e
z16ad64acb4cff194b1ef638e4b6686fab639ea2d6bbbdadc90efd754305b33ea2438d1731b3f17
z897b54db380571096d8d8c8b70f50895abba834895cb64de23c6c7544e05aa9b40a2c2ec4320c9
z802de8843ce1c872a6ea8b3d60d192599e6c883d4c1dbf0fd911e1fb2cfabc91f1c8b3f845a712
z2fb57041fd46a97b94f110c087d013ad074dce1a729a0161554dea3d4c9eda48ee9e17494b716e
zcaeccbf31c9a7da9bb557d042fca60266f61cb6ed7fcaea97082c70058e8e304c41a5211f4f9f5
zd748e1932b7ce1de0bcba88c8813e37bec0cbb272b404551c62197f94beaf9b5ecdfba4ca1c3dd
z0529ac2b7f57920259c85edf28d990a7c23f2bcbdd92a4fe196d83d1cc45a9d5059b854bdf8341
z4df9632723a912caa035e4a1e8bcef290cf0d4743a18bc8599b835cddf4414aae18404fa38f3c7
z8a0cdd764a4f6694e7913b919022e380ef48f273a5d81349edc149baeab4ffd1e215d19cdec41c
z705e4109f36f0aada255dc90b494d6f7e2f5a5113d8478a4d064ea235ac2006f291d3d9f749b1a
z502cbf216c526a8b90896a288fd00a1b2d6ee89e8ca210dc2ce26f828023c02f9cc107a9117d1e
zb9c3e4a52bac370c13208ac0adee118f6dac59b9e4281b4cc561096ad88eb1d11e7bf7f5c2de5e
zc1ad72c38d903c45ac6c0ab295b7647a48a0afce06b14080f3cab0b9445c89f48eb1d20aca0650
za05083dd786034bc901161eed18e3de0fca7d801542c5607b5fc4751edd0c47064534a5b542bd5
z08b457bb23220c95d4e1c05d66e736d8b8e3a0f069d47b76d41d4cbd60949cffe6934a3d79b11a
z49297160e2c3ea72a5c59f47b55428fb69fb01c2948ed38ab42e83dface371709a99cd7de560e2
z6eae8d11842c0b06b51e2fc12b6f0b729a9031b7335b92b238f65f3cfb30a09def7c8bceb7039d
z444ea176c772497246e38b3ef4a6a99dda2a1fd7eca68615cd9d5125294e08c0ca51401328b761
zc2aa2e444e83788d8661b5c111be5571ad69c577973a9b3d3d20c598fcb60223213632726cf579
z97f6a8444d076a77c7538180741fee81997c781a6bbd59cf986d564b79acba5912c511d36dead2
zc36cd4459890f10b1675139beaa69679bb20e09015c9e11fc8a6bcf57a6b38188432aaf595b02d
z0b9eb59e932d5c16954ac3d96678a7e938bd31670b4321877b6a22e81d8476d479bd724c49adc9
z740f988af1ee6702d158aff2aec84cfc0e44b916cfe5950ba5c0c065d44c1bb864f39557d920a2
z2bb4c309318051f2d5ce0e8467272703b7e4f3e8223d25511fd11366db8f9fd8b55ebde927b2b9
z4d4ca541e14cae8003385799cc2ff9d7018283e19c415d103537cb073bbe6f7e27c76755cd6266
z0cf6f35a6c6e9c2f60a278461749faf13cdeaec8c65fce4c1a2edd0a2b93d2a280ab12d4cb599b
zd5897703ace4a43f8ae73e631d58bc30c758f7622495e4a4a5b270eb35661e803f37c961650a69
ze81792ede52b518ae17a6a334793728c9c3c63ad0e22c47619a8b80f28be370f3f43b3b653467f
zd5c34f6df90c87c0e76731b727c55a3e79ac1fb414bf35d17c6a977f2ae3399fedddf47af45f5f
zd4334ddd26ec4cc436dc648d0c86daad0c4fc2e529ac674425ae0864512e560dad9d911ff45aec
zf99898f3606cc0831e26eb74520c62f1c2bd4b6c26e9189b6df5da9bd28c196e0d0bc54b40c87f
z85dcc9b33ff2d6f0900c964f5f4d7b2d1f03ba9f17c73adf72f437a2b653feae884470010c0205
za074d97cf1aa78d780ab73e16493493a0eb6d97f5a48f869436f013a8ad4eedec4530ddb6d6ae2
zb71a684655887c60477c10b994bcc5bee94700cc335a4bdbfcb9be151f6b9e5ea8f8e0bd700915
ze865d2a0f7dd68f0f2c993b65bf6417199a1d8c11900d2be6eaaf3b88e477fbe83e3a9e1025ddc
zc2e52466880912b9959994db168a88f4c2d81586d0016ed26691f1026198225a70d5747b664079
z3519c4d2ccbf6ec197d9fa32cc73d04826ac4cc91c03cb3ffd0db50d182cf17e66331e4f41cbd0
z245ecba2d1fafc937f26054085d35c02f572e933099c1f38cd00451965fcf9cc97b0f632d9d263
zae7426fb8120753e4e4ae21e64d5d3eec6a861e28d4514c997eded028e72bd964d407ffbefd537
zfab8c9c30242dae419717f3da79aca0fe13dbf660b3615977971b55dcb034690a78e6dd2b9ea16
ze9352007cbbb7de3c89591ba7368b1f657fb8c014af498d7b32fd98e9461ca52b2e5a2337409c4
z5d20ee59a6855b0245b1e3de06ec4bea03b5e8ae53c47853c947675db93b4f3d1d42aa3b3ec69a
z24b3f695881af8d04b23f11f7aa710bfca196b21bfd1331010c17d20d622023b2d4b1397ed4a1f
z6dcdb06d93a083d253a40e5b4ddbbf070ab2d02242c363182a76b782e93eb87ccf0b5f78ff3155
ze67714306c7204b7d8f6378743feb5b94bd148182b80b65880ce8d30e7f35ac64e07b8f2711565
z80850c5a6b70def95e3b19ee6d65fc872b7748e7f1b2ad19feb5d2841831d1c3078a60eab66360
z7d02e9de0a405b77fb843e371b20fe476e8e182f02b9a30545ea7db195f30d8f7176ff4dc36297
z9f029ab80183b9ff5ecf365b437e0aa1493fdd8a7255bd6d751620369c05e8b50e6547efee5ee7
z9d91d0eab5a1be1745bf0f1dce6c676f777b41e59f322d9981208e76abba4862bf7f7bf73acefe
z4b5543b438ed0e5bc339d88b2f012beff2db0d46b9cbe4e5ae428480cb2137be6457e2c7d8323a
z10ea3562604c4338aec37116ca32cfc686b5615df7d49c680cbbd135700facf248c5d44aeb795d
zf29cbf8ae5b93cd3b247d1e319212da9209c06ea9a79abca7a4a8e9d0a35ede6884e3f3344ea1c
zd16f7e7180b46c676497b78eb804a4316e4ec9232208b4d34a9876e056c6546d732fde2b3f2c53
z5472d52bb3f7bf47ff0fe4aa5b26300eca2a5e0e7edf9e97ccec9af83190d1156f7baad3cd56b6
zf8fa362d410a1ae4bd3e55bdabe320467cdf50d93af36117bed6f78d6621633c6ae7a555527d90
z5ad3f911e212fb90e76099e76052b6848b25bc147f6ebf72c1e008dc85afbcd936ab5676c6d922
z8bd00c32371fcbe36ef2a599b5a80c6d57b7258730ffcae25da7ee05134ad7cbb57a3c496ef132
z3e38a816d496f7a5d2aec2864d899a732b4c5ec8c107663c8ba538b396721179a5ad90e042fc02
z56af14b2367266f852e65bb28aa900b256bea4775fe2b6f9d228e00d03800c456fb4ca6035b65b
z61c864ac6ffd8ef787182df384eb4bcc65a5c25c6390fa2762c4faedecd29d43cdb7eacbaa03ec
z14cd734bc7fc9add3e0fa42643a9ddb2a43cadf5c0be4ae8adff4825706a601b03c3bf82796754
zcfeb414986b176fcda0b0408f228d6979650b200642aeb29a7c6c8294c02ec8d5b6dd999f10300
z6505181e081ae3d233333741a812b159b6abb7bf256aa1478cff5a8a6d8977017f4f1451053ad1
ze16f9d3cd9aa00dc6fe8baf38e4d3c54e82e2885f8f8b1f0b78756281449441dd49b63f5368748
z7207b563f45b3ee7475036c8c88222f5c8783f933e2235505317e8b0dcaa277e65c3be7e57abd0
zf6c3143cb6aa6e2f4e767ba9ad6d2aeaef5c73734c4d9f8f5bfdd8cb7c170a629a09705f91a775
zf3fb32e30af4777027abd0e34d9c54621cee446881f1d264459fee8509942f8eb567059eb8642f
z7471e3006592c3a912cc272b7e375550ae66065893f5c9e9fe35b6565ed435acad8e2259b2831d
zdcdf19b80cd22210136721f74a914b68348e5b31fc20414a0ecb32633059b908b6d640aa13ca77
z0e590973feeb994dd04caf3cf79cc77874dd55f1a604bb6b9fa99f79f35ae8d5a2329cdb53b437
z0b0ea9fcb4ff0c7bfd47335ac96623696bcb57f3057aa328e5f4a7a4737fd125b7a294bc2a2430
zb95d81ce6927140ab5af12d9aef00773f36d9e6edc0186f22ac73537bc002d76b4593143315c23
zf117cdb1b0391ea3f2cad4e3a32bc6eec140c8b6ff2bab0a1f78020b9650ea64854c0020d4327e
z1ba00863d490b77fe1de984362274d9a58636cb1fbbb7d068120a11ff6d8fe14b4a798389b24a4
z9bb262034765f73c10fbee74429595b28288db9b6101d13a282b55509d17890b0a3e4015f9786d
z1ee122487304531c0fef07da7f5ba0a9e03612e3d06bf213a2b278711e968110145ad881711283
z06c1ffe96f3e839794e4ed2d01bc7bb35bbd3cd656dd6dda7fff56e802d734e87bbbec2f55c3f4
z6d4e1a43821f12f7c55228bdf7fc1157a105ace9516c2719b1a71b77f77fdbfc72e22c54a4459e
z9755bbe38ad15dd2d772316472b90e764b8f3139081f0ab2b5bedf726f527f2f16925f39eb0dd3
zbaba8015560dcae0108be7e3951b7f62f63a9fa3c7f32ec086cdf93a53e9a77436ab817dce362d
z9ed854c5d8537eac1478d2a4403fea0806e746831fad90b34eb8fadd8a6ab74ac05dc2352b7c95
zfc6609e81bf88a7b7484029f6960e84ed843800b2aaeacaae767d8bd97e32e222e53175a531f97
z3594a4b03a38e94ab6b1fbd90e205045574fa82c05c3984d007cd58237dad4a9cf11a0db052177
z5f78186427bb12957fd2598ee6d6c53fbdc05f40d7542ff578926a1c7a1cc40e216421876f0f90
zedbb514e98572357ccea7053d75f5621d4beee3f1022214ef038c4289e33a62c07aa57f480fa07
zfbb2a8623e4346feb5eb53165437d5895b58b4e1dada4fe76d7f5cf77c2fb38b3a6737cf135443
z14604f9552d899dacbc8ebc4881aaec3c2eb886596d66cb6dcb4603d11ab982840bd72157c0397
z50f3455739a70be5a1f3c1ddfa24f68a216395bc46abe01b2d2cb9dc5213c44a485fa764a61387
z57986586fe4e4fdc4aafbb611e4faba68c1dfbe20a07e62074c7b9ef0e587e2799e4472aeb9564
za0b6e50ea9b795c6b952d185d671fa4179173911594cc280ecf45013f6bcf73c5b59689d534721
z8cf542edccc0e42c52f3b615ad6c17eeceefdeeb343dbabecfbb90dd8421d6be459e26ea5ef80a
zd3dfb4246b88ddef702191df35dd00e9385cf4d46ca38a44070ae678b0fc1a09bb728a004356c8
zadb730cd86a3af489637a8cd2d67157bf3fa7dcea216236b2b5781db94dafaffcde49ce8605ac4
z19a5004bfe33294b068674d27631e67b10f228260a3f693de5e3b7d56423d9b04202f4fdc89407
zb4da233a54877920581ede1d336cb5b20ac4cf9ea8f9c456774c9f295f5e703cefb3fe309d5a80
z5165556a9689419005485a47ee20bfb00c0b29bb5ec3599e3c9999cc093a4b393381c8c36dc996
z09e1a65d41b2b691b63c31e8664478385a9376e31cac6484e7abe14cbf725cfab0fccfd36a9952
zf31efdceed42cca800cc1aa00f38b9725db1bec315160dfef803fc8a6777dc0b3513a6c077e014
zd3ef9027c27e1a102d44c1beaa6c2acaffbb5490bc45efc645b56cb12294010eb997baad248fb6
zaeaf8d60ff439e7e8637c5a1a24b03a55751c1952a03f2d40bf999bb9f9c0112c6d01bd516dad5
zcf34980ecc1c0b404eb7dc7b646d1e313667b9c42adb0b18059eac88f26926d7b5aed801500d73
zd6bd5e5edc298addf2906e2786933db96779370c9205e7d3d0fe892dfe94032cd78e56ce76f42a
z4a7d62deec112cd0748802ea73974b20a6e2f4e1d70963f4a0c362b6ded43061f33252f1489fbd
z195f3c9183917ad3584a4af6b1791822903a66d2a6f2a654b72c1b7a70237d6d221cd5b5607e9a
z6151ac6d36f0bcec5eac3a5489a74a2f82b8e9ba004d816d76f1589a978a24936016e62e90edf0
zc6a638836ce824c3de202f57923673136034f8420c869c6f9ecec8502a4d0a66c1e1a708d9dd3b
zd3b03196c12e9bc4069cc26329610aab0e26973d342d30825ded75d4233b109d2d7f693ed53998
zf74afd723d252392f7c1d1a074a1db3702ee5671a0f82fd3c5d87fc2d565fdbe0f39cba17a9058
zf5271e66ce1274e37574389c9d121844266b84c0469290cdaf036d4e63e32311ad9a92baef5ebb
za12ed0c8bf9bc7e3817a2a6858d17491a6b4780d11bb3138915841a96ab2d501cbddbfb81148a5
zf85c9fc606a49050a5012b3b0abab7b8980c7605dca088d08d585222258006d7fef421a6e8d075
zc5062b9ca43a15c89cdcd6b3f9a3f2bc65663f52bc8530ac0f5d5e08a98c9f1d4ec4a76af61382
zaf48de91343c4865ae0e8b11ad7d040a584ec5620f1de2904e3e2b1c9cb5476848ccd43e95103a
zd2c1218626d25c90680ee2f26a6d898b3001ac9bf7d4802a31f8d4e2f080a85149c90ef9dd9182
z5ebc1b3e09f8189169ebcc0478bc4ccbfff648b1b0d2985b4bf960eaedc31ff8eda57a58499634
z1bd210cbe720026aab25089a80b4795cb661738c3ba19d5f21169f3d6c9574f1f58468e39b279a
zea5c446fd732058f58e83279caeecb71fee201eeebd483724fb059405e32f69c14794b15c57afe
z814e8408a8bb0c1f9650bfdc02d5f6e6b3491560c0b235cb3d6a92efdae24841159d01780f2947
z41cb5395ed06c9cc3e828ab9e0d0f117641c14982d29099f8da62bac16ee4a19e505d884d1cebe
z1da605e7c7c2d421c5d0948edbdcc3e471ab9a4c096f5a13b074e03b1c6eccb66e4325ba4512df
z3abac02d69640e057331b363b9dbb71ef3fcf955108e01e8cf7f79b6f91dec0c01edc994710e96
z75c2d792adf18383527b20f9a8c82c7e55f0769fbca51762d2087349c17f388e64e07c239fcd7b
zcda25687d20ca68e77cfd3e4100df47c403fb48d148d3b3a43c743adade5c420833201c8dd49fb
z07c9555f9136abc51a399c4695add1fdf98269d7bbcd724bb6293dad336aa1a585d59a7f86557e
z43a6af3ddc46170497ee7ec09e985bab698f753024d76214ffc6c2973f91497c22d0be30b6e078
zebcce9e4747b2a542e1865a5e4a0d089a615cf675f7de645d0572ebacac754a9a185f7cfccf061
zfa7f51b49b6bd86e1c1d60fb0d08e9224e5d490202bd6ffe84334bbd90260e30578e5e256fdc21
ze0ef50aeb5d907dd6d547cd59d5b88adf226650b605b94cc316d797ee374932d7c98afe1979b87
z4b97d7a4dcb99cec7f8036a2bb4e7a06e6915f8157424b8a0f855d71d803b4eb0f221350e346b9
z75f9faadc3dba157904958848752546877f5278f7ff5fddefee4361e5e4d5ee6e243d8e598d15a
z3c78ae9519f8f26aa766f4914139b3f0a629c2d64b3ac89a4b31a7f41f78714e0aeb4c7f224fa6
z9a06f4597ad1914ba9d739c486cafbace1e0f83d52f725586700daf96005dd822c82c38cc4770c
zfd30b1a3e8fcbc6dafecca0589048a22c7e56bbb76ff274c35e810a735adce790fbb58d2a747a7
zc0ce8de8a9c4b26fe69edf0820087e9cf6182be1e49899c56f97af8a853c0369303dd5110f0a13
zc967641bc5da8defddd51a24c616188849a7be49a0dfbdab2a3aad49409a2a5d393cf4e2c4bdb3
z4578739c953a3b2ddcd20d32e5d4ad6e5e6782a33a11bae0660000215dc9ff102fe15242b825d1
z99a065c720d8774070318764be2ae62bf68857d7b154cb47a8d1b995d2a526db7eac65735927a8
z8b52ce03d58ddaaa295d47b9856cf6d8335aa58f13e037cc2b94acafe5771da08d3e5de57d1a3c
zbbb9e79f06ae125ba772ae002ffe3582dc74453927da3fcca607b2391b3979ba5ca3957ec488bf
z1d3fc7d7d74138359d17205ef7156f14df1480413f7d47fdf346919b32e08d4a2fdb441799e950
z13e5e03d8a71b48202d839cb44c18a5997845383f10fa7f42e49efbc19bf8b367039d223a03bb5
z433c3850497d54277f300c3927379f86f7fe657a221f145f84859a453d63c28eab99e7e856fff4
z5ff82f94a9c6722a63d5e41a35c5db7d0cf1485e8437c80cb78cdeae3c3442fbd3200da6a4725a
z40ea7edd1c23cf55b7a5652473b0286cac16c1227d996c3981104a7de1aedbbb8e2aa18a58a29c
z8fde85753e33b7a978bd88e2e27efcd6fbfcffe3c8fa147c55fad2914a31a876d41c34a180e091
z405c6fd76990ffa97d52931b4b0477a47ce336a11534d6d14941650eddb4131326d6f8ef28287f
z7179bc1177cb0f57e48f5eb01349c8c17fb92c47db2088dd41c5ac99df3d195071040165f3a5c3
z2288e5239e2af1b34dc9ca0ecfc9c54a66df19bc6c9776f0cb5fb048fa6e12c7c4e903f309c275
zab8232601e25da2cc14fc6078caefe57e6644960ecd1c4a04043d42542a9f31c7ee48692e75e7b
z827847b7748e23463078801872d2211bee46f1cf4880c4a92d71ff44ca3139e3da28bf87cbe197
z8249df265b17959b8168930e8f25c4349942001c96bcb80c5beba69cc8ebd67bd87daebb6e68cd
z8060c7d416da17a11b1a17da2f879665e29079a4a1a472677cf1485d99f2eb4c2010612e5d007c
z26bc42362594ff777bc994218fffa262d45a03597dc651476295f6ea946db45c2df8508559ce44
zf5dee04e8753a66438b1a7c2abcfd99f3ae9e9b778704ec1598ba6d6a576f0e87e07789060924a
z1075964fdf75e651da63af7488f7ff71351bd02960fb6ca90829549c641fc2eab357af26e0f1ee
za6dafa218adc5651951c6cd08528291438042668b7c852d2dae73b184114889fa69951bfc17004
z7799e8eee8a786f5c4f6fed90eb0be14018e415358c6b837afc0b0aad79f73f9255740e7559d78
z4b31bfe0b338fa468d1d5222a30c9075e79b079efda12bf0530f9cf4e60df39f5ec33c97250fc7
zaca58c5a2566081216a2fe25e6ab390668b681b75e0b77af8cbf9e62c19d36c2938541a117ec7d
z796289a22e00799523c200b3c2332a2742f0850a0779c11851badf1ec5153ab48cff54e1cf8a30
zc8e1a37d1c112bc2872c0f4a0fbed947df6e972d2cc8c90595886d7273fac0549c8033ff983df0
zc57ef2c6ed0381ad8bc9f1f7e86eaf469ef3a041820f4baee9ff6fd183f6ac9290096630f836ae
z4e9d4401b7340cf5c0520cfc6df3a1320208b1720a8dfa25bf20793c1332c6e912c111a066f345
z593e268d6b70f9e574d688143aeb1193b4bd605704ec9c515fea0a4cbb95b5abf5b4e84a8607cd
z3bb53da2fe96bce01da21613e49f570fc8e752fe2cae4fe82b0361a1764d07c4998ae1ff51d6c6
z33b52861b9bb91dd517795c81b9e528f3ee1d41dd05249c07533b15ffc7cdf88a633f4fb5e61fa
z836bfec45bef5c9c1519f26b6df209fdd094ff40e63f1b2f2cad77a5b9cfb966525f32a1a7ef8d
z05167d73ca581fe9f6438a9f9250ec21b35a7edbf636d2595c66b86450160b3df5d345b0ade7e2
zf949809e0471be6f913074e0a49cfccbf5233cead67f3b1e802c3b04fd703508a09c45b940e816
z20da1e6528e55b77a00597c7209717f0904fb78d479453a6aeb6b38d6289ec0340bbc23946544d
zbcee52678953d1b0912f1decea0e83690331dc20bfaca99c4c980d9ff825ac01f512344c9d1cd4
zf2cdfcaeef52dc430e4ea195c641b44e98f3bcff2e8d4e2ba0caafbd52abf9146eb12ad27ccaaf
zd4803fe8870602a3294b212774641d849b5b5ea5b9a971a3ba678159f4a368cf45fbb733fd3ebb
z9274c4ceabbb26811148dc9a2f4fe5a7823d7b74610c6fcf88b602ca9b38e78a4cbae6d61ad21c
zbefea7e3fc3137e56aa5a4256a42c152380cbbb31f5c26105b7fc218e48c5caf5f10457c93d9bd
z8ade305282f0a63ddaaae460a913422af2d7d260e1954333faec525ff57a3df92bd65dc71dede0
z8c72bdad127f4ec8445e0938592f84dd357f9d140c1b282cbaacde2ef2ec1bb07ae2eaad615443
zc123b31666e618b72f3727292f796c5b5267a73f1db72c9da01470385c129174482d0a0ee161d9
z6cd7fa6329bc765b6cf799cd75121043fe2eec1d7a27e0e7d09647c2f13800ad985617c752ae90
z5f693cea5bc440267acd415f125f5146eff20907d879c50ba210b095bd7e5c7dc82cfee6eecc98
z1581bdbcd255fdbe23a7289c3d14814aeec5151cac17d2ff379dd4ed8a35b27519707eea4983a6
zb244f56fef482bb0cf7cfa36a34618af367dd23596499004d360871b13b4e8bed0cfa40b66675a
zaf68cc18b942e41f3b282a778e76d5f0a41a3ac30bfc8e204306f3fe2c61a5ed0ff8d2d1c82c26
z529b16940f5b368ea16c8a9a285a986a039ce214c11c0771f6545691c8082b4f281063be9ed5f0
zf072e8d2c148ddfb84c525d0509b31954aceb3692a9b3b45601951367ecae2c705ed3b83a72065
z617f00539bbff27e6e4a9dc32efe620b9500dc22f7edf6de4aa697f809985fc49f0fbc6aaf07f6
z7b44657b7528e7d2a0f8fdfd182bbd2eed923c5f233068db58b43f2cb5f0637039bd1683c5278d
z3a3aa97203ef8d7252993c7ebe531f4d8900337aa52227aacce471427395a2cd319fb7169a0352
z90fe05538672afdc4e5dee795ca0697a59664a0959932bbc6fb7d80759408988ae7ee0ab78b90b
zbc8ce34229d42860ed7fc5a7ae7b064d4b02ec53a67c97d82a28f3e3f0179fed5209cab5203468
z9426b7867dfdd0de31420d7e5aad111eb5f344c3d8ab4b9eb8ed3a33c5f51952ce47fca9c5de2e
z1348b3ebe84906d1a50ecadf0757d80eb2c2bda847e76d3cb27ba8e342775352ac6218a74b3c79
z04497c913cd6d9b1bc523b470af4bb3fc7100e5b7a262f27fd837dcf3a45541547a3960b8367df
z86a88f3497b9c1982a048bc03a4c7bc8d5de991ca60dd29619fd86ef8004bd2b8048fc025061f1
z25b2e2e71c16cefc63cee91e3fb1fe2bb17fcc855d3b968f91a9e771bb57557509409064a9e643
zc950d5878eb31947a4e3fd42663d6b8568d8de7f06ae8c1bfcf1fba95d7645da3b4047f489deed
z101e0777324df9fabff0785e9f7da3133d401a3e2c6f71c4ace84d662a4afafbbaafbe884faf0b
z3570933301685fe593061e9047c58af9b0adf03266e1b7c66dc70a6d47433109f8abd71e208a66
z0bfa710bcf53d1421b37601db20b45a86e3e204b9f6be0b8760dec7cc8cbbc0c3360f3fb55a234
z10a71e931a043e38f428cd49d4c412aff4254209f2defb4828f203c4043c4d0a3021033f47de85
zd7a099fcc89ef93b6bd84e808fa32b162e826c20181bdb1a18fdddf6c1c33e8050d96fb1b98dcf
ze85df039039683f127a665670cae8bae7fe04f120243c7f2268b45f0fee28a4ef4be3761c44ed4
z358d19a6bca6d650591919a51cffaa7591295c36eec659183733470f327241427cca386dd8d9e3
z75e5336d4bec15a1bf21bc915d2a6cc2d5339748ca76d69b77da5ee644d552c343cbe664854a82
z8603ba24b9b1753fc2912f021be4e838d31aa5ccca00436f0fff0cd688631647371fd83df136e8
zc8b7ba0458309956ef72e1bc0e14806b67b2f13a64c43bb2e0d85e96adb19cc95d558950f352d9
z16f4c3a1fe187f742ad0baf965790e216cc8ec7028d8980e03eb1fceb5f9f95b26094592a7225b
z0a0d8e7fe7a522105de23d8a1534a5330ed98d93607ef468f542b4c9dd973afa399736a91e5603
zbcf5ea94db7691556c0dd4fd1e57b30562813018ae2bcd8e0adf38aa27b323b80e5579a4504276
z91c6879fc2cef340ec3a1b9fcb01c6a3ee021a39436a55b462330b91f3a253cf0f5885871c4cad
zcbfe2630098408e07052f5098df7330c2814b7d78c07a11eb35281442e27c2bdfab143c45e1173
z9c2fa63d6e33fac9a2293d5b49d45d05b4e3f84bf406c2d1d7e2332f9b32ec5adc5fad9411f6a5
zb2464b80fe670910774bc254ee318dc5ccdf7a6e4208a38d18328ccc760d4665721f9afcbedd4d
zb7664858f843ee937255af0b5ccd81edb0ac139cdf62e03447d7ca60cfb873ca7416e1cae3841f
z3620de6f8393efb6a4206e3f2a05e774b56cc1b19691dd4cf51c5f5d7261b7f6a521e5607c7629
zcd60ca25001cf4e505e5def5f6eeca935c6c5dcc2612768d2fa48dadb1a09c8e3ea6c37109ba23
z750292c549512570133609b62bae5e4210a8838ba47739125d619e37c0f794d0e24adb8b8fcf6c
zb676987c2690994c50df170328295c6c5521a9247cdc49e0af83800bb36fbaad2977fe710cb978
zbbd3833edb841666a5c2966aa62dc5564be57b58ed535f37db0c48ccef500099404aa92ce37d09
zc9ecaf8cb5073c7217754f353f9ab980cffa0cfbf0320bd95a78bff257e4b243c9d5fed7bf7527
zec77a56220b4d77298448bbc57f51661f7dfdedb6407a504176d79f8e50202442213725e52e0c2
z7eb82a3a9e227909c656044a99e4e3991fc61455c5532e14658405aa0d43e089a3af0be7e8df17
z83a3d35a46aa2332b2c741c48fe49944778ea9b1bb30d2dca1b4e1af21037c41f3ff143444a02e
z0cc24ff8c29825e43d294da71fba91879f77eecf7da3dd1089a95978b36a00310351af6c0a300d
z8a4a007e309a2ea696b6488f9cc4a723652e5125902c82da5890dbe3cacd63fdba1a2e8a3bebb2
z0f11f83aba74a39101e303e91818df35da8bbe3d17a814c95353a7856c4fe1b4a73225679a6ef7
z386d43161df3efc6e17de844b96f94a6cfaf51d0dc5b52d7358f4b375c6ec1e38a5019d603aa7e
z9e5bfe64a96d974bb01f834334b5e2a82e514af60b81c962c747f02b1f7a36f304081f30c1a867
ze3b8b96c35fa3b16d7ddc7985d4df396ae8fc67c5b5952e5a6372faa4de141feb1aa91fa1d9a86
z6011a3928234baa4dc349544b4b66a39c6ccbdf227117b84f806cc3dce28a2e8baba1890f8f1fb
z104ebf1b7b42753b9acd69d1c3e0e80714a8f3402766d26b7853f8fb5ae65ab992967536abd098
zcf7fb5b89de31c18a9ce1c22c8932573039c359395de896118dfd360ee3e7a204e7dbda447e322
zc4d2f2ce05379c6572a7a341bb90039544a257e720c800d885c8d0118d1fa77f442da9d9bbe920
z88da2eab3a9866cb63a2d2c942632e69edc33506442b37287b0cfcbe45030d8fdc1f7d8fdda835
zd73126900021b1d25b26aa7d136db58fb06f47acd2b83497e190d1cfee281246544b32e1f8404e
zbb38b124df31cd5ed30af954096472e4d281c7e5d6d408cac4826ae16f94e7877dbae8cfea3707
z86b715a97094bb4ce8f3926861c568f6ce7dc10cd1be3fafc19e83fc909cfa4093831b1acc7686
z986ca74ccf26c78673542f1e47f8b92f0269ab8ce2a029a8f4fc60da60ccf9ba3a20b20a9dd84f
z85d38f392ebe7338d2518e49c7d553f170a0e88430b18e3f7b4a0cbe1e2394b8cde8d1cf6d3496
z2f4a4217cc0ab97a5ee3340a411dff45307892d4509b9bb809a45168cfa8575adaf36daa4c393f
z9e4431b7498279f05833084cba037cee2d926c11eb399573fe0076a0a729454bd150065e001ba4
z0d591bc40c7c12aa14e806f2ed64c7450c4a87637e821dd644c94737401a1a29ced29ac668b63f
z76fdaf2ef50f17cb5ef0d7d8005a596e8ec0fdb0748ed03f8e4626a351b79c9fa96d71935e0f1b
zf0bb63ca9ac042c39018e3ba5d4260dee62cb3df55cd7e994092e1c0364b76094cb486b55c4edc
z4b25cb186a000df118bea9fa69dabdd6d12cb4b7773c2344d639618c250c9531687c5bf29e854d
zdd395fa25ea6cd4455d962c5d33ed06f997f0c44687aba79f719dbf6f693f84787b4d879b5d46c
z0a6165dd4ad4962bc7d9d89b33068a92b668230b41221e75b63dd2f3b5409a36fb93925a580e8e
z03f06f8a8d2cd5519e74ea75676cb50bbd15a564e17c1996a8d97e5f133fdb620122b70fd32f8f
z1e64e5a40b68ce0be835f2e2f74a78e5d0c63fc0809d427e1deb754f24644194511d834cea2c98
z1ed5cf76ab1d4a437929e8d2cc34b89b983c02cd005fb2ae87885acd8d09f7f8742f6c679ce516
zdf512498d7bddd57003e2971f71c1ce3f36781c496a05e94546bd789b997ebd4ddb6bdca830174
z91c6cd19349bdb55d0132938e707ad8987aeed675a21a19fe7e890e8ce9047eeedabb3f96d517d
z1bdb7ecb67aed1f1c28280afe8a6dcecd92bb7b59683c6ca0f9fb01397c6b37bdcf561a6172db2
zef35f808a39d0d39ff9b4007e0b8812f949c715c75c330f7ab21e75b1a5849ac399f6b1b80078c
z875b78a857a7a54b065a5e12eac33752e3e1f23561d8ad081ee0c0f45b7510c752fcbfb19f1d11
zac07a50fdc17c714e41782fc936e570802a6d27ee559aa3fb1a1d410e069ddb4bf35ad5440bcf5
ze75449795e6d3faa58098c0a4a432b77f55e715ac117a4fd698fcd7e3aa58275fecfcacb400105
z369b556532f8ce7bc0aed32e0b53d88fec21569d684e8973a6fe6ba8f7a2c5c5f41e4a64adae75
ze6e366f22653b633101f67b5fab820a82fa636bb4c0d48477c9e3c3ef516478f23efc051fad5c3
z4383d655519ca5aeb566f77d7c6adec0de55a9bed396477dac5b7b9e69371a0d54fa8b76341be6
z435099b4c3f90b11e6228f7df42d87ad490a370d072f9ad99fc12f51164de8199f740a5d1a9918
ze034d8907cb0ce5e7cc4e9b15ca1b9210632fb0bf0b3692610be497340ebc82701c226b94b8fc2
z0aea98e5d03bfb15143e55c2e014805fbe3f5e468c6666c4fe33135fca1b02720feff7d60d1254
z3fda41c8b14ddbb0316ab7135b17f96ac56054978495364dcaa2deab7f2be9fe502db36792f086
ze0f9f19fac74ba0ef7aefb115757ebdd969d03c58908164e9785447b1bd80ae8ebe8821e637649
z794e1f248c4e8e0fab1a6fa5d4d12aa3003eb4629fcfdfa7c280b52a63955a2c038f8871cb3c2f
z7904fc4e29a7b972dcd3d1e59d8eb8bba57296b05e9648b6625f7caa7d0026912fd2c854f30162
z17ff5b4169cd88212ddd9e29b682cbb6ed8b19d773407d7c50f515cdd7a984eb354fbb152768e6
z69a352f6950b2adff315b5eb65a000f84d17fbff4a1899cd83c45566b9a2dfd6d6b9c775230ed9
z148e82621aa890335f46885cef13962d220b0c8258535e3e9ee14edb9a590e8fa35509149e8239
z80ba3d20ede26f736dc51e13d9b394e005c6b6a7a5c7bf6d3e2bcce68c50ce057dcd4589f531d0
z3d122c3ec19ae7fec0862cded05284e8f7ae8df512a888c6eb8542895fc56310336f8a9f2690f6
zb03a9ab3b9402ab9089610274918b34e16e38327d0c8dc725c62cafa1e6ea73c36a67f9620fa72
z305a549e4a690a200c62a621a962ec45bb5ce5e6c13c2ec60f73dc2ac76ef20d21be9d1f5ae76e
ze6b40d8dc75b50b203fec1a29186ecaf8be60ab95a6b9ce5ae1899833591dbe8bcd8850cf549a4
z734c0988fc249724e6065a43bffd5c285cd3166e7e8ecad14da4c842aaaed646641aed7f52a1aa
z71ad5debf5d239b62c63ab12fc7c0462fa2e9ee40c1c70c686b4272caf1edb4fcf816be8ed7f24
z4b5e2be57bf065b01fc050675f4a997ad5c661f53730f8c60292bd3d9487fd02cbd40daf3bee5c
z3c2162707a82f0b714112219bf30c0b16c9cc54b975075ec4a8517e871605de6b5305548531d05
z5b27d73d532e21380a929772ffe560dc57257c657f5e204cd1b5cf8b46d517925b2874bc119a83
z935c38875e1ae34a15cc31c1247c7bced612b06506253db6d55dac5344ecb4883be8626f6d48df
zba2446e1542d5f5f0baf638b77c8823111f0cc25db697d45de87f6d156b458a532bf91a3039e2e
zf4673ddeb7983a24f8bf165dfc8d231b9ba5f2b7e60701c6bebad2ccf2596c1443ae73dc39e4cd
zbeda4d0f4451e5bc86be5e4bc6d1d6b880a07aa2685b377910c00860dd4adb989672b83de60490
zde01321641d7db95575d956c478eb3b071579920658c74736da0519e86fdb9ded69393308755d1
z21c0582f8854fcfd4c7e114ce06b252f4488812d4f111825d90a4b34677871094440d8967eff5e
zb6d34e0c17694323dde808cf2f97a2db4ae91cb3cade549ba26f6edaf09bcd6cc1783e11817f65
z3fc3fac89f87918c1e70d2adead9b1f7038dd6f2e44e59cd7407120614b8d9e0c7255aa74c4714
za25d5c1f77020c52cda733dff34ea39adf5e81909a3d0b56cd64c0758b7becd1fb6e08e8f15070
z678600c1605ce060af1e2bdae1fe9111adfa187c378380e2abf1b235e6258ba894eb350bb4d7fc
z3594089c33b127ecf352cc716eef902e420022007ddfd1f93ff454bac5bf46957e2efc94ed4cc8
z298bcfd21d29e435f61f002d904550bba92717a28710163284be0c2b64764383b2bc0b24c74952
z784180ae76a55915e848aa2f5b0d858b69caafb0ef91f44c3467f6b7df13f6a39b01b25242c9cb
z3d1f20faf2e19062bac62fae50c0540cb56dfec48b3963232fcb34604e25565aa38a120ff90339
z502fdc315a4da38f0b137477243767d914949b4fa87ef7569b07f27ea80fae6f7c685f6d6f9958
z18c182c70b36d3445ffe9e6acc20ae762897c84df06b05f3777b1f4b6fe9e959e5bb7372f190e4
za86aed39014cb906018a41dd78958a2e9074c5e02fce95ad6dec019d21b04a1d7ca6364975c616
zbba76bf13dc7058513c448cee68541fc59238a943962fcd2db1cba7b67b784690bdc727cadacfc
z1c67f2faaa493c73207d283417a1804d02fb4eb001132c98b1b769d62dec6042057a0ded4a0a82
z714e4ee2abf4525e13afe2ff4def7e87fa437985f964fb88f8f64225e6ac985d9f3da3e19b13e8
z72b9bf73f2b702e84e1c29743cd26f571096eb9f12e50e7701c7961de9bf4c5401ee77604d7324
z9926970e6aa91a087068f5691df76f7c15277486dca672a7feeda447983fc536cf6ea320c0fd78
zf0656ef594e62318bc8f49268f158a7286156c068d0bcc97de52440171ca4bd3ba4fabe7df26f4
z49b1185071c836dd44681478c3440e30884dd3614d31b075beea4b7a5d3c33769c700e340035cb
z2d488ad3f20eaa6563942ec2ac416335525b36fa3fa3f60dbec93c8cc3c490e449ba3370213101
zac38492ddf887f89c342efb036d6a7a7609ef8d58a607a894e5a9f4cb3b1723a2cecc6c20642ed
z973bd8e8279e6bf7fd9ff17f4d7e742741905bedfbb0d74627194e712f9078f55f75e2b07e1759
z67b53d52505cc784a4da6914d9b6de0fca44a653fca19d22fe4f5c79f7cc04314c91c073a4903d
z32346794ff0b62837751266a481637aed89831b4c64596b120b4883d726ab569f9acddf12d41af
ze038ba0700487c99d3cc8d280a960679b0f0336b18a53ad40c1e73c923a5ed54c3c47fd518007f
z65037384e900d3cadc94184894ee706c7ebec6f8d200647edd0bdbc023281146e5eb667e3809b2
zb0e1d8d9bfbf3809d30d92f610fcd50d0705dce2ff8809b58861881872f1e76ee94a62a0a7c86e
z69d1f1d1697fb906986e3daa8f194ba19192e95367e2476c54db7621cc218fbb73273e26a230b2
zb58b8f415e709da2c0d4b09bf27f3d72f68da06bf3b7250c4a4844a10995795083c5fde8acb749
zfac6b2d55b931b542111718b1f23d7857e3f99c46b90137c1b18bc96f6b24b8d798362ee049cef
z64232b63bc5228514b3d0fd47df40e156e21d3ee96cffc38eb191584f9d7f00f20ee203bdecc33
z2cae1f8b8a7cbbbd3dc6cfff3f0cf6ee2cf94d39e8cd87c630e9c02f2f319a0b62e8c25cca36c2
z1716d59e199c357591ef3631ef9c0e499598da0f9fdb883208c26e7aaa2031518b9b470034ee36
z83e2cdc70e7de86e915e077eac8664a81948ea1baeda35e23ec054a7468fac6134128c22748446
z6a82e10387d16cd9fd0963fb22d7cfad1a998a419a96e4e3cde36c63a15a00ea046a2b2ed70519
z70b4661d39fb51f7ae932680bff947b51b0b2c346085ab6f0c8e07e015f36b2ba45002b163f294
zf98dee38d93d70082625f12c11365a9a9646dccae9407e02dc578be08842ddfe40a4f184bf9a17
zae14c4861b50f4d4586dd3edfe865fe2214c2d3ce20e7d8913ecc0621e988f45294a83d73b3b63
z0f101c52e09335df9f53c3c9af9da172c0109002bfedd7b56fd10036304091558c35b7dbc85f88
ze0d758afc5fcd7d77478883238cb74d867a07121ff0cde676b2b412dddd94f9d103e00498fefb4
z8226a5717c70dc09f807ee694616a708597ed008bb188659be16f937b4371429e643bd1f5a6746
z9d5b6554ee8a898f4d42805601fe2da49e7ccdff7fd3706c2b39529ce9958bab2e7259b8aaa004
z124060a6d78ddf09d86e756437110734e4a8a302a1bbede4b55300433fa91502a683aa190f0221
z7b5071ab5d949967dc4737cbbe5d8f678c0fef4bac02cc8be13838c7a246c9223fd07e7c96f5e7
z1a1e57a760eab7865b94ccf67ec315a5ae4a14d5bc1635df392601a7d35c6481b3f468834c681b
z26fb88493e8ef67e251eeb5845f73a265be43541c98aec9cb20c409edd08fcb7e583261f125efe
z969bba7de863ca01011ce43525a639d7f91b67820126fa03534bcd7d1122525c16f49dd9e90a37
z2562f7656b9271bafbb7f6e6ddcdde34dc0a23be9d0378199c63ebee536ec775c7b961e5862a1f
zb50e1e9808278955ec7db53514f479cefc9cad09b0f467c0801c00a266ae7fc3218df3923814b4
z137cf6465767dcb5489d46c69ab1a6f7f30869b9a4a73ba74d1fb6ca53d5153517b067745e52c2
z98b16365a73775c19b9b7e12a9f22e9ab9859d2dda07d8d8606a3db6e5fffcc93714515e7b0e33
z9a9bceb33b1349484d9090cee3f09c95b9b566b466cdac6ae54094028d2be2d9a784679dd878a7
z745b5d1972e87f3167c1f4e9a6fdd4cc0c13cf452cd34e0aea3bfd8a51679eedcae4e8ca718074
z965fda7175b3bfb39531ca5648fa62a03b72ed8c87307ef7d8800e0f1346db44573883a9fa3044
z4fc8dcf4543f7b36baf9f3464eb96531983c4175be897c0a09eb3a8a73db4131fa53db4a263c6a
z370f9f7a764c2c7e3a2b40c4216d0a5d0099d4ecd78af1a0ef34863c27bc35688ce7ba2d1f5120
z40287294412e4f948daa69b144e72c4ff5a5bb707892a0b5867bc88600d931223cb4a0d40d5d08
z7fa6b997cdcc6af2218a6e35bfe862965ac10424a57ffb542f3f4940370e9c4fa1483f5721b0ec
z89389ba107e493bc62cb40ef40f2bf61bbf38f69ce3bc58ba8fe8db916acf803657b111bb6b739
ze57492fa239fb5c1716129da43262a573238946e0d9612e5ca59bfb8a6e55ffd2fd423c5ee0758
z604d3d0f1435bc592ebe2fe169c691f408704a60d7f0b0c73a6c49848674c1e74eb485ce11d28d
ze59baef168fa58920bf36e53de284af08419b8f42e6c6870bd85063c584d8d527d1f8402446383
z9c597d2dbec968b4fb641b25e7b4f257df3d500d329e392d3bf6c51facfd81e4691b1299d4ff27
zef189825ed5ba2783ccba3a4482dbe9d32f8b74fd38cb830435da071118f1196dd40146320ac4b
zb47aaf0bc2f6bffab0149e65c328d7f67877f6a7686223e4d7085a22e4a8af749dd8ec0684a26d
z6e55e667549f22237a3aa634dd5d26e44fa9ccbb27eb6a611da523547028667253af2843d22314
z7e3dea6d7a8926e81f793967639251863563107252687f4ad7e5da3dd42ecf59af7353d0d79d04
z5b6d9ec0c6e4f40e1aa577190f52e0a6e7251c7beb0adfd0048564dfb9d85f613168344f8bb6c8
zb3a190ca2ca52ac555e45ffe1a81977fff18a59d5c3d116f75029fb3df79c02396519d7bd64fbf
ze8d9ced930d180d835dc1c486fa7041b33314f81e583455919e6dc9cd8216410ba7c218d1df056
z716870cc3cbb5e0f2a3dca5907ac030f77e46220cc500cff205d033ee63a8b4db3177c73dea6ac
z7e838cb621a6e941f632e8d29e786bfc63c487d13dbcedec5378411a8b710f207bc7f8f1506469
zc99fb2f5bd213f6151d61cde1ba05ab6b0ab901ea455fbdebe6cc3bf5e2ceff85c02b81e401b3d
z7055b840042c2e130808bf2f37cad6b9de6e335abcbac94014bb0133bb00505586d76c46795c29
z6c2703f09053667aba33248743d90c909a017a365423b1dc4097fa93946d06aff69903032efc76
z5a1c88edde64b7ebaef0082ba0bcd486359b5414cde60c80f785215571dad390ce5226cc010391
z42771be99ed830d0c2cc53139ae7af760092588bb960490cc460c08de454272c3b159f6ddae516
z45fe8213066083dfe8eda5e0c22cc98be82c6d65ec0eb068fb9fdee43686378dde46a6b803d42f
z11f2a25fd93b3ecc263931eebaa595b28ac6f078b893979bf9b5d5ff8b1e5810e0df1e4dc6557c
z23c7e961832f0080369e2fd23e028b6c5752d8c0ffd8334b9f6f932eb6f8fdf876eb1815de3869
z2ad3f9c5c7228979187eeb86b25897b1c151bd042c80ab185cd9d86eb64ad24fa81786fa480cb0
za007560bef7405232f121cb6b353ef526952304c26cb3b2376b92557982f767e794b2584734e42
za708724aae7580c3d701342c37a39e677a3f7f597c3c4c59d61beae77776108b600f5d3b20162d
z0803cc45167bf865653e3329bd429ab1dcf4b8d06fd675ad87002d3d10fb54416a8288106597bc
z522c7cd6effff898ee2c0f0b5895e479b7ab0652ad981abaa916501dc7fefcd0a0734da4c9fbfe
z1edaa2d0ba0d9acb49a668b843dde2ce2618287601a7a5989396983a02dc7ff632e8766e203db3
z36b5d1168dbf167bd52230fb6ef5960d2efd9e5fd83df2308bd97b0a012b327784921af49326b0
z2971ddac4cd205c2e86355116d7cdcb0d15c95f0b5b4ccb91c6f9bf8d9a7f63416c96ffbd077b3
z41528bd0c3abcdd536dc9dd9c666bcb24c3460c94acd400b4feb6bb7083674dfa3ed4083bf5fb5
z4d5d21bdded5f8ced4f7e110b9d64cf00be823e730834b3f700ba4603414ae130e48a2405765bd
z21e701280469e58c83f54291d31b816f391e550190d45ab07a3533313b07756171fd0566f99124
zb084cf6e7cd9ab4f807fd49d8899b6de528af39a08f03e3c4e891325c5878ab74704b825fa49f3
z1727c62a803536dbe9a63cf3a88e0317addb4936bab48fff3fce7036137b6f05af1041ff740e75
z411e3dbb770808c8cbba3f89f4b2d4e575195d569945e9beb9bf19af8f85658c64b4219afd215f
zd5e477137a5150744bd9e88cf00aeef6b2629b6058ca910106416bbdb8b0536bb0746474903336
zee2b21f6ce3bf00c27d8b894df4754a1ace693e8d5e809a6722db09be6130b297918a763d37ff1
za2bc49a048ab775f5c48f0e487e058fbcd26fa13856399a8021b71ca337a5f30487993e75025b8
ze3e8c621f7b6f8ff8b1561f1de9dfc3932efd26bc4ddc52a16bbc5c98ee5303275b985372fb8bf
zc4092709d063347f030345e16845701c706d41a337055fd6d595297ebf582afcaa4f339025baf0
zd5786cc15fc9323fd5297bc23546a583b6aa03d6af1ae3a73717e4d84bfdd8240549ca5b55ab1b
zb49c6272ef44756e0d57e2dc9cb7ef27fd78f01f1540580fcfdeb035b1d19c49485bd1bd13de3d
z02d2828caf4d576970de153291796c51148e5b8512b2f00db2f9b16ed68c3146bd3983bc831440
zd486e42c3a0039c9add17101f896b32db4da3cd0f92c868ba040df057f78d9339eb3246bcadd86
z380cfcbdac31ca4c964e5a40bab6e4ae1d416f8940358b60cf60551fceb645f89c18d4c8eb510d
z582607bc09f726f9e76bbc354ba0cc64a547ba6cc53e65d5ef26dbb4c05c00da050ad2f5dfaa13
zb9d83a6e15267b1c4cd4c1d99a0567078b976f210f61cc0a163db8e3295237cc12c7f3ddc02e28
zac57966ba8c826538b2aa9e6e088932567e98fff4ba9fc41b2e6d8737a89bb21177d5e60fc6b27
zd8b86fef259629a3f7a8266818b533133b45c494d2621b649e06be840c9c89a9e552a64106d63c
z287629d0b0edd89452edfaa876344c84a9bc8459d281788d81c2d44806dd2f605c7281239f7a50
z5b6a757d690bcff4b36fd52099b67153f947a4d1a816a54392b837b09969544aaebfd28e3026b8
zb4e8f145ae998d5b08ebfa5caa3b4344fbe863af5d5763ad57d5b75a06e06c202bb59489daeb9e
z088c53b4d566589bb764ac60be41f2d49c77f32f34f76e5b24e52a8d3cf2d6d4c2dbd400c56103
zf1d6610f7c272763e5e2b21690c9c7a544154b516a3f13e0197e92589139709477a82a04118958
z0b54a9e9ecfd2b9253607cfaf173690fabb75cdbb54d9500096f0e837041c1bf49a72b1069317d
ze26767e73e665b1d95d6092abae87d66339cd82a1671918208e11c25cf08673a664258374ffd13
z724d0b371bfdbb9fee97fa4cc92ce74909e8b8fce13f027a26be5a34e076e129ca3c4f92cd765e
zbba98bd065ec5dc73161f4ded2abc1b4d40291a3852f51a466db3c075c1a7773ca66f70e326164
zd05b4f47e782a50cca8631371647920483ae272e1dbf0e452e98fdc421dc67d862a7127e466eda
z6a4b3ecf8cd04785496e769715b47419865f7ba924177532f5477def5f3509ebae0bab4003049d
z3026e8144fc20d4c577c0913730d4b340776b3fbb3fd791fb8bf4f2caac375235c8669f5cbb267
z9233c4f01149a73bfb6db337d3f461e53785fe04027356708f500ce719522bb1da7c1a97e68e14
z72a191a5185726caba251c661d56f8a3e1038e83d85add56430c4a1169c2d7574cfe49548623fa
z7ea50f12b7f5d6bb394bb394df9d556ddea9de154229aa49725753cd16811904307947db4ad82b
z8365e3bd348a102dccc840f636913146da806ff23951e9ff814b828af27ee5b0fb44c909419cae
z9e5234fc0db9eac95d8fe2b3dcd2b1a414891156ddf536700fff706f527a6c0c8d9cb323bead51
z7b20537586061c75730d07e89a8922660aef25c7939478aaed176cf7ab88652eea87e87d0e4a19
z1c507f92f6ac2ba93f31714c06304d789e3350d2d72164465d0e8370c10710f68ce7e3ce35b975
z07ed8b6eca958f11ee4add9705eead08fd612d2f32638b8e3b431469c19904f98c6e0399119fd3
z44228c456d3664b9732f400ed086dd827aaa11194d8431577c483ecbcbb6ee083648021ba0956d
z512653b57654f11f7990097417e2c27feb1168e043b599a422589a3e8fb54de665d38c411ef2ee
z51d50427eb0ff0b78705c0d43ea13778c3e45f4b96cf69775aa4d70d043e8ced730f07de3998d5
z70cc188b58f8c7b75e5f168c2bc79127933589bbb268f18e9e7569ba1a2afa2b144f7e1bf6682f
z948c0e4aa7991444d02160f0281ef2972377d6bfffa793116e6c017d0d9685bb821f543d38466f
z57b35c62e0c2801084c982c242a5f1cc703666e554b51a23d86ca480d5ba19aa9ecac1fee442b8
zcd3129802943fb7d1770bef2497b867f7a1bf6d9e434d51b9ea446edee63b602ee7362ccca7333
zeb277b2fec7e7e2ff56f85f9befd0f7b7d3b616a5a5edfc90d618fa4af310dad14896ea404d77b
z498514da77080cd74503de94f84b3676b063ad460c6c221c8a75d618334c386dac186e3fb06ad5
z9f48b405e2f7dd6b9ed879583d9fdc1795b0beec4a99fe6a5fb23b95e2216c7382a4d6e3823ba2
zb3830f2d39c9eca87353e6a6007fef1d672b1c450ac40edc726963e5512660fc87b9fda2d0b52d
z500395014e95e3e4927c99b36c2ce2399580239be5979a559fab5ebcd4744c83cddbf29956dd08
z2efeb9b98d4d996702e4a046a00585b58f00ff89c612450008ba806c70a1d1607db4e90131f081
z29c410fd2deb164fd944391b4d9e996ec313c41e5543bcbb35ce5acf03de8920cec949b36884fe
z62b819ab84b4b721a8030111b6db60b52716dd3f29d9db20d166f766d2588826276fb9aeaf9601
zee9358a158521be1a5ff5b949e13e8b2b19eba550e16bc4ddbfd3793dfbdadfd663b7ff601b302
z825f01680f5174567ac69e11de7c8a83bb2c08c47d2101a6bd2e909adf96950ae1d300b6da17a2
z1f50ffddaea5fc3a936d316e52fc393b1c626197e0eb86b5a8b3f44a8aec8707ae57d77ab889ca
zb82269dd52bdde1549471ca00c8079aaf82ffd4f247cb1511aeca022f3a5db09c4bf9243b6e210
z4f529ac8fad539dbcfe65e021d5765aace63ed999911b7d880dcb8d720f7d3bf7629f87893a9d1
zbcc6b4497fa62aaa7877396a34730a90836044a47b4883d5cf8a8a3c604ced13d100931bda612d
z4f491710b3ab743aaffa21d022ab05c14f405f19272d184fd1d14ec548e2a5daaad44b44dbd5b8
z31e7c1a38badaf31e43db34c4d37770c8e54a302196ebfc945e21400693021aecf626f3600c864
zc6bb649d3ff332ad8d759219870d6fa77e4eb07dc571505c719b1e270a4e44b35f2bd702aec0fd
z4d2e6fbf822a6a4c25917a63f254083bfde66cee94b08fb91562951bad7f83ad77e8fa40294c02
zc598a44de373c155b01e14c859f481c7ada30e46fb3ca55679e52860453aade9cab545a5401ea1
z4351a1242896ea3b96219c27a4b9e62fbfdc484361d716fd114b2955be6bba97b53d8f6e651ba4
zf03b05cfd20dd8b16151eda5d0273ddc9d61d338116817d00547118ded299effc96d1735e28a4d
z74bbb4b8ca53f977b20424abd979d0cb711c0e1b340cc60bf87c677ce0ffc4dd932d06e51feb2f
z1e12edce4a48e4a19983b03980bce5d2636dfbed70660094cb23d2d0f41c62b90291c19f6dca5f
z3c735397e7c833fa3be2d7afa4dc809d4a1a4237e70c99c7e8ee67d421faf1854356111fffc8fa
z48faa36596acc0508b7d46d34f74d1d0e11caec8d88ff37800d9adca1875c79a8869fe6589b1c4
z9cd797a3be1dfa416f3de3fc569ae8c65993c32c5705139f41ad4f8f3a159ec9ecbe51c5340671
zc9b2fa9f7b389f54e47a44622270b10182a43e657736f6f654380f1886553494f4e4e17e9625ac
ze221da411cdd9d88c8ef92304523fe515e877b7f80b70590f4fa430a56d95a22ccfa4d17d21bb7
z4ad0510684587d866dcdd2c02a93c3bf5eae2f9293294e9f2d86227fff58d7e59e2aa66a872b14
z10fbe22175a85c57350f6e54e2aabf3ebd6ceed18833f5b2887dc305afa4f2bce5ea75298537d5
z2886682205a117160ef185502b5154235f18a13e5a5c2b4863f479533992038c201d72f75bbf86
z6286d1c823b9c2dfff9d4f4aa523f02f8c0e43b207dcefbfb00780ebe73e0325b41f6b230c4ae5
za7e4796e6ce06956d3c48d932619c5e8021ad52ee656fbea284a8561d621e445dbe6a5a65d39b6
z34e40b07b62a6689db611de815b0825ff3d82cf9c2b63ad1eaccad91edec4487093cada1ce0f1d
z158971c954140eb3d4d4577649fe773acd55f46d3de32f49b9cba39a48b79d797740e4ec8456d9
z384befddddeba67110761fa92c41122faa6f91afff56dffffb84f9ed041ff803191ffc8a3a3e5e
zfb6bcbf057a64a0062e9472f656abdfea1a639864ea5a2adabdac4ef68e10a1b7c469498785944
ze048975bf2d965e5d7e43da13fc88f45f74fb9354ed17925483fc0753d26265b05177de48b00eb
z773e972364af6b07ac4e5ae3f6051312b9302c7aa40a7a7f61d0e286acea2255a89b14d5de6d0b
z3947d9a5e93c28f68713eae21682291cf8d5b104b59db97ca55f83ce81814cc7f70f5f18d5213d
z80ae65d69c2e08e4e54fd72c8d2c70f485a010e3ba7d6252b571b210b590475d8e8a3734dc8fb5
z056ad2bb315110a72ea9e0ab041507b1a947baf0541a3ae087dbfaddae3c3f9494b3f17079e72e
z423d7165b5b9a4d24406487cf21faa3e01cd4c123a31a4495a72bb15e76a775042b4852e0f1210
z66a0a74e020ed05ce862e65f720ca258bbfe6eba095485ab082d4cfd107117d1ecbdd50d3617b2
zf4dd6c87bfca805b325f3a0a7cffb0142fcdcb30bc69ed004742d169237e444c0fcfe1f6d9bda1
zce3ac37806d66bf718b6827ff5032914af0d23236d7b91a057ffcc57f0e8fbb40be3743e2f8fa4
z24e16c76cd6b34dffc492e39e98d72c40fe1de1603d0be9e58da2c6fdceea0c08c5a4c48137412
z6ef53df871c751d205946ee23e2c073020e7ee0209914607e9d0c41660a2544ca21aeb0a5e993c
zbf205b9fc33dc76eb4b18a14226b3319f23202b4d2cba4f3fdd53c51f8196dbcf80396ff6a7724
z2bb88380a210e8c918d943df4a9c1de2155d3423801fea21e10bb235173bdd2ef69acb2e419b40
z27c23f4fd17383ba3df1bc97cfe3f76a90776a8e824a5d35ecced40ffbf6c17e7096ebe590846f
ze51e35b8c9121f407490e7d1568d8c1e9e2f9caa8b4476100702ce2caa8307e7c542b604b15712
z1988c70f94157a5c67fa53045ab2b6c6cd51205c34075e85ea61190fb7d2becfc90eea0da8c579
za6fa38df3af3850f9c2bfa8a29d4ceaed30997231f21bd21c497a7292368d06805a922783a813e
zc1c8d3a23cb48d95ac9bce1f5e9704664f48722adb5a5a89b6edefb6a26dc9cfc4a1b4cb9eae85
za065d490b2f58656e1d827bb2bee40bf63f68b4979ad6376d80351a197d87f896989af00cf5111
z7b66e375e0407cda0ac5497437315a4a939279ad47bb06c8815a14b0ef73728b538362a557793e
z6e8fd83f023b75074248a7dd16cb510530c52e9b0c7b0fe177368639a5ed9768ca6e9be5386c5c
z2f73f8d53314b9edeb0949171cba12472384478d31c7ab99b7e308b948fb205a870b236ed24077
z3a79d5d2053ff29b9fbcf021c03c87b0390fcb159417f471bdc6a25201fbf7933ecc4bc0ec3a4a
z6cd820dbc9feb318d323c2e4c76f4a382b2e4f23463912c47cfe7874d283b5d0fe763ee2d3153f
z155368fa6518990dfd8effabaef62b333ca901a92a8109b807fa24f627e9a9851587b3d5744ac5
zcdaeab38f251bae9e6d4a6816f53e6e33c2376af336d3e347ba5e804a24038a2da74ce45137745
zb205f62a96d8f9798a1009ab71f095fe563f47b10d3bd17601f85885f637e8827d188f4a8b5479
zb3528be6dec416ed9785c46fa20e00748bb269775e91594350759cb558e9a598e11e5d8f4955a4
z24b8240454ddcc6aced8d9da98eea7c70117b6c3788700a6001f7c57620d56be5dcd4020d42b22
zde70d41586c321ac2e9347ec213bc4aa689dffe5b15db7f5db68b79fc88b38a23b84068ee02c66
z03ad7f33ee2bd6f02d3231364f546422b1f57e9fc6ac31ffb60e346e808abec26bb63bec843e36
z638884a84c3e928fa4974bd839097e2b898c97707d7e231d6aa07048b99532b41dc6f6fe47da8a
z059c1e71fce8d2a2860489faddb02a7c8357d668ad049a0d6968bb0a4681f2c0a477dc05887337
z9babb5bfd0cdcad53cad1316c6e421bec3db77e462fc139b8fe694b770f03e6d01c8ac47bb0bcf
z57037e4ae2f2bea5ab76c3c395edad065c6eef0b206cd68d13edf9d06042e57492376ef7e25bd6
z3c9a8edcdaf350cc2dbf7b44adfa307c7c3c066d2b56b6a0c070cb409d8ee6a9ff385fd89c1ac3
zdd32f413badd2999d07af088e5cbb07c714ade9b748f20f49fa5f0d20dc750b20925046f4381eb
z2f9acd77c46af38c9d1cc20fec0dba4308aef88779f58ea80aa26349bd4242737f1867176ef760
z0749eba4b0239d8ff3d9f9e0c3f79de26fe8dca4e5c8991eb7b21ce173bfc77009a32629f375ce
zcb097ea67eaeb06b8739f419986b693e7bfd68c26ae95320d13faa84ae170419c64a8ae18ff420
z90c1adba681cd9a4537ac51597779912f561a66cc3d9e634a904082568a02c1587f68bbb11b1a5
zc5e64fd6fc1502a37b5377e8fbfff8f5a9a347247fd3cee117211350887fabb0790a28a98ca20a
z991957dff4042b9bc30884bd9a3e807628472c3b233f02afd5ee56e87202292243351f0b50a579
z8bff491bca994a224d4169a4eeb7759af6c873c0b4fd9e424eb584fdc806104536bb1293769b50
zf7f37c184fcf856ce87de8dd16f50e2b4fe6c26184455568a8b69829407ce43d77eaf3c751abef
za4e6abb0d89f8534fd3146a6519a0755c91a236ef886c879a0a34c05f0ee026676f959d40ea32c
z3d00ff22da33dd1589c31becd591b7db26facae9bf42783ca869b057998c9f69532c047cfcda2a
zc524ab017b1bafb5c4386b39284f5bd5152c199e6862e4cde959c652522420a801046baf415aea
zdfba42526136683169c925e55ed63caf84ca1a0f66218174dedfcd6eccbdf0fc8008a51f3eab1e
zd21fe3825be8a5c966990aae702a856abc4d95b0dd4b6edb03ad1bf665e66d68fa6b3f34031869
z51797a5aa90366373180f0d07cecda1cd1d83eb3b313c68c07cf552fbfb3e9565ee50ae58c4012
zb0f601713367be97ecee53f411a153ba8a5b69e635eb95dbfe51b2a3f1b293ed897f704f0ea145
z5f85d450d9ee1c74e0b4f81d65204a7956028cbb8c3fc86e757d653e3f0309a5b060b8717d246a
z5dd9a6479bf3ffa4dbc109263a2d1375f01853ffda1ef19f4e57260483f0e03022c70523741420
ze2729912b34b344f44d2916cd2592f08b1e8f66ce921e9f225290f1ccc181f93804498303687ae
z5b9f0b39c9da4a5fa41fdcac73dc611f73bbfbc1b7402ef376e7f1289ca7df3f24a4d173f8bd13
z4c58b813c23da032cb1dec71637c529f3f40576eedaec42ef0e53d665f81bec702ddc800e1bf64
z8309919cce1449316333b765209bae7b34cf6589cc9b113907fccdf61ac4a7b4ccdf5da235ecfe
zf402d1ab153a12ae43b9753a12aa9aace55de4cd8ec8f8516180d69e9b5a80865ec4c5dead7ab4
z99ff8b030c1284262ab11d03c192fdb69bbc45cb87179ff32672a8d808ef31a0f4e7514276f72f
zbf471a05a41a8a73f82d992b1272a9d0317b2f93d03388b2d04382f9e375baf5a9ad37653ac7f7
z771c9fde1f51f5451c23dfaa6a1c866500640a8b830c9c8ddb2467b16575d9a6895181b21bc582
zcd9715b17abca8bc116973305c3b4ca431d563da39edc391497efa12d9bf798e9552bf12229a3a
z8965d8d5a7d7dd141b72bfff5a5e9757848391ccc1648957b67685aa361f239e1855ece4b73168
z2d8c12e616dbcbe76f28ba8bb206b1a3c2115e845b8099140a3ef688b4e3293ba578c67949ea85
zf2a419f320052da096122be06258b0a24bbc305ce305ee858ba71be6881d2fc81b53c45695efbe
ze5949c5cf8567adbfb8b3ce294936f1e3115d9e4722fb108dabb0fa7ad077737e4ac273c95a92e
zcd5629b1a588b4f5f573b97ec237d0856eed0edd3c4d6a5c01bec03b69ed74f6f3c4be878d6da8
z5c085ab25642bdd76a354089c70ce0cd6df7ea3da773c693747c76a5017208af37af60711718ff
z7dc1ab7a353e44b78c69b1a4bfce5d16e378d2cb142b0ab59e42f4bb0bafd90af40f8414207ece
zc7dfa62e099dd2a471505f576f4d442485fb13884dbebb2449d1b7efc2c2ba102e530953bcb320
ze5f555d2fb55181f9de247852f26aade0c829edc04464dfee60e8e4ce62638b04cd6c125b723e1
z63da70a8367356b06891c370ed56244b8da010cc2228ef590d59455b2e4f2b76a4e5f5f0fe71ac
z472d965f797439d7f09d967cb7d2ed14da99b4bd438293470cdd5435f8a63f2ae1adb7dff9863a
ze344ac41a6eff03ea3430e9d417d40fd955a28662ce8edf88943508bfee6aec025bbe28996e3c2
z764be0a7b8ae8bbd18266bc72979818b5fe8902f17e7458ca447793de9a72ea52bff5ce953dd14
zf4874597ba580ebe06157719e097fd5b6bdb64cbf3a34cf1fb2bdffb33e0a8d7fc24f758546802
zdab5ddde33dba6dee53aa707123263a1eaa0bf0ae5e5877f7eb162c397007682d620bad9477ca1
z08a03450fd39bb4abf1d4badbac4041cff00006c76b01fb8944fc8e250a37c74944fa0624f0114
ze458f1392a344bf3e78110acc8057bc3a031c37c977e115c3194f747644e27a41d188dc02d490b
z98bcb967bf3238bce625b494de727496dade1778b14f4e40dd85d0e246f36c13e7af70e74a850a
zb4f6cc2b4f5fa1a411519b404744e5250d599ebcc8ad3c01350ba62765a760471d0fcd18a62ca2
zbc046d0147a22b29fa802154cf3d59b644dae01b2987587fbfe3ee5be0cd2bcb904ec63374d523
z5c89bd77eb736aa2dc65d02f29d64f3cf0ae1235dd2cdfd754f39e4dbe04bd9eaff82632a16a8e
z18bf1d8264d0f7937ca33d67ea49e7589e6814a4ba4855e7357067afe89dcfc185aea55b0bd10a
zf60a7ebd6d10b9def85d810303603b50cb90f215f1d723a4170f62a1b4d8ab33c54fabca59888a
z4b3172660995ad4caed707bd1e69e67068ed582c632f2f19d5c2942e54fda1d4319e7d3905df29
z04fa70c009d76bdb20d782e1ccad608c05504ecf9e9c2577178df15a521b12f333eebad7544a1e
z9bbac3ff5c1b63188a12f2551c6135446041d785ab491756b4a3ead6475fbaa6bbe2ec656b4bf9
z2f1e3268f15acec9005edf7a318875400a17d7ff8cfd826f34ba982743659ed32679bd26f39532
ze23066640203cfbe101c58b9f6900435dbbba45704a3bcba9b21f2a80eceea8fa93b4cb70a8d96
z5a7a435708383454b7d9c769a2e45a4c098728f45bd47cbf5c303f83d57a74adaf0dc9968c076b
zffb0cb950dbce7d35aa041ecc920b5f1f714fdfe3aec58f87500b28d37abb9d9278445ed64ebea
z73243313d01605713911107ec622ca1b0b6195c7d1ff4986fcdf3ba81ef3bf0882831609630b75
z485ae48ff1305ae129d926b5357607c74ca0e0ceaafa2dd57f3fccd76efc7d9bb77916bcc2ef6d
z18c7b1d251dbd5f3d80cbb89d6cf70163817d5f92c070977faf13996a39ba9f3006f2e745eb1d9
z16dc5936202624b83dcebf7f769a6e8f6494c834fe246e56b840e26bc5dde02237f2bfaa5db7cf
zf9e891822f0e51dee5b1361bd7c8a936c05b1e486c7ed7ec843d78dd03ea495ad775fb35302669
zfbdb5d544dc296f70007565901d1a52080437c6e719e884e41360e7df9de47722ff58b49d156fd
z27f9d9c599e5f6b99d2ba8a6192886074c059516fadeee597dbbea8e83cf7d65ea87be24e09b66
z96ee1bda2f39a6bff2f27e8aa41b28bb9132c997975bbce1da690be2d2db8c7e88150af6a9250b
z4f896278c3ee117541dd2073d775f8b32647bae1c43403a55234b192dcfd671cf6678dc8362d19
z8795ee7429e72c7787f9015db0a3b058aa8bb74a98d4907388e94c3a5cf864060ed6c1b10572f0
z3790a9429f239f1812d2c2ce50cc4b37154f080a848b3aa3739512a0a044ba7ef64b389c9eec26
zca2dec5ce6818e560788b2f9b97a55fc31e295859cd65b0824de6821e8e771aa9b025b094f6799
zb403973997a6b1af6e8e0bee1427336d89e30ba721cfd31138f1243842e0a5c42755dd1a2b32f7
ze9f665d8042d33a17c5bcae985f155bf1964f8aba14419e81c402f6bc87570346028aef6bb7df5
zc99ac7f2208ac20e5f7cc7e745294545ef2f452fd320685f954a0a1d11c209730245302ef6c8a8
z1bf54d20da6238c569078da5cd45100d51b67bcf8f61fc49c8b8297ac3bb9c1a0158945180e16c
zec29addde33e10a79b0518401626d97ac5315d274da079c666d21c455e8e0c249bb57c431b2fdb
z3d585c39a400086d9a2bdf9e4d396882b9d42640be875e854dd3d9898223d7135bad04640f69d8
zc05090de822038e7f221166acbe16a24ba6e51fd772aa9d208dc89ea97f7b0722272976edf86f3
z5b29651566d50dc96b95929678912cbe197b4e8217e2e72006f096e8ea0c5c8568d25032bae806
zbd32ef024a2046fff1b86c6b2bfa6115deee4cb36599e91f3ec632619b4a84e506a17f4035e16e
zb130ce04ac70ad6ee0481bdd903f0d8ad6728c7993bf674249a9d4e9fdd801c781ba19c90adb68
z42ccf2fd53e68946e4e2b0fd17aa3f9a74be01328e6804892db51b4086c249706dbb6a002bd607
zd9473a4584da3b901a41d700369af8b71357019355450a9c997c296683c68ca9848ad1a8be7392
za616e471c52f2e70f12605cc8f87e591112e67c7656c4e2245dba873b618c85f2be13814e122e1
zcc99652e22dccd28eb22dceac8ae52b3a2249947807b933410aca9916e57b2540b64b845ca1a2f
z9d74d883ce51237b6bd507e4f3ea2c0d15ae60144537957ff4849e5250c297cb91d45a6d85e39b
z489e711e072489acbe65d739eda2524af164f6389ec5b2feeb3ff04fdf9dfcfdfe40027288baa9
z280804755f9ed3b3109d0150cdc61d8e10b9995bb1499c2a9149982083a381fe9ceaab048745c7
zff6a312f47c47b234de6fcea8c8550fb6672c166723c981969bdd96b11802aab571a2b62c7ac10
zecc78eeba0cae96ae02b9eda5dd99f0c98e87f0d14f5e9e20261528ae2c54fffb969d1d8471e04
z1b423a99107c6b4979d281c6c5500a99c7d225ef29d1b250f1e484d4735b4fe66888b9c92ff65d
z73780b88b87e650ab52a79d5334e2dd92e111be1196dd1a3ecaea44f4202729a9443063ecfba1c
z929b440e5fa23b5f972eb128132f90416a0d2b7bdc45a1011a198e5a65f933543a27c9d5a4940b
z08ee95a4ad2eabc3cc3f566bb4c132988b01eaa986081572a527624a4e817fc57ce21edb9f26a2
zc3cc1f230100ac84c2f54d5034ff39c1a4d3add649fa42867bbc5fc8f4e0fb20339b49ca16c602
z4659597441ba5bdec103e3b3ed58376cad18243a2a3ced7b836fc6d93c023be211037c9af47a4b
z3df9d75f644c85fd8f5a81c95fd4792cab882899d7e45efbacd42a902f9fd1fff715e132ed8c6f
z26bc50930bc54ea69a2473f1e8a5d487de5d77f580bc01238d722efc0273f1880a9193f7fd9115
z9fceb626f4b2483744ba99d2e41aa75f01f5afe49c2df9629c5ee4a7d6578bb032cfd4ca671a4c
zbe4ba371affc2ea8a2a0e39d1570f5f89d427553a2cddcb6464f2c2a41a481733cefae9ccbbaf9
z8f2ea261ecec92efe4f9f5866b50233590df9b62ed045a0f0153bbb1c9c548f185eb0d142180bf
z4cae0c6b36e1f4a8c4c8ff7e8f7991354b74a8133612eb50ff1be2c821117e7ae530506ceb31ba
z796337710bca10db7a8b1ebb9f535c21fb9205aeeac3f8a777b9c5b4947af94d1f8d0a35651a29
zf120c3810407de21ac2d46dfdf62600c62d4c1c98d32482ec49095c5a9f176e5da7e3e1b8d76fc
za681ef841c4f9b17d799f69a4e5726f19597eef401c4aa01576860605d0bcb09a138ffb2b78028
z12a0d4a204e3277f90ae6b3b1846c7b9b4e13d013012c9fc94aa7979ec0a4c8af2f9da4a6c71a2
z3e3ed19b0f47cd0f5d1850c5fe7f67ac38db99961340ec778059c15340f8033f49309a60a17bd4
z6544c8e0879710fdf0ae83f5f571e28b192973799d69dfae27a9c8d06ff2cda8e2445199117ce5
z57065c3b6b0f65d43a5f52fe7771470b3ad31ccab883fba9d3d0ac786958196daab3e46bd22bd2
z7063e34539636bda37751d516f2ed66b9bcec834842bee74fdcebb838b18bcb960bbc6f5a3dea6
z0e9c2eb3caa724c3cbb9c77f582616e77129d52e1dc342464f6cf3c7301edebbf5022f5bdde19e
zf359f31249253b97b3d43bab5e020077024627c50325701cc497b88bb9968d966242c49c6de275
z28897d3c02251d3495e3b6a79a19c77d7b6b976fed6a7fa4f8c763b80ebcc7cf400623c22c5682
zf6aa426bb0d9cb8c7207469e87a7b3f4350f7533aea590e0e5a0a0823b39c5dc63a7d7286fc1a8
z1565bc5b35041253c512c4ac98c87c77e16324ac1fc5e3c55e622f49b68bcf699b4498a2791a25
zdd0431cb4bdc5d92c53fdcbb7793085cd7b198938a670b4c13f33b22830adeb98e594d99283fb4
zdbe1cb850fbf9081d455dd962398bfe2b45555c8f9466bd16097ab5f6f0bb6f2872e75ddaec04c
z9e77e49bc9c47a60b7f73a1d3f99b44515ef8c5fc69aac5d9ca644704bd02f8493adedf09e8f26
z5cc39bcb322d5b47b2a4b3bcb48a00ce15871dabd30233e3dffef19c076da45dd381a6f0b856c3
zf669d02754cfa5bf9b58a05766095705807327afcd758c58a0fd35308f24849e181bdea1ea6abb
z36fed06f5e313a5e2646170ffdac926f9c6fce1a850bc6037f011f18e6aa2ea982e886f2bb22bb
zd1c9cde92d2aab0c0b315043f9a211c46e8cbd1a5671ab51693c0769f99f44904d79f7fed5f29e
z0d03135e8bc61581c4e527ef95ccf7560e91ed6c335668724b11bd2014823f07194ada9d8ed2a3
z996419eb1c50ac323d4f6b3c754e290b4fa258f84e3c798d02d0c95fe4d02185e489fe20e43aac
z4dbad90f6a644ddaf664c97902140e1dd52e13181668f82f2924ce30574715aad0eda217d83ecd
z92aac5c5664f1b8253134247b6d2824ae2694246f5a41862f4d50b79039f126fc6688ff4f16c40
z6dd18a1f71dcc28eea08e927482e96083699d950f3ebe2e31c2c7c42d417f8b519e8d624b3e1f5
z0424334d0c3dd28e85ad7cae171eb7b2aeda2c75704864dd8949405ab63465a2e7c374b1339d45
zda52e04af40f227885ec9ffbc3abb50ed13e48c0fc72d08c3d011300396b715d4a956b9bda3b95
zeabdafcbcb3206993a886ba97a97833e559057dd249d5052f7dd1ba687ee821d45007f216f9fe0
zae6a991c394ba6b61b1c871ed95fbf8116c6757d4a4759d0d2d4c2faf0cbc6bac7db98189b1ddd
z713f44cfd225708e8d12432ab2d0393babe6f98907db87aca4acee3c22ad8260691ea3d4464640
z9c1f6efd9904669aef15c2b7aced06b6ce824b815f249b13d5db2eaa2f73538679a0285b08ed99
zb6440b1e2a2997929515565a298b73c8bdd38f3487d75fee3865fab4da7626d2965d8096a47fc7
zed81dd8812e17bb1c7c7dcfd36d048da4d93b26fb2fcbbdf25182c2bf60d01a3554cc35aa4e307
z5c95d115377a4f5aea43aab0bf8cf04a939625e1ea6dbc23129b1110531f78454c33deb0bae26a
zdc3247dd2b0c2881e73c4da73fef7cbbb8915ce6f29f9294596ea1ba9d8d36f2883dd64a1e4b84
z2eac53e2e5ba0bc673ed4a82b9bc42998fc6ed46a4d217926bce57a162c4e642e002af834cc98e
z76c9110922dca241448e97266a835070bbdf2a0a25eee9923524f4d3859088b1fc4904c0e7fc56
z0441daee58cb38de13e7cb4db8483c9ff0b3a094d6995fdcb57548bf6ad4d250d2f43f6d4507cd
z7168246419522909466760781fc8f0bfcbee64601b8065b20b7ec0fc67c86e17580e16ce9e09e9
z7363c5684ccaa5521faf5b3c27094bfbaadeb54de2ce285b1eaa70fbb9d2c70518ff83af8b8123
z4db1f7e19507f6d368cd45e7ad365de00bc0b8ac9776abbf54395853d1f43f2f51d2ce88ceefa6
z3bb315468de302c2d976b1ffdf865fa7ec329ae6c551e8081e51086af6ef5d044156a8ef15ab51
zbeb39ec8ecb10d2a0b5e338ea7e2f35e055d4d7367d6ac35c2b5d7945d48fa664f80026da517fd
z152837e5da131d0bc42c5f4a133f28c8fbd25f00bff256897892c094edbace087875866e0220f9
zdc8af0c38cc25b25cbe089d9373a5d2751d63bdc1491af91126dbe0b94ab9babbcf3cd5d0add34
zaa2fd8e6d017fbe70563fd922310a1e56ea9ff9352ed547d689236ea3550b27954bab5b8cbac1c
z1e113a61bafb3aed3555e28884fdb8a20ec2ca03ecbb9c2c6a20d27c738300bfb56e8fef233d65
z6c5bf3fb12984882f676553713c94d80140a4bce38881ed135a135405cc15062421705c0e7112e
z5092b4298e36da4b786d0dd451a2d564c42d2d6802214cb08ae557c82b0a521e2c84fb5fcda823
zd8bf579831db7cd5662e6925a8349f905ee4ba317a42a2b43245d530de643c25e917d434bd6164
zc84c2941512d91ddf5c6792db8a3eb35f609fceb52e92ce702b9d0e00a6a9b196b6cb7a9024869
z3ea33d08f5ce660fbc33c2a39825495977a4dfb2de8aca99f8deab72845dbca64660ebbd1437c8
zb9b0887157a3bfeacbb1955c1384900e46a51de68a0387f88ecb28141e05e9483ced5081367dac
zee17db90c776dcd57fe8c1a397a177559bde6e090adb6d3c89e6217da008f6051a41d53c8d9871
za86264dee5c53b493a3b1fd97ba8d7c38ddddee174dfbbdf5ed72fb70c97582a60197ed35ac30b
z18661d04acaddfbf355d1aecab0848d5c4ab2a1c49e5c5adefe9a1d07917a26c094899d9798a49
zdeb1ba6f7caf13cc13664544a225500230792d67d64151255a5705fe41f5cc92d6362e48f0e385
zf9d8fb77cd151a060bc87a73b40f3f1f236814e5e6e6623d3a7a8493b11dbd4385804e26f10e48
z9d6c0dec874ed434fae196d68b25892e58508635169eeb55ed9307a3a11b8ca618f59b8bdd9233
z06af98741b1c045853009e70b278dce7acb84e822d362e4356af3949a75fc9c0f1866613d7633a
zc678d30a92a8d502af6573eb90ef88601cb5ad814428377a1216ef6c44c13d22201f26432fd8c5
z5dd8807ec2b9d915263702a033592a6c982b63b9546c9fad29ba7cd41962f321ea68cb2602663d
zef862ab10b610106d69c73de573c13544e42aa50b403c2905ef25a0d4cdcba38065c15bc682c13
zb8bc23627e81c0482b3f35cc27e54ea70298a92a53db3b5b5ff7a47696b9548ed2780c60c128e2
z575fa9145db2f566cea5a27d21f774bcd66cf0b2065cd7e6a32b51401e38efed4083a708dcc46f
z374a82a416182381030b6caf507318f0b691a69171ec5093e1718cc6b6a9fe546fe2123d9aaec1
z8fc504a18d80dbe32847ff8beac2a033205d913e6b461d267f5e28b7bdc2cb3f155c62edce0dd3
z1c2955fcee62cc1a5fed209163e54f04035e5fd1b03f57be398ad6d1858f5f14821b0660676691
zf819577d143034c7e08820e48db6c7d3437132f919f4c5b1bea8ee8d05169eb83214217cffbd68
zcd81833cc781e21eba83f09d12a352941ef046f6bc21803739f82e34418c4e3a7c8b65cd930692
z2c42585046f19ac6ee89bf3d76e52e0ba8e3c30375d1845125cd9582665a206368a3027bf91904
za952f849d897b972fde7240aa19152fbeee6e3b75bcdfe15671e86f261cb839ad661bc7c061cce
z69043cd99b5c17e14e2145465d0495f4aee01abec75a2e2d57d83b42ae4285b123b1e1eaf9a696
zd10e21bf0427578462b72f3dde7bc17bfc620e34d4a1d5d6cc48e20b6b8b638d84326f1a474c0c
z43734d139363cc461fdef5bbe4ed4ba5a901922f273ada245b61636c4243022266758c46b65619
zed8d63f72e47f9cb4425283952db3d2737c51370f189b1852285fa042be39fa09c4638cb7f6003
z08c86351e5af5734af6258a443f7aa709737b07cc068dc38f71a29c0d3f5cafbb11f508de10529
z70e1bbcba8c20de0b6c7ddbe2b9dabf6825c63293c6351125f920c80f4fded7a98c31b70abdf66
zc67ca7c44871604fc106675aab890778ea23189e33bb9015a14ce79978657a8d99b2fe57411e34
z15a4e8c86742a7a1d76b6d1ee8ca374914288878a2b333b6701575b3ed49735d0a62edea19dea5
z0d8ed073f4fec396a2005cf19d292657edcb4c3b792d94e8e7dc5e5473269f51f2b9ab559447d8
z33282a7fa10867630923567b2aacee44c6c93c55e407d145c0b8c08b28aee87ab961bbfb60b8d0
z1d11317d6ac2dec532c886ab7fa5b47e3e1f15f8171374132d608f2cc9b40df89c36c46914e34a
zb0167f6fcd34234255e6c413fc63e4e7a68765ae541719547079a1d1a9f95269c09df64270c1cb
zc84f3df18d79bde2b3163ff593e81008a986f225795327d9ccc0cb842f17eba0b7c30608113379
z2831e0f400b5204a401368494470bd5405d06979982cf1b542685fffcd74fd0c19c73b8ddde373
zfeaa8b3c7ebc3ad496668235bf3144a711506c9a1a66e165f6e803d4b26ea4ccbfa28d9a30777f
zdefb8de6ea5177768170380941d6f38ff8ac8f9b934bf1a696ce9d487f41555b1e2cc9e6aeb8bf
z53f3ece2060247919ad854fd2d8791bfbbfbc0135a7d4a4ebc3e2e8036b9143c4fabae98eec7d3
z71a15208feee6412bf1cb95146bc8a223827999305f4ed158e99541a8d0a4afb49d923ffd64534
z9569aff125ae5932f826eca3932c68e8d8df480fd2095be44281472eca20f70043f3e82cbe48bd
z67c40a0ee597f6170920e11d65a757897a84345db3ad009ae001eff79cb24d1f8a67c056bebf45
z4a615b8c83911206945c719ec26a34658e626cc16360bfbde4b553a88c833aea04a5be38f18d51
za4936ecd753ee72bf09ac80e5722e9ddbf36c732810817ad148f8d009124529806034bb3338c03
zee72850069b3284d78b52808939b10de830e2a4f8b263d5daf7dd75f21f050daf3db52179d4baf
zfe2247a02632819c66e6845b4ef31f6a1cc0c32424339dd2505aa5f56732e141f563ddb91fb5e7
za4d409b3ca5972dcfd22ff63233e4fd1c9ea8e224e8825b565f53b4719db8002794b0dcbf4ec75
zc8ddd2148b06fef887a14eb162a5a005dfc69b77080ec8eb75b23c12d9abf9615b648c0f504059
z26ec60fbbcf77d4c90412a7fe3da8bc4e65c552e94862544cbbcd5bcb763c35646b3aac28afab6
z7761a5aba2247bfe286cfc01dd087de5f285d9c8a87ff845a54a45aef007adec06bd75ad786562
za213f09e70b2f6dc57bd25bda7c09c6e5eac5578099bb9d2bc6bd8383fd107395b1cc3ff898593
z7f58a4a0725348878a8ef356506e39f166daba870f49438ee966dba170d0f9d0f3a45e1d85e5cd
zc8537bca966cd9e60690952a057e1c8102e386d8969edb38bb24d418f19aaab16c58add8c07f26
zdf92bbd0873f8617025e1a3669287f80f6db18faaf8b0e454fb7a9692a3e4623b6ba4033a1b93c
z1bdc81228605d8a3fa0f12a1436bbd28fd52e761b797b2047a2b40d73afe439ef27859c35b3b3d
z227c6f08ff741c38f8fdfae6e711a397d3835d883c3334e09a7e9ea26ee276816b4297e87d7158
za9d1ef55aef5fd4e4ce4dd50c0482f916d41e71e1c1d42684cbff4312683120fd74ec17de73e8a
z1192ba1b827ec5ee1c1b49aaccb2dd4f2097792a65e42f580fbc339e1fa253948077a35be61d35
z19765953b1ef1573e18edb418e1ccf880dccde8a0fb1ab3fe3a4843641f15c9d74f21925685f51
zbd48bdb62bfee0a911323c5aa549c9f770f73d36a4f715b30321f1427e77c576a631eb72acb6f9
zad510ec07dcf5c377a3317168c2e250e5b9f741e694e004ef37e3297d20035c63903bc7898e8c1
za92967b7239497f7fc27a9b436cdd315e1c480ce152130f26676983a97e00ce3223266ad3e39a2
z6d68d09e4cb05fc15d69c5a026793a26e384484f064a2c3e3bec097065154c32542fd42add8a74
z7db0c5f6af6bea329e8bd71a142fabaa2191023beda7a88dce81211dba7d3f5099b8d7c95a7e21
z2e44ab19612e3db99c73f386ad6f9fe11ca40558d92f4ac7e753db36a11a70e95f6d446c65e3cc
z13f014c75201715dff603a88099eb93fc3eb88faa55c6f94459fce44a0c7dbe43e0e0a339ce44e
z27e3db5ee55e77da990e6258bc2b55eb5ca52084be6042abf4fb6ea34079f0d8349ba0596b3d96
z670a1a7cd19423a9bb4653d8dc16e4f269912c5877b757359097b3079495ae65a893c58ff96629
z2ece440e6891ca3a8e52950934b98b639897f8d1a2971dfe38ec61b9953bad7c5bbddcb5527be7
zb9a6e31c27c2cd4c819d8e8ef52b6907ac65ceb38b251d9b25d74356f12c121991ab7ed1e94e99
z1ffb55726ed484ba2d56a7a252b2a5c6ba17be2799504a668d1ea1172bf923e71823c4ef1a1e86
zad4e406e24b5467f5e2e420f785cfc6561cd145a0d3597007ac2c554f453e57294bfc4e1a2922a
z93b86e32edf860962496977cf661e71834a471614029f53cfe7b86ea5b00d92ab6062d5d585ab6
zbaa029da381a94a127bdcabb830c0f468fb155744fd14499e952b5bac288f323ebb7b6a4b7eb1a
z2fdbcfc5a0f6de263a6db69e7c79ec1395d28a4c9a77420f68d553b97b817b5d572b074b8af266
z5fae2fcb4766f084ca469b87bf3956f1935f635203f461a14b31f5b108da2cbbd8beed12364220
zc87888289a595820e21b5d08e07b19596c1457835874bba371b1c14ebfaca0b9d8f9c1a7aafcfa
zd8a444bb34a2298364fbfdbeb9344cc825a5443a866136034d38179c95095d959cd7c56c4fcf7e
z0d8aaae76440e1968355aad680b4182786c0a6acb1d636001a082f96836d797baa8cf90ba90782
z4b9dc7e3893ae1fd6a0ec51b024629a549efbc97c6179e232d85a72c771161b2bf963ce04cd606
z6c639de67c6a596344c4bdffa236c9ff94d3b225dc9d3f78f27e46d7fa1be0924c720c80ebc570
z052aa43a2c661457076815f4a4d37bdfb541ab7da8dd5d158280990589030e02af2d3562a5ebbe
zc5289744ebfb284172480e8c2268f9ff4b82992fb744c08cc944dfa3e63824b88bb4f1953a155c
z04992e8474900363d122ab3e4f791da2daa59a6dc69f801e25b787702fdf5988958df6c86f7874
z4fcaeaedd37395caf9719fe95ea3b318bd28ca57b0d8fbf16ff93d2e2fd12a46694a7216e21061
z17be78bfb17c29aa86b2e621f40ecd877d8fb8df70c670ba88f0997b7884441581815f195b89ad
z5d21f6780bf84a0ce1661814d3af79c31d66542433a72299b285fa6ca73e014bd53f0aec004828
z38ac7388110ef00bdf554969419b941206f1cb072cf5a550d3fb4242581a892f4eb24df4a09ad1
zfd5763359ebba44633a26fc7e65cb297dc0f8c37885c07429391fa91113f8d5fa01b3f19fed860
z8164253df2a26f617debafb221a3afc8e72075a21ab12cdbf87c69c0244f25c266510cb09553be
z1aa4eb313f04a585a403c46369c19a3ccb9acc4563d1b5d127776e4b294442940369f68a3e2d72
z961b3b8133ff56902708b2817dda63da93b64c6d223391e3cc8fb0b1f497063315ce79a0ca7370
z8f60161a8fe913bffdaf3697087b85330a4973ec08edfaccb50034af5381c8368fa88fbadf6c12
zb0e720e517a2b5970d8aa54eaacd1fc3c4f0e1172097a2208e0a1615c43c56b9adea228a38310f
z4b2187a815055eb225ea3aa44e0009910ed3eff1b2cbc98954c68b47a57b62b2f720e860ca8bf0
z606358a49399055cb9e43f7e6feab7eff1a4fa16110485254602977d2b26ad2e4f9cb4617eabec
z0023c2142b3ec4159debf77142040bb6438204b0076bf4a35986cdd4bd0c2288263bfdbaf667d5
zcc65c3e1065d6778312f698d8231ac613fd178f4692ac0ea2283ba2f95551fd6210ddeddb6f47f
z58557b908d69c5d4f11464b58c2241c19969e67e688fbfdd61d7d42d3d9ff58c5c41436b841f1a
zefe5ba4de7b53b11332da3c698c0648863549af049de5b5462b903a2d1e0a9aa27cdbcdb93446c
z5157bfcdb0f8f3d0ff3761ec1351af4bb9c1bf1711732136ff5e91c4d7e73cbad05db3016bd28c
za455d3cb7b652d8a45f1e77530c2faa960e2a41f4da3cfe1c57071ada099a9bc313258093e9619
zb4514bbf002c45aac2d9668f84d2c93fbd39f79ba97e707cad01a514a99f40f4f6795bf397a035
z23dc64d48aeb35d61daa3c9cb0311d147d969f54e6c7cbb36360645816f1a7266a8e3f620acec8
z510e48bd87bce77cff2a1ff31170d27621906e886b6c47a5501690e005fb167bb58a09794c1cd2
z0968fd27f5916e4ca554924f8dbf8aced9c7acb63a71d30cdd4dc9880041afda660a76f703193f
z748e81b4ad7f5db65515068b6436471a889b1fd6f0b485ce95bdf3898bc4a36962dce5d4808aa4
z2dc36d8887c4f0b9c6ad0a8cbf80faf913debc5ca08f50f8172a1b1ae295833cee084fa2613cbf
zda7fbd0dc83ae6cc16a6544cdec9d14f7a2191c331b0ffdecefbb2875d0127b3ad6df21c88aff5
z272adbcfd97f6b737f2a0ddd8d5e8174df27120c5be1c79bb7472df83c23499808c5f8209bf84a
z0c350870ed216ab385a214811b18b7b9492d8913b1dfa495a4ed95862e1592a072248f52ab6d11
zcdce5bb1770da515e08030a66f986bf883d8683d673513d8ac40ef16fe6ddfbdbd5adab05b183e
z7eea7e7fabeb285d7a7ff13a9f91230ec2d9208826dbb82941a1c4b2d7d9ac8ec97c61ec4d8958
z339af7f997faf4168c1a350b4b0a6272514e210a0f72be2306d1397496aef6e546a97ce8394be1
z3b613e8f3a259dfe8867b39b7495cb21bb353a96d7132becae22c300083aea838e3932cf10a9b3
z1aaf3d50ddf8a0a16bf0af1c87ff71c091e1d5a348f28f216d6f4bd7326229a5d26183454e2e79
z63fcf7bf557ab0ac52611f51e9c4c87f38e991f3ea4eba2c06204aa5f3342c96d83c4749ba57db
z275b638ab9134d84f8b9295a17230b51955159269caf097e2d5882452d979542faa65155ff2311
zb57f887a90035f075eb4cce77ddcdfae73db559058374e1d66a70c1ceeb4c391b4376c1394b92b
z8d666fe1358516b9378f4e624bfeaabb1c3991891feebe63bb0c3c07b7bc4284f88719c8c4c58d
z9c9c8ffc05528b48c9ebe6f2a7f4ee9739eedae96e5d9f53b69b68a796e150735a9beae7cc649a
za3c20ff557499866f948d2cb38d8ef2f7824e0be1b3d04920fd877c738057f9b311665aabc7cd8
zaf3ea191086fc0726511ce7d61bd39120315488c6fb0ea4ce5f808e0eb93e1005fbb69009c4f29
zf56aedfe58c204c858fd82a21f080fa483fa784c8295795cfe864ad3a11d2eec152b5dfe1f0d77
z15fe71bd79c2fd8d30e8e078dabd50356026e8285d53a22bf6ee3a91f3827365d10ccda0d046fe
zfb8154bbbf3b046d1a56129bca0a018cd9a56a365df94b1782b8ba5414e2116caf70e7536cad28
z47d3fb50807a3aa623de759eb53f0ff83d051951fce57bf756dada110e6e3a7b5af6dde092cc40
zb00ffb062a1c38939efd2c27043281bdb73aa27e6ea68b1061d155f59bc30948b1de6137408783
z06644aeb0a5c899d74fdbce4cc6a2d1967cdab5d679781e44680a4c6b517782826859346b604d5
zbe92a450e1352bd70f4f19f3e811131d20c7b4229fd4ed80e4f92a7bd98b75d36dd36c8874aafa
z58b9c997013364c7cc5d3aac212a2f317c044f014def15b90f261df04b15fb977066d37c86cff0
zb9ace360672df1d7bff2c373fe8d4bb75fa244957ffe3bec23086152830341a198f9b6a7c99a1c
zb1bfc40c58b0616225eb03eafa9a7c683f3850f3697bf5c950699b9f1e0c95ef75c1baeb6cd391
zbf7ad67e428772084c312414cd8697afd4b177c63b5a608fb4ce2372a84639a10f4dad015ea035
zce3e5b6b9118b4649ad88b0a33290b731fc809456176aef6083ab2f668e18b901530b314580d6b
z300d463d3ae256562934a7ed54802a86b0f10c60db6e8a4a878bff54d7a23d61892139c03b546f
z92e6c8aea8fc998929618c8ef7c925feccf8b1c34383e6c97ad305977ec7897c343cb25de405b1
z436c5f6fc43376301de8f62113eb5ae22089011292b4e243483c89d7240faa4ba2560c1562625c
z4cda98a6b1a9caeea1d0c4492c6f5b0545fa58af6c7bf806b56332375cfce4c8d9e93eb4f0f43e
zb4b52978f60b9a19b97235b42ebd839c52be5a591e29e4880555095629ab37b9319ace040f5de8
zc301e0b190a76554491af74fc0b8dae59539b6091b9a1d28d9c0fc238a9990447e6f414976f4f1
zb3d57124c29fbccbd74fab16d2c54910189eb7169c4b9257b1c73ff9cb46517b28a1ccd6974a08
z4cf7a243204351cb382895b8bff45735629cfba18f3f4bee8377cdcd36061c0a6e776c10e48629
z7ff3d759467bb3ef103d934136c85671c855d868703927d114b9d912176420081e3eaa9aad5323
z838bcc0b91b0eb8c195c5e313be9993c8683dc17779c8be43bb721fa62cc72348d30a8e57e11fd
z83a49e0086e6ae7f78161dbc4e7f2c2eef59b7ec1bfc5571a745ec13dc485d10c0abfc8360b27c
zb28ded6ed7a151f223f689c0071bc6e20f6a6807929c837247b792691a103b5dc0a6a8729a7aed
z5d4789a5d5842d00325291165ebef5ad7ef02ec81239fcc5987374a39ee0622e2b28f0c9852307
z4f9afe9fd05da3f7ba4366bc07a11959d29d712da3a6c476312c380459c8600421e04df5b60e3b
zd00db043d45a38e7778a20ec3f408a195cfd59935e8c67748b8330cb706727cc514ae541f10166
zc71f8ad311276edfc2831345f284fd1c6998cab00fc804196cfbc1605ff2753f89c1b01bc80f50
z9ee6a5599af51cc9619662aa8a9048019ab64cf850135fd768694ab6251971037af943e56efbcc
z47aa74dc83b0a87a5f614180a838012149b09d5f2fc41db9bb21eb6d2785b73feb3ca92e0e84e3
z0029c975406e2631515a47a5889745f838a3bf284be2a26b809848cd446de7258d9fce6306d633
z43bad513c0be9cbf317d457c34d06aa42c9c2fbe1e8a08c834c6c2c146619a7cb350424897182e
z4e6d6c578873670b9e2a514f8cf48f6e0ba7d444df3a40b7786f026ce45e38fe578e4583dc11a3
zb4f80328c24ad3b6291170811279bb566d1306dbab52a5376cee601f1d78e3fd4a1cc0a5560d27
z8ee2fab5e675bab7fcf5d75fc2e080df6a6bc650a3f05bda5e1241867fe2e9b6f676d7a2de4ea6
ze205b64707c1b5f7c1e20eb48011aa04d550dd1ed1b8f9ecd485f43139cf9d146c320d711d8af8
zdfb2ad73562743d3e5e4a18515604a365fd29cd9c385241e8b523157749467a3b61f913c15e664
z5d6fd6dbff7107d2fae94c7507497470d68488eddbb6390284de1306c59363fca2272613686be6
zb05eeb527c2332a9497474a72bf1cc647f0b671fa51109ea6a415be4eb498fbb62b7455ac97b4e
z3973796740f76a55a41fbeec0461e10cca74cb2d2c415217ddffe0eddce54e85396668d7995e75
ze9dc20ddd1b39d32129a4a2774da38ecfbb8dfa75df570500bf131216a27e87225426a1eb6dd50
ze487f22719b3ebcb268a70351728cdb995eb8d10b6d90601d332165c89c34d93ac4caa46e89db8
z0973368b956ffe542d21a08f91aa6175f89715c420aa46c08ef7f65fa5893c38e980fedb26b217
z3c32b69d7fd65659484fa2046abe0597d7f09c7cfe5f387625047a0d30f22217148f385d34bc4e
z02c5fde422aabbecd7d0e8fcca00f6029841b50327d89b3d351a33b60bf482cf4d3c82d340a973
z981b8826cf4f19008a547799c4f620f3bcffe50a99169bda3f7036b1f07c6dbdda3e44855cdddf
z798b5e2e2256beb3155dbcffce41cfbea0c788ba75897a85209a9fad30f7f472dbae32b1bc26c7
zefe3d3e333d04214a7546b563f9a011b41c29f43f672990296c77e078a0558b89024749a4daeaa
z6670c5afaa20304d91f8863aee0acce78ceae6496b0178db99197348a278aa4b5c30b5f305d3d4
zdd063c0eda8f68611a637dae16135b2a991bf3f0769c5c8e01cc47706af97002ba09163163010d
zc2f2ac9bc35f96992fdfda783520ff19cc560562184dc167fb320b9975ce50814febad2c808e41
z992fb5a4b026fabd43b88f7cf5a93a220169e0efd9f41fcff72ef208a5c4c944b6bdf8b173b15c
z97b0a1c7178705e89d66e9e7470de362ae82442d94a1992ddc16690a4d3b9f4098068bcad9cd40
z04bf45b882436da5dea482f2e759fa25f77a0cea670c858b47c71a488a008d89aec9792dcda850
z10ea4b880babf2744d4701d2e4470ee5713ade7106eeb282477aa4e40861fa01a1ec75f5d577a6
z952015dccfd6a0af173e3831c60ce5ae0d5023ea319bdb0b1fb140f123a1954520f6d4a6805c46
zb4d2958015ce96de8a5578d16e7ee7d291407cd008182b2fb46134520de77e2a9079de37345c74
z1af62b4c0e79432eedf36d9637b921fe56ecf4ca862bd26f9870471dbec51af8daf3f4e62ba660
z9306df4fde37ddb960a0a01298115481e6efd3bf8dd6d9b0ac15456b8aa9dca78806865dbbd93f
z4bef62388a0fa5dd115a6cea2d065ad9a82149dd3a9b21f6835e67b4b327af52c35e0f62d11d94
z85bda964f08fdcd1abc4ef845f24354f3ce6781ed7d41bc4b15902fefafa5b336c5af34f81ecb5
zd8efe3455d4aef924b41d2c15b413a577907e609947c11b3061a698a86f72a87c5d6e383e8bf3a
zf616fcbd7f88d530344c8d92725f0adf8f448aa6beba139dec2a4c25700baf59403230e0cb1592
z5621890de77f0ada6eee2c1426002c2559600088944a4b8c260a854a4fe2d039ca4b9dc1532d47
z636fda440ff1c623bc7bf9c8a085596340dd4289619c08f60dc3abd10a8b08a49dc3b6b1bff377
z6be7ac8b80495e6259e5a3ddff22607e16f8292cb1e1b9e9cc48453f676ff0a46cd3c4e87f4a43
zb0aedd2bd0f48e26b063d95c43a73f4d8c1b890c1246fbe6084bc94f260634433a76ef345af429
z3dca7ee577cce057d8366d7f54a5c3e0c5d279780a22fe6cc1b2d7fe12dacc4bd809399b217894
z7fb5e86fa0ddf0ce538ed45086212e0cbb99c7d134dab9aeab8a8098609f00c3ffc3ef7f4c4637
z5648ad12e24a618bc951470ee00c5538871631e56d10226e60174f61044f21ca24169928aece59
z12d40231404143d8dd8dcd4b6a2b2b5367f9d60da83f5b3983ff5f41e7148a262d5ea006032e60
z495907482f9036e707e2a8ae7a9435f73563f24a97a5c8bbc83691a2b68370b903349182a84877
z32c41a2959b028ce81e8ff32b1024ea69c11cc71eaba6adc2c81a5bd42fa28aec380c4df636bca
zec339eec136264f62901e497960265144fa6ee091942cf17ead96bfcc5c6af895bee615402cda0
zddee392a6a6a3da94fe4d33e4f4eb16d54dc519a27fb5686aa67503e08723dfef5ce5788679d7b
z1fe00dc4486e067f13adc9391a3b313b975d48ac882bebb822bd7a3746b39eead8e1502a48ac04
zc4752ecff818343bdc3b636dd429bf82b9d97566f5b98be7985950ff1df65032dbed3ce74e0463
zfe63127f73a13162208f957c346b95d01fe69222d3653b29c77def9d72da7275a3a64b53a2124d
z48a63fa2f3516fb0c37288227338d6239347c889679e97215a9450893206440fbe87b021eff7d0
zd461e844bc833a971c1560623556d4ebac971e66997faafb706c40e1979cb0ed9519ed8348eef2
z707246b87940b1055413ecf1cce006fa0519f9724169032363d3b1308b013938292315c2b95542
z0ed0b83d2760fdc8686a7c57561b4f924bdf4c173eda6f27d5393dbea8b0606c5ee6043901da54
z9213cd11062038b7f06ad1d4691b8d36e614d97bb6714a3667383164d9fb6265d50705620778df
z5441c62a9147139c7b87864bf029d6cf2d0aea66eab70cb9c4619fe26df3b36f9e1705d0b73636
z53501d62b4435026f37b46c038ce1c58ebf5c19ea34546f225170c954ef06f4249f31d86ec7cd7
zf80123b825b463c057b5dd2b81b6f02172170f45049f09195361a944c8de96895dfc8864759e04
z966bc44672bd4d32f14b5e4f9631d6e1d91e354487837fe15b4e846d0aafd24f2026fbef447e42
zb9613552df48265685f9d184e96b98f678fcf690554f4802fb8cb635e38a3f9a3a2e8e3f3f0f3f
zefdbff33b84f0316f5fe5a15986dd9b30d10c14fa44f9319c4280877530cd350bef3a3a60cf860
zac3adaea3e1114e0bf11bc8ff3a415ec92aa37969bdb79e368b21d0de1d37437c437c903a7e1a9
z7879f70fa77dd946ecc1bfd6119eb1abe0390df14da706a37936b94cd743ea3b2bf1da8fe051c7
z0be9b0a4e66184dfcd75e80f83328fcfe3db1eae79252da0cb955047301c484b89991be253a5f4
zf29c5288b55181f61fdaa4648c2465532018f6a8fca133ba6e0675e9649151059cf8ee33a988f7
z5fb942f1e3e7eb11369e1d06ba91401116603b5fb703f186b3a5b691c998348395c3a75fd00914
za81717d6e38074d50061bd851e208deebfa64b7105fb1fb66eaa58e56987933697f8cf9b33cc57
zcc73be2f72a833628e98b50e47d6065fdfb7a7b91ac068bcaad9e6c4a314a9647eab91c4d1dd01
z75bc0f8f93e618ce77b9e49f461bab605825b0d0dd555aa3e67fd654f134a255d876c9ca360f93
z040573f203fb2e5ca1e984de06d52cd4bc4970bfdb134f28b0e78728b7d92c298263c9d913232e
z3b7d87b72419c40c96d1b4c4c380f5f6f53f7bc736f9746bbf46d3d3093d80f41a55fc10fa8c01
z23c7b637dd45320273c6760fa50733a12561271bd0262462a1410a4d7b552a609054746b399570
zdfefcd5e542ecd9e85f61840da52c26dec32f2f9d347e85f1768804494b209b85947b5ce5f73c4
z637df107c4c9346445d41987e547676056848932c79a971b0bcbd97606af95ea1eae6fec885132
zf0c973329a11d45af2de444672d12d17040a459165b3f2d90cd9077925e50c3067803e84aa8c37
z039c4119ffaff654a3f9ee47527dc0e96f5e7da5e762af2d8ff92dbdf7fdfb284494fc81a57d86
z04a62cca9a380bb9b0e0fb45e910fac2946b6b5d7b7e7c142f72082fdd4e145ca2e42c91b1f706
z2504e6e0153e2a6304cf80dcb8bd8bcc58152939a9c60be1a2d067b0114ece464b3af1204b0109
z27cbee089c420bb0ec59610664840ad65e255f280ae98c03c4a10b4d8e238d2ddff49b8c3394d1
z61c50ac644d69e7f7b05218054a2539f71e83605cbb5ce681cb7cea7d787aaf87aed66d99ea2d7
z04db468fd9abe183c4d6cba6ddb2328352ef81ce5dba3b676c468dfac9fdef4c7314ea54d79069
zabb94baf9d60027dae2e29f96ea9e328a56479bbce8408013db55b1f53ebe8d72945856cf1943d
zf4c71ac6ac917ee2d4399f22c3652ab7d678b128e0d375443a68e9ef2ea2ee459f8d913a465172
z5cd4cd609f388fba9898d0344dde31682bc9fcb13f9ec7ebf69bdab0983bf51720e0807e57b066
zaa000a55fc7e7af081f39ca66faf9e6a03040eb9ce616459909df69e9f6e0036558b5b50fe4868
ze19a7b94f9067aff6b6a25f9fd3f386266912dea8f917d9951e9bf40ef268ec335cff4c7b6af7d
za1beda56b8292d413be08c71292bd680f513136a9d406c1bef926293ac7b417c443a9395465897
z993fe47437d326f09ddaef99a37ba635f7090eb062a90408eed374741e52c743324c496fc5cbb4
zc27212a6e2a41347c1b6ba3c8671c0ad3c6e496d20854b1050eb05a29e562f44050b1766edf552
z53063fe3554122b8675fb80e2102c148fcc4f5e36bf32ac945f07836034f4a9ec613f3dc621224
zf30b869513add9bf4195f33ea0a574ccf94fe0a2e7ca658e819fd00e2d3528a59b2d3fde62849a
z3ad698456a7c3b48b9f64154f9a90afe9d482b077f13a4b324118eb9287804414e18e8897dd979
z48a132f6f1c9552ff56efc5f85d801941b17c4b458475e8876ed365205d990020307a4ab9b7e47
zd916d869a914a9825ced4ead56267a93f333b1e48644682ddb363f75dde9c10c63d8c255980a9d
z984054f61d66b5f8a5304fa86f6bf7d96aa4e55ccf926e97bb99c4b42d8070523cbba97e90fd7a
z03be754706cf734553087d6c7812ba711df4dac889d7c255edfe74b9226210c9f695cab2b666eb
z716ebe69d8be27764b331614f61460df046aa7e8940fbcf79d0940875935a7f04fd8066075f94f
z430f72873708c5d7e3e7f3e798f330eb2923794f3a343006373c2ae0d622feafe1ac653029b859
ze256e997dce6d73747c6a3d2b9c3e7179215c3d89a5e1924719cee2145f2c10d17828bc670482b
z42bf36166cbcc94371d4fb5b5da78e4a0f57441adec327eceb618703e6da416c4bad48992b971f
z3fd3f213b0ee6de97fa6fbcb62c887577749924528623b4196de616c3017974e96e2942b13cc7a
z96be9bf2142b1e7f4d30558dc4571b3d7d02d4c56d3943a79f23c8f78268a2899270a1ecb298ca
ze76519a41266fced3158ef76026e1ea54c36728554a691b29986633ffe7d574ebeb9594331493e
z94cf4cba39417109e6d97b1fd26d4ab496c3656b12d5b032e8707d886929819d49303fc4409ad9
zf3fe03327ae3c382186c36b3f6c4a589ed89be6f0f1fcaf777d8be25167ce96dd3d64304bea760
zc03cd15bef703b741db33d41b11a438403e1efcafc17efc1ba4b5e5c89fb9930a80f61a0922077
z8092bc190b3611f9c7cf73a3e5b2ee83d7093022a2d1a7fa7634f4ccc21d4e6a0f9c362c0d3a23
ze2dad7bdac18e1d5e0edfcab6a1e9f32fa2c47f6664af997e25f679bb2b6819d27bd480c050800
z2f6bff9c6de6669d8aa8e6d4174f51d24616766f608b42dbd7b333c3f4f324ca3e02fdfeed3b9d
z43c71d1ad0f116ae06427a907141ad571ec03caaf8a338efa7bb57539b06445f28b0bfddeca2fe
z1d0398155c64a8d3e33ca7bf5d3c01b5d171877b4432735f7bd35ed9fed91861f46bd4c4b62ea4
z13cc3ec922c7c1fba97fd248fbfda10cbd38b94230dfdc0326a0e07ddd4ebdcca3bafc63ac2376
z177fa4b5ff60ff2576b0779a76150039773df6cb7d35eb74b9b82e120f895f0914776802e1f897
z303307dfcb76b6aa3a959aef19ca5c6dffa2356f2379909cc72708f2ffb15480a6a94247b117d2
ze33d2dc93545c0bea841878a491ba55780fe6f38a25eb88b50d7d71760279fcfce5db30a12f770
z3557b7116351a08f42624300fa75c978486d451aa9ddb32f6cb5849b6bee3007703f18c3228c27
z15eb12a75868f12fbd291d2f58d0d260159cc2b204180ebbed74d3bf46d4478ea5da94e8caa384
z56aeed4e57c1c2b4b77abcada3b897fdbb49c5e8b73d112a960b2a08bacdb3dc6fc470d1786c06
z9b2d376b8dfd559a487817928a41549141602c3d1cb45c6e5e40fb91364a7c06d4b5e7268306be
zee9bb5c527449354a96773d08f5f7d4b9ddf0ff82b3fd9602f463dd44a04ef8f6d0c3c52b2eb56
ze734b4a3e15212b2fe9501c4aebc6d52751168b0cd7b87e384b8253657560da195aed96257def3
z2d24aff0823315a8d3721428f32f71b1efdfc1d58e441cab42fcd3e5ce0516a4a88c0f53d1ccdf
za72828833347a02df256cbc3bca521e87ec42e978782965ce59793343b2e77bd69a62d6b146471
z35e7aa72340a13f3f6f1ca02a060958666d7b7800c37b563c992e43487a6922b0fc9f29ef1c496
z77ab83e6a182de9ea67b5a8c17c267e67c544ed3241e6f7db86c0b49c8de5c348969e40d230939
zf66ee4d063fae4ffb01577727b15059a99944c2d4b95804fb1447e2c478ae5c74233519dcdb95d
z83fc9043f51d6e64617610079b83ed839fc553f80b60b5d749560c3068fd9fac0a1796749c60e4
z6050f04923e6907fb8b99cc5ef38e72f133766e225c0e212273c24c9b288068a55b937480d8b89
z085d3219f07fd22adbe864bfc3f675a739f6ac9fada7ad84d855bdbf2200f120da22afaab3d1cf
zd8123056adc82178609dc1440f0b670d89adb0dc8373699a26f07946f6d75e63bbdce925a4187c
z4438097f87f8f25be58e3e75d9fbebc92cf9151b565e580fbd0480c30723a79ece3b1a2e56dcfe
z4370fc1e4d72dce03453a9de4f35af106e334679825a56a0d4e9171d093ece3c3dd7faed43a558
z2526f138c47513f40bf6dfb7ab7af2215ac0d064b8f668db90e448b8c704aebf8baecdb926bef9
z4a43244287f856ddecca9892bf5751a22a3745703e7b3a23c5bae44c39aab020e3d574ae47d4b3
z43af7e4db60aac0b3d6f0cf9ee36ce94c15b8873969ea4eeafcb4648acb636e5c0e39d559baaa4
z3b6c49487bcb5f7f30a636e40472d1b4dd0ca7bdaa41b05e2ddf8690725477281a8ec9d732c015
zaf4f21670d85606e8ff83a5e51bf21b33d0fe90f3dd3175e83e0c7904b8edb8ed17907db85d472
ze05c8d34be4215d20e6612483574ccf7ddbc0324d5aaf162cc54b5c08239b1ed1cd1c08cbdd657
z5f36a2ca7940b439f968d7e2e1a4faa7c79f097266a1908be581d8e7ad4b9feb4d2139511c7341
zf8756c3d4ef88b667035772886c94f380ba5c4f43eb9a8d47aa23eb4ba645d6e63bd330a88426b
z981541c37bd834f29b1e00392b7ec60b3747d8f5ba921fb3d9b527a0c9d137fb9c28b9f2647157
zc58d0da20391258ed00d48f7dbbf745685ff45a82410423e660e1101047c7743e1f9e377cb14d6
zf1f16762b6b968b027dd27ae28d2e64fc1dd9c4729c984caf448ae2287e6e9bbe3c7d9f4243da3
z6c02ecf3435c0c57e23a1f7c247349701c686fd0cba0e50e32b5ec88b6c8c7e87592fa6fdf1723
ze8b3398624f6e3ffdd8d7bcf323b5b616c83b33951e622e547f14432447416ef101751625f7ef6
z81220c6973cdf874fd9c5f2d1c5882ff6e5deb61951d5c66ccee6ccb5a52430e83f8b52c468ed7
zef1cf3fd626d73879cf1b6ab1e21075e9ab7e342e02a20e5e90f834ca7f40591cbc8f9791ab7df
ze63f14a1c7b020fab6ded3d586b3ac642b8ccda74cafa8d77869308bda98d1d8f7c0a1a93fedd2
z4d5cbb0e179954ef974e48bc2a7cee4b9505ee7205b2fb4512c23bcd7f1594f0ff32d4c6843b93
z8fbcf50be17deabd45050e711122006773ffdff375878bfe62a34c49670834f45459735aff4f84
za4fa85b6f6d6a179c4d3f80bfb64b0f5d7fd6131f7ed5597828b36c8e2343d410b145c7161766a
zbef19ffaf9b5bba693147a9bf0dd6c482f93d0b98439fea12cf843b64abb73e4fa655e77650682
zd7d5aeba188ad2673fc9f65f195ca84fbcf86174930cc03f71ad8c5105ebc1201bc7a142320726
z765815b20532f7bdac9e3937da9253749128631243f3fdb3df7be5537af0598e7dcfad9b315e85
zead85d3cbe1eb381739c8eb80a53fa7cfb9864313680bd8c95a0e492bfd184bd82ba1ea4e50d43
zc3d1b4019a75b7c1f27a10d94546158e6b1e3673fb0e3906612f472a137cf351f4bf6177cf3a52
z335368543ae68744c8ae23f7fe60eb12ba7850a2ab5b4df82756ad40f6c005ff5640d36bb218c9
z16721ff1a906dffaf9de90d3794ecf351ee6f72b702725ee3a149305c5cb3ec29da509f94f40a7
z2f065ed73bb7f9e8c64a66720ca329a25375a14ecb25d3aad034b715d8f83ad8b9b2ed8c687536
za4a3cc7ba39865bb53ac1703d736b9a87b34ee373ffb9d3159aea4b3c2620cec0ba7c46729dc19
z47a54644ae226e2e65019f67b9b8d3af591df1b3f0129f99a40f05ef8d3457df931884aad602dd
z9cb1e52cf867b941895ee5829ca92028dc0125dac80b9a5035c4898740ef3bf8d1e9ecfd01c2f2
zb3ed9ffdc611d7c11a04c8da891ece6b41e1530e20ae12129fce1548e8ead890b0fb58914348e5
z05994f91ed8ef3bbbca7952861d939d2fde84d99cd51f22285bb995182790839266a3d63c01d8a
zb93117a106fa62abbfcb5176528013cc6a552f44e03de652a5cc3a996c8391785bfb414320f5a0
z07b3a596e965dacd8b26ea0245e8e9a3a7329a1fc764ab112703efe31404ebc2bc61baaa360c12
zf30bfa96ef0991fca6a12457b7be1396b5a2676d15f5c284306f6b1fe0ce694665e18731c8e146
z4615d2b5d8ce9ea299730c635eaf9e67d5787b60a784813113bbc24c85ec0d215e3e7e0ee83ebe
z4cfe9114d14fac58b03b13262a404e62a59f633e9576b0e9bf915063118df7330b7c16723483a7
zfbb3e65f31ee3a3c112fb40b93469518f06b6e1b08c5cc55e73aa59a28aaac6114e5332d6fff91
z637184efc4518f825d3f6281082fece95c4949cd4831b5e947a87347f03656ff9bd1f323888522
z0234183971269cdbcfc25cf2130db811c7b38e226dfab4771162eb7f80a735707cfe38e99fbe15
z7b3daf95f8eacdd30767e4c5964017758bc24b141e5af5e4ad385a2fec8d1363fb18015d09323b
z54625ee5a92fbb11b8f9e620a67a32dd0ef49e1c6c7b906a031521f70884894f915d329c68a069
z37065b61c5655532d817f01bba313c80bd3f33e7660e507b85978e0ee18c82669600d4884ae33b
z8cb1be211700168ccc4ef58e40594a0383b97f756eca274014a83f26e66b9495554ea08c45d2d2
z69ffa05f1933d5ce784277d615f9e25441bcd66297e3cee092f722e98713753eac71f28fb4efb5
z6b3cd0221988dd72d0754ff401373aa1e606aede2d527ce549b07a6d02027c90e46f25505329b5
z653cdd8076bb9a7786df36bb42c0b540d9b2f921814b7599af944479d6e21fdd20665d6ee30ad3
zef8bd34b24748c72b8c51a36dcaea6b84421ff74a99e8f8eace2e0b2d7f569c8920e6940e9e347
zcca4eb0630995fb94aa8b41aa6345be7f60b713e87ac9cae22414a6cfb8f820f92e07cf666e95c
z681af22fa2bfc6da7deca2a8dfc9c15bfde66b7074a344445705b73bda11e58295bd29274b0f42
z6ce68854fbc22c0d4efe23c1a546e1c278d940a608446b5e6fef7085523973a235a5b631169276
z62369df19528de02f0c14717a36b941a0491bb4607ae93108a8d66d9138ad6d2b819f62f9f3698
z1bae0bdd7bd4afe217c9b9d2cdb8b113169819c0b4b13f1336fca9903ee073a740fe632fa9328b
z183f781eaef56d828b3b141b41224790183db8b4df30e419b7fcb90b2de39bb30624b00f816576
z7a0be900fb893dbf3a473e5c2df744188259441891f770cd94ad04a88929d8f3a253ad62310960
z7f457eeb8a9c9950571cfd988dabddfc8fa98380f28ef616b5ccc62360113b206fb99b378cd9a1
z4c3e160e5ec6001ce7136851fd1bd67d8bc120d322b4bd7f1a02b75b66efd11f6e7d93d05994d8
za60f959019181d994950765d0c5cc8349905b04821e5b807b504ba41d1b0fdfdfda2b0cf584b1d
z3e7ebfb5ccbfa924b239931cc6a020589016ea7033ac44c118b8e4ba9ed33fe31bc586d24f6134
zf4acc41ce1a26f099a9e514582c4c660b9aed24e117ab8adf42b29d732c42afec9c5d03fc2703d
z7f077adde89d62915370a3a461d18f44d7228648b0a93e004c5ccdd067199597554fd1fc5f0649
ze7eca32962c464596b46d354509e7281da03dbf799b24d89eddbe9cc121775223c96527b0fdf5c
z59541351e3695fba9c2240245719b1f7546964c0033a86b4088888a67ec69b1e761f567f0af566
z65c2ecf7c70de7f0bd8b53384ad39e25f404cc494081f9ef0ce1aba28328a0dcf23139732e1e1c
zf8762ae9a7f9418158ccce258ccd9dd50d3bde303757563c4e3482bac5b1d99c6e19bc482fcafb
zd14241c3f6149bf413ed7638b0d40974232dce8249e6d91b56284b07ddcb3a14452ae537fd1fdc
z25fa4eded6b81ea90fea307cddc6d728b74a3a9c000b0e303696e3d19167d53b2daf0ff7f7d037
zcd59f15ced4ebb4e90a383bdc8a675d70abd7c94d9b6d3f992d7b4a3b5b6d398172a01561a07dc
z8842f67f6d02b124bfc3666e99360c6c9c433951876147d1ba7ee93e04daf607182a4330836ed6
zefb8b67c54e46c4cb06dfd8eb6ee698b8c0df5a22adb7c72ae8418d10dceb9126fab346b9016b0
z122993d3cd3ae47047b666dc576ecf481d8f4e256f4f86e55b2a3ccca64fe39ceef0389d8d3cce
zb68c6bfeedb7c7f142d175c8836754bd3635ab85e2e6575944655abbe68cc721f495c0a59c39f6
zeb1ebde4d9100090d5a662a784ca7278bcf0d24a890d3925d4b35efc620cb5218316ef14cc0c13
z53d972918cbe269cb8d50f4780b85d9831e0983384cc11a25f947fe9c5b99437a229e32775ee4b
z7f461c00b68d7eb035d2dca76019efac83b95076aea7341040cc2f45bdd781b95cac9a460be0e7
zc8760a2060e3a608fa15fa7bd63541901a9494da0f7f4213a626a78d862764542ad2a78f809369
zd57ecc9ae791079a8e1d3d57fc812d7646316fa3261ccd1585eaa4ed8a31410aa44d41fc585456
z55a2235ced1885638d4f5fde5262a3d5fff6bd29e5c39f1f1487bb5042a9de8d48b9f5b55af9a1
ze167b7a8bbc1d786b1a5d55398dbb5f7edc973b7de9a63691fd9ef954debc347ecef93303fa55b
zcd296c917e211de4855971cd24c08f5937f69899c157c0696bd28134fdf83048e7e76d3d12ca53
zdd8fa7d5126dc55a891fe6f27c0f2ecf865fb0b394a171d6f1b24966160699391959329668eb46
z36ca05e6fe97da26bae49dcf4f81973c284cca96a60d4691f3cfc8e6f0cade2aaf801032eea1f5
z39696a5c89b3a5bbc84e389b5cfbfa3491c3e10fcf1b6f67cc4f620b75ed7e7d490de69efa20ad
z6eb9fa40ae777270a11e6d14221b6b84360b66c87c478caefd6f0dd8bab0fb201115c1397eddd1
zef1c72a76503fef072d8c3ca7ec2ab965afc3fe1b6eb7fd1f930fc47130ad314e2468a5089035b
zf726ee510e992ba4aa9dfe6bf2d34cd8aee91052a2e40ad80727555adb6f92df34b874c03e1038
zaf18dc0577e6db4de92988394645ee4a97d39c7a222c9968263bc00c98a84a1db8d8832a83faee
zba8ea402f5eed3affce4ca1630e81f5bde914bd77d2595da073da1a7daec7412ac2ebb746cd9b6
z9a0a4563a15fbfe356bb4b9d78f80a3acc998a523b68c3ba338efebc5d03d9f51c6b31010895a4
zc9404ab5c7e417a0b452453e779ab2aad34431b747d72db11ac263716bc78f60386218a5547c39
z4a96be1ee082cecc260065dbeb15e2a8a8b5592acccc98dd24a282b89366c772a28dffa477723b
z0d36d297aba9be64f8390ca977a858a1180e52c545f99f739918536c5a411970e40cae4889504a
z41ef32d86ede8ee8ef1096aa471458fa1d273060504b39c6b4447141ffcfc2e6b6221b8833a3b1
z0fb5ec8596138b4ffe750d6c3f4ee2e847b37793b76405bd886be4cfe7d5d0ea5d3f6ab50ba21b
zebfb420b6eff17a19c186222f97f0ca110d36d9037a5e20afa9c4601f26fc1a26a30f92cb9e30e
z36c8e65244f12a0bad6fa6769271b5ef60757b86f13a9df58811e64c98490807e3f379ad5b9f42
z6093c7b6365755eccc2ff3423dd58fd371ed7ee5d1c958ed9c8f12897753fd0a2d1b7727ce2ec6
z29f94ccb186c23a6215b2af54337415929282f3939d399749eec10aba6431b9728cabc619853ed
z3eed8a8eeacd27a38af225dfe660e4819461228aeac5066a9659e563b04d3279cbe276178ac87c
z0b9aad6c0df51f28f2dfbc7b5d1af860b31a3fe2b9173031a3b379053891bc9e0a20ec5c452d50
z9404619156aba6e9805a354ba91c50aedae68b9fb9f4aa4f604e9ef0c88ed77ec2c6d3c57a5c73
zaa9ea95e6f7f104e773850d6555a39abb7fbe9b0246f8656bb8c5a0be8b0c96903530c1f5b5e4a
z9ccafda68055c7f669f6ed79d4e3cdfe2afab3b111daaea849a3fccbba111687d7b5a8bc62ca1a
zdba6a9b5736b2da64562e2bc045e93bc26f63ea521d00bc43fe8812466c502a41f2f43cfbb2aa2
z8cc3cfe829017230c55e18f8500d1032a20d85e1c31b2df82f82c912f63633906e956feb7ccf3c
z1e24811098b89632ad3a4576b34f4a69d63ee56f4f24ac739676ad9f6081b183b809944523a974
z8ee6594bbd202caf3ec36ba6bf48aae26727aa9e683a7fbcda970ef9f695b4c9c5fd2360338823
z1902bfbc4021e177cebdfa27bdc6782dc9d138673d406b497668d16528789d9983869b41a22a80
zc582bc3c75f768cc82547ee45f88424f4f06fb10aa2cc7f488cb172e43185cbaf33cdf838cef1e
zfd203276c4e8b4a9bee9bf1a40592e7bb1d38b8a00b3b77a6d0fafd0b477c2c878c26ce38ecce9
ze392acc1b3dbe391cc7542531715e1d0e91917f39bf5ca381713a9ccf62e2c256846f61d4204d0
za33d08c07c406845a0273c65c838c59aec379861cdc115ffefb96b1890e8e7a7438702c985247b
z50651f2b56cbe4471914edb693fb39c499e2c85e9b7cdd2454704ad2cd56651c0fc7a5f34e1374
zf7f1094adb353df4e7c3d19dc6ff57a4deb7bbe2af373ed4cd3322e4748a19e5a7b92efd6e89e5
z482529cfb8c9c11d932ecd79996d19e7951a956b5e3056370c280678265b99dd77c9748914ac25
z49159dcbc5e8b2d7698c16fc8bf50f8a6834701617edf1e3d7e9fc9a230d6ee43457780cd73c89
zda934d36ab755a7e5acb4774676f5a80e2ec47b064be8fd75350e62cf2b6e1affc8dd39a8c6458
z8d1a670c56c4d56fed87afb69c581a1b3d48949cf3d584bfb999faa452713bf4b1719bb4d6229b
z10e79f78510129fa8a2c1c1c73c9e2bd27d4d9cb56e02b22b78b00c2431b0d3f1189a44928bd9c
z8cc12d3b00bcf9b46ac432832881059855d45b0aff035c4a08b05430b6434fb4d871e760cd101e
zce72d335dfb81c4934afe71640a4ae8de09e11275c4df0bf810954a620327a38528ba5f6ac24c9
z24d608d0610edfa0b8554d4facc8c1051fff1718024d33392e6cd8dd232540af6fa9fd43507844
z23e7d9d2ed444f3e634ddbe9b45a492e11a314c00340cb26ff760211e29a79806c9e90038ab59f
zd8749efc6cce782f2c70a110154163913a7d52c514cd8294befd61258653daec3f9949a3679522
z3a13aa6507b93586ef0bcd3e5c720abdceeac0c362b073e9195a75be0b340b8b9cd697945d3bfb
zb565d8264dc9c243a9bd83b326fb0495fd9ed205a57c950591fa561c2de106a3d1c034ce5a0fad
z3f86c7e0961c07c77e632c5eff27d7f11c103ebc29ba7a8e0c3917ded38d26997f175003b6381b
z0e142ff56b84dad44fcb4677e4c881ad71bb528ad2e3df5105843bab28af4e0056edfa6cda1faf
z2a858242948c9071e0396c31c87486d5e974e9d90cd4a8e01e92fcd44061519cc18acb70f6272a
z9f9cfc43c9b2573645998105842542ce0b6448d78575c89ce00f9fd723fddcd8befe58eb229e39
zb3c2ee476309cb355db3848a24d967f32883caa530513d2bf89230eaf3a7653a7e928e1f3d934d
z678f4a15841326a057a03394332aa022a4cd02a1c1613e7c88a41e9b6f9febd89fcb1a5d75e346
z8e11cdd1bc56328698fdf6a00e63b5a1d9a24a362c29025657acea4e5357bcbcc529ccd5a443ea
zb8a6fd39942120d7aff4397689f0a78771477fa8181c3c397fcdb75ff19771a2d778b3116212e6
z21c2616844fd5eddbe228b10a107214d80c809ef272e4dfcc6ad40b439b1351ce1a94ef8197d6c
zd0efff570df9c0694e716e281d1308546ee7a9d8463c797da52b020ce21f2d07d9d8bf1e4b879a
ze866f35ea14515dbbb56d6abcd5d78789323f8646f2a9758df423fc7e232dc4d67892a3670c8cd
z7e2fc550d8e24d631d47d737744bd626b9bfa7a2e7df24ad8ae91e8261dc343287eb934ce37900
z7ea993b2511b82f0a2d282641c7baf322eb8893315fc0c4de19e8dc2a7b02386671935a6f64b5f
zb79522310ca6630242c8cc3a5dc712a6da36bd7a4162b5da430b1cb0aeaf6021c8b3207076d959
z5e423a59437c15ffb3d1f850119de1d0a7e400cf2e67f06594fe0df64be27f8d9ae0e5a85b0e06
z5ad9244688246f31569004b0f2a4863aba2b389d53a18dd8267fc06629b6e20fba2073f0669743
z5f0f73615c8cbdd14be356a78fa960c636e9aa1d6ac4ffb9453a21803c6c42c35c8c059d6ad102
z827081d33c007b96f4907ae464c6c27b871b489a4801ba91563e37fdfb779d4789b9ecd8a3cfd1
z0b81a43b2557d2a89bb9a74028c3252e2455caa8ae17e679bf5640262b91f7336a016a83c463b9
z032ff788cd20f49cb6633c05f9f86da44e2def3f665845c3691099daeed9099c06d1201fc4b379
zec76542b461c1e1cb51f629db96e6abaa21f3bfdd67eef53404a2753791809895c6ce78f95422c
zc63ddf73049cc42732649150f2adcc7b75103015ec4cfb07b0f9179679814e82f824715e828897
z93a24277810c2624acf7fc009b0c23186414790949b2e2954582f34576f20218e3530db9a75952
zd75ff61e0bd3b054b0b9aa778ca80763341eeced4fded576b91dd3df91eeabcb5aa8182629d9e0
z6205422179b4a8798e55571a1fe69b6bc043d4ccef18fefc5eab28af3fac0fd636e9ba393a5675
z3cf8cad0f05a7fbc644b4a104b7a0f731060ba286f27152c5b96e0fb6d6f512d1063c98f94f756
zd50ce53449d13e0061204e120a600e9b9c6b76eb135ca4276b13291f6c79125b96aeb90587061b
zf4697f7a523a0ab3f75fb228b15e3e5f91249a05ed3df7615b404bffe7652b4bbd740c281b67d9
z92d3007ea3eb3c3d340df860a9796450bd32000725affa468bd295be60b9e8adb2f57b56c544bb
zdc1eb004f3281e85f7a9ed75913d2a8ecc2105f7b834141473b0060e827354f51b41e504fdb2fd
z4d5d0781488d50aefb0884df70d6a2a374c57a291700019dc4db6b18f5069b722a554dc3b6cf5d
z53433e6a998846c9a8288b31cf8f24b4382d1b3a7af6861bc25e0e49ede078c0ac2d99e278f156
zdf9fad1cec90eee7f99eb2cbbfc60471178731da54116d6ee7496c6ca861e5224cbea57bcdd000
z4d14bc1fa99d846244edb7ac020016b1646acb795da46a092c312bcfcc1e6588b0d9374a80cc6c
zdc80aa140060fb344e42dabac89a82140485721535fea6ef38bacbe408f9ca408bee0eed61e363
zd2434d23b42ddb439cd346fad881b22730fadffe853f956e2f497ff92566c9cba33df2884e2966
z09bb5739c90f932fed2f5402c16c132d7eda520ed6bce4341fb4e0069d9635d0940711ec0b3e63
z325d2548f1d74ec3baada42ab0e52065a34e710313d6df8305cecf599204d37ac2cede6b26916b
zd3a2a58934493bf513413a2f95121c2a9dfe680f8c30da7977d7c7241bd5fc8ee7f7bc8c83c36d
z384b819c84eb82eb658816dc9433acd7ca9e146006cdf07f91689407e47f042dd375e6dddedab7
z1bdc1abb6b595a55663fbaf46c55a1f16b16f93e74c37c8d860a3a579f18f9fab16f63fcc50c20
z513d0bd2fc2319ed0214a794cf20205bbe3e333efe4833e04c88bf2e0075fa531a148fed48da89
z5e6301b3c111bfdc9ba026659d03fb0af892fa38135c5e7536dd01958052dcadd7de41f519716a
z66a7461004d61745c8618e705be27a73bb57def5d3400132efbb93985e94d00073e8cdea74e0c2
zda947cc0afe089485dc80915048e774d8ceccf54a61d438889d07081f2fb2f505d7cfb5580c5e7
z6c8615a60f781e3767586d597c708c7713cddb7958eb1de2d29f128f5876d224982f923192bb93
z26ec5304a7a96ef4b7b4687eaea048e151e7b948ccb9ea87203deed65e0baeccfcdeb569c1eddb
z178fbaeeec5f5de0018d2e9efa6352f622cac8503e886c085868aab4544ae69d843a22df526b90
z8e8b8adb657d2728bb7e98db498b71914545486fac64fa0a9536d4e22fdfccec36b468a9795c2b
zbcf82f1838ab702d37c2db1ef809f4c3e0b5baac82bdeeb7c41e1be8d0940ea035975b422a11a6
zd761b5ef67135dad96ee70fb89acc824020591eb36455f3aaa396500324a89dd7abf44cff56835
z77eccd9668ee5e649e79fcbe494fb3f2f5ddab71a57db3516dbf641b28a9ba483fc699624ead13
z566fadbdad41aa274d55d0c4ea95b46ef936e41766e30849620871d2bbc2014642038ae6885164
z3ae4adf63cb072f18324a89205ad3b0fb8ceb96099d0ee51116fe9aa34c1330f8004cdb9b14ebb
z15c83aab6e4df0c0f150d883356c41c1bb0f15ac3c035704e5b10df8ba7e6cd6558cbf3c96a523
zf50671b1585752fb30caad6c69ca5cf9e019be167a9cd2f8557e2d2cb9397a6e4148c337ee5f39
zd3703a570bb477fd094abdac6dff15d8f71db59908bc875008f29bf2ce2ab2b3cfce772fe2b61a
zf2ecd96747254f512c4c9b26cd921f027d4c54fd41b985c24ad47d16586ce47baddd983b031ec5
z1e143f9b073a704c75f053c7fcbf9ec3ae619db47fd5619d0f8a5b13b8728a8768147f989037bb
zba92183eeacdb2426c1a162a5ee09ce83dca51135c9f36de438496f8d52b25e9b054a9d7fc9dd2
ze08c8e09a5050588ed5f59fbd3f523ed6b5b7309419cc25cfc5f7184eb5e51838815f70b8b59df
zb57ab0373e7dcd4131fa6fd00531af12066f8d31ed39ead72ecd1ba4b681e7d233dad5e9103761
z3786a8c603a2bbb6cc74a7e497a5587fc9a2599f75c9732b87ef07488a61c05d316967e8c33b5f
zeb251d7dd7f02ff72fe11ac2e1720c74b1195f778394040f9df193beb57c763273a8ca15e7fb79
zca4bc4835d5f2cf29510885764c857554091ab0dff47bbc0c2bea75753c537b9d9f8df39436753
z36da5e8899797499b5be4f351cf47e16f1055b0423b1872cb3defe4ae2993f95c023b61b087069
z031e88f47b40744afe6ccc520c820f5a5e78291ee90b114fbc8e70184b9dbabcd39b9b0a398fdd
zc1c92133c5cc79f2c64a94c96c992b5fa75cafc8963a3ccd364b1524cf2eaa2795abc70c4c82eb
z45dba58966e709240fdd9705cc7e8f2e0e373a46b4812b6d48473b4fa83b2b34a84ffccb789969
za625386f66c4167290a2aee8c3c2ad5a7fffdc50f975d87f08ad9e3bcabc89d9137ca314547cf7
z6efad048b689666b3499fbdaa45beaeead488e76d8c794d2aeeb0513cdd4e02a9e41251592ca3d
zbb980b041293b5f09a75da2cee2556aa3bd4600c28b1ca40c5e616e39987714ac817298eebe50a
ze65e4992ff5303939af9141d5ddc13ffe4d451425aac00a30fe1483545789bfea544ce5da9ebff
z644ba49f40a500d701d9b826fdd6ae29ee2963cb6fd637db6abf3a44066908239b2b9cf9b09172
z3c9b5f8481972fb785e916e5ddd677f161e8a0f5762f696210b2a4aad47990232ae4d56f067834
zd0b01a90257875b478b0c9271f911b054f260c986ec2fd3f153fe4fe8b14215b7ba11f6bbc930d
zc2294bd79d509a192c6354c1d8889ec3c394c68c396c0b4d8ab742e5eb731c7fe7d9a28c320109
z832a532573d53e8d2c3913ff5d626f35ed73cd0c716c3bc0ba2102b73a22a1b91bb5b779a63d83
zdd2e1c8522b39c393870a747aeed0ebb3219a7547120276e9b2153712623ab366b9ddecd5d41b0
zd1acd4d19e15ef6b9d1e69a7d5cb57f8d6d7a959ddbbd7409f058ef1e87f0a3859cb7fb1352ef3
z177fc91d1fd5efa22051af1c14d0b712655f64dbdc41031448b1e82caae2a1debc8fb09ab2c464
z2ceea09dec7072a87f69b76d47d492f787e93dc2430077aab03650df08fc6d6e0ab0ffbbedeb23
z69e487e31f6152799f1a8663841b4526b683a84ba10eac9909f289d133c59b446745ee306d037b
zdc5f1de8a24d8837a50cc781419a6cc6a755956bf824c5f99228653029f3d66175bb9482f91f35
z46aa7b11618c713adb58d48bfce6585bc031e440d5363ac69150f6fb3061c2b909fb6529e6873e
zfde55ad3fc97bfb65d64baff34d0733d1b8f89593d4053ac4b11fc20a3713c2e899ba9f45593ae
zb7bfb999bb8620a0fb8a42928b4ff21bdc72289d41dde662b39c4760f16fa11ed6c958614c9f8b
z62bf820c79b95b4fe3eb7dc8821480851951778d4e9549ad3d69ee11fcfcef3dce8e6854a30dfd
zd5bad7acd5d46cc4d418e17b655f6c8b664719dc29a87b543b66ab43975fe6cabcca0e2bacb99e
z1c76bc649cd1ead912ca5bcead055e36895c5f87d8e8e60c25fe478ee900eb68e71f8274ac1109
zbdaeeb5b40726cc84c75730afa4b4f6f01625fb0f55eb31090ce07e9913f4459ae160b49307da1
za91836bb2a962e6d35b9e18c4e9d312fca3bfffa761ad68b5a920888414a5a8df56f68ffacd7b8
z15b054ed9ceb8cabdf80cf7edb6ff2bd307034ce091da0f3aa61d655a435fa39ee3b0313306b59
z11c8115c69a2541f343c4e312eb4b5d809b789ce84ef0b7b0af2f8b85522499bf699802f351b89
ze3f79306f400113f95a4082254478bc64229327cff55366cced1f98f446cf7ce0e005a7518c025
z3fbca948508fb7d33d438fe3efa1eeb93e444b38c912d4e10a5f772feb7180db47bd65c1a96191
z798273c32f3e5df38e5320ce6b478dfd13d1fab0b893d5cf02074eb0912e2e4aec14f17cadc0b2
zaa32f82fd83bba9df673f9af1ccdd16b453fa9a36133fd70f605916145e4bdf777cf7b5199d143
z2b4e403809ba5793599ff9c354a9b2d70e3dd0cf65e6d60a6f555953a5aacb75508273a5094409
zd6eebdf5eeaa87a6f6016437777b102844e9b7c7cdc966bdf0049988941f0bdf91f392a3bf35d1
z6e5a0a3dd974c5965b1d4f65414770d56aaa796d520e39b3f22cc8f44e18efa37cac2a4492b1f2
z20b458a9c24329a2268f92e383b02740b2c08f11cd7a761ebed614e10e991b2881d49dc8a3cc8e
z5d5f7a893f798c80d78f57b70030c2d62721893bbf5e7992db7cdbd495c7c18f24eb3355881638
z3b3502b6a48d9f181f2793df45ac732fd9449e0cccc886cedf4d10d4afb94d90988cc48a904e0c
za4772a9b89b7d532dbb5ba1421b9041b1e5f68890f968d9725cdcbc4140e10d2f4587640b5223a
zb5b72fc059916f269176a85e3682e0c17fc47e0315fb1ae7af0f19671d6817b806f72c64a819ae
z6cd8bdabf1259f0311b325e14227bdcdf5ed6eeea0269724e1c578ffbd7757bb0aef28ec44bcd3
zcc77cca180063740d35741b4520c412a636451ff1856ad373f693fa812a7c8441295253e920dfa
zabb4f0bff90372b91699c6d59b7697eecdb40d8194ac601ea9b80a3147a1c3f1ac065d8fce69b7
zb4191f2b308cebb8932a599ba79320fb01d3116ac0361fcbadf3c6da3d94f8e73622f30efc8b6d
z9cfa9ee526c864a0d17fec8da6c29195490d83059644debe3b21dd21e34fe09295e23ba6965720
z9f38a00c3775ef3ab8dbafe1f4b6d1d3ce0b831db94c7237c85ebb46654aa12a1dc58f24cefabb
zaa3273226dd9389f529fefd7afcfc94a4f2c2041d38ec82e6698837ceebdda3aaf787ba27d78e7
z62d4e763ab7dc2976a9670615968a112f6f11f9727e6bdf1e3f86c007fa72a6a6d7b947723ddb9
z5cd44c08c16777290df258a0327593512227c7233ad01b35ef8b4137dda83ffb52eb89740ddaba
zeaa29b333c709bfafdde71aec9099a7782551a54a37407d1ac749b3a98b0ab067dd04198380c34
z5b73e5b89044864d180b6949636821286ac2808d63561abbeb0750b85fc15f7d6829c5a041740c
zd0899c6b576c0dba617bb5a40677f135a31fdf3c20dcb94ae06ea0133007749a0fea3e09ce6020
z6720bdbcfe062dd7e9674b683d1c20aa38d1bb4065e93950cde6bcc531d410cdfa5d46dd644aa1
zc48ff4f00a286ae7a6a6828b13d2756841d68b3196f7b497e1363b244ca5db03fb72e3c635aef9
z88b78386bab58b7d0b96bbf141c16649a071d2dc36228588ba28a08c347b14239827fb8a155d05
z786d119072c90b45811d08efa28a89e7b6c95e07a86a78e32cf5e4bf11913ce3e04f9f49ccf4c8
zd11ed6f30adcc6da58f4eac075008055597ebd99758ce984f6990bff26bfdc442518495cdafc96
z0713828667e86b5d814991a94177d8ef306ac3de7c6c08e688cf50406a54ef53a0b101962e4090
z459a91bd8676dd60bb617fd639f7e45eb17a6e529071b3a5e2d74e1b330f25469d5abe271f3910
z6722bc53289f85f4414b129a90f4d12f4a4b4ab84334a4e0584835ef9326eb29e4718f8d78f590
z399d876980d571c7b00fb107dd9c9de2981bbc30a6f51bbc19d4d5697c272f43eb4530031df81c
z774a4219c6acdf5d882eb356587c7cec68b6a00a9cc014913b651007fcf37b00d7cbd65f746b46
zc1018a4064a75dc903d9e5006bf551fb31c50999d8039acea11737dd603d8d27591c61115fa8f9
z7620fb00add38c33051b00288fa92550f2f4093b277a9e87bb65f003956fbb682eb45db2a4600c
z36c72f61a2e1bba46fc188ca77d62b23a039967f131a48952ee14ed30d77eca4632d9f4f0798ff
zb2a7fe70ff76df82fd6d3a5e25b9bd7275357f4d7e9aedaefe02598af0db6a87bd5d873a5a78a7
z084a3ab360319a6ae9b4ffd23f1376a2180f8233319daedc655c4e918608bbd5d63f33fbbc5052
z25b9f9ad6c412afd11fc419cf62cfbb2bd91fb0249f941436cc2d22270edfba8709f650742b1b4
z4667313f4d7e9a58a6492fdd53adeec20961d447a89f39b8d3ca6b29ff50dae369a023011a8f10
zf3fe82299d9fca2fe38d37ac35f49bad95d88606478a58f2316b88969fa72dcd0e628bfa9bf9d4
z8f7597569a6aaf228624c2b61cd063ebcddda28176d7a3779a305bf823eab56c2d5db2f0e14d44
z42f26e5890e5c512f3e77b1ff5288b2a397c851a2941f83b2d0342c66327f44c796526dc63e15d
z12ee12ca9d403cb7bf741a350d9bc71c2009725737322e5a54dbd8862e588e879c6768479218d5
zc697da64904138e096dfebf027b6e0af30a4fd516498d81ede8eb4f69967c348ace22009b77e03
z00561d7972c47562dcc69c750e76d92e92c98ed17f8997c48656c6d4ef5adc707e22b7b2c315fe
z86790329d9a24072cfb260bfdf94c41ba7e4ba0b002745004c77c2fc68c7cf5be3b7f63ed5811d
za39c67d4b239588a0105b740a8392f71a2ea1cd5758d1c6d93574e90d2d5aa1b6e66db2e0d82b4
z0f87259c4a3e0121f755aabe0ec71573a86d595ca710e198543dfb4a4fb4cbecaa0bf6b326fdf7
zec10211972dea1e9cd510104d6c94f5e7abbf1978eb20c15e71448a568e8804d6985bfa43f92d0
z06859ef2d10ea29f11901ccb80592fdb3e8554d644749868bccd54e8251cbf55c892285c0f8a0c
z38d563bdfef987511984d2e7eefd137cd161c28a88e7f6576aa7abc4a6ef29f203962d7ddda66e
zc9b2c4e73e125fa6f20575e38ab7719f244d404f6e91305dba5bf3ff22eeaece0bb2cc38cdd0c5
zdd4108fc5e1a1e779b3da4bda7e4d9a41362f1865aa3e25360169011b3c691e898a4357bb77946
z6bda3695f113d6ac736a1f82bcbb4bdf797b3b463e3d9c46421462a786412da5b40de2323a96cb
zda8270a040ed09b0c9f82c6a03a35875faf76671cd9a08eae6e9b65875420bf47179e453ed4dbe
z1932984e5c7e97cf0ae0af1eb80ff4db04a916cf7c3e4cc64a9dcdb53012597ee3f12de0e74e4c
z7552a541c73893b751401ea70d1834dd1863e6600a5a2b81715f5356498ef478015bb57710f0c5
z5b195271e7a33f4b54eaa4f51e7a86a177f2676f937c6a4464c88f239de454fab19021e0ba829f
z393714628279d065ba9f653ffa3a23c0548987434d71c1f7b89c8eea526382aa233457a178a44a
ze431822ce72ae286f2e284b7f27f58fe42c27a85652922de7d45395ccd7096d587c90b48748a0f
zcfc2553e99b3655e4e82b20ac916a87a0d94074b6d51de60e0fd443b46386740bac85929762415
z83b9c949ccfd9ba629fd63bec2baf53dbd3ae32889bcddaf9de81f2643176a8376d5ed86bbfd74
z8a5e1556396c77167b8f38254802b3b2c8766fba5ab69161ed31713c9bedae4df1b260ac891555
ze61403f3dbdc5ecebcf39f32a6f9414d3ee931a10d450439078626fc04260702f5e92f4b71d4a0
z9350aed5f146851cb3e53ff0b87dd3bbaec7501a209936ddd21a7891b9944da05897d691f8c558
z2e2f3c961b0347ddcfb0eb708f01e0306cc4fc8b74e9508354145730a94952a491fb64292c97c4
zb1ab0dbf8d8ada9f7c5e0cd7b7406929926deb65b583e37d728e13fb239157c39631aa4c18be2b
zbf531dd15f55adfea112e1632eca798f02598e9d570b2ec209fd64ec8c432a3f50e58b4929ffaa
z4faf0a8b8c03a71001f391b3fb7962fa3fdc50930303c1ebb2da5272f13a58b522e995e8ed4721
z1193d5d30fe86b8286cf1f122f57a85be922568fb7afba5bf0436bf3b9f609bd009b84e3614225
zb0cea750e4b8f02bccb2f3451c4a5bd96f9ec38c3be3beb992c8459d3e95d187be3c865d9e222f
z4ee5c837994d907fb741774543bb948046de2c657a2688d9645d40a23317ae859e8dcd64a18582
zfc93778c25ee5a701e24dc2dc6281f84ff1a0ffe7b01eded38e14446f24d33c99dcecea223c99d
z363ce47de514ba5fef3bc3a62904c4fd2639d02f7ec64f403347f73569714d624750c284df4d15
z1a965170b1bddab141c25c49ef082cc4ac2d7a3171e7b3cab2ec842fb88508dcd89fa5f1e8a4f7
z36bbcd8ced8bbd3d3f177b7e995448dbd96245c953bc6da4a090572491be95d6291ac69fd73256
zfe3a9f6d697904d0858fe01d5fafd2c802016012a729e5bdcbbfa9a74b891cad0a5ecfbd219261
zf165032a5a9d75f58d0b07a121dd7584721a370907b7edb15f679091218331317ae2f6846a4b59
z405a9febc1137ff0eef063ef083330b6ce478805a69f31582dedd5397f31659049bb229690b48d
zea1fda1205898b1992975b1557624aabb820ea426b4d2b9ae572b4cc9dfca526d869f8856c664a
z10e24c938bd9469c5d86e8c7be71319b27547fc9ffd0516173db35b1f9f0b4d12891ac95b0fa78
z37b79480104cdf46d6957b55209b3a89436c287e2202640a26e7f3b27bd80505dbdde7a0d66c4f
za171ff750ec864df720337957a6051423da9d14fb66f44efa8040b07d5666a99079bc13fb59253
z444e1c8205fef00c23b9286ad9d5a6db09d5c1cb2adda19d8c4e4fcd8cb0743a2d3eb729afeda2
z7fb590592cff5d63c66137343146092384d937f5cf619841f39a03d4d886ed890c302ea792b88e
z43014b533723e8acee1dea70b9e768cd323411b3ad9bba7f8ab66eaa9e627dc3cc5dc800539b25
z7b29808a28bf903498e3cd59ebc78fe05cec414e9f0610b252204e1c24d94a841a7e338c47a70f
zcdf83c60489e2a586790740d384b723dc9204bc4c1305a73eac4be484ef878229df67536672b7d
z6385f9851eea30d2553159347cf3cf96d845a7f6ae7942b901d403bdc6e4e8d48a6c6163c8f269
zf2a0d036896a7472c027ce84d83e2b055f2aaebd80996e3e229444142ad5e0e548292eb5b21166
z5d3f9361b81f85367e4ade9f39dfdd1adbfcbdb1b04f841e9b2bfbb151571f7c78136dfd6ed512
z04fe9bd21ee2a3857ae943cf68ffc114805263917db1c3bd4dbfd18fdc7c471e7a9c5885108868
z9d0493d1c8e82e51f83012e9a133b4285cd7674e0b60f1e7e91af9222486059030f3bb18588e49
zcaffd0897048a3e73e7c3b0a3f807719f96c4d77e67eab77e80c270daedfe1d49cd071b05902d9
z27809d27b946564b7a4a65d61c35979138ad6d453d82d92c72768e621283f923f0b68454a65ad8
z2b4d281bcd7a0b027e3172ab2670888cb29b6fa9699fa1ea6683a75bdd157d5b36b1a30582f61c
ze2d5dcaff17ddc204d400654efa3bcb644eea7312c88bc19479759816cacd3e4548a039f6d33be
z03d6a0b80990a5542bbe5ff4d2bca00d77c8603f1ef8b8758293a13c8ba2fc0cae54731730c67c
zffcd11668f675c1f85a2b4634987902bd00dc88863d02b7b2dc57ed0e986292607d48455022261
z478c56c83be5975beb4bacb0d216917bc6c47672c448dfd7f92530168ca1310624fd1a5be0a9d8
z097b252055da75d648aab249e78f54d0a13c8e1a13bc8d650bc2252f16e2cb76f3af5601489f76
zcfb301049ed40b41757f222f909adf599ad85e36e51dde07a7102f09e4c5a1393184e741ec3256
zcfd024af90a5f3107b37e2f6cd80cbd89eaca793e32878ef44fe8aaad17c71e0abf71820d9c87e
z81d12ac493b04d81d901858f34fb0359b091cdb9b6e076df2ccf4620d43991f2542f4d0ee0089a
zfccccad2528ba0b5db5dba6ca84dee0e385044c6a13884e5a25501a77d5f9c9b478f345d79749e
z4fbe5e601324fc5991070064f8cf49754ff9e7f5d3c0567e89f5bba3c97cde52c615d575c80fee
z29da40dc1d3b6bde641b57530fd7f0bc08da5adb994bd59dd8378fe3d25f417a8eba3bf694ddc6
zcf21777bdeb21791d2f2a5ae807cfd86630febb1c4882a3d7b22f60fa35cee2d4cdd5acd9f1831
z9a78c71ebf8c4d4a25b42ffdecaa51135ecc274b0a2857dcf8aa087f1732b47a0f9d2e9bbb77da
za3b16dff89ea9f59043b95e58f057d8772f7d01befa90bd4463bed4573a9a26381fac3d8e0ca84
ze028860cca3ebe2448efddd69ef07eb489e4cc9cf4a1e29132114654ed63482417f5ae4592ca65
z11a704bbbabe006e9cdfe54cc01c7db66ab38658aa35393ef640275cf88c6c761084450eda4831
z6937396703a181f7fbf5053b6a0b26192ef5e034071500a1bc050b4129a41ac90c16c1736908fc
za0ee8505df8329ac5b2ac512aa66a9ed098b1c07b385ed5cbc1fbc1a4a812e207236e8d715a962
z5bcb3683e49bec2b52ce2a6d4b830e707fa96d4cf1c73fb134d2351bf389e2ad658d9c4b86c7a5
z476122d166cb128673ade0fa8ba7cbf6cc767a61d7dc96b3d667241384f4210f65dfd5b7f6f335
z8120db1ee0b96df14855a82f9b473ecfc9bfd40e8001652832bfd258e1293e6da3aa22d59660b5
zbcb34a36bf47fd294e1c8b3e9296947d5080bb7e5c2abc61cf5299d44d4f761322eda4a5500a8d
z81e1a3abc4c48b71d3d4d0db6dfdaa7e577bc43108d13623091a1118a58df8f0189a730433a21b
zfe53c3303c16352bffd78c1c6c0ab188ae5f009485ce9d25e7827fe8f51aa12d120afd3a2196a0
ze985838e246ac8150b381a2c4e4345ea6299de14826708a803840f1326d7da81c9dfee7f9c9ab1
z74d85cced668770ce9318af582c3ab9034f7c048e7280fc204298ea3303fa9fe502db705218174
z4c2aef0bca76eb770ed2d572c308053545da6258baceef7ac5569188a768e4108dac509ed0d708
z71fc1cdbc890d09207eb94e9a069ee8c7b60b7d5e790072ec7b21ad5697ff7765b3efd611eafd3
z4a99a695d2304e8821bd7b9c51ac9e7e28b3c9f0e2864a7ec91f8cb500b4995a83b3cae5bcdb7d
zc08b8fb3f1ad3cba0e6cd1c596ca6b7f607471ec268cf6b054cb39317dbde9fa16c898b2d11ed7
zfa74113537df2435bc54577fec92269844688b1d0bbfe88549e81a16fcf443843cc8f9ba9b9c59
z4ce088c02a6a1411210cb887ad7b386c56c5c28de403107cd74183b1eb0a61c144a58efc23f69e
z0a96ad453e0ab811cf85d27272931e606083c0cedea1f08aa20b71c5fd6ec0662bc3314aba9519
zfa9cffefa7989b40fa12036f529d772b4c0c9fe0cdb9c73e3c11f617c5294b143d5eaf934b3ab4
z49db79a0ebb698fe930f6a66bba2e3c35b8d3ced90c653d9916f35f2c9a848b7faa608d7356cc3
zb7822cfec1600aa0c2fff1ef832283b7919d59ad9b195b2ea850941c232c8efd25a47e742aab64
za6be98e77d997a23a24b1765469e7056f3cd75d662cdbdda34ba6f1255941e05937bfad15f67cc
z4e54ac274d57fbe7ba057effaa52c16af62382118eb9e2d57173c281fe8db0a3f4328a00064187
z53590d2f329e32ed8a116fa2abd53c70b8d01eb6e0bbfc759e3bf274aad3f1d03874c9dc65f91a
z7ab91489e821f5e3bf7968b4bc4353ffbf1c55d335d636abe7ce9e2c72db72fda5d1d2b01f8dde
zcb6d0fc029dead58a62bf66d0e1162a64652a19ad3e10846e3234b1407dc1e521fcd3651995507
z021233eb59b515ea865127320fa49824b28c09af4e4de3213173f37426912a1b76d7c5ce4f4706
z8a22e05167bddb5636b6c07bf6e142059aed22cb6d8bfbd930c8d77c51c151f1054c9a0a01bf62
z482c82b2b1b9d7cc6e8bc5fc34afbc5fa77c55b053fa1c32299a4ed97cdd4e31aaf711aacde2e6
z016a8edc618fc877c6d2e6e38799620165fb836fab9339826c847955fcb13b5599d9790c3eac34
zf7b62e7216c8a2ad0cdefcee6811e94b0bbb6d4b6e5ad979a100b2ab428fefa0ba748dfea444bf
z8dc4977f76e18d1837be2e82f90a108f938ea9687eb14d9982e1790a5ae4539a5f0f0fdb586cf3
z70d5e4a84c24025f7bd070266de5e2737117ec64b9e5c6d118ed911282d747ec8a4fbb2e3cf38d
z28167fbcbad4fce1033e9bb976a86f21df9025d9ceda811edd1a5f23c847547500c52f244d6adf
z468c2d8a73dc6bae85a6aee420dd938db5ff3d684cdaf62385b0499e0da60c9499d520436206f5
z47487aa146bdad58469a17951bbc19872afc3ef38a138af3688b099b6d5ac0652d475fce68e677
zc5ffab75100f779df189b708c292de9fa90617b63377422b3479a91a78e0b4f3e4b8aab2611a1c
z75075ea4d62a043bdf54ae7ff7686b6d14e0d6e6e076c79294623460e1227ae414d2230b0fd2f1
zaf3cbcbeb64ca72ea05e36bbfcdee2cf974bbfcbd42ea91640cacf480a67619d9d1fc506254790
z2ec8809112434210e6cc0db8d25baf4339f36d8d1a924e49420e3403c2655f0872e649adb2ec77
zdaaf2633308855f4330931453dfe26a6358e858610a0a5f6c96a421bbbe1f497498c826edacec9
z4b5c25fbe2a42864b15bcba96bc7c859586519879ba73eae47b4882c3a00ba4f9156fd91a18c0b
z8a8dbb1d38a9240a55a3bd855d49b5877fd8bdec640c3ce5e5a2823fe93bfb0808c1ff856f7d5d
zcc6fe3228d337654d4a494f37690ae56ddab8e906ef7a3211d9971689fa34abfad48928ec06a2e
z43b50d6213d5ec96356f39806809132368b6b07f3647af2116631e43f8cc70735181a539b9291c
z0672c60d2fa71f1a6990dfeb8252680c7fa0206b41f67193faef5b6e39f90e173f4668b79059c4
z4838f1ed9d2c02a79de0f539bd51601ddf204c6ac02e427a37a04b639df5a651951387061775db
z925af439ea82a72b8b252f5d288ff957611640a081bd9f0b7e5da1214ca0d1ce318c30eb492377
z82b120099cc91d966aea1f00b766759ff961585a95c4c48c36e4020790e2ee5b3c9be2bd882e2d
z645aeda54beb53490b210091fff8bbe14f489e1cb0bff43e2a52bb54974267be232018e62afc45
z2db59cffd4dbcf1ab3e15967971f7216fa2acd0b922aa6eddf3341f3486154e221372981e86a4d
z417920d6392c0f13b881af16f52d9e650b39bf8b87a1c437549fcb59dd7ddc967eedc9e1c215a9
z718138865475ad6cf5f5ab61a7ca8807cb10294d03a04c46dfe2b88efdf4122e5047c9f960fe63
z9ae8c152c3c77a4d25fa6430292abe920ebaf2e050029758ddd6bb04c5055ae561073a5581b4c9
z306fa60f28bb22f1066e4cd2f6beca20454d7cfc32ecfdf8277dee96d8aea6e825bcbc3d6f443a
z6c3897db3098e5ad7dfc78ba41208c9f8c8c86782e19d3cb0da4e96c1771df551eb6cd5b6e4e41
zc4ae987af8a0c79e6ea00aa3f0f78b1f0cc8e5a71a20e7ed3353088de626ea815da3dafcf93bad
z08e790a798d19386135d9a305d874eb5530c569ef6c621b38e48e8adb97ec6a786a5b412d914e0
z4ec470a89e2c58d9553a20e9557ba5c416625e4e219df32ce2c40943548cf1bfcbba3431ca993e
zd18edf60b4a6ee81d9bc9d239341a72078487f6c0c8a8afba4d1838c72ad8fc4ac949bc19735a9
z635b429dc02699adf9889c56ea15c12fc3f8e1b162975010421c2caefbf9739cce2c67a1865995
zf4da8f620083a2747d325aea3a81afb8898cf7485f581910f8fa65350c1bcf1bd597dd01bd0491
zb62d623c8c80b359f59d7c795e0c6dd1ff36b7c39e93e3a95c2be04bd1f6bb5d7beee0e2a00041
za1d662d065ee56f3744ffc5c4c2f60044c38fe9c188cc4f5f31d0f7548b82d267bcef27cdb022e
zd32dd0e98abb42a7f49d5bbc04c3bfb25c1b5764e96b93b1d5db143ecb57822ab36d60f9ef22e4
z784f185b9c3bc326b0dfcb8d01b269d93cd785769102c3543b51eeb860d54a0efbdd082e5e17cd
zaea89155dd2f8d3a849073e42466c95025cf7e613c8c090297c884093db5f91f0574f7c13b5bb8
z3ef8458cc78f1b5707080883bd6c5873014abee16a1d6d6ccbec77de9cb1e144c624054ae9d0e1
z7352c9ed7daa9635c55cb80db1117f10c175aec95d2c5ad5e193c74be80b8c2dccc5e3a520e248
z93775dea6accde6e167180bad041859be9efaa5818f2f546a8ae1e991c6183bbb96cbbd9d4dccc
zd81fa643fe7b9af27838678334781ebad691ee184e77fa4fe1b42b8b554c0901526af432eba550
za727b8033e189814ab6edfeadada2673dab122195bb2a17cd6a56b73d526f8e3efd9c228c8950d
z99e671df735b44afb9aa69d50a05ba54b1f94b1759433904885d953c47a78525e7e84ccb372336
z05187844e4e43929cb30a3917abd39e5dac6cbab61b66c6363f14d1a43e897d0170f4e51227286
zcda62780b9ace7f3eee6896e1ddb0dc323fb0ec96bfb68282c723894bbfb0152d106c845e44219
z7ab7b626d77b6a2f1ffd70e2ecb022a3467db5c482eb04318fe7ab405e60bcaffa43031867f560
zf0c7b2f42116ad04b522c3e6289786d79751fa2e50ece4262f746b48b905ad8bc34c3b04161d70
z0b5750eb361d968bf6eb4d5685568874d70d2daf55c58361780dcfa6372ce47bdaa66d491c1541
z04a42736a2ade374869043e542276db816d5d8a16ae0c7d8c54d869002139f0928ff1aaad61c21
z6e43e0bf5482bbbda65802be57261955e8039ae98120db994d4fb42bce7c72bcbc09208c0eeae4
z218fa93d7ec3c07d714cecce56c9311d8a367d48422b94dfd38e04f91e82661b32a0f1c06ee6ef
z23e5e48d70e22a84698f4277b4a5f4fa2b3a2eb43eb389bdc971e28dded0aa017bb0234a2ba8f0
z2d196f0a06291aac21c5db49ede4e40fdbab6f58cc337e40259282c0d09c43db9e90a9e42425b0
z9b2a7d5ca9d6ee40f4be26b92b81f2b3c78bbd7480d20c4bf447993c859958427bfae6359ecf7c
za994cab3e0abfb7e3dfc9d3b3d90b8e7d44deea5672fc181c685a9ff48b27cc35cc108c796cd46
z450c2df7873edb4da7890767e7581259a39e477fcaec802e345db820fba2395d2e207a4ad7a6b2
zad878da3fd9d9e20ca7a792436798ca67378eaa911440b809d583d5e2b2263bcc3d6fd76479afd
z19614e7d3df87f709d88d960c37334b8c7dd8b9e70d54e2866557d40f9eed556a62af320c249f9
z2911518de069edaccb756d8a31104a824ff4b3a550caa169007e4440e9a1a5737ed288e5068dfe
z294ec001e1bf661b761083c4f48bb6df68ce8e00643ca7d111fea46e1bf9feebe07279abb7184c
z226f08dcb229a9d5c7706f2738b5398b6c6b531b3b046a45da1fe6113258bdd24d92fff7081581
ze52ac8cc9939997a48b0c5a9aa0dff7783767dfec811fcd5940541885e75acbfc486b162b55dfc
z0a68326b0551592c9c87099484fa952dd4029902caa453649f79f52a4d4c1517b304fee1f9d322
z73782396d684465688a063e36ec0a43a6f1c6c5fb9a93be9fbe6016ea656ba66775bc38f9fa04b
z1f926bfb1c41890c2b5af54c640da53b3a2903893ab5cfc19478bab21cc6509974ab0bbbb0cb66
z5927a242a1bbf1567d8fcde544c9fcdeb938ff666d5a8b947e307a55ee402699e5a287301c7c27
zdf23171529073469e7d68177bb178b963f5667adb0efd2089b4fb40158d2da066218b3b9290af4
zf44764f84b556a8996f2efb1b222b05c402aab8c8e0ffcaadfe1b6236922d71d826f226e371263
zb9f3e5c46d9c38380795493a04ff662e6a8cbcf16d19a3decf5c0c8209d8ac2ccba1363a22a722
z032a131eb02af7668af7ebeeddc9aedc639593dc933e603563725ffe6a160bd1011d8f0a6ba66b
z9a65aaa1c69faf07a56fc959ca1e402f0f00ad2f6170b3a90628184cd5d567eb17bfc6677c4dee
z9a084512e315b142b5a6124ec4b48312afcfcd7332d6bfe1ddfcbfcbb79364a7c98c1ff7036d37
z67c984170fca3503b411e7264c64a4739b0f0d1236e33b03197eccfd3aa76985befb522c5d2bca
zd221fb28f1183ed27aa993d4ec065632aadc05a39099cd602e5a0bb74a758e3a23c2798624f17e
za2df42d1e5e519e97e9c9e2d126f7a6546407a87d87f47997a0d00fa9752951abce3ddc7ae1264
z300617461641e2a65a1b1e965004f7f0700bef16ad5aaf4e28238256af21d87e558432692aa5be
z975f8186b5e2c742a7494863955af09cdb94ac70b008292645848e4afe2c01d6b001717f492a48
z94e2d7c36d2290c2fefcd206abb13a731b021b931ac80e10785edafe41bb437a3f0e4a84ac06c7
z42909eaf618764a336ac661a4419fe62a05f9d8c196ed99eb07c7b037cd80db9d2eb643131b273
zb7c6ebf04c3b623ed9cc7b997a9c121ed1fb57e7f6ce32c6c8cdde7b18ae8ca85a65a2ce2bab68
z0144ce1ea6a64b2aa5130476ca38bf2063f43d2e3a1908fd6e1cfcf1e99e46c5cd953e6cdc4a2c
z4abd32c8ec5fbfe46d33eb27330b7b1a6f8ae26e9c1b0d1f5345d8a6a12226d646b77ce51c4b66
zef97162fef2c04bd455649a26f665ec5f117ea66b245e432b357ab6a97022a7793a5cec8f37062
z6980bfc1d62562eb3a83589edee48ede7870e3fae548b7f5d54c3a783a5582a132df4e2408b36e
z811cd6bd8379c559d3d63827f0788be8fc2d3b44c9781d93471128a49f8d90034a5ab0ba3a0c76
z13b2f358f0a4979946d4506c5f424f416783d375ba7edf831eecc2b4206760d3a7a0af572b2769
z01746d9f3edb2defc69053fc2089875c98cc4d6de440af80d0ab729d138cdce1d0f809d33b19e3
z3a061425dd0e3b924ff3cae8236e13be693e08c48f72aad2ed29e2afd21486ed642bff9cabdab9
z7ec388668e190a6aaed7223e6fc350a3e4f8284da3abf2a083a9123372ca0ef9051a065b710cda
z4debfbea4e960fcab94c24f912992cc6d8e9d057327770e36d57c941e1bac40f864cbdc750ef9a
z0818aa31e00ffbbaf92e47b178a5f0219b1156d19389a1265585d93881de8e016cd131f4a0bbb5
z6663d1844cfd597c72048bf415219059b755340aa8e6dea13adc4805b7f84afdbe4f07c70b5f6d
zdf407845be171da5112404c32e10318d64d44bfdb59d4ade68ced0ca1902bfa20289ea6c5d8226
z2fde4c8acce6614b476ea4d39cc0f44727e7092373c2ef3e80d4b27465b671539a61e650d4b503
z03fa6a6f1a318c1cc35f59e7ccfb4a3b4377751a4f758162fa0235aec957c1741e644c93fe73e6
ze4f505222796c349925afb6ff0478a36fe8adacfb8e0650b6279b0758e27f985f3cdb3a8690f1e
z4cb213bd699c3e050a5d0be153c0f4263ab4a6b42c2c377f9b598fb08c645f1e27b8d5c8b1b9fc
z26404c397c556982a56cad44fea6ed34883a8fad498812b52222128cfe1b588a67c4970c9e0386
z4635258a83452ee8e447d1afb3034114b56ecdfaa35c7b77f1ef7e846d3433fad9df26d0152ccb
z79af41a1145052b252d79b9ab4339d0490d5e789ea36587d8596517fe397dcec01dee8971d2244
z5d69a1fba10da75a92ce7293254ef96a88ab82dce7d66506dc90705784266b334e8c11a2d2dbb0
z032442c661a96f9fc9bf11a243d0b57f6517f5288f31c7a4e09aea19c3a7c676956f04fbb6e92b
zf6e1687cfd15c76e1f6ebdb3b0b8576c9164b21dfb2e5bd71427b0035ad5134d374c40ba3ed6b9
za9cdb2ee28d826a06476a29c4c9c0d411004c0f2908f6953c2e7833959084db68a12c6ef304a0e
za724fdfaf78e1139debc48019b1c93cc3fbab8010bef82086d84819b9a9c2a996e87db7ef6f69b
z338325e1325970f226fe271c1355d489b37c42eb28144f8ef75d62b570cfb9a37b0acbbedf7939
z794f178d630fd2efb1d1e216814a004ce7d8d0e02a170b697baa6c05de787c84188c688aa1cebd
z596740bdddb62c6e209ee9772b6ba1eca78506ed55e0f409edc4e4ef155b5f3c854d6da9557169
zd2448f71854ef050f1b9ac7d46bb4484ed0793bd00f3499bbb102a17c9aedce0db1ee7758b7900
zd661cd046d6a881716fb2f590d303b180bbe5459400be4a0106997984615f2ca959c3192be5411
zcaf5b6ad6e065c88977482e8ccc91315f12e72483cfacbeea27c2183714ee9a861ac518cdc4c07
z28dc3201e42938cf4d3abd8b1a79bcffd9aecfe122a08ba877907321287b7b47ef5930ff7f8f12
zb9a09c1e57e7eca92ce4c0df9b7bc206053a30d760435b4b52d017e0528549d49b62932e770e4f
zf99b2c5596b9c3c05431abcf345cb99260bc0712b5c8d34992e07dcee9a025c1c428e770852152
z407789645b1f9794219db017c0d1a27c7439ca10bf63047cc04d7ef0a8d88d44ed57590f411520
z5f4c22e0994f077be17bd0d5c5f40c740b7763565ba23b205d56ed90c0ad64dc1eb17f72a3cf22
z4aca1256cb461838472951128a766c420413d8c76943955f74199f16459ead9dc2cb5c1ca6d8dd
z992d220cf8beb950136e7a2281259a2943e28bb60e43f4d6f155d382e4ec630f4b86a5247d01ab
z63740342c6649adcd91b7690b32e3620b859a4fc1a733232c304a2b16184221e99c055c1bfffe0
z616bcecf5fd190f3ed53ffd71b8d4164604ac09c52dba4a4458b7f80f47a7e051dbbecab8a79a0
z2117e560894808b6f8fbf507f7971a7c5c1554ff488f808a9315d47118e913953163c41d3238c9
z7819350000dc72e4e83f56ee865e9b9517232651adcdd89074267585793e30a36dce12b2f1f12a
za1e9244cb1a773f6a70d7aac3dd45f318c92b6650a4a27a05784f6d3ea2fbc8964017901231b3a
zafa93a26ec407092656dd350aeb59511bebef9d81b6d6acc2cf2e07761089463de38a8f3ed4f5f
z0ee108e720db79c3bb6097efa7d61d94ab34eefa31a9c9e3c844cf146487c236e390a7339f29c2
z9d0daa1986950db98fb159e797c9a8ab718b1cd186834f8bb945fe17c920fdacda04d596a6aa3e
zcc3e5fbfc287e6c1cb63e89a74797212c5cd374d15b21cfb605e154ba3ecbd693598af8216c8df
z91d947239044fd1e6b193cf5eb7e9bb57c28372fb091b2eba18bbd9c3fd1cd1ccf305f490e5835
z1cae70b57e80b36d785f4b93f442dd1caa2d44812539394e3891ded36b24968855092967e6aea4
zf8b48fee4b7dd3faa9113b87fff9f3a6e501c0b7c89e338a6ccf6f0eac67a00afe06119950d11c
zdd46142b8e8b954f7f8f1b324e4bfc99d2a7a029db342754dec68bd34d1a12c9ab4922e3cff89c
z94622e331cbfd07c3cb0902001d2a292d4356510fd6fb42fea584f5fc248e38de397e3d5aff6c2
z948bc0e09cddb10bba993c502e1fe665daa9135e5390d29bc48a8a576ba81ddf5fb7150ea8b453
z5f8850543c3234871a718c2fa2c439f5d184b744fbc6ac2ec3b9ae629098b7e1d03d202af6b0c3
z0e0d5f1c5ea6823c840b381a0d2073cd45afb53ba28f963fab7b5468311ffdc0aa8b48cff78aad
zb52a6f22ccd83bef1ec399a1bb2dcdcc266bbd14692cc50e47501ea7a6dc10e7f597bd77a4cb72
z6b8bdd6c9ce2e80d6912d84d6eb5cad617f97863e18ada32e8b9cab9d34c179d0ade10c9d06b02
z6a19c16c11ab4a0099af2caad9bb05c64e0b2abcdfb9db9e3d162402b1324a2a3e93263aafbb66
z99c176abee82ac478344dac5437a33468942b85bc7400d78619cd893bf2731cf4ae4d5b6b1cdec
zb41b933a63c92a430bf42ee2dd05f62f5028013bbbe8cb37a5e0bdf37a6702de693aaf8ce23bdb
z145e9dc2d57c2b7319adc41f55c0a8f124a804abcc04a7478c6a01f1afa645e57557e4403dcd99
z2ebe9c185150b6edecd137aa8013f3f0ba4b82e6cf4f3991d27e7eb25f8fb5a03cd381f9092901
z7d3472bdbda8e9f957ab866ab5c9cacdd628db71b80a3f570dd661bf80550881aa0d8bdfbfbb9f
zc1b0070527507252d68e2c4f6efbb8905d3a4c92f0888f7f7000a0d4c63b29918615c96ddd8b76
zad7b740abb2d075de2cf5d2889dec1ae01fea174a2cb211e9a630d3bd0b538f14f4f4984fbfa29
z23204d20b90f61c27604dcf0589ec637e77ff5dd57f3ff904b269ad4e12bb284e99c625bf2d1f9
zca9e6e319a09f8f27b0fadc44277319ff0f30927d1057756fb9aff69c0c9b3894bb36e852dd7d0
z91de9372377b272b39f212883074ed4bee73dc39c2d1125d27802788d786ace63495b33e93f795
z22b37dab68e34a0b978451ead07d5148ff6ae5dd6ee009d2d382c3e78a39ec19e16da820e706e9
z83a0a116c7cf9a93def73d29a5484919b2d3eb1836fa34cac3138b3820ea96eefb136e3863c3a2
z4f3a1fedb9cddf7a9c0a65f0a8a62fdfaa68358e58017c88eea82e4672800d69cd25079f3d4d6f
zfb5c377a4bec0ef706f8851cd64ed287f5acd117ae433bf60367ec33c31e75725a96fe8009bf05
zf9ee940025aadb0bb64dfdcfb34a17d033672997efc0890189b3eeb3a53f72839a4f02d6df266b
z965cbec5e25a562d2c416d1cf36155439d9ed5fc2cae0d9700c13d6b3243aded533e66cd0ad539
zf34aea46ed3ff96416b3f80804ebd24760b239074eadbcee523d3468b2b7a1d9682eb2585ea84f
z0964a0dc612497b77c8dd6eab651ee696c88c2ab6851071db5c1fdd06262905176e3f2d3fbfc2c
zf16a1d6b3c97c8c7c5c9a026ff7f137dfc92c648c9570d65c272ec0eca408ef9b026d0263d3967
z86dc4642368a09bba45a05fbdda9fcdce558de7d3a2ef72b317b5d2e0410af5dc1d5c7ace5d607
z46bdc73889490a343ad68cf9c29c19ad71171e1533fe1ae46a9cd6e074c2ea9b41070e39fff5ae
z4febc44d577b00f837ab98436bebf3c93ca2b27192f7cd09048b885b487b8db0434e7be59de26b
z6be39208bcb3904534e6cc23f0bf346e01ccc9960a15cd626c8f5334341823effedc299682e82e
z11d0c17964143085c3a432cd552c05d3cf986c618897b32710cd199fac8a5dc68bdb7766fc3ea6
z75ca2f3421356a15f215c745e6ec06f412cdea378a9a6a29da7b4560aa82ed1531cbf5abff2415
zc4ad59575248b5415c1d3a57229c00724b61451cb25b8610f61f140b6cca652b9663884447331c
zff278d98f419b850032d5b564b8dea692e4d8c8d84409ca522d75b419a5fb4bbdc7eddf4ecc4d2
z2a6c81f49b59eb971418048e3391f2dd28e8e3802f4f31950cea8e7beeaeeed4825eb7b178e542
z6b6536219b44a941a188d53faa012978d3f704ba5384075cbc7966923ee59706c3a401c6944fc8
zb431b05624937f5de762d3ac474ea6e1b4c6cec6a64075be15b0900b0881acfc7a1e515df13dbb
z91c25e6d122686439824da1bcf83b0e1bf02cd458fa21cbc8751523d8165f616ebb37e5ff91d29
z4f265b857df1d2643063e04ad8ad5476a5720e15876aac3e86ed9fbe0dc69ed5fa19a7b852f8f8
zdcbe3dc88da0e5034361364b8c0848c11528b5176ecf4d75824ddc9fc2805efdd568d669c14c36
z2ec76c32d30cca3ace56bcc60d8637fb61acdf4190b59531d9744b7dc7ffe1bf0a64a21b75a227
z1b74c0a24fd271cd00b82c1c1ad12eff8eddeeb5f79490263c6d4bf48a6b32ab3ce2263db4c993
zaa17b535a5d3ce7e227aa68c9c009a8990dfdb591a913fc036341d84f1688a2f30cf1ffffc5c1a
zf2ee1d5f679e818fefac30da94abfc2b25004d4d244e984e4de8abdf893a7b0a962117a82b5b73
z67e8da46c29db19badac3f35ad4c20501e490142287de4f1ef04525e9f3fea6213f969cf549e61
z5bc142525b1271b106c45ffe0fa0697f5a903a01ede399160a5f07343bd5ac19f0deb438266364
z91255344aa339c2a82b9e5b2cab483f92d825671a267f4fb8015371427961ba550d7b24eef76ae
z94010238cb1d1c09f7bbc4d8f093c57a6e9490005f24ab69814e2b5c5a9f475aa592c5a39b8aab
z219d5172539b214a9e14b79502e412c3175f5e95695711048f7a67c958863d9f7b7b7e46ce4b26
z05eaa009f94afeda1720e6ee954b7d9257e5f5cddf162cdb52b11d3606cc1ca2d61b66259d1a58
z5f679ceaba9b722ecdde759b5179c7e1a0cdeeafdfe25ed3ede286f1ac2f9923820d6be36c48e0
ze5bc463880f0d58a0b7e0a450074c8b025b7a4c8198480f71b2b80eb88284206704447ee41025c
za6167225ac17c4f587d33380f60dabb15cb73708e49cc9e6baf699f6a8bc1e4e350fde8d1dab13
z1094eb606f257f3720938ff069cf51a619252b12109c890da99c3a09f0f6e91abab1efe2a20dce
za97fbdf9196f4b6dd20038d38fd2685620312909c7257c3b9c0c5fa82c75386f932ef36d5b9f4d
z7d0312de0dd8a794792ae9f2b0b88c7f3761bb07a473466465d24cfd56962a962b51d052a3a1aa
z33d7378d9c2f7498628d71907d8aef15156b8bc3e6a01c9e8d5c1bb7c4886b129e018aaa79e606
z7ef3aa027bb85e396dedf1d4a3ffd876f930b664574b7cb92b8660c1aa6853f2e39981f4f301fa
z1251cc9c8cd1015643ffd50e6d75c0c0213bf977866c7d29e47e0a0e3840ae20bf9ab71192b147
z822e33bdff803a26e3de9991135dbf101b84d14549f3e1b67a87324a7ae802652e0b14042472c2
z6796b8c59e29b334aaf31717215e87d5c2aca448f0990bf30ff1257e3151fcecee8d69d316f598
zfb268c8fe4c1249c4030754ab85c3ef50f90deca4848dca880f0cf55be2770e4396cdc5cbd3c6d
za88ca1475bdf54f75945e2b363b77310dadeb5de874e057e557821867ca0dfb70bf00fc54d8391
zdcb5af2728e126fc0c4f8b88862ab200432010569d585bad149611e3a69531e131fb16f095ca5c
z5f7c7a2f7af1c8821e8b79ad8a14052f140f24b74bc85d3745de453215912e051b21237c752e6c
zcaa069bcfe6a586ffba4e470656f736744b142267efa9fcd3857c40c882ddb5ba5f97d6c2c5da9
zc30625f3de9d2400611d0696595d7fada3823d973a561e6860ce092fdeb90be934aa6aec7a15cb
za560cb9abd32fdaecd6f65f1977520cbc719b1522412be39e7166f4705686d752d7e7c45b9aadf
z577fd7ea97066d26d2d7311081fc587a3f122eef05a902ff75ac31d0fb986421b308cec5b6c0b2
z882a61fcea6761b38aabfebe45c540d0acd2d64ef1936aa1e95654d86feaeebe62f341f553a24a
zbb93b53613dc64fb990f4f3a62518082811f16d401354a9fc0d4e749bddbeb1192ce9c4188bfe5
z8e95217775015c0cfc1c58fd5af9c0be6a071532929ee38b90072d58f67244e62306cfcb54ebbe
ze638a950c9dca199c94816aa36341341dd3822ae1d8ca90979a786274cd04117afd3aeb4452ad5
z6d9a51b8fc5f776a9be78b04d83eca4810d8511344d882623e05699829afcb4328e0c2563c2c4e
zfdd1f26fadaaa12916911daf9c7c15dd8281c1042aba3b80e7205315c7ae123e61988a1a4aa2f5
zc3be28c5705889ffc7ead5b219c593af186f303d3c2e9600ec525af3a07b3368fd8ca468b3a742
zf7cf1169daae80139a39489ac8070b4552edc8527a5c59e39f298ddfff1ae0bade75cf284e6896
z972fd1cf2e28b02389a5758d67745f391fd545640c28429cb10f68e2f9dda253fab2e1090a717d
z0d66749e79dc12bdd5dc2292e532a529ad369bfe83cdcbcd47a3952e8044d2de2090293c0365b9
z286e11742cf20b0d935aabf9ee79979c029f336b1c56c375fb2188d18762ae8f67167a95414de0
z44513b6f884e9c3fb5dfbc1345d244978be9670ca95334b54fd738ce16e36da0a78f8a63080d04
z925c8c87d63c7b345d7fddcab1b8f665f85d742203173c45a24a8232a0e1940060227673c55928
z2671eb8bb6df3d79e125c0c65321457eb6ab494d4e26feaa33fa6ae36455b40a5437e0519f5d48
z5c026df1dd917f30ff747546862476bd9795ed27e576ab416322917705a86b2a1b6fad80934c2f
z7cb6873cda4520f12f828d760342f31121e2da6d837943b2a57fa125fb1f33a3e379effbcda131
z20070dad87a2b348afaee5f0e34245b75fabdd41c2c8c1a5ca727f75d20ca55172439d6859de63
z00e363505de9dae1e5f025b81cef8e6222afa111945bfe8331c5ba7eb8b54dcfb665cefdc8a3cb
zfc35285f16843d8c9e005c1b396bdfa7fecb1263fbea5417096c984372fa0b37b49a8d1665d180
z4a50cb85072fac2df7af585a11f2ad40e7e76cc97e519b75720c4c7d05b9996eefc944e9cef671
z3d03618fe9651ea596f33ae003003e6e1e862b4d63f33b9074c301dfb55a9bb8f8277b29eaa705
z2427f2872194192b02379b2fc6154f2a16a87bd0a2cf6d62f38eabb9da19cb5691e59983abcbd8
za7affce0384befaba216d04294a91535df43d50dfc8c0fde187b3851f6133d8f58114cef12399d
z127faa8d5bbcaeee29378ed7d8671c3d6e6621ee6edd1b098071936fe39c210fdfe64c1f69641e
ze15f2d0b2e340cdee620346b7290ec9ea91429d42c0fb9318c6a4beb132d767a51b79bf2f9051b
zf092df1f1909b9b4e70ab107e0fca033b37ecf101ddced433473fec4e363d3a257ee5de144092a
z752de4f734b0bb52a6b0c14fefba837731ff3f485b81c3811df0d337cda2bf9c2760e9cfb3f9ea
z35cd85bfefca6be462b09b9a1b2efec2d9f8ffc0eb29b4ce1642301d67dd83d3af4177a3d2d467
z43a7cfa680afd581b6461df5e8120fc1bbc09ff896ac3877fe5530f03774d47ed12f628095e4ba
z36f46e7d697451d9d2400b9d7aaae46bcd29f1677be6a8f68a84c9a6f9b8d6d4fe2fe1c7f9217e
z74aeaa34307c9c641db2769034463224bfb05e8e5dc748fda1616b96f05c8772def6affe6786fd
z5892fe19a57adb55c5785dd0895ca75002c62853be48b61b3f8ee72463d593ce46395c28ace303
z8e1a05633227967dee49563859ebdab43cc4ceddb1c3a6c59e770f6afa14c2bd21f927f4ab6531
z6686d9d30d6bb77a2f663266093d63ebbe87416351bfce9996058f5c17752f58e83562c9b95134
z198ccf951275fe127bd7c725ac1017555ceaf752fa0da04395bb9bb9da423218271f604ae44203
z94bf7c1c9af7dd11f21e7bee79a569e56cb4106d444d2018fa652e7af7aadca42367ea0fa2e67c
z8f4ad82398c6d81757d12c1cdaddb01b9856b60de0d4870c4c1a38cca1e3b4802a5a618b76cd3e
z568c5ad5d272abb4c0b79c70032831482c4564b0456aa20d4e5ed6d2416c102c4f9f38fc4cd080
z8883c3b8fa928f38bc36cd0d25c01650d9dd547853bd69fcb6a5dacae5a7d1429668df725e2049
z32e74f198821160b37713055e7d860b2530232dbf1ead6030a7f23b89f99bfbad304d5dd0e7ddc
zb5b25b020fd7e6df4f318df59765044e8cee1fa8b2b738820aed51d9f278a83bb342f70d2b1729
z93afc04f50fe2259a5d49b92c78d941072874844a3bb20f1169e660a6167159a0494a519419d2b
zff2d4d6129d770377469257c31a812a8b2678bce393e9c5b825e208b5d4cae7e503501f5300cca
z451e5281cd07c54f9d14d904555f54dc307fa53ea68e2d2745e62fa1d49e6e51a8c85306016c40
z3470f9f4c931b897e06e6f3d5751f3026ce976edbc7496748b972c533e26f6151e8d158c4998c9
zd8e50e4096a0c70156291fefe7007a337eea7b24ffbc806723954a780b23f5f0152f03a7af0ee4
z6db8d4ed27fb9d454790c17dab39fb0444d110937cef2e6e4df18e560202bd9a0a62167288adb5
zc04a5a858e0ca85a319593da504264c55cca57905e1f7fc8c69b6af276bd9f1299951340ebf535
z371c74d315d39693f55b7dac78bf4134563f78039228c6761b7931a51902ec61c2d3f653257c5b
z08095c5ea53e6fb88a82b7c53b97ceb4990c542c381e63213a00758ecc274056fd2b59b60d587e
z201ecd89369fed50b535912a2d5d660e1a308a9dd070e17f22df921415898d56507b8bbac42c84
zdf6e5f09b6f429002e541df1e45147542412cb7424070ec4cf6e2e570e007e8f58281d65f8f856
z45adf773c2b83a5eecfa30956527eeaca2758a36099c94451a4ab9ceda06e68884459377a0d31e
zd856d24e074e1618fda66e41b0c2489665c23e6b732ab3eb08bc0c43683c5025513d4b2d55b73d
z8f94310b336722a41f516c8ee49d12221cf4ca0edf7c9bd5375116b79393c6d3892d97c80f327f
z3cb2860abdb909cf0691c4d675e3d2be379a57d5f3a16a0a4bff8196bbc9b8af10df2cdea0f032
z07c6b1684f0b1caedc85cffe36ee104a370868e64ebe926e8e72f22a9494367452bbdea4822af0
zc116395732c98b49abd07e1fa8ad366d4267db00fdb7f9c5a7309a114626efccf6fee7f6015046
zdfcef2d72bf3b8007834ca7c04958c183a8d7d8f987c32856d47f21d8d66f00db7eab1fbd6057a
z97b0b06f164afe55078d1d597e32d982c74bd7cc0e57cd09dabd2be26641b927d2f679d065c598
z1069bca72506c8161b15837c95cbea7de5968f34848f2377fdee302591dc1b70d9e92539e49500
zc5bd5b9b73ef4b1c069c8b479b70fd0bbcc7d97d874c7c6df453ef6e7cd6d6d80aadc4d8e91284
z9ba18774340982273226b7ea57280861572b083400895acab0a2be8167c98485ff56a5b305e3d7
z74c5abf3bc24940b8383d8281df0d4e9f1b50a1e4f6296f34df84b8117d91bf6bc8dc6ca1f76b0
z711cc25901f5055f7d897a4beb7b9ecc0869726ffdf3718d6fbacb75fb7c7c11b647598bedb078
z21231992d7507d1ca3c254b2283e85c4c7fa77db13bda6882fe645674ab2c5f4ba87d9300d20e9
zf6b347618f09d4dc94205066cc534c970d4fdea34e7ccfa313028588ca03f78652935036ee7a96
z20bda39be286ce4fb9e6f6fd48f1ad006258580be5cfe28bb83a477bb59ddc7d6a26d99d116b58
z93a69b447af9378ae142c37cd79503c42bc625be3b4a8d7a0dcd1c108e3bebfbc5cb7d7a123bab
zddb58d40bca595dd104817f586255c93880172b7cfa1e1d409ff95e7f9c15013904e052ef76887
zd52f2ffa7f787c4ca6c70a4227592b5d4ff8a6e4ede1faf5dcf717b0196e1eb9a09ff38a3f1056
zc11d9e3938770f363fcf9efdbd0d67fe0bd28b66aedb44404bf990c2fdc1872ee5251a3d37d898
z7448fd30fbe5430eb6f06b21b483367982d1abd63c53b953a1123a3f7d77c5bfba7fcf855e5349
zb7d77fa50af2fd6297bd606d6be09c41af70709f7916f6f4561d4975c9051cb0b4d69e4b8856ae
z4ef7301ffa59499ef805dde4f47c75c8b8f4b965754bd92037e18bb3bdc7a8d396ee95193b84ed
zbefd65645fdb45bbcacad527adc941758439f46498f13d6e2518bcf4490e271ce443d0bbaf9988
z717bdb83f4a76e8676385d8de86b44b12b554810faf7f5766c88596d8208ddbd737cfbaa23051f
zb7fa56b0c115c0483adebef2894a24b61d0bd4a460e6fd9ef2d224c53ee89b6d54611a586b803f
zad6fef3f785b8d9c96912864cc850b0370533db0a46b21b27988e6f4593fac09e5cbe677919d22
zbdb68f161270e80377d6982e3cd2afa9d53ac7a1a27ac0c91fe68360333d7c3218eaa7c141831c
za1d0477077bd8b760f6bb215a3fb4b87c746157b26f903dbb38a44b617f6cd0c106af993fb0509
zf182d9c9ac498cfb122f6358fb477a984d9ab4b91d7306ccb63017ac84cd247546d2b5bb1c67b5
ze5e829bd51f0b5a92cdb90292b1128c9a1257f0151227e318b6e0adc855890a238a86f80dd849b
zb1d3a2b53e3d2fc0a656e23d82076ea9b5d0c057fc9670d9fa6166dae268e38dff2304a6bebb23
z0e8bf72099c709e88a445eab47ec7931f548cb121d83d7050faec8c49dfbb333eb2379bbcd474d
zba204f8599cf8139321abcc423ed577107b310bec31a362359b3df3213cb59b4ff4e50aeac9e60
z12065f079347974d85683bef54876e00211a103685f30565716542217ed187f800cf26c6dac554
zd3fd213e959730b748b9ce74d48e0d659a408777f882ab27ee331709407ff712ab8f8b528db841
zfcce51b7ecc2365f3a8cf96c9fa7d013778a1a3717208b9fef3d1841501e8d9f8ba763be9942d0
z2ffdbc271639034b383a6e065393e50adc88ba609fad82c5387a09a0d6d2f48fa1c9650b0c0213
za10f0c54f16ded8456b2b5ccc0dd36654a62594e6cae0827c9730683b0e08fa2577eabec59779c
z041f1e141daec7b232f9396c42f4cf73832dc9db09c3671bccdda1030231a00ea471c522882992
zf1a862d47df04adba9aad948e850cc98c334a8d63ff989f71e197895a58ef31ddc6c5dcc956616
z25d159decb2df5124527d9390d96cefac256520bb8cb6ce7cfa0f80964e6002d47e79305d36d22
z9add4b9480be9cce631c13094deadc1b5954e148d4091a64c5956cd3d0f19af4f290422a4343ec
z9d2ab7859c96a57bbe7eb678d510af239156a8b4ac18d34387332f9f1429bb932f6f007b391cb9
z3a6f03aa4853f5d0a988c5949f993c6a16f9e61fda32ba21a0747a9d85a368494d143c87c39d95
zbd5fa3db084a11c9f2513c17827570d481a6bc664be323b75949b63d0d9a93c1e78f2e65ce8c14
z6c58be4294b9b50bd6699162e16e8efcdc06f72bd3957520449e0f330fd625f8bf9f174ccb8e4a
z8b71d8045cbe4bcdd7d988249a8e03708e8606147df70e91a992878882de5ed93d93ae9caa78ae
z59d279f554bf15160ba33f9194c782ff776e5fc2910d848724703ab9229e4b0303eeafd64f5dcc
z1c229c30c984039cdf6301f26d19aabf1507ae5d701eb73db1f15ffe1bcf3fed339996ccecfddd
z1caad5e8fbb1574df122d38541d9b067512da6d12bcc27740c6a3b8c6d42492ea03426c17999bc
z914db015c681f34b9e4552644b92656797a2a3cb660b936c479c111a28c7622e0a415bd5c962cd
z248510abfe4d2441c5a9fa6106ddee25770567c9cecc30a87c9a45bf1400ff20d4e26e47c3a7ac
z4d0116fd32d198c17361d4326a822484853d0ed62d8af14d3e2c3c42f01049c8d37f3cab209bf3
z7071b72bb010133e95f648dde4a7026d84a839cbc6eb12714c711f57218822432e08eb02ced04e
z8e4a2ad80e5de527c840fa04fef8a66a62dd6010dc737ccad56ad9f79bc53566259c09511e7676
z48516493c54353cf912a4b0cdf76c9e206b1e86b3023ea63055825a56d2a667f7a9524fcd5ac7b
z42c33c945b394a81194230228e058077648a22294987cbb1b499477b7dfbeaa6954301e62efd49
zd38366a01921845a671f702d3681c83fcd6c7af3357a63d050edebf9747c11037655d223e7cad6
z4f2016cd7938e53cff3cead537eb61c99b0164ba0734208de4f6426266ae7ed4a67c01abae3f94
z222e1c055dbd727290957ee6e72b35f4735393d0a1d022acbdc45e3b7fc2e91aca95a5552520b1
zfa47c167aec118d327281c0038a40ae0d7e287f5279101ddecf405833f79e9dd6e3ea020fa7c56
zc58fe2d4f8b60bec91184b97cf5f01f5dacd718a73f8232ef9b9ef17d508f0cb62cecb9571c2fc
zfa42b031c80172d32c524471a28f10b59e9f71d0d129efb8c56ccc7db15bc2e6491c46f82aa793
z6defa29da0e7e49b9b32e121dc9ed7f00437839252eae06266f5078174361a9f840a88ca833601
zd03657afdc948c0b79c74f3679dfb3e4037f4ea18b320994588e595828fa45ced55f24216f9e73
z4ee31593abe3e04c862706b7e66ab1cce4cca79dc1f3cb62a6bc136e341c2c0360a8bf9fda1ea2
z4cdadd42b233fd718bcc62be4db903f220d5ac0a47db99ca041f5641e356702e8a451deb2bb7e4
z9e56160c8f02c85ccfaa641fd7f7a63b5d192885e0069648ac110308939e6322ea74e414e0e138
zfab439b5682901601c2157939379efebf33b0e702bead4f67bfcab37054039efd960964c7f2848
z8d277d695614f327feb365fab6f9d35652b42180dcc68a75b8001b0aeb45b09104fa8f6107e4e3
z58ef52aea0be68057647c241fa6462d7c19fb1daf522deaf01ca9c382d592c54b5e5159a276b3b
z123a3daba37683373fa85732e11fb1715f5f7174da1102fb8f13d58428158ac8fb1d3592381545
z3c602fc4371082d351071c7ac7d913a95c647b61383e49093b92ceda1aee8600a4a67f80776cb5
z89e9a93996218fad94cf27c7951dd164cb9c53f218e5e173b1ace2f2f52783e2f0b441b23c6bdf
z058a1316b552cf4bbc7cd1623129fc0c0b36b216d7c628f154a0c21e827346080959d1d1d0205b
z4cfc3b6f935f281e9ed317828fde2d764b6b3d875cf98d50460fc2e46b24d9b01deecb530ec1e1
z1a8409af2fba2deabef3098a3d7ddf71694281b5b1ada823257da05465a2b408cdbe848c5cf40e
zfbca2e85ea024d65c444386da5c8251970f98f50c130db45a19ad6610c8e9c8ed3583ca6833125
z712e1a04255bbd44af0bd844fb82a0e152988a1ad530061c8d0879f7498b6d8a2dcb9ac4623d2d
zd926f70a822d799b138e3f219cfdcb6112afa48c40743bbae675b6b4d06fe08ee3468b2627942f
z8bdc8c7247c28df93909b72d36e56e49716e4cb88111201a6b2d605bad9c4e63d5c34e83eb6732
z3672896d9da4236a6875616b40f779de014586d90c92a35e380e612768a985093f4397f7784f9a
zf40d2fa2de0040d37669a8ab6e7f6aaf894638af5222a5183de99d53a2d87d638589da5fb28734
z89e77c8bf1159693189e9140d9477255641bf6b85260376a47fead5504f8c9508be8cf019aa4dd
zb1d00bc5a8ee99be50a3aebd3b45e5e6f4ffd6690f853f9ad464895ff15428aa151e6d5858f10c
z55be021206c1ccb3f0755593e5b6fffd97ca6a4a17b4351327320fd69ff82042d638b67695484a
z6604da52661d10be8b132288cf4a0ed5ef688c74b6657392fac73c01aaf50f3174d4ae00df18d2
z3fe1ac3442995b4e9507ff4d423bc896173dd3653378d6ef6931b5099e590c814e60ae121eeddb
z9bea6c80e7d12212b58ba134a7ebccb8a7c8c635797dfa657cd9dc85dba26440edca81139388a5
z54b35b2ed948d479289d609bb5e4aa3b98cb3460ebd596d22e384858b7e47247ea30f86017bfb2
z5b8db18624bb29c08ec9961e9d4cfd85e329569a093ab2728d0a031bb2c604a9001c8bc42efe37
z15c8159ffa8e7602f2f3c1bbc35db569fcf2d14235be50f2d3b37a4d2c42965e6bf956dd3bd321
z3fbe8e7a69cf40577b6437f888f35307c7350468602d8163f6f0de69af54568012ceb49db7e20b
z8eabafc3095b4830af6945dda0a8c13a6806272f6299955fd16ca29640b56e8b53477fc537678b
z8471e67810dd81d64b6ceac53e6d490f260eb5ec057e82cab207b0ec827ed043992f7a0307741e
z4fc2a4500be031135b330947eec1dbaddadd494eb80b78a9da9e8116483f2a79000cec847980d4
z77c4a819722f5234fcfa012e4977c068499346cf2caec5e21cd22ecd6ca33dfb1f011508236e16
z6cca162f73ce028fc339090131c4fcbaafcf2a762d75062c25131e810a6d851867ca1057d3ddc5
z72c534a2a1eda4b1e67737643b6f90aefa518767f858479d2633430bf36547f52955f6ec061217
z1bcdcbda05ce03cda3d5e17980b71d5e11712ab9863c37aeb73a3edc582e0453398f7b50097e14
ze2e3542735810427c2c8c1285919e3af6b530263a40c19bf320a49b52480ac4c8c0de4ea2161b5
z8d62f4de37e77b0e8405349bb1c47c7738f799207dc306ab7130e09177a8fd3ea188ae4e93d68a
z9e66ad89258d6422d3af62b671feaa1f93f72b37113530a6a23a87aa6f0f394a130f29f47e1a79
z774124818d922b2ba390c6c06e61a618b7742d4c2166b3f05275b3f0005dbf531f6c5e2a40be8e
zc34a1c1122fcd2177b4da1936951b66f5a312ad3c046bd03338dfebc919d754b8dfcabdd4a2582
z468858cb9bcda7d19092c074a63c2dc627f387a895450e4626c0655bea6c4c25ccd2aba07656a7
z38072de68e57cdb59949cf55c0429d7e0cc344178e0198999d0a5a38fcd4dfbd9ea3137d422bdf
z0ec35b7fbc1bcd235988013d474658cee7f2a8347800c34e1773b39d1441b2b2c197572cc9e487
z0e18928d3a318f45d2bccb3c86095f24237dd95a80c4c787c6a6be0c7a78621e011aba4c7ee164
ze9beaaded796691d1a2ba3e4bcd5fef6d2d3e76828f207861628c20885d5de31255b00e8109109
z7eb705979840493bee9b85ec7fd261cb76eba902ebc614025a7edf509e0bbdaadf6d32846b96f7
z368bb1535e3dd03bb1aa08299ab71639feb9674b3d97946e8009987429d213b2aef7b0158a6e8f
z4aa41b0a4de1f77e75b9e50d65b07a9cda1b89f292c58b551d71314005642b2eab35af6ef28231
z5e96e9dadb9884e96992bca2e8b2456311b232af934f3361fe9868bb0ae3ac37d1c4349cf63790
z702107b5385843275436990c429f293b5cd63bdc091a178e36a55d0e67758b284b9c77b4bc0578
z2d4011a5110e8bf57176fcfca19f7de8e196414433e28876a611d8180c5a4e7d97c1dcd5772acd
zcbb454db814c847ea0d0316935e463d1d0da5108cc46761cfed214ceabc6d67247ecc54b338135
z7e63d2b637664e23e103a0ff55edff41f4af9ee386a9faefc65c6e3638b40b8de97431ee1616f6
zb20046946864b7010229ee87d1211f3a31594d2a375e398535f90df36ed77a0a78318fd74a9c4f
ze95cd2d2b3b91efd131aac8553d99dfcbb995d0924a1857c7b6015c2e43721caeb2edd8c9b43ae
z63f462e70cfb31385d12f52a6673fb33a2c72b314509199a87be5e060bc79ff386d5187f05add2
z5f32a396c30373b6902925f697d20970532e5c2283e319b5263228e4edc8ae078e05e9f3a9e46d
z25fe758a1d4d28f42a6272f9ec107e8f263d3e57254e26cd8a99f0907872a0ddf72aa5a420071e
zfa4874e3001af23c5e923ff15c1d774683a0fcc24e9cfb62482f2d28455dd362edcd8706d5ec9a
zfa06a09c1ea0c436ad2d20d7996761f160102d6eba8f55d468bc32b5ae0826962f08c19f06e10e
zed131cdf5fe757062ec28854087510f867d8cebbeaa21bcd972ff33f7e48f0af806d0360755294
z6c3a766e374a870914f3665938d8d6a3447a9315c55ddc223be42cda8468d73bd7a36bcd304c2d
z925dd2ad96d3b88caea90a7246091b336e3e24b271cbbdfb37111ddd827a4ce1cc751ec0221128
z96db15d47952d6c33ba2c16c374e5a4a33b925642987fa7906a0e078f690e97a2a547cdc5c8f13
zd404d1ec7984dab0310f86a9f13d20fa711730a605f835eee3a6f4da3abba57ce47fd9e27a0a04
z271ee05e544917d2324994adfa308abc7eb9b97f678675c86d913a3fd0c515595c6526e028a14a
zce3676d7ef5dacf50428a502ef78887ef4d5a6a83c4588932fa7917e4a46d52bb35c73b1496e18
z1a0a3642c4a84fa723bbe500d3dbf8064609dd5998bd76097eed02bdaccfb2f179d26fffb400b2
z225810e7cb863ab53a04db3645ddb09c3016bcefad1f3c5b07d3eec6c66976ee26f7f333c89226
z2c9c5a718bcca4ebd7808f4ed95af40c3f923b01448974ee6522c34ecca384fbd1b2f57382dc99
zfca71c9a7a2f752b44666a688ba0db23c1187d8264d11dad079f15fa514b0ba3e0cdff3c750c01
z040bcd61e7e46dac59ff32043160a7e3673e3c0de3650758daca7b712f1cdf8e63cfc2fd40f32a
z1b2f22fd543d278cc351a4fe34bf963a3cc310776122d9b8906220614aa1f40a03c4cfbd2bfdf0
z5710a611772ad9135321b644bf51efa68f090b8caca1909a00145a45616ebbc8b5a12cfe9799d7
zcf212f781964dc1bc82badcae60fd1adc45dd8575d30295553f524f2a4631f4e1b17460a39ccc6
zf0c2ee1b34e8419bde5cf54a354d3bd619ea4cb963ca325967f75e871991becc7e18a7fc61534b
z648ab7bc2933d738200cd371c4d7054b7e5bfe50c41ef73eaa9951497ea1299933796ce38d63c1
z481aca614c5e0e78e2dc8872cf9731a208b0a0b39d7ae1dddb18624530e3731cccd71725277d30
z4946a56191d4f07dbe6ed971f5d8fee0256b875ea1a6a4cf5b9e0e6517ed4f847b4bdaeb3a1000
z5741c999fe7349a871d74bc24c909f0c47a68265df4795d1dc0cee58cd7500f0d4d7455b4cf800
z771cf2467405b06e0210b9018c4af6658d55df1962d0391753069a57916cede38b7d087b280d65
z5ead5fbf97cb0ed7b686b7da49ad3930132c758709d93ad3fb234bda7c91703edaa79d43493e46
zf445bbe953208c05080be4cf5d793a2eae116636151452796a8bb13ce1ecc686d76be5f78accd5
zf92969f48c050f7d9917fc7386d833e63c13c4d7ff7333c93011d5d14ed3ba54102c8dbd6b8c72
z76e4b994f8268af13f2d93547975493a758245deee1d62ff9f2cb45e88f70fe17b77370df25674
z151305159955ea701a907c735b3dc64cea0d0dda73305774ee1b2416e065e07503c937b3678a52
zff2445ff266b6b1ba61928d47b16870cc3260979237cf2cf1344616fb2afd742e0089d6d2ba90e
ze1b9b9e1634f81e808103da42c70dc9f1500a0cebc755f90c5d9d89704d66c1c5d5b3870478b94
zb1b06514f6c806966935845a3aceb174ff466986a27b940e55b00603f17f4b5041c6ed9fe87c50
z789c928ef232f586ec560583174930302dade2fd0ed7d9301e67e9169a26456e125f18380f1178
z600a3eebdd230b96630867ce840441b3a8ca1793fe0cb56793819bbed4919ed0c8617da7e65fe2
zef1d59643b4e096ce000581d2554b1220730003a436475284a38334180b64ddcb6feaac2dd5e09
zf6b5089d32820ffedaa62973b13bb519e4b435fb0cd46c0768404e2b8373cbaf29652cb4b34a4e
z2d4e48dfd4e00e98b89d14b5eb376ddbaad85e42d08f6208afb3d0f3855d2c21ef774dd7450a41
zd1e0dafa94551f9d336e42daebb89208afb3e76a237e7c05afe8b77bbd26bcbd2aca55acb57a52
z2e512df3b7fda7439bb39e5bdca79dc514e0df1ece3ddf1d6871b528ad2ab01d527f259be3ed70
zf6407dbd91c809784018ce47efc6b8843d9032b4e088d781b69cbe06238e339dbd82c107413267
z56c61fa6cf9fd9302a5e6e5106280875d07a9d25870c49e9a2cb4996142be160518ba646b66d49
z5543be79185a95df5adf5b28e01f626290ca5186cd0b66d1e5153883556f20cbbdcca9bf8220b0
z6edfe44cc953b7ac3ab34e8eb448278a09a902a071e122ee5d577dad468edf59c7754a39e74a75
z24e38c7ee1610147a191fa13324d032e17fc4b1fb00030aaf663b48f61b7cb0caf029b8f9b94c2
z7f62c179120f8b9888b37767558b284d112b144681069381a89db635a95e7dd6f8cfcaf57e9660
zf3a535e603058131428abbea2054b9d76dba084da7ca4dab35bb4fc06968dc2969c196c317db72
zc394d3ecc1977f7b459ea394ba78083805d66018a87fe4d06ccad8d9a35cb7d764af47c0b44061
z91e03330251c342caeb82853e519389c1af5aa1bcbf26cbfed984011faf8326d4d1a4e387a3e5d
zeda3605357ec0b1a5811b2acbbefbab5cc373ce38db10452b5a64466c5d55c305f68603bcc25e8
z0450f17ad0d4fac92f032f5cbe357a6d93b887d6d34d2aed21ed3cff6dc56acabffc0cd5a42a51
ze9ea1775d1d83563b721edb83d95a0118f8f86fadf74043659c2dfd5f0cf8d5a7ccdc2d200af04
zb445430c7a6720ec22f935c3d864af4ecbc012473dcffcef0c415fc2269d9a35c4059614c0b312
z0ae14bfdecf53b7da573f2992a4dcf0fa027373ef067054b2bd6f0802883837817d76e07b5b2e6
z71042bec9e1cc29f60f6d0a8c7084cabf483e4a7aafca7fb47cd2ba48c2d916a4b3118a8d500a3
zea71db1232ca38b219d89b3ec7f26655694a4f0444bd5a4e3bd5a3775cd73facefdb5dc8895952
zf16d7a0815c0bdc7648d1f32ec95436a475382929f8d2e60d111081b9861b921f251708a7c9096
z9c4bfc6653ce7c0666febf29355edd940e36c98cc7c92c397e96f8f132c4b53e9b7c634d2566dd
z013096eab8956d568d3f3c82caa40dd321af12a6416f095359fe55596b8c4d623f83d8a53099ee
z186424953078b42d7244bf5a583ad9ad0ef9aada76e6599b7bb37995874f398ec864857e28dcfa
z31c62c79efd32e8ffa3e17d9b7253c1404becacf325258227606cdc0dd12f4b3c91567ddb363df
zaccb3aa1cca65cb2717a9799dd28104dfa50d2f8460d1054d364da0b639aba9dda63de2c44b58f
zbf377a2406fedb2f32cc501bcd0ea0e6568eaba01e860a1c446baf2abee8a6d880ae6be47fb865
z56fd8ea479fe476e1cee31d76a3745e406dff3ad99b9c8f14a12b6f66897c3727f5696d9b0538d
zc193c6ddeba60a299358c2d81f30fbedc7d6fe64339f68cb7185784ee4e0eace60d645a05cacee
za2b7af7cee128b0ee426ef4e684750003a636c2916c696625c7796e7f34b79757c1fd675eebd58
za472d8705920936859a63fa594073d64552a4e87e24b8d3b30d4ef5a806b81ecdce3e9ef4ef082
z81156908d3bf9ca0b2e64968b2efab1d52f5d8ab6c6c62a5c75e6b7d5badaeca9622e034cdf1c9
z19f2bfcfc680e0caabc26c1d803771566b2a6641d0ad02357374f8e1e7a97959e2028b4bce91ed
zd99fe0c0656ec862bf18fb5789306b2861f9e15d71d5aeaf291f43900ab26d015958cbe10b0a0b
zd33789c11fb528311e5b6781a7ba2c692597376b00b71b816b907e9e085957c65caf4bbc3df789
z51e465e1975a1bcb3fa915b3fa1b6853da02dc9f07e66aeb906bea13add0ae4a60e4f7fa1b02b0
z9ae8b4280f8b403e27f62c4b3168b98b790e5aa8d55509641c9552769ee746d9d8be2afc26a33a
z4325f6b06c5f114ae799479fb3fcb77193dd4ff6e05c06bef37a96fdff842bc6e5dfd5681c30ff
z79d2eb116c7ed9e56e68f86fe230ffe34ebbf636df7dba964438a017338ea790de8353158732eb
z03947c87949aeb0dd703207a833f8da4b86e2f277f9cc08ee23910cbf9cb6fe339d756529a088f
ze36f9b43fdbc15295430c63dca6c17041250910ccef76d09d9f14e17c34ec011f06bea81ec1d07
z295ee8d15e5d0117e1494d21d1103787a907b09c7e0f2a134fe0f5511f17e8055cae41721fbbfb
zb36e237f2f6f443af469ef1174cd06bf1093fda4bb2f9819383ba1a3ae0351f1f149a381c6328c
zc1f47662bfe122e48a46ac8fcd88bea99c015f74a3c35485b5e9c7ebccbe67c05292e533b47800
ze61253c5560c84ba5387b0ddb4fedcf5308de9f4565a216221316f50dccc750803c6eb4d83a7b3
zc2f4331790456d458f072a7813b94634e5dc08f5ab7bfc579781f49dcbd35530fa613d48d33d3b
z5d01e8d88ae171479f354527b91bfebb5fd511367d4e96ec2fbe6caf15c05d2ba70c6a45d5f1df
z9f205e2371ac0c59e567c9f708c81b8e8ec67c3d1dc3fa70bdd514d8967ad7c494a6eee54851d5
z4eee5ee00efc43104c8f2cff8f4c98b2f0082ea79d03e1f8a00b71a433e3c58cacd75f00c82b5d
zb27413910c45996aca828e9966c7a6123e3de82a5a3c6cce433521c81db0475e9a01b60b0ec4a5
zfb8d0b9f3fad843f9c5801ac6b72bd484287ef60e9ded7296fcc93dadc6023bde674aaa5a44f8a
z14bd4cd7ddb29566e18bf326fd24ef4ad666618c3333d7756086271040cf6e58f4b75e43a785e7
zc8010672ceffb6ec5e9d1e1492f7ede019c71c2db7d40de691fb1674eb922597650ebb88d895b9
zed15b62618e2058a91122a13737be0bde4e25a1a0288b799a68d9cb161e79054caa860cb62e3dd
zf76da033ec7a05e6b36a4a8fe2edc6d0fc65107612b9454e908616cd452c8a79d67ba5af2f54a9
z3a6e9416b3d422653ca71867e16aa556df45dbbcf89e9b29dc4978fd9a9e0c4038b20aa01f1618
z314fa80cf5419c0b1be8f54bfe689df8a4f34d30f65b49d92f7d3cb63390407472a6508ab5ff72
zcc6d5d1d8d887cffda979b411051e24a3ba9e15376e7bfa3b8477ed2baab050ff9e6ace402ed2f
z41f176c344a0b8067370d78e54ad8009c4cfa0c88f8d3044154e4c49142eca799ab8c875d9493a
za40ca584a2c960b7f8f9f7c2cbf3304016e2a0d2507a1dcdcdc73bf39e31ddf221739f6d5540b2
z9aa929bb1ea969d04cf1c8f30d3ccf3bea8a7b32a18a33d756ab7abd3b33dd27f44531b1db9bf1
z7e6602b7d59f87abd6fe710a3303f44eecc0945c68596b6dcd5320ea8c8e8d7033b047572d2e63
z29feb7113bd7f0eea533288f0935c9d30056b7ee98d891c9c81a9840f32997b326377316157961
zcd29e291e8eb908be2036f4b7bec38383d96bbf2cb648784a7b5a2c2c1609a3841768373eb11e9
z16c765721239ba9b8b3ef3e9f75fb9892532129c00d10d4414ea587113be882c9f5407ea4fa0bf
z01623c49291a7b7aedd41d4755c944f7b44e42a59e9f8f47e1630305cc0e8feb163e13746a87d3
zff27cdf79ba51998ea5a2ddb9738d5f9e3b8afe923b1105d3b7e84dc2da0a2dbac80b0a54a2db9
z6506175694fe8857d0ea27ae59527fff41d61a34756b69e4529d8c75536ca537710e1cf0ea51fe
z13a721e95fa9975a08a6eef7b0ad03c82975165b21aa9ff5db66bdcf8dcc1d237d2d06ef2ca502
z711b5c966e61d527f566e22dc1362b8d2cc76d2b2c44d362f2415eb1fb0625fdc84249f0110f83
z94f48c2a859015f8fc877b570b7e3e787e62e9a129ee456332bc541c318237b4b5fc1b4dca17f6
z7d5fc999fd93b641ad62972c0fab14e04c049762f748f2d4d391bd77c6cd2d468fb67131a028e4
z97fd979ad85b64228daa0bae3b6bacd188650933d43f1b2f0e0608fea749367b1523d3f86dcfea
z2283d75c16a9e655cc2b264c75296e2449ea4b739b8bb58437789f3bc9f4bd7e9d4cdc77bad73d
zd0acf8be1d47ee3b833d43482a570215039ee1f67c9243c80f29a3fdbeb1c0155d1620c7bcdc56
z6240e5fa14bdd1dd28745946e1e14c64ec1faa80cba76b4f31a07bdcc1d12db3be69587059db27
z419cc1d4fa105e76ed73defb5667e6f12c9a5df0871d47464b7c132fe4e3e39b80c6a33f4d8619
ze6e7eb310bacc7f9455c2be55427a849b5f16088469b345937b039ebeb5cd4a49c295c47e8f348
z576d2b522dc2ee0e591569ea4b07c0bb8bd0f6d53a435182d6a23560015e56437c55604d39916c
z6f96315e2cd53f7365d3016cd653824b63ae9fb062fdbf5f9d5c452adc668983a28011cb6d3e4f
zfe3036839ea8eea306ebd75fe448497d014d3f58e9d0caf4c6f85d656a3d432e2b55329c6f6ddf
z377c143858af45c7e90da3c1839672f0260fc51d1eca474d8e525825794d581ade2304a148a721
z801d1fe280cde3c089a77e143c67226e035ba47a39cbaeb1e53764dd7b417d064d0580a0dc2542
z0291f45facf813106f3196691d4853a7f5d4b048b82d33eef963c74da6e00a8c43c7ff839d3a33
z352b6f387300584e54a9e1f06008d9d607a6f56097aa1752abff26f3cfd424f2f6402afdba788d
z40dc2fb5a90073fc8719394596d0fe97ae59f0ffe14d5616941caff2f088d5a4c131480e6bd60b
z539594ffd7420c57251b7233a97f9aadb4c8b8431bf1a5325ae04fd73517f9a4d1a96c7a79eb8a
z4840ceda8556e173cae7b7b9ebcc48b110924b464fe9ce4c2f6fbc0a40345b51638dcf363a6155
z43d8c52b250a19b92614e7572b622cecb12b168b0d40cdfd53ec39abb5c6a39a8baf6710de2e40
z55a7329505867a57779f57d524c6eb29ceb4d1df99f68b6a30ee2799feecc9db22b5d4e1359b15
z744c11be0aac29cfc3d16268997c8f84cdff2ee6d46a6d76c16cf3d2275a0bad712bdfe4a9dde8
zded7c43c892925a20084843bf867f5b3611121dbb1b090612cf25d77534c933d69ea514e162300
z47449de6678ca414fa23b727208c24f260eb93ce35250f6ecc4f9d50b1be183b7f516f8a90df49
z14af32a450e6b6a0dcec866f0dc381f223db9c62f948ee07e66aba7c9a6b92d940c4b4232576ff
za1cc5f8df761d92fd69fa97cd7397022b57ddaf1c735be6833c4ca2cc965d803a48521e1bb9a43
z998571d3bc2f552f257c2bff68ffcd6372f5cbcc264dbc760cc7cbe39edaf591646812dd006c6a
zae8d229a0a04431b818569a1346631c597f0b998f02a3e5af53f7b5b54f9b0c8c3237c71de65ab
z537afe1418678e2229270ee8487ef9391c473696096b7fead4bacbbb9e933d9ad4a7f23d1080eb
zd3f57d800f82738604de2dd39d0183b4b8dfc274734e6b64ed7d71be1808a8ceb635bdcf8f74b9
z403a5a0674dccf21b1ba9586c98a959bd53fa7a1616dae42416b19f14f7a472eb3f382c095c04d
z81984df7940834d65e40628e5d8c2689fae57f376adcdd3fb03ecb0173ec0bbb646cb29acc20f7
z40c330274b46a94cb2c09a66a472c55db1f2ef60fde13f4f17c262a7f42f0b06f75574a8be8d8a
zce20759c8b28d1709f12f7648a32c4d0b76aeca34cc0f8d28a9e3cb1f9317ed1a9ad40da6aac0a
zab3b3e68a2fa3c3ee1c8cfd995cf83d5d2ff3eeae937ea6e39281386ab433df3a8dc7cd93d291e
zc5ea34ae4c6622de232019955c6db65d512206b96708259a2e89407dabb54acc4c6040ce62a8f4
zb201e416dd47fe3a26d59c6d2aaea04e8e7ca927320bae58b9feeed8ecff59b1bfbf85eb8c4fa5
z4b6ff7bde1a2b29703368a24a0de51d85784e86d0a04f358c1ad70a2d39b73628567c8f48e23b2
z78de9bb27cc51ea8e67e281f6790cef6dbce9274c31342232221f76015948ee19f257849ac0b4b
z6def935830bac1a8718e95bf0d948019f98b9713173393c176358b8b71435e1160e2e6829f6be5
z47b59489401b0c3336b48feb8bade338c5ee2df5cc1072a02f1b3e49a2fcf57710b0a6eb4fb380
zbffcbf08ef46553cae9a8abc8b7296c4133cf84f0b7a26b3a59afe17a44cb825bcf7bfd31704a6
z3f90610d8e50da3570d2ceca3e5cab6f250ed39e28b10b0e8e6efc5adc922ed2a9e8512da0454d
z390a3c024477188218f6582309f25572cc6c2eb41c7c0900be8225eea03eef4ab8fcc220d0def9
z2e8ccde82fb68430621ef58f8704eb5a524e04036ca6e3c540d78f5da60e14e6b5fe1f97011a84
zb4f7a3bf7cd753f74b7781e9fdfc3ed4d3cc4c6f9e67e41ed8ece73b0c52290d538ab2104db344
za2dd9d834e9035f9c06502165fe766bedfc054112561463c9e86cc4be70962872e15742f5c6a3a
z9eb0f7baf9abaadb615cccef94303a6c5250f3f8c517bbfcdebaeeae337565db1a406f3d5c6e73
zc6e4629bb08a7b92eb236376907ca7dd5fc512c5d62c521d5892ea8aaa82d99d839e5393df80b7
zfd60e537fd95206adcf0509f49165f53f9a04bded6975cd8f229d435c05f780896a6e5d0c9e94c
zb20345928ef1f7490e91fe01af6f29a2a0771ae72682be9546da74b9bae0b08407d30a2b6c5002
zffcc12e2549d537bf1ecc0cc41b9fffb40f30f389ef0a4a0e42ce53927b3842e9711968c85c6ae
z82f1e75da428d221c6c4fe5c1bd3704ef62d2b555747e0619d7c18766f895a4fc0fd4602fbeb2b
z75884dfe53abdf33d6c237a6996f086b16a20915d4b45e5364ab5f7cc8dfe7264f5c2df240e01c
zcad021a4206b20bc63edc064d9c52db691e8816a8ef01d76fe38402c79a587e5ec6841f58aa800
z586b2a78aac2810ea94fdaf5bc0ce6c7fb4e9e38a993e25dd8d92b6604ea8f587429a3f289b900
zaf8eef2e443462858b11aa70300d57d04e99878610eb3bc5b3dc4d986436f74daa1b2fd32cdedf
ze3ccf4159ec7eb9ebc395a7cac7c29615100d88080ee321d7b739ebcb4ab391cfc0747c77ce8f3
zf0a044df083a3dadb6b7e0fc2aabdf86e310139ed227214c8f8970ddd57a7fd5ab1c944c844493
z2bb8567345eac4fb739166bcda7809e127f41f7110caced15ee5134b1085acef4a3a93967b83a1
zb81b54a21efadf81c8a6bb21c0b9a6fdf9efc4ba077b4a9f82dccef49f7296d0141f70fe8af668
zb739a9d8684fb21fb85a234099051fdd69a71a4728fd4799c6b473838dfdf935f003360eaf90cc
zd195eae8aab0b235102e6ffeb477edc8ab07ae4dda9ec94411214124ee9e09403906b18a69c22c
zc2c59584a9f0df188d63adc5a4896a1fbedce48921a95d395e1ef47d36dadf47edfd62ba1fed61
zc4aa0036090edae35777701edfdf18a6eb650caa8c5591ab50df229409c1718aa6455604cd4927
z0a2784bce60f0e28f225e6cbb7c1a2781289073da66418a95a7248b77b651c405a0e0006cda4bb
zf9a4f0d44f04b2d0411b71def1dd878451493070672a823049060dc48b2a1ce512461294230d18
ze301fbd6130faf5ef6a9a3e13b7bb657df1d09db4ec93b43276bd6ce29b505989ff22b73f9eaa0
z6ef6571a5a14b5e802634b8ab5227460b83211b3841a6cd8efe4f25e5bbc31a76952dce04d3819
z2999f25e23bd3972238ba2eeb6e127fbb8ac03c6156af7ddf1ce4d048dcf4e5212c44f36aa71e7
z145ab18c95ebbac7ec696ba890b9774930d6f7fe8bc3e0a10a0bd953416d57f63bd56d780ed6cb
zda21aab44e795715aff154fbcea0118a2379ac59ce8c0432d114284a97b80166289cfad943c43a
z13bd8fbf48ef885c0fda0d74ee4ee0eec3797ddfd63af9a619317761fbb45b04b7a1b8ad0e89fe
z15a20a2bf0dbd7a2cd84958295894e74b3f3aeae238f2876b85ed259b75185d9e1dcca060f5a8d
zd5f11d7c2a3f717cf373301fe3a22a85bce28e3dfe0a0c28ba084af519bf288f099ba1efac6a68
z1d3ca2c161227dff148d74b07e4142a627350278d9848304f673fe36c066124d4387e77690b144
z33f7396f7e5ba170a5def946bc16a97a0b6b158a143e75e35deb636cbf878116afd466f09631e8
z04224aaaaeb2dd1259f0a433357ea76a97b86375bb0f66f26f5396e1ae773c24fead0abb3b663d
z1d1cfb4b560a108dab3f6a19896b95b701a1c6c6c5463677cd82373204fef14ab93c835e8fd3b8
zd7c1f510344737efda1c633e1624ff0ce46b942b2e6d299a28514d279c500c03b5be7e2bc9bf3b
za22b3537da7438cb6350cb717a2573ad35b3984cd47a8bf99de5efae00467c91188fa391a1a16a
z4029e9ed560b96cb0b542b59206379b1aff9f67e370dd162ed19ee250cc5468c70644590e6f3b8
z1faaf150fcea006e59b458bc89ce52ecbff302843adf81870bfbfccd3d3f4cd57ee64f51fa565f
zdc13f2571540d8d9420cb22eafc0ffc4701f96a4a3f5952499e07dbd3721a93b764f9936f8eee8
zee1965d126709bf53b5bf99bf0a5f115c8ad328a0df65f18d3ca123ed132e94611528c146fe674
z42fb9c9181edeccfa262e4dc5e0c74a8058d2a88831d277c489eafab1443112d8bd7849f51192e
z949819f80043ba91b7705e57da5b7d18e20cc863950a07223ae83fdb87be9ce29006b33491bfd1
z6d5e4576db393b79c23279df7244d4e8ded6a3f33aac7cbcb5c38492c7918a96ec3f669b456d88
ze2e5ab4c00032b987aa1dec0ac432d1a394ff8e0b03de511b1717a002625a0a10b5833f6a3eed1
z62a4e3e619104fc1bb26b56790fcd3638c5ed62fd8239865fff3b3b8cb927d6766159deadad7a0
z6772b2f4273d97a120e8870215e4af30b6eaeef14b384b5ed7773f0b78f68dff197d300bee6efd
z8cf1a1a8c4fb20dd0889be21472064e49942b14c0bae532eb72e0a1a5a7db6f133886ae9c74f2e
z74f2989d4c7b4a3544c8b8ffe3eeb383101955e4fb3c3a2f660c72d3e283e809845ec8a56f07b1
ze72158eae3dddde147ae89cd7060214feeca303cd85ee82d83018ede79331f60f05f3652a0cc02
z0f1c86fa562ee4e86fdcca245741f16b81448882008f0b6c3210dc0819a9ff94c8d639e7ffeb89
z4a087bb04a4d400ad077d2bb2dc5c9cd7c460bc89b4c496153a12734fc46f35ecba932de3e696a
z08ba6b9f10db61592a199bf69def6ecc05bc771a5e885bf4c8e1c1271c9d4c92e61da7d4640de3
z8da7b10c9c7f63ecf24cdd202083dc2593246ca5b2b452366392af995defcae3e6807fd26eb002
zd4568a9cebb5a1a3b21db715fcaa2e270de7d7dbc51d19b55063feddbe38a2d67e07ffe5991a50
z6e836d25a6d4843094b81f2447fe748cbb50339adff6aa3002ec7b481793939f6c1e932a991a35
zc28b6c57b2014eb6b73a911816ddf2194b839a779863c3be4bc97d52898268daa6184768568209
ze52869a608076b3bba27d4e43b20dcf85096fd0e20451b1022c9a51877095603ed00444d98e75a
z969814b9e6f63ed95603a95efe5c2bd0005c696a36d6b5e1c7d493fb9183991d874053af952003
z92d958a7e4d93a8c3b76374f73b09bacd314f058ad16df921f5a208cbec31479d7554f33daea56
z84e8d25e5748fb6c3959cef38f2276ef0c840f3f00434429591f80890b280352538b34438ee823
zb274da0c632f47cab19ed9f2f3461662db16a920edea5427eb02605c774b6c5dda20bc12e86969
z0c4011624ebcc63e9160efa9d42fc052cbcb8ad714ad57413c57b53e801570443794bb05557ad9
zaf9e359a61c8e25dd37a798ce311b41fad51dc3d13921f5a7fd7c19e18b9f5c91edaa88cbd25b0
zfee8a6fca5a8aab508ea90df3a906d22a4b3cf738742aeb41a293b0abcecf107151a60003084cf
zf549b5e40508e7b2c0887973bebf08442bfd7f95b943622e09a465abdffd7d2e9b43c94e3ade75
z4bf3a885db6d95adb50086edf782a9565c22fe7687f5ae569dbc589d22030a1ff96f0ba0b98092
za57a89ca2b84f32fd80a6e151f79363e8104798ffea11b1095a599164d20ad900c73d5d655f28c
z66f13c36eb0786126fd3177e99106ee38ba54e254873b53ae757b40ef273a985af0289e85e366c
z04169c4b05274c0cae061a7aec0ab5b2311e21a0ca6c10243c377e12b78e11e2831035106934b9
z404672418fd39bc9d7396747706c13f715bd85a67a0bde42f16abc13f957468b48e23912cd4b02
z96c0a0f3a2d309f6584182c429c1978d12a125606003f8fd61b7a21714b735cfc2b39a03f3585c
z527ee378aa67b66d83f327b4fdcfd0e35028f841cf31ba2f32ecfe93707567fafdeeebfdeb1b92
z9d24e4516ab1f6d72825155a880497c5ee30a83a9d9d4c3d31c7b8d2d0a5a88d9fb9f68482834c
zfb902f24de3f542f48227a8f1e895269c3b112bb98d0481481f5c3b547fcd8a4796f2722eec9df
z8b5ba3ec1cbe2517ea5a231ae25797a77d052d589a532275fcfa11d3dcdf0d28b8cbf13c6529b5
z07a8d8479751f6ed6dffd0161483cd0fe8418cc33ea08f59e5dbdd5a030895909753fe847423f7
z0b6c38de86de9989c2aaf61b10735f60bf4ce0e8da5d4b05963bd82b50f044950109bd649d030c
z1a3809a8b75c34aeb0691e479fa75fd2904106efa5769091f2552479f8697732ee24b0e0e55daf
za330a85cfc723d9e7ae75fb769caece9ce3fb46a4d85318b6d6994668ffb9ed7a3cf80f7a55cef
zc1007b76692d3db63bcd66178a70bb179dcdac8dad6e1ecf6fad3fdae451834c050501cf8cc24b
zdbd9ae29beea87606b2c631ca0935d8493edf56c2d747ba76f87d388ebc32e051f72967f86bd30
z295f6fdc32c1f201d07a71c04a6acd646ba9fb175817b1f762b2d2dc47d1c0a939436a10eb01de
z8130a4b82b539bda8f16fd0763e61ff5dc425f235ddb76a54938b66a98fadd41e896ac07a964e2
zd461587770d52a9b5063cbc674157a2190b3792b1512eb69f1ce8f8374ec4396cb3743605085d8
ze98f727303c16c0903c6622ab630348a9b15259b63abf7fc89032f7ca36e2c110873b163725a0a
z777b1deeede5651e945520a30c5d8842e734ab0d27e09e248ce260b09de077492ac18636dedd30
z3f48f2b078f01139668d2b2644d6495fe237f64c3f60150cbf72285cac9edf15daedde5b67bb45
zca0f52c93c5a0bd02116913a8f16fbfb7debea658947c17ba8cb3e11cb6a44bc00af3abc26d2fb
z9778d2515c435af7dc7166d8771affe4804f741f00662e34bbd5a67b9fd2a7bc5a925c2e9c21e2
z1dc36c2b5942b49f9d1b3ea151e64d414482abb686ae910a77a05194d2f16e8164d14b526041ef
zc50c7669bb7a2cc9b8975b6fe1c71fb18a586ab130a0dff118b2042f0aa95a2501980d378af60f
z8fd54d9f1e7ca68583dd14c0d8d069c07052f147da1731fc56f4c81b9dbbe590ea70c9f5c5b8c7
zfa0ade2957f7fa71b2c6f847ba1d85961a0f2a069f1dc80898c0895e43ce91705bbb03d644361a
z6aba876aabf2a0000a6d9992f7730495d6272584ebe08ae30af04df47c8ddab94b4d2e8279a3a2
zca117a8a11b49c563bf823dc61e00136e17695de3e760c31bc2db68ca45ea40dc68ab3d3f8b6b1
z24304eadf84b6db4b8bf48f7f06765fed44cc2b73c828bf5d2b5ec03c5f9216f36164dcd020037
z2e5c7550d9f021cbd51b64d03ad59f5d28424905dbae19a5aafd0c4b7862d52ccaa294aff50d09
za6080040233d953ad339fa89f14f439a81059ca574626960caaeea6eeb5fe1e191d20fab6f5ec7
z0b70264da58d99b73ebe3cd3c4cf3733147ebe8152e61ca5aa1c10d41501a01937b1c2a8fafefd
zca15fba47ae6df28a0b80e8bf922fdc3ec47c3e047e5261472888ec5a944fe53a0116f2e00d71e
za8aa6d2c2d64a224a992222d8389784a86cc33050f7e4de556e3d7d6cb7b80a833d81a1c6f4b19
zdee92f536afb26d2825352dceadf0995ef2f6af144e57b6fee2de11817df9651f8481c5b54fc5b
z8d531faa081bd0ec2aa94b20e0a1555a8522960d45fad15f1442e253349ee0f59b864ee6b741c9
z73e4faefea064f843625fbd3198a6cd600d38480883c190517026959d4ca2e995f876689b34d53
z2f6450230f2a6aeff27cc3321365eb91574d2ead75a66d3edc5a5e9ddde4519ca6acef16c658f0
z4e5f3e8c02987cbf1fbca956e9883e28323293526f889808c417f39c1bb0cba552b5f8b93c2e6e
z37d879f79dab86aa9c16d95bf9baec02a7895a2d796f0b7aec571fc232114671b3c4100580025e
z34e837697696364b2ec62587c60a112d9396547874b2f50f30885730fbc81766d2afe830713d49
zb27d213ff43af5a625e20f28ed9f4b33b0ea957721bd85c84019ffa34ea715dc4ae407857d2e61
z95847318c54816e9de8c004f5f2c4afc19c1d58429437da0ca0c6cb4f80e257c357d09ec327b74
zfbecba9ec94df101feb72e5d7a26dafdf0e24005ddbb7bd219dc0e61d49f074e3b96ba0444a65c
z960883296e29ac2a18efb733464b434e956cfec2f8c6e5fe81c529454860149f109c6a08c5e784
z2a95fcda504a0613a68da30067cbf0a7802107f41616c1b49cce70f453038c9509679c487e7e06
zf2691de90ac90a4e0704d163ea70119e4442bb0a9ad471eef9419c406d5373ea6df4b8ab2b4dd6
zee5dbe4186a4f7e6f95ee85c5043a138f20616b9ad3cad75e35a94184d52953dcc810216ad0576
zb1c435c94ff583e20cfe6bc6f20234dd819c00c2e98c3e55a396cc77236aec797e1ca3c5f2fd2f
zf30f40a037203312d5e1e8c2622fa364b1d901112204f4911fb39565d6d1a27205f0d7dae6b356
z2d0f76873cf2960c37722e5617a54370db9bd129fe8bf90c3249f29c0b4066b89aa6abe650acf1
zf3a767c0c207fe2dc66483ef20e852a3d6ae293c43e350f6d6fde0f0e74c7b11453469a72e901f
zec7709267009c4f2f69e318c342924afd37bc375e42bcbaa8a543f24aba7d0015eff4cd2d4dd86
z6e00b6c1439d7b538aebb3750ea4d9498b40d948573c20e4130020c2193e732e6bc77ef38375dc
z167d21ad33ad36e7c4ab20c19038eb055df8f8c1cca1fa5426bbad4f3000f9424b92eecd2b0825
z3383ef5c8086aa075ff450c160cc7d5bf11580dcbe54508381529faf05249576d762b29f9de5bb
z979899adbf0d5220ef291e798beadbdab28b81e50282fd0acbc312e4293957fce29c720b3fcf00
z56675f02f3eb262cc7c544a7c210b1497bba18fe1c25ee794c07193cbacc995cb8bfe8ff168d6a
zfc0da22c288b89fe5c790928725733951239cfbc37341497fd856f2341f25c955411ffba254e19
zebfe10d49dc4060d2b8272a85a391f22c6126efc51290f26fc5511c09f51cff7f51a745b2eae69
z8aaf70d0cb0de51816f6625a9742f7f3d9c9c0dbed86358a5a20cf9f59c51ce6d719f48d96a7f9
z22daee9deda9d6b580d115ef4c669577223900073798ec80552f8c1395cf77ced2eac181f0e653
ze3c0585f7651dbb5ed0fd68cda3d2caf01e0d43f8c50f17e36f6c1b310792bbc08864c4bf56081
z9d2e025320e7c0e09f27d690e9ebd849def11a237c90d7e3dd2191495ee178dd0481b3c0894060
zab7466f49ce2e17d7837592e26957f9f0bc704e562e5c123138c55b22c88f4691ffd29b520ebc1
zc315fb7d03790f42ad1552321a10217ba8d04b607d5f28658801c5af28fb1349935ffe065ccc96
z61d1f7228c468024574431bc3276ccf475a163e3ddb83c3e8a9c4d762c24fc8b7e95f43544252d
z2cf194401deb3690aeb519f94cfab206dbf7237a633b7c3ec684bfd40594be0035d41c4dd10323
zf6c1a854a297e83bbc84cc31d04a1ddf356b22255138ed007ba06f625c7ed21f6d364ea5ed1bd3
z4e97dbf9c0877a34e027cf2a0d844dda0e962b1326725b8585fa4b910efe826de8abc1490a18d3
z5539a8172ba639385d44098ad73952976b16ce9bcbbb003b6e43134705ae49da9590da68a47e0a
ze868c9679cc7425b0eef93be4997a5eed73b948d132127c18277e19179d33e3912196404247e16
zc12fcdc2fa093a39f242fc69ae50354c98721fe669ac4638f759ecebeb6eb0c89b113125f98b87
za1f9da5cfd65037657cc516aa6d73127cf972c510327a65269d95e26245b0bf245d52237543a1e
zc726a7dbbd500f522068749a122d62b954fb382ff97acfa0f229cfc4cd76eb6783eb4741277c41
z152712ed4149166f952384d38db2585d43707bc4684237564faff35d9b79738ca3c8cd600d004f
z76e9374619f44199d39bdf0bf45128e1a1cfe2225c42e8d0a85871cdb95d01aa5693ec6ae36e76
z8a2cd1d350675c318f80e1432c24f981ebf875236e216dc3700410c33b4ed7e80157c29b8269ad
z45d37a4aafbaefd4b862999a0473c1886f8bc463ce01ecfbb43a605df7548c1525c4e1ece0c0cd
z513169985ccc5ae2ca591f67b1dc6e837c4c6dd09432dd97a5568efce37fa1c15788579540bb57
z1c79eac29b8fdac3e939282ed65031ce2c3a581f3862b9f4b7a901703e443cb67819d55c9f1993
zf149c1cf3a502b378481ea9092dd2c40d2ddc1e244378c28493f512bb9d3516502aa6088651031
z0aba0c0100ecb769fd7687efc84c28ede440e69ff8402028fe275ec243c10b316b094786ece6eb
z23e1160b69afbd0e25777bda699c43f1a173e735e3e410127a7cd352bd33dc4d68db1669a31fb9
z3037e10399eea32742bdfd600f260debdfac3bfdbd9c22afab4a4ed8c53a7a7245da3f706bde02
z3b58afbd4de1dfe0462731e3749f0522c8554c122b559fcec72a9c6fef2ce5e90f9a5545395432
za36a64916feeb451d2db450e00179c73b827c624055252be8734ad1b89bd849a6c275781faab2d
z4e1a1146e423cefa6d78fa074e470878783ecf92a12834f4887fe62c49f05397207b633a9b77bc
z0375d9026138b0ce9f09c88ecdd8a9bca49bb9d606a2acb607c9e4d3c3b7f2b59ad9ecd0fe25c9
z43899aac2feb6e5aa0ff53780306899e109934245721390b8bf7510e46656eae7bee4f7f1a40b2
z6ff8b58e6f5cf898b09d434d0925e851071e0443c3a7f4d2f8057870450e0179970e84c071f1ac
z65e60708000b1bd5300df2905468ddc8d1a2dcd9ad5ed07fadddd29fbf7ad6271dcaa3989367da
z814d3ed2933c75516ef34f2d67d511a6e633bbc946ed3da6185cb19f8c969e90e63ba92e95fc7b
zeac8ac38a6eeae3803812f6e3c5a0fd4d6c9667a8d59cee20a31e8527643fff93f40dd5277975b
z4d49278b301cb40de474a13dbd054a8e6e67c66b501c7d6e0fb00493710a7f6ef9cc10d7e676aa
z6e44b9c7f6422784be29ea4ab19822060770223ece0b5ec0b5d71b9dbd2e6cc96703c74688979f
ze7ee849d4f7db8d48d2939b89b96725ea1497841d85cc5426062c8ee94551aaff8a6c703b5b7ea
z3570e648634ba7f5700d1de7231bf380895b259e100744972d81ef039901f0edfba31ff1473282
z8804b42235defcf0ebf1314ba75d69acb5ef321d598bf3c57cd6aa23722eb0fdb009d093c3bf51
z456818eb7a7dc6ddda4d22ba1ecafa5f48f552b9690ed7c8768a36f35529a1f80be50db32d577f
z2017c0a415ec3d6a4128952c0afb78dfddf5b7b7059305d461a8a4863e28a84c7db91838326e38
za09ec16c2245339de9bcbffe40d4c5725b2069b797a77eda1359545801703d5425f27320f59b29
z8a7992485127cbe1977a491ed27b059c8d21f29e75003285dd561f84df2d0e76a38a0bea729e4e
z37d6da0ed99fcc415df8d81dcc2fac36a30980f6a287acbab9fefbaa94cf06510a3cce8cc7aba4
z4309ad6f078d376ffefd5710fc24e5b7241b5845882b616ac294c26effa8050a7407fb58b5c138
z6fde4ab5cde4a93eb448f72a1875857b0de1fcfa0a119f3be102e730f84ccc167afa350ebf1427
z4b7b1817e7b1558cb65524db0b4cb6f6a803968d4b895dc52d92dbb8022fec0527daac39dc6418
z6b4c676a2aa943350176d44055afe93cbb35165404be2e76e4b83ee004d4aca53f04a060c3881d
z65eace854738df52d9be9fb1bc6c2bdcbc006f80495067e2f2428bb08417150e08cdc6bd877aa2
z81087d7fd5f86c92867f5ead5cd547dee00e39dfcda18bfe5850ab5e9c76e47af4d2b4fd7e7a50
z6f2928bcda5fead29a9f80b6540d723a797617d7973d5a0b1466e3398e46cb561e459c2c47bfa9
z9b38578eb4fa780756442f092eecda56e3a06bd46c146bcdedac504c47ad3f4a64726ecdf15228
z631461dd5e6b846974191147c68beb5946cac42923de77a4ab3c65b9d500aa4cdbfb29097d540e
z82e3d02f1741223195f6e7bfb533f2522d7b0c922f4afb92880e5149ca5e5d3b1d0fa604cf5505
zbacab586ad43ca076b5d5e5275f6a4cc5a0859f79271739d0cc5cb051d402d6b5c8761507d8655
z914868c6dc1045053d5afef4dee9c62dfe720ab06e02e44e20e0c61020a5462bf32fd63a8cc64d
z4f07a98161c54820b4b15f41a091fa8dcbf30185c6177a45bc1cd21d8257a2c21e16d698dfe523
z4e0a08b6d91aebdf314af215a5b27dbaa8a2cc78226720e245675d9682237156d48f88ff0ed401
z05932b4d4ea861ced589e44cfa8be9ef517f3e53351bc3dfd2535b19ae7519b1bc525c73768420
z7c6084722c73691889eb0f9f80b1a0b47a26f7ab045e71cf1b9ab992be4287579fdbc5f2241e53
z91bfd05caaba7048b08762e82403ea2b9401dc4ff7b4e10c29f70fa2162e9e47e76eb76901acee
z85bf1e9df850e8d951c058b5fd2ffe07ddeb423146709e40eff322d320bda62b7e4c86f09c8bd3
z8a13e2467fd5e8c95f6ad0b6920b138890b3abc8f0166e6c5b0fa166037d0fc70322345875a33a
zea6b5ebe4230256373714fc7a7e97473c9e4a2ff8d9ea959bd07070ff696c454927dc05a846bb5
zdc13c579d75ad24be4fffc89137c9ae6ebe4235e2e3cb420eb533405a3b0bf7260f36b882d1133
z507adbdcfae5d917c187d45a717f20244b598c8f43a588f08b16955130c7784b230739e1108b96
z1d9f92ff881685885df9df5f87d0e8787fa8239936c28289a613c724399c00ecb53c9f345dd687
za7db0f5582559e5d9932896aa06dc817c0ec19d00b1503e3501732dd01d3e5e3307efde24cd1d1
ze77acf2d00f7bf0a5b70ba5fd9891d34542ca610d7d8f951b2fb2a432fdfe529b67b007640355c
zbea1742a00cc4f9dd69cdca37a168554ca40bd199ac4f1543c1c0c1a41fd7e8abe94e7177c56b3
z87d8e493216628b0252994ca9504e69d57558ac7c04b1582cd74a8ff05b3f56451b5a053bc7730
z58c6dad7c1d8fcb25bc83a3f96bbf4768ec6f4edbb7cca2004333b10a65e634b7daee3a8a59522
zb6340ec13c11ec276d8e7d13ad56612c3b1ebc97d4f66e64a7d8a7d929bda4cea40cda3ddae967
z6172ac2cdd11dca77bf698f746ca8bedffbac415749acca8b01d75f7eace43c275a19e8bae0e7d
z18899283bce39cc7b36829e4b950ad918cdb5e569f9b9ea50534ddae3b0400c394f57e19d868dd
zecc6eec21e26589a5e74e08ae97d033cde4de93ac088d8e2ab9d2215e5c9479f20a8dee5c71be2
z4f49b48064c7cca7b7cadcbbe4da26cdc63b67a743bcbf5fb64482e1047bf90b9998816a5d41ad
zac7510c21dc1de87faae72607e13b9b0c85f2fd6a240d9cb7a8dcf561d6c2d2978aafb225da345
z9f8791fa8e1b24739faf1c05df37f17f30bb9d6c687a7083c47ca6e6e8548552e4d83d2422459e
z78fbee6d907259f16d4c97c48d6bf567f46ccff4a0ec046e3289d2f8bce2355761991b2721a68f
z232809ea708ec86c68a0a635d137aa9de90f698b5eed758b87afa3207910424e9fbfaa9369a645
z3bbbafed15558ef60216ba5c9ef8a7a1dc5a8f33d2145d19a31493255ee7adb330e631344436e2
ze75b3d334ee2ce9fd817a8fd00d3d3e82bd0fd6236f7f1b1b5d6095e89f13125b720d19b370159
z8706a8511f03e714c49ab414fddad945e0e73244740443ab7394615e4e11ed998da3f998d3404a
z5cbabfac3d4a4ab1ae5e104b34705c9227038095cbef071fd9b165ebafe579bac16c4fc9f8257a
z4685e2c78799c15c4cb8fed3383792cd21193e584f7a9edc9a31f2082a759a4c5e8cec92fa94a4
z43dadd63f57e5cc9d74385c155f4d30e0d95c8b0572801beddfee682da8a8dbbfc39994630ec6a
ze3cdf9e6b7092e8562c5885644ffb0c0db86a93fbcd000849e58a94ec9febb503718081ed686dd
z689383a6b6ad636fb81f0d3c793065b14f99439f25df52c9f6ed59ad55930336ece2db50c65986
z8f73e035026abbdf0edbae17c2b39fa24a8031c8326fbbb918db6b91da60f38673169dbe52238f
z13e822458f615c501acbd1390236a5451b1e6ba40211df9c427a81fb11a4a55b5f9c45187c0d20
z052d867100220dc365c31e45cb023eab215bda6a3e6ce9c3f4899c7ec5b1eae5f4618730af2d7c
zc2e5fc6c62f0b500bde1a411a90c8c04dea137eb78861c175ee05c7536da3e2cdfd9e4cb795519
zb3d3ad99a8aeb44366bda3c083c1780e39bb14684c8181662ab86d7c56bc38535b632928459935
z4f533fdade3e79bae0434e92d0e5a58dd563d5c51d54b1b7d7d8e7bfd851188db7069c4ca8421b
z97614493b65a61cb2b88dd8d15a211fb7bc9709fab429a7cae460be1f8a096c67a3d44b2c453c6
z0890641a95a0ec4e906848c2cbf6f2b03bd0134c07c6226c191cd52594a25731a583b006d0bb79
z2d1c0524ad520eee4f60d0735a1916f68b540520b3d5161f6f6bc917d6ee4e2bc9c9e68f8143bf
zda0318faf49ba5756a47e7757b01076fab6a1a9a2ec92e781eb18f7dc9be9d1c186ba67cc069a8
z60a7cabd2358ddc0520b7b4040795185e860d95ca784f56fd1f23f037dc3a270ceda7631351ad1
za32e26ba6c00bfa2af3d4fcfeb9aa5d8836c8944ed680885e6052b6202779b2fd0a8ea759de08a
z7f35ef456c681f411dfe40882232667f32c2c6827cd497a979de778790b2437ab04f6435bde5f3
z651e0a670e4bd965cdc40f0c652a3ea139225fcef262228e879f71c0b61011ff3b00e5fb3341e6
z46f30d3de9b62dd029c1d92b7fd4a4cfeb3165c74df3c6c7fa014abbcc25ad06039ac825960efa
zc7a1498a912f952d6854ace1cb96f25901abed3552f8036c41b9455f6f3a71e9309a23b492fd39
zc49fb07cdaa1b9b1e00d80189a4d6e2be4fd8080dd1805b6f49968f5a492c5012c885d78a16869
z4d8ace17571cbcb498fe0904356c0afeae3a0687afe2073f2fc30a5e7408f1a494a6f6ff2b9bb7
zc286d179c3002019fd5175611dfa6c3742dd47cb467b35889476be060d3da4b5252d26865e6063
zadfcd2f1cdf83b439fedd632cb7adfc3bfaf9589100861043ce8814663654705fa1f712d9446b1
zd5014934c21a1e11527c87a71c0f34b4c4d8f851c9dbae3299611960782ba4fc123f55ae237ffd
zf2398cb6ea41f6bace26bfa31dea48e0492b151d1adbe8dd0b8d7a214e99c5dfffd8da86ac4292
zbf933892ca0057eb0d42b052fd55cf85233f52f7b481e9eacaa70301f48e0e04df0dd7a0c5ddb8
zf0338420003864f76c22a3bc2b1de9fa665efb2729a8737531b74fbee2ba1ee24686f0fe000fdb
z972819e29379cf8713fdd5624e559ec0b6729f0a44182419a2924a095a49d671bcdf9c45fdc63d
z848aa69509f4fb1aa46777c02554ac33784541f819d09c33a1e043c6b41186a144443209810455
z15df7bf6606beb832fd3876ce9dd5d4625cbd2bd337d250e62b22c6a67e3349a7c9dc48339a82d
z7a053c9186ca02d8da600aa4ea9d07fe698f4c49a118d70457e4c8dfcdd3af80c1a65bde3e55d7
z2da43b88fc00a4251bd827c9eae656c7325336979df86094f83dfade08e25a290c305e8a428a36
z669e4953ba967f980178204a4727962dad5ab2afcae69415c575eace3333c539396a949118b5e5
z0de88a6e24867f350145f5c19ad1e2f4be24e3a4e653999093098d2ed4b5942e73e01e1af19a36
z4ce8baa43bde7290526176475cc2e84b2fc497efa0c5c28ddb71f21ec3cf616e0562077a8c9895
zfb9571f97d8a8c96a735268900ba22971988b3b54f27ec06a065bf20566b8ba5a0ce26c720ec48
z34198f1eaa5770c215d1d649cebbe35831bc807049913e283f9df50149d56b170473daaab6f08e
ze843f6b1355e4e9eb939725f4b1058c412272359f60c26b6b2a076960bc7923b54104811fcf4fd
z69f3888659146edad472c9fe949418080a8975b4a0f0eae9042c5a76c53c23715ed84571bf4aa3
z6c920d1ab5976dd5f754ca8983a8fdc98d9ac2ad454f3ad593a43d4ba32a94ff4edb821f0e3dff
z577bbe15cc972c29d1af7d1d4fc0333cd10831a300a43540e30679b5cb455bca445b2c6e96d522
z99626328f4256b4071d10a30aa99cd6dd1282ce1718a90f76ffdbac03562c6a11c0c623fa5051e
z1477740eba36173834338ae29b15ae61b677f3c1efc9c8e694ce288db51bfa3bb127ac527ad594
z794fb89328a2debf5aa98b66ef12af1aafdedffffae0bc47855cc51dadff29dd0fe1f69becb822
z324c3fa6842983feea82467c0cb8cf26a05267821606c2d0f5e6e965943aa762dd30f020286ad9
zdb740d9c8f8d5c03c15d92ad7e96955856be900a99b5ec752451303c93987e668ef53b1d1561f5
zd3d98194c5b2fcd7d8f698dc82fa050a9ebafa0bd8336e91113fc2e1d6c70caf129daa2aad0701
z4304d8cfa22f4d35285c9db8bc23ab02f426b4d5e28e28ddcc9a8f33fc4dc27116bac15f4e1f07
zf475316782c11df056414d8f3424e5aae44fbda7c53d10c1a05508e26280611082f4c427d2b992
zcf4da7da2e30bcf757a25d734e9b80715b4dfd564c5699da1826fff2d613200cec8be4520e0791
z24726a5e612095ac6654ff8514ab8c62620894a110ab5c9bbf7250dab045d8f81b4584bd64c8c0
zdbd03bd9518fb14e3993ea644c9eb4180105222b91bfe16f48da96e096ad4b4cbc7774ff18a881
zaa62c04883dc27aca2fc67011b8f7b79d3710825c3c1486b42ccc5d25b21621001e18a37bb5212
zc4eb1817919f2f642df49533010fa2471ac178ecda053e84f813d260b3dd3047f5b12ec11ecdcc
ze5a77b78ca9a8040de580ae8332e1f6aa17364b6a7ca9efa8c978c4301712ad281ac234cb7c5a4
ze508334c9e06048f47c60508128a787e2a5cc73e863a83e536969489fa509c0910dd11837ac2cc
z1ef4f48333874365f6fddfff1476ecd4fbb2f83d969ac028cbecef27c11aac6a30d66a09879532
za7281b70c9bd18c000fd6a53bc7e2ef7f7762d32036406400a876837677833c90c5e0921a84980
z7f99640b32aafa3d4568875eefbd6605cc015c2fb43a708debd5a9bcaa5d68ae9d560e61a79ffd
z97028a41d2ebf2c5c16cbf1f0a974ea38420b91826a671a371376b7dee74fd15ce7f446428d850
z9b6681345fb28f8ae47a1cc5e61e3896caf60aa19c7904164b1f833fc19060e890c9a4eb9ef2df
z6831c61c27586131c1c3dafaf36fb34b1d1c50447a601d4eb49d02f4cfdd8241960feda3847cc4
z0d41cac1c68fdb67c053737143c5a793d48ac6576c1c54c8225ccb9529ee83d8e0ed211345116d
z984076eae0c6d49ffe5d3359764d729a84863fa2b772637bd9349ce381068e06746d466c4d13de
zbf7756840c7b10fdbfb16c2168d9469955eddc3c62d2352be42c6b834bb7a4f9bae995bfda6a9e
z340d70da2ea0098a4095f31eff82c8481ada4602c8ba64aad160571d6956e71e098ff889c5b71f
zcfcf38a9853562e6df2791cd43ded7da468f5787d130a25779d7424c8bdb48d70ef41b54f7028b
z8aa18a45f976fb844e7379f61684090a7b28f83f26ddd8b0f71bef2bfd2662fed10219f5cdc966
z3426a155cafc79fe6f1d299856d88129b2d8817905aef2bfdbc0063a75ddc6d73c67e5e24de03e
zbc0da8d0c70a714c8995e775a7b12ab8e52ec5b61bb72524c23ea412dd108cc3f1c6c0eabf5dff
z8fac59315a8348cac967fdf360aa84b7bb13b0565066752667faacf827228d459f21b1d7db5e6c
z9c3388b95429ea5634e13b72b16fd2ebd9bb1282bc5ab688e84914021f05745fe6ba6a2b4406c0
z418af6ed88625fdd3a6e37e2893c846ab29985cac84fe683e2d066fc65558d8505365fe66dc380
zc7cabc549e7a9a617151ea435cca166ce4bdf357bcdd4740da9c1529afa8a8991fa2d4f74ed460
z09b480579b7bd4c36af14889ad0be52df8aee4019bed1403af0d04801a3a82a416380b83403e3a
z146835e8d6a577c9642b7454eb3d796a3a685a21bb173c81dff37eb7920c9c3d9271cf7f876bae
z51922acfc4e40ecb431466f51e14dba8c3d8909f4f51f3c775e60e626e0ed891d87f0d7286db47
za9e7b2c3a33fc9147d76c77a1aeb6e29ad0fa609aae6ee67910ac014bd915b8546605a886e3d4c
zb11903fa070ca4f304d8f8cd9be88554edd5daa9a0fed3c8cc66d811acb8b18755f5b113f87076
zb75350e5002f898f5a0b8726fd859ab60855832f91a239302a9bce208b950451af29ec4cb381dc
zf0e8626259330a9d01feab4d185be4496f6a70b6b6c02a8a6e168c84d2ccbf7c7882a75f0a4392
z288a6430ecb4f7e840b1db9953a3f318e620eb376f8f9809bec843a769abf6f32a924db5e9764a
z626e58d0a302ef219f20389f2dc09dd7149a578be29907d59abc91788bc895e6d45ed42fc89fd0
z6b6448dd95c70e724968a8fdd0e3981fe3c47adad76fd6025caa3df081e0903a0e8fc0d3ca7a8c
z48187c3d7282e671073179cf2d41171464c6bf036f31250651986e47e9e4cb8452aa83a501ee83
z3bdd7c327fbdece572270d6c8f545b3b4244fc9b814e43b29d0e11414a3a4295980eb1cd3980f5
z83ac7e88c8b157eb1177ded502c0cc993c37ac97907bde5d43a313c3032d1b02d788a848620229
z3ab50dd07d8b77c087f57bbd11345779e98b14b53b5be66067aba228876601840a3d22581230e5
zb3d499860fd5328cf50a66a4fb9e1e5e54b5b0a1c49af532aeb783577d68b160181113653e84fc
z872ceebbe2d1d0e2e04f3c714a8a2988ef2c6152b0d27c1d17b54d757e73febc58ff36290cd2e2
zf1b9fe8d21607eabf2b5474395df06ec8cfc0176a6d2f80b691f83ec3bbe5cb2d00a1e65dca0e8
z8f99e1e83aa82ab02f48a9438b39fb5cde881b9cd432e4a5254fe42d70a0708f79a98ead62ca7f
z87e0d7db26bb0744706c0ac5ab6fd51eb0639816eb22efaf58d9c98c1ea8a6a3b02bb48b11182e
za11547bb645e01732a462a12e59e572368302c37da59b1a05a1eb77e76b2125386efc8b8a97963
zcb7eecff87052db460e6af8ff3c26d056a799bb9d8d590bc0e8cc364140698ff26e74869081323
z12c16c67af9db15f7c8905f1e4a2ee4e4884f73e51cb9121aeb0ec6737bbae343707da1bca6bd1
z85126fe052ab872d88b4bad9cbdde23313d3643af282c4d23d3f4a4cd0a1e82b74a8f547053f61
zab79b3d38647669e6f71b923618df02c55834e4f2611b5a4282a4ddf7ab0804250639a77ca40b4
za92e3019a1659593a92171bc61d0505584b2c4498f717ac420d4bf2695e591427537d55acac2b0
z7dea1839c314139c6bde2940f628fddbb2d1738b0ffc1ce8fe54b849db2fbaedf4fda82978b67f
z70ae677fef3cf782de907fb9116e3818b8d52ea82b12b4ac14a8bd15a10afe06719162180ef945
zc3d02414a05e3a0c66d38ddd4db10b77c1a6ffbd155a21cbae7bfde08633d015fdc3b1f4e7ab64
z9b7c8a5405c0e1a813e5a65132beb2e2fb58c0e721d19e874b825a135008c89e7730dad6649742
z8b6ad83e7f8b959e0ccfb0d1104d26b8a0602c4d7bfa3644807918fcbbb2f611a2f8316df74011
zb80d37f06f5b17573e909516cfc12a10dc0790fd0b1b1f795ae9d6414b479b4018ea5af2c87075
zddac0a1d67610c64b9853dc000ec7b3daee96aade00e1d49742eb0326145ea50cd03e9e9eb2ee0
z26d6463af2fb23c4f90d519cac4f1dc3077497d9614241102dfb01f90ad82f8cac63e568b715e3
z18ffe78cffeb822d13c211b604bbaff782864ba938eef9dc2ec37a3acdf71d0c5aafbb0e1f8c91
ze6da6cfc6e3a2f8b307b45d983c7b7df833bed3db0e791cd17ae7455251f6147773b0711b4866b
zb96d45d6e7e2d5892c58c655c6525aa5b56c8b2aaf747097ba080170aa58a015bd5f30ea18d779
ze3916330bca9a6e7857dc5cac9ed379a8a345280c2760297301925d3bec95e5c6e7ed4287ce7e8
z0edd6d580932b604e8509b533559d7f85d72e8547b7d0598a77299a57c428dfe190e1ec840fcbf
z04e66f7628f9b866aef846d27cd258c5fd831cc27a895014b44b9636e22da673324f55a0f4461a
zb4b123b6a598340fc10b16d8d9565f5801bbf410a52df4d03563edc5c1370568da87f5dc1e8e06
z27f48b243be415af062abe9a7da5f0de6867bb49b43f6a5bf0151c8bb07770abed140f07272056
z168e8d64fae51f7eb2b36f7415cef3528f637d7f89a4e31a72f097de0a558a88dd136069b133a7
z28873d90c3ba5b8ef1a9f5312e47fd111edc69f6b2d7e999591bd85a2d76fcc5bbdcad4b5dd1bb
zee6c6c4fbcf13c5e0371dea039a707390c9842a4932f4e38e134a12dbb410846e6f1cb41ce73e9
z9c92c95ebb1eebe46aa8584d425c0d35072e798b96ef56891553f61f9cbc895f43ad0947b6645a
z47199e43a3094a6587a8a0f7e944ed3ca12f3397453ea6167a955a4a02feee90723e59e3571604
ze0da42cee133b57da963d376f1fcb203e39aa7fa179151b5cb799f42085f2255f9a050749b88e4
zc62151c9c5f6246ca00112f786ee11efde536e761a2740071fe1ace42aabd33a63e97701be6c86
z0686ab71f29283f315b655674349a48406afc060a5b184fc89063bbae4df73816a6d5f4413279b
z43f7fcbfbd115a28c4781f3d053d6f63f80fe81ad7849d5d23aff4206ccf6a3f5edfb37d81395a
z20a6053d8a81dc70be6352cd93017098bc69af261182af597cec9558703d0845d331f383ece819
ze40bd2135e29834b14dea205a5ba2b5ca1f9405c48ac0b01041432382e7f6319f6aba089a384cb
z734c84a9549486c92b5e23e2e4aff0798be5804cbc139a871cfa5ea454c7509e6bd6b3be9295a6
z9c5c252237d03cdcdb7ba5783e9c1d26bda569a176318bd3847f7a0fefdfd1c106df72413c5575
zf0512b5b554fc4ed41c3ebb038f474200bb423bf169d004439e4d9e981ad236f0c6ba8e748e7b2
z8fea5b74c52fb367dd1b766e9f358a6ed675e8a83b273483c2e45bb0a7aca7b0ba22a4ca16ea19
z557d4b9b953139f86deb1a39ddc95145e3c0632e2f32bea069b5db4e4592480f1c95ea50754fcd
z5b7213a2b37c1d0f8016b0bd588c7e4a12f648c45429f29a7947ac08cdc27228dbca12c2fe3a13
za05cf936edec61881b63681312c7526cf33351d57610c69c85d8b060176f0214383624f7e471df
z44f394eae1ec6f97f814cc7860b549aa93f455883a8e216d8613b5521d2cb4119fd58da7816f11
zf09b739e8f302814096b64414b4a3066cdae707495197a72571c251a84033e78a4ae924555d2ac
z54bb4a5baabb79bb400f7c06a16903e8865e305bc69d7bfaceb04fac1679346c22735fe556fc92
ze08af3107049bcaa2c433718218f4a598824fafc3903e780021ade759e2e7271ccac3c1014eeae
zb93973048d3fc353ca5d5030f3d21786fba93abcd021defff1dca735e9027fc24d31f7ccb830ec
z653b4b671ab3e40ed7249d6f7bf6a07e6c69f76de763b956e52eb61c2d20fe73ee5717cbc3e0e6
za6d819da8d23c9674b2f7805296a04b3e723ce927debf30517b695107b9251c6ccd45b91bae84c
z9137b0d34883a9dd506c94b831dce8ef7c4fd75189d3aada0b35c10a1807e31e2968da2e43d0f5
z81d27b0a09667b0477e2ed2c05797a398f3f7a0a4da00faff68c028d6b0350f7f0c1e65324cbb1
z28fe98f71f2901d63808e52e0c7f7bbc6479c3e408a13c442d99032fe3afb35683db621e58e188
z8c4ed40479815719712a23b079d1af0ba327b691250dd776327450d3a0b3dbd692e6f11827e6cd
zbd2655abbb859194970e22d8aa5e69e05030c7d975f808220e1087471731f3fa1fe71a1336e32f
z1db82b2b0ba83f531bb31be26405e8d92cd0b87194cf25c17b1b5f93f3cc0e996032ac4f04ef76
zf2010428cb4d35cf7f46a5639b02f8f3622fc568f30ca4ce54673615e42cee7738abe521d8efd5
zaf243f27c75cac8ba1ad1c03e8e86e3ffc438a6e54dfc9de0e875b93c21d01f56e70eb111554a5
z227997b3a27ac27ce9bcac7d0b20b726c138ca9d06603c448239cf9c7831ca40eea00848c2ba78
zffa9a8593de25afa3a9727a7007c3e08405c4e2caa342bba5a3bcd69542daa45e6dbc004e5538f
z24c1d39606ee9d5839cdb11b70f419d51bc82ebbc05fe82df322b8a5c3daedd1b60864472c699a
z6c3e5db013a9f1d728c722d2886fb825b0cb2856671af0b559775be2dbb77741064eba86075e6a
z11a307a403ff1d50245f92e9ec71c8f527bcdddcc2c2bf562826b87b6923d9254a9fddb222c069
z9dbc8acc9ff5cfbbd3e49c2bdf53eba680020078fdf1e25a5cf33899e5e199a69c1a072f796cee
z01cadcb5cd0f9e47da58fc3dabb9a512059a79b1589b260052f3a454cb737f962bcd64a99b512a
ze29c55e53e0da461a183b64dfffa3e28ace48fcccd2df9975dca67a0121efd7d0a75b961172548
zf2b0df03d5513ecb1fa64463aa81b22c9b18cf4303ac0edeb72730a1383a03bedd2e46be5f094b
z5afc888f8e457b79b8a461d19a258281c1d788e23fe52be56f99bda031612c8135a53d901a5c09
ze61b2249898c02844201d77673ddfd46356f79f337f5235b14c003b704692a0cf3daf9cba0fd36
z9b4829fb62526f52d426c737c779690daa0d427110ef9704291d937e3c594a77dd05af0e645382
zb2a2bb602e35ec837ed66450b01b8052a6325e317eaae81c7edaf26c101103c55fcfe9c9be0d06
zccbdfbfb09130ea34e6f663577cc780313890af2862d35a0f2129ae02b4cfd2b35466635318791
za4726e4a4dc6da8a91c144ebf124d41a1be2dd4ab3c3faf774e3f4a08637dffcd3d7b14145e294
zbb4f09469f80f3bd9e8e2b08dba0b230c93e1d698f7c71fa872e7940fee314f3fd97fc0cc606b7
z71d9a70b09087821e6326966b20764b20ecc238d2bc86c423f22c2728730a1fcd6f872f2fcf64a
z7459b799286c28c41a35b455b6babbf03dd9cc3f1d6c023ae3234dab66cec0e56575c0c116330c
zb5facd2e730d87ec34a85f2a3615b2b060d267f5d31ce022b4bd1f9b6be3fd0b9f973ddbacc62d
z0b3f9d01b2381f7827cfebdb4dd07ee0867df8f0d925c1b79373f6723b56dbf802c2c0f3b95aed
z2cee1efd13f8c4cc0ae44c0771665b04c1dc95bd5482b0629860bbbd48c2c98f7df9d5458320ca
z2d32cdefd0e3c5cdaab64bef2ebdd0ce76f5ca4a024ac46a6f759dac5b38c7e42f3ebd4dd74009
z33355d25d26ec8ede82e49ff108f495b0d277db05b3365c090d92a2b64bcd48d822604537c00fe
z29e28737f7a335b0f62247c013b4d86b9c565a4019591736db9be4f77c78a02d0cb7d866b51dd9
z9e7956ca3894ca723e4327581cb0098212d0f6204065f90b3c132bbe524383bb30e17ea21c5b8c
z8dea7843281c58934963ec3fe03d31cec0f59c0c3af9080c595f9de4778619ed789a1acdbfa99c
z0afcc5a6a12704d4dc2aae3e9607b4708f113cb5291da252fe4a82f6ba110339579107dfbaf30f
zdabfbaf98e8d5c604fb151e0674a0ee828355fc9fcc29e9718b2c85a61fdc2f81fe46c3c0adf5a
z68a4a9cad08eed3070092f4eb2a162663ed8d2cc09b69b2c72cd6ad468a7752959d1af801106dd
zbeb9c050f4cf0c097aea2b62bb4dbe3ab61e81cee2aadef4618d76b1f83e014a68d09437570e15
zd71e1a14f1840143fc9a7068d2b1f491e536f668b9d5fb538fe8aa4cdeb13eb3e5e26864348867
zc36b48426b4868a5e6f0744fe1176166019989acc173e18efd7aab7d134e90b8877a6bd3c0bf8d
z758595cf143d031cdb217060def763f63a0e529c547becafa64d6ecc9acffb617f197955037194
z865a48e6531e9dbebb2a725ef8a6c6a7fe25c96f30f7a4acb14e664267057c1ec22d37234d27f8
z4ab2991a28834dd658d9156f739cebb072da0bc9f5fb551d98d2241bc70169a807d7a7a0b05146
zcc3e6c95f0f7df68a50283f2d273a357fd4d8e625d1f23be8ec1e62711a8ccfb851f2d0c2b502f
z86b8e4a96fa8017d65947261c248ca56c7c4e3a2bdb93b310f75c22959c9197a309575a28f0f65
z8771d3dd71f9d16bdec6ff1102b89ee2aa0f0425fddd1e0655e35e49dd386410f7268316e2040e
zd884b7dda5f0ad53c3626f002156afab4baa66fbfebd35c4922313634509cd6f5990e76d803f6b
z0d160539fda2ca254471cadb7ca744356171699f4e683e4c0090da3fe602c0ab15df56028407db
z5a7384f39b056fb5bea7b9e5c8033c5f5fce2185547dddeca3681d4b36a0e185f1696ad8f0d83e
zbe98d9cbfd33b686a3654ea5e8a4b112808db07e71513ba30bc10fdef60f47d6d68d36ef5691fe
zd2e9a9fb00f1100f16b97e4ba271b2c25ac2aa31a9dd2728d8dc25f136f3c2569c8201a43a07ca
z5ef90dce26d38baa08b6019ad90391cc9d49c0b863b0492bdc67c07211ce256b724ac80553f9d5
z7373c4585c9bfaa5bfa9fc3bccb764809542a978230d6a1103ad229e63de4c14b1825ec89a7715
zb16ac77205daeb4f1d74f06cee259b08113d0d8c3ecb5dce52555a4ad264c1b307e2d0ae1f3269
z4cae241497c9be89d584df12853915af3d8963826dd9915c5ab3bbee362ae770fbdfb27ed6ad71
z74dba12e7d6bea1b233c966f25d1e6d1512d9d06e93d5a7fcfaba5977343683f25152ceb17444b
za75bc02d1ef4652e3f2bfac47bfdcb5fc68394770940195286a409425253cce12af01b57dd5e57
z7d6d2e3f2c969136cafa6e5fdba38641d87e82b21af86d1ac0620e2794ddbc2aedc38e7ad69560
zeafcdac77cca975e2a5063d0ff0dd4b66541099aff914714adce2e5ff8916307b956cbe2accc6b
zaac50e5de4ecdc4e27f2137f36c68e64bcb6b31b830ffd0c98f1c50aabd0f502f556a3bb35e514
z52257c7140ef8d3e9c6d8fb8e06c7058c203741b55c5a9971b0d86f67c3010d9d697c5c0456d69
zc84312de1159ae927569eeea9dedfefaab738bb0e3c9cf5ce4bc6416a1f530a5263b6a5a85cdb3
zf25c1c5e9734bbecdd868d70846c3fda7fc59d296cff668d954b6f8b1af62b2a64f2a0a01b9ba1
zf306f868abdf06915e1c8d85b1f7876900817caa4acbe92bc752afce904f9df4ddf1e983f06dcb
zb80fd41870169c599aec3c80073a4036ec499f93cb7eccc69337fc673284b185afd9bce5f39fcf
z6ef788e8e290b26fca760322282023df7611058775d7b8c6176e4126f104a2c3395e0be248c0d2
z8ff6e8d6a3f9abd242584829a509c19668f56b1446ccdf7912126c52ee24b09680c02b652f7bbc
z7dd6061f89dc590f42777857b19871a1be342194c137eb7795a1eef93d91574d31c7a987d351b2
za93da971ad42d6f5ba11925ae51ba8bff1b79b1af109d2e98de4aac037fe389b5f55ae5bc8fbf3
zdf3bb0b907ac2fe783e2a4fcdff5a8029dd27e052238eec4d9d3cf879dd4d408a9db69d68e38bb
z16d1e57bb70548f7a81156a8ad55062cf7506e5712b0c2113039e289bee29c4b121895590e6296
z31c0b1d6ad96e23a0ef70bd7782d164a21506ed54e2d009c3989c09eae797a25ce84520a972e6b
z933007cbb6c8d3711a40585b7b78d2ee7c578b4959f45d61cedbd6a37445324e258c2571a164da
z73ca28a74351bf54161583437be6f4361072e8f98d9c347f56dc76749d2131f7b35bc7882d3b80
zd8d328f45f631e5e29b9753e0d8899f5cd7571a18615af884464f66ea893764b688761dca3ea94
z826205a04efccf3057c6ab9cb2d02da8d8b9b1fd190baf7973fffc0aeb391fe8269ad65cd5f604
z0ec76d3f88224fd192ff03a15280ae5d18a671f5e265074c15b91891773f7e3fe6fe81d3615edb
zd8de29acec9b708f274b88406a44334d621a45d6a861ba9647a46b60f346332c129f18d2593bc0
z290f1011ab8f338a18de0559312222fe84064c3a9b162a3ebd23d7092f99a12ed04c382590061d
zf064a260a34176b202bf277bb088cb6199f2d11df234d88d09b7bc8a9e0813d7470ff3d2176030
z052151e8285c70b077e2973239ce63eb76cb2ddb4bd9fb81cb936418da18def08529b1dfd3b681
z8294cf998bc2cc366ee9d97dfdf680df5e31a7ff491e0efac212b4177a8782bed3b89c6f26ee25
zea0fddb8d87d27b85d70a7e78f2588a3c3fa91a1d86ecc673240f80e0d3c2c865e90ce33f43101
z9acbebefc1818e3c22685b1841ee0c11d87d28105c9f81c8a1f510e180c235def745bf9d3b75bb
zb75aac76418285b5451ed75204855c2a7f365ea58c975bcdf5d714393520b9b6c4e1c056e1a366
ze1d2e5313166ba9ec76ec568d94495991223f366420ac07b13d32100fe577574ef98c39bc1b3d4
z849ed9aec060121832723fa8566c70a4c1e6a92966337959c319a1fdf0a679fc7764052e1e94cb
z3b3b475f9fcfd9263a78c4f16d67dadcd49c96a96ce17ceb0acca33e651a53fa90785fee36786f
z739c2ac50b74cf48948eded8713b58dc8bfdd3536357a5172d7bbc1545b4653da1a3b9377f60d2
ze853c6632e6af2617656a9bb37c9981cb4265c3cc595248835c559b5eceaee1e0f79ea66d485b6
zb07aaf136c0eb6eba13b67d7f8e5361b53b8d3a335e0a623eb9e536dfb902387c54cc563046335
z70a20d1d41dc2c2fb490d2c43d1115870f667915336d7ed2553e1e3baf90e764aa450f3c9a0360
z207d662e8e4bfcc54a58d9fab8b0fd385ab5f0e3a80936c8de417daa05d5fac07d91da2b399dad
z7ac45c721d45cbc7f987ba22a16f0c5fec3d498bc2dfa5c6c3d259c6bfa9214edb05e3901e4dad
zf88172d0dae528b398ca0c48297c3f025f02ba21fa32f926f7074fe193b72fef0cb630f65783ea
zcbd99216f3fb11ae4358fa4f9b73d5f39c12337c6c7a482ec1d59c7b5425051c00e3f882585a6e
z4978d8a913fbd04538ae4984978ccb51764f2bd1815706c429089f5e018dad7dc380610c951dd4
z95f3f50c819d2eaa1ed1d6b47996649c38d49cfd93924470bdd30e95667743d6aaee0fe423b98a
z590458434ca9cff1f730f50eabfb03b4839af66e18fe10a9408d20a1f770e72e4b46b71677cee9
z264230dd5cdb62ca137415c3b162db04628b14e19daf966fdc0f32df94ba0eeb5587ae01e4bb13
zfca0acf7923f06518a041739079aeb22c313b070ec58e1c0d174554065fc730579f0fbc4c3abe5
z1af6481254f3e31dc84a23725ca3e8cd87a651788ea18309626ea1ad2695a4da47a2c59c8f52a9
zbfa7ad539b282bd1206628588de6395e28e6accbf6c4e811c1cec687b3577f0e70b888cc3b8b40
zb959d9e62b5c421cc1074dfe5b3ec9eef8d2b5ed8b33e89471c34059f4c8cb3fe320a8f6ee1a23
z05983cc81ad939108856360227c54a8e48e865b2668bca9ea29e8c9101b33fcc35dfaf95be3477
za8ac7cb71b15528c2aaaab5ae4abfd71890bd0fa290a8b257a579d426bc444baa435ef403bc89b
z9ee88285c3d922b07b56273b1921721ce0c24b7831df8959696c06b6fa0b652eba278c1d87ad25
z5702fdeea016cfb70edace2747deea6bd4f8c9c462096cee61238ba7fd4edf8df9e8ca4fb1e1f5
za54f56cb94049b2bbd0b51738f4da1338c4730dc7fab11e07b03a666d632b664b23e6671d39f93
z672994299c714dbca894f2efeeb5d2ed1721ce75ecead93b54270e0bb62ba4b95e5366f1af6cdf
zfb0dfd9bdd5d6c4bccc62a1cf728fff8cf494fc7e4552916df2bd68a7a01d913312f7f7b88b17f
z5e0cbb7d63cd61a5c73d483358419f652a2b7dfb352fd5c25879661f7819913d56ad8b8760aeb2
z23d77bf0c78480a9c8dd6898c848c56cc9e2fcb3d6a937d489af384de609683711df404c455639
zb938e71ed78e5a4e5bc74fc0c313d67791ba6663c58777c0666e43cad16a6a5d8724be25e301db
za224145e5e9ee8b5a1bfb8d200b313bdbe5606cb7a1b9c9adb0fff866588c92049ec76b08d4d6c
zeea7ff4c8ab56c32f7d8ba7225021c743656cb0a32112250dac0024c5e2729daee6c64e292103e
z19f38815f27b96796579e80bf1e53b872d44a44721b1b12fc415be313c2107722d5d5c877f8248
z0d53dfc365cb9963f3637bff08386f73cbb74db02601aca505082aebd71317e9d9961245c7a8b1
z10dea10c82f0300e5cf155db265d622c5f485bad186bc95f2f9ec3649b1986e11886df1d821a9c
z6f5e44e3b83f48ee4a2449657c3c256a1c4fb86d460234526f99afd1967736b12c10c045acc059
zce43f99087cc2bdc78da7be14d152ad9aca80ae5321533a5bdf94c45eddbd0bfcad360a52105a2
z4a754ebc9cdcfd10880d633137fcff0892966a254179d9072af75054053164d9023c8aa65c8fd5
za637be6364606af27bac74bfb8513f4ce0a02f8b5e80dc4c803f33019982fbec7278d67de51964
z472202b51b338083ec905a21cf2e0796890ece067a1d17d4a1444208b56bc92b50572cb5c9f9c6
zc2c2200038b715fefa6b8099cf7c02f9b4044596d168b6ceba05460985ae597bc6d9061b24cb07
z6c411cfe0d329bcba8b935be6af11ee12e7200f501d71767a46a5fb6b6f0628541d4c7a5fd7fd5
zaeeaf75268aedef11eb3da6f9e0b9f81f12ba79b73e0a6061e6e20cc641ed424f0304b362963af
za701cbb344c9a9a37ae36383980f2af88e4bfa248cd3f6927b1855f618df9f98785995c237995c
za11dbec39bf599e36cd133944cf666c9ce02eca471293e32c611949febc87afc8053484aca1a18
za9f647d006a7a3409761a2d6f3522f73d66e44f684c81504c5bae894570c8fedec26266b5f94af
zed98a0c1b301c645c66ae9521370d9099ab14c3acde88cf7c9b26c49f783008d58df3d1987b479
za7d74d8db561a9770392bc350b3c8632c7eff032431f5c9e244bea2f7de5df533a0f088b0b4724
z2ca9c20748fbd787ed815079d8eb46c412d3a7b41f052f229e0bc4b47e77c01edbed6502b42bb7
z2668eae35f53a287d63405a8bf55e9be7d9c5ec6fb8be2762450f7266c56a5aeb58f7f72ca6bfe
za75629ffba2df2abad9b819de95d364bbef357f0f50b64a81ea8b2da4f2b23b8a0a8413f3316e9
z3462cb5cba418261b20d562c1619fb387472dc9acd5ee26d01008cd706eeccef71336c42342e40
z25203b32825bf2bacd2c9a3a8684f6bdc2d2bd3e2820e5c1517437d9fa1c5931fe17f9d552503c
z50e8322db0b342fc3e373eb25dd1e0254340a5b0cbbeb31984162809bb2aa1159cd97198c9b199
z171cb9c3296bf1d90f211dabbff2ee29d8541b291d794fb430e886fe7ba63830ad18e97fc502c2
z9fedfbece0231fd3555fad5e5ccc7a0cc7adf430237df6c729e1b64fbdbf63f435e9e36d5c97ce
zfe047f68f341baeb4d8b30a041a6f30f514ce858352136e1ebce9ca701f210962eefa30898e40d
zf785672c98c9c2e9734cb32e333e53475d5d4c006d24be28a60aece498882705a7edac80179ed9
z29302e9c4eab7ed0965f05483ed9ca1ddd1b78db7262089a471920537dd2b7550a5ea2de126962
z257acb3cd18676152278d8317a2b43197cbfed38184b2761ad9a64e973e7470290cd8199a89770
z84ba18491cc9401a1c5b7731c4e438b74bb3ce29ffce266a687ac927075cb248dd08b8feee05a1
zdbfc29fd71110d8a65ae4c36737cd9e62793ddb821cf897bf5128e70631efcf08a1c5170344780
z34739d60dfbb261580560c5dfaed11e8f56dd6319e2d0c6fcd2e95fc3e1fe89bef7011de525d61
z81d6c659968d371b065eb4ca5d37ef3f11e9924c991409c677a3ac42dc857d0cddf14d6fe74e4e
zdadd46ce42c4256a1ffb40a4f0a290b1940269101f238115d76ba097ce18a25a1f72baaaa6521c
z3ba9402c59983f91328949aad5973d7d9935c336a713b0853fd2e327f882ad25e63a49776e3ade
zea3ff702d691c571358f04a64ae4e06ffebec51b1eee0b3c973584202b8bee0ce46b2399798df4
za48df81b6c329f1b28bb9507a693fafca68db9d59bd42b9bfe28d37dbe90e0f24fb5138b3f931d
zbe58888bdc9d462345505e78a52a4b0bd3b91f06f84268b609c544c9af64e3438bb2e879c7e2d2
z795d572e325e7ecad2259903e1f27fb192ab33a1297aeafa487c001d04c3862d8461887d36732a
z269bc3c24469f39ad165f51b5f531b9b618e079c3f8f4fd7cc02e6c1e1a51ca29ca020b88c4544
za01f0b9b6a083d3fb34327c83e748f063fe6360bdabd61b22ab47a26e57e558a3904435c59fbf8
z5ea582142c80f8d9bace021aafeea8391e9667c527e9406ec6dbae64d4cd84f90d208ddcf93d09
zc56f4772b5fe3ef8cefb26ba4d0b9f343d5fdb5ad777dc7c5713d7f4e37521e379f4dae671c16e
zdc02fd0bedf9ef7666577124980152877be979ff1048e90696a762862c5b4684041e838eacde34
zbfffd0c993731bd3cddec8084fd203e4b1147ebfde2212c35828e3d2e2964dc741ca574676e109
ze7422b7a6c599d7b8a0881636e2e654038fe9e8b107a3e6b285378995b44e4a8b2d58ab4b671da
zc7f953f607f76af4200f92b0e03148c73688797205835541faef9cc3a42c23405d87c5f89d2742
z0d1955c04b7f988d6913cb42efa09cfa45b5da9484de02e6de6e99492923b5dc9a54020aa9796e
z4aaf7fcb5f56a0cd9ea0cc427d98c309101d041cf25f69c0646ed97c20237b4178bc6e67f7bb7c
z65c6a01491e5df6cd66847417cb18121acfb0d23a877e7e1d81197857222f9a86e6708cc3612ae
z27b58d629fe967cb20a90f3ee81359d2c687da3cf081cdc611a1aca16a029d5dba9f3a5c36b3c3
zc014b034092bec55c206f06f06c6f138853df1bd801f4475a50d829264585c8d9b4b6a37270ad7
zd6a27ef933d8dd15f27064bc9a059f303456ddd702ae254e280dfadc845abdc6e527ee01c3c1e6
z30366e6e78c6e4234b9bf0071438c59f0ce32b3b229c1ce8e446b21a5cbd49284ab88f85b3370e
z5ffce1243326bd0658ca91358814c86f208068600aa9fb588da4cbb4f5984bfb39d2abf73aff54
zd96d7aae8761d6d140483a369601c4c827fcfe8e69053d69fae67aac2ce17e3a09aec8dd12221e
z2503ad93605c3514a9687c15b4c78120360c84e851771110045fb137ee228e42bf8df9f1471111
zda6b563281cf29507e06772c311b4d488a648b90d7a1fd5089a04af8a14192d0b2c54298966deb
zca068f62bface2944365acdf4bda20246443f07c26dd6835ac608122318692aba339ce71b413ef
z684175a2119c6478fb5ffb18c4fc3d4d9195b28cc271c70004b9bf7aa6c4afb0b41fc6ef52d97d
zd4e4eb6f2c5f3cd94ef61f79e291eef464efff8621f40ef7558f2f4f2f23a0c9ae84097c291d36
z68537e05fd53a6990c7e8f31751f3c31e9b26cfe9fe1462ccc4d5de6867853a965b130706e4123
z61e23695ecd0149222e82132e22cdc2e230ba9f9b45c7a396eaafce9687020b0a04f930fbdbea6
zb5d40f5e75800939fe898d6496cad56c9290a190f4ebdacb77a97441a5c30785b5d0f63683dc7d
z54db9bff4b3b13c263bda8e20fa9435d1334b34103538ff72f90f7384e7008ad381c629b17737b
z741a66ed2924f4a9bf00ef98d2181c20bd11b35c8ae66f80d78c972627f0744c92e6bb86594e68
z8238f4f223f72beacec566f54b6a8e06d9796856f491849bc11a5282a03c8ff83f03ffd967e3d4
z8cbf5be14f1a90f48261d285e5016186f7fd4b0bad0151b6285a620f848f839637c7742bb0ada7
zf6ed07b1ccff5ed71cd05725bc34ba8b6d1dda6d9688124d6bce0796857d2e1a8e78fbc58a68d8
z9af4bd3c31de1eadc2c58904cc0f21a6d8b14be091f8f9fe26f731772decf8c40becfe659d3625
zb18ab934779479a45c9d3e169e349b4c1626025c4a60038310e2e794d17318737ebb9694e8ea93
zc16357f38ddfa26422a30a3e55f8d5c3f2ede1c9c3f3eb4c8ce7e721198ca53e822273fee0b05d
zac6e5e5cd2a055be1a15e1c14a838a0efc4ffb570a13526a55954cea06f2307d73bd144d2d9d01
z314880962d6f421f52f95e6fa1148bee55b96bf6ce713c3ccf8147c3dfb560c75f1ae110e6e0aa
z744ffbb18f11c54cd1dc1dc2d1b327f2b5c1966373b33015576fb698de4cdb3a16081165f68d4e
z11ada0067bfa628fc08876cc30bc19078bef506fffc3c3da94a67480dc7c0f8c91c62a8301fe8f
z09ac84a29f4eff5a843a798de7cee22e911908a98ee3074315f89be48dc24b9e49cabb269be388
zd82e09163807df89125adeb94988814264bb313950253548f09c81d7efe4f613008711213296ca
z15e6a702fa4979ff6692082d725e38339e0f9aa4f3dd476b534ffc4b0647f59e8c847ea9149b8d
zad9a16324b22a3c879e1b79831d5227e2ddfedd61c6df6d3e8340b7f641d4a5edd9bcfa30e4034
zacfe94ff6967c4d1292169738e2255b87b08fa0dab7a0b2557cdeab443ce5296dce666e4618799
zce556c187f81ce0a0a9636fd01c0dde4ab42f06e493c4faf217bfdcac60be0d5bb7d32b48352f0
zb93f482ed4cface3f753945be31e450d09d07572711a0ea587dde192004d1b73c96c3103f570d4
z51bbd557bfdf4321e5fd6fab33290123e2b8bbb1a2ef9c348297fe6332abe447c017b9615ac9b4
z03531b8997c7f6992a6e0b6ea9be066a16b821f31bcd584b7e142b0b747f971fe8900e906e6125
z2accf2d9fbc3ba269673305b6bc395ea308a77592b770e31b6fae963873f353835e7ed9c70d9ea
z3de7983ad421e36246cbbd870fc4a67f061bee9301c41caee74a463ff3cbc43afa2d62c28f699e
z2a5894cb74728d948836d63006d36ad026ba56576ba61ecf650d4f92a0ac1d918fd1adb8357b03
z9f654a38493979ded06da508d8618fc82e850ade55247c7e93805d0b97ddfa3f46d0c08835f8ce
z5cddf40d18b3bad3f5c55ff08f0581a873e4e9ed63f9f55baaa6799d52e7576732a132106cf5b0
zeac72979158cef6d92b73e838b2a66d6bfad9acd1f3101e33b6dcc6772495a295888044c7cdabc
z94ab6b9f41d9e5e2340f7df5aa8498c31fe761cbe9127e767145d21e02253653ded0d03fe43c7d
z341a91c33ba1fadf20797b64dc8e96323d0e2954f31e71058c1da6b2e63df74943181d441a6c0e
z64a4b157aaf5012888ff956c12622d95108a4e683db2c27b18a27985a5842bb13df1c895c3b046
z0beee1ca02ced5959d9d149d5d975904841a308ab1e4d35fee94b849b37b5c5ecd73a67d694790
zdd2ac1e9f9a545ca345aa7716baa73ac9abfdfa1c18e22a7b4fc7b774629b49bd082483e88749f
zb1201ef69bfbf399aa320fdacb4b4b54caebf6adada73f47064920c3ef90a684ce49c09d593444
zf4318eb8882f0705f326081aa5e98c3e545ce68e64dd6156f234f60e7432b5004e3a9cb6430b27
ze17e5591b69f0cd7f0c19f1dca8ef2632a0a9198e3ea36d5371c3c70543877e0553144e4685e5b
zff800786a4425c1df6511ed2927d4626671fa551fb919d35518114784051e5eb79534081f93abd
z3c21425a4c1abb7c0bdbc3e007f6c4de658291cbdec7ed0a489d6f0a9ea80675ccce34f2d14487
z094b579e9f10c9daff138f8f03e7382f48d6d54898b13ec4c1870658c70b51ecc5382c99bf2589
z5306a5fbc5f534b104a58158dc9ac9233105e3a6a300040babe8fa0b00b86b60d307406985d434
z65c7ada332681220f329136e5ea21b8586cddc5a8d3d01df224ec07cbb98d18610cf4dd063406e
z8d2f23972466e0d15439d21ffc8d9a2f020e18d40dc7b89ab1e002480208ec690bac187963639d
zfab22d657a9ee0f88199c01220994488892f353d0f3e47339f49eaa8119bd2a359b0f1c27b1fc4
z5e7d485fd434970d296a4595c5f7681a949e70a2429294c9e27bc18f3bd098d201c0f9a76d6229
za8f1776c11d1a45d237f7a8fc8050408815c41d010fec37a5225042638938507a6886f4ddf8c10
z38c3bc45c51603b57a166e55f41fc19f7f7e9829a082bfa566912cacbbc3c4c5b3ee07f0cda41d
z0e681d424c0e0f2fa002a0dbfbbda91ac671645c318477ae270c358d5ee30a7762976a75b40ab8
z9803cf96d90d3950ff0fa570551212e6221b4d2c366f2b44d49720f95e117b2d66f0e6982566af
z67a9c0f8764aedb04383b645eb046392d03ea19cac8c1a99ff35dd4397a2352df0564fdf90bb62
z228b86c1033112ec9979768b80d9f733993ceb85666a7246e9e2ca7b7e8d28f47ebab7c3d5b94f
z26c8adef4e3913a6995ce268cbfe6afdfdde89525b40f49108684f423816c8525e752ad716e814
z7e5550b8181c41e7f3f8d4559241ec073b69ed64b9d219d0738478a7d68df3b21ea5e60b2aef60
z7a8b6f79f8e902e25b5467e0cd904a3a947a5c70b40e4cb741d783d4b7b863708455754404f37f
z40d1d7c530903506ff9967c4fa86c3e9c7adc553e2efdcb499f2e15b0990b66d2301d31e2f5505
z72d6e6684158e2fff61524d382aefc2f218aaa8dc1fc0e947d8a45212d51707955da282845180b
z1c66567cd74702ab240ed40753b3180ee5895818e99d283d65a1657653542b6d12cd75a7b092ca
z39804e65bc28e43f25d26067c08b68daddfcd56c3d398f82acdb369d77095e2bb9b9e29d0d451c
z5258c78b40af3c95ae0f130aac7e9c9d92e5ba32133cffcab6cc6e547dc660cd8cfc6f98f5790c
za30bd7f4bfe85cfc9fb14ccbf0e57b3f3ba217de41f9c57fdf46c26812e3959994492076c2dad3
zd22278dc87a0d20c6a397203897089d40535bd94131ccca77b8826880da880b114275cb15980cd
z7b3bd68c628279a56e923047e268e373f6aedbf3a7ade033e03d0c8d17aa91ca5c19e50caa1468
z1649558f52f342f450e038b69eef18600d47e6606b0a91703cf6aac5727426ac466b7945d5d4e9
z076011ccd86d69fe6d5a52d6b14460856ab75959d2ea4b74c81b4d9d78e4df1729b0d8024ae794
z2cc7f171fc9770284741aee2d293b46467100d8d3c438e324edf2232ad636138222d9d8c1cae5a
z809a2e255a9c9cbea226fac1cfa25243df37c0cc57751b71067a77a5e5193b46f36c1921f981b9
za7f9455fd925688174396ceda819393f6dd6df6ee51d6e881a4ef4584fd04675818ca86c4f005b
zb72fdc7e9f9dc3f15208a6878d945b9d2139faebcec5397bf5b48168a5b80d051b221ced9cc8ec
z0187effbc3230c52fb101c69f71492677ed38f0cb1ce5eabd517817965da646daffe48576db50b
z57b33076e3bc6c3db90c4aed1c0aaccc1b08252461ce7a874ef3fa91045d60925e72f1ba445263
zf5d0953055672e47f79f39e94da371e72f2ec5d0334ac6bdb2fd78db1ec7a8085016888b1154cf
z877415b0503136fcd3db8c40e371125b94877cd1841b1854f43b99c802f8c129eeb5a6c1f965a3
zed288de0b86c32bde15eb39818c3abed8e51b9cdb12a4f4077176e6163b4dbf3a2b7e7d9d5437d
z6e8ac60672b1774e6183bd22e99af905e9f4424ba42b9e1570a04b63d3095b74af40ac65f69cad
ze344737ed2583ec4fed3f39a6169ee7382a04ecba1cbc28561428173995f33d4fca2b1934a778d
zacafd143968d35bb327797ed17dfea47f79f781783ceb597ccc9185717bfdcdb1df532a49fd7a5
z023855d3d430f5507122d45bd2b1fc44dc29aeeebc163933876f2157e0824331436c078063bb1a
z6120d28e79ef48dca68db5c1ed44e1555d0e8cb98aa7d284aeede74a926631796280c5bfde7dc6
za3bdea65df5318e988ade78f3bc567598c247f87adbba2510c1cd5430c09e066285c00071eb38b
zee0d30eacf452f951bbb15be7280c248107ffb1b5ddad6587999c743cb6c0de9007f79527bff30
za20d92b4f69abc4036901dfacc3b9ab90647446cbe321f5fb1b6dcb6d8a014c8b3a2ee3ea6829c
z180ae03be0a4ff055f7eab899b9823176f86bbed260d8a892afc2c9ef6bff82dc50e6846dfcc68
z60b4d6743cf8a0ccda28d211702768ca7de9b39b1208bfd1e32a940df68a4b841085ffffaa65d2
ze8ef6921472a1256b9eaf28d8e63a3602b401555c39f176d40ffa54c93a5d4285aaf198fc9cc3a
z8bfe93ce0e51ea217ec32c448412f0363a5db08438c6619937dc433e8975f7f63d7226c63505c2
z9fd3b3a0d0e509e6a6d38776fc1b18d36184f652cabebd3533286f827a481cf48dc3d77956abd3
zc45d5e009f86f622b835d5681ff738482c370fee8dbfb81442fa60074d94ba091afd0477b6152f
zce23257fb929031fa2aa3c519b32f214c353cce061a02586a413832addb1bb49aae4b59df50759
z181b7ba73b4c6b4583a78d99e558d49f518f913a9e772fc923fb7d278a18e953d300e48355310b
z152f73a9a53d388a027635c536d71d17f89f0f0ae2d92079d14ff029fdb34a9f771d003399a978
z31f8c36ce30d68b7f9b970b179a6a02a78f3cc48ac3f7ad915b0f8f7abb2b70fa19d6f2bd287e8
z877c85af1062507e0ae4bbd884aa0cfd8bb4c3246ed7794e1271e77139bc35198a8d4da30af215
z4162fd125df753e8a1534abfb5dc260bf0aa450b83679fa2f270f303f2be5c006fe29e44eefb1d
z3142605a10801b0a0ba5980a2f41ef0e9e52e5564c3c151d838d0d376905f88ab8e227b4221662
zea781c124a596894f63a4c0ffb4681d1faf405acfe13812b6f23b85a34477c75809d4bdb1c0f65
z85d0207e1f483734e5255abb4e17b3f373f5d0e9c02ed1a8aa75c6674edf71238e7f4293292716
zeabfd28cd98cc876b2a3972b2289831b50dc078974032b8b7693ee44e5aa8cd49ab73a842f30be
zaab7f287091946283ff76fd93bc39bfda9e4d5055d238381c7a5ec45d9adbabe76da7c3b0477c8
za5451cb639d75afce2b8aab41bd27b0ae9cdf9f4459e2b088e718ab6d9cbe11ee528637214c61a
z944f9018b0ed8ad3fd6c95a143188515b5e9ba1a6e4ab6fd2b04e0ca375c8db8b3c280fbb494b1
z7d05b5e6acdee44fc7be7f80b0c5f4c32e9893325e6dc9494c7f180e211175e532156da7ecb839
z68537ef0c73744b852bb7765f2ff76257ce59f63df3c6bd394824351be44ef1210208aceafd0d4
z9006dc4850a81298c865038c730c8c0ca8f16a7cacb0cf0666c7ad85c9337968682c4fb09db590
z19b0a4bec681b2fc4ef2d973dcf41da2abf63909c2f8d812d5a8564e62e4c6765db765780f3bac
zf9ec4e6ca4058348b671586c087b1527c628cc1d70e5a082e9ada8d45ab8af5c030fc6bda6cf1c
zc7bedb24737118d64679e7a90389fdc1ae71a181845cc438b7712cca744e1de525baba27cf5342
z027bec68aa60b2324ea40a9030fe7efea28caaf78e896dce25627144fda63b086cec3cb0207605
z96b86e182dd105629429bc5304f7065c6eb41b9be727bf30437bfc9898aaff75e772d9155b6334
z12d94988662514b6de8779b7cafbe6b63d9ec58288f46dfec86c426e7a41a90169785e5b0a2c06
z4d8ce0cd29a08111117785ffaa8d02291e28f450ad28110e2b2adb19d20f38aa8ea091b87ccdf2
z6456c2aeb8df52766a49e49163893f1c020ff7ebfca5be394d71af37726bc4280e57bee59216be
z9f29321ff0c9e5f8a808f22387c510f58775f63fb2065e8e36b05e038a4d2189a7137b1447f1f0
z05f583e6373c0427b6b6a793748d8793be873bdc1239e24e516a2d773efef1fe27305737dd784d
z854190262c444cc47e4c153ad6f6fb1afb4ebab20a969842814e69193a8f52bb6a4afd32ad3917
z86da41c7ec79ae2ffe4073686bd9880847d04843a6d017e6103af0ffcd819244ee1105bf483840
z91cf9dbfe27488e2399e4835b2a5fc7e32fa06d4ab065054fa29e4e08ac6e20b6edaedc1ad9d9c
z9b847ee07c1c7547e1ff1e915a494115534abb71f9b7bee31bc079bb6e91de6a8e73a36ed6dad8
z785666d3a4e03f80fa4d03c73dca28fc4a2b2506625f519e4e0779c66c15dcfbe4b66f35025eea
zb1a446e70820e46ce6c8901fe65d0ccbaa1723868402b3723fe1a3a439fb5044a5aab87e7eb865
z39b431395d32b86bce8841ad734d8dffa4f843e45d041fdc945a816ff0f7d3f02f948694329b71
zf070d91b10ba71a99228e8fe4ce1eb74bb6ece35f862f2f95e22e9ba2f5d80663f7bad7ee73538
ze1932e8b3b7eb175c5e6b7d674ef5c518307255344c920ab2162461cf8a4a389adddf74c1f7b62
z0b908d15a95451e5236075e542ebf58298522ee9d168d4f55263c6acd0d141d6ff721389a36b40
za62198a6d7be4bd27a7205f55833278a66570dc0cc189797db29178fb5189927f22daa37003bac
zd8aa75a334c1e38a788d29003ba02ef38366b3339914b2054beaebb865ac6ede08a1b47a402f74
z486f2e126b70a3b9b82b5bc2b157ec2f7ea13d9b36432a85b8a3abebb945267b0aa16eb564bf05
zf8f33cdd860f2d288067b664e4dcce20047cfa42306ed67dd7007f911c2f73f304eb8e150700f3
ze359c4460144634b085d4bc4178fed02185348bedfe18dd3c756bba766577acc63e420ca7593fb
z0c089bf7dbb78f2161c5659c3bc2ea4b0e4cdc2b9a1c4445dd5290f1555a89284f21e44134334b
zb4b370c17e40fe777768b6dd628e084e91b12ad7faf89d9c59cc99deac11d8d004cd8a2a5ccdf1
z660d69d5db6eca893801261de4dae56f8d0caaac1bb354248ebf769cacc592e2b3656e53c7fef6
zbee564588caf7e964fa4d0bfc9073cb5e70b5acb63d4b8509f4f56feb92b587535400e70d0a6a6
zdb5eb694304e5e191099067feebc50acfb5a70d3884acf14109d7c714e937109b2661ebdb6e579
zfdcf0796e2ad6dabc5504250976121d1037698968698b8f5632234ef71db9e728ff820b836c603
z263761d50d242c5c221c91588391a74a697625037953c44248a33b27620e2d0f9968fecbe6dd5a
z1ba2112fecb5795d2ddc93c6257143e436f48d9281ab7279cbb063784bc1a4701d1796313ae7af
z468689807b38b36903bee08880ed67d712f388de9f619eb07a89232eb5f17851179b612f2b5a6e
z6cc3788b154fda3a6a6f82643b3f79c706eb7918b185683f1a25a9053f526851c9a3157196027c
z1d19ed1e89957d925126aae72d26caedae664514d7ab3b63c6a995cc10d103ca3c5917409f7db4
zd509df40c0b287d50ac4521c044137df36bc03fc74b58efe7bf215d72ab23a8b425f2a0b20024f
zffc478b3cbdb808922989de9d4268822266891f91fa0d61aad568a6a494923449fdfc7a27e5eba
z2b3b3ad7cdbc69d52af793226828d5be1c7e4a90a445734517ce5aa5ec8c201f779cdf8612ec01
z1a1dc66d177ec8ac3fc1552db40e5e27e933bb16c63a490f58bfbf3b540ab037ecb11683c0dda5
z472b1d35ee19571fdd3cedd8790982b091ebdccdbeeb418e625cbdfde46f9a6a2867749c373678
z9860f76feeea7d3c264029976a814308e7510b30c778c5516a7ccb9e0b98c6ee199300cd10f912
z38e6dd9da2c4888934ed6600a24bcec6f239f764164644efc0a31df85c45d835d7e8e2befdea5e
z3c7dcb42cbcbdfa1a65e9688f7523a49d503bc9c7cf2dd26e2ee238f66642f2c8020fae8a09967
z85b70982d7391d9103be61c1128cb4a0c3bc800034d37b27aa16590eafa0c994bea2a6a4332985
z9a55f6c376274dc85662fca9991faddb547395a8393aaf7743b04098df39dc0f676fc8a69ef3f5
z57b8e3ea9c21d74007c77c8cd84274f57326be67dbaecb009b3cfff21356bd04206295762095cf
zeca3125da35286f74ba314b27c7dc1c568ddd36003d70b849655411aa18cfbb08e57c54bcdd968
z6f7ec4972b3ec2816478baf65d65ce371affc579990e4c64d0fa14fd97b70e4adc20668b401291
z441475f76ec5faf1c0425224668b2009391d8f2e5f8a701c590eac438d32fd9ec5dfc5387eefa0
z729e8c4e841c41dd9fa84dc4c25569553d9bf2d579337fa7a179c04e2ae3ed2664647fe6caafcb
zcff64fc9dce29db98ddaf5b10e9268ee0391fee0e23dfc4375b0bb5c890015d183447b41f12810
z066cfafa6644f7bb9c9c50096146523d178e439fdfa42a61b841084649217899baf2343e739425
z6ed12ed2c852829d5dcd346635865f3c4c4a939671032232accf238d88c79aca596e3d343fffa9
z35f19dcafcf5910fe4e2c8bd1dac03e895419cb988629dd68adf7eab0d7d53aefde98df7449fb1
z6fe477dc4ddd73cd71179af052111edf6aecfbc4b6841ad4bc8dd152dd55b22abe3e645eb7925d
z24597f4632ccefd6c909cf25c77e5deba82d065eae573c2cd92e89004ad252b0a113de88eb7c57
z58eb51adc6db47349e074f7ac448010bf915439e06c8a6374c4c5504e45632ed3914b0f81e0d05
za35b9cfceeab99382047fc6efb68644aec7354a0058d92623aa59ec652cbe5c3a039f05db579be
z359a1338da278cf0e57ba54f67e98a651a34dbcd2534572bf9e2b4dda67ce2189e4ee90b7d99d2
ze1813c97c443bb9d193a422620111961c1b1ec7aa9e59a39221112dde64186abd9dde88deb51d9
zc091e27bd1e6639d3b4ab14bb55ef164bbab0e2456fceb44723fb92d865f4802e929a92f3cd2a4
z9a8723bfe4262a97be1391eaf15ac284d321e9bb88881da128244090736c1574210110581b2a10
z62d8804c4ca08e08fe9e33abeadaad9a42076cc2c39526181c58af0d169409a5c0f719276d709c
zbe582d390e21b959e06ed6650a111e3c0068f7b118a62d369633c502e768360f2949d7b2073b89
zd5df18a88aca8cfa146c67bd5bb804825468605f4842a98b6e2751dd2a7164b45ee17eefa3c55f
z1f20c35575d9885544a436b64151a4270e79fbdd7013a5a227d2ae11f45f646e6aefd25a6f7d4d
z724d66a2baf6a7c8cdf3a6110ef05baefd8f24ec8aed66d19394ae8b3c65832a584ac73eb47c98
z9b20e8d62eacf4569980a96aecf1c8ed9713bcad196e7ea130743ca6a29939a2f41fed2315a349
z4ab49a220627e00f185221592eef2bda12f6573a3ac0a74292f2884f9be939792ad880274ecd30
zdfae0d5f74d17a7a0bc84eaee92a7abfd91be0120a035d2dd7f4b529c36fa23ffaaf40e755a770
zbbff812a2a66adc2e5f210a7a720289a5bf06a488b6cde73ff05c2f3dc4a005b302428118612d3
zbcaf84b28ab88ab5694ddaf84ff3e753a34c7eff691b897bf89dbd21ca6d340a480996df3c9e05
z9ecf9e897aa272f92baeaed76522506c85bb527a4a1d757008d924f8c5d770a17978c69bfedbed
zed2625fa80df91944a5a9f199af8612dee485aadaf5f9ccd96b3f8c9404a51a9d375468a963901
ze3ad5677b0cdabced6dd76470ba0a4ef61b20140424e0c528d88ce49cce01ea5ef5b39084e9d97
ze3bfd4f9bf371c1a295e008745c4d29cce8fcaf1ba4dbf40107b9eec33aca4af8aae37277f4fb1
zfaa1c9b7d474a3f95215f75201133a16c5c467667fe267341e06cc58a623683b63e9707fa453d3
z9abe7bbeb8c3951d544696832f1f1a8ec179112bd86e131ba5ec8b77893b55d2b2dd2f5760a310
z8aa9ef3917bb7235a5cf5b061621da6a8846329f2f307a91a7011688e25791e220123a1b09848b
z4c4edb3523b28a82d351423e7828c6125099a028476eceede27484668e14e5efa501fa6e05e43f
z65a71eea10d93043bd7ac8e7d90bcc26bb633c92a4a0c67498db3bc6d378f29dc54f285449464d
z066a1c8e0e9e8c4087d661ba345e41bd236e30cd5b1862e0e55d6b96e6bd4c5fc0095c87bc74e0
ze31d40e61e841b9cdf3e8187473e44f5162f334ccb1c0c4019e53632524a5321d785a1da995d50
z334f8df7603cd047e2f38ccede9e9f920402eff4fcc507c675d84d1d10981427720e2b02a8e62a
z7aeea31665fff7fb6c70a7e1c2c93399568a601968d01d95da3bd1d1baccc89bc74e7231298b78
zb89ca6872e89b5f2f873d05bba5611272ac692032579e0753a00d8c9aefcf9de347f30271f13de
z2e39075b786e1f687a3c54a764ed51f2df71e8d0c680fb99e35c8013fe313c9e540608fdd736b9
z986798769712eae57228084fb9ad3f5d228d808a7af8d05a5b66662ed5bf4843ca395d7152adee
z5eed41c24d12c82d8a12a977f038fe3df2671738989898e4153876faa53096b5330071f6d5bcec
z4fdfe2e124c5e2ec3233aa696df301695033dbd23f5f4bc9f9576faf7f9dba91622f35b1f8db04
zac7ee38a0e429d339bd5e52909c1370124d5e60a87bb9f10455ae86015f1b7c95c2f4cb4fe2eb3
zed79b15baa013e3ca798b2d38753202111b82851889a7f1dee3bfbcc109d07e4c0205051ea1963
z65bcfb4faecb6aa9f0691ab819f001ca6aa05e15082062415e882f083e7509e8e91537e6b76ceb
za48196a608f1b0c7055bced1efc7f36e82fb444316e75d4ec7399b5189b54cfd92ae67970b2511
zbb3da7eaaaec01930a7e945a60721f0b5db2f470743d6609a823de9ec2d013e0f42aee2bb30343
zf5d1e00dc388d89300098d0617c916a288fac7a1379d5e25bb49b498ed3ca5fa1112f12f001ba6
z7d73b7c950cb1899b18463e0a3f863043e40d7a8b55a47ee00b239f89127c5590f5adc0b5669a4
z2e906e3661f129ca7080c1c637c542e5a8426f728771bf7b6ab84b4315c5c6b4b27b14e4af5ecf
zdc60f7ecc9c898b19c89e25b5f5f5e32c20edf57b48495d2cb35210038b8e7668cde738d908e22
z73a92915ab626867e0d293444bfc2244932939cbfa3c04c2f6e21063a9ffd5847f23176b89ea3d
ze06d5d2fa9347cd6c7d5dc9c57549a4904d8214a3f680b3bbef5513dcdd60d15f4e0cfd9accd4b
zf7756a0cee8227b61ed47c665a4b5aa3a83efe3f96fda18cf83fa1fa10d8d902387d63fd773e9e
z8685e80e794cce12628391389b31fb94116e40c42c9e39487699612b05becdac09f1374a93b1e0
zbac72266f1455ef22d4f4c1337d087d4c7bc5649e9e968968ca77b2df82da75686f96c85f32e35
z3c7fca406079655b12640a308cc4bb906116889d5f79a37986ad48b787eaefb995b0813e2cc095
z3d31b4b7082db571ff6235574c6d556236585d9c6afb5a5d9c8bd246f8bc48a5bbda3ee45d0bac
z12c263057918d3db0db82e7f660514a6849e9fd51c21001f3ab7c3bfe7430658f32f6bb027e6fa
z0da65890f7f62bc5fbafaa917e165e8fcb1637059c55bebb77df7de681e15059b6b98c5c774adf
z6ec4d4aac21097df98bebf2d87dd73bf0936b7e7a8f99763253cfb8b70ebcf7451b981ec52af54
z64ba904e8662ccf83aaef74c96e3ffda3c084249d4665e9c947341c570d47f137b6b79fa090ec7
z63582443ea4af15dd2de4726cca87ecf3dec442ebd2fdf113b4107cfb90fe32fc0ad47e28d1a57
z85456a69e4140166083dcd4e68c7c32e89cefe0af8407ce53496d96f416fd12b14fac56e3dc9a2
z1d336df39d5d09898199089f745f5037af82064c14aa94b5e89e2927a25ea96735e5bb54f27549
zb7e2d80c012862b715e0918b82c0dce0b7a1f346b2ab9cc1e31463a07aff49b5a8d731790acb77
zd599e277f5e194d45813565515593bf60d04ba0f78241c6a20fcf7a8c2040329dd25b4410e7d8e
z1eacd0f30cab9df44562e7b8d2be338640eba7ab273e9523064846eaa2afcdd8090f5393a7292f
z816480f50f3ae76d58d0d94b248f617592c3d749a09b30ac3e898f9e5057698b24c13bd912e529
zc3404b8b6df2628ef0a4d95c08742ab20c66e02163e707ceafc9e8c833865d195aea6ed4d4a97f
z223fc8ecdd8369d4cdd440d4060dd307c1576dfbfb9e781f8020523784c7d3deb2951779d50286
z46134f36ed13f5a74184f250017a8d7cc5278e4ed1fd17b91157ec5ca1af8a1cb1590549c75999
ze2b3d5cea1e4213987b32bdb37604d46b6c4d161ce4bb3d3e83111c06bd8c09bd93ae49ed01319
z102efcc848a5e209a025411415d792d21d628bfd1baa0f5c13a34ea991e189360038267210c9d2
zc5b6cd550c5843713ce93e17d4a4568f227ad1118f19480cf2cbe6ea18c5edc402f3d2e420a054
z22c73c694e4d71fbeb9682da3d092b4a28057f268227b2fbd058aa08b84fbab60ea748e7f8b6e3
z83a8d0ac78da4e89638e6eeb11db1f89508669a62c4fee7453e5d5966ae645346f1c529d849c76
z4aa64cc81be20811b4e8d483b5014dd64a9ce67146373c564c4d0f7fb463ddbd5ff5a85cb7494a
z6fd66e6b6575217de2afb85480dda25f642656d398423ce774f949f0f9c1811daea6a8ed84c5af
z57987070cd035b863788fad0c0c7dafcc8bc728005ea874a4c6d94e14ea72b92ea29f21fd8aeb2
zb2ae69e0d1a3d2ef254106d1d35d25ee22b27c7cd4a5ac3734de4612ef9da118225f01ea06b9cb
z4e8f3288025e7357e33921ec91fbb6c12048c47977701baf0ebebddcf50f86ae70bd0400a68d23
z972c5d05154e72a3eee0dc318d2798d0735d0ba837e4f602ed9903266b5c9b68ec12fda5576850
ze5e3bac6c34557f8c6faa102cb550c46642bfa5c885d699fbfb8660032008dd5a0aa878e3dce88
z4a3f7ef865c2ee171a7e9fd13b2145b586e571c898c06542db85e131cc6076e9a780763a6405cd
z64d90ab0a998a063d85d140aaabf00ccf6a2b4dc4f97448eddb809b05119b62d66aa43f6f35ca9
ze960ac3d7e7cc4810d809d9d218b3e9acbd6cf41acb8f3362099f41df2050b120f2b2f3a9973f3
z9edf07f51a14fb5cc52f8959c8ff76472163c61a304009fa277842e25771a54ced9273404fdeaf
z850c06ec4c3a597844e4c069e4491706ed6e87ad7fbbe2301c3dde8f93f1779abf7dd369b361aa
z461965ca5a1b11ae5ee4ad8b9e775f24a72ce57ddeb11d19a223c0da5de536b3b65a95fa48732a
z0a920bc047f9dac262f5f34d7a4a199a6a14224fd6d58b6ba03097301f6432c9219b5c097f2931
z9e59390d4c660fbfface991e64634101d7d79e417ba24fee5f449e30414620a92ce33590c90009
z569024554281c16b0325452d28dc7ae7f7d7121c43298463baf57028a3b388f8c37af3b6676a90
z240bd19c706284e48b48606d748aa60f4cf8f9d1a6770314fbee988c949fbd821e7131f6bef1f2
z7b524a6da85e42d2cd61c1f26eafc2f4509b871de6334437234549d7c96e0b81e399a63a4f3249
zcbc6c4a13cc025ddc0e0c20aa5d7f174016812e288ef67943d0ebead9fdf8859cf675887613372
z84d0e200650d95caab83ffd59c77826a07c689eb6a05fc8705959d3a300fd701f805921a0f8810
z9bb8a36c32e313835482f2bc8a1047b4c8017912a2d9d33bb350af6705c4d66d613cd0aa22991b
ze05b7aea3ec65e5922982b95d30d3a8b05d84cb368f4a3b529a09e98de7cc1cb5f3fe4833192ba
z02c6faa9fa168ea73ba3ed3df08d9b24c37d3a08f160d6586e7ce6ed634cc995007fda9504b8fa
z90d79e4a7a2c645241f0c84de46833b5a1549ce1b09507388ad28610b0822296b1f24bb187d893
z9fe9fe6344e7cbc3ea76c034429b5112ac833c513ca93b738ccae515b1e96ff7e8ac930781b2b0
z1dae649c6b84c2199dee8fa29e87d974f3d277ea59b6896031bb6560e80626c556c0be266efa8e
za24048bcbebce4ba821314fb947b8e60dd3c38b6237b3a5e4d59c7d3dac0f5a66177ef694deb16
zfdbfc5d8458a9977bb9ca0571c381a5ebe3243ad71d43a2ad932825602f2b8723337911ded2058
z032b6edc69ac7d512439421d34c22ee5ada4bcbf0e8315cb7fcb04d8c20f1cca686e17959c4fcb
zdcab6f56ede7f954fad303b3752a44fef622b9a04898fe439e1632d2d8a44dd0f582e2fd25a3e8
zbed097609b99ae6806d1d9ac653e1013dc1e0fb01a085663c83ab5a566f675948bfd9d3af73093
z052ac193756dc7c80c98da1fecd617aaf5c52bd45c298f9ada82fcadc05e9714f95e45e2e46317
zf61ea33c833d87b0c7797de197b29ab97e575d4feecf7bc79bbf1709b9aaf82af164e83a60df10
z582f7da178d773af685ca79a35ea7cf496ecabeb1234a14cd16774f7c07e6183a2861314194b94
za2b06f1aa619fa2acd3e7a483738612023e9ac98d809e15acc57c990326a8fe417d756ac73162a
z3f15478ba8b7d7663936b8d454ca1fc6d9995f9efe721ef05c749c644652d49c64aeac0a682090
z927234540146373348f88a8691f98b0c497955c10898515549c580c48101d45ad4d0d5bf30d895
zf19507b19e45a95f5459a94316a49ddf811fc39f4ff98c55ddafc14a3963fe8a57a48ee73b5f7e
zcdeb5fd30988fd27bc489d92d90af7c7392fca94ccaa330b49e3ed3883b7980a1a6f209850fc03
z6061d22d2a81b5998ff0d719f3c3d068132d12514f5c3c6fdad79f09bcd7381c7f976173054c1d
zb909b825c8f273278fd00af06dd6b7e5866ba033fd0ad02ece048d5119d3839fe96c0d34fcfdd5
z47475f064a3f758293566897eb5fbfbd654e952a4875d0b5426c4425af88972374c0c226a6e327
zb6ba6e6c83dd0f70706cc38cfe47fe97cc90abc23beb85cf6206cbfc003f896eca2ce8644975de
z1288b5d0fc0d8a56c57ae5b9eebb6712286a3a143a2f052a0fc7c7150dbc8624127e29476d5ebb
z7db2478205935d20ac55650e13ec7f21a6d37f5164bebc7918532957431ab3d4be7d7ead33c64d
zb82e72e5114b2cf9b0a44d074cc7b47a340e4c4e39b48a529a7d759d9ad09568895125cd44c958
z5283d36b1b70ad072878b9324c4b7a3b7a9959686479da216ff6b426a37a4acea54b7e8141dc94
z9413719ff66dff9f75fdcbe83384f488548577f23b5c9c89ff5af6ab8a883b193a41615956ddb9
zb443a28b0c59b2e3c675a62e4bc129e26020e41386b903264107f36cf79369dff2f294e4297260
z4218144349e4ac3f5442d84716200ebe51e736788f6f1bcda403d8554fb31c01babe088329ffbe
z81f19a96b474adc90aa31df5519770086124df7e9273f170bec589bfb46f0245b8053ef45d353d
za250ada40207a887c304c80a85b33285522b37471d1b51d4f54eea042e3f07e7aa169034f0e694
z4bbe3ea55ec4bc377d5661af57d4121ad2931fb012b874ecb0922f71c1fb6b489b44cd73070ffb
z807591998add7235d6f7ecde0b845097fa08cc844b870f18bdac9b63d7fae4a42a063df04f5f0f
z3d73f77f24e3a0f3b782f433dfde5d940037caf80fd793074aa6b0a95d27b800fd554b6a98a751
z1ed946143851c591baf36dcb79405e8acb1507b961c38a83b7e00db0895a2d858f83ac9daaa457
za3d20979f9b00a55765fe07fc74355336ecc7ec1c3800d0bc64587288cf699010755d14241e8b7
z8b6128b23b1eb2a6788bd547632e0284153e5c762f8d89756c6817d7e4110c6c1a4819f7672155
z59c709e05eab9651063198b0ebbbdd4233122ca967d01ba51b0becaaf4abda3f3c00863c1c3650
zb611246f8b1dff7f59ba9205d9ba480ef33a0b45324a70c8828cba515d38be8a5a1dbf7d9aadeb
ze15c40b740299137ee35994b7898cc9091e8aa849dd403d01f9e3f85842e5ab87230c4b5e7836b
z6b699651cdb9b47db71a4a6abd03bcd4daaeaf8e231f2ec71982d4f2870b57756afda25263f8a8
z2bfbfecb13e395fd046551e87accbb5576cc3113f2402be279f0c475ea564161a7366131fc94f5
z032b59ba98a1678f6467e02faa959286a1437716ae28401621c62cc7360ff54d12b2e2ce37fce3
z67d6408a7b29e43a4b3c7878db804506d0d2c196aaa034f95033e9df1849effd1f8db24e7db304
z1c22b1df8d654160dac4cd9998d789fb589e341fd27c3b400d287b71e6a9b6729fe13d3e9b584c
ze730d8a80107f5b6e12369ee143f668e3928fe41e6557c8b836113b54ae0f208d8473dac52f74b
z13a35bce07c2e43a68c860b7029f60853a0d57f8b58f221e4e071be132faca7bf5a195e7395ad7
z57afea33ebcf453693061a54013d1a2883dd152a30b9948653f1f89fa962dcd2adef88d5ba2975
zf7f8dcd52767bbd8f67917ef1ca86edc5d7cc6ffa7d76ef9e117079cbce5df22a2bb86635d5d93
z127a81990ce80603646fca235663d415a8ad1164460a2223ebb0944e2878c5a357aa5fe97c4751
ze069ad87d61bf55bc7891b710faa2ea1dedc31801e73e3f476b4c254b2648b9df44c17a67a0ed6
zce482d93be0f57ef9a8e6e02f47a2a034ea6c938de2b0f8c452de3077b9e383556eb2b0c09cbf9
z75a3f7f2aa0dc205e5d72d8af1993f9c3fcec2399fef3d9ccef650ee6742a16226ba5243d4d984
ze3c6690da0926c7d66e2d1dd4897612dd01a1f03294a970e79a6cbf67bb2137d918752612cc4d0
z48e6860dfcbdbf7fcf5c98dde95fdf91838d833a647a9abb78a6705ca5a163a825fcdc34ae282d
z05be0885a2a78191f4958703a494c936309f0df0385176d15ab0b374e64b5b36d8da0ad2aa81fa
z17b436231fb42b060c648bad64ad01c5719c4df3faf89f1eecc38e321b2fbdda8fdfd4278a79d5
zda3e7e8567c7fd0280dd8a4c4470521cb5c1939ee9557dd2a0bb9b998db8719f28d0bd49c9e2d7
z40a2210684ce7dd6ff718934dbd373d54b50868d49809e6e4e36e09954f83a112004bc460d454b
zba9bdff1be2c83b8812fd10815517925993c8e62d367a508284290aae74d488446ffad1ba19540
z4bb20063eda46c6583a161a00ab3e1fbd95aec50445e14824e0777fb0ceec336c4ce2858ad9548
z16995fcda617601895e39d88ce087c198200638521610bd172ba93cf336dabbe6028299c694bf3
z8c5991ef4ee460c8593293b96e7e1dde12dcb4a282af5404cb27a9d0d8378e09af3cca4f630c05
z59f0f25facce908d254c96130c4cf7e30f6ae94633a03b8aff0d36589a99e3bcd806af220b5922
zd87618e7f7d8761f7dea0340f0b536163d5c2d0210c1b9c7890777e0b6ca633d073a4897a275ec
zf4f04f7c1ccb2d5063a5d994bfef49a6a31c287ad0b2ebf06a06c070069246527168282b0a99e3
z51c3f327e94b3de92d3e288caf9736237cf46c2520bc3bba3571ddde2608093253aa8bf15b26f1
zdc399990110a5f8adbf20096db0aacba8c943c463f7aa350a82d2313f93f7de4b7c05eca36cd7b
zd868827cd2497facbbb43a1dce0113816eca9601a54e496b88b20113de17a92f8b84961e25c597
z00c60dbd05121772b0ade6a3833aa8543a4ad1eac0759f2dcf4d1c6c3cdab71ec2c1ba53e55d14
z0bc2cd65745b4ba7d1f752f8d38da8ed20b3e8315aa820d40de1103f65a9a8874028f5e3a9fa16
z72a835200745fca5953c52b189e21afd680620bc015d8a66c27e09b919214a8e75190315f947c4
z24aab30b17832a5d486d3811e7ff170a05f2edf0df2464201635e4bceada394aa4f2953e85eb74
z6a9fe5e979b4f1b57d7cb3ad35cd646a7c0c2607e3d41a46ff0650a9331183f62b1c9fe87221a5
z8c0d49371f780ba52db864bd91a86117149b296baedb6b2166818a1b34c1eff214eec245eb375c
z94314d569f9f5e60cf102218be6f7ceb4877f5ae6cb91cb6b5e2b663fe00cf26d5160273ee9c9d
za18968a41b3be2793ff24ebcd7a9982e0ec94a342a916491698bd800e24c06a2d37d8828bd9d68
z1751faa6fcbea76fd8d05120a2789fae1a311835c73f6d4949d35affdfe8fd84fab5d267cee7cd
zb3a2ada62439ea28278ff649505143ca015269520d08418c6572202ebc0c57ea32c52657d53f54
z98d6f279db11273e108c268e1d2e67b397c1cf933ce703235ad78e0669bdf1265536c829556b01
z16e140a8db865d12cc27255cf94f123ec5f4296320f3810481696fcc843f48fed1bec26a848b52
zc68b3e75e235986ef9c23b05be97d6c4e96f3cccbb50317289d83a1d3b16db0b3443300db7177b
z0dd0870ae0217e8e233b604ea9efe695d8be10b871cbd32b1ba4a45565438312631383d0c9fb29
zc0706767ea0a67b01c05fd2a283af1fa19c9dac9dd2bdc4c3faa9201171208c261d70dabfa25ef
zf65ce36ccce9a8d4bd1d0a46067a58c010f2256b40e13c52e4533ac1cdcf7e112df6f1f174363b
z85436fa2c04b26e0a90ae1d1029e53642539b66cc146e4a5f3f703421044d8f54a694e3b40265d
z751def85b9ec7611c1d0c3c3eb8107b02a4e0fb3b11cfe995667f49e6c82e31f294b6e5a6d76bd
z91ac080adacd08af8cb184657a7cd96c5f5b767fb4a3417541745a5091c22b616ad47b989f7b5c
za34d0b25d866d726e09390433e3e48daa6149ba76a422c0839c9b5acdb4cce0aa480d2d36fb31b
z1ca5edfdefae3c82de2e63abec024b2a8ae2b09e08dc97bb0068e83bd1217f7da8ca7343d069ba
z91624f819a647c00a1143eccec360b52bfbe9fc89d346f95feea509ff6cfcf226db7db59374818
zc2194e283e5c541bbee5b4c38a5c973b811e7c7a3d59bebf118cd5960798134d802a43dd8cf80f
z9050bf238b04f0e6284501578d7daf3bdc22bfd54467a22909566ca427853e22a947f97858ab21
z9a2e00897072b7f2cfcbf252e7d8046368895a6d62fc18ac85f5abce7b022dcd25d277883ad3da
zba2a5e5feea96d2b1fd634ae27c0a3279be795f16e280a8d178dd45bda049bc0f321e15c318349
z46c16680caa8f7e5d6295ea61c53fabc93ce1717bc6adfa12294d0cc91aa1e823239667300b980
zce8d8de1bfad0b6753cc9a81fc9ec855835a18060716b3c350310174a827325988b74b7fa73ea4
z70cf6a6d7ee63201150631c6d5d107686cd3937164a9bce5c94f2d0df1e9d16d846a71786a6518
z87718a81cc384a13ceb27f7655d004505bb913f5543bd16fd02526522d526d8cce4f8c1c0f7a31
zd49a57b3dbd2190ef7e5a9dddfcd01c4cae248e869740d7b6ca33a8a5d2ece112c76da1151f919
z9f1d3b077eb98114b7b7fc4f4345d00137ff523a1f30e0e590b835d8caa5e2570ff469ec923f91
z5084ed9f08af87d80a53bbd2c22a0bfe254affdce7a9a9fcf6d047096b6f8705b4bd36005e8e36
z2fd46020d80d3bf041129cfa484f7d99e8361d6fb65a516b946a6e757dd29534776de6ef7bbfa1
z3df91029a0d508a12c431b9234b7fc3f8cb5e73de024ce200f5610a8699f3165f6f0828517e200
ze9e3f5c66ecb49b221285d7290f8ed4d7558f2d3fd68f92ea32f3f3d1b5fe0463e3727ffa5ba0f
zb88ecea70ccc68628b392e600e316e28e0901b34f824a5c9eb85151d9ff2a03f0f6c6bbc9ff758
z96c114d45dc77ebde713861ec82c2f5d9099a89092ff19745988f1ceefa9658cd0ec1f5cdf5f94
z787e4c7422e94ebcc211b60d610d985b552920a1a885f234e093e4f4d5f9e1c53f80124bde637d
zdb0ef49ae74c63b39e4fc4e9715306932ccc9d1bda7d50bcb5376dd3a5a1b611230fd801ab5d9e
z28ea58854c8f27bd8098f43263f45d3e0a31023877dd2f274b19112275eab977edac0308498f80
z5f536f28eb137969215c006e56c92b2935f19bcae926503467bb92d8dfb00833590b962da3b1d7
zdd070bea2184a1dcc115b143b6fd7dccd012322f6dd1688507f70bade90f280f9baa5b7d7ba8dc
z399c1ae10ae1921dbf3017086dd4f235fdc7c66898c195678045602f6163be916eaca4957ce749
z48b1d596ca0173b3626f360539ec780a5df6d4106bff7f5a7790f86fdd6044996f277217e532fa
z3c1bab657bb939d1db51b4dabb74c053f1b7521491f6a00062bbf0ef8a1b15515caabab53a7ec5
z058ef78a359b6ad2bdd3e70883ddb259d742dfb7dd8d545326206cc636f6799fdb499950bee344
ze2df6f5f2f45222c2d59fce4856c6cfb41aac4b0f920cce84982ba2dac41436b87695b6040ac91
z8581590403bcc9ded2fcf86c29ee9160b955330d4397de0d9fee4c3c73b001443344ec7ded2ac6
z133fc01ab335313d9bacfaed51c755b698e2fc66d2bf7bf4d89fe95af8102c60fade092e6c541f
z9f62505775243512f49e7af23c4841982b350cf315d7ebe7bbd330a8f09934e1cdbd2eea6b442c
zc98fa0053c6d975d9ba48f499c18fda89579d3345a98a12b986d54d7c92a46bcc83d611962379f
zc8f21ba9eeb871135a1ba3ef39158750bfe94d3aa54de418c413d5fa39204e21d3f61c90a0e62b
z7340bd44a9d445dff6e1b9c86d2dfc6fa700bbc05258560bf608d4b0f457e0605a7ef3c74b4917
z6ce633766952092d58d9e71b9ab2ac0b08d027f8b7c8d3d9bcb07cba5769dbcb267970c049befc
z6081994221526dd480385faf10d8e7f47b00b5f2e41ca1fa6163cd7bf47d2315e7e249aa493c24
z234bb5f43a82e794a5147b38c6fcd54b16502eba4d8981801442ffef1e773f202eef49d2977978
z6fc00e01cb562330d87fc781d13c6f2bb75028243276b228ae737784c8712a94c6c87690f370a8
zb238ef95da277d87069f7944c0ab1c33df46ddafd8a0eabee4d3122203dee4cd2dc78fd20751d5
z3394893397084507c7417caaf736b1a6329866a173675428c9f98afc1519b6f85c357b93346b5b
z72fda754df36b1198e8dd3f9fc2dd70a438c2527f5c6f04fa6d05418bb6afa3d0f5d718046d69e
zc064701c68cc2d15368614bc7893245ae51eb9768051ba04ee8ea29cb623cd4cf384b8cd0bece8
z3a6ee90adfee074fed8728be2907737ea6ffb6efc6eef3b85122ccf22ef8cc0b1d83280a7a5ca6
z0b7f93551856026fa208f6872683502851cb441b82daacdc01f182d43b912a23ff9037f6185ac7
z3598d9f76400e96c07b4b98820f7482ccfc5267782702f5831452e6ddda10a5a288c69ac773ad1
z84d47a63762722ac7b321dd61abbe1bca7d71073ca9a79a37b75fa1ff308fc500cb2a75dc8ad6f
zb4f833a108413fd5d01065a3aa5cdab58d63ae04b4e3a227decf0d4d5a8ee4e37bb67145ffaa92
z77afb2521c8bfe92ed2bdf24ffc7a5f94095af37a4b3e9fe4c70e4e146d53bb1bdb18cdc9a3b30
z5e26fabcd125e3d052c96fa0e606ebf0a505efd6371347186e30e5d4845a9ae6fc40a68f1d915e
zd814c2131e7de0baaa4c505f151d752b2481e9d6a2ad6da0ef582e53844ec3c4b8b6c1b77a2d56
z8c29815c8e3e1fc9b240f0d84b73f534f9b6730b497385b821f57a0ec114ae2f3095519f53dc0c
z1da31c394b4b3582473ffccfcf3ca6114d6e2d2dd249925f09e2c2fbd7045b67774a6b816f149d
zc25090de46a9291a9a3e785a45650f6b48a6b30463dd94a8a33cb0263a54523fd8cdbfd5a30456
z8d6fd7ed859d8d34c473de0301158fb808a923af1a5e546fc278d65a0ae603e6efc472bf2266fe
zfaa5f19cea88e716572ae5daa457db5d9d197a6b5f34e0f39dd4a52806317164c1d3f82dee2531
z30909cb39efe951f915b347caa46c2829dfaebc84232b867627a2901eda513c454ba89750737bc
zdd3edfcbc5c7dc81f3d4fc95ae82cd77208fc468ab969c5931d85d91117b1c2d7c879e9c180fb1
z5ab9d2dca3d0b56804a0d8174d002519945e8b00c7738c4d82183b1b6e585e1912bd1e4587610f
z3cc15beea7cefbad0a966629931af05b1729ee005c099473cabf5b365d6a5f1a468009fd0a627e
z0b93a4fe4c75d221b9b5fb4199a934a306e8653d0d7bf57d0a9d018708f9e0f121cc5b0651c860
z7a66efb4bb9d4a9c6b8b8d9f38ffbfdf57531bfdbd6ca29ab33c4c62f4970cb440ec1b87a04865
z8da9249ebde30bf79713a2c2a184a668dce5ac58af9c9d49c61c438de9a7fc45af8a5817c5c6e9
zcc7f5f08213173f10ae1d41ef101bb1ed995ab0e475d819a521b2dd4806c0cbb2a7c884d450df3
z0f54833bdf8dbd6eeeebac4e0e8c9bc88e94cb0034412fac31e16d6dd9f4c56e3b7ae44e0a4497
z24b32f83662d9dcad4ed6c026fc7ed3f0c2d168909f908ffdb16e6192adb7fa9a5d2f6eec8a6f4
zf3966c0bececaac0be62aefe66aabd9339d819475401e005b2f77491d0eb6045ec05ea59f3e465
z06ece23765fe8adb3895806226ee1d07f1f702b30873b5d5b8c5719fb04cbb332be968ee1f7e12
z4f79727ea07a7a5afc718bbb523a5dbaeb0e8bee667d7c34473b4c26df994ed485820c33442e6f
z64f71a277f6d15ca52a8d4d3bc4f7e60b81d1f66e79cd2634672eb08af6d0c41f211c011338cbf
z196a78117dbfa90660c594fc324159b6d869f252334b2b3bdfd3bee07f23a983e8dc295810f684
z23554b8cebb139445158c6c392d5a988d0c298d6aecf1e21c2d387beeddca76f4e8952d44ffc69
z4a79cadc4b6b2a4e49b8ac1bd7555d1d6cf95f2d6a0ee473f46a51aaf1e8a0fbd242e96798d6be
zad60d9e9c25537422bda77c238e8f2f8b4c724b42d8d8f44785cdb22706bc5f635ca7341cdf444
zd8c094a8dda50f501ae5e21acd1554b6080f68053cef7f9cd013f0d5ac52a696f9ba8c4fc30c91
zad199639418d8a6df95b7aac36e4d98de6a53e9f7abad8ceee339a0b362992c4e2f47eccef0fc6
zcff43d818cd74bda0eb85eb67dd9b91945bc25a9bd94e2c1ca147c3215e95b2f0bb4266ef1418c
zc4aa65140525714ce4f45f86391561b381514623062040fbb167e88ec546ec4d758789068c9010
z47069761b21d97a3c1ba7183372b9425dba4eec35acaac3d83ac76af4615ab8f9f4944365a539d
zae463cc7be5efe6c7a4a4e99b20730af797fe2ec235325b528f72e3481df2ec655e80906486ae0
z9fcb6ff71b15c7f7c26ff76275f242004c8ba122e65af127e18427a42bf3f5762ea3a471b92f82
zb5b741deb6190caf7a5c838cb8ad36e8ab58c36e6ba3031098446516f4304db2c3071c45392bff
z0163f9afde956b84ef54730c04b02f8aa0b6f74301752cfb17d6d6d05fc76d83be2c83b9e963d9
z46775d4b57b804ccb1a28c4bc66d13c10747432f1ed47d77c3e102336878c0c793843612417a78
z6b77cd3fcd0e913291ebda3dc0651d629e593f5f4ac5e785c2ae5147480060516fa1f319724858
z348490dab7968321919f2b04f0b643653e6cd326bbe3872533ce3654813aa626192b3a9b984b45
ze0d9a2c9a1f66c1126a56890d3d0d680dba3bd1f4a429169e46efd49a4186a6d84fafa126ee348
z9f99e0a8ae87f39245905c87fd723975e074dfaf8f7a23c2411f5a8f0e0a73b39c17443262150f
z489a6133d7b62488282613b1e02693205753d2d86dfc5621c0953339bb72d1c896fce2f53e9cd5
za672e33d9dfadb2ba8036760b5d109f2c7d7ad3e82cc481bbfbf764c6c1272d989e3ca5c15272c
z54f81d00c83c99cedd090a604b68a1491ca9767b7e699a5be1be1d9b6ce755a36aba375bcd7cac
z2b81893a78506448f44ed2bdd5d044969f4488ce281e118cfa9e83560e7128c3b8b3afd58ad574
z18906d169ad69caee4ef3eff12f094379b3c0fafcb591cbc359b2c3c301447ed026d3a1c508472
z44a4e44ec5372604b42f8b754057a140b02969cead62cc9c71f3b5a1e9d3927f38be6b25a9cf38
z041ce6d543825845d2f5236088f91906da313006fb9925db6c94bbfa926ad5bdd4f50b4cda4dcc
zdeaebfaff8c834de04c4919d4b3c78e93f73f7d8a6c994e18f6799fee83f7c6f97cc6fbc3d3487
ze6050b3d41d75f540d3203cbeeff8f0398b8e86766e27f7d41601659d29c0475c797a273182cdf
z5dd025712db046eb4ab0526b335ca6150346c1e29419a2f8e9fcfc1af445186daae19771238b61
zd9a800651bd111ca453084e456978605ad216cf5fc372f934d0eebd0419aed95be5a6f5efd3434
z6907ee387b90094a94756366b18977836efbabc031103be67f5ed4a86115bb99b7e11278f0ebfd
z7d670985d574591467c99e45a0ab25a889aef8c3ab14eec820943d47f1c9dec56a088ef895f2d3
z24ac0841c084f80ca31b7455f897e997022f8b78f3ea16dce750ff792b5d0d9450a457a5c992f3
z050cb913ade7dddf176a8b478ffbe8085a43fa3e750c8dec5fb4c2df098fab21338f1940da39c2
z2dc924590ac8b8b5c7d448d399dd1c0f1559f8e2f3a465a6bade05a3d3e7e3f5296e47e93e83d6
ze3ff93d909caf9fb9ea13d122ab5cd59f7065faaf76e3cd3df58fd585a502a016b1f386e7e665f
z10b346e8e025e1005d6ae9a2566e9fd9643033c76757807de1b13d0d29cfa21ffe8c88ca2e8225
zbb469c30b0d77a7f1e3b4207009a271f5373e44dd3a02a30c7876beeb88b8f929120bb9543d27f
z20140f0d796d1e9d912bc88916ea5f11415d4ec6e0c6e920429185e52299f17ccf2f0c19f8b290
z88275057952b1da1399c7fbb53e3faf7fe9080a461661f094e8d37f7206b3a385ae6b59f2c29a1
zf066bbcf923e6a3885e7f7c75c485da979c59f038be5bc04344efebcabde662f928dc0a81f69b4
z5e2d007682ab598e145d951bc20146097fcb7f7554cbd7545f3d0cec0db6322e9bec0da03408e2
zc55c269e7ded4c351b4dfe2271a45501578fd9586d330ad425c69e56d2ab2fe4150453e24659f0
z70d1d758aee3830a6ec6d05c8da7e8c1b928b5ef3b9b5641496a2729eafed9a168561dff67083a
z4ddefa746ff3c81623be496159dba82577726bf64b00a8cdd77d8b2ba2ca013a6c6fac360794cd
ze27d5125678dee603cb382427dcef976d87cf9e7c49d6d7db9f749ef02187c7d27ad62e2de1670
z54e666f186772624a145bc81ab5fa2bb6579a45767031c38cbc4297b483b95fbacca71dfdc376b
zd2eb96e04fce8c8bfc48a8a848c60d67b799fd58afa57fdc4630d9a591e090a0a8b23fea7ff7a2
z868241abd22aa5d09fe67da78b9259898de3bc2443409898f2e99035a1be42991ff3a3261f0d4e
zc3535bf498b35b5e22df97c9d33c77c2c9261aa2fdca7e8b7a91174e4e04a02b2cc7fd3c8d0f03
zc415e0a7435d5b3d8f3f06d39b20eb5fd42b816262737cc4c80b9bfb9c935a505b82f2a67698fd
z76515dcc775b96cd17150171bfc40029458709f935e13941c23a1733cdaa6d4e640ff1ad806421
z427c6f73357e4f311c22ebf215564dbf5ef2ecbdb177b448de30742c793010a9c71ddc88db74dd
z3c4d44cc073043af0ac19d33f09f1b63ef6c2ae515a38f99d4cef394d31b8d1863a30a98075a8a
z0f9ebb5e806704d178df782faf7a704118e39c1efbe9a6313f1342112b36b5c55ae126cddbaff9
z40162f798932859acf0e805aa4a535ff2dd64c223657e18a3ae548cdb0700557c9efa493610ff4
z6adc5e6851dc96bc9cf42d234d937b56f3aa678f67d72fa719a17e39b10ec9f856baff910662d9
z161f8639533bac261ea0bfca00dd74a73540e6736dbb6f1d3d25f9be98b43e543a206629cf9486
z38491bca233957b640eef8c784dd6eaf7129b8bce3eac909f29e897d35cdb8b62573c93002d454
zf24176009fd667230a649b86c9024da7690a74c9895cbf3ed63352a7cfb733dde72009c5cbdb88
z4ed652ff73945d6dbfc6e8545fc6660ab8c99438df13bcaa10e76935b10ad58a418d2c4bc4a199
zf467fc4fc14579e2853efdd1a7ee82941bfc3d23cc91d81d6ed12b9e311584d77b966718786750
z5971b7ee24ee40d80e8dfbb5993fabe94b34ba3bc33deb13769da39b3a385522915d73f09d5d85
z7b35e2edc5176efdfd92108607169d4925fe61647d0f6fba26e7c1b397927ac253fcfdfe1ae440
z561ea0116752477bd6399b6f1445201d69dff3d6ebb30f549f5c38af4642a05443d0cf4ae26ddb
z1bcda7cee4a0fb3e224bf018baaf2540c20cacc47fde9653f911dfaaa7be920105c8bc08e80b48
z035277b577209052ea3166bed89b97fb565d85abb83faa88474dac9cccb75bced3c7a46d70f088
zfdcffa63a2de8a4ee6321b5c9cb3820798666cf10cb8d065e845ca9e56f3c73e987135c0fad24b
zd9860637c5381c7c2831c35d8e91da9bc5a19dcacd52d0a8cbebe40762e7ab847840fdc3abae5e
zbfc384c322af329b73d2bf448d0e31257a6230f1878735100824ccd931b2b99a57859bcf1cfd1b
zde66b7a7f363860f18624e9aba8a3d569a5ebca47802605264a72b89c97b1227a5d9e6ea26b936
za0cc2c44fbb1d060be06c0f707deddbcd5a8723e255fe41c7bb38ffd77a71fc8c68bf7e42f66fd
z8e88fd6a2d0fa7f570662c2aebbb4151f0334591feb767f7ee6ceb9dee5b760722eb39035b3581
z513d6fac3c8a96971d831ab0cd1538d7e2535df44f89dc4a67c43d21539b28861608c2d0b74377
zd7dcfd71b2224af6838f411b6c4af9ce83c6ad43a445a1dac9a36f6a3b0d6e54c1614f50f0f6c1
z06d689ccfb03f4ff009f3801b795dffa37babbfb4f32d832dc1fa0be8e9ccb1c82e3d18656531d
z6009eb14d613ba20b0001b0da76f8342a437ae2f8e5e93c5fd6aa560aa15c18b3b41366a2f3ae2
z54f76a33681fded2a83a24a3b6da2e6a07876265933feb973822b62d40b3368d8ffd065f08b0c9
zd45c4d5cda3d2aaef07c79cd4587b2cfb21c835b676b44c3012ec0e6b36cdbda98d7678dfecf4b
z35522edf069202989784384f6655d28b579810fb4f0e2353da2476f02d1d8b16da55c82fd377c2
zb9bbe9ecc28db70d2104526e4d78308fbcac2c3e329239e6f695b13ab16fa144a7d27b66a14a70
z371d5ef43ef640240f4ec13df8f3cb712e840e45ee62fce9353ea3e06cc4f6686cc7213b7baf11
z9cc22df3e3aef77d0529900fe362f94e75cb0b9c5019b3039cd72e76f94f8cbad7c3436ec700e1
z0f8dd1f437ec118132712b4195ffdd852659850f5a3137c4c51aa8f5202d8f12349751e44ca64b
z6d7631feb5f23d36cad4fdf7dd5d96a945ee5e7def795c435ef05de6d4eaeb43c10878d24794a0
zbad7e6d2c3d98007abb431c030eee268e6919aea699e772f139f494de1be7891cc6089ac4c4476
z70bec3e4bbdd02285dcda7c9c1c305263d4fbbdbb4ac07828a1ff0b7b71126687683219bccb5e6
z28f45992281439e533d91cc25cb71fb620f31baee01875f79d67ca5bc263026dc609b4df36234c
z4f5ab1249987d462415131420c4b8d938128fca77145e6edbaae8d8c2949dcaa46f5c315fc5c08
ze565b90c06b8fc67ac67b90518dd27b6c47cba32da2283d289d09170f75d1a0ae13810897bc2d8
z1ec3dacd64e3a10e61efd730f9799453dbc1f06d33d013ca8d1dbd53d7349e132d93b78e9928a4
z4e7045668320ff5420141f403bb12d4995db357d3628ad91f4cc4f760a141b8de98e1f4275f4d7
zf4e6f1ceedb770da968222f5f3b1cea26a09c316f484dc1209f626600c0d7829245015acb6f671
z3c1584bfc906a2db19a44dc2dc56fbed06a6edffdda62b392a4d76c71f069d0084c0b9e6ad8ac6
z7e1598dc95485ae893306506d7f43af9a7991d72b3790318dba7099785d79e63d1908ae28c4c8a
za6f42289d6e7b58e20a0f37f80a05d401005dd0e3b59749773f85b7434efd5a212bded94cccc28
z79b4c5c3a9e08b7e57cd3aff7751cce40c8830e22b142451aca98cbcb4429dc4345995ad7dc7cb
zeefd64eae241118741b4ade33d977f50827d60ec6700d0dadceddad542389bc507314e35f01b71
z2fb10676c80906b1cb547535d44342b6dcd227a69b0c5dcb633834d861d4922a4741bdbb23befc
zd52fd08052e6c1ab1f4a69bed2bb58d1a6ab1dd3a7f894bd6aab2b22172f643b2e262402cab446
z3279acd36ecfddf0d9efd29b9bf9c949c279c89b148b81058f88109daf21ff430527f8c7b4115a
zb2e67cdbc30d5c73d3e21b33d1736106d60b14d3a28ae5ddb71dd853d0cb31ee855a325770c94f
z9202a088ec4749b3c0bd667b5716f45ea2064698512e7a258e3edc7ec2073f628cfa5d10ba9bc7
zce00e75ecb54734230b06de7d8806e0676b832eb3bb9f3441cc808be04829456a5a725c1098a17
z871523e1d1e8160069159b609f14cd4c2e1ae783615e711b0dcac4eaa736c0a81845ce4837593a
z750cb9726926c839fbff7f1ffa834e7179be5188368b3f13abd92f269636dcb995790a768c6284
z983ccf182b1f08347a48305e8a206a24579895b485ca257797ea6cbf0806ff702ae09e682ad08b
z386542c760140b3ae5802418f9f54808a857574f91919679384f702736408db42c5c48823ad0c2
z20292cfa9229e00029795109c4176a788bf8c23e27cd18b38b58d65632136ebade9ffd150fc9d5
z9dbb464756c9b4c6d3e3f6132a06520e771e550760b5e3a44f30beccec7a25d950600e1e238ba3
z0c5f5121afef85885cc27d4cc9d3f2bece2f0b645f51c54b9005f2739cf31acc9c4d6e8d391945
zf6f2722ac4874fa533f0f12b964ae1d7e1f275e253e7ffeddb280d60233ebd58bc8d77342a2270
za503ecf9b0d61e2e72efb8083c149942eb3a351db75f0e52c80bc4ce7d987eaa7bd51c2b5708ec
z99765dc803b26383eedfca18e6db8da048e194e769c5514b99f2856c135bf96e83a05247796820
z3b683d06dcf1e996a3acf69bab89a280a973381cad491f824177feffa661e024f2fca9a4231e5b
za158ef379735c7fa2d307c7397566a93497fcd2264c471b8f1a3c765f2229e01658d271ba91b18
z280099c8de53b9ac337be4953692ad7719a6a02ef948fe64c2680c452b915c25d60cb55840e1ca
z546d1c6a7015d1d7d7aaadfaacc56d45fbd98f23054ba74d05484c1be728d28690bc6db05d7f64
z40f1d569b0eef4dce2ad5cdfe0981665402113a88f440e0feb993edda1fef4afa358e3bae3560d
ze125a91c3e5adf26c07da7276e5fbf298f20eb93b667785ea732ecdd56b478583335c7476eaf6b
zf9b101def49dcbee160f5f25a99ac842a3c2b978b4eaf35b5fa1e93ac8ed33548c81bd0621ded4
z7bb0cfb24b52c82b28592030643aa85ca3e5da831ddf953c7932905faeffa3143be967d90238cc
z65f154ea1bb5567ba205792b1260a8bd4da69e573b49aa54e5253b8c0434d4761c3ebd39ae2554
z756e660b04979e09d44a0f0b0551cd2b5bbcf03f1c7727be8cf52bf7f01b861c2d9346d61d7241
z72f286efe3e56df2e39479ca155da188446676b8e3249334e5f081c3594fdddc55f232fb8726bd
z408b9ce3d969c444b58622510d2af8d25ce24af64fede5cc0b530a7a4ff5ffa1ab50226bf7ee0f
z7a35800923b7a6976035be3c6e66df127b6556c4db5d8213805b66c50ac1c29e2d5fdcc7ef9c68
z6fc0258a6f64f39c1cf7576ad0c730c565ba0a3f235d327cf2a403601ebec26e5f7f3cb0fbdcbc
z62967b5413ed88240c47eb6f092be05feb28ba11029eaf9a83a66fbfa0a869b7d516c09c296630
z255d35aeeba4dda0a781fb1c673f248fb2bb26b909acc214e1119d72cc5ec505b8d3ba8af6f100
z80448a5810e1132428f7a623bec1992a721bd2a2714c58f6e4fbeb6bdc530621ddf2fd5d39fd46
z33ddeb934717c0eacc0d9aa8c3a7464fbd64f75f46fd84fad1b3376e65a0107f60a9a839a0c796
zf056af846907d6c3fbe97958aa23391b973e1a3b7264dd4b266afc428809c29fd2da1bdfa163d7
z4588f921780680311a3d6a45f0089c171cf5ac1615d2b74f5395e5d5c2b63e5c2db98b02e3fb3e
zbf00b877e6251b3c755c77a6373d77c64aacaabfc7aaea07a74ba2752ef2516eb5f47d603ea629
z0e996403e0a93d9799a966acf7ad1ddb7cefc828e4ee1be3aaac388fb4acb33530dd191ae814e1
zd24f7f7ebdcaaef02e0ee0672ee3e85298eda514bcc47f57dce107e5d190c00efa1b249227be6d
z7d3392b8f0e9062ea4ebd8931425b5130c0fe6bedbc8b1b67a816c63480f10f8411aabf6175bf3
z3970e403c47c37d225bee254cca10527bdd8d4b9ba5ad48c763bfd9ac78d2ec4905e461554068e
zd6cbc609e978448f1785bce92d42cdc4484e873ce82913fbb0b1163526b1eea3f8144cb4ddafb1
z61f695941cb85418b02bce0734836a4ab0acc4d896a887ba0d7adfedf9ecda77af500866c5c3b0
z29d559b2b5f1e6a0243d584c8a5908c09d632f0a3b9561f418f5a1852cdbb91569401b6d2b3bc2
z2c264ce0ef1bba24a5c47d211f68e217a6e7a448588e271431aada4f54ef9479aa90661476678d
za8d67b9e5e545a7e4528d5fe3e767fda0e826410ac2576b10c52f480614db80b2e03a65db031c9
za73490ff0a219161d02d39d9860d56a85906ef74b76ddf5f1bd98e447381b3402faf31bf18d940
za02ee0e805d385a13420f8867383e7ba77518701e483db8fb5491b25a3446988d1405fb43de9c1
z692242e46ee8b7a46cecae7be5b238b2d9fdf7bfb22626c908c362a6e4d123cf2164d810f205bf
z063d028c74f7d78c9cf29568166b5038b4357c2b71e8cd45473f60051e188479a5524bbfd84cdf
z03e8086826e9016d9dd9a70506342b90516e37c97260655b4f030f0daab7416364d20a25f0dcac
ze7e2ef0344707e5c6539a98749335cfce783e4ec8b33ff72f2a7388fd1dabdc4968e8ca7743724
z1f972e8a9f6cd6287814f56648ddf4bde64a028436f96835594b2f29b168f351a9fb0f5e6e83ec
zbb83e22f41581257434bef42d5f38b7e668a1f07b0233da7d1bac650e945b4222100334d134bb8
z6fb13b75f78de7e7c91bd2103cb75d5902c00d7e23040bc2903cc92cd94577ae8f7aa53a43b5f1
zd31b7d77cc2c11dac084a823a7b7e9fa666d382f2772a9f483e84611c5435d67a3b357093a378e
z568e7247f0792ef3412fb8f86b618117b4aaee2fac96b7be468e4049e38afa380a132c5f0bb0f3
zd23339fe82f42a94b8590d682e70259d9a41c193cc15cb6562b8297f34e3e57724df6867615ffd
ze9bde579a18ef0213320525d23b79d7abe211ddb9a6e59738755341dffe32a6acfb8fcf8769001
z8ce201bcdde6c935b38d944431619dba6a16cf5b26539ac09371c3b9b0bd2f919d06801dc9dadb
za09a4eea59d16faced4e2551854927326a6ca89d0ec53896ba5a407e7ea2d721416c8666b97dec
zf61edb2fac4e7922017bb7ffbdf82105924e88e972b532d855945cc90ceed93d60b70795f17993
z5b5956b756311812678c7f69f99bc3a5a55d5704df0e8cedfd6f86192935a6b7a55bef34f837ef
z9bf8ff0b3feaef1cf3088c29e40552db7d71a30a01111b034be303cc4a77927ac718221c4c8fd2
z1f2019819ebeb78b35dd93d2a644e4fdc4466f1818723350d040d01bae905abc6b4f8ff66f0f77
zc3009ef87cd41a5c92c32e8a2362ffe8fc7b229c1927558e63750f8b000f123a9ce2430f21d65c
zad134bc8d85ddf94c84135b8664d021fbdb03a964edbdab6ec341bed76a553548f8b8c93a4c56b
z21a498744e9803f7ba49db6af8517eef037d775d50f82caaa7a08b201e6eccd3cd2a723843e2a7
z69013d31a1ca752c60c0e3b287ae2fcea52a7394c9c975b3fa6eb840cc638268ef978e33ec362b
z31da96c7295538281d2ccfbb5dfea4bc87fd72edd63232a2a1f7a441ef0707e252584ec340e710
zf326589dc9c4d50306eea9154f18f2428e87039500d46991c0413995dc1366337086671d5173bf
z4f231aa207e22d2c4302edb525fafafbdb49f53e4fbcd018a403e544873ea2a9dd2f31bbfe6ac7
z59b37e4bbcfa65ff63942a04b9bf9ddc306f8a741fa15806447b0313602cc5b803628d19d21c7d
z15bc69392d698679c02d777eceabdc1c95ece2b34d1aafd5ab2c8ef794c4ab6aecc0f15ad139b3
z385f3f586da3cf98f65366a605d345a5b3a461ffe83c6adac306d8a7b1a17dd7922ba47f8ec94d
z33b74bb2ec1e6abc3dc000b1fec7f6a51ed3abd8e17a1dd521f974671120efee47997647c38262
zd6b4cd997279a7b80e3232877501f83374f91cec3bff589a548d08b80b2f920924c78ac87a81f2
z130f0f14a59b9b7a469758ea7973b5ae0b7c14c76e9f39abeb8995de0889876d48219b3ffa5389
zb7aef580d0bb167819ddea640fbade9fba3fe0156b840790b2f2c8bc4012ff37e45b23edec0cbb
z3a4b757c3ef0277bd6fe5dbf2c92387dd2e15fed23386ec638a015ebf4741c135fc0739574ea63
z39b81ed21fa29d0a99abad683fcd1c5e7e2601a563a9b50a74452298a5a52d39fc9ee2042290a4
z59dc1342418cdbb2dfbcd0c4dcc6fbd6e43ceb68d523fb3864ae74c88fce0d41951f807b1779b8
zfaa67eaeb6a856d19568a50721448da93d500b8ce032508cdc820613729cfb27e0f7e5ebf4da90
z39451c43567036d7e0117d7c6a392d6da48845a4ebc0bbfebeb199f2f60f880f614c0795c3584f
z901c6381c2e4c7ff95df863fae61e95240ed7a4359ce0b64e6808464384ea652c52abb76ce893f
z9720b54a03bdc1b9266fe173c92d51232fe56d941fff4330844d9417d746338b64b28328547805
zfd22b18fdd5fa276f445e1d3fb570dab93893100e858688147b35009f1703b718ea855660bcdf5
zc969b5aea67adaefb2d165d8ff6c58b63cec18d75ef911245f808fc7a07356e3d1bee74c13f8d9
z1886969650da091b7db77de22a953c8b218e04cba40e91ab6f50d9904b35c9e3a5de9b3839409a
z94a3af64ec9fc7aed43448b6e26f1bb0983c5abf369789677253d8e726f7f9cdd60c07dad02021
zf91ff91f6c64d4c0e5f9fc14562825641c751d083cee5b759ea4a54ee27a99c0ef605859742971
z1ee629fe609ab0101d4995e3d544d2deab87b06b63652c04d2ca57c31e2dddef38b8476b8083e1
z7966da915538b1298b99c4eba89dcf5440758d28623c4de87d0a4d75b61af4bb2ddea0bc230269
za33738dc92256b817a9d0f306c135a87a4562c7e8ee4244eb894422c3626c3d6aa37a368af9e72
za7041a0454557bac3f064ba27551cc9726e243fab7c09933b6b5621134f98269620e76cb7daf56
z0b503a8ff3b1e5bc80f856e71a9fd71c0179bcb8d0c9f3006a56d4a8d3acf434413f90ca7a3956
zec71a7ef4b6ec288974b65fa1c2e6b5a758249690519d8129490ba6800d1d996ebeb99eac25b50
z03fb8b0f35db0b17698c11840800e8e90c691a7077aee8162195ac43ef5a6183de50be5cfec75d
z6cd2b047eef8cbadcc8c12d2b66b256f9b9764310740585e0a2bce69c1e185baf3e4a143814b56
z9d4c168f587755d72f9021004b716dbe058296319e38d2a6af7561b8ac59d5d5359cdf8bc105d1
z00753f9d0514966b5d8294537fe5302d79aa79a8739ccf379c004e5c1d4f47551f92e43bb513fe
z9e8686bd26595dd162382e85fe6aefb887f003d678b5433e45fc9d3b5726cc4d6be076532c506b
zcb3ced23266852c7e8876664004c61d74f35a9629dedab7b269079971f94515718af28615875b1
z2418e292792934455238f55d170d2ca64db00213c23cf2619cb48cad877955da1bce9e05c8e478
z2f38d0f10b7fe679a47fa6165da81e0898cc7b5c01b0c6d6e608354d99d8de6b449f48adae3280
z5c8dee2545d4a2e6d6b94eb43a590ff76b78eb452c5aae0a088b22e5a72f2d71d46857a8ff2d6f
zed9538aea010012d04ad3028b509ea543cf02d33ea7d27ef4190de095e96fa8496ee26a4903c85
zdabab65f5f3cf86163d54e3f050549424bd109f77e7df4a8ae9fb3438824b4551d07d0e3bb9e29
z2036c2b6f9c6a29d92b78c5e53e76652cf68787c76dea306337e0b77aea73625e1b2c18a010c5b
z0099d05f98965d067170c9df8a91b6b07789f17b357689ea16adee5e19e5328b2ce4d008c7b9c1
z29f0576c432a4d8398dd4eea3bd48824e10fb5471f3e1d6be42d148aec3fe032e10905cdd9d214
z195f998241887ca36ac7c6d59afe72020a5425cc5202dcc9728de76440cb9dffdf0cc6adf3f2a0
zf312bfbb56a0017df71ca881449c3948e0d555e204f38ee1bad19643a1489d4537eed9126404f4
za09e4ba1289bf40949d42fb14be19ca2df28ae4723676bb4b20b4aa6ae323dacef5fa3a89e617e
z082a81d5dba3d32a50ee799752cc84ae7099bbacbcfe4de40b7c026d52eabcfeb4a812efa834ac
zfc9f27166df98cfd8dbdd9ddd2583f36f35c674717cfc9fe0bc23ae92e3f5ab5b6163b0521d228
z4be954f056532c9198c67e2c38b8f1e3be23c14d7de427106dac1c0ca3a0757d28bea3cf2fa828
zb5d8793c41f45975238dd569d4774e88059e8962e77f90010d7dc7ca97c58eee310c35c36c6ee2
z83bf64b37ebd1b4eec726c995ded5f9f2cbd97c41f82e70552083b3c310890087c727f8c2e7d86
zd01b75a2cc144f7e2e9add82493db2bd45f6e37f1e7aa403c95118d4d951e286f10dbf191bdc7e
zf5bf07b5fdff49e535b338d2e5f1a6497494bd21d8bfaf74a87c75872228f2ae608f620d6fffdf
zce59b01d2b10a51eb691d67fa8abd56c7f45a5835e7f2ce3bc5858bcb53180fca52a78c1226f3d
z158e3b20424750fa1474ae97ed0b391d60e771e67f4c78ea45c36a7f80a43491c5be924c59f960
zf4e71fb6d6a574548b8c01bcf7514187bf49885960c022cb58050e59567da0610a46c366158ac3
z307b566f1159bf58e6a1f886a3823cf0fe7332c74e3b8a6ed765e76b34ca7fdcfae7161df572be
ze8e9ceea7036b173a89147b2801d95ae452c8e2f4c73b029961a28744b771510b02514c0d9a483
z6c3e24e42f3e93c607694f19b89fbd95355aedee75160a50fe7271423983c2247ef712a5763ad8
z00c777fc125f348ca86e4763a6673bb7a0c592a748f96d3ca622e9e56b06bd15eb52d6e917a89e
zbab8c4147e8e1cc6a183317e3e6431bf7458a5dea5c806b6d5eb9db38791c5d00c91d00c01faa3
z2a40ea29788b57eaf438ff96e894ccb1a5e9153b56d126ce8400f8a86a1a796e6e65795b570fd5
za187893fd46a858982179aee80f1ab56182366a9d114e2da9e5473574f58abd136635566bb57ea
z8c802c780d87f082f9d4ce6ca1f09bf1c496c5e57d0d01a3530a5dad873bb5d9b3f637549a620d
z6a6c1814a86efbeabd5a00c4e7afed4d6ff957ccf9dc98c48b30658c71ef20e81e50729e8037ba
zad28d1d09f8b95a76036a32b717fc6f4adae657ba24cba632012682743a3e76a1f096cc5bd7a3b
z2863431fa6be9b3cc65ae143c32bd0db848fc257407bcb6064ec65893b96c3a2064256d00ac5c9
z71c32afdd0f5101e16210f3eabc03df88cf301bdf78497fec7045a126856c6f034e195f39483dd
z748556b6827cf1a0b5913ab44bd10a25db002584777e1b3f995ea11387d62e74630a825dcc71e6
z86d7616c8c70f157e41ba86167575aa7c8b7dc3eb439c21f412a7c78abde5835110f1ab2d5b585
z38f1dd72c02a8095282f9931c764878b19bc51c9a773c19872355e6b18731e06b4f6de16a15f4e
zb6b26d887bbf666e6f1fda6deef2e15260bfb4597a6bf1b1fc8f64ad543a056aa3acb9e75baa29
zb5576b0c1b7f6005fd08d439000e7d48741d6a7d1f16179ddf0980b9e971febda93ea50e7e0f7e
zaae61e33aaf19d44af09e143973df4c026ee31aade33d0a53a8bcc9b19fcc0fcfdb78a3626e449
z610836dfefead32fa6abd414b1f80276568da4c7f1b7a29650886052a2cfc6858664c8511347e5
z9582620e16bce5a118203495f47da3aa239cd727c89acd4736f337b09c04b213e6b973bf062053
z2199e66bfd09352ab6dec8eeaddd5f8b70b3cf6df698383adb0484b3efef632d21d36d6e1e6735
z6defb9d8f0c8c311b836bdf5138fee753d8d72faa6636d435d2efd7879cc673df135b9e1798682
z23bc32d51f6ddec03b0dc8b258146514548051081e24a47ca2630fb60242ed27d43fa1c3228d17
z78afd1ead618f999188696eaae82dec62d3d71746d5652e2fc96dbae1b342d73e0741e457d14bb
zf55e3d5d5079cdfb553e73d299e4a058dc91f0572ca5798f1100361b7b26f7e46b60dacd05c844
z237d5f9d4cd41e60db800f8d73ecabf770a8674cf44fce9b751dcc8fa9d7d5c2e160bd04888a62
z0711784827fcdff295a3a995969a4af9c69877a0c039ba4e926fd82d0e6cb0a93340e1e5113c22
zea4ecfb4bccd3949d14fb91c61a7e120d86032475b750df0adcfa2248f4eae1cf997c03a71cd22
z47a6dd0f4e77fe29b455449c127fe2ed2a4357b0ecd2a069bd1f7d30c146fb06feb6a0b2d31647
za18130407dd7d339024447ca552a6ddba00c66f4df5558fda8020ceee166658d0e02beeb8d495a
z05cd593733b5ef2e5e6eed6e31ac831494522a90da648289413c2420b902838a0e63e9b43a2f8d
z8daf1cfa95b4536b21e1bf50d2f73b9749e2103a4298b34e1a85a3fe503a0c6d0bf15fdf8560c9
z0fd7c3fca479e7ae227dc59aef7bf09edcf4958f16391a8e344c1cf98b405ac4094a198c524971
zcd110fcfec50ba293ac0ada26232efd278765d0ca04bf7d3b43e1c6ac3914046d0537f9449ba86
z627e76c38dc1530e1010024b2097c82045c862b907ad007bd669fda1399a9215a369d355eeb6d1
z64e9ab5bb2aa9c97ba645372159a13164815d8186e5dbdde7a213042650f3dae143fbc12cbfce7
z6b24ff465c066ddbe9e132f549a377e0db7be623319c3ea5f4f1e54a13c631accc029e9851dabf
z7c4c62edd4280b0881ca08f2c9ba3068ab1e38c0254963e35e0a993e193194c4dc93ba14f7e89f
zbe51745a6fb2d2e697be83b2d7100f44ee6678c6af75f4207e423182294fc5d1154de660666053
z230e0c849b87f7d50f41dc00db70abd6fae5314e56c137947e9407cdf56900449e97a3871e24c8
zd87fe54796804338603f58322b234423715c2c193142d2632998ef59971814e3cc5099a83173de
z8f13c4bed20329998edfdc0b46f181f9396f20bfbf01831f64bbeacae6b36893955c28f73b7432
z2f69d5b3c5918e9cd172b3d989fb44e370c3a5ae5d30e0d063179461c09442a1ff113d06f73a71
z2b6a2162bf963de7e1c28a3ab45a55b0449269db5c2fb51a52ac62d59cbd612071d358f3cdf964
z778b04268f160aca55582826114f26f9f871142c3a4c67d4406c38083f05c08dd7fd8d9250649e
z8ded960a278dbf7fc27158a35ecd8acacd5bee940cbf39764ea83287bc44b70cbee21c424e2163
z7b44ebd95505b0b0558500adb79c81244a644889e404863ef96beeb8e1e786c9c8276e9423a4b0
zbe024f773940da400921e768bcbf4cd1f83ca7baf001db8f45a97545014dcbf8390b93fa0337af
z25b9da4b202b5a379688a5d27451d9a4e51055c7f235791727d56debb99b0ecae6170cd18ca8e9
z8ba872eb64e79c2b144390bbd49cd321298902ebdf584a981b8b09027bb1f9cf4ebab93ee652fe
z2094247be2c477ce5e46890b51dccad15e48d13e2c354d10c9e402cddf3f4ef97559bcfc6889b4
zfa2554ec0d266ec32992a741f7a104a02943fa357c1c0b2fb8cc64e38806ac2de14bc26564fab1
zfe258dc67a47bc56d0dea8702af114f125c71e83eeaae1c501d24ffaf8327dd084de61d1d598da
z3a8f58b5e955fb970c1997940fdd048596fbd04fd3e5cef1887e725f7b073cdb38aed60f6e9dd2
z4a72c9970a4e992d5adbb24c18e7db0a8709985abdd9dcf2c10c7969c5e3ed4a07141d9505c986
z8bd547049bedf5d972e1f62c061807a0a5b63432b5326f98f7c28b88f35c70d4b3e7d5b9672384
z7486e33925285cd0c37f0434d08d2e9c8d58bd6e66335360aafc16c71f319521a0b952e4f5884d
z1475f27d3658f2485a1450d88422f1be33ced53c3d816e750f2135ac88642fa7b43c045c66def0
z7a755a02fd93cbfe77bd80e7bc19a248f03a4c4d0547324e6d58755b9b552eeac571395963478a
z6840074adf62ebebe27505c1611e040963e92cc09f1a0d4bf6c182adba1a205be8ac4cb65aeb6c
z6f3d44d6db651a6c88c1ff5c580a0f3e0075862a6faf3535334206bf8b44ce7d2e48b62251d998
z0bc2727037c28de5911f4937267ea3ed1544841205598dac5525e4feb4a2ab1683bea4abde74b8
z824b244006e90ca55605cf8db54ab9ed62ae5185192585785e16c2dc2b3bac4fc1eae0c2084d43
z44d4082bc3b29bf1fbceb313c0b1bef503c4bda71d4ed6eea35a45c7d49b6ee439edd4d9b057f3
z68e0e72929576c120e3a1b5a3a6d9d5dbec2c16f530db314c51e91f58fb977cadfa32d96b03b59
z63cbe2f6d862654d567f1fa600f97643cf081feeed8abdbddabe1500d8c704a4b512e6e015fff2
zca76e64ccc6a61d41e50e08a28e17a5b30ffbfe26667cc4ccbe541f8e518e55ca11082fa836d3c
zdad9e1eea6b2a6e6b9fc47046c04a889f8cea90f9f49cb9be0ef3432fa88694d7330ea4d4f99f5
z55bb8f0669f13c4fdaf1494d14484feb3f3f66e06afa969f7d302fad0b79a9c7f5daffe409e6dc
z0298b47c433ba1565a9457ea05c15cf6125ffe8998842d1f81de5817cf5595439c11843e1e0b4c
z931f6fbbef214bbbd2503d102da482e397e504767d93212da1672039479ef8ad6f9f56946af620
z643496c27421d2abf8ede7a820d34488ff7f8d027121d3cfdd8852fe66e2d9442ae016c4ea69fe
zf44210705e3a260368dc0a1acfcb40d2e57fbe2715b6617458061c3cb4dbe2912ebca31c594234
ze8d871115d93356064b75844647a7b744901294826e61f246c05f12f0b9faea6d6a415d5f3e57f
zac82e945c1b395405470b693bbf1c218233678696751fecc1490b10175301c24bf3c03b0565934
z44a744f59bdc85093045b513a23707c19fa925adfc0c974c1b43c3e8e1c5cb150fd00014e7c179
z4e5f5e11f52d1829bb99ffd8729b7dbfce350696a9ee046c3cbca29fc7edab4e32ed1472a184cf
z0856dd7968990dce5f4d440a45f0b33283b30fff43cbe57c545551ab94c01bb87ca165db7f6b0f
z5f99c72d6a2b158b248685fb17e5696caaa39e4226b821b15a5b74ef88aa334c3ef45bfb4bdf03
z805404474d997034de327b745dc9fc827e99e768cb40337e285b74255900d56849d05ce796d367
z41481b5db06538b95fae68dc27fdd59cd36a76300c70a5dc1e10d09202a6dca29d3a064d79f7bd
z574b41b88ed72dd49d31bc7c4fe6fe32c67c73116607300c6aea8ee4ace33a8a4a7e5033acd754
z6f5946462c00993ed63a6d07f4b319fa5687cc09806746dd2aadc3a278aee6b68d1d97f4ae4e7b
zd59f719ee83a78acfa0f850a09ec1ed1e96b57e73883a8010377a4f6cbba9d0bf465c0ebad0eda
z42a5a90a0694ff6c5b5a2af75b57b2347c73272e1d9a8bf61699d9d715a7a1a8f8cd144795939b
z24c1e01a91007985b795a826c5f903750dec0845ae52e27ce6fd151f4a2aa1dc189f78f91db03c
zf9a86f0469e4137b693471ebf5570119d126725ddb8f5396a378e6456d12290855bbfcf420db98
z04ad63aba81ee2a77ad104cc7dc0baa2107a72b02fa1efbfeec8d00984cb24f900640eab233638
z320e39326fdbc2dde64125e18e4c2bca4ebebab5b37fc4a941b21ad6a36e930d586dd95c305bd2
z9b817a6d20ec4307829f8c1272ce69657bdf72098e3dada08b547bfeb9c05bfb07d8365ec59e91
za458f2754e4723d0f8a8f683fe57f9c4c3df82a94b16b1d247c58a32daf509a7add1e59fdf463d
zd295152fac3c007e5ed6911a50fb9ea52e84ae2ed997d0a0d7ada8698aa02df09c4d66866cab66
z964c69bc593e893861b6f90f7a864532f0a6d97583573b7f294f3611ced351ac4ea2153b08335a
zb89b21f0aea814ccfd900ae17b2a06ff02b5a5d09f1833404a51ba58e225d04fa6a19626d6300b
z2a4a8a4070f9e1a8e9dbd9f68b990685808c7cd16014829c42ad1582c92be03a3e54b9acdd6445
z3f4c217ee2220812198889f395beb06ffa08978b573c28b14ee7ca8cc090b84db3ab479e73e575
z23ba1a191e006d3c7c227a6c068f34d17837f6a2e08f321d58d0d4b238d4cc22fdd8b04212268d
zac5414c040179516e93db07e11f6cc42d1aa80ad4ecc1c29b6b01565ac4d640bddb07a2e92ff03
z4a401df36ade36c3ca37603011f24fbff195f26f46fdb65e3ca3e7c651667bc055fbb2452a71b1
z460e2cd13e2db3f5527f41779e272fbd7caf6ec0c404f025085430aa2c54769d1e3e23bfe6af3d
zf76c9e63570d02c49e29ea5866c751d0611299dc4a511d500f29e080ecf413e7d098b6bfcba314
ze646cb3ea51e6b4b73c4485cbc5492c90af7cdea61ef73401a6a4d8a2ba04eb0e3de3700bf9725
z8f6bde0ce15b220f3b821c499fc298a5361d94d8991e4b7b0b0e856a2ca9930e27021b092ea6e9
z4efa692944f5892ba7eae8c310fa4a360fe2a8659f1641bea1e4a6265672e1ab764f3ef6c0c242
z82a62e4ebb78133d50af1f912e0af363eeecafaf90add280b13e07617436a15ace037b5f930082
ze07df11178790819a3fcaf941ae491fceda9b3654bd1426368cdcdf4547debf9a955ffc677d3f2
zc5f56358f9cc72fb9895428c4f180c205ad04ebaf7fa58da03060542a919fdf27efb585b37e436
ze5e76dbd7383950f4558e20b316e074fe56aa533118a6cd93d20a33bf5bb6e78c73e1ae95a1b69
z04ed8c6280fc70c32d6ffeab31f9b297e3d5fc1779060018f5463163e7e3a3acf0338d95dddae1
za48e0d3fcf5e07b40f49c7fe653e2a4d0a98c9f1f4da2629d3d5b71684474291634f81fff77f28
zfd266189607a8933a78cbd63feafb28c703df2f04c2959cc4437231534ae8c62adb3dc8c588809
zdd0fbad334877a32bfd0c916d1d737e7f555e81d57573ce97f1e63444f1311c0d0f71ae23c6127
zb8e5a29c6ec2b538dfd96b76431595457511b0eddffd3e3d749e00f2144a2e6ec48a8015dd85ae
z8dc42fbe1844f5a1cfc862973d6fcc8483ac26d22bb7d5bdce2b1918f7405cd8183093b984c5df
z6d6b4f7d079d88306e329459feebcac5082f63993e6061427740de9be019fb2870d770e2eed6d3
z30718c7b85c2438e8774d583963dd3f7bdcada9e614d02022aa292880bc0af0f389e9825b3cdc6
z92919f7310548e8754fec8170f373c06e35bd829861d6c0d5836d719090e619cda7df8e123736f
z3cb9fff5d33f94002ef0642a3fa12c398280cda8b3271d2b8370bcfa0388b4db797d06853d104e
z2e8954c58cc8810494caac6725dc4d81cbc1f00657cc091941aa4a5b3c847826a01519cfe07f85
zb95b0d915ce85d096decefa66b5f9b196b1ef0e322d77cb156adfceeb57d4e73cf516ed648e53f
z2e72b520fe067459dd41fb29897a09709d5ec1b6cb21d1a43137cdb3e97e39e6e6ae90b1321dfd
zf347c249a7d404336a81bbf4564e401cef839533c93aa25e69c070dc10586b00f2963926fef61e
ze16a4571b0c86d4d783f6b935cae37122cbbe1c503d40a23e15a1b4e17a5b4e5d01194f311d49f
z6bbf8563afddcad007d3f4ad029af28139d053729d60797ab7bcf4ceec117b9ed8184a3226eed9
zfde188f8b68dbc84de9aef1d95bdd9654e7906ee9a64bdbbdffadc054166b576842e5246ad5673
z821a71835bf641291cd44df62e388785772b1cfd0a2a3a246a84862a24fb2bcd935bb24470bc91
z2a3ec50f87e7320f71cb39d149bd8844cc6152a8703f5ad640999b8d3394dd4de2d73d608baf51
z735a2521e58278e5ced1da8554ab16fadc4bbc0a43d20fdb58231e4fc4beb71b607f7594554571
z38f4d45750a66646374911cb16cd45adc0b41c5f071bdcf162a2506b0fcbd66c278ba882bf1c09
z1454ff36062235f0cfd0b95add8083fb91e36f544752bbfa70855f34e0d54135b3104945fee716
z482d01255b2016744cb7a5aa7fd28d0a371f6347b408450d7b323da3d3431a9417dfc3b478b5b2
z19147c56f8160fd3d04ff360b1fa3ee2b44c5e2c7ef716efa0d257d8765374cd70241c47410831
za6f04a515acd7d019d95af57a6f87d1f7440df0cdf4efca6a84d47bc9435c7293f36c682c78563
zf4d8f310f852f3d1de0f632442efc4fae146279ff1f5029474d2a0481bab94acdfcf8ec82a4fb5
z928b3cacb9da8611870635981022bf2c264cdb782e32b669c91900d39aa594f62ad149401b0bee
z335af50f2df658e2e04cb05c0e0a1fce1c45c7c4d20b6ea11e149d9a5c313781b81b6d3b199c80
z0d26b568542dd6504135c98dd168d6d6184c91b14b6b372be3940de60c17e1208c182f9cce5b57
z1b3ade4602119f85c672065e9c6bc149826753d0a948f88d2c3d5b85dc3aa61e4628f7d8da1b1a
zde33e0bbb656ead59c967effb776d6039300a5c6fe0eeaac11e991a4d8c4b9cbecad5499522c4e
zcac5ce722d35ada12953e6db4c1ada501a07d68166dbb294c04a73e830e3fbcf0b6cbfa986455a
z1beb481d7d73c966462d2121b526db7f4e1311ed89c27743b9fa062b85f1a493619c9e67015fd9
zfe4f8e4c1e51879f022fd6f7c53d679aa225d07e33f97eb20bb21e62a7a3d6e17a1b53e13afb2e
zb617a187620f1d111145649479537e63a2bd35bf79576b0ea44580e6ef865607a008eae0ba4706
zd519aa3bf203913323139499c556662b57108ea94c7029776936e1bdb29fb0265a351b11cb3a1f
z62d986aeed0f836b5b6957ddbead7ae9c69ee7bbfe24eb260febb50c1a04f0f83036c8f446b5f6
zae8389aa54d6c791752c539289a9948ef4624d4fa2dfd2538c6d956c6bb9771799c015d804958c
z79db4d13ca787f32b3993bb1b2f3beb4fc7af5f6df6c948b651bcf034a6a76bbe7648023e632e8
z22a0897df4d8b388380f094da566aa071d7864a6454d2f12ddf694f66bad71e15c6b02ab678326
z6578cbbf0573ace7ea26d746f3a41e62f19d0530dd0345a3d9951468599a75f9b011bf3d1e0653
z13b74bf5a7171028f142cbdc3976d2a679502b1ea2b952f19019be03680a6a4e28a90b82a46eb0
z1a06a9ae1e7faa04870e1254138efa88eb789c58d8e1bd36cb8fc77e6d335780ebc6cebc07d030
zb819a6d04f3d29f251dae7de6c5c7999219f6f356df794372f77043d4cf15e96af661526cda277
zd6eba039f903a77a7dc3308e37e69d32683e533b440037e26d356107979af9980642750ac5ef7e
zbeff91c5d18f47aeaf4905316da7b296df6060de895f1b9365272d742a844d5982c2e6b677b63c
z99f512bc9aff3fb725e94f3b2a224c9c22681af368ab6b00f184c886ada46970585648ba83237e
za8f23153ca629ceca26eee41d3d51620324eb55a6537cca4a6a81a2c5cac3cd81e27f43f3618f2
z05a3de71bb616f85abcca516d959e5c77385d1ee1c162aa66860ddf4ca5695e7f62121570b1442
zc3a77ed2c65035a97ba5a5a77a260bf4471e86931eb64192befbdcf862334083aa1f41470e6a9b
z35a9f3a0eff3da664be86483a5db2309ec759abe6645af81a99c70cfeceef8a13d14ed31ca1102
z0efb38a1f73f5e886059c246917bca8ff97deb66104d259c56be1d937969d06b208182e97a4f97
z115a75b8a45a604d5fea3d9724255e31b4d30f150e685b6d430b933ca71e2b282b8dd9e13f0bb9
zbbc82b68fc92a7a4cae569cc0c1f98c4e9b3ad4df0a0fd60e40978f544167939d63fe0185901dc
z2f240af7f511962873d4abf02b0d7d7b354f44fe479dc37632d6355321cd841e9952a66f6a4d18
z29172808fd9768e4676c6f7d0981b5874d7d9870bee188188c8d4b395e5ea89e030d6797757d6f
zf9ecb951450d501094da4937f128f8b12b38377cce36755c5843dcee64b8a143af79bef6f786e2
z0463d9e57129e2c9a946e24de3335a2152638096671f7a80419e71625964a5de3caddac52160a4
zca413f1963d0603f27d798f73a3f58787c04dd05dff7095990ef7ab1ea7080afe2e8248523ba49
z5c1072499cb66322ad94c574911d60c0e9cbb936663db56f801c34c4a43a3114ac829353216070
z0f3fe2940ab6a819a8dda5e12d4d7016aff89e4e94c5b66450df8ffcc6ec6f876daef780531e30
z25a37b03fd29742f6199fa49e8371231410bf05bc1e455fffebda247a40153b5487071af069b03
z5b559cd75f6431a00c99703c72e17b38ea8db770cbb03d0cb21497a025bb56f2d1d0fad8954c32
z11d05fadd1ea29e220e9b3518631ff96fdb89bb03d9fcad6fcd405cd5251fd365b5caabddb15ab
zcd5ba567e32bdef306c289474c9a9ea69ff04ceed6d5e3ae0eb5801ec47f5c6b433023bf95a40a
zb39cae98d73347a4ce4dea7a65c79bf096fdeeb4ee37e44594ecfe0200ea7f9946b9f3b6a429d5
zc69168e99880d974ee4d6edaafd3bcdcf49c360234887ede40f6844f5e38e1f784d0d18150ecb6
z4b74b6c7ccf215939a747f17f5edfabffa5cd5dac45d22351d83b2de9bbfb20be94e7a8bb65844
z035a21e09823206f70a1e64c2f79769055d7b0e9360ef1fc55610eba908742ced5bc141b734e7a
z11c1eb6db1fda6d2c5aa5f13a1f6b2c4695b6752d86005bdef50f5a2300b37ce03e668deaf78b1
z04b7242c57241340126ac88c1171ae5938dc3bcce3f9f632ce45ea6c3a3d41485f75fd74f1d2c1
zc75bf4793315ba68bac66a0864877b4ec1731840ac758bcc3d8f229b05920607ccff32e41ac659
zb0ac604fe3ec1eb1c8e9291015b5f8075937bfb245e0c9255512c4d6074b69a2f282ee63745cfa
za3219c8fea2453f4ff9a60c0a06a7fc98eafe05f27e4e33badf52f1f0099759601b69f5cd510d1
z432e3f6a6f9269440de25f1195eb6c7478ef5f45f3d1cbe58a377c966ed8b3cdc09dd7224aee53
z01cd280f6f7045e218fa9afd48af89a07dbc231701b4b3d905a5d33c4ff958e92d023b2fe1bfe8
z5c5ad379dce9bead51c5ceaaa3ce1d6932ede6f99896f8732ed716b7fef098320ce52a5ae003ac
z206c9105f953d4954a8918835cdba6ef1e4e98ad3cc64030af2ddfe1ec40f05f4baef9989f29e9
z183c5230396eed814b0719acb1d114c310d59adde6c5e6f7bfc6d03ce3e163581274fa2b3768c4
z573a342d5fb0f1ba5f821da37670e2dfb433ef9b0c7b8d4d8c29285f92f06fe3223a5a28ad53b1
z6b782f93f254a5a3a7aa01fd9732dcccefafed0750fffdf344b960486b28fba69c5080e820932a
z31f2a96b83300b46341a4a1871e1726b9b7e2905e6e885ac3b1d3067ab6ede5d97fe58cddc44ed
z948e46208300054f9b26dd6b308b09a3c5f2a1e79a18ab22ca193462a8f26141c20756684aec8e
zd5c8822df02a0cc2fa89c8989b5ea04a758d54a0ba5b839c81377f9d0ea132838f8373025f0ce1
z75ec7824c79a557d7cfe14cd91d16e8787b38290fd9897a5b7d359a20fb3c2bfc96170eb08f615
zc91185648c0b68c0878b1c0b05c6a1dd5bf2cb574af418a4f2e9d9195b5c55eee1495160a15016
z27d5a305bbf9dae480f9e5450fd0482c9c8cb2832bc21202e0cc4bd16c886c1cf46450e75e83e5
z09b6b4c0692f499c499e1a4c7e8de9a90dcbe7f597d9eff06ec88af033d7c0125287c9b7ff01d9
zfb400f8351e42fe7f01ee8e141f47f34f476690ae7e17a87a644bb59d8fdb24f8e816420565c11
z24b7f9c06256f6d3fe3a6db0ce3b813d63ed1935cbb4a59036a193363929aaa119ed9b4fab8c7e
z9722073e03e3c78d543c221dcba0fa841e1e831390ab8d220a3babb19e6c48cf847c1de5de8f03
z5a98c22ef15912af288da85d4faaa60c77c099265e44d40b8860d643ac4b40914d794d3ec7f25f
zd19322eca3705991cf00b0fefd71c50b52d840990044b8e6f8109e38578b27a5a03c0f9b737526
ze5d6ce4a5dcbbfc5b7911fd24d329e30243f683531e5146c42818240d2cc3dc6e2e3480fd627de
zca0f0a99b4b40247e626f15f7e716c715dbc773d52e520a757d654db86cd769535eb400517ebf7
za25908df5fc03cf71137fc0a5791aeeee39dd31aff5217cf46a61b06c12f490c37694de94b724c
z920741bc24c7a1e10f42b23dd6f312145d68afdcf18549fb279c359f6d9a016aa7769fcfb215a9
zaa679d17ff7098e880089040cd5f6e9199066bb22ac21c9e9ceee0eda4be2a7f139847df13d938
z7dc86409b0cbd76f18658724128aea00ce91aad6a1bd419ed6491d0b33a04744e66d1da22c0bf7
zb7b648b4810d389393ed4467c34b4c2f8673d6e54c7b991a1b3c8bb6c577151288096e4ab411dd
za81884a7ba3f6526f0456ab49e6d93daf375ecc08801d7b9102d836b67e1b44930675a2bf38907
z17eace1b6262ce2b4c331a5c7f2e478185e469ea8fa0462d501c755366d909dec46c3494bba145
z6085cb7074e4390ddef35565a192df48b3127e77fc3818807cefa42c00b086eaafe428ddbf2702
z5b9969bed617fc4d7f88a0486051ea0bba8ce2bbb291dbc49d3820d1c879f9022b1c96dfe7e2c3
z2110a7fb3b22e376c31311636d6fdd3785a9b2f129e26ad73980dc2ce0adb30208a7784213c0df
z50195c141edee48aa77e30288c43f5e1525a3580925cb3942a5d146db47d5a17bd36ac16478ada
z00328e203eb747212bc59e5c61421bb2b4358e844ab96438d8c2e1c6a5ebdaa44a7b9cd9dab2a3
z6f654dd3abbe3d08790bd5c8bf0729c10d49f695f65daccab230e0ee216f7c6117ea855caf5ea0
z1a81f3e87869af1c2c8acf71cfe43c578694d89eadaea11e8054773840e82b632fd80adf1d2433
z29c8bf148dd296e47c4bdc9e629f71e10ab315bea8a7421b04be8014f6fc6bc7ef96b656935436
z82b43632dc943de6360c1f601949550071e1ba4ec5d9521b64a38dce46d756926398038b563c1c
z68d467826a773c349cbd5045997313e974c251624d70de1e10d6c5109abfea4d7d17ff019ae406
zfbcdf77fdcddc807b3e77e070fcd4a151f088e300fd6657c2afdf76cbf59b0ee30bdb1b3928aa6
za2c4cb5d649684f2c7950ea67a301e8acefee9dc57f0a625d97f2c9592981b5b8f9d5fe5ef0f60
z911e34b29e7bad01c30dfe12f88f9f6ec8c52ebbf60d1f30b27bbb79203195d423b4cd4a981ee8
z1b7272de09291c01a5f41c7e31c5c9046283abc8a6ecaa89a331cc2298b185333c335a3cb08918
z44677a0cab0bf7d5073b451c04d0bc1238c6be58f7d53ca3527f4dac5bc61709410ef02b9e9a40
z2b04adf1d773d85612d90118ef8feecced4a21b8c14c64f779f9dea249ec68d9cdf46ee36671aa
z41a1e12a0dbfd94ea6a0129e1dbec0a51a1e39e4729eaa824e055bb9e2dad52dba5c855ab3aa00
z970ad85500092b004735efcc7fbc86b88d839a038870244ebb3b9407cbc196626131a60c6d8a3b
zdfad93d4fb6d2d4545c0a4553373bfbb7117ff8e70d63a0f0588faa474c4f17d93ac0151b1f9c6
zaf972a0dfc5b7caef0c6ed1dd90720bf57754bbc5cb6ad1663f8c00e6ad8e9c53dfac2f8527f6f
z50f1021b105c4282de4a37dcfd464442e75e1ab995d5b90ca73b22459d51547cadc4b15172438d
z48206ab4755b2c27bad0129882cfc565464b85c10d756acaec9d55584b996ef83d1f29fe78690c
zb4bc97dc1833f3f1597ac38c62533a00f4ccb7bad4994dc747f98b09e6bd564b49522e5d4d0a18
zba2884d26c2e7fd9a86f1a65c7372803e844fdaff0531465209477acc4a5df353c9839f3a3a5d6
z97df220e4ad8c383e7709b5c160257b52e9997922a75e8bfdf5218283bf172770d51749d4928ea
zb82fdedba3ff1f057940458cb948247628444c38f0c2984576cc481576c30dc2f3c9a599c785d0
z567127f9392390188bf6432964d6c8c438148a8b7fc2cadb63b7b3ddd25face93c0702376f0855
zadf852d0141102282fd7a187ac6b883551dcfedf8f982cc0268b7eb390da66526ef41c564962a2
z3e8b280366433c6f9ce0ce30656e4fa630d6b3f16522f4449a582cf035e425eae4e4591eb102fd
z082b449877d2b18079a3a666a54920c2a655d3e52264fa836ca31e6c4abded9db7662e98e3a62a
zfd4a6d56a53a3f4bdab2dd7c02358947f4e36b5a2e1425264a7598c5e590451084233c6c67c360
z916063ff285dfa1efa65ef5d27a16715f518f0a5e683b2877e85c1b99efcf739fdcbe42a763951
z4843b4195f2b5a5af5df424d71ba0d4c166c10ad004978badebc544d475a77027db4d3eff61e45
zdc2e7974ec9d5b70c2db2211ae88c689b8f08a3b10c0498707f338d427a3b75b37332a5d533ce2
zd968432c197c51439cc3838033b457d6c142814d8e9f8a1b9324ddd07ce650c83300e0dcfff685
z0b152036d5e825ea9efa691923e86e44da66cbb4ee5bf6bbbb87da562f1e047bbafcaf0c4b2f85
zecb873c4a6d0cca3994b3ef5030081ef93cd859760dbf9b483ecbc4c5f6953664bf9b3e619a103
z65f1afec75220912bfeb9316ec8863312a5d51f4bada3541e7c8b875dbba6e5891048b6051b0d1
z722943ac87721e0fb812c33dfe9544adf0aa6f18f0e3cb9db2420df8bf65c39ae0bbef4deb9807
z92f161a40edeab1381a5b2bf921744380f79991602673843fc8b38fc901afcba8bced84465f94a
zf7d45a9612306c4754336b1a5f476e92efb6ce5d07b3f9d094ee396ab56661fb27020f3e9cdde9
z690b44a8fb5ee623390c20f24ae3673a7fe7209e3ef25090de92209586a2eea79e5d0885463477
z8467a6650e53b98895f964d46c65e58fab37764a877c0ff4865214a3801b3f4533eac7086abfb2
zd352e07f86460fc3538434976536a10b39201f79194fe38c290fa07ebadec28dedfdf1c216cd4a
z919e81b54d21fd5c9ccdfc898dd9a446ba9a3f01e5fd103868c95c266a9ebb7682dbb463fa8bc3
z76a84dc06dd8c0cdc6415c969ed6614ab1cb05dace179e14d83ffad5091072e5a97c6f890339d0
zf97908348cdeaa261d022bd3544e62b5294f28c7aa0b0ea88fb18c88d8a2017e3218de5f23845c
zc3c39c2202df74baaed18f1e5048e5d783d9bcaf69c2b725b5991187acfd732ebcf8094218c75c
zbad16b898883f4fe904ce10fd4f80d0ea9f338e6e4121a73e2431954c04ed7389cd1e02e74086e
za821976163a294002159be212c7f707a4f5f8723f510ca35a0f8fe2cf48bb9c5cdb0cf02593a81
zb208ba4270332668284f692b9526c7f09324f85dddd08b9b5bceccb7e460ee1835b9db19806b93
zf5fe48ebb86656c5625bff1d4d8b65f9fc11e08fd6e0e3bdc3c4c4627f9d4240cee9624ccd52e2
z0705e21b4ef3ffa870c44c7cdddc6f110f2a7bd7bcababf353cb0e1e3b65ff62dbef9406ce4471
z5d8426884e6d58c5621a0d1325e1895dfb7fc3c85e8eab28f2452540c29793f0d6db49c9b387c0
za8cbe2e5e815c4146269c8b6695a44bf5f8b5044e403847a0dcfe9a2ec7a8f7fbefc6eae413831
z53ca4a26485c1276c312e2bd9a2292c8b39fd25a656df19f8cf881552ed7b2fb1050a1ee0c2a59
zba13f71e9c6747bb3e1082efd0d096bc0131209b341997f5b7a78dfd38f9fb2ac57ab3fe71a4e6
z6a9b2faafc3c080982aec0bb3de76024714405e5a689cfc58dfa7c444dd6e276088491663db026
z52420ad891a59dc0e9f833daf88f8982548cee4d624a9e7f8ddfb6478795d75f05564b6ce3e900
zb48561098ef738f0ac75fd3a9040293bc82827e0fca54743f068caaf73dead8a809123c7b6fb8c
zca73b642326e503fe254599978af2b83a9943e8665d84620389467764404ff7acec9f16a93af4e
zd1e05a1e892fcbe58f1d4f834dc7c362f8917bd953e2994398bb882a5567c12ed762ad1f9728de
zf611747933aa1fa79bac7430f1f18aff57f970dc8659eeeb12139a65561e7313f4e9e4ea3a68fe
z4e601c0fdcf7c99b11fae81e05faf2228efecd3b9ba6b816bc334c02b02b2852f0f20964c51db2
z0f6ca6fdff2cdbb1c9e32889521a62a96bd1a698363a4e25c45a45a5c3458c5819a4075780455a
zbe036ddfdfcbea37d2344630e06edf127585c9d1265b5d3fbfcbe5c454d12db8c206c2c45a5434
zead62f9c089ea19f46962e1690591700046bb10f2b1c6e78822188a33c5abbf366c5cc0e85622f
z9a3d848af5afb630bfc6247d7d92e4a05cc414342720a7563688f9e1efdffd0207a69d405b78b8
zc9436835997e4d54cec15036eb979d60471367f46c4ada56d629eb33c52f168ce8d7dd6db2b816
zd97511f8eb21050d8f67faaa0dc9524907e80651b4ee7048b18b1330f13317d9e667dbf82af643
z75df5c621eac2b2fa97880112d1021ec3ff65666373d16754d9e587f7601243f5636c02f252e37
z0405f6e5dcd9cae350c4a5c119e776d55b7f15dcc595a2bca8441711cd4c77406b3d49b7491425
z9160a74a6a36d40ade5d979e164ce22cf5291d44094e82b493e0a603284d7ef6d09288a0f63533
z34f649a4e4bebedfd7911aa9930ce293e8a02d3518a191a2890054c9ecd3f62e6f2261a33eb0aa
zdc5793e2ca2ea9fb03f9a21ec1e608542b464088ae009d67dc5723f324d263062e38a462b87629
zd92262ac06bbed61dd0601e6e3224130d4d88ee2514fe82e970d8c2b6f10f30d37e5cc9f28c6a5
z153d137afca70c2be6e358317b345088e2c8702a68de3f1e7cffb28e6141f34f709113a42922a0
zfa5cb92882e8206196a0d46eb11cceb61b0b3e8aa54f042f630c8a15b78fefe4d647eaa42fa609
z0156b373994cc49e318488819c7d183a21ed0d000ebfa81a795def989600e19ff0840cc10cf88f
z64a7eb2289f5e850b3c39750d9af5c269e7a385c51002033ad823710a79a030371f5fb5e7f89ba
zfd6806fed52741e0f83c934f9bcfca01785e3c357c91298cf17f1eec54ff4b3a9eff8a591353c6
zec2ece2eb182e045dadd26d70b804413bbcd2d35bd16d3741b3dc0fd888abd9d59aba9b8927c1d
z441c875bb4413d159d76a55e291b0d53414728f95027d5ad8299af559d0d47ab941607144d801a
zbbdd4dd0e8a525b49a1e139c5d0899164fa77164a1bd4619629dc768523232efcb9ff9c011ee4d
z7b9a258824929c8530d6a43041a55e14dc66474e581e391fc740050755007b2ae2835c69a58853
z9d4a33c8a94ab66ece8f63a949d3b60d256b50bb4fc554e07c5581e45ccff9ec1bae28f4745437
zb44ec5da6af9dc8bc9ba86fd6fac069589c734b2dafb0ab328df34d79a8df4a695e83352634894
z439abc107fc576a7b58b4808bc879bf5058589d822b855c9e525eb7738a9531e673a2d2c448012
z94e03c13d27c44086b220da411a38af2bdb41983cafe9b6afe95869f83f600064a1855f0d17ef1
zade07a07cc0349ba58104b3adce01ce370c3d6d362cd97d8b4d61e48fb4ed897c9db3ad79782ed
z22afdd1f04630928ddf9b02422ff2f27eeff95f705b8765423d730d7f7116b587b869726ea58c0
z4f3a2962b1535e5d888b2f90b562d11ee4387a0333889d55375c668e52783f346d0053fb7043bb
z078291ef3d7e003cf08768afcc1e1dea5592ace4ccbcd5813e85e8e72320417448669290ae2edc
z89da04e39996edf8f128fa5d73812fe2e584c3574a070128920ee85ce34bf3ebb03cda5e9dba8f
z9ee05fc465081e9e7dc0101840a090543f4c13c43ee08be3b91940469e4262f9bfe61d6fc05d41
zeacce57e527e08eb0523ba4b46f89ad7a3094fac3399f48c298897fa6ce4bb96ac0fbd9312cd34
z21834ad59a208df645e274ccee0c7fa9cb9611c0f366e1561a7655b94382be907ffd521ad1f581
z657bbe31a8aa5445b42901e540251720473e48d8077053ffea9b6686471a7b44a64bd8eb0c42d8
z9c02ccfb035f5e3932602965749f30dfcbc9c8e91a151c6296eb8d50ae5e015b9b5c8b495ce18e
zb3a95119ea67f8611cec429e489e033a244d5144dc1a2786d455720ada0aaaaf5ad93814b9c86d
z253a845f062edbd1caa814d5275cfbfacb2404ea5bcb97393ddceee49469226c0b18633132e3a3
zaec41d81b345c30ce556a4b6ffe55b878c5332f822591bb7d8bc272ac59bee90286c6229b35926
z8c07e44737f648c0fe8b8c4c777d6ff4e93e5cfc15e146ebbacaae80cc0d3cb469647127be16d3
zdbe1da81d007ef48123b3f5488a6a2571cd8c694986b87ac12dcc34997b66f4434ec1ccfe81670
z4afbd6d423919ee86ccbabddec8e3c0b28b552b4610e1d26e22c91bc6d522c39e5a1a9ba5f2dbd
z7a9bafe14265cc512cc3a7eec62749762caed25b2adeeb6db1431d4ed2e07a84a50acdcac94854
z3788c13b671d0b579126022548ebdb5122852f17cb95e2bc31dcce2dd843e82c262a7ec6a6e607
ze5dfad083b8f7e04700e993d056b3abec92712c438cfe2edad7de16e2a3981786267157c5a64cd
zb406e788e4da560a5c7f7a6f2f10993ec0c3e011ebfa7a0b56cc66e959649b9238e827200e511e
z764e3eee5e260a0b9b86dbb63f4632ef8ec388b0edd43a4c39f4423f8135aba999de8aea561a45
z5abb571b28abb27cb5e0e53fd3a40c5710a32550a7ad4c7e24218a504bf916da0df69bee87aeef
z633f2de163b898f60b8247db7fdb65eba34ca3f3c1591829d08afb20f1ad42211db80cbeb9ae7d
z8ad46ad157c55aacd7311cee07a9a378a9474e4341cd6b43afce9718995b908dec04beba3dcf68
ze2f888e2fe9746afcc25df76c8c621b12ed4d906da06bb31cef33254027697e55326f85d175c3b
zc9c5bc3780a7a67e11f5208e5f93931ee570aeda90584c14b71c4d5d98954e5e53c5c41321f024
z8358606c13304663b727989638711236c5b4b1c8dc0fed417ffbba2eb37e6abbd86ba531239c0c
zdf22bd47d442f9485d2c79d102faadfcc4953625de29d23b4e6eb685db5cea0834098ca1eac31c
za5f2f570033b1c1cb496854390ec321d8b0c22b8aa8ab5f50b46086e6eac1b07c12235ed9aefd2
z88ac6f315700f62c3abd15679972b9cfec1db5098960883bc5bc358de2d7f68e45756080ce91ec
ze0fa36eea270433238d9c2661f8e99d8acb7cca371b0f75648e4574024bb9d745b9a0b64a987db
zf389cb2009b59dd6c77f0e8c3be3206d86394b41934cbf8b10e51edce990f304cd5ce127acd4a9
zb6717380371c8c459aa4f82db7e9e1073db9c9ebb6095e8d3601c4a032b76d734cf7ca8bb1dcdc
zcef8dae89dc1f95a947e844d6b87b2aad12279efe755add3bb4e196e9fe4e5d615bbf5dc979728
z7802ebd04d23f354bd17139faefc3115e188aa52ab27bc1d46847f8b0212f950772ba4c69f607b
z8e51e57f5ee105314b1ed3e75d01d99d826c7118e234c8f2228331933f3ec7e2dfe1d64c9e1a06
zb5941600add6868de3a6fedbaf599f467dde27f5eee61c88d2c6921c32c82209095c57ad6708a5
z38f5e380ddc3ea785d757d3335d8b22d0486e4a5d20ac8e1aaae2a159e9e0894a4e0f5f66b035c
z1115d3ba756c2a4a60883727228acb09eb1f5dfcc203bcd16b81649e1bd16fdc54ce8de0a98401
zefa32d31ccd0926ad20d45db5bc6e54f8c48ed0856bb9e7da060a285404a5cb02f981d22665610
za4327f97bb39f8a5f435030ae5eb297e48b82110461dcfed6d44f9444dc775f1f17cb10b9c1341
zaa57cec34235b94d5dd22daa6c6ee79f4cf0ccad084b33c5597e655b6ab4f6f6b08661c888d201
z95435a3deba73d91f1ab039deeb3bc0667b219c5471cf08c52f306024b1fa920d20eaaa9ea1582
zdd895b47625b27fe8240b47300450b95fcf7eac7c2e1cfd2a5bba673d814d0a0551dd1e44ac0e2
zff04c6254795f933ea5091b39bec3c37a1dcabe4cb50dcb2f0bc7e5d43674ace357be37ac7224d
z723117ec49ae65df62a58f9646c7165d8d2e46b7c4bcbc83a86f25ee6fc235780f88beee6e2148
z1ddd1a68f54625d394d2a1b050cc28d7c9fd7b0b4e90e86347ab44ab7a72bcae819f0f4bba1407
zc6ef3fe2c32891aecbe2a4c5a0a587ca32b38d6b8811d9f7f8cb1606e81174def7eb698152637f
z8ffb9ca28225ad97adbcdc3191d389b58455ce935527aaeab71e8e7b3113a51d938b79e54730b4
za08748dc59907f7b871de261e4a6c1c6d8e71d1bc93519508930f34f789bcdd59cb4f24703dbb7
ze1d777bd08bd98c36d09cba19f643403addf7d3966462031cae794eab00bd47c0e424135a6c124
za2f312af23825ded5a894fce1782710b8788a28f2d451b38400a6fea5314cd27902a1b7ed6797c
zbda13e8ecf0c1edffe8cdc91f31ffd0ff3a66fbd05ff0078801bcc34950fb73995bda339f6f575
z1039b4415e0dee680f68caace2e7d10b5f47d633dcd3de10e7c5abb224b8b65f7b9dcf0f2f06bd
z140438aa7660dae43bf5fcbd666b99429636b28265c6b7aca0fd826e73e7e3fabf2e9e26e1e899
z339fa29be493664beb7bc64783923ac063b9976a7c9ceffaa553f41803b5aaa299a16a273b1e9f
z2d4e6feeb3b22d7b70a4e412780a4583b4a0fd679d1b8ad283d9f6829cf4dc3565dae9a376d50e
z561ae69819a020d19f05476a763cf66e043a58feeb190e09d191eca439e36f9e80b0612cc59755
z7b3d0e798db1cd8e0742af1f56930cdb191695d8623f51b9cf082369876b3f73cedea77a562344
z857ffa0b7ff5cf3180fc605ffd3c07c7694dd4f9ad6d51fd6a0862ce5b93bddde526500cea94b7
zf5c56113c5a97a324a201f3ec28ffcff6c04aa9b1fe6306f442cf94a17734acb7ac5711ee48616
z1f0d6de9eee10a5edd8594c887b49a19a3014e92b2a86eb4aebb347099cb220d8a9d32c31f562e
zdf2431ff6731c40084980455deac8d953112226ba61d93d937e98b67bbd0b0e61afc416f17c93d
z922a184c5399468638a298951450bc2940a409f97c0cacef747562df4aff8b9471ada911e0ea67
z1964dae2d4db6c92107de7db184e6d88f1ae258471cd517a5caea9bebb40a5e45469bc85fe5707
zbc49736315e1e7d16d8aa96aa02f3f48db5357ca1bebdbd54b9ba0be638be1c08ea0b069af7a54
z24cf7e1adb71897ebbbfff4921cd499f93313aab57db5938c37fa1af79fe64e20bd4700c0b5f56
z93f754fa1d4524c272347e0078228797c56cdd86414cc6a3e8dceb6c461c6d91220e3cc11358f9
z46c9758efb4ed1ac8bc2f3998018c29101cc54c4dcdb9d359ff5e20418365d3ecbf41e683ba3c5
z980d4753043f32d2b98f73d1693ac8af01b0b030f20dc339055d37e0ef5275ce9edf846753b88f
z0fe7c23fd8a651c009c800142cefda326c68af5a2f8dbad3a7c7c238540035d30f44082df8043f
zdebcb3350ec501f2b74d936c1af48d885b28e4bd8f7eb072da4265af0b31293b97fa3c0f32363e
z5b661e42df47b3ecd5e40d01ebd7860d377bc156e67036ee5e198c6ff705af8eb7da4dd3e03452
z810a0079d6bf367d6d403127cb6fc173324a61de545e3e2e195bd7f9c8d9e25af929e485957070
z23305da8c3bd41055c75c418bcd84669c60e7827fd126e2adcb5d3df2f98ac6dab34411ecee5a3
zf5460ec540eb62bfe606a0315554c928b9660962a614b07f06ba2761eb919cbceb81279ff4db8c
z60efcf4f0bca9ec5cb21f1562888e3ac957cb1f031c8011d076f48fb258bc08d4c3193f669614f
z20b98294b28af3f00a326a105f3619f00132f0838b53d043e214ace35478c66d79a372b696786b
zefa37788d1e54a047c6ed53ef076c25ce7b3d71dd2da25aaef4e57512367a378db8938b48c95ca
zc781bdfc8f15fbccae8d9cc00f80e516e31da0fd1270d868ff04d53bc5cd26444b8728d24c31a5
z778c08ea3318f2405be2d78899e24043621c97c72ba3c2df22295b484272492365e3cf1d14263f
z72aaea5544644c43d1ad1ac9cde88b495ee28a99f19b815b36fbad8e9c3967a1f9750745841cc7
ze1cdbf8728b08b2b1f6d9fae8793aa5e109e851226681473152046777b9467384264178ed46405
z74e9765576c534f8cf8bcd7b9b643a74c91139e4558e00eabf7a61807206033295b68b2aa4a2d0
zf5d771f724a4c616a2d01e03fe95d5e1c0d823de451dfe6cd105ab71fbd9c8dc33701335de0214
z001b818f8f10a73cb28bbc27a12e1f23daca6a413492f1a087d70945910948cc8a234e40e7ab4b
za16da1f81cdf09e4d092c9b19a2bcc9b60267b898d7dcdb50669f6d1bdb9cbb9c70a583edbb1ed
z7ff7247e889ea8c65623a0398081fc7b3d2389e39a6e167d56e25af50f098f187c7eb295a7d4ad
z1c05966a13d9b740570b60b84117a910537988f8843b1b2a2fc3064a75e5b602d31d09bdb3d19a
z9f20070252763fc627e8172c85bf35447890386bd83b0709f3bbb261d3ffb7b128d007e9bd0d0c
z602ddc8fe321acc9b712d11d62c1549064dfd670531b1b1044b7bd126f38f549e0e468cf40fc2b
z55312401c8ecb947823847c0b460e9b340a5eaabeecffa5a2fa0ea2f3599c48979f78e698ff613
z7fe147e31d69c8ac69ba63e6aae03116f186db1ad7d2dfcb656334afae840b53e0855b05245311
z71fe00d834148e422fb1c62fea48010d1a6fee15d782e488d724dadd928787cdd3274bb7c1b79a
zc2599e304eb526a3f4864fd7a11c5fb71cc18171133740b6acb344309468b8964330f99a47f24c
ze18c09805aa9de3d443695454fc41be0be7c6dd8c68ca92a88e85c4ed9ad825e013e010f0e52ae
z24ce9a0bdd0c008d4d9b7bb81de31f5347e418d15414adc12e7374572ef2201f627b71b22a129e
zd35e9ca2b46658a463a5a10c04cdece3ab205a8b1f9fec6e04d785d89fbde413fe233d0028e91d
z3d06b90088e46bcb96c7529f064738d92d127b75cac2620c253a7d84faf47c8f464dd80507acb8
z995a96990c6f5eb4129a69c8833a095a05fae79f92ea2415d53bf99e269afd6e9d04cab452e3c2
z714b53e83c4a95da607813d8e875a8bf841e54bdd35fa592dd37d418f7f4391dc71da27abd5fa9
z0fa509760ed0f618f344d59f976d663ac0216fcc343ba7045299b28e953c6a87513afa1c0e3e8e
z6f24923a6bc5ce8e383b5454a92b4bae3c43f20a85a99f9ab3ae6a4fd3a6b045fde0a7aae19fbc
z3f8d2a22f277b236585fa07062013bf4824dc9049634420c71006ebad3847ea7637b50182368c2
z6d3630fde593aeccc45bad56d38e8a8df48da2b87900932a744b632bfdf332af4b69f2a24a8d46
z554a411559a547f33d7e9ef58647f9f2a4d163fc73d240d2910d343063f1b0b8409f516e385afb
z9e47d7b795643dbd7cef20d4451f34c2085d7f6af5169ce6e8482a4aa4822fb78d35271e147af5
z1d652dff8356f89cea45ae84a4ada9ab812512301c1bdd18ffb06818a62feb84deb37038896082
z6efc189b855ef480ff2e536cd5d1c0acd9580a9ebc9941dafe9436d7af8120742868c88b490849
z21376348a972218b61a2a07000db6b7fa765217b8e55eece3d4272fa82c904ca6fcbb7395fc93e
zef7f02aa40d07126a5da1e294f69b970116240a1b4ae11b3489738c2104f4e474d5fddb53595bd
z231b7d711cbba8e27ad805bace133d0804d26a86a79ffb3b1a84f768464e754f210e6a24cc039b
z14a51199b5a15f19d93cc8a7013152ba65505b24e25f94acbca1df22c389724bc0911ae95ca6bb
zd87fabfda3ce9459c2a2cdd8b54698fceaf421b09503fc0d22d5cc3e4eb829398b93d01ab29158
zd9cce7a6c15d37d0247041dafd51c2916baba8bffa94f685596b541be36c41e9f49dd036418b51
zfa4637755fb51b3522db24da37469ddb76532c50297980c6d530fb147e615be93636075d2a043f
za712cfccf7c17ea2ba1b9dfc32d0d389801f34fd480353271dba2952d7652da569cbd8ff3690ef
zdcfdbd3a576831b2ef1dbcb584320da795562c5f6f333a00de26a5e36769ba202f825536ca7166
ze25d05e62f94db9e6710e8f339bcb94545793256eeafab572c340fe82ec58c2129b3597ec5f7de
z24e73398d801161367443e01e2d974868e8dae8c3118e35ba77b859430deb41b460d4fca855b11
z118950b8ad583a2b9948b20893ebc69808336c63a09f8936c08515bec935e1b10e3ffd900943f5
zc8f58de9dcc5618cd24181e804f291735059763bd6d379507ab2424483bf10eec1859ab592aba5
z392f5a902262b399c05f34782720dd499abc448cd125fa1bcbb290305d36ea12d1fe5250b0459a
zd907cc2b2a212dfc8e116db7930b096e0ab86c411e55bf7ad7a3ca76c3d0d13c2e299d351fb995
z11f4049007369a39877ef7e8f8e256a50aa757bdb530676e15e4c66de8ab950941d4533ff02293
zc8570c5c775fb2ed058399f1fcb28f2fecd9afd262df538e63c631f8bcbc9f70ea5c0ff674ac23
z853a6f62b78ae4e39e14f4b2ed28c73f849b75be170f77289e60be3619b8bbe5f1ad71a45845ac
z020e3055b3496b2b062d0d4442deaf3e04e672b76f498c3bb64471682bb9d70637c60e19c66e35
z37f812c19a1e1bb0c3abebeab16fc192ac6ebe139ad24cb49a5bd26659b0bb731efa07f70fb60e
z1754dea8574a7b3a208f6fbeba44382968e7c0cdee525a26722f25b134130ca6d8838e64987447
za31ee8129cebd46be8cd242ed8953b08fb004601a87d24699325e3d15f38c7a02af3251cb509e8
z0442285d52c6f985cf8d51254d8c0a2f395846b09c9b3231fe64964b0489e0db95b493b844f338
z23292b747be0c62f1b025a40aa951d7258e318f6e0979fe285b07aa9e84ab0c8c54dfd3a6cd37d
zf849566c5f69e026ae1d7d9ebbb2f38cce52ec299352c98f5168ee81fea7d8c60abac7dc713369
z17a3a31bfd806048f73eb3216b86f4a4641e2851deed549adaee5f404a8f80891e9afc423db527
z34e08aba77019afe01d902177758b249093ac27ca5d5ac9d4eed701db1ff6d5e948068576f9c10
z05bdfd680ada91744e3ee10de67affc81ee7ae26194e52d3253bd5f6d28a8cd3657be59c444df1
z64601b9927d63f31c699e5fcf304edc69aaf2c49275d94409e8e7dde324007099354518a4d1190
z442eb2be8dc512afeb35d75be59abebf04309c435ad1f0d68c23eb174925bfd6972996f2916b30
z53f587d0621822fff369ad77f44b5e7f70e2d663d55653679530c1623f64f5b9b17cd74263dfc1
z78e4cfabdf386dee8d6560dac6f85c57ab6853b0c9d33e6df123a4964027227998a2c9675e466e
zaa58b48e89645520f1eceae350cc55c4fa249f964333d88d173c3baf2b4928b038d0cc13b9b137
z6af97d8e225574072337c4bce92d33679b63932576916cb51154e5f199fd9c5a2681cfff9dca73
za20d806cd2071703587cb5813ededc38aa8e82b916b13b90571ae7dbaa05cd891b0d480d1d6733
zed007eb7bcf305aa98094971449bbfe60b68501db28e48d8e3bb922418f2cb6e641d63fd0b3f1f
z9156ad1bb0e403f7345d20e9d641bec70e158f7a0c3784f712997fd8e9ec51273231865e9734a1
zce9abd6d3fd4fe0888c75abee5e2a133cb931446c0a76b9d81d8779dd76bb2ae96ccf95884c71b
z0c80c84c4f165005d3586f0fe8ec4c723fdd25bf01b9dabaa1a0b24bf5d710fe7e33c61efde905
zbd64eda5f66f796ca23a51f337686638ff5993eb305773929fd9908dcc0782eefffc1234aebf25
z88269fd3ba9c5e2a9449889cd1e6e377f622cd0c49bac0d4ca803ff654edfac954332400332fb6
z452c0fddd24716df58624a276ccfa1012196ee467aec392f35db18709e387254e0ba1ce17edf25
z440ef5cb2c0ef2614c77c72596a53b4a684684c2dbf3fa95ed35e456c464e03a1c7c97da41ca00
z3853c0cfbd78fcd1295a1b64cb6594618c01c9104f31ade92360b6c924503023b06711b53e325e
zc64708437330dcd6c40eea4dfac6c467aef1bd57f3abfb26e98cf22cc787ef1d85bde9dfbf4cc6
z99945334356e61fc90d11cf94aac2ef8fa416073a79437f0793a9da0afbb566f3619ee940ca951
zd38740a37b7765a02fe12589c1c9705a8c31bc5850d26244c96fa950e99ce6ebb57c66f09cfc31
z49159ddf8f45b872c4ff723a9b814b6617d40bd10397bcf8d600eae021a733797a66881c91cce3
zef763aa1257703457faa4260ab1e62644bd59e5a71a709a46a07bb0e8384c09569915209a94189
z46dfcd34f9eedb15052a65dc7609027de1dcb7a0a8bcbf88bebe3ec81d50b18f8afa97bd54bec4
zce582aa35ccb767f5111025c5c60475482efa490d63d5c13862b0c905d4fe566190f534ff28d1a
z0a598a65c172916aa87a4d1901dc6a284dfee3a9817acc8e216e18697e58684b136f5566ff0e1a
zaedfa972840b04ad86998ea51376709cbc3aabafe7c4e9813d71c3a2cb7df3f9781244bd37b526
z4e3a2e81d77929c1ff72ad3fb6ed64d736f2ab7ffd32dc60103d9a0bb05fd5c1506bcab4498b12
z8fd2ab6c731b072cfc85c541807c1ba22329e04c60816912678a3c2778f56915761a0952dfdc59
z251abaa9b1d4c3d1c317545835886ef95dfcb70d3ad9166d2f470a80d8ee117d18c8593c621de2
ze2f652c49835eb1893b0bfa403f550bfcf560fff182f159b7955362925676daf0f1c49464def4e
z33cc65b0c4a85641854e81a7e97164bede0cae33cf49230a0270265dede0abe0972c66bbbc2dc7
z2568d82ec945ba3469bb55509a0c7f5cc196758df9d11d0413b0774d52959d29f66cc9256db482
z88d7321fc616fde12fd3bab8b62caa9c9f8eee8918e1a55a97af46e2f267908433bd7e22eb1771
zb89b2c50c12f031b738412d959cb86c25aa286ff15d46f6b72b78819d2ee8d0cc5c8f56f3d5eaf
zb2d91d74ffe3b7c9ce13a9b536b85399e244dfc66e134e598de4c8f7cfa7e88c3782ab6afd7d6f
ze76a8b29f3646a6e34107c645ec13de4b325d7219f0dadca7394c935e7834bd82cdea06beafab7
z49ae5da738d27e53d5339fc2ac84a2368182a69ec62a449fb040bc5e59caa57eb14ce1bcf469c5
z2a6133ebdb819946006753c7fb553ce109335425ae2abe5972426bfac9b1f7a72c77405b91e635
zead3ca67882ba777b302943c124360d386f2401a391fc5f65615a2343d23e53431e7d4843685e0
z5c0f9fc953147ab2f5217f9e6147c7f059e1e39c2cae4311aeebf6021066f43942db2dc447f3fc
zc2868de75de923844a5e366ce5f06569a6581578e5a401d41c5303880953dc8406e239db81cfe5
zf287542ef06f1d6551bab50ebcab537a9e03644a68db0cc70b5d731ded8ec16ebd4e6b5f015d22
z057f68274bfa9d148bcdecd218b3ad00e3c781f48437f33a10ed1c258c3c9be764c673d9f69dd8
zd757305c4d78d4e240a49a8d2e9c612227f9e9b04017b5a83058991d5b02c2af616e4b40883913
z2b458e74654e94f6bb86f2ca8f2d43b79f8f1f22fdb1b4809e619c0ac5f78f459b022cd7d9f9ca
z328555b9b91b679f0a3583ca81c094e46283824bdcf6a5398d976b4eeecb2f62cd9033ded110b5
z22ca041a31e340007af58123ddcb80c787ef6e5ed85147790ddfb0ee7218b7852188e508ead8fd
z6771a13ebf3c24fa9a111928ef9f5c7a62801b9975dfe83d4f5e6f234985855cfe4e46a9d2416e
z113b12dff556bfeca41afb23f107de77634e22df28e44d963c94d6b7b1c1625d3095db9456ebb4
zfd688ffee45740006f8947816fb1a00673de9ef7704ae9d6d0e9337fdabd0d1a11bea77222070f
z93db59088524fef730a5466d06e4d031d0088a54e0a10781b3f04eba0e563f76df3659833aaa4c
z382d49b91dc4aee2050398d668f3cfe00fbd413ff836c45a5514b5179ea1c15568344e0c2c8253
z45fbba4a6789e35e0ea27d8a5855eb9cf5a59f03ec3938dd2b64ef9f0dadd18b6ec6c959f1312e
z35eb725475b55f815b67d18241cb36e1161d4fa818cd30b509260d672e541b78201582340e1ce1
ze7c69248c187b84abb84b27b5f8009ed4bbafb150665857e538a06f783e4c13ad5502a607a5b55
z5edd6b14932d9aec1f7ea74471a81aa53e247b300c78ab3fc60af131d76f01d60bf943a1d59233
zdc8d7b6c213f8fea40d303f7582856fa422f1433e0603cf2cf2391324f686bd269d80f921360e6
zd2ced80db96329c261e477d0403d2ab474c819eb205c5fe34602ba5bf07ed5fb428701a6d893c4
z2448da40662f0a93267442f046fc983536e699d9db0cf1eaa595a73ac3a56af8f65c7a496834bf
zb9539339c3ac25f1a6059b7385638863622e93b0b7e6426e1da0eb1d68727d64d002ea3d9e476d
z3fe6c57d5d223634c7d41d37207b65b6042b0141f3037243e5214854a1988a9256d8b09d9d1398
za94a431ab2a0755f2ca12741b337fae5559e317256c8e975c13117357cb36b04cfba93ef207666
zf91abc42e976095db31d302cbe951a10dd7d4c2675ebdc6c012c87b1ae07cb2772d5fe193137ce
z9fc5120a312452e53f720a4c606b33d813f5ff072baabbd541c15bbc89b7ceda8ed600067a2f24
z9f9310dcbc38c8f76b68cffdc31a71f6be2316c51a4a8145277f18b34ddaa1de052151dc228bcd
z60848125ec62cddd2774895b918fea9a0cb9eb7b667d059f9aec553f8cfbe784810090adc7ecf7
z57e9ae935a846da950035af81ce53a2349d74d69e24de3260128799761aab9a1eff5edf6c2c534
z0d5d4c1c796a947c73a985c81c88784a85f5fa764e3bb1bf3466a89bded93d8b2ed5eb502f136e
zf5d1412fe47fc10e5f1df095e66eadfcbf8a5c3ce5fae1293aa51c27e8a9bc584b55bc08aacc89
z8e1c5a5c61559e627e468876bb3f3bec795f3333f9184595ba9688df595ac9b7bd6d30f342c4ce
z30b7a4a34673873c96c2140fd94c8e7e28018e814dd679af015721d03f1135a9c75077836a88a4
z8966e94951db388a9fb803ec83c2f2cd308f13bf73075e804720fafd202eca09d0e644da72ccd7
za43229e7f23a23704ff5b560bd01abf8bde0e1a1a751da5fa52265a3c849cc01448862ee393f07
z9bb5c9181187aeff0951c46577fc3dbf33fc90a45f3fcb74b2987607600f7a665b7d07333a7241
zd29a6726620244300b7e424a84014ebeda9ee65b4e5f5bb3b18df48354183e7e3510aba4c5dbcf
zbd2c8e896de37bd6158e5dce6f57dfdc8b9939baa91308f654ed24d69edf46539ddef7ce0bd0cd
zf2ac4b093488b688960a517ab109314b494045084014f04ba8e419a45594f4de0ea225f6a4ba5c
z414249719326211832a21b24ef09a7ad00925175a6e3558b206fd47e4ec82dac98d4a17f0e609d
z63e7a240e178ce961bb76b7319efda89c7ef631d4d7e3a5b89e4f90e369cb94c821d172dedb335
z7c65da017178247619329579712702b4c6f891ae6cb1e880623338178b7e7026d610431b214b73
z00fea4070b31a62b4ad8e5b1eed17167f260de4f357a1881372ca0ea0cc055c595dacac55986cf
zea97d8b7df219fa8d8eff808059ad0592c9b6423f65744057ffb7d126fcce16962a3a673c46cfe
z7ef840dff3050ad633faa01118959bdf7c674103eccfb373c3de23ac799b7a91f1e8768e781404
z9581b9854cc21306f59c69b71a58dfd2ab999f0476cbfb25a50facdb6130b1a0155481bf3df100
za556d9761011d4ea221a8bb2969e0d61cc79a3e018aaea5caaf5a9b8e967616f83da3205686b1a
z0389e42c7e070f3ba702151f91f5a13281f51c3cb84d02f45f94271b21c7e7c7c67e40b226d839
z559f45dce649e153e52f6055f04dc51166b605c688fcd96df0a9154e45d5d95861969a831af102
zd6a5d7cf4135fe8a8055422cc6b7bde53a514f8efb344e8f6c804013186bfad34d60b241fa5f1a
zc23d9b49dc97467982f04bf70bf7b302f709c956d98df270796f6098f385ff3cf9055b51fb627b
zbb216db451e734da66b86f0d9f0f6b842dfb4e172c9d1a529ec738205cd736db799e2b4251ad23
z46b034813498adf3cdfec8d18e80ad69a39bc8197bcb42dc365ab46dfc68637f5b71ed05f904eb
ze01273796b53b271f5405a4c0015600319971994bea33db110e98570686ef4dc2bd109680ce264
z5d6b207803cda818c0bab49c53f05d9fdb1e73a0ebe4a36c710693b346d8db59d511013b6b6f1d
z9d2af9fd507e828e3300ecf29f6e0a57610bc0cb4bdee66da0e40694549d73456403a874977dae
z5a2bd59062aa87e6a1cb11b101a1551d4957661919791c265797d5e8ea73d0ecdd259c5dd7efd5
ze0aacc71ac22208f6b58e23716f531f66fe28c6774258d97745f78109b981757847e58c3dd568d
zf3ee42b1678f21bf3a5b1cd3a37db59cc55040819aba67d4260f7628cb725d00efdc9d3446c91b
z5fafe299fa7362ce5cc1060cd5ae4cc3439cff892d3fce62816b816e09c3ef933d79053f2e6084
zc05a6cd14a0728263137288fe3bb2bb30dcbfd989055bef06f16dad116895bd69de7bcad426695
z29dbd6d485a7079f995e26ef5c5936140bcc930932ada04f53135e4b5c712bd8d41e6dcf2494e0
z87b83a457bbf17e3cdab51f991fadc3df3d9260a616bbc45815e55ed51e63b3c7dc1c00353a1e6
za7d9e7f10db572089e1bc73d04dca14ba285f3c1df32ac87b5965bb05f37bf3cd0c414a814b7fc
zcbe2011b9c8dd0ee4c7609c30b3bf1ebe45f358a7f68913612fe229f450e5aa124454ad6d30034
z5a4f3f4e8651e7ad70f9a5732030cb080ba97578e8f9d7ddabf5e55958c4939df76554bad50846
z423e5ab401e2631fc0233182d71dbc5e184ba3812b134e7890db32bcd34d2067dcc92d38c7eb3c
zaed8ca0bdd8abaf07e0a50ce7da2bd35c9e3df66ef0e23d1be0fa8cc3f5fb7c66dd0878516c900
z75064868702487991fe81ef7e252d651658247c4147e319781715220c935f1a27fcc227332bfe1
z08f8dc30d0ff907e0a7ac85d4f6931754a97b5fa04008cd62426b1c8f877ec43a1472ecd3c4693
z1162973d867f853ddb669a9a7556a175a186fa17de758b4f69fd6e2de93e936100ab85773d6edd
z26f392bb70084f52425c341dfac261209ae252c84cb5656c7459733e30450b7d236741bcca7983
z8d48611f976a2781cb2b63f076bf46771417e0663d905297f88398fd9ee4175c39651ad4e71778
zceeb595f9da7918846d2649a1dbd28173830c7d70d50e943e7dda37021b34b1b1fb1b5c31971be
z7420dfae0ccc938752da6c616cdd67a866f1efcd1b0ccb9b960683afff5acbc006525486133037
z2574764d763c01616de1a8186455e904de62fad77fbc8a31ee423ab719818ba221b7d04a78f297
z075b8a674900713cba8859e8b97e0c72c85e43f6337061fbc0bdaa08c147aefbf428ab9cbb9878
z3a6e0a60ae693aab449a8dfd749cc683746164c93900754b6436f7e6335a0342d657de1737a6b6
zf5cca90a0b40a3954c0cd15aabe889b68d2d840c485c63a51f1c5269010e7099d22f6dea1ea71e
z8498e271f0cd03311754c98a7a8c161fd96113e9cfb8ecdc0dbeeb0fba5486f34db5ca8ea132b2
z6638e0f535f4c8faaca5af40ba6de129358a1c54310840ca8336e5bc73dcdee10c84bd7f440dd8
z73f966bdaf71113bf448f3dbca244b1ead70ddc56a459342442e338626113850d330cba791de11
ze257e16e9e2563824e9523f0706743ae096d0d598e43e43ed790a2fa7653918a2d5d84e2d7e243
z9e23aecebd21cc97400ac1d9a79f75a8b412e1aab9cac0f6dd8f94378d5e003e18987d07d87e5c
zb479e5394f69684a1764d7c95a253b0f121d1b96b3379c2e52ca1307fc8c9c326aa8dfbbb5ea63
z7c06c519f65887718fe4382deba323f88551fb6f245a480a9b024bceda10bb705c567f87bf865e
z2e5f6e784d9ab3959415a0b861c80fd8edc5a08e49ed52d48520395113f045f45396f39467fe59
z9cf062d5867ed796f44091b16987e3c502d48cc2a9a7f028c3f4071f463b81789982c2b4ce9304
z41ab3f8288d5e920297c5cace3ff79a8a9c4ca0364dcac241add1e1cf8b857db96cea5fcc45bba
z50676fd2e0b66eb4e9b70ffdc6e2d13a1a5acf38111132bb941b5b118281a822d10428a3c416d8
z2c25c9b20a9fda92589f738ae5cb1d98e26f9b200274bf332f8c6b7537c395f0db8560e0caeff3
z4bac8f4a5385c5f404d44c5c794b35d2ddb26dfd4e4baec7c6108af0806eeff79f50f0d11e427e
z362c9f626e52d2744561aca0388578d8ebdad95f4b0b56c0f19e840caee043044036c6641b4be4
z9a633cb3517cfe363320c6bd356892405d1bb0938b56774c7d46d0407d50aa9246a3aa9c7f6a43
zd845651f9b01a99fb56eb216cf85f9f40730b9baba27e9248e9b92bbbdf75e00476cd8be300fc5
z04b4250c0d4b2dc68b2c5db95172dbb9f7329d72644a7b5a89dcad599810642844a7fa101aa703
z03f5c00d4b354e7a3f452321905cfb685ac69a3d253c64fea03be1afab2fe7ab2c746df323c177
zd2e9e8d726ebcb17fe58558a3592eb61670bf0470e44cfa0e891a55ef22e62125e979510ac0d74
z91c0d7f3e567e283b6d42e1a1aed1e7fd081669ec38e8c5622cf6ca6f443ae78060fc329e61fce
z14d4cfa27d61cc33abb99c23ddd7d8b758b3b7ee83ca4e02bd9a5716fab4499a65d3d6398b1f59
ze35f873d821dad7b1a9488ff40a82db488cf1d3a274d7e6ecfbd428577d84766e2ddbbc6bcd0b2
z6bd541757bb5c11594215f4d8ae185f5b9d8ce8080af5ba012fd8ac462c1e174d25f829d534af1
z1a53ee8a906ead31128db18e9260c9cf06ebf69587f8fb4c95568343e4de1e03304582f379f5e1
z64768a6d32dcdf365845de17ebab346c9c8e4e6268d9e0dd3718d6f43e3cf54e4705d35b672b38
ze1025941516bdc0ff35f72529388e69474bfa36063964fc41785654d74307d9dacb3fab938b043
zb90f2848774da56184a81223a7e2a3494fdbe07d7988ac41e26ee8bed75cab55c2b19d68d5e8fb
z2d693d6ab392a628400e2a40b8cc51f31cae2f5e50ac1df8b52ab364b533eb5db4c8aae5f76130
za9374cd4320703edb3584f0a561e5b6f3d50ff4ca480701ec5aee1ed95e3718194057dbdb87163
z80029debcd2f9e006ece785b6fa4825d43fe41b18910bdc708c9adc4794cd1c0f12dac5db4886e
z1120c6c4cebec1ce0795b057f8f2a68092dcb6e86f54de882fb3f05ca4d9c91bb8cc078651a578
z87c9c62bb129801cdd98be482bc512c523bf8a0f78f442a3ef272f0a1ebaa1dc931c886832f911
z41791d09fc4dc2e54904d7aed8e905d2ec0481d2d4097d6a6fa33ddf2c6d8f6c6e662512992f65
z9ca1ed54cd810c4997bff91a6e7487bbb64f562b896aec9e02bbc22b046eef52ddb140ff56ac73
ze5f08fb8c26f390052d192ff53951a6689695d0803dee90a2d0cb4ebe3385f15fe7bdd0bf05459
zf88cc7ee1aafcdac41f6485f6393c4fd6986407e7f0281af66ad3dc5ab5d222968d55140ba7c82
za571f8c80e71fc6ed0e5fae55f33012425d14f257ab0fbb10ac2e27d698772471c375dc4179d9f
z052f131e22673a3f371fb86382b31f7c07a18fe4f38fe7a7e4f87c389afabd3181026288991334
za7fb5032dfa427901c4ac9cf6e5f7e27677f71eaea6c3690c9ae3a4f2c6b2db3cf61985dec20e6
z3d3ed6a381a21c371c7b38b6595edcbb330fd967127648762346e5b97b2d37104c5707b59a83af
z8d18fc6fac83ec8fb80df3066c255bbee44ff13ea3e018d99f8a3fa793c329c510def347436213
zdebfd16193f70b8bf341aa24c7d9bf2c11f44fc8681d2d7695454f31516a280744cc4727cd12e9
z8ef46849216c67ed058d1d056e539ddb6f596cb759f45b43754bceac7fef2532186556c28c21ae
zfc24b026326a222fb6a60b7eb9f5d03a1a418f86d5a97986b983bdd17ddbcf6a657b6a011807aa
z7f61d45b10c91b98732a258a81b08cbd59b0c29db17f267df62f589a905ee7e66aa23c8c82e9a9
z95446055cfd5e957345ff34f63f896176cb75ed9edf97c0b6b7e317e83543c8e2eecd522b49adf
za3ebb6599f4bd1d58dea599b5557d626add0d24c32ac10e1f806369f3fad847348b9fec72616a1
z152edeeb7c2087297fc96d3f0481ba8f30860340c29e3e819b4a539ce6647b4a39a7adee054122
z20f9108d774c7b202ae358dd62553921afbecee94bcab32fc5664185330a3e43dcdf3922add2f8
z8b2b6ec86e9f16abc707dc42e56bd8ae5396aa140a8d1563149f0be6f4d29a7eab00b02bf3ac8d
zb47f32e14d13c10fa82913791b8eb5ace5585cdede4500add429ea98cf969b78de6d3065c2ff5c
z1b6d61d622fb6b74e1048a3db8804e6134558c7337827e5161f7ea687d5234483003a0d061c17d
z6d7ce26cbc84ec06c7982aa6b764f645756cc0e30439f53ad21d2a53f27e960ee36364be1a5a0f
z0136cb07e53f4be93990ff96687a82789290bbdb4efac854b6623085826f4ba3fc459ad922b420
zaa95019acec6b66bfd678a7482757dbddbfcfca8d45c6b4a2ddee4ba6d6d4ac53c46ce7affe3b2
za31e9da33b2ba354d6bf61f3d728b827de2e84e2bdb449eba4ebb5ab20e17dc7d479d70f592ed5
zee02162b2d4a07b4a9ba110aa8f739290a736dced77319fa2a0f72e5ed6fe428a4d01059a55768
zb34dc565c6bd9861b2ffc22de7c96f366393e85ab1518d4378d6c0c0e5d67e66fa730f50cd1ca1
zff0c60236fa693b8ace4bc54e2095ec9ff1b8683b52ac579970037b96510159b170ee6bad69f87
z160c948adedbb97f59420a8f15238fe8e2451bc2ff7d7085337554f78171c092b2d2d907d297e8
z478d8e714e81eac6c2aee96114f5d2a01dab6342e1f51dd7ba5c787b1e37b138986fbb09783d1b
zaa7030df968ae01284e904f8f6cbbb2b539f5e554fd41686a3c4c799bb307ccc05b1d43f0cdfb9
z4858014aa87d81cb5ff50c6dfe58e6162812703292673bcc25a1c984e87a760d3fb3ff34f4448a
z84c87e493e25732b8790e1f352993a5c13d35a6b5cfec4567977bffcd5f26b4cadefd3d8591b63
zeba85d4035e39759fd3cdf824e802c77e3b31e72c35318ffa3d38f42350cfd96eb6d31110b7b3a
zc1dbf1483a934c42c5675a91b8bae9e08e9c13b045fa40353b182b7c06fda293d4d46f4f7e3fbc
ze40e0b1872e19b2b0f363a509caabd556a443ca83400290141b8f4241e2a831f294fa5cd2e41e4
z8a50f6528345e26b66b6d5da38ff8d7963f40522588afb0010a64d80293ce3a3a3dd1673db0573
zf08956f8ad63342acc58d498cc1ebc557fbb99360185f04c95f700ae058b1a02a25dbf97c1a0ea
z1827f092b1911b22d0a7bdcbaeda983d47332ab2e7bc96068e506cbcbd9d8e7d5db204b8775db0
zb222db56179a9e781c74b1b0bd50a2527c5fa534491bce17ec24e225ba794fd3207581d94fbce4
z0fa672ce24005fcf1f24d330c3ad97e1211bedf3d7ee9e012bce6d2951cee25b47bcf2085ae941
z505559e2ff3fd0f06e24cac4d27ea62964ddd5dc209e16bdcc039c3e64aec70fec72ea90836f5c
z3b1fd6bb2d794e624a071b914e696c0936f8411029292aaf73ecd7688a5d282a0e979117db5a93
za7d9b01ed9ddc6e5dc48877bb100a9d3d9d54d6dc4d1a0fea19ecf4addf49d99775b555479ea9b
z60445c7e848754eb42748b4604c92d1069b28076c959cba9a007aa5b6629259f676bdd6c75b956
z7167c41d71d77954439d09c1d6638996b7cc84037658accee61066c27f01718783328c3c8b794e
z1bd16b387ae2220f0e9cbfd0477f5982eaae7060e4a241f06aab25a76c4b912bae21befdae7872
z3a97e6db0fd67983f0f817f4ceff79943e453f6698f569c39ec784d8c14f1b329ccdc1d960fa9c
z50403b622265cba3171c9e1fcb7d4fa2d09aa07f051fb779f0390f74ad96e0343a0f88b36335c9
ze45baa640eb47a1d2f738b34fe628f9f194b77707f5afe9ddb0ddac399361faa569f8d98f2189c
z95c132aeb5bc0b7ac98b87132f9d61bfd64c4be9f2c0d08481355b4538d4768147dc69d3d2223b
za53c34a707e2bea7ffda3ff2782e50a05e37d5320929759885f988b71405131077f46fbb7dfbbf
zba139c6679285facb15111d9bec9c54b62cc116f80df7c4a1576d1530edc0186c0d7ec4c58168b
z6d10edfb458612e971674687d9db9c697613b02c717464e46dd9a58206655d9d06d82165d76a3b
z51952a28fcf221b8a10ac0b6a377353d0e26bbdfc8ec5481a633952256c1eed9fa11c1e63798a2
z8e52d7b4d80549f7bdc874302e80748615aaa6a57fa6acbeb3c4ae1c290f95e80cc780a4c03c3e
z7803d68160d0f750db3642af1c1a3fc64124e6af18cb084de796dc11fd4729b85eca06487004b5
z1042f61de724e4fb44a6174c6b8f08160c090cad742d61ef19c82561b7905e8e2c01f2f601a663
z656b725db5f9b6264504e9ea5e5d31a63d361cc60058d22c93361b1a07e74992d990d9c7ce4549
zf83186e44c6dcc38f4293e37989785607adaf51286bd0b5d83b3d09a1f8c0de0e51c3ffacf140e
za83a210db2af00699526595f68748da448d4d13bbb720f109747c265134428096630c7d788ba57
z47a9c6b969b5153e9497810e391faf6a5426c24d8b65f4b812a068416513b6147949af41f6d722
z543bd3ed9c49a1b410d1ebc99465ca50a0cdb090928477e64336792f0e780fe94ea63635b7dd44
z12037008c467317497ce77513f05ccf1722584df7a7bf4c03f9760d396a3bb000b060d66dce367
z27f734d366beedea732d776e8ef133c4a319af7a921a56ff417a7a8764f9a9940dce7bc341d63e
z19066985808b8bafb43d900675c0ed55cfbdda75e8585f6083196ee804fd530bd28628028f6318
zb27d34571f3fad0cb7f3cc8497a2674fe80ca50675a7ab84cf73bb9d3291497b94ed404c93a3b9
zce6499e7730abfcc9dee326e4300c7a864fa7f74240e59022883aeb78a82f047641ded5ebe251c
zc03e1d7fcf3197a23ba0e18b3dd42c10ccc8d4240ba90e2df8760f0ffc97f945377e09115577d8
z2df887a7238a31ced51a6cbcdd9724b4cca118d252625376578fd705b77e80f4b6e17c32a6beff
zc96d1c33273c64aa9ec0870b27b23a1cc0f270d06d4e61f9abec959171c2e6d3a515b484216c67
z9cc28b8a47340f06ad197dbba342b996dfdfc4859654825f73af71231826383af31dba04fbd6e0
z428829eacd71aeda3ae7ff03b7ccfb83bcfc8495186e8c1a72185e9e9d885a7024eb819cdc59c2
z1c59fb168df1a393089eaa22d6f1edc1ee670470aa809fccf1d27f1ed9db711b54725303f1dac5
z92acbefd1e32b0b933553a17cc7dec26a3b67a908c6f507b694ddefdd1b19d7239f919cc86b29f
zfc474b76f081fb9fcbd916df675f3ea9254827dfac67be7ee068825f98aec06f98d9eeb0945747
zaf0a41e6aa31ef4e90a35c2202304756c9c1c4898c80a22de64c11716a365b4eaf20cca2a7322e
z872e8d65fee1ccdbe02f2c0695aef29dd2b1accacfdb6e521e24f53b4ef7b6a4586c5f9847b838
z088a4c6cc1ffb13bfd4009644a5acdbc8030e6220165256378a06585f608579579df72e02133a2
z627e33facc8f48c57649d8f071dc1ffb0cc3f4962e8bfb0dc7e4bb8240a3ea1a7780be9beeab1f
z07983b5992c9c2940b3c1753bf0dd58d5bd5fd5d013658bc22b036d4bda030067f2b1bfe885fbe
ze31f5e505728f9827a68dc591315129275e515bad9761b3a0eb684e5411f578c042707e3265700
zd4589c04d1a39ea7a48e218bba728f0829ef70c1a58c0c0400fc7b9dea3c61b63185afaabbd960
z63dec8a243118d6e5c16cd24ce468e4ad3e6ce82bb0d8419325c346400fd1f769c7cf3e0550508
z7a835538ce88fc49bea76dc3253d7345568bd569d1686bafd18c6376a1d2b160c05cf3d3af2b15
za7536e0dbdce0d60bf89e76bc27e09fbd1b6d18f353ad3c0571f6184495f3b1a9964b5ad073941
zc0da0b7d836533b9339cbe38ad5834c6bd8ae5ed7cc62bb13c83930ac2fd5b703fe6d56aa295eb
z69c02c73b6a5e9ecee41afb1fa3f4aafee022fc06dcc3ec446766f03129fc8ef59f270f29a9e46
z222e6c364399be1ecaebad6d470681c80107e7059c12d46be387f644782256e61a00d59cd73916
z5b7ea487c81c815c118d8d6af874bd8d36a4105b4d83bc799c93c0de9354d026d63e22b6ad6c45
zf106deb5850ea489ad49bea86942374c69412e02478a6d22841a4fa866f2592a871e074df37357
z72424bf3399b2fa7e3ab9080214ecd87d86fc85a33e1697916a2731726b5daa124ffb7e569a646
z570554a6e6acdb7f47cbf4f46faafeb3604fc024522216e43a0a29e403552de441a6d525fc21ef
z38dc6f8426e466e7eb454f60743fe5130464aa005715dd102baa8e29b07fe44570c36fff3bad89
z3805a58f59669d3a9e8ed387d79b74d1dd7d02761d84be707b67efc0eb87812d2066f50446e0d8
z7f9fff60cbabe68bc2c152b9120a5a6c2b7db4da4da2ff6966ee44a6a4945bfe90d0fd49f89019
z3ac08a920d79d56ee9c32e0a44187459131d4f5c5fe460c1349b77d72b2ba56e870a31af00e985
z1a4bb99b0b0d9aa940c23433e3e947f643198227d50739a08129d174d32518aeda0faeb65cd4d0
z63fe8f083bb07c6e7961c2ad0ac5f66de537ceb3722351423115d2743e872c3e551bb5af8e8ed9
z35614c75d444a33211e499d36cbb465eaf8a2b2c7a3ccaab2fc84280e866a68825279aa0836bcb
z09e80e3b693489cc94a2d17afc6c21e3b103d12498459e061c80ad79a762e9c24a93df2377320c
z63dd837ece9d752ee8b8ac014e614b57a34263f75ac77d12ed6ea2fb9b5714e437ac7ce8a25cce
z4d5bef35617e4a27c543d1edd6dddba2010f8b9c961ec6d93d6e64ff3a5b764c773ad796196ba5
zb53a7aafa9fc86aa794710fac64e2a811db4c61b13def123485060eeac9e476befc572c0e932f3
z6035175b11ce2805cd0f05747b596ef40a8467a8856e107092d1bb478dcab2338bff766a1a53c5
z951757882214fdb87d43225ea9d907d28038830ab43feea51aeb4709bc2365b4caaffa618738bb
z3b3bb798044c758b91ed4a9318926c6edd14e4339305dc957b982ebd79903953875860bceb29c7
zc7624b3dc88ad0587c8472a09867bbe3f1e072fa6b4969ff3e2f011bd1d66ddd98c691af41347b
zc7ed0ee12c5dc41f455045beeb876c0489441dd7454351fd9c6d2fcbaff402d822f83c3ee00b49
z47b8bc414af192a5e06fb0d5e58c9ba8321cc8648c365c2167b3105b4a71e7b18ce9403a60d141
z5b28f23c13739e03f757ca583bdc4335496f4a2037cae4fcb7e7d255bf53e5b6c64525536f2a56
z5e6671f275b59d0a20dacd8c8b30c2adb5963319b3d894dbd7d0f44e973b96532ec351ece596dc
z224c8a3a4af8bf636d906417669159f6e7fbde11d85920a5d774c0b50441af208a688421ea0323
z85390a28e136f47b776531929a2f4a97bec1483dbbf79be4227e2b90662bce4daa4e9e553d415c
za9f68d9f9dcc389261d2c648256ee03fc63fae4e7d97cafc55efc4a12155ef39361bbaa0392079
zaa1cee27ec44a3962b87fa85cfdd0fe3bedd475f64c839da95f8ce5d2a0dc9d94100f3b97581b1
zacb693699f216b288dd1c7cce41990f4104bac8765fb6d86e1ef544a8b888bf11ba6e3f0fc493f
z557c9769a30cfeeacafbab6d90da206b6c1e0b1f863147e592ea7541e6ee90e88e424570b1def6
z7219cd6e1e9fa3ba14c5451139a2f73a433d21b675dccd2c9908febca9357cd3179f1ca0381725
zd73b391a11f2c29a9b459f32272eb32c118b2c08890e7fa5411928d39e23475a11c469213555c2
z5d29bd8fa582ea0312b1b4b375cf76f8c4b128a9b4767a10a2f227ddea805bc12a20e6db5f3735
zd4ad306ae6a575a8e7a45d4e09d65a8c09948994a107431776ff53fb130bd4b5dff8dedd533af1
zd17ba01901fcd893a0837be79cfe3cc96d4dec2f41fbde8cbd0208b9d264a838d86312f195f162
zc74ee15d543164db7c599a970738b01e0e41567fc2cb87f57f8a258c64578f1ecec425a9e82ebb
ze0b4a54b4b9725d8d9a9e4b1a0aee27ec82ba657562238e60851de880660ad1778c59959d9aebf
zc10fe61f0ffef85bb8b376815a65862aa8d2fcc4118d0b9d9c64e183a8dd4fe793dd03f8bb4170
z01ffadafdec92a0d6fb3d5b58c55964dcdf2384ad1195656fbc1fee8f7f20bea95cb8bd8ff3b06
zcead23075a94e8acbb88016af7ec49369b0a3518f58b99b979f47582956c1d973484096270e98e
zfe55f0b60ed36a330315fdd15fc5c605527f4f9d7b0c21faf82707a0cdc86d86697cb4204d5e8e
z40c92133356f46efca518186ee13a453b84c85d9384db658530d42c9d8b153b407b33dee89041a
z2e74f5cd6b9c08ecb8785080f452fd68b250f30e63a65bf334d0fe793a1621370ca8e09bdd6622
zd8093b4f69069d31cda1ea51b322dff344cb6b85ea517d55dc34569b871b1e6edfb8151805c95d
z84afeeea212ed3e77f7f6b29b8b2668b1a6d929be5fac61c57a1ff1180232e75db97b314306a92
za911f505da3feb097e90afede5ea1d21bce8c256160334a3d60b306cbd25bfd7bee914da625f99
z561c13fb9e902bcca56e5e69e6c38581f18f5be27f9669260e707d3f46cb20cd6724a52fbb5849
zd7b5adaf7b609aaf9bfb6e8f078c82135203bb938544de58cdcfbaf20d2f8d88a928e89f98c8bb
z9bb6d000f4152571fcce7213e2131202e789b5f5b79d384d7c487cc91fb6ed41daeb62d5e4b697
z62db1c5cdfc630fdaee890cd87bbe3c2a21ef207096ce63b93034cc5df22612fedb32c18b14e98
z9bbb8204437938368a3f21e521516a6738dbda898c0edde00763ea5b26febf2dd42ebee02f803d
zfe3e838198194b680a057485c746718bd712272e8fab0e3c8cb38e45d4bf0fee67cbff09a494d6
ze571b518bd33e1fe409925e078c74c044aa8a02e5fbdd50bcf7f6733ef56f28ce9edb586bccd0b
z4e07140544f84f218228b5700a06d30dcdcbaeebab8e7aed5c23207b39095d9f26ffb61e2ce55c
zaf6b96e01b8dde33b9dbc17807a4b9c84a589c1590e5938cd4d14c40854e2bfc1ef69888024181
zcb14ec945ed7ff1ca1646b28110de7d26c8ed9e2918a5fd1b64311f3db200021bd9594c5a2bab3
z4ba0fe63d34d43168f3707c107fa75b84e8226eb1ff7426e089eb861ddf587d89105e6ff69f3b8
z4470279ea878fc92070c81b19e9fea0fde03f64c89b6eafcbbb36364f7497c6bafa8266db47122
ze6ee274d39ae8eff6c14a6c071f5215f0ab30e9f5db68ed527e2d274b23c49985a373c45dfd87b
zbed56802305d48e779c3750cd97ff612eb1f63d114ae79955b300a7931eafcfe6d7f78b2378d84
z5d24eced2a475eb10926850b0b5019d486e13622187af4092da30da71aab04b34254daa09e0abb
z1ee240e51fead679d2fed56a7a2b6872e7dfe65bed6ed209d1fa7191dd9a78895b127c89f00a95
z949571528af25d50b716f8998ab326e34a453cdd11d73611fb26111102ddba0db274ef0295dd42
zd695a57164b734bf4e8c661ed08cecd01cfc64dff3296e9fe1a7c29a3ae644f1c83fb4c6145900
ze0ccd20be8b083ae5a78ee84326a7fc7310deba4e33118c076771f61a68e9156f4426c0d8861c1
zee54a5950b5270264c8aef47efe42a6b75ad7f7875f5fa590c8120cf12ea264a0bf5b08039dff7
z1cac275a78cf4f6ffd425ae3f695d94e41bd93f2e36e06e4ea817076713be4ca4833d6345040a2
ze4a40c257f34aa5ac402cfeef05f9bc6d1746c97a12ce4fe35213c16a001b13451e1cc41696596
za197fc0e345da3258d2a41cde9eeac0fe7fba214e1b4b6d34feaf9bcf701fd4b6e34204a9a4251
z6bfc3a6efc2e46a98a45aac02ca9aece9e3080e2b14f5680bbd752fe52ab8cb249f8a6245b20e5
z2c93863b34c9c9d0df1f69cb5db523f3e0e3bb83f7e51534cd79bec86dce294290277344f74185
z83d20fcf1a95914d422608b229c7c50de5b60f30c5e71459231b8e0574d9651d4821baf2595f51
zf513f00b1a897393d09ed7282faeec82c4caf092e79b3923a97be2c6e1564aea91577ab02d5f0b
z498aa338c1df7f2d50b02c8d24548c5cf29c187609948e8a9610dc4b0ad75241b02b686fcf372a
z81614a385e9bbb1ed58e90d0e91654f5c17ed689181d624e045f4c841c5a9afec41384000b9836
z1dd7ea63baea8475c3ee6508972957f4cccd04166d103fe9f54dbbb75ae690cd69b89c22961dfc
zfa3b14d7454b85182456618f9505a89804b6123686b8e8b8d4c542ed46f529eba35dba40e7be1f
zdb71d564826a82464ce7d6e844ba78ecf6472df3540f72ae90b3d7b90184023da0b5fa8df81f3c
zae01acede394bd46fe67499a5738c51ec5a37f3bae948616ad86c9064d056214c32f00dd937631
z68666f4ebbe584a9e47a3004363a430513e96657e0b410f28fc9a33b1dcd027d32e4c57861b65c
z2032a2e5374b9742467a1d151dba45562c58c94d32e665480a9a648aec23470dbc8475a059d5e9
zf494b9b240184aed2a051c3e9b285bb49e7c7995a4348e598dcf2b4150f4fdee5461e0b9caccd3
ze3e81f290f82a6112f92acb6ddfab97a22f3c59051686b25bf2458b31551edfc67916e6d65f865
zbe4e413001357509c57ceacecf15a69a354031760598a8b3c4e34e5212f5f30a89c1007c48053c
z5d3f7da40956df18db381638de95ef14f7d90ec9170c7c9f18bec0bfa9cd8e7f3422b81ad4eb11
z429fecd228e4ceb6a619229881c62d38ed6f3e149ea33ce45a62534c1781ffe27b550a2a27e922
z19971f46dd2f0028c6806dd98cf84bc3bc83cf1f39eb34bdc7689e3de3e6fcaf059adbdac4be00
zc3de5762b53b0ae6bdc57d0ed814c5dc7eb28c0327b6a1cb5f993c58a9de80508ab48ef04f0304
z5317eef450750107f6c31d5d9d6fd842331191eb11db504b008aa0cc0c2c135b3242c16abbb00a
zf5938f12603892588ab2132c72230b1990990ec6605f9f5eba28432f6c6f9c9d40b2eb7b72d50b
z0e3ea71e720ef6e5e441069c1bd065f1b42e84555123cabe966a7de09a4b3ab901338dfedccd61
zd134d285776cb0c03d4f80b860cc116ac342b60bf36e5b05f523a7103c41ed333c276bdf26c796
z0db44df35f18941829a76b5356a277a96416dd2c6a1f40aa3ba6d9b641714ab7996ba06d0d5c0a
zda659b0915779289df2ddf33ba1210ae15ff60c2d2145dc9f77016d2dcfdbb5b7cf46cb6ae9f38
zfffc28f1e6e9c096817cacd3982813d8a26949ef891e25f556c732a6afcf0e9d6a7ee5f931983c
zc7685baa0fe8b374b596c3f98cac013c3ca136b734eea91e69026519a74a8d1cf45887b522f95e
zdcc55a7e93a8d1448a81fffc2ac94a29b04e101b0843c50b2f0b3ed56aa3a020e376e4af5426fd
z6bdccfe148ef4755156f89cfc698ea9658407ed9b970d70e7f93f7bbbf2f4da087a3f07aa367e8
z7ac08b99be1e42376f91f9f28e3d69005e2385f4d846f19247b8b4d3bdf8c2884a7b9c3b4d7c4f
z4c217c565bc9d0c804b6dc00f919e864d64ea4ebadcccb6c3db9df954b2a25d39ede981d98253a
z2b095bef64abcab2b01b0a4cd37a2bfe753c41645e385f20cc5542607935b48619d1af9a3407af
z8d4e26cd62945506922a778045bd95283bd6956ffeb62fedf6b1bf021b7a2a9a7088674ed59c94
zfac49884923422dbb0d7a8541446b3aa2e7b1d9d1576ecbf1b7baaa0acb8193a2782abc53f7fa8
z73c3eb693b1298099a2bc3e8b1e1435aa91a7cca60fff645c178c7f806486c63f6344ee7fe1719
z944fb1f6051181acb6f25605ba66003eca6c7d2e1f734c420d05417c9a2f8a09eb45d4ae3c7173
z59048f74d8e405cd6f22118b773b5ba3c4854c34aa96b19100def2513a1f122e176f742c20ec9b
ze52c008e6b2e27acace8431b2c4f9de24c0c5804711703837a66cf10d1425c5b87f12e41770219
z36dff2a765357bd5c0b8aa4e5b89068ef8593c4c91d6861f030d95521f41d776776ad242c5f52b
z334636cbad3080cd56fe6f60f35e7a94ebd73aaae47a257c47e7e260055e1a7683019eec9fcf41
z264a6588858964d406f8557384832ef750710127969bf08497e11602e250ff7c650f2ecdc9c0dc
z9be43f278350c53dbb7796b7a1b75c84d8931c4fe5ac5b2642051723696c412ff0c22eb984df3a
ze867c64b1ee902a55fad86686d973c8d2e0880c058a4f60469fe5d971a81710d9cee5dd9bff2e0
z06b0876ad3c5421d37661f5a952e4c4c65f76a90370e1efbf9078171920614795593115aa60835
z092547f468b3f3dbcb6bff40257996dc45208dd641e54e16ef66126d0007503ef2074bdd88741c
z50a665d7c3295874cc136370002be183493bcfda3d85cdb63c3c51a73d1dca79fd4193c0a59029
z71e695edf77f0edd817ffc489248be95fe192ac5af0403f95075182bba38f5e6f9f78803af5044
z739600a5b061c4981ac7aa62eaa4d3937d8191c76e0997d5b35ec05c1dae2f052eece59919c6f0
z0d549fcb8fbc4abb78b4fe64faafef524b63b4569c22df4819207b5dead73730907b0f8b5319ce
zfa7cca70664e2b0dc2780832d63e567badea074b46f733441e7dfde931df83fde4ede54eef2f3e
zb188226bfd6c37f74278ae75633b6d153bef4c491b2cce67690f570a96e906e2f0f5f506e3880d
z0583671b59c860d0060a4374e55b5d2e42c0789be844e87bf2aae98f76919ee4e36ff5b9769fa7
z052690ded8228e532ce28a064d9ff6302f7757d81e262a1166a16bd2f04e5486c19bbb51af7535
z4802d19f10660a755019f361f0a85782e0da6c86e21a9f05aa26413802697116b22a64de54d868
z9cc374c5db98f8364597c71eadf743b92bcb97de8a3904276ce3f40e3d3866b43355b4acf6ca2b
zb7050e8b3c0d503e4e3a989fb91eb9d98e47e25841dfbeca987613ffe26043eb392a0135f24efa
z99b0dff3b5b147f4d47b97f887ee5d99ee316f17a45986cf04f38cf6556a2188c03f4195bb1030
z171f52f7d8c040f644dbd5157297d5727f4ed06d1b2dfb99001ab615fc87efbfb70aeed56b31fa
zcbe7e8fabce0c1167f0e615a315d2a6272aedd13f92e231aac47067fdc9052a88b9fe8a723993c
z0eb33e43a0d4f8b8104c3d13bab5a98a76279a2c28cd6d99dc59d45305addeaf675ac3261c160d
z2aa9a2c4ae21bb5936f285d655efbc0475bbc7484d29e83949b77228b86aac4b21c892756d6cc3
z9ca8402416bfb14b87594c6ad7c511c6cc4a7f549a57345dd72a902eed4830027d7e53305a809e
z6fe9f5ab7705065e9f2b7528b7ad14f012e942d5af29e127972354e715423f1da2b39d07fb47e1
zdaa21b60c924be88e46f2e330589478f2ecbcce7611b927bb4c3f4c2144f5ba9349bfca5cfe53f
zd6e1e4f94a8182d055bc4946e8547494aa70e913b981f47bba67c99a7583643c3a1b226a520fed
zfab18509a4d53514bb3974eda8205783d1adbb346e2a5e9ad5ec1c0c17d464936e70f521b5c05a
ze76e0d338a5566ee4c1cc0826c197ca5d8089e6c417c61acaedc7e9741a9affa91c0aaf7860e38
z3602b73467595839e5997f3b6e20ebf7c5a486b2b665cbecc0bcd970cf8b7c7b478ac8ef73b656
za5d2b65d828aeee68714bc0211511f14974db09e2f9a4a10e9374a8f4600e7f0310f02e66973de
z03efff6a9fe1c4d0c4a106bdfc7265f7843830b56394e5dd4dff83fa38995e3deec688cb45cd3f
zce93b6030929b11d60b9076a266c277dd63023e7cdb6df0e747422b32572007a9f6b5bf0f60a49
z143a7119f6c81be5109b32a0fefd28497d5234d11e9878d5fbfef9c48d7bfffd7cd79fa2a1009f
zdc76d6252ca5683c01c4f89d2086e9869855b8ea3cd54f68cf358b21f92288b1f725600d8f41e0
zf57dc022f1596bbf1533d2cb4176cf5c06b98b09c705c774f9c9deebf02fedee6bafef64edf802
zc1408b8820f3f5051363bf0cf5bcbf98f4b55251d6d5096784a17605a0a76b91223197a45e9721
zc42f9fb7b3a285f3a078fc008b178d92e9f3620d9dbef28dbd6443aa72711811722c67ad65f630
z81ef05b548ec22107fc9a0d18cd1c43be3cf07a8a637043aed6a48a0024a80cf2e89568aa404eb
za995e438c2a583cf204db6b51ca94098dae1bff345ac31a99b1e0ecba5772f5dd112e5e26765cc
zd6838be35d1b6972917a4be813f19a84dfd5c18408d014007b4549a3c417e6321b8b151a87f805
z7c32f46255fdf01c29e64970237c4c184936fe3d72190a8fa50de7d84c1f3a06e7aedb39dcdede
z34abd98268f1d92cb4ed3ae64876a6ee3e59f040dba1dc79857d5518b0f748ac8a70949f7bd9fe
zb27c3c45031aeacd2659f54ad06a3db4e3a8c9425ae12a609fa745c55906773be60947c2c84294
z75b1b4672293d93154878bf681d244bbb775e3b4c6704182da6e60f12d5055762085ffb23340e9
z98abcb9a8f9053212fcb40438ce4af5a7bfca3a1695fba3e4a8cab20dccacfa346bde9c0130ba7
za426d89d01f38cf1bc900a5a7819680bfaeac7f5990dcfae21546a2914f2b426c9afac075bfc00
zbbc1fcec5cdc1a95326d7c3ff74794b45b9fa3a40c0c8803c0434cceadd1216d0a46d33cee8390
z2a1d65f1a39bda61aa272c520bec3d4d7c43391b0ff7b63636fef1710bd1ed340cf1430ba8e4af
zf81aba6cbf1e0234847c5f8bf90e8baea39213f286e338c07b01f9519bac6234ac41f19a85185f
zb31f6e7c992c2747db787852e43d49a9d9a644ca81ae3c83ba3003fd5ca499af82cb26d65a7ff4
zbc58e26c05168c0f8973fee435375b817674ac35a243424e562c007c167fffcffdc018ca9200cc
z9861803be45bde787518f2300c09164e3a245f9c8578c6a5bd700959d3ce80731e033fe2ab1178
z814ebcdbc137a4e8f2b773ee00a4cf417824f756e46d63139e5e94bbecb2cca1ed568519545183
z1bcc65e15d152407f3ec36fa2001a2ede992dab66d6a317d7cb1dc907a0ccad624052670bc5a4a
zb6d1b8e0b6c085978728e8c75947c10977ec886d516f860d961f6cdbf7563ce509dd4674a7ab95
z23fbe9629e718c604196cfcd0cbf64f13bec7bd33d1472c84afd420c2da81bfe263234ff806c73
zb16b8d39acc0a523fffac1580767f3b51afe7df69ed667802ea13f3d9b30327ba6c856a6c4c5f4
zb055eadf63c5fd303b1b5d84078d82c03732b34baa8f5f6cdcc663d15279cbc9b1b0dfb9423f06
z25b2e03abc35ac61fd4e40d4cbad638342f35b633b9d3ffc9d37d9bcf9e146b6f35d8cc6a9be46
z4c850eee0adeb356b0a00d35e7a61e1e0fdb387fa4656f325fd13351e40b678f0c5c3d311da454
z940438429c242169309c8fc5a5e87fb943595f957e992a608c47fff843b22c4c958d6a2b7ba68a
zee29f90327a1976ee3978965475bcebbcaf10be31b380352fcdb768e83e555871f35ae78681da0
zc5e60c7582135d1c0f5ab4f0fce34258435e70662e22a51128592f26a85f66a43eea04c1458808
z4cf499966b397e30138b68327e343ebc8f8475c7c1b85146b53dc1988f833d70d75aee0421f969
zea0c437018030fe74a84a2ec859412ad322450397bf1f267d5d19206567bfd44927dc7a2ed2bf9
z17a05225c05df452eebf53f2f6b841c8ee39f83b6e9e876d3b61a7030088c3ba04190a64c9f925
z5de4fb4edc6166d4c6f21244328817d6cee6b69dbce4874523b22dec15febd1bf0aa7a335eadc4
z6cbacab220f54a60faefe78a0b984406ae8b112476db33b16166400acb6866f22bc2efb3810829
z8d859d4f9b0f0f2c9d1faae53232b515bfd0e13e7aaab94e55a5a357ac96cf84a98da5966dfc37
z45a66efd854fdfc15d17cc3db45ba0b7180303a24c1895034867a890d7787444a1d042ae757157
z95330c69a5f303d548e1ac7700c8a83a1e89dd07d099cb6bf6b18059a1302a94e96a3d70424667
za53a0aca96f2402cd1dc30e33373beeeb594ef743831d48300ae4d09850d9c9f23ceb5643606d4
z074cbd1472948452f4bfbe38b9813fb4e20a678868492cb9b50efdb24d7fa3f50df024f69d2079
z6555b0a90bc42e536bfb7f898a9a737dbf1a6b84d0447b85510ddcae88c11208eba025ae64fe0c
z31eb52f94c347a4470ebf286090c79a40f69818a040e37d9c70d46087b91e09f9a9286d4d925b0
z05bd2dca54ffbadfe1edcabb0dcd1f4ddeea27a632a4bf6d076ecca4914c95b7449e140d408faa
z40dcf9dcc3a606330554643f5a7659638fb1ad9f455e9c8e23b67f80d6a435961bebaa95ca30cf
z30af33933a1d837837c74f843224d7cfc7e8b8e243919cdb7a033def163a225bf05ca345d9d80c
z8401325c95988f28fe4143d9280adcb9821a6284b19787aabe007c6f3037b13f74b20c58c48283
z730195df0f8d24956a246108d05b6f6303010fb8a30a7dc8299fcce6ce692b6c54af5579f203e4
za99ac73c9b1d627675b4ada731d299ab1043f9d51ff5f9cb1c010d81bfdcf3f643bbc94ed5033d
z573627718156c6127d0e34e7f43930d885b638bf1d2e956dd36333f44048d53b77dcda4a3e6115
zd2cd26fd3d48ecfc5247ac98999eac0fb84555f2b932cbc93d553492648f91b5818c53a8f2b5cb
z0eee255be15ef91d568233f0719a65f6012eb5759013ff8c4d0199c1269a86e69ec71a372012a9
z02f570e0ac172f60d44d30f4e51afff3029c780fda31bbbbbac65e8a81c6ccd75a1767f9b1c4af
zbae113e9e3ebd450081734d0d3677d6640c5a33ef3f3885babca29dd999b010fb26a1bfac2ca20
z79729f960ae659f010240ae5b17b9e4a1fa605480b5b7e3b5481a86558920574ab0775a895fdd3
zb7b0b29b76264688c5d5aff4b1b81e7db7016b5da89a556a9b8fe3121e7e7f5b7e646ef1a8f235
z5dda3dc20b2cc7db2fd4a1b37233bd657d1c53e83da9f6d5d0eb6205da2d03eac38bf33295faae
z8a207008d59e9a50e43f0f9a215311ef1c7bcba83cb93c4d35a73a969bc45a5dbb52fc0904fff4
z7029896bfc400e0cd8c199154acc9fd980f1174657bb7603484a8e0e7c4728fd08dbe43c85378d
zc8ba818cd76fb5ae51e44b1ba952a2cbcbe6c9e802f6b8caaf67ec297d1dc5ba36688bc6f9e41d
zc3a29086cb1ee8ae96d2806b3aa59f521473fa23189f6d014db0b9758a22d3e2bb80410b133f8a
z3b98110a9f72d66e3d20cd62a574fc1798c970d861687990cc149a73b54be5616382eaed83c83d
zc2df8bedd94a3a246f94805a626f0580a824f07cf92a0c3faff81a7bbdeaf6f35efee0cdbc2a22
zee2b7c6c33c91fce1e6bc7a8153fc4a880e6fbb96adb738f5eb5e13794249bbffbb1aaa7437dd2
z2f3e90ee15d255f4eb153ff68ae7ea923a82c89c925874c38a1f3fa285ed458fbc952141e04602
zcd555496dbc02012eecd6818b48fcf04565f30388ad88258470c2581c202a6e090c578f01bc3ea
zd72bb5f8bea1474a4f0bf7b5e31f49cc1021bd294559a7a47e04605a82e621258bd881602e3755
z027052b6f0e9e729c9b818373e961fe407b93ce1d9536bcae31c8e74932f8624eadacf4747fe77
z4d17dd5919126eaf08ebc10c09b9a198b10618c8b5dbd263b9c92b48f3de8362438f32da471645
z9d9bd017ef016831cf367035ee6964007c25e458f3f6e3f88a2413d98c1f0e5ba8b73833c12354
z5e2777bd5d635459e6e1a9dfe2b9de8cf947cf2105c7327890caf56aec65461a7dc8c660e8b04d
zcda4b793728114aed748d3bc850bfd52493d3365640e37d9cfc107a09cdac2cf9272fdd9e89438
z5866c74f192178a9957906d1f9b706d42db2582198e6df66379e89dafb8af77e7e6c32c8ea9b96
zd5dae7c3f1c5c51e0be17baf7e92adc27bb4264855f8f984f17fc01842c2fe847bbb694c84ae13
z31dc4d4bec43ea1a9fd92edb4f31342edd00d43d90451bd27e512d9269e017753c159ae1b0c3af
z068ead0dff18ac4118580ed9330e888c1760d871ebe5caad1cf99204721322eaaf3df549c8277a
zabc923b84c05ea83768ce2a7d83594d25ce49fa143a8ffb0388bef5e8f85371813ceab0ed0ca15
z419250ee6226777be1020b2313027a4bc2bf88e6a37d441a5e77e01aebf3719c00e7d0448d433f
za548912e190135a778bb90d5be6d0843542aedd5b544f95564ba4ba62a36bc41e15d04b567c2d6
zc37d9406077f24128ee575e2ee2d4bac287454f23d52f0ef70e65c75553f3f2864911a742de052
za9ddc0d6fcb2f4b28c35f9803e5da186fb83406115b73fccd14fe5c0d3ed334f60175f34212016
ze42873f95bf7ab6de0371440bd5fa24d0f17d795548ce4e883a135037cb23694282c860a0a79a6
ze1a9e4687f0fde4008d82329b289082d80357ab24bc5d15df4d28c0465ef90fc9629429af7efa2
z871a118ee00414b6dcb1aff39732e4480e9503dd21927c0f14ff8e9a1a55974367c2cf6e9565ad
zf3734af20e021e4f9b0acbc91b3f4871310eaa98efac57042735a47eb095500a49103ba9a5045c
zf13b25c6764d094db6b08b1853f1fdb57733cad71d377caca282130a0c56da851d5a0f8e4a0e67
z11f691fe3cc3137e425d43a1e9b461bb066b5bcb4e96497daa41fa1fa08daa76c6e25c13320441
zd1b35d9a7bfd07144f0050cac8d9d3bd669a1d8f68fe1410200da09ab49d0a6c443769616143ca
zdceec0e55ed98c27d6111be4e28001bd31e4a4a8286aab7ebaf548797149d155ee21392f3167cd
z40a2cb3b918a8f05707ba75af15a8970349e8b2fa066b7d7c6ba4ff5f56009b74246ceea6ee865
z8bd572f4e98814604ac6c113094ed4080d81b4031794236b3b3ee17cee7aff8b2db1995bea9450
z01f264031c5e01e848b64b925d7434c0d0e9117e9d6f5ef25d1965c9824ddbaa385b9d4686dfcf
zec20ae6ac7e4fddb933c94bda7ba4799790bf7f1d7ddd101d34aebe94430932dd1bb5565a59763
z81003e30ae39ef25a50c92c58fbcbeb5eef86b4a2f5c5d3d4285474a338d1f95bc9ab1b12556ce
z7bbf0c76e95d99a5aa9c2d344ff2a17745ac2054d5838cdc67d937373896f1bd88892aa9edaf8b
z3ac1fbf9a9efed6c355013256d755aaf02020cbe0a26d280e9cc180de02c7affa95c7fb76ffebc
zd5013749238f9d0053b732b00c941baa3a10d3d4e536f51d93698bbc161614f02800a95dcd1758
z76ab526d9f34d748c30d0686a41ac38f9fb9f4154ac665fb135d22f6c43ec27307cbc725cdfc04
z519a5da12dce7f8a8c1c3d3bef1440ab25fb2d113c071bc80a0665407ff6971158803873769c5b
z41c1d722ccb3f4dccdd8ba88d1e8fda43a85026058a002b367abf7a1c0bab17cff51d8bc77b96d
z5d8f2b1d90241b9ed2821be55e1ed3d3233a401dfe871dd440c6bd1cec33edf016b7f2ae7f94e3
z9c24343047a03a025093b07c76e58869a1dbd0bfb525b580a95e59c39d63696eecec7d7f2c5509
zc7f79413f754e0eadec3537693751e7d6626ab893c011f52643cfe305da5814146aa2668a3bf96
zb8a2fab8b813bbc01e4eb5b7af86b02ea6826161435a74b109dba46b8326ba7ba0e32f841002a8
z1f12e00baaee4b495531a49388b91a568c58ff00fcaeb86ff9775ba690ce202374aae806bf39af
zaf59b32316dc5be6fbf5ebfc92528ac7b35cb9cce7428ed2f62d4fc18c4e45c6c568c7f89860d5
za4789b741f5ab28bc1a71eadbac6d1f4eb4389e5ccfa6a23fc94795e9e1eccb079f3962226ed52
za83acec65ac107212b388b230b7164f9619ce3f9b00b7b201a37bbc91c1454f0b2d7901da74d03
zc2fbbc6a21ae55116c8886af26946156ef896326b309bc8dc1b907771b7e45b31715fec119d18d
zba6cf6d686f7f025c538a0afc3cad8440871829ff38cd14e7c7df7ce4e43f07415ad0ff2912e88
zc32076cf41dd9556f2666c183afe158846afa8020e51adc5a0edcd7e24282611378ad8e80fc22f
zfc7377a65eb1146b0f93fb6b6f555d0a2b07681fd8e7394fe58a27b814bd855cea38e5fd3f2bd7
zddf9748d0f167507dd0816de5a671844b5c36033affd066fa0d7c23cd0921b4f5d731c57cd0975
zcb34272e7ba1259cee529da99a634392e2f6ae97db6903c1e667ee68217edac9f50ee30cb5971e
za9fe663ebfe186e9ee480c1e75303f92d3be3c338bce38af68b11d1d8acb832ee100a14f11365a
z8cde285a0a8931ac3433099bd2c8f1c50bd3006ed96d90cc227435b5583006725984c38946610f
zc715c1040eea72fee5c74b1809366255b036639cbde0b2b07d68814c6ff2ee1983196d9c9f4384
zd6a5f26b97f0af77a63ab93eb31318e5ac5c1d051a0cd21cdf3d9b3eb710053a8b7c7655ffb561
z51330b642ec2193a65de025ffd91c290bda1521dae5e9f3ca6a150008f3fce96c9f2cc3416946b
zc5f7b98e2703815ffa1c9dacc432180d3be519c9ef871822cec91177bee427e0512d1302f9f8f4
z298dfd9a8bb686c181422d6039b077ed065dfe162fc9ada79415db955e06690b6b948b2d2ca057
z0891a998123f2e18d59549fb230da6292b91edb0f1d09db0cdc404b05bf79ddbf5a51ece5983b2
z778ef9e08900d0f51e2706cc6cd1b38c7dc9722de22da55cca35a1a090d5bbd5379915d55fe110
z942e908634980a4139731665b0798b3d7ba7075d46a66253678ac43b8c0905b53e2ed6f651807f
z66a18e3f5c6f8cf7fa7ab9a92aff438f991cc53bf87e31846d33fe8c25f80689d9dcde08e1363b
z90e1711b5215a9949f1a83cbe730daa2ebb8d418abf555ceb7576ad782435c31003f1debfeb5fd
z095da02eeebf9b5e1aa0611dc916f45b7a26dc746075d586fb63272ba05077ccd35937acb77cfa
ze09aaf1c1604bb19e4f38bacff743a6d31a8ec5e8caf0b1b7c4195801646c12cc6c046f0da4c5c
zabf4f858d842eac1e69e8cdbed764056cf81e1b43dfb88a01ffccb521545f7cd7f08dd4dd074af
z004141f4850ad09c18130271b0fd792a5f49843dab2e7fb67d634c030823557bd2f3c18bd3c42f
z534b3a22f49f8d003be1ec5c6ab6a593c3a1c207b27c71705b59e6c2ff09b40a09b6023210964c
zb5fb86185a879e37e62f266694f1febb24101f3a284d659d19239cdf89479486da95265902f5d6
z9274a76f2620cfb12466fc1d7dfb599266cf62f315b1bbb25b35d8dabe871e6828eb7922152c14
z2ffef82bd07340167c56f225511e75874e40b21e59dcf61784c6fbd4d4a13f808c496ab625177d
z53c41728334b8e93b3187962fa613801628ed8ecc0fe6a415b6f01412745e5694067501c654bd9
z7db2af37482da85c760cec6ce0ad818de14757bda09f2fbf3fb8e749dfa88559b035071086ae6d
zebf7e5ab91430ea43ac80f9fc93047dadcd1ffdce0fec227f430cf534644713d6378f98a813372
z4018c95a06d1399a1155fd097acbe40f5b1087bdff0412c9e2e5bdcd056805114c37e7c33c6ddf
z6fbc8886737b2d51a5e29e2014c15bd54de149a17051a12c3ada87974307a1180966977132a30f
zd0a15e2a6a95c4786c095470e1287b3decc1a4026ca22033cb7a49dbd86f1f47be3f6b5cd9f9ad
z9f6f830346b2d5456823dc19cedf5357bf8b2b02c324126e34246cc0d7b580a7b152dd6ec6f100
z7d4f2f7a5c85be6c0dec05008eed8396c5ab1d22ff643284fa92119000c083f896d51df2d13fa5
z8e7f877fb8bb3ebef6db2881c71e16c1a648718b98272f9b69848c80de1a11170b561d05b7bf61
zc9f9297e95daa2b1a74a614c4b580b8f16a581588b407ee0cc29f8ff0f577bed6f1dc627b86e69
zea5e2da0cfa5900e8a435d7c3fbc9d16676a67803e31db79e2248d2db49123e04519802547fe49
zf6455c06376ac4a7301e51175313b214e1f448b62b51afe20518852156adc73c10561dfb5c6ddb
z29c6fdb575ace2e628f9f9b1fabaf453e9ad17256c0d944b82a52fefc929ef5eb1f58dc3c7f78b
z670d049d4f42747f8248df660942447d6ca44534a8d5826d5c2b3eaf4ee035e9a58d5e986ec939
zfedbf2fa68828c9e96b274dd3d75413c8740a98f4028fe7188df621962a15bb4bbb9c09b75e3ee
zb253501456ec6af3c6ba88c153e4dccfff12fae03857ff612a89840837e1bbfe97a93cf5c98952
z6196d0a27dbb0532855e95dba2fbc2533a2658c45b53ae2d3619238bad9b4fc081e8f5f65adc64
z3d4f689df3361fdc73d67044cfb4fdab539b9be09809a049bc6d16ba851f72db28334896ae4693
z24d2d197374a4e8c217230afa4828c5109ab188f51b1bb2d6e4c2033013bc344039e403a62c947
zfe5d869140ddfa77e936297a3ceb118a53aeca603b840526e9b48866c5681135698722be0a27bf
z63cd49adf94720312554d046d18642900377b82ded721bed542eb955a4762c6b1fca4d505ef775
zeab2342add2b39b9e71a2be3ba50de439f6f679ad7468cbd0142bc82d85ad80cade7fe6903a6e2
zd09d803d39b404c815bab112c2f975179473a25321ae55ad96e382399d2526182a0816b3b7c82f
z846c542a4d95c7583a304f6b77b27e973b025a53018ab657dfcf2d3ee86b9e332518e1ea14f2a6
z8f5c87f7ec85b44ed69909b4e3d7e03e700abf91517a3bad09a8ca9b2964dac949393f708d7b10
z6a5b4119efbb9067237f671f58407409c9981808686d94224d4fb5889198c3e6c6e1e93ad08b7a
z5ca4571edd9baa960f31b9399eec79150d27ab1d14a702105a1ce013b26637d21ad2caa82f7f0b
zafcc8d92eede059c67228ecf5e18eff88966525b66233b9aaa653e544a909bba41760b979a2f36
zc018c638c4a551f40b73de5306335b0eb8bbf29a9eff186e1ff72744f71d310865f52767042d18
z893a141b225034a2500bf331d1637aefc9ab446371b833ccc5c6930f92a766fc47b4114fd89740
z374e2bf1980cda1df227dc0c677080372e266f977a3006995b4da6f463cacb9a257e208d424b20
z9326a3588e6008e38dcbd23e0d8a0c4fd5f29d8ce3ab2da540de00b57e1dd7e5c856e1eee81829
z5c680f096bfa955e58373e4666894268a8c4e9b01b96c6dead96b8ffb8b5982190f552ba0dab6a
z768589ac897dddee34033c0ce4a9eb9017808f33273e36891ac02a685fe02c25b70e4d51bc1911
z90fc489c297e2315a07ab9a85d683c0934d726805f121ba9fc26e6f4817be74b5df4e37ed7cbc4
z14d6ad92f10333bcd820d555cc5e3b78d8390f9886ca0fdad9e0e6b5cd75cd21751fabe6d88bce
z04e055315824a694a6ec280b6ea6e49c830b93554fa13e5dd08de08967c40c2edd224b4dcdace4
z5e8703110dbc6aa521a4d911cce14ba7b8fbebf3df6c99ca4775b433a987c4bbeef7cdc160cd3f
z1e732a521810baf6489b6c01604c6b69f8305854d0616d902762d49e2707a5d8a4e9a6380097eb
ze59225fcb210d12405c494fddff51c5c5ae7a333e85aed0a2ebd919b87ffe6393ed32f262e75f2
z4d540964b4c24b13a6966c495341e7436ad0d36c1170cc47d0fdeaeb87480b11fa8c5fa86971a2
z77cb25bf02faca81c53383405122d26f581a52b67bcdf81fd34da39d1705c297356e7561f9de2e
z1902de7ecbb65f898603f85302d1e214f77324e03ce5ce0cd4f3cfcbb7aaf4ea9ef7becda5f6b3
zc8141195d01289f907ec5a3b4664df2a7984208a162d88d087538bf1800544c88eea6cd45a79b0
zf009d8360d75e16735a6c17e2ef415aef8b1a37edaed8aee96933b717395866e7e4b118552830f
zd5058a288b85c8572be43e944f59cb2ca0ff1ba1c71801e41982c52a1c526725cdc814c053d7a3
zb4aae5d9904341158e06a826fa7d5fc83d7869775d6f9cafac12cc4998bcb4fbf7230fa2a93f84
z8285fad1519dabf6892f20d97b47917e99e5b574f4edc4578a7109e03244f36e3dda0261f2a2d9
z57e08b9757063b9813410eee0eaa68e4bf96c80126576bc6fc634846f22e8f9acf1d25e0f1618b
zd8dfd40856bbc69122f7cd3ec947002dd273e49a3e1a9dcc47989bbc9b01e7d6d94de49b941b07
z45529bbc47b9abe712099170383b7306971b67761c4fb0b072f2db88a9f0133c442730c5ab6377
za28510c2b68a5ce6240c4b97f8960d0ac250024731b2086fda5010e5b12c1c507fc29557e4de25
z7e07a984ca9f5a8c5418d7f69da53aeb60e5bf0668cc978e75ab2f2a4a73105cf50ab59cf4bcbd
zd4137ec3710549348d5984b47e4be3220d281673516b7b982bf36d6abb623fdcef9666f51ebf11
z735de9d4602dabed3bb8f432aee0196e1712b1fe177b4d9cdc734dcc76c1e613445bf4d13cad7b
z3e6b911b43ac902d9271a96694eacc89d32eec2e3f3662f74e0eae85b8fc9a4d909de00fba7e55
z25b79421443d1d65e32b5c3f526c15bb21075d42570fe5b7e7e8ac094a650f8ba10e577663d114
ze3911eefa7eb0476c3f336e9a2dab63c5cc0063754119408a96de648a06dfc970a4ec89e7105e9
zdf50d8ec225d19bae44b51b3dd713a334c6d68551689f21877e7061a2611e61af28d4474200115
z1146493b3456531ec21048d4df5c57703c1db5ec946a09bf0bacf0aaeb9afd7cf9d8f8d9ff0062
zc51af5b635a86bca591ce843f07071ff13d8aa3f240d76c1b28ec90c74c24c09e416692b6f078f
z3400cce85a0664397a42b17c2ae0c41fcda6195c6b46dc743f37d39f9812bef2cdcad20b63d32b
z3282cfda04a15c3390844ee5731f6ee80fda46e7d86fec2679b44e2c6f17ea98b612a19d095201
zd44c84fb156faa1b2d1610618b5dfd35df0b7203438d25ed2c5b4e024c4929fee5df51d82ac614
zfd5b1a59cb66b53c68493bc08dc6a5f67f20f0f3cd96ab5e6a7e1c735bb5d842e161ce82157fff
z48345266e5241d9ebd0192fb1b1e024401961cbfe2d0d1581142e80a1bb3e9261e5c58f8107801
z780eb4fbf05f1ac7b5f8687fc39f9586731b1a35b7770d31eafee865b3d94c498d2cbd7a2e6af1
z42ee1b5beb69e7e30fd08b0af1219c87098474d549e1587391d30b78caeaddec8c6c4169d26275
z2e4b1070f323b609585f16cc0f58013eadf575527b24b958df35adeddfa9539e50f0e88ef46738
z895b0b36fa2e1e246ff4418d5113bb4f2d43b40eeaabf1bd4023f47d7770b468b8126dd4c8899f
z8182aed763218cf4cff13cd9c48ece7a00ae729865415a8e01a736e6d2ec49a11db62f2c699017
z76b2905b5daca09d6a41cbfefdfbd5fff93a135afc34f123fbb9e6647aff8fed45d2fe83793fcb
z798bc3dfae05ac8cbbdf31779d1899a600f6b1ccba43b5e23486cbb5cd159301019371a600da95
z1e82227b8c60e5213b25cc48344fb842b3bb11241c98545720de598a746e2ec74d9c837bdd73dd
z0d826e4fe5ff4ec3339fefe220ff11dd399f3ba5628231303b4c25e909f28b2ce9c35597eed2d6
z63ced8e0da63fd86740cbdf0469b4bac95da534d7427005b3398f4ad8e45de11bf2eaddc0e205d
z37edcdd583273d55681ead7301812f0617ac08e6a42f6d7e6dfe4b62253119c0c4b0a12deb0d12
z4c7d0ec1cdfa9fd2ff7651492ef40ef56052d7c1e8e7f52dbdc93d1d139926dc6b8308a1536ecd
zc4deec428510e6e418cf0ac24a54745b1419ab875f441bf11e13fdeee9a69d0f3a974bd77f15b2
z53b3f7ac2c24e260680d5f70f8bfa093a16c8262411ffd2ef95ab17b10665e0eb99895a03336ec
zbffbe950ba953437853ff6403abb4b039dd57398c4cd1e35270df86eec17ac62c6b5d512aba814
z149c2a09738222466b01c3360c81a53f1db19e65aaf76d7d651a30519ad0a474b82358341bb6ae
z22a50b1dd5a366b7803d697239e9afe4e9a05f68eb0a1cf99d4800886de80124ba71c34c92e095
z30022bcf9584381b511d929373db7f6002eb4e2db4d9029c04a4f53eeb8b3d4a486ed7d1a13c21
z1f14863562b7e48694906f8e33594f30cac71301616681310a0045b8bc9b49c31da08ae9d8b6a3
z150393fb2e5544c21ce44d91ad7be99fea79dfbfdfb303969eb76e9cb1f4601acb8fac9691ed51
z301514648a13e936fa46d9ff0a836f7e3d29d2ea8a0cbc553a492719c6bf5d6ef712461d401ebe
za210c4dcba26c237047a50645cd48ba48fe720172ca48801f58e3b7132cf31a6ac6fbbba83ccf1
za44c45bd12286ecab7908c52487a67075492c15236ccd32a352d003399b9476c9b68564084e005
zc1d1f0be74a352b679bf695e81115f4fa8c5df2c7160fddfcd3b18a6f8af009da6b2f80f66b246
zcac7fcc9ff96b8b23ca5caef1e33d6ba756efc52387d771ab3d52f1bdbf3b4ea4cd14dc448ccf0
z3e7e2dba1d51678f9aae484eb11db6b82b1b0216a11c9eecb3316e278816b98d0558e6d9f1b919
zd7595c51e41ba321c9ddd4a7627f93d6fe8c99f0dc6fa9b9c8366585b6961200c69c0d862ac3fa
zf3bfe4b9754860cd4dda80aeb1246a9a17e928407dfea18f626f09d23383b117efa2045e5ed2f1
zdd329e74ae8852651ef095eddbbe2c11690d8d7d62b58b964f511c67727b55365b3ab95993d601
z6797cd8b29e405f49403bb92064462326c5ecc80c98e800165482e08ef2b9c7b76998f8f947845
z7c6fdbbf64e63147237c69bdb32447c0ff157378b293324f57d12e085ae963cd76406d4cbeb41b
zeff601b38f18982c9c32a3a5eb83cf1e5a93a53202a50e6ef21e6fbe3010f5e67c2030949aab83
z2fd66edf165f721f76356e2e9f153685a3bae1a0388b58ae0236ab4645d50497426c0424a0fe2c
z37ba461d99abb5b8140b88e68a2fdf8a08dac535a7391bf1e657978914461b636a36c9a50ed0fa
z852b1f9574e1c3f032fd1d0ff06561fe3c960abc05b61bd42b49c5425e952033fb2eb4039c0140
za39eba57a5938160113057ccc4448dea4458413cca55093418757ebea40d665fb88ef71c635b76
zb586c14ef83c635f77706c616f890ac3a0780542af2c6683ddea406165b93833c9d0a4c58f3d81
z02ce525e03e4a16df3928cd10872851e97eba8263b8e2ab493f26841c9771877e6df70b4479271
z2acd3e918e3b8a20290a49c805966851cd97407f84d443d9d2f8262125a8e082a4bd9a946d4228
z70b4f0be525cc6d7bf88d1a808c47fda39c9d81774c2f9d713666decf066323081652bbdedf86e
z45667949706ab4cc266fa443d6d074a785e2bc4b28f3f66ef97365e2fa935807a43a42ad683f59
z07985fa0ee0954111cac1315304d76bc1f53158492e9bedc56ab1f33b96ba2442961b01d271591
z2f6c19d549faf652f491713d3f712e4b4717aa440abdabcf01460aefc6a0578253be8653e9bb49
ze205fa4401ae1cca33c98f804ac3b1a1b4b79b95ed5b25991a35c43b238ae9f954d3b6e0f4b71f
zbfb6156322bc7cb5b26ed75bd1fccdfdaa1c5692c3456012db275c706bc91ccb24813a1508587b
z336a90fe6046bbcd79eff13a9a87814ace4f1c5f025247066198c344e85a0477002d81dee8b91b
z29d50d3dd80899e3969a0d00d5797bc560cab2a943c6a4b2b620761ab303d887d6d08f38dcb686
zd5194cebfc97975901aed50140f4e49ab8d8c8dac666650c3ccdd238e5a0341fe5cc218b87ff59
z89cfeaa7ed1a29ee1b6141d36dc8444ccf2a9205761348b6646c651472ecf8f0e927085790e132
zc0b373dfe2adf1a3e483b17ed50052461a0364b239f4272d6f485de1f4003cd72213bb18b9cc78
zed8f0a465592cbfbe645cc9ec2fd2cd078429b53f4c2b2705596140e3d149991e8882507892c70
z39c1075e28fb59c9e4ad9174238b956be98df8784bdc3bc5e92d9c67f2a85b371ea5acf74dbfb3
zde5398d281456d70f477c8fd726e47167f628eabb2b213322332f620e66f902b97988cec145958
z410a4f17f1a13a8d4192e260d3bc300025a7bfae158aa8092404792873bb7eaa2eb55dc43227ee
z046ac3b27aff4233be2fa2f48d1126e037948f656c9bc8325a230892b4c9e91d5b9f299ab17d93
zf02ce73c70a50e1f744034315f2961830ef2d58a1265b8763e6911a50386514edd1d3234df2153
ze4778ae9e0fa3651b706e0a7f61973214d34d545d7da14ceaa90536683243def53e60a3cba9130
z442bb6b6a0aa798f6a50895efbc0eeeedce5c5a27b2eb4ca306e69b80a97801ded89c43939ca01
z710f9bafc65c1fa11f4abaa886b024b45a4e624959fdbdafa268b8914d78c4eaf25897dee1121f
zd7ae06b1798f65ef704e950ed9ecc522a8e7a95d9d22fd725bb35757a2eb2c2a8a60b9b0342ee0
ze39910fe4cec0f2c5c0f9d004a10ce902f7955311e2acd408b7def55384687660030422305550a
za30e5e8f6bc105da2a50380b11d9a5658a8a20290ecd62a079435042f437e6bf1f59c776f2279b
z5a5da1fa71fa153382b8a0c484b48f30638a1e5ec431e039e2c9262980c40f11a61c468e83dd4a
z421238769ff413b3a0ca62959cd492ac15a265386285977cd788dd4a7f791027117d8c69b0446f
z7a3b4e4c6495b3b515f6e0c003fd3db39f938f94dd4b63febba60a34ab6bf1c3a1f7799499f11f
z741944523ed7672027dabd19268658b70ed3ef159f129160051b990f27273d93b972f4e19213f1
zeaae16e527012a0a8142d4e22e89d2d40a8eac57babe04a1b3945239e690f46a968298fc867dfa
z267f3342aa7da987be1035186235a4ab9626a9f82df6127729744e7cd28f88f1bc9176f1dea8ad
z2f4b4cb5fac586b4191da4c5eadcb7a43c8715acad21c6dbc644c6346ef30454ba6873a77b01bc
zbc4852c830cb83dc4bf9876521365a62bbe2b8e03e39ee016d4e4f8c311a3439dcee73e6915e45
za62fa826a65cc0cfbc32ab4854c15f9e3aea792025eb130eb433293573add1734a9278f3db9532
z97c62ff87f23c70298b1a13506054344c51b677543b442e796a5263dbe9fdeab46f6d757b9cb08
z98121db9b464eeb1f5c9d1c3eea2bf61f9301f5a39a331d96f0d433b063fe5e8020fbd7c4138ab
zbe7c0d0c530cda9425ba66962049488e1a1c9e14b663adf034959fe44c36e2ab4c5e7ef8285922
z7d331ba75657c0099bbf81f01a77ed48843988f3a058859ddd21ba5dd86d033b62c6f1adff5585
zb9f230ec96a0a527243e3603e1378ea41759f44ab3fbe05928502f7eb311076e986c3e5360958b
z170ad9c0f0f05440a3b3e067e3cfb674af5d97e21faaf3b0288b11fc6c10ed52579288e4a5776d
z83912eb5e9ded795ccee9677244917084bb0c2adb3ecc6e90f44ad0331c97e0d4e3ff173808685
z8def85ca722845693e038b1956524cce06ec4128a13ba888591bcf512954dbc0d0bf6d78cd8212
za4ec0ea7b3f32bd9b886ca2ec1550a5a16adc3fb952f446334312a8b77fef5bb4f5f70238d5112
z53f39e29f8724268cd3fb9f958ccb7efed69b4a2915658231db56c06545bfc0713d646fccaf897
z1a361895722bda42c57261185da2cbcdfb378f9d81f446510ee669c3645ccd793e43329bf6a3c4
z5d32c25d86bc1df9f09341d683bda5ef27714ee5d8aa926a26970d2cf3e4d7fee3f84fad444136
z6ee500d73a5ed24dc8d484c9a7b10316c4bd1371e336a3aa32ee0ebd58a23c992040ebe6925553
z305866e1ae856dc3dc0ef7122c55190bbdab9efa6ff1ac1cc82100be2dfdfaec7a8ebc82a9cbe2
zb6fa1cf862d2d3140378b3a26cbefdc4daf8cff9ef0df7d9f0510df4f4cdefa99783120a1742bc
z89d635a39c1cdf0967a539e0ea8df8ff1f8c88a6761fd61498f4e8860090bba3f9a5193e27de1d
zd7081698aca74cbb852a6e90274898086e0516b9a0fd8b6fd4b7c8efeb3ca7e9680b98da58bf3f
z7dd6ec3a211348465d5409228666a651aa5f359f6a87d702e08908b6e2b4c1f5ab455d8f4fd423
zd1d87dd1d92c1338508431da28934177f19a10b395ada90fbaa057142527d16f8a79928deacc5f
z9d780f34f93d69ae50ca7be9d4b7adca09b313cb8edaaa4a137643f2998c267e74c30382379fe4
z67338f1f7b00d0d221a534b791db6b32bdacd9eee48ae694012dfa362371a69ace73cf0dc61e83
z9ee98eb138e0c677c2f54aeea4809d7c943b38c0842e062ec46696f26c4bffc622a7fff33cff82
z879aa19b13cf04425e4b7f2ddca8df1332c8abaa030ffb1c30e75d680c2bda3b3aed357030baf8
z4d330adaa2b03d70cc2119f38fe8cb9484f2d26f9bc4d2792e902832f96bcbb58a6cc955a958bd
z1b5c67cfce9b9535ea64359ef21cf28ecbfd58d190f42cfd28f1c983f228f69f0aa2dd69309962
z5a4d0c0a378181a4073cc069bfebbfc677b55c1a6940e0e519953744c259e8b98abed04b6599b1
z333de9bb87fe78d869c497dfa6d2932acfaee884e80787e2818b441db7909477036776f3940af6
z3b9e9b61cad8c6d66eeadb80bb955ce4d4e5592049faca9b31c2d610ece777584610834fbd925b
zf21a023e5355741bf1fb72ad35d9c33bcc85dd44ee29c9f22e3fe5863ac3f392f4f71a422c9c42
z9f425208da8d2cb795efda837857e7f829477073f85a2d845bf07ab096d563ea51dc6fa474d1aa
z90625e8d8295ea00e303608fdd775c04b1f324984d72c9238eaace7c9e2540fabca777cfb70c27
z8934713b8282c14442b56fdcaf36d69ddaf7a0727192cbd448e9d5b6a97c6e160e7cbce0ace225
zb89ec7198ff1556d3a06f02f9504b01d8c479be43ca9bbaf0f78053f52931a64f8360f55658b3a
zd708ef9b291cd85e7414a6a20dff7d86f8d55c0ca2e9bb3ee7d88f90880cb1e0a5d49cb0301db8
z05f4886885954e3e10f5ccb82328040e7392f81ab9cfa3304157f9d36355a8b71d04e9b6dc263c
z1ff6ded6667327c5f261cb6c53ac78f8379f73bea9bd6165b7f1992fb0b4fdba590f33d7cf8e40
z006fbaa0fdc59397b1b8548e14c4bf8627d07772058999fe6e775a72d1e9a6d41b792af4d43e86
zd4a79f2a4d7615c89f90b5a5888714d7989e794bbfe4dac71406cc3e0695a49eedc573e87f1918
zae52c3f6f4c410316289b69770e20be24e4e424ea1db43db95aa59ee8b5bdc1324de198fd91603
z75362e2668163d07d649787ceb8acc761fd0f7ad4f126eb3ad4e826626c3f4232022218da2a0df
z63923294cf9499d57a64249d1c52a9a03c96fdd9f940bbcf4dddabf088dd4f94033d299596e652
z1998fc64cc43b9cc942281baa15d56290bcf6fffca9122b59b01b2ad73d045f7410165329de042
zd9b2676b38f833b285f2b85d6d1c833f1003ff9b4b639bb8cd6d32e7a014793fd3d674044972e4
z40a30fc77c9e37cc01baa66ec1b0b9d4b5095e8052916ac89354b67074bd57c78665cc03f0e2eb
z069918f966ea68e37131c80e424137f0f281d4f4c60a6d1f2b18b758739d0cd15bc0b82f43186c
ze398eaf1a3a28348150b912c61d843fec18a65da07ac7998ae163b88992dfc01f1f318b18acda0
z8c9f416e1061aeb71feb320b8bff46b88331319a77404b1493efc872eacf66c4ebc826c565c0a7
zf99c846569a3a6784471f23566aca22940fe0768816c6326702cd7f0837d9b29f0db8bb4588675
z9a7117778eb25825ac4335473697a2cf284bae41ea8345f4f1a7ae8c09610d4ce2a636e37a3f78
z87a204cd7b00f56d5001642e217cc0b8f7d213d8219219d16567262ade480dca16f2d8421216aa
zdf308bf6d3c9e5d1eff04179888b3ef0c77c96aff160883db19e641331fba013c054df9ed4efc7
z77b6598e0b535898fce1e2a55cad7705168e43694b18f98a318385e53ebc36a93e81c89ec8cf49
za1a33dba9ca8e1d4262de44800b6aa72e57aac2180e3501272704b0214672b91e90746428695e9
zdd14d184d3d9e6c0fd7dcfd44c3f244b3ba54210f0e9d0655e10db39f1d210cbbab5c80956e6ae
z3db129cacf8c97cef30c99501880092ffd62cd8d015e0475042f100165591c9a4f2789ae6542c2
zdc5cc3f782b1eb9680383fbcf2901810148f8586c4629b3ca203ddce34ef49db37aadb91b2e0f1
zd25b74819bcde8bc6bd48577375348a8d34e3e6c8329cd7396748a9959f45ed3d2303870e5a685
z1f5d8c23e1e119397d0929fe2eb6c6e73c901ee417ca791ee2eb735ab8e79c61c45555a699124d
z11bdaf53c59433fd8595116b15bb93fc02bf2e48321d45818b9c73aa3c1ca81890a79a1427e455
z04a2fe7f8a59390bac0c42f1f3c7b1ca9df0081dcb115bc8a1b67c135ede080e8d010b2945adf6
z55fbad9ade7a6f3576626e0700940aab1817113fb1c88e03505fd37ddef2813c2720785ff8415a
z23553a065f625e3f234b535bcaa7c932f794f143b8e0207472270ee9987d92383c2873180c0a17
z9fa4a3ec20497c4daa4ce275612a88035948ae69465fbb9d24b765016b0f22dd79d3a22d0f0485
z98aaed2eeef8d8de621dc5ae303aca0b0fbb8bdeeb32194da247d04a81e5c0a89cf5604f05c577
z9d101505837703ae67691ff3f2fec935b4acbe8f282e04891daa2e74ad5d5f485b8d503568713d
z22103295b8b07b57d4d7896de8e62fe37909b68d9ef3f1cb147697014a09875d866958cc6e6d52
z6252222934825c1e89d136fbc72aeca8823104b3d14396f3f13300401af0cb4d7290ea799000e2
zefa39c865249be74b1a309a380952e995f24884392daa8297311b4d9ca37ae38bb2d0093ddfcf9
z67667ed422040b4542955390993b38e2a34c9d6192ed7e147f745ec04561862b5380780e9b1a03
zb7bd1b97149fd44b4326e46d36aac7685c80c9b25cc511badd04ee1e765c1df0894a6a2651ffd3
zf32fc35b5e5c3b37dd1073758cac2a80ef3378fba2cc843a385dcaba158327f2c4c527cd4db410
zd04b96f05f0364c2cf63c575b6d8143b6e06ba545a5b2b0bce1fdf2b089b36e25afaced6903240
zcb83e0e55457b8266dfe15d263c58ae801f1132f4459beb5f914e1bc740c6a106800a4aa84467d
za3117314088096ea5d375a53796d13672abea359c3947536189aa87a0ebf15162cfaf6d1fd30f0
ze9bebc168decf571ca5ab4b66c5ae8307539dd9212ff43fdd056dd6a33af84d44796a3a67718e3
z6df306a3779b1ca4bf7ece573b0edd74804f230c47b7e76cde94a74ae289e1b616c6aae3a43336
z62d0de01460cddc258d2c733c37f390c1492e1cb9dd305a82632cb0bcb0ff0fc9261f53eb268d0
z8729602a8cdf565a7af673db9e86bb3b5609e44c9f1a42c8065817d66a3b8a3425644cd860e37f
z32d64b01ef481a62c03c6b369aec73c3e63569e09937eca2613805ab2a090ea53114b2d40f8644
z6a360d55d795a97daecd4cc1469d1aaaf4dfb63ae4cd50e55cd3e2144483e1af06025454ecb653
zea6502e3307a2e76eb607da6940b9913b3e162588ac72a65188bafa43a0cab4659f5c37fb2b5ee
z0950fe7e6a789515cd4c9f6dc3f48faa7321d35597edf0e437982aa6fe219486419b7cc01ecd79
za096c3d9d19b52c1287ec2d42e444b455b981b3ba67a5133868a8fa68f116cac9d4bfacbf3e4f0
z1336cbb0edc929a939c4112de5fb3beb69f78a6c1b195d0a1e2fbd6fc64c6f5bdafe93566fbc93
z5b291c6071ebf41d82cb596cb2b4e277cf7fb3c9d774a5d28a6e5b0cced5cd4540fbe81eb80c76
z6dccd085e7a077c49f39f42da37ccdfd586a6fb1a658f3acec0907bcd2ab9b625c949cec6f8145
z997680e9b73d7a0c99826adb3140befacffe688ab7a0ebcc8eecec977cb7a72ba9b6d343a4fe22
z27d15e962280f5cc8653af7728b1009ea94cc1702aa00ab4dd3e2e30d05eeebe1770a6790e5030
z54698426a8923183e160e46a713c28b612c3bde47b7c763455a2e0734fcd1638cfeb32b680f697
z738b06447298774b0dd4c5bfa4081580d6ad91aef9b4f9a43533e0f4ace1a4e66e55a624ef739f
zbe4e0dfd2828f8c600c907e5e52fb73011d6a7209fb9afed1add67f3bffb70470951b8905682bf
z6b995419cef602c2da48855a3ef2b438ebf89cb9c5cc388170e6be1c2f1b52c1ac64ab1ad52487
z14d87334464f9077de679fc0ec38c2afe3e08a8e3e4f428d6451d1bc3bccc46e250b62296608ad
z0617634740d441eeee4bd92c33acfb96bb5eca873dc369ca95415585d92095162b902471cbc1a4
z2f4567cf10718d8d5cf52a1a2d418bdce17ed8c22ba7fe9add14a270edf7f062c6f39ac80a9664
zeb3a77286871df6968e8f9500ae683a8f6750a0881905ebddb252b83440eb7b9ab6364c4288eb8
zf031dcb5e08906774a121d7f3af57df697354db1dbe7b5f518123cd536eddf4bccb3b945896918
zcbf148c25bc100f54769e1f319d9be5913ff870188bc5cb067a61de5e50f62d7dd67955319a529
z504a62382a2dc1966b16da88ea2431a74242d1b0203f557c0d307d88d71f1711e0d565a4b83b29
zfe476ff7f125f340b64ec99c196e53c9caf6f3d6490d35a7e90227d6eb664002d8bcb2205a03dc
zf4998a8cdc8a999839e77aaa204a1108ecbad2a397856259a7a648e4f38a0e5835f66b2f97f517
z66590ea1933bb740e88d3045b6fc4c1d971728c24c51b64dde2f3f6fe009f1164850e073a5c98f
zcd243538d66a01cf6514e138461fe978622e328e181ba7b7f7234a656015d3c82f4c1b590b521f
zbea2fe67a6a0d77f6faaf894c19a0b27b37cf61c82e0b7e5b38c8a50bbcabe56b7382e7c7a7b48
z35d62a552e078d5c1d256ce3431709fb657944993504cad595a2d50e8a9a7444082512ae53ba7d
zdddc6faec95c2981ac65623f119677e6ed1c2dfa98deee137653e0f63d0f17e47b9091279f52a2
z021a407803cccf63fcf8bd6af6bc905f2e7995ec5a2ac9b7d062d85b8edc9ea694dfad6e7555de
z585f2075d48104e49dc9a4af02255558473ca143224cb6a4618d5af3bcc9fd5a28e91e27e0928a
z038d99e2592edbc8c5637bef88532043eac3f4e7d31d6d57a70a7822d6ed0d78d79a945a3b0796
ze1357e3fd2a90937464054114eca13caf5b919bfd6432c93351b0113484b3ec75549322c9263dd
z4472eaaa42f3fefd7ce9b731916df8c5b0a5cf8805c0f1600070fad38790c185fbc0736f256a66
zb8c32f1e55aaaf548cb13748a21b71584159201837a131c6a113c45e836052f25f5e829b923515
zf27f66deb0eff48f3bc153170d50f5762d6d41e0c2a9c1193ff359a92516680f5dd23d0b4ac4ec
z6b50f1e3e0d52c204b56b0bc4f95058da6e03c8be61e3e2b532cf68f88b214034190dc5acae153
z3496facc9cb3b81037fac21737d43c1670740f7ae1d64dfc20455c7b30a96c2a8b183fb73284f6
za083756d98410e30eba0119682c61cd4cdcc1fd55f3e6b94b110e70c1adafea315b51a07f470a8
za21ef24441cff83742c5bf933866df49da41766c7685ac9964ba7cf3ebdd61bddd86293649b6f6
z245888e53382dd14f74ee8ce4d5dc31c346c4a5380917fe816d40669c6eefeadf3e7de5f36de89
z27e07938be3e5b6fe90baa86633d0bb762cec92e934542025b42c5f62f20fb8c98acda3df6c3d2
zdc97387c5b725c7440cc9403851b6f0d3c5851069cba93d3697c36b4cb59414371156efbfce52c
zefd9eaf8b7ef861d2b5f12748330a6fe39e24f3699397812ad23e9b8172a1aa017cf68291bb44c
zed5ddcc4735059e62a38da23f11a83fe83fde0b565056fda328a27e280bc525344d8c2f6db857b
z0c81d3d9240b3b0c4cc80e6dc4febfe0455b27858a0ddc5ef4c9f9f4cf379cd628e7c7709b25a1
zb7f09a2d32b9ce4d05537b504282844f1135c5a5a66915ae4e5d29757eeeb132eeb54145f60a74
z417b817b3b591e7bf74c6bb5691dcb2b0914b07f5f2b51c5bf0f720701f06e5023dff6e4af6b52
zd48c7c90227fd93b98487dd84b473fa6218c4e476d3d6eca5271a2861a2cc5afde64803f93ec79
zd4f0b290bb4824376b75f373b001b40c6a53ec567610248454e22eb4b6e0745d0b2fbdec142cce
zd89db350b2ea810944dc37a927fb9995a0fe30576a210dab5c7b8a24d82e3b7584e4834dab0419
z268cb8302a26bb02a96d310c5c2d88ca4a0ce35ca42b0f4236e501e663e129b63a1ccf300c112b
z3996a12cffc3c77726d8845f82127c65cfa73e9fccbcfb42885357b2bfb131a3489b391fe9cd38
z5836e3a47abab9f3a3940bdcfc48ba255c6e39a9afc5364ec379872359c156b7f4085d5dac521a
z9eb20ba018ac02392349b1b51db7eb17be5c2156d1d51294e1e6f19ff831e86f6e42d76396c877
z4fd76e0ac26a657099d4f05b2682113a02f84489c9b2ba7918aad2f5662d4cfbe04ff681b82565
z8e45a833d3355fde57138d34f76775475c48253468c5ee0be01d718cd490967431de0292eee9b0
z84342e381b4587ba62c548005ca8fab85b0d96157e995e32f81e7ac57a6d7ff8f7ec3c113d05ea
z4df67a239d93815b3c2ad672ec56eaae148d281efb502b231c06158aeb01f656d41125f4d0e052
z866ce8fa7723f542d7a04c0299fd43a1e9ff9efe361e556782af882d413cd90797a4813bba6b62
zd771532e61c15961bbecc1db68ced058fe5aed8d5106e7f5f2c54170938864ec12ccfa869b8190
z88d952a4030cd4b5b8356ba4695f2e75504fc68e0bfdf61f2df79ee447f7b6e53f61493557a5da
zdac4b479cc19ebdf9c370a1abf58e2ed2cf427901c06a4c30d31c92c373fa49461ce41ca9a2cf2
z605a2806708a2b979d99c3efef0c7a502eeec7b06de7445b505247b38ef5c4baa9499c297031ff
z74b4f9f5e99abcd581cb176252b2b1d7bcfce10ac2f23a8c3d8294bc4e49b64ad28ac4dcc1feff
z8a825d4c06a022971552089ac04c1ec6a41de42d26cbfa234e2f328162f460d384c98aae2bdd2d
z530aec64670297e3fa8334bb4d70c6a5da7264a594e4b54e8854ba36a5a30b0aaae19b81c766b9
z5e47e82dddbf088405e4db96ad24cd9afb8490ef74e5de7e8125e3781cb88e5128934d3c6c7aca
z9d25fc1bf18b4b1c759e3ded91e1a0411d03d06e8a8244dc8aa6677ce726325dc8eb1cae55e659
za4bd503c8a6e8a5dd61d6249ede06459f630235bf039a963aa6dc917fc4a77202bfa3f0b834105
z914fa7c5e2d9f4620fc18e672d809f92f385881528305ddd4a54d6f8ffdabbfb74b62b0cf87bdd
zb70bf8fda96c8ea7cb839fca82077adc548999a3273b2cc60f85ef5e29912c23d6d3cc94dc8c72
z9cd194c1690f114093462d0482e1f07f221f1331661fe7cfb30f9c272ca868084cc69013476396
z281296b9736f1646a94fd5c0753a976280941ab311e1796936fd20dd82645829b1dd845b245bdf
zbb791643863b22d2be96f867418fec5f8efaa5599e8d9d0f7cfd485f4a6ce4a97769ebcb77fbbf
zb4f40276eff375a44cf06e24ea6225df2dd0e7c5fc15ca2f2e28cacd2aa12472f7b30ac5553d0e
z59fae6e7ba1469eb96fc5927cb52f1983a71b29c8c5b5faa05e2a6d7457f54662b8d35bef661d7
z5cb65cffb9e264dd96875a13228e55a72d2615f7cdaf469833bd1d1b74c39167062202c099dc55
z58c6acb2077b4c96547d644f4511118f9900f4b3d2e9626b53ec47c869c7fcfac76d46e950c0ee
z73195ac01297fbe879729f43088015cb4d68f11fe1951f8fb462e80fbb9940d46ec17a667870de
zea25b4cf6782667d63890bd0037d843d17e075a5d62133b18c787e786fa52a013dcdaa0a3dafb6
z1b8e46530f2c91586a228a6dc2b66230f5c9fe11b379ef72b18e435b69d43eafaff9533668af88
z414f5c2368f2703c82999167be6ba44fa1c77d07e10cf3c328560e563e29d187b5cd108f46cb94
zdee904e41571e8bb4d0428c897ede072614f4084da06868d7bb05ee40736615e124971fa42cc0b
zca80e8fab674cda20bf1a54a40ff017ecfb366b52ea3027c3056a4181e09d22c22ca64cd759a51
z058af8346186cd6de3f0c1e0fd75f30fb7532a545d4e0ab7b8837ad71240abc9a6c6d18b259551
zd41750dd54cb38ab815b023ee422700b4664582a2b338ea455c0d1e098e2825b85e9aed3de46be
z98bfa9298b3d2d85b92ecc30cbe8e239db1496f7c6754d256c9a4e6c8847292070c23aa3bd2834
zb4ffd6b7420635b961c4145e9b932229a2cd932026bc8af384808dbb48974751a3493329863a4a
zc739e90a4a59ddf035ee56fd8011e6a18e89614db28b81c663e7e526abc071b19ba345cfb6d30c
zd24b44def0c0f79056f923a1bad0edd357287ff2d3fef31532bc8080b6233ffba3efdcf6add8ce
zfb8f6374f2fcd06f781127f23a9043291d0863c56699f82c56025c157d8fcb3b60f5cb219586a2
z6a5afd8f0f1cecb7b731f26a8f504095ce1e98324fcfbf809b1a02739499adb739fb063f5e534c
z915e24a37f8e029bda240d27b19e4f78f31e3ccc5febc51ba20b5cc2206838a713ec27353d6330
z8264be65f0f035833141b6c77a6c13b7b12b6b683be40dea157eebf393148c9477d05f1d3606c8
z1035440837d08d2e0b005446f0a44f7ca11193410fe84f0b2699f772f8732f88cdfc1e77ad92f3
zb7ef0aed9e1e8d7f964962542b03c2373ad2784f8e98cf3aff1b352926fdc1aeac85d8245800d2
z79ea273e239cec464ccd039694b3d195e64b39ccb2a9c21aeb487f4f5653c90532c104033889c7
z60052c2e7f3d4910e9736b68b2d3ac3f29986b24867edefb3b61cfcaad19a6dd1cbb87152a4eb0
zd53b943b20baef7b6bc46c3699a8628a1d5937b681c9dd13c3ebe3b17e768f6e1f222ae2609f2a
z37301aad6fd32320d6b22a7be55a64fdcad8fb5b0639bbf87b1ac67e64ba13c45a9b8866760c59
z8609ce31725e8edcd496f8349c36c9ec72ccc5f15e4e4bdd9017d0ca225eec09e583c4343c3328
zcebf4a1406f957a1806cdbc7f01263b505c09f9cac5a740a2e13a7a9d77ae8c528c3298c72bf45
z4ee4d1bf5745afcccc9961dd756da73a87954786edae52f1d6bef48263b9d064957f1f3f3df507
z54f25feb03b65c71ffb92647cd40ed00bed5d52a21d1784f35d266d049b726421432f69e4c89e5
z576c6b02777444bc8b860ba261f735e9e04cb35eb4b70f9e14f91e3626a289dcfea2c2cdf5d53c
ze5ab62eda2661afa56838b8609c325bc4e6279b3cd974e62f93dfda15b73fb316d17fc0aca86ab
z80c7dd0fc2e58c0f57fb239eda43d4f8217b4a93e429a3b044576029714ffab87b44bc13824fca
z34cd47e608005469769295c98a11337f2bcaa47c54feacd53a4ad9047eaea8ff205744206b2c20
zeb3e4ad3d4d47b233518d1c1fc7da5adae6f8a617d573ab429ef23aebb27563c69528d7284a593
za49dc629d57e6510158aae6f66871f89d471304bcfadef2a84e0bed7a6aec098bfd53f607e608b
z38a1ccb2c0ff8baac2377ed4552cd92865b92118a165141839f2788e7c025eee152c1618caf1b7
z9b35fa9234e4c78262519ac441593ecd1529e9b36ff0d71597dc0191dc8ff19c4effae1f158096
zcf790f047561ea4efa858cf381e273f69a224685e679c465b83a09b6ce50ee4322c4cfeb9cfba8
zb41ac2467e8a8ac57bb46b3f3d2940fe737f33704a95a76abe51cd250a489e7e0c82d80a482ace
z4ea847d73cefe39f31482c17389b53ec29d73f12f6795aa2f6ff55bd959df0d6c3d23545466989
zbd2bc0994ccedaf57337ec22c21c348a6e1a8144ab3039295d88224b9f979f2bad5b8db3bd7ae7
z0d109c8d7d3657c58db5cf55d90afb85ce2eb83fd87899b25110256ce23d776d849b0aca26eaa4
zdc552dc3336712632066ca98db7462738a05f9ae2de44672d81cd8cd200f515402374548ea91e5
z3980732d4fac4be0d172e3a270f575ada5a492231e5cd2d2d85a849ad518f88b0f436fa742868b
ze8fc81f48ad20fed5a0f13ff634ee44bba98bf69f62f91f336091a9987de253cb593928e72727f
z661bc9029dd41db424110153dd6e26daf8be522f209daddf71fd234de3a3283a7defe8c560ef86
z87ad5381414c76acd2ecd547cbec7e8cee0ece3bce72a6ae045a64c5da70204e985bf7a80f29cc
z3382d9f6d20317fdc85789b4564213bba7a8e79dbd5db7a27f9884df0991d74ea938acf04b86d4
z60696cc2789b66c4e60937d6c8907c2d24bc031762f7502900c5e527f6b785741a245d6a681760
z3db65cb970a7ec6e176f1c572904e7de369f34d79aac5a965a9b96b10aea5ea19e56572cb2f999
z9aef32f377861fcd0cf10a1d66e0b95b5c846a3100976ab39ac75a42352b1b4275da5330f95c98
z0884e9829ba6ad7ca8818ec2d6e7b59ced3d2087fe5949ba6ec4b30a1f8ece22c45f729a832078
ze9bd6227cdf1146f2052293376197494c7c73011c67c63dcb7b2bc09ad857e3592ca6569cce9b6
z46d034199681a19a2117dc4c895f28692fbe7d8326242ea63b94d57fe590d84d7d3a297e33b740
z53f9b49aa75ad428f0812d89d4631f328629a91d9bba634783f33687c3d41f64722a6210a86ec9
zffee3f02b8f88342bf311a957e52ba06e6466f2f880b53c7c81a04ad4919f26b95e64b32188c84
zc63092c5d2ba6fea67d6422f26cd486e8be5d865bf5194a13b5c19bd7799dc7a33ecb5dcc1fcab
z985d493c5281d0afe5fa3828170ca7a42f9f883f1b9f5c7710257f60e477c318889dbb7f14aee7
za1c688beb60ea891d0f40f51cfa77aec66f514345740bfdec38b7013ff39a465c0835aa0499037
za6739fbcead49d8603941131befdfd58ab0e3f28f00b480431a3abc50c1007f97e8a1ce2463d08
zec1e765cc46a126665e31feaf4b8edeb116786e7939b11397af5e392aef501bea1219d1acc4f96
z935ac705884569e0726196fd83c236258bd0813cde7f7857849238ec9812ce908b224cbe6ddbf0
zb54deb961229015c33b82c50afebda7cf33a4739d890813105e3973d9ffaa20dd945374ca8eb7a
zc4641e34468c4e71ae7ccbb318eecd75468084f387a18dfa1c91598b4bcee9b90e1c9411ef2034
zd9691e98fd3864b253a610a55271063f186b8c5aa51c7806e3aec85edda1f9d462c661e34cfe1d
z3dfa427f8b44da2057eefb148b81ca55483b20e7eceef4b49da9f820fd453e6ab9b74a0ba45365
z73436dae60da136cf43031c839746b35d7a49e71f04c332c1ee705b3ab200c670899c9e2dcfb72
ze72fbab0cb898b250b5944d80a367939fb2dad8be03fbbff24b39630b764bff9ef65a36d2621a7
z75c4155d271de42141d2f4c537ff628d4acbd88078fd94e89b45e2b3210310cc48a067698635fc
zd72da5df2a10a277487de6d515222b17cc6387504f19216dc8b54f8d34390ee9c240e0b6a88c76
z17dd72a7c40b8d1ff2e531f4736cd3c1fdabe76567d425b21793618e9da6d371fc8dba08939b88
z3d31bca9f97a2ff2d8bc72a6056834e0c27674f3e1bebd0083c29af4c5bdc02f200e2e94783f86
ze31cb0a5ac4f2c116022c8fb86d7c7388f0ddc917c537afc635ea3b3e1ccd1c7725bbb8c14db62
z4514849c45dc6b9f885b4ae0c92179fc6d8d84b14102feb0295fafa6e4b7ebe5834d0191bb20d4
z70607bab37807e7174666fd12387900e3af03619181092c3749d0779ad77c6af4839e4b7f80f8f
z6a1108a6f4ef829b2c68a15fedbd5b4bcced5bb2e8217ddb40ab57d9cb14e73480dcc4e9d92548
zbb6ad351b30f3add36a5bb89b93f1471be7a70fae2303d75ee8258fa4afd6a792ea8da2306bf1d
z0d7f436ee42b015dfbc9506cad0c7bc20f5e566d385595593698791ed673eac7f04a363b56873c
z0e2a543f02aab041431563a1274bd465a19a168fd0b28f0430ad36942bf69fe73908d10a933528
z32d734877b3a2cef2dc8051f4f58d57f553325c5e75431af3fdb56830a218abbf769f130687a0c
z61e38fd27f3e67fdbf10666ae2daa904830b9da0cbb56008339795e24389414f82ceaab9f9d689
z0a91c5316819c137c8263dcdb171881610b79fc988a6c9ee0a191132d02d3bbf287457cea8374b
z1ff7c45f5d8807151e34f47b375ba282810ab6d636e23cacbdf199be178ae3e58df65b2f449b4d
zf6bf4d21cce76159326409d4e75b6eaaa3ca9ef42937ba19ad0ddcef27a05646a492403d03df52
zf2b9464e73932175f97e41f2aad7288a0783c8c6b750c932cfc93901109024dd2e6e36a63c3fa8
zb1caef7ea0a3f6e7d9699fb7b756158f6fd211d8390ae97e60cbf30528eaf9cffe3132a5ad547a
z3397616bd7442a2594fd183957ef2d71febae55c26653e83e9c3f88cf0a917289654cd73ddf035
zcbc7c1de4690f72edebc25bc2c859ceeadf8f71cc52df3241bebf9f9554166e5f9d593229ec74f
za11d6dd4562251fd15f433c2892ebf52311fcc7ada209435121556f23614bc496416de7d44d5e7
z1be557caffe903372d0accd6544f2a6048b30034f6f3cf5934ff335de4dbab2a29f39690cc71ef
z8634d0d412fbf4ee7b3c2e729f790ff82d8ca38479f0c8a4b96806c2febca7a09a1f172c59ce90
zaa7de7033f6052d6fe4237a0881b7a85b76a6cc43599edeefcca4651a48743f43dfb25a5ecaf7a
z3fc7ec765ad0406a82ef7552757a6a7df464e03315ddc91b99b7f2d6ee5a9349993de728db7c4d
z517879e06b48e791ca1518c16ea88c9b6c914515fe2b4779d6bb2098339379dfa135b79bd5c97a
zf78256d81c2533bbf87cfe2120efc3bf367906d0ed80c85b4312b7f2f57f01553366e0db0dcc87
z7dbf68ec8f110833ef50dce963c286281bc79b53834e835d02b9ab526a07d8836b372bb26b14c3
z75488bbf3992735d29a84c33a4eb1251bc202575a8a7dcc09bd6a3138364dbcf4f846905ae7320
z9ad866909e94f8c89b843b206e05dfe78453ef42e4308094c862b2637caa2b31df6f0e817c24d7
z84e53aa8642f82336858e99df54eb1ba227c4cadfde0a28d0bfc7289078e29f5d061b83fdfefb3
z6a3277f63a3586bd1c0737b7076f6f191b787e8dbd3812bb43c674d51ff6f05181768b679c8ad7
z1e8d4545e27adae80ff54203a4de694912994dad0212f3138e42f3643634f6972ddfd37489b8fe
z08571d39e13225364aa137ae44cfafcf67de2693e6d0b4e311ca2f4007ca50b2e864bded9c39f4
z849efdbe03676da6a945c3f27a488ac790d0a78de57ab96537cc258c89fe1681edfd0cdbe845c9
zcc515db5af0b41759dddef2b57ed63807328d42d976306042e918ad5e37dbd81445405b6c8af0f
z97d4b57b1f7f807817b5f65b606805829d5e60007e541c34dfd4bcba8d988b48c1dbb5dfeca7be
zcb11acb75020616364ad2aaba846239eab39d84605fba3af30fc995ecfb2b475c5330bec5e299f
zdfafe015b11ce9dcd2e90e211164f06e1a6f88cb091ec3463e2319bbf3fa9bf0ce1bab3de95188
z02e4a2ef5fd137c6aa0797ac7ac9f67bdd367d00c1b65e256336a4e551f941f50f7b9bc6ba2dbf
z032dc6440d98edb9c893ef31367213bf08dc717fd5a08ade7cab5323d1168d8fca691c328bd7a8
zc898ab37a306c6606734309f23752925c37666291e140800e93aa2b474e3d962ee8b1838202740
ze0641959c306884cce5f1104f8dbbb9cdec60ed0415d135b9ad934b75e618ec48eaf6402320d4c
z5887c4a71615574137753178a784e921a83f25c939ebaeae29c65242a649066561cd6f75bc6454
z25c8014dea2af21fd7bbbfdbddf3f5fcf26412e7fec2c4710e0fe8c3aca281e0478b2b6fcc48eb
zc07cb8bd7eaf3ddf2653d1013471f272fc9eaff9da79f1cc2c91f09ded8959eb3d4792d2e6692b
z6e378f43b0c87745f8f156af82a31b59f0b05c973d8f5346913f1bf0cd5f3993ecd94cddb86d56
ze504777b792e369dd2200b53aa2915dbb97d512de19b6a21ecf0713422206a395f956f3ca30965
z9963f84e5bc3df5be4dfde406db7d14dca421d36cb10262c7f74274bd168a0e082de762833f024
zf2299bc639d16c0817df232257881ae93c50f6e0665e2e36ef193abb6815275ff7171de98bdb36
z159d38cd6dfdff66c113b69e585ca19817ad9bde461c687d72a9b559820603666e3f0d714d8984
zd2780c3dbd9e5b75d941329c7b5478d27e86cb414d9fcd14c430f5807fc726faf247f5c35f7330
zc5bf086890daefedaa693f4d0fb9847c1fb6af8b99f006b452442b500384905cb863122e5b3c1d
zdfa981c00e8e96fa80ae75eb4c9589f2f31d86672dba057787b49707f988076ad0503f0676df93
za245513760233622988db1147b97211ae4e4e9a34391c741dc7975ed1f6206014e7bb726faa567
ze27d1de2a02ab5ed9785cbc062e5788bdd7dddd16696f8abfcb7ff19f729209ff02a17df831947
z5819c19fafc59982b83df17450a6492023a3d5fbb896525302594ef853dadbc94429e42988c845
z796ef9a3648c9780d95bfcb3954ce6b10ee56fa41a5318e7794b46670c5a3e528be786c785875f
z8fc4de51bf08bbb30ccc4755f11afff09d8bb71cfb2b77e0d79122b803849d6749406337af3ee6
z7628e898cff5f889ac8264af517aa3418b2e438c1703de685eccfb25d122eee3201b9e282804ef
zeece8fb32bd63278c0327efab6d4e629c174eb9061e8e3769a81954800e7e703d24c709f292729
zf9561d3a426338ea475af6ba12d7d23fc07df5e559aa96529885c7a14c6c1099ac9d1ab3197f8f
z65b82e183ada2e46039b2e946a1b1d9dbdd475c5c05d3c0d5a271b83d717026749fc9c7dddfb8d
z6f62b83a4af448d78ccdff410bb83ccf164045ce3a4d96dac52dc5f6113256503b285bf6e277e2
z8944fa186935603b40cb7ead4e69cc2bc6a5660ff158a5624a2cd6cdd3a79f640cc0b9928cf1a2
z8f22620e216e363f9d4528325e184e984670608e1c09c36e93c5f26df511679bb910c315961b25
z66cabaa9c0cf525801419314ddc1091791c8b2275aa8e2a68ee79ff45d76d95794e5f91e44fa15
z7994ad348ba5d402714f920060393d3f5d9dba3fab7fc9db5cc9c4abb1879dd6e23cb043c2173b
z712364f672769393bec421ad1fc0e9673f6f853896251d1cbbdef2b091c9af22cf07f355083c94
zde0287aabdd6825dc08c5e2993114c4b8793dbf3c0d3b0927e70a9dbe93b200c60913e66399abe
z9019d1b1b9f1cd992491abb817b5a2a1dd1793b0316708e37085e2c38eb5651a45bddf9ca44141
z7416670375a9717319c3d45ede23f13a67d5b7274cda612874cc1a6c0b0d53f60a7a94a3d1a619
z996f56c4669b2af3a65d68ca20abe6c3f32c427a53da1d10ff58cb092ce342cb6a13546c063435
z2ed03e54a203cc7ea293e91bba058f954027cb46b2ab88d16d346428df25fb8a1c8c9291b68700
z93df9d49a46d8b0a10ecaa4d9e3d380449d9341243b41fff0e2f0d721afe9ef05c3c7009c719a9
ze80bfe32d16254b4522ba564b2fff049064facf7ef6a3202080cfa482d5a839cc22ec4c4e20426
z934e156252723cb555f4c8eec0a605ed525c1e269f0b3b8200a712ab5385a64b59fa2f03e9d395
z78f109f36ec05232bf73d9c68e4dae94bf7d4d564b2bec9a969fff3da1012086d4a69cbe432ada
zdab746085f979a1b8269d177491dffb7a03e746552ffe246a5d198cbb8ee9dfdb00e8040c018b1
z7d63e5b65e68f2d78499803d57adae2e6739ed271b363977f046fb15eac78cad95b5092b02cd70
za04434bebce80195b355caef8c469369cbf8ae0d49db4452156e3728f9c9fbd565e4a0affaefca
z3afc1309ccda760523f7c426dd8329a489ad73f71d8073fff3d62f26703783f8f0c7c6a11398fb
z0318f0d47207fb831e7112b25b24f8ddedff0d5ba945512e8afd983907ebd3ab38d8e4e8045be2
zf150fbc91b3f2c371d681b29f00f5b29da5fc53a672fea346077762e4617b52b76073ea1f59b76
zd80773793e0877d1f88b030dd177e10f2f59be19c491c4b87817b7d8550502db650f32ab91b122
zaad628cac9b47ef91048cfd9268ec6ab067e55a95d99e4474cec6e1f126585edcf6479bb018fca
zc51e42c018b9f22b9138489cf10aeec8d1cfdadef6528899f13098af3504f1db4a3d5d8e904b46
z9b87dbddfe68555c8b51ea7e580b358938dffd5320988bec3c58da1d6d9cd2fa576ec80a07b6a9
z4774cbafa7323031b842a118b40440866fb21c75c4a362de58e3ea6ca4f94f3d8fe94d055e71d5
z099cfac234d9f603e88a4a6c3f065da92d464f64a7e0beef364336e1c598e3da41fe8dc53c5177
z3434bcb58cc0e2b6e9b0e659eef077bbeadc3b13b624abddce39a524d6286630d557571cc7f5b7
zedb39c7351e3af59460c8e69f5e68c1e25c74d33314ccd2c8dcb9e33580e3a425152087f48bd6e
zc5e4866a742581b7963198d152c1f8b26557e68a761f2207fcb8ae6b08a23a139eee186e9caa71
z2e4ae92c2486ebc6797032fe64a605251aa206f43e8c25a8179e661d81ccc51aa1100ed3b74ea5
zfcf171af1bc79b839086c4762eb9d125e1ac4412d2a65ce79ad1643dc3b9fd7f09216258a92cf7
z7dd1c5123b59659c2872bb326205ab75cbdc16a88983c9360baba557a7d25f064294530eb9a590
z2883633aee413b496c0b255df24b4e2ce1e3e9772200ed225c9facda19bd001e874eeda249187f
z669f263fe157062d5b81558b9af15fab15f85b23b3794290141c047f9e37ef9a14854f9d40a928
z680c677cf82fd1136ac3fb53608e9c51ddd9b667febb228751506b756836fa4db3fc2a1a69a458
zba4331eb5f88058171b0b18f28549464b03e902e00b5c2160de7a22c6c478d6ad85effa66b9884
z94f7b336aae71347c05a93fadb3a92f996d15f8c0a0e76b629c9112314c815047bc93578ef19a6
z41d1da4856c8926b2383d2536bfca01b45e49b176cd3f53bd8de3e16fd168233a41f4565715ad0
z05be0592d2692af315892faa0dfc1ee9ef9751e25eb2fd6a8eb63de3e8ed784b3eb9cc784e89df
zc6334d396f7123d49e91a744ac25ce97aa0ef24e14b747809cc58acc2bcc3de1be120108ca26ac
zd9fe3c8480ca0e8300a0ae857fd2b16506c2594545f3e0c10d3f481be7097ac18389191467c30a
zc150e57c54201fac719e09fae9e954512c62cf521d1f746166d204795af1b886a8301dbf0d2d61
zdb74a9010c318a8ca0f5e0289b2ed42d10253287b251d9e1bc915e63df084700932d8bbf445019
z99eea2dc575f1312891dd77c3cb5f4df643a40041540e744945273c4698d0291690084b9d653ce
z35d33a7a5d1eefd0a0d1cf1d0d2919ad2d9a01a3e858a8a5830e4d1fa97f14431eb50bac7f601a
z9ba283e87d11db9e1db6ed7e80a6854f46604dd72bb98ef70140b7b66b6f245a6b9a457399e222
z7232ff5a77046ea71d31b7e60a9cd96d118940b6412d66d6eb88d94ed22e8b674a851885b279d9
zae494a9d65ea763309f664cfa878eb87d079f7d1905f9efe45ef6ebbf7a8cc718c800b46de6039
z08db497ed847e307434a8004f31eb0b668ce5dc9200a3daef1f05286844ccb5a10f4852e7b9934
zbf2367804ab1da063d3c749f9aa286f73dbd4bfd5723e874fd80f2b6e7b2702339c1a88d2354b7
z3e167a507fc4848be87c252c5aafe54d9c2e55028da2af92cdf69ade28a90a2bf57d6d5ace93d0
z22cbc6fbebbd56edaf19e0400af497896f02f6ae62caced82368b1c938e8d0d447040b40948e57
z552769fb51a4ec643a721496fabb0fc0ea5e1902298d243e0de0c26c4a5eca053e8c8f115c4e18
z5cb843d773b5eefd43d988ebd4ba86222935ef26137e00539f363ee59c0f69b289496bff5d3a6c
z630fd3ef09d1804658af960c17c5230522aa1be562f3142179613b5aee6b6b1378fc39c1191a0b
zc35d42a60c8ae4267336e7cb681592431c18649e82fd708e71c77c5424a6b176a0d6e62417afd6
z84616d7e857ecc96c9e8f08b06aa4bffc91c8a6f3afb485ccb5350da0d039a151c927134bc7462
z739d32fcfca61ffc6dfb4104d50ed7fc11a47f8ae9b3bb9393194d9e9a76152eb8b009b5593c30
z4fdbadd43a8c1650400cb1f7993a4ab448a507d85e1958247f30111cbaddad603bee97fb418bd8
za3398c5576b12ec6dd32c33e5389fb16d66bcf9f84e31c81f5572d4d2e5fb4fc5b286cbd9ddb1c
z9e7932afb950d0f6eca78fddaa7471a8356027ceef4960d542996cb55f4dfe8c89151488e4a36c
zca04756ea6003a7be9106dfd08c2c2c18242541bab21c649d01d8f6f62d442497b535c134841be
zbb9e30d4309fd470d9afdccc2c4b2205318c04324fd9f473380e324f710ee1ac8f06097cee209d
zbce2f620e10b62910f0027b5e59e01d94046cc87d674ff63c1ba1a7b1a6768e7215db61c967c52
zfff0757406e2df9df0b24a3145fe742a520b1a0ae89d00712c679bfaae92c01be1c2d2be3920fd
z8d88ebe081e67079279f944b50b7bb807a9ed4467e3193bc7333bfa952123db4c77a9ee228c50a
z9786fa83d532035393e4fcc0c8cf1bc25a2de09d7c8869372ef80aea0a66213dfc9f3c3161b72e
z6d61f98748b523bf50cf308db2f28821c5c9df5745b691b06c843530a01f92d4f341010932fdae
z76f029537f64e75ffd242b2d22c0195d6023a67657f742612013ce81817da43002816c10a30781
z2a74a7778721c8cc513bf24fee0f427a2f312328fc17905748222084bb6b9b33b408308bd15936
z227c13b2d29b398a2ecb9c35e6d52995fe6711e743be59e9c226af2c4c7e6fd04185b1146bafe1
z86d80fad322da0a61b39a4dbfbb417cf79128d592b1cc8579330f371b76307eb4ebed6690888a7
z6be8d1e589a366554866d9ae1e7f1fb54f40444483df423ac9f368bd96e560eb10a61d645324b0
ze055b193a2116a08d8a218935519d96a14ab6172124dc876f8c74646477759170bee12194bb122
z592342c092a222b45ae4b8e7fcfdf3a5af2ce284109dfc3c1a949e58906323f14c56294677589a
z83bf7502ebf425b447f8658ab354b1092661eacf016993621ad488b79cadcb8fa5a682ae2f5d10
zb1f27f97fad1cab87d2d326be6162d62cd3326bb6f970d5c2c15dc5ff647163fb01914f56b4a46
z11cf81ead0655223513f25804758675f926a0e9d26c2161c534b88b3903914b541d688d2b199b2
zcecf13ddeeb5ff367263fd6ab5437436204c801b77fb65a808a358c97ba3d26f139d76231a100a
zdb5fec8f29de21102fa530c56e5296c535543133e1b7c400841a4a6da981c1691507cfff44b2eb
zd771b32094b241e1c26ab424899b827c6f02e369d4fe0470d995458b4f686de68d2b4ffbc96819
z8632aa85317ff705fca001dce7c96295c83f42e3b84b2b6bf4def03314f0177c59bef7f079f130
z891fcdf28b013519a60f121f19ea302ffa89ec5f505014f75c0569bdf1a7f25ad4b2c3d2ef313e
z6c4e2d1ad183dca9581906975de233f82d724eef6b27c18d5e3339441cb68f3a193856b73c953a
z499f3e5b18e363a9e06ffc97224941942bbc975908a7cd8791de9a347532575754b13215ae1d3e
z641c6376cb1f8f134568d54312ecfb4fd61ced8938e47ae18ba7a6d255aba48d293f8d13d84dab
z81a2940ac8e1d12080813bc6af57c987e72c2bff246c4cbb23c17cd76f16df24cd948d94beb96c
z3693a795d732444593ca1080b8e761619e231a6ea6e10c20d3770a76a0471975b15ef2088afc95
ze359b5adc9568d1a1c95ee765c823f1808a83ebd73edd7f78342a0f4ea1a037673664c41a8ecfe
z4cad19a1d8cee74d8193d1dacc18b113924f8495975fd0139f40a1025d9df0597e953a3e1e5a14
ze0736006aab9fee4eceafdf9099733e8818549d38239447097da8361b13a7eb6efcc736006c460
z6f587a8b4d66aecb1c44d2fb5cb1468ae4a7336bbaf2d2c944d2fd5a5a1bd1aeb2267576a11961
z112d0cb0618f87810d092d6558c34f820880e60800877f0a52e2bfdc4c1ed9a7ec0d5ec5d2bb37
zf32c4cecee56a9f9a510bb915392126829c5fa89ddd8446989cdd0deb8336f2933cda33d16e7d2
z98dd7256e709cd336d930245b2467e40b29c4014c013e301fc88a6faec5593f02b09bdc6cc0601
z9c9e8f4a5a78266428e3ac124ecaad087d790509394fb5a9e3ee1f070e2547f20dbf45112d1db3
zb339b6a7f149c06c33682fc47a6cb911d993ea59bd53c9acaca2b86147384dd72a1ed87a886cba
z617828f015d542052f76442c82ce4c52c1369b7cc47e6aa962e2e37afd4529703bf06b270d61c4
z23f3df86802e9039e87dc534e5efcf4cbbecc2a6928f083818b4bce5ac1b057eee468c6cc3b37c
zb0f6f42451843dee91c75f0b8bac5341cb4815cdaf11a1b1de85fae911300f73f46f05d3ae0c9d
z065e91479257a732a7e0c21af43f529330d77e8db9725bd1e06202785b1790b4259ee09f062109
z8b4e00543d6aed216470ff253b971dafae3eb5a0d2d9993c42ba41f0143e6492acf560835e9886
z355812181f51b1ea2e5b730140f64df3d870671dafd916e601665519367cfabd4ee7c399ecf51b
zf03079ca7183df23904ae58f92d440301f63a356aa293fc69b907cca0e3d1027c1a056215dc0ae
z7b1dcda65d5e51bd24001ac4a8e0f27c02cf98e72534ee4c81ccaf0f59bb7a3298375ca9fa3b4f
z09e1b3df54e2e9a5e3637b5d235209a9386ffd70e685cf0987d09b49314a99bf6b933018108f84
z0f9b255addc0f74b0b3dd4bb1e985eb71d67bc46dd30bffc3c0baea376ecb33cf317d097001383
zeef74bf2c45570b700521155ebeb32f49d3736f157b094986c2c386e94a059b118a9bcfb4226cf
z5cc8ab8b0f204fb4918d69e39869ce5eafbb2446b22e7df333cca79d93aadb71dc91b4c0965092
zdbfad695dc095ab7c89242bb8c801b410d37ff8394a5f8d4d6ff50b40cd76433fc86ca1a65d94f
zc9f47345e8c19312ce55a71f82dbef9a7e40b1657439c256931ebfe1504d3ddb2c2b68784c6e4c
z77fcf057e102c44c32410a2c954f6e8b5c9f4e75fbce660d25414d4c658aa7e2e87d4721206a0a
z13fec4d1198ea1e6e049676b1c130c745bd72b0682e821113f7aa8043c724d7bad55c232f18503
ze607df093c88f5bdfe8e95679b37d8de785c8d0eeede2ef0d99af2698ebdb9c599f66f1a712308
z2d45b5d8a50c904b525a45e507ef0f57ea45de31d87682c747be8528eda9a09331348ce13ae846
z51650e30825bada9845e93f1fda623ca8e1795c284889ac881d9814babd17b21b0a271d8b39d94
z5c2b93fcccdb555c76acb20b6ee82d3471c84be70c5bcacdb33dce1595c7c8133032653b13964b
z2c514ca8ab75750f51506546303b30f59d7d7f74c91e9194e1ca63ee163ec05352c7c050d3f69e
z1201fd5eb0dc7a0f6fab3e996c9607dc89d56b13a75f3d89ebb56285e3662cb36548cf56d5d161
ze0bb33784126f3be1aba60410f95cc1e329f38b4eb364ccb1e32f23bfc8f4f0182102d881c34f0
z6fb5449332ef2abece24cfb3bb659d4dd980d1a2e4a97de29bb86d48a01a285fc26776a422a194
zdce6a3204b898cee049dedec5d364a42b8d529183b3a66937d9931c24b30706323f98249a699a3
z055ece73d125dbd9e4fd6c1e4aa0a99e7951eed0abf1231b974b86678ad63ad8b1d1b26f7e7dc8
zc6cbb5613170c3e0c74bb0099c8f4828baf95e6e7b1e5b8e49f895041849cd3d1d71eaae027d38
zf00cc6c67afdde247dc5431d324a52b72d7052954363c3c1cb3260d4accfd381efff18b1f10f9c
zf3a6a752b4eaadd338dbb236bb65e14ce3e9f81f6d6e25473dfb99c37c79233284c226e6e70fed
z932b5bcb85743bf57362af421f9f4c7e0d16e34491c5c6d5b26e92b72b218b7c117a29d724a9e4
z3b2b1b7f353811ae5dd9450a2a98e7a0b022820e1c3d14996c22e3475dc7523e007c587f799cc7
za8c16103f84179aba991efd239f7d8c31cab0c06a66a662901f57f670bc9b5d59ff8cfdcfb4df0
zd7acaef0829b7b98a9c0d19146fe36ca12edf0d935de7beaa265e9bf90d7ba97f9a7b422f613fd
z530212ebb77ca36575cfe9612b9975349d1ab066f3454c5ae6dcacc16c6920f7602ee793a1670c
zd66d80f1336b58b367e97f2d4b407fedea1e876c477c57b74e868740294d9245620cb40ba372c2
z1cd29fcefcad355f5bf6755819d71eb90a15550bb03dddb8254e3a4e0685ba749b1642f9fd9583
z7df6b88132520133b832cc705563a7d570288cdd04818f2a98c04494e9565fd001ab9a3c52f9ae
zbf362dc89726984ba9e27462c738867ce1c2e3c33cf88c2eacb39abd7429f369661cfe4cce1857
z7b0a294e8b5556441b0d1fdd93361c21b881a931c8b7f721a8ba969845618285a0ab2303358125
z90ec5c18ad19182500cd391fb7ad22fb7db0e8dac0c2ce0a461ea9fc49b8fec79a67abe51b8551
ze73b50d0f251405687c85d89c8ff85df30369c09d2c2393e55415c332ffa78b7cd6dbc08a8bc2b
z97fe86e049fea2b5e7c38f9dd7d45a0c9f9db29c2526e6074127d34094f6d77a5f539d1dfe85eb
zdea92176c2168afc3e13673bbafca984d712e9678fbfabda829aa9d298ba71235e97208bb734f2
z3968c2bb67f162d5e9a50548f3b3c6402373258bf6648dac2143b1bfc0a5faa67a29e60f6252fe
z6aba934d7332428a8dd7cbac1f5c83d65ff57b0cff22293784bdbb017ef6309df0073884a361b6
z19ede7f33474977306655b01c1290db33bf1fefd977ef68a60e39741da3933ac11a3ff6246b7f4
zf44967cedce6607a97f3a5ce920f41b13b22a9d37f26962f4f4340d01950a30b8e2f2c054a7b5e
z91b887d959a51188050a5de51f5a2761fcedb0f3bc6bbd2009297fe8e7c8e153cb45092afd1959
z83e229f7a827fb38f28c32d8009ce38d778fae6e41d0a98eb1a6a997601c4f8f84c16f0f341ae7
zfc05d9cae284f15268c876f8cc2d4dadf314c2469021bdfdd335d886c2f65a9c7bd367c41b6215
z3b78a6300c7736da40459f54822e645b3eb88a5b5a06ae6b50656933ccc55be16d31a26dca9409
z99c870f9e35c399070287e2c1a3fdb0721a623c511bf0b5d583dc18c78566755679d94bcb44796
z06012ef7f4d902c7be1a9578a15d69270792b75c132c7e54864d415ff1abad80ecd9105919771c
zfb575a66840abbde9d6c28a384d2e39fa962b43b34a5c87b7b01d06d7ac89e5126fd7682aff8b4
zd9088dd661fb275a414729d60150fd3d829a0224441c8932a199aed8d4bc0d28a2ad807e6b1774
z3d8a6c5fe0f210f2b6d9ccff294261cc372d967af10c491d9911d744506c4caf7e2769e7c88af6
zc4e686334e9fc8fb5286959209906c456e2f4f4e24e7bf003de190b01eaceeb3ca196df2dbdc6c
z08cacbc39b0c3e722ddbf41e83b29219562b3aaff018006a19040fe0a7644f5c8e8c9d4687cbde
z58988c9aa40232554d29ffcdcf108d6fdf8d81326a1acebe7ef23432febdfd1f10afb8fd07c099
z5e24bbae5c59a38ee19bc14334042862789cda8c58e2c1b0a8e56af0d2b2a94bc0aab5545075c2
zaef11f7fb747d6d6a0ca76169b1a6c389165c5faa9da536c91ddb3876dda70a79b3a3202db3cb8
zad54c4196fa023bfe23e9fb82649b7ba9ebb995b5dee715ed20f57057a4f02b60b01d621d78347
z27ba008114b5f77a4c89ff238a6afdd587609583a689b16b54ec848e7b934572c0bb081c664367
zf46766f1caf68e9df6e6c8853354d416dc0f6296e87b65e807be5ddb497fc49c631b310b91d021
z5747f9131e789c447109dc0f312c8dcfd15e8a0a4f588498d8d5291117c6f6fa84752ed3ee450e
z91c8502a2969f7b4b287fd45c126673b97d07e92258ef7e42091166ba0a260ad59eae5ac4b5b31
z5d8b5f080f8496ead4215a51a34a8b720aac5fec925301f36d03e1caf7b2581f39ef983a08be2a
z6c757ba6c5895d3040ae8e65c93ccaa20a8ed60c3451b0759194624582e716bba71ddf0600c923
zed7dfa117255f7ae30331e1cc288304680bdb2bb0515152e541b3ade7f7d092f8d46bed18461ee
ze410e74bef0c4f03357c8c793a27e9e1df583a09d306c7a0f687d1662425a283405215b3fd4cf9
z2822655ffc2b0373a342ab3e854eca247f1cfd2c54ebae8f0e0b3650c91a090ab7d5a43f4d8264
z2c0e18346226f19133a9880ebae74cd7f96d41de1c28370354714fe433381c0581e73f7d0d2069
zef1b269d690a92179295d96675981a39d0730b5ea02c0169657595f4e36c05e159fb4f55948f5a
z8c67cae27ee0eb04d8f154cccce3bb75618815767c05b7cba5447edd29f63d5b1116113e911821
z74168adeaf0864bff820e80f6d3bf666677ecb2c0defeaa2986eb578285711cd0670bca33b8699
za8b44d6bae8e42db7700cb0c5c419b816ee68b69086a0eaa165d8401072addf710b9b7ace96d14
ze7523653ee8ed0ea2bad2564b32ae3bef8cc71250d2602cf18f78ca948529b727ea65d4b59f5ea
z23cdacbf9973b59173bed6a3cbfad358a2510d3810f4e6b57a5b17b4a5cf141b03e5c11fd70a55
za60217c3e4e88fdbda46dea81118de3dbcfa377b3ee5c98d4459ac208ee4589a2cf18c244beee8
z1382bb4449edaeec712ffcea07b0a8be70c8aef80962fdc593a24b04a32dbd9ab9682ef9e74f74
z8d9d4bbb301842e7ad06f655656be4e2f881c22febeccf1e5dab69b1fd24c85bb0e3ac649ee2f0
z19790ea8b3b4e780f72118a0489581b0db01c25720fa3178e57037995e0a4072e032a62b61cbb9
z11f4667e7bb8b86ee54abd8a58484b888cfe8518d58a4a5b326e2c133b
`end_protected_0in
`else
`ifdef MODEL_TECH
`include "qvl_ocp_logic.mti.svp"
`endif // MODEL_TECH
`endif // encrypted_0in
