`ifdef encrypted_0in
`protected_0in
ze74c34e226135848fe16db9ffd31815111b6d7fb642c521a3f628cf6da949865580b22efd062a7
ze90adae0e65e66a2c36a587d0a790699161455169ed55a01f2084f11770a774ec4c588039b380f
z6de9c5084882a40b79a175f5c2114b2b6d78b070cb806e1c0aa9258297f4687ab308bc470f0040
zb0b1de382961eeeaf2e279e1462520fc31c119af8f2b214846f56c2b3cd2eadbe4099496abff18
z15cec83ec4a77b868344aa20ba7360908f5c0de2a79abf8b3534b883bb12180f68b5d4beb444cf
z3fba8f13afb0abfe8fcc4294810f75afe452434d2d0f1166236c82f76edf1e12979f04bc35693e
z32ae028996dd85737a8f5adc1ebb94f39c940246e887647b64782cd7ab429b0544c173176cede7
z01dfb26b1f73408344a52b7e1f117f12bb9c8077b34876c2e6fdc085981637012dc9754765e1a9
zc512ce062e0b8fb16a214591f5c81e1353b900a611fe1f4886b57940b41b7f2ce99a7b84b04b90
z916f717e73bd10589c81e207ed77ec660a8cbed5b487fa50acde1b055c8870bd8676023f21ddcf
z9c98cc47cfa2d654ff1365d1f45035a045a66c5dfa827905026201628cee5aae21fb892db766c4
zb5b1406e11aebfd6dfacc9da5ec03b70c276807a3eb15e28ec7ab1dddec42388b9424ea285623a
z248195c9f894b36317ca6e59c86f11031163f5f5e0af432ad71a370b503d5afe29967480e0ac49
zcf7c756f92650aa81b43bb5505acefc12a9333c15090c386c323f8cce4e7934214caea9fd9c42b
zdda79bee782f6c797ee18b17b0c257e45bee7908de093c385d7e8a753e689ff7fc8a8c9e7ce08d
z05cb3d56bf84f1fb3473afaa2d473467ed0a852501771349b43fde42b4344a1328f0b9488ef772
z0ab2e71ab13ec995ee041d04202d900d95c299a1c207aca6e4735d4f3857211f278f025542d047
z1120c7526d7c7aca9b4535ac2a7c89914a071ab6e28ef5a017369bce3e9ab2a40b1045e640a03f
z1eac01f38537c460592b18e6569eeaf3cef2c2394144d0b4682b5a48720ec74e4d0b2c6180f2e3
zb86b55096a5ef9be48293937fffbe514105bba4c72b420bddbaff7c98716faace082ce2b7270d0
z082943369f9adbbf070172be89ab7354b521930c5a900dc87238b1766e67b7a0e1191854639319
zdf1223e075dde8a5cf288060271fb236b0645c68e01c0ec3232b83e1cfa0e95b47ff1652160747
zecde91b28ebaf7a1a398cd45bce9bdfb59d8a39c019333c8c70a92757f3498ba94a1700a22cdc8
z871aa793ad3267f5ff895ad9188610226db47921a6b2373776668a9b2bb5daa92fee02383d142c
z8b55f881e25ed88fb59ba9c730d78bc55a0757a3afda6902bf697868acaaf20ee3ab8a85200ac6
za186225ff0211433acc05f5df1c2b0c330e70a04bdb8ae144ddf093ff61e1e143a2dc7814f5445
zda60f461b3cc96c31c3ffe91af592ab64af298369479c6402812a8f0aef1298bf74b9348aad66d
z7096e30f35ea4205e6181575b95d59b1704055c6530760412ce718eb5b1e106fd6a179f4165d39
z8b30846ff76b49c610f1199062e473940596e20516e2a4d93413f9b79c94cad57b5fab211ed856
z7548faf36b57164d3e598195148001d10a1ee6944d21f69599b7b4002edf2846bfb91c88304bfc
z7c2ef11e4a5d4955d82d2f79e0f61ce32e3e1a32d73c6aed2779ce5d7057401c0b53a1ce86b67a
z14dce24a1141fd5577a376b61629ae692164d11b92077cd1cf211a69967e8e2507bbb7b018c668
zd3a4c8bd78ccd7e3256918367dbf654b6c0c31f9fc3d170253249aace4f7db3b1940d44f44c9e8
z4a1c5b5ca99c3087c8b889dc4e453c650040afa921ec3bc79711a8afad1e6700c6508a487142d6
z1b495436115e5ec58141e54bbb74297e058d57b8bfe505d384b0857689cd22076b5212bd3ea481
zd881d2594bd9829b0183212fdc49fd49b234b87dbaacf31472edcb89d34babfece7ca2050259f7
z9bba58c8d989b4e472092233d94b57dca47dc69c547969363949ac4e45dcb38c20478ad0f76e52
zee812be562af73ed06cbbd1afb19bb37840e41305d5169047d9842b7f850acb1cc71924aa55fca
za56ecd97d5d2fd19bad64f8e43fe3326b6e2ae877a910982d87bd0d607ebc539576f81096838bd
z032f50eea83ce5060df70f577ce5163a92a2bef3b59ffa4aa098c7a00b39ed48748b7c232b4e43
z1fe32df17673251debc24f699efb28168714094231f3a47a9cf70fdccef91cbc3882974cb5a59c
z9e3e019bf96b1dcb63c025425e149b13932511123c2fdc1b697818a84f23c4b899f717dc37633c
z71a63f60774e9a418056c6156492e7fe7f8af18daeb5b3c81a2bb7263f7545eb66317a0b216bdd
z1d7fda29344c9dc228f16f133333a1c4e471f1cc04aef3f90884acefb698424bc6c87b09217bd5
z868120a3b350c3742543ad1b3960b15b3af67bacdadd7fe47bb8fe41e96d14524b97a1e88728ae
z25bd8a4f76309d1ca4ce35f4c4d8d78ae5411bce4f761323b91412ff88ce7b34795f25e9f4d30e
zf4133861f84353669d9a81c7dca7ee2b306a62de23f17632d7792479c2d5acf9a6316e0d5d93e0
z765be2fb1eca748c2a6645205af4c8d9d7c8cc9a840ec8307d02118facaba0388f05df3223d6d2
zf2defa5dd5796e268630731f48d471fd9f16a9ee151b5825bed1562dc5160424ce35fb74015be8
z80db3721076d61e2ed644ac939344ec61a33952e45998f621994ed20760b49849ff1a3deca4abf
zba334e4ae5dd7d794496b458e2e9ddd582a41d0ecbe5e45069072a209a08cbbc5ee4e5e6f5512a
zca68a86293df4bf3881f737a33d8954583ee4fc46fe4e7ba3a8867ed88afe153393cf470ac4d67
zefe5cf87a143e7abff710ac12309084361b46170d540780dff3fbf21312bd3a28048e618cf27de
z9f1807d2815755af6079fce1c2a5531fc98f51e91092bb8dde3f55e9832980b40a0f7c0875fa25
z61be7d40d9b4bc160cb8d3cb144d916d25d3548123059a183d79a9a132af804a02cc548b06452c
z63b3aab32df32f3e74e1c677e54cdfe273eed1856eb8c5b033752423c57ea0c4a22367a539d0fd
zdfe2a4d751a91c0ae87ce35cec2e1c8fd636a3fc922712a799e9ce96485d9dc975d64b1f610c2e
z86aed5cd184133dc9c19c446fb2d293e67a11d04d84fa9cfec363992da7d601a362c43dff8c467
z4e159cf9d05011d57e18051dc44689d8451d40d1c3df36187feb3f77a08643779bb6a11068ad81
z47b4c6ee2d0ebada2ae266464ebba1e4383f6731460493be17493696aeb992ab5b8ca735154a4f
z58a3bacff7fcd22d75970d43a1bb0b1c2af32768c979667ad2445198ff998d16c50494177879e3
z1a7d0e264050fc7395ef8206b590b8ab6cce2ca633c1b2f123d227c33da2761f99ba8b83255075
z4e658ded24e3afde7f8378d2058bdb094dc9e9f8262121fd556e616255ecf65af21a134d41b4e5
za221a31670ea5a00a43772533f91d1e4dd6fd2b007c28c5a53351960febde743ab7c70b47a23c8
z237ec7eb3f584f34abd35a42c8f45bc822ce2e891bb5d9ffd43c6de71a4ec488b06c558ba64593
zedcdb0d596abd40489882279abf38933962072aaf6936640e20714196331915253e92c8b0827cb
z7751a3a4c6563783a7cc669abee44fab4e178ba0e0ec87fffe5f8f36769aa528668bc37aeb2072
z120f0cbf6dde0591b0e334392e6da44df36e7793244017c2b8c7b2585d3a8d3cf9f9ecaacfee1f
z65e0f131f4fa0e943a1543499cbaf5cf4b63749fdffdcd757b154eb9cd147e020583a3717e4e08
zb6ed41f7bf249bb21843904694939075655b0608c63dfd08d8a29ff1cb3b0f46d96cbb350b9872
zbf2dde0c225fa45f242e4becf4476649b54a78cda685c5ad86f5c5d1d9bff7550fb2e508ad8211
z7ab7e53540ef3a15a044672dd652f6d6c8ece1e7ace5cd49e73de7decf4442f9257d459b0085f8
z83bbe6d5f6f3edd894b57e97d44188653972c61df117c1245db4a22a39d25f210590d078ae28f8
z633952c85bc533201dc7e96c4e8b257580c2e6e50141eb926470091530ad0469e8bdc6f6daf9ca
z01218f849e1cdd8632ba031e7a27b80a793672d6a37798548fd79535d518231b6efc99de64e112
zf2325b5ef6a821abbb71d3a4639d677911f4381fbd73660a415120f4935c20e8134af24fd7c723
z3a341669186acbdfa50b066b650e10515edf29445eb172b500f3d2ccb88d323a28477334d5ad25
z0d3e63c306d01df2b67a07182602858736b5d2dae0d2a4c5d463eddf0607c3d52fbf97e15e7b47
z67b07a30ad33105c3e8c0964ef3c3243b7760f251ecaa768cbe4856eb856ddce46d0f43213439c
zacf5d803ae4004f6b04afb777ab5f063f70b80bb6f5e6cf8e8b0536dfd2138366c7c3dccf22be0
z0f147884d0b8def890cbafa609482aff6fbc2ebc40784b56701ca796d1848537af4b87f0dc65f1
zd2d74ea1b3a6e3ee87b92296b9836a1022c7bc196004c96adebfaf0f87ea0fb52af1a56e536ef7
z11f1dd01ea9e1b696c3c6186884697054a2e41208164895e9ffeb47e7e613368d17b74ca396e85
z1c7a095b336b22b097777c1c681f34d0ab22ebddc6b0da7447dd755d7c941e541b979fcbf91544
zef74c354750498fea2a61dad8d39041c91aa57cf30f2f883bb93ade04943eee32f942758678424
z6996c64f043faf459443d2c95d5a628ad37f9846ab230c6bd07c4c21561b71d883ac58c651ff5c
z4c1ef7b6d031da343c3e19e9801a98c98eb836cb807bbaaff743e7c2a6e31b24353b19075793f1
z4b44d53982beeb7882fd6aab888bcd92d7a93469ef9beabd07dda7c6d3bbd0f929f5cf97b88029
z57cb87634f33ceda3485c798b1eeb89294d74b103ef55c716e9a2c3bc05e86bc80086ef39a6233
zbdb0ee3ea839be2e7743c815d6308ec8cd1aca4e7c7f9c4dc567a092bb66a14a6072f7a9e76d3e
z37784a1c07bd06e9d34778de2676821a502057f646e0170e3d9933c963c5f67b4e632426c41b48
z7eac3a33a3593fcd4ed1ac70a060c839e3e7a2e1f5d71d64f7816a434a4e905898cd9e1542e9d4
z3f7cd9970ad77d68dce25381b4f22f649dffe6fced267d2408493b191df8e36d05a9384874c681
z4a4a0a7430d77f0e57fb1d40fb328082985803b27383405cee11e10c32763506434bdd88094711
z5b9a351b652a95d06b9f13737eb7995efe1075b9b06f89a7ae9367759c384a25a91280e439057c
zde5d1e72425f9eb4f967289520d1ad781a4d4058bbf25f74d1ab9640e7b59ef3eab0efa984bade
zefde8dc5cb9c003f79e8a266c8a7f11e5aae3e9e3126c3bd85e6ed92869b07c4ebce25f767581f
z1d9afd87b6f0bc5dff30f3b838abe836bfaa073a8f80d25bc00db4866bf7d6da72cc2aa55d47e4
z612a03a26d491b0f60d07b83616bb3a73701c69060cd3f6dd1da9e13b3c8d04a379038c64a4754
z8e284b1851692d4cdc5fb1a1e4a4a930fb57708ee599b9a4da4e45e840e98197ce870ac3d5cf33
z0de1a920467c7e423f66179e0c6fa242bf2bb20b0455b9759440867bb5699121b7cfb119e3cc49
z4667cad81e1b754a280d3cec210265240e325a2abb6adc2468c5e00bcfffaa0027bfe7edbe9e7d
z8db0963d9267e3c665e11292b4c48a7b2e80fe738843317faba854e0f6981041d9f8c9869370c0
z2d11c603294a545b7e9ef1507e108f8a1c396d0e73493760f6ee75fffe2195780dc74cf64d1c85
zd66f9b4ca6d9b854508f10bc88c79c19cd319ff2507bdc78702511403a81309757352ac28fccc1
zb9569b1f0a07b6790e6a83d17a7d8b699adfa9caa8be2c3c15cd28796ff9e3ad7e0c4a8b9755aa
z7f7326322d1a7784ec70ce6f808435c358921499ab4d309d28976ec0e728b3937e9f0b18e4e1bb
z337e114a6e0b2ca68c3a1436cafd01d95d16522ac0c74ebc01bfff9c3a1c1737400ef4fb04f6d8
zbe456f37aba562b35b863507cc0a622c72ca1b2d2ccfed546e3f2a42e88a0c792f0d69a10fc52c
ze31f0ee53f0d6628c5af61b2953df636eb103a192b4abc50628b475028638e2b833785e91de59b
zf76097c86c838750530b9fe7ce34ce29fa17fdf9184ba52798507633ecc79e3138381e08a22c06
zd48f37b0acee2c60b23f423947c8f37f9cece8712bbaaf47dcbc9310ec77d2b36b6485b6ebc963
z3e9105d8cea29e4347a32757af5e75467a85dffd54a552924a3d4063acbf011e4ddef67873d3c7
z0bc898091081fbad39c3d7ab8e5925b55622e640304dbf3eae9ce08557d944be2e74434a6e0922
z5e4d2e2a98209ad1653de62ded588d481e9b1da422f3fb6e9194f4191cfc530cb0957b33db9538
zb740b362b98fb780d8c65ee35d3da9db269a8317dd88a5264bfa7cff8f0d05ac023810c0e8a2d2
zc4947b4d5da75277a2439edc649ebe52ed19576f114b5bcab36a6c2e3b9ab72459d8f2df4743e9
zdcdd5a78b051e4f77babdd7bdd0ec9da6d9b1de33cecf1bcf11c3bf66c213fb745288268f76bdd
z9eece9b67955ef3fef806e3e405ca5e048309eac80f6b2da0a41ee3894a054ef2a5c75be6a7d08
zdd2dbf7019143fc98f92388a8a071abe6c0910884b7961b527b440b39c69a65db548974460b29d
z040ece13dce55b694facae69a08f66d84cbe71aeec55fd3343affca7b6f6f3141e761f89f70d0f
zff644c1e4e38d0a70e0663118a7770d0edb3f806791d39e47a7ce166e2c246be9b189d775ef0a8
zcdb50bd5a9da5512646627f831702ac539b9214db66697b0002611e274bc981ab63d92dcbf6a49
zae70024ed43f2337cf590672048ca30c6dce94e771e7d60f8c7889374937f69ae7734f45e587c1
z88f04f9f968b684e63041a065cb6e7972a0a8bc3e02ca13a23dd7d7a8dedfd562a64667231ff38
z8faa3c433885e8cd45d78f997bf597fee5057810b4b2e7b994779c858d2c49e1ad53c034dcfe13
z9b1b975ff24b8a6720fc350bb71558675bdd6bf7619152595fa169ca038c0cffe22e824a69c577
z836723c4701a6002af964ce6797e88a46d9606bdc86742acd1e73c17ef462d21c7655dacc0f9dc
zfafe30822dd6e655b4a98cb6613758364558a165b12e90701c0efea488c4c15e30622fa6cf59ce
z6056ea96e80b1e41777401afd733ec30541e80a24d561d3313733abe23ec63b933f41405219038
z389a0f7afc5b06035f63fa4e8a1ea94e49d4b14f2a3aba384cade3b51620e3033af22977e4b577
zc4cbd8548fb89b5b6e78667ed86e9bbb0ea99feb88bb6dff5e05810d9d84deaf7b064fc7c3e264
za97645ffad44f04e87101f29e36d4e27573b7b2c347d3c29e414983da85a96a91666aa93b7815e
zf38496231cff9e0a928ef3823c319767c36740e552fbd7cabdcd0b16ea6db08a73e3bad2c5cc3e
z71c9cc3ae96f482aa930cfe3f49333a9203da56eb22f34bd1923f1e7e480ef3a8d6d8b1d745611
z261415a5606770cf14f1e5524bcd00d478840d51593a9e07c0a595bffa952e79ae02968d83d00f
zfa9891e54e4c08272c3d405a0c34626adc13da038b7c55647d9d75a614e91d045d6b22b1c3d909
zb1e76dc3fc0d2ee8bb65713c3bec546b647e26b054556cf0553bce8a5fa0bb509191db6a202543
z84eb408ffa731207b2df997b64f2f027f25b1c6621a56557d384138564306b2c2f5434f79cb34e
z70f5aef74d6dedd8e5c54a421dd8eadc7f1752c8d279ada75eba21dee9090155b1018dcc27b8a8
z458c0fe3d5061cce3dcf8c2ba52895955adf5356d079e6b85d1fd96fa0ce658a5bfd1a5b674936
zafd99e01ad6647af9fd32d6de3717cb0fdb2652b0f8899373803463c004397abe0d40af82208aa
z2e9d42946e312ec81590de4cf935cfb71105507a339b1a1ea6ed6b0946efd6b022f2de01557414
zab255b9947eb244d73b8b1dec99625573c6f56db7fc7d7b13dc79ddfb8ab63672b280db9e2cf21
z37f4ed773b8b9ab5aa5a6dc13b72aa8fdab9e2955136af7f3764d61b7446dbdba66b5c7d03ff62
zf8d1bc2b669f60564fd32c878d0d8323246fc584942bc9a9177656b9c33cda39a9b7b335e1e927
z0f26b0255afe5a00f33e893e215844217d288a09e3fc3154924d56c3f56cc5e76a4313d675e958
za9a599cf77c526dd85bbf3cd6d34a561f102a8c45fb8bd00aac591fb8781d013eb7c15d846b4fb
z1958f3a06f475aa1e066b4a63d29051727ebe4e6f91fd701651efaadb875b308af40c161ae068c
z7c3bffbd2f062aed0c21b0b1a1d54d666bcf940026c317d7cfb103a55cdd9fa65ff09d0ab89007
z595b795123dd574e152b567b57e5e2626836e24628df9d6d7adacb9b9d86eba4f9eaafe385eb5c
zd9dfee0bd20a097ee14541c2ddc1867c9b7d501f5a5402dc4cbc69281566fccfb816cada719e05
z4ab2987d7cf7c8f83a32e203b59abb60082e93a7e45a9a54fd6da37ef5d42b41147a49b3a53359
z21897766d979bb0586217573d40103075f1936b477e607c3f5a8866cd30b7e7848051d286d6496
zf55e1a575e3e71ca4cfa3e6e8b2e95810b9ab2bbdfba06125f13fc787d50255dbde32aa2ca9503
z23a72912f0b42df88bd38b535dd4741c1012c32a1d1ceff444cd17db005f2b52e0e4b5ff048ef0
zb99ea892bcb811781a0ecdefdf4930400f6e3e4a9204b7006af91cec3184dcca2431db0e9e33f4
zabcc061eac145d1d349ccca8ac82723dc8d3cae3cecab10125600074dcfe32cdb9fe585a623583
z4536502a2fb42ac12c339b5f9b1bc93cae1b2d0c3a8c0ae0eb781c763b8da70be4c2ba47a74f09
z1700546cb7d86220d16c129dc135899e102af4a8a06aac56550b4e1c26c2655f30c79269a57470
z840fd2aa9f53b1a32a96964cdf77b25a5a03704bb350806cf1f25af69f5aecc65cdf9ab3ac7d84
zab87ab8f39aafaacf1ed95e8d73cd9ce53d5e872e967d2a6795601cd6c17bb1f76c7399af7c2ab
ze0f360c6363561d8b1c2240e4d804e3763d7d1a7b06fc886687a9ec329aa2017f94a0ed13ce51e
zdb5c5edf825d39a45afdea92b3660cef890436f82759b023fe433703a6e9ac2a3033e92d8c9dd9
z1ad864230f937400d88b4de86d28e6ad207681a134a5e34fe91f8a110ac886c17d549a8af79080
zce39162d1f1ffff53bb5f4f2a8b0097d7c4676cd4e134bb3c30e88c16adc4c98cf4a6bb66629b2
zecdea63e8ce90bf53299a9463ad6bf44c3fc75f956295eec4b0c4c930ab3cac05d44746de1598f
zae693efc2734b52d1e97a6bff2b3570ebb22fc80566a2ec9e604a4511113191914b8e4ed94436e
z6eef0f5ac0969c4cbb9c71aeddf044b0e26a666450ba46cc1f3c5cbb684e046d82d8bc94598178
zfaf4ad2f03ded80f8556afa5609252a87e87e21bf1470ba3d95a12daeb76e6d64df9cc60e711d6
z0787190a3211a76f878863b60f644bbff00a88f2e36328bac9bc5b8a045837ef8e2a1ef141c5ac
z717e55cf6b3a7fcdfb61ddeff4f88821371bdabb1141b0e198d153c391f46f11ed798a34ff65e5
z76f008b37e1752ae5639d0f3d9e0975ecd32f1679e14e846669e3e6cf7f101676a4ee7873a75ea
z3d002156b8b38d05c3a4d7a694215a8a1f8825cb1b3b1722eed295ee0da46e706cc2d54da7efcf
zb18d2917f6afcb2256976d34b8a977106299e157dc7110e401d0f4500999c2bd6c7dd290e2b315
z4298e81aaeb59ab3d705699bd10e202a1141d9f4fb0d04aac7c21fee8eea913eb2734e1e3ff302
z249a8acc6f9084bffe03852a0736bcc50a6f93f556ec134afe9d9d118f7a45f8f2ce84085a8c1a
z3a2c0999dd6730268f9716ed73476d4aaad712803a7a0901cec8a8cc9eb82e740cbc96a8148fd4
z0b99e65cda27fefb06db42e521bd7a913df6d3a4590845b0775be5faff9d21f836c03e8222530a
z298b028b4f9d7c95f72f693fe544c80d04756c25008f9e83790a5d9c1907f4074c6b09fa67efd5
zddf536fec0793b5e3a536df3bed844def2b41f10f475550b0e9f03d0531cf42f4c6616ef16e49f
z5c92fcb709fc142a082bd378b7e882e731c907cc2e3a48a2bd3308134845d5a9853e1408efe920
z6795b6c21e0753ec7af1c948b9c834e20b30157bde5db912e86bcc03a0ebbf42b44893382fadab
z2f48bc17c7c80ad781745e4415b9e5312271bb9b29119983c26782380331c54a5eb6cb28a3f80e
z5a9ad975be7150b9bdc15e2b0094983df333712598ae72c4b6e36d0431b5c983f66232dd39c213
zfc44c0874a2b2f64832d0c3e1f46ec679b9d9192bb0f6ec391ebc83ead05358ea3badbcbb7f157
z47f5715e53172811c288351c7648b1eb58ea9098923c40c0fc944944709cfb2c8c1726c1fa8237
z854d9708e7088c79090693a51367f63bbd066b0ce4e60357d6217c47e86850c8d9a3830a3c3361
z5b953fa7899f8b62f8d68aa3a1589c5afadcb03b3562063c66d77863dc204807ebb2ca5ef0e8bb
z169918141fef0c162046e433ad2ec428c30fd144d75478655cc7530394a6bed7e43b99ede3e31a
z70dd1687528b4886b70ecc0c4490f2921a62d0c112cf6d9809a2ddd9945d31f37f91e0283f4992
z6ae431b9b94312ac9065d25587bff2a264e6a410941d7a894dfdbe01d35a6662869ae936c18457
zc1d55700171793a8c5f9eb4606843f1a0df8c5fe2bb773b40b45c5688abcb674ab1f42564b66e2
zc449c86e31ed0bd9ad1eadbb99b8f8ee1e2ed2d8d9fd2c75653144dcf5e6e308f5e4b8d9cd9132
z65ba0e552fc208fa48fab922e13b794f845937b54a73c62162357a190719c0bdb5d2faa5abf729
z465d16744be74efd6976bf1f8b646348e64e0dc20d63c19d693514a91745379d2e424fcca0503d
zcb299094aa50afbfb57642c4a548b5aea46af8ea23cc4c4c5168039dcf12a3996186c2c5ec4f8e
zcd02136d836b219726e465581e7f48f0ca62eb1b2c2ba219b8c5d937842fadc89474c9e5fc2f88
z14c6a4203ab3bd8a23a121e17be33e8e622afdee558c10524e42e9d8dc2c93a8797bbf049c5a90
z400f5c55c17e1e656e1aa713d388b2bd87669f8a22caf63ef5a987a17d82fa634d8fcd0cfc3492
zf1386976882acf88c812d4ddfbba8f8bdaaaceef1d9ecf1b18fd3a8d632a9591804f624ebeb948
z08dc0235b69e5fa4f38ef41cbf554a86e7d44f1a400073fd2a1e416193b8bda706d1bf64b5af7c
zb1042f9e02ffce6be90278356c334e24f43232bb9308bff254a8cf67cbf1618484956368d97e13
zdf04dbc93292ceebf87401660523f31da9df40fa3f6440a329f11b05eae9938702833c34682d10
zb487d9990d77c910e3f723967794ba588c2afd4a61c39331b7be00ee76115f39ba756b66012591
zf95117640ab8eb08163898c879ba79bd534ec209e6fe0ca26752201d1a2b58dcaac5419d226707
z5716b701a9986c4cba87995914a8eabad6b256a28a165fe871889a5d3351da22610e025566e7df
zdd6d066f9fd36ded65e9a9588bb768d4b9f1c96907fd553934e30bc8e5d32baeca784a1fbbcbf9
z05718a8127bd3067c1a09f112dfd2f3bf4815f9a113dcfa2517a0342fc5474011eadfaf646eb9b
z5b7783ea550e8b475b8ed925a3115e83cabe8d3d72169adae3c013c6759051baf43aa474cae0e9
zedac68e04beb0943630924566b42602e744ea0b2e06b2def1c244ab42f28b6801470e2f7d4a9f5
z133eae60e0a4f489e26a95383c14e5a7d930fc29f93a2d0ded7e1ee1b6d73cb6ba887979250bd8
z6d9516cdd7c3c89d924c8bd59d7c131939d6cf76df58d7e9912d74e8b72af47ef710a5fa9a0e59
z128d2ebdaff16d95ca3397390e4abac9d6c01ffb857a4d5a50d5bc36cfc35967deb189a3b3c3d5
z8b563bf0975fc22c6482aea09813fdb126f75b2ed575e94094b23e460bdccc0ce3d4ec5fefe207
z5e291337598be9f8e3e991a66caf78d7c665abd0105edbd73e0a71497c77d9747de4fa675c1c12
zb12af253f0709389dfe92c9c36e011a1bb7a0a2a3d8bc48edcab4745b35133e37ad9201bce66c7
z6f3f718e815204314c06d2aee96946b201de92166054d6d820959d4df97df0b5bc184f1d7f3e29
za1866766a84e8abcafcc51525f78318ce1111cdc7b1e43decf93c423143f6e5f0ad6c7c6604bfd
z96ce71b7ea3e1d34c3b3d4109676add03b2539bf8a31e99e7bf78dbad9039cf0d064ea510b1a2d
zf5c14ee212b6e2d9de9a75ede04717f9e21bb52afc984fbbe772e918928344ddfd142c1a6f3bcc
z30274993bfcb035879b7441b253c8fba656838a2f104cb5191265a0d4069f098b88a02e8ca7582
z8df76489b6ed93e25e564cd6bca2d4eb97a8a9f96397b84757dab8ca17c699bea0f081b1d9f27e
zad86b64dce8c13a1d845ddf754f649059bb310fd6ac2b9d1c98c04078d2fe8b48c990f16a88c56
zdfd1994d037776153808994724732b883e52446eefa6207a5f3b058ca1a25631c8df07fa1debde
zf97e22bedef574bc6299bbb6718b02e9d38cd26b1a8174c6829d71360106cde6a89e1fc47d8199
z784fb4241703a2f46e2b5c826b622eb41ba97d7f9eb3b6d3c4a737b5734587c10f32d91e808310
z59c8f037bc72894c40db63dbbbdf148504d8bbd9eaff4ab17070ab4d68ed9f35d525e7b93b430b
z06493794b5502e186b81f496bffa5113fde23167ca47ce9156d768dab290e99e884e7840de4cc7
z8a27e9999fedfc00f7bd7a9067c53b6218318203b3a18498802a7c81b6d6801682305f61a1dd88
zdfe6cbc5f43f39e5fce1edc34fd4605c9a3ef125760cccbbb99af82271e48858d0c54d63f2d236
z7ba20a950f3c81535bfc3123a0b63442a07b0941234e12a0435e6752325053e0c11dc0189dc003
za59951045854d574eb6974bd4022189b7733ffb901eb5d87f8bcf81b74b061683e592b473c977a
z8b30d74c778be13abed668779e4ca39f555e74f095b9cebd0375f6ae2f78951212b143363b9008
z5d4b2aa2fcbeb7476245bc5de66176ac2ceb406806e651b397d51a192a12c3fd8ace83aa00dd58
zdbb22f94b41d80173b1fadf9a5e8d90d6572447039805446965017463649e203e2efdf58b5e629
zab74fb9d7a09036ab6f7f04c9a3b825659d5791cc8c42ac091c0b7afe09d27d0237ede8e2bd186
ze74559ee71c0962ef03f4e9f1b61c6c0fd4a9aedf28bb7334cf947bd8451dc46d667290ebf5a41
z6f19fed3826a433685d9a97109b0099e8a7edb7c1a36bf8e5acb88aaa862c5cb246f97110b2694
z675375bb261b453778a339afc35baeb77a8427edd25d7b7c302c22d46de910cec6f323c6001b77
zd8d4d4522f0fd5024254d875cb9e3b64b9ee24fd17464c5ab32d8f75a2f41075cdc20ac694998f
z94029dcf377f9d705137471f088df6b13ed9c68043af0b3c46bc875cecc8759ee741f1fb48a227
z75fa2e557b4bc4c94cfda32757de8352bd76fb1b703daa4d7f159991cc9d5856816d4dd101655c
z245bf64661ae203825698008b4915ff93981ad9504b4c69cb3575a157b7a2a6abce9ffed20f427
z600f109ef38e343ec32c0ef897eed1f34364bfaf664efe2684222d4fda54750975cfa5ac34a407
z62c00dd3d24a8849477f2484f66fdb2a8a2aa36176687d90ef6cde8d14d66289ab0f19340d3198
zd0249f0d4ebbf4813d3b96a63cd14c47e7a37d5034afd772800c89fe8b4c3f08ce95d76e4fada9
z6933d7936667c1f62720404da6201349407e20df115b0e2699a0b030f84ba51a06208122892645
zd38ae220ea22688eaec2321bea04b83fefd35c495cab60aaae7293a742d7a18606a36f85b5a4f7
z97b763063aa09dc4f982972928fec4d231605500cd2462eeaa683851f729fe364815ebcde90b35
z30aea06cad4fca831e6699909429422e69669e9747addb50cacfb16d700b68f7268de0d06f638f
zccf85aef173e077f4906d89e95b6b59a8e569f751dd9c206f5e763c1f9394d7a981dfba35d6080
z644b694caa7f9a1fa01b66c05e3fb6b1b16fb068e17289f2430ae1befef4cfc3197595c409b90e
z42aebf8ab09248df02c4294048e282eac547cfcb3c8bbece1319474f22742856cf7136483db9fe
za40e5cf5911151d6ad033374dec6cb1bd9ed8cbe15ef792883d8c5ae2aa0fd211f348c5001a0ff
z23bb19ae54eaa98be8b381fb8a292ce4f6fb7d79c180e6ded0db3196d7e76c093b4e03be1903b7
z33f163603e375a9a6a9e8afcd845834b76763a9d98c069b7af4ed4741cb6d41fa6a2551357bce6
zd9698baf84768385aa9bd9bc4ef62daa1ca93cbbf993ad2ae850556cb8cdd0f956a8b26100c6fd
zecd86e73d78f76846ce1b108bb29ccbfa4f5619c113656182d758b7e17614f68bde9d7bdb8d65c
ze0bcd6ac3e300a1803bb54064dbd488cae2b97d3811ac5dc46e94d238499897e3a8b572bef2411
z108464a1c597fbe5d71b939fc4e81d4e8a9f890224eeae15ef541046f3779991b16e39d0a946ef
z7db2d7a20c7bd173f6e53653d8db58a84cc9595a9ea0d5194d53bb52147f66e7f284ec6f4d5e34
za5686096840989820e0707c8b70b572e82c681be88708132a7991ad54c0fdf9ed3c1b38d1b1e45
z98de037ca899e945a922062ca1f8bc8d999d11f427200d67c8246c4cec938c6dc2f04b4145d887
z816cc50e1199e5f7cb2333d02aa76150b0ff77332fb54f6fc814bb036319fb2e88c9486c2b3dd7
zd957952eb8f61d6c1a91c3c9ffea2a52cc580b00271f957c991d329a3aeadeb72bbb82bdcb1df3
z18805e0b168da53d61764fac9cef58b6b3464a45477d60902d66626e5f48c536358bd13c0d7634
zcff8a0ee1399a93ad3c86d86dca7fca460b7d6547d197d43ba4ffc11aa424f3ba79c1a87b6d0c9
z8ae3a64957c344333b1497eb4c44c189b60ddaadbcc15cd817e16c88d7fb83f31164450196c053
z0f568b9546e43a883947fb172d865218e63dabd0e55bec7bd07c57002d164b216e04f1beeb96fb
zac939050e3c0366cdff05df02df943cb2abeee29098912f460f5bc414a81da25a17e780731e3ce
zf379646cc60d06fcefa624be72deec1e32a2ac11dd78c2ea21acf06c1d61a99badf3f522c4d6af
z9ad04dfe8d74646bd247286e3058db950281f890accd5ac53df6a6925de94de5de8e4f3b23927d
z4a13cdf2e2348d11e1708cb13cb4beb5487459738527e0110511cbd68dfb22d0f5ff7db48148c0
ze08afc15cd9ed4d98eef12a8f0902c83cee6ceddd1406930936fe2266798a28dba309a15cc163a
zfc63fbfe97896b3d33f0bea976318c6d9ff88dacca793a4d04b2a5511ac467d4dfd1f1ae46149e
zb23cc4237cac4552f10a01fde21953f575e5bc2343a5fbfd0b26f270cc9d36ac26077e8cee08db
z564bb4ba0b0a59c29562eae0268608e02dc01e76c6b96f1ab521f3dddacda76bdf5ea1e7524d6e
zbff85e6a1f6ad35ce48f20e1cda46fde34e41713d6743ac51e063fc19e700b4fd060e1da5f8deb
z91af2b6f893c4b7595740185886d4ff369a88a29f483db0220cffc63ede5ec5cb684639d342054
zdbf61344197b77cdaafc266e8582759ff3f0ceec6a806b2764392550cfc72f94bf77d6c3356405
z9d81dda1057295479d90a9e398461d1674694aa50f9f7ba98e6ae409edd56aadd3d07823eb2be7
z394f9dc5a624ccb15a17073a1c26cddfc5b80d442bc37a44fbc4997ffe52bd28d08357090bc554
zb1fa6a1ec99dda23ad65827c4190ff43cd0f3f8a3992d9944177ee918c9ec7b31bc99673b13f79
z970331dcfbcf8a5a7b1523771961d8418ad368f0195e0478dd5eb477ef027cb01de91e86c7c0c7
z059c986a989b305d0f35ee53efd5fa351ecdde30468cbe633f45a2f687f4680f50904d02a4a699
zfaae7c802120717090fdce74d87b33cc80ee58a85a2a3b2d1126c33d2a6d897c72ff2e9340808b
za895103caf46c96ae1fb177bf94213860f4fe0649aff5d4b825220bc520fa64c4164741e915633
z1cbad830087e9434bba2a90c9f35205984ce501a057c28d835a7158a33dc079132d987da22985d
z41613babccd89801ddd768b92e3ee8ac1440b982c2372006f06997d1e66c3d48a46ca8e8b9485e
z9a9d5cf43a0db6b62bee29b77009bdd4a7c0117f3a711af70e7e02e5c69a9c7f57d38ad9c1cb73
zce82072fc8b6821cfe4283d286c8a7107734c20e0a77801d00c2aab70b559c5b932099b7b445cd
z611bd9feb24cd62a1f5d7a3cfbcdd9b497e6c7bc3f722e1de0b33a878576c874a1b58379d3da21
zd52e3841653e5566722c42e94ff409c24db463f341348306d6e10d98cf938b4a2abfd07ab849f3
z923531108e2df638e88bf8ef8eec237cb3d4f0d3eb898599bba11c28636f7b5cbfd95da35c098c
z5484975f9a1faf3e0ea51f9c5841443696d1fa2102132653a70de3d3b623c41d5116e08352a1e6
z1a198ad6fc74139a64a02447a894e0129b9de705d8132004341edbff1b8512fc4855535375a9b6
zec1b034a00a62b4ae5f593ea71451cfafe8783755cebc8096a2e20f1a88c2443c4b39372e94ed6
z3a60e78cda07a8f3623c4389cadd753195aa6d2420304a6e622d71467a07b7e57343468df72966
zca743aac799b24d7476947a92ea248396e7d93aa7acc87b38daef46cbaa26333fa69ed51545cb8
z71ee2bd32cb90fd89dc54b0dd1b91788bb3f8906c90c1aea0c35b96b562131a133f3779fa34dbe
z25031796e8a000ba556c3cfe09493a47909b42ca9ce0e1af56702f92e13e876443f4de44b6814a
zd3167aa1b3448c8238474aacb057276ba4272c451c3b1992a2d58b13d449927c2e02a55eb72544
z68bd0ce03bfc9717a8b5c95ccd6d208a2cbabcaf31c0afb0fa134b40c1bced188d2ab584070537
z4ca84615e0104422b06a28b2e429ad186b35693d86f3093ef873664d43c3cbcb46a68b685354d2
za8757b4bb65b85b10b84c0c743e76f578dbf9d2cef92c356fcf27e0acaf0caa711ad7801c7dae9
zff4745c053f8407ffe2b5632be0917cb044181edff18282c4a71cb3be20167a44de76b64823252
za028d9985954677b340eec60e2dadc6dde1bd9a537e37f5f20a7f992d75a903e490c5a76b803d0
zcbee1458ddbad05e9c56e816f26acca9ce9481045f61b1dd73cd9452dab26ae1206b6bc73a7da0
z9b03e0e9f3255e93f88e0f90e3b9143c1be26501d67601ff5b9c626738949e3f2b7dee43be21e8
z6730b4b23f55b041ee5ce5a2a27cba03ee18dd6d517fcff46d981073b34fa08e67cdb6cd2ef4b3
z8deec8a0e5151d93495087b32f60368c0e4a5c13429ae559edf59efd8b9b6ed5dffd97d3adb418
z5a180da53508ac9abd0363786af292716a43a2170af11552bd516c2b74127adfc276188a9b8c32
zcdfd3ef396c3b0269543633ed0b9bb010e702d9c72b0675b2a43ab412b381b999423b7a647c5af
z9fb71d97753e7010bbafb0db411babd8de0fe15f8307918b13742529f03652a057d90d22a2fa38
z7b2fc880882554c90acd443a0c534c13b04a1622f4562bb3d9bb6d068172af06073a01387160da
zc56615c7d4d24fd76769a80a8ab2af97721ba902f37406354a2de5f027bd7850fc98c029eef532
z329c404830aaca84f30c44967745cb052eda7401f8ad0399f83c4b3002fdcd7f19df5747e1927d
z5f23ac0aa1adda7928d57be081fd4feefee659ce2c55d7761a07286ce7b2c82b2cebe03ffa5963
zbd30e3ab9fc67abad67578bd1f3b545ef946f945ceae51c84a5d34e29d98be0061b69088cc5ffe
z3d48414c9a55bcbf2d8f44a3c6ed6301b706781fbc9063956f47f978d6e7f65488dde30f66e5a6
z79ef7f561859841a73134d9065f62da40e5fa2b58b9bcb58c4659d72c688384cb8c8f1633ef4dd
z3205d2597506140397d50e5aaa2412254d2ab7af67d79b3457048880660f09aff528318e4b2a9d
za0bea55f3fb4ecfe68ec078b97840e7583d3663c49e542211e9906736e6abdd1ace2acfeeeaada
zad534d4762e010f88ee779ca590dbb0f53854a0af7c33cd4b36c9c495331de04144383fd7b3db0
z3bcfe23f0e5563c09a6f45173a1a567ee639013a4d39fc6190685ea0dbe677b91d8c4ced99a776
zb23c4d9f08165764f8e9d998a0f6f25702ab3e47e43bc88c021775e1a22f8453728c5ac34eb234
z024b0d21f20375aba138e9b7427226085702f109e722769c79819639bf03ec56e189f3fa00c4f4
z7cbe8e0980c548412e9b498634d2402b9c0f01e658cacccfb9310930eb5ea669ade96b6efba55b
zc082bf704a7bb73bdee940b002e367031e850a60d94d02d298e73dfbcf522d05f4e67bececdd3e
z8d0f8e514f177b231996cf2973e437c47645e59b8c9f71eacf8e6cb47b45247f3ba2a7b0bb5c7a
zcaf66ab78d9edd7df50a379b352abdec3c6caa65468a9b111abdbf7b12d65defa900ca49d956d3
z8cfaf7fa2ed815fd32786d4817e5ba0019750203dbe38613db4d4ac214a3040674668b59585f7a
z630eab2f591ec750715b172300b55bf3f60ce21748963cb196ac7d347f52b490740649855c7b61
z14a06c6b7fe590d3950e48dc80ac1fdfa2bbf07f46d2b0f3033a089dc91607216e9eae4df44c5b
z1025a0c91985f22551ba8caf034ace717eff88e7a1e843e844f297fde352f3e67f4741eddeefac
zdb06dc1c41251dd757cd291b0cf5c1c672383598da20e02ecae1b5c14f796221f2fdf675470d1b
zc5fdfd7f29e29fb98a6f20bbbd32b830b39d299f0936bd350ccd079c47649f99d80a398da5952b
z7fa1d7b90cea0c025ee6863bcf0d347e23ad446a92e1c3d46538a2697fc84708e041277e373ee5
z7c39c800db4adec56568692ba7fa6c0b66a0cd74f7a67f3c3e2cf720566960d91a291cc9e0e3d9
z29b8ebefeb9c9988fe83ed8e95d53920bebb20cf43b3bbe4760e2789392ba32f052b59fa58c851
z100c47a9abf4e4ba67b7c238d5c187744bb4912d1576d032c7e80e21b250dc48594312e56e9de0
zfb5b180de994a14ad0861951240b81ea70a856d574b13ae74d486d16372704e062f98cf194c94b
ze2465ed4b827919c7dfec287411d23636de29332b4595d0a8932b5a75c79598b7747a647c7b73d
ze2c0cd64d820dda3aacb40fad5ce977e33dcb07c04e1b09686f63693e755178a77b263f1779e7e
zcb8bee8b1c8b549a15cba464740e758ec0c58cd92270b10f857380e88990c22ade0713faa5a55e
zdd3d3928fd3ed07a25d87b3a130760f31384a4448cea8d9ad65431a82f7a07608508fdaa28b840
zc4d9195cca3c6b7152c6594a17aa7c1fd622d3a903609cf7b4f6c9bfae7d72c7039e7f08540eee
zfee03e7d88496f633e9be2e3f14c8fbe029b7a8ea658ad608c5b8379d9917ecd4a981404b206de
zff1b046072efbcb6f9fe2fa7e6c1dbf0c1dbe8c10ce5d6961f5151b6d9016f22b901142cb3c99e
z3fa4759077bfc42d2648612a13a376d3885027350b546f95878ca706a17cfc55b51d76a3408f69
z0f365920840c9a109b3384434ca86912d9ce1d774655fa58d043e6f20c19fa572850a76e6cb79e
zfeccfacf6a1ea9783df6f2f157aa88022aed7494b3071b79d419405617f8b9a186705c5d2add2e
zb0ec9de2c2d198ff6134ae3c52adb5394eb061c83ce2cfb106d91ec60a9794f56ea7b5bbabb411
zdf408fe35a06bf8d7cdfd5c8c2d1c65b35f193fce584a98e0c7b7e1cb295ec6b1f461f4c1fbf72
zb127104d4aeeb722ff7282115ba0bd5f63496350817fc399ab05a1f02d3e8bd55239f6618eaf44
z1bbd0885109ad10985b47a494d16ec980d3454a5cd41c45dfa33b2a314c56e2290de375750c98b
z569ca0ffa214982cf125b441c5ea674c84869da02f359cc015c126073b62a6b7307fd447ea60d8
z01fa1e2aa22b69fedcbf8cf6403d64674932f5d498f028b4918d31991b6d1524e51efe2707b5e2
z412a4d210de1da27f9907cff41056190089a44bc687fb63bcaf921951ba24f09ad7aa9a4c1634b
z3624aefa8d4745ee0043a14a8bcf3d75276f1f45c82f38ad10df987fe21a2a7077cc87da3f1f24
z47f5cf6a2caaa631339c877c35d5cad1a5a75918396aff9dc2e88e5e368bc40a7673ade00a8db3
zeff9f09e223b58b978452591be8188e1cfc0f6b627233b10b137e5c321d2df3be2914614432b07
z3c215ad30edb0b3eae8bb44c6acc974e1b4d8178e1492d36c6a17546ce820ae660c355fe379eb3
z108f4041f9f8d8acf452bfb6aef3d4af6cf57bd2a3d67502472c79ad178843893adb385670f4ca
zc5df38b96afa669424b79fe0f32f3ff72e19059ff712fb3309be05c1516a6be0251b7e7b7dd56d
ze897dda9f1db54159cecdf4b5d8eea23175d46563140012b15df80b69d62d43f8a5ee58cb4cbab
zb33db1e9b70142c465ea4fe2d0e36f1d028eca1c738477c5031fa39911d0ddef0495888c7312ac
z0d5fd54d9df3d517d3a22f69dce3b35ab85135a84faa49bab7b3fd488d34eb1c937c150a766b46
z327b470909a32cf249364287367a5ef3ba49c0253e8d2fbfa6d94869062e71e604d59260c1bc6f
zbd8d8bb3de24e0fbf97877befa41a799b27d887fe46f549412b2f9e8b2721410d346c06286da15
z27e19f4cfda6e5aa2010cb87f7294b840ca6ec792432d87fc582b3da60f112235118ff10e34c14
z1b8e360e2530ed7208e35c2fa28c1bf514214fff9b32acf4b3ed0678982b3829e8173f56bf4ad7
z91ba464c2360a4dbe78156aa9b17f4c15ad8fc776c9d2fe7641ac74e58cccba9e5debe9c735d28
z9c5cf7b81946d3fc5311d3412ab90d1c8172f989438d183482cc9360eac183b50b090a5f8eb6f6
zcfcf9c20460e421e29b8f0025056698da31133f91d0e6f15fa6ffc811b8e56a577a7a6531db71e
z782e351efffc3bbc9de5bca86b4566376ce2256ea43fcbe125f465f71f20131adef0c14ae3b6b7
z266585e894a8e46e726d619791a4f95392e9127e740059c1ec977fcd8794307aadb50d6e504336
ze6413fee24d73fb48a47de6983c691c119a33379d70d3bff7324ef6405e087db96cfcda5271767
z44bf7ce8e2651ba581e02bf6f00b01be369441c7005bf9b2632e30bcb99e2d0c1ad6ce0cc96522
z05c48da64b5d0501de31086727af998a7274e539be35931e20b2f53bc03e71bd76f466e9aa5736
z26463055009104ec89536fb3a30dbcb4d157b95572d9fd4329cfcb64150c79c514c567b4360a47
z658670426bcc11f05ceeb6176634f96ba4f94191815673f0735c633f9f23908d661cee93752dab
z0288e6ddb8f980fa61562ca44b396f8bdef18ead802d170da049ae56f9e18ffb5d5588a742c31e
z734855c2d4a1406abf16f3295409a4792d3633e4ccaca49c014e741a416758d51a648e05c41169
z2030840be155d5cf9307aa2c2a279f11993365a597048f103cc89e059d091a249fd74930701a02
zd5bd53c5fbd6e417961aa40eabe378c29702ac9d72403475049bacc05c99932a5db81e93bf089a
z3037aaf737493434fa46233b32af2036c1e13406aa7070ae1300ac7cf21061ef4b5ff54b988ca7
z22101b1b934a208ab18c2a9eb56217ce9624559cd5517b32dba615c570db0c922506bb9f077486
z63f041adcb2d71f65ebaf5a3155eacc4b4590c865c7980735a8f96f6ca489bd9d5932d259584c0
z5fe48a1f140c943e2992febe12fe343068e4f53ef88d48733d58fc1401ce62e037edc2610a2719
zdaa248a0ca66b9a0c26a4a52d927dd3c6568c412900cf790ea7fe2f8669fd5773f8f217831734a
z85dacf6f44b11d565cb10c8fc559f11146e4590ae39e8125690781a96e4c383f3d8a52ee769cbd
zcc2f032a1a19f9faf0bff7cb32e03d7c04550bb5cd946a3b3ab551b9456b51522e4b6febf0365e
zad404183be92ff4af81bba0317c4abd9792218214ecfcd54e1759bbb3c1277e2e563388727a831
z5fd1b6a1a7aaa678ebc518f468f0275ecf0844cc01bed1a5b2733bc02d29ad8169469cc43d3664
z47ea68b255d85078d7ad14e8476ea9c3780f2fb39eddcd8cd3f8521ae260cf915b24ff52c00aac
z5c021775b4d38f85eb0d188c643a3e1fc35902acac833362db81691b5e972ab1141a02a9aeffdc
z580f0151a18d6f34de4e8f81e809a1a56fed4be9a941eb611c21de4796c67c975f638746763730
z8c0bc8563c76f31f7b7522c889ac0403ddf628188f064bd2d7180b07857698f2ae055733c1fd55
z6fbac720db76f3feb2fc6eaf827fadaa51c5cd49330d0e4f0d2f27e5390b17fa3d26e54153b65d
zb3fa88411d73ad0dabb82c31e16ad0223d72e5f3f8bd0b97f78739ca6d2ba1a5c506f8eaee9b64
z86562789d2e8370646995a6af430c606b5be4c92e8e559ca2d93c7b82f3fb558959c396762a071
z6f918d2a67772f1751ce4296bc9921dc58c55976ba21c88e1bc05fd6bd4dac83d7107cc6d08bb0
za7780809d306422674a1a61b672085e2ef7ea2c7121b51f47d6321f1c2d9b96b506dbd89e4bddb
z35167808fd428d08d6b388f3ee06c82dcc4f675c68b8da49558c1e3600197030d064ff93d9807f
z23ecfa42a648f01933db25ab3a39a9369a133daa46a413ccb11192749a455613ae51bdabec4d51
z871fc8311b521dd0e59f4320be42b6f1ddf6b0e81ae1686301d7bd6cdb5b11d34106d7c7f5c040
zce32f743c7f32f5ffc39101d139ed657962bae90383b5674cb3b543996fba759d146f37bd1d54c
z2def22d2f40326903317289a53da61c9cb11b9d0a4dd1c700de43823bd76e01687c801236c6997
z87585c7b1c69382bc7d31ff65b78ee0588844d3b12f572db98a268796f56f5aa99e7eba199c857
zff03398568f4588f82684661131b6d2e19d56008f587001394be287764a1e572d0b06426edae5c
z1de5b1892b2b5121cb41d7f79e1fc92b2639b1880f96400c1c4512a09e8bdc1327b0593a31e666
z581a66c70b6bbf611c33709831ab436b8d625fa4ac73ab85feae2663e39baad949b24f5af47970
z54931253865548f31a255b5c2ab9c5a91027e9d9d30c7d450e02d1b5a4a70fe0a4d6b02de5e526
z9714cf167107b80dceca2f2a3d338f699bd806479d98fd43c353a43222511346815330cf34586b
za982dc7f70d90f3477ca6b70833974f5eaa7c9014c4c2e502dfeee05e35a28bab09fd4755e8e8f
zac557e786641f778a5443e6c304a450d3fdcf9c8647eb24ec679112815d264e3920d55df801437
za19d623f55ce08ddff5a975d8e2b4a1d635a340bff3ddee01fe0a93cac31cd3473cfd5df3e934e
z2abbb791e5f33a5f186cdb1301714b9ed37e95eea7d792bd7dacdaf513f0322cd4814ed5388789
zb29a926f80306aa4d54e7f00de980a30eeae48a87d563fd42e96f3b1816f5f831bca2a8fdafc7e
z9562622f94904e0734385c499b7a6d3657971a7dc8effa4101304a43444b3c8cf85a90fcaeddcd
z5e2033286f915c0d1c07f8d3d8cf830bc8c3787f5ae1bab70991aa82fcdbfa07a5560a7575c907
z5a50e62a82c47bec0b294385f1280ac77ab2a6fc1e7b202d8ad079551064a5f46e7ebf433e4cf3
z731df0c2a04c5243b9a36d30746e924c9e1095e00c2bc1e0760b718ac3427ec2541bd796898026
zd83cbb5b07d162654f64fd114e4899ca58c1a482d8b19c4d1d3e6ba4acb686db03e7f4f9485320
za303aa0d8013d07a008a38ece4012c2a5b7d6eda31e5c7c0bf62832fa310e14cfd681a5d24e800
z3135049a5654161546655e8aa3b99932fecdb8ee10bc7d0d44ccf36c27aa6e7e91f7a9bff6e73d
za0138924969821da7444fb84827b64d1a9802667b11ca7bf36f6769f7c6764af9db2b2b1cac67e
zd17ef18e2dd85504fabe43e98a16adbe09cf03d8ec4014ed4ae77004f4cd0409bdf5dd16958f1d
z3d7f4273b33ae1fb2e9b87f4c37b2e64ef817a0452e41d9dce2818bd2c8ec34399c03b2b4aa823
z14f320500096230deb3a6b7989dc1265b507f975a616013880928046ab54ec1a1a3d244fdb39fc
ze12d1e8d2752d47329f20ca3925318d04a4f787389641193b1c7bbc36d0642f6b01096fd8aa66f
zfc7964e19fa31e54de268d6dd28f4b705f6ea9696ea4648e15ef1025d176fee18a4cee01b1bc17
zb2250f8c3a94001ed05735f1c182eae489cf8cb3b2972eec66413ec18db4e7cea009e5e893aabd
z526362dd511784c8dc2577670ca969cbb0c010bdfdbd16c452cf4e9068573836364b1b78d0480e
z0fb414efd981616a05d3f034afba5f1a4576be293ff9e224b3a15a316ba4089969dc940bac7353
zceca306d0c1b4e0b07167c94fc7614bbee4ac60d7b2374f71cd96ef2f82804dbab1426d0546378
zfdc72e2ad2c678412826244d5f8d09e3bf50eebba5538dbbb131c47b322dc0611446fada80ba43
z822ae3a9917d09b8b74ab8bfcdc662b138f762e680f1ff4fb8550cc03b94e1bbef37931e15d589
z6c2f1af80ef23c535a9ae50145401eeb090654b8aaf1346adad8cf5eea910b45910878b14be1be
z1b7873a8e7c1d761254d6f67b8959abdfdbb120dccb956b7566fc577d96ada5f5661efcc6e40e7
zd46c492c757d24b04fd415c1442ba6fba841cc4893e1f1c84e3a7db9d0b3c010ceb868883d4db7
z9375db93830b200f9821c37d84079570e1aa39b760530b219faed3f018f82ffb3faa1e3f4ffc1d
z90b2341c342cfa8968e514dfdbf416864c5beea27cfc0b6241dfc4bed07f116d2b486e40d0b3fd
zf772b89fe463d7a6ea2649b89687337e67d0e9370cb54f9dd148fd9ef28c5d9a76b2a25773e146
zefa20c5cc89bd46bdeb7522eea0137244d1c3b032a5322515c5d4168113e236188d9d0985e8b6c
z3bd0a2fcc1dd0a22961593db35d94c7804c32f5274862bfe81ec5ab876c4e7d9ccfac2e0624985
z40a62f057b05cf51fabd81861f21df3e128471e75e77cd9450467ca1d46d691ad8a8172e5e635f
z339ac76c05cf16e898b3b10fb6fe2ec669e31ec7b0e981268736c564d662cd41fc978cee7cddf2
z81ebecf6bcfc4422a75a783a5d78bdf638dc3c8d53e0b7e00ea3f8f12eab16a5c44a5f0b363fe7
z476a18e14ad32d8b7ee3a69674eef67a81eb792244240194f066ef0686eee1b1776f8efa8866a7
z31777418b6f2a4f86337cdfd513eafaab9f8daa38902f4d554dcf75d263d77d77317a380568f26
z60031ec1364fb8199396de255ffd7569cbb46169fb4c78b7b5734ef69f6ce6f17698d7da0e7e1e
zea6699a0f1c59fd50d2275ceb578e8d3389592034abc701aa36edf47b99d8abc13215d2015d8fd
z01c0db436cab655c6ca90dc48fb2e0d99081b2d1ebe2bf0417dd827f7b6f02fa569439a881b9fe
zd7be3388c5c2a04b42d1fc84a03f80fc3c69b2d0a75a2fdb525766906847bf4a76fd4bab30f31a
z76ee3f34cddf0125f706324403c96dae26e94e9e44c22d6061bc44c4e3ca09f0b60708b6e08cff
z8f27204bf6e045b7d27fa514b7b1190ba4ed8de0eb3612962650f02713f976ea213197be64ac37
za213b54a65b5930ecf6d833c37204c3c3dff5aafe2b998bdbf6e8ae5300b5aadec3350bdc68f6d
z146241bc9422e50fe030b90193c85e6b9f02bf54aa83f28371fcd3a96429c8a8ee991ccee7c798
z6da2c0ee464721c7ec0f3754e235a91d64c1606d245283b64d7eb0d0ab876ae95b9da39c27ec84
z32027af494d70345f9c83e239e858ae2017ed642304124140eb8719fe9da3d86823bb21769e74d
z659a5f40e0ed9bd78ed8db906922970422fbe8f5ccabbccf96c8273b8e4b5a63ab585261541008
z925854efe58a4602fd4a20d30d944f1a193651e565ec2548bb654b10278e0a3b6a5303230b1dec
zd50bb73bee924d3e2b3b0f8f3bb525d7e06c882990fecf7c6af1c97a352675320f312c9a45bcd7
zc24d53c5c3a21598971407397a256a7fce524d22a9fb80371b1f0057c7de98bf9cc37cf163612f
z9d83eef384a2aba9d915f7dfd0343976d2c3e57fff2f3bc9527bc8359589b91fea8774eebe9023
z966595cdd27efc9face16d7a32a228c33c2ab5702e4e50b26d093e65878086ca4de8ab148d09bc
z0bca49b991ee805274ae3e28748953f0cf2bed07a3aa2b11be45003d73c7db0debf9733d72f429
z4f59ad27c323dda7239dfc70c74c8d2de40e2a4303e64eaee748d02921dbe4071880701eb8c635
zf65de0a21bbabf1f83c5172042029626ae4996fa002e222f2efeaaee66f852c54098ba2581f10c
z8394fe71df70f65c2f35e8a676e94e23125bfdb6caf244ce60f13e1dec39171921e317a7d81f51
za1f76f33bf3b866fa88666a0a2d76183abb31787964c92e93bcdbd436113fbab5c1a0ba5ff6af4
z64e35c2169976b00aa982f92564afadbc56893234e25b54ced2eb25cddb953ef61ed12f96f5192
z3a8db325184e840d86d806cbad278c8769bb7b8b83a8b5c81b4428b8750b752b903f9eeeecf5d1
za991633b6b27c83988df8f65242c933af422d800d693e109f87a3ed02be7668c73eabe90783f35
zde11803f5d1d0d16c5d7571f0b29ce17bca62cb44db7f43b0579d0335d4b63feaeffa78cf0080c
zc4d5face61cc9a06a8546845c3918fbaa47be1e3e761d7fb55d691b5a3bb4f6ee7691dd32475da
z2e191e01f1a5c236cbe42d2d44fc257c2b3967c726cbbf08e3a619cc10a154379f2f3f0a0cafdb
ze00fc68b4c08ef5132138d8efbc9140cd485eddd54780d3f7902fa05e5062f1096980482dc8dfa
zd3f6d4cdf7522705f15bf09e8ab35ad7892295f558ec63d747eb16b1840affab622dacfbfef47b
z78b040a1ce93992a467351fcb90f092061d49ea94d2a20cc896e49fe06d0d8f1c6e006b48479cf
z40af8d1d60540762baa45570f2a397743ab202839e10f86461813aaeb4e14b5a7028badb44c80f
zbfd1ffab0fd2f79f40e577288737cd0d053a7a167ea0b4c431aa3c681b1eab459467eb6941c603
z26e8b5449f707c61028cfa5b79fb7db3cd52154eea731f1eb2541fa9107183963b19577304a467
z0f99b91e9066ce6ac3e34d436011280b395c40c9479e54a588dc961a36d48081f5350e80e242b3
z9c270ac032408d1f980fe7fa8c6b8f22fd2746ee69d998bc43f39c22e96e187e85c707949be6f9
z638fa6adec7f6a81208cd5f86cf0722c201451ee991bcd175312e388711c57b5ca150321006bc0
z575ffe13bb3def28de1d65b6f1c00a6a5f6bf8f26f1c026d8381eed2eadbbec0c0e03d5f62e8d3
za6df654429f7d70684adcdb5bbfd61d5c614ca85cdaf6d803e35ea6de59d550d4ee36d83bdade8
z07636d1d4cb95607233152e3ed97ace05ca2ac1b3e7a24de47908e747c7a34f1b77f84805b678e
zee73b5876d1803d187744e14ac25a13bb2dda712010c9dbf96c4c3b8384145a664923e60e320cb
zf947c89cfb02c2ca6fe3ec8412bad9496fc5f45c70344d3462adfe15f15d78c9371bd99137b90b
z6c8180b4e490900d74884bfc6488326cd71102851092749522be5450cf22727904832f1e3678f8
z2510646cf4a151a9f32172d0301c6ebd48383d3b7aebcba0393b2f0d23f1d9f4068e471ba75509
zd261327de28b8e77fc3030bc1a6b78c3934b51ad8b7dc786d50e183ed8f527163cb0962357ecf5
z177f0180e1a404c2a305e45ccfded248e58153838505c7ca16d673e8b05a05d88e7873a092e9f6
zb8051acee164399516b9c2d5a65c61301d3826f67db5ba5da25381ef9ab0586f8c27c7fbe23ea9
z492f81fcbeabc0a09bd54798a03acd446055f33bf8cff7be8733b1c431abbee88dc9eed965aadf
z6a691fc90df60e4e6b07723a61c689e03fb5d75bab4d5b860d47a8a1edc26804e5a12d463e9d23
zabfc2a85ee7666732b43079f2699b61e8369597eaaad3a49cb19ed1691494dc68ab90ac750092f
zc21c2f39358229e6184dba5a03135eab997c18565bd0b5cfdfcbb58f8f918297d7e85e6721dd25
z678d6de827e284958445867adf55d50681cc81f3f896b4a720cb1911678c02b9d843c752f10cb1
z550dfb8ffe8d25a0787a3a60e82b6e6c29bfed10c2d5add28e41014b255aecfa6218d515e056cd
z55f42e4b3f9235cba6d118bf44900ca1eec343c4b6800247397fd8dba19aa709bf8ee3444400ed
z3a6d3a995e3d290465cdcba9714d834848601b4c8ae081aca754306e1aa5d516b454b70c198421
z4f6e9f3396eaba4bfc88b12f627f32f49a50940526fdd1d8791f0bde031f103e68ffe11e7df3d9
z214c6c1f2419c46a7864d1bb82d103544497bdd7d2a44bcb5fe711220371699f3093b1d6497f55
zb424d04418aba5a7c56382ac9d94e2cacf01f593c8c086ca8d6ddf4091fd87288a85ba3db04fd6
z0c54da3e57e0c0bf5b6a3356422ba8c1f5df3f9f2a2e83a6e7d2455c64f9ebf43c2fcb76717ffc
z6ead2e7fc847c39033151e72b493a3fec2ae0ce3c825f484498d2bbf8e97139389389b2c01dcde
zcd9e20788e8e3bcba9b4bae45cbf58e653fe2506bef97bbebac5b03cf01cf88cd42b0f71817f37
z99dbe715844f727238c82159922cfc396d8f287b6545db3b2d8cdc333be639170c4a7709eef01a
z811baa22d42158e1e1b11b1327a428d00a35d78e7c4645ee7d24d3b3c9bc33b83ebfe83f288e7c
zbbaade2f6d8c2913f0b173088788fa49ce45139f180c2ce2d9514d831f96b11f0a2bc425cf3c63
zf0cf46e57782ebc63fc17a27bb9cd547e58035d9b6b03c588fdf8e4e75cc9ba2ab69fab702b453
zfaa256686377af3e8ba1647793066d80077877076a89ff5abe7c06e43a2e16345be73220f125cc
zdb9710d55bf4aaa8113ec92974ebaf558cebe563904bdafdd46146fab3360bc7d9d99211d59376
z08bf3a263e14941ef99ca1e6cc36fc46216e4a54028adb5200c0b80150cec8391969a228926829
z79d64b2b86e463442cc90c0c4bb41a3528ea1cf10dabb093cf595cffc76f9cb4512cfd4445a0ee
z2f99c4627fca50acf16584bdb500a4b0d40a26e775b29d0bdcd900940189ebfb12bc576cf881c9
z4dcb93f06f86001f38631454170b5b6cd317faa568dc1a9a94e8a95868355e83578814eec8c86f
z41ba3e4c81b292e94956e9fdc3b074981679f39d86f069fe252736ae084052d97c79f627f81f47
z48c96d6b898893e4fcfa5f8e2fe9c5f9011c211448d4209f58a693dc7d734fb700ceebb3d0ef36
z13c0e38e043ae6e0ac19815cdc2e68c2af9658286747a21ae50a2274bc35fb4b356f346b81a599
z5d33b57fe88195b3f0a51975515c06763fb06f804fde03878eec4879782171b7edb90375d648a3
z94e0407ec86ddf868907080564bacea2dea5e05f8f386af062d9cb1e504efff88981b848ddf6ab
zc400dff978897b69c5dc935f14e451453018b672e4a6ea86dbaddfa252bc06339457383cceeb57
zc9560904f59340d916f2e4d970a57a0c70079b9439b4b194e761e49a3da5dc4f3af4bddfc9c34f
zbe29f92b6e79663c954fe235874594f4d068930cc885d39a8a60c72af444e829c844b629130ee4
zcff61a7eda083106003031e41f4f346a39c390cb65cc45135ee342c86cdf7529b11b2d2576ccba
z16c15ec4d76387179fbda73909e923b83abad6997b905f762d2435befd1ddf3c7223da6fbae340
z27f79a8a9087c1df0f38da0f70efac4db77c25fff73226654a512fd95111fa77df53556c2a33ab
zb5488d8d4be7e8d3a41985e7c169887be2555a4ad3688f2fe7ab9c58f60835a7a75d4f4e04eac1
zf789e89fcf8695cc5f2d722a5611cf342d08bb9b63e655188e66215e508ac6264d38771cf74532
zb787e3423342ba66a9ab988e3873a748ec4b55610bdf0992589719463d4b563deefb5af243c8aa
z39cc9f94084976f5155edda73966c96be542bcf6b1f9ad0781cce2d0f527d9db73d9fd137b0efa
z8f4c4deb7855781a346e1ae13868c2bf6504f645a4f9fc39ee861d6e791a91712b0fd246d3e223
z365bed2362c1716ea6b24e8adcdf368c7c6cc4f66f4cfba5d8d9635709c074383a3de94baf5288
z83811817e815fca12a73e8299a52407d32b8105ff7a23eb18cecbc8595567a58effe9f9d745f6f
ze0df7ba773037d7827ded9428eb1786b0b950d1d3c78f97134a6e07dc2d09e37ca1a72f3856e81
zb106cd07af3cc7cd16b3acfe5ab1f3ed905ae1f561958ad72f02f156d491ec708ad38a6389e493
z73a18e43c5ecb8449904c49fbb1ea65de34e6e01509d67c9267b17f771d6f575ac16e658ff9b8c
z58f4faf7e4b8f8aaf934ec11a9d63e85f595ae4ec7199b9f57e276aab699f651dc57d00808c8c0
z60bc8a3953a27a7751a2759163cfa6c4ca1893a20918c54f6099375d6177200b697f2d2939cc77
z9d7c93b6e3eec784d342c7bb8b7ac3b8d853dd222df58acdd5b0d4d10e74266953e3c09745f3bc
z4af32b5c621d57f8f0921b0a423cd24ce3641c474bb72865f78417ce526e7266d679ffdbd908d2
z002489754a7c720c10beae995a51200cc051eee35f1e5bc22d6a9b5fb1bb2cdf167b6a7265ea59
zebf77539336b364187a090faa9cbd6921aeb1b48e05864c65b1e64b8e0428fdf3eaaa4fee3e81b
z5d9e9586d0580d44e9c94fe697d4f1edc7eeb30d8f14e76f2803963a71ca889c49817b1cdf805b
z94f995dd2088195eed9986ed73f6185df60689f91ac3c34e335da9d220f7de049dfe3e240247a0
zed3d642fef3a307d94a3d0f0f49d069b657a395a0f26b57f5b6dfe875ca8dbc57702c340b4105f
z75227a67c6f86126c4d29761a223d8d49c513afb28d1e074954d3a8650411d3117532d6582dc71
za92db715a60d5ef9f8dcad73f64e3d040201494209de381df68b3adb300374fb86d18bcd6f2707
za5e5aa46ac05fb39003d564e34e2ddf08df7e1cfe58384d388d324e4d0ac973c1b4f492bb15f23
zd318981e051ce43a8fd47480ccd4c2c5da46f83eeba5fb54764b323eccd72816f7c7dca2526beb
z77f7204f48e9262c895db567ab8d1ecc5bbd9929718cc80aace48bdf318cb26df882d7497cd21a
zd8e960955de05d03cd0d33670106b75565fd82a8095b559c74e9d6d47416227e11e5d57acfdfd7
z6134b7c9bc8dc8ce71fda24c7852b71968b5ab585567ceeb688f61f80b311ef153cf454ff764ae
z42a199dbfdb80e14733aff28b6a85a514ba0e957b5eaca3134c35db1f78bd146f3dec40a4bf586
zdd4053ba504156f65b49406d499f8dd020ddafb1dad78320e1a4f3f2c7f98d7cef8e4144284179
z3c88adea808551f8b43337b1db6516101258c8c90597dcd0a725961fb1a13298710830f5ab5229
zdc2c5a5b464d31fd5dee7f4d4dba01e2697050b42750558acfe272d368134bbd2f0b15b53210f9
z5d6bb573285601fabee5238056a86deab122d37b20d5fcb2dc23b6cea9916e801c9d021b4a31ff
zca531e71c9a60f3f1097c53eb96a53ec9596f4f2b0abc1a96d405e29deea7530c2a5b3ff54de04
ze711a0ea0f713f8d5958552696a9a424bddd10acbfb7a4602a3d1fa48a1f5df37368d1a8316f17
z95fa218a4c5ae303f644b4153a66892451e6b394c4295e3a8188ff7672e79e9913dd65ac91cc8c
zeb3ed7a9437ef6c7b5f972db4588eb7c02042247a06c49b20859d580f74cb59fe00e447f00a421
z175439fbaaf0552630e0502802c5da7a7a10999d561126a62e81d1fdb39d7987b4e174b047feb1
z18f7478288c70c35a6061ee46cd3bb93d7cb558bcb8790043be92268f5f50b5781063b6fa8dcae
zbb010e87cb24103aa2b53ca83a217c5096ee94f0fce002d70faf7a8ce8c8dbb952f384b17e50aa
z7a409e3ec1a307400ae95ef35f8c38774a4001ca4497cfa908c9dce723dd35c4f274931aa570bd
z41b8a854354f7ff3c4ff4da2df1313584f16f81e86947b3d14db0a03aad84ca2112e4d356c9299
zf6ee03fb4a2215b077b50679f6250d52ef9e9e2c55e7e4043e63b46f080019d10551a2b935a765
zf0588c433e5fe75cdf3d3ead903b32a470edaeee0c831751c74fe2cbe0273ff837a99796a8266e
z4eda23ee1ef3f817495f57c00b85bba5918bad781cbc6ba722e0f2ed6e8575057a8e8581377a75
z5735321a5ecc212189aec78c02a2285e3addd0279c8c3ed911054ff953eb7d5746762d5e89a0ae
z9a13d99225ce8b0f28291a689e211490e1c2e912d4595d030f899c481c20c94bb16b1ec249b2c2
zb0502acdc33469b1036baf387bf64fed11ae33e6d262ddcfd65cedad5271be9bc3881db6b4ce0e
z7d7ed2665cef9e2f7d7e5d74d57601a12646e81e234ba0d032e8882265a59ae5ab6209a20048c3
z8a15061089330951c5d81bd3b670967e02f2220828afc8465a9a5685805176cb5b2edc1b32865e
zb6203936409489b4bf8c9219d04b5bc0b3b65b0a2b328df42996f0fb31f8066fb560ebcd12bbb8
z0ed1ae60df0d24639b6b4ca6afec9f8ef9160dece3998aaecc0cc523d1d6610c464bc9ae1e8296
ze6e7e909976fb37b0c14f4e1f2d063f5180df119bc34a2e7e8326beb40ec816c5f1f01499326c8
z6e0b80a8e921f52cfefe884e7b35d7bd0a41548709b53e209405c7506ee80d24f8d460d4418a3c
z2325677020321c3ae5e2a446ff6bfa88372e231548e9858b7947a1ac7675fcba7058956a247d3d
za9581ea0348f6af1046e051de809480d43bb7c9e8a19a8d90ea75da5aeffaff41350767d3d4996
z86033b0373436ac07ac14d75113bcc5a1f124af18b92ed09f422fc3b0f784b6dea247051809ea6
z0666b44627eb513176e5e764ec9a901615030000938045dc4eb556b16b21bd1e5c3ea44e2383ff
z1e0ba3ed71f7030263a9e4dff4630cada0bf761e07e7e298d6401b9449a66fdea9e80711d8fad5
z6309a5e8fd279c138837ab5bbc9ca60fe40f7f3d312ccc94f7ef4229937acc0dbf7b71716d51bb
zadee65b84615cd1157fb68bc962d11c5d6838a02efe9cb3e294b4f2608cfe3b288cf6eb1f26f2d
zc4b103a9d9637670d2bbc63ac6af6bed98c3efaefc5f4cbe7e1cbcc517da0503898e442c747906
z57a9f0766a764bcbf1faffa7445901ec4739016375c63df2a207717d314d53591cbd87e9c8cf84
za86b32cc6b7c8574906d81d0db3b50667935e98bd92f99bb8eb32d633db25f381767181ad8d072
zb1a8ede9480113889e2022df769edc247c3bd6faf62420f4aef17574f9f670ed2fca5297dd2d02
zb6653b3572fe8c872abe94bd970a6762b6fc97cd51a91556e923862cc0e20bed836b1ebfaee6f8
zcbd4ea1815c59922e372bb93370ed290d8b9cf43375c2d9859a66e77247fa0e10950ad4b552c24
zb2711656459b7a41901c211eaad9379ce0d95a64a185965f61bd6a434be024d98776bbe58c2345
z42ffb7c6121625cae01727461e9051f47c62d1c16e8dc8bdb9921715baadf680374c18e62d270c
z13ba31562d1d312fd0e1ef53d86907226b70eca4549a2101fb1f10e78191faa09d97080bcf2e8b
z8891bb2694c3fd18983e409a5126a634b18d19a92bf5a3fd7b130edf571aa616acc17e0dd3f077
z8a67ad0051676ee20a7aef779a0604339c954d548fa2bd03e89fe2e7d778fee03d1a69091d1f98
z630b0fdeda4f2e7148e18d45fdaaeda77118d27d94c83404b6237635ed194b9824cb332f665fab
zb17a20371d76709617347497e638d1dfa417ef99e23cdc824c00af9f7b2be349abb1b6babe8fca
z06e2c10becf8cf217920ea08605b0280d0a440b7bbc1df4461882d2fb309e44ce228d5e69c4788
z685855681afeda2196dae82dd37a14375bf699998caf856e89cd66e5ef3a09a364234c0b2764e0
zdc6f87be3b3f12f1dd8a20f21d5b445e05124c186b8e01f869e9f4540ee3514bf67631ee23d1cf
zc67ae25d7f139380e3cd5ea90b295a8f07b159f1bb896565bc136edba5ac3b26c30971ee040ff0
zbb7789902d3d6d1e178b349b7f179ba49f9ce1721c42c33d134ede38fb2eed86a7b6e45b9e265f
zea79467d680d90357918ceedba806d9e1f3fde5468bb12297087499f265fedfaadbe0514c938f9
z7b364aa8cb3cb8fcb3268b5e45624f8af62f90bd98617ce62afc476943bd36849bc7e430dd1aa6
z91be7856940307e9370d1dcb45e0496bd4af39e67417f3d0eeca901d6722dd2fb0518cac92ec3a
zebea9404e09b7176c5db973b20d04c32811d7f3239ae82fd2b20285162a975b0d73a127071a047
zbf805f6821da094845e354d4c423e091d412c3604fc03d0d0039fd3664152c1a568f64bd0e730f
z509074c420dcbc0c3ce65962f99cc1a352f466eee958e643e25686ebdfe9aa33aac98151ea6205
zbf435d028de6037c50ae6d0a31b677133d57503dc36930484516e624d88ad8fb23f6c1eff6f383
z6fd72b45ae79d075d4a4eb3b4e0b61e09418360201de7aa8ba7dd1e553603201a19eb485d35a61
z22b733ab60115f0c3530f7273794e3257999b905d8e76389ba3153c355c7d07ede5391a5ecea3b
z2eb61e47ddb859556de87f9106d3a7a3b55d9158d94220ff984556218e39d989a5972dd89adbdc
zd2d0f6b48505129695120b7ee5e292441e3295aea054d39f0496fd83f907a872c362a9755958ea
zaca62e05f55c347cce916fe3ab51cb0d02339120a99cc75971a8e8c03461da3c0ab9a601596500
z30da8f159e954b2c86d948cd117621f4828718b74ce0f32e549e2a5f52d369fb0aeb5b7daffab4
z1dda62322ecd0fdd7d52b73171bc7abe784fb0bc011b0a98bb8d9cb605c78af740d64813b7c714
zaa5d6ffcb2452da89e9abcd47cad7cde3b8f31c1273447be4a4109fc94d6dd26efe4f6c8bc9aa4
zac44b3738e8a2d2966cdde3c2d313785bb9e4af742922f810a17f2dae7975404e1379afe376fe4
z015d2acefb3d4169ed556e6e5573839f3c848b4607d1e052045abbf7ad12a98f2ab35ba9bfa26a
zd372b38f590fb73a68fccae68a18661c39676fbbdd9852dc3ce1a86c7ed99e4a3d700ba1726fc2
z7566cf79075f61c4d9337734ac00ac3f57af13e364ea7b264b0e804ca713e98540ce6b002c2c72
z5cfd43c4d3f9a9276ad771c1df34c38258ef0753bbe83c8549fe58500977a8614dceff0ddb69db
ze819fe5627719a9dd60cf63cf6f3af1ca8486b180e09dea5180f7eee981bb40f8e8acc76161d9e
z67f97a81986170501ffc3a98126ec01ba8eaa6e983a833546c22b63f0c0e6072a78fc20fd0f8a0
z8e93d2f4d25d7282e007ffb944a1b156d9fa7d146eebaf17d45fcb22d64b4fbb9cfabdd0ff2a22
z21e61d861ebf2e0e3d82e3b760bb33c6a54e3a3b176c58e6d5cced340dccb95f6977e1cfb17a0b
z25f742233b0d661566482e2c6a46c2463c4c2d581e8adbe6ba41c0dcf00fdef91a2b107f3b6fb1
zc90d1f4f33de3056a52de343be70280b6a1da3ac9cf069b394cfc49a31ffb2d63d97233c7be441
ze89a5379faf066042846f7144ddc3dcdc44c62c9d1ae255a121a9c7a50b1eda4dcf815dc6df8f9
z09340857e1d24a73d3408e05133a139870c077fc26791cc16b1e59e1d70aca5706ddb7c08e4744
z762fa9757c660779b1ff7ebda807d62abdf347ea2f6b559b9be832af0def3fad119cd67a45d757
z4321fea0a696069c26de89489048439e79847fd1ebfbfe6b27ae8aec5f1695dbfaaa6ef298aab8
z1287c09b7102f19dfb726470b1acc6ed65c1962d54bc871d04e5a597a8d2382c3913624623781b
z33d2841d9391fa2aa385890f06aa79e3c497ce960463a90aee7e7cbecd259e385061f177229496
za4ea9357121c274e3ab349d0b12c369d3e66a6544938915802cafef7813cdc94b2cf8417483df0
zcb51f1ff22ae67a0db854549e0bf97e038fd113967adda0ab07802d4d3abbb20c0825d64e0ebbf
z6375a388c2f9f46bf232072a9b3185e29f496d8ac7d6b87c23864cccf39434100bfb3c8b2792e8
z4af32ef7dba08df69c730f2bee4ac185eca2a454cc19f736ddc96f90bfa4ede22309b1ce981435
zce35e4cce3678e8ff972ee132c004ffd7441df7d51c120d8e6100e80880a50858dafb1af762c51
z1ec642582889b4be84c26249d2798ab04a6633bee516cac42a8c3ba4aba71b6e23b4949834fdb9
zff6ef1f5b215b8ae525b57cf0fa6f1f5198d64b2204ef371806f4f5a1b3a746918a5e9133d7f80
zfaa0c788b93b6207a6fb964f6ae48f3bbe49260968cdb9623c3dbf3d2b55ef425da706a5ef2723
zcf08fa0ab108286ebaff23724e8091aaa37f8f82bb726986cddbca894df4e89ff87f2796cebe2b
z113eee801d3209ff7da382ed8a0431eb00267e793ff45733cb5d8add74bd8694be2ec528472b8b
z80e159c0ff351082672cd940b87110236217517cb741345ac54a77311239222749b50885ea70ac
z2d322e22c80d9fbefa18e929ee35ec32efdeb28da60e227dc2e64a0392511df8d640198982237b
zc3b8653e6a1b4a66ca0bed29bf09f0eeeaddb641c4e22f86dbc0bfa89153fc858eb3410391666f
zba150e4b63e1ed65747cf9ec412bbf92d3d343f0be248be39d8eac76a1b2f091291aa7da42eca9
z1d7a46859019070de047f2fa4ae6958d88b0b345aff32498e43bb6eaeef431bdb5edf29577b493
z5b671a4c2f6ad5aedb660e1e73521c2e062437367be12a2a35571b402de7ebe1f233dea0dc5c2c
zac6e1349a8017e73a79e7c4f4b10abc5f96eaa30a210ff4811af15fa7a24b6c66ca67aadb7b19c
z4c3c2aba87a8853826c2f9dd2d0e66dae5a3437e42de480db7b74571ef16d9970d62e4910b28c6
z7d62dbf8109f094077f411af5fa5140d9dd25b06a70c9c2f7f9099fa8dbe94c53574b5138f5b15
z34b6905d000e8e1479424a20d1374e65dbf73bd4baef9c8418b7b4c6f327e68e2955066d73b315
z8385f5884eef68a90dfda52f531dad73a188ac5faf0fb4911b16aa5177c7337c67c4b2b6b9f9d0
z3732214e8348920d2c9be60cc8f4b8e01898ea617f8fa47ebb16dfa0f2a1f01b19f88fcafa5e5c
zc30302183a3a04c5f231b9d442130b0360d4df618040228b2d212d559d663e0728c15a0a0f139a
z4e2e01d19cc48d8607bd878e228562c90cd266f2b813511024abe94e865733e275384ce2be0af4
z6b035a9bdedbc1e00d8e242f53a9e7000618188afd7102effed109c4f80ce6494a2f4510046e54
z4cf19c98c3aefb2f4af8008d2ca235428c5384446d7782d469b16cf5442a895b9b9f4d3cca5a7e
z6a9f5cc6ddcee155a20e86cb3b02b5d52a2f6ef007b64a4cdde7ccdca0a1f372f6f4175faf8bcf
zd48e87310789cf7f3bf0b7e8676d97e32218edcdf54aeca399d9ab4bc3cd9e326f3877d342c8a9
z3eb6fd239613792bfae71ec71e42a8e01031b157bbea1e6cb72b727d19465a42d208bb374181d9
zd3423f2ef2a2a084c70ad3fad7eb7b3a3acf580f126110b0dbfaa125eb710b8acb3b20794c3954
zb13787c14d7dc56a492a2f5989c4117ab75fb3224aaedb0473b3d97d29ce00dcdb81c337d1b585
z4c3878d5088a965274f1e32e402bc56c1e021c286ac06337ccaa13252081161a7ace294bf75d8a
za76ca3502e9ac37e437d4147ddeb416d9c57dc14cd5f55a04888fbcd5ccb384b5d5348d2ba0c7e
z2f39f6a1e4a285c95fe7b1fceb737f654fe7c5b1ad21b421537cae86bdfa223ae60f7f6c3a5a0c
z93d700a544388b282a192b2dae7c4409641e4487656247c9b06a9af182e3a0882491c6df243701
zfd42dc9117a9fb22655a8195dfe0c3223b72f0690f9b00db83ebb0487badb82e88202e9b2fb9d5
z634a644e0e867688ec6252417c6a73aac22e42cdeaa84dc08229b65c7e7dc3a33f1c167e161668
zf4e664b419c64fcaefcbb4c72ff35d46506e6bf0ef50f12c942823cfd1a04d866f54dd34762ec7
z20d3a23dfdcf48b4213ec481870cd5741f59acede658842da83a25f6fddc0e88cfa2313d67487e
z90b3d19acfea1d44415e9c72e682b1125f4c6097be88b2040634284451667d9701b416b7e83e79
z8ad92d306ef4797eb99de0d027a93d30636562193ca0cb812991ea3b519c0506490c418d1ab46a
z96a22767984c832bf32877e0946a839a81ca3e64d5b5ff864c02c44718930263f18f0ae4bfd7a1
z3a5c4c11e9f5e77c096025a6fab9c397c0876dffa74af87c9566a8c078b92efdde334f2889627a
zb613dc8d7c63234c0b2076f4111858850418d9baf6b0a549b3f12f0d4a24a8263c006c7fc6c894
z42a548d713f8823d2557be51d5fd99549ae86f4355ff8f92ef21270868caa5545c7317a03b35b2
z0b5773829fef4c6a051a57f7c26268c0db612e34d99a059acb71fd09918324ac1f3a5098d53f68
zc0bfdbb465fa61d323205b8f78e26f99ba56a9181fcf466682f7abb8927b47b11b3bb38e39e582
zc91498ca77152d5d94c838b4157bde01946c8b559dd11d83737a173e3c92ad4a010ce9040a583a
z0defaacad6bb0cca9d9095bea0a9df87c937a5c86cf3f2cc7b9ad208779cd8f454aaaffa5dfb93
z15c986b40b75b34eb682b4cc58748dd628de55a3397b4ffc4bd714e4aac7826df4a3fbb5d23c5d
ze5be0dc5e46b825ac2746a01b26aebec1dadc9f3e13d361ade5a449ffc3dd09d623e84c132121a
z699cbf00c86fb5062b71944a03cdeef2c996426f619d3157cc767013faa23579a414dcef5f89e0
z9000b9950c76f8852e6d03cea09be7e16c57d76a59d2a65faad2b93b6f80b387515f056900f8dc
z9b07a0988b8edcd324b6251b5ba21f8ff15c2e8c0a441a616f301be2e19844dd61be9fffd1b123
ze140477d7e0fc972973e22e1a79f8ff473dac61fdc1414b20babba8047fda91f65f18fa94d6f02
zaaa3a1299e68b620caf25fb322c39887f16a64720cde942de8ec28dadd909649db667c6defc85d
z695fbf8211e209a2ecbf1430f0522c17aed9c52cd791c27aec0c8876d55a3de255701b67443731
zca6827ae7095b5c06b5665d4be42e8b5a54559895f8157566ac2d508496090ba4e343a3fe43671
ze91f0169adb41c17226bcd7cd405d9f24b111b93b3339267b9d64d49f7368fa1547a91020abf8a
z3384047d4fe585411d6837eaa10c8c2a4fda2a846853f4d94b73a093e3c0ff0044bab5a59ed3f8
zc0a6a3a18fcc56e2ffa858f07a44b07e6841c82481680d6974670ce81b8117f7fc5be03ab4b1ac
z51673eab4e761a99c5ca519af55b95956f921de3d5153aae9d173d999d2068518fa02ffeeff44b
z7f78380d39e393545270c40f4be4cdb3c328ce15f5178004e36bc9bd342b36532f1e3cb2e02134
zd468a8994a281975d4393b16e44394cf81cd75c0d7b4209c01ea652d87e1e4cc9b7663822908c2
zc78e4cfa81fd9625b9f109d56b150b52dfc93209569d232b580fa34985ee90eb9a7e4d92359f93
zfb19e52822929d0376f30b3ce4999d768bf412dc8c74dfce90e7551a17128d64e23b9db74876dd
zfb288d116a9b5afd055056fcaef56f0a839148c0fd62fe484f185b47198304d7deb736d8a7084c
z1594a26e59de3e643872b38b454a3bff5e81dbec06dead210368c1c403398f8f82ab521f6c9005
zb27bd503039e932377ba18cbc10192f3649997b8794cfe55bb85c6299556e26131bbd05d32420e
z99c95908094513d17d56a1fcf1755b63143eec6383311dfcc1a03b80bef1c4ae4de53b195b82ec
z62de38a0906c8fc64dde006b70158f688ca8ad7f778e34febf08bad9fd1bfa9414bf4c64718518
z0afebdf05c39afc660ba7a05cf6fb6e4a780c83716f966ed3085fef23674ba93cdeb19b7c96d8e
zb49a19ccbeb460e7769e0e5aff952359df4345204f0f7234c36b194bc337679f8b4e24b833b4fd
z1172efb7b93146f1b14a434bf85731d5264fd768ffe6d6e46da788af72c055af5e1285a8006e5e
z5bb0f168b35d90ad7aaade4324efa4406586fd53f6da38b371ba9b80439d908825b7ab50a37608
zf622a065919b26dc3c2a35964ab81110d61690a81b365986384a03f7187721feb4bacf0ae4a19b
z3be5c2dd8c5de8d98bc8ec0a631900f7bcc7d69310698e7016863e72ac63fa0512a0ea56f940eb
z7a326b0f88e70aa9cca8ec4445fc4e4fb90cc56331a4f528f65b770be550f04e3811a65fb9ac67
z3a18a7583ddcda6481e0acbdde239dfedebbc057b9f867476f01c2939521d88b852fb378e1478e
zfdeaecd2844b28daa72bb35e61f3caf3ba06f818503442a1d13497dc9c4fcc1115ebc5812c46c1
z6c1e5585e72dbe1de3220426261a5c8d9658a5e167d83c02aca88877961869862994ae24f246ec
z567184c6da0c1532821c822ab8c69e692c16e9eef22ec3619bd87a6405d5e91212817c21e4e516
z8d4d87078d8a7429e480cc8d29853e40b94de8ae906c9cddec27dd43e70a809f0d183697eb3698
z8720a880e9adad51710ab7afc163f4e573a873c18fd1392607d012906e68dcd05371f2e3108c6d
z8dd9119f0ebe12c0925c2c3251b404ec576dba00c30ee8e362e872eccdfaaef4096c5c3c8c35c2
z43438d51833df581ecc48186f2bb4d6d804785887d3776e167adae6dceda826a0f5e4028f370d3
zc52ad96f49b09878a3d307b27e328a48831386353a4a6e5947b31abd25f0a596227df45ec01503
za2386a23946a78a534a0f5ab052a5fb564dafe689a158e82ca1e020cceb5d7b4152b3f10d07d3b
z69061ff5648302a9694beb41d596176285da4af5bb86ee382d116b70d978cc7e9aa9e7262518d1
z552df0368841d67fd4dd18578e0015db6bf7d5c5d28fa0a6fbffa5842d9154753166a2b8f419d9
z0b3281df2ef827cebe5169051abc658e3dcdb9d055b5159faa4130cccbabaa5a0a311936d72718
z80efa23b28087b27663106fbf36bf6ba28ba63c2828761b8b71584b74e8aaa3a6a5a0f99088254
z27eba50b4c236ddc3e8997d1b75ba6357f1ef74b45d7b37cc09e81b0ee3766e0f1391b2df7b78c
z88a01e33af441606bba673b750c6e4d0f46c8fe497d9296f31b288b3c1dbd84a2a4ab2b8bba644
zec78694f85be02ea4fa8169d86efa3bd91738b19f9af7df44657638ade968d3f7bc0127c1f0af7
z0460e13753d26003bb02fbc5adaf193d8181346626d03b3888645605c7761b5d1c893455109fc0
zaf846fcf253e242b4273e26cd4f10f9c8e6568ad36053e47834509187ab3c04ebcd219402fb892
zad84380e51991690065760a4a40730746bdcdbaeb8e6c589bd2905b6fdacddf63e202c388a8eb4
z6c8d9bce2b66039eb4051ad444d62e9436efeadd43dab9215d3c01d570f364b30b5b926ec6d053
z2a66742f6234f45e555cbfca462e6401b5ef4913110376d9602db5d87df5adf86cbaf5886d378d
zd1d7489f516e27e25393733f7fa5b4a89041ad5229490fc3066034e6b14df063faf9fad38ad07f
z5d5e61bc5fbde5251df0701473ad733f8716bd3aeafe52ef9f16ae1482fade0d92ab44f0f8ef8d
zfce917715c32dd97b5d40a22579f96eb4eda948ffd2e117d12bee289dde97bb375fe8b32b08b52
zc334db30455e2b366201c2afbeeb91df4902c7c2ab52870fe280d854a4960cb25de6fae94dc4d0
z9273b5fc754c3f1518adc7f4c2a06568b0e0381cafbb7202cddced8f0605dba545f3df822e3060
zecbadd8b136248935d4153e7b32012790a4eb19c69249aece1b860d902b9585dd04638ccaf1ef5
z24e60ece2f9026880f489f246da48d746aced3e7249ab6876571109e340aabd935f0d66304e01a
z54d07c9d71b95e72db079d443fc8c9c4e06d6e156b3ba5ed1c53f87abffafff6a871b72ca7a782
z65200c131d65a555d44c4292fcfd0f4d9a15e96ee4a291f89eefa002d414c74024fa8fb62403fb
z685d758d7ee109dd711348a67acc965f521961afda6243173c65022d08c265785bdcef23bdb0af
zcac561b2cb2f30b04cd7692555c74c3779caf43eefb399428b36d4dd4b4161bcdf31b2f785e38e
z966c545bd5c54fc566854e37a56dfcc72e9d90aa32f9f429f7fe5f35d333be6dc52e2085116eef
z6694a1e29d1516c80c0e25e9d0f4d3d81ab0b313b6d5ed74e72f5a6e0c85b6c53c5e603ddef93f
zebf429e5c0ca9659d5874ed30ef36fd8824ad7e3b036f6232deaa3b67ec4212d61a77e29d0a7d9
z984f49eb2b6f630e2d7eaf69f256f3c0cdcc43444427646636cb68a2487250b449023e3dfd7512
zcfe285194a0f6487a37eca558119fc22d99be78589e4fba36186234ff7f332402218b9ba2b7526
z65f05bb51b8a401c50da4a7145b8fc80c2702dfce701dde73f53a5d9b6ac089f3518c542d4e927
z88627f9ae24794e6aa6f8cb7d2dbbc2ce3bb38938c5c0d79037462c617923293f1860efd71fe7b
zdcd3dd8174f2225c4432f27d2e8b8d457fadc71d20fd84a29f43da68eb422e31ea9559c2116a81
z0b4165a4f917762d3cceac02fee99d77b6c18af6d081c393326016f1f26ddbb29187f182766fa5
z0b6336c0279553bcd6c05590340a4c73562da20cf95f65551681a5b1476bf981124ac96b298995
zecb0ea5e2610f20e162e92f966da780f03c3880195bfb7f3064a15a2b1bf1f798ef7a496459fe4
z50e54f23e888d84830a6ec40a6e51444a483b452274b78a33fc066205044435519eddce65a8c04
z32ffa7ffae2c260a57ac78fd2983e713c91f21b74b94361c9996419def1e6919b1c3eef80f78d4
z25e1ae89a5a1d77178dafcc6248b6bd0f490d5dcac7516a9c58547952103d8e3c026c789134704
z602b5df973fda5d8a883101f409360d0e23b0d002a20708ab7c5fbbc2fdf0fbe1c221adb4bd8e3
z62bca2adecd64ee42f76b9b4d10a1d4b1019a085c6c07fd3135babf468956b48dc2389b311ee96
z0a498f96cb04c28612efa973880d9ac1021077f2f2bfca58dea6b7d0076a5542c51497e6249619
z334c4b9560788039d0c37996ed379970bc7e4245af77c2a8dd321aee670c97625d8e99c18ed5b3
z241b5d3ebd83e09cbace7cbc648ea2adcd6b2c38d4c09e5c2ba7ef85bd71082c660d63c95c4dbd
z66707d626aa52af6b393946e8d815b946880459a960baf2dc950bd5cd4b42b974e6589eac5ad27
z2fa77910d891924426cbb4a87064ce822ffb92d98d31c0ff1c035a4c1c4454c2e8b79afdf4661a
z6a870b0d63121436bc15b845e83bd5ce66b7713efd305d2d9f790aa6c13869c965db891ca21f7f
z634982d060b7004e3768eaa772d48792f08906cef2e5052d164620f140b82010944a8c2da478ac
z2e0ddbb5297f53f5ac010d74e6a7322af1513cdf4390d777692d03a36d026057d465773175c084
z8d509ddf0df53cba8a08a1053e2bc2ece2ca8798f65a1a74e4f860b82ff2994d0930b890444654
z635c78030d528baa29519396cc6d776f3a1b2518eeeb2669ff300fb154465fcf89d887fd2959cd
zcf2588ad223f3debd2f8188590379e0b8a953a50f672b67c3cba9695dd49fc441b590c27ab0bed
zcaeb3a64b9d331c587301497d11e83952c3cec8aa5aa6b9c4a82eb3124970a3be427d0ab0ec920
zbbb0f1e21b60c79e4a58f17b49f2faef378b91ced304a4f00e8005cb476f9e658027bc47b0d6cc
zd1d8bfbee14d27010162b5a3a60ebb7663987921450f29771a61bc9a347f4afa5d08f7d281f3ba
zbd2fde9487f0e29d00c95b5c789cf2be472b9ff1b278596b349c3b80a1a2f847b00b39b421155a
z57a16e9af6ad7aa68ee3bfb3df3297579bf1271da50072a3c35475b551d7100c8102ea987b94ad
z0969261c9e606c4ecfd3cd3140bddca3a64b97c5cbf16552c207e2bdf432fdb108c7cf281b770a
z53f11ec057a824a46f9debf7339f25d9035da5018ed2297a336f77ed07971ca361fb281bc8d6a5
z524c78b98758d455d718517c8a29de0c92e6aa9d52e3a1d7def0fdfcf20d9021d60f4adf1678a7
z37963a7cfb18dda9cf4deac58495af3901923a2d07b12c7f73578f19151f929029dd7b044299f2
zcf05e3d121292b2045d0ae4049ddd878f5f11ed77ae5d781965191c346f14a912edd0f6d9da154
zd755767f08e78cecfec71fecb8f02c8be4bef90bca809993fc40c12971a6dff925886c582e69d2
z1521fbc08b969ff2b9b106e07638baf639c20124fae8d080b0bfe3cfa7637c8366206b88f82ff5
z6fdce24fb803f08c0d2c56d8afb623112c27400409ad024e13ae0f644886700e997bffc575672b
z437118240e8b25ba2c02fdea764eb1f323524d05efceec4b897bab5c028f77b479362211ec1305
z3428e1c9d040cc4231153230e3ee45fab9740ddee37e241c8e7589d50c52e2aa555ea69ca32c05
zd67376485122edb44fcc403b14e48b32272e314738b5c690f87260731d7bf9f0c5845b6238c6ab
z5ad6874acf2b5fcdd2b02eb9937064198f6c3e7715177565991679ffd14a274c4be94db8013b52
z0c3a2893101bf8242e2b6fca6bc0297afe66da4a6665b84b46652e51b7f87519efedde1bbb8b74
zc3d297dbe4de93085e2794293b47352f13f771e39e49d4c91502ad5cbfdb050745b57a95292f71
zb32751b3ead141e836b8182955a9672ba6d48cc725f7dc43e29b33112a254c7046b889304728a6
z9be1c5871539a49dc64dfec9575542413dfef90c92c804598541bff78ee67b1a85278d92682f7b
zf7ee5963c85371a21a46fe818d2ebbd28430dfdecaa17f7b917b4e972db7b2e53d3a6f67d98b83
z6beaad94df3edabd04a5dd9fb85460de41610fef3de6f14388b146cb0870c2e255bb8f4220560a
z7fc1af7d604c893b5667c4e493ecb8bc7695498a3322c2e96e4a6022a5dd9789843c15da1b31fb
zf025066293df5653fb05d22425e5b8290985b0cb5840872df8098eb8e18b97fbc901c6b141a47c
z14ae44c2428e04b1dcefcd273ffb8e2cdc3c187fcbd48db0b11e649179333824b9fac309d37287
zf0df8f248be7e1534f1e5fed0ce14dadcab14dd7dd99381da35ba3d17a4cbee4775763a4f72c46
z090a711f5f784dc4967647d94b5930f0e07aff7ce2fd5c458ea37045812da0afd567e20309b857
z78133aec2011af5b84bf261d4e87be2221f4574e97a8ee3e248eb6058a01b9ed4c8abf867f470b
z7927ffa993932a0bd2719c632fc02969838097aaad7eaae3feda8f9670d8c217ad2740c0f9622b
z39037b63eaeafec07ce15e61b9e23ee7c51a517520fd893e3e5f19da1b63d98e4d5ea329dc6dbe
z452bb151fef73515b9fef4becca403fcb4e0ec17e75cc0107abe7ecea40c7557a0d7e6d4a14915
z5bc9a1b5dadd618ad96c6b98eb891625d87ceec75a243e5be003c43f98734e65af9f51760e0455
z10eef2e3098d6882a748e75d396fd3c6d028bb044354ccf212319fa5ea88dd2113e9d078d042b2
z85ae73a7d19782c71da67fcc1de2f560db39140bc747b03226d437baf6d9256381168fb9ce7705
z00c0c7e4f6860c0067f2894c0ac211561023c38a17639681e697038cb993494efa173a54313e59
z51507eae4a8074998447244fa01bebbd0b49905bfd92192f535c48f6c88327540f407f16d73bed
z44f26d36759f6a9a10e694323921ffcb19c6a30c6b70c4ca309bd79a44c65f31e43013f1e71256
z739fc59a4e3e903ad2ef3ac9766c38304f613a594ad66c53e215ba04496ed7524be52de58d27da
z2febdbea4d47d62255d6b25ca36eeb77a8bd162aa62fd6f342942281a3314adf69834f3f9f10a3
ze97ce145933cd764fe08845da38e001dbd53810bbb12a75f6e710dc38ce2d7b3726032c5583a23
z1d187baff32bfd137a02b7faeed4c5df260ef601b7ebea8120c05e451108a8c37d7c4b48f69520
z0ca32d8d91e72d4bc75b4a63cece3143602f216e8a082394992990f57d39b12fe763123167a7ae
z051f9c3e96ff8ed94c348cabde60acc57844552eb131636f758fd4c1dcb80bd1b5f0b85bc7e9f6
z9f8e303a2317590b3b55ce91171b616e264944e6f6f9238046465e779035fbff9fa23aa85a75ff
z4958382ce30c91217bd078c8794db0e927cc439f7e3df33f8f8f10cd56726c57a25a7b35d5478c
z1d2f0ef6a34178afd8c5cd9be80d66c77a4182d2235300fdefbbafec0af1b1a7ccfd3df61083ec
z4b4ba15032a50d692d444cb36345d714a851f6c31bd518a20e5e268df6a551d339bb0a87588d8b
zd874e8b8e6e6f6d08f412bdee1b2cbf57390474897c67e8b8381bb065714f1450c35538680b5b8
z2e37b96dd57be1e3f22c93939153f2130ec89964358550dd97b21a071ce6f2f005488be77588c0
z2177590cc920afc6831ee7db80e10a9480b496404942d13d183dd1f1948cc0ad4cc984b163f07f
ze95ad7ce18b32d989f77ba0cbdd2e24ecf97307a52ff1aeb855a120e46cff6c0a1b4d458c27a8a
zf71514e9c2b5a897e726a21ae1f71cd29868744928bfff2d01b3625ed4e097758ccdcb7ca060f7
ze5f5b7423a8b823f15b6689e504b52d226640ec6d6c7c9a8b7a45e6aed430388e898daa524b78a
z5b8cb78e28646af018efa26d0fa5d0bbdc2c22ca70680d666c1f043ad4007136538305f9e1b22f
zd29bb39ce4af21f73a218580443d179776c1950f9acb3b4287fb552eef28dddff9798aacae4756
zfe8796c37d65e9e745e223a3e1fba89f83830a99f87de758ab0972f786216e5acca51d503c80eb
zca4f2bc05acc5f0b765c9091a4b82485f7b784c812ee682b9b8ff2a64fe1f31e791b6589834c86
zf1c6bc654ffa64e4e984f55eb71e8eb3c7203557faffd82578b6c9aa5eebb42b7a96cd7955d6de
z9f0323e8aebde761fa0b6beafd36e42d269b364aeacf059f3797bd7d6b052d16d4274abdc8ddd2
z43494e1690e898a6d2a4a71b005ecb7c01abc911aa9c7ebb0f871594ac616bdcf3ddd2a50ab925
z44d1ac974e21e563b92f1815e4907489f7e67f463f7104cfc97c00a66e9c69501bf46c1a87adc0
z4ef3cc044c935a3ac8548c93b6754eebaa157a1f9ed3c91597cd5411b4610495a57960601e27f2
z5d51dc07f7638b953f1a00223abd6d3f785aef4789cb1fe92ba6241454039b7dedcd6aa74099f2
zb85484d323c3b775156156e5dfb8b8f512ec46a2222d7aae29646ec75526bc508cbaf74e12c608
z30ef86f885033c998c0fbf879d880dd5c556a85a9adee6fd3e73512de1a772c55a1553e6ebe23f
zaa89f978399026d9ba52cc99bd8a116000f970163e4842aa0e06609050c7f171aed87d72c99987
z94a315cc7753a0b3e3959481766ac5c51dab1b680204fa73d4dfca80f95ea52e44ca5f973f1de7
zc1dc59b13e8a848d0af011ef2129a8bc579b55a9fc1882e4fd2afa0312454318f7032ce1a9f9a0
z50aac461e0c2354117a5a3f9475adb6c637aba709704f8f8549554a33ca2cc81bd6cef18239f1b
z725f9df3ca98b986c7225ed577d3c6b81535a118dd0fb139366142c0f2c54740e22706a7af0fdb
z960e3531312f9a02d2bfafb5b6f4ed57b41c613f60cf0f05030f1e9f75336713e9107c04f22d00
z063c9f6f4187c14f2d8e51ce211315f6b3143d71eee279701d63689968678a22baa7ea7f806620
z9fe681cd7bc3af60b0c2ede6a9547ca78ceb6f4b59bb619c2d16ac51122734248bceaa49a68fda
z612ed8c1e5c2f05126633d88f5c3b4d23963e464757e5142b57857b50545490825fe348a140354
z498fd1ddbae37827af1ac2a32b0084ccb28ca3a3f026994face11751a478b22fae479e3f4baa2b
z343c3dc76f2775bd92ff00f3dbbd228c4983a2fbff2e90661456db7f971c3d9b9546725c41e829
z05e2a0e656f0e17195008971a220d418c295c0bb47f7ca97ffd98f62897c2e0b4b659e37f830e1
z3e431187447411fc82799ae8183e5c202c5216b2c9f2626ba6c309c30beb120d25ca20cf544f09
z34f36d19c52e27329f63b7a990329bb915ddf8244ceb7b698d1067f7d7766f2be86bcf13fe2920
zab97635da01d61337bf1d65eb72c2a8bed0aef25cc46ee704fd351fa9675a077ce401fd54fc0e5
z3760c70850ce42bb75782a2efb0e0f957bfcd042b7489c9b913f27c7643cc25fb6d73518c1b9be
zf97657496ab1bd90a7a632611fe283c2f84efd2538fc728e717b4b104f107762da4dfe5304459e
zf82d19d16c87cf04081c104d688953d285242905e5f3ac055247426a9ddd96fd29658516b51035
z3d48bda581f59dd9b59ebcf39c3d1514a0d406546007f6083077555e142e7aac2f6b29d8486c66
ze00465ae4d9ae418fff47eb362026a595fd9729eb6ccd9f558d673121e87d1b9d19e7f4fae1e7f
zd84318c16263118d59637e1c577382bfe9fbe96a0e588cff300e13ba5e1014d83c9f01b68090e0
zf3fea9f6451daab77f1894ec9baa06f65eaff1a494e6c198181d9791fac61745d0462804f0de90
z7128200da9cb5fe7d8ef910662058afd902149568f9a716125d48cccacb8b8748bf849da2be567
z8f485c13f22ad3ba607fa4ecbc8fb63f45e364c23e5e8c224a58f77b92aad005be81707e20101d
zef1eb5310a61962803b7532d8fea5a1419291bf8667bd642a487ac4a897c88819457d3b23a7f77
zf1d16fda24cb4207a3694476d949a3e8f8082caa94763272b401a6933ab896bcb643f205973b80
z45eb5c8a370875d0f363a8856b4b9d8c343f1e8108ead9d8348e13eceef6ad7325c265849a1b30
z50c23ad0038bcde166e9f018e26fa0d2f046289aae9aa34e64d6d64ede0c7efaefadc90bf2e2ca
zc739cd52358d8bdd8edb2f0bd8c285c4e7ca9e68ae5fc3592f992b763d1bf3d61b53a89591f3d6
z3c1d42eba51805d2f1bad9f6e04384f301a655116789c5a0a98b17f48690ee7b120461d940101d
za6e596aef684bfd8c97654a60dddd3a747271e58330e65c376b5bbccc2e190d81ef542aad7f26f
zb599470d9cfc7e4760488e29db51ddb17753b3eb6bff0cc318fc4c68c500e24f9c6bc3e5997a59
z37bc41ee67e9726d3acab11a9cc12cf2f5cba6b1c62c5488e00a5b01360deddba47a468008a248
zcb262203c71e81bac18a4c7950e9a578ee71c59785d4018ce1e219935d40dbcb24c3808ef967c8
z6a21b670c7a24aa41d5d4528d0b46b8d848809c88bd60bf32981d476ed8fa7c1021ecf17085f13
z285a4c9ebf65e1e9d2368b104365d9cf2ff84279c41a9715311dfd6781e8aa4aab103e9816b699
z07e6eed224348f86dfe61c591551ba19b6556a458589f40465f5531840c53e37d31ffe99c3bf29
z043299e8506d64760e6a0b2312574d07298eac2ebe1ffdcb8610fd9569e6528bd08e5876dfdd42
z268a0b224ec6dddd21ff0c710f84337ebc17bc1966f8a4abdcb9d04bd8d7c2f826cade9e949f40
zc63d3817955600264a62ee67615ff80989db51ecbb52d6de6d262b80a91cbdc50d869484a6a6fa
zd0f62b52d6c1112780b516a2e841604fff850ab9add74549df27b4c2c93ea6b1947cc0037a2f19
z4a08023ab4ff42417a3a5d91e55dabbdd0209af0bb56c289b0ec1b8c8739683d22b2e52d46772b
z7c4b13cdc08f08a50db49fa9252c1dde263ac8c259a0acc878ea74d5a14a76040345548dd7e3d0
z56920529e431458cd3d6ab6cb575e00d63ed779c1f2a61e516db3211f495e574bda891f70837ab
z1f3ad0c542c77028c145ce153b8d1ddea1f0bc5a12e029ee436fc327bc7f3436648000546850b5
z48c68dcd80fe7f368e5197a00cbcdc90ae8f0bc8b59d572739a3563695b1e2caa8b2de08014282
z99be6cefb7e2db5984d8bfe486e8c193183b20f3c29d2717b2d976d7cb62da9e3faf787a65e21f
z82418042bd26e49b5692ff84df25b0115ea2a362233a3fc13a3949ab3f3484b363f1de074d1182
za92ca1fa330856ea2213ad2e45af0a2798eee3a49af32b70738de4badef64d153c3701a9deb981
z56417eba7f76aefaa20b83294d82ab1709f9c29d68bb1377aea8298ca55c0913e99551d16df123
z83d039d8a9721076f2cbe8b38dd0385cc83707ddebef573ec1da0161896fbb4af257291eae283c
z897d2a0e55766d8870db16ce359e64e8d12407407370fc0c614771efb4ad25f4864f0428903b36
zacf471942618d0f4602d21569a4da7a8621b0a155f48ea91a1eb29dadf6f8ee31b7a43977779f8
z10d847b13599ab3b48e7603ed5992fdbef704119157260002268690f3d525974994addb91f489d
z105086e46978dcb6b54a0c51fe5a7c91807a8518f36b7b1a81afdf0003b6d4ccac10372d727d6e
z6057821b7f7674bfe5386107cec8289e48a66e87fe25ba698b242bace8bbee56a3d0da2c3c1726
z2472b6382bdab195437f513549e973b3dbc6fbae4be72dbb6511a7c586082318a8bdca40496f8d
z9d89e9fad9925d93fcd74838899c6a3257df2a8da404b47f59cddafee982e37dd1bdfc07929948
z55cc44740bd1ea5cdb79cbbaba4ad5a157e974fd9fadf6e2843d8fea0e8681fbf3baf3718b1371
z26f7697942ae49441cbce130c1b97c888693a2493c5e6c011ca119d8f8b758b3c8493ed23a925e
z06244d97e7ee996365cbc4e7e1269d0ff6d2a7b357c14492c3357e4b48414f8b33c51546d57c21
z38b4256625cf4cc30d21f30db7427d58e34f92ed572af3f5458ff4c7a9908f5d4f6032f979e746
z16ff6104a8d4b1ffc60ca44cd5a1cae8fed1bc54c4af7b8f26e1be23839990936f7e2b9dbdc72d
z906b55509ea6547d20273f8671ad85d3ff4737fe62581ff14663218721c83b692e983dc662f8d8
z1c07dc4fecacbfc3c603b1c669c503a072c5052629657b492052376b47c24bc6851d4e2c7e49eb
z19b1d26eaefbc15c
`end_protected_0in
`else
`ifdef MODEL_TECH
`include "qvl_i2c_master_checks.mti.svp"
`endif // MODEL_TECH
`endif // encrypted_0in
