`ifdef encrypted_0in
`protected_0in
ze74c34e226135848fe16db9ffd31815111b6d7fb642c521a3f628cf6da949865580b22efd062a7
ze90adae0e65e66a2c36a587d0a790699161455169ed55a01f2084f11770a774ec4c588039b380f
z6de9c5084882a40b79a175f5c2114b2b6d78b070cb806e1c0aa9258297f4687ab308bc470f0040
zb0b1de382961eeeaf2e279e1462520fc31c119af8f2b214846f56c2b3cd2eadbe4099496abff18
z15cec83ec4a77b868344aa20ba7360908f5c0de2a79abf8b3534b883bb12180f68b5d4beb444cf
z3fba8f13afb0abfe8fcc4294810f75afe452434d2d0f1166236c82f76edf1e12979f04bc35693e
z32ae028996dd85737a8f5adc1ebb94f39c940246e887647b64782cd7ab429b0544c173176cede7
z01dfb26b1f73408344a52b7e1f117f12bb9c8077b34876c2e6fdc085981637012dc9754765e1a9
zc512ce062e0b8fb16a214591f5c81e1353b900a611fe1f4886b57940b41b7f2ce99a7b84b04b90
z916f717e73bd10589c81e207ed77ec660a8cbed5b487fa50acde1b055c8870bd8676023f21ddcf
z9c98cc47cfa2d654ff1365d1f45035a045a66c5dfa827905026201628cee5aae21fb892db766c4
zb5b1406e11aebfd6dfacc9da5ec03b70c276807a3eb15e28ec7ab1dddec42388b9424ea285623a
z248195c9f894b36317ca6e59c86f11031163f5f5bfdba36b10b435d36514783bc1c6e60eaff7f9
za2b8eba90f8fd9a9cd7c932ce34efca1757e6b27183792db4eb9a2748cd3c1199fca3ba95d5fe9
zfcd512e30a61f3661d6f0d353873007808f9a77d73b67c394cc2f534ef756c1d0cd29586c06485
z670933b76fb2f10496122792af3f824a49802c7b02e68a1ad5a452206cd54f492e3ff59765dca2
z526a26177ca69f1f82d5f8faa94e8b5d822162e8931eed4f257b39c3215947f3875ce2b0a82765
ze348a0c2e5a63ef3af742684d34d2a4f066392e77c57fdb20cad55670edde1f2f1285738af78c6
ze274689c0de830b4215adb8d68d36b8f11567a7aadf92d8db968dbfcf256716c7eb73b8831f387
zc00e2b6c048c23be913bb8796eec895fb1ece84622f6a5a0c7db801f0a4d1b451039f9e3533b3e
zba59993f316a38d84bd15702c1971105ad28d5f562e302e1e92b0aadec0c8225d7404263872a14
ze9ba482676ca81103c10508b0c603b52c1974c958eb8a6b0f83efcdd6dc70cdb3f2a4035e8312f
ze9040a5f83c1e4032ba8005e9ad0c9dc46d706f9485067761fca056ef0fcd152d04bd1729979c3
z6e6de056835eaf8977afed310d977b39c509fcbec10cb09c2411528ebb6d935cc4f14cdb98c268
z35a3a0ba1839a9c17ed315abdb42a091f1687053fed1ba612befd7cf83e255975c35b59a00d90c
z4e8f704c4321d9375e356f24975f384e8b1f81ce1912f75415aeb675f57e7317d97bb5aa0bc858
ze508d24ae8902efc2fab06a641f220e5b38eda3ce0deb0cab29e3fb67ae61e2ea846176a6a9690
zee78c4f9777550988dd7210b49d953566061dd5da7c4eddf51e14ba8f73221fee285837b98c16d
z8d690261d61f901c7599f720b7f3ac3bb7028ae9dca5579dd1ff815ed92a0ae50c0a1afa03ea76
z2980f42f950537d9b6fd34db07444579cea81edd3907dd493eafb5592b1f64bd701748650b0c29
z27cb424f8cf392396dd08555bea81ed4a9193027b97e3f5d4d9537ea2131c36f7d940046eeb40e
zeb23de1a290e66a1903223759b5bddf8ead4290403599529c59d05739bbac6f1039c86c3173476
zdb8d882bd7154c6f811b012c3934ba35b8ec6c32602432531ec1d57f89cbca61d8827c069d6778
zd5c718462e8551932c7bc585d19cd2767bb96aed7931617497aa57aa3a095566b48f36ddb9c068
z25d66a166676e4c390553fec9b840757c74431feb3f8cb23a82615d1860c4a10113d3f8535a891
z5544344f30aaf7d0585154e95a9a0b7c5940fa079e719fb7d565a454932880a217da8d40e35e71
zdf4f124459ee721afd81e1541789701d9839681cf0a53834af86f75b531aec0b37130a0056411b
z4aeec635305627b80f3b09e256c4bd73e9587281dc21d73fbb8bebcae45cbd3dcb324bdb92a045
z44981b6a8e501a6a0d1e5e093b1f12dc69f80dcfb15c2b58a63998139f3b6bcf540e183e3db40e
zba56ee2ef282522e1b5c2125c15219f63979c25f917ae1a1b125714e3298126580d4b8185ebf03
zd081fb7cf40e81bd2116680d0b1bd2bd39e82a577a7f1d8006995de8f52b2f7971a03f5a11d143
z974db1695ab68160e9ecf72ed346b87bdda69a86ead82dc94f894bdbda77368a3981a1144d560f
z998278bab273bd93e14467c696ebc01aa07db7d481fec9203a0af5c944d6ae34707134713e1dc8
z56523085a80a48e3d6c6fb82e5ebb08217b2d2cd1887f9aa9d39f4b769ee627c4b2db5cd06de29
za1572214689d8e0e98895beaf818add53362155aad885a759b22220310d21862bc4e774cadd315
z85d57a2e2467688474f0ce1aec3b05537783e66d31da0d01d4a614db1bc70a0af1a013b1e519d9
z2bb3d231cf9f66730ba953041d323d4e68a5f88c75145153165514a5e90e316638db0bfc6321d8
za4a2ca0ee681c0eb6053b1f5bfb07aa76670a9e023e68709c3a4e084da4a6374869c8548cd9514
za94da160870fa15bbb75f75484918b4b893946060da14c13c13bd0600014278532cd9723a9c808
zd590f0d9a2d4628663064160b3b2d6f00265ac25d47eb1ead6ddad53b2bc8eb781dae5605b8e91
z036e014eb5d895d6b52f67db8df625cdcfc510f9a19048f394edb9e88630cd4c3c07d546bbbe90
zd96d07de7c5d594e5e8882d446901e1a94eb8c742303a100be8c5eb0f68b329cb9d13baebe4eb8
z5db34f9bd0817aa852b19e55c819246cfe6bc76f67e23f03073da0831a30b2b3f539111e09aae2
zde9434aea477a2ee17b6de7c1bf406e583b9d3719f55fabd68b211dfee888a9c311e0b80f97ca0
zbdb9f9cc3054b0271e4883f2779a8f97639853dd1f9fbfbd5187d655f10fac29a0f72091f3aec8
z8ebbda35f5ace96a12db426518104c9156156c385ca9d3fe7a93f45eeacee5ed8be04bec34c2ba
za7f77163444942e35e09385bcf227b028c08cde68303392d474e25244d091fbe65e00bcfaa258d
ze40d0ab0eb799a2287638dfbaf8bca6c961152dffbc611596c3458f5ced1893ae4360aeb030b53
z01b46c0cd9a314e231e42e455a7b49a0a05b1d4b5198019afb932008cf206fe69e50159316c1d7
z93c0b68da91dc7dbc75a171d11eb4321a2f70adf709e7cb6761767799f76b725052360bb8c28bd
z18591514a98b53e98f509058a8ee8cebaf1a7d5805d01bf786f015210919bdc32e2ca55ea49fe7
z5a521c56ce8abb2021e096b4834190348233b4edf4edd0fa21d02c4904cfd8f6a7fca16f784831
zb0d8527d203271475ea9dc80afa936a3d5127b8222960c367bece0c6139708f6f4585125c62e70
zff368fd8400f0813309b89f6a618e4f94366fb55345946483346d909b20774cb8e04a4dee88c98
zf1a33d46eecdac32811f39c94185a5d3f6ad6c4dd25fc55c4ef79f64c3c6e9b1cb64f3e32bc1fa
z0d8d483a756f1aa2b4695e26eb3b1e5b161b1699832cf9cb7339bc69ebdc29f5f27bad23d128e0
z19ceda397330c0f483be504e09a64136497031b1215209935eb8153c4aedc7a8e08489a06afd48
zad37904f9b488d56bbf570a14b0414e79341d7f36d494715f63d47cecf6f18ff114b3e410893b7
zd4ad76be5133e961adda2333258c27f3b0bcfd261af40d75c80080af2c969276f72eaaab6424ee
zd8d9392e7212d68657e51907af1a5ff91b83f7081362842060111095744c9eaa76b14f6de5110f
z305cac7c7c954025fdbc7e704f19de48ee0fcb5045ae1535dbf3333fb5ef7355dfe7bf6930986e
z712493f62f186bc7f92f6b728ea49343f170ed78f0b60b40abf01ccfe4cef315d65822f4dab8a3
zf1d21f1223ceeb68c221010c2a131b06671775a1df9511cd89cc8158c6f3a3313a803cda59e0a0
ze4a3fae231f3daaba30106a55cced47146010e3fc42f4f3a74bba82f6828083be59ccc1e5518d6
z7868758e63fc86d678b3fe9c76b29280c3ed6a2f64821cdc25d683547883962cc9d29c6ccad05f
z64e6113f6f394ccc4189fd2b064dfdb095219bead02b74cafeff387be57cb17a94023ab3101719
zfb1b907ec56377383d052c872ee19949baf88c4175f2504edf3ddb9395f350cbb3bc025bafc44c
z4a801da4a686d5a7d8bf0e42a00bd632274e55edee8e15729d6357ad3dd7a80273902d5296c63c
z574aa6d7b51ba382b086e145ce8fd4a31cf02ff859c2736e20b4840dd5ccb0a11e66bdbda73f91
z524391dcd983cb405d24f1eb7dec72f7ef0c48b7dd2b35665fa5c3421c22a07e127d260fad689f
zfbc4e2fb44305e74b61fd10b87bc2ca4212093a31cc3ae9129b449254b90cba5dea73bc325a241
z37678abcd6afc95b6129f31e619a1824b432453cbf5013b875488f62a27f765408256c7d620a3b
z5538a1ddfb78334620c554608527fadfd3d5586f3f79724a0a64a5db32ebba05b47b7fecf7a45e
zeea1480e773ec9da11ab9586b3424b1fa90f7c919cde454b8b6e047660067753d996e6e95eb8f8
zed5ff8e4a63b0b72acc0f89831f5e08ad76b7ec8680881cbd3676e9f5a9734c1c90dbde0b4cc29
z431a0ce848943bd5b4d43e8566392cef03c59ee17c636cb9418b2dad413cff7d2d6255711e6b79
z85e34a8c90dcdbd251b4d0f1966e4fdd3a3258503d0a91188aa0a3d43904e5efb2d1b49d0eda24
z79fe284b6f93e36daf195905c5ebbf3f8e9994a51b14caf88e3b86ff3dc487eda6004e029ef49e
z21c641ea799d923899063b2ec1420a8ad06c953a3736238817da9c60efc9e23da9c064645765c3
za2cd09e1f1d557062ce8f7e60afe8562da23d348a6ed9bb6c5f533a0753a11ac3778d2006ca8ab
z796ceb0850816e1a34e1698f481571bae38beba885dd1a21b193ff640eca3c8acb9d6cf15a67c6
z4f6d7325c04e8318cb100dd70f0219476901b3e905992b80b6e2166866ba9c108b9f59da51ab88
z7d9e36ffcb2fffd9bfcad40ffda3f570b511c25cd289ab5f6d4beb6c01f0c2eeac892dd8a0083f
zdb410db4aeefec7e7169f0c7e47dd4034a6991ad65330bb85ce4caf0f04c2075e95e199ee3c250
zd9e7a9ea77ba8e7267853584a2e7b1dd952b705bb64fef5a4b6a40b68241559c39c27213494826
z425d3a699bd6cf5ee93c34174690527210ea37467b43a9883d6680b419e912fec62ad77fca2940
ze68f0d67dfae508334426e00b8c2474bc44b4b77483551bb55549853cf8d14ba28dbb5d65faa23
z5769203e4defe94e6c074902d027d78b3d3fe992cf480f22318aba8dffe720e66273a13054ac56
z99253a54d087fb42ff4f8905cb852178d43d9453c041a72ae7e838a6e9a854e3129ba8a727ddc2
zeb2a113d7ffdd3783fc0f40e5ada1382383a6283e933c9587de03698ae02efa2ced9f87d3185e5
z68655133d4a16bfd522a72c676231d76c28d71c7a3705fb90fc1d2361b88097c104401790b01e1
zb1a1d4fc1e2df9e68442f416712840cc699cd1b9d664b7e38ab184212eaafc64091f8959e520f3
z5b648cea6da1771a67c806a51b0d5ef86ad5116cd2d66d7e1f2a433af6da5ee2bdb5b5de41243b
z57fcf29768ee742415881d1b3c333d12ab10a888d7e41eb79d05dcd1082ba04162a49b1301a277
z433180b6500fa5e39d452971105f6dea0f9770c7a07fa020b7b98f8299da16ce396b2896559f42
zdc9c060f55b27536aa8fd1b157aeb5cf734a2fd3dbf34b840618673861583b98c953dacdd6fa70
z94a81b9b86ec962de35a801b2e870fe80817b6f1b7364fc8a60da563b3da1f0b3176de24f437e0
z1294e009602bfddc4ab713182309216d0ac6d5dfb1dba74355a5a919f6f07431530cb85a86ed3c
z09763f3d8f8370caf49eaa390dc0577a3970c036ee4cd9f3240e65e744bdb7f7c3bbc7eb1fb31c
zdf339b40d6eb4ab0ae0b021233cd61ebe1ba9054a197a08aaeafbf5e578121e527bb75369be3d1
z23616781d1612aa39d0b28115625de8150874237427af091c000cb2974db185237d86bc7d2bd44
z146a9e37103de4d3e3acf7a39eb0b45036718ab88d7c26670666b1534830a2037c24617da32fbe
zd682df0f8a4273b77f2574983a8b5f188816bf0ec08a1992f913ae5baca3d193de8908f83cea71
zb0624d0118799b2c15219bcd4006864a8221ba9bc416fc1e81ddae6405121b8ba4de7f5f3c7034
z5efad6ff4fffb712bcd4a8a0ca6894e51cfc593ef099cee405c347821f02361d241637917520b2
z3680438ad3b59faedaae87aa4b474c980d14a417b93a7fde27926ed795c64436b1b1274024899a
zca13d6f4322bdd0e751045ece6ac86b16a575d8c4181be6fd277e10206fb77fd51f522e9a675f0
z3a12715fd5a8bb16391afa272f019e57f3abc2716ed52556a68f22aa3e62aa13b83c88015fc3d8
zf46477c92a28dbf22f6c20d4bbd99b0e73a458ba0e89ea12df9d4a89c1002dee19a94b1d463fa5
z7b31515c31ddc73965b32664957a4f5e4d32de44cdb33723aef622fd3ca8138cbf246a82198adb
zf5d83a11320fcaad11b3be6f1a05bf2fcb11a179db3c1dd23999212eaad301a243176fd6e538dc
za1863641d761c3d5930b540442040d99e7dd111c64a82472479415cc3a53d6267fb3293429bbd4
z5a8c916ee756ca2b0421d450fb80efc88cdd0a338077b9b775fe8b2c9b261aa8817a5b958452a2
zff2033e9f64a830d82a9ed59980ae65e855fdc7af592ed687ddf91da7f09548ece99f2f841d2e2
z381ac69398be8327de2a0d03808c4884281ddc2fa303851da1b32663c53d2598ab131f619e27f3
zb9332908a69b4f745c5f69bfa3edf6aa76817fea3f1fbeef17547728a88fcce2436d2ca5a5988e
z0518d3dbabe3ddcc4d224ea7a9996e12bf43bc44697cdab03a2764a50db65b95cf6abb4e5a0bf9
z4a2e32e9750603e0c0e42063a82b412eab4a65b04a34905c114017209f8d6a596f8b95bc913da7
zaf0952735d699120f1cc56bcb6392f41d79572f15c38ae639ca257ad11bd258a743f6c9057fe30
z6196e030ee4beabe3703a2b78354990d964f6e27353163f8602a56bd8cf566221d59ee34fd8c98
z5c0db4afe2776d2c362c420cfa32b38cdbe71c93a98306d784d6d1015c329fed7a5e98930d34f2
zec2314a304911ab7c350ebbcb339d8b5f045885b0871595aac957a331efa5f3ad3cdfd10e082b4
z84b6f9bb38c2bb523fc4ee2e2fcf5ca36da1f418dd88c68e9bc634975604a6c1c1c0787301e79a
zd5c6ac24d1cabcc5617539f4c2f8f266b9b603f859a3f743d2f55cea69bb6e5663f3acb77140d5
z17a5d8c908e6588599793917db752a5c009e068765c2116a4f3a54a0fc75bbce45de63e8c788e1
ze24e1a4d858da726bae7b24d632378986516c7f5e528cf08285bb1d733747a3db85fffe5b84079
z2499cc631e6c0f8f38c01558f05a941cfcdb4a616e5e78ee23ef25fa511715494a9d39658bc0a6
z0066c28615658e0cc4d1e81640d8895b200d2da9e08fe62b8ce2055d9de68f979247fdc478e49e
zc56b84bf5c1f0df5b7a4ba15937a041c1c1db4ba2b0e20140da52750a7276e7bbe7d342f035444
z3a3ccbeb44a58b14e44b4e3b440394b8335aca0d1798d95fc78651c795b1096ea9f1a3e3caf37c
z9c3b8e1ce94f92fe9f454c408899aa7471f0e8973bd678bc1f9c191bfeb07d8c6b00724219d149
z68367bdb3dd1821e5f688d95eab3779faa26d8b8e56b13414108fa4a25d4cbfdb3646f28f4063b
zc2715fb82325ee01bee069180c38f013df80d1e928c7a2d674bb58da189c43243318ee6dee1387
zf0b420428af8222f131f0e9256337c2b0d13b35c96f336c5da122fa1890bd3e36f2dca05aea253
z4c9ac78993c39ab7adbf5e034c1649b4bc3212a4f8c0e75bf35a961f9cd99dd5ca4a6a2cf8ff97
z9650d87027e33253d400db5ffb6d41891bdbfa37362172a454bf333726da2c98ddc0547fbd185b
z676470b427db9089ad7936c3117992b91820b218fe96007b5fd76b7109df27a1d97252e1565460
z83d5fdb92ad7c51fc09c4409d242bbdd27cb92c81e47b12ed22904c689fd5b469f80ed140ba2cc
za92b8e7fe88b8f3bc93c566547abe309550ffd0175e109550e7ee9c836d8ac6525fcec3b2891d7
z94f4d345fae1930321989d2e6a363fe6ea4323f2a7dbafac1b5592e9dfeb9ca074b86545b21144
z50b987fdff5d9a7127e808be185b9ff8855fa9f37ac5b5112d1b0ad6fb47d1fc445beca1544d09
ze88814b0d32fa30e765612381e44bee0da6a2ec5cbd5eacd46ee01f6716b5608e9759cc84562b5
z9d8e7fb33959dbc5e436e3e6d33a68c85bcbca987896871e2b495c5343d2c62d19834ecd13667e
z1c3b406b9e187b692f459de9271e229516d8c79fd124e9b263bdd1b8cdff0dcf665a73fa236e0a
z114c6bb9af5dd0db0569db0b8d224aba291d560bb873af6b0279183106e11ae1aa9f8ba7b78f4a
z4b184e0874b9a2e89661e32e42faa48e4e28af4b80c0ecc13d8a419a6ddcb77d14718612848040
zf7460d57db8ab931b00c07be34f7a9607737a4b07595912a039bf83600af884901c66c7e38235b
z5484b979af02055c193b5320d8c6d147a59fb1f2ef65d02d31d95736d5b7569a2f3a8da2f7568a
z8de1b474307fbded91400987a03c3d45602feab18a90b281ed9ec48589d0a51f53fc4695bed4ae
z388abdeaf62af9dcfef4932315d474f35f4b2f4ba9fc2757cc8e40a1f287672e5b4d9e2b6690b9
z1d65d0ad6732b847ba308e809c7025a76c05b7c4ddb3b7d9dd78be761edbf6b808bd8067eaf620
zab62cd5bc9134ab935177983101b02651b8ce23eb6024580bf2965ef86f4717e7cce9f1d701f57
z6cf118af195c5ea1432adaf8f7db5507242688346c3602b86dded40f309b0ba32617c8ac45c57a
zf19f6d14a5e9e97a2ec477d74189ff98b94ef8aa072db0500c0b20b570bd9bb2bc21a5e39d4bd8
zb3f3ac0f124f3f7d7ee92f70ae5507675e7a8764a87e1fa787d44af89f18ad50f745e7bb708414
z7dd7f98110023eaf65ffbfcc957e3e69a50b1eac35d299299594ab358ba57908016a5eb268c7ed
z387c1d7e81d133521ed7cec737977215b78546e48ed7f0e2b5c294f04a852837d015bd1280b0db
z428227c673c951cdc786631e7fb25f00a5a25c3a7ad86fe94b725731410807671aea0ec60665c0
z979924e471154aacd032e6d019a0f024b5c6a6b51ae9f70d2147a4b71f017454b67b541d38dfce
zd240ee8de1f0e6f585680629d332dcc455fe0434e2eb05858199ab2a55702325d76b1656ad3f15
z43a48f9d9c35ffac516e38163d7b9618e4b62911cf31ba575e8580bc62f6fac1f1e02d47373006
z227f0e665be395686975210d1274f1a8f889681873c93c18a2db28e18f46f34bc3ebaed3dcc9e5
zc56e7c3dd3e97e55dc7dfedbedbfeb0f8a8c3d1c83aad25abd3f3d1159769c5d85081f335a27de
z849b56b2199b6e1dcc413e47af20e82018f18f7391630e3022698aced3973849628ebc1f91a6a0
z81e1b230cdae32b4358c7d188e288d918e7fd3d94cd50ba27a50726f2258586408d7beeeba42c9
z63938fb42fd37479df467b45e91b34d082d1b8d58b84f1d2dbdb9e4c15878e8d3b06b56f39291d
ze7734bf5afafb10f0e8e1ae2a3f0a22065f7717fc98ccf360a0fc4d1d6633888c145f2222e4b89
z6f7da98ac63a1f89044de2f4b3926bdd4f0aafa59cb42358e5a59c89c5aefc1745e2380b6d8574
z644ae843c6f9be0177fb3eb8374d908ade25b0685b9fffe8bffd8d860997675ea19c8536209f2e
zefc13422e6f8235f36ce6ad0d9ea4571af064444971f1836f7db9dadb1ce02769a70776dc59858
za8ab30224ede3e4ada72e43ffa63849284195b95110c69b615efacda6bf8aded529d8a2ab4a9c4
z6bd76e4fd1ee402fd848b34938b168a300ce6729020f123b2dbc43739b0412b145d779063417fe
z8e5c177b3baeb7dc05982a6c8114291b1f51cacea16d04931b1090fb92ef5835a035936892f6d9
z659f6006e1564b171c78c217abfa6e46bf4d01aa7bac8e7adbcdb93d0599baf8d297adc7ab5886
z0f7560a790a64e9a50ce5943c08548d0218d6da0e2c7207a1035624d2ec5b056019b72dc1804ca
z7da36b3d6991df00a7bd7644308dedff2426e562e9dd8acd739ab9476a9509708fb231b73f9db5
z6e7720033ba358054e83c7e037bc0d84d3d3452ca1fe05f1846024938ad75f804f1694cb9be8de
z20395116e3b0fd53ed5cb6bc7d40622269e3f0c7c19be36c9ee8a7c28c9adec4a9f9d40696e46e
z1422e2bf2a9019df99cc35386c5bb4918c31c204e51a678494c53e6fa892a832a8fda3cf8e9111
z2e71800c1a11465313e11989bf2a34dbec13880367bd0fa6ce379fbc5739a81a2164cce0258fd4
z8dc20037764683eaa8f769613d625c337ddfd41f8ac065ac71e51f7d3f99164cd9168ea3765459
zd8059b4473b2cd765906141de86a434762f343f830fa5aa26423d43ae8a86a0661e1d4a8600514
zc7917c251c0d7db53a82bb7de9bbb83c857c10f34144cdf0f6fbe2cafc1fae71e399dfa11304fc
zf9f58b83f25997c3a6b50930468bce80b02b92c0ae034a6e9ff9f16b79f805473363d12c2b92da
z9238f8a86331b28b6b601153cef8f4a19aab4013391a78b92fac43b4337e3ea03c580811f36b84
za38072e53898c94d2a034b6adab55d161ff1e5c76b1abfc477b055fe8032caa37b42ee3bcec42e
z7da0ea2c8f8fd8bdc611d4c280754bbfc4b01271e670e2df689af9398332e99c94950a90276f05
z23f8e261fa79de8b775a40c68dc3d81f6771d1b8edd2dfb4a49f3f8ca57d9c90acc74b92ea7b50
z113d1b98665fa5218d3eb4943d4b4377ba0cf2c16b72540e1cfec73e25f963054c0129e7f23cd3
z13c318ea254fe1e2ca862e0a8084ed3762baaf2f036f0b4059fc5f4686871f57d40a7931a19009
z2e6ad71a6e5a96ee7f722008e8494b59eeaae3e44ef7918c677def598175b3357d3802c034c5de
z0e1dad23903ff2a4c05f7a7f46ddc1740127645080a81aa5cbf9e8e95c537b0d8a9d088e8800b6
z247aff8ff1834f4e119cd8a6e85b2d55732ec05c9781582a39c90da24395f008e1647adc1f1f17
zdfa9098f0b9d22b5b97f34b6296c57c449b9b84681af35526d587d49295fb2eb141b6399858d6c
z7b3e71743c546651d07160861abdd1c5c739f379a7334c5beabd53914ac6d4cb01196fd8e72ada
zcf84d17141a5309fdf6df45404852aef4e7caee7bb6a35e84a72dee71547c7180029f6b951adac
z641961067dd2c255785cfe3a51f8a7648ded908edbbe3fc5e3e0545be3f151090e136f55ef9e15
z1b10b14da83877b8b909c90f36ad51fdef269f6e2cdb6bef3b7b2e4351f3b19075c16bfcfb8180
z67974fd424094ba050aadd27a14751d3424f714b138fff687f8f3b805aeb6c029a413dda8675dd
z8380ad502c30b41b13e943e1ce0aa71bcc8e909670baa7c42e7300ed152f040dd6121ef6f4b260
za970a5db71632485c5a89cd76981d53e599d21b593deeccc6b4a6384b4b56bfdeb71a691477fd0
z4ba6bfbf7db61bf09b031fd8b34afce63bdf64b3a83b6cee38f4d0a5c770937026400466fcfc67
za37051b71d836ddbe3a59fba4f3da90f2cc450b7498b1f8e357ae7468d4131b712b62019d0c825
z334384bc2649d45dd1691d7d57e3abb1df178b39b9245cfd77bdf65a5b680266a557c683b794ab
z97d9abfca90dec914fd84caafacd5bf15df908daf5f6671dbcaf224fb4da4dba1c8663f228009f
z583ece654b91d15735cb2912b19b82e2e4df1b58b2c6e3e5c52ec5905d3e1ac7bb39b87fae855b
z176f0f587e118075aeb80716f8a1da16727f5d01525bdde1d7d827b0fd447f4a69d3d3ea2e3ff7
z8a72d295922bb554b398d02f8dedb526dd3793992e0142a3724de5fe9bb0c305164a653828db3d
z511b02b1d2285adc0e2f1d07225bda0b29e7c75b448634d195357af74a18f2e0ba904bcc56bd81
zd4ad153ad943286113cfd0432296fd824b9359da05fefce95de259e54accb8dbdc9c9e59808022
zd593652854ae61a4b622a6bc874317a8da8e85a4575a303ddb7bf1010cbeaa216a21c208dfff5f
zd5082989045aa4392f1129b151442b3801c4fa52f6eb76c8f4ed3b901aca4bd87f3804a552fad1
z2da95f7f50b84ebde64c1c5865447a2f35c8ed70b16a13a2c20456b015f3191538577e000a9618
z3161d37a6f7b3658b1de1d7e960339d50146a34229a3fa4fa7521b155d5cb188d5848ebd8c4c0d
z497a3f0324f85fa7a80bf338a576c98289a50af21ec0e3ca9ddc285e7899d0fef948956fcf3e8b
z4f00577ce92ca28093c300818a05915f14aa6cea2cc182595e5d07d17c7c553d22eda1599e411e
z0e4800c11b8167ec1e060915e55db5236a97cf6e35894119f73e74ce865aebf953cfa982cc1623
z4e47bdca986b91cbe403b0656b62d436fb0dd1f7a6b27e86feb4aeb31933c6bf256b6dea957be4
zcf27547987c17901bf64c0b01fbf4cdfe2378d44d50711757e1703da8d1233c1de4fe8de1b2396
zc4bde567cb0c6f54f1ee220fec896193bc01d6e8c22811c42526b8cad61b81adc8ad38ea3a46b9
zb71d50fb03262c72e1c317874cb99acae663b0953c8ada880db75bd5a3c2c54027ca955d99bfd5
z36bda99b26d8111d94579e10ed0d8b3c7663f28fa1e4e497e37c5cfec8058e641796212606c17c
z221425171073a3db4d9086f35ea01f515e2a7efb722ff91579d7688b5e83854a44617636d12e79
z0395c4e54dd26254444be93ec63913b3724846617e58ab606c17e6970ce2da87a0863850587811
z68963cc0b52cebcc514cb8a719f747ab02d1c63ebef92c277dbe3cd6a6dd111fb0aabc7d65d833
za148cf39259417fc4351e0d184693a8188e58df2e428d36f394177386066f65959b77603fc8a1d
ze643ded78d90625823b11ae4d335599474bb0797f39b4fe6087e250de0c4f7c916800a1fdea74b
z5473afb6ac568ad5724ca0181a21bb6c8d6046b2494d8d3b5f04d4a42669929a089940bdc66027
zea3add593f7c278fb0f5d8592dc2749c26a79393e1060b12f4e548ae38705d6e409fad0c029bbe
z6b8ba1cee89d6dde789ce3148eae8e8cd03277753618b7992c94261db7b4a9b66e5458c6a8ec0d
zd3b5884042141449c0fc726d944b95e57c4544fb3b783fcd356fa5e2bddc0ec4819650729bc843
z09cd35e08b161332d9547e8bd216ed74112892520c09498159245c4e90aeaeac8284732344eb13
z2764a8c98372834c879edfa1a427f0c20cdfd7dd8a862bd1305b9cf5c775dbebf7b8707aeff5ac
z235f472b794ac99a5127c4cfc7968d74c0c3d83f14e5b9243d2a62889140c43fb1d3f024e0be96
z0ce1ce542f498b18e8509a33d64e9b02f27ecf12056540f5482824bb606b8179ab56a7d6f33d89
z3d11015c6dc2230defc9094f7e80277357b69ed1764beeb0da7041f99cc6296f6e9c0140694c2f
z16704cd80cde36163b5702b995f643237f938a2ced60183e1911ff9060c735c57cba76ed6a7f61
zad00897c1cb2968ea626c8ce1c032b827cec315be9ddaaf8d79df2d2f8576f76ca0e5139bd1a70
z6722f50b6aff4384a65b88eecb0555443c2101cb2efa4778541b50e17ba37d206bf03fe29c4fae
z57aaf65a716fb267d9149d6353be994e245ce6a8d8aac519baaee4283ff8d608a9084cefa452d6
z67d52792103709604f1096111ce027ffb5fef742b02801f4268f5e386b60387943d0c2c15996d9
z25a6124c4ef452aa89c995c33c2662e757ec75f339674b2410bfee6ae839851a85aebd3520260c
z808fbfe6036f7f91d1fc7d8fe5d0776512efc232b9274509c57c63f56075c908970815d32a37ad
z3af016ef420bca844e665c2516933f7c0e6d3c690ff08d54f87c0c0e2e61fdd1c188bb5b447000
z88d6235909d1d8587b0531e1405a032141f2be8659a0ee915d3043448c24560e50c74c8deecfa3
z3247342d91b07316657832c8eb0e862e0a28e58baad8b457961ad989d67b90d24a7fae00181ef1
z12b8e80b732af9999ccfacf5127d1545ddad541b2f836a488e63d665fdbb1ecf7b360e9a6308ae
z6c689794dd88e5609274eff0847007e9288a4d887da9edfca979980a43630435b13172bd61557d
z2aed88c7f93e62b11ab538ff572e9ae98a995660daebb44a18b3ae40b1972f3c65e754ac805870
z4f96cc1b3246e8551d79a16df46b84c6c37ad062954b0d0fc0748d0b6027fb6fd168b7c876cfcf
z1ebf2ea192d3e1558396cc4545961c65f385436f1b59946d517e458965e27946ccb8a5902f909d
z41577346bb1a2888f5a4d46590444f3a13e29045d05970bd011b06927c681e8358d606a5dd2698
z020f0d6b0519bd85d9a9c5752acb0b6d689ae8df860a3b1b15ec34229ab7faa4ebb5623707446f
zea343a8369c537da871d1d04a33d83e6f06b9843cceb61d0d91511f3f8468fdbeb8871489ba34d
zb49ca30f983f7603642025fa0436661bd8b61c3e51ea3c11c773e227a7175fb17be774a98a44e3
zc9c1e06acff8ce78a742a7f92dc50bc0e74f50629e6b037ea76ce07b8cfb2078450f8c9e9d6535
zc0ce1bf171565cc097baf4ea10129a936770a169554fcab0baa67e2897526d5956c4f983b2c394
z5ff523326cc4a0d2a8b611b6781f7722ba66fc75aaa6f1e2e0837f45360c6f24cf9fdd142bbf20
zf32f8a55cb2ef70d3fe4b1f38abbcac0ec4d667310f3fe73452cb9016f5d0df62e97275e2e3bc3
z84df9dcf40217c0f34ead308e706e5c6bc96418f0bc251564332ea9b27cdeed3ba10425c216a8f
z71ce489a2ebeb6de1f34d2a685a3b9aba5ff23572c891bd14623ca0ee3689f9847f7531c8cb286
z5fce5d26a94757a4a087211c6b75a467a3a4b7398832cb8e8a455f98f00494d8aba28b97eefd15
zebab85f3b1dbcf3a6f2cfd6e4e4fead033cca7d108f1dd345ac6e99556e1aea58a46e80fd1f9a4
z8d27009632b8cc0e88b09610123bb9e5c2dd7c44f7d31730ba99d39ea02024e213a9c53e0e9aa2
z694a4bbbc519f27cb2198adcf48d9bc9720cf54023377059bdb046b6e759580d4a3266598ba335
z5744e83baeba3e82744c54cd85e80ac0dacc2d3eeb5ede3d9006d877ce1950d9f8299f070aca85
zc1c5830a4e94858cf2cff3ea252915696feeeb97416052f0a96557f84212f797ac89a30fc4efd7
z680ba5b82ce21bd2e4c55b55f002a68e7acced54c679183763216c80f3830e36fb1ed244edc1a0
ze32b8b4feb93979b631f882156b4bbf1c5f8db4275de8ff98a33c512a7e365ed9afab473553075
zb7750632b43024c40997328f680332dd0271e05b1aa2ee97d0b804fa817d0e45c2ff5c6df26e69
z311daaac9ded4473e39b648cda6d1c28bcc533f4b696fb0c79c0e3bb554544dc33e0f0dcd326c2
z85fbf26fef6ccb32099691854766cdc3e2cb7a3250eacdbac4da847330e6a986c672257eed2588
z9d58ac0d6e189f15cab1b02498d2c8e188dee1e96ff57307d0356198fd4f449f4d40aa87a06ad5
z110623bc93410d9d21e532159b0309b6cf71ac9a52039726648736395661c4c5699b3eab595607
z7c79208f02cc75235306be668553a7dfdc380958478dae8a8f325ba3560a7be03311b017931d89
z162cd3a138bcde6950ee145f5196ec020c50b8712ea48793de64747c609505a95155d72c415fa9
zecc5b7cdf38fce7d9387a25aea91362f3b47b361a0ac7855f7ff998d2af4f1c95df62f574e21a9
zf104b741cd15f8125e21f6bd7674a260eb7872f375dbbbd1a0396a38711ed1f7d6bc4a27806931
zae43c59bb9052a6f4819e1719e166bf51fe6d9ffa7c5829e5b4980d8cd336998d4151e5e95293f
z1528278863905add7c639e67cbaf1be7d375f7db34a76c559b796576a2207a2eada1483d78f1ad
z5279bc9e6c70eef2766b48d6a77f8a94ebe5979b886149bf7551234274c007e03ecd8acc8e61ba
zaa4109896c81caef56748d3b70e76e6e9f3606b7defce8e0e679fa144147bd30510951e6c8edcb
z787a13add10f769ccf3a2da8fcde25d6aef0c28b3cc980f63bd7967332db896df86aa9337a4d7e
z15dc5137e8a4ff01129672b69d8f5adc1374beb5e9c32b0340f24d7ba5c2191b5dc3020d736c5f
ze6770b2dd6fd44b9e76fd1af8495e218579766cdf7499889493424825153ba6ca0bbb0bedac086
ze8f52ebee6cb17561439eae22a417ce5783aa1cbb8a86015a4f77de018a3c7a51928a24a18d552
z35546c048fc395db30b925518b6d391f829d304de6144d4db1245afbb2e4ef0fe060165c9be23b
z80066ffd109b2ae23184c4ddc2206c6d8b9e91b96cb28f4394e8d8bfe8867e8acc724a624c7dc5
z42df0d700510dfca84d8be7992419b6801f1d9764d0524fac7850cf3a32fe9d17be34c31d07b42
z8cda4a2620989ccaa02e6f427994cdc71260842a76db45254cf8392678e67f8e836c765b47440b
z76df2a9f88959c5303120319d117e19c4ca223c85c9681e810dd5638e8b2e4c273a360d67b06d9
z1f02062672dd3f91ebdd5ce7c30239003abaf552142061d645b1698434db994358cdc37374adae
z5badccc3d69da67e7035a0fbafad81ea6b961f3e8d77bc0854367fb21a85a9445610a1ab3b37c5
za9f475ce0ffcb11a2f9bed6ff22d0480efa2cfb3e976cbf65d8e45a1ba1825fcd17e5ae5a28e1c
z4521995efa465ccac0295ab8479cf464f4d08b7caa38d12ab8805498a62aeab4031f6899292762
zc18649a215c63da1aa62845f8c14a798f84284bee906b26a38501ba088bb49a1a410af75e56451
z8b433f10c9d141d9ae42f438a62e552b610dc51e939fcadba033c400078e1be905bda056c191f0
zb87b78ffae0addf3baf52898551ff46594db53d93f2b4a58e03f855db60352a4a7d20aaae8b5ce
z1024fab49cd11fa3d6e67d99b7101faf97299d5301d7588ed92b324079c30a32c66bbb807de714
z402296e589da00ec0bebce8e5a6364fc7f350629047ea7987d05499d44ff1b89b494ec8d44834e
zd9dd3e15bc2d10726c288d9bcd95a7d298edd03641b44baa97b328be00c54191c1a9ca75f6b58a
zb0542e9c42d86cabda3274b143eb5ddb730bc4880a84db039aacd7a91c184df188875b428ba30c
z9e4f1a61da36665b2ce04305adcfbc850a325f201b24c9868a6d355a34c2a74f34d306b8f8e00d
zf54ba2f300a0442de0ceed92f758f236b147703107ccb9074372c7285a4011df393a8c9dc29b58
z14fbac7720be3968e2c1e91cdd0dcfe77205e4725c800ba17551b33d03d9411c5ea61c64f06e22
zde1f5bbc31ff3ebb6475f00b48605b2133ad9535f362dd863ac73ae50f1ba9ee3609ea3be4c254
z99fa64f6192e6ee25cbf6fac2e33d9577568a2e4a217fdd19371dcd18137846620372082488ff2
zccebb4db154dd4181ccda0a4d4e29cd470388efb16271a84f0f0029a13b78a52e47e3c106e6b94
z7e61377b31d131a46dac2252d323606bd6d29707683757f9ad5c88b6a18a00a49a60b0bf119161
z2721c03381ed0d7b6931f36a5daa191cc90d87c17b7340383b948931f27965ea3442005ecdcd20
z2a9aa5680ecf12ec42d884159edc52229cf5beb408e7b9ea97a14ba182c3c2c6a9e0643236d27d
z87dadc8399c3866726f75209a4c3c817872b14f3a2eeb3f3b803c50924dcc0d86b86e364657088
z73bbb3b69ec61d6b3f2b85155765f8ad8dcc225a55906db0a8ba2d9513e22b4a4acba01f12f9f9
zc4fc554cc3520735d481c2c0309b6d1c1ea30077420a3a870e644b905ec1b94d69bf94a353339b
z73f41fec30a1108ce11fc84fe1691cdf733ecd43266bf5a244f7a2d68cf3edae67c455998adf48
zc0a4fdc43f0ba68d85aa2b69d4f0537b6455999c583ebb16d79aae456cb59f212020fc643e9e1c
zb2a47885cd399bb7ffccf160f46f49171be12c3e169040238a2bb91681bfd7cc78cef6fedc74bb
z9e26f70d464b15b500667fb618f98accf1208082cc7347def9458cf8ba265596e11aa09f524a69
z20dcd8ea361269364d4ec06ff0bd5d0e828df7508cc352c1b7437fa2a64ea7314093a01d22e6d2
zc53e32da44d2ceacd4223df029e4ad9c5fb1527a1a9ad3dfb614dc07d6b11fac015d501b234523
zba353ff8803d41d587cc6a8a9502e51bc84f0c093fe80fbe8a3f4f7c4d6cdb781b07c5cdbb80e8
z0aca40ffc7e52c89c4f8c121aeff981cd4f60ec249f1d13791941146e7f60dba8670d390111b67
z8cfc79b2edaed17789c7b31abbd5f43fc6886e5e8e6342deb027525cb57b30696104233db64cc3
za7f1730a1c0055aa3915f84f23393cab64b17e5cd4bfd082b6ea5a467b45ef8423e7e4cf4b4ff8
za3697877b60e6cc27a4bb4b6122f5af2381a920f1ed456058bebebecff9af5589d8d14770df6b0
zdf9aee1d8d14392786741d1a623a2b0ed3426453ac0d20234f2a55818efa55b45276e815f5c21c
z2e268dce408cda0a878923eddf596bc727329350b9324786f42199279e85868cce8c733910929c
z3c1544ac582ce12ade23429c9e164ee83cb4d21b9879c27a68e73a5c20b9e8c0d293a53bbfda74
z6339792a7dd3e10d388c9974c3c3027a2c8cc2c8ea7fd3f6b8cb669cc219f01c0b81b11c08de35
z16b28b9abe96b92274c9d782d9ec376c36b9d113d7ae92083e11a23c88184aba154e2ecb8e2082
zba6fabe32120f5e50ba710272c2c0382d8108ff628e3312b22247b1a5257564fbf4ab0cf124df3
zd2b45f3342615af688cfdb104b308f5eb836879b93f9243e3481a27ebc2cdfb1f013ede58be3ed
z3663627448e324c5a3b936ff271239966f9cbd207c58784825718e9da14eb6b5cb70b598a17e6c
zf1c0bb1699c5eaf179d7cc91d4286e4b3d92d44d3e78e46e0eb0e5cf02712e05a98e266c78d2bd
z6b536fa70f09cd48d34e52c486d68c2ed3cc4f50ad59fee2fd44d0df34f1721ae46a90c759fdfd
za6de09b3ddd3ed37112608df0ca3109c77c5cfde17e61e1f60e80631acccb044b4049d0e3a38b0
zcc3e5c5ac5c29438d80a0578225583859b9bca6c4d0a16645e7ad670d00ad9cfd711178f7fd788
z4aef39f70c7c66066428ed75994055e155b81346ce16e9b7a39baaae51855d9c8b1e07429d3c12
zbebe7b4749ba055539902f958b3540d08fa934b2e9b5235c29c073dd08f99c0ae54715e13cc405
z36d0d0a512e3a4919fada255d7f8de08702e00e646309e8a2b462c49ec2f90967637d81964fbee
z2cef2c97f34110cdb5a76694310e3017365cd3c83e406298d85aec9b98388bf7577723d8a96ce6
zc7a3ab430321815ce1004d8b3cffafa62631c6911b3bbf9cffc00911eb7e1754aa928e66760bda
zab32db1033b2f7e1355ab05d1a5164ff54831723bdc330d87ad852861cc3959f4a47ddca147c91
z3a51f5db7cf896dc5a0fe5181c5e003772a5cb43b0461369c8d383521ec88d594a0990f098e7d1
z8871b19420be863dd17ef2387302c3417dec702ee4d8c933df238bfa5225dc50de3e4b94468c7b
z968c464c77bb678b0ec3265b99b45105186c1e894b9f295fa1a26b2aa2d28d48c501cdc66cb680
ze7432bd892a400ef6ba959c585e078e214bf0d63a179388d20977101f8d9b538e87b5fde4b4e13
z20ec647de1b8221540b2edd4a891565acc8000c7e29843170911f1a1a5b6822c631d0791abec7b
z732c0db3dae261cc6a4d05012d2a87ee2c93f54dfe4697419c31c77a38978fa2db1a835e6ed7e5
z7a54c2959db4926c9e5ce5d9f69177276870e1a2078bb2b3b4a2dcd5a8e306461b365f946cd8b2
z512920f152298f473dd15d694a80506f237a57e580b27669d5737a3fd323d798ee45595e4fd963
z2a252b2e849bd1a62f60aca6a4cbab804e716d6a11bc5e706cc6fd3dafb49bdafc29028850a578
zecb012f269482fc45d8e1d01b098deed01e0717992ac3c02539f05e924666f46f818ef05765da8
z2ca4763d2b0f85be6b6731b97279aadba1442a549dc6c2e9da5deb55f17a57d391e009f96ad7b0
zc3a79feb3c2f40cf857c022842c7fb5f5a676e4ba5bad9a7a4cc93410d88e0b4c1695e02104666
z3676c3cf2f23ef575d4dcea90375d1b93f38ba272437bb336f08296d143b1ad0302849960b0081
z931da3a7502934258d3c3dde3539e2cbb27ac6423b2376b57d4d2c1149e16633cee17f1b6a5510
z5028f2c4a7a0754d5387c0b566f4993c54964944269c2bfe0c63c840bedebd842523d2382cad7d
z3d1b1ce717f3638551c219946f840408597b74a32d84ce5c74895cab6d78539a6ef97f83df7160
z6d17fc9ea03321dd645abec1e34913dca859f15596f7d84c6114fc04dd2deaec05f2eb60af4b9a
z7280bb0d0b8bf9c26ea956b14e1dcb6e93e0d2218018dc79f6b03b30d9e18be58053f0c9802a9f
z54475ab3a24c364afb9ee3909a396c683978913c1c497d7ef3de4dfb7ce2fe1f01e951f9afcc43
zc29b8659f1246f626ded78616336f5c4fb88d5e6c516554054bad8a114d5d6090a7ca544da23d7
z85493d6fa8a129179e9c457455e27230535c9b768d38d5b02bff0220704192e9e2524bb5e82db6
z39322093e0fdab96c28a41b02705f08844beab9030d0ce08718c4b0323236dde016788d8be20d0
z8494fd2ed99533b5df4140f4289064d242d0adecc883aa3c034fdb2dcf32ff7b98ed9aa51c4821
zb5c2f04e15b2eb134f73f869e17cee4ccf2d09c8d2bfe79960b49253e2b3921154c91e44639c09
z08222e0eca4ec6a04dbf2830131e44eda6cc9f0a4aba12904d7ad12792559621036855862666e5
z2bf23e5d016cfe7e8f544f46010b5cb8eaeec1f7ffd8bfd40724fc7672ec102c130c31bb41f03d
ze3174b7f1e4dfa29b66656d8c3507fce61817ef9c5e8ef3757d7a0cda7531bf6a31dbbfa9ef957
z53bc3dcf60c199477fea4b3cc303d54bc9ee47fff36a2f25f6e74f8f48cc393d4b41a957f71ecb
z076dbc58fc560c38b047cfb3ddd51c0296a4256f657f7ef3b5c68da5938a7a065e446d2afc6fd5
z338f6b2acf1782fcc0d993b3d338f0f25f0be666bd2c2a5219c9bf3d0080f98afd6dcc0d14e4bb
zca3cd4aafb930800efbdc1f6df7c405cdd7d2b6a27f8672adba0eca72a4ee4b72d0306c657c09a
z0ae92ea1d0525c8a0953266f5672f2af7ff10c269918dc6aeddd53b2f88444caf58cb3cabb2f70
zd18c9b50ea23d152f69b650389c13ef7bf89a927536725f05a2e12f7ebf224f4e4211841d760e7
zae9da580e9476bbbe4ca76157df09c61827921d2412b8f507f175de05183f3bb3d137a9319777d
zee030a5769a339f062a097566aa6ecaac155faecf9beeb0195fd315300749173492071af42f790
zc90310efd07215d3b985c5a9d7209370de44e947c6129fcf5b442dcb47bec4f83443a5f094cede
z444af6c9e18a29316b06329591a72d150d0f07d7cdab61dacc5f18286875b980a3351da2c6c205
zc8af24512f4c0b9777170fca595d3339dc937a548b525ed510df1636f1235310bd454e485943d0
zd805dd38d341e197eaf3a8238e02adc273ddcef8aa63201460c5498fb44103402fc0cc173e537e
z14ddc86de841991884192277678e91eced98aea93acf6009443d44473b727a08a4a04cf5827073
z58bc993a9711b539eeaf12d365c300437c0167f3629ee392ae587ad40933bdf598ead0e4c51d03
zdc8ab19ebe3c3d8e8ae5f89c0010f7cb9c45b5d9135c7b086ef9b512688abb8810f6a9fb1af361
z456e456d71eec715ca514b88d366f896b0a704e8b75e065e4e50a95150934de583587ce6bf9dbc
z690f006bf5365f636486ecf87b59c57bc2d455bdabdfc7a55ce6301ec64089df2a7feaaf80b92f
z903583ca916df6512cabe5d96f40c2c8b2b2dd5b776bf304efb795c126f4d285ddb75ad2f9e175
z1efb98f3c8fb82eacbfc03008f59354cdb6274569382779338e23f508291e5cbdf84fd4c80baa1
z1669a1277b01151cc4cbec745adc66411ca25e3dc83e2ba5d8bae53a67445bd7536a33fc030919
z07e1c736e5f4df65978cbb2e6346eb4b7ae84251b51df55939706f838e0abe04db69b529f48f98
z2f701b3cb672a875cbe195e707970cdfb7ef50ee56fc53d1f9bdd6346601c6a622620eda0b55ad
z78f16d8b315d7d19b22c7f22bea0cefd502fcd637fec8c60563a904de40d8681d17ebf05c227d2
zedc22a0f40761d0a25bd1123f8b386613a8f245f092242d44739dfb95d4e46e56ffe3033d4ecd3
zf93017abf2fa58b517c62862a8a8c42ec348d019b8d1ac5d2c6b0484b2fd941f9b1cbe7e273543
z2df6482b21de45f15c2af9c46711a8fb5ab4645c2425670828a75d5addba2a2a179b92eddef3f8
z7b059a49df3c325b48368e4f969568c40443f85c0a806199a6dde4bc16e64d67111e1cf96ef753
za1e52989f16c667080139db75f28c68f6e7f278034378f631240623119dab29eee759a8bb28729
zed31cddc9f1826306282cfbf02f003e55b02b20a67bf28aeb513ca0423a2bada157b386a82c2d8
z6d2d554857cad18cadb406d185b9c67423b17724b04610e93b69bdb25973cef61159322d779e15
z402c768c53aa28286f52feb1b9e012e851cba257109cc897bcf59912e6e8962ffd96c0afdd176c
z18d3c3a64166d951adc3ef475c3ef8c8f68a083b6ca3691de1120613c4d94ceaf9f05bcdc42bb7
z00fb2de03de9a4e06ee022b5493d10e7a8f9f105f100c7aa4e826b7368cbe6c870f3ecc27cbfb1
ze88e879e745234070190de38fd4d5f036c30dd6632ba33f4bd6af4806924a752b388d9b347e478
z13de087e55ccb32874c29905843feff6ebfd91e1400284597112350e50ca238dab5c5a97e97adb
zbe3d94b0af58ea8bb2c680b265c75d7843b433e8abd0d92118ec5ea9ce1f7b1809c55ff39ed8cc
z02c96560a84f17851130f97cd473d8e5348deb750185f90b9429a564dc8be3331f4499ced60b1b
z74268c83f923f5db72b0933226880d3006354584cdc2c1a8e035a2feae25ad218cf0549f787e10
ze6c7c6087dfaaf7530ab6517d1b36cf025a5167100893cb0f2ffbf4116d58d7d3323cedf9b520e
ze5e4aab36769a70527dd34dd33ddbde114c08311159fe40caeab9c8b27941dd3d5be1d5b00bac4
z76ef06dd1319f77491025e0904b91c353ea3e0ace63b3a499ed4d8282e2191b6bdcf5cba038c6a
zc07a6ec6c1825416b167a6d2eb65fb769104141e9b69159f8596fca0b02eb4d26255eee7774f03
zcb22539a672ea3aeae9c9a7af367b1e02a8db30bf8908ac3f003f7af665754e66e826c9d804e15
ze4eedc17017caf64230ca9234cffc4000a5c588cacbf457fafe0db5fa58b7d22406dfcfcc5be34
z64cea4c8439574eec0314e581c0d77cf61692e6c95ebf222f4e6259ff6a78b173b637067ced4b0
z585130695a70b4eaeca480f72c22e14814c60f055e1a355b08c23031c91f12c514383a02ac9e92
zdfe138b2b5cbaf2b5cfe902e69ad486f7fff34e93c02a68c483155936ca48b6d41cf9600f48c12
z6fa002fcb0a42299309eb4490e88f8ea1755d2dd95570d1632ca3ea988c450eea6a261474743eb
ze7e5b615cadf741a0454a1723ffcacf117a3eba4e7029dd2a5ccd8516f384f82a277663107d434
z2a63d4d595eecdbc5da7667f603e19113f276c470e69162d43bf8a685ad37c235eec799ccb2dbb
z2a42808bc2a80a663007eae2ab6b34d9784991b9ab683d1f6f15d1a8293013238efceea2018f33
zc2f16f5546071945f15b196094c00d9c4c05aa8f3e22ea545a56817afef6a2158eb14573a997d8
zd10a83b098749b4fe4d630900dbad8538c662d25a6ce9e796d3a862e8a77c3861dab5d4a0b1c2f
z1ade0e80dd3ba1768e1058def5f553db86d64f8e81fc55ca10acb2c6f89efe8673b4fcd209b68c
z7f6e2ec02851e174a5ae4cb8c883f6c7d772a9b03df192c8f83b477f29fecd097a2436b6345235
za9adef722d09e6fedc5f1ba4375d60adb2f2c97a4d7e2dc98dbfbd9013ea5c6fba08168dad76e2
z9976c6ba90648dc27d1dd8a257f93d4ed1d7b689cb5ce976912cdef30d44c1c4a3bd8720de0e8d
zaf8c180c4183912e45f00ac91ea4ae792b8b84d45fd9579341005217053e7b227752c9ef80e5e3
zc60324f7eb413bee8bfbc6494bb9ef4276c9b5c4436a711aebf3171512036e37dca28f062b9ab2
z113af24ba7f4b67106f254f6239db538202a399033e67354fc4906df9fe7a1ad27d5cf9b0e4bd9
z8b68ea859796812a34a13666bc4ec7b257902fcb4d6614aec05634d017f7812610d3266dc5e3c3
z838cdf651fdca9a2d9f413e55e470e02c64424369fe0e50d38b5d749cb08932fa8093504cd69f5
z9eec73bc705c236fe55c415a81151385d51acc1496660f11f0564758c255ea0611aa2c23beebcb
ze6cdd7de15bd45bbd5d02cc6533c4af0ec624403360be3b527b0fa92b369cdc9245ee40f4bedcf
zcd9992833a005bf08c555b55e2234576bceb3a78f11873c2fe4221818b12b19fa6842bbfa2a908
z68e348d39fdd77ed03ea8894194c06eb855b2f929af0b99f677e5b4348e33256f1ff66c4205ade
z4cf8c80054c08461fa13e22580bf649781a44428e842e636e1cabfe1b58a97806dd53cea7b7c93
zbbbeaa1d50cfaeeb009429d6c975d4f546ef6e7f838e951a11c43e92a04056444fe96f4745bb39
z976fe4cbe32ed5eb2deb5e3bb1a23353d37dde6ab309629d5fa87a94010467927086b4558cbf2b
z962ecc6f872ad100de0952d21a395ff909a266a1591719cf99158c338ea7484a821efac4d2c22d
z9cf8ccbdffd540185e21b217e8be11de902be41ecdd23040c4c9930b8685bacc9ca6186404df30
zf29cf4ce21917788808dedaece2db7d279245df96150644f4e2b47b640db562d5f377f38325714
z6bb5eb0c4aa9d34b99b85d619543fb3c4f4773620c299c7d2ccfbf7dc565d2e6dbf819501e4830
zf755215a8fcb705888f6306e9379281dc2250e7bdaa35ca3622c2fd3167e12251ddf3b09c88a53
zc4fefc1b1a0e879aad713527141415ac9652637cb85e93fb163c932ffcccd3bc423cdf24d273eb
z48949691bc8338b83a6573494f3f1f564137be78162fceb8e8d0dfd734bcfb38af9014b64e1b23
z631f1f2c9d7f4638cd5bb81ecbb51458c55c1a1447b6c6168db2d74aaa87ef5f92899b6fe416fe
z7b24668341f47e375083b67055a789909a731f477ce1d6335c303ddef46fa92d201a3258e75e97
z3658bbfbf2f62f3f69e55d990ba1197b2000e98f201cd9d2e5b6b8bd4cc7bfdded7d2ec00aac9c
z914e7041755879f608dca630107663fd4ea03bfd6b3ad8660c2003f748c9baa6fed32abd395984
z2222681d34308be5f9280480026da6ff8cd5360b7b6cba1c16c2c2f79cde55bed9ff3061604a8c
z8a854807990e570b8a781054ef7f3ff6fb59d9b48a79526ab1898d9e4665ac9e31b334aa97fba8
zfb94a1078f31d6da7357c4be1f8db19a73d5331cf824ef7c242287ccff14b83d85931d2c1608c2
z762a5df6e678008b3cb6452d8f520cb930f0380df1548fd88010bca20482dd4539e7bb64fa8185
z2b003d0d9553cb9546fcfe40ac95fb8941adcde7ce6fb840aebd7f187bd927441ebc84fd2411d1
z1eacefc97cf80c29037c019dc573f3d1e158f7202736f758a97aa1c6fea4f0f77ec81881807d2f
zeeefab8eb946e35a6eb222340a219488d9c1931638e771100ef73b827a7432a6ff25b5f213dd27
z541dbb4e6a35dd8c95f6b985542feedb5ce5af1c89823d9c33c0e4afd3ca3213be69daa51e79cc
zdea2e410b15f90de92a2aa0581cb4022b15dfdb3f66b19211550300432f033857b980a347d53fa
zdc7b9c7f6bfd358ecae09178f5028cab493cdc7671304ffc1f82f28ea8833cbdf5292e90136a9f
zc5f73523be637da472c9a73efae769d71475ff6e48800524b4b434b35932254efaac7e58fdb298
z1245f6ea2a3c53a8854f3b1e0a28a37ccda91f4be75169a66f5648aa0231ec55d857dac0e68f67
z9fba2bbbcc2f27a3a2aa8689e281e144f98a2a44dc8e6d5b7bee40ffe35cfcd1a7bdf2beb69113
z8563c74301e57658c94e2f642d375d0b4d5ff9338dfb92c8ca3cd7400cb62d247047a88a687eac
z148c83f2649bb04281f78e91060f2ce75ea3f2bc9315c3cf06e2664300b9e884542f441b87a398
zdd5154587e1a4b1f6a86252e98556e2e1a68c4ee90b27a6aca2ccea5c52294a6ba5853d7460f0f
z00b9f68ef003e7c37368062af284ce3014f74d3cc22829044284662dfb6e4118c996c2d9be54ab
zfaf3a64b763d1f5a64c1985baeead416ab9f1aa392c7753034c40ec6e818b2f849e9872d1dcf08
z073e9c65d529d348f092b6f0e4754de4fd618cb8981cb5b173d1227e4b0ec1ccd60bc0e4f39f5e
z4ee886076564df56b750b4a7bd097c99630298668090304e4e8ccccc17ff9b0a0f4f9f47a19481
zd0c2c619633a93d6348293d69cd3ceb3447972215fb4d061046d680abce4e702dd43f61436564b
zc77a0098bec696b5ae4e58c34195c50a360397bd4f3fc5508910edca45edf6e8d92c376c77b295
zb39353357405566cd67d96a1471ec0cff827d073faa4ae2e46f9ccd5c43eef138922f861f685e9
zc077af186fb3b1d3fc654e6b5001674ef7ea9e5142460d2fc384d4c90b410d7bcf56fa1d3cb73f
zcb10352d5eaf846f1e7b1bc2ee3801adef1445a253101ce37ce9fab2059a935c2be30b7d984d09
z64b850fb474d60230e2e811c907324d9145e456248251881fb5a1f9d7080c208d44fb212f4b547
zf8cabe0068163966768d90700c23a4bd357d43c0ae36a00c697d88f1aef46263382466ebc2014f
zde6c28988fd642b3fe5d0761c83e710a84b0a82c602548b702a1a5fc57b43a162e70c078bf555e
z11b7937b203798c45f11c16808529063d440d784bf3d205d254b539974eadfde50210db317f2f4
z495d229ddd557fa8b0a8c7e7558d190e07c270fcb0c7ec707eaabf72b2fc772640bfd35b32ffae
zffd0a48119b863971226682408c395506d3d922995811f0488653ab11538e95cdde45e5a2add32
z7d2d72231ec15065570f828e81d1631121a57d16d49c8bdfd68624d793031b535f4f96a341dc8e
z3dc6283f39e727c16fceb0b97da025d6de9e7cc71742b4df279f16e8492f2f1e875112d2cdf052
zbbeb948aa41ee5a9f40fe9b788abed81327c8e9f5e76934c75a7830f5c926258c89412a681e8bb
z0418f73f415bff952ba4d8dba3693f0e9704cd703b1445ff17bc7abb9b45c0c8abaee20760995e
za1f37ebf0ea4586ad493422a4775da3f65b6a2741bbbc5142eb4acc5b2ceebbdd628fea1298ba0
z2e5dc5072337a2b00949a9b1eb444e20993c5f14273f9211fadab86b837497881db082297d998f
z281d25daa6b6bb064a0cd6d50e54ff888e45765375487ac4813114170a7f025203d97a4f4ed9e1
z35e451b6356570dc4a16327d85ca8e832983c58478e2de295e20a01df11521290176d5045a939c
z176e180e626d8b95483c6df1d9f0fcf296e5481db875d6875be96329a925f9cfc4790dd0d6cca6
za76544691cf89ffc08431d30ada8413d47d3300e87bf791a28f612e4522cd3600ed71cc8f7ab22
z7925b2e5204fbef7e56bcdbe531d6f6c9a056b2b66a8e02b67edd0b507258cdfc9f38c08b42bc7
z8bc1b762a4ebf5bbafb91d0d86d0d84c396e5f94d6ab168bd6b0399d99270edc1623c3b69c91e9
zcf7112440c276d7c29cbe007923a3308dd0ed3701c99f7c4519a929710fc03fd5d230d11e49e06
z919aa3646c7b844456b116f9d244798c89842ffe822b87ffd635e8f97c50ea868191c986936cdc
z5365b2a3ab42c361e2b416f424eb42bc464b7013b1f1f2f125ca5d8d8ac704ac71ebf64737542f
z28dd5f6e090adc68ca368364087a4ee259d1aa01ba6ff1bb3c0c02a64ede621708f0cda847fd7b
zf01f3017c4b261278200d20df8a09bc23953ad9ce5bb81473ce57d10a6213e34767ac128adf559
zb3ba57c406a5be36d4bdf1b5a46eafe5464c36f51fab44d7752e65ecbf101f14e48da4edbe6d2e
zc4a1daa43d77fc4c78afe3fe8577a99842fdd3ae7691f7bb8f2e1faf138cac033bf540b350531c
z26920368927922a5333139c64d0d816ff9a6534eabcfbe0983f5d0a5b11034eff2afca535a8600
z9de911c8430e65c54c1a3325891dd2554e19815499b6fea5fdc88ce6d666ece81cdeb26ed538d5
zc3b2f957317584213b3fdef5236f279b2cf3eba3ddc4d9ad5c9c25ed8ee8f61c1245ab3624316b
z7f2e8cb1e807a3480d5924e42fd10e0e42a9add251f87273e276f7b04a5c11eef6ee49a1598fb1
z6be9c424d2b996ba17eda59ca15531a01bf4bad985824454f43196795fa50ca9edf1539c651ac6
z3d5a2710848f76029b55c39ca3af415d34d49ec55339319824176b0ed9a8b3964c1d709ac59066
z922bedd1fd0e042558dc515876a2c8a9dcb45afe4b94a1f03fb69b42b6b1e82b31b22fe8a584a8
z6f6d44748b8bbb6c0f0925a67bf801d9f018a08453dd24eef49bd3aafdbbccecc356a05ce97a0a
zb09fd639b764ab1ac9be82ac7ce672c7e0254a4fd20d17d15e2374753b68f3adeb88365ac72d8c
z8052bb5a3687a94c7b43c54846f721b3bde96df09c3c439e9628e9552fefbf508a39ba09c2947c
z9ac32ee15c2e9ef6831d2ed2a77965cdaf03981f30dfcb269453ad98074838450746f0ac2d7b64
z7b44818ea80077c23ee02d42f42c88a30f17a1227e614684b482edac0537b22167412324d00564
z2c39eff75f18d76813cc1d9f8fcccb6abd89e9f2731d875aff43d888453180c0bc3b394778f96a
z3a0c5bd38095d31d1da58ff6a106a24e06d2684e656524bdd834c980e0fa4444b2c6e02191673d
z9cc030223a2001f2dd9feeb5e2766f5b9cc58ea4d2d7d8f4841f05c7de039d6704fcb7368d753b
z05aae2253e7259d5634e06ab9e46287cff41d6a3dae11cd1dc091d9121a46dd796c35615e12d18
za7128bd681fc3bd011d168c2e2a93916b82c1fb82d1cbeda6f370b391654500330e1f1595bd5a7
z94530c90ce4d52bc6925918c1d4a5de930745f6a9c93d03cb259a0a384e5ab99739b532b0a2e94
zac94f21de88cd5c49681a00cbea6169c0d126775ee95edeb23d74515cd8e17b4658abd990d04c2
z949dcef5636611400a79dbbe279c58db66380282bd28c2f22239b8ed2ecaa7ad11beadb2dd60cf
z58edf835349f8a70da381bcf7577ff368c2c011b54be0d8e1d94ab85fde5d24c13372a13583001
z6f08e1a413d5f870f772c90da2ab68cfc0b4402d643172a20b2c54b75ae0a002998b579667d591
zd6995dec1869443cc751fe5f9b8d63ce35136cba56e9e312bfa50f0dceb30ff7bcc9241ea25d72
zf10b74f78265b760764d58fb5f5b702490828849bd52150e4c9d9899ba1f05094696235cc1b6ea
z83f7bb3e33f7c18c8a21807c3f52b61f5eb3b311186623df2914067bd8e86fc0163b31baad509d
zc6bc0566db8acde78e95542b800b6d7b5f792ca24ef059ac8a2c803ea920542d95a95f0b5145cd
z05e3be722cab8e5e64e0f2ba7a92ab269a07ddbc3c95097373a6874b21cbd52b91a196345f462e
z2702093573ba60ed7daa8fd75c6536677f024382a0ab89425eb8fa38713729474c1d205749316c
z07ec957784da1ed954b72fda4febb619ea9d2728f33d5fd4096e11618183d0e859a644e9d5ab0b
zab282c98e59ff58dd3c62ee107a61be405500dd35ba734fb30565c6de52c961c396fd81fa2e2a3
zb35087a5e88859c3fcfce4272da4786e6eb7f802f4f3a094ace85f37d2dd1f89b66d3c36719e2b
zca4f17a294907869f13361c8ad68e44eaba74a491e14ac753ae33d92754a8ec0875a251ec9d755
z82340a90313b3ab4b3992f48017c06fe1035f99b2a07e0139fb75350535e80f75036190cd6aaf8
zd5fa0e9a1b6b02d296cc32bd712bf5bae20547200b108ed762d1b65649f2d14a7e10e8ac0edbf1
z602959075441c60de8cb53717f63b2e7c4870cf8517e06d9b4a8c3dbb9eeb55b9278799d32f535
z1b614609d37a5053981d6be3a5354cdf41d86f922ccbafdf81005ce13cc73431b0399702bd6ce6
z60786ea8ff0beea125e9650d8a19e4ce6924579ec55cc01048d5ebf8bfc969511ad6b44e00d1b6
z835f35fb8c2dd47b3da1b89b784e7b3838a0ef4a0fc156f0047b057674f61684d904533ef12eeb
zcd533f6a9c8998fe9abb90ca4ac6083a7de065b3e6d5a63657880c5fe2cd3174ee661628dc8cee
zab5b9783900b416ada75a0af45b9973080f21aabc40ed5962f2b6a574d9bb813352662873b5d7a
zee1688e8ec62d63184728f7a81ba7f00f16f4cc6a3cd0b76ea78349560c36762c75653f84524e9
z70a84bb2e5e2b523a39dc0a3e17fa5df06d2c8f5908d52489da8e73065b0c8adc409afec7f6d71
z311968ba407c35466e3bda08773a6c71e4d21b27dce5854649439553e32e5ddf5caa3b764d06e5
z9569d3f0e903c60fb04181bc47bb1b2d845e3ee9b2e1ba87710fb4ca85b4af17516d10895ee893
z92502d2bb13c121c1909c9d7e809613e3145434d7e0f26f15824fbb31c262be069caae690dc65c
z7261dda632a9f94fedacf03d203f8875cae1ccd389d5fa79ca8caae5df7a0aeac3f49a809d70e5
z5c00824f1796ea363cecdc610373a68ec0a4146821dfe4207b2748ce8476924ae666b5e86e9366
z530b536a33679ceda9065d55b1c45e903414d323441282d932f7f15f57c1eb85df7036d74c7bdb
z617479e7ac009605128d012e2a3582651c015c2fc90ec5cf1895737e938d48fbf32eae7f88233f
z93d38df41323b03dca426bd7cf0af90c211bd917fd6cf58c998976929770844ed34af6d132bad0
z6ad97f23cc7cf380bddc3a1676b5680b53a829a2e27fcbfb3bbbeb405637bed02a0f61e8009e39
z90e524bad3bfa7ec04068bbe22b25e45a80a31d2c70bfee482165eacdb8e2ea8db476f3ce1a36c
z0badfe70fa6d5424f8402b6acaf5f14b32c5114c2daa7b20c53dd16504e4e135b59cb1a8aabea3
z111f1af583927f315795c3fee6de62bf5b0043ad7ea61f0aad7e6752bc96899cda72a35712d6ad
z1494f509ea8782d5a510ad394abf52432a8683e165f60fbd17ed775d4bef8112cfbef5de7e3aa4
z5624fd6f0cd692bc7bd8ddf0d271199025c08ecbeae7f2ed41fe630f7c3137d9cc06da585178b6
zd291bebd2563e55e40a695b24d8b255ab8bf99262c0bdc0a3f40e8ad9aa744126b20f970f73188
zb48b1dda244dbab9f422198002f5cdd186ff3111cfda606c01d2b850b05d2b85fdb79adbb34484
z847a24e0d73c45d08f107afa67effd5aacfe1e477ec20d08195dd12142b7f83c13846728f12165
z809d211cbb987ef3bcded0ae62d4dc89d02307161367722263f310cece1deb2b6103fba3a6db2a
z19f548c68637d3ea3dc69932f9a442a677cbae23bcaaa89ce24dabd0fae13736087b69db3e21da
ze5dcfef5d2d7b59a46f3a82248f88a9e2fe2a27bcb0df20e4289d07c0d3bf4ea1c6cbce48a6b90
zeb7a2adf61093a069ef5ded246fbca755c46c9f5c824bba38fb7c0eaef8cf829c4cc79aa93e571
z7fac8f21e74f6ec64b71ce3aa8db9fc469d0bd6fdf7cfb1ecd197621b5556156733cef02736b9b
z13af6a95aa0921b2910b00bf4c2d6a3cf444357e5b81f2fd4580a22413c5f8f91530176188bde5
zdd4332b807ceb7f355fd006da704bccaa0d8a407932a705b8cf25e3d5052f6f0cae710f63e8bcb
z23a460ba6488a151da93b087ddfb86ce69db9966261bac82fc1b9f82078e9d8e13adc432152051
ze489c89154ceabe24210cddde6074f88531e7f931ed85bbba107bb938151a8e5c23036aefc0834
z571fbe0915f0723f93bfbeaf6cf68ab460c753d981c6c2e81381d7256d9aa92dd4d224eb82c118
ze5b4ad8920a757733e3f096d033c2def468ede6b7cfb6986e853301da2fb1039532098f0acf0aa
zaa1e6fa74f572c8969774f471512d732a9abadabdded3d417e9d97d7fd4a8b6ab61485a0669547
z5ab3ff16f5c9f9b8aca5da58f56c06d3afc3ed22f500d29ccd73e3a3aa7a84b39fc4f76e443c9e
z871aee681505e8482909737277559adc1ef0ed2cbe4dc49d16a4aaaf6dce0fb733b5979ed01692
z67fb1946bf0076f35d17f8dc93b2655e4ea12af1664d381f6a6c2277ddec4b15ccd86be4cb987f
ze99aa4d0aab5d74b6643090152c4988e33810892fcb442656b8d24ee152b082cac156be6f7f23b
z86fc1e0423eee8eb8ecffebbd38de81fe638363507a1ba289464ccecd715c270ce3575c543d333
z98a59e851b6c8676cce89f1f0cfcd27a4194584469f839941e438cb1951458ad91228360dcefb1
z10a96262d216abc3712ac567bdc17e15e725521e0b656a866a2040b018ab18d3c7eb1026dfaf2a
zf71491a7aa6450ec930f9dca83c752eced477b8898896e96ed975cdac4a185e45b1792fbacb779
zc64ea15e30ca0f21ce2ba5932b1fc894c7dd2c7b2aa09a5258f714fdef932ef7f7585125be47d0
z6c7f01c314f82036d363434cecbf16578ff0ef9afd9c0d2ff0dc0988fcafa0e2de6836e04b2efe
z99d7747a144f8041b0a0386788872b59e239c93bc71aa5bd59a39113bd7fd84616e2349831fc7e
z535d376b85da72d6e4ab6e4345917848040a4cd132cb345707555cfd306109d85485e07389d535
zc6c685729e11e65732d85bee197be283a53e86cadc8102b539b4e206241de60aa7893544b56743
ze80e9179689677373ab125835d6b99326543e3c6b6a4272557cd1aa8b4975a81ef9cf3cb42fe73
z01049d4fbf27661941c4be952fd89c67e638d212a6d94247e707336625cb7b57cd34b6b097cfd6
z374308bfa89c198c18b791fcb0bc33607c83061de936fcb7e4805937b52f84000dd4698042833b
z565282b4887a8b468651ea9a1ed60312223d3b80ae48418f236c5e1af89da83bd38c3b74bea81e
z577d20ef01057b5326f7c1011ea65da8374bc0194e9770c9d2da5aa7b4677d8095c8c3f16a6ab2
zda0d96026f423cf294ec9f77fd4a32f9bf6871b49a9e3a649c742525405dfe70b18a42f14ccc26
z8dd88465b4e63d5867f660dfb499cc883dc370fd0f4d2e5a3a9baf2b95c9a443cd3a9f5c0db390
z86b37ff022662e34fc4e182f64fa6752e93be575402afdbe34593953e2297f21e4b0ccb37d61fb
z8723f0021dc1275b43cf83b4178c40c673ff029b8448d65238809b9ccc5150b8c8510f9249a9ee
z118310fd8def73a9978445f38b0e15787835023f9d2cbc0f7bfb87a13a0ca7e79b9749af807431
z4936c09f9e0c5dabeb40f16d13a76811494701518e3a6e63bcc8f0c2f07de16b64debbb0553f24
z837dcb85e9981ff36ce94bdd15531a74a32fa229c3037b99ff3a2b1c9913d81d6dd3b48fcfd8d8
zb690273a88649d0d6cfdc72c44de7022a999279ec409c597c3662019fd34d78e4d3d01e8fd1deb
z476c81ce1758bfb25179ea5e0f684a59dcbda78ae74387604bc8e9bc4ba68eb9ef666a9d47359d
z26661b468c764748fdef1f6ff1d6fa949f08bb5d45f806b25d70da8ac9a99fd47600a866fca7ae
z2df3582d0f0d94497d157204d24942fa3624dec57cc7313c16d03b47ce0b594618abbc3090426f
z5a458c22350a46fc38ffadc1959da0b9d6cfb80e29ecd05b9df60b9fe6d36098e220397883ca98
z2d0451a9b9fdf519e9383de94404bfd9e0848625ba04aa1c8cac6584432f1dd10e96556976add4
ze187906d7dad11a26257cf825d47a5d6270c8509e9913c99c6cbdf4a3133939637781acc3a704a
zeb725b9c894e5e46b643019b6e41f3402efa04ecf25839f7f95aebaec6101aa945e3b9d226f246
zee736c232a56ebf8a52fdf14fd3c3c13b79bf1a97008995a614e1bf1e1bc2e3bcbc051b4afc107
z2f9af1761142350e0534b562bc906c025dd13b2366f8e4badb7509f900bd5b74157cddb22ffae8
z408c7a639716eeaae9bac18fa89505882ef085db7133f42f823b02f67a41277bdc8c01e7cc0846
z82d88a1bd399ba362891edda3766d9ff315dd794a2d2db59e2fa8b002dac1c600161e1332cb07a
z0c3e56c0228d6391f95d11c0ea757d68753ee4b7e4b54ede0d8397fe86fa1885720d2969dbddf3
zea93ac48e8cf36be086bca8b0ab2960e33298b839cfadb43e2bc9cf9e93f4a7eb8ed8d03699dbb
z05c2135befd62c1463adcbecf276c7a2e7ee69861c03240d76d8607ace0fd45e5b46094640dc94
z16cef253bc41db0f8113be30a85ee8eca6065f2ac94d7931e792850bf985c9a4ab76286246f4fc
z9f169c2d51c3a89e5ffad9557cf5fa12affefe9f88918b3e5e0777208a6877f09f775898d9a0c9
zdee5198ce1051c991e201a89965685e441f24cab88542c40aed2f4afdb38bded2d0cc69e5f37c7
z11cb68316a952041c6223e4b3fffb7515ad1f04037cfbb85caccefb33f27ef2604ff75d4ab6c1d
zf14de3d7089ee02fd0e9e7db31a142c001ceb7d7b33dc984fd1ba364050f59d60758435f936e90
ze356dca56a777ac039ec44bdafee6255f98cf8cac46088aaef51817a665ff0c90818cc84c3d3a1
z2064bbc53c717fbba8480088a60f8f9044aa1df9c0e5d28045c15fe2fd8ead97ba364bc5d51cee
z0719088c7700d8a2b21d54e6e5863674fe86759ddd7bb653fa8432e2fa577729cfa953d12c0623
z28e3430694201a60dfeed4c8e684c8cbf8754cbe9b310f1fc51f1b94b01d65ea8f37755f75ed86
z6cbc0c08e075c48a71d69f0823bc5444130db48ea56772f3277f6a5fb0730886d17fc1a70113dd
z97d2110c97764e259de35d53cca1d4eebdfaeddea526df332858bee2c1e1738d54afcfdc5c246f
zb81f5db70f32ea2bb843df812d8e69b9ce3c0ebee2f8dcc59404ec8b4f8603b5bd45a57d3a6dd5
z131132f28b972df713c59988330fe71f3cdc737ef93ab7fbba7fcef315eeea58741dea85c65f6e
z3acfb4cb09c29d355d4a26cbd55650ef5b89b64e451b0200a359fba1dcc19ad5960a1fe88fae61
zb86f108d7e06d367314445de2aacf94665b3f34262070b2919c79f655c774655d71c9decfcb86f
z6fd9f530d2bdfc20ebabb6c32304c6bbcd1f836fe1c83b28a5370e4529d2d1b2e52528c46497da
zc12b587660208e42c427f611c1038a308f269bd3048e91bc2e877f42d9b671685b86c5d14f7e81
ze8e24d7eaaa6cb036e9d3fd894d55d57f1e92da41830f2a884142ee977ffd47e234679a6a747aa
z3fb38d2551724b40ce7237db04af892be9c6c0910dcc471342083f794f06649b8a276257d5919f
zace345a562dd0e4c162bc6ca65e574539515ee601de4e76e0e8a125d55a0d06a76d81041ecc54d
z6e29f7f8eb509edf893f09594d9bc3bf2bf84485efb90bfbfbb23fa52f1976ef3e736fece01535
z3ac2d30a3914ee5c3344298ffad4bc7a52d98f5656ab0c0b0af1553421e40359a0a3262b0d34e3
zb04a5c1478d3e7ba9b4f06e1bdf20a0d022d5e30e2d3890fdf61bfe62d2b90e13b32dd8e059d3e
zbc1b7b4520eb675862025af1dd84b855fce3e98e80e0560306a79449fb3b3f037e4a4eae30d561
z0361990351b93854f0d9e9aa7e9cfb308832ae6dba18ba49097edfc91e30eec8eb290fa70c0958
z562afd5b602ddf48732859069f97ac925df490483749085b3ddc6167255d196cecb91ec73af0db
z3dd0c30deff46792bf44ecec3ffbda34a6b2b86e127f01cc5fe12632cd318d228b5cb99049be3a
z40bd82a596dc0053474cd67b6cb686bd1419b027fa07cf59da24070f20d4b5d59fedcb5a05a781
z40e19f07286c8bc850e1672f434aa81c13c112cf38eaa20aea58d48d65b9fcc2203ff8f2cadb06
z2f79fc0d954ce88ce41022f9707ed53b4d0a5ea7163269396e80e5ec4d028116e550a05a8a1e9a
z46388e9c911d02ddb2206d946ec9d5ccaa8630eb61a5d0f526d59a339df79405eab5aa3b7d7cc2
z010b634631c83894894d5ee301138961fc8850597a2952921378da5f4861aa783029929c4de90b
z695a2461b1cba760c0c1e47a4f2fc38adc5343f985333f98b580a1099152d99c4d7985dc66d379
zbc102090db9240c3fcf8ef1adbf885e68734a995af293e035989c01f6f38a8895114a5e86fe65d
z9f68e382c4ea40ce90cf882181ede201f736349f53a896117f68e073bfd2ef690759d24a900a6a
z75da280a162e1fd45066049d9b067d516d735c72466f5003cf0eedd70e46a37db04a58f27da003
zb9c364e4e2e5428c314578b322a248b9c942e4bdb50e91e11984fc50e4a7ac6830bc7a6be8a6a3
zb720407aeb89b5749c745f46807543fd5acb77f98c3c77ad37db7f642eb083fef7b7f82d001570
zcae3076f6db541aa6c25b5795a42a6860a32892892cb2a717afe91ddbe6d8ea7f4cf7ccd2b20d1
z411b7f0f31e9b56323fd6c9bc949e86e4f1a36738bdb5c1c63501a6f328a8243ef4b5a8af631b3
ze4b200637c7af38dbc305e327350d4f4fb0c5a3a3e01cd779fb061a8f4fb170808577b112f55d7
zfb54bf2e7f4c9e7a1da02d2e1607fc08fce2ce23ca832d490b27bef3f8b7845858fde368eb6b80
z09f76af853ebcdb6ab29cd2777216a4e1c7daea15e978fa01560bc3a8dea5198418d2d9b2ba6e0
zf55eac79bfbc0cd5a70794d13c3fb3e4f6d5794b1a4cdafaa36b9f82b815830d759b72175bd329
za5767f867c5bc3e4df533539c94b3804cc6237277c0d75a6a5d04a3734cdfca433030c0946f369
z8660c8d91e25542105ed2b0537a74f842375fced5f46dd90d3a166a8e8d5f48077820edf298447
z4ccd108300cdaa504b37c7e057bc22e24c12765a5cab05279a127bd1ff27139abb89365aa36f47
z1a9d7f673ce2862a49651e3bdbb7886beed8011cad06a2374abafe1811c098602ddeb423f0fcea
z6c0a1d1c2c8c07fcb97983238f93d78c0a9614c218c2a912a40523d5aae895f8fc4e75e3c9abc8
z4ab118a252a2b1f8d86a33e162276f99d70f4accb0d3c1eb5419ca96240979ce4e2299f31a4807
z0024f88cd37094a964ee20e84eab432471410874cd5d3be7586e7b930a2f46ceed1def09f8d960
z8d57e64ffe6d7bc5d7a7197014c9bd59c931cdac4ea3ac025d285296496827c1870e21542fdb58
z3ea78cb4ab54597e0279a8ae2fb72135fbaadd154b4ee48e1a8039bf742e995c6dbf047e0349f9
z96973b91bec0a7ffbfa49d2381d03a531a2a710130bfe9a3e0befe9cf7fdadfa31105e961e4bb5
zbf4e41bea47ba8e8a1bf15c84b559c1b033a0ee3317c72b442ccfb169c82bc27bd0496777e757c
za3b59658fc52c39cccb25c5965c121ea5c8dd484ec127296238aee633fd1bb8feb2d6a5c36238a
z07bdaf6a88729bea5ffe55c5ea85c7850fa40e205b4d81b03b4604cadee97c6a69f6f55c3f260f
zcffd9b0947e6b657126b64b5bde936276a36de69d86e1dd9a518656e0b8d094691f97bddf47f02
z8b7461855c424ccde4b03eb57babd8990d36fbba51f9090706a3fd26c3ac1ea11fc8862643f71d
z351d857aa9bc3210471afd0e49774e37cfe0de47a77e391ceab04bd1c6fed863c82f95f513534b
z5dbfaf95a36f88f3904705a10e251ca5e0c05deb93cf9e79e47251938e7a6d9c42706e7b584099
z47518beb249c5b5a0721be53fdcdbbaad4e05dadf0e801179476f0475f2c53156630e696c7fb5c
zcd7946b9dfeddcdb3c837b3cd06fe27a2c61669e93443fb5037a0e844d924202450a89465780b5
z8d87a76bd311e0c56af031d2e4da805d37dde8ff21aa00b528ef1db795d034f3b556e2c272c22f
z3730101f4a28e5f4b9c18ff776c7cc23b9af3f1cf7858551360478792d1fe1788b9e8521ce06e5
zc2eba2af3c5904c1c5befe1a68b2afd40d78a171065fb1ff34905546efd9e080351064420ec533
zc09b2cdcc5b2bb621943e680cec201dd3105e16d95928bae71b6a3a469600c5cb4ec96653a2d1c
zc612787bb66052852052c9675516fd3f45a2ab54ba5c51dfa8969715fef063813e9793fb58e336
z2359baf5d9520669d8770f9459ac819728f24a2099ebed74ef70c4b7eaf85c43f3b282b4e7bedf
z277040a637c4c05ca0efeca2281fdf0590a0c80b2fc4784e4e06dfe040995847c70cf4157d5613
z2a4163f74d9e5aa1fdcaac17e6c04907ac31a2f23dabd6852f54163df1fb085b521e402987c57b
z9d9b79ededf73f93d3cb01d7bfb80b3b4112a1a9e73014c3c6b656dfdb700298a9f088f8aacf0b
z57425df13ae92a3d77ca726994ac9174f09cac8405d69e3ca9c0c53b05730cea80cdf3bd5f7975
z6b7adc7d9e6afaff50e61a9620a5fcd458854b08890682f9ca5378484ab2b5f3cae1f5097c4414
zae4366cd8a2639f6dbf6b74d1815de0a7c52c8a766aed0dc55a22cea2d574e416a44e368bd8c7a
z4317490cf7f9bb827c462fa34db81c25348bc8e2b987df5bf1b22ad3b424d41b73212b69e697c7
ze02a8e1b67e6fe82810b7512085b07df81410f7f8c6cc34e79835ec9f00f71a83144dd9afe592a
zc0ae0bccda9763e9ab98e55e68a943e3424e26fee04a361440ca606f8acd486d381d69dd53de99
zb0cd7f62f5ce5bbc7254471815db696b5c7e57c4deb0f6ab104eb96ed3283493f37879bcb15b12
ze6d6c49f893a041993b4f8d2a8224851c2536c0ee7c45f0adbcdf7edd7bf0e2fe2a1d31840dd4e
z31586ce3882d8e44dd492000ba5da4fbd68bf2c319771d4039f8fd791f61435817300f765aba85
z57ea9a866a136613dbddb9c55c1bf4d9d98e51539ca1e7a5864093ca6eeb3d8a9913580207379c
z80a409da05c0bd17d8210959208de53e80e5ceee2d612dbfac034ddade7440450d16169feb6053
z669f4055ece5e37cd241ee588014ea90562b11e94fddbddd411d185029f3f4bfa1aa0127cdc108
zc49d72c5084972650aea53b1c93a20a19f6c173723933e150577859aff5b9ac587538bfbb17e24
z0d4e07280a99669c40b7284792d55a8af812fd71d998f1650866d691b118621d413efdba18f9b4
ze0397ceea500071fac081f9ea6ebc736d4d7c2e240f81afd72e41dfae8c76389407fc30339549a
z582f22a52f260b8ca2afab07a67bfac388d85110bfdc09e0a53048af6f461962eb0793782140b4
zdac263ee03a7519e9c1ac3ce1cb0a40cbc519e729950753a6c081a7ddbc5e31f3547567f87d858
za8ef9c7369f18b5857afc2cb802dfa4bdf7474599a84e9ee8d17256906a34ac979fab7156cc1b5
z07a0c36f13554f99314c0aea69b86896aa8d2b62853257751529570f026289dc475235b103b9ba
z09a3efbafbcbcb23170fb6d4b76bf4a8c0f3aef9cfc5384b670fca0eda102599dd2c096812a446
z911881420fcebfd448ffd70a7b44045f2e134909a81481b4012e0471067efe9330429a2fec9060
zbc1e2fc77adf14397e714b25379edb1460f723e29ce1063e11e05e0c5298535b64b9cc38f7fa19
zd93ff4e3828e7f13be51ac8b9c28524fe08b822091c9c93ba297cde85f0bb61d193098afd17b8e
zd091688fa29af04ba007a711effb81cd639e40d9de53bc2bd2944c1d576204d7a9b759fe3d315c
z3c4197d625f8be946ea26b5eae05603669025eddfaaf1a83e661df96f6ae2dd74d16a44937ecdd
zf50a933236256adaf6fd3c0875b13979056fec2b5bd8c55d4db1d5f19d7c71aad48a62a748b897
zfa418a89fbe959979872025e559b6c95fd6b4c752401b11028511cd016044ca48359fef12106c5
zcddf4c9026e16ac4bdef5d17825caf84efe71e6b3e62a16f4a32827a750e8a2d56f101c65d2e64
zbe350211a7d0fb3d609e2e2e9684950150c7090fd048f1f7abed15d8308257a4f565a854dd389d
zd99bb120403cd28f8ac3288076f332b41b37c8074488c7aeca4edd1f8e8279d153cdcf624f9fcc
ze43ed4c06376bca157256b69741d5cf365a3fa57fa52281a91217f6053207306add0f654fbad7d
z38be9a6bd40318ffee55dc31ae476b6d26044235b3494dbaee158848b9efe2b9321b9dbc5a8f5e
z2945ed5b77242130ae425bd21c3adf284048a8792a20af10e82e0860e70a7b675c79911e9ee715
z7008f862f9625e9a7669bd8eb64101c40a073030758b9e49e079964b305f57f5278958e05326a8
zd766bd9c80b7415666b2b6278bf2ed12d4d6b0e349642faa36b6ce1d05a6f2ca4c0e53e7ff1aa7
z19b7f99fb6803c2b7996251cd8280fc4606c6ed3ba04aa7431eb7534cd56603f797c36aa438f11
z24378e145830c9f32defe38f35ed60683c6313516b35ef72d4fe78bc0279bc204a4d75a8c915e3
zf1eb23913a324e2e0c1b0e713da339e3f638622195ddae252f1f8226bad7afb4433818ff46c60b
ze988aa2cfe1f4129db89948f69f76eef6c9e4d2a788965c8463a060dc63f02bc19dbe3e34d8c83
z9a017dcae9ee17f0c381a916a26b6f81a22bcf79cf119863f32af7ade54d13f7a9089769c2dcce
z37e845c09feea94cd21eaacd98675370580d349dcd9ddac899473c73acb2633872a1b71b0bfd32
zebd7d07bf6050b26725abc5d7824a98221d7890640610808f75a4171cec68e39b322f779f86e83
zdc4a0d9ed0709a66f12254033e352b330346c484a4755ec05cab765377b5c2b784d131f46c0ece
zfe20687b16af31e4168dba11f58f7e6fbbf3dcf5275b3aaaf90c7fbc7786147709f2f559207036
zadd771a7f4586cd0dc05c3da3571dd1a5ebc0d620fb8e4756fd2a67e976644257cd66b772ed8d1
z0eea22e1e7611faf3b4832fd2f8cb733007d3fbf2e9c30fb64ed007a4ef1c8dd0918bcd68d55b7
zcf49e320a8b6b4cc624be15ff164ebcb8f71ffa926f38070e0610575c2c7feb597db5f1bd03116
z64cf3484f718d5c1080984e5ac922e2d51046f247dbcd940c0dac0dddc991743e27f4c7d6f548a
zc9a5450a51a51b2703b5b1816994856c16333644ba9c98ca9db83c30991abb63506da822629b2f
zc9b0bd0ea2948e8fbc0e36daa6395177304af32db509a6f59ac0a8c8f3959e6945dc65219e3321
z601712148af59ae6bfcd1119a38ae3d3e989a386b2d53f16d636fe7fee3dd50aff326a9d895207
zab94152b51a38ab2ff68f937422921b667b4d5104ba9f7a6670d893fad40cb416adc734f2380e0
z3523a2dfb4a4d625e718582d83ed7a9a3a91cfec4d5a6586b59d99c839026b976f1b480d29e187
z37de4dd69ca8351f8e3b35ec1f496c8fee99d3740a35f729fb3528e17c48f276c4d60aaaf331e8
zfcc87e115386ef0c22b91f313af4eb01d66245828c77046f409630567c55ed5d48e22616987599
zbc35b9ffc3db4796aa2d9646a49ace72395dbfb4cb09afc2b0e20b88c4fbd40711e2e692a1d16b
z838d953e866880b6df564f7ea7dd09bb4dcdcaf0480d27d5bc0528c7ad16506a0170a6294f3802
zdb560349aecb60c77f5bc411b914577370ec65b0c2fb0889f8395ecc925eb2e8adb6d1891a7a3a
z9b4cd6e0caf0ef0a779ca5cf586f47902ab591396941d3903b6babd266f498efa5605e5b3d2afc
zfbc3eeff8edcc3cfcd1d114a7ceeab2ece7fb6ab94e278a3e674d76f3b8320ccff790113241e92
zd76262c6ced5c628fd5d409b2417ee177d9b67055eb1377ea1fc2dbcf027eb41512fd8f4b09aeb
zef69beef6d011368ee80e0d7057f81593856ebb5fe2c706498e47c1e4669eaf3423ad51cb7fb4f
z91891b8880851c6479a95e4647ee85d4a7ebddcf29067ca795408593278ce2bcf1748460a81253
z7493dda18f53bfd28c8e89b16825ade441039b73382af93fc628f68d371f53015ec57b455d9a20
z9442595ca8d3b5b4c7e27475577d70071f154678e0061eecfd27b8eeb1e8150b7329c8d1955e4e
zd53ff583ede39556f3a8a66dd7bd0a4b3bf9f0c5758272570c8bc04e99a76b6fec5d2b59032387
z1d305685532872aeb78a544898705ba5888506c10ee8ea304cfe485ba5dec9b06ea1b41077efc8
zdc239415a5da64be48587f427a38cc551a1fbdd24961143539780b41b8288554d9eeed43c1d349
za8feee1992f86347ea0d86e81124cc3b95a49a159874d8a4d64e8cf065568c03a9387254bbeac0
z9ac9907a3c8f1f479767cb43c78b70e93120cdc07c3a056201ec1a664a7f078c2324cdff0a3655
z63726024f274316994b5746292e975cbefb13a4a89df6f166a95787e9766c22c55d7fe1a9ce7a3
z76acd00a2da97738cdf46eafb31a6d432db31ebd1258f8c142d47039f2ae5d68920d445604e671
z270fc4116429f2725d25abb9ba9323251467a69e4f2edde74b8d547fc7cdc824e5dfa79b3c4574
zeb6e70a729d93fad6f522c535321ccde5ffe82f81b61d8d287b4d823d8e5499e4be20c79237ce0
zce2c461c9f0878f210ba8b1405efae0bcfedef6a820a86145aca2d3879ff65fe51733cf57c1de4
zfa8c38aa5f97599ae58f11258a8fa467c56a4c53cac52ba39a9dd513f455deb3105475240495ee
z30e8537132898053e4e596bdc6a3ef5ddb09b26f1e9f23ccbc049c040919878ac81dce94b1df10
z7e57251baeb0d5bdb32c64a6e3d512958c7b3e66f4765733a82bb6b2b6f276a950c549e3e98a7b
zcadcc4ed37e7d2d1e639b66b855fa0b53d0f4508337acf23c5eb76ad428f878d08402c3954b109
z06c4dc661054f38734996e1ac42e4b21a5e138b2f2e359ecb27e9866f822fd2694895327934a81
z94a140adb33ee643115f3b7d7b9c6e3c948c9599a6fc77cbe3ec9408f6d18485b3aa44d106cac3
z85d27abdb0d03d423875943214a6d09ff89a2a9021a6e737b94d88006c9b37e64fccdf78fcde6c
z06616fee2053071be3543470e272f0e5bcba6317b4dc1898b52e7f7755a0cd60e89c797a331450
z5516f4298a488c11a313a46614f17a94d416592a318cba256a8dedb07bdae726ac83d2217c2a69
z3d562b141e1243fe0f425eeacbb1ac29735344e9f3b2f8049b5a5e1c950c67ca7b135722686a08
z947609bc217f608154fc00e3a635ad33e2063b02ce0aa310fb95b3dd125c390fe947e1a2c45f2f
z36d10d08f2abbb5e06468bcf88aaf0611af2b34d10806df5b542cf85b7480b0ea92a6291a1600c
zb63bb2fd2e8ade1282a0f31f3c62c83510b79ba1cac1ea45f21d5d314294fd1658997a3434d215
z340c158dfa449db79a10adf18a787b5d6016613ab1bcc68988ed55a098441050a3db4bc27e6ce1
z963b1f5a6517f420cc49f5636a3684d45d5e45f08d04177f8c1cb8ab25e399fec9f68ef58332d2
z6b5ed753f887f16c6746c5f39f508f191841c6ef61964eaf3c119e6b294182b9a0319c9be79c71
z56276bc4f832bfca0dfeff189a150635ba484bd2ca7f17c17962c4bad562cc3ce91a6445418a5e
z217033625aa617fd1e18788b99b6c07f1312fd8d3764e8efcb8a91bca505ffa4581a7a92e842d6
z84e68e34ee6260ee7bd0a628a80f0cfa7174e8fa290f4b2409ce0c68fba478e305da724e3e5b15
ze41c4adbdac9392ef3444f70233bff016b5f820a830bc904efab997741243c39a776d2d5e09812
ze433b14115ce520f7c9c01460c9f998a44436f3308ef8cea66d1ebf9d7fe65a3eeeef61fd064fc
z194267a661e2a33e9cdaa22393df8617439c10afcc20faf066293d3508770d9a77cc01545fb6c4
z987abc29ecee1023cf079921f405fba4a7fbf2c8e45d8fbf2e8f6ab1342767b5ab5010e4ffb933
z1e178b4ea355067f36e3cd70b28cee6277a350848eed98d1141aa260d225518501516819af3097
za6f1fb3a7fc0bfca99e19aed92987f6b2ee6fec5e68afcd7d0dad0e9e38694b47df19741553cc5
z3620fa9679bfa61e5c750ef90f92d17ea6e525672af17fe0a711b8f8aab49e5c6a6cebc74cac29
ze91f7abcb27935251f803c5338f49b6164311d11c9ba3b226943d40015e5825e51dc5ba26f292f
zf8c1681ff9fc8a4f59369a2a480958b0ef31ae39a91caf53064a88379e6170a5b9c284c84a58a2
z610176cce03236e73558826a8aac59ab5b3b79b38d1c3109bb7385fa10d88425886199accfa79f
z591bdefa07acbbb7fb5674ee8ecf4f32d1187471ee386b2c8ce8c99d4a34cb913aadbca310da4e
z4907169c08e30ff1f76bbe6183068a540475a62de3708b83da7d857e350fb9c80a3911c64883c7
z1dd0650f6abeea3d6458313097c447839c58d3c358eea759cd0e5e4b11835e0b2bacf2c0a0491e
zb373873e48faf17758f93f8bd8c83adc20195b1f7b143249cfa0b64a65b5da61995e9597572804
z78b8a316fa3c4502a45273bae893f63f3a92ac109612410294013d2c629e44704ab26a22dfdf6f
zffdf7879eb1c52ce4e83f7439b28648b31c1f0be94eca15dbf8f6bd8adb6927190b61e39cd867c
z8abf29de29ccb9992bb7bcde270ff7b2ec4fa68079d89536dbdb3761441d9c6ae11432441e53d1
z6939885511d0ef1d3313e1572705b018cfd612e5de704fe28de5e20a8748a2e5c329b60e957357
z3e400dbb5e925598ac697c519754d8f2000308b4575cfe20e2a5b4aa08d50ccd15573fb818b917
zc03378dbada5b20377421961dcdccd061c0ade98725f8d9c9a473fa697e2164824133dad145c8e
z15a11e4e6c608767e7b812e036630789782ab36d8652ed1dc2e688432c467078c32825b80fb198
z617a1f673b69e15c751b00d814362f3489ef9fe523317b04fdd9600e38eb0387bb75020cdd4a65
zc067d2f55cdc1f694a1b1a429f2f2b76290b572c3965cada05705bd573008b789c9f821640ba1f
z6c3248a302a7bb2645c061cd0cdb090dfe08033e52b1a1fd3d437670f716c129b48ae7129d5b47
z70d23e4eaa888e9310814783a025b084702fcab6ec9e7f55a5ba216c0abdbdc4b686d14bf14b01
z28cd3f9fb6a7c056b0d1f983162b14bb1fc715f6887e0d288570181c77a11819faa2d423af27b5
z492b33db3f9e35d8d696be2efacae223900e648cdb6ad120f88204bf4eb7aa722ed33c223545ab
za95327efdc549a3452b7ae146e86fc563816791aaed9df17b2743f75fb93537f36399ace70afd7
z48f96010faf0d0918f8d34aff69759d05a18dc8eacafd35da8ab1fa089c021ec601bfcd730fe16
z89ef705ae9d9a39ffb19c89f3f4c1e5471446b77e62c64e6988e8c106b0a93277835514b325018
z94b957baaccad1d5fa1bd5bc499e8cd2afa6aeaa5a9157708d0b700e998cc7dad9dd881d0e831d
z909f4047489bc7c0c2d0177e7135eb5a2743a291873f6df3000feed2c6bdfe5e29079e2df6c94c
z1f21d2400b7c0f2b0bf7fe4e67942e753d273137ebe0423d850a31497e4c883949b365a46f6ace
zb9278fafebd79863a43ad3290dbdba4a5c06077a5dc68b75c2ba5d1f7b538a25db542d54ffb794
z6b152353f57e180bd5df7a8cc4c0a2be464bb287d7aa6b715a0f0590be34ed0cb3531495a66516
zfff1fb3e8b518e2893ebccb6ffcf98a1d0ce9338f0623bada29d87d991549f3d9ef8b1006a9f3f
z752acd882010aeea9f9f90702ab2e82fb406743696aaca8d5ef0912f8ee921598115d1ae78bab0
z5c4800a6560d55449fb25733fa94994e4ddb06409133f19becde453868a1a59b9a6394915a2a0e
z07ceaee787abff3e76654e29666724563b882008893d93ae0a28662bcc2cbb4af4e182e9a2ead8
z5f0b8925034a9e1e66d1e11feff131a2aadbc6db02cff871408a8c8e5d682ce4ef6810f1ff80e9
ze04b3267abcd8f4bc50898a9cf514c6488a251cb04ef07ca4dae603aab6952832264d810145fb4
z95490d78c479bca835954b77da19f092de413a94c9f0cf34d6eff757efa80c0771ad5fa54e5bfb
zc17e4ecb026d178689d6695a47fd21d35b33a1b270045c1183c261832d6d5b3878f9dcb84bee07
zab6426fc7cb6966dfd06fbad09018ae695c35755de766ae328052db2e30206dc21c9b56c7b9086
z7d3ee76a440b52c4c02d21115c8ceadbfeb042f7b4dcf2d092b08dca32b3ab248efd1d12303555
zc8364a4d3340f2248dd02587eb58457b17c64c56cfb8bd081130309a04cbe7126f35d4cd94c12e
z8f4d8e76d8b8c8ffba412c855ae7618a8c6a5e46d448ed84137843d64de4dca14a7ed7e1cdd54c
z3649d7eadc02fec4ca1423ceb36d0d8d24596a5ef7bfa7331b6d89afa213382e741c1c05396513
z1312de42e95f15d2ea41ba30c627e74ab17b50ca6279853546e6ead36460756ab9548d231db177
zeeb7fe4c1d7602de36d9c7c51aef478aae8e5d8c21e7f128d38754d1311a2d37658ef8361ac4c7
zdf04008665966eff52ee6ce375e393f078816d89c9e9e12f5c09c676e8ec385f534068d4e51ff6
z7f2319e7a2129f949772c855596d426f793472eeb1cb1f1979030f0add9c0fda5957e6adfa5430
zd52451292ed0b333015290b0a1475a66230209265fbd9b8215777a955190213824a8aa7fc07f6f
zcb0c54551458cb30d0eae87870c14ebc1bcc946ff991d221a8a9354c7dabae379019e5af6922b1
z41440c01aa6ca8f7c9c6760d62cb27e8b28f3e0343fd56feb71c723859f92cd6959cd96aa4c24b
z9f991440f932d819d137f6b3a267de82afd249ff2a1667ca868e684ea66109ba3095bee9ea207d
z3867f350b2b7971640df333f2214bea2e987f2cfa93ed5cf2ba0c4003f75a89747f377eedd2cec
z6aeff547a01751b9385d9be6abb8d34d2a98aedec71cef363348fddf5a54faec30d2e8ca7ebc90
zd3c19d75d7f7e8b9dcd2f18596177132d3302d86688b8b7a5c93e9eaab4faeb05a9b523e85818c
z7325ea094b5f16fd95cbb68bd72e325b9a2c29c91dcaa35ba2cfc283e6c1fb1f7b0690c64376ab
zba09271c0b1e783ac6670da81bde105d02814dd9c67b2e141d29237d56864e48dc32a39c78f31d
zc0184bd947dae38193a68764640865ee582040cb4e9308c4397bd38ef7800057d2115bb9c1d3e0
zaecc6c17093404edf7fa5aa5c9b69871b203613ca77455a7cd1f3f487f73b1dba315106eed6e44
z5e2a75967dd3edfb2b3df6d8d9bebc056ae8e1fb8648951a23315f2c094f33f952ed6c77a87309
zbbe05ad2bd0460085d627d701863201c70bf7e2f7f350830d7f343fffc387f7250c40df6fc8abb
z518ad7214aa5bc75129b22092f22baf8a3f1295eb33376b46f0588d825984c345d2afbe3c018cc
z9dad8aabe2116aaeb825ffa2f72562f252876a7c0a491d54d2287578212d2223a6780c9dcf88a9
z12ba516e6b449ba826ee61066ae4e11273b0db517e37223ca73284be08ec9d3c12776aae6b9802
z15094ee2adc20014d038a9ea859abac9cc4340e8cb24320585e4335edb4ea2decb111e494c9ba5
zd64df2fa05f3d60521e78a1811e3e52e12949aea734cd6d9a5bb4ce4676828d2a94f7456d140be
z6b289ed77c63d52f1206978d69a7d41e1fcc01902fe1b40d4077c09cf5ed3d86e41817d4272a12
zb4d15d631b45e4083d899dd20bb55344815850cc69b79ce37f0244de2fb662e369d5edac48f60f
zfc2559902dcdd363e393c2dac7292b4d6bb6f22238d94eee1b02b66169f7dab47e092af1e3ee5d
zce8f3486b3faca00f15878c5d594ba65b0003b504cdba29796227e681e51360268a730945f6114
za4c811f171ec67087ce82c8050ccae6615f1d5c0c0580924a37c2bcfa38647d0a8d4ca7c7a8e02
za354c0603c96439a898e3440e1a061e4d1e2c9537666579d1257f51b613c8eb6bca4e83f988e29
z41139bbe4f4126a33c5b8f37e8a26c815c7aa8f051e48a1de169b1359938024a5c92617d7e6dec
z29f459ce33d1f2de89ff4eb6116b2ff71a302beed00ee704bedff09610a58082841f1ca13572a3
z791dc04ef66a1264907105ed2bf53a49216b58480d523d45515e41cd4eefb1adf892e6f6c6515f
z92b7fdb61a2177d823054987391c735da352542be039532254eb67d255ab3f00e7b8077773b3bf
zf86e819360f4ceaae3352e15d8086be766d5a09136cdc004bcb8f7357d9ca5b2215234229ed1ff
zb6c5d0ee4232ece56dd73594b6d902eaac71b6abb41acaf5116660b8e6b3f02e2085caf80917de
zff13c64a7a7f75877de15470d3851a098f2e5eae2310b5b9e62ccf478d39a507fbd54b066cb9c5
z0241817051f5c01b980f68c57d35cfaec9dd21e2401b9e904e1da89a841c2c0032b788fc6b0c2d
zb77994f18d3a2f007c0ca1c8ac4140b21794b06abff4ccdc96b9f1e915d9f6e6a000c7512bee9c
z10cd4239859730df3ed3142fafe8b9b0eed10b6e3337aba0f3b21c346e275d9fc55c509b338774
zed7865257722e033e49d51678a6994cd7b5bea39d727d5c43ea48b6fa583beb0ad08848f72ace4
z8da2e1e8990d1ae245098c356863161924fe9624f9612747e82973f522f6c6f78b6f86370c02e1
zad28b15a4fe37fb2b0b116a509aa672bda72d7b4ef952d56e09452c71d9bc59f460f7bbb5748ec
z2c5eb8b548ff3552c26df604ef5b738f81c8fb7481fba7ebeceb71af0381465cd7ab0f55ca49ed
z3ae12211317a82d081d08b951762670a6119269618621452640ec2f69358871c4ec08aa7027e87
zcf675f89265ebfd269fbe70cfa80b79c558a76b9bf2fdd45a3eb7604a13d72c1a2e611f5ef6c27
zd72f02dd7b085284004755dae9019a3debda658e4709fadbf760d4009ff7afff9108a64e49b338
zd0f51ce677b71042dd78d90a0b92b4e138fc492c1c92d3915ce1dadd2409269919ac4b7e64ce5c
z5f50efab03c1202e2835c6a53861a8488634faf21d6349bb0014214881783c50f5deca5a11ba67
zee8d0e9ef9a1b2387a911a28b37b900ffce7f4e07cfac740021e78b7d369cc220fd6e0d4f15015
z7a08ea072d692807c596db50dc00c6e24fb021711990e8faca9c343f25aab574996389907bc5dc
z59960fbe9181a744db94f100571bbec79a3380ad8871b582e58b3e734a8653ade870bebb7b933c
za82997ff075b8fc5199191e6165ff7c584fc1da6143aff4e368640f3c5c5618fb89ce77581e56c
z37c84073c52a5c490f08957a4fce7d7250558318ed61fe5c445efdef11fb9bb3707ae94ed03464
z665ab8e83a77515037e009f4e90e24a67fe1aae299147f561e7fadedde211342c954ae0c79d387
zdbe87aa9f6c877990463d3ddff4f01ff5748bd5bcbc40f62c52453b894cbb7c94274d14d80b2b9
zf12f77289fbc0ed768fabbdf5e080846b70d3fd2325fa78f41d39b0b1b8bf9e67493fc4375af54
z9743c63f5b9dd0b57976e4d6ecf3e9b2cb19a26f26ff7b02be073fb832f19b4507a0caa162beea
z63c3c104fbcb2fe8666b1a9d0371d56a4140dc62af6eb7e8b5b32df90dfe637e4c5e5c7a398a27
z1e76f0f4aa1c80450afafb373589a1130ef9df85f32aa0d29920055981cfb9ee87c75d0ef217db
zd719d412e2cae5b7083368f82487ef3c7ebcede5094b3bd7ee454262585137278ed5400d5e911f
zb64fc797287189458cd7eda33711063731ce80c6976d3c2084ab2d8ae0dfe867a211b6cb5f5f18
zc6baf92757fc06cd2eb2eb456e74a86d9b1b3e9af4a9d7d4def14043695912549cec6728979ff7
zeeec0a1d9810c0fbb555d8673e4eb234807a26c61477d65ef111a43e5926298ba117e005eed3f2
z58a3e717a28cf2ce555c5d819529aaaea8725c7a70e1a408727a07be3b5ea2dfd56722af8cbffa
zd1b4ac937ab1eea9448c8f03ce8dd1b36bc89b838a32aa973909bc531d6a6e62d57283d56ba95d
zb6f3ba8cd7f9545513bf4d69320396dbd78f0b6cd5b32421e54582795f63e5dbea73d3728f2eda
z5c2e8c9cb630d2533ad50450ee9cc106c5960d7b1a13a8fbc488e4d233faa2d42aef3471bf1a09
z9f9ea840472005e0cc739bac82b6182ac039ab66223dba907ceae14e35b28ce90c17a48115a232
z0abdf96c4f150602c40aad9d1c26c306b27703e07edcd5958fde45d1b7c4fe64e7b518a999d75e
z81056e23a02950555b955e28f55f9288557d9b9acc8ba7646d4ee4fa276c24d71dcb0e728cff57
za1d7164dd64fa88b0d7e66810b33647ff0b416518fd0859697611f7e2cb81e5b663302fec02422
zfbab8496ed5ca30658c8afe5d5ce4756b96cbb4e4438adff1f910f57dee82a9edce8c8ff18c271
z408a6264df61d10483c746d697f7f5708db330c6d6e44c95a01c94f4a7e4daa360ecca79df6fdd
zc7957e24202e60855f785cc81d12510fd0071c68348aeb4814367990402389a99b6101d42ae5b8
z2b50ed31507e7f7ca769f51c1379dd7f217c1fd324c21a5e8ca33dd763bd2dd6f36a59693e4a4a
z35ecb427b6f3863ba2994f9416c27a6148214655ca5a4d7489486e4ac67b0266084bbc4ef2423c
z0c1acbf4a3d09820ba139e1d3e79b1249a39b141068d7207e897261f10b01b4925ba01a9419efa
zae4cf9205f964f124a705cfaaf5197ffdbc4b6fe1797e2cbbe9fdfd466e4a24e849730e5f54122
z567bcf497517a72a55c1439089ccbe69b4539a41d9d6fc37df02e674191bcdb30d48dbb89f96c5
z603dc60976b4601220c34ffe72a2e1853da325c03712136af089e52de559371ade99cc5deb90b5
zf0f4121ae81197ef4b0cc3b4f0d933a59090c16216ccdb2bc94a7ff107ba8ab6c48920944fea87
zfa0ec89e9e11f8eb5b15a72b7c5f4f067cb9a1931ba023fc424ad101b686628d27af19587a94d7
z9a35413dc9b56a2383557325218cbabf25cb8e4b36247b6dc88d018b88aeef44bc4d201f7f46fa
zb61def5276356a33240e074998f0e0f10d31982e3fc266874eb488e82b55653b3b8d377b056599
zfd402bd17198a0be138324145fc3292d672d329eda719f93d44a461a4c05bbd2869a433fcfe37a
z71e9805d0254b60d45580967f444406b853699ead6dff4b973c8e6378de697785e5b28bf9d3886
z96d3988f57a75919340f2118fd520704082afa2b4fe6d25e0a8eb05838af5c08970361afbe0f7f
z69e428cfa24e7ddc1a77bc055c295b89b2ae6a9071a738f3430d8c36e9a2f54ef185b57bdb3c9b
zc8755516b8504f73c9d4c5d756ee1bb30e9c710c788749c6e72b951e7f65e26422a52ab924e852
z1752e0720579582f33a003577fd516c89db4275677b1aa961af65581c8275eb9de8f5fa8ef6bb3
zb2b697aae5cfcdfab9ea8c51b4c8245986deb4150ed7cafc12c00f2ef1c3fb76bbb031d6739520
z12041f8965737bb6b616014d67362ef565f4454c102cbcc2a065d5e8eb6f46bbcd6336c40787b7
z9a2d01634ded410691ed0fb043d966503232c7c8df0c6950e4a60bdd6c4e67abb7b07393eb9c1e
zaf388306708e67f64bd438ebe69b259ba2fbddd32288e2de442526c6b12e405d265e6c6e44a74c
z95159d03ae480d9c14194164cb2003e0805dfdf6ec6e26e13f5e8a764d83ecc2bc37420dc59721
z9fa62accd7bc43f31e8c038f65bbf230fb7d26a2675b5fa4b9e3e18da4d2225963711f38991c59
zd612363bc7b303d9c8f2e8ba6b4297e8dfff203ee34644f6b480461cf14b91ed47ad009acce5be
z43317a79ca39c098b47a71523bbf2c8821a7da22a1498de8f83bfa627894edddb68523f4efbc73
z8bb2a8b3f18cc04c265a02ea2b2664a5ac1c3728c7fb8c5bdd8e7616bded1cbc8eac801a96a657
z4dbae3467fc65782972e198af26cdfb7254e3a2f1b6815d602308e84dfd202c64747e48c51cd5f
z35210fdb296644ac100b2ceae0981c202bfd4396a407ec3492da1cc573297d2999ae6fcddf7ca6
za649441c46352e3a00f57f885c54c71f6085e5baba4a32a8be8e25c1b526f2ddc7cc0d70cef093
zc28c619ef7ef2c3b8656f3011a5f1320aaf9a9afe27a5eef86a6f01ea6feafc4cc9cabc3931793
z3041c54446c65219be8f0304bcb640f9a1edfca3318a5e8e8150cf6fcd6e820f9f176a934df5a3
zfb96988ee7403092b77694a675168b1f50084d317d2bec0faf7aa4776f9fd5e6e34b43968247ca
z3229b71685a716602c17c8dd897fe31d89b017c259285623dc37d737c558ecbbe75872c4b7f06b
z14fad3ab2fe8123f0e9c0c826fb489978108eba230a65cfc9c9180a212e50bc5a895a05c16b8ba
z438cf5f658ac5de346947e50cfb1f2adae8e155ed50e2953f7e897f53c7ca46ea9e968fd77b928
zf64b6f10d7563e951622a4554ef6709d472d45cb2ec3fe54a4bbceb9c30f1eba1573c8ad4c5f69
z09542cfe76c5d20d815c0ba3f51eef4c2bba38e0ccac097f438e10e7148030830774aa502d7456
z6e4fe5037e76cf7eb00903091e7c4d2f65dff48d95d218a218d661db8b45fa6d0adef55067d33d
za0300a6869f8bed3c28db8935b2c996828a8af96337ddcab9099d95dfd86b51849315ca86c674f
zd95e75160629ceaba262655e0b6fa951d8f7f1b875ea417866e94a8f03a4e67060b479e8eac14d
z0a6351156bde6047f0a8c5055f7e063095595a6a6709f8fe4c9064da27151d8794b5887fa25383
z995f744f806ef6551abe07fade576fc6cfde64be77355dc8796b00e595d21da535fb5757cd0173
zd1a5620873e26ecb4d8137b1435b09ee1af87b4952672a3762979cc684b20685cc1ddb3d3b4d89
zabb7dfbbd6ceed3dcd9c656f23daa55dcae2a5a432c3849eb5090884920f9af12e69bdf2331aba
z3ea738862883dd63425420fb21d0c6a76e62c07b048197335dafe8d0737c76e3aa6dcf768d61e0
z14938fc24846e1caad61c60ea864e11fbdec3f8714578ab48e9f50bac63de248f6d3e747d610f7
zc724d15cf339f1bce04b438308efb87b7f2247876c4f886e7d87fabdf5d7d245acc9bdfe736779
zf49ba6139eab3db18f5a0a78270d130a0bd28fc65971b56ecdaf936c9a438840416914212beb12
z86abb41843bb0d9e6403d952826adcf2d14901d905b814636721617c6d0eba02308c0f39642477
zfb4a6202800384f6be56076e8f256ff959a1437f8549e865dfce258881bbcf8d475ed455b79b92
z47dad5ac0c0a4d6ddff86789af638a8c9f74999efdd7089a3f6361dfe54dffe2a63aae9e39d59e
zc2e4153b5c281a040d7a7cff9e2b697eab00e0bf7937bc8ec2d167073365bc41be64498aafd6c7
zc170cd0391ebc3ee7b6a3e9427c9aba8085ad099a892ad39fbc50f25673dbefe03b61657a079b4
z29576935486421f265170ea724575ff5651cc7af80524f551000c2ef36090736e8f286bd4a628c
zfb1c7041b4f41cd9e20b1ab59d4f4b22437d154e18d726cb6579cab64239e92f8affe9960884cb
z6dcdd91d52d1d393535e85ea2f9cd13cd4e936fe00178bfb16eeeed07b43bb54524532e2ccff76
zb86cf71f7c0d296fa8307439acafbff08388bfbfe32efa133f24f5c30c1359ba0feb442907cb9b
z677df08de5e115a0ad5beed955fd5845d6e0fcea89c1f4e7211fca27b15a60a8e01e115aa1b5f6
z56bd9cdd83229a564a8215603c28ce995e6170e41d7e4f2e1c5b0ff7945fff8aa96454ff87678e
zcfab2ccee71953ae4467f2f52c3663747c84efac83490eadc5d7c9b4ab925b7c2457b08e416a61
z2c882d27a28a0d768170516f93987339dde10eea18e04d5462bdf952bcda723e9e5494e36b13ba
z474325e41d3ad6dff4a82c2b83bb8bf6a118dc8e171102770dd86c51df8de635b689891149c588
z762ff21683a1658d850700f3bfe519d0ac793f7160432f92954436293fc979020efdf5c51799ad
z4a0ee81e4d32895743ce1e095182f74f23bf725ab2dabe09df232a7f21f7e26e20c80be8335e01
z798b227beaa9d1311f89e1443e9a1267cb892cb4dfcdda8c6591b78354caea48d1273de3ed9ca1
z4e0b1ac147566312e0ffba646c156f75fa9e220097f657ef958dd9abe922473cabf61b75c0b018
z6b14e97477ff010cc370bcb2489f39355d29aa4ad54168416764aad891ab5d6cbb8e399119f372
zdecba51dcae6593e03c89325168b679489ac2ef8b05ad389f4dad1215bdf1377524005658e6931
z001c1e67b89baa6260d5bb0f706a0acea3ce887d630fd66b489b7c17387fe3801d73822ced7079
zc7012fa653ac187034dd71065e8f4d7f15bff6d0d921dea707f19b4b40a54a6ff0e9b95116e55e
z0a3acb40f3fe9e769b12e9544301bdd459c0ca8f37187a922b73102fbf0ae8bc0c9e88f97c7506
z295e20c7272d82913d71d2fd604765d9fff7ce09ed1b1de256594d62dde45d12ec6baf06f1f455
z2badde33ce410338c9542d754f76b4354770428286c31fde8839dce81396668474a25048d8c91d
z25618b446d5a86d024fa2ce6b3593cd6a2dbe71ac1d721127b77229c4ccc0f37d5d0a2e6c79be9
za31fa88565beb02db5dc3b202b1931dbbc45c8ac1ce991ec27647f533bb48eb9a6dd84864d2e2c
z47d0d5d7a4175f6f14cda18a5365c97552e30b476a8bffb218e610c7c92107035d0030ffd42a73
ze67f88128685fe3f610a4bf40b8e56092b8618daa6fff48713fdb2e33b33e6c9594fb994570ede
z9366884df0989488012a231666dc94a8e045283873fed392c0b012dfd5cef467e48dcc49a79fb8
zf634ae20ba567c37ae31ec0259908fa9afdbf16f3ace3c871fd0d6b155e818b7d059517f3a1583
z91fad0644aede6e253733160dac7a2f048186e7bf4164e4ced7341dbbcdf601f530e17ee74351d
za197cb5e9a361ce68482404b398c47a77be36e3a65c17f47ca55e3b6ba87a77a524730834326a7
z1dcfab5fc2107ed290f633cf0bba5aab23adcb1e1749a5ab5762742876cf691c3d8d5e8973078e
zce312a91171927dd8bcdc92c4e685ab83e467c7c0d7e43a9ad29a65415a55c8d1b77aee6c50777
z273d18f1ca3fed404f72ea552738450539cd8338ae1897130a52ce0b4b47def080ce1818e9d92d
z66f5b2c138e8f28abf1885739e3f1fdae533cb49d088d5f1adcf360e4c6d42e4cc105656eba81a
z15768f22e34ee646222e39926bdca63ff2eb434529398635c8a72233828e6273de5d9c7a457ff6
z37e9c06462c707d1b951c3c1319c684696ba0974aa4f314ba3629dd293d1fe8cd64523e3631ccc
z7f824cdcf0ec42dd3ae0d984a3dd704d33ecf512aeb1bcafe2cb57f7330b68066bef285b903f2f
z64124a8d6ea8f1a48700aeb8c8fef0a3523f220c865614352b3ca5e1240a5d5f1f54c56759dd35
za88b36d9d72c904db7ac5ada1a51dde025c690b1cb8eca3af6d3946f7eb2cbae500b90292215ba
z0ef18afcb1b5fe1c6de00046ea07d4b1117d9bfa35ce0ee4929b2293080623bc358b242752cd6c
z34f9a1a9e4a1a0e78e129a51c840e366a00467b7f3b90f493dba50a6786422d73d03b765dff976
zfc630830425a72593acd45e78e7da0ef590de80860164b6d9129bf57fb38260fd6d554bb5dbafb
zd03b3fc8edf6ee8eddf7dd03b95ee070db75d32f6d720001aea3840db3ed1de58a3d95709971da
z6be85c8e9c8a9378cf611c578fe55983b6c32a0ed0e15c3ef19fe294e29cf926b03ef2229e99c0
z4f342f732c06ad78ad20c40f26493a2917cd9b0c603d4a9dd0da73468a06494662051e2ddb6134
z8b250afe4811273915dcca13d90ad44cf6157c8834e53174ebe308830df869c95f004ccf0d56c7
z73f461e14352faf682677ff0603ce3d2a9defe9c7b66a79b14e03437370c2760e0184b80c38ca3
z127e532e1159e131b0c20df80ee83d705e3772e17ae62ff606744a9e9794496cc9c73c9b479684
z46bb8e69337d3aefe27dc6a08a2ccd16017f8952d85d064b2a79d26fa259a42aad313d2f69f7c1
z96c28647adf7be14485fa2de51ce6f3b1d02337235628e8b0bfcb335cef052a6b63fccbbd243fd
z28800495a3ef7f690b8994d4b178863f99b39f4c427275a2339d7216f3b1259f75829c803c45bb
zce4c6d929166df0852a6d0c74fc4e91a9938536ccc0bfdf22f0f97e939d36d1233f6d6db15e32f
z6dcba0f1cb518afd61fa9c79d1e4b77d7e98fc269792030ab54ec458c49c296bb4c659e6b92a2a
z660dd7b21c6ec7b9a8d87d4d8b6d6e2b34bd5788b24dbe07e079ed0496d182b13789120e8b5627
zb64f7091d186d7409d6de863ab798e79fc7a3029290bf61678a4024c87e5eb976e7fe862700f02
z44241dabf1784a7c116760688100441794be286d6a14a907b6230f0cd1fcce5ae8f861b4097278
z206a127d99061a45daea8f5927b0984929d4926a7c0fb172c3536bb82b600731aeeaca95955a99
z07587145fcca3430bb700eeb30604aa13e7e7876ff98aac822602d78039c1b04c33e22ed15fe9a
z96e6c21afb5b06d69f5ca728c74841718b6f954a25505c006df28f9d1d54a95c227ccc26b65cb7
zcd049aa3dcdc0734e92d91e05c5920bfd6e731f74111b528bd682f6a3de727e00a752b145ccc96
z103a4407090ecd8856be3c7d5644a498139c89c46df4bf1fd310dadb560b5510de9c9f9de98832
z5df43cf5bcbed9d5878c48b774d82408777136239cbdc99283fc90afbaa31f8c1f92113d94e5a4
z964ecfeaa35d8b2f8238315dfdef9441db1caf56c8044d12fae9b35c2d4f21c970b321217c05ce
z8ad7d6cdb1866f26aa2d5b7a3a98d194f3054d251de47785ee9a971d4764f64478effb2185e73d
z548f9154d6282c8a65fa38c448e8eabaff5ea2e8f04c6941b7111c57ea12197a9b38d0a9415372
z8256d75abdd00f703db96f506191f0c061e53cc432a862fafb86ec1fe9311c6f4fdd4ec670e9e5
z5e01d6bf8cf217ecd000a51aac59bb85d27ee541d82307c70da16bba432c34d56bf769692913da
za43daaa76d982217091e85dafef8b629c023dbe54b5df54aa163a1aa1d3b16c5cf40f64911f684
zddce4b59c80f4a9b5c60b75f06aca5470632087958c77c59399740b1db19680a9c3783e10f3f41
ze7888eea2e79585764a6b5bf96783d5323a92e099931c7a1ad692d7be17999f154bdcaeb94a6ec
z61dfa47ccd959fe022afdf2629ff9cb3836d65356d4a9e2a173eb23e1c03aaa96d751c5e81faf0
zfa21bbcd12c2fbea2ebc37d57f60e68fbfffba1516d348b5a12e2ee931a49417b8eee6731facde
z8c012a0deebb5ce6248b055603e5f707472b4dd00af9f48e31746a805d3513d3c95a170bea1783
z69263ac6ff5c36a4020447e8b081e9e70ae574fe23b4518bfce38d8db60406c82e02c72f91859c
z77601dfe478d26676144946e5492d20d5db6054f342f927d1f1b520418dcc806b4b5a4d74c4dae
z05aa178ec36f2e43206cb07894daa31c23b9f4d86154fb21fda773654b8fed0a5c43ffb7060e7d
z41bffd4859eb30c1981346c06edf6b0d9358aab634d5fe34e75a3a28da3200b201ab20faa6e945
z0236e753956aef3239c2091459cd1c39775d81db945de2cdc9aeea4a63326c5eac8a51c40167ec
z1adff46afd48532b68a8793471d8a79985eccceb254ed24fdeb520eac4c2ff431d0677fc6f326a
za78e01fc72349abb25fd2c90a35e5e95171288dbd3266a601a5d93e53d3c8669b8bba74f834c6f
zac3e0c1f90eb50e3be4b020a18defd4b2469ee42db58fb0e36b3cb84e349265991e8f7ede3582f
z39a475745b26529915d40b50d2b3e27ba24388d507c192cd661e948b6851423af0bc8834a3fd2a
zb26a4197d264ad6b03e68752b71776c14c49387ecf5116add9aa9a4493e4e5d0ba890e9a003d8d
z32c4187b481a00af61f5cfb166b9b15bad3a6f2ea9d61c9805b69555730ee0f4833a784d967da9
zfd7b2add2fd8b18f5d481011083b4a34b2176a972131230df592f9bcb34fc1a521e7c3c4cee38f
z69098b140d2d2760715c994d0887fde39d05babb04f82fc2912736478a5a6193a506e2586081d2
z943c59145aff9936096d627f22691993d6dde1812b255c6164932a6e0c21d8c05e5cf464093f1c
z288b0ed3e500b01b3c927a33a4c4c78efdaa84d9ccda9bff0b490746dacb21cc15184b3b24dea7
z15221b84d48397bb8922b2702a2265f0358eb240dca47a2e5cd94e6a9cb28286454cdb57e8a058
z0a90ab0d9194f49af0756bc395dfbce77986e667c3cabe2a47b1680cbd153bb359602403a8c8e0
ze7ed66f6f163f1e3a7172e35d0c5c909750b93f5856148d74d803333a5999a32e40baa6524d9bd
zdd19fed2741dbefd2b1ae180ecbd16217fd3912c77dc1a277a726c6a4e1f6a689285b37da7e198
z58e6862e291ef829629abce9a406945914b9c912bc2015c0420197b3a524c0bf7c7300ab50ed64
zd68e487d9af26aa4dc8055e857a89ba69313484c2ee3a52afd2d59c6e60e44a884a58b0e4b177f
z9f69c9910b56229a3728fe57f5a7cf0dc552286fdad087c9e8013194ad3efcc87b9af6b9701f0f
zb5e6cdef63a1db97b52f3f641e49db17fad82d2e2cac4078680b5d36d84fc0b0930ab3c3060dbe
zb68adfdec574011bfce1ce2e08ab71b0612b77965218d865c157e112aa5b97cbd4093e2949ed08
z8ca81f82a06ad02182ec1b9379256a837a17f340ed2b12ac34a7e88d9b052c9f34b447d825ceb9
ze6800ccbfd0edf231459336411ffbca82e3c6a503ec11803c4c51a98fa19ae2f16b3d2d6c5fb95
z0a47cb80646caf3d0b09b3bfdaf64322c66edf302f22bc91e42e1482e6d6efcf484c8148614957
zff4875fb77fc5f659dec68f1e934fa48c3b9ac1c4d2ec102109be31c7a104ca7348edf236abc47
zd554591ff9128a76fd4cfff09c2fa3c853e805fc01d4ba67c78dc666e2f9f06b5aa884e34c1dcf
zb0f97aed2ed0218e467da8dca243ef6f24b58ae410e714d7438baad572592e92db376794dd359a
z9a614928684aa90757ff51fd668a320ce2bca6c93049e9a8f38439e16dd9d8136cb691dfcf0486
z9320133ee314e5d502f20927b65ebe079b7c303f3ca3fef4948f0258aad255c51e4ea4f32fcf8b
zd6f23b011dab8a87eb9e0233566d740c101322f8f39589e8955719670fa0afa66155b0fb1e7236
z08f690807ea54c36639f8ab8eceb0b620743bb040a9a97ec4068399e000b090002e347f032b4c5
zef948470974b1b61f4d0fad47975b3d869ae6496352dddc8cebd674ebd3dd2de4709e2a2689bb2
z496fd98c18bff9c63f3f2abccf4e1aaced80c7b4d21f2467c5db7c109a76ee1af195e17ae59b03
zca5e3fbab570f1184ebf0276d50f7a907cf7dc1bc92fb68e273009487a725eef80345225061d7c
ze062fae073b48057176e3ffd53172aa8a6b6d521dd645f8a7e6218a672ffaa9de330e29e2f81c1
zb43e7d2378d75632c5d87832edef781bdad150647210b78394f76e050defae834aaafeef2b17b6
z1ad88eaec2dff1bba54dd04668b59b06771425da7ba4ebb230a50d81a2e98ebc260940c633ef9f
z590e8f4a8ce6792d65c6b9c8189785b150e5d4e58efa90afb5f5beea1f81ba891ad563fcac0455
z2add16a62bae8b344253ed3643773e192cc0258b004f5a2edfe045fa01cc346859babfb7bd3024
zb7103b27b51d4fb5cd0645ed45054f9d8084a0a59611e5aff4eed248973d18b49584a741ee60b9
zba746f90a5ad2b78a1da8592500a9a19386d778d00912200cf37b06f7adf7a2f07b5ba6845b81d
zb33fea08bc179bbff377aecd273f88434c861ed3e92d75edc4888b8cc933122ba088229c26a1cd
z9058f5e8364c7e88cc691a3702af94c6b37f7891fd58f1f54d61caa7d3094e8d1564b5295a9ac1
zcf44387ad504132f856bf3080ca32e7c31a18c241afc5529e1f1573ab1ea3423fdf09c72f071af
zb3f1be6ba90535f48d0c17aa1760b1190653f7b29cdfe3e2112c66356c17cd25240456b49f6acc
zbb4e9d9f0522397616d666d0b645f4e31c986d2c382cd58616bec0d7d7facc225bb23c2d17a2a5
zcbb50deac525cbc24e87d87e02a1f89ad160760e720fbfe90acea75eb4dfc6cdacf10a21656334
ze5cc5993f062633069449021a299716e3118764383406696701623f929173bccedd6c9df74740c
z168ef51211aaf0ee80f196c19843594e151875f0198e782cb3a1a331060a82e7be6e640732280c
z5b56c635701476ebee032b847cc0d8456bb035ec74f462c3ec724ce200593f47ccc9e2a2cf47e1
zc4edcbc5a4906d8d69058f9ed758c763f21cd32bd872ea3e6dbbb2bd398b6f7499714b1ed15585
zc209e9d04583fe58949569d62c54397b2d1fa78d020eddb8d187553476834447f66ee8d30b11d6
z56c0f69ba3b131a5d20ab4964b78386a8fd8f51cb4acf1109cbbb7096444a6dcbcd5c6b6f78973
z9648422531498f707b7d1ed9e75d3a90fe216f507886ac921e150c44b5888318fcb77d76581935
z0c66e655a8907d7a2e19bd0b57eb1c6327ebe98700409de79d353e7ab72d4a29ad1c83d75ec1b3
z6f1921ea2f911f428d457968eb4b6be00866674706457034807d10a6bc7cd6a8656c4ab04cb14a
zed9b2c6d00edd37279bcad9c303c9d1ff38a88811650979cb54bd4a1884d5cc535d96b9adac6fe
za871037aba13bd6469e70ab88befc054ee116af8fa04d0adffad7e56e148bc8b369f241c5c1647
z7f61bca7dfee8631a1d8df3528fc220272251f6d31af2a4f4da79d485357798f19731fd42c447f
z783c89f6cdc36b98bab76b60b870dc3cfc0b9e8c76b9cfd9d28fa43e83df7a23082eb4d3376524
z751a73811b5b1f6d55d8d1b88557dca2d4f12fee24733ecf4707bbe6cbcafcd6151c7af9ed804e
z246db15a7ecae197491ff96c9b291558714d20853665ebcaa779db287e33216620fecd641405e1
za937c59c012ef9d0a5d7f71a6743fcd45edb2c5d47ea4165c182da362e25e64c286f8036b69b0a
z3b2c79ab04978b3362ef875f84481df4528a6926466b015fe71d4e9f60b90175c116af40941fec
z3a3893e22c954434222bbef04743e1d85acef748d8c7244345c53e7b147b7d33d1b5d57483ea62
z43049321d191e214f13156e7d2939589c114e06b93550d92b0176c5c6476e67e482817708618bb
z375b5ca5ae50f09dd585a3dc4fea0b677753a7492403eede35e3573f0672fd5c4c6962121cb155
z0a08f6458b2df92d023f6c7eee0b9cfb4584216dec46bcff9dc0f6ba5bb34f3152c22a8ff641fa
z3b7abe25dbfa1e8f89914eb2027b95d5765aed6b83610eca214b3b845ed1a546be8df5d71ebe54
z482bce44e4c562bd38b551a9261a6128d34abd23e5264351732ce2b5ef7d6dd620ebb1062e5aa4
z257fb880f9cd3093691c4ddbc43d3567977ab64ef62eeecd4fbc42938d558a46b8e0e73b6860df
z6e1825c1bc99fc687a23dbb49785d4e5d708b713dcf58b7ffe2b8dc080d1d875800de285282997
zabe4d46b1d298ad2f98cd92228af77b562d264d6b2fd101e79de5cf157617ba9f0267ca2548918
z0ef308032398eb709834d6db8cdf2654d1f2ababe04af17ec102debcbee41d6de3505a70d96c58
za5a27167f72a7632c9be6460741ea8cecc5584d5345b12de0aa6f9b0ae76bcf82e5627a04ee774
z66accf74763677e1d0d80f33a8a68f6e3b48e3d1b5de14eb7db72091ca3398121c006ec21e23ce
z823015d4c99b3a40010a06f82b202f883d1385a4e5d19dc58fc606725635bd2b18838dbb4244d9
za5a2c7cb5c66aab22ba83ac84d2fd50b7c547d76608a6434bd5657aa56ed039b2e7d36ea988760
zdd2c76e00afabd91b59a3064f8f51f3d6b79ea4f7802a8fb17b96c6108621f056c3bf6729b5174
z601eb104c8e07cd091c390945c798c248309d87f09d5e91222b6f51fc82788c434e169fc506e16
za61ca352cf5ccfdfdf917745773443692a761287fc54e6ebf4772cd87038d71d486a53e226b5e9
z137e78b508f8f9cd54b6355e6cac032bb42cef7e3c60100511f997efae0acf0e772158ff71186b
ze9b493e69b0071af00430317caf8ab2abbbb853e18253d22ac3997cb4d21d0e5b52998cba1697e
z1f061face6d36db1bb75b46dc7bfa814a09af0e5ea575a90b9547e6bc8fcd4c2dfd814f9762544
z30d25143b6a4c302b55cc4691313c55395723f4c6b5d5fb7cc8729aa632c5665f5398a19655b7c
z2c6c477b093dffc917d62fe6f26baeeb22124b9b97d89ad3925c810345737d9645fb17a4920b0d
z620544aed2e69d558bd0943957ba3aa7a1d7faa2010828dfb7f012c27b7ef723af89f1306111b6
z0821bbc10f292aa39e66a8f560e57fb54d6214506d2bcbd561c83ae7e1dc6d3db0c9a28584603c
z3a8c52ec9f39edc3bbcfc4bbd06d2afbf65b98408826ab216e24e7eff8a06f9c61b848f819dd47
z7f99b50ef27593002481aab0cce9b0a7d208d0cbf85864cee55ffef7fc53ea4ca1c88afbf81d29
z6e60f05c0d0f827d47b98e8e389d118c5b0ff5470d83a2dff342437350825e2577daf86f775db9
ze986402533c5f37c5d791ed1a6b8e8823f4681b79055495fefc11782851f79b4dffedb7533106d
z67fc6837f848d400179208326827fe758a76b49800fd3d7f851064489fc70aaf59cefbe1b4f45c
z37420f52d85b1ef618c7082881399774173f65881a9c4e71172726a7bbae356249b101b3f72ada
z6469d5dbbf8376dc3f91b221361f599eb30182e0559bdeb04b1117b2cf34f3b8d5ed84c019d9b8
z9484a2d960ffaf4bd3585901abf6c86fbbb2023fd9bcf5526b90e9018d078ea76800d2a31fd87b
ze7c22d917d91e2af1741a4fb2188baf85256147f68f664e278291e93e408d040ddaa9148077f92
z5952c6a9b08fa873b256a3693717b361155ca74858cc353f0184791720b56c39ae313bf13e48a8
z4d588de4e99989534269c69ffc32b72a5ea12eb27c49d870e593b53ad42e126c2417d5eb0b2777
z194990fded1f9843286acdee3cd68f2bde3352ae5824464423a0944d87d666b838d33504aafabd
z868c5634b251c95d5ab0cfeecf9ee6bc9a5b58c181ceff6e1cc52ca15b58ef0ddc9d82c1c6427a
zd4a86fa2cafe2c9c17525fb83717922ecddf82791deaeb2a7b573eaf6a5689bcf39c735bc6be99
ze3d0e85821f5bcbc8b4efdd3f7a294abdcf1e93b63db8656340e0395b2ef482a0d0eded0389d0e
z85a4b623a1cc2126d69215bda229fa31c738ac7a2909fcda40e674f2b837d5ec2a86722b6f4c76
z6c59df129e7b3f0eef7bc2102f9dafd71f700f1482d162401f0bd5537aca96f144e74d269a52cb
zc1bc5568a70c85efc14082e2e42894f55fcec00687dcdf4241a1cc9094d60f29a877c3bcfac0c5
z97f943c01f64ca62df85325528e938d1d726dfff9d8031fb106da924e1de3a90c6b0943fbd7c39
z4bcc2ae1136beaf6c5b44a8237d08fb2ba024d92e52b14bf6980e593681925b3f6781965d7eed2
zc5587fc00a130c1f8cd8f5bb486d374cb77c233686e5ea25b3f6e2055886e08e0a3200b54dead7
zf51c938ca5ec07846ebe4311fdd0396024a92cdc558c0098bc610e19dcca6da7f9c4166a388b3d
zdb2f0f7df018c5949eb0ccd88e8af8153d6896d0d7fd1ca6f6c08236657ff9eed4c6488cc3d27c
zd7d722b866351154390f67b51dd0feefeb756409d2647a1dbd2f44647d1866a7a43031a1f60fcb
z370c5909b35f83d90c70b357abadff0c79f2642bf5da22735e85b5214b47834881c4e37b9cf40b
z225ae2b11d692a90c99ff19d566d999064d1ba4d0223fb521e30e904465c81c90a7861157e77f5
zb4e121ebed01dbfe635b5a08633503318368e63daab4796e2679b87c8d91c05103089c1bbe6792
z56f47d998a7c063b1eee98d1c48f525dda792dba016eb394f58da191c5f8928af7f8af1e09f487
z0aac0015049eab9444a3185e56f56fe51c75f9fd9aaa852e4e2d9c5127c864002538e0cf048d04
z2dc222b6ff2a6a952132d1e02546b960331b974a77c2a5f4208e606d831d95c827b22cde70ff71
zfca39a762294d82106ad8b8c2665e45dc381a7cc77ac5f3a6b7fc89b288b2f8d4e7042994da6dc
z4c95ffebb4cf9008bf06e72b18a891a8cade20a39da2fb7ac60c193bc9f277e6873b5a6755517a
zc580bcde3b7e77b15c90b4a7346674a605c9a027481b24d17b22e95dd4bc0f9d729cb8682d1613
zfa1cfd45ac1707b14f83985260bbd7a4e929ff38cd481414e5200e1683d3e26af3cf31b8e8ef67
z479e33d722ff234d8fd6ce38022707eeda66c70d21cb4122ee8b5c5b5e0f6f140536a255429bb3
z0e97acb1509cfa7eb4303ef81f39650bcda920054e9d845da8b09c895a4ef2c6565db294552ce2
z6624f7bb7741b737ff95d53c595f5a2aeb2f93a0ad2ddc1e469afcf8607fc9ef199ce6d8fc9a76
z976b9fb56989f22024e7ce97c73c2a385cd1fae9b936e0d1e44fb6834fe87bb2f56d7d7f4e808f
z754d482a3de180903259bb4745518f9fb2e9d4684660fa07e86cfc34634d6bfe8e1f8dd615eef6
z536fbc421db195c09b16ccf4acdea96d3e45e58a55d94011456ae23c4ccd2bba32dab248cbbf22
z21db94ae53e3f19205fa19a67f532cfc780cd3a78abfc396e4f8f9d6e229625f573163c5d175a8
z82e5ed78590f1a4f262135586d599a1331f27dba075b8fe70eae16e35062297d14a27f1a54ce41
za04606df5e78d425fd5cda13ae7d7b3d622d2f366139f59e23563170afefe777a6da40a9cd93d6
z8efd236076d6d5aed8ad86b620dc823259c70995ad3a18f25a0c5931b9ef7bbd41caf996e01e8e
zbd692e4646c44ce53082e5f88247a45d2626b9036c84e219aa25cc4d4d971c3565323fdf8bf2f7
z05a7a75b92c6cbeb2dc5211edb5dab26e099511004454eb1cae397d9df29259fba50eba60fecb2
z73fea581c7e609b8246a07b1597ee20b6138649b3117c4d5f5856e515f1f7ab85eeb6a6f287454
z718464b1ff6ef634f577b13a14b8a2e770a5fc1c61b07539cd3df526a4cf9a33989e5b25639cd1
z5d2adcaefe896a4cbf4f4d858a0e8610b96ff3c88e1b5392b9c5d5bfb1761a5c1b73d1a67e5955
zdf537426f2a481f83fe06bfc9a3435722d49286cf073f39240ec03a80165ddaafcecac26f4acb6
zf3d8789b2f0300b6c4e4822ee6b705cffbf8d06ec3854cde65b3cc81be364256bb6c18441dad52
z7acbe27cda46dba0479b8bdd0f7460ec9d873abcf760bb5c3a299795ac60a6ac5f7c8e0563fd4e
z1bfeb3acb586423112498c7334c4a10a516913648030a898013c44fa120fe5a1e84b9b763747b4
zd3fb2f29afade436d00882e0681821439183afdc22ac8902fa944ad205855cb12f8a3dfd6d4c88
zf5eebabc18918a9825ed95662fc79422cae87ee6748e118a54203a429629e5ac32a1dfc7ec14c1
zd0c2f5158b1adc3c190a70861deaa606a6228a814c8097164f6aa8b7fa3f8fb7f7e019724412f0
z17735af5b8fcfa1d22ac3c8b32cd0c35ec69a40f745f4b07057d3e9f01cbde6dc9579ab5928c8c
zbaadd892455aaf186f9a932885d8bc5f60214a61c655c71cfbca880f1f8f32004a1c5ff4b71933
z9b7843d232d36d11d62da102da0ac6eae1cfbaf573cdbae7341b0cdc94418cae9092c276090940
z1813b95186e4a2b1867b576acb2188c15c36f7b9950099498b11de0880c1deeeb9aa3337f0c2e3
zcacd3cc63acc2d6718d6e8700b72922a50d1ea8313d5a8c6286c6e0af669039edd893d9d1ffdb3
z70906cd8dc0cfb9312251cb5d6711364688ee1f2678d8a333647765496a97009c961e932002f4e
zab046b034526734afa835613c6a0f635cb4a596bcf9ad274b775a831080242f43659220f558aaf
z7a53bc8a841ea3ea2eb41fb727cd25c5b02fc45d3ce7b24bd2ad0bef577ecc2dc1331223c0377e
z2ad6ee81ce1950a90dc5f252f830afa3ecdc65269b518e6b72de74a326439ddd7340eb69de0c70
z1468458c146fd24ce75360c27c0b3a8d71773c82e791d18a6a8674d9bfb88b4917b06b784d6b52
zfb55895cfdbeaf8fbaa031c01ab3b540f89172ed7cec1abd65a00981ee11bd66b2faeab14913ad
z8795d6f3d53b07e954e04d97b20830219ae161693c204a8726c58376c842c84796b91181505480
z58455706b294125eabb4458aefada1988546d9bb2b650deeb1fe51f98351dfeccd957acd168727
z1ccdeb343177fc4b879dcfe007ca6a2cbbd972435ba212b34dc0c2d25391bf0e39a8b96a2d912e
za145f938ac4b95a8297cb101e51d10c0a040926a1939a4d2d51318b0b285b28ba16b300fc75910
za024169a8e2fc72652d5eab5fc657fcd502ade29cd20f637c66ea85a8342e674b8c93112eb1f52
z1502d8f6697556e08fb2992235b646135aa2f343e43dd8586495311bc26ac271265b81bbd1cdfa
zaf246a56f44f7ec707fe481d8ca11e0dfa8190c1593068ce5a370b8498d531aca51d29aabf4d21
zf621f1ba9f8ce9470f99d4dcf98f3f26d9fb8d1d673faf031ab306aa2c1e672b96eb026cd677e8
zdf0e7921b71f8a0d632d80ae8e3238645a36676f0899f5cafa4b72264c42133698ddd8501565bd
z233c95a29183c178f9575a2975c1816f9912d643cae64b480d2502b5ca369558606a8a2788c496
zb774c3568c771c6e556c964e40a47d7c8b11628a0686f2b0adc2755e842d3743dec2fd49010c90
zb3e465eef57fc6685f11689484117190b3b10b1b12a6f04a90ae104f332a2091e0322773661be8
z2ecee2064673f57a3e512a2bb6a0f135810bf50529824260a0a1e031da373bd921c8e01e7f14c8
z93321dbf7874782aca7b660d35fd12be4f05cbb92e84f2a1848214cbbbae9253b9d67337ad8cf3
z3485efd6d7f5fdf609eaf02511bec07f62043f8a0a3d1c44ecaffe308bee0fc21f815a93008cbc
z9bded2f3623980b55f500b3ba254e38b0b049b7e773e5262991e54da689d3ae69687822ee658f1
zfdcfce91338df7569c2cc321e37b4ac99b70bababe269f540585e33942d1a5dd619f238ebf3e59
zd1f2f72d2794a2a20b098c380a158d8dd39772ebb4beab551124256249ea1043bf4ab2c4497c5b
z96ca56edfeaed902504049169ce4e6d676ff0e870115894463f0b102aec5396e9f2d73309f79ed
za5a66e4bd8f60fef45ff386b609c234212c1182ecab079ddae68aba8348b9e1d81915a22b4f4b1
z3072466c01b094d31252dfa4a62e72cb45c03f1ef7152290a361bedbc704c7f430673d443ff9ae
zabfecd42ca752494a3f342bda7adcf4c5c04d1d2cd75a3991b262d18949fa11c363f6f19e1e922
z25652a40d4ddcd8f40ffb016fc244de2893b0eed8b5ec55627cb011ed8f8e506790e99e05dac31
zdf6db59168029ccccc0156d879206551917660d4328d073044792871ccc0400405b2aa3749c4aa
z29ee99708b28f271875d5ca0ca971a8fcd0996ac6ff3cc133b9f962fa4a13d6771cce6707c31dd
z71f3240561e651c801e4b2506ef02e44af3f6a847eb3c9961b5793747f28cdab84f67a8b3701e0
zabcd6e47595ca257fd3f41e57fe41c676e5557577d47dfcc146b9d1bb33857f0765f083b55a73b
zfb3e7e9f27a98fd1fa35f72685ba7816f89fe7bb563295cadeaa2de821dbd65885c4665947ba00
z7a44102e1fdb23212ed6dc12afc138dedafca3caa0444e46d6769eca21f9895ea35b126d52bc2c
z91182b091b77e9298856bf1f9ebd4e96cd2d6135687edf0f9d97a4a71adddbc64a1c067c94b8ea
z7b3494e425cc20a9b1d4ad3f3c98529efcea897a7fd643889d6d63414b81004f3377b7e701d8ad
z316e3b23d5a2f0534ae45dc2c36de6df1de72d2430b07cbc0970d8009cdc37640adb6a26fbbfc2
z1aed70ed19d05b258a2e4c4d9d3b99f29809b992b91b260604957550104424424a2813ae2187be
zefc5849e84a8916407c959e3a7dd938c045aa95a28e96387e70d419d54fa260a5594224fab1887
z308917535d6c8769c2ccee21ec74a9aa0cef09b4c8f8bf65f5067038a92a97197de361b80aedf8
z1faceaf9051a843d69a381b3de35b9b8150f547ef7d46b05cf0b91b262c7bb253ff62deeb006f8
z84bd03cdd59d07b6d4b0666e6be5f97965650372a19be125a744164e5d0248602c927184daeb5c
zf0a0647b694c69a302a37157082f871b8a4ce96b69d49f8cdbc734e1f885804d06f5990266b18a
z9de3195188ec01bcd3d58df6991d6372802c5ba1bf2f36a96c23c238d232f25f5fa47e760578bc
z3fb745c9fa2126f64c495826a8c69090ecf00c6ced1958693ed72d27d912348ad54af02aca3bd0
zdc4ecb668327960b3869dd75988afdf45a8d143337b825a6c931a9c1b2f79f46566f9feaf5bfb5
z641de42cf18b616079ebec1c83514fbe50b1be7186690bb3a9077eaa7e5ee53dbc6ae4544b73c9
ze9dcd4dfe16eb3719431f26fcfc41f96068004381e27be5f59e879a778cc7058a75508b2785709
z17d6d17d739f20f50ec1d60dd62fc163cdfb5dd8b77c9c4830ced7e1fd7fbf8192ee47e44e2598
z6ea2dd45eadb54ae93332d6dbd6b0334b04fdabe7b2a7980a91196baa8e3d52dc882cb7ca01ae5
z71eec08031b95fd5ac14f708a6298b62990d07fa4920786941484078c8785169a2b20063da53a0
z9562b3dfa6e64637d1c3b5eec9dd8bf73f1ed77ad9571c6a9599164b0ff74a17cef0ceb518c2a7
zccce13c4b052f55504889f27c21a8a5876b58bcb1a2bb428be0eeabef9d48cc81e72a443cee493
z72f7a5e0f650ba1cadc5e6ef20decf9f57433ff4e08b1a0889c80eaa932ec7942525fdc48bd40f
z221df7c427efd553726f911788f41256cf8d06856fc9b082ac7edba0f7dc059c91dfae0bdbe7bb
ze03cb2b2bea282305244cf015f8913600ffe1a2cd104f9d0fad01f6bc623e3c420e4bd517a9254
zedda9bf7b1b2d0067c427d4a7805ab254e91f95dc1f6d84c6a6118341c5131998b05c51c48b2fd
z47e8e5f3717aec21062e4ef889634a3f27142d093abce744d3d89f5f4559f8e7e47580cbddffa1
z1d18b93b3e5a67fc9faaef93c6426cf26668f3d931435832021e5fd219def14b0f46442bfb226b
zac6644dfedda8ff47fdf8efe487dc179cd3b96215252a8b127b10f9f8c44fb468d711400d4fe1c
zf5bb39567b437da25bf29dcb2b221c04c7aca0d4948242ac85943c11c935e7a349d031a032992b
z1bdffe5ed537ee601bf64f0c6ddf6cfa25ca6fb98d9686021ee57c2ea6fd62bae05267e2fd2ada
zb0d11fd0d22ec094cf66b6fbe7eb61e24ec787afbd5f9a804562f770fdd95e7b243d59ee93a54c
z0b8a62bbcf2c91006293e19116fc6d0c49c498541887a2247b08377b27242cbb4cfce84085924c
z4fa90e57d78171e5642b2b7e1650bd0fc95c36ca9a37018b115d17c9ae8ed5c20bd6b6a4e2ce0d
zd18f6df869c086dd0c6f8dbce66d5263cf380b959c02fb85b4bd33dbf634e67ce969cf573ec9db
zdc19b92df185b3c279dca78352d00834bff1927a5367485126a03e42a6c81292c6ed609ebd949c
z55c655a8bf920f7df9a80a327b3a1711a7aef483cf1eee74c71781dfe69ae96363e6934390e2ed
z5d8b10d363cdf8cd6ebb48a00d77b06ec9fcf2e7420d8226f738690e0a1d07bdbda5d573cadd93
z2d1bc589dff008961ccbbf4352820a452d4e6ef357a1f7b38d2cd2fb0b226b6a4b2e23bc642464
z18fd276689ad7cd49d0a222097bc1880faffc583c8dbb9626c7896c2e5c45ae4feb94cad45caf7
z20b04bf1dfd68af5faafee28be678673d3906bd7cbfc40ab18eea0be2878125d21fda26ee2ca21
zd8c743ac69599194376bd3b9ba4fe57eb5be1e5edfec6fe8c57d69b05b2427bcd7e0557b8302e3
z6d6c885242d6f6e4c101fa33a1e253fb7a927eaf8862a2c7e70296140f230acacf167b06e524b6
zb10163beda84f93a96178d93edca8dd8d0b4e5200c8bff112dab8ce8d70893060599eb888f7c10
zf9234ade70ce26f30b2c5f9d5aa8cd2f627acb53d833878892ef6affb9d738153747deec00fc34
z26382465fe4f80246b120f9d5d40e345b7610dd2b1b0cb4ed9c79385ff69ce28d155651c1523bd
z1991d6897c1ea4964adde8d8e300ffea36739459e1b0999316e85d34952d8ae2d1f89e36e4bb5d
za060af31ec0b84654095fc50e0769329b0596082964d5878017cafecc29fc9b2835aac8de37b10
z598abb137e10fd7ecb29f890aa924d0174e968d7529d8195a2f2a264e7fe0abcef231ededecf2e
zc3a55822d661e891902d264e622d64bdf8078f24715647f38715b3a04442b251dee2f43701477a
z65607108ca690c017f36e697d85cc17df002b9ef01d853fcaef0470b54809f9420fbfccc54027b
zfcca7dd4a4bda83c1c939619b46104645e8a952eb9c57b1ed24877d4f9cf2a6834810831086c31
z827dcf0db177816f58674bf70c9974673e4bd654cc192029cf7587e7d7ad85b7545b6084489486
z57adf3936c019bf8340b592a9e9619a571e467c015c18247cae3df4fc85e4a3db779e9b30284ae
z39d91ad181d2dec2de22994addf3260bf98724f2a617825ee63a58cea41308ad2ff4d0d8c90ea4
zc2ee6d690ed2b657003ba26f86d025fea521fa2fc317012ad5298d41092fa5e2819d9ebb372427
zc4649982fa151c6f8b0d7c5610c6ac1a0b0c30522ddba25c80c5a965a6f07fcbf32afa9492beff
z686ace39c1da1621e13aa0655d2321f42a216179626802e023e696a4a7f3a4994f7752575db95e
zfc2ed3f290d9d79cb383f32d5674f65cfba11293f82ebf170146e9be52df8592678ceddf40c96c
zea1084314b04cc3f182aab8addf33d03cf6a5da109fe3d402f48cd132137414964fc465492a5ac
z3e1026233dda609ab2aad4b0a40c20e3415d5a8b5da36febd2429ab6a48e2e864b07d4613ce04b
z728c6d222046c25405096f7631cd2ca8d40e9b9025e587dc4b379b73c1fc20b04dadeec3e6b145
zc074574a2f3b2562346bdbe7ffda13d30875dd46c87894c6fa35be090de94fae0e1152513acbbd
zba18302eb63e87be28b2faa57ee2820da4a83c6c0dc26697bddd309c24fb05763fc0a9fb230a1d
zcc2bf3932556f91ff1248584b0fd4bde9ec54773eb2966322666cb040213115fb2692cf7cc0851
z4c8b0d1e9ea6a2f7a9882b61d0375fb2200afa2aae262fe245f38dffb1967e9399f053907d86a2
z8531899937683a04a81a651f76ca696583c5cdfd84a2d4518ffd2b13efed2583cbca3ee5ec760d
zcc2087fa93b4bbc18955a50a09553b92599fbd9dae18b2e1bc6cb73fe37d4cf286ab6c682b9d1a
zd0eb6fb36dc6c7a604db8077c345df87860b4b899da7caf80a574548334f1046b768e7003ed91e
z3aeab75b23bb6ec107cec82ddcc0f0560d8b561f3ca878d0b1ed96234ef8a0e5b97e1385964265
z176f1e51858d65daa8e97cacd56c1bee5ec6e60c4bb51663593bf7230c12d6108fbfde6a4201bb
z1048f19f1322e218a3f9bfb71f075220a8acfab7f4ce85c3d01ca9f37f473372a48977d9b931e2
zffa4cbb80c1ee90ae0bc4f931033cd3bd26f010337f29c429b5a9cd4b53fc42d150442c779906a
zc3166654998ac754427a8d14364ad7657f7b51bbda46a02c5439c951685f9d8c541968b7a1d15a
z0b96958c512e2af7ee14f3b64e5e6a1f6da4214386df2f050d1b90b32b61c907428a4813d3b93a
z06c741388fd6b79b51982c5cb17492347492d26eabd72dfb5faa7b7a84e6e3e5102ebb8deb3afb
zd5d9c5af6390866ff89073ef72910ac3f075b9e4b8d7ed799feb824b70ecf9795d679d07d598b0
z230559252fd2350c22b4d0f40d1a9613917ef4d4109bbd81c252e2dff5ed4907bcc560d890fd86
zab38a9d8400ed8fa8d6c37555d00001ddd23f8850ce3cdb888c0c2bbb480c3c2df5ae90e293738
z1599d1bf6dccb2557a6dafbb6e58566313f19e815336c5f5aefa4e589e553c370bfe8e4207c057
z8dbc9b5ae4668726670ff0668cd759656f8c44c3c21b03a319db19744d7b8f88c0f97a47f35814
zb4cae520c2b2bb6ac295c2618381a47249e00aee3b9acd576f0efba4d0a07edb0de711c02d2fc0
zdc14da3b77fed57fb499d6f45ccf3d83ed253a0420d5937665692a5b3d7ece010d4e9758729358
z25b3ec388dd1cc0782f2ec71ed41e2e5735006dd9fd11216fd3509fdc75fbf0af6a3ea6995a621
z95181e4a579a26db9dd8dfbef33c9721933715f216f199b84c7868bdf51381f410bf27ecb73891
z393f4b3cc137998d0aa2e99ef40e48c3f47ae8cab368224692222bc7700cc7685ef73e1b970014
z9e9b261044e139ac9a89942a1881fec21fcfeee3aae4f9b736c35389212bb665dca1ab264c7ea4
z13c7f5c6c3071b8dc5424bfa0cccd49b80b562e01809c9564c586267958eeabd42c96f3258f183
zbf760a1e42f5465b6a1d029e69fe1a4ea879e95519bc2f7cfe3cb6f71970481f8a1307b13eb396
z62a217b6cd7f13b22efd4fb05ef119abdbd2427b79076703b4e66dc007ef3ea896210d0001b307
z757c070799a07f8d7b084319e1b943294042012b6162200be24070a724a4fd81c7f894787be3fe
z6bd2bfbcdef14f929b1a442ed590ff7bad1b5a38ead52028e319ecab3bea9a4643f6aa7be67cb5
zb73e5b01e66cd4a5b57c1592d4a9b45069b5acf631549c1db320d2d952a6d2ad44dece3aeb6693
ze7344f08379ea76a47df5f7b4f0d98dd2bad9c276731b90115f6b41fcb65a59349a08cca1dc410
z28e3041d0f3e9ba62d7d2067ee5862121e79c39acdabcc94293515614617dbd7027e8732b48083
z6aed2bdb167874455c8451d97c5496f24b5eb3336868eae2114f074ada11b9b9e3d4c84af0be95
ze2d18df81aedf50e76ad15035dee1386ce9518de3220bbe237a85bb1e1a516d300ebad68feb4b9
z894590769317ab464511825f8251c390b42bcd8dbfcfece25536c6c12a25104cc617901fe6182f
z6a99c166dedb48fe526bbc3f79fc9004bb80915e89e9264ec8dd8b4edcdeb7b71e83c758e6264c
zd95aad54da00a5762ec902758ef1706e7374a7b25d32f7edeb89352a3100505e2d4b9453ca9a96
z6ef97ed738637d5488a2b3dc156a392ac964a71d8f61b1057440a0034b52addbf08de96229cd39
ze990396cbcdc99b29577227f4a5b36802b5e6d647476b68bc5c744e78a0f104727d631a95383cc
zabb0387b66ce153d24d568fda03a07fdac02a2b82c0d7eec1b77cc98ae6f2885f0a2590e4aef75
z32be587e637693531035819352bd2a8af219a8cae02153e7c822f108f4acf9411766b5ac8fa749
zf12caad228daed6d0efc97036a972fcf6cd2632e492258c0d8643906f211cbe27e700464c044ac
z3166ea6f8abcd3473909e84dce0ea1ce5b1970b3657d897d446c60eea5ce270101e0550aa37358
zbb99d8934e8b6c7b62477d3ace289a28ee8780ce4b37f196a9c7b5d68ec9cc43755b5e40f50d8e
z4eb15a4b204ecc20fccc29e66fe8d4d9923181e42ce0d93322d39a959d57bc996545371ca69e79
z5126e79ff384c9e319aa0f91c7e12c46886b38c538a1ceebd3ba8366a8e91a37a24a5645448783
z018f31c840829ff53d34dc2a36732b2aa91a6884b4052d0afc25ffac51bdac56e6b270e746c20e
z474039c54962734412cffec31d7a1c31ca7762dc8baf340d010560e5199f3773c9b6c4510feb62
zad23bf7a1453482395d43777c7dbfc3f87e0c5a52e05794b32ef6bb17b9a63ed06342229a8effd
zbae928e3aa42a78f48d6f252eed5c68295fe8fe55568742393a042db4246e0dc7b49bd4dfba190
z24c68a0c8663286403cfd19ca4fe431889c91c82e7df0fb11c866322f2e948fa8d35d626214c92
z8264c0d2b97f8b9d45580a65c601ba0a78e69fc4c0f88dad993e466f7ef82c300e9a8a37a3f37b
z81531843004fd66b397f2b0e67baea0deebd11b0461fa7a3282fc15b8b7edc5ff86438c7c1ef61
z0067833c60f0fbe1be485f38cb27579804639270c1bf8ad5ee6c0d4773138a23f6fec92335331e
zbbb5b36bea931005c0a656c8144b48e73fb8b1c30ddab0c4d109414d492cea97c20cd00fdbe1c3
zdb43e9102c5180b5e764af80e8f585cc56c4c97d617476f3f9cd76a3a281b41e6582fd613d3c04
zadad5ff0d88c2411c00e913a683191358916fd8f9f90b7b0fdf79f24c080f77d708090351f8c07
z8c4c710dd6915808b8593bc3e38ee58989610d76d324c871b303577685ad196db7453c7a1559cf
z1a844e139d712bf49555f8208bf2eb315149d264b4eb7d879ea31925a0e4a0197649cac2336ba2
z754f9308981be0529e463abc09f038d6b932b88216325ec8f65a0c7d062eccbfcbd7a175069984
z3a42ad71e64e6827e12f290a29aa620e14f10fba73e8a0fb49b68d413174374d9a1b241d167a87
z207bca7aee842d15ef2feaa186645ac5c34ad62f26acd0fba82c9a018857a18f35463b9c1be26c
z4add74d0b3400e91f60b01a238d9528ef11ded6f40118b233f6a057b8e6bec8ca90f479c4fd24d
zc0aa40ab4bcf5bdf8028bc0a4cf09a537c21b81db60501dbeae2bedf3eae64bcea8ff3af3cffff
z525e1fea1bbca2fa8df5cb054caab77081b143d414be1c9f3498b16a0a9db8256788d7f1befd81
za55d3a74ce4cf28ce3011792c5a062c34914a9660490039b36a80a8602828f1238cf0dbd36b75b
z71c639a596f618bb45246e6aee8857f85d9316ae035d45d647a8cd2433ccae5a9bbcdcb15090b9
zd7fe458889b186168557129042f66ff2cdfa3f9c7c26cc284bec2b7af5368d981a2d61630c0303
z8805b954e2bf6593ff61d75446442d8dc2f662dcba9c6161e92d6375d10bc33c53c208c93a8ff6
zd6fd651f0347daddf8deff8b9fe688773c85a21f7c080704042e4b56b52a2f9599399f24f36983
z31bfe07d718c105ab749b55280e8902ca718153f2e9bc1bcfdc8bef908f6753554dcdc7f55f9b0
z57c64a9e5f53fe96912292b50b34ada75b411f6ca8aec87049bce4aa676d3c26ac5b9bb7932b35
zbf6d901e77dc57fa594854721887665c66162add1d54978cab43617f22a01689b9836db2cce21e
zff42ad0e9a2e1bcc2e881847254827489b5421dedecf9f8403f94a28afe71104c2d1d382ec48e2
z7d39a57c8029103b3567bc38d0ca9e2fcfff6752991c6abaf47dbea75694dd3be1ddb89950b1ad
zfbffe42a7673321ddee0f578bc19ce4fe70c0a34f87f080759223a66e169f923ef3f73dcc603ee
z82eb1108a3cafe8ae7640f2a4016d0231e9101cbe1d2a8c89cf2b3b69782371cc3af999b7fb7c4
zc870c61851114240b39e6aca0efbe36cf630e3e338285005e6285a3d2c0b93cbda6066326290af
z0deba3e9c5621873462e51222ee836047a7b8962abebe3ec9dc27e2e6f05ccf83db17ee3ceb178
zafc323e3ec131632fc82935d583f48e0702c485a056ae5f60d8ec0c2a6641fd73f9aba319ac9cc
za9302b4684a458a7a23942fa8d6ecf60aa45acb0717da453a519082a20242f2eeec70a54e94f8f
z962de68ecee47a0afa73c2f1d0e99440f7beccdd34ca6f7eb76460d0118250eeb0775475a789ea
z9b9b8dac5bf2f34b270b1f752ce644085bef05bb55f1a5c1357666e3e22d8e22aac99fa74c49c0
z4b7557c4f70e5e05630fb3fffb688f7bb9b40f75dce5a64e4ecbe82199ec82bcdd30c4cf891253
z0882da43fde8ec50679a740baa2a5484b8c9bb486fbc628b6ab2b88a6ac1558545000b40d16161
z13209661dd2ffe4caed93036260301137f541fa9b129bbc87e982779261fe998bfc90aa588baf8
z16421a1a9f50fbb9964688d8b4951837f3d7cf82f7ee0608a8a1aeb7cf391e18e57f100083f070
zfe4776dc94de5f2cf68d6cdd4f7beb5f2ee35d3f37732471ce64af34af0b6f66e99b5d2a59aefb
z498684209a32201bb483fd67fd52d3468f64bebd766d095b09d396b46fd34b583f53857741bded
z7bfab05310ef7a0bd431b23d4ab5cc7149803a686a59204c9344181c56b1dc3f44b722603bf410
z8ab4b7ff8ee83fe1e33ffe6b4ab9e4dd267113b86ad7409671ddd70230233c6991a3cd8b12b762
zd28673383d4accadae350184576c92916ef880723d7a9a856c96b78507f9ffae6098f3904b383a
z55b000321f294a9469e40014ff97f222bfafd58e188ce54da82e4f692be85e0277fde1d0916483
z9c625d170205a3f4f8f8d92bd38118b46bc906a333c87f09d96b27b6b31280e7db0b22308db270
zc89247f6db5ef2526ac3d1830870c6a4237563adf452504c7ee3359af0a3855e5a9f67376cf9a4
z9fab8d493355a01322a8e14a7d55930a7a73c5c107d9474846dfeb12e56c68b3da91af17aac96e
zfb3fb7a1adf9d49ee103ad4b20850ae74ccf4ac34e42c2ad9575fc3aa270f96a0761b668ef5ad3
zde14fcae5dec953833f67d114f8de2c403aedd4d67274978be7de5e6f3f87999f0627592ce6654
zb19012fbe978f0da02bc609be87043580c8cb3f2f81b9a32077d4e455320aa4e2cf2397af28411
z517dae0b47662c6d33d6f5ebd7cdcc21d614cedd27be99ae316c4043a2a15e412719f19488ea2b
z48dc38287506e382e0be8d4a7a6a40f409d39bc74fdb97cc64fd36b56be620b600700ad2e6f34d
z8d51c77d14fa5c354c55db2db0bf81dfd1de5c7f8d104972c443bbae4016a1a64946edae82e1cc
zef6fc32565395a3c432ce664267e2fc9b7fa860115374abef2056ff06262b3555791af0670d804
z184eadb8d31336b7c867624e40c4453ca35c7a71f7c6a15c4913cdbf80b414df14c17e27b28428
z21aa615f85073fa6d4c6b4af3b103d2deba0e998daecca62cef3c6d684c4c3a69576ecc5706ccd
zc3790ffc91234dc85f7df7b17a7bc26cabc3fda4a16123de73615ca193ffe50873033efcf6fae4
z75f5850807085a6c8c6a7c3ca66ee44001986cd9c670c5065b10f18559c63cce3ecb4b4037c50d
zbba1fe6cf34ffcf9d9d5a05b22528cbbbda7d587e5cb439ae2f1e80a16aae7a13163fff1d50e2c
z0ab07336cd1d4abccc77c6a30ba8c12ff7feefdaf7dd72bd5ec2c0185615468a58a5fe5b2b2eda
z5440cdae82bba0b740566397a9d2d4dfa9affc0264ec0a1dc04e1eb5d9526cd8bac08794327765
z65065ccba2fd92f12c153e191e9c7f9856f015eba4e50f7f7faf0a3d4c01b6781860d295f01fe2
zb488dad94ac390db335b3dfeb838495c3e181bf33dd973303a6d1f8855aa4bfe6e68863df04ff1
z75f23d5d080a183ee4e57ec1c9bcdf4cffbe838963f4f027ba2d8fcc8506f0dc449fb39c9c257d
zb5efb901f75d28b5be859770bc3ce572bc066ce97beb442d97155e655a589a054b046e7171e88c
z25a3612df72bdda0e75e82d849c9b18da28b7fa62a8829c45972780bf2e5c0a8f80dc4e9be0bbd
z02370f1910960a17b1504724f6ef1e72bd13c131dc4bdb916fea72a5cf9df6f57bb3601a2521c9
z7194f5bb63d474f3746c64ca97402a16b39d5f5e1cc3aa62d472097bc153ec5091632a2bbb2abd
zd8fbb0a645e073c6d1f0ea0e36de49b24cdfaeecfebcec764e42931333e3ddcbf39030ee706fc5
ze9a2c9b774d27481d0fd8a655b359cd84950c07cfdaa84f52d038d66473b35d68e5eca6fdba330
zbd1e2c30fbc6025bbc465522a4916c93ab9dd420aea86aa1d055f85ce4564f01b590592acece77
zbca5eb527dd80df365901243ad3266d5965e81954d3ed0caa6d151b41481b3770c3fdc4f1a37aa
ze1565a1521654086127b9b2abf7c2d7b44b70745de1d5046cf55339056ba29a9491a4b1e16073c
zada10873938b00942632c8d4947feef4957c0b066f09daeba9cd421b7c2b4c73ab5f274199528a
z08b2801be484fee4220a1d921ceb7e64fca91bf06e980c13a61768d6ef606d1a65766e7ac64822
z5a93c08ec9aa8ee38ca47bbffcdc55a0f236c7a392e4a7553d159afd4badaa90f0a35837a0152d
z504428ceda80d161440b6eba09e394325623ada0fac3d5d149165c61274080e61b57edfb978dcf
z96756350291beb4e0c7f6b38206c5c244932f33592aa4f0f1fa5701ebcf4072cac44d2b5fbdb28
z28ac784b6fa1bbbaaa4cb17e0bcb9d177a5931874152bcb6f0f7586015674b8de5ffb8f7062fbb
z1aa431ff16811e00caa7d203e282b8f612e5266e73bbd334189be95950ad9f2f7e27c7cbd170e5
z0d8be339c080af7157f7e21e76228581a666064fe0aeac6ff3fa196636fd0ef5ea2c916e345b16
z8bf18223b94d38341f28d8df8889f89138ec5a1be764367f34590475da45dd75a512886c7a09c9
zf24fdd0015d59be8b3b68c2d0956cc523dba04cbd5ad339f3cd72b16202b2ab63fe60bc9f16023
zd73e476935ee1e3164a6b011b61e6f4eec1c5c914c2594ed4aca22adf58b1fdfa2539ac8bf63e7
z734e3424b1b8c192c4336ed4cc34b65b4b1a9a9a3b900c7c9cc1493149f2c191658b8646a1b943
za823341fc979980c960cfd8dbbb0bd16b2da2b9305dec37f9e3b6aed3d09388c63767843feea62
zf29fe89e095ff4ea68d37d737bc0e80467c90100c5b97b13134f1b58afa591b214643a45855e85
zea14fa50f7b2592550995675df2049c8c621f4fdafd8db651670365a54a8a90a6632c81461ed8a
z702897ec009f4f54220ddd095a4a0e2e57eff22f7f838cd5ee18cabd519f33229ab746c0d7c966
z6cbb7b43f0bccddb260bd74f706a54fe3c7bda3409f7f353cbe6bca5159afbed117ea1f0b33d25
z20a6d1032deb1665f934c20599c065a34a33cf1cb46aaa4b2f9e8d8e973a6aac9831f77f9844f6
zbea738fdcde12515cac6e88939a58b567074e82d19ed8bf843b64dcab790bb947208ce2b953274
z12f2154596c9d90885b865738244be4a0cfaa5e579a9c2b2852904e00f2a0accc21fabf5a6d67f
z65f27013f3e0e09f409debc7d98651c000472b8df090329023f1809ca9d23604e03305f0d8e892
ze088363e25a295cb0fae9002eb037acc60db1fac690fb755bc783b378a0d61ac074ed3bea7fe67
zf3c8ab435aefba9db2721b6a78cede7bd510c627c7097db0767267aac8c7ef007e83ebccc35894
z662d74adaa47dcf935818e82c2e25e9e9d3bd4ae93fb2a6e2f317834a236856089cbb0654f6eff
za79a0ac5278cf190fb00ab86f11d0c48a07ecebf16676adac33a52e58bccf84e4d51d94eed1993
zcc2ffaff8990d431386dc002cfeaf7dc67d6100fa37e6449081d7356a3c073a81b91dd183536ab
zed87d7dab24cd9d1fb5d70c9d6e37dbe4af32a3ff9912832fcc1d1ded60b46e2b956b01e734f3c
z30c2a9902a68fa1d1f7f053e0f3ec19a7ea41d1cbed26aa9d3d48751ddcf02a4a107105ff00b8c
z2fec7f8f49f911ed3dec1c69c56984bc8cab76020c122d2e8dc65a1a1dfc147effe7d36787e70d
zb0d52318188314de2e0622c2ea908ccb8ac9960b89f5828c6b6600633baa9ce86ef362c644f0e4
z7e33887f4b6d08b9a11654a8465c0eacc2197cf0160ca1404cbd981007d7932381339a051af4a0
z4e772ff80a2cde1b956441456932be1f7ef1f74444e0cbdef8fbd75875162c090855e7070af42b
ze6e0db85956a9a230814088823dc7cf692db0465b02e9eaafc402c3a3ea47c480032a89df320bc
z61a767d753b54c75435f54b4ab968bc2f60d34e5030ca8fe6b0ba90e6fee8e734decc7b897ec97
zec3cfa5764a6f380e1fa10f3b0ef461c3a3105f1b6a420e9d9efc238a018d61203f3ca886b83e2
z11b9adb060949b3a374b80f0af42d825e63e01d3604c4a286c4ae14f4a82c5a6ad0802ad651f9e
z090c8b366ef285cf341272fccfa59c576a23e82096b5d325f6bb271c51c463cf9e18a5293374d1
z8ec7cc867dad0495ff51365b5ea47050d7bf0d9e06d9cbc6e1b56dbf6e3ed5495f0cbab2b3252d
z763bbb06c6ceb80946bf4a46176a233fa82aa34da96b2d1632f40e87804ffcaff8ca76fcda33be
z7e367b5491da6e7ef7eacdec8ac017676a5016e33ffe23c0d35f051591b049c12f03b879f1802d
z80fc4a2ac1ea82063f1f297082c0af2c8e64d3ea1f73139f12858dec6e92ea38cf50f77594ff86
zbf565324b1c419fe8d18cff15eb01cd153610add9da5e0a012f91d6732dfacc3f956f075e6a093
z6e81a94c7f4918559343aabecd8bb8e5cfa9fbf7f303a957a82936c1c6bcbb64cdc05399db4850
z81ad7d08be819a6efcf00fb57e53111f03d0326e4dc8cdb5364e5967a437019e1a6451f4bc9d96
z8fbac3f4c01b079e29dc30278c25de1e94c49eaf66899858ac7a4f5c7290d3fd7db746540d1a34
zd72931c4dcd6b36cc425f0fe808e1aa1070bbd92b95b8bdd722899a156e426c809a59f88928716
z6097792eca3d050e01aac4960f8c51ee370e593420c768657a2f8d45750521542e53ce243089a3
zcffc33d9a09bf4d03d4de7a4184e199c5874b1977ff25abea01282c3b6a51fcc78a0de6159d916
z15f4659a6d9d2142c1dfac0fb60223002c89ab03247915c41d9d9b4da80a443ef5fefd766fcf8f
zd9daf1d1119887f5ab0e3b2f50097bb14401bf62e36af764a933692abc9b4bf7148309d8be808c
z0fe83b8c0d5feccfbb37407bf45982c349ad002dd84b3126d84c876daf77b644da8267ef316a86
z7f892ab9304a185562cf7f09dc9c9721f43772985c591315887ff1b1054cf127f24f570a5ede8f
z0fcaa0f0888913dddcd038104cc063466de6bfed8447d04dfbb514847ae8cc13082b92a9e45770
z1237de5512a2712010607ac8501e3cb21aabc4110b44aeea179ba98d9f07557489cde6f679248b
za8eefb53ac0ac736d5d4c93fcdc073a312f79dbeb79f66c84e7c73c15d089d0a22eef3c3043b53
z26566c618414f8790828f7cf4b18e4501b32a4790c53bcbe4e6f82facd417e185f797677f31b3b
z9a431f49c48166d254eb96c62e34007e0e2779ae88ff3205e340f1f1c8b72c696546550265ac45
z671f32400b6a511c922935e75f4711f7dd04e3cb9f500a500fb5c67083e36fa6cbdcba2f59a742
zcfdc349cb95f9e04f1195001705a9a02514f37b73d950ccc5161027be89f8702e4f4e973a65c14
zeaf62cfe0b917b72098ff02c0755f47b7c96966cf753fd7f8fdf5547afc2681232fc91b2b88bb4
zfa7ae0fe162d6ab1f7b6684ba107e3ed0e13af00ee2d1527a8936daed16fe436866a12a64c8901
z3b90acfba473137da75d8ecc2282d95187a326dd0e84569f9ba8e142b50d39546df0d8031fd4f3
zd8d4673eee5f553398c05c795e17867fcc10e592e72bf32fa9c1bb449539ac6349067ca984acea
z0a9e83b56305b817fda34d909eff07eca1acbec7a541302f03c8b9b7816c716791b7806db59a79
zde929b1430366baebbe620ad7c47da3e93128c71bbb46e64395a92eb0a845ec3daa6ad0c76a964
z800ffe261168edbd86d9bc1886c3cd2d651318b7e381f6bdcb6c58bf57b7f355007aad5779b56c
z3ed53b9de1db5cff816dd2ddcaafbea1aad387daef35a42cb58c35f72d0f6be089a8c0e2daba86
z21fa926239c8a8f5bc5ed0f24f56998f1410a430fbb8b8d002834a5cbdcb6562e4a5e48a380356
z4828ab3082818b0cd38a7edb899ac1871491900768e1e6a9b55f5776157ecb1c8babdd48ce12fa
z84831ff11c138e3048038d5d673db619702419b8422b1a26ee9eb7a45be32f65d0adce510d5a0d
z1416a1b5eebbbec91e1f3e599462b36d6c569ebc0ddfb045139a9eb4e9d861bc93cf66e51427a7
z6d4fc3e3219527520c5393d82ecce081e0ce4b54849a74686e2df31756e8879f583ecbe87efe3a
z717861ee42b7389f46c4e018456f970a4ab71bdd2d1164dca0a6e901326b4469b4927929a55f43
z7ce1613c7dd9a9d61205c97b5da9082d6addc0b5d2c86434a06dca276caa46fc196ee6e4406c1f
z7ac18e28e6f3037683a8c00d2c81a9d8876042104046eb0a514a6284aafbecc32393bce9ae5d9e
za0a9a5068f6a5b0084935d2f03b561c9ea1a6f6fb40824157d6cbc2e607cfbe0444dfc055b6ea4
z4fc5f13b187b8ff8ec940166ca9f542f3c1600bfcdc7b20a0399864eedc418cc47a955282c847e
z1c28f87ee8ba079f2c34857f7354b14ef85ec0a902cc3987c7413b279341938b9fa1796d9d0967
z66f1e162a3ccfdd70efb0a240df92506641dc0025b6844548bde49acd03ce7b7b93a1d0bdc6b47
z63ed9bc65e2592343dcbff6bd96e279dca44ee8f96eb827556ed7a2e5c1cb76291ab75ad0a8f87
zfc8572eb208739ad4549aba22e1b5379dc7640d04542afe26f53eac8d597456b5c35c73c869281
za52565c437fac30fca90ba5397ff6cda0c3442030afe248558c66264a81f809be90960a80de794
z708f1d96532d5da031a39770890b1ca292d81492cf74b7e2d4e0b96b098e41adf5e1e02666d932
z7e642e9e307bf38d09e7486d9ecab9d1c345f970299d5d7165da54b44f0001ab59e719fe1eca3e
zb9e8e56461ed8ef2ba63bc7c1b80933228462cd02941daa0eadf61c003da90f84a0b69fb1dcd73
z6e79a414e94d7f8b261b481d27d75d746294147f157756829b31a3835370e8472e181b67e46b42
z433e0d6a6260cd49fd1252244f94c7987ff109af2fbc991d3f20ed9481c35b1f0d5f0f5e3a667e
z1b6b418ee98ba0b060bc79ad2eac3bd8834cd76c5a42ffa7496f2f29e36729e0522b365d61683a
z1f0bdf1d211f23fb8c27f77f1fbc1e354bc430702abf66976d6ea183c52c94174c0099a59447cd
z94cc8b9acdfba1f08c7fcf286a7a9e44764ad1902b487e800479e77bf3066bae6c6bf81b268da2
zbda5fd6e9ad00c10bb532ed6d3564fed1d1d36d36fcfcda72aabc16d4abdbebd87db48b695fbc2
z2d54488bdf5d81889d8ee5dbd063da61a58487a7b678f8af0b0629b39cb0d74d6af4483e3e4c75
z5ead3e1b3fd71b34d8fd07e1f74d36f488b63725c6574db2adcf4052921f42a1b2291e347f84b9
z3560458d1b8e704602d83bef7b720fca2675a9ca008ff5e96226690eef3bf206018c89c24de800
zec42ecf1b36fe318041a82b6cd2beeca2afe46f0c4085bc9101851dcd789a5809a8224c1c7c657
z7075bc943641d000338d9ea40981dc0f75d81eaa844f31587ed8982f071504b6f84d04d484374e
z8e7cc1d9a55b46d0cde9faf4c14dbd2af49a1870751e0e56567d35f7d24f98971c22b7d700f714
zf638bba5e69ade41fbf1a271ff770840fb46d9a2c9535444f3fa134ea8192904a86a726132c490
zd5aa3194bf2ac15bc90d46a89f6b733d4103e6b25c0e380c8881afdb5a813808608413c4136a0d
zb58ec20a074900cded028705d7f55e020b270bfe5813012215742402e6ba548699017faccf4808
z8103595ce0355861b432d34067a84875f12609f97ee59345ca5c11a73a11cfb47986c5d4b601f1
z64a216c3a0cf5606fd32c1d4c1b9f1aefaa64bbef3ad531fb16f6cb9fec94159e317f344d2b298
z03e5dd225021dac8cb07a1d24980c6295a92ba09b4162c26f539ea55196fc15c42e11ca7734f27
z17e2aa1708cd37baf38de726f2e1e3fc7641e76942432c7b087ecaa0dc97afeac51aaa09c53b49
zf7070e8ca4617b64493815ffbbd55fff7e58b9a25f8e48580a289aafc06796e29a8ac08ac4de5b
zb397942c8674847099411bb5843926a6286fea32d5e2eb207e7a198403bbc790ddb2c4927cd3fe
zdb4fc928eeb2a2ebb71b17886980b9d956d42aa8f042c574e7a522a7fd36bb62e6913028858ef3
zabb80a48918d246b7207e0f40c146276a3ee1d66875324227c40047bc70f48dc9fee37cb005725
z981b5202ffc5569d141b785d2995a4153a3522427388e6db3d9310e9bd084b8b1b972b23deb9ee
z5d8136168f66d39b01cf8b9fcc842e3ae491c8c33a6c6964bfba5f2c3baee233a90235caba0dc2
zbdb9b81bad6061d7fd5f00328835f9ebd7388a4ede5fdd39df6e3a618e29aff843d31d3cf39fe8
zbb21cc98c258806c804ce5604ce1448fdc1b16147a5c9cb8dc2dee5a65080afc8a0b8b38d0ebd7
zb964e616c92ba55402942c17b3c72c6f93800794ba41f30895148a3e25edb786c0fd9a2775bb59
z8cc8a754d7ac88c7ad375630e917529687df4b0e4e1c07c6337a600559cb2f25a30c7f26017508
z545a0bb0e35057fd7c08543c058cd7d0500b3aaa5bdc428971055923f0cfa352a971926a80f724
zd6aa0da7e8ced599a22bd0c5c7a8dbdb3a08602a0393e417a34647f08d5ca9848c254d2ef5434f
zda1e5d021b517ff6c38b142b22f3ec2624e0bd2338ba3296a663b5d8df24d96f0ef5af35bd01ec
z90dbfd01563aad1b917edeb5f27b9a26e5c825c5991c01923a806c05a54ecf98a11136d4f29e4a
zd16f185866d028683949325395b8bbf3c42670ed59775f57107302a1c9509586b5e5366b6344f9
z00a8020bbfd100e9e542e97c5c0a69ba850c1c998adab414d75de2cf732cd3554461d5c3caca31
z19755377da8b07f30e7896ac5ba55561d1853eb27deb54ae7ed31841a1dd724610439dfe2fe931
z996f46ad34be048cbae09325ebfea02c2eadb7690d306bbcaf47b230ffee20102efae8c922da8c
zf2da7ec2efc349bd509ef9a5eae452249fee4adda6f186a14411f80d4bcd5bf92f35036e1b8e06
z0421c4fda135aa4660ba401bbce2c48b31adef5eff7af3df3298fced961b07f21b4b7f0121e766
zde7905b1f6814e458eaba08a5c99064cdc03fc800dde8473b24dd5cf503b81a2f2dfbb3ef159fc
z806a1a838066e238a1b3e958b93119fa5f0cfeae64b03b8d933c9cc24f41a9ae6f554cc8d51042
z7e38acd2c492dfade8fe1013ff8af127c0d8e5a6c5ab25182c05d16d92c6fefec7c1116693be2a
zb4b705bbda507216265dcd4681a6c333a70cc3bd7bc4b00bb9c4d8e019c034ebe409ce3b218c71
zf94412994362b2b4f716d585b232644cc1f7b3a2955eaf03de7c5b918a8fba1f52b6196b234ab7
zb1052253f86c526a3432cb9196eeaa777fda71b7b9b6f6331a7ee436dfdf035d7a1344fc4bcce7
z4ac8d86876abe8b2aff8cfb4c88f4c2f620aa3b2d98ce32a07b9a7f529b556a30a219a3d4bd230
zda2fe8fa0cf9ac9d0c838c3517db1c0927a20a31d6bc60f481a31610bd6b5f0285a01f9f2b3c9d
zbdf3dd35587013f95aeb6c74d0eed7aec6a3150af4f5d1f3d8da8317d4e351116ce9223865485e
zf795e9b123591aabf333e89720bb89a37ed9ce3ef515d11adca4a906d0d5fa7fa86f2daa79b7c7
zd5be7e8d2062ac1099f38eef335abd027854e0df603602ed31108a2d08cf5b7169b1faebaefbfb
zc11dac912dfc6ae5bc1bd60b2378fadc0cfe1a1bd93e14799408388dabaa43a63eb3412810e66b
zf931db5ac4c9847bfa6ecc8610499be5191639439d2509e3ef452b768d7b0377f747a7857f7278
zcbfc8b7db2be3461807ccdf5b772dfa6c4972e4476f186d6a6cc56f6e5f744d4bbf5acb03affb5
ze9700e25896b7552cc65bd37c490f009f71636dfbaa7c7b2c4ebf413c37174359e038daff3d1f6
z8b415fa2875aea2f1d4dbd27e469ebacc5acd5a7e9d1aeb531fb03ed0169943fbe189522c22a23
za831219b29e33008828571965330d83c46efacb0b28d743b640ca93ee91d2bef1936b38c7f0abc
zb1436a7d65c032704007501d8e506234981fa03dbb9cfe8c761f356a0e2b194fcc4dee37046dd5
z965c2d01c112072a42b0a6c99e685c80297353e50a580c9c9c54b1cf38cae0d10b4987f4bbe0fd
z1c10bd6333309c599445d41632e534bf91c67c64d79544bd42cd93c748d570ead9f29205c9cdee
z6e031f6306dcf441e098d22dca661ae1d3442a51b85f7a0aee6ce077c7c625a2a418d9863dd1c8
z10d78273a08a0635123a9a26606ed990be0ade6a4b9337f13ac7db43b11b329701a21d1f3e499f
z50cc2982f3498e7548e8923da0150df883584feff7d4e2d9d2b8f2139848b7d7ea9f94c494b7b1
z53803b6e09a8bffdefc62a50d475306d5dc0ab05f89bcfd2c1af9e7c421b1295ebbf036b41eec6
z591bf0acb68019ad686adc49728e56fa8153f5c40fb2b58c6452fc624bc8e2dc28bb4cabc3db5c
z8454bc83105042328bfb6bc26c4044c802705670c8cb365c5e68f4da23ce3463b971adbbd2fb48
z16b08d263992c925fca1ce02757bb9a2797dc1159b4780ff696165c4dcd297081d63a6ad38e612
z89a949e1b22d04805b2debe48863207b1766800e824209d30925c724ab3b795718972bb56f7dd4
z7968581fe02d8e31f7199df97ef4c4cf04d5088d7a4d4f44bf6ae37836238a381095176512b30d
ze83a6908ceea98c24a53255140df559b9f4d23fe8ec344d1016e65d2e00c8739640fede1028b72
z596ae6d61291c00ad54026b141587733817806674e97a56f16667c701ada67534f1f1163a59484
ze6ab23a3d63c6d47297e833cae3e5c5c9dbbc19f90b3c871a02359f915ca637d2b28192c813359
z811d17029dcf2218c9f7d3d6327738547b733600d4a82d136c7aae2614555e5a0e60a5751c9c40
z439f6f0e299c7c87ea91aee4b5d63b23ab0fb872e12af50aaf8c2e636b0668bb96abf387aad520
z90848fc801654d6c1bc5380876145b64c2c5e46708e6e7a993c149bf51e2f8f937221dc1683bd3
z460506c5a1f809ba48cebfccc2a3e78311e8357c839101bdabe6cf6369eb873281bdfbdd0c270f
za88334efd42b94a3c355a77e9870cb75cbee74b0ea8d3ec1adde637fc104ec0a9a541f908234cc
z60fef7d53c630c200c3ec9c80d1165e97762f331c46f930104c701a718e5e11703c4d4896904b5
z7919b15529947cecacfa1e5c6f7b0cd630459d0a4068ec1c2e66b768bce3402fa3e61624bb0a1e
z1792528d434a427c4edeee798fc97b1d93f353d2e18ec01a62bfb22326db3d2c90af0ef9f5a823
z5d1d1509689edc288cd0453f0125e7398960466b38feb68a4eaea861088c3428108c8568535086
z874c70993de2d95af7a745c516965ffee214b53724861f196b9184f535e102b58902fdd9a2b7b6
z66d23298829b8d342b975f0af31fdc6c409917f9916e7eb53f51d454e09a7ced5e1b57bbd0fbe7
z93566c831220bdcab43eedfe7f1fc6ec4990c743f67d889fe26ba40afa59372b6a8cee64799e2a
z8597ace5406cc9c5ee180be901bc9a1ad3e223b6de795860a16ac38a8b826e24e1f108313991c6
zea0a1a43fa6a3b776a316c58ab426a34a1ae76b69966cb0d33d625f450d031089fae4908d140f5
ze2f8bdfb3c78d2121f86eaf0227bcbfa1702060aaf1990bf17792f036f0cb95e75715105836059
z95a7f5037226535375fd3c94c14a71df9f1d31958dc0d85520f4d9bb636fb711a55e6a09cf2853
z3d1e6a1d4f431663030f1b9a219d4cd7bfff6b035c83ac0f5eb28ef10779ed4c45974e437d9578
zb4c4788bf1bb60849b80350edc5e52aa3aa3f7a423f9ec08f7eb1bca99040420cfd50d95d608e2
z00dd099fb1ba5e64f940102ab8954b859bd50083a257c145a77a32302724a29af32b8490412218
ze80d816dde05a120d1944c2ef55768d9110df71a27ee9ca9d3f99acec7902a6da89ec13f734ee9
z64cf91c4d02c20167b6252d22142516d0ebc1ceaffaefc593370d5c317230094192eb8b71c5ea3
zb0e801c3e6559d2531592b93024c1012eb83d8185cad78e8ea499e4d4ccffbd860e944bb507a47
z035c406b08b595cd905715ab26a539408b47f29729b3b838ea341222c6babf1842417fc1725265
za49a435e7a08da04d453f8763d8200ab8a893934c0c8b5a9a2b32b8c91a12f76806e4a14f8903e
z753cc19e03453ba1cf658d5854a04c995c6adb504b8ce3195b261c0d32615d5905c5fd4b4ae7ad
z89750573d588447373de6c4a39eff52c4bfa73f821edd9faf91334fdc421598bb819cd07bc71c1
zaecd478af590e7df0c3ee8ba79435189db44ebb077d1a55a797fc2693c22cc2f1bb593c8635216
zd0e3243629e3e44685f81387e9fded3eb8558500972800f3bdf5a64fb33617954eae4fba1b1e75
z4989f8b5c5ed933629e4dd0e67f9c90a21cf4bf1a16e92da4a08cad3138952d402aefa08ef9654
z47269430132c639e4f8dd6c53e554f8e43ba39fa6c3a868cb1e4763a5dffa2f225b18d2cdd4a1e
zf5562de3279f09695ded15e0924dcf577a035a16cabf2dfa115e948afd7266996baedf9085f9a4
z80aa2aa9be691ab3d75e6e1f9796d41dbe5c4a69c45d0d141320ab67d55ec8ee6c9ee9e6b3459f
z5e09e6f65006cdadd9d6816f5bbe8267ebc1abcf94381a753b12f96b30a70079c19c64440ac124
z3c4a9816865d8f0aff25b3bff8da8d2471863abe684c3a4841ced3f2fa367003043dde45b3200f
z5055a5c535fafc34f2a253864d41b7dea50c0c077f936e293a63648ec2f413ebdf2c3b89f66ff6
z9518b1cbab3d04117ba20868ba580cdcc800c6fe71ea23581ddfe90157faf488d55e74425b5e98
z0e32385b5ee8a8a96ffc8c45c7e4416524bd64ea371bce9e4e6edb3b575950398b23d176a994c5
ze9c805fdff10f832da53ceccc3e5cabff6bc887f7ecd7502d5a7aa33815b0ebccef62a0dce6cfa
zeae17d75768f825e34c5a17f276af624a7966df125a8648e1dfa2a1aa357fad707382af2cb03da
z0c8bc8298e5bb90c871c9ddd966ca541e3298855a3345ee631f3d3ab089d4ec14e0ffa6675ed39
z6da5babbcce0783e869c3496dd32a1ea844c12d4c50a0847e492b82abe58334b63bd93b7af61cb
z134ffb7b87b7bae2d9b0531bc88a8ad4aba833cc2c1cdc543b2e7ef1ae7803ebb7393c05d4927b
zc2d82d3acc8759b1ca3760ad6d328a35ffd7742bd33c10b8757a291c5eff4a06a3127e0761c998
zb323fb3a2712b6ed0b24f80751d4b6d44689f92f8123a475b87ccfcf0d868e3e9c7fe6b2d0361a
z65f77fd48d21fc43a7999cec1323335940928f2ea683941f4b830b8fdd51f9f205bbcd04bd3d1c
z00bf5585f8eed0d4531a41503a427f9a0b767970cf427e36e1909e3fc539e93a0ca43e6b497857
z6d89090a5aa8fd57304659d374fe3a6dc656452244c5c8bea6ec071b8fdd321aea0ac961375f79
z27838adaf914e40e173c0e2a4815a1a8e6709d4ca12ce6af4b4ff436eecd067794d423e1793f42
z9296cd41cc50123b1eda2e1c67c559419b57018cff21202dc9fa1b748861cd7c9b51462ef97a84
z1748bed791527f85a37dddbc7e9ac08b926bad2442fcc9e010ade0e3d7d47ea70411dfabf8cf73
z2d4c7dd30cd3aa93efb428f709770aba4f2ef962022cc611bc6d7043c5b8bb2e08e337819f68a3
z4b5489ac282632aa3463273b51d3449a44683666fa1c036b80bedaff53ce912652f7c23c066744
zff177d9f4047834a083fc2dbcb1a0d6e93804cb1c41bdc9bc6f28ba9aa41c35cc45dc18316866c
zb58ec24a582e6163bb07b30213f02420d59e6a02a6572ae9b90f108bb3cae957abeb990ce530ff
z1db51dfcb6f46a5b797bbf59d71f847bc04b76381c21cc7827403785778134857d8f0108a863f2
zf7bc2bde702ef89feb1066743e4d6f753996ccccbc6c6966302be9b60907b8b2d911bfa86b4e36
zb5723d72beda07e23b3b0ac4a83e21766dabffb80ce5615c7961738f4f3b7ae83d66b6fdc0ddd7
z646881589a8f2d5a3c3acd0962927cfbbcfe4402376f45e6435aa16700b7b196286c5a7a4b09e5
z59ce1d8ed547da21bc60aa566f6bd6253683ae46165cedfbd1ad9627dfe39f66f6209ccd726c30
z0bc7985e3d95e815566f96e686df1ef42d3f5fbb7d8559c7dd9740c070aee749e08fab2e0858e9
z774204aa4a7a017f6693a0053662cf7b539183d5d05a40400ca41f0210a5784fc2958fbb10fe5d
z481f238581a9b564138945169bd76882ba3d3d4da7d901ec3cab7bb37ca01f9319a3ad99ffdcf1
z8b9e4a21f2a2fe90c2a31ef0344b339f83f1a9ce534d421f5f39c506c913223e39ef6aafe3efa5
z9559f7e9c4d5201c92fb54ab686218b75bb8f87f48f7ded0a0fb63111ad2a2bc644ee990053f3f
zaa7e8c41ecb896645907e846764e261cb12d061b90cf83a06425ce915b5ba5a3412548116a453d
zadd4805ebac2535b1adad5d030cf800e3e12723e06319d03c4667b23a902487183d220a7be3d56
z2f98c2d342b35af29980d11e82815b0678866fbb9237538d3a8c3a736958bc82a27f65d56db0c5
zc4c1d760e14bd2b829ea2dcfafe7e67c036874c0b5f439ba68dfcb149ecd7589ea3d737a34fcfa
zaf984e6085922f30ffdf9f4f4f218dc2df30861cded373d406b801665af2b56b5cf62444e74549
zc2766722951dd4e1fc57db8aad2cbcdb0def6c1c9654bdfd126c85fe7a6106d0850c320161a823
z101cc109fee73ce1f0a83d958bf19970b451e8ac74861ca8820c420ebe78d88073989660b836da
z1556ba9124cdeeccfc73542d0ae9684af1a43a572b2d54230d7f47bb1714a55f9176064bb593a4
zaa58fcb7044ddf477244d37194907b68d645028df3ef3bc39415f8771cc4538b55764f5b8a75cd
z13e6ad67a2cff411f4b6964c64b9adc400a63e08796e48987ab402008455d0fe56a33189aefe1e
zca866d5612e5e6fd6a889df43424a16bc2a0a9541e372b9e06727403e6c668a0389cee98ceb1c9
z73ff42330b7281c4576512a208c56b41caca3c82183907d69ee2cb6e4fd665631e097a5b71485f
z02559167ef56fa1efe34ef6c6d4cb4c310fb822475db2138d00acf046846ef8c584b431dcc94c4
za9b82e8d1e8b2d5c8970e376bc7fb18a2c341f5c397a8ad719320a4814de1d8f20b2b57960d2c6
z21b060d3ad7fe6d2f20c87e72c4f2eea39646f046383de4404a33a1095d9f27f58a43072764891
z68c7df3c658078cbd902119741e204aae44494cde111504bb499312fa0f81e7310e8822fab85b2
zba92fdd213b898a592212a4a593fb488502d47a2ab5ae4fe75e3953ec5a1c5f00739e6628dfe95
z04b14d8fc40924243d61467903124e0a19fc64c5c4f77faf00a6c3f2a1ea6e5e7e3077978de4b3
zd189f822bbd093848145c5a4af3efc7bffb669f84933681fea2616926fce27d9e2ad2b162e159b
zb482e72db2e2453b2bd7cc1bd0e06eea049c76e7ce010d01349ef3ec0e2d1cf0a761b8e11a7c4c
z8416247b2c51cfb3863030678a2d75f5ab21334c106e2a53c4c119f6b7eaab85b5087041bff665
z0612646f4597e7dce23a97468d072369ed3402577b1cac379fa8eb5d5a4bd62fe17e2edaf20773
z0498a2ad69c3e6de810ad6e24d797f6198be965ac34cf2415334a6a0f632fd295447d79d848566
z53170fc4f2562a714e73d6590cd704d4d71b09c6e80ad285d2199e2204666dd7576bd0438bbf42
zbb6eb56466b9f79d35851017c422c91ea945b22eff235ee917b1726db068c398e9a518223356fd
z80e7bdbbac96e224fd0d76a5eb5980da4012cc5121fe691c08a968ba69231d41ee41ba19c9fcf6
z517c064887030752d36ec4fb39e6e1157516b3b81c9fb0f6f001754e60059528ecff23f23ace20
z5ce2a289e2e6dbee89f9d78346bc3b84ac0530f09ecf1e218468a2a0549e0da9cc04b1a12115d2
z60b5fcf497ab65959b401d6b3c6a21e327325f12e0421c003fe05adaca83ff4bcbb2664b3609b6
z0fcf9f082a12c244740a9696ce9274ce8a03c7ae1c65dbf221d7403af6236ce91fc2c117d1eef4
z971ea51b10e068405624abd24da1bdfea3c67a77649135a61eb3658f1b23b22092ab542ecae103
z37b582a0b2cfc3f7b0d51cb8414b4a6aa3c578b8fd5fe9fa56019d27b223cd518adc78e666c085
z8ea65200370da877244ed9ff724b4988f49c21e64ad8be1b3fb04aab0f906a81b6566085a07af9
z31c1db6f2f4f9844541a18fdfd2bf6ba2e626414a14f5c5dac891916411a25deb68275a3d2f840
z87ecba8f7892bd0ccc9b45a291234ab51c4bf1f27815fd61697bd3fe300b9ef1009b0ecc65386b
z7df0aa8157d1c38bae7977ad6ad82b0736c4ec1e988d95f95bbe00482761269a23b623d2fb5119
z0c12202656471aaac3889390995685eb61fd8a5807aaa9ead08fa4198f7faaebf27cfb3c10f50c
z39ced6c28020cc2489fa8d5251568b92739568b18d46950850b9fcd4c8a9922e28bc27986f5990
z0008b987402c19534d7f4df94199ad40bd333924570f73afa203366644fee155334c171461bdbc
z8377519d779a8b1998f3cbb093ef44fdee17419bdd489d7ecb040dd571553786d7671fa92da308
z345908728de1962ea2d2b93039325b8e9d17c12b968b77c04ac1e83cf6b765b2d64f9b519065dd
z0695e64682d9b6b5a2719ba53313219ad0d92315c236b725694b68b8720af5f15ec681ea6af954
z414b46f8103fe1f1c738c08cf13a6a89b6827601093ebb25d205bfe27e5a2905f0d61495d88662
z9929ff67081e8b465cb63481b38205e2806ee6472df54dda2fe678f3f7e3668d82df9c0f9f8cd9
z514741e0e49ecdb6c8e98805e97903db92e95f7f3993212990798b31ad141f4d7bfb15222d1763
z5044df9a54110b24a29a158ce355ff2b23301fb3007138a88164a623500958be8644d6c854bdba
z0bec1db3eea8eb4be7da515f44412749a698b868e5cb83c381e8e73b648c223feb84bf3e0a97df
z9bf40677d5c53ffbf68425843e26983d9f241e7dd9a72fa7daa89f00f9a68e3587adaf5543dcd7
z668a8444b7bc23e89b245fd5065e38285aef64d35c2bf856222fe22b868cfc491aa0b9cd75c7a6
z134bbed309b2da3e410ee6586be6a8a28d559755c4923f66ff6b2de779e95f474a315076b7f410
zbe6caffc4693ffaebfe453541ac49acaf8e9a3e771b29176157194e904cbbf2cc60f30dbfb929e
z268bc2a29db6848f4c85205a81cced6fdb2c2d2af86c0261b8a3e0661f076841d7b3bb781e955e
z0c8db7e4fdbc729fab75049a6a876596168eda2eb44a568c54b8ca95fcf28aa6fddbdde1101dff
z9002519696d85f3d3ec2c8800d1ff87129cb234dea9cbc314242475de3914c8f7a051b8acfb80a
zc213b42dd1263c7cbbb33f32706b31d9a80b7fd5ed018401f408caf7a3f92638a304788eb0178e
z3a20fd7c23a8570e9702f671bc3dc50a3e6bee2441ab2ee880013166ee9854ca89775a4d085511
z8c77fe95bdc7012077a1f1d202ba2990d4a50cca8869a379d16f9cc6a222987f3f8109c3c83d47
zff8ff600e307a9372aa5b70001441b094a3830906611b15d5c6ba8c5683ea71ae1bcfdcd560c8a
z71aae4c12580b5bedfe5365439cb37a20c152658a0e5a73ba281b63aaa7f60719361c164840583
z51d50fddb99cb1dbb34d7d895d76241b4fdb46dec15608f1729e8466cdd5e47dc3348376948664
z916f1b56faf6e55e4f60395484647660c3b3bba035f15a11162eb3b99e9099a7de252c2f6b4993
zb26f02ccf72e2fb9d395b78557a3ab97f7b361a17892d94d1b534cf7cda623bf08a150e3dce5cb
z52b8173a2f35847a6fcfe52ae1b1db4f35b752d2bab0992fa302cbca473143b8ba753faba3b6b2
zfcb8d7d4fefbbc9ed76dd00ceea2d94fe3bae1f9afc1a132a0541e73af3ef83566f6e49056954f
z03e240e9b69f0527d4e087eb3688d5db92775de3f4292a8adc1efe9b4f635f7c416d4f8aa9bd3b
zb58786407c31a0b76a9554594e151ca2c34b3d7c416d7e748e1c3135577e01433cdf71b646a82e
zca9b934732f9f15504f9bc140cfbb2595d5de4fe7295c6f72155baaa7e8660fe3a0a8ee6112c15
z65f5992bf4995bf49d4ec92087105625fc3df53b526fe7a2f351f44c16f0a3aee60b294a32604a
zfe101176c912a577a82c77b3629b0f0ce7dd95e7ce482420b65b2470b307e56b44e0ac5888c7ad
z77d2d5bf8940862eb995d066c591825bd87993681fd4a1845c27aaffe6e03446316b0bbb987a4b
z682bfd38600a164c51b1857f78b7a4956196bbea6a7515ac2390cd37f67fb8373b1c10659d52ec
zbd4df73a2bd8fa9416c57a2fdb31134c9b7be32983f19624bafb1599ae0b7008847de1fbb09bd4
z70a0a88e763a0f086b7fd132a31428fea5ef4911d886adfd94ea8650cf08ea07117f3a4b872b0f
ze149d2d8294e0ffed975e0b3a2a1e61dc5f67cabdc8318db83479b89ac7616225bf3491bec735c
z3744bcd087dacf8afadfe2a332cd684d714dbca1c9f87f7601f10857da7d49f90c4e978e63be66
zcda2ca3a074fbfc498d497e6f94cd2ac2cf90743a9a42f118500effef5f9de6f48a37eaba81807
zc6b7759e91aa4fd3c7945d1f98683f9d5df37f6d2f21a49fc07ab7c7553d20ab685b574c5a0b96
z652b92d9cb8535e3f2cb92e2560f45fd365e48de060f1227194fa424d8262afe84c0daa57cdad4
z73f6dbf58f30d893bdec458a3830a8ee3a333793536fe352b93a189f600fb1ade5f8aeeb8dd6a2
za90c11d8324fb5414ec66c34683e6a60f6b7fc46e87874e173a26badcc51c7d65acec3b556a1bf
ze9f0d0dbc2142d38cecf7046f3576c33e869559abd29924b238c1634560440ccdb27110e3acadf
z98cfb3ff87a8a0be0fad9defe13f6bc9b9b7fcf7f6e7f1083365bb73f0feafb3e62b1079ee782e
z75e0410317d9ffe9b69290f0d60f694a6140bd506f013490d2d8cbf8feba4c2df84d2b07dbdd50
zae87df6e6aeb3ec51ebd86ba2e183565a566cb1bcf4a17dce23faf0532db708bb5a3ca14188634
z6b2dc02a819ddf656cf50b9aa1eea41b6ad27426522782b2e8f4488c15757cd9697cbd0756dadf
zb961cdbd7917a29cdf882b94334c0a79c6a9aa1219add6b29c752154be0f6d15e2513b6ec28ab4
zd46b481ca0f5ba1cf98f8f06aa7adf8a0ffa2b500f6baf2296b71f7c093c193b8cd144519fdd6f
zb626cd2761322715fa954ff1d3fa8a80188fa4f9e261412eaf28cf070e79e617ddd248f4a70cdc
z7e6b4707cf1eed4033281edd56a7032754f5268bee89dd989e063312dec44ef210dcc688d121ca
zfe4dca7c4ebabd757a76135a9b51d3b2567fc38f68f5b147c43d998e79194d8896ec893d299a87
zb225a1e5f704de41ca43e06d2095453da749f3c4a10723c0b17f889b3398d5632c3777a06095d6
z44cfcf6b3c70e7849c12cba5b5aa6139b5ed49c2b1f42b2be080c07055d80b799cc976acef0da1
z80e5f587dbc517fb81f93e6a19604bad253a5f6e2a025e1c166d1f3914e0e68c55269388864dd9
z6a12a1bce359d3b408028ce103b27a56e13452cceb90862f85c57903d81668a891789a6ede3148
zc01f21954883ce006d2977fe1c9edd6d82feeea8303df8475eed38cd15151f0a51d56eb883b308
z10760e5844cb575544342ee404555717f62b177abae05d9ca537f7ffb7bdd8de402d3474b08977
zc17be3d1ae8355b9b0fc1a19b1e1b890dcc7d08c9424b15936664eecb5e7c4474fc97080148a3e
z61686a9b9807eb5a717710f575ac944d8ed12894701fa0c65df39e80d6a950cbb1fe97418e74c4
z21011d78189c1e178ae583d929cd2a037a759023299fa412af5a23893527a44b72145d91a25275
zde7c39191472e2f9292f91e16e009c2a104016032c34a770476ca5bf65a86d4baad00cfe77ae7a
z3261c4df134dac62683e2eed5616fc2bd321264a9c03c65ec3227684f0909655e8c8f317be82c5
zdf016dbbb6cd109590526411108917f8b4d49d74dec74ff44d0cc139745121c51ee2a4ee746248
z7dc5b1a2e76620ee41b9ceed34070e0c1256aa076e212921f567498508603edbfd9d63f7fb888e
z8a58a59e85abfd8ec708ddace8b112f4783b17dd242a653e261a20e1b99a60e3f9113f26a7c2b7
z2e33aba2c3056578c0e33a21899c1e1e155e3b57703437d77a5750eaef8b36928935654fd33a87
z10d1a395be724fc81b0b9e605a3ac75ffd80d830f31a6285b9182234ee2c1a2a79706808cbaf23
z05f7c6dddf59e4ad856896396ce93c7f3c49f4f74a8778914717fc40be39116b5f83e641fd89f9
z57ac526f6e759afbaa27a08a06098a0c3032b736d7cfc4370960bad33a33c090089cf36307abcf
z9700ded4c7466d419353bb7bfd935afe742395e3373aad7bc40bc099efd7ec5d98b38ff56d80ec
z57fb37150b3d2f930966102e95eabebff1321e4f84a9d974ee5d3fc91ca3d130dd1a1cc4bdbff8
z53fb671247d590388f54974c9fc05d85d81e9dfe6264e8fee2b407d60649e9304cf5e35992f4b6
z1e7a472728ae202c4ebc0e3ac2302b067d137f25a92850c1d03dc4d3a4bd23677bbcab12c51d9a
z0dddf42a9d802f8c5ce6ec1757824fea6a18c03e70a805ed08019dc906715a9cb501c146a196fb
z17f5acf89a9267232a47056f01fa08385d79376b8cb28d82aa31b70143422419ce4b3ba90b54c1
zdda09dd9e1632db3a885a85d1dbe1bbb6954928fa37657286c5108d99a1fa624ab1a2f30cbb99b
zf3e4f57f3b96b1ca8a9b4f8b15a633acb90ebe6b4919ac0b566108816d9e18c30c870a25d34fbb
zcc9172bd346369fd779f5e49b9a4590aa31f9cf38efa99bef765692534c5272f7adef0b6db4e22
zb31d9d7bd159ef33ef4cd3dc16c0cd1feacf602f95a60081906373a7758763eaa421630a454b8d
z85fcf17db56c4d43d817ecc8ecb1c5d9597d5015c96b950215ebefab7d8a0b7d78a8d763eb758f
z86d058d59d1e0eef22e53a47b6f0e38f291aede1e21dd0aad2c240d33e853f32780fa83094d4de
z84e8c4e0dc5ddc6e097c5965d1e22f7ade2c486a094d8dfaadb4b990d388485ac27b0a1f0093ed
zf4b34cc1709a536255f6f50618fc760ce32f0c33f6d3bad251e93fdc3f57e1fddef0ad6967a634
zf4ca7a1e3a011393654fdca51b69ff4c74ad2863aa6cc25bfc7db1ac721fbe5e1f9d7c86377ef2
zb8de41ee0243684ea06a70aa426aa8466b4be23bc491236eaf51e1a038a61b35a35adcbe719d1f
z80881d31ae7997a705a255d674bf67b84f32cd9d65baacd85255992b28c27234629e1041f49121
z6e03364952b7f769bfaca19de87a43c334e0a6731f30520ce603a5428def605317289a8e357297
z636c499d0da08c165f5a87724f24babb4bf1763b4fd2af062d6e13b459b3bd04a2c38d6d18afa5
zc536427f1d7524278925e16e078977ced04cf8862bcedfbca1ee1a35841babed0a2078ddf30b4d
z8f00ebaad5e60b371f0ac90131c87d1749e06b00b204510aaecdf7080908ca59ecfa9682e59853
z2d8a86938cec8761818b9a1b0e4f6f3ae65c3d763c5d046924b725d9b1404072f931873f5423a3
z019f224db2eca8018267f465d5142856e68fc0e9d5586fe6f5ef746b5c1c40afbcb23149fa5fba
z5222332bd66a8cef1900ad5c2428fbc521d58de6f3dae97957dc26f840edba848e0c9e3f022587
z227ac5f62530de63d008dc9e5eaaed47e2705d9acbb5d32ace3c6b4d7d2651724f3fe00db2f23e
z6d7a96d502090c8d7b1e12db34a24b8a084fef95cee37098f10d52b1747dc93a9f6a41e4a03423
z44d9f0fa2cea0bdbc0020a807fdbfaaf729f35d5603022a940a85070c1fce8b679c4f1868ee736
z2a70155a8a261b04301509c49d4d1517f193608ac4c3c2a41f38638057c918aa0f035671cfc75a
z4fd7e05f3da1e05e88a4513ffbc54d12a4ebd5fd6a5b1a373696314a8b237fbf67068cfc48ff12
z5726a267bb82fee2b46e849203bb4394b8f097a5790fe9d0eb4ee858cfcd3b22765b690dcc29e2
zfd01cf5839b056af488432b534db77bd34072407e04b71544c02fb440bb326d8fba4f7ea5cf6db
zd884fc342290ee5c5fa0c6b560daa293b24528fe2a0620fe74d4648cd1d3b069adb41dd42f286c
z84d580e30fce2b914202c164f7e558c36d36122ff976805ef43238078f0e7abdfe75c64b593ba6
z3fbfd1f04b23a9b1bc98fafe8f287080a68f12ae10fe6dc7e53ecc966aab670915338a4933650c
z3d51dab9e61407482b2a9198e77beb2d5f845636b9e04f7c527b7f050f1d12e26347957a972ebb
z339206b8b576b461da32ee12a466b232417333680796ecefad43599d94b8bd6265c4f2defc49bd
z3a6b65059d18b31438d26fc2eae926b568c677e6ebb942145604b5934dc91745b8ec45a67a684d
z4114b0570c65eb4c4b70fa3eec7986120f69bb4998ead001814da39855e04cfacb8bebb4e3de26
zbdc0aeb553d974e430748f1fd59ee772e432f2b51db5ffda88ad0baf3e0d79994ed484f8742749
z736b282efa916de1d3a6a2cabaf968b10cef2c761baf20c04f2faa3ccabbf6592da924ef52f8d9
zf7c8e47550b5e7c236a03b1fac0da62c8873b8a78d85eef3424d1f6443ba6ce7aa8e62697b7a6b
z79e84ae6098b0b30963daed74c5a90feb5fc8e2d0f37dc57da4fd98f82ec1b20d3c1823f985b99
z4098237dbd0712076d60d077f8d5847fa15361813f829992127c4d65490fa299cc889ffe641b56
zd051363d9d4b49ce9c0be4ccd184866b1a7d53aeb344b922e9e3638ac709c8c653aca3cd1b7a67
zf21f937540d6bfe287e15bbd8a8abc9311159f6b665f96d4199d71aa5a8121fa1ab893e0fd307d
zf2058977f77e8e17cd07ba4bca468210a051f1fc81df524119422664e776cbab62c924f7de574e
z2c8cbdee0e6f402da421c4511f1c0cdf573f026fa9fcfd2edb28568a3ef0dd8a483840dc64d2c5
zb7fe297ff582eda7cd39dfffcad7bec095e1afe5af90dcda1bcf3a90cabae581cf8b75dd66a99a
zc0955e194477b9972c81ce3784369cb2e5676bb1444cb50c95f4719ffbde29b7b8f5c3157603d4
z07b8ca9172987339c527f8976a857092d1f8a55be8442aa76712660947c6855bcc6aec5f3c8db0
zc1e8744eb358fa44ba1aa8cfe7e7efdb27d07956c1ed95e99a757b2d98a5bba163d0f71fd38d0d
z13c26de89d91fd74697697259ab3f3a821bd76463d06ed1d53e6737f80f0eb3ffdb2efaab4becf
z107ed6d8b26320fa46d8c46ee3511014106df5f4fd3afe2634845ca58415d8715ab26e641ce13f
za1a1d58b4ee8623b7252df533fd3355982c458bd6a519279605a7afb793e695eff8b276b2d80f4
z9790f1bcb8339a45198d1c55b38d2303bb489fb0b85d02bb3b75b8b02b097060c3a23651e902c5
z1ac7f389ff993c1da9bf1ce485a5a4ef11187b9e43c41ab5546a91d61d88a9bad27521ceebf029
z394c51a215d922ea134bf28bec7792cfe7d406915c6bfa89d493a81ef986d27ce8caf7ad23576a
z3fecd46aaa0a4908f10f35e075d7925be4e7231b65806c80ff5a0d5a7353065ebd748e4720d703
z1c388a6a1a60907014d41a7344bd836983b5354c8e7febf16220f87a88bb79072654f7d6cdbcd9
zcd32e1985bbcf64820b905171ff3be87d183a474724fbcc032ccf1ccc8b188c81bc9293f4b66fc
zebc9d45c58e015407b611d207574e5bf42598db5268559da3f556116b6d8b6f89bfdd4a2f631c2
z0e18e9155cf9ca9d13e92af2cdfd3520549cf79934d789805960bb630fddd37b6383e5fdabbcd1
zdfc97ccf88a6fac8f3784f89ccbce8d04d92b4a76384db4ec4a0df0030c073641836d41134af0d
zcd7e5e98d3b506db094a3d9cfa0605fee5249601eb8089de05367b9f0d8d693aab7b6e342d3872
z4d9345c17b721abe35f35e5be70eb22dd42d1e6f68b512cdff3aa2edbecaaf6bb51ce2034b0b39
zaeaf441a28170e27015d54cf27283f33b05836a4b6a4332d3f3d6549c6a5e30c68540c7d9553b7
zb1919291e88843eac35c6cb2f1298a45bd4114362cba12f6560df825949add48799a4f6613fb9f
z856451130f23372f4ca525d1a6f408ff730974eea672debf6d7f3a542b704acc0b291b693d4617
z8f42aafd1f559502753ce127ef71be053476a96ade093af0727827f6621fd65669e82f080e6ff1
zb116f8d46e71e6ada67251c787e71af953c00b45327fd63be9369b09e098335dc649e7f4323461
z880dcabf46088cd39284e6281c3d6eaa8fe5e4dd7f9342ea6400c3d5e7304cc5daae407350a086
z777a04a3602cb63fc3c10344c9f8fcb7cfa168508db13b7836cad6e80d048e2da140057123e9f9
zfc387629e2535ac5fe580d0b217ffc0c4fb4470c2a9564ab733b9d44893f1d0c9ca8d5c7639d58
z450fe6d1b7ddeae79f1310c3d35b19a2be4ee7b7db48785591eb51f55d679579d36fe5007d6570
z84eda37684aea4d95dfab56b3408c81c161a53d360d2934e86297d6e67ea0a24afab27ee6d05a1
z6a7dc97cb133587f18c947aaeb4aabd05e2cfcd6d9ec28e277903515063329383fd09371b16c7f
z8f598ef8edfbbaed3234e0679ada1a9551940c19b9faaa96a1359805d7a3ef34fa26815c9d72aa
za73bce34694ec60bc4db6c6dcabdf23dcc3d58cba7adb86d4d26bfbf46b46685f96dfc4cd71759
z854f75e39241943f3a945effde846067f4d610ccb9a361dce3d83ceda65699b195ea40c43b16ce
z766081ca56cbe039509750c074b7deccd5d976360c244e30de0b0f05395391657f2115fe1da52c
z2f99df98ffab07c4ff6f738b556fc8e50cfb3552bc55e18a31e28e419eeac1e27568421b336d69
z12ce4684a09ed3d6e94466720ccaef8536a9b2c735d40f10be09563d394a911ae2b42e68a97cc3
z6c06d98c3261bc3fd574d6bc20a22bdced868c90940ed1e4dc2bdd36c6a3284aa2033a6c7b782f
zdc53ec6ddc373cd89d2e07aeb9ddee7148010a93c5fb14e685f19ed147af275e481b44d50e2237
z84697063ddaad6899b8f6cbb51f3658dd64d25cd776442a52d067d6195cb0fef78445a3f5e50e8
z66133b09167872a243d6426daa4e186f109c49689c9ba9e33b79a73de3851bd3938aa6e5cd992f
zead20653fdc81fcfa902e2f476b813bbd72da0fcd13f5d04e33d727412775a242944bc6018dfad
zcc5489dc2990656062dff922eacd586318ea7a91df8160e331b3db2b59277483f9644bfe3917e2
za52373a39b6974aa15dffb37ff3a442f82ca57439841252574a2e11b95f2468ae5f23cf1884261
z35cdf6714505076958ec25d9f99e7adc30da51a99d6d48d21ab53fb89c13dfc23c005722f88820
z18b47db35ca69f0ba0c7200d82b838ab20b37628deab8fc74364e8910562154804efc985b06485
z38dd78cdaab5b0a22da13339600a87eb81f1466a073e927727a3827cdd87c4d39d9e087bb33d8d
zde0571151f4ac51012490c67427d87e07470dd534945807ea613951a574bbd77ecd896bb7cf22e
z32c2b3c7475840b4a6b6fcda2e4155e2f4f19327c9e2d1ab987b4c5c4e563163276a703fc5800f
zd425f4c44f20eb920952ed47042cdf795fdae9c7eb7b2862f235ed6816d972d383d715c15a46c7
z21a0adebb354b2142f02e83734d20164a7b98052e25b11b9d866a39f54972e1ec50ccfee5c3f3f
z35fc63f857c87a2028c6ddc47c240732a127e323b4693c46cbfb9e1f1cfb1dafd96f006687dc9f
zf022f9b2c46ce0bd529b57d9266a554c3e7dcd95e5c4987705a74a590990c267f78318aaaac18a
z21028d3b351f48f75c33fb5890cfc2adb3138a4fa5b21fd8888cd21bcad1a9d6ae72ec338aad6d
z53c19e209424cd556e1d58a27bdb5b2049fa39d71f524c7030a66c8347a90d4546ab4298c3596b
z5bb65ff119b38c8d76e6efd569fd15d93400df187d0fc1da6323b793370aedb7466449047771d3
z741e14abb58c24969ba4edfcf54b691ddd3f82e92d828afb2d27b8212a80ca6e5c9872d3df8e24
z4d29debe0138aa3850cc189a5b065738f720cb981bca6ad325d705ee182b5345109d275b073035
zd400a5f1fc4a7d1be90a3a6a10b13313c063248ea969628f4fd0498b327cb26cf303275c239f9c
z141e09d247cfbede697fc35ff1f29b843fe16fbf20bc7e498f759eff5f1f186f6147b5a216c7b5
zb742e21f0e64099bc3c2ce77a7338e70bda8999be296afcf9000231366ad84b659d9a82a003d07
z5ebbe081c88fa12239d160c19e14aacf41f389dac2e0eb6b3840bd1f4bc910990d346a5647f858
z3d5e1039f3e937765d696fda3edcdda595e3a37e8af89984de00544b0bedeb7a54cb3346721c94
z9678772e6a9b92aaa2754427c7b2b7b8db8f698a1db0571c195d8da7ab1df03b04568ac4625700
z6033031ac3245b29ab28c83800951f69442e428dda4e3df234795c4aeb58f143ccd97e896b2a9c
z2b0360e7d41a03c39cbba3574b7d1421a9c5aed4da11efacd495d2403f47034a63f2b2152f2655
z0a2b5e628a244a956d1020655ebb312e815d53393092dd7e4a4f6cb38269f08986c3d4a816e9bd
zccf053a7c8842ab123f72bff49d4f60f1df4c921bcc35fe2e75c4e78b05e81d77062a84a0b3704
z57acdf21e4031178d681e324f50e48cfbbf6eec0d263da1528d8ab56df712062273b538410e3bf
z34b6ad29e7955d810f1e567ed34f35881e6ff24cbcb572ce107c1ebd9bb66c5a96fea583a0d373
z8b58e81321889e2c54108498d72b208e7fbf77a06876a256e05934349b3a88c1ec09fec61b09cc
z91e8236532e409fff9031ecbcd3c267d32fbf19ee57855488fe149074619716503de1ab027b6f8
z82f1636a65ba076950a465e562059f950a1853dee544dad39682108b4dadc602424556fee4c70c
za25a2b863aaf3010aa36129ffe08f6a6e3ea39693bd53f6634a0d45a4fdcb256289c2a0e9c2539
zc7032202d90d1aa46a471f2f4fcabf8968ede64a936c02ad7db3eece26f7946e2a813b95ad7a7a
zbbf1332da308586c9ab1b731b321b2cb424b80f2078fc00c8d051b622bf61b685edd28fc7b7621
z348e0901f54a3ce9cda8068ad9c92550377d7f2fab1cd80c22f33efa40cd4fccb7cfb802405225
z82d57bf24d73702e08cd2c0836ac6008384bd2d5da94a2844d8ef98bf0d8a1a2688f7d32a54034
z7e5813959ce3c015e352b3d2e701abba9ba8a196860bb22026d9edf3b0f05a55dc9c1402d92541
z6a48b22c9be23150cec99fc8e4b2e96541bd007552ef5b19c8b9346f84875d190b54886f32d309
z654277a70f93c5bbcab2bf233a14c522c6bf97a196352615499eb21ddb045fba3e3c97d579d528
z9bf48e72516f64d455beac5a9b6b98f00c18422a09a4eb654818c5b7473e978f82cd66b96287b2
z526fdf4499a238ac413b6c562d4f61843b754f99f12e50fbbd26b930c5762fed4c1618fa187d91
z0a5dd1456ee75f189d4312087d6dda24e4e45ba540ae9610ea027ba5f3f6deef4c27dd74ae4c90
zf86024be5bc1b66849f74e7217cb390401f19ec4d85b44ba56120231c25986c380c2315559dac9
zace8316ba0848d45c10f3928ebbed856c21a0d820343c2f9fb1f8456b3ae43ef6e397653e8c85a
ze10fde6753859d9dd053e40a3b12210494ca432387a498a0592e960527adbc6044498d11454e73
z0fbdec8bbcb6de1ba3fd294b3ca6b9705d3e12c00abbbdd2d4f71c68d6686beb6f3e0bfd3d17c5
z8a29a00f0c1bb52f851570d252a5e3aa717faf23516785e990f222578302bcaf9a8fe589f574ae
z3a3c42c7e21983d2bfd01d2b293c5e93c84c93921d39259560460c173e176b40001358f47760ed
zd37ec2c2444b458ffca9b2c71fa0668d61d3e268c823c383fcff8e28afcf190d19e839d269329c
z9bda89414a48ef8f055a16cef4c3a3fdbeb2b19b67f61b6c888d4b84c32901b85ba907bac2a84c
z56fa3060cdb4307ab8e0ab621e66c8831292ca89ff0fa6d5675b74375ba2804ae58447c9af4e32
z64c5b431ca74fc2d52b6af4fa16e15f7d9bacf5b859095467e7cd9fa5e4a15b2425ce10efa0353
z299e518961b142cafa075e2c095b5262c89db24cbaab2a3b91f1db75cbfab8a842a29fc6adc847
ze33283896719675b62af076d619e2a41462921548bdf84377512e9c9691ead835a74553e2a0eb6
z3e1aa37e035c37a16d50d3f56e375ba84222a19c5495c13818ac57de13119523bbd3882d9d5522
z1e27c649b3a058399f8bdf7a663991752f82949fc78645b47bda0760cdabefbe9a0db52cf0b912
z92490c51b6cfebff8d2d5b3dd5cb80b3417d24fed6dd3e0155c26ec0f323eb33bf24db3d4ee381
zb0e28f4fb982fad3b5ff36dde80d1bf68f0890360539b73a035ed219ba5842dce6e5cab76deda2
z64353aaa618fa8b517d1434dced7ee178a32142ba4ae96ee44d1b72ee362b9526f7074ca095d3f
z4b5fc5004d1f5f06a1fd7edb2a6cbb42521913df1d7f05bbe1456df957c072f711236eeb935ee8
z6e32d097f005d24416076ffb55a21fde0edcba804286a8b9dc3497d7d265b1e102fe5c3465c79c
z5f069dd99608325c4e5ba4d03ffd9070f1ea468f049a1391d52750d9a53f10e3c3e2380752d556
zdd9fbda8e30a3d4f2707e149d983364bc14f5cadee45b4bf803f9bfc77730c8ac7dd242334a9ed
za4e41d515925f6bc09c1234ef6ab3b740cf05340bb2102ee2f929c0e304399de3884d09d0c410d
zf1ce054c4353cac961e7c8a8424a66c707768c8746433992296a57d99b96c70946bd7e0d08097a
zfc3cacd9f44cd9e6cfc773dffed3c0dc25c270859a23941c09b1369b7d5b654b6f0fce8d416688
z03f48346204ccd9fbe79824de93c06dbbf2e8aa2161386746c24224e6a26bb12dcf64cd3756281
z188a530dc4b5fa93dfede1bece50075f32bd8e90d21da9adeaf28b12e499858cbee8855452df13
z114e8d60888c2daba9aa7cad9794e8262e51fd1954d88ba7d35d3099cf415737b401842fd49ba8
z7a3c48995da686605c94a0d00cc5ea973c320c0acb29678ef311344cc0e95001183f1e4080fb11
z7abc9abb43e4650593daaafbd5962fe768feaa2123dc5473435da31433f30e8cc14bcec57d551c
z641d8dc5a765c72db5a97d34c87421eac856fa30df282958ccecd14ccb080264d1ccabdc1a6f9f
zb130963133002d02af94788239b87344c09872b871e643bb0bb196e81d8c7d08bf90cfe89c1b14
zd13c23b0a09014cf6b64f0da5b2b43ccc7b7397c96731c8807453e6be81706b2548095e16e94f8
z3459d7df8b5bce7164e53715eb56c9ec9542a8b6a60e358627c69d0fbb373a2b187c84b02a789f
z48af3bb1c9f3e27e9f1cdcdd32608e877ffb06f577cb831d580b08e8386a580bff52499ffad872
zbb1996ca0644a6f67c8b70be7702f9422b66efcbe32a46f78f4c3934488556b202d914354d0ce4
za3c0e0428d76962080eda1979f1f37b45235a98fd4bdc8741707fb529d03a2dd35d3c17531b55b
zb51d9479906db3ec9d606ff30ae67bbde7bf6646d20761a0bf0797d5938c543819e024d26781c8
z7425a677e0c2984125f776a750d3caf33549daebcdfcc8fd0fed22b0846c8cb2c7c5d9cd1eec4d
zdbe76b47555bfb8f23d7b91522af25d537cfc64f7eb25c2729f35f40b57bc93ed484c1be646e23
ze6c13de7df68492eea8460199e1f34a9c34144cc4e9f08c5ddce483a3bc7c8e46ae7d491d05724
zf86ee5aa80fef784778c076c8017887808af9e292ad0b1d90a3071269f757cb83334d0ab167c9f
z3ebd2fd3de83edd01619a1e42539a3e771a91668c8f6c153448bbc2e24fb00575589f31586b694
z2ae01283cd2daf9f8407098724dba8ae17c7360b1c2e7067e2faf96585d00ec0ced1ef9774be04
zd7efc97dedf0d1ed00ead1795f19b457bb77f9cc426c6a685bcdd446b8165742fc02069acfeb79
z55587aa67368942af051a1b20fafca08549aab1bad4ea3305f3f9ffa0ed8593c602b9ed76c93ba
z729b8beabcfc6a2e047992a61a2e8aa435a325ea5d4425032629c7eee0832b3993ce198db9ef56
z568bc733b4579f69c3a336a208870a1e5de05a31826ff5eeaa190a5ff7602587de5cb939004586
zc26a9cd4f30027a1f5a01db2f588efb44e56ead86a2a29dc15b92403c619c3bca2855a02501750
z9398793e1dbbb56f7feb8c130c081fbfbf9948f6f67f33fae00d93d72e1bf00d5093c79565231b
z8f62aba3412e8e46032c5ce19ac9456821466c37ec5eb535066048c53b2587fa7e6d3b2201db04
z18b35def0eee5576064e9521092fc4533a67c50716a6dd2b6f6954c3e20ecf4fc4664456b6a7ca
z980cb6e364b96d8fbb1dbc3671ec68c675f876d2b2aea4d42b65f44abbb365744619f93e97c215
ze37b59f79d286b9e8128685bb0944777620adebf8b8be71e16cfc776f979aefa9bd09319708171
zf0003012469126ac0c143eeac50727112d09adc386e542208cbb4fc5ad8b7a857a8115451884bc
z504a725d32b30efb7fb3688d7b20bb750775bdd0c3a80e2c442fcc1adba2856c9c8204e86903e7
z0f5cd63c7f7b0b5090cd3fa07218cea8afb3f9b2b880345467dc508d9ddf54e88fdde551b5ab14
z0686fa6887d6f7b8f3fcb250e76c5dc90ec6ea3efd0d267af3a20c916703152bac2c8552daa4cf
z84106a7d714a0fe1484dc38b5f3f29dea9819f6361dd72d6a6aa57f62eb649c7f284a5c3caeb26
zc6b5881eb7de3a48085375715e7e9d0bbdd8c7f8dbf95ba47fea6e44a4a3d337d63177655273f5
z24aba6b04078d06cc372275a3a35ef2480865be8b378491006c5b8421bd253cb8ed83b1be3b019
zaefff603cdd8f38bce54371726aeb10d1141cf15db815c56d74000318dbfb43bd114229cf9d4bb
z038af932d203f045da07b6b0ae8cd89b8d6ee46bcb1b7c06813f7472ab3250f44c3f77a8e9da6c
zc64f0430afb8ab143eb5a4804468f190845e83cc7e4d0955843515c390abf6ff9ea257d0c00fc7
z8589a79348d2ccb4105dad6a4bb081958e99bb40d4d2ede4775752d3a8f7ae5925db8da5067d0d
z39b2fd34e9ff274d5b0238225bbf8799ff110ff01730c519c3c3deaabb8699afebbd2304176490
z345ba6420d6ffb482ebd9ab32cc8c159c39b250858462fd79d55f3af6fb7aaa9f7fa46dd708538
zd23b1db391c5fdb5c08ff068d383c64399b522c4af4588556ef17c3d93e4129d7bc42a81d2c00e
z92ba6bc7d7d91f8a9725a086fe79c720ddb22e1c6e0354cbad664c4bf65c541ef40a39818bdae8
z4efbc9d6f540f1860e91d0c18b4e66cda5a034caa7702540af9155eb8885d23c9b581d099b2bd8
z1ca68304900de1dbf9a7040c4d4949ad50fcbe41bdc27515338c0fab7b25ff0191548b863625ae
z3680bcb317e938d886aad49e281ed67dfdbc9ef5584e6be49b330672f401a69e04981459a0d372
ze47e97c0f5c547217498ebe12794883bae2d71da47bbb21163e3f83c1eddd0bad7a5b891b1164a
z56c01aeb25e711b2d4370687dd4fcfe98a0c716a14ca0e9850190ad46057cd758fe55d952f99e7
z44a89ea27752fa030121c082662460d0a555ed89abf276331e1bb0859b81c2e01c933ad6d37370
zc1428541134f689547ad8a0dac7cd45a69af116c1f2ed404d18db0c484fd721e132541c4779982
z7c26348d58aef5537d8637560aea3ae0809c8879f73ffcdf8e8c5c2a09a40ed4bf194d24ffa95d
z8efa1b46ad1a1e05a8508e6a5c515e813780c7475b81e68dcd7b8a9048e09c8c5d68918416ff4c
zd5178868a6f03f9bbc195ab70238ef9a2e19ea08efc0aff7a284b7645cf2e9b29f3c0d597efd46
z2f4ccce45497c2c0d13ee0e3a37640dbb0b399caf7ebdcbf0fa32cdd151987fcb96ac9be20c349
z506d05143bd01de7ab065edd023ad6d62366c4879b4470e9f3a96b3d6d68bc3968bedf7d5750bd
z886dc2fd0da5216cb16658d54f5a2654c2fcf95962a36e43d5265498bd741738cae61495e090d8
z081bee40fe2bd4c05e24c829153644a41944bfdc00cf55604dd702deb8b3f433e5ee87a6c727da
z53be4fb72c23d875b2ce0e406140d1192c4c074daa24c8643e64c5899d947dd970cab3127ff79d
ze5962f29ab72a57f827b9eaa9d23e937f27e0579cd44dbace428e5d68948f162580d9dfaf02d72
zb9d93ac12ab294a76bf65878d87075a68bf53453984958554723aad80b302ab33ac4dd588e52b7
z0cf72a49bed1ca71601421ce1ec95442a613a07371b381f5158427d51b31adc53d44208ac96e56
z764162878a5ef12f7a21433d57a2aa76c1d2561401f97c7e03908c277fa6b04f5c0e3a92415835
zd59bafe70a8b58eec32a1aafaef6106081553d9f04414611a93cadefccf4da401e44d106d3cff5
z78d56723200414d82496e6cb33112375bf928438f02de7fe09c853031e85e3d788a3fe1f901669
z4e610f459ca03c69275bbebcbaef089e4ef64cd45081bc6ba67e3fcae71a384e96b627c460085d
z8dd6d2a9757d39e743e58dd38e6d75c962c7066919425db19dfc0fd28591e06da08bb58258af2b
za94c023fdd02384b256ed39a6447988d558bf9d4c7ab67ae6c2ae2cd9de49a7e26ef5d5657056f
z44045980c664b6f022f90ef50a8a67798c7d55087898d7ad61e1f5b1d668a8c4bb1e362cf6d325
zbba8d934862cadd793f789921fa003b3511c488b51d53c70228df9fb83b38f3f773c25b7bd7cf5
z76fdd84e0310e1b67b33a71d389e93e1eb6a1fdad3efbe401258e39cbb2ae8702315d00cbcea94
z0fddca46bdcf2f20c63c5d1f8ce53e76a132e0eec3d0e519a222c516d17a89739b2e566c897c46
zd9e75c451d7d5f46b8a69193377d386f28dc30c684a3352e35cadea02dca39dd3ff38294b1c898
zf64c59ce8b660da249f63f0495efea049abc4c9248b81749d462e26241b38b1f8aff0363f78c37
z9bb1397dfd3047c62b6408a2aeac0a0e29c943768b6129f9315df5ff33177c57e7a8fdca05d78e
z7401afccdc6009db674128b22c2b873d5bbcc79a1c9ea1b7b7916ec9b4ec885f4013fc37206f78
z3968364400ee1dd76a704dc2b6d577b1941bf88564311f96ef8b4cbcc8ad2b61aa022d76159e98
z21c48f27afb159c743620ee29d96e1c8bfbb4ed025065150061c117cad139e72e022dde28ef18f
zd0553d2dd401c2afec32e68c1c44c533c81b9d5dd22861eea23359c0e049c6ad7cedacf0a77a29
z40610312ec426c30b3afa591d9cb28a45ebbbcaa693185a79a892afc605a73cede1f45cec63636
z57415519c830e68aad3f17c80b56aa8c3490340f9a86d6cbc22aec0e3180563a76414d3b957beb
z673bea6b2fb11fa7f20bf05d787c43a8e1511a7e08756f38c5d85cae3deb0501baaf55cc3401ec
zec0c2008401391b54f0f5f7473d11ddb8fa1b5fe155dbc8ae79f0f9e4183cb042a5a9208c3c474
z898ae54e1e811ce04b2e7cbaf70520f5cc38fc46fe69d384c64a19a7e0e37d6174bee19bb594db
z5472ed06701f589d3612b9e55e16570edaac868e08cd475c939f1f3b01d1da26a462182be6770b
z01dc5a7a8b868aebf679b9af561f138c6364d7a481bad060073a88cfe1516de9e9721a282121da
z2058e6eabc353e8f9516b38bb4b5a316eb0228e7ed5ad523b50db988768647d872ad612cca4025
z1e6916115646dfcc50f48b01b09b5bc25e2be192506d1574922860cd0d36ab3551c2ea883a6af0
zdf8b3287a1d165ab0974504fbb10a67d0cdde100981fd29c1a9cf6e1cc3223ebce0275193823f5
z94c1b88b9cd245fc08f0e418e3df48bbf60d9cb4ab09d4ec53af81a17acddf5780f1414787ec15
z62875b39aab4206e472b428c7070e62aa1cede02afa5d6d4e6a8d2c21e32fbfa4232b0f92e944b
z3e06bc6b35c960f60156794f1c19903a3fbd3eda5d1dc47d58a4d4eeaa13694a2c32765e1da896
z8e50d604490230d3e688ced6d33054ed5f455da19d7e1ffa9db87baf9ad0f116cb4138b4eacfe8
zcd275d34ff484aa7079b19971d37ff846745ec25a47071a8fab944dead6a27daf6b9174455020b
z2c57c515c1639819ccae6f8e2eff394e1d233eb578631a0e960610f27582f3d59b6ff7cc014a5b
z6234735337809d89d6a17aa41b5370eb1360bcc048f6c2d75a57af2ee42133187885b1b85d2c82
zeb135d70e12160ed08079737b45c33317ce8e8222801fad3a6149efae25a4d967da35917fc375d
z3eaeee23a0ab1710829795e88cb1be661c3fd052601dec271acdb8772d44aa00c725662a947097
z137b71fe8818ceeb9609e3ef57f51618125702879901e1ee72ac7d7c2332384e3ee3a26568ac3e
zadfe16f8bffcd69fe0566e4d99ad18f1e9a36afe39955d8832630736ecb347ec1e7a6da31548d7
z66ea22b78d321e44492396dd7ab97441e7abef116b4b567cbed039dc4ccebc3078cf780f3aed63
z2bb6e490f2fe428b55392087da384d09cd3070baabee26ee94c89f48c8e39c5e38c40061b96862
z874ad90280460bddbf45b49c84aa6b06e33627f6062679c204e20880a3c0dfd9ebc58dc6c4d408
zeab251f7b405a42df80c5f7eb279cf7a5cf6016504488c45cd411b52bc7fd3ad2b1ba5176a287a
z14d4f87945a61d5e26119b9d3eb21f86b30367f9711a9049fe0939c7fe66ccbd04036f2ab340d4
z7b3c6ceae1927464ea2b38980e540f4cd82e1ccc9b3c9d2bee2760d4d3aa8229895924be066eb5
z43e9eb4a201b84854299d8b98a9c3ffbd9a80a01fed129ddf51f3bc63692c1c1f7c6fe151e5cc8
z2aab3d7129db2e1de35472e4d98b95100f4eb2cae65d8c85cf5b90a83634e8fd88e1da3feb3c59
z7c472668f14d49b2d6a03219b6b4bdb7ad873df955a34072a827f10468d2160232b1670061d969
z527babe6c6da3c7ab75c0f591c9ebee4a887e36060d3ed605a811540b5a81349da10cf5cf582ec
zeabbc4b0e2b2453566e4c370efd4e49414c6260cb32213cfe295df4dc31681afdb18c81a740ede
zf2a82a98498c7eea892b4345f41a224f3d99a51c8a61f22922308f23612462775fb982624033aa
zf833ef27d1d61cb01490ba1ce1306f6acacceb547a97267eb9d5043fe86cee6740d6f3ececc0b5
z0ba5e97c713f81632ec75ef187e7f311de8304d320f0002c45fd173239a974c4159e0ca6be2c3b
z79268eec16a01d04c5d8b67d4c75a29275cb4e66454b014c8a1c043783c0d45288af84b49e1808
z28743f1127f4d2772cf3ae268dcf9ee1eaf0b46aab896a939ced9dfffcfa0997cafa50439f425a
z1812658bc419520ba8e504dfe703751e7a5c681eca3a5c9912b6c6a10127ab80c773bf984264c9
zf61da414f5ccf0faca6c9ee0f34a61a307871605b867c635cb171e3d30fbad161fc69535e9df17
z77744db2718a400bd3c383c60ff921b5b4428ad3e8f830630022dc1dbe0e34311d38b3fa53ef4d
z35f173af97a9c355bd532fb28fd373cfec8f6cdba8e0251c120125a92de09e8b219d808340e7b7
zfeac565566cfb86d015e154a43d5444e7de3466c1bf5a48e4ad78ef4fdf4772d63f8aadd1db682
zc6fcc52d0488911022f6679bce4a4a68a7649fe1b4c0a5eb1a8fca1e8ef17e70819e2907882112
z41b20d55cd32a9b1916c8956820f426ab01939a6bb5540d0195f11edd761bdbd66a43d389a113e
z01deacd56b603f50c0d34b7d08122086b96bf6dbb10d0c63e942f07e19959ff408955fe8d4d579
ze5d439bc19a2aa46c49a5a00e3c82ce345c9cffc9c6ad0c77a53d0ab3a4c581a946b912c02a8d2
z213f81f5c04e4cf307543129ea3e79564bb238b00f44ed40180f63c9c80a87857206497bdfac64
za02bd1fa8d74d2707918b1b4ede034946bddde9fd3a280ce4b6214d3b8ba7c0f62922c3dc75ca6
zc46a4d2297e295d9e1396461fbc54c86f7860c20ead7692d6584021f7a27e38cde42a9346c92d7
z8bf2b0fafcfcd28cf216ef9bbf6c4a12d68e209bcf4c78ba567ea21c0be08ef87e6584eb9b8a7e
z1c01fc055f91133ad0563087183b1eec5f45753cb31de0f8181aa5d29659b5a8b079ec0301c438
z7f5ca1f85f9d51cba490a8d5bb09e646cefddd941bfe70573de92888c47d2a8c34ae6c7bdd104f
z0589eebc1b263dc313c9389944d0d3254c1a117e0613f59dd8b19525de7f70c2c7aa97b6ca15f9
zc4cedc501b3abe94d73e281a5836145d1e0db269741b954febbddb73f41a8c1ec0d1ed92c029c2
zaa471efbbaf462f806a7cf8821531ff83cb4b1d6b987f03419c93d38364c329fc68062ea18a1fe
z4e40c2ea73b84cacef8cc2667b92abdbdf025b9e86bc0cf4f20458634044d71af76b3462903c57
z70fd2bb0beacc16d839adcaa899f3281834785aef840a0f3f6ab75639a65f44ea18a0f3b50112d
ze79c8c7b754f818b7febf59a2db32d878a7512cd9a67e09787818b281b5b888b6f21889e6ff200
zcf427c25a29575238e41cf3b1597357bd7b6b0277b1d5b2609381e67bb773cf9bf2eb69146398e
z6934f5ed86e5ff2983b7be6b96700dc66bd816c273481170d3d965180a1960b09748927538f2e1
z87717c45795b4fb2118d0355e321721c5b5cee5d4dc5c76849e240d31060bd461f00cce2fdea9c
z4f8ac2e69b0bd8126d08169b769ee9bf477392a2ec83f81b932a2bc677001da96cdf2c30f39d94
z017a7bc31f83c417d9448e7f200e29328e5b9a35a5fb308a172893cc7c342841de8ec92e6e9527
z46c5804e1c6b33f6aa195346370ef0c9bc762e42fea9dad15863bb31490b3095061d00717a6e61
z59ef16d29ee50d048f5f726fe6456cd2fa3fc89d6de2a7a6e0681f8ad170408d91a03ce12945a3
z998e9adcf0116b4a34e61bfb3bd3b6db06b41490e076b00ecca5fd7d9e8a7a27581e7975aa575c
z8056f750565a26503c87788e5a63f0706f30dcf2390f3ca9d3e5ae0805ff4dc23919e3cba9d68e
z583e393540a9f1f23fa753249d83076746c1e6708acf257f008e838684d919985904535aa04b53
zb066a5cf9ded52597df6bc5aab39314d03f193f5235cbea4477f1f928773a5d0fd1954717ae00f
zd37b84d127db0eeabaca265596da6f8e62023527bb004bf39388e53846f6a98ebdc89e53930f58
z3af3b04e65f02285b0478a97cfe8777dbebca4ee824a45c41297cbb28b386f8a0d2fdd4ae17199
z0389e5354cf54844ad7caf93c867600229c50be1235a8334a0ed104979da7ec2bd0583fd6b2d67
z518f4e6d6adc65f6b7fd2e67b480002b56ed3d04fb289f29f59b47189a022471b1c97ccf647857
z17404a3781d07ad9fd11456f6b65fcb9ab6b4f47aacbcbb2144394323b2ae74ef613a43c7e07d5
z1de2f918d1fb15c2ddfe36ba77d830f8c01217de29308ef779d7b783e0b2f1399ba78c7089447f
zefe8867ab113a084d0ec3830fe40d4fbc0e84fa7f85e7d653df2193bfa857e4d1f103f7cffd0d6
zda2b21313b958d67aa14c24c11f3e4c652c990cb453841dd8fecce151047c6b6132cedde846cdf
zb0236b48c15dc5c5ffa97a3f4edadd0e8c696f59fcf32159438676ba227302e74461828fc1a711
z4e8df7fa1e860379b9b7d8a1a41bea982a5609ab2d373cb8b45cd96f371527ab6f09fcdaa41c8b
z38297e27ed8a626932c80377301d886672dcc6815ce385c565a00154842102b7fabe2032bde00e
z8610464a977a69101dd198c823c3bc657eb92821fe3ad06ec62712c1bb6b69fa8f8b8ba24bc101
z9220a8dbfd941f6a6e1d0de4ab362708825363baa6b3c9c625583098ae88853e2f03e8618db064
z18966f5c745044b5321e39da48886cd6af260b04f9461fa3ce4fe0588f246a995635a03e4f53c4
z0729d9a52b4a4a9c6379df7fe4cf00ad9837f1c565fbc425ede9d655d6d6feb6097cb7d18cad37
zc2bbe8e3678713f2815da7a06f3ef24c8131059cc0056d1f0124aa0f5a996b2dedb4f710d7a25d
z97249ebde294d7f4c6b853b39229306ddf6a1ef40c00aeff2468a99934375bc13a929a9e6373c9
z35dc6fe59b22f7f658cb349aab7e180174f913cdb8c9e3e54e84688ecbd465e1921c873c574212
z63ec716bff897e805c0d50735227f9887e4d0fa0e6e3c5e24913bf62976f04cbbdbfa4a1a02a83
z07d1ca958a1e9812ba4806b3f585405a1c3a97d790d867963e719cb7886410a490dcd9ffd0f333
zf99e909ca1ed6b17fffb52e4a96f2dd5bd216c9c3c4458e7beb70ab6bf41965fd3672ab622a7f9
ze2215acea671e856b4ac1d8756cca3142c6176833d9b22d73e3396329fd0f82d673242c503cb68
z2696e385574331e0ec8fefb9f4dd7c7b59e516db89ce7e30db15506d89c3305599ca17f9406116
z05f1f23dff7abb52398c2454555b3650f144f820c50bfd966f56e4db6435c14229a7c7c570168e
z883d54bd7c069e990f14877711e8e23caa387085e3c494d35a416c064a768fd7bb55903b256e2c
z0b3da3a7845b054480a4749fa0ba6802eab7b36cae70cd7070ba6f1405300dfca49cfb300203be
zd9b002c5667a6ac0452f53baa6b2fda9d8a37bbea6fb517f189692510d9aa9cf2f25e1bd9f9525
z614367490da0fbaa7bcd0ebaff614db45a893acb68c56efd549a467c814201b435cbaa5773dfec
z0e5af277d721a16dd7baa9bcc265197062f16dac5715c40b0f5faa2fda4c114ef722a474b8c4ce
zf0d74dbd1f9a8dd1989d553c77edd90d27b2a8489f103df014f0c22c32d71946fda6559020737e
z05dd218aab7d52292ab7652142f176c570ea9db47055a1b4fbc42c95c1e7bf528d1029cfae8d77
z99561e4f41baa246f84bb2dff6e0c443c4bf0e37538dd73ec4a48d1484574878e293908fd2d47f
zc9090d314c881e2bb3351fce896b6a23220004864d7c16a9de699a17edab546ddf08f34083c201
zb67d6ff1588d496434c85184074c1330e5e2a86ada6bdb25ba6252b848ba79e3dafbe209a026ba
z14783eb4f258301c79affcc19552e68e486bd77d78c8a78cd263a9afe2c684395fe1250e4efb17
z3fa624e8bc0e4757839d63d003739ce0d2d0444adec97c0f49353c2fa8f4b7311f22c89b5f10d6
zb86c0627d5a38071312c33c0c9dcefd9b7a3a756fcdeff94f03eaa13f906a996b9dab9e9206a40
zb21a37f9d60bcc6520e8d5a3bfd246705522c90dc631dfdba1ac4970f761e005d53f58b6aea1cd
ze2a71fc544e2d4a3b4986847b61167114664bdb6016832adcb6c83f3668b4288198a4bc80daa20
z96e813def94807bffb93d40e7cb4f6958c7eb26a0e29558af09c6db3693ab6af4b49b3784277ea
zbe370a51913581aa1ac4ec8fd1cd65a456880ac5784b2e004d25f9f17c3634cc61441811e90b7c
z3d88e13fa85bd75fe56667343709671e8735785f69f7f235276a86b450a20d178582a8023da7c4
z1514f4b5d40afd9b0582a814441a3f3865b558669a66d4b6a9a6c0689de90ea738193374441e3d
z7c09def143089ec74e5c6dfbdd5a9cc4237a44e8d838a54a989fe429010ba640586ce703247e0f
z5c8208e0d2348885750415c8f35fc6a2004b778b598e9509cd384f19f5f7b3fe15f73cf7073a69
zac2487596a48356520099cfe9ef881368f79276f500085cb65675b1a6fe26be72f06d5e84c9d6b
zcd3f3763243aa920a6519759283eebece9331cbb6b756fe8f55567b7105daf4efdf69f37022c36
z491df557aa009338c08e893579aba239d1a1a8c31e7f9a864d555ad8dd8b386de972b2f8739908
z4834bad86bf0a0173d5c876b26bc7761dc26b57d57b60c89112164da5a28b5595311e0eb33ad2d
zf5f9a4bedf956a4b913089ed64fbbf3d581c51f3b941d59192f82db0c34281fee38b8d7036aff7
zc8b89636980a9139a6ee2cb4cbc244faed2e0bef59938f6e7fa7fd09360bf411abb1622035758f
z2e0ad7c165ed1831450eef213d20123d04c862044387ff4b8078b6f8abfa2ab5f39fbde20ea3f0
z182cf792af69041a8add5fb794eae15529d8a8d023c069fc6f9858fc2437ae4f7f97e45385ec65
z73f01d4597681e296074fa91d54297c507491d5b4e9f0c29ca8346a9ae97378aa65b1298a95573
z7ac9e405965157116c41adb3793a050cc57eadfa6b6d3ea00434fb3c32068695de6accf1bf1bbb
z1118e2803ac4219305538ef76f4d5c9f8dac5a30e2a873eb0362427956e2fec60759bd7c8943ef
zaaf4d914f699819e8c0c6f2c7087dcfebb380591b420ce4e11f8ccc4228aebd6f721f74b1e201c
z7378563c080ed613c6e2b7d2e7f6a3329db73374a559791c6368822d5b04450dc0d23847382a0c
z3e92070ba70c09f8610b4e7683b742c8f81ba928c7caa9282cc27bd2d47018d10a3be4347713f1
z092cda38ea6891b2964f66183c47ac1b4ca2a9cba7a18997e47c57fb3aea9bca1f42cc43053011
z0d9466487bb0561ab9b7d85979289daeb1128b23a0635a1c551b6aa1d104ac8b400b8237d0d109
ze8da0ef802d56d4f74bcdb8625b95d5e055bec9e0631a53be0ef34315af34c537576016ea8f5b6
z662189f0e1f437906a35f61c16bae9591d3da63ca5d0962f8417113fa82c7d5f1db83a68489472
z79a1e22292c6ffbf5de7d50650869318e14bf00760da8f3728de81769f6e4379afeb91bbe47d78
ze2ba3ae7b3d56784bb890513ac08189b6bdefe1a291b054a4dfc62a08defccd977e603dc7d15dc
za67e6f77d95653682824787457c8893c309ba0056f81a72615e1f641c5cab03da09456ef94b408
zb1afd23a618d04a6d1182242deb54fe47d5573f016604e40b346ca5752cc398acafcfceda24a5f
z64f14413d23bccaa7f7e59e664ff134377516ddab5a7512edea93f9f2f1ba30e10703911faf860
zd092c58cf2d390f993b295e6194d17c3b3aebb16b19f7871b8c1b6742485a9ee82af8fb7c49d34
z1b5f8889cc8502b898ad18e8fafdd1a96d945e25c4eadfe90877f2c35a2922e8093c5d7c0e5105
z04f21c9050afcea0289d374120774155071a23272d7b4f544b119f2d557414a315eac94a0155b1
z84b639106e6c355d70844e5ce06df19084bd128ab28ba70746b6c0cc2c50f9919e0ba733bb169e
z973ff4f68fc5bc9f1ceb78e3c1f688586cc9d5c4169f2516d3d2afe9399ec53bea1bd85c049a10
zd5c2ff7bc818c271626eb32b0a5fec840993672607e137c04a07d17706557c7b739769d766d2f2
zd6cdefba3840cae2ecdd84146d1e163f53d84ae2425349057f90c189f2f1a4639029964d2b0bf9
zcd8c9451ee29772f7d690623e74073e567716a32f57e966a0d39b4f4853b5528879c409eea65af
zc385f4287b31e49941123a9873e4b12700d4872c59b1f34291ba8461841e05d6dd3a32e5d94fae
zaf7b70255bbdb9e86cdb8f33b716e15b86c08f47b325b54e01d67f13681deacee7a99a0013a359
z5538836d19bfcbf67a54f49262c134b29050263ce6bcd855fb585dc0092aa698c0446123bc8cdc
zd84f41b654180070b9215b1cea5190cd5f0d5bddb698ce4c40d8f5b6255706337f479e5ddbca30
z2ccbba213d5b3ff73f1f8ff2c52e80575579b22b364019374cac71d542a27920f4665a72ca4604
z1ced9fb15daaec2778dc32e7fb847e686decb0e33cbbf27fa8b851314278398772b74fbfbf3af5
z9d502c5b5db62b5bf812a250b1e761f7b7356f3dd7d2677ab82654ffcedd3a6713a9f3e6dda1ad
z43a9ed8e6e1526e11ee1454a1b2b915fa8fc03cce75c3a8c8ba4c7583bacc63db8813555de5f01
z4c0bb6de351d4228ad42cec13cd107e949936fd16d2aa85dc5d992de914631ba1186399ed32b41
zdc4e9e7e204a7c46fa9a53c05746d07705a35ab8fbefdcd30bfc798a89c801000368d54be50975
zfcb088ec18e0269cf6f56a44dc0bd4e48bc6d16dc27198e52ee053bdd3abcb65f59c4f86a93771
z784a7ab91a5b6d2007bd7f6ef1c99aab76730b3d2fd156d2b13a4e04c1d1800215779813e8946f
z65a85a62fcc99bf0c20b097dad1d7a8857975d253d0434e2a27687d2391f26899f6a3b61da7c7d
zf5fcf9923b6d588c46595b0f3c3f60fffd1ba4c8de74949ec6e3e6689a22f4351ee1032e26a693
za38f1d99096690e278317c415153cfa1b7c7fb4d9bf77c548a45bfd2e18d40aed79e13088511e2
z82ec493d56fc1cf498e5347f2eea3f09d9bc41b5a82a1909b4c921c401fdbb14869c8c93917451
z1aaddd87b541ea6c0fffcdbf49c3abd081d1d428c11ae06701cf5ecd82fcaa1477af7ebc13e7e7
za739cafddd21508b7bc14295cb00c48eb668d9daf3cafde5b3fbed8c53d4598caaaefff9ac3dae
z0d3489771fac83d964a12fd89d50772c5b83d15c86f0acdafbbbd9882ce49ae3c3ba85c3c12ccf
zde697450526531d8d855f7feafe0f34eba4963ef8d9b1b2efba6ec5db72bdacaf7e61fdce2c95f
z15d0b44d3669eca117d90b9d20a9f4070f183ca7fd833877f480aeaa04a73368626576b817d071
z40def831733554334f19173796a6396ba6d3197fcf7e4ab0b21451bdd1f5799f99b0f0a99f8655
za11c6ddb598b40d2b02939f8f70bd20e3ddb0841cd9cfc56228699f559e6e9df87c0674b6c0e3b
z74df45d7b22a2b0e258aa8739abd20734da63ba3c6dd5c3e6262e04e2a32b26cb29bc06815c3c5
z46cfd6d41871262c7e3fe8e3785b0e1f661f459d3f656f23bdb3db93b37a2316b340ada3f93479
z0c3b28e1daacb3bc4b9e0aaa0c601c0aff25b8f7f9f6ca34c92ab799ca8679d388a808ae246de4
z2564cab8d297d11872d6d2ee3e550ebbcb6230e365afc394160fd891ddc971053b1fe01fd89404
z0cfa28c43352e100406094a0f40709ad4f55db253f510c6a513394aeaa06a9a76616bc607386b4
z3ccda0ce3b93ebb9d05d866484de03129f2c009e9ed36580842f5e3ffd7a2c9cf0871e5c0268b6
zf646eca92ab0fbb78b929d387ffadb3da64080236e9be8606c2f7587a1f8379a28d585685d98b9
z90abb363d1d804553f2a81f4dc8dcb0b5febec491f3335b565360957d509b77d7ea9f881c50eb0
z45528dd9627fa97d2bfc6d5ecd3de5e2ccdbd930c9541871bc4ee0d32e0eba46bb8b4b58b41065
z86dc2c9e77f7a75ed32dfcbc2c41b94e5520db6acb97614211a3cbd0197ead586bdff6437084d9
zcd44935b7309f69067c639b6651d6f4769d576a6487914f61f2adace7f6f63c5eeb2bce439632f
ze2d9c020837c4d90c2e94a30e43e592f3ed3eab553d6fac4200622aae41ee417bb402906305180
zb9dc0cdb6997ede45100bd99fd972d22640fb8dbc8b5bc73118076ebc2898e6af4e7e0c5bffd33
zc4136ad1aa12d9a8874ba5be0c990d47209d4d7926a24b5c2a6e6b7c57262716a3837060e49ba2
z62490c00a4ff8d0dc23b47a32222c124c1a031c2a6cbf1b14808684292739426f0a593515d3f04
z0fe3da19c8cfb7eb6a2dd80db94611c44ea0cee0b804a65ff3fa658b1e51b230cfa3bdea3da8b7
za86906730556032af7dd88010afa857599b8d83f89d518f9ca5405eb7fa232994fffa76a2893d0
z950b1922fc5290bf7701ca511236bcf00239d1d02213b36597a8414885c3edeb2247741a55617c
z062896e96d9c2fc5a6fd5cd15d6458822a0a41e027c6550613194d61a2bbc84a22a32e96e684c2
zd66a31e0ede5155fddcbc7516e0b5d81cbf596bf3452efaa5b5ea39723fcf762cff9ac5cab3bc8
z8dfff783cc5530d553f67eb31a9dd3539c333a52765789b6d80b89478b2c6472b785040abaf5b4
z6d4f98d1677b2d2885551c43b0a57ab191ee0dae68354d3aaafa7320a2827280a5b95e90c2a8a0
zb5a6ae18e12e795020efc9b03584a356c2d091161f030df77980231951cd48cad94ce046df76b7
zab97ef19e2aa8704de550e3f9a54640fdcd62fd9b5fb537dda100dfc94f5f6a315c65b1d136810
z687dbf1ca5eda309b267308ac3c687d9585ed24063ce5bc74ede54041b82437407b5c86cd52850
zc732d0f540c8e13bafac4c3a510051ab75aaa6c5602c9fdc5feafe6cf3201aa69142e3276deb5b
z84f670bf70065990150b24a05970abc5c666c6dc92b54a4a69f4da9c844c47712fc17c62ea06e7
z3cfef8f58d95ffc831e7a8051cc35fc555ddfa57a08f2cfd355f980dd9a791ce2fe05b3ec8b5b6
zad94bb2d7bab379042a0d70796b68957e9780f92536ea3ef34ef1ef99fafd7a2a82098838b94bd
z1603232a1ab69eeabfa161419df655db1f282b35166336d505e60c4b4545b0d95253ccc5368ddd
z2c9d1146d4f2381a52b0ad99fa78ff5c3f89c73fb6e3695ad1ad9c5f5ef155acfbe0ccb04d6c7b
z363951da3052af16700e17196de1d0b1e067a9826db86b863d2c8660081639216214649ca1b681
z815f3c3b054fe0a6741052d007a1fc25a234dffb30386245e04bb41f0ad9f7f961fba3fcfcbade
z2d479f7909f8bbf8a31e2805212736dc4b01c4b8206cde6b14655edf38bb7eacbaef7e4956213b
z7285bc6b9c403f7fe6845a1d46325ffbffcc59f923104ee6615aef4b09d432d82a6c414e310bc0
z95b69d3b465c0052bb677229a7c73f92ca7234dffb6f44c3254d461654cc3ef0967afdd24267e3
zb6d0630d2471eb9bff538b2ac371ac6a507d5441294addb8ecd7304b2d9f9fab82f3fbcd6f66b0
z7fc2a2cdb332f254f84e5f7fcd9caa4eda376eac23e3ad239c9ae588cc9a304e7f0abea19e1803
zd466ef86b3238891678e4812334ea1a2eb69e0afcb92e522c6ccc31bf13bc1948d12012dfe9688
z744b151bd44c7348e5a9f9bed1ffa946be7d29ac76b9f236f906e257958b2fc64d4b28c966c5d4
z953be97f11a02e192ca2578b34b427d40cefa3ac2ad349d510bdcc178a7449d85416fcfcf735c6
z2c931c32cb0a0321c92669e859150fd19437aae0cffdf75ea8297125d245a8820bcfcdb4727830
z896399e218114e63a25d9aa681ceeed4a0541104e16d4662678d672e6f53db9d34d110d8c1e729
z418257b8b9f71f4d77397c90ce5ed7bd7f3e3e6a606206aac7f74a2f02a707b7e6e67e8c5b8015
z1f4ca076ea7a21e85a5e027db24ac1be4f9c76cfe6dd3868f648686553ed6a6660edd7a90fb6a5
z3f1388f766526e21908dbefb5729f6cd2b0e8b550fc51e8ecb8e609914be9306cf1374e51de524
zd00a6bcd7a51a92fd2d6833c6b15d5c8f43b350aed849b34cc80ed2963b1a424d3d0584875695a
zcc936a434546d31c9319e168b2009284c2299c408a8acd2441cddaf6b92f2bfcacd7b2d00fb59b
za8779a479acaa6e8a1f08ecae6f9c0b87e36dd69bf4e657bc99684643fd6ff283d275b4f778176
zb48c41202575ba2076f7046c33428c498cbf7a2a7bc2952135c10891f5d158780418b151bc89ef
zb826fef4cc677b8bbbbd6043b5f08ca65fec5f24334765b5099a4e33f2efb4bb7aefb449dbcf6e
z9850fa09b832f0d9754db0ee51d130fc6abdd5bb2f2bf9051e70482334dfca2f6864e81a972f4e
z60311928b723ef4984af059ecac7817d55966c61595fddc5bab10c806c08cae04c94f0d8d98c1d
zc053898a267d14525bf97630f5094cc66e1536b62ff83a37c7256d123591c0128e9832ea55c634
z23aabdc55d7ae6ca70bdfa3585dcb94c518dc5c234c5fb45b7b3d8413c821650e662e63ddd8c05
ze80cc643104add30ad29ed4b8872713a105ea2d698024745bf04e42cc157be8957781adef82b08
z1a27d5ef4490b3fd8b2a264cb559318319f9b5dca49b8709d7b4ae8ec1b889da3c633fff14df72
z7e11fc79f961e23c1098d923e174a498aa7c2fc2fe93250d22d1fd1670f8825f153f084bebdac9
z1db8acbfee876f4a3ce8d93fda4e825ba102fde76de2324a63c4665d25381fbe616906265b9e52
z797b78d7ed664d18917f450fef83ed2fffa9c4aabee0036b7a8bb33612babc0436e5c04e80376e
z600ff0fa1528cf0133134f7dc3d14cc1e6ea9398a303a5cf9a83a92fb32a3f64d1ed52deb0f16c
z65aac345c2e52144ccd6214d3332fe01ceea0b9cb9617d81b4c5a24ce10e1ae192ca929f9e9463
z58d4086d5add66096dcdb400d2ca4881bb87c83f6a9fa368b93ccf82c5bcaa91094d6b19ee2bf8
z261d1fbe0df55e59bfe59756a3a1e6dcb0303139d8554e74604ee2dbac36dedb04abf7eef4e514
zfeb5c85d9e76ea2dbeb3b441a8cc0f807166c8c6b5a35ac142ce00b4d3e75b2fff708e7df391c3
z8059f3bc44089e0be57126916c37fdf25db90cf0d3a44c5f33981ea3e3e3a293f7b07757d45806
z3bd81e2cb85cc09525dace39351dc4ff493aaf18c9d5a8a72c672833316ddec4d794e2c03af683
zf29613acbbf6892ca088b563a455712ee076f21adfe47df4f1bc412e36fde70be7bde75f14077d
z0fa90b0203390825fde5f6fa85891691eabf707ca379b46adffbeeecd0404bff6d18beb35fd0c4
z890ac575ee02c0e045de2645dcbf6afac2fcb426e3d7cb88e7a2b2403121929186a111b984f01b
z3684da2609d13bc5d1f788f02bc860db949ca2e642a4f51d4801155a8115d250f894ef0e3d200c
z6143b863fe3eae051dcd2ea0058d642fff57d6d57978fb71dcc4e4a2e13daeb5b1490cf4db75ad
z53acca726bd5580cdaa68b25053b44c5bc22d9455592c2748390855ccf5a10eac72442b4614b7a
z0d928c1773008c06d3064fa6ecc8036e638419063b0c346c79ca9d260687d202bc0847af3c9236
z2d45da94ff968370005960ec2f8399b56c4f3b541cb88767d6e1ddb69d1b1722cf9e2142be18df
z72ed3e744af4d3ced37e56e67c5e447acc510f9a143955ea60abb3758c95776397412d8dc965c4
zd03948d38b07430d9cd7b69c0b175f6cfa0061738c3a1639819ab24962dbba197a9d8f2d743bfd
ze1a470ca1b48def4e9bc83d6f6b22aec60d84daea9e421174da218cc4e745bc72089fd84fb87b6
z96b20269cd9a174592901f78970d24fab9b657437dc99a24b062f3abffef7ec816a96a44f83c2f
zc5dd2d88929b1906d133f903850e66129bbd7f084b83711ef7c967c6f68cac6964f03fc1a9f982
zf0691b0ed547c000cbce7050a06f971628b71abe56089d41cb128af38291648275f11f8009a537
z525a715f2f9a4cf5bdfa8d91ba0f4acad467cfe62f768e81385957867cf12c64dda234c42188f6
zdd6e07d24df3e54e25655c16f2ff7488b644b0a6266346f31acc586f6383f384859e552fcb467b
zf53aeadbe77d2f1b37efbf8e7521135cd8d42256d0aa4eb47fc147640bdfa386c4684fe979d3e4
z13fa3d033a3efcb6e169121734871b2364897e5c1b57b1f1bcdc918ddcc7e051f1f752f2811c4a
zcd5ed3ba46c746174185b29490547a22155cd40289cf6dcc4949acd6e896185b8e2fae9d11cd3d
zb4001016ceeb3654b6ea414596491e1f3b56f22e658e277af78586bab822334ec988c8e854e138
z94cfe382342bc39ed3e170fa6c72ddb9363bac3c032972d3834d5d314a19e92918a47ea38c0732
zfd6df1d74eee39cc36117d38c404d83f3a4ca8bfdec289b1e6da3f9c61ab5115f352136705573d
z82b8b37e34ee5a061894e333fffa45b1159c2d58b7d3a9a831235db0b20897c91f17baf6b38de2
zf7f61a5a37101852f8561148f947cea3aea994bec5a503ba77ba1fc74ec5db433945adee254b45
z9ae2f6c0525ebd6703186619ff1f30eff2c834592eb2f8f23a36fac13201c2632c1bbafbfaf420
z9e885b8fbe557c6f1e59b4358deb23c5983652a2d4f4263904b5e7075ef88847e6674069ceebbb
zbfaa5959270ad3cdbe3899aef6342825d1b35fcc6263228435d594d63d0a03fa397987fe7e1dfe
zf796c292630b7c91a96201ebfdc78346af25845b6c32dd32a15e52070d0a4a66918b6bc87de59d
z13311fa7cdbe1186b6ec3cb17a6836b1616f7541a0bef84f9449cade806e9132dc00475e67c263
z95c2c6ae49da1eeff6966cbae74df3b6eb1d838dc5ebc3653066cc87f6c9757dca439367ba68f5
z2a6ee7f846d07bcb62e4bc0185cc46047fe52035f8ac4914e9d9cce6e1681803a9b7883c522c58
z77d1e2de32d4da079e0207c96a5daf4d62d28a2efbc33e540870d21c82e46c71cf5da307297664
z4aaefd65268729b1cd630d622da73ca8c1a4ac7524b0812a7d69d7b6bb26346ab751a4370393c2
zbe8f8dd52f0d46c6326a5ae662f22b7c767f26d882c1dd8cbd589bb20923aca441b02beae139ef
z798f4fef828c1a0b1d377ed1b2fb26b5d1f1ecce4706697932e90c377b43e7212332048a6cfc29
z1aff441396f279136e9004b8a979ff04028292ed918ea8409256e16a25d626ba4d7b9e17ec625c
z463f58ee774b0860d18567bca1cac9afca973b1a87d036ceafdb4078a938861dc461a0c1a96194
z35652d26fd9cfc51073c4bab96ea778ee156432b36554e166b763b2b9a6eb3e7e45f30500abc08
z4131ebd9499c558b0108bdcc4bbc87500657d6bacbfa575eac01891fbdef1898ab4d1aa57a2bec
z327c40349ac96769a71c8f890109f0aad44bc0e7230401dd075166cb3501e3403faa35b8823245
z3723b73190ec82e3491b3d0d41314259b431a48bb3161d1186c2483666e222f8e82f414dd92249
zcaa558dbebff2d860932e848c9867291403fc0e929386c871e1a56abb8fe3627955ef19eed2cfa
z229021652ff9f95d0bd07b4576c0ff2e033b0ff393b706a291f87e10fc178e3b1d173e3d3a9920
z985ef40eb4faefab12b81cc56e2bfe45d54fc420587b64cdb763f9f6f80d686510227a7d5ae711
z1b578f2f5a03815760b56e51af62ce42251d8272d9384cea9546534edb91c6834156e8648ef05a
z3a2546bbf62d22d13cf2a712bb482d697e7b406bf95c87073a01077caba1b24b047cf4be6b1ce0
z3b6a6696112f1d4ed47531d9bbff784511bc07eabde1a57f6c7be85bc24bffdc21f79f58a20c4c
zdff210178c6043ba8188211a226d9de370c87e77e0e71b22924de47c780459361c721ea1729832
z64943986f1f44803e08fa77eb565f53413ce858446ae818cf5c5f8c608530c2f0200bec53a4cb1
zdb4d4025ec6b811f3bde78050019e65597e09116530604ce41d3ce83b5b4c70db7ff6418ee44b5
z4826a2b11d71dabbeb9c6b0aa66e25066f377aa473736aa2460acf336e8595bc65304f949ac052
z16e9ce140433858e516d36debd72dcb979bc860a83fec88003839018923dae3399d5c38e9bedea
z63e8857df5fe7740000d00a2db33bb9cc2007db482070f9d6c48dd0c61b34bcc1829d835959831
z42d044c8e6a1ee9adf241f9c39f90579b524d7472b6c9b8cf5b961137b242579c7b16c1c6a6495
z24277a31fd4bcd0189d1329295bc7ff065d0e6a05a580185b667c0874964e0fa7eb58bb1d3c03a
z44eed367c4a1f371f8b13f8755533822d6f86bb731ec570b45bf3ef2749e5ff951d014a7f4d9b9
zd9f854535e610f3d2d4e66548f65cbf57868b905c8ba07cbd9d8491c899d91fd2a4d207f703ee3
zf94000a81c8629801296dec2ef3f6f249042b83d5d32b3006799fe0774b20122989b36da44518a
z83849c13ba8eefc8a7435c85c3750b7895d258ec42f58f2009960666723e90bb5dae9fd48a1204
z4351fe7600b26cdc40ae60c3cfab94d21571c37a384e6af002690ea62e445686433f1b19543331
z5c958c040c1ff0e1e7bd7bae9fbb2b88627811834c96ad7acdfa2baa55a40f94213d7b7821877c
z744420a408353e5b2c72ae9a36b97b66522728f8e0320c819c6a0db065ddee0c8389e3e36d9c2f
z4c6152c0c24f60c64c32a56c3b8e89caa01022503bdac16aecaa15fb0614e0fdf0e96ae67e4e06
z12274bea19457ae949b462a28d4c882b5a5e5c1490ba0aa770a0bbc51934ed73ccb845547af9ce
z86a793bbea7605ca97033ea17e10d29068f706902032ea3d1bca3879cbf65c9cda578630fecf2f
zf43fbebe98a6cf809415372bbb4c5d7240de0fcbaf8d0083d7e937c9b44d0543c367eb3e503821
z6a07d07a0e02145ebad06b93080d717f93534d60b49f65af25757ca83afc6647ba9149fa0017cc
z0ef48214e3e28913597d2e9205df81beec46a4c03a16f87028f559d16f21fbde669b461dc194ae
z42064251567e3b0ea932e5c117977dcbd098aaf56cba7ce839f762ab83deb74b91935c392dcdcb
zf9e2ea71c699d5ea5f0b9d28b62a75f1f5d8efa93edb0cdd3e612740a8741e97daaf658ee2bfe9
z25d123117041f1e11f8750853c1f111d2bd33a8cc4862f6122861c168748eb098b2fbaf2ce0c32
z9635f96eb1691587a32908196087ce67fdc2236dc7bf985e189b1211122cc21b52ccb53a8aa2be
z69421cf493373b3ca9a3bd373db304b439b746f11c7afb68b15a1f475909a1dbd24106893f9146
z6756ea1b63ff841188ca0624327bc7ebd6562f1b2c2b7028788151babb8e2a77748b4f7cb594be
zd1e9f87c307c4b43fda73511241571b7163c1e9e6dc213ac0f3d633e81a8a432f18343a4f2d6e0
z1027809ad881dd10112f30aeedadf883740d1a3388774f30306ffbf73c1d9ceaf37b70041cc9b9
ze42d24bdb5914716683d8694db3509defd39725b9cf908105f05b5ce301a01c54199522bb2f28d
z17c8569cf23cad91857305baeaa8fb3d4776feda9a008793d82a205e81b231c9c48ce2f2a648ff
zd9cc003df0809850a41596a543261ed0781d168b52b51dbcbe0cad96da4c6a0ae59524a0138a85
ze6d1162748950ff4b1cc434012a07fec5036033d7234bda56e7842d7aa5e05c2b82ad0e75be9b5
z867a0f2c53efd8ad5458673d01859a744f61dcef0856fa53854b0e80e416c359652f0006c14343
z605e2ea793c88c48994cc94732f3a8cf5301eca6c30b9e3a522d197f58336e0f31a8b1092c6edf
z97978a043ab02ab2723b4f3d0d35f92f1740a127e56aa4e063b0c3709105e8adc17ce7ae6fb9bc
zd20073cd680acc0422e7c5b8c41ab1739c27da9a352e4f70581afb5afc78de481e26087f7dfccf
zd7152ad2f1695cf043ac68e0f51ebacd00407d31e0343ec8e89a3be261427107b05475166bea13
zbf11705fbc7a1d0af12f0d96fa8cb827024199349508395ace0b8064c37d9eef15d99f221098bd
z84b7f79b85f4384a9e4317c31a3665b352f5fd397ac1a5792ae23170a2aff68e2854fb8e468748
z5999028de4b6b98d9aba773f42dfd504d58a7d2ca42ce9fa3957ffab63e8649657af15b369ce9a
z664806dc445d012486a168c11769524ebb9eeeceddcb82ca72f043a92a95ab61fdbff522ec8811
z2d73010335a0919bd4b9c1fde981021146d14c9d061a4e6ea9692f65cebf6d11e5945ed1ac4770
z070b69a507d69cd90335fafc000767a2b4d6095ab4c76211f2b9ab0c57cba98f37525d6d4a77f7
z879f0822623680d351ed3da3c77e1053f24b83ed8546b1ddc68885094c68cb5ab1cab67ea5a9c4
zf0cfe5c22f65faa21090737072388c81122c1d213ec97e227be36e4f6237e7d86a0aba8c19ad4e
z2cd45bf6c3da45cc06314c693be572355a190f552650dc34084837a777e61d2254c5cc626031cb
z86007b2aa9f14227d3a825b260d214aa7337c806e648a7f853bd3bd3896e46af78fa46d0466cf5
zed3fc8ccb0d179ca2891b862d0e5ad293146542c2003575a3ac78a8412e94180060e45fdd35c4f
z26b2b163f13dd77f40de4de884c3e96c6eb16cb3890b2c9e97ee12d94363f14cf6d2f3be4c1521
z9d44d50138186b183b77e93631cb1358eafab94cd346859560e106f1474de7ae7832963694d1f9
za8c6d2179f9a0eb3b39551ec017c36a87dd7f2186a15b1a620adfe12145f9fc35b2086d8c778c0
z70c67f51fbd4944d397ebe31af8adaf829c8bee7b7ff8d28d321977eb4cb9f22886cb2bed31eaa
z3395b5d9cf8fca20660ae2815478b754d9598ae57973b66ce929dc7b358b69c4eaebb540cf8c1d
zeb80e3a90af400cb190789c3ca59262eeacade69f8768252ac0063eeb23a0a150e25516f5fc4eb
zd7b5e08211a7ec51d86847ed96044162ad5fcdb800997d56a60559e195a5a9f0e2311e0bef387d
z9fff6306a89b62eed773a3053a90536b00fbfb5e913ccb30760d7dc61320b9686a3e325b2b28e0
z3dbbbf1b738c84db101443441d29339fc9e77b811f3a143e0f78fa9e390b317221cbfa682ce8e9
zd0e0ce944dfc1d8083d2a1bd99963f6484ea7c6ffd6435f1c98e6e979e40a39b6b2d8bb84bb2c1
z1d8b3db4bb1b82bbab774a97c026c1cfd839985622e62ae2283216ffe6d4f265f1b0de3f9a1904
z630465c6e0335940e44422dfbaef065b5ae34b73e2eddeefdba67508776b5c5638b34a2c31f01f
zd1eef221419c581d394279e0abb7f8429a245d222851f33fc0393db3b07b40ab72a63034e81be6
zd055ac4e60f5e4737f4ca20a741f115eb1030cd4eecf59669a989a76abc1608f7c8e3192bb088c
z80b3efb2a1a016275a875d1e706d7cf2f64d8befb3f7bd52543a6edbf467bde4548e49aa9d9c59
zad363e2cf8ed34a498b30f3bc53ef44d9f6eca5caf63ed7694e1cd34eace1a340eb8dad59cf4df
zc5587df6ca2eec84123f58292441ad5ccf8e019f4277e0480d0a0e317328ae3fe365f65fa650c8
z058e227fc5d91b5e8371d9f4cb7ecbc7f155fab378d8488e1d7c6754021869cbacef9ba67045bb
z86a4f129864a77207d89ac1f7d642b21d546c4cf72ee0d0357027c43082218f4a0f79ac9b9379d
z5b2b2f62161794a12038b65162e16f34090f720e4ff65b1bafb9181e7b630523b4ecbab0be333d
zf4dd189a296b8aae90c5dab3e9378419670b18a552d5dc0c9996e3fd2b86b5cfcd1acda5f162a3
z5eec1d18f4f6a8f7d3fe2bd6196cf796844ea7aef78188a50a8e99acea183b847c965638bb00c7
z6e8a6c9f7c23ae2f94ff954333a6545ba5464809fb1743d2074eb99ed99bd3f7c36ff3dc5e9470
z880c36c958478787245a85ae828ce0fa8c1d8d3c8e5d606555938d69c259469e872a6a712985aa
z2994c877b0afa0bea03e6774abe69015b7a4b4bbeed8f0987571317a708c3a9ae357be0f600ab9
zc0e92d2260687e35886a69e948203c2cb5c4a408608633ed57be52fdf7167d6f5a47e24fcbb7fc
ze52267029e5039056f66b9c347f7d3fca21c7152d0d16519ee75698cffa090473de32d12043b37
z845c01bdcb3092396ad9e07ad428e14a4bce420732bb32263bcccc7a340261d27bc830f71b1225
z88f5be8c586d0fe4fd079a59463a61e1b28e04d5281c360fdc9b5c35e77cbda7ed5a5fefac856e
z849cdd2968932d024d53a5f2bc2618ff01c9598e07dd318442978f5ce6234b3eecbf110ae66dcb
z7d83961436f08408032d10b3d8fa471e48af25ef4b771188ea252efa2953c2efefdba719da185a
z664c421bd2b57d0ec50218caa0f181d7dbe545f8e596605585162b450f478388eb9774b3d3abc1
z212eedb338163a70322e47c90b58ae1f9c16aa97021219ebc5dd6f6b63186db86bd35e5a33548d
z95a122538eecfa698f1e18246fefadad2d10007df6e5c9284bf1bc33dbaafe3d50ed6843ac4486
z0594c249b93500d904847f7184fe7aa2ae0357904869b48c4ab2d94fd3bd22a262d8f32439bc45
z7a75db61f72c0b420b74f190c47d5db8924daeb04d01133ab25404b88726182abe736b26fdc765
z827725525a413ee63b487e8fb482a07a8d16a6895bbccf0b2e2bf337de90aa3fd1dafb10bc3014
z9545453a3a535614d554cd7f814c5b3dbca39e2acb57649ec579c1c4d37e663ff8f3f187aeb724
zb1400b7ae9a4eee852dfaf96c64d6c76dbf29a617811ebd8d66091769591b45f3e6b2aa38f6d56
zd287a412a558946c1c8bbe539e4b4729165f3b429fe5536e2d7983e40f1151e4c967d77f58394c
z9449ad8c655cc913ffb203355fe60c33279d953e1bf29c0e6866e84acd29d3c00230a1dc167a6f
zb32c914d91835c851bf2705aa79773c9a2b4bdba18f5ccc4c0a54e10322645e06896bba7966317
z7e7bf1b837a4874396020641cedd0036a5be148edb992e38d01a4ecbf32b1603b4f0fab12d546f
z3bc872a982b86d6420df13dfee38fe77a13fc3136473645f708c9d4bbef0982417d460c016ad0b
z40ba3f6047d5de42d54edf6986128c574f09de9cbcc44bc077c175fddf64591e30d06128eb05a3
z7d47919bd05e4d0fb3da47142e0a459e3e52e3d3a37e139b53b02befbb1a8e1565317f691caae1
z3173cafa95278fe69e42f4cec1852d09f569b9bc8175c4b32e942ef7ec213ba76f656df54a612d
z1d4b6f74a39b5c48ab71e2a0d6124d5e48079b8b60d2478467873be02f9932d2bb6b8e4e9d43ed
zee6bad106d36d37b2e0e24a401e9e2db2e5ca61331225583c882d7d14559ec89e687950c9d3ebf
zb38d7f7de121b8604c9905ec089e01f3d70cacd77b92c836345c4c85f95d5bd0f4d91d5c570b88
za37f751d8cbba2d4f50cccac7ec99f3a4b5416d3a099aa18132c025cf019879fb6f67a5d0b5977
ze2121f52833e1715759fd94744c89274ef29a4dda613c969d3cec4ca049e38315d947f21341a41
z83e7dfd16c8d6ae05e22bd33655a55124ab7e9ae50bbff7f72fa2fffa0c29fca8fefc295d09374
zf1f07002a31d4c0056404c54849608a70f559318c62d4958348e821eeb44f8b6a151a7f0fa6696
z899f70e413a87c9b99ac4653810ef6416297a945f1b8d034c60e927313ceb453f13ee6b28e38e6
zaa092dc56c125e1a04be13501f3f3a206c22858b6239683904c6be93287d7339dbc5f44e2eb378
zfe4c95eeae35acaeab415f2185a543f9535a7630467c01e535cd29f72163ef8dac06c16151680f
ze183515668e913c6ce66dcfb9140fb77c6c0e333c5a9d86617c0f72c1ecf7014d41e2732c60cd7
z6baa11a2df862d99a90dd4abd6484f7a36cd4b9dcb8f280ab20cbdba8b4feb4ad8e98800e427cb
z07e84bfa99e6ff72afe236f1daa8cdf4ae7289afe216a6dc5571d47d39e4ee76e3d17a46bb161f
z782ea8042e8d5a651d3754fca100df847ad39d508f54d51c74416ac46bb6da219e7d4676637a80
z6d9ad5b7deef317e144b2bd10d1bc00afc5b1b160fc10e3382f7708e584e6bee9648ccc97c0932
zd3378490c22e440fc3241e7034d979fe2674f384367bc53f829f032474a87f774ff69e23237fc4
z260519de28fd03173882e0b7fc786c4a8cf2539aab7d0b27f249c72c64a67e09f854a06cb0605b
z4fcdd7d107a162537493459a31156dcb11b7b882a4ef0287f9f857101c9c64d6cb1bcd17fe5cd1
z2da25e5dcab0d2bc4e5151aa9e9e37d71b85d66f4e442f26643361eba6e12c371db34b76006766
z45ec72884d8634d512f16bbe4c1459ba68701ddf42201e4c167ace6bde6f82a4c21669753dd63f
zd9b8798a265681c53c4d22e047f619fbfb218a6614b48b1694b2158b9e2d41ff19f2b41877c43e
z2389bf9af45aaf395da3664658a778d5c5df4aabfef518a1a9afcc69859ad3cc7b73c0265ee240
z5a156c6e82ea2723a3a669dea8694019102e271d65af199ff47594edf5e252e43465ccdc8f798b
z7320167466632774b96c2aea560c2e65b90fddefa3544c088971f09b2846f6b59daacb2d5fc59c
z71da9980ee216b8b9894b201e99b5f1e88162d555b85239ff7eef3662053b27e490da5f86e901b
zedc2d9653971a1f2ca90df75301e39f3a780e2c826fa05a658051973301d84419f9afac84970a9
zde0fd9f6f594b6bbfa2adaaade6cb58cde50329705e63fc6e6cd8e4d664eab3ef367b157f30722
zfd45590e6fdb24733ea90c671e6fb349b7eb91affa938d31102f64f58a475626696d9cee7d94e5
z74dbafcc669f109f877a66fb4da8172c589607852fc3224c5b0862088a3f17fa4e37d0bd851e83
z71caf98c933fead27d0477d562a51b1013ba9a090740ea121583f01ad9dfc658e7ba471c2d7df0
zcb9084f9e33da7f9bd3fada9458c68cf333b44f32fb3301defe1fac5f74afbd8dfeeb6c4683827
zbb39eb058627cfce7bc0e7a68e38eefbcd5532fe8dbd0b5ae0df1d8e337bcdfc4cfaec0da3566b
z294773c79492cb92d87e35b918d6e33431c5656346f6dac34ea699eb5a027941bda5ffb6705d90
zd55d2ffa16b1ba3a4c6733914b218819659553fe91a768e7924934cf34e8356489e450cdf9ecfa
za5163adecda2b2c15ffc2b9898435012a828392b52ba25b1b51bf3db7513f517ff2621e14a7499
zb23e1dcf5ad0769d03f68560b0b149a1581b8d053302e2c3b7c5d6ab6b275cc9a35794fb84b295
z0886d42d958a091e60290c809d2bc4db234cce9ffa2516bf10d3a39c163b9ed2e61ff6d6ab3af6
za3dc729a305dd615cf20361d6827654b722bc3d7572f41e38e09adb8934a24acc51f944e8e8a1a
zcf6880ac16d995e9d6c1d7de81994615b93510d76e0791ef4cf59e2d9a68ee74381a626e4a5757
z6a51371c14674cbfaf0395cc43dd6deefac54f3454777a6ff8878533dd9fe01edf5fdfa6a74a38
z3cc0c83ddc8f7c6bad4bb857a88eec3ced3719c1f2c70a703368f8232f7a6d6a7a04e40feb70fc
ze4f56c46eab994b866b7ec71ff39e4bfd44155cec1fcd5e22400269dc8ecfdbd8fed4bdc2f71f5
zba1bcbc79163c8f2e5fccf4b3666c5d8265a29ca1601c3d68a1539c3fc9969b4ff2e02a8b98cfb
z406adf074b153256a03af4a7312478320b2f12449e8aa4ab6e6e5afbebbed159ea84ee628d22a9
z3c9bafdb81cdd074b13062e1a839e21b9ce602d3df168dcb4057e80108c91725d07c4c395f3dc2
zd3bbbd24cab24aec326bca1ad53ad36df60d38cf67fe02c75c60a4c4b83a133e65d215be8d6745
z972c77a2bffa38c159d84f0ad9fa40a5f3a1786b7d2dd3a380a9db07076f45b19c67aa023e6a5e
z9938e06ffe5d215f7001007d98bbb43f159604cf18b4cfb34c10712f7187c1b76411b925bf5497
zbcfe0f6b04f3156c2ff10d0c472c236f51bd712f4d081588494ce46dcdacbd700cd15ee5f89900
z39bb0981aee33a8a566798ea8ef29dc33ad1222060a7d83a7f0f4b35fbaf7673c06a06f8bfc05c
z906af63668582d4b5ccf6a4523afee70a1609d8f94b76fd5fc820649f112f969615cdd9ba4d640
z2bbe02302d7fe10d16f8eebe0f0fc7a9edec71a873d27c33b67b9dc50849ac45dddec554ad172c
z226bf00cc9f297b64b29edd4f9654b2b2c1548ea8256b04eaaff90c627f4c7ed97a82d10aaa810
z6fbe97a9819263b01abb76d718e1b1e531ec03c6dbdce413645dc056f7ba3f2aebeb4125f779b8
z01fcc0ddfcbaeda0fb7e25e8b24f2c6106888c8bfdb465936656b5edbc97793846746807a09d56
za866fa260547e26849e1367b3d2f3d7debef1b1f062776c8474fab2c263ebc926b3a41bf1f4000
z4d20229bf554f6e827ac0ec3731a11bd65180e33aa7254ce2556adc85595a3e1280c505dbab9ba
zba45d0056570254528b1bf22b1a8f94fedab43b0b87c08fcd68d8a5e77d0e0b2b42f3c94d35d0e
za9b88e751b7acc5bf7407dc1821b654b82ba8faae1ed5cfa4d784b8f71503ee1fd5c7e5ffc1ae3
za1d0ceb08bb925118f05db3433b8c28a56167bfd80909181b9e5cd3bbf5597cac20b86cf717e17
z234df58c088abf74b0f8eacb807a9f647c31f482150e539bd9473c94587f4d323a027ac2fd0b86
z8035296ffb5c74e70f2b36eccbdef7f208f58022f28a97837a669a74504da0ebd3cb02262ef76d
zc9c26fe5baadbf5c149e28899ca55c0e3a172b0aef2d156f94dac1413bb38d2fa94016ddd62fbf
z9287ab69f4642ce91dedbf81476fc096cbf5708de669959d844120624556d81ac820ca255bb2f8
zbb4f437e0f4024c5b6f0c1191328031be45b3f699cfc99bd84a1d97ee321732d78bdbe3ad1515c
z5c46f03e7982dd83a0010380f1c2c1c058e03fcb9d655184ca59eedd2a240a3298057aa6ad34c8
zf29e289a69adc1a7c5b6ec08c4181465e352de419b66187577d87c9814f58e08d493b6e486d8e2
z7b0a747bfe1a5672f2089e5d0e25f950c8a8714cf6ff671ab0a7303709a7bdd04b652b5a1db98f
z43ff4653630c30307879a3618b8e4b671fc56a26e225d330cac04edcb404e746c0b8469a704ba1
z301c0fe82e9fe4be299e5cb0b5a871b65edf7768a8a8f8bd54fcfb89010d5c9223dc3577bc71be
zf9bdc5d3ecf6b92201c45057c86f3c1cf557314fcadb2861e5986ae5de05a27b4a66b716d4873f
z38557a7df6d289b8c565ebb833d5da04bc4ceafff3661325cddfbc6765096407658af8717b78c6
zacf3c1ad521bce1c46065624c12fddf10ec967043b41c708bde43105935b71aad9066f2029a566
za53a37ce990e635e0d96d81f468dafd5f3f23b2144de5de98746f775a31c56f3626329047a90f8
z97ef3bfd809c310a0a41ab790af5d23f171de07d4aede62dbb24ac9a987be577e92d01dfdee5e9
zfde2851b6f919eb23e62c33792a4d8c22689e39d8fadb7a47f350c49d1e567187b5b9bf8a050bd
zeede5054113f57ef527e31a5fa323928088fb59cba4f8648a243b10a18ddf2eeda48392721d9e0
zca3f5cb6834c537d197d0f1940caf4aa676d1d5bb84be101a2963c647db73264608960219cc52d
z533847aa0a2d78400cd4dbf47eb776b6f003142176560435fd80a61f6b9928b27966e075201a7d
zcdaf9edcdfa163252247cb12867a64dce816e1b325f8d9511ac76178918dca3cf64d97e0fac3c4
z9bee4cd2024f3462d8c98d5ecc1ac53173fc663ab5d6c83f7f444bd0b5ca6db7ec23a808a7709c
z7f742175d2ca610526455edf16bf54ed8a0b1255c8554fc856f8e2df2bcddd892939a881351d2c
z62d1f03a1d03af2ee7d83eb5f1503043071382e8c5c579bf4379c3083a27da3ec49f3b94aa4562
za6b8b6379b31c79b2aac0d308d7c54821f811ccaf4dd252c76327677d2a4ecbd460890587d1c68
z5ef8e374eb0a9c4cd3245722188250dfbb5bba054110a490fe6b3bfa0e8d8daffb0a9b348ebb90
z57ad7f34caedbdcd5e93ba420c6bfb276ea3663b4fa359167a773d910e33df5892d54cc56d634d
zd1d88dc939fbacddb7d22a1d01f316483a3dee41132ddc9d9fa807266e22ffec3e416fea64ebd9
z205c10d7a8612a55e728d6cb3e069f0d80d278addf7457fc65bb2f0fe86be16c1befc4b81ff215
z5a8861e2d2987bb2ab369e34f62106fbdc92d0f69f13e4dffa702e24118c5b6c70886902533ab2
z8d6e6b210e5b9202cd4d7e5d09ec3e7afd0b147c8c1a935fec0b65e6b4df7e831e13ca1a4e1737
z5ef38cec29123fe2b7f45c3cdb85732c950366d01c2db35002ff8a3a1fa742b34b1fda02dfffe6
z576d881bcc08f63309c9c90b8f40bed8e645b10946526c95b9d0e76975a47bf64ad8944e70a076
z56d12d409ca5158fed4c4346ff327de1cd322fd9e79c1a9d6de43adbf2bdeffc738ff84b58523c
zb545d7fef919f67b79f8d007d553a587e0c592667d698f78e95ae0359081c726bfa03572fea2b9
zee864ab2cb943c0e8d2277432f21d4b4c1b4c11a936c099016383adcd553ac25fa781ad37759db
zf2de4e5bb35aa07f6955e9e1a97b6e6f974b9f3f9da41e1b949dfdb52fe9f2f8246fbe811513d6
zb5886133bbd2c507b017f871ea4be92a395b18b8a3957455009e5b6489edde940108185e92a86e
z6ff57ffd0f5135a1552d4b5a961be3de0f77f1c6d1c6994038b113fa4c35de7d539734abb05b8e
z0bd57fe9eae1d63a07127c23fa6c595dd0c4e1c7e2a6006f0868965c008f7549d83e44aa27e404
zee55f4a211c2a0c1ff01ce7c7511ca777c4a03519d9eedbf5da45cd7110dc4995122abc6be6244
zade5fb3684e8c8da80565eedfac956c35402f225dee7900b9d60d7e714efa0fa8307a94d931537
za480b9eb8f930b89e45bd71b9868add0b03a014ec3655c10e2e41d018c19a6938ebdf70c49ade9
zb0db893847402bb86503ed708e481d2c3c35040ac6e84ee0e099b61d5b32d3b94e3c6290f6cb94
z2a194f33bed81f29717f8f0bdaf32a664fb5dd6a18e0e0b32a9907af9ef62087105c707485aaa6
z5a472156f95194872e8fd44368a9c27536bc51115906f5348bc860c1466b2f7f8502e54989934a
z4903221e127579c9eb669287810669911e9cb8ab285b5c92f68526f5cb3016bd2785e1e10c7161
zd01b7c8a0c976afb87807122c5259ad91178fff0c0396c94b4fb97be41ad221c13d09d45b48603
zc9224705623674018f3ea1bb66b91cd93a1e7dbc14b2d395eec0102743ca9db4d6a363c93e75ff
z97469395e94b6b472b6570c28abebf487e6d01dbdda7a547d8113fe53317ff82095af52c89d746
z621fe6a2e93cdc1d1999a599de279fc6427d4b348847db8d89ee651a9a7332db8ff8bda0cc0c39
z00bc57d769d3f782900437639945192eaafd1a5d3a098ccc14305c840d3952c9a9047df0f226f8
z4e213da58561072399c5c1567dc8b7382e93c2bc5624e922f70dc87ffc8fd3e72ea77d5dc3de83
za906bb5e905db7e498eb56d17257ffce4a5be1be7a97a642809a2ac729641326097896c0368913
z461c5cb16cafddef044af57737a500eb623a71b1382e6eed672d4c458284af0b33518962c7faa9
z893eff973c1cb742faf1d8175709e427f44b712a078ef49dced02b18ba9923b42536fb625bb003
zc00217b1d4380e30503c42d600b7384ee7d1f5f96bf667f5381962541a7d2d85c3aa879749f80b
z54f5a717a805b965fc0d5deef44e708ccb8bdf76b03ed82eb088a52207b744f3b6862048f91abd
z64a6b3247d9a4038378031a48a93a48bcf7a030b6a7b8b122167267612f0e4578995a741477f82
z3e28958c4be064d1757cc45eb1a066b3b31a5d63629ebd0b0047fd77affb99bc5b5255941edce3
zd26a8ded69dc780e533ed8a72a155e51bd1a76ad2e039194cf86f7b3cdeb1416b09cf3c5bb9920
z5459aed84010896e6ffb1b4e5e3ab4877d5063fc0ab29abfe5dcaa067f6615802171ebda023a3e
zc2c448322ea80b50a3b42ec7720e109d6f4b03fa6bfa280e65804c74b1204de2a2d11555de7d21
z3ba4b50867a7a1871b122661b25d42933cb9c70ba666682340e29333b681e06fc574e81c9a7ad8
z11618a267718a15725669dbed781f82ba1a4f8c68fce365f2812b2d695bd946b42544d90be4c64
ze29c923e8f9e5abc0edb3f9e9bfcce2646972284a2be411e828883f915585acb70099729b50a11
z31b5be30fb0bce958e17c1a556f0ad7df1be51dd233382e227093859b4c3ebe2701aa52555eede
zbf2c744316d3f89cfda28f549a8112e04ec208d4b4cc4f48e6a87631917d24a66772929bdafb8e
z9c91aafe09362dfd4a5920f5be5103b044b06cc832f9a2979621d3639b5972f31c3b87a9121e95
z7635afbee81142c5a159d5df75c4dc52399332c19160b9ffa1fd94ae3257065158d9762d1eb66a
zfd8a885c06a40d4c727916eec7262cf4278ad19857ee64f1c2537c285765cfc893b85fb572b40f
zdfeb7037c04f23184ab959fefe0bddc90cdb4c094d87393fa4cf0f99c8e1bce4bd32ce9cd52d30
z3a1bab9bd611b805cb02c7535b0ca6a075fbac89830a4c12ed9cb19b872f06112810a8e131fbfd
z0afc30b7587aa5ee6f7a228f385441c2dfceb9dd0e7465ca6fd82e3a677f6f73906ba27925756a
z2b3a87b3aa01623c10ea05b4bbfd0b0f5f79fdb22e92f7d05370bc370d3596064a2acb1939576b
z73445a2a304a6f14537ee39875bc68e5685fc17280ea4d9b5ee4f9aee164ac0e8aea92852c11d4
z2ac5422489470d8cb272d3600753f159d8b04b2674bbdf36f8ca63df3cba345a4f6a30b28f435a
z9ee23eb832a47808cb9ee020cb190f3e73d0aeb7ff91feb04ec916b751823bb4448eeaf6d34757
z08eaf3c6df0a2be60d24c3e0233c0630f1d219085d1ddc42d061520a5a08246bd541a353c41be5
zafe76c077145c98f978a64b50693ae6493e09dee76c6eba23e792c59b62081c5c5072f658a60e1
z7cd28c057422a739f026eaa3159f4732afa06f14a8b829a7aa2291a67246f61be72094902c4a25
zb89a496f7c634a4a70a1d919e790b859fae53c2b575d094b425011ee5c6e5ec4c172478c4ff405
z83d0ed319a986aa6b63eccd0d235f7e7fa3ae1ae2f1a4045b33228db4ecdbfd97cdeef0337fc3f
z1d28828f60917aacc869388585dd86d633405af1ac4dacd57ce15c801282796e2f24ed21429d85
z1cd4a8c68f7754cfd9089e3943846fd5a42d854e5d80c11eecff830a2208c47c8afc72ea0dc6db
zebd664c813d6e4e8272d670f16df9d59113ad22c3fa9b140c816749aaf5e08e802c1a7cd54d620
zbce828f7ab2d413cb698efb12956ef032fa6a0cba64dce90031a79c296ee5dcde7af23c89cf91f
z188d2579c99aecf5a3f1980a3be1837494f001e04edeb7109794f78e379267c7ec7bc8d826b5a1
z6e46b07d360367a94734f20fd05560b89b6962ac71e9bc9fe35b8affe8c40c99c907e327ece06e
z5cddfe5a8b3ff3d72a24e5286742c75eefcfcf6f7b41552692a61da051bd81d90bf3d42deebeb6
z3111fcfa14cafffb8ad2b6d63b1e28ac5c086b445c9c05a7da9dbfbc9e82e1755f3fc4c0abebf3
z676f52f7e7eef51b8b8526373ec5a163b56cc4585cec024235824bea83913a5fb09715a7a7016d
z65196373e8b2dc0ba1186d7cf2ea4c716029c58c01c0074f886e7e8d30385ed229bee4f72ef3a0
z559529c1bcd39d174cbe987ad094a210a1f91b9cd4460cf1b6cb59d388a45d56767dc0a9d8102c
z9fd1f3fdc17472d9e9fbded1a739bf16889aebdd45294ac72272c0a60640e39136122383abfb12
zf0501852c8707af0ad4db25cbb9a34312fcfb601ebe8a00c49019cdbbbd8f5f661314945f2af32
z597e748dffd1f22d35ca0646511ba5cc7ccf732571a3027bee31ce0ff98b56d9982136a7d43741
za6381bacf41ee18b8e02acec3f54b5cd38a43ba4bf545bbd9b3c57ca5deb85bbab30add4b83d71
z596f5c16d5a3df8962be17035834ae5684ea6976c967b899b59ac717220c58c9b5a2ca1e1b4bf7
z66dd7f9754d494490250d19f09564158ae5990d9d4521a82b76235959da1138f6f76317b143e3c
z92c78e64c34cda119f0ac75f0ae9f0f3f7ec2055d0740c13101bad691c79754c1a1694f728f42e
zc15901a5242d5c354a2bb6d27d06eeea55c375f2c4a0e3e449f87b3b891b95c985f7cadbf96130
zfd2248777ed56c98b39ae95f2fe2b5b3329a88e3e573572a9dd59862859b0c241756e0845b193a
z663d84aaa72b82639cccd493e7c2f14796389d45c93499cd8733901882ae4f05ed2297c2f14709
z11334018eadf550ab47dec15df027d65e3405284d4d4be2724f9a04872cfaf99965a8d4b967cd0
zf6eaac7aec3e73567036dfc6e1f93be73fd6b03a13e9ce10aa1b8fb8ffcf3523f95840a6a4a4ef
ze52312d3e088124f1955ad5d10634d33f0cfbb1f49c78957732054d2301fabe406bae381f4c02c
z42a16cc55e56ba03e4af0cd7c0cf9c19cc5da1d3810eb1b14cb7dda1923a288eb9150ace6189ce
ze0c7f6063c4c1fd5350e1f1aae6a28e257baf6ac0fca63bf994d289c74717e3ea3bc41797e24ee
z86259271aba9f84a7f3b98633e750b58ef87554c32b866dbdb96f853a6cd3d0c0bad7da592df0e
z406c897a28087c4074efaacbfff02c78fb0be415cc745926629bcc87a6484b3235912f622068a4
z026c21ea63a62ac4789a7ac6eab16b22d27727960de5f3a7028c74b85887d80a5b635495660bd9
zf686ddd0fe3656402e0c0dac72444c234ec8548e90ccf392062a2888457c6d148dfce18f9f7ac2
z00b7e1a86d414e24639df025b2eda08c91e180be9848ec6d9cb1dc22c712dd3cd3d31f3d7d8af6
zcc1c8a836c7fc2c8368bb75bcbf9848b13a6b159fa74a263113cd90d3ff0b5f1fe092405513e66
z5c873935eed28320ff3b1e40f8c69b18b2361f84b2482ad5dbca203ef93289ed058c6459c139b0
zdbf7e203afd7a9c1f654e939d57a02b693402b93c933c5691a3d459fc43295226a5f567e7d8c2b
zff7eb35f2a87e5cb75c0a2544a1507cfe1801d349a5004c11d87314d2a453e52e449108478dac8
z56285fc530c8e7dc353de55d15976d05b990b2a775111c9db068336baaa6202c9bbec15ca73dba
z696229f55855d9ee91466b755866f02588684ec9ae3d1edac77127cf67bf70d8e51ae4288dca50
zd0cac2e0521e6a711979100f9645075dbc2e4473957462b51d019dcd86badb3816a4ea83e99596
za79f553b9f4e1f5556d6f54282e0b9b03c58d2e6655709564a7cafc2f41d4e465edfdf4336d39e
z22ed96036c321a2008917fae7c4f94cff192722665d4e526d243a24a4b81b255876492590e0907
z9b00fe5792d9565d37b1b24b20ce12c4087b294ac176f43d10a0735d2be0516a7de888e28a2e7f
zb4e127bbaaf1fb88ce7214c7265940eabb9734e82c744b347fc09c0215ecdad016820248e4a5d8
zdba28055a737064ec3eecf5951b058ae27fa5a8c9f66cb328d3d780c72a179dc5acf13919a5f86
z6825d3a0d782e6245e0d99ff167c7ada44bb29add3cde46d978787d3ecb481839f49eff946f711
zc667d787e1986d44f5f6dedd58c386ff6ffe7d4a1c482d77c5a359ef13f40bf8a8e59d9edef572
z8b946280be9a1f33a4eab2bbe2227f809997b4b3418f4c19f8e8a7d3bd397ba3aef75f3024e377
zc372b17e9a866d16c8ebdce01ddd05fe11344ecc6c8dea983308b43ef681540fb334a617b082d3
z591704718ddd6ef5b68890bae82c8a19f0e4dc06874637ae078dc8c611954f8268909190921409
z9a36c13c8974ae02c1c853b32e1a0fed02d684d50d81a111a2281d7eea8f48d2ac4d199e5b3fba
za792a3be2524cde3d99f66b9721231097ae8439f96976418729c2243faf8a406916f7ae12bf3e4
zd6d91e5af1f2f1a36e52c8570d4f0aed869ad666f279fc4eac443db66ebf8493deade8d70f4d2d
z614ecfa225f6a7c4814553150be87e1c17b0b082b1caadb9688666f7a82109fbc11f1259846a01
z0db7841d6c5789eff2a09a819a8d5329b73cd5c8485de9d9a0f2ae265951feb21153c1929890b8
za0a877e2ab4cf52b82eeb3de4d5f36f5e52e459309461e3421d5d3ad606418e0cb3c9a89b2d4e5
z2a602fa6400d4e44780bdd1ee64d330bcb4c87f4e348f92a9c94a326a2347f055a3dc9eca02695
z14a8f02a9a2033febe2c2a924274ab7b06b06552d3261030c2e92fd8b15d80cf9b27dbf1df7819
zff6fd96c9d79d5e22541487ff08cb675da0aae8b9723843926eff09c1329e6aa9775d3c8a5b45e
z479db4e3f6aba3d3d978b1e5ea4c8b4c8b7ec019d07feb93408c0cb1057e63f61e933d7066b867
z1994a88e9f8688e9ed0e296b136d00539e0da8d1cc48ec940bbf56eea0f2de298b33076d75eb83
ze3404f81e271f8849b281a518ed4befd5d634608fcd813efea5154dbac01d4432773618ea64e4a
zcdaaa09445454eb4246313d3fd10ab7e736f6bea839da737356774c87d80b08a872397528c26b5
zca4ebb3dc6e20fc9d80c9a567083127ce04d474b696cef379d8745573ea67a6263c6072ec5fd22
zc1c9c59bb03cdf212218d503187c0db4fb6d08494b478d15c8092f88ba5ec6b0bc71e60f5f84fc
zb9fcba8d56fe7faaf13a0488f62c96bfd86ef62f7fc456ebe2439b8efb14cc2e178d080996c894
z0d943a9ba19688b099cf67d5d7928c929341db3fd86449908928326b2b9c39790df7eb44c7c6d4
z52eb18ab058884973621d80afb58456d627e07c564e523c7f43fb0f6b1cd555c42e48b43427429
zfec8de794b66b561213b3a59d6cb9238ef2b08bd7a55e56b4a53742b6ca0f795031261b471b583
ze5d5e53d20499ca2530435438719e6f417bb3c0d7082df04bdd01b187d3973cd1bdebda5b282c4
z04b0eed70f4ef2fe4d42a5c3307ec81e2e09960e0e671f92c8af9976bab96ac4b1479e19b9ccb3
ze21e999940c5ecced9d6d718135274e50e3d3d8adb76d91ec5b73ff27144a0b812ca4622439e11
z81b5b6c28ef8ccb6dc47c28ebc16fbefb22f748764e3060c4a1efdf09e9cc05f04c15623e27dad
zbf3b67ce0de5bbe65806be38bf1a24568c8367dcc23b4b0593e283d1f71be41e0d6c3ff6f49bf2
z1e767adff2fab3515b30492707c2996e963790fe067a3fd6635d6ba23030db73db4533cb58c198
z8125dcc944102fe1ed0dc4fe9b32a512091710d087f58f8cf65f4928ac6c90e0fbc98cadc16dff
z81318e00145af4980212166b707f2591d39eb1645507c6a82c99b826079532ab964ee20a9540f4
z3e1121c4f011ce32eb28217534a5bcb46a59996142d37bcaf5e3b8e09f63653f6e1c5b76c71e98
zf0f376177acb44d3357c8eea201a74d834417cde6cc2eaec25f5654afff99f21350c953dc62854
z6503b526c146fafa8ea760cbe1aac9719d81114c8281e289ee27bbed29f7f161fccf1eefbf51b1
z150d6679e1ce2cebbc8aed4c86698153a8082b888aa7cabbf0bab4f7a3d5b60a11199240b801f0
z344cd999167da2a55a24df4703c7c143c6be511f22c61590e13cb6125fcdb261efdb1f520bc42a
zfabfd061b05f79472bccf0a62d1a3e6125e7e5cc8502d8068eb1721e14376da3d1a3cc04ea70ed
z66e6e1c082b51c811db6665b4a98cb333db67e2efc86a6af5e1530a5353ee53cdbdd51054630f6
z709ccd186402cfb40e2eb3143570520f5346a9f04e2f4e0412a5547440c151b414e4b7200c492d
z413091935706341faebbfbe349833c4f1460e51cecd6c5092de5834a8ed5da6d8e49a0975904ff
zdee1517b6e04eacdcdd68eb39f7244a0eae5abc4ffe5810cc77e52121515a76676c76cbe435b0b
z75bd1dace2bb60022a1d19afe019f82ac73196fc22830c9d4aedab4ec4683dcf68bb4ead9535ce
z7a2f5fecbc0d4e929bbbfe59f31d5ec73397502afb31f9ae527315d90da3e27e11a7d101443e5c
z0fd8cedc772e0b9439a33bdb3cf406da32f9f71bc77f376f8c55c2a5818114fc96fd55e0a912eb
zf1ff5d4cefb1338879f2d58fba30f2634f066fdc5a61aee010a11fd8000157016664eb2b7833dd
za3bfc1735717cefa4708b14ad17f21bb2da11ac0bccbdcbebfeb5233c56603ddb1f0773d545554
z0c07d7f28819c280045f4519ddddf5db14138bc7d4d097b0168627e9bb8b1380baf93b98ba4c64
z629f672a13abaa73c8ac3c3f0eb469017fdc14f0e9aaea00fdd364e9c8026e6e69d2fa9730aff3
z75748dc1b35e9b841afc92fa1d27e843c6f280e8301203066e40e47a71742fbf214fff2839cbf2
z0ed2bce03593fe8109b7b69ae20403ef82f95833e41cfd90ebb2285404992d4117ed485aaf1c6f
z364527ed3f33db8339326b5b14f7891d861c6e64a586814f1d931924e8a98d36cd402ce7df48ba
z85cdbc6b8af46d6788580dfdeddc0066d928ffc84a935dcfb92758b6be9f6880533d4c33f7fe43
z8b381b8774c82917442a9ff985d67e613001a3230937a717c036feabd838eb5542d4448154f6d8
zbcf9c3be84e747282644299078959a2d2de098cecca1e837d882951cccc934c27c9011e114f0b3
ze2a5fe46a23e280cacd7a9fa963645f50705092e99049865a301034efffec8bcf65f40fe8b5666
z0c6dce3336fe5743552f90d4731b95c3749b2225c5a1f755cfa00c9974b4916a34e7318d987808
z2c4a6147a8b7682f251bee53428a9602db7c6470d180ddfa6c110bc0a18f0f19d20e4612094bb2
zc8a09fd06813e2ac69cc64c76a2d9b9b660e088bb6f853f5fbfd7c4d9c99c5080e62e6de515944
z30e80a00aa544eee289b973550a7d40c2860cdc1466aabf4fb6b022dabd222312d838dd245a9ca
z506508503b4361be29d372799b2889072c30644fa7adb2558cc7c37ee7c80dfac613ee1d0899d9
z9cc034292606b57251aa2edbad171676cc3f1a40e0dc185bedda19686b014e66cb8aff0a805273
zb26ba567221249a6891b00553968af1fb66d5080e192aacc21c2acfc72f08b3dabf143ee4c6c73
z4d6a31e4ee8b9225368393b8d75cf7980c4d35ffb1b39ccd6ef4f1ba4eb0d68f60fc1c370cd352
z1b46f5100bb20684e834fed9f9f8a8cf876033aaaaaec531141e82d7efeaae58545ee4fd7442a7
zd605418b01633f1bf78c383467a5648e8ce020121b06f608887d3aeed007573b2ef7fc7485674b
z464d9c40ec539632db97bd9a5877abb245093ab02a37dda5e8dba25ee299b313a731b6d354f1e6
zccff979a041672cbe96e41ddb468dab067533c5420b5c5a32cc83e9c20358277e72e9b2d63e748
z750b28e180a78453e0cb7797580a991a3db65027307ff5dbdd3499bd4a9dc6a31be02600e7b7b7
zaa9a2f96d79be18c52a52c975dc65b9d0eac544cd58b26f29ae5994a731abcc38ecfa7dd90c484
z2717da89aedb2fe56413daca1a2b8fb9d3702cabe567d62588b4bb4977f1991ee7a1c6c22a321f
z90bc0d2ad5f618c9b225326ed87c47fdc0feecef5ef93bfd003272a2a042a07e610706e92844b7
z899ad52c4be816d8dab67f05c02b95ae0b94b60a2d291c2a66d35f260074d56904da14d2abb545
z49c028667e01a9f5f1824d85bab99a1800c4037062efd1111fab9e76e7e9c6cff0851ecfcfe053
z088b0c5084ae2b99c880c34935c2066864dfba1e58cc3e7ffaff9e95a541b7fe78f7b2d5f92c77
za016718108e5e834f5c5327c6329163f523a0ca9ab9faf899df6502e95901880f3a4402e25b9b6
z9abb5fbdf982e8e316e2117dc66ef29b9d0bd1d8974ebfd9dfafb0203c2da860cf55ebad66a0e0
z353e8baf8803e14dcc3ff30612602672a176ec2dc4ae0980362d2ca1c93eb7b7872b54da6477d3
z4cb4065e8a73c66ada5d19c756b525336477447af1fdb768b23a50132884a143d2fd7d9360f7a0
z828c73621b05e7564e6e6e3a9888146d5e922df8645b53183ab3baa65013144a732389ef230c7a
z289434a3673bff63d5d55ff2fb4bcecce9dfce331a76f8c94d1868789254e2af3f6366ea09f30d
z4c9f25d876a06ecda15942a835274e953ef18ec5f2c900e7ab599ab96e44e1865280966d0b708c
z12b0b2075b2e24549ece3daf9f2374ec7e7720f7c13e872b1eba9fe33aa3fc89658c88372933c8
z7730741374d8cc4309716b0caf2c95ef7a769c9d1317835ceb362f5589b04adee0b41f818a58ae
zfb35bbf0446bcdeb281f2b499ca6d118ff0c684f914838003e5e837d999985bc7a99a166793b1d
zb5206d9e4da95da9eb8f31bf6db7f251fea0c80df68dc31a17078d521856cf7b2d27c82bbbb5c8
z8b4372c53044308662d8cbe307ea72b25177d852f336382512f4c5d8e39ed29993628e6b183fe1
zf8027cf7068665c4c92df55ec414559d88c69b1620071a232010c626f62bc4d69b3c93dca347db
z8be56e218d115cf62a8e1527b96201997e8b5c0c6b18b852114caf4bb7aea4614af78a7c1cd649
za62d1aaefe0051b145af1e3f3f1f419f82570cb371ec5b18af8aa97785edc926ae3376a0e167bd
zc6245cbcf6ccb16da7811b6ac17d2e13f6d564889a813a4caa4de8f10caeb4ca083947eda1098c
ze7fee55e09924129ffc3becfd7a187cf0e6325b52eafad861974f7fa5458c3ef9cf4f605b69f6f
z3998ca36a49f0957605626e6844e755e82d0f5ba1fd5495a21a10ae5bdfd979d6a0ff1bb65a444
zd1782adfa2f49f5eb191f8d3b41783124aa0c6372f7c6c248c62bd675c4973cdd9d501051aadea
zc0eed14e14e6de8c88a6d0d455c5f6493efc4a87383f7626a834ffa3c9e8690f217408df35097a
zd13d5a137c8e4412765a52878d40ac8f79e8ec0ef13c37b523689ceb1f7e39e426f66569c18dca
zd2dac3653ebd4aaaa3c2d525008d5f372abd46446e5f021285ca6bd7cc989b51a73d7cfedc9414
zf15e07a2eb37b65962b8b27b74230aea981cfaf1aa22f1deaeb037b80d30b25901995c15d2c640
zfcb40d1b3f75b835b353e9bec81fe141712bd0d5085197e93678d41042e222bbd62f4c2ea0495d
z8c31684b82b6ad2d04366c650682bb7e056b3953feff83cfa99387547f13b17f61f88b2cbd129e
z166538b84f692fabdaf23591abcdc7713d0ea22428f1ad0462bbba874eef4eb9835cb06466fd38
z78b7e327e6fb83b49fd93ad8afeccb108add34b73c842277a2539e06eb88f10122dea21d39f286
zdd35f186942578c524000f7650b2698cf36218255a0c144749b07fb8484fecadb28154dfd6137a
zcbd97a8a2dcbd01edb19da21f5b8193ba943acbc02fac02ff8e291d9f772949f56fa38a8398009
z0ef6144c0f5b9f7b7f0f4a42f1526859bdf883f6a3fd0814c6b7a96a2bf3c7cc19285ccc8eb33f
zc575fa1809b4b2af9e785a4ee07ca800373554e9220e9342c96ff99e4e6853e7238dd435a1e772
zd7075186fd506a816059c14003787871a1c7fc081632953dc40b98eacc3679945636cd443596f9
z4854272b7f3f0f804c9859e1a7a4a94cd01dd5fbb1035df946c50f8f17aa9280005589cde636bc
z5fc67ab56cd572f3a434f8326a127f141aa81c79a4c314f08814ca63d2887b3aa70bd4cc50d8e8
zada0f3b3434cbd90bdc685ff316c29089c4d80837c31b3dd04b3bb36d9f13dd97ab280eae0153c
z5802feaa45266b81d885214ac256c823dfa26cb1ce45890f65a03a96e6feba731c7a294460e939
z251bec9f713616855880c3113c5fe499dc4b7fbe75173f23df1200f8ecd8ba9be38b86386cf14f
z77e3a4c5d5f2a26944ae5389d72cfdfa0d8c3d2632480770cf46a555de99b58839bdc9ad1eb6b8
z59943eea5ef9da34ae66ad1bb837932ebf4557b9191658f05d04c3752fc8293b50b72039a449b0
z167bd122da6c77aa9de0eb2c0642544af3e97272317d078d4979f95aaab98a3ee685d7de33250d
zb968cfca9953924a4ad8fea45b2146f78592936a0f9dbe496d2e991687c3f59b1561edb4f6c216
z3777b6178a2ad3104c7434768ad965b9123484f1b2a126d21c47340db6d8fdb3fd984d9367939d
z66f5b3771158d4aaf236a5f9d36082c9021cb9deb3a5f43f1454debd2e4e45a7d5c14b3e1679f0
z7bca5b1d02cad2432efb7a7f66ab415a827b81d3a9e5d04fa04e66874a4cd0024b832693606490
z54d8a5ecd2388cb3891adeee2d0354b8c56eeeb7db234bd1b88e69d6d05ead5830a20555faf7d6
zd88050aae64c252dff32d6f4d7f6c43e14cc82beb1d0fa4c325c74e6a9a4ed318498b359de4ab7
z6c08bfa60ea7c0ef604fef8a4938d9fd4b8409a09c1f09fb61c2a36190d00df88680979b773cde
z702cc3295e192f3949d8e5b5d1226a0f966ae8ce84919483fc4f6fb36ddae08fc00bf692ac6a2f
zb6f37ea217b15950024ec0447473693a9349a8c7d5ecd64fac85063d94872f747d3505a2e1ac59
zc08ea223317119eaaed60dfc07bee372ee6df7d422682a1cd25bbeefbb1de02748e71b766a6571
ze8463ad8906f004de56356f2f87db4dfddf71120d70500c30435a4fe199c568b878f0785bf3c89
z5a7bd5d50391ff63b9289343d224365c76ba92249bd44e5002704d494b534a66d7919bc4239e13
z173f0f29852e30611990357ffe920bb8f245182d6805a3a7d50497bb1c2e96d16fd1352b02e3db
zdf9388178aefecc02be7a00ecd5607878da2c1d688f853edbc4b54cf6b6f7f4b4a06d6274011c2
z2211ee299e58cfda90c0c6bc2998a30512a60db81313057088842ec8be00be425c17aa6b98cee2
ze3145861ff482146ddf7edd1bc283a7050f26e3eca9cee388d509b8e18d1a183150585a666e59c
zca73a92a1c0fb0d69cab402bd058c7bfc68fc3d52034b293ccf714be9742c6a50cc178b47dc6e5
z63048daeaa9717f8432996e72c65c2eef666158976225f49f12a1501630037b76e941c82f652fa
z3ee6a1198bcffb91e38a61d643285f8fe3722e36a796ed90bb0f388c95e3a8c4508dc9134fcc69
zc6e7af2666338d2ee020bb63557d7fbb54ffd0842970649ecd3165734725c605bf61117daf34c3
z99dc9451209e237eef039bb6239b1ec77774a21c9b939fecec5193e9872dd6e72ed4a4aa6529fe
z25dc7c2d310e1439895da027be77d60a8d6b1a429d025077951d9612880b29802df6afefba0ab4
z4977a8894b08e53762cba9adf15f0a489c9dcebd34c956bdcf88e3ea757df09aa1bb44c5d37fe9
z8459ed109922321cfac34b204ab95ee3c1aad4e1c76e64dd08d86109619b2b743705f694a55ec0
z76abe52fe6eaa746ff72e10f67b257850bcbef8db9242004d1a1a5524e00e1969ba0522bb576e1
z8ae6a41441d35ef0728ab36e392f3421c1b8bb3cefad9d251b68702f8f30fc24d65b133fade34c
z64eda90350dc9a210a2e39cd0ad644133dcd64e9f4a7920f28cf086425619997a520cf812ddd93
ze85c3baa882ba515d5f083044c80fc6e2b8f4c5cc9f6dd4327d158c76d810e8975f7ef7b9a6ddf
z9ee0b879882cdf324743d3788df5596bb69a1aedd0bcb2abc62c976dc381dab5c795cd4814241c
z7b7c29e4be946efd92b8cfa0f1d52ba570311ac87fb3a4e425cf5e4d3d777e784bcac8ac4dad87
z9f2a2bd5d9ac9e8ecd57df1cd8a7e81b914ec44a1835010b587423ad76fcd591de242a7d53b85d
z824d86aa2c843169b64449566f77e6bf0ffd5956935d1919e8483bc0d8d91529442706b49d8f94
za3ddac6d7911b044140b19940e58d54881088f7b132681979061507edbcdd0e729f98fef0edc7f
za1b528f4c53592f99671ca96125fb8f9be9b665bf17c132884ae3082c518c19bd923d913a8d3bd
z506e06d95f74613554ab08ee654972af969ec84f6b020bd22afe7c09ee9443cafbffae840c11ff
ze9cd615c7d33d7234035f449af16d44b0ae4b6f0ca2a755ac519e87ac2046026c64fa701a1cce1
z9354f3839174a526396227db4047405854666c7620f69bfe019e32c841f6413a5847e56e11cd97
zf4ca68c06f2ee3e8ec6c13f4af27470fed414067469a67eac2fd06d25b709f3423858c0a14b756
z632597e931c640e746d311f6f39bbb7ae9db4aed2a0db5b9c7b8de23e1c5aa5b446b4ff4a1483b
z9b5273c74f87ea76f2ad0d0669aac81f4dea50e6614f7efe475af5ab7d2f46e618b97ddcd1a4f4
z57692d3dd659d13d302ceef42730c88fbb0ec2ddcce58955deb94ad9477522c0ba49214e7262e3
z0c302bbeb2d9ee82401b7125324ca644ed7e7f30f731083ce394a6cb3e6d9a92a538c7e511c775
z03d6c46de084e316a8d0f5c2e8157be2422ab464ef0db3ce511dc9cc713271b8ee69bc0b8ca50d
ze4629d34390e9f4d4fcafcdab33d76b528dbb7310080138418e4dbad9d33ffd0f1e8fff71f27d3
z03fa535ef47a2647446169fbf200365733dfe73e6b5c3f9436d4f9d542b405a6f70464043eb211
z2e06c020bf3a97649a0fdb63a3b07e12342bcee371d84cccb7f7d21dc6935eac7b294298357398
zbd6327d2197c4f814d6c08778ed402b705f7d73ec47bde83b9ceb81cd13225e6635f6d0eb82545
z63c5c3762a8108883ca5ce44fa7dbc1d250ff4ca45b057d4d0fb42b0151f8e94e05452f4596332
z1dd6d793af0cb6c85ef69cf7cba33870f1e0d581907a1be228a9e2bbd60dbff09b9aeca321c210
z10369d845e79f011d6cddda7532e9b452782a402294e8fc864a83224e2f278ef4d2ec8581acaf1
zea64c6b036c4abc2ed1e194ed4681b58aed34b8e320c58fb2281622cbcd65a84138780f343bebd
z098aad7ee3a085137e620429dd46efbeae0101892a038e1593b7960412caef64622d9b222c5290
z64a9a8206a6cdedbafe5526812ccb1096cb88cbb16555a1d5a333771928b239401f232231784a4
z8f1bf5e0718223f1031762c83c3709b50453bbeae867d70c400d294a99ce8ac3a37fcc8c453ae2
z6c16976a3bb86f00ea14fa3b7f071baea70d4fe57efe97752121d9d671c9d8c1eacb71f69e10cf
z0ba0ed3426d2ac23b185ef3c60fb0ccedc504add259d9a8229df6855839a091edadf465754fd35
z9ecfdc46199c2f7331d6bcd586dbcab1688131b24e01cbd1ece81cab9620f1cc10723af34a6ade
zd680ed623782643e646b7cda82299115c8a7fc40ff6c4a772f542ae1dab834f160953598fd9297
z4df06898ed04552dc146e58696c4faee72c0dfaf5600e38402bf8a7c5333d406762b343827f32b
z68dd359b6eefc933eea0452a5e6e044c57b962e4a7fc75a3b6954acb1f2a282cfc3ca6a57fa394
z7047c1d4e2a3e43d04fe547f3e526388b03b21c4992a9a39c571cbafdee5521293d1d64dae3c02
z9897caa9821dfbbc26b4e6ac8a06855f2358f75a4bc8e758fbc4650fba9eca9ab47b578a2f8a04
z3d40d185c8730ca596bfdde25b5bb7ddb9333c39b61b38e88f346123add94035e21291812e74e1
zd5f20ce0a3933515e0dde3e58b9b49078a9d83311e64b0d5af1c9eab28d795a668d13afbea0b85
z8f6b07b0ca05c56ba359a1961eb9297b0faeda43874977e09db99879b459e143d33cd3026cc2b5
z7f70996445c2c71485c95b3c39123fc609e12e4d636b2f4f8534967d828ccbec284644839d4434
zf196e3438973457f5c9b3ac94caca97c5c746bebdd768ff8a816a35fc889c16db1722dec45e0ca
zd749c4ca5f122fe8b434bae0b472159d5844ee9ab6ca9cf0dc2040c83b574775bf239ced533aa4
z13c807d5b6427b712e94878873a28286379039183bb13569a8860dab391f7aa689954faa8ec75b
z9c4cf102a4fbb63f2f296e5f093baf87cec61910534d04daf6fa378d12e0944a40a9e293f4ebb3
ze69a0a2113931c4e6cb14c7a2f7d6286d0888fdfce48ada9779e7e84cfa060a9806709fe7f0997
z5ba598dad4f309350640f7f6e336fac54649ff7813aaad0be2717129b8446ad339456207ada0fe
z0f865754e0a46a3c52b14829d32a301f3a74146752b0de0b206e6b5e80bf9ef34ef59ee8ca1f84
z0d584a037d9995be155a48c57d7dd004a66d3d2cfff813913bd31379d461993eb555b89852f0d0
zf52fb757e6f6d709f8a527bceb099a65ec952a218f5e4664bfbb253dfd0f9dec11f7dafb78b406
z624300fdcfb6d136fddf81416d7ebc3675daf5aec254f4dd0cda5bcd5a33b4da33b907276e00fc
z33f845cf993a3ce795a8a264d557f9d560588e5f57b4ede36dcf4e97a154763b5ca107d2dc7e92
z38b8a96b35a9d3afe205fe6487031f857027dc6d355a3d8b4cd1750e61232ae936ff6f569e6c74
z2461f82edf07456d31431cd853b127bd9e18453a0f5be7d384f8ce8f07db9ae61a3b1abd066eb8
ze9a54d10914fb0b77fa94d6d5cc5c9fdd819af8d2afd50404e5ae9032d49a877c0662f974d54e9
z98d25f316621e5445a7027290af7106fdae8019494c6accc56f99de87dc1e65d3456db87792992
zbbe949251a16059f015e66753915ef998662bcacca24e8ddb1637f3a0853556a07e609a83d3060
z9d94a5be998aa7694dd68b4ff3984ae25c27bb1ad749e179af64e22aa6f20b028d498e8f05ad31
z40aba32ab4356f1e259a2bae33feadb997b61292ace329abbdb7106b413c7ca74f7d9ef473346b
z0ce049195b94a35837e8d0fc2506f4c62868482a02ae74ab60077ed6bc8d319608dfd29117e11f
zb4484865ada55a7999edf465a28dc7edb38115d70eaa6ee6323c00f971989e731feb7b8b0a18b5
z185baa6bce6c62c32fb8222b8e5e8d2fd0a62baac250cba392a944f833e3f2b2cb60f395ff4f6e
z65aa13b47e4275edd9d769a8eae0532bbbab22be36bf8e811ee1fc93b631d0f1f8c9d66f377924
zbdbc32b2fba766cb002d848fb8ebe24857934a6ab3b69506a50a73dc7115faae50b806b69f4a7d
z2443d16631e0e87450bc37787bfe12db7b51fc2c2196ca95568f4bb348a955371a4f971792739d
zc0899eda652fde66297331ba2fb4ce5cb674f12a452b49d4606cc81d2ab7371fac2b82a28db133
z3b1e7deadd10970bed683c4fa8a6cfa21556fc130633e645ef5405a00ba030dcdf0b706ea7c39a
z888e5554f1affe7144def071ba2f24c2161322e05b09ae0787fa59efe3a5ed7612810142d14800
z18f3c7a1791320a5b2f552a999a2db061c848a4fe28ec3879226d682f7bcad564dcd4f457a931e
z44802520e0c6b7742cea0f6305534071767e17351c56933f0364012f2994d8a92e721d4b119ec0
z0a9de1ee1f22c8293ce13a0e81554a103fb3e8ab2c910aba6c13edf3af5ac7438575867ed39268
ze853b815473c7a7bcae40806d13ecce9d6f3f21c8436000149489c26ef4ff051bc61a920504875
z04ef59d959cc4b7b88a2e5b68ffa90d930db8999c9cd94a5051c1581b7629621ce97a1e2e82d58
zf40d55d8e005554f6042e4a99adfac8a8b578b62c84f2483f80df039121f4c2390ac251439316f
zb90a46e4b81b724e931730c60a95a626bbc6da86f03cdaca6c335c9e93c49108bc9ca32fa877f3
z87cf7d3793b00683cc6582a8e150d53050bd386ea32cdb9235801091c676e103ab38f84e421311
z60f9c7f2b067d4d8ab5ba84623a29d76a7f0c54a2fd36bea2ce6c63a828258290e5637236f645a
zcb64034447c1108ffce82bd445ef8d3633a8142a31f8fe4713e6ead0a53ff7d4809099b6f7e648
z011d728d920f06da35f7dfa9d9a93f15d1aa91072c52c7e2fff69ef26419bfc5f1af895f348d5d
z645e13616e86e6344c51890003b2533fde6fc50810caf2c162e762af2018188af3a435b67199eb
z29b9b3d1a4a9d231284132e2f9caa6dd0cbbc116d3727b6e63b8ffeb107df8bc4eb9f9726198f3
zd2e8af5c9c2094bff375c4d456f6c60e266060637e1265f89d39f59ef21fb8c6645e2dd959234a
zd47a005cb5646c37cd4028e7bead623cdee7a993fdf304cd444ba2669a9e9c5b9e5f939c7a6766
ze53218860a8053992adaa7ce9c7da9e947033df0b66a45b7dfbe576f1489077ef503a752d9c057
z35048335667590e8c757d285d1cfe01a79401e54746055826db0a3f0a0aed8c50f76197f932f3a
zfbcd1b70a214440772feafa0d14c5f22c0316fba4ca0fd8673ceb677ec364ce52f8ea300cf93d5
z6b2644ec0e67b67be64243252884dcbee07b20005ee9ed9d21c2c0a41677159e97389327c31427
z08c08999c6c077e8c7ee77613ac292acec8ce04a9ba0ff887ce2dbf1b09515406cb33035adc943
zd18b9c6b040998ad2ff1f10d3ee091238a36760cb918eebfde1c5e57180af91e8e90627e16a626
z93f783387eccded8f6225c3dcc1b84633a4b1071d3b97a6c5b25aabdae4105e0e0b32ae5351b8e
zff2544aefff3a3c34c3b9f9471058eaf85993b570a54e225b975d731f36d5768f269c9dd0079b2
zc83a0b882502b65da90a231760e1cfe2a3ac34821827bc034a00707f3cb624d49d84582d378695
z28ceea1971bc2225400f5275bd2296977b54efd26e279ca9fd99b91d2b84dce6849f259694a5a8
z3b3ebdb5e19db5a5975e11c77a771ee3ab83d541f8fe84bc0ab3d2f5e7eb461bd795803a62c66b
zbfadf0cde85483cbce513d4277ee707db7d703bc34feba462c42edbcad625126a92016d6a340cf
zaa25b380e4718379229d02aa84e737aaac1ffa2764f24420ec75817a3f2b85f1b0685da6e41585
ze5b421c978010f0cf02a7142e04cfda50df2c1221bb8b950943db0c1dd256b3bf203b0680c33f3
za10c91cdaedc7be0732af32f66b0af3581aa0aa5aacba6821eb689aa5dbd53005a42a03600e7b7
z4d5a7ef4da20ab73a8e150ff94182164d9879b9c196218fb9f67ffd03fdf9641b247f74306827c
z4eaa7999f94d2005dd8c5d5c8b8534e9656edf434b5d82cc1418deece3e6d0294098442039cf0e
z5bd6f0ce032d1f7e678da390f2e7e17d956073ca5f5e39a810673e5f83a0bbad5b03432ac159eb
zd2f640aa8f9d39dfbf63f35b9eb1b15927a00da0bd79a4b08c23b5ea747931efc0843a7fe5a01c
z9432ae82dae197e9cd9f506bb3d9ace8ba729ec28ae09409f99bd408cc9c6de652b2a058d23e74
ze25d433482f1598c6b68b4ec7e5b122c8efcf6ed9ee45f84de90485db9d0b136e5b73616bde183
z97b16ab9a6e1dc07e7ac8ba0b07a6372ebe7f066116e28ec988f2e4b34467711f973e95398ab39
zb7df6237babb43ff4489ac5c30da73a5d3dc9e36e756ca5a3aa8fd2c74353141576c24a90d6502
zc09a2118f8f09586a25ac3124a74c9647292864fa40034c6718db4a7aac61ec30eb000337ab82e
zf2633c923816ea026b2e36253683bc604681528725ea1c662a450d7ade29080ccc4926d2005f32
z0645ab374415587648095d5ecc9f671c75d372abe9f479efc8e82647d60c6737be38b40d39acaa
zaeefa22935fa8fa7edca3973952741d6de96c21884195c9bf91eeff392f65a1bc7d1727afc41f8
z548ed422021ae856229436883ee6df77222106046508a32d196d03b42025265d57cf7e6d219cd9
z474b3f87a9e72001ddfff9b03c303d8a45a6ca7100bc6973fb5d78aa129062f21a49fa7cf5f391
zcbd3a350bb8fb4f7a062cf2a793cf1a0d17d73cfdd348af82074accd49a301ee092c891d928f43
z4200977de9949025e7beefd9c5e2a43260d0a6767e2aea8110f37d18946a61c1b9809405b97a7a
z9fcb9cc95fa971acb5afabcba6bf5a9238e7fafc2adbe04c810eb69b5da9cfa254c91e223f62ce
z31752b4e2c8cceca6125770baeb931c4dfc81f878a4bd690b60160a5b3c01d3ca83d9d8508a3b0
z762012534b90ad22a721946b8049bdc7e3119bf0a5a847cdb3449c23992ebb7ecb21ff02d35e03
z2d228bc1ad529ef19cba6731cb0edd34252c0458a54695dbebf33b8fca1d81c3dcb3e84bb5399a
zd46f965abfd8c5ee7083f5599b5888f8493220a6d21bb7dd3b05544bda0798f39990a5951c35b3
z4bb6ee18fc6863aafeae0ce4cce7b180327bd11a48e3c785058744bc6b453c6d95702d6a04694e
zb9bcabd51dc01c8702e7ca00f883dbaa2ee6bca0308ae6e540e166c346baf8530148443b13ce8f
z5e532c745dbc2fe9eb4f49dcf43fcec59ce0189f42d7f0185c14d47b65610d15decdb0996f4a5f
z595469d70f9789a4b0181eb2d13ffd432c9cfdd519090f363279cdd0adace57f70f3fd12dbd877
ze249d2421fd8869b3cf4c51a9830714d7d11f3196f6a5b8236b9136717c0e5e0d92de811097262
z95fac4f7c040095aa2cec24174227977fafd3fa4405f3b9e5fafc1c467877ea26111dbbd266737
z94deeb3b66277fbe792c3f242b8eef08879f46400a442972904e3d009eff3257e3ef7d6f5e72df
z0dd6e442f056cec1b5e728fc7f73cb608071febd1f711e2e470887cc7b0eeb341fe9f9ed6c2611
zd00a6b021903701fc689ec9cb3c6680fba9728b1dbde66d2a6211c82ce317190315fd2e7636224
z8db522c65a542224fdfb542111f8daa1c4ab215c7a85f3a12fdf66103a241680dc2d6bbda67750
z8229df6b6eccfd9786c49b3d7d0ea7edbef96d2c99306dc1211a9c328c11a1b24b5188dc642d1c
zedff4f6a96062992096afb24e9c8aa4514eb753f775a4a01c1352a0173f8e68b5744708a23a39c
zaf175d7b8e153c20124ccb2e751543f8fc9c24a421b8b8e5b391113b700616d5f673d20046f867
z7816902f30df1d4e1661cefcc768be068c6602ae2a5137cdab53c65c67526812394531962628fd
z795e5f07854c00db546135b33975492b1dd18100ea5345b3f61262d2e0a03cb751ebad2fe5d92b
z221b53d0311ea979359867925a6f0b8d3beaf0270fb599fd3bb973c070ff2b6f920b0005093f78
z8eec15e1bd53dd1c457258f7f1492f50e4f28f2494fbefa4baabe0348980f640133baf1a96b5dd
z9023153f137023c94fd0491203ff9ee69ddd2aeecf801f953454bb7ac0767ed1c24337c13340f9
z56a990d9dff68826ae64a46e2934800179793b48937a8ba2a91d5362ac52162119e721d25d4f72
zd7b3eb0310dddc1efd101f4f18a0a77538bab91656672f41d1e13467b81f316ad1c9982c581395
zb4d60e53937df64e40f86f770b4c28c562c133fabd55f80fd36f1922b318fe9a1db648f0123ab3
z7efd12e6107dcfd80826126b07d2ba932a63c5356c37bfe6f34322894394ea6ac1feb990f56099
ze6d59ffc1d7bf1ec2ac5982c12e1532e5692133e10adec39c9e5a4b8e06a23e6ea65457e54bee0
z9a87c0343e4720534dacad4119a820dc174a575f8a3a17c2059fa60da3cc02d8ee8a17b3b5f6df
z561ff31a80349a3843f3cabf234995118476b0ad940a644e4540d0ca410b933079b386579cc83a
zf62749f731d8e652852e1f34e824b34a17d005d0a8d60d48b67c8c08f2484905cd1d99191e843a
z581b536b1a8aede5f9e0fd82a82d24d0b8f43c1a632af362274a4f8356451293553b766f4e3fad
zf52f3c2c2711239a8ad0c99bfcf5902b84837f1c8c8874357ff2c3ab35128dc5d807807ca990c1
zddbe5a9469dffc18888857ae900fa5d57499d45d76a26d23f6ba57d1e30873192bccc49d42ae58
z78ee9ea9ec007887cca3bc04d5ad604e1511628d94acaf732c4ed220ad9a2ab1d3b94ec0d46a88
ze7d276f4a67505976659d16f78d128c44dd73618d85b043444516072a704f5674bdc3a02199a08
z44e1d1bab4ae510e3e4a59d5da87ef6f78359ffe5a828bc7aaf2aac1d76f51d5646d3f523c653b
za5fbe859f36ce30c0c2166fe52164bb1142018602b7635bd44c84633175565c6cdacd8d5931517
z32bb97127a3fb91391a68cdd6e9d5ec3c6c7ac793248d4b3efcb4a4bde012986ce15ce8bbf23fa
zc8ac4a627721ac95b3b15e79ef49f2d61d962311fc462117306da9a2036e15aad2a39289e7acf6
zc28441daa50a95c4abc69f66ae2afa579ecb4f30ea81677879c32b826a77642371252c7e668863
z3c600313c420044d5db5d8653e7021ece1aa3d7062360c408a727a22fb312e4b7bbd67fe1737da
zffaf86578a94b11dd693569183a4e7204c7e7b0fddad495b84f2170ad1bf019dc3e2c2a8eadb6b
z1d18f727f1e8ef863eb94348c83a01d55be117fdaee26bdf0c0132f363b58b3f9857a753c7cee1
zdfd2f857b547e55bd46569275528942fe44e3125941b8738c43b895a1e4670fca499421f43c1bd
z48ada31fef861d67de883676478771edc74fe04e0581053dcbaec35cd4d2ebb3754f0cdf5f6b05
z33e3e7020331ba420fa3de84643e1bf1339ba1fc3bb67dc1cacea46137fcc4ccb6c33a5ac4e460
zbc26961a05843dbc27cda3c01e4c9c69b94e2602bec38302aef3f864d3a9b748077e298ebcda34
zaa495a7914402c3d64c23e31711b5cca38aedf0e5aa0de8a1e6df82049a59b25fba9f6cc4f98b5
ze4e0f239a69dd6a13ada5af221dc637416fc26cf7ab6f60458d3144b6f125a048756209c382887
zb136b544eaf468f318fa9ce73d7c2c2d99449f90d81d9aa8d1eafb0c80502e589e9860f3e9c3e1
z5d2c558702657aa47e99da4bee989ac5a81d3e1fb6e1c8bc72374df0d7efb5d43584ceb29a1cc3
z3321420d13e0b6376fa3922970b8f1e6584dcaf7c0e13a9096f9418c23a3611ca108c4a2dd769e
zfa26e7947244e6c033224aa5acca8a360346ef9d1832b8de84cf04333e11695d7d0538f91d7f9b
z388d676b31816cfae13f4608b97848cb176183f26e0fcbbc61031feb93533a50efa5b98d8f5c52
za8234be4af153b231453a94c821e0f3dd598f2461ca093582696ae04ce2df1ffe82b0c7bbc1d26
zfc3e01a53f63329b955be443e9897b74ec01ebd4e331304d53805b724dfbb8335e9051836138fd
zc826f08ccb4237ed1583fa9301a1db0c5d4afc3131a05c3dcd9e2db37c0e3bdc23d9a22211f4e5
zab8989a8f41dbc66b94b2c91fd4f57c91e8e00e538154bb11ec9b9404728ed20fdca2fbc57e3a0
zdfb340edf055ce72ae9ef5c98f06705466a17866168a7d3c5238288dc483c396d29ee48506293d
zda15243d477fb42e44423c6caf822e1dc685ee0879fc41545bcbd1f94c6303ded734c7aea90a58
zce0ef2d77cee2097ecb5002711825d4d64900fc25a241140ec94b6d69ff0c09bdaca94a9c37f5f
z65094a2edb7bbd81f51872181c42343a605d1129ab474ecf3b075e67c6577fc921085a0d1cbb61
ze2887bd2fc0ce04167a01f3ab4e31c4ca9d5830a87b8ff995e0c0d296b2e754042112447239fca
za6f1233363abf6b1529538a5291a582138e804e6071271390491db544b99c483323d71e3a561bb
z23301034c1503d7ebd5c63cbe3b2e58bc4da0bdd615dea5f990c38c2e816c708588237bc9af519
z00fecd3fa545d7640969a1af724d6fa02a6a6fb722dc630d0d6e887ae4dc83613dfd7503c50f0b
z634c79f1756ce14decc89bd0c66b3f89ce8a5e9adfa710c86825c9d2834165bced54acb88bbccb
z5fb89cbbc6cd7cc86bc5701e71b6c29a228b116e8fbafbeaf6b9a11982b2634b92620f1bf4cf37
zb79864c8569a22d742e32ba2f8948ac30a148666c690ad5a4e5ddc2b4130693d3ca468c0981da2
z3a96391d3d1e7d04c085924f06283fbdf17c297458efbe8ffe0b394765ca4c9dc158e20d581555
zd3c2b6925d302e284129b3adb70296feac8f1dae3fe93990ff023d55eac7b1798aca1c1dbf8c65
za573f6fcba67af71426f79ab99813ec6ad47ab97b9a471bd892bdc508cb91c72b9e323d0f278f0
z9e7a5a3f2571d7eb0f72862ccbbb58ede527f64a4d9521856ac4274d441911ea6e0af05af451a1
z451065f39054c926d3af046b3b83d776091616c753e6fc8796a755b1a0acd40e9d0143d4c833e3
z37cb212958ad106bab5ded31f27a8697bce6455b6cc3c6e0a248f1ae1d53198b8f48ae08b79856
z352637a9f914149bc8b978e1af77e287bdd7559205f54c311f31422617ead4eafdddc901b9f93d
z20b48af3b704236cdca9030ea77cd658cd0a4cc8f5709e880e923fcf17e9de1697907a78d89dc8
zda4ee109fa15342665b28e48dfd5c3a3918e7b725a64ef710c389db5b8ece45538ed0f69966f8b
za51ba788cb79b94d0e04f30e6e88d0324e0ccfd3a4aefa08201ae92d27cbe3e852ee0a54c60c0d
z6781c546698a9b48b4015b32115c91d23ef02272877d56b687aeaab792ba829495546ef123dc42
zfe15fe4c3cbe269c410c5e8b8c2158b531d14b8d34b475161134d6d4ae01424799ffdb3ab38abc
z2c52b86dc013dd438eda6f3c2658ddeebab3c2895232ff84d8448abb6ac712af8d4afcb748ba90
z9dc6952f7ffa4a64e98e2aa0d103eb331e4bb446973da330f547ed196bd0b2f15b4a6df0a863c5
z014ea74b41aa96d688c22c62aead980213c3ed667f57dc0cf48951c4048ef51a958ccdf38ae5cd
z16b543bc83997f85653e0b4ed6ae2231184667018b191a04f773db78a0e55ff0979d5acc1a0ffc
z4efafe298af6d8be874f7f551fe1780d28010990d5e908bc03f85faf267b472825996b9947c116
z808e64466ba30629fad8dfa9585cd0c68a7dde2d6686a9e7fe874dd9d63896657f20387aaf5b2d
zda853bbda04ec59a089ca6960db8b0f2facd85c525349efc5e31062e8c4aa726d96fefdddf0c86
zdcf4c8c12fa3b4f022247effaa389432b1df990d31cb24ada42db50b3f2004fa637ce778b2022f
z0fdfd8e8b4dad62aa006944165a8d2b3c32268774c4843034958d7b9ae90fb1a6fe1ca8369f68c
z181283bd087893d8bd7b64e3b7531d90ce9bd7f95a925ee0605f5413206d36016c38c4e613752d
z2073b53f7d6d795e535ec22541841a0f2caad9cc83fa2eddc7c1dae97235b94fe7f03a1d2b9f0b
zabb631e53b46af8b5864ba0552ad09193db39382b3d04844799fef8c6584dd38c3801d608714a7
z012d37021640ec65d5a336f2550e4822f7bc8411e5de271f8fe21020eb7b2c8c5f79df932c3774
z139378a56bed33829f79c70ba9bfa883c6aca2d5915df320ce7ee0b373e1bcb30adaf8d0cdead1
z55833e11ba4bbb646f58165c04941d0557118ff1b6cb8333757e77aad88ac32451a8d0a14c8564
z8daf10f04a89145c2238f11b9ce3a6d0303295f22e40cb1cde23e87d7ac7e3ebfe1e382e776501
z3e21976cefaafff28c1b8737c6067cc427173a40400f40e142e61ec5f10d0ac1f8738cc4542105
z6fdb0261d687aebf9e505cd776713a58f60434b05c3a85901434fad7a4d7cc0b4b66272e68d9f6
z620cbbc59a34c040681e767d0b6328168b73393b6f6cc98e57f8471e013c1b8914aea749ff6a28
zeaed92a004e12f30f258482507f63d77ae158a16d978e33b8a4e4f58e5eff00e61f757d39704a1
z3073bbb9cde3e5b0db0b03e06324a37c9c59a93a02292ce22d71cec9818d60d47933fb7ddbdc2b
z4cfb321afc896955bb1a4905215c4fbb9c31358cc5603e39fbd6ab8cde37b2d7a7093d2dcf14a5
z04ac80ed74ab69f5706f38423b32a16dcd872c3142a49330b59a0eec3b4271b4d6dffe2c372edb
z93a3a133d21450d4bdd9be9963d7e0508114f3bcabbd891fed468cdb9edd0f1f31a2026cababeb
z5c2cea8799b68e9b624ca0ed8d654b36374e67ad3cfc24fada34fb0f8889323700dbf2ae71c770
z95744685dbcd55433d7070e8dcc0485ff0b37a221a3cb9ffc0a33b795ade583c54aacb21f6dac0
z3396083a1a75e13f57380e0242adf93685a87464c055c5c4c3afdc3e705eefeffde341643ca6a2
z2640139d9170a3849a12f2c33513fba9c959a0a3ab6c27a58ccc396f39bc75d210366dc3b15c05
ze8d96e9c0ffb84dd6f30cfabda06da070051e648a150af5344f4ef39a88c96ec41768fdd4414bf
z830473a6c74c39a2aff2b40bc453a7d660370e24b466d32ec01459ad94ba85ed6d0fa32dc93a11
zed3b438d5849828ad33f13cbe43b12f596512c7d754aac10878d23dca623e240077b5b459d95a6
zb6f742017134753ec123511de5fc809ebc010715ffe1c8a456dda089579fc7da57dc5496dd7ed2
z3d847919e4917a590e182182487a275c2e7ec3ba99ae7f4d49f3009d038ee2ac31ce0c629611ad
zc051a20c6d47ad2254a3d021dc48ac1ddc930f1eea10a44bea3c711801dd0c5f6fd1f2d764c5e3
z4633983655ab2449bbd969a1f64baf4cc93cfdbb5712fa37c30a6631f9f173e8ec801043975381
zb18ea58ed3065e15a00d94685d370e9cf12bfb77cf6bcbdfee23ae023c78eb908a79b6e89583ce
z5ed1d02560f493e374c7a7ebf00c6346ea6881a1e66b813c2b65800fe150b1564c6ec6ecfafdd2
z916ee8c340f4d5ca9bb689238f3f2e230528ab14b9b5e97de5e0bb8a14d26ac36c787b8cd8b8f0
zdf5bf9ed8f66afd213bbd4e829929a822b5f262c066744497d01272de4950ca7856de5597b113f
z701cff14c8c2053d67b5a0f423dd6c4c73cf3f0c5e889a76c81c802dfa179b8d7500927ae6169e
z9cfb729ec7a06e52aa3e76a42a4ed14210d3b6042bc05906e996b35386c9fceee20eb71bcee69d
z9b734887a8e6752cc30f10278a0a9b730fadc6d480af87703026f4e45e9e5bc5876372b2fc5e9d
za6f756886d93ea12ed602726a4df2155e2e3ce0a0bd6007a1ed3530cc4ab52c82c3af7302d440f
z0b81e9052dbf9195b03e3ef3b9fc94e608a3ce065129eb6a9db5176c34ecdf6541c6e39605f29d
zc641bf58e9be2ffa38423294bc19d98cf82ca84e0aec05b9ebecef31cf8d619d40b83d1f2270d4
z5341598f34378f87c27d395e4b5e702dc5b410bef07afb2264bf5b15cb3b802e85ebe42265b10e
z28b9c236c1dbbb917c68a0c5d0d646e43716df8d47e3350ec772a10ee48dac6d133168721241a5
z1b1d0222e323cb5a1f2c800463c3a44c9b111e8dada8e866ef36616120af08fb6d11e191c7d3bf
zd2c76faeffeb61720fcf2cc93c96c305a2991703c5b0fc0fdf799faa098250d0295a25fa2c3dba
z1ec9454e0f885a07a781a860bf47ec3ca8c6c0ae4a2665eadb1ca4e977054748311deb281c4b5b
zd53bc7ffcffca758d4d50caa0c005bcd2a336742496ab7d7d84b69dc223000f169829266898639
zcdb85234baca80e7b34952214843d29c3718b780201033efadbf524ffe9b2de2335b4119047888
z35c56642be976a0a11c2f9203a2da3f99dd0992ccb8a1a88edb4feecb1447facc8689c5ea0a940
z53883b1af0254628ea8180159a2f2980809fc8c9ed75fe291fafabfc89630629eac7ab09c1beae
z7cfba15f796742cb5f3696bfa98da76b581ca51a5d5b8f636a17e3d71433e9fa84df1d757f2590
zdaa5c131a07d0a94ba3c6e346b93ee4a4747f8aa7a292006598d1c5b6753f8ea1371d8ce38f463
z4a39c68e801e0ef51bf30874c39243ac3d16e776b03a5e7cc3c7f9d8ff6aaa2607d4a19b927484
z60e12d1ecf059ee801f94b86002f9eeb542bfeaade8e98b04edd609e45ce163bacfd68302a2e25
zf3e277fd6893b6a2371c970fa1627acb9ad8103585fd5b71e4d8bdb2af2ea76ba81bfe407f54cb
z2d211acb096d1713b6ef033438df79831e07478ae34c6cbeb5f481a99f28fe16c577bb12bc4474
zfc7fb87cb01a533a8505ba2f4379c24cc310d84b1e7fd81d21ee927066f739370a9881e55874b8
zf4d7d5c96c65dafdb0c3645d66d4177536f559589a9a83c508d786d19634ea3979320a998e9399
z2ffdb9fa137c6c70f510e0d869439a66fff2284d78e5e37fee54ba69d0f7a5264c9ccc298c7a54
zfbcaa4e54a2621d1b924a414d3d3263bef8ecae2caff8615e2b537642a9178e6c7d3bde95924af
z9ec7248815bffe69113b61ac14757cfaa4ec5885c2ab7beba9aab2f58184c0ddc5044135933389
z6099d0a09150fc1979a082e2b5766460da3a9b4ad9c4bce37f55e5a57a7ddf4969c405ffe9311d
z30c79e699b40c5f1dcda3944763e8baaeff98760dd9edf2c67065c9dc731155d20bb1fefc4b4a9
z794ca3a1e28a3ba5a89a06eaca9cbedea40d7fa1b4b9fd820d572cae1879958c6f2225f685e1d8
z958e9ef07c1618d4197d47ef08a0271e76fbf4d0878521826971fa04085462a8f03ecb8e12906c
ze54e23311045923d806779915f70a4b5344acad997945a1d9177c71faa88d4ca2a764a36b0c4e8
z79fa04526c87d6a323cfc2af4400d27833e6d4c0e196e753c8524fcacb00923f8eb34db9baccc0
z067eaa1212d6dbb9c68ee4aeab910a06bfd2a39d50c73c929d3f5d71e26693c49b00c805767a14
z339d8bd63bb4a55e2310a2d175a5fa6985ccc4d83d8a5111b4ff79f57156831bbda806e380c3ef
zad80c92999c1f0c80dd73b371f5fa6e9e4f277fb31a98140050ae5b464c71a03235c9c593e6f58
ze6b330b58d89db69c66fe8b85edbe289b0c891e8e049baedba1d98f2f8413a69ba997aec666c85
zd6b745841d32e6c53dedf21f862014a910a5eeeef40681a7440ade0138011ea7f8f55862571e3c
z0b204a361979edd941d6605095146d895d90c53cf32d4cd5c9637a0743bc12869e52a06e3536d9
z14ec633102bc49909f8f1e3df00c710be0cb8f2bb03c11070a5b23566962160f247460890dc370
zb6f31f665f3eba08f3deea3e083bc1594456c0683d0f1b4f3f38e7e69f2b59e46f889255052b1f
z0083e86f7be6683136334424effec4e1fb12d62a7e8fc8bb6d0a72049d57b57f6b18e03a69051f
zbde2056c5bb125e7bfef0ac653ec971d51050f93dbcfefa1ada831f301fcb5b1d0f7d02f427273
zde731f60771533c14bb185a7d8b3394f6071525e75735b986ccb3410eeefc99e0b0cb941886d46
z065c179b73d9912d71722becfcd4712f0299fd5df176b0f4e1e7c6b79acce59d9096e91400a384
zcc05ac3a3c57501f707eec61ab3625220277c6ca71bfa91adc684dc34ccc1bdc7fcdd026bc08de
za6aadefbabb93b611423015ab109fa5bf57665c41a7be8deb6956667e5833f4bf38c1aafff363c
zcaff9aef5e3b9ed2a81de5321533d275569941b9a6e5d4ef68367ec517aa6a95afda621a39f320
z23fcd9a2460ca9f2b8aea33f38dae0f1bc4df20f1820eae52d5f8ab94f17a4dacc4f33f2f3ce85
zacb26345f5c83695aa2e07d3fdd0de4f2738dbe0a3d1fd8f388b322cc73e875bddd91ff45a7680
z13c227b8f3efcdab7fe41165269927f352da8d22080016ab93e5975aba293ec96526f6f0c7fc16
z647da37b8abe222b4e446e35114bb750330edaec04c250552800e8c1bb0615e97739ca1e151f15
z785de0a9f7073590824e3dcf65bd57e9a500c09a014c9affc342d7bc09595fbb3f89d58e41fa88
zf801e94b0060d2835e1dd5e80b06ae31a7355f4cb92c3e95cd9661cb4f6ec1c12f2be0672ab2d1
z462a62652d85e2ce75ba973c98934126312b3790e70a4bbc35fb542dbdc0d18baf7a26a9234a1b
zf93bba21fc253d7c6783772b9d6530505fff0143adf61b0869c5fb73b087d2386a6ec20d58a2d9
z341fde88c4da9ffab852f3f136d72c8b64780e250d9bc2a56208ab2d7a76cfa115b2aa30b0625d
ze373f0d343cb9e5c68cd8f34346ef65dff98551437d606c15675565183aa41176b31b05edab6fb
z60d6eed4bbaf552dde99018866d828951e714f6c4cb732e412559d6242a0cfb88262059a315382
z86ea035cac1e56558b8a2023fc31c65ffbc971456ad12705ed503c7ec98a8b6dbf42c3bbb04d6a
z29e6a58340b8c5719ace0e60a55d127e143041a3c219f290fd9e1583c9910a41ade0bed9cff4c4
z3f2fc79303712cea2812bb572281b53f493f8045cd6cb59c403ad5822f407259c687301e16c731
zc92973682a067c5469c70f0263aac2c3f4633f9865aa10ebfc61aa3709b9f48fbcf89447545fbb
z64ad004f9cbcb1811825cf59253a551cca7372bf865359071b5718d559c6835403bfe63db18fa4
z3ac87b69bd44c26c9171d439b8056c243c0d6e35225aa38d0a4454219fbc54107f3ccf084f775c
z794b2f77501b80481523a54ee98350d038a046c74b717afd7e5a6512573818f725d70a42f34811
z460217ad2998ce750a354d1c9b5afb15776c30b4d268cbf3011c1008eaae2155b3cb06f71153ec
ze5a3493e2ddbab40b0864801588cd4ef9f96bda68bd6fa262a99f0193e09d6509e381cca03cb21
zc39564f7854224f80a95ab95d1517bf5feddfe55f91eab90d3c2b1f20d7d523893642060dcfed5
za6ef89cf210501ade1b8a7a7166187f4cb5386ea5619f0a7f9b2a25c6a6cb6e444a103df772b30
z0e394899e8cbe6ff0ca2750726af19071faeb5cfd8c6a49e8aa7d7b99abe9ea03a5648286cfc98
z62d2e03a4e3cb50260619d33cd3e80162dad837d61baed9c93dd7062227fa1754d75269c36086f
z5c2f0e19a7203c941934f80fd8ce64ac7fb47c0dfca8b16313059367338031e7eba4de04983545
zf2ce8257bdcd89ee8007985f9cf0442e57ab646d0c295c5bd0abd118956c4b4692261363b777d0
z8eec1bba09d668ddf2f81840d19b50fd0660041fe4f2c46a2abb9102306c7a0ca24c9b6b226fe0
z103437e46ae8ca6aeca8a4a4a68c88d93937358a2111ddb2ed6434549fd05fbe30c5c1063c4750
z902d5c26d114830d4e0b13edc7800cf185ff65fcf603d41b86751d329e2f98c15b973112699b46
z4777ae1c738f9197a987fdf5d48486fee50392031fc6d63f2a7ad4a6b012642ad2870a8774ddb2
z60f47a957a735487697c1f8c349bfcda2d28201e3369dcdd7fc3b1ed7361d3c665711518a1ea87
ze73a5049c0203d75f73f805bcb978ec33dc849633624be58c564247afdcba6c7a9fa1c7981900b
zbb04a46453a40e632c8f379345e9d045c45c6140d5a86f77b279686ea5e10bd81eea8713772c01
z3df6a0e1b651467950a8e230a178612165ded3931aa1d199c39acdfdd9c5c7b532c7ae07c644e4
z677076d662a16df3bc2a95ec8114e99674007d5ec6b9f0726519eab1f634dcf1ae84243b5321ef
zd25d3e49b439bb757a9890fcff42c951c7a9f93424e8cda744b687b101dbc618e5b7e2f41fe0ef
z196859384f4038c4e36589e602c43a83be580e3277d47a3e9c16a748e66c4ac80aa7c9ed27e0bd
zdc876bff7bab3b05f58574d2a8c176db675485efa66f7fcceec8c32cad7a70767a96ceaa3fe733
z3a0c9866777b585d624d8e6546346b0393492ea132ebb231bd1416b5fefdc765d53f6d8a8eea3c
za9a929527bbc94bbf36d2f1c1f6dc992db00f5cc567c9e2181b2904a9fcbc048a7c7309a63656f
z8b51b011e1e207d701b9e5052548b7ab10a8b9f03f018df35182e58e99f4ef1e8b90b79317e955
zb1139fad548a1a05d026199ea27932a31e310287cb92b3be610881590a15e5ca2d88595bdd8750
z43cba276f2b299fc47719b149d89f9b22f98484fc4b2c145d83ffefc3b731cf5fdd141c59b1924
zf3e9ccc497e2389ef8ac7a28af175cd7d9144cfa2828a77cc82bbfb2dd42e6a31ba3fa28c54b54
zd29483bd4baed4837a513756dacf3e3d481ccc973cf9bd29eaef59ecdd30495f891cdb1bef81ca
zca8ebfd11b28a92d61b297d1113c24c5215ba256019be641480fecd91e72e82fbd42e06e565f09
z12a184d02ace9eb92fe2e13a0048519afff6d837555dd4c67617132d628065322a316bed43c163
z1d8a71214847bd4a88d2bcb34d9e4b5bed592233686917072a380a49540d859aee4e34fbb1819b
z97ebe66812066b8fa68859d54115bd69e87ac93948d035708d548e5600fe3e5dbdc3f20326f1f5
z0fabdd9edbf979c9554649bf00c84c4463e15ef20df2442bf5301aee73d86363d09ef6c4f930b9
z578ee68ecdf096a970e0165e16d1a7f12b815168809e4632a77be9a3bc3dddab4ec1e6005879d9
zc26f1916650d1c96bd285ad4afa9da423cbab1adb9c4ecea98b483122b4521f396133e35d89921
z70c072a69f3519caad1a22d1200ac31aeaa6c68f0844abe339819b6ccdba876c11a70e3c9b7d5a
z382156be1adb950020516652290c48ebf7bba6d197d66c23a665a4fc5c26870de5ce9f590f0d82
z1cef017e1db9c3ea9c4ce12a54541d4b19b09c586b99147ffc1b6654c7b20ce63b93a1246b8887
za9b1dc6ac82752879e465ab78857477d5f128b2f2b742a649da08145df61df7a8676cfdb632bc4
zdf63cc2a0f913e50a3badded9d3db6f195c23be5d673f74ce99bc49b8e5aabacb5d4dffc341d36
z8f132d9703059004df31cfe9eafa2cd387741108e22bfd6aae9040987a817d3093ed33e57eabeb
z14231346ea62e3df7fadefdc952d6e8c2c4cd6a210dcd97b0fd447b3bb6af8b55e519a4925ae6f
zc9e95915fa902256e7c46c22baf409fdbc5c217f7dde764369a1160a0019754deca6dd34fa6319
za81feee0e30c78b73ed5bac6fdd0cf96f7faf34898405ffb1b769835d7364eb1c795106dcc53e1
z895b2f894c736eae8468a35c15826e9b987d67b860590cefe1c7ffe4a67df085f737d0afc83584
za3baf8276e00a6ba48e8aecad999305fb1e9409182862428ea9c5f3efb5f41c8642079a55918cc
z1c26deb9ea81c28f491f5160bbda7901176d9ec353bcadfc43197c773b3f2f579788183a5b9f95
z61ce66520b1b0ea5c869cc0c9035bc564f9b30677535b4cc1fccb930888bcd5c4898022ad08cf8
z23854a0d1aa28530f608bc3ef6435a5177689e40bb8eacec9218818326758027b66f77319a5d62
z3226f5daec128e20a5d8b4b359220dc4ec62deca4950d7aee7c4ef59872b39d83e2ee912f949cc
z739c20e378f6b144e04f9e96978fe8748c8d2bcfe1a38b15f4cb04e277fc332f21b7e2c9b41a69
ze91f4045464c2b4a966b2ad591ccd0f61087ab0477ef82e0053c70f33f14c37f23cf39795bef41
z9689612e953d1ed94f638193b73323fbde694e86c04bf02da30e4e9893ad238aa25f41d66ee752
z0810272ad7f94d0e447f1eb63c8bf3b730b0c623522baaa16d1ec514cb890236d2c4f9b0ac1926
z825d76522e81f1f6eb2c453684d054db2ee1df76c0c88cebbd962c0c1a761fb2d4430153fa4cc8
z2edcafc36507c1a2090b56ac2cb1b713a989cfd689dcc3cfa0c9ecdde3faf75ac982face70d7b8
zc363759339bac14b6633be082014423d243b61bc7d917f5bd3eb6237f1fa9a88e00191f711574b
z62321ea24c3b582d0a07bfa6e2840772b19b01a65f4d68fa89474902600dcd73b689c1c8fafe46
zdff0c0073fab661d26bd365af181d4a78a2aa0368f99c8783cc45c3d6c89058a82706657cd94b2
z5d084a075bfe0370924c970ca02f99e21db0b7118e1acfab072c24be66b147d51f5f75c2e6ce9b
z56404464ab305b5abc10639ebbd488f5c4a908fa223e184fde16efe8822b1d102c83281db0f261
z54caeec40321e53a446b5399264184cfc2885505c5306b2afac6fbe09d7237d1d881f169b02095
z5af9baf60ae123a2edd5b6985ac3f7920cd3db58c1cd316d8cc8f8e226575d28f5d0e12f6d4f0e
z4eefd7c5d00c2aea75aca05291b5dc5927488f7c19702c713c8e352bb2a330213a5232da864e40
z7ab408e834bfe79a9fbb647d2147d57895725a036c1f55f207f71d1983491cfdc30b05c411369e
z4e2f3af76531ce7726b5b8185cde15a0aae79e47b35fa6326cd64838b1604eea02874e6d8c5b8f
zedba19924208e11a500b4543412923e43842dc6738264b760973dbb5c6a7b027cd8655d77918e5
zbad4fdbb85e9cac224139e0e01070fa41f723f4922140da360143eef9a9684b8c62f6a36dd145a
zdc8e6e3aaf63ad349bb9e1fa6c2193b58a420a50986571ab51a7616ff85c734b8e6e74da236f67
zf4b507b809cef6ce295916c0c149bce6d619b1474b67b92d35a7ae9fec84113de93150a6a20e14
z20307b25368702065a4597a3dd5243e67e3faded698ce71c5f5e8e5866a81ef72f5304b66fcef5
z27cee33ccaf4c16f4886f7e8f20b7fb64aca52d5957dec86efb6cb1086ff5fbb0ee57842f61cba
z18feabc4e8e154360f6fc0f502382434590fdaf7e6c700bd3bbe38fc8b99b7dcb44d128be38991
z178dd7802a7cc01c98e994052e092bb671e85b6fcb71c530e107c1117623eff2296438615ba7bf
z674ee75f0904979a62643b383279e68e7e21ef6a0b798b155b3671c1e3d257ccca36ec238ca0c7
z11dac1376f8c0e886a8269a7a597c4adbcb9c25a008da8ceac47fd0f582cd50e8c022b5e4e1fdc
z7cde8c6d405156a72f0a9d065656b2b9984257d467efcd5b31c1054b551beb6a0a2ccdd3f87876
zd0c0de7fa69dc3be06e9e472945a09bf153d65ea12e22525137deb676c97c2613a603e2419b5ab
z97d20361876a1918b6e7f54966af99d38f82a8802b2ec8210d14d523e785c2314145de5f2a3c2d
z66a941ea8f432a649166e664a0d6fd515e352f6825855756776c08766c3e2c548117aee8e18d88
z980dc774e955ce7dfe2f57adffbe92b11db005ec7cb1ab89f1adabb42df1ba738d66f1e26c4cdb
z7df3139575cefe3aa08d882c0fea8da03138f9a33732b48d137e1e0c00828c8d502996f00d040a
za63078464f379fe9cc4912726015523655841760725f508668327685ca0438104a2092a368f7b5
z74749b9241c80fb034363ffd55d1cc43ff3bd50e53350eb1634ab602cc1beb036fb9dce9713995
z7a02af6105ad1597ed0791381474f43e326bf8795762b8e08346b9dcdf402bd58a6b210595f69d
z1770897204eb32898e02171b60f3735cfff2e746be59e6cd3c1471acfd35210ecca832ee3e622f
z3db59f7c869430669cbe1fb4beedbfc1bf9a295645ed1f003b3bc768d38e0daeec37393c00b968
z6f39f893d922bb9130c5f78970fb9380b744bb66fe37cd2aa483eabd2419e0fe31ab81d3ae118b
zc2cba017ab6230c648a37e500e6e2b91e7dc8966c78bc9532bb324270b9fcdc5879ae038fe4731
z7d1d7fb1e63cbb7cf4c082ebf4b8eed3e1f21ae0de95431aa6301685bf876c0a72cc9dfd8d5336
z60c7c51d812281d526b1d8f858bec64e7062a3d1ba88ca68439d634e5edaa7d0ee2c79a56085aa
zdfa288b11e803a3f708f93ed5f0ca29189a456e42848b5aa057a02de2519b50465f0d60e9759aa
z1cd3199f599e71cef6936413476973a8cbdfee46aa8c256b37eaf5970d2546562239cd6a8c73bd
zf01ab8029ddc32500bf540c660ad3d5ffc486055a3f30a503ea6d7aba709dc1720326816e00a47
zdb9e36edd3d4e2e42ad15ccda3939b5e00f7d9e897a444c18d98473d4845f574c4cc2b66339b13
zd4f61ab8443803814cb4c6aac5679a7adcd8e9e061074057084bb55d8d90ab8dcaeb6c0eba14de
z8b74d05bde4445315ecd7163f58d6896302939e6cee0f1efaf40d5300c5c361b57c0b69de02856
z65a339ed9b5e696158bc774fa778087e39b2c4e222c5a01daa3d7fab7173a867d486100857da3a
z9c080137125a7720012a96d31acabe76d9396b0aa7ae2309d43438b4b8d6f09e6a7477dc6e99d6
zb5830c5362d3754e132d876f3e77f075898b5b8c6380f360c981eabfe1be2480092bfb84797ca0
zdcdc8f4cccf566407c12c558a9c151240bd70fa2cf3bce7cac2d523e45d50314876970bd412f14
zd5e718eb12d479366a23f4fb18131a0bbe8100ea42d616a176278f9aaa985d6fdd2ad1971fe032
z5d154af5682f42f650f8e0c1b1a91d9497c1aef80240ba466ff7b39dc8bf1a3d571cda4bb25186
zc8669609c702635143b845f692f611c58d5c302ad87b60b7167dfd4f2b8b94200a27e2c15bbe9b
z0befce7ac489c55ce4296acef68462dca9da52230328872ff88b0b1b9a97d51310e0bac8903d51
zd5312a3260b1016e81eaf70e5dd94d00854d86e0f0e6adcef7b0ea6c9174a55a1086667e5702ba
z961586f44a16776aa64aa259864fe8f5c7b9403e1b8141204c0dc605978fca8f062c419032d04f
z03d4a867049b784ac7e1b5d88a0e42ba7284a511f30f4ca80dfd56bbeee497870acfbac16527d7
z060f9187b9b88438a090ab5060dc66f42ba7bad7d0ac44334321aaa1c36bf198413b7ccf162b76
zdfa958ec3133d3bacac860183fd61b86ff8d568fcd568d0a95298cdb03adc2aba666d9022040ba
z18d2ef065d608dc81dadc6514802fc402ed887821d11e4a2113236eb1d4d012c76924427f53919
zaa06a2769c5a341bab3d6b4fb3c0ca3b9e8af75d4d4e3764192386ba29f2617e8d82055ad532f6
z7879510e173d36ead15fa7a2863ddca7c46ef62f4088bb8c76e95d975014cbda5481adb8d8cb46
z2278c968ea823b51a50d6035491094f32a1ee9740fa92a7333dca73e8037fcd82f2bef5500af0d
z3c2fcf099c663e5ad0f8791bcba0e842e83c7114f4efaade6819cee6a5e95a9ae4f8b7035e01dd
zd542ba56277d15cbabded4bdd54a27b54f654108b4b4b59976e5316a91b15252a71653e49bdf86
z8a039ffdc933946db6ad34ac45b89900e38f7610d69c13dfeda6280bf695bb2c90868047c89198
z0951c3979c9dcd890a64628327c19ff88d6ac09d7483e02b7837e102c36d88c3fe0fc25d906a5c
zd42756e8882cd55abb82c6aa069d5da48fdad7027943506607b90e0de871758b7a30e3e0a5c500
z69fd4931772db8ed459342545633435cc5205d003c3ee9988d0780bee0e3d05e49af208a0f79f4
z3233190346f95b0ce6fedaae23056ce8d673f35d7e14cedcc057514bea3b5084f8d89c1f187c5c
z15c4af05ae2dce52646040145fc0abd70e4469f2870a2f3151969eb9200b8d901d687724479baa
z0d811ab262aa9b46ed1ccc3fb6168615843f45f546c86265c44ee700e780aab2d1d5d31e4ce8ee
z1ffdcf20ce01a568ebd80b35292bba28a0a8663e8e34fbf2fcc3d04baf61c296138497e0842535
z6cd4e13a16d0292e8ebc22e8494895c13d34603044021111d48a0178829e910cb8f1854141b906
zace0ba42e13173dd7f0c372603b9e2ad437b0ddcd2867af626f4e9b93459fbcb8d4355c4635f3b
zc65b094a285f7a486622784b8ef364e86d93453d7e23587544ea8ee07ebbdf1cdcc7b93d82a566
z37de5aa16bc520660227132c4cef70b0ab33965d8cd5d96ebc35447c3a9e74c3902f2a322da40f
ze3559b186bd82216cd70fcd148eed0bd225768e670c64e7c972c5a2964fbec851aeb9a1ecf3a99
zfa10af18026a36576689e251e88bf7d0097e9231e1ee86d876fd857ff0d8576104cd7c29512da9
zd59adf73f378e5cbf508d72b4ce747bd066dbc6c3688c41a7b729f722b646d131b8770e4cebcdf
z81cc4e2d4eb02c501441c08ce36b4987844b26a969826e85b981a92ed97f86334e01d1f509831c
ze54c040e1d3cec6384a1721160418dc04cb61f39d6a5bfe230734b7b02cd7aa6098261d5e05737
zc006ea9555316622ad5c43e3753af93a2ecfcd316963a4087e5f95cc5b75fe7be65de0d6fcdb40
z7e12eaaf0c9242d5b87f34a35b0736068b3be90bc785859fc5c9486c32f29b28520e7f6b88cdfa
zc75792ef1ed212873f190d11ce9e090c2b40b28e7c82c9554b8a12d36e4ff8c746c3b32395937e
zbbf4fd4408b768e7887e67159ec4758653788705adb7663c3c708b33ac42a5703bfe78e44cf51d
zf9206c8c858cd73b366ffaca8be7a07e406cf1cf8ef06cc2fe5b6f81990d373ea1c226b4ed6b39
z2928bd5ec9f7ae9fb8e5efe6bedf77d80a460c625998138c7028b2298fbab67dc04902f0a4a3d0
z776809c7048df460c9e940026a87d27ec5662eece263bd910416989df5214b085df2c5ffabadd7
z206102889af8de2760047ef47751dc7560a22c1120979b6605906ca16b6a7b9a6a4035de3d98a6
zdf0846ac4ade0ac10e392dffa3494fd72a9d64e8d7cb66b90d1dfc0696305dc5928a4aa0b0c8ac
za7279fd4a9e64e9127a9d44b47cfa107440c9d00c36f2fa123e920c0632f04d859678814bf5409
z5fad76dc82a9c5355d05b8dfb213b8a2e3307115688b99e91a8ec3cc0964348719625c12d1f786
zecc81d00c5714e882db54a0b91e55475490e7bbff1f2d4258cc6b70681505a336ac4c0bbb190ad
z18c7a2bf88daf6bdd5e4b66826d2be809691c56629a44606f933ab87499da1364c6961c4c5be75
ze3343fb39286d74ab994a86f8f19ecb677980cc759fd0187fc766b99e20577c74a41d74d6288e8
z859268246d355fa7ba7a6db29e687141eca66a839714e442f3239a2954d093a3dfa1b3475bf60a
z3bffe657530bd18638e6c737c4c54868ed317d2c8c8ac2cfaf0a0f35966713a6ceb6b8fb962e60
zfea913d5a230e7946d1f17f899c39a8c6005e1b70ada542002883a44db2c56bfeda5b660019035
z75e5026149d785f0c1fc322ef42d11b7ba83b97e7d5757029df96a4e3e2606200cc80cc194d190
z56858cef29f3040a91f5b5bff9c9073c52c5f8ef3d33d969298e8ba97a81d43b347d0ff81611c4
z1f8519c619b791e97d6ce06203a2e18a4f0e08b29fb511bf5abec90b50943efa9da9b52b1c5f28
ze082d1101346b9bdf2875b23f1c5885d58eae4508dca62a7530777166624f47bc66eaed60cd88e
z73a02bef7371b0e84294564e95bcae538af528b4b12cccf2fb1f15ef885e78300b9ff50fd69da4
zdd4d11b05c381c0901868d3972f0eb649efc051f17ee3e3833cec89d18335bffa8a8781b3df20b
zf76a1101631961221b6ab78d4e030f2e824535bc5e30da5a638581d1b421f2b60dea75fa52f2fb
z4f6b00664aa078afbe9285314bab63aa9e36615244023fcf1e3cd0389074034b4de75f0b701851
z42f6a8f3e517d9c2d3f26eb28ace2692ab685d218d6eb637e446d1998c7523d712523271d50549
z2963fd0188dc620faa76fc66b60a24b870046c00d0481df1d43c41398c732411a53a88475d1e83
z79df9d35b3c7e475bfc8f773ce32498c557c9ef9aea0e61fbc4ea39d069b1dad963c17e2844991
zddbbce1cef123df8c3b04b95d0a79fa72edd3ed41f42703c2bf14fd1e2a40e279173509f1c97b1
z23c43c6847c387af4b433779855ae3681e7862617d90710641d06ed48bf5aee2c3aaaf127a9a92
zfedd5c523f2cb5ff3ae94da78b7632da0335a8bc083711e0560f33f280692b7bda7a287548964e
z9c5821fd55bb6a9db0230701c074212763a0d4ac22543e800c274468c451738cd49d2885cc8dd0
zbd9395cebd05e3813491871878a3214307e8d9e668cf0d749263c514c8144fe8481f9b20f92afa
zc94410967ce11c2918e688749393eb5962c7acc572488d76748510e50381a2b255e96f90301797
ze7c19842ea51ba6d4fc74bc54a754045dd870d815c21fe075b7f70dcaaccedca6b8fec1ff2f89e
z5917e4b9ab51e1b4485372f2017b897badff185b8a2f8385dbfa03dfde14f05f173116da4680cb
z5e7f039b0d02007bbd1159e13179cb6bda7de55d5eec746d0a1ea31d1fb3e9c5211966244631a3
z691b5739903a92dd897a88b61ea35d0849008eb7b7c9966a079367c72627edea1e70b21ef466f4
z388d5e2fce0956cda0ec36823bb342240fcf8a0d1a69d92dd15da312900acb12668486ac38f235
z846973bb5919dd16ed6647591e9c9976606308d7ec11b591e28988988b7bfc5cb336fa7f682ae5
zd9dbb1957a2f8f121063c2d26cde3573316d1074086e3a55d9741903ed7f3b32f7c92c2f6109f9
z7de7ffc3fb798af753e6152a612a8d5f1200248a54bb79eed892d4de46dea07c2a200ca5004183
zdf31a2c225341888bd5da62c622022ccf3fa0ee4cf4f712c05db141f14f0af5c9394236d277564
z28788be0b9a4b158772a7070a56ee1fc1d857ebb7848341544f20489dbc9a3fa2e4e97572e6c1a
z623a56a440eeb4c3231f76efb68ccd222004e6ec5769b416934a98ff715edd4dfe5ce4b3caef5b
z72dccb0687e3d11bf88228b1506a0ab450df0a0daf4887df1374535f097e8b67a905f9790abbcb
zb73ab16f5cb262285932ea679fa69d0ac789c7495d094f3bbf26319d5594cd7e75b4a09fd080cd
z9b04109d1f3a3a68ff84c524422ed5bb35b76c6fca8a6eb6f71ff5eb85a727bb26078648519197
z6f2deba17f14a7feb9e8b4194bc136257ed13f5dd1c54fd2d962731de92190cae74c2d2096baac
zedf859ee533486ca70f55a1fa7ea3f0b1a6284a47fec4b1b956047303b428cfa385608ae34cc2a
z698fd1586348184cc6d55f5df7b67b38e0e4c767ba1c444cb9f9d6b013c83dd8c2aa8c725485ee
z0807bda18bea47a126d977da1353270065a565159b238d6de0a009eb0822ac1345ad5ad4a8839a
z65a1e8873eb7dd6ab1f09d0dbcc4d36357f08dccad934df71a1bb53f69959e64019c5784d561f5
z120f0af70b256c9506a81615523e0e34da3008464848e0a058eeee41ca69bdbafb950906bf58be
z1c0c50376a0553bfee421efe1e878b43e40c20e386b7e4273499149f52b3e6366b3ece7c83d1a0
z860ac9e0ff22d17c6f377a2f68b264344abae3e4aa1c847134fd9bf1256b35dbdc36f3ba62b020
z0f3e7ae8a169343569777b57e1519df4e351d2513e08079f99484a33acfe7716a39784de750b77
zfb18c395ac8c0be199b103b78f79d62e41a7b87c8079207843bb53a661c8d0e852c866105fe455
z476c2e9399daef22e34ff2c3d177d5e4ab04e0d3e4128983b8e02626b1b9a34689ec7bc3499a99
z2436a4406d2c56a16f53cfcbf185edd15f1c96380b8964d6f35c63341e575890560922832d3d85
z12bd747bf0d7adae7fc6aa7fb001cc11215a0f0a7d5bbeb902993afe3b612ac4cf3a2232d508a3
z347d9c606c06879b348fc55553db1a5246ea14e8bc9f3f82a593f382a8eef8d871254d1a75a482
za8ec549a39facfcb720c77e2f10154ad39d0e71da4a44c2db8da31fc17f62f81cad03f7b08b8cc
z73fce0f12b9b6e628f2693cbb323009e09dd8f5913c649133c755cbe33db4c622ad0e13f16702c
zdeabddc5db85d034694d63e1a2fb8a9398e383fe1af8f87b122d05219641770d06592858c4c6af
z1d7d303e9d24f270f82fcf7e0460a656c0f79e65058b8c30f84fe50b0083adbabe49e82c97a61f
z1b7680982e6b16f5532e25892025f237160c0badac90cdeb14c9f321693302e7e7c3d2723ab700
z267363adba995a947d2fa428830b0db19bace0334e2f7a9c5d22fdd03010457c89ed1b7343ec6f
zae565722a4714a77af9e879495814e6d8cdcb5761549f525dda8ab0f724f39fe16b90929b37f2d
z75adee502c4189031ec02d45f10ae2ac01729adb5daaaef889897b3b4469b15cf98ac7dc0c5247
z2d940e96ab1501f5af1509443671f15965cc8815638a46cf517f771da104f681163e6f85581920
z9bc57a382d93c672b2443c50a78cb22573b53abe072b1bda79f8bb70ea3fdb61b8058f1ced63d7
z9df43ce307fab088a819d47cf848513e9b13bc7a8cd91f97d23ba6f34748ef6acf385d77f38387
zfa8fa93349bda4d107527c000f7029d3a3c0248451130ffa3e9254d4f110ec8f12215b71f290a1
z431175b73e7a846fb4e5471f36570e3c25959cfebb078650504155a08c15056f5b16dd0b23573b
z289bdb1fd8f478c47f613e48cf0a3b2a2a222288acc2a4191195ebdd5159212e96d87f112e83af
z3ad537998ff3c85d9c10892edef10eaddc1fa1bf3c2c3149f58fcb01aa43f26909823c70175419
z03daf713aad3838172609dda4a7d310a9bc2d991b4b426dbd4f1a14f69311eb38ae1a8467178e5
zacd280cc1e77a06900ce50cc3005baf03112aacfa3dec37cb74f197a5a8ccc4ad4920fab776522
z155ba8a24b4fdb9de6d05149a8e1fb24deb0483f14d016ae37f6b6b3ab9616c9b89c0f1f23c3fa
zae97f5ef5d552561639f9ae9ab960a05695585770128896faca362771fddc5812f432c8caad215
ze5abfcb36da197aa90556eff06b1f4eee0a3e2ddda87a4da7890be1a868898bdebfec05c25c64d
z490fcca7571c5d9af401fe9add578b57192400dd92c23b5c72025592b71762c629005b26f45d91
z1301b2baafaa3ba018d5c28df933c3a908b03a11707f3a3c3b22798312866d8cf2c9485a496aab
z2f28178cc03519401c2382242d8c4846ccf8b7dae2fd6d74f28f783120581183db103ac3446772
zb08fb9197fb6d4a4d03ad3a4aab0ac2aa6dc601698e3d541f8aa0fb2da5483120ce74467e4fab0
z0dcd78295c38c2a60201a1c46da684e1bea2926291c448158c8d186599f36de75a18adce9469ba
zcc1e6a9a4448ae63d9131ddeb658f84101adb5773facbf9f5b96fd043f57486d23ecb7be873b3b
z0285280f84d921ef15c30d8c973f6e39baf96691ba6352c362db1c4628fa298fba6eb531e86550
zbc161d524e6f55355c32c9a48f8ec0111a434ec860393abdedb84a0794c4aafcba151d3a3af873
zb67b172166babca425b5c0fadccf7178da909192f6396a4e083483b79ae3c812f4e7fdf4263311
ze9e5e2ffe4899d8d8c1451fe34ae0e21c65c55c69bedf64b45f2df3f272d3cf34d1f120878932c
zce29699c41e44e80f3aae120e519ee994424133892ab667d2d8943abcae74d017565f6920ed30a
z41c789485e78a219247e959ae9be2e3f1cd1e9af5fe1166061c460e256a70999671e1f60e2c7e9
z84a97af03b1dfd973e26f4ecc6f62e341e8fb558e93d5ac5ea6872c8f35609543f2bc5b332ac4c
ze7e84277c084ae276bd96dfc13d2ec03348274acb8ed164a1ae785d380441a98a1b01c15ff0911
zcab84489832d6542e240c19a58d2c5019e620bf48181b6a2cb5a2d2bf1e3db6d17b40e0c761607
z8937eb604e716f9b47799fabd5bebbaec0ce2d149b2d5547cc020c7ec30024d0c21c7bdbae56d9
z3edd36728533563c24181cf918d44a9baa2f498e9432e15c968b3ff3468d9bd29a1c25c1c4651a
z5cff1676cfaa660a996fd9ab17a93d472c25fb3511b2fe8826e4d3c43e1ecf118a36f3114c2f04
z26d40b105a3d62531b5e2e83f594a61b6101361cbcb9a6269e2d2f124e5c515752e6bf20a05f6c
zf3e3e3583f458664f0fbfd604b1002d72d6dc976d78b0aba3b0c735e6f60724d99ffac89b8b874
zf17ea5fa4af1fab692b22b6626219d7d51d3bf9fef82ee6b60940d9b808b32697b5d9da5a9e509
zb98172ed7123ea1c2e58bbcb64d0f5b6b29522df51b6e7200c0189f94e0ba228f637281decaa7b
zfae84d3c8cb41492d252f87825bdb92c974477f400973f1177ed0cf69c726bb0cf14f4d09940f2
z738d82ad11f7a49c3cc67663cfa87bb7eae665c4bfcf3ec42fb49c2ff64f9d11ee0db18f0269c8
zcbaa71d830c3484343d9b07139cae9b22098c0e3680218b8e7295647ad8cebaffe8bc7796ea77b
z7b4a81701da8dfd6af08ad8d928f99b4c22dd09059832687aff00d4fa501fec231b9a25b43b09f
z4b692f6c1cd6f09272e0397f7b932aa95f56c40392335af05caffb7dfdb46d3b0f0850afec8cac
z2ea5ebe6b724463de85d1f4a8445a60dbfd2bb2b32e34f79f318664ae6863b4e44b8bfdbbd0d2b
z4472327280a786ba78656cdb0ed2f77229c49654860cc5e942eb8ab1892a36b675c0a93c02fcc4
z7f6d79f6d9e61b08ade3b91bdaebd4e3c1dbfcab29047d57d963b052e0979fd34d7684737b0aaa
z863c850557209f3f218694788b8f14ff570cfc802afbe2aac01c9435bd8ed2ce0ae0e392c9a7b9
z5493996d908266c8fced6e60e866bcd4e37ef0c2b941292e4b86ba76beba58f8463e71004d2105
z33964348a1daad191347d96e1d8dafce9b32654c97837303251b44daf33a0b249b6af3e4b62dcf
z58ba5bccb630c805547e6828f6d1b9cfa8df54af1585415c767de51e2cba822b788a0894e665c1
z84e68eb3ee3954419842365b1392c71f86dd2568545539890470a8daeb5fde995213ce5250c785
z4f8f65e47701b24110c9b29c5dfd93980fbbcfdc8986d9c357031e2eb9e795ae2710bf8a5526e8
z65055a50a67c363845d0fc4ebfa6eb9487f0b333082ee864340d46b2a800833df672ada8578f24
z857524c85e4835d3f55cc362bf0a414efab726165d693b0e437e74c82b18399a3fc7078dfecbb0
z29a48fc2ffbeb892dae405b5db24623e59020224bfb62a2ba29342375790673f1dbdc6c28bd7eb
z16a2244386835c6868f1b13c1af5eaee1c0ccd04bf3833beebf35c2d5bff2b76d3033b5889d0c4
z2b1e7d4eb13ffef29985cd0f4c55be764c7a18029d381bb2d58ed411b149ec019cccbdbada6126
z2f07faf7183dd871fa35f7b37a1728a363540efc341ee6b1fea3d1cb73facab41a6d00a6f36af7
zd37fab51fad458830c8cc7077af17a2ff388f5f348928d547edcee740eb1dbbe403cc33b9d4fbe
z22a001c80c795b62d841384ea3d2322cf6359ad57a705b2497b09ff15a03188a54bc6dcc89baef
z0c9523ff0dd1b90542299e9d29e20f7a25cc274ba5f362ae2fadba2c07d5d476a5e08800260ad8
z56e30813f9fdff1025e39217ea57d525caac3e9df1af70cbc97817b68dc61ca37eafb35994ba66
zbcd384616425bc4961dd3d0be7a85423e91f728bb085af6cfb464ec8da228458f2d0100231ba22
z848a4c6466bbab92b816ffd3d876dd23d9e215a39d53b9778c64702928856b713c2e6e28c236ba
z6f669659fc59dfe4d7283e3add335291d89056d08a6cd2d4907cd6d15e78fb492f0ff1c66eb785
z58ab1de9c325f4c5fa5c72a01252e321502214e03501ea9f4ce8fc85ddc500e6fd90338145f880
z6f6b7e43099c6795a11135c6a16f119df7f9a05f01f6c4b34b9697775d6d4bfe423fc09ef5c884
z064da127d0d75b56c5578dcdf5fbf0e54b17819f3ab8b30027ab0aa0226a2ef5d6b8127288d0ef
z182a08465396937dc60f3f7a78af6f1460580665b4a3ef3f10780b6b5b7e0a02a8afa9d868901c
zc89c94723001df240cd9c77394cb416948e3a66adf7a94c6c2ed328806c970edd10a9129a5b2f6
zca860be46b328cea58d1a5095560506ebb821860141b3272dd137589a096e9d7498a8750a8c229
z0ba8feae5143c361ccfd49291f06d28582a827235bcc7f13fbdb85dd1cbe523f44d66158434e58
za14ed9bdbea687276ec2f4bccd037200421a8491f669be400aad4d135472e24254bca19b427b7b
z74b80bb2061e28c995db5c7997cc3b67bd6d96417c74b0b87cd86b01d6cb55edcbd158cf301bcd
z2b0cc3dade2236555a9b4f5d9fe037808a12b1c0043ebde2fad7b16a09cd365008d10ca4beda95
z54a156824820bcf2e81ba79ce30e76dbf87b05b052f0499d868edb8078a5ea0d94de5f129a9cc1
z922ac9ea120e8e7fd9937a4a0856da358d969b9ed48d4e9553695437e3087329e00d873d36972c
z28c1f5cda7d1210d027c71fb859bf164049ef62768a7b45c496c90bf9e1698564de0c6f6e276da
zf0b1a9f2b9c68cdce6861b2e5a960ef6c67fa10e728870c20459b9906cc7279f0976ff55c86bda
z19e37422151b7ee886223629bce262b7db25f8a0951f8d06ce946dd89edbb9dbaccc65c75ef79d
z41a7ffa22c47e1e3514f5ab0d16677acad41840637dd79de539b2fb3c255aafc429a4e06605ee3
z057836bb6a69c200ed78e3de745a415de130232b2e308255ac78a58c0adbb7363cedaa56d75ad6
z471a7d32b38c398cc2e28370fd86a16338a901523e802cd25ab20e899190ba15154b98e8bb2d4b
z95d08806e56c3fda821596f3c1c1be7cd7b6904956cdfeba1c2c07dcd3703dd5b5ca948e71ef7b
zfe35b60195fda2da46ddb2164c942963b89c725dbbbd5a3c36d5c9192526b8c84437c16d2cf4dd
zc69f0f5cd88c4b9001bea91860aa523f32dc3414c2f2eee51eb628b470bc4a272c18a57ed453e2
z4d477cb49c6f90e62c95234f8191b410ffffe70c3b4107
`end_protected_0in
`else
`ifdef MODEL_TECH
`include "qvl_usb_2_0_utmi_logic.mti.svp"
`endif // MODEL_TECH
`endif // encrypted_0in
