`ifdef encrypted_0in
`protected_0in
ze74c34e226135848fe16db9ffd31815156fdcf5491ff70c3107000761e07383f2d117f272b520a
za48ae13031718d9a985bd19583c36208077cc8dc63aeffd55531981c41c4cd970589c21ccd8acf
z0de8a3793464ff56ad357b3d586e151ee48ac551aa2ee9df6efec420d2cc03817a64db22c7f362
z7143fad0c91180671b7851aef40147be22aaf8ad53772f5635f2d5c103a0905d8acadc54cf18f8
z66eb3f0f547c36147ac1f1262ba04e73bbbcc2e483469a8ebf419e16b597ff069b2101015ce3b9
z5b1c97e72a5d7f4612f06dfca0710d0eab09c9c98a36000584237358a2e41c49283b4e0823d1ad
z5fa29c0d6a646aa4a80751a35c296b990cc03e5b6611824708077dab2412d0a18ecf9336298816
z3b8a441752544e1424125add4c9ab9a217e837fdc8395575227965fa939daf8eaaeee3afef8cc5
z5fc55644dd4830b8ed3e46a60daa10ce721d35952baf74401afff81236406b03bd160ac1c957e3
z555a4f8f1ba36d8f79623eaeb8ca31e9d9c3a76335453149748525415c66ff209e4a3414f5d7a2
z4afc6a65dc72e80342550f85f819105788307d7a21aac0e07b5f6ea6b818c618826b48a823e61f
zadaea531ed040f62f1a7772fcae07bb8afdec9090343893c7500e7618e1a3701684c491062422b
z77f7b009a04f0a0015cbcdae72369c553956e0a388572339135e12fd997ac85872415539eab5d6
za83877dbaedc1a0e5f056f4d4c41536dfcda0b124012ef7e519fe52bb33a1247b5c3e92177ba17
zbb3bd8118c790cbac30f0ce36f03633c7b364783bffc53ab9ff6fa48605bfe01eab13396c73551
z4224185e91572a6842f8ad36da7aa81d96cadb9ddbfc02d20d0fc5ac11f6f7d031caec6f21c3ed
z698c19392fcc82fd4f5b1b0326b6465b6b79eecf41643e426c26d3b0b9b02a9ded3248c35200e3
z7bd526b6745760b8cfaba14f05fc5df18b70689648fef2617d7bfa210b66b3970e2c3e3ac9ec14
ze1c20ade7039280a0765cbbe956a9d05fd5448ba38d847f062dd3fcfd74344db6c07be450cadab
zc27582b13ba8d433e0eb0a75ea05c7d7196b7854ed120e8783eaec14347ce540b08e28f916daed
z1f66e0b15cd75e6c8404a3e4450fbee903318f6a1ab144a6699bbf0488568f73b509d2d105c5a1
zb55c1df59d26c0fccca9a5d14155b908d46a40c64c1977216831946edc8fa9301094a71fac9e8f
z4d0633319e00158b5c4101253695f68655ee3970eb1a57f660d2fa70550bd4b50d36bdc6bd7864
z452f2d400e5fdfe81d45a33823c6ad44f35fc0c6ef7891088612f048aa6de9496a56cbbc032da7
z667c5263c9604a15650f290b62f7f60326fcbd3480b71a96900e9dc681c3a0a346e0850b07a35e
ze261775c655ed8c9b3dd66701b1d1d01074815a9f96a67bcf8d8dbd1750fd4609e3731835b299b
z205ac123bea00e214b9f696b108e6563e1b25250e597267586922793fb3e0ca9ba8fac1878930e
z45469fcf93b6b4aec234f0186026953f41e8c69e3e642b821bf803e6726b24a01e2072fc7b0c44
zd09188083853a1e43b11c6058ca9ce76bd389aba9ca09b2310223abebcd5b27571fd05dcfe30c3
z8a4931b90d503b62140511fa4f00f5cb2e8cb3c8ff967c51737f91461334a691ede1af7d471f9f
z6b708c1d7804fd13c0aa0fc44eb4e85395571236c3d0087d4d6ddd8b4aeaa8ad7cbe3205dfeffd
ze22ffabe5b35b544b86365e28b7b7d82e159d1dc3e5ebb14b1dc7a72434c1de621464d9e15ce6d
zf6ec97982270497922ba385768c34f641aaf7e4da7b718f408b02344d312f8144c5403cb7bf196
z620e126401a2e58a57d347ae223660a5d09b18892b99e3dcab0d35ba72b8f2ee94fed5226ac4df
zeb0cb95e0a75c02abbc368e67282c6357f8f2655ec07cb59f60d551dc271176da4568316833e5a
ze802a542b8499fa93817408f50724a35e2e5552634e18418856757a171a861389bb94e8f3e1967
z4c6bfc8760e18c170e1eed7b78c7a19623adc48a4895cd54da0d6cd9d1aabcefd3e84bb693c381
zb52b91f35515d99410e882cb4a7144e4aeb490ab1e893588febbd256ba6c426afb6fe7f6d9517a
zb84ba9dd6990b892575bfc9fe689fc9bd0470d7c02fdf28fd9fe336b410636de13e73107bed257
z5cf9df7587f7cb982dfdebd2b59d85e67c21ad710d5b8f894daf0890604f46a4b7f905d0929084
zc3ee30bf544e42f14e30fd8538ca97b94c697003dcabae6515111e8d60275cee60c80e4dab9ce1
z8429fed08b4005a74078021a53af201701560b2b9fb38a13bf89691329d325aa8abf3990b95348
z21e2d554407e6deffdb87e0265526cf3c2b5bad82f6d3d34734dc6467f4676d1e74c9d94bcd730
zc1f79484320e302ce91cd8327e06df89913395cdd3edc790f3753b4666231dbaba893da2c84490
ze315c7c40559354a8f1a95c969662bb1fd9faf6c087281e1f2366d2eb0df814192df109dce7e9b
zac7d55788fd366e385a90028bff09cfee6318853ed87baa2b72efd80e0c483233012c8b03b7971
z6324adee0553bd8801e91c09848f34080a318145d257648faa7febd7de6703a6283f336def3ed6
zc94b46148e90c1546e610ba3d84c57741f92f894ea083f29b6745bab24df67995829d63233b2cd
zdcc25d698f1dce97910000578784c0f48a371e2c442158ae1412f449ead58069a1a950c1f7bb2b
zab5378f7fd12f6e59b051c5539e6c091df48e0c0913871b9626babd06f77be9e1967126d7f1f96
zb95c481f5aab1d8f7a160c1b8ac871a38a6018e1972d10050ceda1fc24836d6cfe0c96be1a579c
z45c8071163e773519528c46e4b6853a0cc293829a90f5924847143c41a3bbf146bd331eae715b8
z77fd24fde80ea5702a15c88a1ac106628507eb8fd9912613a048087b2a572eb674de04b686adad
ze014889a56e7586a58fe5aa23187a1a0b01285473e9f1691150178047969a4f8828473ab14d6f4
z8a56dcaa6eaea4da2ce6e49ec81a5a8f981e4efe012d95aed629d397928938847283bdbff85de8
z2e62c4d4cb6f9b3634dd8bda84e33a16e0ead3722a85e648eab604a9cfd5e41c785604b46159b2
z7685742a77ff898fbf1ed40894cbd55bd4b64338478d5329096639688492868ceb235135a46c15
z189ec7afdd04822c631390202a2b2a686d73073a4be8b1458ef863025b7e1c3e8da0ab27efe123
za4966f9339bab63b0ae8e82bafd19a087887e685718eeb46684bbfed6b07e5cfa25359b2b0a3a9
zb40dfe29d4cbe7a0f952b7586ab59a5f08e2101f9ef578879c7e495fc852ffb2ad7dbc19492a62
z45fab0b89d3b5630bee0fcf7d6603987b729ad0b8b53c5254311ee62f27fc16e03dc681463203c
z30b074fa2327d45fb1ff54031dba9d6c70b57e694dc63004c43d73a55b3b6eed06e81028979b08
z942255e5d90d6550ab40d51fb2717413f03bbefbf2ece5781441d0ab7e54365cf9f2ce0497cff0
z15a41f257159c801083b0ff1ed7c6fa3413a40efa342c0927da92f551b8d596f03a6c68829ed7c
z5a730e7781e5af816fe0e99d50ba136fe85464de3433f9167e3e6a1fd5c3dd2a0af797b4efcd21
z542b6e6b4f5de782e9ed79be0e85aaba8ce2b480928d56be79b02b09d22c472ff4e9e783171a85
z5302186cc00607f299e4e56c564911022c18fe2d5e0480bc879340f17f072b3f5df778ebaadd17
z925b8aa5920442085dda097f64960ad5d881841697a02b16c7deeb72844d9711416f618d5e07b1
zed32b5514e5d0ae7d23e11807f26b0e0b99505d687306a82cfbb379a5b9bfe1637d72bec1ff69a
z613fac20374fbb7414c13e19efb406ac00f638507f953bea09230ec517ff178ca6d0db991c1f66
z70434441bdb0969bc7f5214a3848a52afd87fef9aa2b4890b77cbf771b4ca29413624f6928898c
z5f808818e1d2bb43993632c798a1d1e99a2a9c221460b59f80626c3bda5cadbe8705a94cc5f440
z1c39cb200aa559f6db35f5413b97be38f81ee931b4151e74dfa4f1aceb023bb0b859dc7788e143
z778a7ce4eec4b51ad6773e2f4ad61928e0c73dc6bdc0f0b7432179c225b285374ca7bc8bc1f1e8
z362b8d2f67e69cca11f3baa05210733bd4b6121c6dca44dc90d7eb82c1b23fb04948bb0b415fad
z13f4c38e29df0f8a03b66bc0fc03ab502253760995d5750797724a761ad8dd3c868eaccc3070a2
z0e838673a167392f3bdb6bf1cc9ca39fee501bd94805d7a2c5026a304409b89b323e5d78734c47
zc531a1c671946e2abffc063eba78fe780b422a55251133b0736eb25f52071b8af1c3f6d1d63ff6
zaad29030f6af7b755fc8ff7f9b39aceb207af0d152f6ac96900a1a500c8fb331faebb059692698
z7fa08f6edab3b1aa94e62efe69ce5f6b8d27edf6fe0e9e73b1bf3f5b2839ce7e087fdd0cfceb9a
z420c6d268a86d08556aee459483e60c0ab65515f77d61e70ef049f586aa5d2e2168d34bf4f745b
z7d1e8d1be72056e077b65dc4579506d42d9b68ab3be733c75f34796aef75faf4378f545b5e8c45
z99b44408f29b6063828774d9a7005d85ce192fde220af3b8315b5f5d8a1d5d5b0b010766a066b1
zbfe555274dde4b4288abd8c3c4afe83fbc9b31e658c81805f6c6a76d2488bf01bb076c27904e6a
z8f2e3c54acd12940f2a782891512ef1173b1534bb2d636e989c0f5c0585059b2b13cca65437854
z5cfc49e0ad2d5b0452dfaa7526810d4144b70e48241f08dfa682a1b7224b1a409706673dc4a4dd
z9fcb0e3021f8db65cf207a5f99e8375258ba498f127714d6e705ccfc26b719e7631dbb3d0413d2
z673b38d6b33d18e786c172f061114cb2063c1faddf232f2a048f0ae973d88d4ec048950665d29e
z236d367381a3307c4960c89c503929c3b336606c7adc9017cca1cd8265f8f0a7dc2e2a8e2be88f
ze9e0542e393cc937eab89ee5be1e80fc839c28dc9fba459cf1fc96503ecfc81c081ebb307eb764
z84c7a1583fab9dc54fc1f511052f1f0243853ae374552383652d558b774648f61431e686cdacca
zc42b320773b2c699f8682a845984dfdfac77da82fd5c2dbd07ad1fe4e8012576f4cda16455021d
z21ba7ab4f56484747379192680660ead03ba34980c9129acc875df04ad61c2d32770d820ae5277
zd2ea50f2b7efcc964fe52b833d04066c6fb778e4aeb4cea68cfcc84882f9eae3842c98c2de864d
z73c51b593c90c9bfeccf3c0a367ec08323beafebe1d1f57656909ac53ecebad713e60e1a479fd6
zae63a6212776fcc62b44537b1a41922ba58c898ed4619d9dd2cca9957cf15866ac6a905283dc0c
z8c5ba749910bb470ee31dc57c93bbf10198d77886a313f88a363c86fef268479ad8b3b8274aba1
z4f903e77c3e7c7b88990a6b9d7dda25825f5f1be1b49309b7a14832d1ac19e8b74818523fac1e3
zebf042b9962eb116e8e44d0ea62df9862bc2ce5dfcd9b1b39f03bd604b65154ea8d84ec8158f71
z11485c57c3088cd602560aa6eae04104fa152b3b00f941502f094ba407cf60103275567f616013
ze6cf5f23cffe7314ccd1f0fb1dff49d0d0e5915a9920ca33460ab24a4dca5cfcf9aa956f8c6c24
z0907f0236c26a9b9b8befdd0f2b709b7b5edead47a3cd60f8f6d06362cdf3b25682ae530ec081f
z6411ae48be1579feb91fbce4c7e53c1d60ff03176a86a1cc3bb6bd3d862c1c17cfa7dc5cf52295
z40cbc0ac2969abda5eb528f122611c776d9384c5c27cda4693a22b1e7589814f16214abb8a3436
zeb1948f172991d1b3644babe1d40b9140a179078aef7c65e7de3b007b2d6c812729f627f246e07
z9d53b3fd1f7edc571d40a028de1b1708b6cafc757a591e9201d4aa65ce147a592efab1d00ec12e
z782fb874ad764292f1392c374610ef974eec896fcf34b495e151e7c8664a1aba508d0c3b25d3cc
z2b8f26f38dd23ce372a8d39624bab08dc46f29a7e12585e1ebc945e8bee020dcd40e1728672c4c
zaf4ed8cbb6d38170f5080ec84e269f31ae71e5e45eade4d86e055558b4db77c74aee04a7600451
ze0842d734750b1a7723459b3dad49040382097babe586c9a06abcafd764287e9b5ebdfb09beac5
zaabdb4958828e9ad948998b093a6872d2ecc15bb711646bc88383b5363d9e2979909f8d5f28ab9
z84c1c1363e6e98d7dbdd00b98c19014bbea25c8add5b4c45c392258797255c2e7fdbfe913789bc
zbd5d06fc6396ffe81ad33aa0fd1bee21a09a693df268750a3b4659c24012c17e317ab5deed80b3
z1e0e732d0bc1c0eb66b798b090639dd2fdc76c2b17702dcd71ecc483d3c639416d52929d642f35
z3dcc2a917205f7249ea83ee8a1ba3ad19bb206d673dc512665ddff950a5bc2f8b1dac46510048d
z04d202565386c427908891b6c514f239cd08f89c25e7d3ba7aac61fcdda3b14728d8dd22168828
z8352e4e1b3dd79480ec8aff65b7e531a48e6d0bb2e0ae2b94288fe06e26e0feaeb33e59f04defa
z5090918c65cefe86f69704a43b7023d778a2553a119340fd7938037622bf1c9c1293cdee17ad07
z81c11d89f934e6a1177c51da309b186595804c76530a79fa7f18bb79cc0f2af6d2581c7c042aa1
z5fb6f10cef2fc59371664fbc3b4f3512296879221131ce363480c0ce6ecad42fc9df6f58f2679f
z9c87d525b613c8af5e247dfc5022202b5caacd4fc5682d54570b3987b9f2c88eef606b42a17e99
z7453128bef0838bb24d4edd38c7e02b35e5f86bfccd82701986b66e6181e95409ab71804faeaa5
z0f77bd773e159908b59bbe6cf7334ffe4e2d4f320019d40b6f5c51e8b837c19652963744962166
z4c397650b10f8a295e7f0087850447c832d9bb6ac80aa9e0ba6a968d9b4ee74aa1fa93d2405bfd
z1d70e383eaf82176c280a108e624104deb962f12a894e033507d2965d1686f248526caed686086
zf0b4dfcd1f9d57b32f9b1319c82baa7c52e086e6d2f0d3ded944f0fca75bd0602aa303ea10f0f6
za892dbb60b0b7479013655104dbe6557feaea6e604050dd9a4b1bd5069ce88e4c71ffe188dd32e
zad014a352a08066b6ab78df7ee64d294aefa848bf5617a250042791ffc41a72f3382f3f465dd21
z3f05d11e29989715fe9609a4515f433832a85a00848165f2cbcdfd89ba785f82dde58e291eaa96
zf39ad84c7251b7b1ca04bcce245f02de6516331beadf34a03d48fb1069254337fe9d0937d95fa8
z65c6c2a7143c1aef7ccba81df606f86588a026e49b912f09c03fbd84c0331041d2f19caea75144
zb2583b004c0695ae9127c997f0bf787e1bd4d49e44f05c0cf070dfae2c87d57743f8fe3de8417b
z1e51df8a77fa23d55d4b0492e9aa1576fd1cafa63d703af077c6cb11e5ff3a696a924b7cbb42d3
z61b9487c9dfe8946a9548bfd132fae5e6290ede228545a18f27f2cc3b8ea477d25552c2a37a29d
zd9f7b9f96f0d049939658379ffe9281eb17f1560538bbfbf3b671eee2947584831f92de46e7877
zf9f290d0469a8112cc27454a34fb7ba1c6e3364606f89a5a5955f4a97439defa4aa62de3645567
z6e64f380710c7a93ab44152b7e4270e7ded208ed9aa6227da5307b5e4264c198880fc243975042
zf646698de1089d52c496d68401720f266cced4a3fb3880e69da1ba88e64f7f0718280f5666acf8
zc23ccae6bc39c251832ef4200feb43dbcfe34768682328c46d8cf05d6d51868938404ead3691fe
z4ef09b20c01157defdcd9f0c58ea3631253972668c3312ef96ad09cb138a09a3014a6b0ed0982d
zb931e903cc879d8bd4d7698808c410b4a6d159e6d7686e62da10d499011adfb5302ac293e974fc
z67f506dc1f706b675800b41a825aad4a310491b7f0511c63b6b7c4b7276112bcd08410fb7ebbc2
zeb6527feb81299d2d454ab9d440d152ffa55215adbf90041c91762b39bda53b684831ac3e2184a
z149c8d51774da6ac2a587c9a8ac706f85704cfba161a53745d969d449bd15398a30df0282db3f4
zde6fa20aca0304e3844477bc12447f51e39cd302141036725e1c40f7d5f419a49bdd40e1bbc331
z50579aa24b6ceedb4c33bf00b48707c6bfe2767ed299d0cdf58581320bf9e66a0349a30fcc0594
z7b54e383f9d239c5a47eb988a3113e44f7b344e149cd4bec818281ec7de0e683971882546ca172
z00c8dbf92a0aebc9b46958f06e89b8a63c789a4ebd2f13acd2c81871e50c4b3242d4fc8acd2bc7
zc68e5f05f12e1c3eafbf3a1999773c883fffc9e540ebd06dd943b7e745bb9e4c623928e40acc41
zf3c05209d167e71e93f4dbf211db189a847d3f441601389567daf0341a12a7e5ffc49450bb6498
z9e96d2479cd14f1fbaf1f1acaff73319f6b78d30633ba445422a1b8b2c38fb0207b6e27528cb08
z84d6ead43aeb19c3398aa8ed95caef3fb23230670f40505f3ac993f54450236763c3e3c2b8739b
z50aaffd6a926772d395e704c10658b854951e622425d2dafb28ffcae72c4e509130de035a0cf89
z35f83232ce199a67b5201558f871064916e492c15aa29622bf9cb05352e1822983fcd89c7393d9
zcbd12ee52c40837d221dffadf8c74f3aa38bc6e166c7d734b3bbd35d648dc27493ac69314428e2
z65667b8906bc9f9aed179fb67e9060138c5f1d28de4922a2212e4f438c4b585f0f3b1359e053f3
z0ce6f678c124cc3dc69de5d62078dd87fd7f64c8cdaada9b84563867ddd962f5deeecf788297c2
z348193c740c404382b5676cf22356ea9af4761e4b9460fcbd0ea18a83828bc5d70daa6dd120ffe
z3eda1853e0a1cb5ff91135cff163235a49cc236cad0fefdc0b2db2503a0258afcd5ec917eceaff
zd6dd47e6d7093fe8024c0b5c98b842488c1fe3fb34dc73c035a830577d64113212498d7b65e8b3
z99db9dab9c33300c61d23dc13da29b637679eee835e87eb61d7ce1c544fb2fd326f1fad558197b
ze1c9e424142409debbb3c55b86d05aaa7b1d777a8492071b64ab6d15008c8854938b493d04c116
z831b31673edb04ef74b53d3c6aec6cfcfec8f9c98423ca6b177e7aceb393df0a06d6bbb9e6a3b1
z4e347ed29b541049708d1f4735ecee75b5eb8153b9a9ffdf9e1e5123dcaecb3556c1bd287ba5b3
z10ae8e776b9bf5b6b424ba5e8bdb0ce2600638b4d5f96617531eb3ed8f3cea7e32c25ea3b943e6
zfc6ae89ada286c2c4b74aaffb136c4518f765625fcc39703b8e2ca8e79e9e128812387b6d5bf4c
z790dd292fba2500cbb8d7a62ab02aa5e0068f95e0cd6bd11964e07c23cbf3510bdb175079dd44b
z9d3f92c9ef7efa3df2ed4f0caa894addbf873b39447d46741010509e596f8a69a29e807e501a89
za00706ab578e64cb58fcea6dfafba1976c76198f11c64292e8887eff5fef0268fd9b966dbbef80
zaf7d700fe9cbb50f14957413adcc5309f90dfd29f58be3ddbc99b1ce4e01d1b24e0999ac5e57cd
z696bfa1df4de2fcb3905aef2de20e6449951db5afc880e001eb7f1ff860e2d557b876e1eb2937e
z62e478baf647165328112c31f382b9fb525286a8f89081e4a1ca4a26e038111500c44423a2a259
zc92dce480708299c9ff8737b405dcd84755900383b508f53736399bf864d6d0062715b847eb98d
z7d6e29a63c217a21b248106debcd13be4c825d7316d6e52993c317c24c4b3c9eb5e9e04fde6b44
z79a172d2f8d2ef89968af9ad5793b7c6782fc74e16edccfcc49bacdb52ba5d746f36acd17f7bbe
zd80c6ead3e20cd008bd0c72e43275ed1416ec4d6f182a3528472ac09d9e9f73d8fb3da670e4403
zd1c054e177e3c3b870701d3536c7a9e5c339d914e142e91e2ce50ca08b3a6a79c8fbba1047ca5f
z9ceba91627574528f986bbd82b3e8e9c61a974bd6608e04113a7d3711d2e41ff4eb387324ceabe
z51a81f1cb39c984cc6796d14a92b2b3eab6af9c23a0e6a04b077887504e4248466c96c8f12e4a8
zdc8bfe4efcb167c159b6bfb3238bd4a48e8bb2993655a64e8650915b3b118913eb8e7dd5d61599
zb1cb2815f7abca43ebb70b838141cb3eee8a922d0c99f3d3dc8825b4bc761687ffc2aa358da8de
z32a338106b5fba5c2283e91eecbded725ffd9ec4dc92720011080d62a4bb513cc8b6bc105946ac
z0af41a971fb4ef444952f3905deb4efb30a835dd878e656717a141768ea236da205e61413a443e
z91d675883854dcb324291dc3fa78ee9ab5d4b01274bbc2f6f214b39f6491b83e77df38ef00a60d
z34e5c4163777ade5cc482943999d9dc29cb78f9108ef32400b6b744f9bca602948d2bf0300bc73
z896c17da89b9aba6b35b531583bbdf051b61692670fd9f82edf300a058daa426e987298cef565f
z0725df44bc713b69387a05567662a53900c06f987384e69687d9ec501576a98f2202f73d46b14e
z1017cf1ae6fcddc6e90b4a260ab3c9185fc8cae9e58892bcc2e4b3b11794f0fc1b73bb58e055a1
zc15abe57a1c5928b3b178607bf578196b2b964ba498bf592227e7ae7c2548132b7d29a1611868c
z27b9fcba5d71cc58689a366dfe8a757953c714d168e3e20bc73caea547d71785af5b834275899e
z803dc669ff167c3b2eb620d7e23d5272e5d947fa2900f9740b581b6f561e5bbc5f75da6dab5620
zab5dd0c05f2db1d9f7c688c013fb7d06946876e79a61614fdd1d1304432159f49e5204c9805ddc
z10b6bf85fb2553b3a17dece93d4bb62cdb3481d3a1b03bd2744b6cc57d90d169ce63890ff961ba
zf96239407fb22f6dabf2e184361c1e229d51817de0110ee7fa809486765c20f466fd40ecb1e926
z6e9fa5c9c74b4d5d23d586a43dfc89e2142579a15ffe41ca55b31acc1e581d05e8c09f01b3f04e
zb7bc711f21f259b60ee3ad8db5adfada119d53cb4dda8830330bb92832f0cc5cb4ac6f9462fc4e
zad1afcef424f9230e1fa7237c13c3ebbd1e8d04ceb77f2490c0aad83445034eed41972449c5d29
z8e18b206bf891e332816301469d4ccad479a8383f0c2e792975a41a33d47441831280d2257ada0
zef694194a9b83a8f8426e52c364348a03bb189960d2d201176843d0af061c6513d8b1438aa9658
z9ade920a1c26d6151ce05bb3ec50dded8b38e637f6ab00855b17257b3acae5ece2f7798293a5b1
z162cd45ea69241d373d980e3300664a5974d79047c57d3f7c684ab08c3118a040e8ef3dfaf021d
z55ec94489e7d6979de64adda1f50f2e9387c16c24311c042d22f2c32876fefe619c21a5e8e7700
z215c03a7ee10d231b13a8efa29e127467fb9c4620c4eb5a26ff9e4871314356689c1a4d1ebf9ab
z3a43afc2f6e7d409c8ffa961a4d9a5b2c076a9f2e058fa4f5096e3c1b80024afa869e24010a2f8
z946f444ae0966223dbeb9dee356f7b8ae23f6b70015c2a2c1f7c55e109d739cdb2b2b96b2f5c50
zd3a143d23ddfe6b265dcae69508b62a223a83ef50ef1b941a62e50479a2b608fa72757b410e65b
z6f0d250d7cbb7e6280807284c121fb478225bc584d4a1f4ba7d39641c7dcf25919e930138cc600
z41d6bbf7e0cd5bb3394c5ba41cbd96057ba1281fa301337aa99bc5e433bb562781b404eb2920a2
za66be152e77c06562bd5346c1542e294443c5df7337c95953d158595ed9a7202aa57d66a9d0912
z1a126b46c3a47006a1d9dc23072fe09a854f0f5be2b908081b57ce59550699f1842e42ad1706f7
zde03852fae549c2640f3a779503a68a37fecd5a0f3edb2d4184990e229d7cd839dc60f8bf385c2
z0fba06d134455b7d9f9e7e4dd6ba506c21dae14c1c3539842769c45b2d4dd3215b328c60c8cdbc
zdea16d5e7bb599ce4c50efac518b600d813070c424d867daa90d5b9f595813ee41ab14670aa332
zb50faec7af335adf879f684976e33cdb361fa009e1c6ff325ba4465b9fd4e3df14239d28481363
z239817bfb2fe4994233d2ef967f0bd38b2ce3755879349c239139a33cd0f61ad0bc162dd47edd6
z1a47f1b7d6269391437b2406f322b710c24c78c91876b930ab58a8e49fbc4dd25f28f70b141c47
z50453e67c523126c99a35b23a4328a7888a312e6ec532c2c2770e133a5823df3b1dc1f23efc7b0
zcae77fa954dc772e73cb1086d6d9c8fb87b1320af64f0e8c3d50a3529100a63eccfc58fd796a79
zb410f177de7a0765745ff145bb431ebdb143158b564222bff9e3d854efa763db72ceb95dadaa13
za1ea3c0df0c494eab0bad8d1bf30785bb9cf2182bb0f2cf90315e5e10cf32fa4d13e3ae6411b9f
z8d28addc3a89c93c18b11a5619a55af37fe576dbce26cfbf24c9c68a2fee770f910d4839001ca7
z74422a811e3b69ec20ffccc9403c43f36df05dc32aac8d429f94dd8d711e20c9a6c34da8ef76b9
z8ff3b8fb5a1697a28617c78e5a33986dcc1d826ac132163ead573dac0856612c8626bc0e94826f
z259929dcc74faa522a5e8466c1093f799cb8407c923d45161df78598f47910fcc5171e9bfc612c
zf8809ce9ae6ccbf69db61bd23a96b6ea2ece448f02e7d3978a13bb519bd8edfa5b5b6678a9acd3
z991627815a7d988fb743ad0a4a12c562f972d195cfd5a66098a8e92b4f0012fb90fb6e5c4d9ef3
z1c9f299228fd5ab9cd2bb989fc2475c4abeed8c05de6de0feb97c310130efee8859ea70db60636
z7e9e2c914e8ed166fec0bb6c7262d3e201e38fe1856af59d3a525906e4f9edc890dbe041e8f980
z4b1eab3ec472b2d60accc27695fb5db0a7765ad9909156dc4dd2486c15e0fe7737123d0610d92f
zcdff3433b58983144289da198355240753b493106ef45178cdee3df535785d1d6132fa4172cccd
z849113f26d41366ffa45db9601706d1709076db61f0ebf8f2b1c2e50899aa613dc56c948faaf2f
z1edaa05cfc7471d3d3c82d9305ac99a898f9c601a9cb63d126ea4e52d60e9deab071ccbb131ae7
z0d141904d51a18dfdeb3d72fc15971b690f2eb9aa3eaa5a2278428387835639a7edf2ecfac2dfc
z8005c21b6209a52c4dee192aed2cbb2a755cebdf8d5253e7ed580c8ae7b11a30f42c46841aad2a
zfae4fd862bb2842d14f109a3acc26cd8ef089270627bcf14bbca856a5b92800a92c5bf69d77391
zf20b3ad07fbaf839edefe694cca9f4e60653f40d6c39cf7dd53e418aeb0fc4082d82c9b69b56cc
ze5f20a9b2ab0df986241292820e5c35e5ae8dcbe085afa23a03f14a99ff039f5d9777c71ee51f3
z936b59cef868eb80081f94fee04c7026e98f1a80c407a84878521583cd44ce23021821c5be9327
z2d37f1524c805c736eb5de35186774a72650a25ed700979e0e0c74bdaa04d6c44a7fa2e789ad6b
zc4b6b8464099dd8373410a189f42d0995c97c21cd14d5adad09e58aca5a03a6f7a170cc38c26b4
z9399e0e227cfa9a12161154e2ca1691816be44eeb658db6d7d978452c46789fd65109995640ff2
ze74b89250460a2a8d288fa2d6f599fe9f8242b0f49c367c1646f49a9fba8e391839939060cd63b
zab40e3b018e70fb1769b4fdd4ec77991fda51fb4829c72487cfa1e8e0c50c684c42a35aabacbcf
za58d3ebf0015f86bf9659ccc5112724661d188f78fe2054a762877b7eaafd2d9a04daaf1a353da
za41de730112db329fb9eae580509eb8facf8e26cdc1b05b9ca33f5f8d907483b100a56ca435ea4
zf128b5c00adfe7d2a7390cc6dc9cd7cf2a5fb16824d202b2c0a3e14d655738a1664f21de833137
z0aded8dcc930fc3fca0804f148e343c4380f58918706d018e4b02a2c8d4b4d5bfb08697205a899
z0532aed113bab57c67c225a116395fc4c8811a9351a6bdc0110f5ad8230f96f6a8b75696bd3a14
z42481b1dcc9248700482b6f6915253268e2ba8223e2e67fb4bdf81d5cc7d19a84a1824de47b06e
z6bca62acb05087d3495ba74620ac684f3f03bc9cec7eff2e0cb9649cf3ad6f7f5567add857a030
z8db924906b750d943b7abfa7d16d9bef8abe6f787c465001cba835b2575f321c4561bfb141d4b9
zd40de1511292f07643be5419c7cd884a93d7b3831878c7f0fb19a9f1403c6236c5c06eb7eadbd7
zfbd6993f8b9f34f10cc1aa619cf7cda24633cee1650d95d3c0fc4d7e0debdd0cdaa64430e69f4c
z1c1c155979764eb7b510a136ea051f2f509cb5f0102d6a5b6649713a95ad40b6cd3cd223a3fe35
z1d53cee1988c27a625141a00d3d03e71c263a3e0814c445bbeac5915ee46b46427adf593743409
z15542817ca857a57e5068b966eb68d8bf68c4ab049d338f51fc3ebeda6e8a15fc2a5fb6ea7883b
z24a8a87185b5512db460ddf6a3143c8a0c90937a2307a0f59e9c013a2fe6bebf70cb0d20c45456
z16d9231fe098261abc2f1054757fc1177e18dc1372c24118b32a33db7d37f0ecb99526c0a77539
zb7ad8589b21617a809507ef8eaeb63f006e39e67660878407edbd69ce8d9ae81cd89c0b3b5401e
z1703575bdaefe19cf74ed1979058851139d41b3a56441c574b6bc809e21233c3ef4024e8ef924e
zfc6c5782a564f3e2fcafdba082cc25938b72e17116a615ff9b42663045f6dd26790bcc6c58d11b
ze969355460b241229f9eb68b407f5d27b180aae34b45355f0403b3e12b43ff39b93753a8295075
z9812cd79585c371313ee30311dabe74ef8a98a94b4319a2b50e630df12562205a9ab2271a54b66
z169040928aefa741657d37ce6933932cf544abd09c070b5ec93d6e4903f1e8770c03fadaa0b42a
z8569a84e53318b61472d4a58d363e2775ce53bf78e71868ad661d8792c7d336008aaf5893aa658
z9a0c061bf07de1bd023b19e31fdeaffdda1b1f12028c1b038a239bf52d35c1fa21b12a23dd7b11
zd81bfbec659ec583a6a1de1aa95bc59c8d0fb31d678f09cb063c7bea7cdd1d45d8a41921ee59ac
z25a5dc69d36702d53c31c34fbdc3e877f09fa79f9495384c859dbd263086b26530137fc3e087da
z22b87f6ed8dcb043f3048b5df8cee21bf39ad910c17696dc88bf4305ff0f197a86ac97460c7790
z75718949d9824de96625173f83e99b04c188bc637292782cf3e2565323f88e9497a1b5f4f0b296
zdebcdc450d8c0fc6373f90615cf80743dc356e19edb4355964d7b806f1541694223780cd27bb7c
zdd084bbab72e5494fe6560ceb3f1da9bdc5288f155fa20c355ed997cb89a25fdf546ae01acca85
zde19abcce118e9831b94042c8f4b63def0e9e20eb8429e894b2b75d2f2bec4cb835835c6d37a09
z97aea712283b126afa4a1ca3038351595409cd83c4d7eb87a67e7002f1bb94b3ce32b300f392b2
z8c1fc2bbc433d48631c2ff654580ec0bec04d0350bef0dab70634b58b62626428c261710d914d3
za72783b0eab5d50959dbc225374ddccb14eca15ea4fe1e64e0b203b2cfaf5bcc5b87001a0e1289
za85320b3d851eb5c68acf77def8cf71679e6d6359bfcc1e2ece11a2864aaee41ea4360aee25560
z05ed818c83b49700c32dc387394c36c25b46715be573a22274a60e3cdec57ebe1040a632ea36be
za594a317c21b9f0a6c4d516b46c9e24e896249b101c767882e3d021c55f2ea9cfbfe9f4da79b64
z123a6d792a84fcbd4e27c58c2865effc8955e21a9735e0d877d5dcb3c0783621e00e4887ad684d
zc8011dc641eb2f87d5f4114b7f200d23a5c8128fdbe257195fd62e9cc35a3c66175c9b2931b8cd
z578c7b3a6dc1ba33624264fd4d803359e3e66c28fdcc9c6880409e9cf7035eaf87673f900611aa
z2675999516bf0ebe8946de3bef2b6bb4b8b6cbb2aea059e8817818a11e615a895b03d361dfe28c
z32c731b4b4f98055a35b3783b7066665a4d35e031ef9ff0a66c7dd70a963af77cf680542611a89
z7d32430e0191393bbc563d5dd18e84b87176e1385f4ee5afeb2bfc3fa78285dfac877af122f839
z716353d4654a902750db38199d393e3db750a64ef7a9336a6694296084071b75a051e8fba6fa92
z508390d08613a73be7e9ee258f70739ae6592723caf00671db275154a0db64f3355c14db6ab757
zac8842f7b9ab951d7bd717c01b98bb7e04ace0fcdff5c75a17736f8620bc492b02e0e7f14abcdf
z8840c2882bdb4fc33488d0b1e482400f185a911c3494b99cbc69d38bea409a519193bd93d488a4
zba8b8b275518d87557e8866151364ad0f18c36954dd30bec90b269371357b09de988b1811b3ba3
z755dc669514f9e76411207d7fe0ab56c1e41bce7b67bced30f023fcb345f2c60acdcfe59f7f153
z25c7eea50c3dd9802fbf7f42e40d50d92f4f3e859993d398f52b530c3efaf2fda0b738bebc7975
z06cf961261fd00f75fa87a7637e00c257250bc29479efcff0d41859c4847c13ea3f80615fcd5b1
ze0520b060a9dbc132eb43d297c06e46f2782aa652e3d294b13d146202fd2e4ae46ec280e4902b9
z9107a42cd73f505c376cd59b7edad7c86e7190b87ae3e3452c78217c407fa5e5bf8c595d43da7c
zddc6aa6b881d70b7a6d16289e2ae4541d64867c6a280ca0d65d2495e64ee10428533992110e8c5
z7b54e51d8f660218522341cbc22472eff443873a3c2d5890aa8aff30b9acd87260bf0ca584cac9
z98bc83cd5d3c7dadbf0b0afdc2dd718d752b6fce5cc23cee209ea17fcb2ac047d197c5cbeb6d68
zb11aef929aa581975bcf4eff99cb52929737e51c20596433f7f79bb84092e882d111b9bf7ee8f3
zdca41e16559fe11c3537b6eb90ee52b400e0bc892f6d8ff33f19db6ced8529507a644f1caf7beb
z743657c8d8e307df3c8dbaac6eb69bd5964519fef00e9e0f18df099d0c3be959ccbaf2574bc270
z96264b913bdb646b8461906a624449e060b72ee3be6e69f8c9e944189d269f77b018339e624f32
zfba9b5cbe133cfac9ea36fe0494bbf0d1c97e9e100dfa2d7b21b63b2d0cea6112649dd45acb3aa
z2963ce8db4fba8dc0769be749ed9a41a6cc8a4153c60f7b26fdec9645ba9fb3f6100eec67d2217
zc9b9daa8c0edf8a5c9820c2d9f372c8aa6aba8e97799ecbebc01eea60c76fc787475b42edbb6d5
z8bcb564442ded1ecfa332e6a86e5f8b7879c536646d8f8fc6995e7214edb14978ffb59c5b3bf3a
z174d6fa676eb2ac9cfa0d6e9170c80328f01c73d95b397946263ea72837b11b3a7576ce7c6ef5e
z095d8ca51eec473e76c4e652dadff710b43dd250931f319b46e14b1180244b0766479fe0b02213
z65d6b91e2f9051cdcaaedca28c14fe1d3522b3064eb5db6cc435a2255dd3ed857281d36770296d
z9da44b51e5db46231b2f678426c65a2f082226243a479c5aae6cc3d7fe11a9f842fba401438e2a
z0a884f654cbbc488a9fe3ae5723df48f51f027e6b0dc8290d5d3b0a46e8feebac682670a8416fd
ze675a24ed7a184a3c4601cfc1e5b047a843102e60e7bc9bfe5030bdbfc9dbc8d437e2bf4198bff
za70f2f791cb20a15f8206b6d145922640940f0eab59be83482d02a2853d394ec64a61b37b275e7
z20ca50d6f0bffbdafde3a68dc8bf2ebaabc8de7ce838771febbe3119e97b9af72cc13a55bf7bd6
z05adb270ec6e76cc63a16df92eed82f8a2e039b8b71f69923c2b9d9dad2dea9fa98306b4315c0a
z6c41c46cc96d50deaf741fafff24ca65b7e020a2886beb5a5387c41f649a030689eb9c433a8394
zf60b3c7bedce640a65b6227aa0f1c1a9642c00fb8f1184bb90e9591f872bfdffb4e618cdf94fd3
z3ef9907801e0c17cdb4a0a371282e588f7754cef0d46692ceb6afe111feda6bfc167a8a8801dcd
zaa11dfd0028073e483a371b5da98856703bb63eaa3b4d8d3b41c5f66c4ccf835f1b1076f27d7d4
z0da77e14b16544739c46724ba78a04a48c5f5bdbadb32ee23d13316df3402c97cb06bf0b58fb80
za624ec31e68e2a668fa1bd7a6ded83a66b16c99056c322f8e4fe4a0c9de75dd6323e42093387a0
z48b941217ea50787d5b5997cbe849f0c8db35220ffd5464c0447753c0e68c23655359ecc064812
z0dc310a7559cec0451dc1b2499592040f8d258c449915b358a9ba7cc10341bdd781e795639112d
ze3ea9cf06a160ae2e697ae123f0554a6fde2a7816d13728ef44669c1b6f0dd875f2a57eb3375df
z8fe8d509675a19a863a47dd56433f2728aede42e6484e33cd415c9675d41b91b19cc75e7b70ff6
zca2ffa68594ad9f32718e7d709a71812ddaca6476b7beab41a1e08aff590ed9dbe2aa5e36e4bbe
z81e90b388e6db4b64e88edfba367ae0440f65fd40c328af201900fdb0792c064c26cf349e10de6
z98e6341e7fb18f55fdebb1ebfbbe11b7b9d1855c3f6a5575033ea810d14b266d0f5665bf0445b7
zab0492157289c8ad258e69f8c62fbef143c76d31cc5b5b48c28c58dc79118bd1fd57240139cbb5
zf7d1f37e02c706f86ca9640d05c7ddca050624a21fe78f844bace27dfd014f00b9a214b02db47e
z673ae7e79396105049a6281857acf774bdccc5b502e9ef131fa3240d87816cc3f772077b7f2a90
z3ce7a331614ba6c6bb394d9f627be7d7391b515964512cada72e5184e51f39f0e7b4e6ecffaa5e
z75b6d11ce79481edd351e9148ce975c74ba5fbec27cfb1ec3c58218c6c71c64e6b0b44c6f102d4
zaed3e0e3badba5d0e07b93452d0f3e152013dfc88372fd0610220050fabe63a4015d4236668491
z3c82ec0467cd92cd03ef1fcb053c4c8060bc6d6ccdd6fde30060984495c5d9296ad48ccce6a7cf
zdb7a8a086132eb496022e4ee05066b99d5873934f67105a64a203f6cb132d79df518efa92a3b6d
ze8fe0100760567af371dfa87117cdca1da4fd0f906526a9096f226ad53128d412cdd0ee3c5ad28
z2563d96570c144949eb23d9f179f9c46dde041291dbbeed7789ce412f5a0a3c230794050273930
z7ef8a5a1ff3975cc591e131c5a283d1b9ba7390ac6d53ae73e233dda733bb1cfa38e356f6eeac0
z2a7eb1086c0a373b3200358d4320d2ef68213167b5b519980f2edb1270df094334ce4714c57195
z330c50177e864d88d6e48dbba4ced1e8a35864fe0c92b5593d1c0353695271f4ae6d12f77350e7
z737dbdb519263d60baa05fd3d7157553849553342a703714c2dc9469941294fc97c04213f16e35
z7bbb2490a13a4571ca54134267b3a0ecd31b27ef38f8792830aec756c755a5a4bb2f58e7c6807a
zc85d17181cf054d1959e39355fbd823f74aa797188927d1256e46be21892e1f518a06577215417
z0911ef94181337731ceec04a3bf4ee9b224b6618c8e5674fe91ee6337f1811ed6d65f1e347f912
z22543ca7bd75a24f333131747bdc5471443ef5078566c052f54bd5a771195abe36242d6814440c
zb98514255bc0730332a94245ceddc72e1fa500eecab8013830e763be8a08a5d6653817ffb548d3
zccc6d10e32f6c1a1b9f9433a25a3adcb10e09a03a25e87374bd45657e6e7bb30d1953e7b5d7b4e
z926594729796f50a565247187362c54d55f726976b48a43ca0d5c22cf53dcb4790de807ad2a0bf
z9dcfe937b8022c8d56d1f39afe7e098d6a5b03c5f60bb4ddb68b362d9d2430e82ab645b063fdac
zda11f1dbb2f58d1f1fe70f58a4bb9e40df9215ab409235bd15cc3ad2b74a39d362d41eb8bb815c
zbe559d17d6ca082f68b62ad19f49cc71ac6ed9b8233a31b86a8c781dbcc3240877b84ceddf4604
zd941d7e95d4f2ea8520151bee8002bb5d44c87e4b136ec9b29e459929982939453fdf0fa8a9881
z28efbd037d31f9a7a8186d3e53a8e8280500623948445c760ec31be640f51b8244b4c1bae6070e
za4077e024364a77dd0a5110413562318ec752bc672f6d823fa7880fcf99147e45aed1c04fe929b
z351d485980644492f689ccb554e4665dc936ca17297869732df6338892bac8f12efa8fb76234c8
zf09e5ae4db85b5d1f70ba385fa7486864a30489655c198f51eb76d026d1e911a28798618eaaf6f
z35dfe9ff636e74b0207edd5917a44d60c9c74f192bb6b3ff5f9eebeb2320cad6a143eabca6b36a
z68ed18895fe23a31cf51c7efa4ff95a1c582536e508ff7d6916f628f5fd119c0d78dd173513dca
z733c2c61cf8c5bafc65b2a2e017b5da5a81ba5ed8f6c711d7125a076d13c2470b5865feb142627
zced111326513ef364782e4527aa9141bc5be99ffc289c247b77edd12887ae05a00f52b2927e9eb
z6e4f4fc9f8dbc309e56c88a8ba48cd9cbfc81f491ff1270d86d7c2d79f3e4889eaf08ea3861a24
z52516e7e5ec7bf58bf3dec0abe0209b09816756c64bc2d6e760d64d07ce571b9ac3476181249d3
z445e646ef136a9d9068d140e38a64f5399a568a7bd05cec2f1b5646e8b853aaf395009b5612947
zb29d634cf922cdac8f782c979656103f27733d5dea0166abc238f1f9f2c2acbc63c8e02534ef73
zdf6354e98880c1d3d7ca1ee76dececdf98a1d89822cbf5d13b6240a75c14b2b1b825ed1e609611
z69fa279c3a149715d04374f50a39cbf8f85a6f762492d2cfa082e71cfb28fc4252635236212990
z27e2d4789a81a972d56e73b6e0536573d0bf5181af6ba067dfe6567f9625f688681a8c34b24152
za6b524dbd5de4869c7b3b40391a51d6a805839846e727e6bd1171a911d03183712bbff985f417a
z700aa22ae3ff11772611654abfa8ea27e529346dfa8856dd0e0e563a5e4af70d9b4aa261c8a253
zb45bde864b778a78f70140b7f052ddfd85944e05b7b17c394c7ec8364aa7c14a0edf39ec045d23
zb38025b6d4324622208166eee25dac6e404cddb783addecf955b4bd726fd5c7431d19e1951c447
z20fac53abc5168231e0d8b8828befd5dc905ec9c1b3db3f18eb50f48ac04aaaf8f5a6b02cdaed6
z4734f5bdbcb3c045182302dc59bdf43be069929950f6741894ac5fb24c5a6facfa99fb961eb9a6
z50ca34ed78acce498a10cb0c259a58988536d10808a7d5fb202a7d785d5d1fe80f779b5471e473
z097b1b52e4c2a4651df4c23e0ace4c8aed02db17da2acc738d0a05c33aec565d640a35926108dd
z5f3bb14f058d02c28c9672d52e9afbe83d90ed7eebcd8669f3f5ef4b5110fda821edea5dd3ede0
zeab850b99198eb50b6e31671eee5f1b8a8b967b2ddaf6076b9dd09d39f322c5d5cb21bd5536ce9
zd12251dc31311af4acbe92b2dfc48d92e9b59e2283a109724be3415c8702f673f775337e9f11af
z991dd54866f48ae45c83343125e7dae00a808203bfb7d184a7aa745169155a4163728c6c5f0cd5
z82c645975c8a67ed3a88cda1e1906200889f75d8d94aff19ec4f48e69e8be94dc9dbd8099d5d96
zcfaeb2adc6804c22396d9ec65f23fbf7315163d391bd74b58e5d6fe812f9b22c4740601c4071e9
zbe0c2138f8cddc8ecea0ea0f7b77aab2b72be96ea72dc6625ad9a565095ef41cfd68d632770d17
ze1ced7c9f236af61109ef2282c3d8a0c9e723eca2c8064f8c0e29551f15eddd963b94fb3eb6578
z91659ee6fedb4be7d5e66e1d5fdecf1aa6f16faa423b362dc22d80013a2bd919bba38af9c2bff0
z607b1e9288637546ee75a657f665264046f10d2ff9a700a0cdbca43d0acd30a2a6bb4fdd4085a8
z371b9ec82e1c98303f66e3710ab41a9a0a6260cf55058ac22557224ec10bea21189b65ffd6bf4b
z72bdabbaaf518fb040866085f205a968e09f18140006bd6409ca4c4533b17818fdf61d57d4e86d
z43c847511e1a104e582e591889b17679278d8adef40ac67a36878cc18dbaab8c3bc3431fe8dab0
z3be6ab380e6903a3ea553be0af4083420824f7aac344b861aaebc4c9189f1b2557ca3937c0be02
z4d876ede4a558d5e4f2962885ef47d085b6380e7dce7bed194966e7473dc87dc55878a535f8acc
ze237ab904e96bfa5822262db66224c48d63b4f628681499466a7e55a6ca5737e398d4ba4e9ee53
zc8001b31b50dbff17b518829bf3629bd6cc1a398ebf249129b121e78d17de7093899cfcf6650a4
z02c9b3192111872c80d28e447dfd66c3c58f3fcd242a00cd4770171988014d453a9d0b7e918030
zd85bbf14ea318eb0d58686ac354a505ac322fe0f4b541553376c9f0e9b940eb06978b979d90430
z025faa18c7c7ec03628b370a87ff5a2609dbdab74cf0b8ca86176ee32c2b20bea700e8d9fcddd7
z8a0678a5351b7c4382d617d98ff986a1831f21536b6abb1ac09d1d7a458158186aed5087c47d2c
zc42c90da92fd94933b4b9483ff4c73f5d441e4d7b0c8d5d8b3f7cd909740e2fd1b987076cbb103
z897d2cf0f6634c0048c7008d5fc90f079ae9939bd6bc888de1b703894b85f40850197b9c6f9802
zb9b4a3dcc4fc9246b4d3dada43f41961aafd769a33c0b3d1b4f610127706c35d597f6b364e8ab7
z12240f95a43ab951a4dd5c21fe55b657c272cae38fdf421120dc23a1efbb4c6a4e5785a7877856
z359c78f3f74dbd1f49a127421623092936b9266d4bc3df28cb3bb035f9869a4ce8c94baaa150c8
ze1f5a9d1f47746862a0df75ae08278eb13c046fb6265d4c7c7bab1e9ecd9d6ac6b0249b25b8eda
zefc4fe3bfe927573ea76fd1b344130d832e48cad9d3dcd0e04d3e1803a0f9e285c1c7f594c4313
z35bcd44d7e24bbc00e03c0c643ce1b017767874fa765b97b08c476f12a2f9aec0884b056479a65
z4ce389b0ab9bfcdb24db7c49bd6ce5fd4e7e275c3b5c41ab50e55b9e50d9237be8561e64bc8565
ze0b016200dee81f49224c11333c2723b1edea6b66c8945310e3c4489db2e9b8492382306e3c937
z5040be3fb9afb9fe9df8ea57c5c7b95acc60564da6cb9fc059cefefc85a1a12797b31e00a8ccd2
z87b145e3c1981ae447066d6a92bc8af5d2c762896eb8fd32621df42d002cd70e2ad7e4046c8a26
za80bbe0d41e06b07b6382cb96eafe6ab7e95453e0017ca9acbcf1a9f0992995943dceffca5f5e9
zffb3234a904abb9653db7c054190a8400a386d48da637dd5388562a5f55936219bdc9ed184c7d9
z9d846c783abfa225bcf489a4f1beb07cd9773d2ec895a44c2e115e5f9e4b0a0e0d5d33ef827957
z0d7ac4c33fdff53b03897fd92df4ba937f972b3e58f49ac853b3f77b5f0b8ab99d985d4722eeae
zd17e3f6581d68e3870eda37011304829ddd6603fb595fd4d2271ffdaec73abd5666b32b689815d
zac4e0ccf8341849609d4a3848adbec0f4a62de53ddbcf2615afa7b2c6f39af275636c03562a21b
zee93dea22e0a02e2403ba3d403cde5dd295ebb3f98ded50602de6bc1abc407811806de3a2671d3
z1acefc62d859f53a2594440884dbf94db9e40a372c2145915f05d9b8cdeb44dab32a1176d20919
z0339e3db94b99fbb0f8ab0c1caa000dab7454252f2a704f91baed9c7e3b78226696e522ed322cd
z88be4633bec5fad12c57146620a64e9bcb4df76c77359581386a7fd0428952ff8790547e66aa54
zbabef77fa1ff8613e8f2df79532ba05c61d36ad317d785cd30df523d684caf7890920941d8558d
z020587d4e1377023f9011875f5187a4b8c50b8f0aea1a1d20f59debc31ef1eb42e845a1fd3ea45
z56348a91386bfb5c3c5bd962f982cc77218f5293da2a36031fc72cf8aae36a571f66bbbfee813f
z2a7c60951e2bf93b7a09ca8c26c91bfdffcb1811ca46855669031da48da9d4bac7a7167dbed163
zc3323f526e0c476086ed9360b09ad199a2aa533322007912a38c61847b2d16f835f659283e61aa
zeaf28b5e79f8d02301ccc0da5b90bcb5c9ac4e3edd63f58545536da3d476c73d6b301c893d2e44
zd6a58058cf9b55b7240a0e8c30cd0920ff90f4935dd0b3e87c08cdae114d57fcc5389d2cd2cbb6
zedcf81ab833269b2518a6915321c5b2c712bffbc0f763cf1e388490666ccfcc06d5bdb6a5c1b20
zaea03b5e78eab0b68804267958bb8d983fda2cb835abe6cb2fa2da831c2a75d4c5301690763b16
z6604ba417d178bac9d79c337b38ed31a691f04b1942b221c69e998101b07b725a575f0f14bd4b5
zdc7d81c55fa6c5fd0329ca3d915ed0c00de3ddc6dfdf0cc74dc97cb1739cfa718362b98c2ce783
z695312258d25cd7da226b90058af646844897597db18929ef551a303066af88b7b5db542c3192f
zca8c540a518a10057118fbe0d8db9ed94654f90f949d351684930c0412a0b7429a901d210787f6
z7c59a4205ac170d6cddc0f813b65de8811cf66f3b4910aeefe0b0cfa5b37243cf618cc2643844e
zd31b8fde6db3b6ec535b2e0a4ec7c8a743f0be35f73019116de5614076393b7c7c91272f5339f4
z83de0d7c8da9b7d3dbd08628798622872bf0b12396985f8750fdf7ea52ea8d0fb9dff17d3a82c7
zacfc2edc6eee630480cb41cf18a67e654db1bef19bd3ca1ea3228a2c64af8fe7ea3974aa5128c7
z82be60f2393b762ab89ee33fb15d90596ec7494ad48728124bab01e8217a1dce2b728aec0aa543
z03a1a2571e30987647f14cbd38dcdc58d0a33cf313723c2c1025770e7fba6aceeb836d23b5b4bf
zb55f115e69f54aeac17b1606a49587803978dfaead4deb2dd0ef8d386f92c9b43c0e986f78a49a
z3eb371ca0682378e501d1f0859f1b5660f8503c61a731beaba763f383fb5f090006d0ec29103f7
ze915a6b609f35fd32b64a9ec609a87ed3e014e2906d578b1b852f52d175c346d5fdc24428cb8e3
z70ea1e112719c1000fa87b487a05519838431f706c6dd225eee42d6f532b286e9bcc53397b9a48
z096c27ec89af9b2f525d2d238720317e4ffee8eb257b981f9f9d42b051c42467b9685b2c8f6fb3
z454c83509b38e1424ae2f8a79812b49c9eb0d1ffc656fde1937301a109e63c78471e2d0cb1eada
z253e07a392ed13ff969b59029e6c64ef4bd57288c0ea5d3222c463719148769f67b42b0a6570a2
z584e4b57475f2119969f46fcba9e76afc8226f5c3a8edd49b191461beb4a35e16fac432ee2d7ab
zf7866c5823eeef6ab0c7fef19547bc2d0784381ab02f99be920bfed1a3abf2c8120aa2c5af357b
z6f27a01b7d446d84f22b3e025be29151f9d691e395fd9737b8c0cfa9fe10035c0171c83610e609
z9214318cc831e0395212130617ab7833c1c27617a915258c50a2357bd0305622de3a0415c1189b
zdbee65a3259a20c2bf7a2cdc1583cbfbce772c0515fb2c50a986fe1eb22df169e180159f642de4
z595138a56fca4eddafa5abf97c4cb89189864de58932e6bc5ea9ff7eaf5c2e5ff6b5df5b0e64c1
zdd50c080aea675641609e9e00768a9ff7b25e7626327deaec97ff89646b4a5201e8c40cd001003
ze4ec5d807640fb0cebcafb6e4019bd376f9b7716a9bc85730cd7e7e98334d7529ba1ac5b8e1643
z7df450f7e8172a04f787c5fc7cf31f8b18c9a1d4b91ff6b6d94fd18bbb5ec1a3ba10d73c2048e0
z18e1c73904ec0f21b1bc8e191df4c3bb583d80071d57300a78cafdcf4a7df54c065de1ebf6fc47
zba2932040608bf0860ab1e9119f989ed05041db78fc5499a565ec0850554f25261cdf0323300c6
zc592fb60d176727519f8782d83df7381aa65887f362411a90a8b84b930b1401bbb4fee18e700fd
z708e2114aafdc63ca7d4e032faddbd3d87b5ee458be608bf8f4a33cf905c45350fbb0e2c19e0f2
z78a42d290e8231d236eac9e20900a05240bb8df9f29d0938fc98c191d4c4dfc1cf21abd0096f57
zbbb17495db9c4ed14a4ca6abc5bec776f4488286ba81253204d63603a8a96e0385c3ee458c5dfd
z7c9d153bd750a9d6abfca2faf5eebf57eea3535b143bbbb24b0835f591c0dd6e21709b491b83d1
z7b4f4bd9e50d0c0cfd6d244c54df560c644672ba7fb5394a46269b2bd6e08fd60061f34db27da7
z133bae21c08eedd070d3ead169a9f313a0ed55e7f983ef8dbb9d00a744b2de9085c8830d6ae51f
z6aa66f52e034c69cd090b6b6d8df73596f49091bb55305ef3a6321ec4c13da38bfb246052b1871
z81d7fab3934fba4eeb743b1325af3ab17faebc54d5319c6b399bb21125bdd0e7fb88925ac4dfb1
z7c5deaf3224f3ec529852570e73852149e9cc28edf5c3300b863820045ec5a4845e7fd5ed8948b
za3244f1e8749016126f1d75c3e5a6b2fb8c590f192fb2d6cbe6eb1bb55892b61e3d98b35a06677
z0ed530c910e6df0a2fb53a4f4cf9125fdd19a953162ca035ede0a2cd4bf7fff3b8c49c75e43eeb
z8b0eb769c29bcf6ac297e7ece432ec364dc6320dcc0b074520e8e3716217ed976ad14335b4d760
z240c60d303942c7615a1956b36c01e24bf0c66d9d32b40a6ca0b7d7429ebe8f883f29d5f29b0f8
z2ef2cb37cbb209efc1a45d7c376ee87f5bf6c23bf17a61b6dd58efbf6502f4ad99386ae84f1e14
zcc46307f15fe04fcdd53c6441022151b692009b679677cdb5840d92b3dce8b3368c7d8b0750da9
zf10fd53bd135cf43c160eaffb82869400f6b8682523819b560e11fe789bb04ea4f5dd04799e2d6
zb37b789694c443453b4d9bcc9b57afabe00a00db6b819ea04c09a5b484d6dee4538a63b183f741
z396629f1d17cd4a7e66d46864bed6158a1a8337bc08f4667a40672c04609e11afc0f9c4f36d6d7
z644939928b5fa8e873bb52fd4be8069dcd30f7173b77c58b627437257ba9f48f1c3760c5d4f44a
z9e5346fdc70a68fbc520794799db53366bc34e5a6f74df6590c05e59d67417524d45fc9dc9e10b
z56cd5cb1e9f334ee7b546edf3d982b99c4e85c4789a25496e04e9bfd843048cec58b7a8bcbbff0
z2adf2e029fff7dc60656a307a717f963142a2ea361ffc5651f1fe35dd511d16a96556e86cdfbe4
zca2c1dc1618a6ccf9a2b25e3eb0643053611aff1fcb9bfbedeb02e773defd1c9ca78a40f93c26a
z1d49710cde363d69b47fc81ef2040041941cb283fa2cdf2d0dd9b5c45a50944a7cab7bbd3ed376
ze6d7132dd462a9039221c00f1023a61e5a03364636bac45b952ff01ad99eb32e27d4c17869bacf
zf30add56be8cc9750284060d1349a18e5f83846c60a7cca453f5f20f47c399df566f9387ed8d2a
z92116233e225acf5ebf647b9d878f91a01b1fd43c31cbbebfcc9068778c02118fbe367bfdd6a27
zdb20c82bb8b3ff0a05c3de2a8f2829425bb207263ac5aca0762bcd61b9c9a6af357df476de5087
za7b07d0a828a7a8a1e0714b91bbab74f308be106f13dff0039e0fec921f5192351fa67a1ba6bb1
z6d85c09f5a41232c183307511d0fce197ac1da2d15dd03886c5c558de8a1b067917e35d4a3965e
za05ebbd4d6af04a71403ece6ed37e080aa10759ae5440263854843fc12d6550ca714b97e0a43d8
zf3864db3c4e462cd578ed3eefa63a6e8f9c9b37dfd042cfc28b78fdcac400547a43ee2c1831f81
zc89078167fe26f18d47c0b13abb8e5196252129566a455843e862dc0f00beecf93d7133bc756d9
z517fb53f46dee70ed9ffe563523f03f2e084fc64e4c360b0c00420d7f97e6dd9eac0f3c4c0ae6b
ze5d3d7a79e475b8ca581209703690588ee3652a698f02286a9653a48651762159681792c0f7b07
z85e700554ebdce101f32ef8115e9846bd0294212f5cfc5a0ef7b959176b9cbc370e455455e8edb
z4c731353559cd0521ea7ff3281fa4847e4b6b25ae928ceae25a2d5aa4b65ee461018564db4f7e7
za42eba707cf8a4764cc5e6df81eeea5f3f7b5a1f08f0972944192afe70dd9591c21dcdb1da2355
z250a63d07336fbb840d4a96f4d61560de5360515342e50de74532d5b0f8a6811a8600162d71fa1
z12a4f8ffcdeb88c70f49eb8d178e56587951b561236c0b2cb276754b6182ead42052b835610b2b
z833eb60aec5004749ea1fea34dfd27a5e46bc27cfebffa3c3ae4edd1876292a3838dbecc2c469b
z20235f46cbb0299efbbba88d74192d030ca09e20a26955183e51df55d7013cc735b30313821d22
z89486e05e64aee64f69ea6c37a97b5cd4c22a03a2ac4b7504f96a28c62eb78b0d0366e5fbb3d49
z149e25c0ed4f3bdac6838a7ad586047adc1a2dcfff417ebde65fe41c641348968490de0c48c6aa
zb425389930115658ea7ef38ba6bc437b81b4a1ea7c2c7d31235a27a14bd1a0153d1b27249ce053
zc97aff8dd8472d0ff1298d9dc60ef23a285b8962f09b4b0edcb934468f7fa10b169c0e013c4773
z60ab72d08fa990dd81a1bd489384beb7c3464356e2bac0a11328ded9c7eca52a785706aac1cdc9
zc1cbbd71ebcea2801df86deac02f7de60f259abfb23e901c74ee15c9af55a79d5355e8868d257f
za1170f759e7c6e318c2a1279342f6ec76f186a090b688f946261fff910fb1d03d19736a376cfb6
z421b03888ea041728dbab6cb65a62f4e710f811f8f2118f81bcab1d8a1d3c56cad5b12af77ee43
z39fc1a0348045c4bf0cb248891859d3e2108c09f14041681aa177fcf26b9b8c324578f2a13372b
z2a01e0301720aa1352b246c36699635207728ece2ed885ef969e89fd9640cc68c56cd54c8728d4
z3033317917dc091bb0920121559e31a40e152dd304436d7fd59339ab08b3c5cf7047909ae262a7
zfa4fa0d05a05ba023e687737ed03f4c74f95ae46737aa95efc827d1e786a9d1c969393b0643724
zd2e82ea0623af49b7b96336c0769d0cb6f2a55f5c3fc6a9b4f6efe9a0429d7bbda05629adc1d2f
zad8ce49b0323a86bbb6d09e4d416d2b7815efca063193ae7a69a6d3c9452391801cfbdc7ea92f5
z90db1c06395b8d7d98215befdf6c3919846a42cb1b3e0fefce272925f2bdcfa16b5dc525a6fdb5
z06019bb85e94de4ccc76a6d408069669b9a45951685f193272316f844f48f431763592e1d8c05c
z44ffed2bc62c552bb3fad0399e0eece5c14cb6295d2bc47685ca315e1373af225c9bb3e20c6ee8
zaa9178d2a10e369054196a1ce3e253981ee2fc2fb785f7afb8c0ef693e55caf34eaebc9014e421
z5d8d93b080f585e50a4eebf9bd6c5fb06a4863f1e1df2df5e7f32540bd165e2dc303745f004c77
zbd7a8c8c9417a99fde07fa5a3b5621a7056ecf093e84b7cd26e14eae1a9ca48852d18a0808f089
z39bac0b1b2cfcf82d5b19836a37b28c955989ba6c96f4ede5881e5a9f42c56a610739ef6ddc6b7
zf61be0a923f4b665e99f4ec7366497aa50c21051bef4162af14da07f2c96c34b9c8193cd277e09
zce6423d39fcc2e4382d4ca9c116aa019c028732dab18b88d3a063a593da74907482d4af63a763d
z2b8681cdc4691f9b566ac7b073601c84a412479ae8b0ac9335a3105346c107937c215c410338f8
z0a8e260263cd66f872709b187676cfe02831786402fb4da3cb34cf6b332eadf04db5094fc6b6c7
zade4b525865bae3d2e5080486bad24c06890ce2c57413ca9b90139f3ca688a20464f876a023a35
z6eaafd96b72a73d34a940cab83fba863361f935823ec2d106e70ab01cd9be9657b4851794225a6
z408998f112b4f0fc8f620d4639076a4d90bf65aac19fa0d8df157bfa3ee0732a412740e055e585
zb2d62527dd962afc16bb37d948d368b81222cdb29e9d994e94153622508f2ee418847a3e973d5e
ze01f251213986cbee544af7a5f60c1c87984fe2a9acb3d4ad3ecb902f89df80105c07ac0ce0c66
z4952f49a337c04e0e634cd38f8173b5901faa946681e021c85f7ef9f975f0bdfe49cc260d4f144
za289ce8362ffb19bbe920b4ca41685eb028afa5ff1168c2195aae8ddba1b6b1e09f8e739747b5b
z0629b7e1185cbdc98dd02f350a04fed59243a8d908c8583d1b9b617f8b07b22eaa46b341281fbe
z62bfa77d9a78263e000f6af080f89cda8dedd2ddaf21f473fd4f4cc05534dff0aa1f98255242ef
z1d54e0f63beeb945706cff6a2dcc4169515e7cdcf6811a1aa041e198dd5260ba13710db6339ae4
zafd9eba7efac6b45b4cf47ef16614392a78b3f230a134b3f91fc94cf07f5b83b17f92f086ed981
z647a1e199d76cd24c07e72af6f11c14abb6b5196c6dcf241447f7944847d22f95561055534d221
z7a4ebbb0cd1f8a73ea82b6e0534c4c82213d06b40f07841f3db1337201ee4674478b5f24b25c79
z81431a80a13ca628aeb873c04a0ac47039d44a4f0e43151090b6c656264c8eef78c129c09c34df
zb428796b940d556eb7fba284deec215dbedaf8366ecc50dbb7697a626f47b780fe97a92b11b295
z89ca4c71232484c9920486565b71823a940a3301a5f5275335439ab70d3517d91a146744590a7a
zff4658beb088d92b2fcb3b45ed47b56f9418e6dc0a6e2d11e70e948f771a846ea55b646b92f31b
z3a146be9b1f1c454a08a4691905137af3bc8faa59463d17293a01bea887ea6ae69435d5bdaea3e
z935d36eb8657db8c5d165e1896f51017580cf7249bd55533ead4ac23e2a4e7307aab4f5f888aea
z5c6290433633fe857b7af9a38a924842b36cf703220c8a45c1b0509672526c667d9be2eb8865f8
z5405f6f2623cc35fa29d35b049754292c209832507954a3b09ad6166fb8177dd75039b0d1656f3
za0015ae2f34d5bd10249dc785b9ea3f3d9a0a432d719e42e08361037cd37c99e6bd05dad026dfb
zc92f079c9911b266dd7a84729a6ee30c6544bb987f263e78ab370bd87572d9328cb3eae66989d4
z910f808471011b99140db3d11f0c352a58b5632210a4ae3dfa3483f004028a59c9a6c95ea6c159
z4078e3b10a1bbe2e3e003ee9865aaab42ad880e05d91bb0935b374cc670c20de509bab8456a218
z0d8dbe04b2ee2bd0c1559dec6d676b0442c746b125308cd2dfb4f4c5d5680b58e7364e767a9cf8
zf4567f2a7d5fc66876c600b48856f03ba2d9e59ef67bc8493f46b4ae421d84f0724e875c818f82
z6be231df008a9f3271b0f688b7b01823aa65b5ded96c6f9fbad77b7f9b5372105cdcc90742d81d
z3a0731c6088ba78265f1efa52eacb99581090db319ff6a50424751b915ca3837dfd84882a6864d
zb2ad1664de88d83a3ebac406a0ef4cd93bcacd0668633f29f298bbeef16aa5e0e57204749ffa7a
zfaa5200223b2713828f9316edcaa76fa20a8fc88e60585ba594d45007e0f78bcc791ce403b9ac6
z79964f6e02d439271347066ed0d0698628b250bf571d3bab6ba052a1d639efab1ece4132d41969
zc91390cdfee1cb7257337c2494538f88aff6ac037b41a5e2f2cc1d2d5826b04e0c11baac913292
z597c101190c671f403689b43ba1c54b60799b5e0761a354680c69b30811f51a688f5f23af93c9b
z8a02f842dda67945f0dd2b0c1a4aa4c8fe0bb8a455b239196e6a11bcb8877443b824d0010f5d27
z46476238729044b6cb3dc6919110d5de8a506e06e41eadfe20a0d81cf59ddc9633ea95f71110c3
zde4636f95eebfe6b2385b7d50b962c7fbc1ad541938246ebad63634bcb1873217173c271f08b73
z8f2fcb722947b65f442d64f487ed225d7c8343838908f50d20b735482b0ddf6734d326ff20c7ee
ze9b6d98275fab084f5c45c91bd16dc96ad3ca0308ef36ed297f973f09a5372d290c9b7b99650a3
zfdec3b6bd5d59f9092a67cb1d2ee5ac82a276a9c2c33337594c17e7de55df94350f16949460e60
zcea5237ef2fa68b7fcc99ec1fce4566c0d6229519fa261ddb3ce5c4832dd965a21680a4e455603
zc303dedf37dc75a8c506995e4c2c737b4fae0f511dcb243791eaa3a3f1b625f5ad7aa03d1a9f09
z57dac19edcc83795ab56bd9cf9ba51edd528d1eb2980c786476279d55206e77c61584c9098c678
z32dee5c755d427bc4a9821ac544ea410dce514cb965a5808250117cfa64ac5b2c2ce8b1e838248
za8e39471de0dcbed4e0b4759db342cd8797bf7931ab0cae5f9ed923f93a371fa7a0e703f3cf302
z11be5f16e7f0d14a5262ffa42dbb944df569c2deb2a8b73070a1b080792ec40cbc5b708c172406
zbf3afdafa1fc7cbcb16d0d39034d9e5b5bc35934e339db9793791ce65c305ffc6f86bfe65cf165
z8a731e3764146da51440d59357f6a007104633b058d0c3f731de8a2e222a0ced7d135b21dfea2e
z7cfd5cca5831a98f1b203ddd8d7d7e31ac1926337cb9d046451395c104af52a1d7031f64b4658e
za77c2171dfff11788c581266f791b18dd02d2fb8d10714abe2bfe6a1fd241e61ac49e28c2e8c72
z18bc44ef414fd9fa2a0e65c4e9503cb94f16a4743f68b24bf5fac8ba7109d71055a6fc13ec2c16
zbad1ac8fecea6dade4d082512d895d6886894ced29832e40960431d2b7e4da7c87f19e4ae52046
ze9edd3ffd7480c67e73998deca83391442e9865714af13bd14624d12b0c472ba5a727ce7db65b8
z3c74a3521f18849a071818759ddf84918f7469d43226ce2bb02b6f1e025abb92e09e7d98962ebc
zaa5d77359423416a2185820e33d91a289b395fbd33ba8ba17fbef8284217094013dd0afd72bafc
z894c59923628ae9b882573e7e9db26ecc52ebc262da37e0f54abf283802a4db3898aa248949eaf
z7c46f665ad606735262f3c5bd22015a3aadb9bdd9a1784e95bc81a550b1defc60a54fcf5c27a74
z6fd4745f95360303b528cd0af471851348648e98fb75accf0d138783dbc5644f8a69c0016a6eca
zf2f4c6acff0f6d3d6ada6c44feb63474597b65349a952aaab11897d19b58bef0a1cd8069fc041e
z85385d6c9ce00f2ddefc702bd6c041e918dc704415db9446d9fabfa4640b66ef0c4c21601119c3
z841cb81b47eee79f0f7b6209479c7d227ae0d171c9b60f2d937a5c410e35782756b6b0b3779277
z0f0ce485a912b5923c49abc4abc3ce7fbe7b2ebcd40b08ee2f0fb23f38472df80f80402bacf5e9
z983bf8d1d3974611c9ddf83ae6bcc94537598d6ce1c1cc3fb2fb95fd6bbd2f77c95bd0fbf02281
za1ed89fe689456bf89354c1ffc3d296fa34220af18cf98e5c6c6684d62554e791a5bb18515460e
z6cd2cd007492c39e5c2f35840aa6b366c93af6e22b39a325a4943c0edd048cbbf8cc83854c64d9
zebcef172e6954c92aa443b2221116339528e078679ef732d3e63b58e1f0940a9a38589a50ab700
z50c4b2a003bf1bb0658f53d587615afe48f7a6474a920ef5cde714b79c7a95f87a1724c7374d6b
z31533bec09cfcc24f60a63b032c2ea7b92a7db496a8488aed04dc80f0a710ce35ee2d55c7fc8b9
z0ff4eca47dc255d8f051b0c5558003575725cb0ccadd55880f4d9b04fab74e5407967de0994401
z1b9e75a9e40d202233beeaf77d57a7d846b780256552d95388c1df720b1df32867b88064d385f1
z56875792018c226618c989f9059ad93b9a19606d938fc39b7d4cc479f068cfcee95a1720171432
z4eedf92371ae84881dd1b23371c4e135a60281fc1239d24f4d953ec8da2c9630cd492a93066733
zf12a57eb1e4ab1869db82898ced1cfbda935cdfa5356c11f5df99228ee3e7284d185dded6fc8b8
ze4afc078326babedca6820817d892a71bf959abab436af7cbada2ce4a11508d972549336699cac
zac8fc6b2545847c5aa2ae54d7b88bcd42addfb66f6fdcb9816729813364bd447a8c7bcc6588b5b
z86e5c35c89addc17fc95a09000de6221aa41afa9b830153e9b57508ca6314b2738049e8fe5f8b7
z9f01a25178b4aa0c19d0a619117703112a92534d460caeddfb48657a5bd1f978d83dda23b1dd2a
zddec2dee9d1b532bf499cb3273bbea6c588195e9dae4eff2d44829d0d87b9248d41fddb0a49ad6
zb2c57ba3f1a419c9cfd23c4c824decdd285603fa1e807e74880b4d583a5e82c7642b79eeb63c30
z2f6fc47fc1e95223ad9713bd9b42ea019e8d98135b991def8e7d3073dcf49545ca608bf0ba5d43
za1322e9b09f09d6ef0de742fa64087d97410d988a3ca0ad3ebbe9500f328dc6d470ceff70760c7
zcb348f5e648dfbd9a89f25def05c1e849eca82dbbf7ad85d479c7dbf7792dfdfeef519cd07f953
zf883644e2089e2ff7d173a4962e3a2e89c23e185a766a7a6bebb4417ba5caddbd988d2071757c2
z664050dd9f9ef7090fb38e7a16fb5f9b84026b37bb6ffe203249f72dc4f443242a957e23a24cfd
z12385933a2252081c126e608ddb77e7f837b397a7dc63fdfc439231035675948e5dc1feb4a2fe5
zc86ed9da08674786c35f77d0a284ba59d5a4192145a0c450ae50222d838f71746aeb33c38d063d
z4ad1c60018c4c81e0b8f9a341fcc2ace68bdd4e6a3b635a6f600d39caf3b14fbd55ba5e752aeb4
zaf3201ea91c8f3e7db7c583760def795f5c7a03016b472bbc02879f0fd2215c42e05871ff45fd3
za7d7c7693a0fe7541343df7450cde52ac5f4825d07d943bfa30e60055a07032244385486989907
zc3354d5a6f7d1e02e1aa78c9a13df63479ea9f283a017fab6d4afbc2c399b54edb26c664e45787
z9108997abd90994d5afd8767b54f2d57c425520ffefcb94fb42728e64d508f2d2531f3d457e97c
z2006fe80c9cb21e4fe75adac0114dfc70155bb5efb5a396099a1740e75c30794291643874d8840
z1c0b89db4d0fdcf7382b8ba88b530aff38af8dd1c584094f80baedd8bd34d57ca9332737088e59
z2cb7bb07a6f890e689267eb1206bfdb30088b7c85cbfc2df9caf05b9ebb5ea77555a48166ee39d
z82cd7a8f67107b76cfccdd94ad726eacb3c00aa1e353f6cbbda7a6160cfb8ced86f5e80ddf7c16
zda1ea63fe6c137d6c216d053100fe8c2ea6e0b59a2737d9a1430d027df533d63ef34306ffcbada
z4f04f35e65b088894a6a56ae87e8b4ea46c9dc9f33f6724ca6b43570667a3ed5fea72f21bba5c5
zb4731fb8830d71109b946254a33a19343104f5e194e110fa14701a52eca9ee45190f6b91486a07
z88102a930bfa8bb67f0930a43f078ef6e9113f00e0fe141797d1c4f74dadd50776223f3e868bb3
z02ee5d4ae61fbdd9dfe60f699201d62bb29aaa81637e66b2fce183b300d2c602708f9f45ac6e43
z00068528e1fda5e3b5b65d148b0aef88981194efc628f2e65e3844af9b7a4d97b6d17f4d27c73a
z0e95b7b06d83e1b3461275de2b4eaf55df5d74c4116b485ead74333ebad6d5c24230d85963c81b
zddf7c7d3ca28f2d33d66383ba80ecf3c02bea34050978ebbe972cb3d1e718c660fa3aa85650029
zdde4509ff4cf80428a5be64a95b3f919818440a5077619e380e549e6196612b104a94f5f8635b4
zd7943992dbd7f5a86406da602a72f497a9cfad9bef11d98dd1121148fa7f3792a2b7c5f97722f4
zdc5d5e56e08c897bd9f66a7767c073bd6143f2b2cb0c4649c46388f2c5d544eba7d96f9e653b59
z53af400a01bb1423c3bb3a1afc2f553253fb0bc3dea45eb6530543b908789a49424e86bb6de7ef
z3f992a4b7c25ebb0a468ed70ac92cbb6e79a33d12fa8a7dc84e8bdbbff4d95ffb90be50e5f8d9c
z14fe952c538fe7f529a569ede9e16e2ea77a2d6fa68f182d8e92954481bb3f14d707a404c10c00
zba93105a62fb0a9ff0da1e7dcaa665ae3dd46f2c2a294f07acfc672043b7032ea2274078d25af4
z714e21f7f9672b96ff8015da49bd3ee9d3e3ed7c184a4c844aa3f6294ff283216cf73ec78aa12c
za9ac492db6f21cb12c511d1af911434249c51d9a36cbaeccab433b51f68b0f54c30997c09198dc
z14d1c7a624f3de39fc6e2dbdad7941d173fd7f7455d1a5c674160a48c78e4f552454542b72b78c
zf787f6039862f2ef75729074b123be096053697326090bd57340f531e14d72fce8b93e90712f21
z26d3eac8648af8d269c79cd2e8ccbd3f2d341b007cec34304a7cf260c6390cd540f77fa6e516f8
zefc328672632bee0a295670dea9d3a357ebb6d674360f11bb0ec0a224764e44d993e034adc9034
z28be99a1845334356c5d394ec9eca98db2c7f82106cc8c847a7cc7d11f08c489b3a0a2150c5fa1
z707137093259e654ddf8bcf90a3a8b48fcb6f8849fd8277f8009eacc5cd92c921f7c948048aef5
z1554ff94a63b49fa86adaff74827b5fd8d723960db0528019c8bc48d85d795702531a5c41c2298
z30486a820b5e08cb14e58d0f6f31dc40c68acd8a7f3bf700bbe08c0c52668e28b6bf011a61125a
zd285cc7f746a4169d2b49f3f8c5a0960b9b784f8b922f2b039c925375cf20c4e7302f84b4aea12
ze7c779ec10e8d441e59852b12c641af59a36662c17754e7258e3c1960b83ec7c307045ab0df412
zffc59a58f7b9154f989d6c5c45c08660ca2802ecc68229df90076e685211d4c6e3a27e461aff7f
z20f5de76b007e51104e0e867800cac716e5dd542d53ec78d1447c3dde738ec89d362caf3a7860c
zf5650335ed6b5855c902b55ae35873c01e83b466c98ccc3968f1fffa9046e907200f4b6d9f7e8e
z405f72edb312f7a027770a5336f7f0596b61a4eee612c1e12c60b56ce2f5cdf0d3ea279710e3e7
zaeb55d06a047f49aca96a515a4427e0116d4965c6b86ca24062bf035cab6be57cf3069a14e7c54
z1979b4fa3496a3763fc469aeb4420d9a328c4c8f3f28082900314e3b2fbf8036fccae8ef5e19c7
za8394f66b48ab53dab34916377456c47cb464e1810959ff9ad6da2dad8c00e39ec0ed339dde1b2
z92c22452e041ae10e4f30f17598d2ea8c1d29c6deefd03056316f0c205dc067dd6283ad74f6a62
z3c87e58d4ccbdb733c1121bba8ac47f6e0321f9c36f9a2e8de4a0de37f7058a61222e31112720a
z74d42fd229fc7860f51a8ebba605338bf1c97240c5b1fcb0e115de2feb4069b8393ffcf15f1bb5
zeeff9cbc6bc520e483b4c112f6309518394357259e47516493929b41f245cf79b33b211f4a4414
z68295169c9b1ea2e0bb6a43ffa843a9ceb09e2220682638e56d1a2eb0cdcf449bea53288af2248
zbe7b9760cb3f41724ed5f5c14cfe19e8b876bd0b13488cff9b63d63bb73ded7297d155a8aa7ef7
z67b03c5ca0934fe22a0fd64524d763e0d0eaac00e80de6d9aa7041c9713ec6e90b3702c031b191
zb7643b5959a2d729f2b1eb0a242407e809b100254e1d2cf76db5fe00d4d5802791e5f69dae15af
z3ed806ec9a25618407302ee8218582deed4d6fd219dc322d674cf75f3953cf449916f18308f7a8
z2c6fbd626f11446e67711f70bba1600c8980daabb2a77ca3dde04a712a2d195620d5a4f9779b31
zc0458a94d7142a0efff6f37283b22e28bdbde5f0b551ef8b357ef8f112450a76f00e550e286c59
z82940c0bdefc17bc9a02f46e7533db6f57761526beb4853e8725051deea231f25f9f5ae8724a77
z2050a3e47982c69e44bfbea02aaab07112bc2d46c7ab517764aa7e85684cb939d0def2fffb9efd
z23eff9e343cf2e5e17fff38a4ed75dcb7430f30ab9a7b817e561f26533fa22b17ccf4ba96da6f1
z2874ba8a222c435af3791bda8e9ce5fb1030e13a93163937e69ee53c9cc9d46a5aedf2e6844990
z660e4f61d4b8274714e8b0410eabe53181aec05ecafa21764f5a0254d070fa37cf2e84f83f343d
z14f6f5d21ed59c124f0a7a71d66f345fe36e3d94ea1b25ef619e58bfcd9dd4b712ec843adaac76
zef9cfdc43c471561a2c21e5eb043609b835d82023494006737f59e06eef0c35be8a26272db89d4
zcc1cd8ec0e569fa3ded99a665f4e4661f43d1d069341229c5c4726fa6b67180ab35821f303e1f3
z1cc40a90087ad90fefea28725fd0d5df2f29867e520adf69e2accd863a52d6ac62993a239d2b14
z6811b1dfd4c299fe69bc542219252985ee43397210ba75a86cc211de0bce180e38779d1c468812
z0074ee6c436d8f4fd875750c4b0f65760bbad74b51bf074c501fa7a9dbffa57d883a0e3841a127
zdd1f56d50205842bd0225671ca1d5add7f05f72b880e011236c805ed769f18d7fc6dcd8da0711d
z36b6e1fd70fb417fb615c08e4832c1422dfe99fd4ce0883bddd0d1d01f15ea510fe5466acc16d1
z4fee0bda0e510523d6949becfe36ee99de05bcd6efb0b0a3e1c2ba37feb971586299bb8623060e
zdd8c872d526d7817d657424d83270fc8c5ea168473e87b1eea224acc9fb03740ee94ee3ee171dd
z3be0d7369d134449de74d7d180112c198907a4d3b6d0283d100647edaa74803f06476bf56397fe
z79e2d3adab76ebbd94c542296431f0edf81e47c3689f4b6b6c95a1a6fedda51cafa0f87cf0a0ea
z9d44e1a3348dbe55a13c18eb3afef326b7124c04cc226a874e8cb1f478e3d8c16abd7de42df30c
z7d7fd5558b47fbc0123004653c22a418b64704aa9b9179e36af15d096afdf9a4d616b7f3ba5d99
z43cf430ac808f746a4e6cff268b77b02b5ed5a1a6ea88f02534dcb61e0a552af7a41085611d8b4
za57cefcb672086a454f45002f5c7414cc9404f4e4f76aebe5b08ec4af26b83f0eab96fc446f76d
za00f149ed9f5f66c1fe75b439116371b3aac4e40a4976a6863e14538df058b56d21d1f7e597a8a
zaf505744a0555056f64d09d770ca69be2beda24fab2d0ad4fdcbe222585ae025ca5f778a59799f
zcc2a0f3d42470cd0de46f902b4672b2004eef9dedbbfb20e87ed427a552db93d8b4f5237745cb7
ze0b497ec757c5be163457a86f853b195c56ec96b19b84054cbec7f9e95f0aa8d5cacaf312754a0
z44aa1390d87f0f46f7528803f8f26f6ca44f273b159e1fd2f697f4bf621c8853c9c15a2d1f914c
z87a4cf72e2a9109fe5640b3f4aa3111615b25abcf5de0a5153847286d3146b4d9fbe9eb9c30d5c
z636fc8bf7b93c00a889ff92fea472277bb4884e8024eac515e13eea832ec676f7de0278f8adaa9
zcca5bcc1a72d65f6d4b1bd5787c61e4d74c1d3ef2eaa91c50b2f5b480aba8d09038fdc005a1dda
z88db0919e8e11909daadd259c5e881fa5c6a24fa6f0033ddecc25827c949738755ce9c1c8585ac
z21857a44d8cbc3cbd9cfc4173fc4be9c8e3e5b885a641adb280511db2f3bc1799910520b16345e
zedaa263d2c823dc896f8c1ce5e390dd611fbc78da55ae45182a28126f682e6e8b876b3ad00cba0
z7366e410d08a64da6ff5c4e4d6a6458c8e6922d44f6e97fc1a49d3a4b757ec1c0871b7e55fe2eb
zb19088916f655d6b6634daf0e0f1c5c312f2a6ab2fdc066656724e5b7be2de1f3cb65eedbda972
ze4d24d9ae1abe798ee0d5af295df87e6066666acff1f4420a68b40f354efb7950892244954a41a
z80f39be1fab22dc275f15694d5a759076f088a2e986d38ffe99f8cd0cdf35b26f64f532e95c2f3
zf5852477d8bfd4e9fd3911d45514f0a7f2345520ed262b3c0d9f35a194ddf4679f324054f1c02c
z0c00aad3d5559d03f44eeb6a1db1a5ae26fb543e8786ba27e805a403161fba869e474930cdaccf
z68a33f7d174a1fadcf4cc9888f53f6296119dd8b94e2f84313d40b3b5f9432bc2369ef8d53294f
z374565fad07c7bc07601b0a59e85d89275744cc7135d2544db7c4220c0545350bc88337f668c50
z63e949b539fa175ad62e443f1489084535430df65bb888092e5463ad1ebcb9b0c5a7a77bf2b155
z5c7e1ee4780b38687d141f9bea230f2f10c50906cbb2bda61f99d6f6b3c6170e114d228ecad3f0
z3ad791ed21b5779cbdb4143f6ff2dcfd9b6ea16b0e0bbe6ef09fb005c94d52c41ad79392412b52
zdb9f42af52eb3fb7c4e8d4ba99df5fe19be4895e321f8af6ba2e70cf875df4d7cbf6b49786be2d
z7c28411453127e46524c58c6098598c9a661c792b3c5cfaf4c66c344e73ff08b9332560a6a4e8a
z642462db6611e293a9fcb3ccb64dae5492c0000660666ff32936d7e1384c17bfd79e003231cea0
z11eb5cb4b1a3c08d3f5a701d6a28d6a0be4f62855bdf0a850925a7e405f2cedd625bd2a7ff0ee9
z9a193da8abe8b61c683a5646c4fe0796636338ac55cd2ec46efa0ae4e0a9540cbe3578df0a4a6d
zcea10683f856b71e3e5154716310e9fba78dd53fa5579aa429674071f8d48735b0138395599c64
zba4869ddc37717e4963992b89881371684a616bd86646f1f6b1c10768b2f90e48d8fbd7b615f7a
za4a4c2205fe6e6a664eac576a40c677b18121c532869a7996d4c1206a8f90f3586e053ab7e349a
zd754952ab5c046c7dcc19fc6b880d9df9798fe4690e9e5271d57676b6a87eb0eb809b4f4c1fa98
z720a05746e9a8850a2268f7e81f5d11ca14e64527daca269890e481175072e142bca54333f7d7e
z4d6ce2763bf8a6eb109ea90904aefd5b847fcda3056573058f7b5b4e84ab002e9ef6fc5a09de1c
z7271a7045a4fb6f733cac14b81ad5385779cf2f44fc1c5b907207f9f03104a1b522685526327c1
z337aa1eee4a6b4c282667978703805200b1ca8c82fbb4dbdcf2295a4e582e2fd711f4ec1a7f0b3
z5b8e30a9021d2bd780f3fa9a69da327921184510ea15c73c8264d920104e6d242499cef8a94b05
z4707a59ade4615d76d4c8d8cd63fe8842e717421b1a1911bffc0136c8eb9763791f7a875527710
z28928a0bdcab4e1cdaad8473014cbcb70b172302c6f91d216e0e5cfdc8347643b254d112feb82e
za9ab5bf27e9648cb6557a331089dae09a3bdec68780c0a59f09749a34b188e5b3006d588df92cd
zd32b694729e5ea3f020a5429e44d0c8195a18d5dd5d40999745842c5c89bf4f22a378b99de1337
z63384d8418927063e1df399f0e52e1514b3e3f5d661544f9786f986982db37d558f87de3311f24
z45101d1a46ba9470a2bc8f3bb0722ac72c36e6bb34e705c80d7dbc04dca06cafd222c68175700c
z2d5c59ba77d90aa752b9ecfc40708a87dc9fad86525ee2bc0c28fe3a471ea32c8320c36e457210
zb35d7f24154372b4296dce9e016233890c36f7ee96ce9f828939e166327b4b5a641eb892f2cfe5
z24b599e3ae52cb7a312c75601563fda080c95783a6e1b8abd87c8306e3ad93a3e8b24a4630b2f7
z7c2b85e5892d836b9d5ba28fc20f3fcf5df88b70fdb69ddbeb75cff6802c5dddcecc9b8f18c711
z5808285edc7f82e5ba564063b3e9fab58aef1d8cc5d41c1e41b3f2f5b82a7e11e347993ed21a94
z6b05d861bc798a2256ff272bd2695808154e84b53762d679a355392d3405fd6eb7b889ed0c1fee
zc5286ea7d9f19019565f62f7f8d2862210f67d755930904300ed45f9522e08bad7dec44fadeb32
z6c949999ddb3e016a3d18649955d0210ec16179aca0814f1a88fd39b70ab55946004e30473685d
z2471e48661d30f47de4b457eb38f07d5b7b2c3aa7cc15abd523aeadec31af46d6a2a2ed62ee509
ze6aac09ecc11ebe463f9e80f49441bb0b0f7c3ed49d6724d86486fa6742d17599ffe3c1b33f90c
z2f2e577a1390b6ad266df3ac8d8c13ed78a8993607ac491256332e7c4bea71dab5b3316b8b8f12
zc5e68f4374e8f4cef1fdde3acaba7511cd1658103a73d000ce6d42c282789b83f5991f856ae8e2
z67af57a88a98767011610c014130b9e473557bdee464fd72f89164a7d9eb1af5bb0e04545d6896
ze5a40ded7aebc10df24c53d99cb92bf3dce5a9728d44a40c3b2a095d9d31680778af52ca3e89ce
z3f727905241b9e70465d4b793a196475c5fd5edbdc2d0f0976e3dc9bb7cdbfaeac556a0e7eaaf7
ze5230b05456731d8388cb491f924a53554ec93d2554188a8ae4d2e8154ac806d813c7c0695a1cd
zc206eeb6fbbdd818ae39e3d80783b4c008b2e2882abf69dc6d08cc383c7e30ca49b32aec7e92cb
z4264389288bf7e1afd4ecb9988a6c8f452ab65a23cadb7aad229c5f7a9788958f01c95d0a379ce
zcdf62df0b7b7fa0fbd452ff28bbd4f96ac71111458198062837cd7b7959cf8d9d10a7b1719b48e
z246526ce03ee766b74c7be6b73e6773f12eeb9ff8d104c2a2d20253d6d4a6872ece67393524d27
za19e27e40b3a98ce97cf58ca33be752d110fa6d7744b25be9df53d3ce8c41f3fc18b2a174ba942
z3f7d019830522bd07f2efcf4b94adc760549be942955cb89f167eb77b90de8a5766a641a87838b
z645c0f510db95bf1f62a8c402a5fab4de06370ca32c58e7e4d77e2667e07b3169e464801ac8e2a
zd0a7e515bd578e8c036c27ee8c710d3d2b743f9ce8b2fbcf9d6a699137722b53ef813951278b75
z7eb3a113a531bad22f72b486153a8cfd03b0147fceef178a3731b61236bec0f448b0468804039b
z7919689bb7f519bf8d2d6d4a665b9a0e7caedb8a29c12a22dcce14512d551ddc8e12cafc9168f7
z9e61b4d0145abd56e198b84cb40f505e0d77976117d82fb326756c2144edef9c9715208eb90e85
z8e0d701613474dd551b2b02801be322699dbf1e34a2a6bf0146fabb4df47fd42b1f19240d024c2
z4480ae8f0281ed9ec9f9a0b89e98817c377c2784d32886e7b920617e32bd7e65314db2873dbafc
z6fe895ec4e9450a7b95ba229dc2cbc4f31d0bba64d1aa80ba53e212ec6f9a8433c65ff016338fb
z411a759d5d831061f9a8fb8cf87cd43ed994a29efbdd44bdb20bd1e9e8300777b277e82ba6ed3d
ze342cb7ee7909262c2cf5c078e4b23013a2230da9af4d4ae221eb56b298c9eb1707f8c28e5efc7
zfa02ed18df4c3dcffa88fa162f357e0717f33710682b57bb2591bee7e3c84db1f05528206808ad
zd1df95ea4725dbcde3a74d07d213ec1b24ae6f3fdf37b6686039735ba5b3495088dd0dc37c5d2f
z2824ac684b02b17b0408a3751e9923d42c0f732d0da7412057b284b57a639a7c213b02698bc421
zad4275387dee17ac6eca550a6bcdd9bdde6c0220c38b47fe4689384fc4e9258f0a89d5633bcc0c
z27b39876b8cd521ddce48099f42c18521dc6e93ebf217ab705ff453ce117471a0bce3dd03cb5f2
z2c85c493d2447596e784578e73a4b6a38dee033a8f93edfb6e16b71f20028ca01111d4609e35be
zf05a16f9ba5b228f585b819c4df67ee1433263f3aa32ed358dcb67e7e52092a73485e2fad79199
z6ee747029669e09d788f6d760f2f3a664da4a09eeb9c32fb0d53ca2b4b843614203a1b83546c4f
zd03fde02c2cb17fd675d224b97d2bf75f357e2ebf379b4727218459dfad2d9785f2b33045c9c2a
zd2d11d35ad17ccc4499c661261e1d710aec7b63944b5ee726cbc844acf14596176481925cf7785
zc5c948e648c680b3a1566625446a641c659b759e4bc77b2b95e20802a6771848d03db457886382
zc8b9da9fa3e06546d63caff9ce20de78d30a59e50fb291caf47c1f1421de187a160746fbc7c273
za8fcc164720d9f487e6c676fa0c7ff7e06de4c256604a1b7fe071851d1656a6b5999ddfbd5c33e
z0fd138bde933cc76e1b5029fb59c61441822c91bdcb9cd15e0128a05ceec693611df7862656c4c
zd1ff4e5847e879f0606edde48a8ea29c897de155f0db5d907abddd45857c46ea8ec168cf7679a1
z58ff2cdac3e2e4ad598534f02dd45e4fd99a2e6c7262df2fe6b08f787f4f731c073c0975f0cc27
z20c24480e8037953d6e84bbf270a727ba2afc79a5f4a4459d54a4391e4ec610063cf87e528e801
z81033da341f4ad2810ff5452c3f5ae68e4db78d391d5e707a31d199546025763103108f64d2909
za43b130bf1988070d4ce469e0715191f195f049ffd0a0439e8e7807ed224a7efdfd56a4c2d59e4
z5b273d60464bb6f30b6944355e5ff2cc287371e0f7cae403620596455abfd94acc3881e9976e46
z9d91c85912cea1e354644340bae1fa0bc171f92dda3fc51de04e51e20a895db0dd173e79ea7705
z7ff2633908ba81d69ad3bebaa84229c67fc4a66e8753d0e9ee0e4ede1e07c2504c785566d86b95
zf579151a23ee243c294981be2f3ac070da95fe6627a9f848c7e75d7fb355943e1c3d2e8eceac3f
z5746e46e814b3383e5208a975c043668d36f7f180918bae498525ad58302f6baf2161f3b2deb6d
z88a5e58e20557b733a132dcf1d1949cef280a00b43bfdb93aedd2cabdd05ec036f9a94734d0c2a
z9c7b41d2dbb90e7da20d3706491bff8a48f6e43cb34903ad20cddc794a48a9b66ec7aff547d4f6
z9b72729c819b014d59191f4c17526dd9ad4e46eba364fcd06b01bc8c5dbe05e2e20184886f1828
z9d2a9042b9c0f8585532577e61ea90c8df9881d4438d3b1dbabf8cfff131b2c81168b0b8867c6c
z2c77bb3ec4a4f514c89ac56a49487ca2da26dfe3757f493ddd8dac5a60cfe34f18c4c26827042c
zf1c78f672937dbb336a5e8456201467cf29f761065a60caa500f9042e7df5b5eaad678c043a852
zf251ebf9de48c461cd58a6f8b282903d68dda516b25716981d139c69005344f5bbffd24527a764
zdbab4e2cf269be6af3b497b1ed5265f23866f90eeeec522ffaaef2ce15e293b8324af2bcef38ea
z9fed380dfc8a03bde05b52bce6cfceedd67627df1c222fc7322fb690bbd5c6c82eb0c841594160
z6cbd43ae006911eb4d9cc2f36d0f864eed707eba9c8445a2f36a2d8be4bfb873e02d8c90fbcb6d
zce7db5be76df3643710b07498f4cf169ba835e0961f0f06644c4a8a483e1c7c6286dadaeefe520
zfda94560d2631b4021b5bf9ec291399df8ee5d19eafc7853a578e3494bebf14fbbbed56eba186a
z75659738fd98fc65587eb358a66de49e1088c37948dd9112b6151f5adcacd63fb2200b8a2e5f0b
z9718da6875049b481c51352dc749d65229cabbd79e12501953038e93b35557914bd2e95cc79abb
zd6aa7ecdecdaf883ae99254dd6f5b2cd272cebffae5886f382cfcaa22b040a9eb8af67a2c30077
z1ddc82cd40d00247adec8711087276a3251f87f094fc1d695eac68fd2d76e6337718bab1bf425f
z38ae56e29d0698ba1467fc2ec9ea091dc72670cded4a37705aabeca1b94bc009c9635fa2742633
z3d5e6f0e19cfd1578e99e9ae0c4a3ddc0b1484e23cd2b2542c67f37a08b1e9c1a7183edb019495
zc6ecee9cd6e657276af3ab0d2f42ef697e1fec8cc7ac4b4700e1f7a99acfb0c9f148e64b6d7342
z2a12d7cf48e3250089822b67888f546c57c730a67afdea5c5310d4b05a53b2bd1d892e5109531c
z882cd23968b80841d1391a805a48dc036d2de7c20b43b33c24dbc35045a9053129dd42a00c7928
z6c897db35db4c3c8730625057a20fae0cab3bec0f4a057e33f8376eb216953f7fcbf817d3076ea
z84e552ab614e377489e68f0560aa90a420ce9d61e2c790720e9caf9a9e9d8f641c2dd5092fc785
z0d8f38053f51e350dbe98f400599c479de8b5170d2e0a460c18533b9cfe5c9c7aa058f77c46dba
z59504e0325816dd04842355f5e31177b0e08a82ed10260839a9d791049d1b6d2e36187cc0dddb3
z36937f6009d5d53baeddc3dcb382c52f44ef963937788ded6dff65f6a8bf93521544fba1ee7a3d
za723c2aa8c33d91265320d40defe0658e667f6c85f5ab1b502333eb0307866311d58e81af9c969
z301b3393f415f134c8b85dc7910adcb312906809089ea75edb9eb5b2fd1fbc92414984b3b2b92e
zf94645e266169071112eab2515f489e560cba103216f18d92274fc02f3405bae8bbb2e2d8e396c
zb60835b44f67701532f70d9548296062e48df87c9ba428cf82543e0ee5ceb706a70b0af9d8c001
za533248433bce36d9d434d2b6bff25e3becca00cbb2078026dd451651481aef1a92744f61740a8
z5188ad5a1a35d7b73091753cd427780a08d911976613cc767f8e7c2e473ca173cb3eee35efc9cc
zce262ead9a99e75f66d453bfc8c6b1deafced074ddaf366a585b26021757a7eefa20cf7238cb98
zb84eda14ad7adc0701cdae3b6df8d54d66e031d2c0ff3807a1a3a50a3cbfc7b6efc8f709da24c8
z98b2bcfdd3bf15243be33dcb1aca1626582abbd451bd795cf243fe22a6f983cd5d40577444d4e2
z8489f34af2eb4f87e70d4ac39902d1753639389c321e7025cdcd449a965e001db0cc8101e450bc
z506b54109f5db73635b1993c9566ba28ad04e1f6b60431457b951dd514d1411143fb29f68d6424
z311b0663bb4169dfe44d5c268740890a519fbcda46996801132601bb283e001554be24cdf6c3c7
z2b40828d973d42b28d943a32e845ede776e85987cc2c15a783818446b5e17ba628a2599b7f1a72
z2100b1faac7f0541743b059eff2fefb2e87f5eec5569bca0496eeaf982753be418419078a7c069
zd929559acbac18169e7a55a3c07596a5ccaaf602164f26bdcc00b5c253da96a667c85586c932fb
z975bd13bcd93648fc263267f01e3cc813574768572fc2511712bc958801a02be8c0ffc4aaa27d0
z6bf3aeca7aa9a86d41b3206d4da3aaaa977027317c8cdb172c329804ded9f65d5412e15675d26c
z9cc5e050325600e3115d2f1ddee9cdd4fb71a79958559e504e5bb78754cef171312869f2535034
z80aec72d72649e745a1c24ed769be215730f4621c84b6182805859b6af48a57981ffe468c1a5a7
z8fd1bf8519529ab1f2c8f712f23c48ecc2b7073fc2c082fd0d2b398ff15cf1a82f918d6a9a0042
z0cf3b6b90fc8af5078fdebb48e127c6e865f5e37542ed41b535dbd0e87b38d3e4bd3be33987529
zcaba35d218daad1ada10239bfc7e30427805f263216ed53a10eff5b91fd7221072454dc7f0acc0
z3f12dda2614b0ebea4cad6a09142d7781a850b0bb39e934d96b305062c1d2e8b7b4dc8978a21e1
z9e54ee90b4b9987514c75394ea7760a257514090d1c9e1b14dd97ac2c61ca2d6f44d3865f5902f
z678b54715ca36ed1f25187b8dd05d5b5c16c606f0c249786dee452b1287810339ee8b94514c5ba
z32f30710a671cb6ab403b8ff13bff1d70a468a243a64618b4e936241e4e647a194c3f9bed8dae7
z4ffee5bea3bcdae496db808919832a5fdbf31d6906fae53833f7f56dd38259f6ab0c1cfdba0c73
z3b16f28624291a5a2bf331dfe2a48fe2bb2f6ffee2c40376fa6ffc71a906fbc58f79cff0771cd5
zc6c9e3e94c69dbb5aa4e3775e3a021ce39a7251dcc9327e3cce7556a1facbec533c280fe79e914
z7dd9e2770d4c0893e3fb57ef2e2e94da5519ecfa7e022bc8af04311e32cd15d9d731ebed89a27c
z56e36e97ba509456b9f8dbd19dc07fffa61f358c9bb39b747d6c7a7c7fcb9f86c6b21b5c76886d
zd2ddb33960409c5f521db55dc488411af178ca5993204b53e562e1c39630bbec352d7215926bd7
z12a01f87a7ed04b2db46ef3739675072db612eeabc3e1ce5ab5b2835de5acd9dc86c01b12722b8
z83bae4356bacd1272a51ca97ae54565b48043a3c6c016f6adb4ab0a5b7031e8ac0ae3061cb28d1
z793dffd565a0e0208631e95f237eb02332e8f2d8f41b12e48c1c5efe75e7288c6e219832fd161d
z60d37a721e3483511e96fbf6cf538fc8f4da24f59816f9c3c2f3e322355925bb98387696892734
z8a2ae6e92378fdc1e5f04d5305ababdb939b62a4ab270b870ccf345fb7dbc200e6dfbe58b47c95
za1c1eea130da1aa2077d36a9c44d56ecc2036a83357b29fa4d0908981a646c3f412698e218e187
z03cfd4ccf1525b8a02017d5c48f74af3ddfd9abe81605d9cf03325e0fae08b7192280a1125012c
z7de473f95276b755fd82a62bdb12a0b336083c216e5f049c3bfe1125ca043948a2baae225d0c2f
z70fe32777aba7ac463510c172d7c56684024229862cea913e6a3a2ba1072251ab6c8520e5a3215
z1fb56553e40d56c367252b75794e9da688aa5c04b888b536fc4b2cac8e061b76df2657d4015119
z6d1fe0d3970538edf28b7d3510aa42c822dcd7966d4300591583da29d212ad50164bed72fb6ebf
ze0e18c712719457e33f7cc504cc6b7b529bffc4b7e4c4e9e6f58f52b82b2769527a9706110ed7d
za9ae581a324411aa2e6e8812dae633ca1d06439a12f38ad2f631689334d0f85a7c0836108122ce
zec50e9111461dd4a1bdb10e065fb0947b58b334174426cb4cfaa68f64e9ed1724d7928872afa5f
zfcf2c8219efb27051b72502ea9f8924435ae1b42ab532683c1d6c80d357c2c0a600b66918e670e
z328f8dd837b9e030e8da496c9ca975fd8cb1239f1670efaf6d6fd1d34c19b8a680a9e15d18bca7
z9682e7c3c54073ecb349076e86de70f3b7e89e59281dfe5f3f0b2887d98f35c9e63cb5669c9596
z2bad6758f798227b6c567d08babb5d3f36540aee8b2023d5334eb9f8205decd17d90e581b16617
z9e832d1e8b11f710dfb33d200df700302d6dd4cbf3fec48f3f33ae9294f40105104aa955744967
z58623624dd5f9b42be6d7fe93203d839f34575951d56d74d637893531747b09f6b34504d1c010e
z1f8322f6604e90829d5bf2a9181c6f2bafa3f77c4ec6dfe4c26ecd8d4fda58124f55f1e5d47e3e
z7ed93f05e3428e63d3e4e0dd6de4b6409f8a3a9bfac6135929c11db2403e03a132225ff771dfce
z62b4f45ab2a521954a5328b87894ac556a4062ceda2491d2c0f251992a41c722000afdab3aaf24
ze5a9cf91925539254d65d34a0b5d02ec61a9bbaeb903674c1c727f4ff8f236fdfdc9a8ecea5343
z1dd8528631bad8d5b737047c9de478c6f3c79f8a402a85610798ba37409b7c47011e137300a2b6
zc004085815aebd0b4eb54b0d745ee50719aba3320259b34c5813b71e157a28eed5e1f06ea50c28
zc2f079c160bd5ff186a61bd546a458b128b8559dbcb3eab2e13a35b299b2de7455ee521e534c11
z20e61ecdcf5da80d83cedf8f6b5c83f3dce5452927ebc8754e2d76213b77990f0755cc3a190118
z090caf1a114255c748079fe38a4739aba6c461870e68458a4642e43ed853902fae691805a11b15
za7257012e13eee2e6a208c9c8d4f87ca4c9f2b1f1a8c45645b76fd8dd4cb6f8f03afccb921da35
z28925fbf3ace299e0355a86725bcc9b6eea17552603adcfd69971c7714c77ea4d53f289562a465
z2147ddbaca0befebd4c12e716bc3ab6581856e4f07b480a682d3313b816a717257d8ce586acb55
z57e71528b65d2565f6d946fdc719a0f84a9e31b4ec4dad13cf9f0b108d3b7f05cb1919f35f8f5c
zb6e972201a169a54e86ad69ecec4d669a2abddcfd91d93af1ae41b7eb357af523e04e662e69685
z42a8335c6a3a07c8e3314a8ed7dc444fb1142a1460406fc6eb496445b7499fd88bfb11f350947d
z8279d62532b08a4c375c6e5cccd982054a8ad2001125bc0fa40d798f799f572b6498073876285a
ze1e59ceeb414df7d238de9590e56e5c0527552836ce83b16d3b3b8a2f60e9d6f441f0813079244
z6beb478707b9ae827bd8d6c858754d6e1eeb5e5f1e132522bee08623c8d9638b7a70091723248a
z1ce3e55640766bff7bf9a93abdd5047af511dfb7565e4f09d151cbf4d3fc830f680e6fbbae73ec
z3944cbbe6a6fcc3f46bd9974d58775bbb17a5018f407fe973d85e4d2ef544ade4db0f010f6929b
ze61abe18ff1b5ff7bd09980f7ccb2bb502afa18e9a353dc7f3f93829f09a105a1bead8332e3395
z197ffd1fa52ba5a0a0b52df8cc2c1bfd8040f9c46b418dfd41bb2718ebddf8836d8d984bcccbbb
za7b0100a60edb6fe4eb9a850dc3f6b252fa4bb0f0a03a825f0383cac8ede8b209a5cb29c36981d
z91675c20dd9fe45072ca9da5cf6dc16192b671a353fc116e7c2755cb9426c5de998114cf41ac77
z6b35a6b5435ac98a601a0d8cd7503e1b19b593176c0042b1e784f468b66e5bdbab68ab1bbda80a
z5a5234ba7fd00d62acd87e3d6917e84a61477b9871fffa5730267cbf00510b287cee843e03dd48
zb6e357abe0cc59c988c380072c7171dfaccd7b4645f8d2d1e74e192b51600460f9dc975c8a7a4c
z73b4fea67e48adfbe4f89a54f54adc31e8225d96ecc32b1d0dcea308a0bcdce9b3a03a30f8a877
z552c15b2e6074add63d9eb96d2953d4392d221aaef82a858d97a94d4b70222bf35953418dc496e
zb50a64fbb96b4aea450377767bfdc06d2b91a8977757601c1b995d0037bddc4b446acaa5d5fa20
zdaa234201467606d5a38bbe3ff43be06c6ed042e2ab61273678095b8515bb4f87f022e108c729c
z8d09453c888e66ba9720f60fd6169a9da2c05e6dba9640b56ab228df1eb93ee33e21eba735c28c
z5c84bc5b6dbc0adfe0148e7b29104c562cafb39327aad31a8647e687b5709426e0bc664f63d4c1
z5605b08830f87e3add692d9a263c7f69f8494102fdfe958123ba3b2aae5b92feadfbcd77c01ab7
z8f2d2446869268746482d7b75efc86e88ffaa33697eef95d41b0cc8108b610877210b624bba32f
zeb7dbd096362aff8ad3e96745da548baf47e8ff2d6707291ade1da6e72b9b7a0b825d5e7f824ad
z3fc7181564e5134d9d9cdbff0f296771caf6025a28ac130cc5ec5f22c65f45e011e79a9f22831c
z353d448608c0238e5249373cec8639d04c57b66509cdf02cea26d9948f20ceccec30ad5b0d35f9
z79f7aee201ace7b8e207f77a76d9b98fa2bdabb4dfd43a3dccf0f29fb96a2d994135fb3f346594
z5ffc9f20d562d2793913919e88d6bd5eb4a903bb340a94d1cd83bc350b5af0a64c7dfc37c133cf
ze08651497d350862ba0bf4535c12978822844c3164731a96e652126b01b3025f1f5aacc0b84196
zec5fa9722b8192bee518642edc4592320bd06ed47f7532a907c9484134be71c2aaaa5657c37cc0
z64aa1a9f9810f2a40ea0f8764cffeeef6c89e8244f4d60d9df7d488c309bd0109b090febd6321c
z487410f13f0462c08bbb84076e1277b925a9c8758537bf63e9bea20f4b62cb8fbeef92f990713d
z99c166c975d74bffae4e0775c8709b462895e437f00090399b02667eab21287ed7881e23cf1910
z749224f2db8386363e86ac5e9eed9796b325586c9b42435fb2aee73422604c0647542fcd876ccc
z11fcc77440a13b4b6f85baa9f9f3f6308429655baac1e7af9cadeb35e3bc63dbedb1ac4e37ec88
z5fc894149f11bd0d39ce1778d1f67eaa7405d40cb7c12dcca5603d5e0c12c761174aa348c89089
z00f14cb80a11533a64921f38a5bab669e4652d037e7a9a29a1a553a7693304632bc95ccec17f29
z9f167296e2bbb691794c95d6d6f901b3c77bc0ac0912cd5105e1f19ac75c16ac5631065a7c005b
z7fdca54096fcbb7b35ff83b2d70b311fcaf505cf9cf110827d2ddb216e94f539bb8c2c4a03969f
z4d1d348884e0861e5267fc2259a4afe3738873b651222cf8a8f63197ae3b5e93946a64067c00be
z7bcab8acc7cf3378b10862fd6ea5b6b16a72127cfcafd7a4976b17b3a8aca31f89c4b552325423
zb405a74452d9efac7175a8093fc31b7ca1e76aaf59443266fecbc94e8819d05f672e71774bbd0e
z2aeccc7a40978c1c06f093b02f53b452f1ac33664accb652cc2aba242af43c4ee102f331745ca2
z4c83511ff631e85e61607ab45e3004eb5d2a33b2b95c5a2603b9297c3e939a0633bf8564743ffc
zfc0f59688dc592589658f45e5fff55b8e6a34f01a72ea3f524ab07febbcd3445b639bd2ab557fe
z5d8c95ac064ec766a7b3dac342a2c82b0d190310a2d664f9c362482a29108ab946e049917d6b3d
zb4d62bed869b25e477c06501b1c25524de25e463a64c194227e05e9da724685aa91c6195ba33b5
zef53592867199764cec89f593cde1e84c1016ba1851962f385b525a7d7b670e26db3c745483eb8
zb7fcda64ecab15e880bebdb8add542a33d01aa83cb5be593aba8d3f6f97a7ec06f84b47f26973f
zafb6a4302ebbf149232356d5c5a73bc02f5c2ed324505adb9ed10b9ded1eb5ac2be336553b6c8a
z866b6480eefd668b4e10f8a22097f4b92c5360ad8b035172d3bbbc27606e7673ae042aac2a01ae
zbe9302488f989ce00fa18dd2f9895828ff9a0df8227fd1657115c7310b80187c9dd9a9a9b96c46
z874c0ec7bc7e581b4ee270c98dc906841692ceb73218a67de161ef41161bc12ed14825a93cecd1
z2059aec00610af50c0ffcdb5de36c3c43b02df183e4599e2a029b0185ee20746a25e13f6c00549
z9a363cc2e123c055ab09b4df4b78e2a12fd9e751b34b2c8b89658b72ca7d9e18119f72bebcc9b7
ze90a8df2639686fa88ea35b5c529c3f5a12e92681b2129a7771d956d44222ba2345ee53c47dad1
z06d5a15fd38f065132210bfc54b2e97d4892164f4013f310429b617fabe76d7247e395afa3715a
zecd6a228dae30a7c99e924182bd150b954e516a20683e74b8cd9cbcf956f4ca51f3b665780608e
z591fa50469fea32c930b270307d57a8277454c27e0c926429a205b9c67fa7fbf3ddd6fefe79f58
zbb160cc58a29b3b3ae63832650aeff9c7ce554e6601b8dd25f88b43b8f8c9be54052f0b4746bed
z7a0cae2242bb3342b4769b50479566a9fa1fb32549ad57b6c52b3524214e2e9415da876e3b720b
z6cf85f16b4be87586f936099b2f983ed6060f0b5572e48e2fded194242fd2e3a32b2a51165f2aa
zd2283f1f074ada831dd4815423857baf3ff1c1127efe4716a6171318f0404e7a5e4c095b16b429
z5f1e3622e2b96f1f0743ede2db12cc1b41b305f48bd9c9a47bd2a9c0b6d159926ef049ec4e1545
z5fcf20e5a145864490f34f9f126f6375f36792570f2d0f8dc0b6cffe60e67a53321a2d28cffd6d
z130bca7d7a0964891b02e885c8429a523e3052615b4b7791b05fb9464bad2a5770e216b52411c0
zc26d458d40f5060410acced2a4711a76f7ddba667fd192ed1bfe7dec177d1e342165b1fe6a5d74
z909656e0f6393e4c38524ce5157977520e9862d34a9e378967115cdf4d8838f1e381e165aab05f
z1ba4fb21b4bf7139d51a11cbe2828334511220bd1666d8e6403102a0388f6e1457824977c87cea
zd22a07390ce168f3b1abc0be3659b7ba5d6a085b35272d6f2cacc99d077c5a68defd27d94d3e9e
zcc70e1e6390da810842b3d5924afce893c0e6f2866a56902468ce8c2b7e2b2d059f5bf1eaa5313
zca7999a07c4a5525db96356d0524dae583dd709fb77367242db003753c69133223f0b6199620fe
z0f3dde989e7b9a66d4b869a789713ec360308e6f15c7d4383d0114ba52a59bc7acc17bbf973f79
z92ac53e46a74bc5e94a33e1ee29de13cc3a95a13a0d025c5c646b9a7d49f84d005ec85de0a9bc2
zdaf6e38d689b07845da6ee219bf130d7846dbedde03476a9ba4afdcdbc136902e2c1150f57be40
z617460804c0478ef540a1edee63b99945f41623907015085f648e327324acc739f03fcc0014ade
zc748f965b208c69b7e8fd8de69c9a29e7887ef4b1b61b152769b6b904d255764e14145e453779c
z27f42aa55394ad8ec793e587c3e3154bfa02cb5caf9b6fd4b70bdd8afa7a2fd3c15861ae0e65eb
z77fef8ee482a034407edd2caaade1c3c8eabaf1ad63bd2c20bad0d5f1453fc135a77b5f21f7579
z2f6c2d6f7c6c793f986a0ba8ec421efda9f81a2805cb10893f1f6f8963daa957f37a8f7276bc70
z81097e7f5c51c1528995284582ca3d2dad64b5ea2ff4876d310220ca28e77ea308f47330c88828
z9825eee8d8725103c064ae063fde4df61a0755b34b900424170b4ca3610c0e356863775e6a7eed
zf0d97a90e725c3173d3539ac298b30f090447e11ca11373e970ff629d56f2b86a0a46bc5efc83d
zfe64d3c3ea2391571d0cbd53d2e99327909323d9e9f8e32e76c6d08580b1b4cae7e5da5e251c3d
z3faf20e9519015994ff20d5734d2fc85648f7f0daddcae55581ae9aff06d6d517e651084cb708c
z6375bf0f26a3845365c4d0b6446c75f97d611241ed3d8b39fb1d0e131ea763523f102c53142ad5
za7b07be4fb538bffef764518f158b8189bc20dd37d266584d8724a614fe3554c5ee77d782cb2f4
zca012d134222855dd6bdeab8caedc7889e2a0a4f9451aa832e1cc258da3cf7a22b7f9fe703852a
z4664f22fe0a2f8b20c8b1fa619de480c9a1a6f7435d95cb27e9c83c0d804f1454e7787aa156eb1
z874a3beee80ab595231be4cc3ff475ce19d8c85af2348a8fc0e6cd83a6bb7dfec16b2b624eb736
z172719f77b5037909b86a0a4495a27963dd04093988086f0416dbbfb6819c4662e3032d8344d3f
ze7cee441377a805109af6bc02aa679819eed1a1a4e62132bd2515d3ee58b8a041a793899eae29e
z3cc0d31b4a4f64d12c65c75fb507f0f196dff3ae6c9cb41494907e191e2703354c828546184373
zf2a7ed054f7aaaca4c274236629a1028b692ef94b045dc448ec89a5e0a95edfe6b23daf4a961c9
z02f483a4de2c799dbb1195b4a96852cbc2b09945f43e1a306c6319e4d1bec9fc0635e6d6108d19
za7045029346e9466bccb497a1c1f694e600aca7f77b58fce73a50590634349e2ccf999c9c7d93d
zf14c808fe74bbfa1471ab87455dd7f41c0df331d8cc04c9a852feecf3c3436a8c5178901ebc73d
z08e9db16ecf66d309cb021ca3c1fe1a285f86d03bec6d60bac035d1eb5fd12bb2c9328dda910c3
zf8280637786a69745ab03c238425cf4071d16da70de55b38acbe332d734092121c85782982a36d
z728587d7006e58cdd463446d684cec6156694af6dd3c7819388c82e60532509226bfa93551cdc7
zbc71d1a4e21c88c2ea4cb504b3953d0663c7967377169c11f225c975ccc9bc3a17408d053e0324
z895f017dbf19a1a64641bbdbf55e2333610296caf804517ae47bc133abd7879593c36529cd1288
za5a61d5d8021ac7729af53d00c328759e6b318e2a2bcefed0440578f100a3ca442a8e8ac6f4617
z78e0ed2b43e27128e4bd52bc35dbe77e5e9233b5ab64913faef6bf4541aed9c88f2a588ee7c9cd
z008f05030a4524b718dbb13df131eb6700ab243b23a1b02486dfee9f57af84364f8e8a916d5f79
z38d790ae7362d08e312b4f794fec02541dbc909f414380ba13835fd80601db62be473c9b3c9a6f
z084b4c5b52bd352f77904834ef202fef6fd192a5aebee90bea0fe51adac9b490e51f38267dc546
z47a5ac7953a54c479a5df12c35ece81c43ff274ba3849ee79627f9624d8157091af7dc3cc3c0ba
z94d9d6562ee01b90d52ebd1b6bc703f4496cf5d59d211347b68b360caea09342a7a7e2c724c702
zc6eefef9cd144f060e2d2dfbdaa0b7f0cec620b57218dc81beef9801771b7253be3111003bcb2b
z45e2532b52e388ba48d201a68ef790ac36c928a03e727e733800ea9f9adeed211f139e6fe460ea
zb03bb3ffbdc8f3db47ac57288fda7f8ee66b67d1d4c072798f8282962842b79c32c134ee7b25be
zccb67fef3eea11b44227ab5df26e7722f4df79298026c099b67c9d9994c464bc6d3556a83427fe
z4d27700eaee53c39dc69e194f83cad25fb33044352391826789849b990a8217e5ca672e6d0fb81
zd50e93fdba409e0dcfa1c2e715dd656778e42e3f27cdf388d5d215e2c4f36d1c652f4e037f1dac
zf4d2cdc2557c931ed5a3b213383d88a3628b0e52e18961e926a4633d666c05b525ef543db80401
z8913160517f4a90873504640dbfeb555752fb86f9e328efdcf964d329d67597fe5ce5acb39fe79
z01ca44dc7b8ef183d5512fef1c8a2e3b0d98427ce883262fe0a598b0243eae4164089beefa9534
z50e8e8d75453543e5a00e343ed11f8f782148c0452ae9db4822dd6b3a180f7f6d3046910d4f0dd
z62b4d73162f12bde82d892029ddf4acdb106f3bdfb426d307459f91e0b5943d8e51221c6154da9
zfb41198529ef8c181e240a0d926b09c40a3ba94e4a0ed756d831d5793c46a21d51f57524c98caf
zab753f52aef8fbc5a703be56e90d1f9c3160f5d3475ccc5d66ada325e5330be13cb6ad58d2d467
z5ce09a000d311d1ee40268ac3f1a6e7f4b8dea59f17a6a6eec64bb1f8617135abf9675e8a40d0d
z04ff50b4ea78379ab5d0dc5766288e9df82b60a1f30cede613582c28b056de16b1874990fec4a6
zd4dff4c8fcaf6093452a3dcbf756ca3e23edac35a9e5456a58efbd2a1854e56c5d14f3dd0b6f9d
zb514f7a7142d4e6bee399dbeb2db189fd255f3dc0ff5d2accd3eb58d370e4a4f9fcbbf2fd5a588
zca3f1766c8efd7d3ad0a6eb9bd8e3db23a9e8f3620abdc4fc130b1c3292ba62858358caea929a2
zfe4ecd06ef08986d4c7dcdf2c0bbf96e5549427eab22f281965fe653ef5303188f4394ece7e521
z3522378e0e4efa14906623e68fe2c648526e7164e060f1ac864945930cc9e2e2631974928425aa
z0ce4df089f988905a9629aad283f9b1a1872e621a6692f6677f6b89c3ea3b96319db7764064c69
z4f8f0824a27d5625d90190289798b6ee14d97f51b5e7fb74595ce0694bf1d6c694a81f90c5654e
zb7bbf32c5a8b350400662cdb747fb162946078ce110d47e11617d7fdaa95a445f18c7d82e15b99
z13ccc4bb22bdf3da4b27824a48f8d65172691185c13fb3d68d99ed9fe0420446d3191e93303184
z836d39e7a158e9485a916777ddfe70eecf35c7e430969c62b6c6cda0b7651c18e6cd1787fc6e1a
zc08d8fcbc214b0a0379b2160f2fa60d0138f98db440b6b94e0927bec348f04a5c7a22543ba5911
z991b0661054b7372bff602dc3de04d73eb730b2d2ab065b6c3bb7154ea71ba748ecb867a452c2f
ze6f7c83a11fcc6a6b6529c7e6147049a263c993664852535bcc9146151f7a903e5640072bad63b
zb000ed855a13e9244cd4741e2657ddd1cca14220c04c802a41f2460c94da2f261ba9c1fdc268f5
z98ddfbc5066b21b38998a157aed06f48a0c5252e93ea80157499bcda0763f932e0b1e0b77d373c
zbd18e5816a01c7bca03da47fc6e69f4726a87db59097563ada97d92ddd2c8776fe5702f1558d54
z54bc0bdebc0e09e677c222168d1b5941c34c8f294ef9ede9b8867d854b3c1d1bb0f9f12b9b592f
zf2de4973a351fd1023b7b04cf3c51f99bec3628a1a0600be8ce251cbed8735b0ea6b1a868f3c5d
zc316e855bf698175aa1eea68af0f9730a939c8fc1d3370f2003b5b068088e27bdd93e40effab31
zb28d75ee1403dc0ce0ad37b02d720bfe3c5bd885a9b83b4c7b1a13aef4668b4996e50cf07b377a
z93ab66665e5e14fe83346f63a80698924345371ea75ebfc7f6aecd4b53c765971366eac018022f
z18ff33dc984c17a9e12e8e20e1dff280f489abb293688f8cf4f2b6091b3db8bf72cef3c17a5704
z200475253c570e72561e567413e6eb947700cb27af9d003da4c941789749d8748fecc63bc252b1
z2351c08a04f351c5170c4e1312a9c917ed45c64d31e27d02e36a643d56ef94ba14b3f61ca5ddce
zf8e4934d5fda0635f145051204ff9ab4f7793c1b5449ce2cebcbc60e1b320360d7289374d48ef8
zaf134bfe534bd9bf3d3b9dc1b1f637caf3610d81debc0461ef8f86397ffbfffe21512393d80e70
z54ea706b97fafebbf776a296c1d3c6bce849a5d308dcc9cef03f5137b5f902290659b780734e51
z44c8d0ef72b3b640b1d9583758f25c6e996a581a7293190a0e178b810fcab3228264b8c9f05e32
za61163a89c3a6eab3ee598defaf3ddaf28662fda1aefc0b8df1bfbe6544297e323b675aab9639c
z4989d9cdeed2bc09bd0887eeb071f005a5a1cf1756d5f4582a7ed87afffb70f3d54f69705842ff
zc47569bce925112cb7612f8d40b363880ca8d1bc26a8d0b15168abfc5793763750bf4b80d6351a
z81a0c34055c15872ca7546d8cfbf02a3ed141685e1a962a50350dc304663e111fbf25fd53f255f
z0de00cc1483477039e9475d39a3709eef03abce4c15e983496216a88662ebfaa7ab81754c3bb2b
zcb3b2ab1799cd1ca1235bf772573a4af969af6c3c530ced03bb0161220eac7251649f707681693
z0590c2815f5d7b7ba62f09699718c8c1adebcd6d35e449b018aef546afc5ef851584295c684151
ze344b954b5ee15e1eec604edf1811d81688b4671a52d8f75dd367abf1c13e636681e0e6ee3b142
zd5534edd6b0426b6dddaa73d5d948b89d78759d50f3ac3f31b407987f805541cdf0211df103280
z2e9c7874ed28e4f689637fa54615dff2ead05615e79bcd03417fd96415ba5c4b96776be96068e4
z59f0a714aab176cd536d6003fff6d4576204635adf3f2fa2b45f03f6046cc8c20fffbd1c2be058
zb7f3f0a99251a02548db0ac17b6971be1085fe881e9a84313c252ae1c0c00b3975d1599d0b69b6
z051b878f77327805fb4edb1025c8320d1eebf1cfd03dd211a9d8c0fbc5ee0f144ba3e9f068bf64
zb578380d8eefd0b3b089a788b8d430de157ba6445a0c3177eb3130b3d5206936e4f6c6402cd7b1
z14cbecdc7beb35c71028d2dc6595c4cb2ad83867757512b34ac1bb7ce6dfa967850f9bb30767d0
zd7629563a518b17db049ef1164579839464b7a84ac0eaad503e3da6e027114a4d0778726da2e48
z39543bf23f5c5fca9af62ad59dfcf727318499bd6be89f8d55bb389924dd3a3f6cbe5af0563210
z5638207b9713443cc480111223f3c712a03a5bc75f77ae2ef9a272f23add9697e7df12112f980a
za0f49eebc8e91843334108b18bd6da308373c33a9472690af45dfe61a4159a6e7bde7db2950af1
z3c03be8ebe0b3d11ebe0e6b6f9de2b534700211ea33534b6e64a499269ecb7d1d00058f50c174a
z6a2321fdf7e7a8b4eb569b4fde2c53e44fdbd43034a0fa0a011a224a1a4b3cadc9ee1d64c4bf8b
z0fa8beeaf51e20223677eb75d74c9b82aa5b1cb7e8dded18ee08f738211c987d84fb3eab9a8bc3
zd96cfa619a7f729dcef67270f8ebe56e94ccfd0b9364ecfc0c1959b5120d588e2d3f7e0075ee84
zdc93a430e718057ec3e53e6b2b6798ace53c63b17da9f32ef49a2811aef4ab0491c3089284b26c
z32388f79acbf402094b6d7aa67a0ce2ad1c956e1aac9524f4d62649309f0aaa156b867d80b9b1c
zafbd7462bdf1e7b09029de8c49abe5ff931e0ba65ced1561a0926588048f10e78ee6cdbf0cfbcc
zaa4be09358c2470bdb5ae683a4b4399ea56baaaf0209f59f5e75e952e0fb5fb375428cce3cbb89
zbd560747a39c0568259a35d1f102bed756e39516166c310a2c098d55a16291e6bcc29cf0497ea1
zc3a873d3fa42fc92d5b4e7a322e55b88e0edb050e187b49284249cff6f81e6e836fcf00e612be8
z5532bc3031cc8635240c0b4fc840b22c5e2e710f3cd6d96ef398db09f556e5d92fcbc1a1471c36
z567acb59f5d0985985e6a6d46387c2e920bec12e313ae2cb414edd1fd86bbdcbd5103b1a6598e3
z424d33947ff06b7a7c1530718f444e669a7ed8f912f80cac956bd88f4524dd2ee3337196799d08
zf5dccefdda34e6eda20bc87e5164e5e2d61b1847b833452bea749d778e3040d998057c67d7278f
z6d331148c852afd013572fedd6a317bb4c982aefdbc1f25ca42cafef15cbd1350c6ef68806a9fd
z9e78e84ee0af2f9da72fb6091311a43cf56073ea630a0f93bd549a7fa029f71f4cf1072aa918c9
z04bca4770ba46b240c5a858480beafd30eee6e42a85bb3f809d8f726d85b6db866dc00c3b3de23
z891fbf8ff18e9a654f01f7aecd1cc787c1ea5d0b94ba33230d31a234b3c04282932cf06ed91880
z40e54da1eeb7d6b76249d4c0c76bb8b7b04754b2f847935378a3d90a721f004b145f1b0e79fb1b
z96978e1d3f673f7e60d91b440e3f5e633f9f9d20e4b629bd1caef7ce7da2e9036551517c207252
z373793de6abb0c129ea2614d8e6a81ec4baa9e1c7e376e76aea4276c8dbde6b07940fcb6939090
z719e3d764f1f8c614f3dc57e2480ed4069548aa37a9c9bb4d61553a443c8bb237714693dffb1d5
z148b12eefdb966ace07574e8b3bc6fdf7cc262f4055d57a12c91611b401ee8e767cebf09709886
z7b1fcea2537240f6146c3da8f053bed42b80c04dce867a4f34f928a25b424bfd5cc3bc6cefb042
ze497a3b355a69b6a1ad1589db1f25b1020840c4f643d3f48551b0a8db678858912777d1a90e99a
z2b5f74a13fc9a37ae9d227082acc78394d589eabe77059943db61e6e294bfb89655f7a220e9651
z8d6bd6529fbb08b429133dfcc9c89e55ac5a8f1ab7f6781b14d86b34955ecff6bafcf8221c70d0
z69d71080fd1d3975c30bb8d71ffc689ee593b1e24113876c9fed46e5c82f4f5af9de43107bfe9b
z5b20a72a58406285ace804c2915a3f87fd617b846e1380a7f3039975e0789fdececbe049a7ac12
z8ae7d133a33c5b0d2c885566a43aa36af22b322e5688286c10676b27b7d1253d04ed5a0f19ca46
z936878f617e15491063efe3658358c4b43b19d4c1b934b7e5c42e04ecee2c5175b8417d74eff7a
z645efa4e7baae8da3cb327abd355e267e1c83674e57eecb9f9e76db84b0b9545b9a2939b47e44b
z119b0c09e2271b8becaead7b60f4578b30e7245cdb0eb2e65be2723bb3f32541c66d266c6da186
z9c9badcded9c6eb21fe40cefa125c239ffe9ddebd049957cd80b2a774c9037479f39a8b1b132f5
z154f87f404b7b890b466ae098ebdd9c0cebd44c740ef7a0d37e2f5bbbcf2044bde915bb03dc160
z833c8aa3dd317cd452800dbfe1d2b7f3cbc64fa7a384d31d6c2948503a3b67189569d68dc1401c
z8a062c9f067b4a5a903962d6789a41d8c8e0d8886141dc7d2a9270c8600ce578ac1950747cf295
z58ef0ec10d7c58dc3bb2f9933b1ab47b445523f20b758a2c68b6500ade1b9347d6b8bf756baf8e
z4a4295d17afd6b110bb935e50ce3340d849df5c4bf0c6402549e3a75373667241c1bdee1b7abb4
zf7d3e2a429d112ab53d406740c781216bf5e82b1da0e51cf0f355820840dbe5fd577d181bda78b
z1c86516c87ad18220b4fdf322f7bc9f5af499538688012a2152c75d00de3da41615b830138221c
zfc3befa7ee086c33600715ca8e60580e15d0f82b06c41db80c017362be6047a4e2ec075d7929e8
z44b0e03edc2875f6641e0c66619fa99d582a4141c60e4a5d92d9800873e2b8d64038038304a86b
z29743f83612ce329c5d51da25582325b0c1c2e87d4bc6257597ebe032cecba09e5853619e13944
zc199b3e379c5fd58d6e465d7bfa0c04630f42880e34892cdd76302a7a4bc3df54de7709e58909e
z4567f56357598a15694069fbd8d5075fd5e7d8087c9d3b46cb4617537c31b8b9c544448b7dcc93
z99cdb0e0d0f62ebddade321e0fa0f24f0ffb638eb4441a718df3bc9d77a761669a261c817fb535
z1e7709b775102505df035ea73c3a91bfc2b8feb4972c7cade206fcf8ef769ce8760ca5504b64df
z631e95129a404295597a77fd8ed9e13fede412795f4dbca9adb16a2478996f0349e9447c1da8a0
z7d9392daed8ccdcf767fe15a2c6a78f92205731f56ba691e80b7406053ba539539dc1eeb1a2390
z08d88fb4b1ea98a615af0e606380a0030a96ac38ddf3b56c636e0ee93a02453028398466a68178
z89aa21bcc42a898d85ed6c3a6d22450dc3b30ae1effda4c007326225ca29540b15dd08f2f3cac5
z8f9858c80d6a5aa3b5f88186b3216321ad2ec7cd0c12d845450e5c9fc3a8f9c6f44ccb99fdaaee
z696b1aa1c0bfc31920c297900fe35ca3f5b760e64754c36665d01c5e916cd15ad93a22b7b5ac05
z9eaca8bed028777fc3d0799bd9600e8614f6e92c9eb5bce91838e632d8a7c3f92f488dd583f4b2
z3f961029383a76ac8e55637c774fc3f9017063bf39583e050bfd61f5c359789448ef9d62241adb
z7404ac3ec376210f3fb4b309fd922ed99902cd90ea3074ace1a5a8e9646b6109cbf9eb7a73ae6f
zd75110ad9f103e8e681ece12f06f22e729585b8ee6e441c89ed30efbeaa8a27b1684a02147ec53
z72dc4c02a7a7b68157305235ffac8c3b7fc0c17f1df8628cfa9d2afc3f3ad0bfc6a1fc45b0c63d
zfc65d4d7847ec064dd5d7da2b366f970c5c19edcf42bd059519985f2ae96f3dc71452036219772
zc26eb4c3c8be69055f0d123827164e254be06302b3b993678b2e9c32e3ea7473ff46c8cde48f28
z831193b0dc49c44a6f363158a64308ed4a419bd2b4c2d68d4a0b8ade0d4ca68fde48edea5b7b40
z3148af0db679bffb8e648c111323a146d7ad9bcf891a6a6ca5ae427f6c84f7f3439ac9e09f7fbc
z8090324e23a1c7d61b34b4231bb8106dbceead244fa1ad8ceb977f4e80459b0adfae72ea4a4218
zfdcf9052894734eecd03118e88c135deca3f7ddf55b479f7fef7f888a946a63f00a7fea491e436
z089b59330499bf56b6dd80fb25a8e01d438c944e72e0faa4c4c601e765583753f8edff03ff275c
z1c2a7ce7e1a2c373fa2679229bee9b203000267aced8536421a055e58c7f2831740b186b98d8f1
zced1d8f7957e3d8b2fb71fe8548308047f71e8f970fe05efeaef92e9c171a7c74baf66693cd92b
z9ea491aa5b2b4fb343fa12662ecfec35022346e341f6dcef0652d0acd85a5c1e6afd02895102e0
z1d1f693cbe7b62922f89498714fb83f334d2ab6f497cb2f6c39f81b6ca6c94030a35128d81dfaa
z3e76987bbe039f355cb17f1a6469305e7132aa83dd9fd05905858daac2cfb4ce2279b4237b182f
z8da6bdd5739dbafa458c0e68f60005487da503801bb3a5a2077f902ba40d7fb61c5a1858b60e76
zad171fe1afdf5d298ed3f28b94b8bb3d5a279874dc6a43709444e360ab7d76972d1d2e07816b61
z5ca50695ab28b37dbf65ac566e8747ef4699a3f6ad5651b4d27d68e65e6bf449102f81798ae893
z6c8d6f4199cbe6563ab29b22e873f160190ff66c05607e769c10196009345a84968cc261b4f810
z0008d287976e85d52abbe34b9f001217818b6047249ba721c0cb0fb3cbf0bc4630e6327c27d532
zc7e9549cf74b8d19ed645c99866167bd26ced1202da67b1aa3f53479be7b7b300d0aa7c09be899
z774f5ee488b2e4595993c68576b908472f98709644621cbafaf8d1acb092a38a235b28cca9b298
z4c6f9c8cb916902a55dfb2a6e9a604c971b40c60ef7819e07764d48e89327761cb4546a404e98d
zed97d62972bdd9537d5dd15dc415d484e883f7bdcdf4fd7db29a85e0e60c72ef16d51a65f9d89a
z4f2c3ce5288db327f11599dfb05a29efe6f008a6de8aba9618fb26cd9b59ff144224b0d3a27512
z67a533538282da3d2a7354e1a441f4066e413dbddc79cbbcf9c0b6ec0a2fdd86324a97d6779b75
z627d0dbd884283c4f8d0676347b072bad0a9538661e826dd34dfde6eb5ce7bf2586cee89993ff4
z6f3fdef05ffaa9f7bbf8a43c91bf733afebeb7dbeeac6364e5ffdf547441b0ec5b8a0cf10869ff
zf5440fa207070f81b4ea0979e7290141f9b8ace53f6683c58901b986b8e9489a3c30205e4024c0
z7ec5f4128ff563b56f0eb204b4b7251291728d89e6a08bc551d45adb4f93ef8318d9599fc244fc
z9353d8457c36c83ef98abc7ab35b3ed854ee106bb1d185dde59d3013b2bfdf5726fcef85d015a8
z6d28f9cf2389757d644a37b9ad858c6148f283f1363d43f8d40f5b18ac8438b55509d3fdaa49ba
z11fda5efd5c26026466f07aaf16393f7abf9c917471c3e8bab69ed56b4da5cda9cb62fb1e2eff7
z697e02e673d415ebec5ad9babb407c877e3a960496c5226b97b490229d2b4881055fd843b95e4f
zd2b2c01df6f9d80d87754f353eee5a3b5119099ff5348db820f0cc628423840ad1a7c5891e06fd
zcc2c31240b459dc377199b705f3a64e64a8f3eff0aee675bcba80022136e87dd5bb8f7b1810e94
zcbcb48845e8114b8253140731f819b4118d8f806eb3c0f2bdf484f89cd903074cef8c91f803086
z548aae4d27b84b4df697328de408ccc9fcbb3ddeeb97071f7fa12da1a6efcd97c4be6728f2b52e
zb02a34bb11dda2a5cb6b173425dca65014a77a7e9baf85ac9759c2a93af7b3999b5e52a9a1e9c0
z4b52b4a74ba76a93c19cec632ae80cb8128f6dee42c3989d785235220180111909a5ce90322e55
z9776a901bf1fdafbc48b7911d2883230fcf76d84f2ae06a6f2397d1d23a9eba1937715e3ac3374
zb4f6c9dbdbf9e879932062d48bc8dddcbf14cebfb046bc1f8cdd18ce4274ff5f6efeb64bfee678
z239c1dd22e6a9925650b03d737cc704641ac837fc06c430c3c230bb4f81c76541eca8732aea8a7
z2813ead0f4477490d7ccc9f7fc39510d3ad06c07eb842b38df10f71afda1df04cb6bfd96397f12
z9d52a0f7fe570d10a22e0b25e6f30531bf872e7745d8cff085d55ab04e2dea2d0fc552491d9501
z6c806c4e5fc05693cf586a4c374dd34de3c25b338d009112dbbc278e66ac7c363eaf331d475d76
z21878801857980a649b93f65dd3e07e9647025351c373f5e90b55829293614c5c572163f212852
z5334b4dd09feaad8ce6e008e952e9ede2154c6da856cc0b8fd63feb4b6970258da13e998c37339
zc7c2c96488616bf825f3d077085590d9dd7c25b9cc9aaa4ab15dd9679a1945889ef3b937f5bf06
z3d65358acdd80cc92729fccd5e1667bf2424a6b6e8884a4667e5c6663efb811dc3702d193730aa
z7647a2d3bb9425cf5889665fa866611e252e0f5f821e97d2d0b47b8658d551a83d6263b41f673d
z8ae6d22f88bc22a54d1e5d4cf021ff8a87934e39fa18b48e108fa397c147cb19595a5eeae2e25d
za20c5670c7f67e569bcd51dce79db06ff3d5de0ad700917d5aecf0ca466e9096fe156f37bce624
zda675608f8a003cc1b40fda57a35480a1deab7bcb0a85eaa9fb19c0cc2c06f64480b733fcc1801
z612822a2845147b724ba3ac79b582e470377f1eb0eb19384324088f42f727d521a61467345bc45
z5dd1694ba08caed24eec41f2a256e41c8904503b1748b7fbf072beecf6a276693c9c7f0f66f3c3
z15645b248100011868b36a921fe82a92e91941ace85a7dffdc5024431141583212e9bf752c9c61
ze40b32bf05d88b6e783007de88716191bfbd77f882eefc726247dbc71b4331636b6513cbc30db8
z0b9d9db66a7cbfcfd6fbf703677131f36a67890f9f6c6188d2652168706fa735452496957388cc
z850983eaa11ab90c3e48245e8c75abff6dafe448a6e25827a07e6523333c92c13c29ff8b471085
zd0c32a6be0eb1f2455354a1d8dfd132e1227d42b0b9a3bddf7351b26e4b7edc7c552fea5c4c784
z7b660c4e7bb73a748c068da2e9906dbb7072d125664fb6bb84411613789942a964ab065144ff77
z38d915d70116710e0f8f118d0d99ab1b988874d9d553a90323f4202921c2d78c0690fd62956810
z9d6bcc81beb2c58a551fdd7863efb78b6ba2a7c465d789503d7f84137531f0fed53c8cb0971bbb
z15a34041e917f05b705d9818456c29f018a055df626a59880f70d69a2f048615ee48a7fb4f96ca
z319d0c1e8ac97399eea8c0596ecd1d7348cf1c15762505f1accca1a95494741fc6476275772e34
ze3e59b32059129caf920ca5c09cad660687b50626d639e41878b272ecc4148f30862486ef22b29
z299e09a23d78c814e3eac2e7d9c6e2dda028579ac0dd387f21797c391d6925525559176772c87c
z8672f5c1b09547f7ee5c725903ae02da2f094dcb6e6cdd2a25a2b3ddb6edd171e2d2861af7300c
zbfb5a6209c87150130a3023905b17ca910e626fddf848fe26155b446142764b5bc130b6fb6d51a
z611e2f99928151656911ec5698cf7afabd5d36cdcc25b566e6bd043543352c265fe0b99048bbb9
zd94115575ea04ff79e620fbb2659e488019ba5eca9adaede66d0e186902890f1183f2d3a5c2ed1
z1d24d14c61d627c49fcbe2354abcdf63c7c6b1543086547fea71293eb4af5597ce97602594f95e
zc54ddd92f18d788219d392208b6a5958baddb0db94159bf2a3c21890e0e0d59c5477d5b39e3e32
z6d3d9bbf5f8d6b64f9cbd16adea553dde056f95cc2627fbb1462a4973bd8dd75ebe3c7d14d5ce7
z95d10b725d28e4f49c91979ce571532038d6cfcdbff17d9b62fc3761e17e3f0cd6b11eb7e26380
z7cc3e7519790661f27b1ecc7a6b391d4cae3d1351221eeef4b7a604449906157db5c289b5e66c2
z96824c9982ea0ac5a8b0a2661b682dca5ac8db8a279da7d32a88f4e8eeaa77249d189b2344a1ff
z19ca326b32ea08e9eb214a9c60499c248a4776622d9304f52b733f116291fae17a66e4b6b720fa
z40c9928d1d26348a4eb962f1d25449da9e0cbfcdf764b8356d06ab12ec44c54f217ad0a10ad061
z991f1cda9c11cc39ef5aa9eef6af4c0dc9ee3963e7919dad4e91b6bf18f73ad749a29fd580ed33
zb8d21b30514504357a0033f837260090ce12a5eb9eb30f1be26710d2d2b3cbcaec978fca9bd8a7
z6ba95792e9f9944a27240fb818b22b68fa02ebe0e4f5411009bd4df7f77f86d4310ee908132954
zfc832ca481cb41f1e10bf9b51dde8d08240a2700111b6cfa063a5fd77e24a2f1d5a01069a3ed27
zd3f5e035b8b122df5f8cdc0c928e95a2e9c59ece983640c59694ab2abede00945a6dc5018cc0e7
zc4960aaa1e2c0def3e9d1b0f83ddafe21f51b43baf3710e4bf76f87c4c7aaf393d966d17f64616
z76326fbfce40887c3cd015a74daaade27488c41a892b85704c96c8c8c0486dd148e9cbb242ef46
z7bff2553b6abe45920dc783f8c8a02bb2744d2f7bc6d45ad81a9d8a6e58a2ab9e536020f829d3e
z4ff82c5f18cf4b65850bdbbe66927d394ff8781255c57db8027ca731a6e225ecad91da919a9548
z83188d4d27586a56b78b1cd5e467f4eca9ecfe11da002119d6fd913c7a71ab93a4f51ec6d655b2
z677497e46b7328e6ee40ac6bc4b34bce70aeed288957973aba82f0ba15f870bd756e8e779883ce
ze17d6c76230c69aabbf31c5d864346fafe722bc8c1ab3baa38bb76fdd5e648fe00917d4f6d359c
z134cfdd96a0487870e0922915e9b5c041d776036a72ee21bd7e340877c36648b7671924f573168
zc442dd27072d243802fe4f6e2dbfad50ca83cd34f3d134ed68a77e6e5039e43f2efb9e30b7303d
z1f186f6d7c8fcb852948afae79ca0a7a1c2a21517b6775f3571f212b1f0c27e05cb15d386d34fa
z29159dbf3804b808900564f1f60beb6ef5c22b6e32e72bb83da6f6f9799d33180b77279d15ab6e
za0400d89c3d2b513ef0e29e3ae8657703936b09e1c8de9433d368632db32c0f4a745cf398bc20a
zf2d158e943d5d02fd7ea31d967cb80a024c0652c1faf8354189d9c0e214d4434cf8213781bd5ba
zd3c701a3035fbea2953d05f93e528f4ffa26c38e4e906e644087bdc77e17a8c02d5b1d1869f613
zeb0108dc798feb78c145750be35c09e5989a384e80c223e81fad694ab462266502c732a8d7aeae
z635a74ed68ac852824371ff08ea32d427dd0f7981262911f517bec37c680363f753d4374bf1be1
z756b554da55347210c0f6e0fe7925eca5f5055da2de88b6f1d8adc13fd19b94d200f3b7144d135
z05679c4d8c66872d4e468da279810fc6b75b97d62eb18956541c56af0602b88fa65076d83f197a
z34663b52238d6f8af8b7b6d3458a59cf03613d74c9f78ebc07168fcfcaec11e5731cafdc98bea4
z60d86f16784aa2ffa37e8aacfe3004bdada6b050bba96c5ebcdb5060f54e9e72589d67bdadd11c
z579e8f7ca53014bf709d09a61215d7141471716b4ef67f17305eb405893c7d79c2785e1ed2b0c7
zfba5c11a7765c82f44ce1be79c8057d2717782768e63e736eda1d0c766b8b1c31db9d3a6691a56
zd1aab42bd3a181634286bc4fed571b80a4848f78baa3ca676feda4949dae6ebd3eb15364371dcf
z6512f72f3854e2b8c0ab2c19a67da99033f21517813cd9e188bed92bcc989ea8d2fbac9a881522
z0be9fc396cbb1d0e87c1d5d9e2590dcc0f102fc5f08c7bf6505e96818b65e1386bef42b8dcd21e
z26cd18884a83e746585dfe44ecfb0cc5b2c408056fd79abf18a1616cb4306b98c962d70f8ae004
z4d0bee2754b644f5850ebf95f71d94cb46af572bc558091709c92f662756763f12f2d6bb481662
zf270f5e65db1f93d9115462b98d8992d35c12a4acf085c2eeae2469679b0be52271ef73e51b6cc
z56ce41c56d1a652fd3d0b06e1eccfaeec01143e6b84d0a26383d051cc815ac7696157efe616a8f
z8c959322d17514624020a66bdca53d51845ed655b0bd1772514348b6c03a4a44051345f0183845
z38a4fbd04c9375d90f9ee974e851ba9a2c5549c898669d8281ffb6d093028f7658f6e9cf2d8db2
za163d3814d3c1d54f689449365d2d1282b9204b52e91f09d3bb5caa1fc3dc6327ee18864b7e54c
z1fe9599691cf4bac8e8b1ead1500361270ab6fb2f48f24bc5ada01ab041560e399042baf557a98
z69b3724fa997ee144a5cd529f118857cc74757fb459034f8c0df2c9262befbf69ec04d39e33e52
z22a9033fd48ac6b92c2591e1c37ad1bb50fe42e6c31b9a8d88a255f3c464150f74829f3b0302ee
z8480d33f6a36d355ff9596478f8193297d6632f19f846a8d21209c893d1fa1e3e5b7f46ebaa789
zeac7d4ed9947da67f194a0df6a3cc59646155bdca6473dc2e84f039fd3ad4ce8e44c590e358a6d
zbdb43a5333505906b57eaba061c8304f5d4c8215ea7dd60c27853d0de6bda78322ee4fb8060c1c
zcc9e7f1312a07ad9ce963b4e59c331c6930060aad9d2af2de69d5222f58f18f2d4e5dc5dabe7b0
z0bd03b5b0f6e500ddf6f98d61823fe0ea8652a8bff545e6dd8d609cd7a66f5395e962b5bf29401
z13e444c3c65e296ee30f3a30fc97a9b1bc6c688640eb5e81b60f8fe549a98d6fa22ff18ec863f1
z77d8b108d9bca534a643a03ae08dd780b1582217db9843226606e5142c816a93f0e74e5edc693d
zc1243a9da6d9469125d7d6aefcf31c293536968d527311a26fdb1c947c4d7b788efc426a74e3c7
ze37745c2585ceed692a5657775540fb69a87d7598931181042017c223c0bf1f4b46e756ab47a20
z22f3d31524a640deb6e2c176e5df9223b955a3fe0c0e8a945a09879f7f321706efacef06f019cf
z17192179b6b93dfeef9544180ce6500d647b43f9dbb002b85e42fd9e317d46347f0f79b40b2855
zfb6524ad2aad958b7a23b93222cd16c9e6d6cd730352a2d0aa6969b7b1a15f32bf24fa307237bb
zb0752e831ba1e576dfefc5ceb94126050b81ff509ac8c0a18083217669742bf9739af9c78ec829
z50f6f6b70907f88ee05bb3d1b7f85c311519902466bbffe757ff6225c3f3d9d1eb737baf890e08
za0531b6575ce5fdd1194e99f9fd4bde123dc0df3d4aaed6d7981c1542925fb8944cbdf4c139b54
ze0479f044372d6cfcda1d41f02b1794214be2ab24fa5213e6d42eac5dca16591627e19036056a5
z8369544c87ae8c11aa3583d95f2f03aad17e1677e65aefad7e8e351544315d5395e1dd52aab73f
za8f55560a3c786df38bf9c3d602913556609df6cdd4204754b5d682f6e87833ae6a5a72ce7652c
z6c7bc8b8a6fa682c7437eb97075b8409e9c6c2fa030434e9f4e280bb98d64be25d0631c1cca86d
zc1eaf67ed4810e27cc9fbd563b0fb17d4638cbf84dd1b9583735d9000b76cbf8b72d81bd30e944
ze389414d37934716a1324b48505e98c8e2a63b43f1ba90ac0ed96bfdb9a0bd1a5a2ff9c549811f
ze8ad6e3b31160bb5a6f1f54c0b831f7e0932286171de0d3e63b33a1da8d343265701834b1c622a
z7fd684f0f223f49987d91f014ebb2e916e3222d8f6ddadf1cc2b7aaad690ef5bbf4f48201ca2d0
z3fcdc29e622f492aefcee8536c6f8aa0a6b4e5a849936ba23d08336200e80675ffa6aaf20d2204
zcb436ab94b5dad02ec6b88a962a8e04f8a8b0598c585151482b0ecc0fb5a5968759e92b0bb2f4b
z6d3b63a1ee131b7e3a45ea997ad688a5dce02924159499b4702780c61891a1af6f254a61ffde91
z973d7aeb05c08bacc1e278e9217df2f30cfed7252dec1ffc1e7703260b325b70b6d1d40bea6f8a
z5cbc2784068f3cd3d72307dbeca8af5af5d6590e705668fbf6c5e0994754a84022c2b5fcc62bd7
zf5ab8827d62d1798d2239dd11bf104867899c7d2dddbb931bf5c8078eae1926a71fa1192294ca9
z66e0fa92b984a3a3c80e2acf57e560e662ee4d234c262688b6ae3256c6b4682e7b35c14b1bbe5a
zcbd9867f57f13c66b8010baf1536bd4cc0f610602d8b123e0821948e280a238afa4f9ae0b0b91b
z538dbef6afb561d047bf9c379c32e92133b9689c5a00e1a8d148d199abfa5bafd29d73572731c1
z5af033531a4db1ba2b392bde455d712d1cc7b536ba8e6dd5a8741df36e418157618c6ba7e0a0db
z3582d90457d84c19eedf0e70f0984c220dbd1ebbe2659e71943cba8d47b1e6dda9ce813e6db3bb
z5360e64cdad82a0d9ef5311ae9a64631e682eb94becbdb3376a2f7408feee0830d71d8d0442b6c
zf58eed8e8796a68d3c69980c30a958c528df01a9d5b244ebb5437963ae2d212ac9a8ed5b27291e
z71bd1c084fc93f9246ebf10bc4411d4c7608837515bc23966dcbabbde0feab2c0666e0d46895a7
z4e4dc0760a586df4a751fddf26f44bbe4ab73c905fcea74f0adc6c393aa5a2093fcf9b35f71c57
zb315fce88c56d7fa6b3b36dbcb3276a82ba431fe24c9a5507a740c5930dd7de90b7982cb428ff5
zc1306505c0eeb6a79fcbe42cc7aecfe6ac3d87feda0387c8dc6e80e6554dce1907f7148b465429
z2dc4b0c3453e42b203b688dc9ab11df3d9ea6dc2da87a4536e98bed1cf75ddd1536c5e811c717c
z11873dda0b212fcfc91044f6361d26f8ba6f5ab61e24a2022550951fa95dc34e964572b892ee1c
z42b9f96476f9feb936203951f70666a79268a7cf33dd71e88a1347473a191191496d1b248d1e84
za83185b035e7a6e33f4a166fbf9f913adf90af104601289b387156ec28e68eb3e5fb6605bb653c
zaf4524070bc9f14495ba98a9f7def055511154b7c67ff5b0162b84926e1f9b3410d17fc354c5e7
z783e9b83c4a078a652aae1a85bd93f7a26beda1d8988a735ecdb20fa5ba43038cac4d7658da982
z7ff156da9d79d8bf9d1d2200cd9c43fa898971a52a496404f597d8705c1a2acb1e10ecda4ede29
z285f2aa412a8c24d7ed0e5a1550a2d9f9e03fad345f552c65b482c9820dfb332af3a20aa7aecfd
zcaf83bbf2831bdc5186de3138aeda2a93358ef3bfcd5a05c5fee63d9682a392ab0d49516487480
z26f42b1f3772e42bed5caf37d66db35e7787405d5bb8b56f2a3cfad83b1f9677321df7a9b80e8e
za9cbd36490f722ce255548008884dc5d1dedd774e3888afbc81137ca87002cae7f3dd42a63410a
z7a4ce5d08371776c42dee975129a423e0934649652be17b14829d767c924897d342fb05d98c82a
z0da75d4cc9d4f8736fb4bb00d65ecdfe1936c70371395fa7c8aaa75279221ba3504a5f3b33869c
z8adab15b80884f7265377110cb8d0f1c7f7f020347e4cad0cf3e7a080ff37f26cb82b4105894d5
z4aff13ef75671a295c0085166894d1caf94814958e7e1c382812d753af4df32ee7ce65439084a3
zff8a41e240c0fab430a5d383d8d95e88373b452b38db2e6cb87037df3de36afbede7276ec2544a
z5cc2d788741dfdffee0cdaa049823a0ae78e18f2aefa2da202433ff3582542b2170fc6d9ea4254
z68cb4a849c319d8089e0aa4b1f8eff3e8a28061d50717dc3bdf511438fe999832291df861166fe
z1f4f86e12cd90b7cc4ef597c9b0540b9b3b221bcd99544282bdb386d90d32d1ad7f45cdc6c23bf
ze0a22fc401b27da52bd9ddcc2eb37d6258c1d3276647bd4336f90f6e2660f0c21ae7b61cc4794f
z4380ad86a9f543be07010975cafe2f41dd0ef44e09d41bf5d8a6c4f3473906994932c60b655a26
za8564f9f2309e7d0921095808f249a5b29ddb6738ee8f314e75f5704cb219fb9ed882f6229ec34
z436e6884519934eb63d54aa2df07c16de8e4920484a69f96b52767160d456f8b7af4c08fccfe09
za757c1e9a055ef706a2ef727b897a44890f95c741bf281b03fd07fa3532d09a34c640c924dbaff
zceb9b4924fce55de1319ff3e1ef82a4f207044fc6c465d8d301d7845d64d55e667e11edbcc2f6f
z3e045c1978c11d86fb0c0c665cec469b001ea9e37cc3b677ad6204efe7b629e0dd8da517dd509a
z9144b037e5ad4b8de04f9c6fa065f7e6e610ea878ffd674111af4deb0fc439921f54fe74c8f53f
z2ca261d71f4a55daa740431142ff6f0b0508da2d259bfafd8c0f288d85ed2685c664f9841c4b79
zdd5371499d35f3103e6316c970c385cd3bb7136b28ef0d6688e35a75391d4a7a6b2289ad622172
z99b6330c4287aae19709561e1755a74eb008457c4f1aaaf18869814289778dca2aa588cb405ee8
za8c8d494df2f8b01b21457191e9cab5a9c7c2c41d6afcbb768a3ccbc9854f080a385fedde56d59
z0bed21e9c08dd9ff72b5e5d9fcf9021403e6696dcf68fdecb6dedba7eae0aee70d37c768e571d4
zcff5b1c6d9d65818e2858e851d8af5a3896b6797b76541ac921cd4040b2741a3b5366175d47af5
zaedc078ac3ebfc52ce0cba7a1f89bda2e83d63232a6cebbbb936834371482d063d8badb8415e59
z68c9bc3658eb37bd046e1aa10ad7aa8551f5c175f370cacc1daab8b0e13c98f311b763d0786215
z7cfdd70f50a6b246371e7d1d9238949c065fb112e9b367490c753b4f0cafc290305a781260d91c
z23dc35bc5be187273c42ef5a6e8aea71eb0ad9ec2791f3e05a624575fd4b90b0de870b55b45cca
z199f574fa4d9b39fe50d1eaa6ef22ef17fd89497bb5a3f871ee592d2cfbfdcf5fd7bf3ee0f3fc2
z06815ad1ab021c19937e165b1180b862d814114e7bd4bb42f819f6cd117e35b3a3a41a396f5cce
z1909963801c396a3dd49602e61084adb615d7c96a5f80ca4d2f1e09d392dd47b5f241ba5619be3
z554f009121100a37f8649540dcbe69dc8d4952a551589f9a5d3b3efca825927b0b6c65cf76759d
z08664d2c1be39d4f459bb5e7d9a99e03593a96215c0b1d61988d4ae45680613f0cdb1fc634c492
za9cb0b166663d512c4c29bade161ae3dae426c81fbb59b85edcfa2f634d6fcd154f267b6dbbc53
zddfafc69dc4a4f346d82867a57b2745c6d6f3c1b6fa4d94d1be2c228c8d592e7bae058fe734c64
zc529b852068978edeae4d6c9d0ee8839f2300b1c12b30d7c27591e86171caa176005e40defb6ac
z1b499456f40c32098209fa22f389ca29903ffddf9358f8daab4bd6c50056511ce44972f5c8b696
z84141e0a4413525b3264a7871ef354431399db088f3da5383c62cd65ee87abcd9ad7c5702d4e5a
zc07e79272c45461964713622cfe89cd7aff247bdbe654f960e61debc7124d246102ee559726543
z2f88c36193efe1ce418d9ee9212580a90149e85b26489d8eba79190ae4eb03d922422e6e89779e
ze4d773084e4fa4f5817fcbb5836a22da84e3e3d2c68fce2123c6b7d9bf20b1293e683a50673672
z53d718b65ac151a3f8eabe3b68e53ac386597f10cf40a52aa3c88dff1a46661dce076726c2e58d
z34fcf1ee51a235cb73782055f0e0ed8cc7d5cb22104817040f07f7cbffe13a805fef079422c974
z126688566eee28814a35d38d6aad9782139b9d8a7ecbeec605666c0045301a424866ed27c5188f
z2f9d6a6e9283bdaf56c87de8819ebe3a954aa95f514f4bc3b3d3c20c1e1aa00add28e4f89ce15e
zaf73adb293090e2558fdadfe245330805f5803d964493aeb38b85aa0fddb936c039c473290b14a
za53b72f87570745e1dc067f11da40032351d499696ab8176b9f2478c1621261f30afe0c28724f0
z2427a63f69035e2c80de1e32e4947fc00770f5be89f9aa8d03b8dc1e59f15de450e7d3c03a8858
zdead9663fe678e0e0258dbbc0e6192c6da218c8bd9588771fc7d94d1572a43fb87e4b2112bd8e3
z1c8da1c5967d85920844617303f06c694ba85b5a8a34aa1c7e955c6edfe93ed77d6f7c8d780843
za8f34b6ed54e2d4d8ff0968d89ff23c3eb9f088bcab000c9e15381bdb3e351ca9bb359aac53d9b
zbfce00972adbed9990c89b75fb064059feead4cf7bb07761636985456e9175ca7e8d56e0d2e946
zf0dadf8e6d7e2ebb365e7aed8932ff9415b3aefe510c4ed10682ba99f92656b334c7c615bf6d1f
z48eed3476116a59bddf83459193ca047c1db7fd553a78542daa6c94d97acd3016871d3e4b965ef
zd0dc67dc73f6239a34a53be8927cb944533611b6cb9e32c970f3a08e37ee20f7ee0e300777d776
z531dedf66a4b6b16a9abf4761cc7071f386b75dc51feb0811a54d96f22a0108aaa7cd739819f64
z245beb0a906d216f18c8b0a5d95fa0fd5406280c029f86b49898b58fe21f86ca72a07ff9f1911b
z5e70680e319a489b65ddfdf42ab9a845ec0293ba40feb824a4b2aef7f8ce061502e0a4666a3479
z9460c826fb2f3ba203ecbf7215f8f2a609b9c6ec4d8d5ee3062b47fbce1b7b4050ee9183c813fb
z6d24b86b70e4a39b164e40312f087b3e787a871094ddcadef71d2e4154dc1f22e0a2ccd010655e
za996652c571d70ffeb895c0212d9aeff6bc10b6b1ebaa0b44efbb5872bbd66c87bb3f83761734e
zbaa5d94174eeb7d7b8b0a46b882e7ad8a1900b91e8c09f7e16225228a20d16a51ee9b45c04624f
zcade4c3082d73ab674b723edab9befd0bf16e2c7a2834f1005d419862652f90b14a948f8e07b34
z2e2eb2e19863cab86867c3031fea5ab9c728126b12b6595f391246016741e70e2febb5d0a135e1
zf2bde58014adbc15efb090d1a5c8bed4067225fca1eebaf9aa2e8c6d62886d2815c7ce10a86220
zbfc4d34ed57961191aea00579f544e78ee2e36a24808036370257cad4281fd0f21bb522118fce9
z00781b053947e8aa53613c5d8a9f4da5346b31796caf99abe7fd43b2e19ef123b5c67adbce6ada
z7a84c098a6e9f82ba62d95e317cb3e0ba2f96b35854bff5d9bbdeb7aa7e9938aba45d7ec874d16
zabe6bb87a0ed51c9bd92246bb3872dbf86560feba6b6b1f983e99c836b9c4cd30871603b114f70
zfafdf0feacde0c48412dd10f4def7d062c474439c8bca0142493fa1122dbdaab38e718915dd4fc
z69f3b0ecd31afade00e0947694a1367c801ecf144eaf27f53999728cac03c55d3f13e199476cc8
z8679246d6ead419a800f26c9890a5706830490f86059cc616e6a93efeca4fc3404aae816801217
z39754110f8d4ecbc1c6014d8a4de043fd91234d7914e211b91c11147f75ae6a66b908aa4e5f7a2
z2b3defc2f675292e48bffbdf723beb450ee9f7cc413d7f84befd5349ad5523609b5b52625a5ebc
z3ccd9ca94869ec05ea7beb90bf108a75e2d3de649d1593888e49103c66876735303e0e9c1c3894
z27d334e622992c9a7313dbddb4d3f3a389d6e4538adf2527739151e19fa16b8e1ee7c62d122f25
zf3336339077c912b04b6405231c7acfe5156b017a5ccac91a99935480a38a19c468439b7ec41ea
zf3975fc0207df609ad5652edd3fe8600c31c5e79adbe522300768b3716170269d814682d127abf
zaea2b972041df344600458b93d243bf216e09098ac9f618e0f047e5c888763e8195c41080f8a10
z640d769fc62532001244af2c490762b823cfd344cf07fcc44854f214f1b072eb0bfab38639d842
z2a54174d1dabcd7495b448214b3bda211498fe2234ea6f6ae1e446de9992bc1647188df258475f
zf11b8f6f42b9b6d6fa33d354fde5ac033026e925bc4016f0c18dcb71c453de0913e501dafa67b5
zc7c968557d5854fed1f1870a422e9e633df04c9454e197f59625b8358e375642847bae70c83ffc
z573537005a901c7bc9e639cbf5effc7a20ca1a4b49cd51f07bbbcac153276fd52715ad28e2e61c
z3144382afce2d99339a1a24f3825889fcb669f61ad903c6e4b774506e3fa665f4b901355890a26
z9da80778b434957e7828f09772137d676e84fd812384382dfa3a11abb80e9bd22b44845d5fdae5
zfd95c418ee1f8f78f420e2eb301c6a4a6c7fb865ddf180b7eac428509896166fcb16d63c1fb2f6
z77c6c8b1781738083b794cd5caf7ec61f16225034c86fdbedeb239e23920f5cb63d9f925349e73
z8720f010e893163d586a8e5be19dc1d81687e8110505292bd3ddbe9502636bf67603f5c0e379f6
zef8008503641cbcd3ab6267681406e7194f7ba92cb4f38009c270d43643e3512a29f6604e151d9
ze2088adcc88ae846e14cc3cc9d6d558eed9b920123644493668f198e73fd33905c2af2c0706c11
zeac178c6631bfe14d660c5ecc6f17e23393bdff6c8cec6c2d06d98fa6edeee6593aa7be1fbe316
z27729da1b1c030fa08810868ff9e3375a827ec26086ff21b4132b042b040e708ab2402b6442acf
z0f03264724bc6b84eb7b536db50e726451acf8fb64c2a85c586d06d0f547a405462c8b37e0b6f9
z5b9cbebe957f639dab5d835ca65ede9a41e60e87a6dae7ef2bf18b880326afcd7756ed02f04fef
z59a8c65b210b1e135d2ac343690d87ab5f6411bcde1eef4dbc1139849cfee49085d8af5c9dd28f
z40364954e8b75f61017709e90bfdc9013806a4d9e943b2f1756f0e9261fcf3e391121f12d3dc0d
z033a706ed786fb3e933bacb41ead2aa14a5e9e7e111759d774762ca53545cea4a632fc58c0febd
z5cbb6b0f3e58965d2c814f5304db6ff59ebef1835f292486dd0b05733b9265b4519e31e4decac3
zd720ab22cbd6449c63ad6217960bc691029f20f6911bb8f21b0800fab08aa475611215bd33e1d1
z8cc3d1b92eb6b7a5a41e33dc517f6f3ca13300667f8b6e8d73084aa7e69ccb812b50db3120f72e
za13879d18b182b8d6eebcef626de28466f3180dea526c8dc1222f4c3bbde98b8a6c28d1f19e9d1
zef359dd5d2f67c507dc5e82f01ddad71e9c8510c70d6518c088be411f103f08bc73c5af6330da0
z42261814feb76fd221eb54880767e030553ffaf29d2b9a8a17b32673198dd704a55e6173c0ac7d
z4b48f401940a0cb46cfa2b1f476abc1cebbcd4a56e4749c1615d53d67f1421ee5f88e32a481530
z46f0ed64a8da4c0df932e86114123bedb1ea1064a83a70ec7dbeaf754ec0fd256db09a4e4b54b7
z87d169a4df0b4b583863de1cdc6f665ce370c9c014ce04a25d5e526f41665aea8ae20bdfc3ac98
zfcc4a0a254834b3e17fd7adbf5076f490131ccd7d5ecbc2f14199732208939be6a37b02fc8e12a
z1a63e009baf4c1213bd20d31f58b417fbd0ae0eef67efc5014053dd4a2e07ba6f06effcef7c833
zcb4c3a0e4e984b4a3f876ffa5eb3e8d57b2d122511c60d798dc38d8270558fc5dd19e3f8dc36cf
zda7cb35408a06b1399b43355f994e4bcb752c11d74dbb985bf7852bfe0093edfc139e0b8fb955f
za66e5d1cf314cc28705bc50045a2cda444af210d0577a8925cbde8e515d00f80f1f95296c6ff32
z1dd96a2bafa4b64c1bf4722655e2e1cb62a2161b033825dc459b1a0e7f0789493d519717ac4f3c
z30222e83cc77ff6f2f71f08f8ae5657c788cbcec252d80bb93892da9d44eec63822be6d883535a
z3a1d4ad453b89cfcff5fbbbab2535aa04a1d6f97431ca2c578813a709488c29a8b46e678b77c8e
z3a9c58524dba28ac492a57cead20a3b3d64a3f35390232d4464114d7abf5d294995ea24ea76323
zba67292cd44a872bc81d0823618a074bbaeb3a683d4730861aae695039738593e0619335dfe9a8
z26669f8cc39429bc451127c00ea4e38ead310923c38d9ee84ea14468ac14ef187612356799ea9c
z7c1b4dc0f3415beacfc450ace234c7490372a9a0c50845722b93839756c7b3e368b09bb35cc0ae
zc30c5749a544f8b12002031cd44d1d6119ae0e3326ecbaeb307e9da745b1a7da5689003a6bf54d
zd86465f7e98edd565e28451c1f21ffb0264dcae6e3dfbec2b424d058e4ab9a46b6ed3019850d7a
z7825259be9186918afa5601914f53076cb6db518847de6f9ec79e89ea03f5a68742fba3d4cf554
zf40088c7aafddde4e47d5f6ffa34ebf201962132dfa08abe1fc13d5bec7e690a978c3655041834
z826c45ea131d1421b036b86b8e4060526a2f205a06caddb658a2dc84f4c77cdbef5e1ea2afab84
z13451c9dcb54de345d157c1a90161ecd56207582024971f8edcd6b92e3925d260ed3c08bbf6032
zee8ecbde6aa7898d4d96524d97a66bf09f14fff2d03ce14c9f2fc52019009c9a67f936a6ac0d41
z9bc1a6a106f41cc40b50038d3c58a51277fba871803b16b2372d54a95ed1d56c8311606ff46562
z7145a95a405f55fe0be072a0c509f81ae2369b52d89c9a0d5ce85d0d455487dd787a0e1fc55c24
zdf5ec86e90d0d3177ec615fa553835fea6b5c033da33bedb539d35009f463d473142ec59ef1804
zf294c810d79998f8fe97807e0f3b295ffe5318cdf14af6ac824022919b4bbcf007485a2c4b28e6
z2ae415828c01e9a6987d3d0c41aa70a9a8dc72180e5cd8d6c7f6ca7920da82df9c5045e073988d
zf808cdfdfbee8721da756de0bbefe4074483a6030903b85bb2ac562e7525eb69e1cf4542e094a3
z2bee9375319f71d2004d632f838206464df52e7bd20ed6bf7b2415cc97b903909f11d496a9fb07
zd1d2c294f6638412432c2cf8f99e088427bf8f6cfa09c16bcadc695d5ef82b36f5ff62162bc360
z27fc252e52874b36382077631273538019e2ab8f7e46a17ab13e29a0aa218b805c37f315c4e394
za07add371c1831571d22671d2583066050fe31a77d820f1dad2372cbd21d8a9cfefae26f789bbd
z766de6bd8a3a43af06cc0dcb3f8b3e9949de97b1cbab8b11d9bcc18d80bed3ebb49c6ab8cc08a0
z3402b0aee8d2c62f976a5694126c737d65d11e0606c216f8a959cabab6a14eb7ccb819c7119ce1
z227b5abfd70a8a987fe841b0a5b672e3489910fa14a6ddcf7f1d801ee1ef2a1b8832b6b6ebded8
z0a8ceb523e35ce8f62963c904e1ad5204c83a8f4255accde795e40a8889a00dfd17ce925b50290
zafef50325da76343fe55fd974f6f0b1347c568cbde4b7f7d8e8d12de23cabe5a22a15915341e45
zb83f912ad1cff3f601756816750b27ee656d265ca109ddd879672a4cff2b7652a830ecff93722a
ze888606ecd463835a06e3a48d7dfa10b46984eed5d496dd6dfd645e0278e590471f343af3a3743
z6b9c893d71d12e09b28fddbfa3cb5435e4a975b7e1d912ca40b50a473cec24b748bd4bea6e7fcc
z62e95a1f847f11b3be17bf033ab3e5f5d8e924030ffc702d0c525518cd6d7b57c583855927410b
z708b73a46bbfd47ebf9c4a7b8c3c62c211c075938349a03f655e5221d373998cfb2131f089013c
z523cfb80e5fd2ac1fd4fe7fa6eb0a68b47de9efec073eabaada1ef8800c3dff4e2e29ecc1c59bc
zd52b5470eef5768870180728f0330e14828083db2747b10b3d8291f3edf77d3f8b0ab3b62170d8
ze4ed5b58b55c13985b31e7c5c24eac372f49baa665ee3f984852ea4da4b19326edfdd26ec68485
z32b0d971b61eee3b5864912b81a14cca33bbf6e1c982d70087108af53f7bec448b6e0ff465888c
z1e95498f08455173450723621dec2b0c84322a7a281e94160ce6258ae990426d20b28e2c6212e8
z2f5a5b02bec9a71806c0780f1aab5ddf2361f10ea008fd3f4a22e3b4affa51f874bb9b39a4fc98
z37982c540c251f02790e5525ad2fc5a2c4b9de2abfbffa5527f6387e424de35f71c583c02139ec
zadc99a3cb74411b899d197384ae99689f85f38c7d6c36e738c86bd271957c51a01b584f72c9568
ze10052985a565428ac399e2a4555bdfdfeb86eea38b32fe06546ba6469852a92285e109559fa80
zff008ac64dec539e88fab251396a1cbccc93fe523fd15e4d262315534486f9b8d21ef0e91e4ca7
zc33ba5afcb5e93373b6e678b6dacdd7dc0790d65b393a186f34469b0b1223cb37bc19ab785e9be
z5eb2132aae5539a9c7e6e069757b10c913cffb14934ce6a043cee733d238e02e0dba19b106366d
z30d238afe639a692d94c0abd65d2636f0015b5ec14deab4dcc2cd450e6e8d957e92baae384e5e0
zee013ab0d64619ed98a4626a64993081b65ccf849d6a4022baea680f4d9817f79ba91f24bfb5e5
z3e52bb8ccb2b44a5955e99dee19c98b00902abdc297b20cf79da2a6adfddb847bc1304bb699186
z196f5af24e165c39aafd9a663a3477e0a7cf9f5cbc1bd02c692f6d2bfbe97e83a7da98d94bcf62
z62fd9585d12767f5fed5d368394dcd86cb6f95c00852c304f9f4471af0f75404b38c85e81dd997
z65872eb7a588cf99ee4645462f8a024c0a2b754252f7eb318e90bc05d8864168e619875ab329bb
z2f48146657aa91d56bed014a8d5292542c7f9e9b551848f4e122ac5d2a1186b40d2dd8aaea4d57
z47e446e5c88d3715ace20e6720305bd8cba01c64a4d91f07ed00cf462b47eda1cdad4d2882acd0
zcc66d594714cb07821eb787095d6b296d43c6c84b6d27466d7e37cac38400260628173d40a79bb
z9d92ab95e2fffbf3b3e31206efe82b959ddc4538a61ecaf2d9c16a58bf5adb20fd593b5f2ce05b
z51125b0a0d2ddf6a37098d9db57e9ffd2f20a3fcdde9c2f9639d6c781901732cfa02f4602f08c5
zdaf284f089baabc5683543d988ef3ca853e67c6d037c99df7bc83fd8057e26b2d5e6213bf33aa5
z2a17d1ec3ba9501da2b067fdbb44ac10b2f869431e009f3723e02705df583de7e5a6d085df360d
z2c3cd082bbcd1d0ee64c7a6ebc7aafdeb0e247981be9e06c1fa0f9abf14c508abb83b7bbf2b04f
z9bbcf5b82b99a8935813ca2ac65f67231662d1a98917712d18f504d5ffeda05c5ae09438d4fd9d
z840288ec70b625056ea68a42fe19f9719b4a2cd8f427a229f9693b85a4eb037e4fdc17c722280e
z179036012029997b8f1cad8f39f7436af5d32e3faeca4343bcfb4a72a250afa560873d5933be62
zcf7b9b1b387122c441faac0405e5717e83dfd8c17a2430e200f2ad4a7f5f54001517332be1d0f3
zc3293ecb12cd2e1da6adb9ae72e5d56b5a33a82ed2739fb0897ca131616293e1d4941c37ee561a
z0e566b93f7053b737a966cf78699624b723d2d872469786d4b8297079ab255bd97febbdd210d56
zb6b0f566b1a98c63691c55682a9e8192126a8460c548cf41bb63bd9fa1782ec25ad1694fdefda6
z0288e7e413394869de44a5efd77578e58b5a2e1d268f7af6e4c7e90ea13fdfd3d0c029b6066404
z7844f692b4e0191df0f159af363014a671b2693072d752e18fe2fec451b7173175a9cd9cc029f4
z4b83c10627304c30665054645d2c61ae40cff5f7fb76e0a0dd91aa329366df7af103c72eb1635f
zb6b6097c2079495a25c03b4fbc29dfc834553d51557284ed0cd68493e7ad47accfa00008e2ba63
z5d0e44bfd2f083fbc0cca7c406236fffb4c53a495ea69008c67499d1e9262ec3c83f20d906bd09
z7cee18004889de06a52629c95113f1a3ab2b4577f6f259cb0c609fcccc642c5e0e64da27154cbe
zefa965dea497862ff99c9455c92c3d6355ea75e36cb4b0d89e0ad317aeb134cd3afa7c332fbf77
z559e676b4eec2df7e22c2aab6a3e6df03670add801114480766ce1315ab23ad9ed1f2298c04a77
zd0a68a4f49d0fa7d902c53b172879f5577605cec3b9451ca4ca1445c0f72463150283988b870a8
zb793d65a55719fa1b4f259ac70a3446b4f2c65f341e7383fe27ef6d0e8e045ef3a482e25390dfd
z812ce0455da843c693855485bca2e47e9983c178f3ae457c5a5eef06bdcf85329c29822442a1ae
z2c02c103869f4fdeff66dfd7267b65137021dc6776b7451b9360c5e8608fe78a7c9b72eef2ee31
z6afab815197499c16c338963bb11d866274a1f1b7b6f8cba268cc125ba396c8887411b06912e19
zcdd8468f7bc70b8e34a85f22e760d20da4f477b7aebe26a1f710fd46a3a114487f39058f4f0ac7
zcc3055294317fbf53881baf82a940d94c59e70a54ae331142ba9b34f5bfb75654eae42c72d9797
zdc053d3c8b4ce0081e00eff993610b1217206fd580df3ff18e32058fcb282dba74dd151e06ee6e
zb8da807de00db021d8e03ccd7f94698f7fed79f7fe1ed65bd928d56e3fa58071ade75117b42eca
z982bbc3e074228b6ce9e2eb28d85898ae7dbf112819c3a9acd17b50d01d94f7feabf9f376614bb
z2fb9e5a72c12e1c28bd2bd1d1692e1a96751e0ff4af151718a29f6af821c1891cb32721e5d0e4c
z119da68dee42991cf61b9bda2cd7dd663ea9e68b9d8baafe7e3f469ae49506de2699168bba22db
z46710e4335289ee19f5dca282122b3a7bc1d9942ac51aa1b7b6c7e17110db45e9581842679c061
za999535284b0332db831a5ffede7c84667544a6294cf8a9dc771843c2c5fe6b69073fdef59dfe7
ze4cad7720f1206e2747afd960661cf2eae0d65c6f7d9d0e7f280f1dd0f4b1f443791e9e543bf95
z54fd237dd05d42a704eee0e01c1cac0955c65069b385e840bf2314c38c577a31c7109fef0f97c6
zd721c095fbbd553dfce45adeecce81f1663adc0174a567d43b5d264e8d4f1bbaed6e22c07df753
z2fc8d62a8c816677df7afa1087c0d2b0de7111f69c01558a5b21e87c89ecb63ef50088546b642b
z55ad11086ba243d26ecea9cfcb8834b40eadea1a16901752e16c95a9828d0060bbdbb4df517069
zffcb6e16b08c5ee0d467f723b582f7febddc10ad1acd3cb2ffbdc79a520e602c5a1ab02701305c
z22ef701fa8579802d84d4515342b3e195bbf0f0043accc92224bd3b58361dc922a128e5dc7e4f5
z7362df8cb9d2680fe0084140dadaf9990888801ede24e896ad6cedfa3841d8cd9de0ce175badc7
z49a03d090290cc21bfec4c4b67129a120f097c3df3c2b68cb2437eba1b3d1e1a7e0d26630695cb
z7406dcfcc5cad5d596bb5802e80bd28ab68f51abd7deaaedb1dab274a46c7ace9f05f45a3de12d
z701a0f25a5d65a055f5a63bd71cf4d222ec220120dccfd6e878c553275e9e3e756d8844c26c99b
za248d049e15ac77a7ae9c43952554091fe9091122e9e98a07692a5c8787326340996ad38bba900
z629a436021ae27e4ae72e9e20cd5a927b0d952d9c834151bdcf5416c35689696e8e52634f70341
zdcefc05b8a953c6a91a9235f33bd69c00d67d25e75fe30c33ce58ed3248687c1b70ec86aedefec
zad2185ad1dbe89ff6ff4f636913177c99b3488794a4e40da8b9309d80925f35b5dac2deaac6ea8
z693195f7ec317ff394c31c83ac25fcb78f5839605218ac15ff4372b2b85fc6323498732ac3a0e1
z25610db892190284ecbf9931b8f29d203cbeb7e5ddd58dd5a4d4338b7e7f868a83ccd25921f75e
z8f1e034e51f8426794378b3940792fc49dee12347be156571bb6b7f5dcf87e20cd565686c4773c
z177517f2538152b5390cdb158f641cd1838784fb04d4478c430245c78947852f32228d12baedfe
zb139ebdeec5fc15ccd3cee8ef98f4bddf63cb541171086b92fce3561cd919c3b4b8025c428cf62
z56c4ad409e66efbdae7ae89aeea0dd008e0ba357065a2d3f3ac7d3114d590f076e4d539ea5b8b8
za234bb5231b9bf6d2661fa28c2ee21a9ed8f54ab670b5492dcfe7e6c824c5456b7b768f68f54e7
zd0e66a8d0619784f9f8b9b3266d665a7c33f2ba7430406782d4035663f33e227a6f8abb93f253d
zaa486e58b53f73ef9f658c1a4bdaf9444e88d56681eca62ddb14679a15cfd0594643908f50704f
zb79bf820c6cf0559205e0e4f897128fc7fa0ded2313a651d9d40b95abf3ccd27cb58cbf84e8184
z1da83f726d9819b53f0bddfd98e8c98ef05edb6196e686122f1dc0d210f719482e7f0bd90e1e65
zdb897782f0c3ee39b85193ea84c2e2f6cf154ca13e0abaf8ccabe23fe4de8dc9f700a0d0beb229
zf5cf1c65b0545fdabe5211d9135b10d3ace2748905aa65eb38c50bf73875ee4c4f034459ad7cf1
ze38af10dccb14b87ce63fff383a99b21dd922ec915618d8b857ece36eaa942ab1345cc9b7964eb
zf0aced517bec4e0b93e45891eecc9ad6a33fdead269e28a0cad19fac38f919fb21a2dbc982f9e5
z1911e430338f51f36d603f10eeee9794c35a4d429a4a344e5c6e6774236984549b9ecef36aaa79
zbc1cb6b6949768b3df312f4399344e3a5f72a135b7667c6c199ca0250b361096829d74bf762f75
zfe9a6fb7eed452117971b6c1e7fab09b4fe30b8457d8908252a99e3b85930191099cf83f6b6185
z5073232506665c1b1b0457c2add649635ff9ed0bf2a1f476419b588f0433e2bdcb5e0ef5daa982
z1652f507dc6719d6ca9ded2b59664cfba1e23f82b7fef2d8a77954b3783aeacfcb7911fbc6a62e
z99dc16809630351116c7eca49f923180869e5f627e36872311b8fe6ce4deb9c1a038665a5a7b39
z42e70b82597581be78703fb866281ad706fdb82bedd6e2c60a6ff1b258355a1efb84ed408197df
z9439a06600369fd24fa0d2815a48dabe928c6483a3d400144951fbd8346086e44b3fd5845e39b7
za09d375ff31ad6ca6c77770f62a555ecdbc9a751294f53c1346d33db32471ca162ac825d82b17f
z37dae314bf185422882eb855c86e1d57539d073b23c381b1b76f76ae1d0912bbe5a6db0b55ec20
zfe1b95dca06763c3f15c806cf7af7c7a1ff81d15f641ca25ba605f37942b976a9c8d9975e69307
z81f3b4c75f1e72a7f44fac7ac77e0962c5246b7435d9ee5c14b3017da63a1d9b5607e481919566
z8d186f00a305f87962da1e8b62ff6681458c09f60427dbbd8cbaf36601a85c2f09255203c4d94a
zbb76e36dbaf85eb445bf64159bd048514d97e77ffa1677df2e28490a5c891b317f7330ab8bc016
z479c765e1dc989d027e2e8f435a6bbf1623c7b6a1d0974a152a6d1aa85f4c2075328c08af4e61a
z33bf8d01be4bd930d343cb16737cf532d0ca82be813e83c7275af2f2d75b6ad71ef151cc7115bd
z09bb493a5d2a2fa4c9f7c5d4ab1ca39b7c65ca4e6873cecc6a278b0c25f894c71b3922ae84e3fd
za00c5a32b316520ebf055005ff73f1040d8e49e5391c46b918dca23e8e0125555b2f47f8807a91
z89263c49f96c1e3511ddb2251248bc3643a75845d491c034b092143ac60260c34fdc36e0f1fa70
z297e46dc3e0a284cb38852c56dd1031c9e45078b35812ed7fea236783cddacc31421fb9bec74dc
za61249a71422ec0cfcc1218c40bf325d59f340f6aff813f473b932f1ce7dd5cc2b456ba3e0e562
zbf5dc0485cef35a87c986af5582feeab8c0c7be338c831574cc2c0dc86a7bd217a0c65bee21391
z507432ef7718fd9511f0fe0687d7d71a9e9aa0daeab78517781aefee3c3f5822236251cd9ce287
z696177351f247f4340fe3ba75635296b7e8dde351b1d267f8a29dc65a94124199f1aa4aafee463
z7de211b53aa2558b8a20fbf7d9ecc32562b388f12e2f0940e0b2656f2f7823871b19df4d18dbbb
zde342598dbdbf08cf828706886ed7f1f35e8b4de3bc300f683da378ea8759103ec56b6b9af37ca
z4dc937beb3324723072a04c455fc6ca4582666f8017dda839a804200ea1d169fbce5e087e01634
z7b47852d38654ce9e7dec200e4049aa17cd4cd249be834cdc5a186b7cc2dbdeff963541f1ffa47
za5a5f0fe4e7cb4fc204c57cf1b8268a2421c76e3cc050aed34de6c5d840a1e8273c8f647cf055f
z4081fef9422ac31e3bd7308beb425551c90691d9269876872da7d1d4cacfbd1c8fabbf901a09ab
z1b949d424768b1e6ba31b2e7c24f793d036c6b9ce2920f9c96e522953603af5eec7a6f2e8a7e29
zb935ae60dd64ff4c6098047de9b5dfbcb9aa54ad5f9b6f797b38b02af181c6a26391b386e4aa5c
zfe3bccfb688b1a76dc9613bc0aab036d76afa996063544331078f46bbfb17ac24312e3615be0ce
zdd9c6407485b96be7600199b5bb0691f39c03231492722014209a9e5acd46c667a6423d1f16a54
zcbd76c25ff0dbc9fd3aa638ee039235f3507d1efd3a1e8dc180a9375bd39c0d61c13e0b9a033c7
z6c42ed37584e0d1f52bf1a86730b12f6cc0b5882959aa235188de40897b9458e6d8d0710a02601
z13ea1bdd06abef24db23f5dc3fbf9aaeee8c88f50774146b45f73c9c043f35a0d84c454723b105
zc95ce8da6f7f7731fabe877e940f2fff6dd4608e44e0ef8c295ec6fc0354ff984baf966315fabd
z92f5bc0357ecade0b3ba3afad70d3f08a13fba1da856116685e850c20b44879f0beef1a701cc21
zf75321b8ad28817fcede56600695e54cbea4ce936aaa2df8a8d344dc83d35122a7372fa976fb71
zac80a2194945b48417cbe6bcc06dc622147c23d75391973aaa2e39361f39d41ee49c995217b99f
z5da3c8ef5ba6dd2d7f5fad4e1a0a1326323885fe44e048252d56899652314cfd7a965e7106dd97
z012c515e20e6fb13c1e2521388836352cce4f5868336fb34c5318d4cf06ac9f5eccd015672e5d6
z693596520967564ea6c5d6c5aa77b5222f6dad03910a8cb9a8e019ba2f69a6fab077ed1b4e8ea9
zf1b504f783a5e257ad06ff4a3c689c6a3d741eb4b71f6bd9ec5e709e670cc6d42a2b78e67e00ac
zc88de514bd6bd621d09b6fe78822d9ddfb62ded5ff1d03fa6417b34351268e1a8a29ab059bf65f
z28d7bf656891ac3b5a7602d929fc420676e4065e28f0c23d59ee307ac1a3b8a0a2c2ca52a3f7a9
z862f978f708a0d7d9c76f7dd79305738e80d67532bfc5957e81455350f09e4b3f2ec5512c5c901
z5f3932f7358690fca4cfb3f844a7886d6f03dbd1e334d51ba184a03f5b3c5eed4ffb6a517031a3
z87068abba8dfea56236e7e38f5c415cc49c8bfb6d025776beed6a9c1fc37149eefc3d343f1b6f4
z54a2066265b24ed88220f53d2db914a1e475053c4bf9b3b2363e40d2663ed209642c21fcb03392
zec8fd01a02d6198c17d719e6e5f3ef6f69da7e6a746161cd6b60d6feaf17593a796ddf6b598ac3
z5e808fc42a5c67e675735091c386d2a1420c521d985cccc229903fd20816391d5a0190263e4515
za2edc792651ccdb13a9abd2e510f2a7ff0dd243104fca17b4a5315f60fd5da3606897562f0a65c
zc19121b95b7a85080500cf50efc8c7b9dc52e4d4eacfced0a1c0347532550f4f2ae848a71e45ad
z64dcaf280042c0543bffcb81f11445d79576d0046cb5acd8dba201650114c3814f4ce5d155b882
z48d586532c2b2647b872f0aff2df03617cfce43592f3ae0796dbdd174f7cf10f3a0b224d3f3705
ze48efdace27ec27a910e80dadaa34d74c9afbd93d95486597246cbb12a48bafdb755206cbf88bc
z9cdecfa9e79950666acf31ded6aca89c33a63a6ef4d7ecb36755965714ff2be477109939331ca9
zbc8e3d03d65ec9ddb29418bd48e890677a2ec7f435c0721555e3e8844f1c9bd2154142b0a08dee
z531f764079d76f0b617267e4746ce1182a63573552c565696d3380dc5c65ae537d3da2ad24aec9
z7ef02d9c6df9ecf83ef51c8c4a584f5e2ef717eccbe46d528c72f80695a215d8c9aa811002fdc5
z4dc901e4b44913a50f803f87dd52d402723810a6f4dea35ef73b2f1bc4761cd6f387493c303d18
z916c91392edf2fb011e4373b136ec942c1724e39c0390d6f5460a2d2ad3030a666749430e9d827
z1bbc15ad229b415778d9e5448fc07bcf7b1573c4c2c22254dc833ccc9f9c541207b151da25c9b9
z691a849ce8c1634a152d7ea0885359100f33ded73a1261a06b5566985c4a2554917dbdfe69a8a1
zd3a402f89465c2062dee22c72990536d74327ba7cf8c6884ef121600ee0e824dafc814651fa498
z6c41131525ef376eb69945760ffa021a5a6cd2c04d490e11f501f8d7d6291674e78b59001e5c8e
z011adf36c5d1f5faf4092d82186e463ad51599210ab50191f9d3fbde15676d4551d6c8adf141b5
z43caddc2edb6c88da68de2ac5f3142816455d6c15cfd3e0b3096d4bd33a0ed80dd8cab80181389
z822cda3b095a958f8fef138480d64432035ecc13b460da9d071197ffa33bf2aa9ddabf3417b509
za2cdbc119152fd74d0083734ca97da4f9431bd6c56cbe22debc5f5a5dffe08da9f70769af1fcc1
z74c71a5a6d37346bb147571c7d7df522f74b1101ecb73f1f9ffbac7ad72d11b979876d18fd76b0
za7af0f303e9828aa0a4e8bf4e4a573178bcdc1f0993b7244eebedc64cdcc713b0068457ee97bcf
z6945bbb81ab5fb90e88ad3d8f671eff05191b16ccc06c14a2047f077958bddb0272cc4d89fab15
z5432bf240c91060733b29ae26fbd958f0292710a5c97b8f6a0fbf4a0e2246ac14a061bd6ef1875
z88aa78ac54fd2ae2d80c3f238cd7eece2f0ab93eb990cc55004c5320b9044a9817b3c1a4f11a7e
za1e001a589cc4accfff2da2afaeeabfe19d440c7b0c6212300dbf742884c582ff6fed4e79f601a
z85fd44b6a07cc06660a7c6b0256892ec87dee153fad2a24267d2ad32bfde26a066dea92053146d
zf31210ff69b8fcde39daec9e40da7d528ebb29ee93596b859554242f80ac1a3da8d762a8ef9fe8
z356d6a4f37f68c185137c5d8f96b145e231889546a439010d60b751b2178b016df714975477251
z13ed3962d7d6edc1df768ddc9750d730959f93dc8ce9dc3c263a5adefc3c71258a2772e6ce3de9
z7e1446dd96d48ba9579e308280af0bab2a423ffb2eda30dbefc087eb33df0aa0a09f56589f2d6e
zb08d74b1905756f621c7c77ef67127ec9cd9404300f2c0ceef2a4f15efb8246561774395bb3ef6
z8343363643283e793ecae7860b3e705d6af44fdaa383bd4fc179e61e94a7b153aa4428a14fc391
z11994d8476db042bd8522e5f8b83454fb91ee18c2be5204ee041b235c56d4fa8a251644c32ff28
zebc7e1b673e155e54b16797c19e69ce0b0454c6ba60192dc01d9519ed54509549d17431f82f1e9
z8dcf622cb1d0345eb0ca4a23480db1ee1fcc1c7bf2d0b1188b7b745300e6b6a2058d283ee614df
z605e64c57c44009c0bf56624eb6b7ba940c8e963206007e8138f02e919071a3e33c5375b0b3df9
z6d3d5e5802cffc9c999fbe805caff87388c44f005bf14c6a31dfd8aa42d3f86d2bd4c3f3ddb549
z2e0f44681a7bd17992234ccc8bc8e9a68e1c5e42842e9ce5499be01cd32ceedf48cbbef4277c59
z9d647f74624bf65cced8b393958014df29cd3e05f4c87a951a56ebd7b88130afcae071fe6f365e
zeec891321a2220811c909d9af83fcd5a067e9e9efcfba76a957c086fb15a92d3f9690cb4eaa206
zc2b906933a9a3868cc932474bfc5584c701545b2cc4441e62c3b73bc007a41b55a36e66e4c6260
z5c205abebe8111c74279ad60251fd595b255d23a98917c38fe167b8ee3f6f1adc035063fcb5563
zec25948303055c9fe07541085b1f5ec7531389259dccfaec9ce81bff1447d9acb4fb2852be79c1
z23ce5c90b94a832a376b7c9b8afe373729eb18319e947270f9abd8e2ac73d79feb85074a9a43ff
z9e929514dd25b34440353cb84fa982c5aa1620794ca3503b60c9c1fac43b1c5a1a76a355bb1bdf
zdcac4a2305b6078aa0f00b71d00134a37eff44b9b7a5f71f1553eb98721e8209c524d88b1b4606
z6b566034d862ab1ac9a6625f20fbdc266fefa164bf34de80763cb8139bb773ca1736c4f7d2e59c
zc286d393160b89140d82ddb356d3c40ea9c55e290f0e016b689a83e8fd2932df8582ab3e16c721
zf74d35edd9a94d3e23306a29a5710d76b86e5c92c8890c7770652f9778c7b06e447c1ff63c1e65
zc363c42e89cc0430d508482d5581ef7c07b61edb165db51769879e67eb745e489c1859801785bb
z7b7270160fae42c756d3274283321129ba0d5aa38a0c28af087a111feb9ff2f5d274f908819179
zdfc9ba52126a6dae19f3bfe780ddf98288920daa1482c9a0f5d38e052e2dfad56086065956a068
zce3b7aad9da964cd63b7ccc92f0c90cf9e09f69e461612403639c87e45248602ca5d83334c0dee
zc0c84a844961170d9a607a13e13ba3d7d0260d2245a88094b9095fc4bdce6e87b6e4b41052ee77
z2b78c53bfa176e80ffc7066c4c509d6da60525345132f86931308dfe18d5f12aa108e3ebb242dc
zbb79a19489cd4d817936eb456dd10edb5156e2b93efa7471c31717c47da18cbb0239254deb7e9d
z4c9b3105a969064ea1fcdc88a5b4bcd579c21875420c730f72d0fce1852f95f9520ca6c2598dd2
z1f364df7b5a0c649fe4390d16cdd8b3b121176e1cfdc6bd1638d879774f84c0f52ee192ceb23fb
z039264039084d918da21ee42b800a9e70534a0406a3c0cdf0fff7265cdad1a102b839424a7f709
z2d4fa0c6eb437645aebb42cd66803e36a6cc7732667c236542440976deea8024737a306a1d03de
z58c36828253edd7847b951b35f9d363b9ef8c6b519c63c6136fa831d19b05e8439df1d0f81b640
za086a34e654d78e72c7bffc080b771bac396b6ae6c3cc703e08c0c4eb1b7938f012a8702866cd1
z914caea80881fbf41482b744fce9f4b48db9d45a185e6002e345a16797c507850911090e825bec
z5f3ac8a8626f824628cc07585d6f697db495530bbeacb06e5fa2ab122cdb0e669ef360387f3e5e
z0e9dbc14768419e3a433f0a69396c78fa5cfce9b89b7e126ac2efb38ee8752dc872322652c1eaf
z79d838f5a20f3fc00bbc88bc28d0cc647d04b3a72911c1e760538977ece126c0f547780a41d8bf
zed97cf6c94c37bfee06829b0dc587b3526b6dcf3e7098010ca8686978c6f23c5afc2725662d113
z6e4ec1f04a644efbdb09e86b6c0eb91e7a73c2699866b26417feafe25eda58cc33afaeceec5c69
z1d1b2b0ef64faf7e7466c70ce2164704eb2892ba264c2983f6cb2978f2daf89cc7ca5b31d776a0
zcbeab63d0c381b6c2689b50d912842f419709f0e8c177105a2683d3af8a28a3a1bef03ea85f70e
zcf4998902febada2a73f77e76ab0abc89ffa44a1faedef64389b6fe298f7b50621bf8653bbf35b
zd2f6d3357a7f574663a819cf4b7890357706b575626b44edb01540a8eb1010618675f83881b841
zfc68e39109b5fb49ef9c21c24016af4846d5d1c1e188735f3cd518faa9893498f4c7c886498348
zf8f42c8875a5de68b0017f17cf819dc79d9b3c17238cf219d30f922a78011e39a0bef17c37457c
z3afa950ce176c52d7f194b4952fe552d87b13603b6478cc9e8e501e1b4f67c964d0cc63dbdb517
zedc3d0b98f61e6bf7679e4e27d5e88fc327350ff7302a1092c791a68ecefbb4eca11c24fb39abc
zb178fa4732c788292f72d463c5e2859f3f372cf8739198d70291a40ca8807356303353b27950b6
zbd069915ae23d7d89aa89351a6dbee42031dfcc1f7df6719c12a3aa7ef411a4ac0eff44e239908
z3ff6a6fa00a0fe0a0c4e2508edc4fd31d54da62ec764501ed8fc7d1773b5622b8ddd7a5e0a92ad
z3e4c6d0d02e0c305af003cb8db7ce5243cbfe1ababc071f455152f806e25058ba1987159256625
z2ab3a3a55d1421b0d451af139b65653f2b97987754a6e8dd0cced801eab307fd7819074b858d0b
z56858b48b9966bb1897dd0a7b55b904769c0e7376c725e599d00573ea401584a847982f2c2473b
zc83e8819f66178d321ab28e58a77f5f5ce96d31257fcbeb3aa11d84a23eb4828668597bfd0f090
z10bfa18a1d201e188a2dab38b6ced78e65654dee9f1b6ebc2857ed7aab8f2eafe0e6cb732435fa
zd1930387a71a79179459d29b0f58181c1daf64c0937858e63249ce0274931a875f887260d062ca
zb593b7985df4811987877bfdf69c3229b1cf071140ee768af847cc6b3e434f88feb7fe06626c33
z03cfe605804363193cce61ea2e9252ac29d78a09666cc336e16edba79e23481f09b215ed22e020
zd6dcb9d6a3085c6a22fecdbfb00d3fdb98faec332512106205d54814c5867e511de6f18a086ffc
z08816fcd556fdd5f06b8c3fc28203d56fc3556260d45700ba365c11622e1c5455fdf99ac38889d
zd3cd365c8f2f6e48f149df2d9d8553a91ba0100c8a4f3869bb4cf0d993d3397d289fdd80235d12
zf9fc97b20b15135e73fece60c1342814f03f69d65d92990361e9befa166f884048b5830ea7ee73
zcc368cadae3f5a4e10569677ddbec72f842b2447c9d02d4d4989167347005302f9eb4153e076ab
zc4f5998e59aaedca9b7380a019825edc20299f0051c2d68c653037e640fa3f8774d1de38f0c420
z371e77c275ce80912c2cdbeeb992b373b473f63accee96fef4ab1cb82686d1345dee1354a6166c
z13bd02622322337ef9eb00b282784adb36eba319078c385811b075da4d39fc13d25bba7549c910
z785253496cb22e67777e0020ba733268db9df26a122808088c50310d59a2b801854f53e5df8f83
z77031d02b1681179effa30e37ba52e26f8aa62982764b3fc76a0658d6d140bbcdda6f2e7052f79
z5a032bdd921770597172ce9824c403910b9d684139c7bd46f8b5412718fb6ddead8fb85f10742c
zfeb6674f4371aed3cbb7359d682b193f019885f63e398d14decaca0bbe206199393a9c74935356
zcfd716159a09d2d7b64b058a16c48647a9641787c74cb6f5e15b943655f217588c1fb27b1c429f
z1929e6958f861857decfe7ab79945670fa837f3487d95cfdb5c284c43216e4e7f001a80d76518b
zc89e481c8b284a659d3cb7f8d1087d008ac796076f06d68402803e68dd5f2613f7945dfa120530
z5bacb41e4579a2ee13e4023ad25b287eb6104f976c8caa82a3984b2bcc046f25c1e94cc7b86346
za98bb1e1353fbdef2eecb7fc19ccdeec9fb12a6bce75f11987f17460f9119d524195b0eba1eaff
z9f90c80360b8eabef693b07e368a818fd40b149d4e660933236360ea491edab4a77d3b92e30ff0
zcbf7f33670d8f9a6bf3c01042736ed02645e712541ecd2be72a78928cfe31c903931704f915e7e
zd97748c403085ac7e2e89ba97404984d4e67d80de1883ed26c42099ef717517d96da0c168e3bba
z6a00ef37bf63b896bc3ab6c092cdc0c3f03fa2ce76663f1433dc73b3e7884a2642cd9e73885eaa
z989e56c0c735fa28c122b4d2b16d88c6bb1049410f3a87319e501b02b87f83149d76a6455a5c7f
z6a4bcc71a7e1bc5b3537894a33804f2de195db280bf7b31fb477cdd0f76b8a6ea2a5b7a4c6f017
z2931c69eecd7fa794c5e713a74a5b34bdf32e88c0405c599a2d1d4cc5587a3fd112fd891442154
z748f267aee9aa6d4592419f8cf7196e0e1db1dfa4f45a5608e099697b484c68e8c188b0d6266f7
ze4ef3c13d8e72b057c35009508e7894fd21f83b794893c4823810bb04d51fa5c1ea15736750ac0
z588d00537777d1845770c4b186502b411a2d387d17873dccc9cfc55a3b56129857eb5827e8dd17
z5c81f6611896937214720cb4e8d1a9ba75633b630ebf17eccf31594d5436e82496ae4c9b1480b3
zdbbc604f717d37d355237b0fc9685412862413bb8db7b9e4b0372be6437e51b3e53cf8bc978e63
zf74a70d68962ec0c90f5444286c454d2ceffbcd47dbee3cd6b35891b81878963cf3824843a6b26
z85fae49100c6b9364677c53975798d4224b2a25389a956506af3e72e1fea1fdddc6d4fa27b1e53
zb55546665552067d2f667fb1aa1e4261bdac55d9d4da9329d1fac17a9189d559f01cc57aca9365
zcb77f8a57d2d7479e07b1ea94c9b8520bb6972547e3120b645985d75a8f9902fe61d3318fb39fe
z789e67e55c5728f60b47970d6cef287f44674ffc36b82245ab39aa65e6bf36459af9bcc94a5763
za2e23219208a2bf7b723e7b93bedc377980e6d56abfb243831f7a7c7a81d4679d84d993b8a643e
z481f88ba2fa9b14ef9c3533bd1e6efe552b791eda2fc5014a4919850a6968c05a751f75f265e9a
z5f7c40f4f8f151a75eb7ce5c4a5851b666800fbb1ec3df46991ec5a682de0a08a0dfe4ff55c2f0
zaffc4dc5b2e2d86620baf990497dd1bd3bb21e3d8440b7845b34b462d001ed4354038c8036f02e
z0f6da8315d6de306126f2517f238c4264898c48d205fb585e3ea439b182273ba23cd96b1210435
z3bc244357b93290310773239a1b78d643b170f0624d56a18c58dd100e6f645a6353985a706d2cf
z122533c887a5dd0a7776bd30ec17340ca87b2283b08368c6a29007eac3c23dd90d6e548cba9432
z761cc933f027d770d0f0f95406b42d8543b040ba213e76c70c343ceeda9c4b6ab009fce1185e0e
z02e9ea91fa564a6325b2f7167cdde5c687a052ea11367f4d43cd1f00a534f7230f5a00fc7d8d7e
z0c79c22f3aefb65c06caec7b63d2f64f4b40b9deb5fc80a2bba7cd381f4d25ed779e0dc1c86a37
zd0da64d25e828a5fc43a78dc4dbabed43fbe0563878cbb576c70fafc5a0619fd4b73e319e08772
z1146a8ec298a34a86d0f6a46165c75a22c8951d90fe028743c3b23227613550e45fde483951dc0
zfcacd65434b4280cd76c4abfd08de4ba81ab588ef80d87caa9711ba4a8b9d9762113d5dd2b94e5
z2f500b939dab03985362739023275363624805bfe265a4109a0f9265542bca899cb1b75e372437
z693998226aaeffacadd95f36d7dd45db84c15e9cb494fc27efec92120435528665eaf4a50c55b6
zd4d901a658521ba4e8f726a22ece7acf171cfe5d449ca69355243550bacf022d5c5c6bcf526830
z540f80caeede07f36c99af672d65d4c6507f0e65c6246386d47ba3cb2f723e85a9e236a8582d0f
zcac4fc5c0a16ff4e47a698d32a5c997d1856bb7010d3aa90b32c0a4ffefd66e7e6147f942597fd
z15e40c1ae7f5fdeb78973913e63c63364ec546b88dc05757264b6625c50b6640b0491e78f08f99
z4c05058e81d7fd324d5317e679e945c8848368cf3426ec60a8028757e3119f1d3e5c2710267752
zc27a1a4eb896f286078f66f87ec48e013084a3b9e6b2318583cbe26f68a8b05b1f6bacb4880bda
z2ee56f3ecddf78337db228428165cbafb956b9d9dc3efb41d5fb6e5a58daae31e30f294b14a318
z28a50bec87d068a7c5730d830cc28c07dbd4b4af511771274ffe80dcfab0a07c59c2b26081fc2c
z30e5fcf21f3c71cd811279fe48ebe210c13e8e1e088b547c2969b1300d0fa73d27a365f9f339a1
za60f7c799a4055e042c9a51d66674c2047942892d9257bf3e417e9af4bae5dd05d2ea87c159f4f
z2d2b1c05ad1bb5c56f4bdf9bd69465367d554872de4a48f0afc4c225b3c288dfc145e8ed58faab
zccf672f42fde66c555cec83cc43f2b7b5ecedcfa3cd796d07b688ee72e5dec1df493a83eaf0930
z9cb77060561ad74963dcce636b21cb18668de41ac3409f3fe3f014cc27ac424ea693eb7df86e89
z9af7e64b2d0c6ea37421f0f6903966969f886bfc4ee7086f480e02ad3d69f0baf77f9eae5768c0
z15e899a04fb5347cdfb0cde1e67ead186656627f3c963adaa8d35c9e0de576f39d90c9afa78c64
zf5269ed3c7cda8e6ec27f70e80506a096b2eaed761d633a129346e32fd13de092f4b767968867b
z419de7b350b884871f46de80eb82cfc00d7fd27dc65c66a399be560580ed30e780c7b48e47051f
z6eebb85992d038cc2fba63a556a9df3db587d06d482f4ce85b671a538d563ce77d5d89bd3c4b09
z994ee4068f7bcb3e0c674eede9ed1130ffbad24cfecf455b4cf3784183c96187ca21a9d37c81b2
z8bf1653835e45030db7f8b44416da0152dd60e098a865928f729126e1df3ea7c878a8c0f2307af
z8c523be9a7bed3ba388f47b1b2d52cd0b5dde61bb8501abc3f4d637eb7f0bbb9607d2224343ac9
zf21327392e4bd9eca07717f2241772e018bb916d027adc652cab17bc8541df1d5baee6731711a5
zac57da30a5c3882604db187b916369f755676498be889b3451f29ee1898dc07f1928766a897b2c
zfc4867ef17146ada238b808225e1120f5ba08fd7ce8876d08ef689aeb637b6fa9d67346c97fa44
z8b27d13bd43974982f3e9085c9dbc3677d6913410d06c48df9480af1219a7f15eaad35f771b4a9
z20f2c323300de5d065605a0a8e5eca9ae30ef4a4fdfcf26a42c84bc9a3c08d177c1ded0a098844
z9c2532b0a4488fb523b53063cba1cf2f90af3d5790fbd66533d776c7818b0541b87f24936c8eda
z532209a93bbbfd28a5744740cd3e4de5c11670896346c040a7a3b6b19ea6cea5007d0ba265a393
z2da715a977241df2a77f07afb146e724c3a64e2f47eaa443537e8b82ec937a62d7c0767550f7ca
zd72c15c6e482f1b12fa4d39d2034ea35668cd983aaa734ff041c8a655f2149a1602981d5ee525c
z1402a271f321698c2554da654b876e32bf92ef18916843ea08ad9031b815d79a685828c4f701fd
zb2475765e4fd40b18370dd5f791a48b5629506ba2ff5ac8a7a987ff39256e6f4f5283862c96196
zd9b12db531f3981a1d71d4bda8c4b41be824ee65b76d4cd1ba810c9d09601f2a30232e3b03826e
zfa12e1bf10725b78d0851f58cea5b2d0055707db774ae808933f33ad7da8e2793d2e4277acbc9a
z28163a5dac6c1c7ed3752486c9af933c5ac528e5e89e6c4fbd99e7acda0c68551e87ea52f384f5
z6c5aafc6df9ea441113e488607906087c51050c1efd655c8d5dbdf078f991de8ca27b4e4dc3673
z39fc5158cc6cf11f4131e848f1e1821891b431cee2a532ff3a6ffda3f1bdeee0eadde4312f2f0b
z7da805d764329ce814bd00454547b8394c67e635e856bbc67be6e1032c05ebcf10db76c465b825
z80b2b71bd88a4f5b9e6657595c6b5a47673bad76a11e323d4523461fda75010c3b2d2ccdb0aa52
zf95ea1c9d4b2023b8362f2306e776c5deabd2a5581c4c3f75dfece48dad8a658875176d536f459
z99752ad8443064b5956c97274d897bec5b040cc8b73c53d5e7587054ff0dd4919fcfbe246b76d5
zde0c280ce6c3c63ce5111523a2a58d2c7c2cb792988f1599c3eca65ea4b3b03ca17adcdd0c3de3
z63c150de99062ddbfc08620e582b6f08f94a33c61af542c185cf3f67795da1ceb99e2adee023ca
ze220304956922c6972fd9da0e6050430ae20be0c6888ce2c4ffb5538e10af082338f00fc8782ec
z674b33888adb04bd30520feb39ead333bb5b735f3a62757eb6650b161b36d68ce6cbf6f32743f3
z46b600d231602ad92566102e1fb44f1bcef82c266a2771b2144e9fb6639891864a0ed1eb9f4698
z3bd273bd3cf9a96604ca982671b0a65e7faf67abbc9ae4c6b5ca04e16569d327c3ff1d91675163
zcd1bd7cf6c839713f4d035fc02d913dfe094c021f19be672e93cf8fdeb65d7751e133df15a9fb7
zd6c0075601ef0c278b61cf951887aef5ea83b14950123c35725c46426dbd5c9393853b11026ccb
z2bb785c2fce849173071d8cd0dad8dc7beae127457e8d9cb56eba7ac2ca48fe0fbae2374ce5e2a
z1f609fc927454e75a41388e3e6d89dab481faab7fe1088f13b0d495fae86ca164e0058f4e6016b
z97fdc8f281081497079810583886fb6c929ac62f9d11f35848a235a63ddba04cc8872e7882de11
z08f3fa6a66c5cb5fc1c18846820d115c1aa7e1c0d09b646339bea1562ac15f24fd4a678cc3b731
z534382044376cf28db88c87d16f325a7fc240905967fb78645657d2f8fc5283d094e6a9fedfb02
z91053236917de2d2bf817dd6b071c43a5e6108d6d97989f4abd1b2716c2ca9706aa956ba0a7c00
z4863d7600a8e46ea2c6a55fa598354d3583ad7bf7127efdc2753a9ce9eb6172492a1ac7aebd0d3
z66e783836b08296074b368325c4dc32d04b5897943656f02c1f31a0b88cfed9440d1216f2d91e8
z3ba81e88811cd1c60bef9a56029554f4ab1148a0fab49f572c8cdfb2b3d0337cd37f6d24ea0cf1
z90ed910d2f81fcad296e80b4e8bf7fe3bf40387edd362af41cd182c0db3d91c5c05fadd8a00dda
z64331145c6bb062a9dd6854f31ec38ac21574bb0c5ec813b224ec8af8130e293ed80df88b7039f
z24551d39804b28b7752ba18f1a2a83fea30bdc87ed9d9911f0014f6febed84ef41fd32148ca18e
z6db2418e84be2367ca703ea0dc4215175632528d07458534030c30b6988b4691f75d420aeb06e6
z5e967045728b31b475a52393a9bbdbf3bb7699b000056eff61cc7bb72121e4f14da7e45128a6b4
z60cec181d69da536ea8faf3ae28ab150da888554b42d9d4027e3494b141ac1ea832a48e01ad2b5
z4a151612d3ac616369f29065ddafafd843e40d28422267b0829bc4c15c59bc6903f20437366e45
zf146406cb835dce145d287556e3f003ec6ba1ea3d241d3d210410c008d68b1a3ffce501b61f156
z9e2109d224decafff5f506c89325bfe692407dcc4828cf13dba5372a033cf7c1e0079f2fb8bff4
z881aa5c5831c8dd65b62b2bac5c3807db4b9561da08646b6da81e84c9cfe58aeac6d532479a078
z48e4ba836dab9add324d2c3fe904925997b733946e23ad50b1fd6b5235bced27c28715333b8cc5
z5e16ff24bbf278ad8fc5b51bd09d579af693bc08051de6e1d38f75d1bf88d7654b08fdcc76d236
zec4352fbd73ec6ee6599470f224b2d3ec236a57250d1c2c6349ceb3bc76d6ae5d6344e5d306a7b
zaa6717eac5e010ef420d717e5b366c9de082953904760c15ae2ef32b494e5ce0b6bac524b9a5bd
z7ae11c0d1c393f1a01d3e336fbc87f4d1ceed8a05f313985fcefcb4ab4ad840476428632b3d75e
zcc9d62c3c1eee8e274a2e9a2860521543bfa170033a8b3e5e640716c026706c975f599737ed927
zeb9bc5250baccbb2f5d9a8207cd6da3e709b7101212b44fcb15f95d8d71cb67b13296552a684df
z19608c4ae777c51a85f21147d4cf9da5824aafe440b7720a30c866e8bdc2ec5c235ee7ada0bc78
z741e7eb50096d7afc5ccc9b5d72ddce78fba1cec61050f7753b55b6c0c6a0cbd7bb3f0dbe7ab2f
z39879df6b1f804aa5bb5ba299aa6cd4b21bf41b790f1c983f7e84b654846368e5e092ab77d6b63
z7028db7031e8aa319250d28e70287ae4fc06480747a59707299667e380cb04aeef4139a49e9bb5
z69c79910fab961770851875ef4b7cd3bde2532744f96e728a23bde82e4441681e69dca901b7bb0
zdb05803cda49737231e295d020fe1625452d1ecb4434692199bf4dbe0ed0a7d3f0d4709adf4a13
z9d8df3a1b7e841252b2ec48b9ef0195133a5637d9691e17c8d15f28bf8070f7b48c8c738a035e5
z43206c3b32050a71442ea290bfc84f0bf2a14ab4d2cd8b60ed9096719f48ee42033bc41dc7bb0d
z3102344b65bbd796b43e9a98f231878ea71c267c05ffc9836bb8a526707874787445dceaa45a82
z604bb77d714bd08ccbf9e109962db6353f846e1b9c2b5fe611e806a4bdc8c4be9e307d5080db35
zc519ca12c04a56e9c5be8f810e2e55d6bd6f79e68222fabf8e7129d877a4512abe49c3424e59df
zf8a370f578b277b83b0a7f4f37d2f705e1ce4e6aa01592b69803c776785906708fd5ea07eaef02
z3ab12087f5e2260332dafa28c860c59969b0ae4956381a2f65aff725e2fd7d1dbf65de4144fa1b
za160f497971e0d292ef767cba91cbd272fd7dc3035e7d5171dd38f3da62370ce1a4fcde052ea24
za6b6e62c456fb83fbc279a6e0fc91e18e10666bc24b41444e45d5c0f841107b886641d17c9a683
z439cf436405c59515a1681b12977974fe5451d2a5e075a766cdffd64cbc54e11a19953506070f8
z1e90b73d0c912150968d4857d294d42686f705911846f4a267327c6f48880ca824e333e521dd31
zc7c5108ce1b4edadbd2541170e3e3641ea76cf9b4bfb3336d7b0d074a59fe40d091358f48ad0e9
z8418ed19082266b2fa0929cb2563849afbdb026386f70d301b2f39923e17c61adfe7d26c6ff11d
z85514e53f02cfbf926feef99aebe06b612a43d91a9f4f8214b60d0b19ae8946e26a7c613510932
zfcfc5d9a21aa11f1d7426a652cea680be0872dbf3218a35d5bb94903590f30dce8d3356933db3b
zcf0f5259a6091cbe0c04852d95912eedc4e7acdc42f731d85955b6cdfa204170cdc5c9feb3d56d
zbe6ebcd8325c8b8d3d7a861d0f35a71439f882ef47b2fb8ef918b5d5c4783e4b16a9c5ddd2a1e5
zdc085222083cd3a241237d3563c318649e8087d0f0c3a4c5245f224cbe4df752c0382f3b640aff
zc8df39c9a0dd1621ca9b9cbdb12a9047d70899c82d85c347b15bc756b6602a4038f83c67739659
z1dad0ff10bf6cd0b5e8dcd4a8fd5a29bdf2b359afcc7e2a8a4b12905ac38866c1e024a88179cec
z96d983c1bc3b359df0ad07c12acfa8cb355b9b7537a73945fe3ff38b412751b9aad1e50ed463a3
z7d302287b53afe1d11da8941e46aa1b6acc106a50ecbf5503581096ae857b4e8f06f8c01b9986b
zbf804aedf3a8dab60da02480bb37626c87cb6432e36f801e2da262e66c82da15b70df30f397ac8
zd4e36b10993ae55386ef54ae28483daa111e0d05817fc510a51e56382d26d3e4cc9e76ad292749
z868f2f8501d7be375e458906826c0e6a39ff184b62ebc0ab319af6d27c2219937966079ccafa73
z0096b06cf68b50587d4368910e5b1f6fab8bfa9ae355eb762b57ff75a845c089ce0be488ca09ca
zaff3634ae149aa1eeb0a3d88575e671669239578809df695a49860c4ee2fc1c657205ab602a463
zcd31699a0d8d5cd947dbc2a35390d4a2d8924e537b519387838a66ba4ffcaa9c9d7d6bd19a30bb
z1a3ba8bd960e84845896ada1e9b36c7d7ba91adcfffd4b07a199ffbd9a247aff525ccd7dc75c28
z163fcb401c314774025f923405eefd959d566013a018e9ce361259c5d64392a3b37495d8b209cb
zf8ddab0fd031c9ae550f52aa4df1503e982bbcd036bb2e56d7cb38c5b00591f7b2fc708d509546
z4e7157d92dfd2712ec830dac1cb02bc79b682db39fc6309a317b607f27f17d77448eefd16ce1d8
zd059c00f90cad1e7ec8afa12be6991840dc4c2d49093fcb753c0694fa4ce1e121d076bc948325c
ze8a7b4d9c188c407b65e0df9eb6f582d3d2683717c4113b66930d41e8caa701382b7cdf90c99f6
z5b67b397935de3eecab248d5219d8cda8279f5cca30ac710c575239e2c1e2961f3cf904e179a6a
zc4ad19da126692208fc0da5305e6a633f87f54ce1e41abec5c536e043252ac4fad02381b2e07d4
z0245f7987534f155207938552df3bb48d79903d601fa7d3d066f9a734a67f2248e5c3610ce51b9
zf799be53f08e02ebb5e2e1082bb2b451597c959717d2487a36ab5387996ec50e75b840e7f0f653
z266e8cb037f3ca6f956ab423e86b53a27b5a6982243527aa9d58a50db93b90ab55488889fa3f4f
zc9002baa86408fac700a1798c7ff48313b7e576e5d2d6b695e107c7f52215e55172965e0a7c1c9
zda5b4b128b68f3edd442ceb8cb95fe012e49c20e5c7778575d99dedfa5fbe51bf411f169a13ead
zcd3765369811ae12caeab5db6ce98053508b14929e06fe64084fea835ee1f14b6a5c2aeb3c7d88
z66b44c6661b3fbcb7547c0b1a41d3f532e56bcc1def4e2357cad6f9d1cd137034997009078b864
zfbc53f938846d8c90782b6de1bb071e2e5632b40efee97920bf00d1ac4b6d32de6363158f68466
z4ec30ef2c65cd682d26946245082ccdd35b4fb2f1fa59ed1a7f0c54a50cc9ab594405004592350
z377e0d74dfeb3c47a3276873e9452d118277b8e76ca6da9e6248b8c2ff6482c35be9ee93b6c391
z4bfb0b147e6fc7a27d37d4c084c71fe87d41078b730776907e0089e7e5c2a386fdcd3b1921234a
z36961f569cfd84f6dcbf8ec8fadfc90ee5fe8559a85feb27c0d40121a4f9c2d0b24decf3e7ee74
zdd4743af98f76288219fa1d6f4ad47e98102058c5d56a8c2a64f2e1891f6ad6975a46a62759432
za9d0f60712923a8260039b50fb2dabcceaecce97bd080114e9004ed39b8ffb671ef68dad8f3255
z525c2f3b814b2d113ab0e2a06d3d2d592dd55f0f6bb8901d2685a000874248f03335af3ec56b82
z10301c560ba9a169f69f6a402a5d5beb7196700fc10f3eab3cb9fff60dc1a9b7f4992237307679
zeccdfe72edbf87a98d736a2a934a8351471016cc7545cad97529b67273962a3977c85a38a8ec88
z66911fcbb505aaa400746350f58614fed391a6c52d5cba8bd671f66602cc3e5487fa05a6c1035e
zbb6b3e414a17cb292e6bc4507b7dfccd39e40b0316f4be66a0caad10be87c47d0902bceaf50ed0
zf43237ec05006b26bc926e71942d287e765152a8e9be78a5d524a4867eebac1a94086e75709159
zdb1855268a5843bd7786e6c135c6ba53b2e698e31c7eda9a2793bd7c94a0891505cead40757867
z394522be8a75190b861f9bf5629233705511991d3720c97a6587d568e84746d6badf4ac50f215f
z8102fbbca1cbc785c9c0ff0128a5784a03ac459f45f088a961b59a8eb578dcd4b7ceb3829276d6
z3755109ae877021c909d270908ecafe3a8730ba15b8f71e9eb93d8abb1c08b2d24272642f56a83
z6c5953803edfd8f0b88f21fbdbc3ddc3cde712eb2b386e9c71ca2d5780e23838b9b464fa6293d4
z3df63cf4f1444eff27ad57a40fa31c2211698e6b3891eee13dcd0b984d5adb2c5a7767b47f1673
z995c8e5ed5c80589772f0009ad60d0a8823d0751b52d49ec16de0e5d5446a42580bd005843a489
z81c6013e2a710f6763f0e31f61534b524953446a5fc11489e91481275d3a76fab26c3d20c9277a
za3d53635437ffb33e90b4cfeba3ca939bb98bba98e82347179e5df8e3478cfb7701915417bd957
z11987adee34ef20bbb2cb0375406f6372667711441a29120d92f433d3d7bb08feac4f836a122e8
z41ad64bfa048740f4927400bc9b8ce78bc19689378261b972afbe6ab32cfcc8efece8edc36dc13
zf753931392bb6c304fe2d09d9e355b3c5f8ce63c9757d16f3e911e706cb56cc142a29a0e520883
z3a4949b66d274d8a11126279442b70647131b5606482fe0bdb18e7ffc8f8cb231c5797a54585e7
ze3fb51877f74310613148fbc40de19f2f03583f7bd1efce275b88e25df9df4c0fddf9381382947
z3bd32f1d08e23529ad4cc4624ceffb6140e7adbaa7ffb628c4cc9b8ab146e862b1ee60d8741ca6
zddf7f380d6ab94f546ff5a3e1199b540e35dd4979e925404cc1905a4ed537346be1c0636691848
z679aa681bcd722cb97a1b36ff7f6edfd8f7300ee9e2864450b7a4c13b9d32dbced09cc16980214
zfced09dc5467de851c685e4de68c79bd9ae1cc9995be9f8da8934f9fca80b01648098976b027d0
za38530cd4d91e4762c0b8d0cc7b99ed37f9d9027d1f816232b3a2d6fe3742e63afcc2222fc07e2
z87856f5da6a9896820e02f5779b4528ae5e3f7c092c0bbd926a6df02ed7730eb028ce825968a01
zf28f573a9719dc3444e59812ddf0220cf737dd3bbe31eef2dfe62cac2ad55e30af822f4e7abe5e
z533dbe19033a89315dfcda5934a615e1ea8e64b16e197cc9a88732269c502fecf4e32c4097b977
z0cbacd1fd719903e45e2b3dd118674c3c0e247351287c9ebf013ab797f84937a22ab3dbe2f2f59
z3addbf2c4488d574e007bcae280f670018c1b4dd8eb3fc8579a214ff53f9aa352471483c32f3b7
z51186b51bb82b98a94c98307e53fdf42a6daea3a96b73a5e05e85cf0111b690a90e94f896a1bf3
z568eaa905cc12985260a6d15a37e945905540a1a0c3f1b99f545cbf45c47f46c2a0cff2c9f1409
z62de1229e3460e5dfb161fcd765a709059a25f353a1941d20f1f1a5fdc0eda5755b5f9d75f91c4
za13f4bc01a0227051c0a0add75a1f1c868d4296c295d5761aa73f2d1ec49369d7cb5f8c1da2574
z3c1b02d6864575017aa7b41c9819453f7b91903782866b378cf0075739e5b971ff912c6e8d2aa6
z7aa99eb9138dac7ad85126208daad75d1591777621327da09273e90b6aa73827374e5bc07095be
z2cde33aca579664afa93b78fb7a222f4c00e7a800735034ea5514b6b395a69ee258091dc4290ff
z7c6bd148d795268892761e018a596cd15b52f2269f6e54d32ed6b03abbba8e068f7b9520d257f0
z7456e3d32d969815fca684009389b373da72e8f7e717f2a5c2365c537995c5a8115991bb832439
za260199f6e65e00c21ff56f1c788f410840714878aabd49bca0f7f602be233309783446d7605e4
z030993d21c8507981b2c8896ba3d9f17fd82714890bf8fa001ecbbdf230c42fc20e8ff0c5aa65f
zcc6cfd14e2199a81056cccfd5ce818a39f3edb765e540b2819579b290daa3e86e451b7aa005be4
za7ee7af13a1f6519c5b9653eefb57b2296b652f6d38b9f7fa2c9fa3405ad9a0161c0f05f67f0af
z3fe31f5884e5d72aa80324513ae5f6da9cb9f2dd7694d6b5bf9de35ab8d46493c198396f9509c3
z4e9f0e2aae99cba75b92847325e7c5eb72fc7623fdf681b602ad0a26987fc5bca3ea37e133c881
z1474417628eb3e2775cc4277dfe1f43e70abd0d1f0e0589aaec569f1169e491187b753b605bdb8
zedc4a8ad15e9680f03625a0b901b174eeb45e10549478c639072d4981aff1ef73504ba64a6ca77
z14c8ed1b04d594976b30421a39243e079491e8c740bdf79707488d2ae469ee2ffddb89e88ecb46
zfef4393dd15e8fc5301e7aa6a4160fd9bbf2288e5deb67bfcf442623af030940b1d4aa8be48097
zcf454c3fb7fb754a2ea8e01f86edcaeba71587645160f81cc1daba959aa561a392f77bec8806e5
z553e2ed03ec0d21bf63c2abcb67761df0e01e05409673e07d5fc48ffc70085eb6c760833c1f560
za1dd116e8249732f615e1fd1360cfe2e4695e627ef724c33f5c70b80b2c311ef55821655e86510
zfaa777f4133739f8cea460bc14cf9728a19dcd923bd3a078db20bf90a8bd235ad16d1b44fe3d6b
z8b9008352c3cdfdf83a29781c82d64717d3f709676e3e72f6cb854a432ce89b45d0a2100647601
zbab5be3b43dcaa5bb664f0f91f1801d7def90a7e4098d2bf75a3b8cea0dc21defae976e1a1a9a6
z9d5a082d5896b1ae119a491ea931395043817d42284a8a7d85bed5961fc9b0bc2bca1518c089b2
z6702f0a7f9d0fd73ec4773c1d28a29a28ef973ab4cf790e4fb155ded5ace5696cfbd9d57af3184
z57a3ab4af91ce915d7b2348bdaac73b115183f59f4e5792a257ba279b21727f82c6e71dc732cd7
z112eb810809c681d1063adbca94a2aeb46186c36123c3e38ed1f43849c1a2bd4f9cd410885e389
z7d0db7a045ff7cfbee776d5fc1150b323e17ddc68c9c001ced8fc1a05138e1acf8b2c1a492874d
z3b07eca236bc8e4a9382ca9fb4f13ce21bb36f497e8f0d9d19a2c53879ec0d898a4cadf4dddb1d
z2b5e9c1e388bca7cc1fe2b9a4e64d5c2319f761add59770590f09db8c3d7b28e4717afcd265de2
z000e0432a9cecc61b1fcbee4c45868bb350a7038a4cde3aeead740cb364fb2963e07f2719c84ec
zeab7217c8c38d25c62a4235a1540b66707d1df6b328fd4df64f562436b5f1cb4a6c08b91578127
zd6340f256d0a3a9f86349d5f29cc3aa02806143e80a289f98b6ae621cc4ddb024b23f8617f6227
zaf62eccd9a9a4c3c6c6d9414ad46d3f80387fff4e161880126454839b9b2cbfb3d10f960e85584
zd1eac4d98b220d7045bbc88840fca6456f36803aac7668ed4ab59212abc203c2a83ca6c41752a7
z0c8dfe1a2aa1b3007da60d8c077a7900ba8acc01fbca3544d4b978ff0239f9234639d5da60a42e
z1109e6bb50a5dbef006c9a8f5c6bee1576faecbb4ebe55a4259c763412c39b87b64ad140e64868
z438cd29964785e179ee8b1f20f617cc57cb617f64c83d96f4e173f6904053d20bfc515276c9c87
z2f87f409cad02c3241bb53eb03e1c549a09f3d5950f7f4f83e4a46871aa7e842acbc87d3670f21
z57656adabde0a3404b952499cf36fa89a099d839803dfa385dd89299ce5f03c0d6bddc24b53d13
zdf4526f5d08e7c76d0511a717b7520b0535670c3c1e448c17d4e1f7d714597ad776baa701c9618
z390220e15be30a5d8c4a5efd507fd67972a4b71a937af417d4c4eb962ee55eba715c29c3a2900c
z498e52a20243d572b669c119bb17adf4f0e8d7ff22db0f535c6b63ea803bc883af1e8eaf96b8b3
zdd4762f6c4da71ddef8d048e33aa06265435f4be32af9c0aa9b20030d78f68ab875f0d64692a9b
z0e6dd5e0ea559d5b7b685b9f1e0e16b0917dd475d98445f3a67fa6017ee1a229aefbe3b1104f69
z83595bf63f5068474452d94ff53060676628e408a064d4b5726afdbd09f7086c11892d538a839e
z8b7c1d208f164434a5f4e30e445a37897a0be69264a8360a6b3d1dad6f4aa3ec5f2bc6055e9313
z4ff1b4c09c06a480215ad91de46ee8dce99332604b4a0dcb1d72719c81a5e1d97c8707d9ec470b
z91ff27fd909d0ef74c90e80df36cfd5e1fffc4d32c5f3038073ca16df9bd99c7ec90aa4757b684
z7a23db6348dcbb3be0c8473fff8a64b054ab242a9e9fac37d54f1f82348575c9fa38dfb324a82c
z3ffc56ee25d4d1f3973043f7591ec1294b9eb6e7c4c3340f1f931667bd5f14614ca230a1e6011c
z81d37e07cbf0049fe90a8c089abea7016f8aa3941b6b8b56cf82a47d6127caa81753b054612e3d
za23e269e9d68833c141e9aec0cfe364c8a91d5ed8fa6908b9b5af27f4dfa915e03171181a20fb9
zea4f2bc43ccbcd770354eeb1aa8a564371fb518492237c3fb38dfe996012ab5835c4170a528d13
z57a8a4587e905e438438a178dce56024ab63bf4ccaaeeb02dff2920c64115e07e5ab86146b5010
za866f8078e9999434fa5ed762539a64b3f2790198ba349199154dfcf6a9c4b550a3eb557d1d2e9
zb8d244e11fef9e72c2e0a91045f4141e68da9a3cb621c6167a8e1ba341daae73316eccb4435560
z87bf1f2e3a87f57c31e6c59217bae9c55dc85f7890bf46a98a4d73b68be2d18057c7faf171f3ef
ze15b219745be398bae81d1c04e819a6b582f6ec2b8ed338e2c4a3643446d5b502b884d8713d89d
zc872edb49313ac40b3454151e09561527ce0deef7ee5ccf4e94628c96c21c6a8f0017752d5562f
zed2b51f596329494f70b158fe66edf355eee9c67d1ea8ed58387eb8644f94a5f2e7504d27e4b6a
z3857f393ed3478446e8b1033504c2f280aed576cc9d0bc78b211b493484abd37b649b8e62d88df
z3202a74835fd619d4d959996897fffae7ad1dd9c71288ebab350790a291dcf8cfaab5d77cdaa4b
z188c86d0b6f6e57d497c0fc4185fd84e02492042d9f15e2fff386ef4908398b394cd9d5df9ee04
zd0134bf2be8406c7c08294a15bda81def2df1572c2a072343cbc959526a432b0abef704931541a
zcec2d760fcbb95584b6210828c149902f1adc9f34b11da114a6e373f59c8291bc3a1a7632d6291
z04e84b23ff06e5051ef4a07ffc516f214d978c7c2e18046e60d9dc2ca5b9e28f229a7756c8450b
z0db620a6a0a609273b29225887ebef25d000e39f30dcbfd63087ca84b13553d766df4005b241b8
z0af14dfb4c59905c4d863a5b09675f03b89f913a550a6a81a44efe04eb9068e61d1667a60ca257
z693ef5f142715fb2baab9520c929036eb1546be4e5a2dce5cb7d7f6af222256516d1676f079d58
z22873e49758a73e7cfaca4603bfb1de087674fd617237946c62bb5f7f36bd54d23a97b1a5532ce
z40f6e22dccdae6a22349efd1c1b85155ef97d6703c7c8f03fcb33528dc1a84095a2eaeee1b8898
z3d8a39dee141fb6819228ad9b7dd4c5b74daa425d64151e37a0d7457961d4888529c083065d7ab
zc3091b24fa4ee2579e71d073e68491c7775bc124e8f9170e3471c1cdeb50772a7a61b40ce9a156
zc48426a67acafc970a0c9e679a3e3ca80233521cff32f13fcd1c2ab691069d8db0d2672e321af8
z541db9a6cc70cc40cbaaf73a947732f35d4707dbe503324c64f9665d17c7e68be2d1efacae49c5
za1ba8a63796520b6dee7ce1bec8d26321c30f1c7a4539c91b96aa2df8657f0180eb1ea837f3172
zffaf48153af127c59081f40a557903f271f998c1f9d864f9c6951b9887d6d47ed4bbafd43c9f25
z040ef9d6f1044cb0d3ea3e77a6ab7833b965a7aedc2f15ff490fecf5c2579ed991e35858014869
z548dd66c620b6f25b2bda11a5a817d912f92873fcdeb08308a101ccfde1938fbc9871d16578401
zce148a9ca6321ebb5c0d69056576a4e154722c65a3bf9c48bf5f6985d36b1fee469c76b2e62fbd
z29ce69d5806ba4713bc52ed1cd3f517f867a282351c4bfb3661050dd63a56b5e61232f3fb2ffed
z5dee071f7e44ddc7943d947766811af4b51ad6b57beaf01101d874e2ea71c2682db8a68ca2569a
z2573897d434b5d66a8f7ea1c708e51a922f2b6360b331d3c267917bc55b5a87c8ec61c2333b910
zda537b23fb9fbd349ffabd4514197dac6015ff5c04b9d8e1745f30b681628cf6bbb453b871c894
zb100a9da547e349f3809eb620b20b5983e8b2a9c1709b0a34240e7db27eb31ff5e80da7b29da25
z06f8d787ce0c22571e9acf0fc0ff4e4754dc800a0e6b9361b1ec3ae6f43b34ef1b20063eda782d
z28f161e692eff3a4c5c2d1f1703f6e841bcb98ecc1fe7b88ae04c1376aa03ab67b19f8898d9788
z85456b62c5aee308954c21dd8efbf256da938a91e6902811327a1fab951c231cac8f9a41f33d21
z7c426c0dc7f0885d9e9b53f3944f5970d47eec1e17292a48e5bb6f307a4c2bc3697df19011fd8e
zf0ab9c07013c5dbb29bc6830e5eae1e7d04192fa65850b0a54b14d044f5e7f11bf0cea23198203
zf76f58d246ce81f4445ace92eb09956f2aef6707f6be2977698757110543a66ba1d24ba2c78d02
z37082f430940abd8fe9bcfd085a8e6d3eca05fc4d9806cf29e2702d473c64bdba8efeda21b846f
z783e4f996a1fadddb08ac809b3b27fdabc8530d434b2cc6cedba622a6a074f897f9476ff275887
z02864a2f282a86ed5b5ddff0af47d3edf31e34d40f188bd75b3b67f12fdd979e46cc111ae5f57c
zc22169f0c913b171774c71a2ecd99c6210b47de97208faaafcca8030bbe1247395ad8a52caaa56
zca75243d02da82cb8b4d217aae169014e8bbbfb875aa5a03e9e73e10d0527a63f501c74a1d01f8
zaacd6646a79a969427d66762e7b78580490ae9ac4cc9ff9499422be7469635b1d7d902f313bb76
zb26f325861ddec316d82c522d76da491746f926f9402477cf814ab4f7d69d275450eb8dcadde8d
zbcd4afd74d3ff959b5e91de77c5f9e27e8b2fc281bcf55d06060397b3bf32dee894ac0e6b30d05
z00508b4f9010a70bb5ebf54c349d2e56ecd6f098a6e96e68a46143c8f99bde251860f50cdc12bd
z1d4facb80bdf05aa24c23c05f0b0d546d255923db5cfe4b621ea3aed142a2d4efc339314a8317d
zae71cb157e1ce4cb3ed8b6214f5dc5b73a37fd2ba4f1fbc7a4d8ca127d27cc9dad96f8b54fd62d
zd0d07bf91cc26ed66415a0551baa7d4cddc45ffc4d784a76e540fa8304a0f620fea6d92dc6f5fa
z03b044491b10b6bdc15666ce0e4c65fb8ad602962a666f30c68846876ea95fa92b0bd6902f0771
z4e2989932ad94aaa0832cf8e1bc74e37008bdb4bb1bef4e1ae8da21556f0752e36c9b90b1a53cf
zbd315fa7f413b6901dc3b23a358346b9bdc22a380964b68455293314307c8194f4d786dc6cfe82
z46f9d3f27607155c40e1a37aa32527bdbb9aa8cf9eb43fa49e8bdd430626e74b43429e7761f7a0
z15e0e42cc96f9c5fe739e9e59e4a7db230f12f6b8cf8be66ba5b29ac8893cce79efff3a591103b
z151c316d2fecf4d921fcae44a8d2510560839263a318600881bfb1856536e218d9fc85435c3801
z0657783e8b77e8df62c2d4b7b9fed9e4cf250a83188d5b9cdbef4bf74263c4d657f2c292824701
zdf919824676d8b143cdc0471324514930d513aab13cf578c879f9a10d4a2739d755caf776f68bd
z8f487b0d95e73f42a9bac6ab630ec9db0b7ccdb2c2ea0956113e67ac0dba829b697e709eb80014
z78cbbd5cd7486b243587e4f82869483e1d74499a2221b24a1a70a8871f3675151f307269ad46d7
zd0b3855e43eb8ae257fe269d2255f3571db867360865935a31543e8403379c352a83861c5dde19
z55c344bf7ba5d2bd88788085d89834f5b6efc8ca169ec7377ad5c90bc8df416dfdf93d4a5155a2
z3fdbb66b85724467bf0485a638dba1bf66ae8a00e85914295b2f2e866cc93396ab7b623a7a3769
z5d01b84df6ee8ccd0bb4d934a1dbba6933983ef5dc3bfb44fdf426a5165379696610514ac3eadf
z0fdc4957325a069fdf0bc9ae529d070b8d6bdb3d89c74616f5c2dd3f677643efe17f44df5e3d34
z24612e7a041609e8d7802aa7bc8e697237c97be2aebd98eb51fa699d65d6a2c7a7e1b02c00d660
za89f84c02922f62e430cf963bac6bc86d399958afd90a3992f2d3f897154a45923d3e437a1e0d7
ze8a921a66bf641c9a2be02a0efb823743501f8ffbff3e6e3039381de60ff83f581c8a36fb12643
zc187cdb8c5911b1cc7121ee86dc60f3ac57cc1e679c54e4580fba40edacdc3232e466d489c5098
zbe67cedcbe8b5ccac50ea63baefcb2334744329c63cd1db3a00091dfbc4d3854d493ce267248a3
ze05e6931691157d456e50392e7cd5bfd2383b4c6c98fdf87a8b56d1cb7ca1c56a4d3b0aa306923
zdf1a18c53ccd756e10645a1a8e5ff76e7d68c53396e7953c55174fddebfb4e28a3359140366d08
zb40678226213f24b7e902c9bf36a034773a91751d2a050729bda3e2e4f3f1d74ccb3a771f942bd
z1a02046d03e31e59562dc172ea4e8a7df3f6d642019944aaaa42b9855e6dcf91e25257f91d3159
zded08d9c93e79c8bf6a79df1c7ee4829012afb6ea61b30e4984143249eaeb8bcc896f4a7e7e3bc
zc5ffe9cd5f68792d76cf1173e83dabdcc85179e096ad09555453d12e03c952ff6d3e6f255000ad
z425551c86d7d849ba357299e2f165fb6b3600eda2a1750ca85e11742ad3585ef557a577496d012
z2e7079078915de2b0db498bfcd162074771f5e4a78111ceb5b8a7f5b39f970f30b89f912ff4b7c
za511659781a4fbe9594b367c3d3b40d31e389ff482125c13f070c450bb1e27d7d919e29d75191a
z00c1ad4a9a37fe6c8e963b75fc5ba424a84dfc51d4a6cffb943ddc64439de5232770039faebe44
ze149dedd1e6a6d13dfe2e697b97de18a901dd232bc4bcc5a70da2de1d0122e07169a024d2de4a1
z926b1f61cbb11409094f52db9af304649598f0c86743fbde46d84de9d32c19a6e8a1b2659d759d
z1a2271cbe653aaceafedc81b9a5ae65558741323fab09ea97666121a14770e575e3671fef2884e
z47ea4ac89a3516a8f671edbdacc068ce3ce0cd24fb97c07fb2625421888b7c973411591913ab65
z25814b78bab455a189bd9b42d712db0166408407f40bd1a22a57aac484b1f2d8b15737bb21c0f8
zc9a9f38e8f62d18cc61c28275f8b0475bf680eb828cc4cafdce0a00f56b30bc334a1190fc6ecf2
zfbfc8308aae7ad86072dcb2eaac7ffb07b7faca533a978eee2ac506e4bc3fa7a076a589523dc98
z44b114baff75e9086aa2d7f8c3ce7e58466c7951eae8e051bcf6b583e9b02aea3a7940a5aa6ca1
z57160aa19fbca7f9b34f64d75df2bf8fe0d2738d40f7db92c5772ec9da7ea0802a9f8259d09560
z36f9ee619c59b57b810dc6a707006ae6a735b5e942c57fbf2978149c32226ac3bdf184420cafa1
z0502f84d3e8ea77d87f6d3aaf71e86e4ef09d7310e39030371ff26baf7b2f11c8d5cf3c46ca32c
z605b2ad096e86bc1d2cc292442a8d30d770f09af9e51187c087ea929a00ea1e71b35fba2c5baf9
z3aaf10ac9a4c2c597a8358cd8e9a9e8af490d0ce282fe3b0dc2f1f6ae36776fd170d01d56872e2
za3be9a8ea9154c385daa6391365f14936c32292a404abd307fd2fe8713993be154bd32bd2f1d63
z965c565b8c3d4b2f59ae4ef8ec73a6ba6fdb9651b53cf9e6aff3208c8288ec863abc553ea315eb
z3a4ec35cfd35564897ef9eaa5c7427c5e697850c52cc2b15cc072352952b9106d310793004971e
z3ee7745dd3170a6157a6d7463f016026989832648c2cc2f937ea5552a1e336ec2db6f92cbca105
za6be6f305efc4b569ccadd6507880109f557505d97f7ea85c39ce411ae58de9d83aadcbdea136d
z479675e5033e6cd2ef15f0c7017944b6fc5ee5115ee120928bd2724b4efaf5bd394544c7e67b02
z8e1f821960599c4289c46624c1d1264839d9be517be32cd82dad3dc55c378370a6e89444d89c27
z06b99c13225c34ddf44e416bb2fa375ac17d176600458dee07c314442b8e3898e6a5861b27c00f
z136f2d3c194ea3174e122953a9ca4905b4ee19eb4c9c9b1fb17f34f1231e57dd664bda3a903482
zb83ec38e3584bf17ae9009529d24e9918de1c545bdb94463ae6157d8783ba9b362191668ecbca4
zd394c405a2502e90581a11a5366160d22d39516f1ec1c7cbd731ecfa5833f4cdd4f4df57b82481
zee12e660dbf6d231b57c9a227afb11ad055a0193694d0e32e5f5e85da93c523c22c046b9aa1f29
zfece7c898579655269f2d16515336bbcb4bad13720d9483358fcf748ad8548d7cac6f87ef07ffc
z5ab1e99dbbd4be6fcee064c8b30bee0e7196317cb6ef86e0a2fe901d56938f8b05b8cc5dd6bf3b
z8dc940876df80f618ebffeb9d2bfc84a5c9f460c9d0e774da96e8bcc5c2a70b2d2cd659ec62ce4
z464b0a3ad6c3049c50ca88b7f7e82a0d6806e85864089d13dc972ef92b4865b7772131964f4d3d
z71ffe0b7303c2b6a7098e96c65c27974e7194c4e63ab78925c8480dd9f8ab0ca0551495c8d8aa9
z1a467f71d845312f8eb3fbe22a0ec951f353d87f823f34849c8568a6cf365df200db6de9ff6a6e
z48422393e12c5f0a9680d80dc67571b095ad5ffc7c3ebb3816293d5fcc06763a54811df3f5f415
za7f490ca9befdf919cb8abc0de6d8025893f1a4e4c809a596cadcda0749037f2cdc620a283ae45
zdd9f85820c6788eda0d9e075c3bb25b0c7cd251e9d5c3befdddb967996026ef4ee7da4b193f9d4
zafe42061968dd23ce40b187a2040f21638bc67c67bde198da1392d8ed7e39e98fe1a4dff39bfab
z029b3ffcf5390e5f406fbf2c88ec68a805608ceada3969a4432b6a9e87c75389cabd3854145ea9
zc2852fdb96834f48cc274950a31fb84a02ff309713a01d60b46301243f2a496a59902daa40a299
z4bd44985ecd7e7cfd95be590dbfc0855e6bde7684733fde9dd983d6b0fab261d7beb94f184e745
zfb4f8310e1f100eb8ace70202f81b2aaff575c7a19f911423f57a33a28ef1061f1682866bf74de
zaa9c2aef6f5029252d785fd53ede34b6ca8006ce53db9799fcc1ed11448eafa10d2e873c724dbb
z210089a1c6fbb5360d43bad5f98420c8189b9e3c335ccd6c192f878775cc899151b8507294d4ed
z4eb2b5d849b3dc8db41965bef30c92ce777bf0f14f826b2afc102e8956af1c01ad5fa776cab2da
z668d4a0d3741de39e30837c8333a7b629a863fc4d543700561a5b24b0051387c00f3c00de433b4
ze741c8ddd8515bc2c8b7db13b27cfe3bcb344fb59b5607d357789dcc30bd231a679953e193e1a9
z9574596c36d5d5da538fee5c94858982c3789e9eda8665487e55ad0d6984605330ac738cb97aa7
zc852a174aa8972305103f604268fa9403732b6ae348df65d5c34e4fc10fecfc34c6c2b8e45b464
zdeebc1f7ecad51e89c365b065c7171075eb74c7fbbcb888942fcdd30453b3c29c64d54a917472a
z4eced08fb61730329e7b5922d1b29b9359c3cc8201f5157046a73c1333947808e1b0641d9f428f
zd58678dc6640f9913e37720403172576647cd168798ec25627ac299f87bd04ed1dbc11594663d6
z4a4fe44d500b6532eae482bb69e544d1114c9de4b5c1a2142a68fc0eed2b4e893af95ab701e1d5
z0b4e8396652e50fe7cc90b71afccf9236f55f007b199036f74d53173e52570b0f166c41e6c2208
z220cb3d1fbe6c1c046975ae4cb191e9dfd95e4522aeec95cdef6e816d90d79749e2acf0fe5e9e7
zc53a803e21ed9e2686eaf8b219bb40d486355002c24609e63b2c75b4049e81c58e2f4511a5ed49
z33d0e900b2da3e6edebed632c6a83326c744db60cfa21a96b5629cad16d17c16079960f92e07c1
zae4cdaa11f38b74f9585abd73481e2cacfa309a866cd05d059ca3e8155a36b14f90e0f03e5701b
z939dd3a4a0a117c03ff03e0c0e566c1fb1020f967b7907f958bb9201c3edd6ed62d68fae5b8396
zd4d8a2c8dd3bde756e18d50d4aa9d122f99d445305a888917be7bc708fc8a226f686dddbb78c2f
z704a8c4bf06a0916d9642138e5d09994e1fb90555f0388e3ddde7a3f9e30b7384df972315bd5b5
z36a41c304fd2cea61248235b619be14f15d5e1cb7262221dd8e9adf57175e13d5b10a27f803cff
zd17e035ef970fc86738817737ff740ac2bb85c34a1d60c6005f1a64afc783e493769547ff57561
z882f9cf567fef3aa82310e44cb07a97462f2e1c505f76939aecb620f8dcf0606f99857091e4797
z1718cf521ca8a0b7346d3db8a9431df07421cb7401be3c2104b29cab243cf148ee695242f445b9
z945932102164963a1ce5166e1aede8baf7af97b26ea8e42a26450d1f321d92fedd4d0afbe93e31
z75e17710c1374f6bb17615feeb36cdc092a106214e52f38b676e92dd873ca7742855616ea9c5e1
zfda876ab7a4e0c876c80da95d495e33968953846b19d8fb0585e517ad6c89b45bbd35c9654efab
z476455a22c8c74c1d2ea4ccab59a5ab781768b5d582fed0b0ddf8cde362f53f6be6786a67460f3
z3f7624e087daafad261d4ae6581b609538dbd90e2230b8eda8b57b299669c77fb4ea37e7213d98
z8851e5a2f131997f5fec466146d392852d2ee35726aec6bd161f63f8a7428aaac5cdff323446b4
zeb41ff9485ffe7f2f29cb3fba4d2b8c550aed93dcf3a7cfa8b389fb8dce4c9e57213cf07d91719
z41f4966f41f38d171e9be505dfe12c03ceb33991089c72c60bdc43e920172dfefc003244be5499
zea867a05d16e353e90ec6640605f739b672e459acbd89476c2a3886b7d7840c736565144197d9e
z2bf816c5da5e6af54408a0a2493fd78abbd275c84b27ab610e1ccb3c43b4ceb9ef38c8e7dd7380
z9a9e5df2e38b158e24ddb85dce91994abf02c95bd35733fdfdd0d41437c9b5ac614b3abb180a5e
zf818ed53e11c72128dab7c3b91e92e0002257960805583904e64742dcb74151a59f9520d6a3698
z25cee7c083a51e65df807925acdf88b82784646ac80b94fe3ebe6d3f068a545df6761112842e8d
zd1378fc6be53ea477af7a2d5014648f1f875572512f3dc14dfa48642b2c4ede647c44e3a73d3f3
zaf03c7c496bdb509ef44104c36cd37e085763a24da22720c6fda66aa4ef8885759f74dbfbe7684
zbc3aeb559ab714dcaaa46813c1b86d0b4993b28d5f115806fb61dff705a2b0ee3b8cb3fc81304b
z460d66e7d9816692455dbbc9b12ada670068dd0c484f2686f683f1165156a5ee571ae8ce891332
za4d197b7913f3943deebdac4196337409cc62bb489219d934587a3cf5a701b55853720de3a09ce
z6393a12fc9db0c9d272411ca143aba3109d65e9703ce7e7420d1abcfeefb9a4e96bbaa3156a195
z93af77809cc9e004dbbc4de0a15735da108d7a9336be7f23e52af695f28dc91f06de3dc0cb5f6d
z8bcb143cb761d050d721c8f4a80b2203612ea1c74d762bd1d453c6a1a09894775c127cdb41bd7f
zdd5065b8b455e91daf51f768465b169e293684e6b71e0b269388404d9bdf6e4b175da082f06fcc
z7e5bd1a4ff73eb9c93579d01a16476c109621855e3cbcfb918182bdd8788b2fed1b323162215f4
za76c5732ff83aaa6cd8772f5a23601bc619d6df55f67e8107254fd8211fdd5e9d49c39b2b53564
z3b850e1345d12644583e92d714ef6fcd6c2ebad0c0e0449cbe8401f7eea6dd9860281145b2792f
zf0b2fde95813eaf53cfaae7b5ec713cdd17f6a2b06ee10b17f28cb0b4306b7d636d389b4da63a9
z0c8ba0ded0317615d31a7cf4e8a339876d15917251f097920f348401d3a6dc9727ee20f86e0b81
z1a6865de0394efec14cb8c50e0e5daf8e9aa8623bfbda40fac3d4539dc4212da46756c3be0a0ee
z41add46d4fe7baaa565254341dcc3151c2d51761cdb8ab43c9c1a4b4d5f17302f10784ae0219d9
z855b4cd6f3ed7c81d5fd38cb151f794a99c88d0a0ae9f7652fbed23aa27c3ebaecd2cf722b0a72
zf59285c30e6c8a6742458f57472dbd17319e19f5c1554d4c29895332b8c0a31e29d22f8a07c447
zbf606927b1c12055ecdc8bbd69c08d7d9b4e9272c292cb8fd487ff22f9b5dde87c1fb89e69b2a7
za8c9e3a4a354440fc2bba69357d61cb33132798894cf3be971cc981444f667612c5f3b9dc34c9e
z45527db6e6aa679d54f2b80213a826cbaeebafab6398a68cb6272ea765e0fcb1ad76dccddbf976
z0a651879b352bc19e6f2c91940492a106b30043b6c43cf2db8182e569278c31eb88bdf1b496c64
zbdcd5b6be1b6fa612b767bfa2d1848eba0bf3329851088827882527afa46f42f52994cfb2c2a12
z501a0cf0fa465ada84422d7e1720d13a1fe9d7353cb8262379cbb1dbe815691103f8bb62b540ad
zdbd477eea4ab3504a1ceff5605b7bbca0aa1c1323b06e1a6492b03e927b3f13aab505e91fa07e7
ze16f56aa769ff0912dee7daa01bfc5b8e2615ba68e9918c8ddc86ebd0c0b53569dade5fce71edb
zea866f6ff530b053f02c4f44d606f28b2cd21d8f6a70354753851df6cbee2af6dc513521a3c038
za9834f6da2ded014b7bdb88107919085d43109ace13e6cbf0b329645d590b1339334f26028e8dd
z3edd6dbcc812e6d346ee8bf92ef9d62ef0650fe5a8cf92662d0435338debe50ae01dadcfc1eedd
z86af9f9a9098b04fea87b293b72fa17561283f17bee33d4bdb51c4e22de8fbbc8485d923b35d9f
z17ae8f7eba788ff3fc624320e8a6419fecd51a970b455bca296480d5a991f572fd4128038a98a7
z658f25d7442103967106266095b1ee713777cb3dc7a6d13c3ea50c9b99c0df1c9dfd07a3e77f21
z8ce047b5cc107182ab283802f669229fb45e333f909296605c442c36c8107183a724ed20f4c879
z1860dc3c3809cad4f2d0534a44d8c040ea746fb3e4783590400fdd6a82eb7aa95a0b5c1e18c77e
z3aafb4e4939ebae7aa95ad3d6ebbfbbedb3315075b2fd730ed935ef756f4a615e8c9ca20cba9e1
zfeedf72dfd54e2e2a26419f81d8099f398ebbbf1e836fbbb29df6b176806f077ff2eaac3aac909
z5f34b07e57d405c584ab58d37916af76a9e9d7c46f5b4d0821605d0b1f23df5089a1b927f97d51
zbd58e20da38c7dfd1c35c2ff936d9e09a41a73e5762f60132ea50126663219e18f21c42a3547e9
zc3309a3117699b4d5452edf58ae952d0042a9e1800f876b804cf175a9bc6d3060dd998a587a91e
z733227ed6c9a57f95b600f5bd8313b3f69d4210b3c5b87d347522f71a1a7d6600e47ed28e313c7
zc8b17deba7db2ce0096408cc4c0301d18bd9d48a08dce347a4680ae4fa5d19e3cb832c92cf988d
ze5acee43fc7ae70a8247dd55c8499410235a50ed5c6585a6f1f06a4d06e751c8acdf327b083454
zf3266113e6220c33dc2e366a11a897b53e240311a13b0ac76b46e758ac12f8f795fc620ae0937e
zb8b03377ccb614c0d476632c4182919df9bd62b2a8a8169d19aec2a4f6473314da220ce785236c
zf68df2a9e84e69df6fbe20d7ea1609a6d9248f2887c941c20436c2ab73fe98dbd78c0f48da2aa1
z2d090aea00f43a31f7c75ad8637e1bf51981db0f40ac037686c7333bc13cc6bbca6685ac79c5c4
z03dba851c9bcc7004056d88024af2c099bc82e58aba9475f2385c0e3130c7b75904e113f736920
z5830c1dee7c21c9e1dd0421af37fdb12fb6bfd3a2b99e8b1e9ad42bcd99340bdf2efe43f2dd5db
z375bac77f933a97034151353472cdb5bb29e179d08000e2b5ed5728d41efd0dbd44233e43b32f1
z42d4928e13a4aae2ac603a993f6c64b81976a6abd75686d17d621091fff6a39f9b44ce8ef0f122
zb5308afe19ac4c3329e7f758cd3e60a26c414b7227e7c9270b0a2d64c0e21aa556bb58b3b06d45
zf5d0561b5068870ab5fe27d414be358760ad47926180243db968fe61c9c4cfbb426e873e5f62c9
z3ed4c3848222098bca50fee4426b5c14b54f8e3012dd61ae5c2f3b24763ffbfcf463ed3d217a4e
z9d62d4ca1b70ae4a7e0610382aed5a3076455d74b90ff49267d6b85d7ea1d781ff2142362a195c
z67d332430f5a24a137785e8cfec8a1ebb60eaf5325967868036f9badc6253d3892effbb469e5c2
z7627caf1933961abd98826667bf8545106446e7535cae5bf732767a0438a091b8836e5e1f153de
z83960e4a49a3011318e6c5b3ba8ef8a1320090443723c7f760e83e2a0c349ad5cd1003df1d75d6
z4ce4add781bf44ce5c3aff98a76d97069119fdcc8a0f9361605ed83a35221e3340501b159304c1
zb2429482e118044afa327e6a459dd1cc4ba0afc1d91c5ec21154706a7db92673dd7f5b8565693a
z105f6676fa1b16ff161d6ba9bac8fea4b7c3d0557261d5f6aab3a60e016cbd14d1f35d9e571ed2
z6b736f748e8bc235888d1828590e506966356e37c388dd810689d6ed2236f3b0685653a6992320
zf69355835f837736feaf5921b720c32f8f7880568e9517473c4d84a5f7023d6df084410fe41244
zc7169fbb455963e51d6fe4e30875d9cb32e3d1074d6df6f534342c6e66559c909d385d5714d291
z0312a588e3d5fb39dda6885bba7469aec0c2f6042dc27cf7188c15cc84bcd106f9146c36d2b2a5
zd02b064b5e8cea665d05a9456c3f08bae09c384f9044318aa0518b0384d0fb4cd8dfe5fd7a2256
zec2eda0fdfdd71e4ee23490cd8a8c7842a0e67eb590b8f9632c543493d839437a464022523200d
z9255c228ddaa6324aaeb98aee62100a358c1b8e6c37cac96d2d0f04ff966073b326af0727f7d99
z93d9d484d3c2109c03c1da04650ca6cff875bce98d3f0ef73f9dc06231def963f9b691ee0640c7
z144eb7e2791ac71be28ae4cfba3d080ea3c143f20baafd2e5fb292f212ded907656c87a58433af
zfb13cc6f023bcf5a454f59bbe12e1b2458a343bdd31bca0a60f0a742114bb88d08a0e88357201c
z1cd28173df4b637dc8d657297b645f226f305e252b66632c3cfdf266c3014d81665ddc7d104674
ze42ededcf0c09d8936524b759be4b0f48ff32b78895c8388a06593dab42056533e09b7287ce726
zd7c52c9de7cd5c15dc463418afbc6995ebaa0a7b1944172c1b75e4742809250374aa383199deca
zd2b26ff59d1c3abf497099b4124365c75614586e3f28681aac1c6a01f9cb903ff3d4a433d274f3
z38f4ca42ab86609c730908f31ac66036abf12d239aaec7b387bca4c47b4edbafc9fdadf2a72f84
z3284a1930bf21e78f0f6a6470a4ddb8cd57a9da69f32c491fbd0972f6fc22918eee30c53fcbf42
z352f34fbd1291f80d90741ed31ba77ab1d1aeb425e07e8e761a72be6589fb6a0a81993382a2029
zb619875a26054983fa457a5817c179b8a9c9b458242b2e27db60a33b25ec1ccad5ea679541e4a8
zdbf068f0ba461d6a5bc627a792ec3bb8be0dc8455a19457bc4128ee473980abe3c63e6b7cfce80
z2b3a8bcac4489629c44741b01d2b4b5841afda30d73dfdfd615c3722fcc0b1193b8400b3a05898
z6f63eef1c6c96fed0121b35e882d9c32516aa2d2ac4508d2becfdeaadd41d2a11b0abfd3cf6fa2
z80216d5a73907259de63786b518e1c98080286395ff93c821f30c0aa14af3485c110ccded95211
z77654137e3cb944d3b63dd5fdd7d463f211bfb858bf1e8a52f2ba52ac1303941676112e61581a8
z8420cbb916732a421d13bb717edda058042ddebdf26fbc38ac78b2bb5ac66c368322a5bceaf24f
z3763a9a75606aee14fd386d8bf38a31d66bc2e9dc23c53ff473cbad8acddd7c9d5272be89dda15
z85ab3923cd8dafd4c48da6704bb2bc347b30ea90fe91b01bb48f8f2cb2dd3e8c0173d1348ee4e1
z57b7b4731530a7f0bb976ff31f6ce3a63f9607af385ffe4ed0b741ace55bb1afa94153577861e8
z08476878e0ad19deba11c64ab4ec69638dc535c2833c7216073952a97c832bc07b8ac60842562a
z6c54392d8f8d16661ff8bae55a08e4d6738c571019d1ba56d8b21ed7de93a60d6fb7b4f929f938
zb54c13911f7ad2676e2b01a76e105e05b46133f759cc8db8907f761fc41b7dc369fa5c88aab9f5
z79f3ec9fb781ab5cb0e78cf3a806687842cd7684ec8ee6c57f49aca539cd8e0333f897a4d4e367
z3573fe5aed628ae9ce432d489c1624ddf9e7869e71117640ac1b07484f3bd5550ee6518694408e
z6dd115464a97cc1920f8d43241a268d715c73384176e8f328246d481e93df4074868281ac8a305
z5d50be6903ca0dd98902cca702d5c4288ed257b5ba5011b65065345f211f752b8f869c8087eedd
z21d477e78a7cc07ff4dff3320526bf1c1f44b2deb0a048987b04adbe18792f58884f35db96db85
z21bbb02533e4a7577ee34089837a786c9181c5bf20c279961a22ff149953abdff60f31d104354c
ze0b0516c4ee093fda0ba44835d411f77ded1e35187a8b157251ac1edc0258e8e414dd703f26994
zaa861aa01ec4e82bc56bf321cab59b30495165a8e09bea09edbda6d6d7329dc23257bc745ed7aa
z0d1bd90fda88e52de5af88a3da2827cd43a01395e0b9e68e78f1d31d6a069783abd944c0c2fd15
z99dc13edaff96b75cab15797fcc93b4953feb42cb222336551ce76301596646ea8000430e475c5
z53452181c1dee6c814576c9a20fa2b1f0407f71e4d256bd11fb0919f1788aa9f845ffa73160c5b
z7c3991a8475eac828e7f6a858fb6f279a589ddae51a359bce0d98c38a5b767c08f28e9f652429d
z22bf8109909292d85608a537b7bfdcf8bb58a684b768932655763cc3d43a7632ac6e0ae8e84fd8
z3663d38197b3748b1450fc6bc3eb2fbeffa464f2aff2c164d9cde07369094d37759058377f262b
z33eb55aa43105f26b2e7c1ce30c82cd211bae639ba653e6d9dacb523fcc77340d67103c0953c21
zcee3c68e8b81186f121038d426fd28d5d4ba0506134afdbe9e8352a1af62ec2a63ded2b4bc4fde
z01698291288fa76bc3004d26bd6ae64cefff504f349f603795fe6e8caa12d59fb78f55957d601b
z8a209b4c9cb493eeea061c8bbca7136efd8354d72d4f32304d1affabfaf3e053bc2c7bfcf6b25c
z1c63d11aaa7c097a24ccbd1ea55c21cc5f9579d314e12ef9d39fe96da31db96bff10fd7e65c3e5
z17f07eab1ebef250d7dbccfaed2dbed28de2b96a84847aff7c04ec94fdf8d162bf9880ee3986d8
z727f69a39c262edd6b8bc362fa8edb70269a211f3472208cb394f170ba328dd75c61a7239e0b30
z18fa52816ed9a7988968cfcd5505e028d1e3983c18ea76ecfcade9737ce0a39ddeb65784906386
zeebff559cede7fb7e6c7cd35ac58447ca0b565dd14405c3d75e69c063f42d4babaacab9cbfcc9e
zdda0a7880b007ac0a3babf115394b0358486c800796bd161ed2e841d878a1c72d109a26dee69e6
z20608b398093914063ad4920adc4dabe477cf0bb2a08f97fc5d3fc4d47d90132712c6fe4857c0d
zbe5ca719c8fb857f1b9b908fd6bf37fc9e8cfed8f6a1aa7c96e6bb94f9a1d9c7206a22731af6b6
z21580b122abf85ac96cd45d1769003e449b89524a48baf92478daed1931ae0f969774fcea9a4a6
z08646316be9c18197fbb0e65336b82859d55421d12e3db21b629c784cac6dc3fb1ee01d47d6374
z2054e1c3fd69a579892955523aa5acbac75bdeca88f55e67e4609d81e8044e959484d7f2c020da
z4391d6a47b96101d635cf5fe5b42f7254d9e2d2a61650ec855e1237b1936942d9c01dc210ac73b
zffd8c71ecee7aba24b9afda1f8529173fa834e4b607e0e5f8e479c9799f99b34579c1c2ce4275d
zfee2c0ee4bf18e3252f8b1d2de574fd6e3c4c0207cdad8728ff611881167a8b2c6c5fc62b69488
z89599b219cdc2872b70e329ac4e9be4ed3ef9e8894a8e83484da4f8cc187358c58fca148a38502
z8466a554417c02475f05ba5ba076ec6a03ccc44b43de3300d3e588a0c7c55d30be56eb264685b4
z41b81514ae5f53fa6d259a74a41c4dcebd0633bd351ef75ac949686114ba8fd315753568b517d9
zfb742caf78d74d8d5dec7774272a6c2ad22ed02912079bdeec9e473249a8034b99259195177c14
z2b7ea071de991adbfb7a9be48fe3c27880b43bdfa61a1405903b4eb4bc9aa7c677589f0a62c9d8
zedb38e3724d0a563ceb7019e9e8be030a0a34a132f6b3c416d5ca3d31bb583256ea7da63a3998f
z3fbcef8111d5b09e34a096dabe032eaa4d9faba0bd4d30e45292b26b03593cb017a1c9af85ec85
z59369571f74a515ad4a3902ebb3da5af1ab086263a18a28a53d2b1e0c50bd1d535767a2947cc5f
z6a61a52af8bb5f70a63240795f7704c2331f0bbc5d1a4a9432e50e112914e4425bc557e379f805
z2e07e09dbe4757054333c9a1fba7a51392e3b6ed9326d5779e1f9c78f8ad911cff85ff9d044ce0
z32595936205f2f511541b695eca9b076c5bc27ab6cffbef1696ca72566f1492359afdb7f22d9a9
z40e979853c7ac2dcc045d1146f570cabe17cc5ca60a56ee305c0f869ff9f8745be34895a241999
zdbd4558f8b3c344934354f4bc3f09dd71506bd8d052ae0676ac477ad5aa526f8d92dfe759d976f
ze2b5dc076fd08169bda2aff428b7483dabc7944bd9f869392372644d546cd936a01fdbc61c32ef
zef27bc955fe7f45951e3647dd8d54ff762c116abbc6378668c186db699ffb2523db8c88a4f8b4e
zf04729268109eff7d4f352518c202392127243d19156e448072034b232280b395cc46e3589f069
z863a3307b845039fd02579297e3749d6b97de0fbd08e8bde4e6f827217b160a69c8f961b4e12b9
z50406eabcad014d90e61daba1344c59f7fb8d7939aa5d15a1f5b5d21749023eccc6c39dad200f6
zdb5849611036ad531b48ec748e18b21adb9afb16045fcd4a148ac2d061b6694635c53590cce4d1
zdadb36181d3c9da8e3d1a48aafa513bdb55bd20e93d4d2ef4145cc0e7778317d13eccd1ee88263
z4ecf042db9f66b268b0209606a3ed7a996e432d968730c1923afc0b2e2e49374e4d9135b1fe44b
z715e929cda241c2fc317e10a2e8b0a759f8c10d74330c0518ed455d37deed8d9e6db0c16dc7fe4
z7f4a79639b4b4ef688d70d17f33a6ce201ef820b037ecef4abaafe2b1482b218473d3ae86fc94e
z0e6dd1f4e652958d0007e668c054d9edfce07223738125ccc58213198200116a90372c2e976bc4
z9833182cc088298d70e1d673d1d36959ed735e2de44ab8017ff758c05a8fcedb35d12c293a5234
z321128f59a4f6a421a3f4e515f1d44ae44519cf45ca71fa8383ec958c9b231f360cbddb64b8595
z86e479e2cfd2bb8559a4b63664507227843333e1a612f52f51e1a3ffe6d70b7d1ed814bf8b98bf
z56e92d8e22ab477c4f9e7b55a5dc72e1d9f3265446610adabba59b1f8c724873cd09f1548a0958
z7058b993e1cb0dda37173951f751625a8a8a7fea74b0b71e6fd68afc881cf08d82ad384a7c6567
z5e67da3a061fa28758b29831afa6646e03c687e33c5296d3c0ffd1002808dfd1219a3b6db2abe4
z3ba3418c7a2abc39bc7d6bd50891b324f5769a6c3b4077be01bbce6843a9266b2621f25c16d70b
zef8b4e1a27d1770591893bb865bd046f66ce1a0f3c2f0173b23f1dfdefc7987fddfa587d0f7d19
z8c86ffce1309ba24c1b0b3be15987d746f3493a5aa821ff6f36292f2c3032c4380c6376bc2d128
z367318f41bc167b66d3b2da9186d9c577107bb717862b108d8956717fcddaed4be2eb4d96bb544
zcbad8015197ed7f031cddfcb112327ea26c6cbf26d120f2db279ee138ffa79c688f6ecf78afd79
z40487e961bbd60eeb9cb5f72aa838ef3e4178dabb69314b4c141477d2411c4691ca13da69e83c0
z097c6d3cd87baf02ded494911ec2b48c52b51e816f2edc7d755978a0625be31a65aabb9f06c111
z589286fd4c43def1ca2e3350295b54aa1aba670db850d51315b3e6ec9c55828c8c399b0d0701b2
z2b6d94336d12f32c17d07699cdff0720263227c7f217f8fb76def6fba6b1421b83e3db4103d702
z30e5e374e903a35f48cd9da9fab89beb8633e9abd76d9c193546af98ca0925872c7e9a38496831
z80996870141ae95a343ce8416f53dc5af27f0b78ff760c7952886e4c74d4a15f9a7a20934ba89b
z786c3e3936927b4c36a8fec28068f84d89223d368af9ee4e618cb9cf99c7e63407a31fdfba90e5
z9f27a72d151d474dcc514131484715c909acdba98bc58f7f7a1f177342a086a672152c671960a3
z875d7e89722e3efc8cf4fa82d5117f48f4811995374a79ba064d579ff764ac7c627fc3bed183ba
z0cdd2cb7aa1805252dcfb47e6bb53ccff055a29e973b9a9706f420c27d0bdce6efcd69f44c1a40
z88399d643293bc5d5e5ea00e10e29aacdf2193c03c7e8a0a750f01dd37ba168b2c9218d151c5a9
zd8f6a3ba21200435b958ab6b53a746033bd5af42542b279db8dcc1c9a4424c9f71d4722568c054
z8b283a924465f59e01defb5121f0c87b46a2d94621ce43360e19812b7dec33c0f3c3b306eb100a
z4a0f32c8db75891b65577060aa7c68ecdadb311cb660ad68100d3cdea1ab7e8183096dd4c3142a
z0aa93d6544e609e81130e1939daef13dd6bd16b1e0df6f906292ce0bd33c7800d1365be80db85a
z570413d81bdedb7c9c2b46360acb9e9c4ff2ca9e77d937e9389958fc690294620fb412ccc5bf0c
zb88a4f2ce59c67115b46e1e35503ddecb00fe36c7679a0921974c1b79d5d5155247399dbbfdce9
z005cb2b4c8bb57122da75e2980ea01200fcb4214e43ac9dea5e5ff1d761366afad4032288092a1
zbae4405db01390c668d7c098964e53057277503707fa491d4d9493f6c279986ee2cc20610b9d69
z7696e538ce9abd35b8453fc16e95455acf2f7e3f90c4d1b744f3f00072fe517b3ef5b376e6fed7
z91a92a734ac9337ab8b233b0922353ea6d6fe9372b199076540d56289614d21d094a225896475e
zdbac32cedc4f058faf4b9adb192a03b46c22085a95926f5f5697e5edabcbbe15b411d422177a18
z273bb847820e935a9672c1f44cc66ec2d265d5cd9d9e07dc705c0a2c91e7de824dc10291931b5f
z3e95f0f66a706590c3643cccf5d1b5bea6f420720c85b45a578030c5bd8799c70efacdbbe83123
zd4c2292b93133ec0fb7647469a249ba9da380f9e39d0af880db6eb1b26b1f8d7f64d50464a4b7e
z49559235e27939dd645557260f7fb1d4b1b3f6d96b2fa56b5608eef0a2420e5d589676e9f86c03
z8c6e4a69a7e01441e0ffe46c7f616cc0dae6d02940bd043d97b3151282dc24a045597ee3bd89f0
z113a93c362568f0cc1b28a4ffa2d826d3df8542a518522add7f55a901241dd174e48a5a3521b4c
zdd56c448f1d13fbfcb641ea94d64cd05cce4e17ee0987d2bd3abb548a230d0ee2f601c72a540c4
z08f971f572f91f8a8b2758d64879e8967e0f86094c04f2245bc10a5e41731138960e519e512063
zbcd48ee9f5f9a49a1a692d48920692d5e0b60e0f280d9d4d9a3c0495b3e5461db1531b566199e8
zd16deb3a6456c2771625876d9b399d25dba6f01667a9dc837b3ae7e5db4fe2708141fefc445a12
z58d8d75d7ad98e3de0021f2dafde21828ee073a2e7715f3acc46cfa5de604277fe87985c6aee5a
ze2f3754137adc5f79c146fc27619e184d78ba06943a9c216ee47fc4eb5960ff45d93f8d709e594
z0a0561f23d4b5745f5c23b765cdc1c10c85d4794b5f93b8537ff2030806e58027df66fa73362ea
z6c6d48a538091301cc3331ea64b1255010014b77c95a9feea743a290a2cda0971fc09313e773ce
z9687889b363f292ce75db5c525cf899af3431e743fed76e9320454600c1b1afd1541137765c48b
z97e477dc0ac04f9edd5aee9f45d0aa8237db5ac5519995194ad08175e71b3e0e6a776c38c460f0
z59c541b00dccf9d886523af8875845582c8a1640a2c3cdc4c0c6106c40274626e28ed3edc58eaa
z8171ecc5d7adce20a4babb18f5312fbe0ddfa6fc1c09f53fa035124a3afba9820c54bc9d8bad8b
z42f9bca4d75280a26d7186b0f537c5fc52645bc0ad3838976294c7cb1142b35dfa97fe6a110af9
z35bf441918c6e48fd9aa8685e61473491748a5808b41fbb220c1f36a7865edd89667556f36f148
zf2c502c2abf15eec4adadc770606ba2378a8d494e4acf0e9a0c0f6a078382fd13e33e3ca4aba56
z8e04d67ccb64a6b649f321bd12ab235806d218cbd6a6e870d36cdd99a743048a977b055bce2a75
z1bdec34be842354a4502b7a090e8069c293370e3819357eb9e637f2056dd7ca0d760694161ae2a
z8696a9b741a478f6a2dc04cf60473b3292025ed8378cddd57007ae14778030f65e5495eb2beef6
zccbb9c3c0856fab65e4fee05f8e26c0f96221d34fe0d4be686bf634dbfdd052e26b41769f21d1b
z5e31b6db1db2b644bbe9d229c578e54faa7a38391440f7beed1a368455952b24f9465e691f47cd
z3d8b4390cc22203dd64009dbcf65d8840241eb3c8d7eb7d02330aa4164a08b364c30f93bf74358
zf8f1c993b475af7649578d6a7420825739ddf62f7c5a5df925b1a705c0b675c6d3c5ac7148abbc
z57ab53374f410e95e0ccd9a2c87e4355788b20ba3c8169a36c98aaec20979ab23621297a6172e9
z975c0e648b1e11a36e2f48d254ec071c895bbf2989c13cfc6b71ea004d917277e89f2d120b4894
zf095a8557007a0400e1ad819a7a07def9e63995d6f799c40bb93ff9ddcbe3d268719de781441f9
z6f900240515581eb28ed32b214f8773ac0124dedbca3d3277d141ff01137e6dc874f9931af9db5
z82681d2efad065ca3d80f693f7c65110690c0062169ce48c36e5e8cd0a80d2c1a6ba19114bbee1
z6693a08f30e77fcb7b7d3d77298de4576d2d67efebdea9f558c693c3cafa32f45f619287e7f466
ze844f54fa6ab37ca00dfa1a6cd8bb9ff852a85aaca0624ff517d30c896f1f7315ababc1dfec278
z4c1418a6cef74aebc9889e2de6f94e45e64165db41039739dd2481201a536b6bcb98de6716d0da
z682cb30f2750a40fd7ae57ae5a280e7b3f839d30b2f57a0816c59871d45735b1872dbf3d1fe98e
z627d365e3c50f72b865a1ed286e9f5d5657a3ddbf8abb51a54bcee9d0a631e698541ff461a2168
z3c3d6529766d657ec3821464933d0362a7d04bc724e2f2955d447c9d69b83319fad21af5132570
zac982bcf2a3812610222745a10fef077b2e039b9cf24a19e97403ba386b1dbf31191e2c12d091c
z19dcf4c72fccb116f96dd627e2bf493ceb4aa6bcbc5b2a0721a90f7af88d1c4d3232a5700458ee
zb117bf667c36594f149cd22e433b7367c1061ac0989b93ee17ebb83c65fdc1ff304d363625f9fc
z5d0cf16b5f172a8406024ffa9ea3995acda063a1957d690471cf0aeaa9b463abb1a35f26748acf
zdc7669b914a20e1281d713e7200cd1ad81dc987dcebae9558833a838c386e8b4d7b373e5d4bb74
z8603c16dd9f12acf1a71b095ca43afb27e073e3a129b8311cd29ef5ae59135cfdf74846b2f18f3
zbc35ccf30744984383ea4d7a448032c56ac4b165965ec683e9ca718350dabac09224e26faf97b1
z05703dd6f4606b11e51b1cb50370c69f6b0ece13f3ec2d140f71125d2c9c798c5fffb1a13eecbb
z8b55724a0872787c794c21ae091fb54f12de3abe9ad0a363dd08700f6255c831a40721e4777a06
zfd956e64b1153749b68b2ab40ad3c1e526b9550ca1b9df3081b07210b12362dfe891d259eab2fb
zef464aba9d0bd16cf2af1e2e9e25b73db74920618ed4c7716cbe1505e08f0c4b6e3fe1149e4347
z42fd8ebc70cd3040abc8a729027eb0247c15343bfcdc7acaa76cb2b002becf5464b8f22e072e2b
z9801b2c801942d845e20021fda2ea914fa89963d7fbf1791c24ba9c907f3154cea4d06647ef0a8
zf17c6315f0562b03076d991055ce2775b65b27290ed6fc39f86a768b87b236a781eef41599893c
zae6295a3b063f07b38caabe40b1f0e0a61be6b7404c8d07a76a778fa621a36500f3bca1ff3ecbc
z5282eaad987aa71e209465d635c637c9ea2cb934d54df9b4bc169815c700e43d1e6a3fb77e934c
zb87f24aec0f958ab4fd37e7c6ae05745c7a1100ba9240b2f32b848acfd10183fa481e5572b6924
z4e4e6e2125acc991c98ce077554e6effb27ee22ea2cfd2ebed792c751d6d3fbbe8d736e53b3f3a
z3b27fe3d90e23824e0ecb1cd603bae64e5119c8f511d40f8bbf65e9519ae95f166437bae70e015
z3fe5e8f6e1245fa58741d725fcdb9f219941a11711248b2d6108f2a0018b5024087bdc889e2c04
zdc878d67f8ecc1a2a7cf04884d8e07cad1ba695d031314b9738559978df98e6b96ad1cbc84029a
z7854bec61f872d4a4c44ae58307ac33463b8b5687f437a02652dc99711319322779d8b6863215e
z2ee0703eb20162443334b9309e338bb38a63b3eeefa70fee5276935f6e2a377e95a811c5c0b1ed
z34abdfdb09792798da3a8d5c3ea3a9f2128b94b2cd83b8abd2f1395167bbdb0653e41305d35f3a
z027c28410c94a085faf4880ad9c6bd262f34b7cb4e746768d7f1f200f79480118cbc38aa7ad39d
z8e55486aea37f294f211ec2fb5657751627fd9a91c26bc78063f6493a5fab3c99d7e9dd4bd8cc1
z6e77f53f06e53454a890c42da2fa0a1073c3fe522d2769b9e343dad3e82b46587e03db5b99073c
zbe210a58e4a3b04336d30f863736408c3addd76c682ae07dc183dd4858bbe57fd48da7bf3129de
ze98d145fe4b3a175ca9f7649c7b529105927c186e62f24ffb4b98896b81e236d523f25c09a6d6f
z1f17227e8c2d9c51f134f5978c528cac0ed5548b0ca4684639e0a831b23464cd4ed96a89b307ad
z967645bb50b04c71a9b87cc29e8fb2cb2337ccded5ae887453c6ab804c2b11630f8ad3a03d0627
z41fc369a0c6094d925e08b8f65cc6aa0dee33b2b7b58db10ddea5df2c2f2d87a6ba0b1914e8a8c
z30e89b21c053e881302a197a39887396283289e8129e1fa9be928d91f85e8e86a62cc079eda3dc
z0811555545866e9a2adfc6132ac5106cfa57f43ad2b973df3ff5d593ab9ad8ae1d553eb1cd9b8f
ze1aad315f468a5ad88594c171b8c917fa79e6f89fef8e57f50da017c4c252aef4e3c7f49e0ddeb
zc3502de584bcc8edb9a39f0a8ab6e55fe770d8a93f6801416c7ab9d689ea669720cfbebd5868b5
zcedfce07b3aa5e176040dfbff2732b1cf7609323bbef598eee8fc5bd6e95e3462061145b270d76
zb0a841dfec8539840b2182149ce1e2b1ddf6e77b0eeb2621ee3c0a6e4da24da46fe9dc71c8763a
z93b6bc4074500d3258b9e1ac0a793535a6ddfc498afd9e73c8364fbd18d6be22650f7cb225c06e
zd71e00cab488a503bcc5d4c5a70c0ed3d582ad6e1117a913e538abe76f5ff6e80e54afcb66d552
z1e17097fca5e0feac05483b7435fecd8790a08023fc14b5d3c996f941f58270964306f2f2a498a
z338aa722e666696197e1c47e49dafb0577ce88dbf6f5591783c3fe86e00aa5fa6dc865d2cb1907
ze153a1f1ecba1ad56d8a922b8692dff8bddb2b8397ad5bdb6cadf621f828aa4b0b0c0069f8f99c
zebd7535c87de4ec88ecb95f1af9ac8b5e4f009fea413f88829d203b541a5efbefcb0d8e4a7292b
z6be3e1c6176eb39ba98f9644b363dbe07da88a60537dc98e6879478e333a8cfb481825752c62f6
z02a62911e13baea5613accc3f2c51132ce7272a67b246745998b4f8ee85522f9d33843f81b89d6
zc7b889d893144578061d175fe50ea207c9a28a495b9cc5d23d7c168fb0d890500bb84c5dc8c5b9
z86ba65c86a6b4e5fee13379b96113e51c9add820a7bffa7f86d7720da859067cf6d9366ad47328
z3df15982791346143bc0bc91d41ac031a5fec386ed12d9c07d70a04233584902a145edf8369af6
z7247e0af6f59361939f51a5c966d5d8921e51bbc13b9f354d6b3d922a226770b754ccaa3ef2971
z92a50dde6bfe34f53755c2cf80a2d82cea82da7053e0ed8f4a49fde8f79c884f5b8bb4af405a4d
zd7f5eb02695e63e35fb88c8e09a556e8ee7c66979c0f39fe6278273b33c916a31e12fa7443736a
zfc336bdc8179036f24f6b28dc364454c351bd98fa593104c1ad65b117fce11fd6ede58c12c3585
z679510ebd76b94b002d5109e215ec4621ca7941fd2bc53c17e3caca1ab2ecc618cba29ae168898
za1a316ca141fdacbfbaccfff8b16ca688ad43e01c4581e1371d4bf313d6ffc5a37ededb5717462
z1774ab6f63a3a2ca2f4da3da144aafe5a8de024e60e7f21c001f51db4991163ad20155442d05d1
zd3a5712734c85bd461b9d37c7f1fe68387100afa875d0b9529033ee7c1a80d0314b15317edbf23
zfefca957477788b7c0a8382ef55abcc1480ae40c4f411ff44903fc81e9d016a27832d8bc12b9dd
z958ffb382d08612ee0c12df3aee102885e648b690b8c8a91486935f0f80c646f323fd76bcca892
z70c27947bbf846ab0913483782fb29a8629a8b55f3404df8abef38ff15b1a526e458c7006e1d74
z8b67546035119a04c875a3f9783db44cd660bd169e1c00b06c544c9a8f8cc2aa6efe376a251622
z40882d420d02aa47c18cc2910f792c7b6a6e99e92fd5d9904d44b5e8323fb57aa7077513430a67
zfdf2cd1375d67dc8275b008045e0c6f9b1048e5a0e04c1fa170fd49334b5b1165dc64a95c31013
zb203a8d40393da86f292f598f0593b8f82b862135c32884f672562d9c41f1747791be48ed667c5
z968237119af3fb7dac734f24dda5133feaffad8b3f572828397ce55d8395a6b6727044c0bb1539
z721cea9a28f9bde11b9cbd245f5b8643876535ca62563ce92232efd71e86b000b93dd3e0990575
z94d6644f7926bad8e47348924e1b273a99f7e2f9f50c508e6263db972b50401f013c6ea7a091e0
zc739c50434c14db858fd3df763990b6a10f009c84b72a10832d9fbad680a3554475bfe6bdbb9ee
ze2f652bb7e3e671c3dcb69db789a253284ba4ef55e918e97a98edb9be205e3d91890a775f29443
zbd474018f8a00bd51a1164ff0135f86cc8499037d698c5c68b5a4ede0c1042e1effa69227824a3
zbd04cfd074c56b27e646d403e8d134cc883ca003cfd61e7f71d3137b3e250b0709930d4a1a4416
z871475cbe4218c19249b57761896a8b84a2a7bedd718be8e6d2acda98be4b83ad6fea87935ea00
z2685ca4f5f63d67bfdbb375d1e501c86c30541b84b3ea4d74a692da10ffcd8b54ad50c6ba0da44
z7d440a16c610e2f2be1d55a7e20c6f8a677d85e1376a589f902a4593703dc4215ddc350955d088
zcd0161b4da2b4291cd0f6001d69b058c6a989f3a72618852aee14119d130f303527f40806dd20a
z8955d8a4434964f0039862201d3b13ecb0872ff9f4f10639b1e1174d8bad8055075ccb3ec7f640
zd5b081b54d64a7622d3f64977811e8b1e9123a7cfc7a5d0dae3d3161180d94f273530c7ffb56aa
z74584da378102747a95b9b70ac562441c3e8b374e3377e192ba2665d63ee2e1ceecbf7af07b201
zd799e633fe9e15f5c24475998eb4c5cb114c7cec94805484c4587c3e26c338b1aa22da67684f9b
z413082ad2af21bb79be3b895ebb9c3dbd42dcd551b2b8339cf450c1fe1466c26ac422334030207
zd4588e96af0967a27c72cca59588321f73837ff9edf91a4eb0dcf637b7462d9a97b94119fcf275
z4d6f8e29800ab60edc568720865a9b01b135800b0c55a347a960bc936cf8038a8159fcdc2838bf
z497077ab5b0174a7243761cb8485afe85a2ecc684aaf9caafe97fc0fd775596262c9497ef8a425
zbc0486f350a455ea8a3e50e8a1f51b9f9066c6761c9caf128959049f821a76997d5c3b7f47a659
z964997c275907f1d2122d815c2adf37cc24f0ba676aa1bfdd229279bd53c7f60dea4d6a9ab28ed
ze72fb99e284ecdb3d131aa74d94ee2a6f7438c755a1d7b1571f9a7aae734e2962da3b2de74217b
z02f6f364cc137615d163881da53ea7406ca98f70a28dd7024cbc04a05629cb8f6b2b79d529deee
zc3ae3e1157387119dae7b6c27f6d42fb199057c5d2ba114c9353eed2f22e918f4368dd4cb11f30
z9ae3706ca658d3283c1307af93014bc20279ac8021528fb9932b8b68ff6f087f7cd4196c5bf174
z9953a3a1e47c43422e982435ccbbf31c4b6fc9ec1aca0ed72a6c2a2ee56509f483ebc1988f171b
z2936a97af757471f3261f03de226635a00041b8285ce95a6881f40bb155dc0c2b26c9bd23b430e
ze093b55272d43e3d5b3af1c6436ec4f4a2bd4a03ef9a8094a01c7e4d5038e35b4e893d20235a0a
za0eeb9e478ed20f6b08c88f625e9380d7f84bb792b5f2ebb10c502bdbb66b305b30e24ab37dd3b
z3f9c1f8d34cad3375eb27242f8a2a575c244042755ce12ae0f9ceec592cc184386e593e66a93df
zb5b2499bdd08dda7fe8b2f9acca55b7829b5f667a1d83163bec06cc852db13d7d32cd58d8ca7e4
z20e80f13712c037fbfeca0ca00c4b83c29bbe3a3ce9090cceba871c41b8a2b49ae2e41758c5024
z436bb824d5f8d2fe0a3e4a71e7af9eb9f68d96fb80ef2e74198fe9e158fc3a97d76ba549d204e8
z5b6c18cd2a8e732b3f54e29e0404be163ea399835a7fd9b9d8d6de66a687e01226b5fb3ecb84ab
z0da104e01ae39f9c5808973ca60b74ab49009749c3c3984dd2bee9d7deeef256998f77faa31b6d
z20c719d08127a8eae5da43b1e429b96202dc797e8ebfe8475815eb43903e5ee50bc0e1843d37ba
zf93578b0ceb79d572d2aeb61204210b3b7552d4825a5583c6f41989110eed6b1797dae3f5b79c4
z847ebd296855142c1454bcd495f1e4fbbf24d5ca77eed57284a8c284a5cdb0585b8c970582a45a
zbc189dd9e22d471d9323b8b05d249953b72dded4146e227c4b01255850fc6f02a8306f1c25b49a
z58d6d249766fe266c6e8ded3241ce0293e2518dd20305a711e8a2baae0ce9e23ea1ac29473394b
zce5df2ac928c904ba8fc73aa6edc2571448107bccf48802fc0d89dede03a03e08b4a62ec9fde27
z5d4c3be91618428f711801e98a2300bb3b7b3c81045c8fa977742926302f051a0e71599aa3f7ef
z489640d8507800650c5086fbc384039d4aee682c453731f677547f09bee4db92a05eb93238d3fc
zb48242282abc03987b2639b041e27424391de65260e9e7578f02b7897b40ee1a87f8094e99ab06
z3a78c1f98f95770afb0e1d9ec674be7310605d189bb88262b0726e899bd33d45b0ee77c4e658b3
z389ac609b0d8179612565ddd2fd9e57720e45097b0658d5ac7c5c3c38131ba87a0064770a104c3
z4ed1b38413eb9b9dfe5a778f1918bcc34cba59f76e612bbe10309ca10fd8d721624abad9d8b394
z7d52309eed998a1c8ddcd9af6a25f7701790373ba8ae90adc1c0e79b21884b2753a8e2b97b3339
zaa82b099815783fcbb802782955436bdb2890da4628c20bde1c23f8a151ef50cd4e0a4204fd5ec
zf179918e6a260076b741fc90c5038810d26bad3389e11e70cca3575fb090bc87a68e5fdc74b7f2
zebbf8473e831c71daf64a94225daef860ec297e9990c31f7f0cca83b00ad6a39665e97e7c90741
z98c60a07348f0493be11e2b16cd2ef51fef4ee40cd899cd5f1b68b0fa3fe96eeb2538e4e4a5a06
z7cfc6ee507e4a4865b51cdd59b63175beb5f1e8e0346c3b4dd4b1267e27b80160ba215845a04ac
za2e218aecd33ab93d6939f677be226572f8fcab25dc6e35a61d5a63303a43ea2f62a808d698560
z7f6668a93279361b27ef25a79ec19b1d5fdff1444eb95a5957fa3ba12593ccda17c5ad3d1b9d9e
z4d14798f7a70bb781473eec08d14ee2ee9a07b25bf396cddfd05382eaf04fa694f18530f8aeb37
z3eb3e07794228362ae4d0b9b0e530be8301b01e9236150a7fc055737ed6946136162fd339a7064
z414bdf8601fbde371c2d4682f3abfcf12a2c213b50126e0e2fcd4e95d0f1173ea71d07898a751e
z8c349ad6666a9d86e2468833f1f9dfa4b2712c7371276bbf5dc6ef03f345e6f77fe60fe9794ee3
z491a5a8be8f0da31f00ca7cd2ff321f6d85689599abbb31710cccfcae5f3be26bb1515aaf882d9
z9effbbb56180d2c7fbb30c9f8a218648a73aa576503a1d018f5ca836275cfeaef539978293fc1b
za4ead22f67885ee7796d550a6fa8fd20d6a01fa2aa7dd97b4521335762100b1f7e65a6fc0c3203
z0d3d3d931b2ca0e97e1ebae78eb9fce7e4f6c855df62e2b3297d0a396c79a73001d476af3ca666
z65d65bb27bda7707e8b9d391b2cfd38263c0453611875dcecdc9f19fee68b5f3879a9bba2685a6
zdc3d90b0a4ef3d56f391879c81765b82439c4f9a650e209e873e594a8ff2bd35efc5790767b4bf
z4950186cecfcff8b762285d926de48b29be93b6c0b3e7cbaa5c2558c7525cc11abc9c6725c6d6b
z3eb26631ddd18efe6985d7a17b1827a25fa352f119e163795634cbefdd5e5b799d3e3b7de5c4ab
zdf8fb1e16c13f9b60ffa70313376e5c2b07dcde489eae9c0606c2176e99a7914a41c0c80639061
z24ff9a17ebb2e8f3cfe9db827094f2e2798f2eee063f1174632f59c7e54bbf1f650f0e30de9593
z8f733f1d7ff7e04b93e2aee7ad1e569491a5680c0669239bb5c029bf0531c59c69e5001c438deb
zeba6d1af3fa5f418ec082a275bc87fcb94acc3db8549b91fedbbbda8bb31ef8239e5508c10e3d8
zc387576b3b0cf017e9d2a91ae4e23af39a5c78d7f33ed2e7283a80c08a9d221c9a82f9f6c46da7
zf2cd715ac240da4e677ca32552ee98f414632a86d95604de90cb62f9a78e2f6af955580ba6cf90
zcdcf6e7d0dd4924c65230560beff94d33214c7ca50703a4916fa0fcb3d73a1fdafbd600d5048d7
z31ecdc816eb9feff953fb0cfbe0ae9d30556dc18a9c8a1b7f9c483bf336ff5293e40e0872292a0
zecf58cc2eeca6a8054cd6f15d41d344b491976779f98d6ca50ae1fcd1a6196e5b14e5a042cfaa2
z0ec168a5a1fc44b4f25e8807ae28b199b97af17eb4eb65ccb6112751de80481d1992266c04ebb2
zf9071c5577f1363bfcdc99c9f797c35fc559f1ed5098c92ed7b9a00cc04fbd273e054d380206c5
ze9c69d379473458830b5a7c3cb0023af60530cd846bef07dde2fcec9f0786f16a973d6a61c9679
zf8373c1b6e46d6c16e5bba58160a42ad1747c442a75f5b8f885efa241d4335a53127280f1d59c6
z1e0460cb740c59eeab5878d90c5a33471ed898f9776ff09aca69d5de6a8f06bdea17755e2a41fa
zc52960e764813d884ed4bf1f6b202728b8ee423d6d7e02d468ec83c99b3e464cae8ff9cb1a0ddd
z183a275cfae577cf9a052b6c438f1855115a7b1127c020a5d740155d27425e730f9358e916e2bf
z2c1d197ae37cac1d0b9a34ba5d6e121fd9bc8a036d368bdffaacef504544aea8dc67d69c9d5351
z0d3d7a4ce099e0a17c19323737c20a4e4eed4cb8ee7a4a16725c1ee73c47191f92fbd529a530e5
zaebe7b981e912b72619a4632ac84b0c0c6bbf10dc6d19c01a5396859b21a68b029085568358b33
z07b43ae9926ca9c8aafa5a2501d5e9c750ee9af3b64ee9c256090546f72464d17714a06a07746a
z50a8035f08066f39ebec867798a95a8607204d530ff785f853015cdac4ef620159f35c827dc5aa
z8353a868fb692085b601d0eccfac4164e19bab86b98a85989dad8899c0fbc3085ae324b9dc2f7b
zf0a66f1aa9b5dd134d528dc81ebaee9f63b84f1841154ad00157b2fce77a4eda00b81d2267bb21
zf6cb25c1c20281a18566c2d3a15e5b275af7eb6e51e48454883a6e1c95e98be6db4a84a24ebaa2
z816a77baad8b04ac6488c1342ce6731ab2d21cff601353e015ab9342f7f2590fec9ee5a399ae96
z5fcfca16de41b71881c92064cf5b345f97792697d6767a579d69086550499bb77fe1c3e6c8a3d7
z7cbeae947caad0b5cc96122c4d67edbd019014b25e62e1fd42aea74c7f5f94ff94916d9da03a46
z825f602c67d6af0a362a70601bcf19711b057c42ae281cc2bc24114bb2410e4f563dbf35756636
zd6f37d642e4d66954d8d66f61e18e7cd336d076adc065af722c0cb14cf5d5786f5de106f5a8ef8
zd9eefdeafd0b8d79f39731d882f666a1624ffd38e5811b1f82f5878375b25e193a0c9efb45adaa
zea5076c0b8a12c24cb17ba1ae7f2ee6c38d5c9f1cbd9ff8603fa02b841c97a7cb6de656afa96e5
z21f9ea07b7dbef23b003ea8c8290d951aa4fd16357228f975ce28e3461faa508b3599d5611c159
z3a7a5505fad64f95eecea6673e2b65553863b9961ee1a2bd111b4106bbef5a912ac41f2e6f5902
zd28fe5c589578c7a49b3d79379f163a2075c1a722f994d6a2460e55622bc9f7b0eebdf34ef1e80
z159d841600ce6abc4648d0f5242f942c44b589b77ca96b2fb5e7ea5b8cf8a08bae9d0c61850379
z28048410287bba99d1dfa30d5a3d1cbf0fd90bcdab06501d46e40df2e2ee52e8b3a05a3afdb882
z310cb1e8d85c97a5485b4631417ee31dbdf1fb844d3bd66d621678d10f687b697c1ca129a53615
zb760d1fed6195c11b5a90faa52366cc5b0dff4433b74314f67c09600133790dc893cb8538de31e
z13b1679c5537392ff8f7e06a35b2335ad585bb19b5344fcf7e800673de8e35d443ae435f6a34ab
z3de14e3242021a9d82ef9ffe3d44b5812fd084fef5083d588f9b77d0a402ec25dcb03fecd24f72
zc086e486d9cfbf969d7eee692e178c57b6a33ffef9dbe90603464027625297ba72bc3a8c657ddd
zd38b026b7cc2f686a650e74298cf674c58c8b048847e539a6e836feb3f6cc9c0f54f2cf8f44e7d
z91f3dea1d261197093951056cfe64ac60031bd74c82e05b60911f1e5651c92abd335fedfa53911
z378cb9e2cdaf83d68a8bb3db4bc5314f2d5511810813c472e91e73398ed93956e5745709bbd925
ze9984d73a5d2c661ff9b9d22f69a40d4be64702571d85d0398c8ac29039874d9bd94b1420b62c8
zd1fb2a1585a3b8118f6746c352cfc18bde19a8e1a0eea2451fdfd09bd71c78f8ff5871b56fc524
zdcca22850e9560a698af149601686f2de21f417db54749a5d90a0ec23594aef7c446dcfae23a86
zeaafa6388b77ac746b524d420e7dac9f66736aaf431b035e9e4405d65b626d99fc0e1b9fbd4dd1
zf18437444f64acdc04e200571ad44e3f45da68cf9988bcffba220cd71fd124fc864d8718fe5807
z4a718ec39a501258fec2e8715d6e794fbacb1f26729b35347390e462ffc6f1ff61e8f845dec7b4
z6c5ec9a966941021df86b6530accf53921199578bcbe1fe9c87cac9a1635cb40073d3847919190
z429ac61177a1e755576b095a99b1038636dd95e7c2736c7e983ca740e93c4895cc8d0b3b515997
z33949fa5d5b8a35b9937e8580b7cdffee445672df2f8dc7bc94b58c934ed9068d891c16329f789
zd00df78492672b4b95284a2af3b4fc0f9e6647749c352ff0fa31f026d0f7e42b88ea8495d1b80e
zac2e68fe4848cba4b80f0f7cccc88fea0ed328f726b14fd1823405f4f6076ac79e4c05b1f4403d
z358ea576e3adfa065d8eb429b04672950ba85072d343ae1f587361616b5b68ba349d10a4fe576a
z4820bf13ea0c5c34934417ced59c067c3498395df8451f2b260b32e119d121556f8dc02fdf1f26
z598150541feb63e9990db6b4d40e7e349ce14e95223d54bba11a44c2020f17a76f19b159ea8e54
z4b2c50f8175b9d10e969e6b2385573566a578ccb96fbb2e9fa05af6b9d8716687b9aabd9c51e37
zc90f96e8044af772244e131e331ada68ae61d1602e3d5999d83e6fc111736fbc99ff0d8b46de58
zfaf9d2c809a2395b533d284e23120b61816a1a0324b258bf232ff4afadfcb95e46e964dedc66c9
zf62afb46606d17d250ece43ba000ab53fa5f227ebb819c7f33302a67eb45f0dabe7963106a99c3
zcb8dd86863458bf827adc1138cb643381bb831dcc66e86c3ae368b68cf9979baed85a51b2a36b5
z6ac69cc44819c7c63c2405a0f490f8b2857caf757d816df7049de7766b58803ae6589d99a71ac5
ze119663c6f09a377c54615cd37ffa19e558b51626ced3907d64b6157117fc34409d39cb3c12a23
z42db5741b03ceabbdab787c92c8e17c51dc0197de6bf2b1e9ea61c980456f92b89f83a3cdd84b0
z9dae0881b57365d43bc4c2a732d577f2aaf3252ddad22ab620daac7904a48465226beeec656b42
z84ebff3d53074edfd16bdede79357dd7cdf577c638b10942efeb79d86ef3c87d717e962609de5e
z7ee369a4df4eb756467b042c84bef48519a20f18d64edf5739c17322382dbba2cca81413376aec
z884df2ab11328dc6650d2841cd97e1de441b6e2f04235c8a80ca7cae2f0f9c3e50d32accdbf472
zf100b708b04ffa7b7c157bf5b4300289550f7d16c3bd06b12d008cbccfacb58f2f963c10c4ad9b
z6d3b96d47b899a436eb2f50dee48f81fb583e37ba38fb00e316e3f3ba3ee2584c8c047fc3a48f3
zac342f28d749f4b1068db0151252be5298fedbb6996bfbb04e040a2eaca1327de9a682728340b6
z5debe10f4c146520be43f6a290d2985de00eeb39f5cbc5998a36d48786893851214fc717b10645
z6f28721ba31cca372c52d584f6405850e0fb9343d16c8c0b382e3557459532d48f4f8f13fa7606
za30b107e40cc6583939c856cd8e2b77b0121287a13a65369d7a32d79e82904922d3d00d18d3f00
zdf35fd0ef8351350d00d368299051368dd2d41e52913c5093f06b52829b375ffbd95788c997aad
zf8d2a82acc0758b37635f79ead4366f4fdf7788b443b0c7cf4c43cd5531f83d8ebb3463a93ceb1
zcc3af0e7d8f2c38f9923ea40684d184b6652e5a27f02e1b7f2d16c4c2dd4d595f0a953c88b7cb5
z8e44caa7889673c8d1b78cad9286cac9d34f01e6e074037e9ab58d37a020c718d521111a425316
z77d410d2f9cc92b84ab9c32c0ef8eea211b9a93b84f31039281f39954024d17de5f148a4a5bcd0
z06fb071729204926fb676b7d7de176bee44f71c3649a4f4cf24a588b7c64af3028765c6332c131
zf65d8a31cb2664bd38f837f0bd7b902975846093f4edba648e54216a4da22b68424af3e4da384d
zf35ec04c63f0c92788734861e130be7a56df85cddf1930726942b5cb3211b4de4d15e36b2f4632
z31a02b282832cd8627e0bf3ff95d68fa8fbcc5dc7d64a124702ce715e7b2c70fd7bd60e2939f2a
zb299dfdd14677ea6da711dfd6388d6a373f0932e7c578c96c37aee892731d2aaeed54c2169f335
z665ca38af9eb9924e39cbb445ac141c03c282c034ed4ff5bc26dfa42ad3a4f7d8ac32ee9c90045
z1f96b3a62d9cf5217118a2162e41114942a003a2bfb342c0a017875338f97946ea474da05fadac
zadc6b2d7351da48d9abca752ef6de5d9fbf8b487ee377d95319d25627130515a49b5732a6cc250
z9ce6a4dcb6e1b3fb4101fa4796d566c4392ebd85e82ff3213c7a5e7505de402029c329c5aedd09
zfa7b5b04f8f818b4758167f7aebea211421e52cfbc754eb3b8420560bb7d8a33169c140113d3b4
zacae1d53f80dfa80fed616c60780009aa859bf64030cb5878aa380366577083ca2c27cee282871
ze44f06e441726b44c2712bd3cbebe23fa0e42f588ae6a256c5266a2300c25705b8d4aaeb7df70c
z730589aba5839ed62f73cfd2c4e05779cc9ac5b6f0eab04c8bbfbeec642764fe56f77cb378a566
zafae2e911f6a099028fb8a1efec1036acc64e6f12ed6331acd0ccbb562f950e78732bd124b70c5
zfc0489eb1b94e6d7e177d8c891cecfd23c68dc215554b3a8c944fab79e8ff461b0f30cc669b0b8
zff849aa287dbb2856a2541c466ffa40c11173a8870e444acfccfae3b1ea3eac0773e79e0181ad3
zf037a5b2c076c58550c22f503e4b48716e688f81e366f8612abe2e0dfbca713a989336a2486d54
z363132802ecf789c0febf46fc3def732ec18f08c1dc40a46cedd480b2020cf99674f8d13a13c9d
ze3f4ae64491fc1c72339d9bbc63f755bccb0b1a08da31c77d83ddef046af3caaaffeb2dcded2d0
z6249e22a96d278a544b6af862a0f71f0970bce1410221611fece79da0387eca6d228eec515528d
z813054d139a85e1853df564d33302e47d0b7546fd9955c4b45b329d6f84d535293ea5ff67d55ec
zab0fa461fc24796884732602b68cdfe64e1f891bc3cc6be90f0240e73eefd824ca22eb258ab229
z45775046682dd745753e3e2ac96dc892b799bab176a54b7048aaaa1071a84b3579a08faebdd88b
z17429696584b0275a4dc27e93718909d2178f4816995f4c63353c317907a2cc1bfb23ef2feb57a
z8b15a599cb7065de95405963a80434d3102c119cde43535648d07423000599b4fec3fcf4f07288
z04adb214e7b2f2565e3328288482db058308a5267706e556c43e81375152fd79e8ecc8d5e0ab20
zd755ef3a1e61cae9db105ada292113fc13c7e33c6ebee61f886207875038caf5bf3e417b503b6d
za9907786e7342a4908f581bc2f822b35a32938569326d2ec584927c483743729eddac6608ee745
z2d8e3c85b59f064a9236905326e9847eb3fd1c1371be26f5db5132ffdae57fd1908e072ee093c1
zffec5e359c0e7da2d8b2660c8baec05c2cf66cf8fc06a03744397063e7af7e7ee73d309c578b65
zffd51fafc89c1159887dab320dbb65e23df5eb819223e196dec1c1de6a025420da3f5fb755e9af
z6d6204ef02fcc23fadc0b8a433dfd6747db654aa65e4c66438ade19a438c1d13cb9755e72ec5ee
z73f5c560df9ba7af3775e1674514dacd332ed2001075b689277a20efd451d4173eba717e555560
z94a83c6ef92b0bc3c58d12b4c6d70d7a6efc7cce71dfb91be64f1d717837100aa667417ced1417
z1882aec22de098ff2f5eb9e6910f83b3ad09f96ba4db98d64500a7e6164f54ad8e97834a686c9b
z4a7cb2af41a8838b85a3202bf90c392cffd3feba3be38a9045dfe8d1150ba119db0a304f5ba125
z0008736c2f448668a8de0a9bd7fd63b9b823a632120dae6245f929bc15c01824f63204bb803037
z1405b8de78c2000452b07d763d8b96c7431f5a3383b2e598f96c734ed389c53d5e13a4a32b272e
zcc62a72f10ef5ea5803311623e8060a9d29465a8381eef559d14645f76c1693adbd648dfa21a59
z0bfdc453cb3c00040b96aa4a2f8697c220815d13b36bccfb7580ce071d1bee38f258685f168759
z7e4b192f04c693ccedafda8a20be1d2aa642df6deb5c920757047e54185b293f218177d59d300a
zef891cf09bd92c8190e69dcec7e1ed0c6fc1863c3579497b2b385b6390dd16167f82fa61f55377
z69dc6e28ac48fdabd3f4461e35dd08b8e0990deb76d188508d70a7182f2b3212af77e69bc4596e
z9532ffbf932d8185f4770ed91d4b84b08d5992d6d46445a4b8298c98c571c8bfb6d7c69cf5e9e9
zcd098ed216bdfdb095764aa4fc1d4430b4567e694bc86e49abd899cc2129c2208a2394cec6c0ce
z0111f81d679b61ac63ac0e919c44c4d8cb8b7d0a038cfc0f0d6003cf2efc079d4c13a24b987ef4
zbf87522d1ddf42f6f6a340cec160a3af7f282237d774b9a941232a95f386aa395f74cee68f8c89
zd82a34c13f4364cd3fdd589e41b101885fd8d4ff0ab3b200603f7143cfaa7aba0a12e480e91fd2
z9abb810bb5ceeef4b38a4a8d23fcacf641c9fff30f274848facb39262777de1589393af2a14d11
zf4c8b6e3aca332b1d3caab1b96645d3c411ea56fff8b09686a1128cc63e37038de88e63cb32cd4
z0c4962345ae453a3dc12b25691a08bd168a17601b9309c2b95627bce053957e39e87d452fc1f66
zd7a4f65196415e72e7a40f88de4ff2d1c20807fe59076a8817dee9319cbf212b3ccc8be14dfd98
ze9c87a0ba30e1f48c8947b2d21ca2f7d748878a9271cf469963fc06a162eab68e0969dad0c4c33
z58897202497db0bd9324003c6da3a037ed25e54a7cdfb496640a85fdedab7a90714eaf90ee9f67
z42b8f53daea9d40a77a4fad99ee7ba64b1333e34b619465d338460085172bfa2b4104a9f7214dd
zf0eb68d50976cc98da133b8eec2ca4d4d34a9537d12c73134a74863825e5eec43d421064abb694
z1d5cbcece8e265ea44fafcc666a6fb244b990dc19e3f0036ad0393e3cd99b642ec7c87c8328828
z506a92ac216c0a0a644c811b12ed70b3ba5b96a03daa03503188eb8899fdc4db550d0424e0d9d5
zaa8ed9d0d49403e2de8eda10b4914bd20e8fa80268d9500c7fd0c9616bd3168a0c8a0d6ee1ba6b
z093f244cb9935751cf7df89aeef73fdcca3379811f78f2d02b852b7082f51f5e249ee700bb5851
z9efbb0f8d75efb9364e29f51635f53c4dff96afe3fdced19d0295c4620715faa2e7b3c9f3bb794
z25c3034fd245831968e9160f6bb47cfdb50c01c3ab6f3f885a02012e5fc7eb9880c6cfffa5f1c7
z766b0bc451c7cc547c15c92b0dfccc311ad634c166c4ba3f78a28ef1827983dcc99173a0395c50
z9fbcdf08f1fff360527effb5d9cb8b90321c978d0a7d8c991d275ba19b2d25110d62b0f0baf74a
zac1a5e8f3297a7dcf02b9054c51c815ecce03d04a49a476fda2e969ca7257ee2f496a76db5bd5c
z0d00b2645ed84daa1a9c49d804a50ce5bfb09c880d306d9dc4f30e5720b29aa37e47789ea92208
z58ba7b8f834b19ba1679a410ec156d9d4f0ddf4fedd65de475cc7ea2763d18e229ba3217075be1
z009beb0aae8838f2ae74160290385ca5ca3ccc0a1c7d784da32464709d31bc7214b5a8738c41d6
z598f7dc2e0e163de4a6b64769a30952a01151e251425efd2897728f50e7b7216de46a9f0429e7a
z59eada9e8fc667643e3d8ae6325dade506cdc469ea9db8c75c2f095897f6f6b0bc5296255e48f6
z33fe44bc6690040f9dc65f9cec1708ddfa1ff00a7e5f2059fcfcd8fea4f2211ffea69efe9ff869
z28d0d2b175da1fc57fae1b2f12946c187206fe571dd8ac57959c694b12f0edab050f5c41916f31
zbaf59bbf7793fd352fbe52ad677ec82f21484e170bf5a12d1bfdf810c1c8d7703d06a1f29c840d
zfcb3be9a83a76468d97abb2604df0adfb43666c5c06803a29fde843a7830ff74d8573a1f6f4bf0
zc78b9a8370aed6a48fdcdb957661522c5a700ba3eda102b0fcfe13b5af9705c328c28a0090ea02
z6b56ae7331926e7652b65892013934422e93db8c694bfd1dc9b3ff17ba3ed38bb653d7066a0d80
z6ce42090129a0d2470d918f51b8f98b5783435aa557fe7b2836ff011851379f00813782e0f9c8c
z89fee99508803302b300c7e99b424e26a612e71ebae856142a7e6f3d3e7a56781a078d5232680c
zfec6a3427a554b9624630e8ac0c7930c3c48ebd0a33f361bf7ea770d6b568999f063895c81ddf8
z108b2c1f60273e794d023336fa364aa74886339d84ff76e87b5edb270bedeca77c73e492afa06b
zc9405d4080e4ebdd6507a086a23771d6b1012764c043eb86e2059405f05dbed6ef92f754f3ae04
ze7493601aa2ec807ed5ad6ecfdc2acb42b268e32b875490869907d87dffee4652227cc18baa86b
za0b248537aa459bee502603b7eb61d7b0bb1c8c2810077161e3d01f8db725a0eb85be5442a034f
z989381d2a1ae621ea387da8c9eebd139a31a8884a705051efc00d65121df4378fea628bd5d22c2
zb9ba003598021a4155ecb054aea4952cabfa416052021d383eb5e90ab6f250584fecf13b00c566
z1d3f20062e65dd137f9f72dccd07796f31f637e1f84ea606a1d081477cbc897e920a73600f1c63
zf4eddc262a64df8e81852583747b99464fc422546282a733c2cc120c2b04e5500b9c34a0d6a738
z5677ffb9fb4a20c9ae3553a76412f55e9e15e8be0c8f9ff86051ddebd5b6a36979629b66ff1aeb
z376c49cf1c91f027e190afcef3c5578db4d31798a89dbbce5129c8dd2f23861bc5a5e4f86b9ade
z9535c84d696c63dd78ac4968325ae6db55064d650ed0d521c6a606e706a7cbe90d4514280700ef
za22bf566cff4e08665fa75b0ac630810081f8b498ee112da1cbe1c17ebd305dd3337689f8aeb50
z8faebf1d62532255477800b2f305c149b96729419512441998c492a78685e7c02d0b9ab83e7118
z83089ae2126b4c678f6a19e54e3c169809ad7e191464c2d7ea99883004179573fde47111ef87a1
z95453081a5b1fa6005aa4bfb243d05f6ac572b2168e85f43b5d735ca39aafd388b97542ae1eb15
z0ca1a0277c767d1a44f7b4a411c7857310ebb19bd551d5b83ca6863daec895f24e46a9d63ea6b7
z15805d9567f795ec82cf4d03a57785c77673ad840461fc341b02643ebff0240666c253d3b28d87
z0992c59ca91eb7efa82a83cdef6e197e74f64121117996788150916d997890c9854e8582e75a74
zfc314802a0ea309df2bed33c34d329893af0bd6f726052d7a412179743c37a39ccede63ac70ab1
z6a9b521362f1588652282201a30878e4aa326b1e386265fdd12f2b5470ec3d5c4f4c3fb543851c
zb84f1311919d73516890da92788e33d64b5a8e36ba6478f3ef4e335eabecafeeeac1d3137ad3c8
z84ffccd4aec8e01c2719e1fa1d88b55b0345f9d99251a130b9311a958ed3b6514c5b39beb0d166
za110a231deb0a1e0124539428dc4933daa444516f922216cb6a5302e84627aefcb40b3ee6d753b
zbb39e942fa0234e41788692dc2b7bea92f114c6d90b1b48aea3718e95a97fcc06dd2b554222e78
z7ce6163931a524346f6107c75445ea9f508d2af3aca8b6dfec113cd62ce8e007bf5562e7f43a36
za73a5b1d71cab58b8f035a3b78b2a9aa1bc0a999b1860b19fe50dca59b16982871f1c32f9d123d
z963fd115e627821524cec7fc5a4826f38d8501e2995c8a36ed5017571c1a3839d50a7db9a3c8a0
z88a1b931f8c22e47c536e2e8ff5975268dbffeea7e2c5bbfe7330df23cd0cb50d10c008118a684
z05db224bb7521007f14c90b51dd3bc4b34a3ef1a519ac5f5bc912f3f51e40d0f8ac18bcb38b4d5
z2f2f5252971b28dc80b2bf750b85d50d786cf453626a362f20d2c4b47128b6262ee77a97584929
zbd9210ad40b7880623f6dce38cef668b11e7b50458a0288a560ce74bb106d1e3b6f7c986cdb5df
zbaca62f9543843c84077a0076232f30995fa0dc6b5e20f5586fedb825eb0b93f8108ff45371fd3
zc732e0fc11ed90deaa111ffee343b74749e3e7cccabd90f13e1f2c2876f9bad49b652a2fedf000
z170ef23d38e52fe58ba2e53b4ce3957da064645e9906a64e6a050198fbfd22f440d3f69284b306
z4cdeea3ab5a9ab8c6bef11ddfad511f6914e971c367f745e43ac4c1a17eca9049a8287934aa14a
z333c1f8b7b839a603a452d00262fce0bd6ced5f143c57fbeccc8df689d370dec37252f3f6ea0f2
z285e79a37f7eb22932d57e592e76b89de019ad71d970f3faf0e2aedc136bed044b25ef984ed729
z5ca00b03ab1995864172faf3ca23b3e415a3ab52066f2f9957cce023fca388b4026dc8fa96e102
za49e89e28fd1594dfcab82a4e5865eac70c5473fab9b39ed0d5990a65ca11c0539109ebd41b93c
z84795d77d153b15280ab5128ce6c954227cff5c93f8f8ce78d4d5cca4f5fe4907e54fb8c8b8bec
za3a9a5d477b47cdd8bea13e9755133bf25f767d7ca9ceed286b2913a9e9aa7a21afee771e4e2e9
z8efda5e202bca03fe9e78394da0e4afcee9f7c6403de17cb547795a4f0edf865e828e624ddcb07
z656c995aa34e7efd6601e71b5e285f1f7706d5b7367c58a7e64986dfbd3d76235b6f007e3f4555
z439dcefa89029e64d6e977d8d59446cfb902bac5b0ad89f6a3add087962961330d009573c24b09
z9bc9988f12d930c7bf04ee33ce3724f36893be237f4bebf4720e6dacb8bbe0f8feda2dcdbfaf63
z676d2d5e85d57785430e184a8fdf9f97083b28746b817e469202567ac7846cf63d72e46bd53a86
zc0cfc1778cd6cab5b92005f53c19554e8f23160b8d97444ee376a149fc09d12ea75fc0f29d42e4
zceac9f9a0bfc2942a9cfe8d59c9a9aab1e03be4954f9c7a1dfa19155bf28d0809b2351ea3b0f8b
z6df407e5e1314fb8854ef68f38a1dc3765ea6ce91044be60c1d28f3b75ae08390f345b828d76dd
z77eb4cbbee325d96e89212428cab9739f4dd58db0985465e79b93ef4e5118f1bb4f4ccf93e3480
z83c0e54b148d75f74036fd6afd56aee574b498e7d28ea54fe3c6d1f2462fa4bcb2b602b2712e3f
z420d5597ab9008322d53311f558c264db86af078a46ec721cd2e2e15bd7a06c0bf1d45be8e7baa
z9aaaf5ea1dbafb7ba66a44125fb831217d4ad7d271e7789fb67fe8797f388a2da5f08eaa282561
z244a129f339b4acd83e7feb7db979f4595bb59367246587ccbf351c69bcf2268d6560d4214a5e5
zbabd917e9d739ba2791dba06ffa2d67ab5adbd7e47d8122678b64277f8623b46f340cd7a5cfa52
zb60a950995ee1921962fda70b4fdaa9dbc9b1352ef9da222b48c6738ea5cd978dffd4401b7551f
z2f0179605f148766c218de28d7816c6a44b65c1ccf0eebdef75d533f5d66bf5bb431ddfcf48337
z525098cb80dee94dcd641889a9f817b54f47b8479322940606ecf98027f65ac8a7a23753940ab0
zc3c60b5318c7c31a230d9b7d456e4cb0257d1f2e24866f67923019c0ed7b96d10325960428f83d
z5505d9f14e2ce40653d12fa2c0c0601421cfa592c570e97c6d04e07e5f8a8745cda9269874ba7e
zc9ee6ae2ec60e0ae511da441237e7948d503be4cca704905b02db801d1adbae75dfa81b2e66bde
z7e6be1d8f29c1d5131ab6a3dd26e2aa7e9bf94d2be8111cd59f2473d5b24c6aa9607a006eb96a6
zc6923a1c5e72a1a174ea94a768bb0a283b1ee5724df288587f72f2456ee9a315325a14a444b6e3
z0c783d13cc93b6475e17e6c991111e4899ba16a3a1664d978b4c3eb9e21050ba903be74a5f02c7
z3b292cd3017eea1bb5d9cde4602156a00af45b023453e226d6bebb2bbf094f508599818df361d8
z8e18fc91cd29bf2dc22a58a7774562923b7252614c47c17f65c1733fbf8d12265e8aedecb44405
z92b77bbe4d65a3154d55305f3db2bfa31ba58c2983133046333332956b2a25e355d2deb26b0c6d
zffd069f2f041f9e5586893a38ff22d1b0b598166fe2401410f4fa9766d886e34eccbf1727a4c36
zfbb8aca4bf6ffa0418ee6eef4a938ef8801007de98a311698f7107c1c5018f5e043a7d46df3b83
z0524f6aacac33a6c4c7de089e415ab0b134cfdf4c9250b237fcd55f12074629071a8d0838f6155
zf43176703bc43c606b32a32ea80475c6239bb34c660134b2b76d662b27884e877fa837ad24951e
z20180fb4fb2415ada6acb2ba34933bf1cb2f95b8c6fa592d407e5af30d5dfd705d276296d7a5cb
z3c7ea6c8bcb2757ce7b6b63023ef489e890f6f7f0a60f5ceba44aed8e9b216990128062c7340ea
z12e06270f054d4affa56391fd908b4c25f11c9237da9fcc547bfd54b1f9e9fada0d04bfa2d74c0
z558eeb99c3a2566c417c3640383cfb3910e25da1417bde5c3ced718b7202a0645e2ca14128eff2
z44a1962cf40c786f965e30bd27844ef217b80d1ebf8461f3328a68532665e6ebd913d09906e86c
z351d8146cf46bb4cd2bfa19621af4975d74c5be6ac8df670b302fe03b34687f6440f8e01d2415c
zf2180b66012846b3a74b90ae3221aee30736452636c2bc48b1271a85eb0fc2aca2296da10490a4
z150e65683016cdd9060de9d68dcec8476e437e1ba3c46a084e3c80bb0af04fa2c4a658637635ed
z391867bc75456a2c090e2d2a9245f2440c4a881042f0511f3d0c144db8cfff3980e3d844689c04
zc8aae76963d0724fb43605d55c13cc5077feae50a07290650636866490df16a1e37c85f5278afb
zc1648c5676c5765d3e9584c7f6a8523afa019b6bf2ef7a06f574f38fa9bc4a669b066d79f12668
z53ee7dd1c75b1d41896c03a0291f6d0f67249a42ee91748557c03f6a4305e7f88963b56e6851e7
zf893e648105e1b9308f6f92f60adfe5badaa24be8b1cf927f790427cc1accddb079a08d036cb40
z1e19dc56798ef60a783daaab030294048717c239d6906904901909653ca8fafc8d70a2732b0f09
z2662bce4d728988518b7071be3789b1f5fae410535d3641fbf7b32fbc22efe9bcff513b334040d
z7c7d33e4954268debcc44cc2414dda873e4151ba5d361384ea2c624c1ce7a90e956ab2b70f9fa6
z85ec3a0518fac9dc65919057b044625c9162f56ad2f6edf9ca65944b88d93af6607479781caf7b
z8d4fbee9b7c53b2b319bd3f2ac96958b54e17250b7f3b071cb146eef6e8f6225d2af4e08b2dc20
z0d0c061f45415fd68f27baa48e6115de435c90d5204a7af6a0a16771a51c4d437d6fd0c7511277
zf7f15e9855355b8cc889364b74a788fdaabb94f6a7e57833e1ddf35362f0a0b5779decb418164c
ze704dc5e6478ca8fc61a72fce5de4811333b4938bd9e53a0b77b5ed3ead17c322d69db9b39886e
zdabc5336b426b9974ae4cfc91089ae83fd7fcdd942bc97661e9d8e8b64ec69acf92636c7873b13
zb25168c3f8770fb73fccdd18c35fb3459364cc98ba08063115e3a26a27fcf8602ad356cbddd296
z9423cc9e81f873ee7f7019a621ae9832e384f44df76c23669776a736622ca8b8543939652de15c
z255e48537a42bf0b7492bbb1cb9beeb963cf824fa8335987d162d0cfbb0b3e30e2cc62faca8bc2
z7abffb7a496295ba5def359ab8a672ec52349d9828c765425c7a592b06de2801ae47d85bb1954c
z9a0f1432f37a8b59196643de7788162da029f14a7f86276b6f2a686ec170b9fdfc74b622b79d30
zbe63f66b80e80427e45e9888b672ce1546190149099cbff532df0f71b446fab02b08bd50fcc8f5
z528d6db99f41051890bbb899a53e640871fbf96adf1c0973ce620a500a78ff4fc18d1946c04a43
z12a416bcf5043dc4d161dd8a191d4b016ab34aebeff7892a6760a68a7a9f5991874582feefa46d
z40bc57e844c88c6df2683a1c078834a138a21e38f56c7f801c1db2230822ab9fc3dfeb0a79ae9f
z90c168cf839f6480c2d0a230d8903e4549c27c23908cb4151eb836e867fe2298e3479fd09f83b0
zdabf29a3052b3b2fe90c3cdb79173f604e26c82973cd252544bbfa781211a39786ee9d6ae1666d
z6db27bd762a01cb730e3da589e18930679e4c1f524cfebdf49c32d1b881b4fe5fac6ac5994779d
z59e8bdcd81ceb5f35ac1b3f3ba81b91124501ba7b3d7403fff317037e3a816322d73b299e208a7
za047894c086c018c67f1f0e41a3b05cc99cdd2a6bbdf8cca732bbb63b581fa253734f12ca4cc1b
z3860be170c60d1f254726ff47e515c012effa387dee626db7530df318156027c690bae6d3beaf2
zd292cedde3b70f6f13774fdb11c9f117f0a4f9cf23baa199da0a337e120c7e23876fe27542083b
zdac3f437649c8c191bfc7bab988032c0d2961b8190d7b76625a2cf8e8d2ab3734f454507deb4b3
z8e6b3257b69b923dacbcdf7e699854faf1e2a8e2f5898e1d1cc2b6d96d0e736266a1d9da002f4b
z6434718c22ad518de692fdc2c15e3dd8de1624889fd5bcc57cbf866d892a776f3aea2ce99503dd
z822685ed304529f035059ecb191e2b01da9ad6a47a7c77fd1388ffc68e010a49749a6c41bcb9f5
zf6acb468a0f05e73a8ae9c0b7069d33ea475e3f75db9c2970ed488fc97f3f0a215b93075f25864
z6a4ea10039032886a7eda7f9707fc26322d33ab7633efb6324a96053f19e46bc3e366ae39de1cd
z95ff782c08de10d6f73095bd9ef07d92154f614f665d3d446d95f7f98293286fc59a7a9d89b6fc
z431555038772e0b3307f78123acab32b91dc1d7ab25464909432bef03ceee5dc8e56ec91c174d9
za8d0e75701677e61160dd3ea0e1a47e5286a7e4ae6253a28104f4672e32ba9e05cfee900249559
z44b38cb0d4d83c5c570fd3e0be33be69883aea7839872119c9f0122716e6528a0a407f16484691
z2d1fcc0d1c4a3960f34c07d8aeae3c07af64dfe3a13c9faf471512fea13cb0ec677d409cf860a5
z92a154dfcfbd9b9531cd6ec2632d62231d08b309ff2f672608560e2262e74f8ab73be593bb87aa
ze3be8249108e811e3d9d0835e0454276a6e2817b10f0e2ebb6d5831f2927ed4cba5c13224073d6
z7de9aed3c4aa14783314718610ed6f01f6d13315ace3d4fc1399eee5454aa70d505c59707d71e9
z28f7b24ed013fb4d7f0b5dd3697532b93f1447b423aaa2c948a8807278ca944e0256fe48c3d499
z4b260709364f8ceb7a4cb4b855176b308aab219967dee4a202bf2d70d12af6d676f5fc67e418d5
z20c23d675869ff7741d82bcfee8c2d774040f8e35fa171d14c6422dd59a12d4d4766a825190654
z30363385274514dc111007fea78d45ce31155a86af3bd6715e40c355f8a6de2199ba6e1c25dbe0
z600f6494a4dbfe8a3de759523ba62933737c52610181b61ed9df0e65b729d1bda12391a60df80b
zaad3c38f9b370313a9a3067d9c4b27be66ae1a5eec5e0dfc22419c90c0a3223ef2b04ec0cc268a
z65672a8fff1bdd9c3c898cc89dba656028e856da58884e60f949b5
`end_protected_0in
`else
`ifdef MODEL_TECH
`include "qvl_ahb_target_logic.mti.svp"
`endif // MODEL_TECH
`endif // encrypted_0in
