`ifdef encrypted_0in
`protected_0in
ze74c34e226135848fe16db9ffd31815111b6d7fb642c521a3f628cf6da949865580b22efd062a7
ze90adae0e65e66a2c36a587d0a790699161455169ed55a01f2084f11770a774ec4c588039b380f
z6de9c5084882a40b79a175f5c2114b2b6d78b070cb806e1c0aa9258297f4687ab30857016fc53a
za25afc8341302f0c829d94450c399b8ff9b0386c187cb854ee330605b7b59da379b1f26f488e1d
z36e675f0b1336408b3a1ad87d0723054f952fbefc8d5a33eaca6ef5be8f42bc59870a29a5cc9dd
z4fec09ce6e44cac279651402e7e1f590df88ce49ec26ab39f12b4a02855703c6f03b1e85c797d7
za357087d98e5b1f45502e45892e5823d6fa4b762932009620038c05d74efcea7c3fdb38901d620
z36515d0824367e48d1bc182335f158c262d396cada6b0ad58add4f945eee634c2dceadbfb5118e
z14969c29a743830a07124bfa78707f3952b96b0db7af7c9ff36f77137d8c490c4f79328328069e
zd7d5280e4f95742c9841340368b9764f0f80413adb175ecfbdf3c40716abca7b8cef6f7fe92ab9
z6bd2453f1aef7f7899c5365c5c83793cacc7795c269413f6cf0dabad14d40e9285afde8c01a47e
zb61893788ec5060288cabde8fb553f21b02eac61ab0b48ad3d54f4d1d76508b22f0c600861b5ce
zcb30ba708be817b1f50f59c0f6fce449203e7355c1be55b662fef3f92ba58243d81537761af8d6
ze27d7864d2dae99372b2b75bacdc0437a4f7e011d68c3487a89759e3625548fcc920ad06471ee7
z2d701aabf726859343208b0a543c73eeff8406febf277e3babff437ec820fb49d6b78e73bc2353
z884917487d35a6cd06d7d73ccff5f05355122888b886d178a03d8eac5505df521c14d1e332b234
z86bc1de9891c0fe4654d9d65be6ba17e0f35eaa0e5fb8d4ffce747c7530d86192c5a60f63648d8
zec2b11ca4783a37281db3c8b2556885556aafa013f24449e0a06d5242cb51399b3e756b814a7f7
z7d2f3363d024adf895ee1f4c57fb3048cf14f737f4f7878d0d0c6b48a3aeecf0d16f61ec999e70
z8673047544b470019ece6d4e6f8a1469b42dc3022d4e7bf3ec62c2af4cfb08f5a5de608628cf8d
zd4665dcc3f4867d0a07a836531edfba94cdad9d90730ba8b6b2364b0eba1514c0246e78124c617
zf6a26bec02cd6601f40650424a431a340361b2120bfaaaee24cdba68de41a962bafca77ee84e80
za2da1ab25b494bec121443cfa771b7300360491417b42658f3967a20c16d3ac0978600bf5db91e
ze42f8327318524a1e54cc36e7ad8520c8c816f80b84c9ff0d9479576d7cd1672ef64238f1abe32
z79ae3fc34e54474d5a8bbc35c838dfaaa353c658b05d461cd2c8f49e720db95e635eeea7febf6f
ze07bb4999f7223c3b56cc588c86895b6050939610e70e427d2b96bbb9ff98b45729947b56fed80
z5eb57ef463636c3b8fdc404f4f8c82fb627d1860efb4331021037b5512f7c8f3dff2e029a05125
za88736637ed02999a0466d8d994324513e3ac1dd57e28a44d1e115b3c27890613b828c4dfa8f3f
z731dc647ed8b84655f5fbda340c35ec5acef1a86178b53870689f3ceb95c6d43f5206dd16ab0a0
zce2cc6bcd032298b0ba041ff22840187131dea9e7c588ed951f20df7f24b4afd1724603f49bdc7
zecfae5585f41d6ca3d3a4768ef112060eecd07d667f2a7428ec6aa07dbbf0cd1f19ff350791b49
z68cb095bc3b64b0899fbfed94269a621e6edb9b15acc6efae28251dc93b2086815a1205ca8522b
zda5791a010281b6427ff8acfa83cfe83c05b0e7a86f55b5f7684dde1c20b18fcbd656d73cb41d5
z7dabdd6deb9a78ae8adaf9dd9a35ebb4a2b93c12b050fe05e02c1f9d685acc8d9b5c6b322e8ffe
z6965f5f5343a06a3378ab10f093855f0a7ae05ac67c1edc2a2fc1df3f57e8facab1b8bfea73051
ze0f0f55cbe5a1775c7e4274702430c0b35df624ff0efa60bc7464ce777b78d5c96851509db6462
ze7fba17471421227f91ac10ebc4016eade39bfce8e779bdb84b5b8b794532604ebb7137496a8b8
zcb9103ffa3381394958c11a376e84ebd5a72ea2fcfc0aeb5e0eb151acf9fc3858c954483af8ab9
z52a95dcb8412cda704bd43ede3eadea729027d71db1510dc3653251b071d86faf16e7c89d198f7
ze6573cdf9fc0ba1dfca0ffaae25e55051e51117ddd236d4421249f87a6c6f1876b677a98f324a6
zf3d784ca01328b251bb75c37516c62cb1ead4f6e1698654c1cddb7118c6950ea932e0a26562cc9
zb310e40ad20129fdc8d80837cac1425ea8f79260fef7fd016ce555a3835848c701c41a92de24bf
z7304c407be20fd84e9b93841ea37d54e14a6b87c057da27106472e88a0880dc37dd5c9d9e38baf
zd3451bbccb944a5b7472cd101803bf4aa30cee5434912722f31c47540ec8fe34db95f596b253e8
za2f3d093b34c62c27337d5c167b58f32e4f8384bde8ffc05301de8ed24271ba3a4a10cb4b494f5
z4db61538713e3f8dd765867bffaaf1d89252021fde2a05d657a4bf44a73ab3cc3b4058f594d252
z7bb1dd175879c83d2abdee24d73f2b8148bd03a95be581789359a8aee237c88d136bd92f8c3007
zc262e585ec5afd07270ba5942459c97775ed2af7c9dd02976e760818d3af02391792ea48494987
zba4a3974345dd2b9a5c9c2c38a96b94e07c715e7e2ddc076bdfbbc2baeceb8bc633e5c12947ccf
zd8c745db6a979520faf3686da3eb43567a3841e43a13c75448c7dfaa2e2095d3f224d271dabf5c
z31a3ff5eb59b14807026ee75d0a3f49d8d23c90bb837d340615835ea5d58f808a9aa21fc270ea1
z241b60223759ae7d5f230963890ec60908db951073a8c4babd75ce5ea7bea0808d67d930b18e33
zaefa0b9030b82c34a79fd770fa1c252066925460c239715ae18f8088a1924eadef1861207268f7
zcc55136f981770af1873478ae11e656ceffbc46310a0a5be59496dfa0e593850600551123acec3
zc759d4bf1d9066bd36a4b887137296172f2cd32109140c45c391ceb0ba7067246ef6fe4efa7f13
z3694d8fb20cc55386911c32382dfd92db1193697dadaabef9166bcf6749653b40114952932e2aa
z727511cf0d908a675f4281468c460399c9e8233ff4a16f5830f9e892349e0f6f932b13c3e1debd
zebc26240809e5d774a5de8d6ec583c6fca7413a1968f21a82338d1724a9ea1c194db3077399949
zab071a07cf581d7d6192d1eaa061475b0413e3a952a8e3e221aa62c60e889e17da5313ac6bb9a1
zaedfd58cd996792d0d3776546087efc07082a749633be520e40238067d1b9b6c4cb05e384cbdd5
zba825890feb942310534ce5c37b54624ce564bf4e58ba5cfda5a476d3a5ae11e9cc29f371215a4
zd0d70707ac953fdc6fe90d80052f28b47ee6758f15fa95718b6cb4347ed7e138dd4462a2491be9
z8b7484134891105386e2904c64720bdf9af7ed6dc230d0be256df98df34a7db0db7177cceed7ed
z854800162a678e725e4e265b51e8bf87d5b59c686a67ec7ef0912836839a916aa4fa0c68f2f172
z637a507d3b92f95361a0fb0b09e244227809ad792dc9d5ef28e9555b1744466a67c2c41f89623c
z5d35f9a285152b3c154065f2754cbdff508c0c76a09c01ddbb804505ffb7d0181de53121892cce
z2a582ac9e8fbebafbf54d32af1071fa072ff8872cf57b7927cf5c0829853739ab9ee714ae05e3a
zd5040f07802769e941f4621af57b204160a6f3eadbe9e5d29943fffa200b2dbf4cda3eb8960de8
za895dff9be9c64dbc38eba7cc5d4216aae7b9e197dc13495280ef167a65d200b88aca95b961c18
zde6f55cee423b5ecef13328364d19a2f6f32835ff8503e84d7e0452144fe8c5cf939e0405449ef
z2a41519b7a9d0ef01f556ffff1f56c05a2480abbdb0de9760aea1e06d9d03c7799dd2f86456f81
z37433d721b24f27d5e774eb6abe45b5f5286c229f4eb7f872b693edac30b869592c061c2b650cb
z1ac3b0b1f922069f3e062f4a11a27497d11094685fcadc8440f0652e0f138d5feae0b762daffae
z8ec4f42c236b268336508119d07949aafaa5c86209492aaadd6b246970053fb28dcd30def2258c
z7d9b17a9bcd2ac28d6dbfba2b9352f96cef667006df764dbf510fa43c7a6d7c82b9d1b637f72ac
zb9962441479bd6311c6587a0e36704f3538fdc1b594be6621d9f23737cdbc54d7c12d9453aa20e
zc514d8ead4d7d7c0b6dc9b926690b0bb6c32cf1d2b471c7e6c3c7a12499ec84663e4705e1964f4
z5642ff46838f95f4349d872253b0c9d2b51ad3159e38245bc12c112cdaf7015f3ccce8f1259048
z55ad84889208c067b6e7cdd98403da820c6c549713cb8f623fc98d4f19d0b0c33f0c4504d716b8
z3053a7b96df572008dda58438d533d34d80f17be6d04bc6d80a89ac7bf4acf6f4c95c1dc8e087e
z45f289707059a2e4b00e73ca4a660d23d7db68ab3a60f9dd39816d3c695b2625e73c20281c19ea
z5743f68592774e7e7bea5b763c21a51ab2271245228428595ec147550dc372e5539435909a4814
zffd5270dd979bc4b021af020445ab0a25b9a987399e38a8cdca6e45672be15a39602bf69f97c75
z90aa96e6ee04af2da6f418159f5164f0ab96144c048e8aeb6aa0e6ae8a5c098fe881d619fec47e
z52c9a85caa63cce300fa60a3dc2128389a1c5d9bb85d36952f43f8ed4b8fa101081aa6a3e8ffc3
z477c5f5caf08e70a38ba3e1a10981b2d1e2a716b96b63efef363fcc7b281488e7799a79bf3f13a
zef32af924787e33097d255425f1de88c09ab4ff2dc05b84b8f61f37948480081ff406f1ca6f3d3
z0e5d6ef26015095beebdc789a24b2918198fdb448ea24c365825e532d5b4470186db88240cf5b4
z4a0d136571bb101f3682e50d53ceb016f47c05a864d0bab24546365a1738c8825a1241e475f4f0
z6312fc7fd87ac0a7c6e4721b0c2f1e80a82b886a3726cc7d009cb4f41b3618e7fac4f4d766c9f3
zda047020764127b0ce9ab5d928b1d394058461b5288218b7dc5914abca7efc1a5e34d8dbfcbb38
z3f58ad291a4fe816c337184eccf30ebd256675287dba88d0b603da79feb9dbd8c0a1f1cc9bc141
z8aa13677dd02816e1aac0ebcfad060b125176e76d70e6e17f2b10655fc13c0770da6c97076136b
zb44caffbc11ea894c914cee4cc989da9ede219f82501a57f16d08e6a352d5af29405622dfe36ac
z80c23baae50921d95092c08b78e90abfb4c5e5f767c6281644dcd2ac0b7fb72854fdc6cbe02803
za30eaed0d9ca13a464c86dba64945092f73b73c935a9beee019728bfa2fbe700f0a57301ca5cdb
z4b5379bb4f7fca372ed4240cdcd7452b94797e8e62d5df02780159e2b2976b3433b5133dd451e0
z29898ae912c2f21e726b649f2a74976c312e6cacc68da043fac33fe489c6c87e06b3330312cb59
z28deaa6856a9b869d9ba2cc5506e916ddc27c7c3f29b4a2a6b257335b4089c077d3f33325dd157
z31b372ff35cae713b9b67fc4fa57726b63be6715b1ce716396d17ff7747a85c40dc3189b43005a
z2f9627cf7ded26614a38ba6f11ad462354eec27d566f101616b2259336aecba86203a3ab3f24a9
z7773ae1df1ccc0b45de2117fd6075f53735523525a32071e1c5a9dc439434115ef6ddff4105824
z1c41c5076771abcbc98830d623082687ceb19930a8799d67f9397c491a5264a96ba5bb7ad6df0f
z381290249972c3573e7a630d0434a1b3b4885d84351dd0b20f6dddd625be88fb4b0c021e4b5126
z9140ec6a40d41ab42008f4c967d54c578dcff9c8a26a79a34d6aceb3c760c1f3eac723bbb61515
z819fa20f42b1298d2b4e1d0bbbfda7835be817a505272b89f6f8f9d250dc685674e7f72088dc48
z192359006e2b1d1c4fad11e496bb03e3f4db8854a546fa86628053a1984fbcf819b80c0c4fc89e
zccd7e1d72da77af44a7555a07e7cbff0ae909674def772a2fc4d4b8b03a570276703a503d7e95f
z681dc4cbbd825a0a862b1d0f494611b2a42cad1aaa7703027c6e8e5b21c90fbec8c947f7db1f0e
z935128d10bd9e5e660cb792ff0c83adb6a8bc36816b7319534bc733af725f02ea1ded7fbba012a
z3fd03bcd26dfb1a87aaf2f6058236685da7230a6e422036d6df477c39734f9518ea7baf505fce0
zb2a2824df48ddf2fd8c24c08a999449874d3aec528d2326e87ecf24db4f83f9fd0cfdc8dfb97d5
za950f7e3d81391dc5a661e3d463d1cd5188aa37368d98aeaec093d511583276211802361f5ee75
ze4349701a7a1c903eeef0b1e36df3f905e2339b5ae40f7f3813fdbb3ad5c09c2f5a937a4445987
zc9f7651845d8c7875ebe76a268519c3bfebf73cfd85d7a06315edf1370ea0d395bd0b52f2d0a5b
zb7f666c303c70b4d3535efe081b1617fd51861ed91a82e44f30720266b550ac1afd7cebdb6dbaf
z2eb19ee3c39c437747b57a71adebb2a15c304da527a31124f5574791b7ef54130478450d9ce2cb
zb529002c05a40ed6d90599ea10ad42ff4b5f639074402f4c7ede53bf8875b09190f1f17f6e9318
ze063f590313a89b822c6e9a257cd6692c1e1732646b3af47cec8822a4f8166ff656fd68c2da8ba
z5576f1baa3c1b0c4e8e3457cbd60fc706bf94b058a8eb6e08033054333e59a2752be5add6ef047
zeb3b8177bb79d724cacd823ed0d2ccaddc8e7427ee26392514c3c27f0efea4e9ad59c32a9ec1f6
z723ddf1e5b27e7a6a584b9347a4fee5e913439c49a3fb137205f6b65f2b8b6f642805f2e769624
zf879a91d8fe277af92974a93e7281a4a3564a32138661906192034be3223c5738342c468c092eb
z8728ad97717da6c3a9fd19785b6d44958a067c69ff52c6c01ab40dde531ff83be90563290573ea
zba8bc78e1ee50092b0ee138509253c66335cb60310dd4da644ec158ae37f932697c7f8a7846e18
z03acef342780bd4ee24a6023f73b06c71e240b10a3057f606256ba5e012f2a08f4f01ed75fdc94
zc76baf339c875bdb36039701c37abdf3cd8c255a48abd53865f80572b73bec025ba91b62cbdc7c
zf7146c328107f9bec179b4034a3682feb221564906df8c3c24e82320782104a1911a7e6fd84326
z9fc54daf77763f7bcd43d33e1a31039b25d3e0e491e74d06e450ba7fc8823605d77b2fe6e41b85
z80b0e028a8e8fa3289d1c240f22817f2ceaa4b584d2b20011819a0ed3475e0de71d76f4f8c5eb9
z77d5552c81abe2da34d825f635138a958ab0b9eedf89c20206ec8d7b9833eafe0f6b47cbfd15b9
z700953b9e7c797ba89baafabad01a1505a1df24bd7127009f5564110a3e9f2684be0dcedc2aa15
z4adb7ccd79ff9b239ea994e9664c385c9691fcff693a27f2d43d1a0e483e7cfa97fb79e6d89439
z957731ccdd16b728c9b3ab1c3bc44ea0bb6234193adbecc1b98f347fd568f9427db8f754bf8e50
z93c947f76e55195b8d7a3438f2c8f74c51a0f5e0b7f2aa0021afdce37519f154cb5195458682d8
zc0168832c3aa6e9fd66f2beabf61e46bf4899280ec8db5e4e882a66bf8cde55346c9f6f2972b09
z6bfad79195ac97ef2c3c648c50c69bb2dde9074f9e7c206e905ddd858d0e402ef1839b8b2783b3
z89be9e0fb34c8881e74008dfd61487ec5f41b53538dd4949819fd9906207a1c190aa33968cc246
zd95f82c62ff761b68d35d997247605400d9cfff69b5da810ba4181656252ac7157f10ec8c7615b
z63a2556f1d8a8540534f30a3ed6403267c1656420a0f7cdfc7d9e59cf6f10250afb8459dd065d8
z5123c1a30118112038408c1411fb6311f7f2599d05580cb9a957bebb2b845704ee8f8a9767a708
zd815dcf6d2e39ab9d36b3a8d50db0a1c596820bc2d2d9f1706a6a5b6a1c0fee1b1203943e4e161
za5d8afb96588b23fc82fad2de5c5d30b37bdba8084b80c25782c59e33630e2935f1e7ef740c761
z494f3c38e2ebcd8d04b70f237cdb7c9df42a16165e55528fc39af05fd8472d625d2821916e4055
zcf8f5b340c6a73e0f42c803095e3ad1f96a8aa73e6d80c34ecc6b71df21e4779a77051ceec24f1
zdc365cfc50701d1739c9c08d7dbe21dc9b833414d0e9ad306b13c602d1fe6be529efa342b57b8f
z9a1633a93a4a330747c186c66b681af05dcfa1a617f6e5ff1f09b3579ea153e70095c723173bce
z99b2e1506eed847dbc164f0c41ac74655b6b2d34a27b25fb84d7c10667a59eac1ec7dadb015171
zf5f04a6e613dad902d8ade2dbffbbcd389dfc52177dc6fdf7136d4567f7662ffaadc5b5fa02734
z9870cd4a1e0fc3afe7cab6c74b9b06f357334ac9f8d937370eede8914dcef711c8c24c573d7d4f
ze60a4ddbc7743d2ad0678e8adf625f24739c3203db4f4e50017049a239a49ad964396cdacb594f
zd80e1c173043ccc490d84037a852f4b8dcd7a28321c557c48e78642a5a92121cd34c345d860bdb
zd9c80438c33d50c20188e49bc68cef0568f79333f7c3b2f0084a7394eec5347cfb150e412445c0
z0d4ae4240f6f5f37851cf5778a4c6c6e1965da2dbf3552dd091d91adc4d970ff5d7c3527681416
zaa6b97b288c9f039f50ad48dfa3119419f6c2c7ace018fb618a19357d5d11d9cc169852c17072e
z1321994e8f4f99ee7be2d781b3112ce028e5d453c160dadd8fbc2468c1874bbf3e54d656cf4979
ze39e1f79d7ba5e0092dc70281814f27202bd33c9d5a6bd9b2dbc213d0684902357cc32f520e8eb
z7cb30e12130a0e96a8f297b67650320cb8680c4bd41838778973f246ce49ee307fdba1146a9569
z0c63ba97950593c99ee72bd0863fa641cedbad4147f0bee4472dc7f260056d61f553ba40392613
z226b759f14f01bbf140a0407d7a69e3a26dcc69d62d6fa73f03469091537e44367670ba1a03878
zc443333e93f30a900b2d9a72c3d7fd85104b0532a95c912603df610b7c2c4abbf5d21c48ad0c42
z3cafb610d0e3cf8e9335d2d7f29db141de55402a3d657d501a6cb804ce70ac340ba82bb848f726
zbca381b0126736e994442f0f7abc33688809be9b15dabf6da23aea753a6edea7751174cdd8c7ce
z0559a5d1d291307c84b18e6c51cebfb5be9bb1bc0d151ded7228bab4f3a96276ad98e5359c9603
z09356c4401743a7a3458b73faf45ec7788b715704768b9596703b70e4133ad96e89ee8ce10fd5f
z68fb366541f7ae60ad82e5425c5fc2054bc6901dad23456ffd5718096cb9bbabbecb92d923c3d9
z942ea771dccf72cdbe1c9956e788699e6b3f4b9dc25a5d320e71980a9b79ba9ffe597b7e84bcd4
z912fafb91f2bd38ae0cea9f8ee4c0b09a0343fb2316d9299f9b76f40426a5f76cacaab21998fe9
z262742a7291338d92e5b4a66f97378ef0f14baeb77cc30787d76a85c34b63f4f9a1d0e6f03908b
zfcf029e33b105ab3936ffa4211ad39e38d452a452f9056f8850b0ee484789bd228a8e9bee013a1
z281b63d38670fd45645095820646eeb8c9fdc5f2d529c03ad9dfe623b28fbec2ccec1d2e6b94e3
zc5ce4b4ac8d1cde8ada6b072a2fc49646765a4be53d728420f643c16990ad833695d2d4ec972e3
z2671f59d5a6751cc6fe0f2eb7cca636f26f5df17432b8cd5cad0e4a559eb3d20bbf434030184d3
z4d638433284b980838d8d3d8b6ef8967b37c57e5efe530ee2df15f9b1b93dc6cff88c0b5901c00
z2df3d6bbce8d6842b902b103cd73f79703f101771ee6b098c112969a7557a038ae72e9b5ea7750
z337e673349c4ccad19c7b59d1abda8c38e78d0e9cc51a280d7021dfb0391beeae99bc7339cd2fa
zc5a29fec7b262218dbf83b9a0f61cfd7806351b317aec1dea9b92132eb0b7188e7059afa8bad13
z8f87ff6c5163b9125a07cc8e102edb001c7816cdd5c5ea08b75b71a0801b0945c289bd3c420611
z2e49f4b87a63825df3f887ec7c38525d7db94a1f5e37235ea25dae2ab6c99ee7b6b9133d2727dd
zecea735eecda203a84c90247a54e54a7d0fa5873320674d981b6bd1a4819de00d5b4c480bd1642
zc4175b0258534715f6a9bc13d4f078fef0a8c6807923dd83c11a9ba65ef913fb9d68464f9bf5ac
zed8e36be4455a906a3a62ea00f87095ad29e9fded683c623b1d889cd3d3e7d4fb148e03abd0fa7
z1709160f2ddc4154bd2be73703e4d79c6c2a6db646693d607d8a5c377756b310d5d0ae665c5c1a
z130a9553ddf2dc10968b1f782a350e53eabcc9feca3f3f652f21d88bb67151357ba3614f19b6ae
z22b0c1be28aa154adb296a207b95d3f02439be06f76a0e2c6300d58743022516d31065af9739e2
zed0dbf89d05d59fbfcead4346ec9f58bd8c1dace661ba8a0ea810b4513a2bc36394ef05911f0e9
z0721c0f040d3b0a3d7dbf5a4dde1e394e305522d8cd5ea576fad75a6d219674ec28657e01083ef
za45b5c0284af9e97ae2ae1ed17e337276891f0e11a5de34afc0df65d483a48544a3b1139ef0563
z9bccc6c51907260861faa9dfcd5ce2ea715b8037d648358e6cae00bb2a23da3c400bcbf71c59dd
z3c9a0a0594d83e08264f3962beb85381d89465591292fcb20e0e694a1d474aab086e91bf424a6b
z005d2e0aae58ce74fe5253d0218cf642f4d0cbc273d7e4107d552b47ec021f9202ca2d02dd89a4
zd9049c4910a0f34f6cd7301a9a746d4d4decf7f6f6e86f9cea64a2d98bf342bc777e8f602d60ac
z8272b1424849271c27b346419c3a9fbf97d28db59b967c86189e6a0a71798add7e13e5555cd76d
z0d30a665f42161f3b3bdb8b9745645225961b7864dee1c7ae6abd8e87d035bb4473897418e056b
z6191a2ec4344b6e472d6397d0a365c220917c46af2cfc01364952ea488777bee06b1d73400b850
z9b1473f33758b21d90a19dc262cb8e6b2a4631cef2d8bb051058eba2a0f03352dec186acfbb6ca
z4fe55669aee6df331b0b9ab914845a8cf8e343960ac2d49c4aa3b153b988799d158ffeb1f3c8ab
zc9239401502d9231d04265d2075882c116f386ac65b57787ac574c83a0b4f659fbb1c3ef155de5
z85476bc4f30a474919d0b821d541549cb8baa2cd62a408eafe4fe836560cf4d3c18f2d565b36c2
z359b7b905d03caa03075ae40137f6894bc9ac5be0511b5c51b1545343c4a3c385164214ba57877
zc3f9215c9b52e9339271db2f8c9e94827bc0db3e53ed918084d1f7ea194d9c10f6c2a5aac1bad8
zafb5a5910eac91e4f4d1bae6376b3f3c73be3b1f9c90fcd374750804fb217ce6fc03407f67b95e
z5cca0caaaabe5b30925f73eb080a9c07f8253d2d52042098a833259ddf0fed38d0715b49cd5b0f
z604d1463cece11e8b214905df4d75c93a3a0a360be79d8caf2e13c9e01dc2c78bd45b6c8ea4f9a
z4071b6e4419ab682daebde36684707eae050da0fc62fb4741f9010474453bdfa70ae4ec7e85188
z4143e0f03f25b70f3669c43e74b0846d8848533ba95b21b607b831bff0eb31d6d76adc29cd7169
z1cba6b6ec58db1fc90e5025c67b82df88de959b99356dd067b08518a568f1576df3e75db0cb9e7
zba91b27f9f3a9524422454e4d8ef01e961aae8073dcbce16cb7d1cf85d2df637c7c1a81e3abdd6
zb50db77eda22c85339057267b3508ec10abf69b01a59a4da9bf52d31a6b4e98b3c3cfadd7b8c99
z90a6c47a9528aef2e8dd72f3d9fdffdaed2b4daa3824dd6353b121731f37d6eca3d6cc365e4360
z9dcbb3a19565101762cf96501e005fdf52ba840b1c2232755da0ce09689e0aea48b327f2f1c746
z491b42a3254ec075d651f9b8cf6c66cd36769043ec7316c6f8269d354d5a1a553b1db9cb97a2d8
zaca62b79f957b3ccdd5f4a5f7d4e47b0172c854695d6bf8a9b5f4fe08e7c805de39e64d5ee843e
z124e317ca8b0b911c706bf9ccd7b36837febe293b09543b0c495c78fa81d78061d3a58cd35442a
z6fc20abaaaa7f2a591e2fd3eed4c146d42cbd92ec66941bca8cad7690a70d929db9833ab4ec126
z6277231ca0c22e845675f23ca088d85b42dcef7f735362dfa4f5af4e268211b8124cf7f1fad1cd
za0e9b28d796f34472ee5b9453243c797d4e0438b1eca4b2cb0ba4610dcf93d3818ed23582dee54
zc9fea80eb76b23fad471bcf9acd12b7e2d10ccaacd151153627361d44d0525ef1871877af97597
z5593e602ce1b8bcf1fd6f81d717651801e01ea09aa969edc3d9dd6e55ce03919efe6daf0e9c558
z2a0b066b069d3e4c92d30eb23324952a85891629f3c324f47cdccc31b121e06f60a8ef442aec1e
zf5368d2de97b87de36d5abf1483b9b50b4c7cebc66cb00eac669336276546d292c57f5467c22d7
zce15590317af2d9c292d70e36ae84250761fa69d4460cec5128370d2f0352b4fdf75d19c166649
z938748101727e24e55a7adb783f23af7ab37399a06b21e6a9a0e1644165bfec44869dc11bd6c07
z9de8d9ab3df84d2d20667fc729175810a0a012b0ca7a4b409beb2961270698fce51168647ea8e0
z6c5ea8466209d42423c629d5b76e0a0f6b107c941d4a3053e301844b258e43b6c4711d2acf5b76
ze3e29363b2be07052065c6e1a1727532c169608073ae9da03e84be8565c374ab1bf1060450857c
zba606cb3cf3435d50065deacd46f761133ae7bb31f1279625a1ca8fcf152d2860ba6e2e08e982b
zbd4886be8cd7f6f0ac01abde2ed59c08357085a56e2eda6c41d206a5e71bb304a8ce541f177ebe
za14491efdd85357bdf6247dd6bb3dc1fe24019bc34fc80351f68004bc469b0340af4d5c2ffb370
z796164e2fbbcf906f09086381f276d0d1e453ad2f44bdcae7c62f9a286348424e3be0473dd4242
zfd968387e36db7cfe3518b4d5011e3c6e6944cdbe3b1887b3a97002756edb6dca1aa03149ca807
zd1974940d65b8ec26fc2c80aa43a98927f0d3fea30b1439ad7eff2bdd14129b1d4f93d4cd3462f
zcc01ee58ef2e20d633ccb17aa0ab863eb4155466d2fcda0db39913c9197f0e29543bc66553c5b0
z1a636e453cc00b81dbbafdfc85ba7a2f2278e0c67f58674ca62bfd5d0bca6d577507d081c986ae
zb70dcde16f1323dade5261614185af4d1b34f08e4c8f2e5bf19c2e641f03e5d4e67a9722dcf8b9
z3dde4ea1137c232a9da9a66242d6248c9486b43b53ad27a5547a263a94c319700cdcc371fc5948
z698685bc48fb38894f46ebcde67cfb67035920d3e307760c3f8985a7b96c4a40e85fe1eee2e664
z766559c6475ac6a479b240de6a5ed780cacfbd93d129693952c6e3f0fec5bc4eacf8aba0dc0f2f
zed30b716b049fd9aefb7dfd66f2b023d2e721535dc4d63531377f5102f46c351f9fc3dd66a3cc8
zddf95436908eb568af8cb75794bc650e4d7fa0cf75b77c49975907410b5e7bebc281d60a4ca7c4
zd5876d6709382d38f63ae5a62b5f268997bbbc2e5cc0e4f340e8907728c816ccb0368474b4c16b
z9710848870dcc7d87cf42d7f20c5e1bc92994480607e1dc48684d099426bdd2018d2f636cfb333
z2e64e7c4fabaede17d5b3a3ea765b25fce6c95245c87f5e1a5e95ba7a1f5bb0db207746479f0f8
zeca179ecc2431ed06d46d5a74232f6fc17aa0062ed8c31436c1952a02f44cd7a3e60e06fdcd7be
z3af0ff9f32f2b1c28c22a1963e483f8c5d2328a07074eefb74df71c55c19ef522be1ee0b863c59
z71f40dc3fc72b77fac968a46dda50b1601448d4e3a23aedace8f03b1dce17595e251779ee5fa81
z20268cc5da37998251832286df4094cda9928b1503894bb693a609d022d2ee27a4fef0be6c5bd2
zef69fc8f9ac3f9736068fad2e6efafb172157e5cc57c0bbcc47cbf09336de33beabcf1ec3e7e7f
z10507fcf41bd2321a17f0e4b93532b121e85c573534ef7cb1d3a3b67587d88e797080892da5ba6
z67ad7e6ab5a80629a6a6c8564b7cd3ce2b65cb909c17dfc7ee359d915a4a7a09f2a934c57a948a
z04c9be5be4b65cd7ced72a1a3eeb24c92ced453236054ddc3d684fe6fa8f69518460b5ecb719c0
z6798b3ca73e6eac19d5c1f7f9167e30a741783487daf0851cc3dd762692c3712cb27bbcbc4ed19
zda29c2c5f23749095feddd6d8fc96afdd42b04120c2a94f83d547e0d70c079de09d93d56e56c60
z5baf41673a8c499b4e0862053e2cda4438f61ad5c75fea49427ea7decab538b698cbebe6fc1bf2
z9da7b1efba429f45491c1d4a0370306816aebe5d01cfbc3891a14bd9be933edd65c892f38bf186
zea8b47ab0d2e5c09f2ff49538c135688584db3c4ccdc290c0eea6d6f368f253e76fecf4bc05f66
z896db30f5d60006d18b30bde4efc0a0e1a316ae975f3dba262ad9e2af0b80e2c24deab76beb39b
z6573e655d4a199c78f57d451be7e53cebd29c724d45ca9dc6ad2ad1c35139685465569d2efa05c
za16f92cee2b6e4512cb8030ab72ab6725b284301252bcbdbe872f5f09157e1d017a923717f7e20
z92712c3fbb79e6c4b347b8c1b57c01ee87ea5e7a9309ba9f1032f78a03afeaee3cc35f1ae539d2
z391b5b00a49fbe1203187594f01e1dbd7d53d42d775d639b65c3dd3b53576364a7341cd21b7ba3
z716f66d665540844a35a687ff07ec82cd09622ced80e39591d4aac93780fffc853a0650e96eb6a
z330abb62a43ddbe1a7f3d5afc17ea7a8d999444ecd65a158b48f38025739f0795de64e0c3eee8d
z3c4a9d26dac10ac2e990c18132fb787ab108e9fcd171e4f301cee97f180c694d6b4c03db76c4d9
zb83a57b003f0303924c84f5b745a9fd9253c5f12a3d6f2efe2a9ba8d02398b96136c18b6c60ff6
z8cacaf136d9db56328d683badf6a7de40762f5e277100ab103d2313b3db2787ac3f01446873581
z925d6f599d594693ceaf54d27bd5c6da77a1e897fb1e63246aacc2825628ccd6a438194a194097
zdd092a911dd843a1aced9b2302a273e2805b5d31309ee60151074e0cfd8898aa2d559768f516ac
z8dc6d4df9ffe9769a0c3808a4d2588ab941540363b846aebc6a464c82212874a47a29bac4c1991
ze968f264f11457257a8bc0b87fd15c6a03c7883e16cd46cf85ed6dfc5e4f30a169b09585fca305
z6c5515702cf151ddeb8934f046947a82d57d00c05bedecfcdeca5f9988f6382e960719644f0dfc
z24fa26a2501427caed355e8acccc1efa040e4733f55638fb714f8ea6d4b353768fcd3fa2f54a7a
z2712e95ac5cd1653d80be79cb6ca892ce2aa79d178c46f705f1ddc6ce90e009421e3dd58ee6baa
z475071c4f3ce39ec995d678ca7d8371f2ffdc7d2dd72b1f78c14270f42415b74e37a2cf3fd595b
z43686167a36e48e770cccc2f7f1340e020b4698efe709d3733169e56992861997c7231ca101b85
zcd6f50fe5781d8b35c45f282fad16fbdf59201472ba6d678c0630fb29b49e9d4ec8609a855952a
za83468f4444ae96e5e42358c5f7ef432318130a3d49fe73dea854c2cb027e97b29d2567db178a1
zda8a91ff6080e7780aa1dff88fffaca529d777ed5fb1a810700ec43568758f1a53aef3c9c9fc80
z83ad25493afa6f6aefa7d1ab0f2554d1108b524b98722a4c903ccc2bf0e6e2185fc552b65e7a20
z2371cc4493e41f82c68014b8baa450328621b353606c1a7e7b25e5295807430aa0d4a39261b93e
za6f1178d9ee72876ada368c0ba2b33dd8f69341fbbdefa2f14ff253c99e3c4d8b0543bce027c56
z88d87725daf3b6a89a50d0fb60f25fa32ac22468657a7a3b0e28f41a1f43bb4005a4207207d8c4
zf4de49b78a839ec16f2a04702f0e34978926ab45eb59fa17484c2c1e20a322517862b516ddcefd
zdbaff80fb75214d6edb9654acf0a102010118ca6486b937a39c69cbb2560d10c3cf3706ef686b9
z0ec7eb085b1b67ba18b9680ace4c0a3b845209de3e7ba74a4069c3e180fb981e9143e364d51d4a
z8ea591a58d09b2ff7a24bd84d9f43fe81950dd1c6c51ecf618aab8c9bef6a5a9a4e4e7487aca3b
zc8e03c7c8ddf05e8db7e184fca218e9c96af3a454acf470ddfc082aa5497c512f1ce1afacd156f
z68b8e4b1b50ae36338f8bb2b8893ff9b1b183a1ef02ecfd665b505309ca909d6aac28c5b53718f
zfd0d6985a9a31eec808808e7c92ec377c290ae439bfe0027aab6aa57dac0cc3918a719b434ade5
z254d35b82018b1330066da00908e0a92d3088c6d35ad59eee72185756c50afd7e9132bf6c08a48
z27c98f1828601c01a346f899049fab80346b4c7be194ca9e4e77f4a68ad3a18cfadbebac8dbca6
z40c97484e736d796f1668eb4a1e39306622c8320f75c8ca41d64ef993ae079c64a5f1bbfbff8a2
z16c92119cd256d2c8586b3cb2024c30ccbb9667287dc1de72848bf3dd0060894379a33dd0cafca
zbff1dd17525c606a7fbb26e4805a7cba03eb39b324dc1434fe4a9e83f87c19e20b18fc9ac4f6bd
zf7c2bb53d077f99e20568503783a48f36870889a83edfe32bcb7b5dc309f35b70cb04aa94018b2
za7d86848896f6e11619a7ba21fc813d1aba8e32f8cfee84209d85a57f885f8a605789863bebafb
zae2dd179960290f44f420e273983a7af4fbc940014cc7c1683ac54999dcfc5646189fad4e3170f
ze2dd6a172124a882790f11d96edda2854eec54a85737a554771a968657acc691783d39a8f92f3d
z113f9a21b7f521a0d3b98ee7c1b3cc6e288928a84b206584ef5b700b434cb2c606cfb9dba8d9ec
za8157ce31681d2544a0883c5cccad1924fbd8b483c096d23280156118ff03ed99328e2d41ba81f
ze27dc4d372fa5b366f2c7b0160027980d88c73976ec0f31d9847c199c9b1433f0a5e0d2201a9f9
z79fac5e226675a360b92d3f54add3635006e2b020ead1695c6900ef49172e1ebae837c469699e8
z09c7aebfaf5219eb56072a11445d1edf52e3a59e2ffb1de7b8fa52b36317f3e7889b40e872684c
z35f7682d636e7f5da456080c2332cb15b7b3aa7c31f2816d294b8de615a6945c0b389543073953
z839887c91aa08a0fcf9258bed2a6a5735ee3bc28b8a528b84e5bb2256c20a8321bd0a66aa82a3f
zb82b5f755eee1efe8a040874a4634593c940487f106226a4d2e65558b9aa1132ee39673491bf19
zda24e9d6ddd5f6093e5ff97db5e81508cb337846024af54ad1ed43580f515fcf539c730fc47984
z6a57828777933f91f3717fbf48b48570ec424b5da13c0cbd7289cd6ce26c7b1535b8743bcfbeb1
za9a0dd94dbb19801a59d2eb813ebb660328f09441c69387219608f4b6fb1f5905780b2c45a2181
zefd329783e60a3aacabd441420678c1fb272967acddf5e49c67f7fa16748f1df36e423ea5332c1
zb452ef0b578c0c40c9540796b79a6e76493f06d92d5ee5033287de912187be9d55f774603c0b46
z4f60fdc107f563c2642b54a6b5a864f770d8b6c753feb00030d641a368dee236efe6757386f07f
ze9881ea7cc87649ae8acb217f1fb78f2f1ba444cc41a092d4ab66f72d06be6a542ad9c5c02d131
zab03a73357306d893e2a77be284f714937fed0ad2414a60ea983a4a57804eb5d10f76bb9541707
z074acce87c981d3f834cbe8a3e2ec8840dc1539b4b37a6a0918af1da03995a3799782af4fce70b
z0b62dfaa8c9c4c3a596e534aebe019cf61642ea4452eb8e7ee79795495c4a26e63b57822b47e75
zd10d9a69bf5ffe998c74422b84883223978feda2671152810e64f13730a159a0b30c0e4bc107d6
za72304e7caa5b0a5962c3db4978df95682b3119ffd557f3f85886d8319fc1329606ad8454a3afb
zc91c1d1097b88bbdff2f0838f3e88f886287a474f888d6e357c38e77fae1ff70395d5678e571cd
z1025dc1ebad05a727db9cceb06297481d88263fbca26e30fd42af52c62bfe5ef5ad7973fc2514d
z5db6def2554479781883c6dabbb521a7d6aaf0c52599c0c4edac6c9e6038b0a5e08a4b4986fa4a
z7e7effedde9586bfbd38e03aa3b7df7bb9d8ec1136563270930089468139a13ac08f1d7e63b090
zf481ac4fd256be1caaf6949d458ab8f7f843d29ad07d03e2863ffa804846849474a9ac99c36113
z5b21e59b2e64ce7c88d23af5d3226fe6147a7a8826a5fffb1417e55b70fb437308170650e90b00
z9b1cacab0d68e6d8d1820be1b1632fddc9a2a5f326c58655e736b0429359a135d2437308d2d5aa
z5d0551990fe48b2f7dbaa884386aa27bcc37e397ef3c01f20aba7ae564633c7ae239143dc20a28
z1e053df6674be6e6be24cae769a3dc200d843f32d03bcd58ce4968c61e6b737a69e5d039a96223
z64cb983d7183dc8fb4bb157feaf13338222a8259d62792cc8880d04dada81671523cce54bbf445
zf64a7eff692d87a59e54d937a0f7663608dcdd229d420854c37b15b8aab110cd4b85a12baefcdb
zc7f64a19d8dc910cf01433214e3e93965a35ab69e9f227b25dc320fe66b7488f38e25f49958edc
z0d448249e6df14cbadfc136ae9eb4df4e54f7d54a04d796e10fbf2ab63c1cfc237bd5ea6b499e8
z882f33939474d2a275c3a6adb81a7abde350b884d20793a1975ff4ca6093a2cb40a10470d4e4e9
zded67239a00431626281829196c940bcece34c9176bc729bb3d0d0dc37563a7ad4e02f146d4b5d
z3ae4819bbcfa2def5bf261da0179a6140895eb696fb2df7657fa74099fbf0ef3238d2523ca6e9c
z75f7f6d019a56c5ec47b229386618a04137ff3ecf2d1e06939d7a6af9acafaded7b1fd3caa7301
zc67b3e41313682f8ae68b0665b952d9216f4c575dd7e7a0f998ec24ef158cfb465c487777c6727
z4768e3e69d28e9f1eef83e0ba6ed39dd997e17bc87359fecda4a2373f0edffc0f15e0d16e3e476
zf73b87981c7caf5afe976d355c532eec8b64866cabfb7d3a076d05df94eba67b27e9555e4076fd
z6fddb2308282ae65f6a9cce1b633355db72f7053bf6f559bd3d75cac5c65c76449c5f73f4099fb
zae9035f3fa179c6bb6c4292e8ad3eb08776b85d9fb3857fd9de5195993f596aa96d6cf72bd82a3
z8ecc9991df25f99039a6d1d55ed8548e947303fd47d6665a5cf9690316b563e7c943551ea12729
z6773a6650a677febde1af885a06c79f76818e9c3dd91d51f554911c90ab347ae316a3f7ae56c36
z542a1d0d1ac74dce7337a716b42008787afc5b021666a9f58526990eb94252bf00e226e8c84bec
zf27cf05244d3af90176a9a7a789031a8c319f0973d4944dcf48297bb4a6ff4a890f691148f96ee
z6d23ff27ba055820471137d70166561ff82ac57a9835c291b0ea6b6ab88292a83f985a64b58ae1
zfeab1b392b1afdbcb697f6ed311976b6e1aca4b0154194fbb10fb4b9e44652ebe38392acaccea2
zde83445a1d73b280db38056d2653f57a2d179df6b84dff94dc1de87b02a78ddb5b00748d63e5f8
zfe82eba31621661bbd81264622cf253683cc841030adf7e48e1a3cf1fe6e5ec102bc8a16fb2a5d
z568c0ebb749e29e9fa85c73b8d5282abe25d332603bf0af1d878487c6aa4d6662d9503df1910f4
z0f10f072b0b03675812cf6340b3f46a5f39f993c676010b150d869e8b8b7676e584881aabaa306
z11dbf6b4ab2dd437569bf4a29befab1d4c05bfc1547568215ec193fd8456cb116fda04fad1fb6c
z6b5e0f7a903af0c84700c2ec6c4fffb6d559372b3260687aee863a79e4595708646fb24b0bcb5a
z1bb1ec9dc5c008289de7e9a80a62e8b473f30d6df3dc9ea56c64b9ef9bb8eb52fdecbeb699d621
z5ca0f03e43f9ed9c0ff862437383d7a67f5531740d7e975f18543d1c751cf1ce07b0dba94c0555
zcc6a0ca6dc8c46f0a846291c60a14397e5808a50513dc50af469282733a5014a2f8b519e029bea
z6b8994871719902ea1ad4a764d8507def6f77590f499cc1b497b6464b559b602b39c98f77b5942
z05be27afab94b9e67ecf7808ae6ae51b956483d28db4e14f6072c6ebd1bb2077beb23baa740a1a
zf416156ef44dd375d772a2a23081508e73bfc16e087dbd7409bda03506b7158cac87f4090d4eeb
zb67f563e21b1fbe04ec44dbb0eda59bb20788f468ea98bc0cfd0d2f4a8d346f9860e89bab1b668
z983c21c575300e296a5f1894e0dab780e3e8e802a430c7a130ec3ee655c1e6861d77c2de7d758f
zb334a275a28a7e42cd7d4198838742978c602be5e928a433597c24da1e5b4b58a7dbf8e8aea6e3
zfe067e0098d416372d28f5a40d160457cad7e82e7489325d65eb3a190a3c1678263b9bb11fa7be
z0d8af4be5a9278e6bd55ffc41b6071a67a8524835d3d6e5ef3e33567feb7ab4a3424e6114df1e9
zad34e6e2c0ebd6122e35246aa0545aa0df3d0e758aeb833381deccf0b397158b7b5cfe22f67052
z047e34088459cfb3026bfc34fb2b156fb8b158351e733767b6eb8f288907d9092aa9e1cb2c62a1
ze4b3b9d749e53a05ea8a9ceb98cc42af9a58021f466c54e012b838c9bae3a3f5b0293471c6c0a6
zac1b441ed8225d2fda99c245e5e3b9b86cbb2047ae923fce4deffb217783903a855ddae28fb4e9
z8bc609d0dc565be32d4b8747f77ec6cf6f4dd2bf18eebe833f0d1fef94c7ef9ea0ce020afe5c40
z756bf9ac1dd8f5bdade87b6c3b7afd583cfd111cc193e4be8811dcd88aabd699ad57bb659be293
z4656ba982179d9912d62393204279d94ec453b19e714da20cd46018b3cce5c76e19e6cc479588a
z842456124fa9f2ebeee63dfef70f136c59c6c82c8895af2f8a5624e882c355e540cf7910739cf6
z1df33ea22a5e96f90c08fa12f49255baaf26d8f40da3a4a06831b914f828b55c9f8b4475a1398e
z96801ec63009cd8d8c7e87a0416d7fdee502b98da3bba4bc0550e79b12fb000d91764e7f74864c
zd4be94ccf44ab6e7a500033395ffc673cca23407e5140c454be20741451d737dfc144c1f6e9fe6
zd04f6d9c924b00b0f8015f85fff48e1c33154f3c4798171941bdc273b31f8fa231839dbf578ced
z2ae2a8231fe1108b68e22357eae3922122390ff41738057772fc6e628e3fdd3646a093929c1cf0
ze0d61070344df87400e199e949a8e048bcfb56524987b789c9e9f86d259b36adf10d7c9ef9dc5e
z5d0ff4ac85ace91a95138a5f9a4798e00ecc8131c4844c7e7a6acd396d243b9e103de000fbdebc
zf9b20712db2aa9c05e9d2a9baf8c05fa0a1a75dad5b90fca0cbac8298df0ef05591fa21b2b89bc
zed4ebce839354e6dc32ea9bec80558de926553270b00728fa7512a1662ba5e0cb8861da6d537c1
zcc4ec86831b8ebd9f7bc7ce56d36f7e1ccedad40cd7a4e83a8f48e1150a65d7864c92d7ab5e6af
z271a7fa45943615503607634d7eaee28bdc4b111865ea94ac4d49ec16b2ab34891460e4954ff9d
z2ecfac6d7649f8ec89e6000323cd2ad97e6639ec758f61955ce246a674dfe0d2366ce241e44e6d
z339a3246b0d7135119351f7cafdbbf03876edd8431156dfaa0df28595ad38b6a1ff29d005b5607
zed6ab20912e2ad296e9e14a004202b006b9174ad4704ee5d256bea60733f0d25641c00b95af038
z8cf9da7757f0be0b108841454fe9f500ceee093796d57ec37f7abd63a0f0b6fb87cfe2b699374c
zdd75be0786e9fd4ec37da360bb359b4411b188fa25b97368075be49f5c99223a10ba1c6dc92f07
z47f5b22f145282eb5ff4fb962f4e41676f8c94476f15b88fdbbda908c76a3fad8b4657c18044ca
zf1dd793017c8cb5dd67bc9976dad9955cfd05cd1607d157d101a0eff51a1f398cb68a29c27d85b
z472ac4cdcd98cfd1d879c932d023c08103f664c48ce82d295ef9005ef3d011e1c64d87fb573bb8
zed5415512c6dc3daedc9751b393005e8fc444276e1dcffdc18952458ba2494ed36003d39735aa5
ze2854dbf1805f8de16f3df6109744b508c6b4e39d3bbba8e2dbf61ae0fef8e650e48aec879641e
zbe61ce7c52012c2e99487e9bf17b853a9175d84908401c1fef28c58ac0e1ffcc90f70f3f7a0ee2
z5daca68561fddb936b7ea192258370ae22a8d8766174c12d6edbe82bee66227929becb9cc9d376
zb5b26f0c354d2cb6e06adef6a177aa1c6f8205028ce6d46d094e27126f799ccd4916695b0323f7
z195b0b741f4df8c3eaf131c4981001d50356306dbfffb8664aa12f97ee810e16ad93ccdd0ce95c
zebfbc070d3b72b95d5624157f39d370e9f382c18d9f62f88063dca6e96a2c7ebd650d9a4fc6871
z3b5702e464e525b926750854cf275be28154b3fbb047ed81d01be5e91c9c09b800a6af0fb8bf8b
za4ffed5e98494fe7fdb8447a68ae526fdc0c258983bea3eab2296904243e153e71bd60889f4599
z0249fc9baf6e47355bb0a1aebee6b67cd8205fe30533b8ba2e99d3280b7023b449dba5346c5814
za13233e4c8b8edbeb25969f8c9b84cb12528a7ca55bb3364b82bc85834f055d638c46776425b58
z204cb93d66d91fb01997bd114ad2867febd88aaf0cad56ad93ca580445c8469fce820011da2c75
zfa97244533dde8a57786716786dda7bb1b26eb50d1acc3ef5f81ec779facc5485660e343589a0e
z574dc75721c327152dfd259db7facbcb1f8908a1aa6a7a83987e1d3606ac28b80a55375e7a5b3b
z18f2f6baf4e60e1d9bcdeefd3cd713e744a83360ea836f502dfbcfb0f4c84e4211c9a0d6781899
z0ecc3397068cb936fd289a4dcb4637630533709cb426f2643657dda89e9d49ee6815dbb4516b2c
z807f427a7b6cf4450b4b3200fe63a521e07522ea0ca4bf0323d069e561675fd271b4e5cda3136e
z55092706334469af9e703bc2dc515e49a69e0dcb57f16673d549cfd59f90f4182bd36207d6472a
z64b960b8943c80e0677d6aa2f505e210a6b9eb2e0ac99010a3341c1703c789089b9251eacdae15
zfcd1ae809df24d1a7060d27d6ac1058c4bf22007a3af5ebb80913f7850d642b163cd3c937e10aa
zf7897b6b5c9585a5225e35a439268659986ef343c6649c5efbcb7ff08a876172c0324eed25ccec
z0e990e0208739472edebd7a2af56adfb5b9f71dbdebcb4f02abfa2f39ce2bd79634d75f8aa88c6
z2192a17a34c5f70340d4d0caa707b70829e8da4c7011865ea17a6dfd401ac9ac19dbe8e2248c03
zbe76b9fad3fe6f73b4a0e7bedcf4db1c25c3a8388fb0deb70c174035164653948e6313c6abff7a
z8ac7d60646208278aad06a5113276ee7b7e67113410c1a68935dfbaec6588373ff5d989ce96f1e
z02284f61d930d4cd5b1d8ebd0e287ec3b360c671b0dfefddba518209921dcb77b8752fa9bd90bf
z369e24db60b43a561ab820e1f0c6509df8c02aaacee0f1631c05da8e718338d67fb75d19e8af55
z6f4d7d1ad712d73cb299d20a5c81f7b34c05ef786970e4cdd025a89c3418250c9f9deb4da06ddf
z82ca505d4c5a77feba7cf2a82af0cbf462d3b56eca976d1ee34de495a66cf3379020f2eae4859d
z402bf06e895263c372f1469244acb10c7a86ce1f6b88c30ae1a553881f9f7dc16aa866a0df825a
z62aa0263a6e20cc21be29e74f6b38e697d11922530cdb934945be3ab5afdebb3cb787d65bb257b
z6db76ba3063cc673cd42d1904e0978b533dd8c5954a642f49b89868dbdef8ad3b49e7ab20fdb84
z6e6d69e05d72f366a1cee22a727d2a3db7cca5c24a5e3a9e1cb931d2c7720316c889fcf3f38f2c
z63374c02514e9d01167957bfb6a16d01784ef19600f34d7687a9b6de9d766593ae7e07e393f73a
zd3c9dc7fc26c95f12cc90cdb30cc1f07d5289b4a05f61993bb11c2d57c4ddb8670443eebc90298
z3f84c134065c64d487a2e85caf5d5c2bbaa63c9716c0a2ff2970ffdfcf35acdc9a16d7af9b0a1b
z32057405888db540f5c7d4c1e28105017233e74eeb3cbf37ec020c24e8fc762ac82d930deb0a81
z9aad1c7d635fc30c0f0e7067efbfab05d435acbe8f22b0e7f3bb88703ef49ffd3c72a95f6f98e1
zd0dd80b2b6495fab5aef1b65280f4dffd889df00ad8047ed9cefae921cdbc3b72c57c775f6f758
z1cbfa61b5466775037d242d72dc41e92708bd9872c8ab139b2fbe516be7ccc0c5b4d809733073e
zcc041c117ef05239735f98836398c88bef26477bf4c28f8cae6a2f9ecbf9d7a44502e879824d
`end_protected_0in
`else
`ifdef MODEL_TECH
`include "qvl_gigabit_ethernet_lane_deskew.mti.svp"
`endif // MODEL_TECH
`endif // encrypted_0in
