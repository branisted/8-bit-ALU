`ifdef encrypted_0in
`protected_0in
ze74c34e226135848fe16db9ffd31815111b6d7fb642c521a3f628cf6da949865580b22efd062a7
ze90adae0e65e66a2c36a587d0a790699161455169ed55a01f2084f11770a774ec4c588039b380f
z6de9c5084882a40b79a175f5c2114b2b6d78b070cb806e1c0aa9258297f4687ab308bc470f0040
zb0b1de382961eeeaf2e279e1462520fc31c119af8f2b214846f56c2b3cd2eadbe4099496abff18
z15cec83ec4a77b868344aa20ba7360908f5c0de2a79abf8b3534b883bb12180f68b5d4beb444cf
z3fba8f13afb0abfe8fcc4294810f75afe452434d2d0f1166236c82f76edf1e12979f04bc35693e
z32ae028996dd85737a8f5adc1ebb94f39c940246e887647b64782cd7ab429b0544c173176cede7
z01dfb26b1f73408344a52b7e1f117f12bb9c8077b34876c2e6fdc085981637012dc9754765e1a9
zc512ce062e0b8fb16a214591f5c81e1353b900a611fe1f4886b57940b41b7f2ce99a7b84b04b90
z916f717e73bd10589c81e207ed77ec660a8cbed5b487fa50acde1b055c8870bd8676023f21ddcf
z9c98cc47cfa2d654ff1365d1f45035a045a66c5dfa827905026270f0d55cdcaeacff2a9a621a2e
zad9d2af0fed53751e72de9a2364fe801bf0b44df415b0cd8c966e2140c4ace0f6bca24916c79e9
za4842f4b48e7bc018f2dcb1ff0deb8c32733ae18960ff67f75bf42dcd9d5200feb19feda7ea5d9
z7ee36374a28d10a6be7403b733bd57efcbc3e2b99e25ccadc2195f641ced7b4d99a8147e92cab7
z13d94596eeaf1e2df1e32966a30aa2f9ae4fdfaf967dcdc01225eea6f5317b3b83a3aba60ecbb0
z580ed4f036c6fe454687543cb2c699ecd601c5a00ac413d43448f92656346397b9ff1711d27dee
z6839eb636c4817bca8b72d87b7740646d21c37b60bac74586379812a36446211b20a41af4573aa
z6c03fcbf5469b77c817b0d6b904d8c43f4f23f30894010ab731ad19aa8ecf96ec5cfbf9b32c1ed
zf7b1ed41df4bf415bfd460985cba8af6ab25db1188ab3e3cb20519cd0c18c6b6225c8619c7d5a4
z46a5a669b278d4bc2f984ba4db5feda90b4e7c51d0d1ba515812abe1484468098a980b170e5f06
z33321afe854effa15188b7342819692d94fe229c0ea6b7a5e83820c8bfe6c8380dbfa4f3d2f992
zd510ca3a59394268a35d2031cecbc5b790843c2499f135a9e2922c2434347f2178be2ec1efadd4
za7338c206e8bd151265927fb37cb42c6ea41c097901ccdf201bd36dbd469834d5747bd690b881b
zd56bc96715b443432adffdaeb684f4ee8f46b673ceacc12cc7095db8ef89c516e46b1e1a984e5f
z46ef56a9d035d879963b0983011a71970e476094e9026359e53cb77ad76a2bbb3879ec27c63580
z1ac7dff7a181a87c4293d4ed2e30c95cd8e58ef452ebff386a6033e786f79f55238442c28c31c2
za5311fbc88fee68395e0800a4ee28ae8b97f76122ec767db548d0619d02834011d2456a2f315af
zde8931d6c53be0b616a64e5141ef167a5da62dd4f53762404c75e9183c4752700380e2553d508b
zcdee7d2816f6f87b9bc07e1e8e1539601118ebe309d4e9cfcfeffd5186922b52b49db03c228eb4
zdf513d5f560d09f577d5e903cbd3fce0cd246310adc12a57287969255acf4559b0b2479351680b
zbde0ef7934a6d28a58c6336fa9ed4e92c0f955672d1c131e293ed23239191151bbb952b4a304d3
z00a8cc5ec93bed0828f42300edd84a5607d410261278101648e1108b8966f8397907cecf4e1273
zab697f6af46a27bac93346864a69597469c4890ca93dfadb18942938de9990b2ead7d5b570ee5f
z1f663440b5e8b634f7aa0c4b86c8488f7f214e98de636b505e702bdfaecbf8dc8b8b1563907079
zd5093e9ae52e5d922e1a432f6dbb02fbcae3f704bb7c9c85a82ff102f29cd9b23583e74515eb5b
zdd55e9e9447bfbd7405636986c92c5723071c1a857021741a3431390460d29c9537d9976564900
z213034607589fac72b5d793e622d83e105524f3987a189dd6f9a2ee1b889ef050eb1b4caf088a9
z6071de29e455e924ff90dd89c9ea6bebf9622a86d59479c70ba41947302e29157f8d81e995361b
z8a2eb1bbbe56a3feef72c85833f574056f2b08282a1c731fe9f226831e9d04dfe5baed65cee44e
z6638a430523baf4295b26d28d676d7f96dc5ba0d66e4896942dfcb949139f37942ea25ce7e8177
z7361e8f2fb7cdc1da45c81b95251829e8c1ef7f05b461bb01894b6d03969e052bb299853edcc94
z9ba97f65bce9988d69a3ab07cec313200980e511174dffc6fc60458af7136a8472a115965e153b
z6a019e64fadd03402ebf067d085b56a9d276fbe0fb8eee90ea1ca79e7567df243272b8f1190cee
z0775ee2dc9fde09c6d31eff227daeda66a2d58ac7387b9e835f77edfe1d0d9eb553b4089617ade
z531f5356a41a9891ff396ea16ed568bd56bb3be40838753b0077db730b35cc8cd39fd4849f0909
zc537eeaad5ecaf061d1cf895f7bc5d5f1f8cb6ffa182121466d571e09a509df2e2fd20fd58a638
za4911ecc2efbe1b8e674fcbf58c5436557dc61b67c18e984858dbfb878e5f6b779df47a5b4f314
z4c5262d87616a59212de4583059bddacb0beb191eeb489a6fa9d9e1eef1667bbeea7f218cee4be
zf5f513f47428d2fc7d723ced671795b62b7d7e15110ffae9e21b4e18b598ccede32886b27b179f
zc74dcb391048e45d1032b9897eaf7571a0294ddab741ddda4f89e841a6f5c7f8e4b4f285d8dc94
zbe44a47bf6982735c872c1b53e9a3d3e3a6b770c8ce8dd602be586cb036782c7ebe4cb2943150a
z20a37f7c99204f372c7211acda61fe3309679b17cd87edc8130acbc411f7484e3e8a7dd6651c50
z597f81d00cc84920c351363c33fcee82890f896383011a888c0a76a22b0a855bf12c5c1e5c7725
z222b264a02864f50a2d8c06ad9b931e35554d6180221e069fc23b253d96079ace97590b216adb8
z1a6bb650aa425703d759be8f4ba654ec8ad40ed6b80c18f4a3ecc9d27820dd2f2c53b2c180054e
zb80064903a251dad2f6266ad58be29fdba8a0b01669f8eedbc6dd63bbd8da324a996c4c5c2ffca
za8c42ca1b47a7a25966e6c4ab83b752110ef6cfa926b8707f20a955eb28f027221e1155ec6513b
z86653b6189c1772bc64a368021a54be7d8c94e24df52b130b87fc94696e98c44fdae57fefb80e6
z7a60d521ad13461d4aef74709e68990961118478e2244f2edcaa37d85ea3848387c25e1253d8ea
zd05a173983ff5da352b109a8d2f619501dbc79faeee8621df09e86094c558b645a25429f765b87
z349f8ddf79ec34837a52433f27decca38a1f28a0395cd185529e12fb18abc3b0899ff9d4e058ac
ze974db053cbdf3eb04f03e29faba9b8ce09c32e96122164bfd4a5aef885c5ead6849f1d7a05386
za0d18a70a5fd12741d6ce3e58a89c3f7c8ae949d33512ef18209a0292a10c69a9e992b9e12d140
za00fb443ec20b48466a4c06c79fec1ed5cb1d3637cf256ca6d03f239f8a677aac938b7793d32d8
z97fcc8f3f87cbced3286c3b3dff20149c3e25540ebb0bca514fa43026649bdba0b29e00223f455
z0f42be967166dff1a625248b9eed377f0884203d8d63b7e43a5aa5dac1a4d6935fe10654f1ea30
z04c0ea1f125506db1dd489d7e3274f91befeb932b74c9c05395942b40693ce98dfbd3e72a6b3d1
zfb45b81280aec61393c3111d5b63e1cc834516b489a6efb7ed598679158e6bf9ec16f8af1e929c
zbdab117bc1319beffea9eb34b2828194750b585a6bda6f8c4c71064099ea1d5cd770f542ba2ece
z930bd01846480e1153a7f4838e5523e79238ce6a58f5b0627f95aa99e1c7bd19a19f6da6ced734
z20e873ae174a3b732dbbe2136706102dfd215f5f809cf637504db2316a3dd5832ae640a1592826
z9a71897e44cf84bf1f627c12fac2012bf3210d6295a9a28736a632e176f900021dabeb73226bb2
z5df65d633769c19a706e75881918f214457faf2c846c7fddb79e7b033e0e6d276b60b421cf50a1
ze53ae98f6d8a4ba5e016cefc41960bc57d871d0f642f823ceef51871c84192227083c5e5611f43
ze1171ec40db0f5a00d2497c83832e39afdf739f537110ed7ccc22ed27896ae7192cbea3e0b2391
zbb98230b756d6c9da0e8203606f9fe5158b33c0b2db0823963378110523a9a4ce5a76940316d94
z0547874680c2e0c28dc5d0753784ae9f359e3783505e1004c2b676ad2a22fe7c8bbcdfa3de3294
zf7c97b1445153cbe46f864f7c0becd7955f97d98ca2749885155d6f66437c8364a469d7b90c55e
zb92e0747b78b86fcf257fadf1a1b997bb5a8111b7e4e1bb95b2c4a8124ed4040f75003e7d16f23
z847378a1ebbc73c1d479bac828ce121f0f42ff330e38b7cd3247c430bc899b125c1ecff28821e1
z02472d4bb86fb39e169d67a1a3614df3745622434f4c06a1ed7ac47ffe6e80a89a038d8617cf86
z16258986a68d6b556acc50494e1aced7f13424bda180c95c9247effb9d29e1628d35bfa03a2750
zc35c7c71b0f0350ff5dec3ba60bd4dc2a2d87fdf1ab528e8dabd85a66bcb3235532ddc03c977b6
z384e526bd09c3efa6cb0f0388aebef806a4ac3cbd25c3fe4df3de0bd6a13ab9d986b9100c9058a
z482d81c161873fc717e1a2094fcff0923ccdd466b169b2fa45f8dab660e6a10e249b693139dd23
zebba93fc66b36ce1e382e681648418a4ab7a86bf7d7f50f2c3708554906a8938c44b6de0c790ce
z6ebbe1feb5347f7fcd538872b4b94ef99f48c247db9e6da33086fcbf0172147a1b7fb6b6a45994
zf8fbc8b1f8fb6e9056ac5c96e4e8167a758a3c709b60f172ba647df662c64382269d361f6eeb8f
zc373d88482f6d2cc2ebc42af2ba6dd2056c2b4bd03d53f21a380d9a11eada37bd0145dc365a12b
za1258a2c2d3f59464d1aa441ca70bfdb8c2247d574c0c0be378d4ee47679126e4a268e6b4b7125
z9a4d048afc965d97de937269c71b9e93a0f2ae821ee0dba6d06ce187a995c0c54d488383fea7f5
zb538759d7780fc058e1d06b90c638723ad4a094e6f9ad86fe6140ebb873ad80c0106649d51cf0e
zec7b41c96249ce4f41cdb1b99eb745f073df280beaf5d8a0ffa200ef71ebe008d6b3d193a04554
zb9c785d996313a909b9a7bc731b2d27b41f3fd5b47ec7258f440b5a5e0afaf80ba44bd8a39dc62
z48a9d2b96c9558ca10176e6fb34a97afa94805c2709618f8903134db91271405c089ca2f1d55bd
zdbce25548dd7b954e1371eaa6ac0af7e23b3717b07b4891bcab90d8881f02648b25b1ca1e832f8
z4cc361df529684fd5411283568618730540216a0fce01bca9fa0f622bb588cff7c6025bfb3a60f
zb623d97d0fca7d6febd1c48105a03092900be8f609cf371f9a3b2e20c09c49a566331c0837ba70
z6e11014eb4f2318e1adf7a7d541bdf8881904610f5699198aea52ab06f1649d7a88f30e5224af6
z59a798131d397c189b084351b69534c8e8b84935e33b13780a69b18b24086eb36bdd1a7eab0cdb
z9d3a9b467a909e6cf390437729629f9c7acaabfe938799186db049be8d6b02d366fce75eb1ff64
zc47a774b3c2f630e1f4155b483b254ab8b59cbc245e25d0aa2e1d3cde4492a52ea8e9a02a94582
z61376395d660a8ab392f38530e775a41bc0f7c76e175d62f7f9f8fe0f47a360b616638586e6680
z126419a4e3d83338ae4d6cfd496ee38bd7cf172e8b3f74c22828869ddfd965c5d8c42736ea4ee3
z888a3fb2dcdd590493bc73b542c91827095b7f96857db5eb2c6c5b85484238ecb06931ef8cbccf
zc43c2410400cd0b93d4a4569e48a999587b46e474f180e3823be2aceb75982c9351a54e51db5c0
z1639c58e3e0224647a03efa8da511539cb1e40653e6950b555cceabce36e260fdd2885eff7e2d0
z903d77a4bdd4deb05391da6c8840bdc073f0ed40730b25455ac17b152221f5e0b353f4595aac0d
z35477bd41807dd3b51d246bcd6aefffa32ffc53c2a4f365d838d2ca3654a8017edf7213da44cfd
z6024268177db9389ee7d0f2edf9860092fb6177fcb9b43d32c626722019ebd50c1ea36652dc42f
z576f615a0302ab95f4c4af4cc78d5df0543987c99a3b188162f5ea17cfca44f9f0ce23f6c12cb8
zddb69a8ed6b0ad860b085f1ec38cc2631e917397079d57cd0386b1d09cced6c765cdce79167c48
zc9b7e31d45cb0fa02d881f9b99bc121d270c1ea44d941beacd194db3196c772c51f76afea616c0
z66b4e3933873f55ea662859f611701ecb5e8b773598101a5290931e17acfc18c96cfe4c9896fc1
zbea24efb2a10414b66e7ba2e7458f0643bbf99e89282bd4ad2e4977e57706e2e6acf5c00f4a0eb
z9d12db134d7e8af1572639bb3a59b004c70ddde49196813403b394c40e51cbcdf8fd8d976bc33d
z111cde053a42030a931dcf111aff6e0f9fab8e02a721dddb2b9eea7c402190b32fac3f6cc9d8b8
z8c0e0f52c179607d515c3d2866269e4c197c52fde20339aae3cf30a42f41c06776ed7e9dd24246
zf670a7305974dd6669cbccb596e8f75921469a210079223a6439e4c07c7f37846e163b87b2a4e1
z71e953dc540d4bd50083a75a531801199589afec8b868445f9cde01f5f3694353080aaf2b4a1cf
z4a9a79a6e6a82e1cb391b45793926c08050ed18818d291077563d072f0d18122b2f7f09b3e8acc
zb0029d03aff4cf0c7f7197d8045a79e6153721436827fc74db3f684b9024cfebaa69343c14fbcb
z76d31c495a311922367cb17f7d07d6e3f98479d15652d23eec34624c30993bc1b2c77a5d74c6f3
z7bce2387acb9a8d2c921d951a6c98bec54dc8836ee7929ba6670cdfdb45ecdd6d73177a9f2430e
zaef27f5cf1976e4cc7e9a6a8933b064a57fee6f58b4978e46cc9e43a1329c332d6a65eca0ac623
zf5d1ccf6e4425c6e013a6cc48625bd26dc2841054951e589993248b6c7e1dd6cb3d665e15fae1c
z9bb157431cef73e3807972359bbdbc6beed3546058bb22dc3b73e6ceca61b1fde5a5093c47d1e4
z30480ac38eff4a9f7af7d4b23465d57784e2094981fe0fca92e50a80c232dbad09f7a6fe3a8c15
z141b6df1fb85c6021a74ff8da819dc3ebb4737d1917038be5b3ede55be8ca68bca86374f99f4e4
z8a67db6ff73ab23306c1f75112ed58dd7efb9538416cd6c288ee48ef7c81536ac5cb100d707ac9
zade684466418a1b4746846a531e2021aff2a09dbf752564bc02c08e377118b279f00eef0e733b5
zcdcf5b9caf287867ac8f78d412b6b6c7363137386f464be92b36fca90ca42fdc0869497e623b83
z6adc832e7dc388562080135c94f92905e8db3e7c1865028caa68d2b80c062261712ec12ffc2054
z491a6a372ae7eabdfd42d94da5ad0d96a006b6248678c7f42b949312f207af03070e8a6eabdb3c
zbea1a1680cd222245891a0c6e147a1fd58fdcd79f043b48755e98b4aca77cceb5df5b48a5678a4
zf82b7f7a32e8b9d6509b0cb68843e02388339a564e15ca2d9a74a664672f6adcd009080e436be0
zdd097187e14ca5ba444911f35c84d95ccff9f09123da3b50fef73500998b3733cb8ba241fce330
z8cfa804fea65867e5008e8ed46c98838e2d35ec7f0fefd3f68b6bc17642d5ac039735f3189c4b1
z64b642595ca2652d5cfca3040726d33fdf6fc2ca561b7e4dd6582938c163d9ec70a1a2349fb9d2
z7c7be74f5bbeacc1cb851995d9980a84fd5212acc3f635b72cda12863189100b66c7e113a54c0b
ze814dbfd5392502ace308eb9b0ad389024fdddb8bdd08b05f03e4a6efb7dd1eec2588bab36c830
z9239ec544588c19e51da093be876ee95f1ad109b42d979136f59781e36ff1ac23c96a8ef0b5b03
z5b30b2770604bf1e548fa6fcc3c6de3983b53fd9130fc2080bdb603b435b48a512d2cbe6776f74
z0b243234319c202a75b60dfdfd38b57307fed7d841a66c6e1d85ec88574b2f53f9ca5208fa9374
z1b020b1f52b35d0f20a9c3fbe4e1d07501646b3c785d5ebc56640b60b86dd728219a1aa21d4c30
z21432d1f60d565029aefae44cb80d2faa02ee1ad2b7e230bb6aaffb21a6199a430c916f1aac3fa
z92b1dc947dda1005ba0b71a349f148896ed32f84da92b5379d250937ce3afb90f39338d96da144
za2df5013533c0a27b2e6132ce6958997e878b9ec73273a88fc23388266108b6ce2a47a561b0dbf
zf9c84239c86587824471e2a966ea26d917f59aeff1b0950f57da4ae47b671284f12f47f804bbf5
zf0def8aa39d55f52e63d3688c7a96056c8cb9b6b046cd4c88edf9b4b1d38741fd906ee47e81723
z2adb2b86840202f53de7a7d910f713eca174cbd1c970ace1488c0c3cee1d7d9ccef6bb421a3776
zb7cc15c7ecbadb3363d731273b1a37a32ce11539c2d6fa5cc715d44f06bee7624173aa683dee1e
zc8c2ab832cd96ef4a5cc6281ce711eabd45c6abcceaa9cce879b6119839503beb866c114f32afc
z5184ff7507308aed8f28d83e34a2d7bbadeb20ac8f6df7699fbba2b85b69e72f65716a77361c45
z6c14494a080823940587dd690b5107aa54a9f0e8202c99c7557b8869cb4b633fb3e1ac394da9f7
zed8103924f4348caed178d7abaf8376372a6298db5e55abc965f230c278d11bb92af7ddfc5b639
z61033184
`end_protected_0in
`else
`ifdef MODEL_TECH
`include "qvl_assert_together_assertions.mti.svp"
`endif // MODEL_TECH
`endif // encrypted_0in
