`ifdef encrypted_0in
`protected_0in
ze74c34e226135848fe16db9ffd31815111b6d7fb642c521a3f628cf6da949865580b22efd062a7
ze90adae0e65e66a2c36a587d0a790699161455169ed55a01f2084f11770a774ec4c588039b380f
z6de9c5084882a40b79a175f5c2114b2b6d78b070cb806e1c0aa9258297f4687ab308bc470f0040
zb0b1de382961eeeaf2e279e1462520fc31c119af8f2b214846f56c2b3cd2eadbe4099496abff18
z15cec83ec4a77b868344aa20ba7360908f5c0de2a79abf8b3534b883bb12180f68b5d4beb444cf
z3fba8f13afb0abfe8fcc4294810f75afe452434d2d0f1166236c82f76edf1e12979f04bc35693e
z32ae028996dd85737a8f5adc1ebb94f39c940246e887647b64782cd7ab429b0544c173176cede7
z01dfb26b1f73408344a52b7e1f117f12bb9c8077b34876c2e6fdc085981637012dc9754765e1a9
zc512ce062e0b8fb16a214591f5c81e1353b900a611fe1f4886b57940b41b7f2ce99a7b84b04b90
z916f717e73bd10589c81e207ed77ec660a8cbed5b487fa50acde1b055c8870bd8676023f21ddcf
z9c98cc47cfa2d654ff1365d1f45035a045a66c5dfa827905026201628cee5aae21fb892db766c4
zb5b1406e11aebfd6dfacc9da5ec03b70c276807a3eb15e28ec7ab1dddec42388b9424ea285623a
z248195c9f894b36317ca6e59c86f11031163f5f52d70922c037057ec3eba50b955600900b32628
zb2250f2b4fb3ed6db7d81b8ca05e994209e236669db511df2c321dadeee74880d12dbd5092819e
z312f2e640fed00f965c7b0e1d2007d987dd08e1042332719768f689f95a8ecae54578598cd4014
zf52c9aa29e5602a0a7c0b59ee67317c72101e7d1c45c07570c0683c158486b6e3157427e0a2514
za97901c629a01f6fd65b5a7f6f7538b7ab683549194b5767ec9f9eb38f388669f93633863ba210
zd15b4f9d05bd96c35341c02c93752c2344db76edf8c697562b3a09dd9e6ea71115a107694a03bd
z48c4beb95a5fdace643d8acd8693678fb3c10dbc716d343185d0f8c8b090128427948cc61f654b
zd79e08af23d1f841dbaa5dc1936e4660e1f04efc36d203629f18a16a4829e3b3126751fa196d42
zfab93a2769d0d4af5366799eff9987e0ad2be0898f05a8a7fe7be72a09e6e962114c35e028f985
zb4f3db4d71c39b999c96003b9bf32fb342a15fac3c4446676fc11b463a9620113254265646ecae
z71d7cf3381b7e84b560f223855b0b20038eec96c1ac4f1af8cb0110cfe327c79fcdd2413920852
z093eec9cf19ae3cd8a67022d07fcd7bc14320c1ce4d9db0e528514c98a62b5d3ec31605cf03599
z4d6eb850c37fec85cf69e6b474e171d53ee2bef5d245d9cea5c101e34ebfcfa73468705933e98b
z1a22aa5b32d9f8d3412392ed7416ae93ef2762a663e61a210309cb52001dcd4a952d8799718756
z65c1db60a4531864be9bdeff4cefb56beffe2bf29fc5f3345b63d7f8ab90e88a20287661fd01eb
z5e716c090119d5d4c08ccdcf8d33e906a8990d677657f34d4716cdbd43f372c20c4a03b754b7fc
zd09a688dec478294aa8052d341050720e84add185bba28dced0c27c13f7c8c7cf2b793b02369da
z080bf6eff0124e7ffd1e395669b8e0fab00d0bfbdb7b4de8907980f17ccc6a990eab828e203546
zc08cabef41d95483de759263a68379bc58694349f4d092ce1c8cbc4d8b1cf9a2a993a7ff3c5dcc
z09f2675b286e7c0bdacfc3510345f25f7fb48b7e6c7f9ce1da3d69c5c34d4db08c56127a25342d
z438ebc9b0fc4b41f387865b25eca0c1c664f5ee46d631b1a7b4d9f584843a2492f0e6a4375f36a
zd408f01e8d60caa0c7ece9914b89550d320296303dddb38ebdcb4c0e7f0efc8acda6e6b587210e
z71b5deece77038173722b7fc945257e2139de2f2dcbf3aadc1d4275bbdb85bcb926eb21d7915d3
zb4505e7608d3cacfd452b687a6788d931c6fee286ac5d74f5c9f498cc7bf8e2d6a6fa197c9f1be
zd7a9bd147265b94b25997659e046511eff70d0206dd77b5e79fb7e3597be5514c639de1d19ad0c
z05f2c3f18ba55f3e7c2c8f092141ffb4ee0f913cca02e0bb1f8f8095244c00ebe259e435dc1712
zdc483bff00a38f281dcf7256310edd6ad95ddbb1c63d82d04456f834dfce146c520a936516a50f
z29a39addeb72adaf9354cedd5aee8b848376fcf1e0930ff8e2955d5b97eac946abef96dfc634c0
z6d65c11e15339bff5a665cced0fff422a2050eb221291d0a204f573861634a82d46ebb13a2e7cd
z54a1d8766affe05b30f533b4430aa6b644138bada310d7e9324ed7ef40e05343d0133ff335b54f
zd0d1c9cf7af527f1fbc9ab345761975776946876b9996acf2b0a5dc1c7ef3a01b979d3c8335fd4
zcf1e2afa4711a10ea38eb5070315628df9f656a8facdea3cc8fd85bf05f0efba585907a683e2fb
z271f5adac55b7d0cbf1f923dc6d77da4ac065b2384eeb11fcbe4e9c4e286b3e0c8397c9338f4f0
zca5cb05d0221de519ac2cdbdf7c08e1a0d16dad14ae8e380d9909c159557fb377b8fce383efad4
z45ffde49c2a441c977ad7fa3d21d5968c4f3a81a3e92e97006f07e017bf15a9ce2ea866c3a1266
z726f8bb7dc1de780ca7405debe14b37ee80aba4e7b76374f984cadaaed3580ce6baa3b3cb72960
zbe04c1b7c04cff28aff46f7e3f9b9bcf091f352d657f97c0a6ebbaa0a3a3001ac19742a265e178
zaceed05f28ee4a98d5b7ca9524c364f47bf2ee066fa1c7b24bd3f92a37fc7bf54d05e1135d49b8
z5ae86802077f20b120dee2b5f8b0ebcfc182c8e312ccfeb7c5565e05e0d92e9b004e270557636c
z0eaa4af7fdf69fdd97f4e917e9286879d6a905abc5d3189863e716f36baee1e21373197d14934f
z200239586e40591852f3643e60624677f80b662e95948a9a41e900d5f6c23f565dfe90df61c04a
z0f7d290023a9543e70690da44322df955e5018cd25caedc3f54092054eeafeec2cc984c8520e86
z6145286c957ce85aa0acd996cf7e5d5af3357059038ffaf73fbca44d913ea5f60761be04bab3c9
z2478e767e0241bda4cee164052e43967c4534469f54063e9bca3b2811d694dc45ca7dbd9937e6a
z773c817a1b807133773e5db0d2f32e689321d06d57ed5a963dc83e3a30211b3cc8f052fc82629f
z119b3a5c9feea68b4363f0f5bfe3725d9c528b2e9ad558a81a9e43ba75ba67931311ed351921ae
z38cb0fda266ca34c98305f40d92421b393f8fe7658cc3684827c0197d88a62e7aea055ecba909d
z93f23d1cd6513ad88c54c83fe93b13bf48352a644055b0115da01c5ba6a14c482bf8d8fcd7b35b
zae4ca8396c69ebe6e229164108d506e0632556aedebc0256e06b028bf00dd9a70dce66c48acf25
zb5451026d6249962f13a15f4a1c215a4f24bd044fc1924dd04f5fc5a7a86b8fc01103fba9e9f17
z5a4b7d916bb85b5bcf91fe3f255906acdac8cb1860eb79ff5032983a578f89a934027ad5e4a03c
za0d64470b622084a0de73abe83adfb0d2e4b41cb5d929de63cf88e7175bc14aaf7bb3abcd35935
z92d1ff6e72e6a77c13b3b2934202d1dc5a371c42c2426645f2c5920af881ff7ca22c0e95d135de
z70c0a78b99b03829ea8edf2e441514347de79056a1b64d02529d6bb1119b515d321b58e739eb1c
z79e74828cf8e2a5379ed097e60e4259b854c2bf84f5af00eb38b920c2623885a57ae81182a602e
z78467b72725a4a106a09a53bd6cf4b69d7b3cea9406d35103b52319b1a26e2cf21b2c2b4321302
zf845a8dd882acc1edc800f7e3e8eb094e9ee738e95fd8fefdf7e58e0509aa6b95c4058c5056748
zc2d1d30f7defff1e4c88aea9dbf058bd92a8d2784050cb4bcb54b881566dfeef527d45154810f0
zcb6498ef5eb60dadd09047339b2bcf92f1b319cb663b708ce0229f187bdcf988c166ec3c72d3e2
ze7eba3d158c68f7fb02ed169d75bd2620e3ccaec149b03f6ed11d192671affcc6b40511bd2ffd3
zf2ee0900091e62d9cf1592b830f40ddbde28a928b1c483f6f9a52b9c3dab361e30aa7311606c36
z808e436d7e7a968e5756ee057eb22c8e2c00c96323a67e8a8e8a2204d5ee369edba6e62286add1
z3f485bfa08d555f9a0f19ae9ed796847f76ac09181af9bdc18835c13c5cad793bda219832ad956
zc64c22d20cf88fd9bb905083011610b8d2b97910ba9eb2c37a73f546e04cd872d3092e4b301bd9
z2b659e124e6144acb1d75c1f8c9a06b5254ecfd9ca898681b502ad6c28c3f39dad1e6afb8afded
z76bf60679879d0519fd3074134254c59eab676eafb0c7fae1713d07996eb58a73058ede0181190
z124b68b7adbaed52348dd24e48e74cf6441ff004f50abcb25b17ca3af2a45d6cf9e84bc3081e0e
za4112a64b02b2fc67026f7843271a401be3663a045f57f151cb528fb20be9986e68c771edf09bf
z1022ed17cef9197b82ec780f87eb2bd677db2efce79a61a6c8515fd25167cea226541494c26567
zad1b87cd50c89fe35f95db2fec6749426580ebc054ca76a8951a8d35339aa4038a1c7c45abe63d
z6dcd95286b0d8b597c2fe08020f10963a518110af9b3c553aed3e16fd6a04b3493ac25b4dc2870
zee37c992953bdc7a72aa3e164622f4f0b4e0398efbb7109010e02330d0b1a60ba5c32e8b6b29ac
zf148bf37d2b7bf29c7ad7a39bb3589f9adcc41b55080ecc05af85172e61abecc619cb7c2b04fba
zc4bbbe5e6eacb2452a3af7c9ac24c1a21b049b9a68cfc54282777f152a15a0b5a5e66a3272ae59
ze5f5af9af996426238d1e07ef601310d1cd94d3baf7985b5f4843ac075234eee28e5da50e880d4
z1110dc18be5e6393d83ea0fe5858db2deb4bb0022ecf4f56aaf0da9bde7a3762c29d27c4d5a78c
z123b51d2ba5ef358fc46c99a28426bd2d31b19ce236c8eb822a4ec0888440a259b70a0fb16213b
z16dafbbdaabdd02aa7aad0b44498772e72562b453dd7656da6a96a9012d4f82739fdca30c68ca6
zd41f02ed0df11ad470316fb34f8b347824293fc3d9c091152cc02d7153b3dc45cd35000917a18c
z2ee48018df46aa59ec64005a343f3c7258f4c22f49b07321dea4d966a6def7147212c2be0f192d
z9cbb75e1392e4ff063adde20aa3f8787b5ef9fa5cffb2b03e55b6929530a37936841ef7a2e2b9f
za9aee566c5eda2b48073d63c3411f0b958b53a8a1f8cecd1bede7c415bfeb4082e2e4464d9c7e9
z71091921b90309d175f21c2a3bbd6dc8b1fee922493ef8f80de2f2888ebc25fdef6deec7b7c349
z210568912611aed3f7aecb456cb0ed5ac4a91e37e5fda1b7dbfed3bc0b40f3d6f06c887a390154
z97eb62f77f6d61b54d7ae41b7778d7f204853fe8e089b83ea420f8d8186f1f5dddb4561b1ec303
zd34f256ac3e67ca9b76bddb7353decd2d13980997a3610e41e2343d52e10ab1866e7243a87057a
z6067dc75f1ce66680f746b930bf448c9b067bf8b915d47f4f9d3915a49b13c42df0fb142eaa64c
zd5eb26f2b05161a938241224413315425a11a1e90000379cefc46eeb83811860e6c26b8e7215bd
zb3c153f9abf9fbbeb7b4e3a64f3238c1e4c480a6b382d8f535190a65db1bb227114f4ec2acc78f
zbbb2f26c63950ff43a491374f1e50aa138c12a5ba0de4e79e8c9cea452e0a6ff8fdac33653b5e0
z9a61890192b0a1d79be66b34eeeed898ecee8ae09c53558c7615814ad05e07ba8cdfbd5f76d09a
z4ae6f9eef26c98e7620f765406fa2b9203ddaa699ff313de31b90ab37690582637ed24edca8892
z75935bfb701a14829943d7c9def07f2027d00504e94dc8e63111f3817570e9d53bf29be385364a
zd25c2d6a3f47f7d4db272c772d9bc4e5b0cef6653591e0bf7ce58e9038368334bbb9fbd1501fda
z29902451166f844e29bb1afd4a874dd24d0403db515092b7aca0cbe7dd4cc0c0b7c2a0e32704d8
z265959e14a780410aa2dfaefb8ecee689603cba3b9e4ac3ebeb367b3cbfdb7129e50f1d1b70ebe
z7c44f25c43541f318402480e85fc0a461b07cb8478d2d58a78e6777f230dd2e1ff9c312802202e
z8798c26540cd1c0deeabc3a62fd94097f870e060232e35ba962305536e6dfd0fbba3e8d75f42f1
z164caf8c4dc1b316279d3a0142f1a9b8ea37e0750a8cecb1abd8ec3ab95fa8a81f086d410313f5
zca21c016096a994ad08f7c07b23eea4140bea18010f017153fd9260f572ac582b37dcf3828bbbd
z0ffaf0cd8f4f4c3547da830bcd8da649883c4d8813b7db5d7492342f9aaffd525e9149663cd431
z1cf6191c3b1f23a51ae40a852a38d5cf6ea46a0cea5ac9d4bcf1e00c95b0dce91f7679b1c9a08a
z33128a48932f5dc6d68b48acb903003dc0bbd84e29e2326780b80984cc546f73829b91175db960
zd55283b862576e335d9d6877b173cca561b0717a1922e6482b789ce93b3bbd113e12979167e182
z7ca03c73ccdce96e049a236708317795c8bd529645b2603eb969dc5de780c26e4d55595b3b3c7e
z399a7962080f0811810db5aa0cbd3014c5298c780c34c69d9007ddc398ccac7ae5f92d770a7525
z770da69e83d3c578e740f74b00fadd7e10790d1779e52307f47e38aad600a9d790590b624cb36c
zb10a4f2e9b57025b1da9e680ae0a3f18a0020d62783fe2585869e6b3f57fc3e92635d414ef9389
zddb01e2a8a562b62e082eb530d148b8be38e6372f5ae62b4b1dad1789ca6f9df373f8efae9da6c
zb6243ce139e015f038932929243d2ee8f2dcc7016d44166c8524f9beb71e4156ff9f990e78c4d1
z1b56aa03db243f91faa1b9f35cf1905c3bba8b990a6777b4ad14b46712aabbb6a3d4bde4b52dee
z38afbff02846942f6a8aa960046f26c3034c35cf6fd8d141dc62b2ebf7cbb6749abcb2c3a1dc5f
z6ec1d6f8e89f5f3c25f81d51cbf1274f3e65341b9bf2301698f5dfe8daabeac4d4e9678d86bf4e
zc09cfb928ba328f389eaa4febc1a8607ff671f0ab9a5af1b6dedcbb72488f57a57576c4cb1e817
zdd010d573e2de18fe16171ef50d32721be55b3f25ea779a9a0dc4eb7d9c4375696e47e3fef7c25
z3b9da0b2868c34d78cbfa5567db50fd2d55b43bb2823e7f79074ac2a3e4d8a96196dcb923e27dd
z482f183e2e0c41c154c36db329906153441585dba5bb6d52c169ffa65cf81aae9de0bb4d5ecea2
z5c39525c108d2a7a495780cc365b7394d112aa6adf0035c3c194546fb2b5975cf6ea71654c61b2
ze6c7115edd7cf21aa3109660e99ae1190980846617ec14777892f2342080384a0811a72f9918b2
zc1e888666acb5c677f0724caf05045efdaaac246d949480a7ba3affbb759ffd85aad296388602f
z615d6d39ad375c32143bdd22c5535004d7cb09e08904bceafcfbe7543311bff9bb12db5d479cfa
z06dc19c2c4537f72ea2e62ef5b972ca273777ff97b75080aa1ff3a7729be76d611b245b5f7df51
z27993c11ca0105a254461d27367a830e85cf9d6e63dad20e30b3ab61c82f6ecfd4ba748e523522
z635226cc82749986ea944bb1bfcc6fc3f9978f0515bb94c98409de5e3af2480d530fc9a7060ad9
z45061f716c5dfa64b4c2c533d07263020cc52df902b986765085b1f1da5ce8fac784e6a98d8afa
ze2311c11d8ac91086fb1dedb5d3d6c15288fe7acb7b73652804a04fc7686df5ff6b24470c0eb52
z0bb8deffd5dde01b1349e0316b10ba4265795b55eac938de14f85a96c99ba2fad6a8434b54d317
z3d5b15dab5cea74d448d1a6098708b6f4e48b77b4ef44eb484a8036414e9d44e03413325897320
z5cbac4a6b10c14cf1a2035d6dd5d95f876266cafa255d2568e24cb9e36dd6129363244618a252b
z1b4377eb3ad3fd825e19e73f3233837a33753f28d15ad8ff6137ae69edfbe7b9b059187604347b
zbce30278b4916680e9b532ec1ac703d2c9fbd7b735734b4ba2c32553ed235cf37c59c77bc1b9e0
z64133e72fbfc8d655a5eed04c2374cd537a6ff2055509f1fc9f711a5ae34202677bb5f8a6d4fdf
z6e519b0c6497eb3965f6a4be3072d046310653dc212f9bb361d81a9ffe39d563b3c2fbe3e419a0
z198b660b8f22fe45bf9b9a16f4e37fc0fd937676cedb4933a7f91fb1d9cd076a260fade608d880
z1551809d8be5037f35abb4dc41e558fe91852aec95f91f87627be35eb5de72ef1ced5fec2f58c1
zd300a0cf163c40ad6069dd23e34539bdfb59b94a21c59cb37e4bde8e5b94d64544d4ec7ceab38f
z526fcaa45f33dd41c92bbb61e3518419b823a3db683ac9c82b2961ec3d3f357916be2a300d36f3
z7779f4a6f3fc206093d0a895a92550eb49d52c24f9a1b13f25452130045a7ece6985790c1ef0d1
z6824e5dc9f695260f6d300cb3ecb2ca6dfdebd6e11b67ade1935dc5dca0869e7308d397b067234
z7907e8e72137f088c300bd4f99d475b35dc246c0fe50faab896fa2845147dc0d9f0ae87b6da567
zf97fcacd18d429f9c0c8a1ae140377061c70a48fd1ce436bae77fd0a9b95818fb4606ec0afd34f
za0763d296630564466ddc168a931fcec83f17b11b07b19e54bbaf2b9a40002c89a3b7f5e94b983
zbf1dc5fa1b0f6cd3a17db661073ded5c2bb3d983ec4ddfa833feb021019e808c4c68eb2213a968
z20955fa88f134c914c632a4ce57ed983fad41ab47ef633a9b67fce5168433dbb5ff6cf99d316a6
z57ffe6c5ec31cf0ee07617de6b409f6330bddd29120451c46526e1283a402595fe59a1fd1d8d0e
zb4a3c450156a478fb68467e4006aff2806688ba86f4b08fc1d9fff9f5a4b8325b9e99ca221073d
z93200994ce01245edb658047e5d57349c037c945b4a975fe0e3c0e2cd48a1693e103a13475a451
z23add28b9d7fe6bcf867cdbdfbd5a50f2bb9a2aa8bb75289825e4f5c9a9899bb0e47c90e5c3586
zb5182520f8af998482f58844a5c96ad4ea1f67aab477c4204574ba93588e90a70606bffcd39917
z999eafda755eb9933c16d40233e1026ebf8051e29ac24bb81b18497caf3df739881fca5c00eb80
zf873d8212e3b9b4e989c92dfacad52927602cad607b7fb8d8cbe190ef19a310d6ba15150b2d9ef
z8d1c16c8ceed05c7bbc1d5a47e839581ff80eafc260798d58dc515ab1af862c2958a582bd3b9d5
z38c095b575d3109c3ffbba9c881899c24a6bc5729441accbbc67c2a7cadc766c50cfc73dd2767d
z0d723cda9eaeeae3735c2d4e335a10969556b2dfebe55bf1761f235e11de5ae7bd8f7858ceb011
zcb7ee941f73cd0385bc2886ffde98beb30938ce26326c8c1b58bbd3a8bcf664002010b535b80aa
z0e8da0dc2804468e32ace49da66905da960592889554226ab731264bce3874e3fe3d8817e73091
z3d18472dea0bda6a9fe1394deb4f8f4ad2a1989537f674e8cf59b81ac32b2c54a2e9ecf1171eaa
zc93d082a4e8dcb65683939031c2d7a7f0e04e562c6e6f5bfc897040ddcdfc897a1124e3fc6c142
z30024d9e3cc6ddafc9042538708546070e2c888ae65c4701db96c512924348f3d5862a8a5fd093
z17e87be96002a703d595dd97a0978226f323bf94da6e7e8ffc72a2bc2dbe4abe4789d6dbf85b73
z96342e58fd90d4534ae202cf995e785ff88dab11becaac74d726a82216721f61b6751bce372e2a
z8dad148f313bd8a7376f56c12b973b3ae138e6549ff7c18313a2666ebd71cda4af786c287a81c9
zaa024c5cfaa072a84ab430f42b1732c4f0fc37a4b6fe0f86cb2d23665ab92b6f9cd92d3ca9f4da
zf317ad8da7e110a9aba5a1c663ba4f9a867cd437faf019b7b498c1ed2d1c6ede5c4bb4f97d6f5f
zc1374d6d0540e042bc18cc93885a86363783cc36b8fe7672e2817c83adfc816b7a4e3b3754add5
z46dcbb1fb11b05368bcc79f666c28f06fb264d0e697a038aa9078e3753737a26cf401fe5c48b27
zc1fb167ee1cbe2469abd6255df0c59088ef0fb30404727874184e35becf88211964cd8c0e59a80
z48ad21c86d82cf3d1eea5e6853a4bf593f3d062a364df2b61e04422707145ff75a667432dddd70
z9dd17e6a61457649d3c8513cd24223d3a0b7effc380943a6fd583e48f084894ea4625f11283c81
z2535d64795e18a7b221dee1e485b93538590cd4c627d786e7aeaacb3b16eec8172992621f5303e
za1653d6308e1c8786ec2ab2aefd5574ad6c6fe26fdb6859364d2ba7192968d182cf1185c0739b3
z46b8582b5d0566fce20b7cd53f16c57999dd3b18ef926cb037537ce06e437ddf71c792bd5e043d
z28b046b2c46bcbfda7c89c6f2f074c73ec002f55b6f990abcd54235c7231e2b8a1ae41fee9a26e
z801e6c9e03ef9c04094eae7aed701c86ecabeebe9b39934c806e8a9f9c9594f53c83455b5c1be2
z79209449f6b4cbc39093f3134df810e721e80b8f5f8e75a223b02d9a8b9212fea28cc4f41804a7
z43da40a810d89dc244eb2dc9b3e680f32bcdb015c9800d9cec770b54855a18029d70ae2e78e957
z745624086c1fb72b6ff16a42e26b2ca9a81432acbe22063284d28bac7aa7ca4f76f1ca33c41c76
z8d898e9a88aff954df5d910f804277aef35d7eec3c0a5a825a711015629db8bd220084850e9519
z5bad3c20a04171baa3ed1a68b7465245b889c50f22f6a2bce1276a25ea5aef96f9bd9d32727313
zde409380a108a3a80c6dd2a79b02797806d7f4e8304e99652732e21e1a59b5dac6ba6952960f29
z0dcaed5b10075ee2ab27017aeb2105d8189495eeb5a7a84567b1dd07fb095ce463e843ed53ffbc
z4afbad323c80fb09ddd04d4ae393fb1317778f0768683ce53117e03f2da0397c0ec9552f4b9bdb
z4cfc5614a182ce5b0373798daf57c9d0f1e7d7db8e3a2007036574cfaafa4d0c56ffdef4bb79c2
zddeb935f3aee142fd0799ffceff786def0b2e2ed549119d2345e3b0a1caf87460f4eeaf95a0262
zd37846af3230133e348b54b6d91cea765f04421c25ee828b572f79a88eda0b3ae64a87eb40bc1c
zeddaf4243aa896e1ecb90b3a672a14cffc45146658720022480e3f011bdc0d6eefab9a1059e749
zbfb41354ab72a01364d16db8d7fa628d129241755f32c5c98bbdc080fea61a4b24138c57ff45f1
z8d9d1caa984ed30f3afd69189954dc481e3ce6bbd63cb28497683421a52fa4e07b5983a9156198
zd4749f2a46c4297d5847d8c702e239e339cdf31ca037beb8b9c6aa6b085fba8ca962379606ac7a
z1350fb9d269db4c9b199d14fb07f7e594ca702381c90ad385173869e3291a3b275b309f58be477
z887243643c233570fc8589862d521a766c236e65f91fada713bdab71b449bbf65c103bbe519955
z56c346e1b9bc4e4fcebda3a70dfc87f3659e483813cc1b94ac2384b0d0031c9e0353d4ac1af54a
za6cdb277b09eda11beae529e6c4bc9242f92bf0c605d72be615edc9c025bc2daa2500a201c3e5c
z303c069c488e1cfec4cc206ab3ee430f70e2d700730665069b33b08686c586fc9541bfcb7c21ed
z0065788b5e6c3cb9729c9cb6ddb0afc5fc85c33555455e081f8ec320e9ac7d4a10ea9d8d60db65
ze6e9cf2101e091fcd749626099baee73b93a88815f5a89d06325a1756d997caa32c46ac8087c6d
zbf1cf89b4ce4c25b2111ca31e3f8f5a697900e825874ad4298f0d02671d74475798c9fc0d5d9fd
z4e38a8d87a548616cfe41dcd79bc36017d7a08dc8327db54e9b776ddc1c8c957082c930cc910f7
z97094d1a8863a0e16b0b1495d2c8f56771168338af9969ef806e9fef52b5446929411316e6ad03
z2300f212b0b08f6f9b12824efbd048254725f182b1b825155c185efa1e9bd6026a68b08e637ec9
z6c841bfcb3019cf29605d02bd79abe12aea37afc7a08987083e6820b44fb050cce58e66cb87925
zdff0a01c0a735d7b9e1b070bb7767d7172b05870d74306ce65d03f34f2a2d266fedb80637ef0c4
ze712ed76b295b39aafd5ef0775f884d0701f78194ced9945f40d53f74d5e31b5d42fdf960ce711
zbbfada87e85a4ef4821cbfdfc046a99fd28757386d3b3902f71f93bf4b70331a4afb96209b3c19
zab0ca56ff7c57c09bc5ad5777a6fb9cea2c66334406b0a9241c1af450ef3a3427e80e793d3d06a
z7cd202ec707c09eadc95e719142d1eed30386e98bc9984e50090ada079c7399ad52e95f3425703
z4b71c9a87d6aa22387095945d137c95ae3906934ad96642438df7678f6f0b9a3d5df817ed88002
zae5e5bb3ae1c4c655d2cd0b10d347fe7b4b9cc9795c902424dd120f90555637d416fda43f5e8a7
z815eb00b6ed2914c37b57b33deb10c4aa0737c77946469a6ca52b2a51215f0ac0fb5b802d61ed9
z75379d8803dd04566a25b1e7e647f98723c87a1af5b566618d45d806ec74874b80ff71ee3e9155
z79a93b5a4f822c679329df0a7f3f84933be1ed99c0e7e6cb4a92ff8d78fe60d0001653b03481b0
z0ee04ab9f038f43280e2b58f74ac4d167ee17deef20c81169e7e3e55da580d74ce4db5c674a468
za442ecdda75d086a9109acc2003cb963e478a736813be7ed5c1c975412382d746a43b38f9969bd
z23950f6bd3cfcab411b5ab88da0b3502d9c42f9643461829cd4fded2e2098bbd0972bbdac4cf00
zf4728fd5123aedda6de2b7a90781e64b5a5a628c70faa117a032c21502481cfdb8acaf54345d43
z70251cef018f005c82b1004502c61c017fad0e9e3e7612b97059780f38b849ae649f698276c14c
z5972a453336029f70d08468d6376f0dcf299508a6ff42a94dd01f0af24fc043724ae4410b5971f
z0dbd5c8bec7d7b322f2930efce6de377094fbc85eb6ee21d712016eab332792ba1c2b036862f22
zb9a167489b17414971b7b80cba9e48c8e49af3964230586bec912442f0ba04db03b2d77c90d6ac
z3c820d9abcf84cf45643e1038ce638a89786856d9b9225facc670c82dd53407edfef1e7cd00cf0
z4684e686ff48943979ba3f3e418dcac812d39f0de55330bd7f5d8791bd2babfde00fbd958105c2
z5af5b15e41252c0341d1aecf289d7a85e9a134d90f42c2dde46f9e708bfa9c132c39dffcdb721a
z3bcbd3dea9897ae019cbad25682567ca80b0bd908488f293b8916835a8178dc444eadbb94515aa
z916c8a636c7d69f2527b8e1c85f3e1e25036c0e525588489e01011347ad729340ac71b697b819a
z19bda71104eb5ef90f15811592f2a8f4075b4ba952f0e81b659e70278f74c27d83ac492f992f7b
ze99492616eff971735d704b23060ef58aa4e96df13588f3fe858038e33f7220eeb92f02a3da5e3
zfd66f0ce7351783911a23839be8d45c99d969f3cb92314c7772f804ae060c313ed06f340caf0a3
zf645536ababbaea18ed5c3ac5d7d76fc2bbef904e9cb8ecc6e58c091078966ba6c98b6d14d4c6e
z919184eae1d4b6bd114ab706729f8e2bededa24406f9382288f964f2a6945de4cf21fff7b62d6c
z3e240bda66ea0d235654f95b3f24a894735aca12a1c45cb54f34fd6ae14c4b2f50a2ba0ab0c18b
z490a41a015f8c1c982dc1139ecbec24dfd6264d91033f3dac4ca896bb0ad838e1c59181c835f3c
zd31b76a4af5bc02fe683c606a6667e57b0e71b9ff2b8df1b19223f7f4141f5aeedf73ab28f3846
z15b543bf42d2045bb2b4c6adfec61c1647f33f181db898e462da75f1963db96e2d5f5180fa2da7
zf202d034011409ef011dc8c125f0a9a6aa0873b5044b31012b3576a33524cebc21a0452153
`end_protected_0in
`else
`ifdef MODEL_TECH
`include "qvl_i2c_slave_monitor.mti.svp"
`endif // MODEL_TECH
`endif // encrypted_0in
