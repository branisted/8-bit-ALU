`ifdef encrypted_0in
`protected_0in
ze74c34e226135848fe16db9ffd31815111b6d7fb642c521a3f628cf6da949865580b22efd062a7
ze90adae0e65e66a2c36a587d0a790699161455169ed55a01f2084f11770a774ec4c588039b380f
z6de9c5084882a40b79a175f5c2114b2b6d78b070cb806e1c0aa9258297f4687ab308bc470f0040
zb0b1de382961eeeaf2e279e1462520fc31c119af8f2b214846f56c2b3cd2eadbe4099496abff18
z15cec83ec4a77b868344aa20ba7360908f5c0de2a79abf8b3534b883bb12180f68b5d4beb444cf
z3fba8f13afb0abfe8fcc4294810f75afe452434d2d0f1166236c82f76edf1e12979f04bc35693e
z32ae028996dd85737a8f5adc1ebb94f39c940246e887647b64782cd7ab429b0544c173176cede7
z01dfb26b1f73408344a52b7e1f117f12bb9c8077b34876c2e6fdc085981637012dc9754765e1a9
zc512ce062e0b8fb16a214591f5c81e1353b900a611fe1f4886b57940b41b7f2ce99a7b84b04b90
z916f717e73bd10589c81e207ed77ec660a8cbed5b487fa50acde1b055c8870bd8676023f21ddcf
z9c98cc47cfa2d654ff1365d1f45035a045a66c5dfa82790502623b57a3af03bf0f0c0d35b51558
zb8b5f2d29acf03737a9ca2a053b7a8f06800d50b465c41b30eb585f62f3d0c2c5a43bc3787152b
zb805730de3316985848c26d87c44af9a794398f1795bd9da2c28340a68741f8d884b83d4e6886b
zec146fe538fec787c36679503d6f9db2bb7c583cec391cdb97277cf1cc1e3933b8105542f2d4ee
z0a416155017e2b77f6d5de8301c6235e763ed7c1ba8551768c422d2829fcb4a87babadc6a6fdff
z0ce6ad846db8e40ab84491c1ba576e63e070f5b22606a1d03093a6c4a0873e490cf0000ee99e5a
z62ec0ed4ceb548b7ee261e1de33608c752b4eb896fb3368ef711d0022dbca4f5fda5ddc6c23c02
z81eca2faa1dcab6fc65692a9dae611c6b3206abcfd5da9237d01258a78fcdf7619ea63d3fb1c01
z807a74bff5577b0fad03e9196a849616c17d6670376d2f0768f573aefcbfa0b43ae90f39d28c89
zd07b2f3c13f5b483a13d3dbdc93502c66ea6d44eb0c8588e24be9ab25a95da025e2fe5fff8d04c
z896bed381d30d532b98ef423b33dce53c1b98f7f101c8729ea9eb519dc93811a02dce6f33079b6
z327c10abb00d083b0c37c2fe7e57431efb284cc808199446059eb1efdf2cbcf4dbc1a3e9353e88
z8bf0132cee6e7e52372ccc65cf5cd5a55b7062ecbec2ce7a819c7c76ee2270b413c808eaea237c
zcfe4bbe0f18eb3680cd810cf5996c9495f62d4acd608f2bd9f4eebedb460601d136072e13daab2
z89b59d9b953de7c970a3cff3fb68d007db50217b2c737eb77ec2168720a21fbb67c692d8df7c79
zd9c91f292eaba4bf8fe141fe5edcb990609ed34763ec928c8405f57e1dd5a39a6a3eac77d3dd8b
zb582187dec7c4b9813225419aad53f885e4308b07df8618756ce893ebae340f696b803bd413326
z81779ffdc8761a2a4c2ac2f96961587b12c6cd85e74f2a961be7cabd206b1e61091c00eb451661
z5269689a24184501c4fb5bb323604c03321a3058ec1238c9e0f4524fcdcc31839a1d043cfe11ca
z6ff541110cae56d33151ec383de739bf0415356bf65bb069414ea474bb8ad00966d915d3e3b00c
z946361b3191019b33bd750cf67e625e9e51c7464b612c40560a911f4266bc2fb44f351f17e8c76
z81c05e591ae44bedf52ae083ee023108d5466021916e350160330e93f393359a26832ace56ab28
z18e6c7b3433cf41a02d6fa3f7dc6bc019fccd321ba600b3c170ed6278bd0f21c3ea01388879a39
z27fa4b7671c1ba33f81d7382611282a6ec70574380b6bbaec60e652814ec4923c18c1e1477aaa5
z7180e0c9491487dadfd41f4bf45d293bdd499ba30c9a977eb87021abb4a67646034b0d4e258060
z5fb195ce83685c4b8a89cb1e59aaf117aafd7466e61d59c62fb4a65b101f15080d4536dbc45b89
ze72181b0786f23c80f0c82bdc52428e03b99b1b6ba4ba063d20b5abaf4bc901fb35f371d6f6fe2
z7194345d237f7aa27e5e621f05b5c2cd1b88f57edff48564d8f8316a49b90cc98468b689f06147
zc9fb092e6ac1df12df8d7c722556321f6fe2460a5ca81195db4b7b66eb70fe7c65b3d9a2346e72
z38a397688701adaba0d3ba834d7b6eeba5d9a1238bf6fc5a731564e37e4293e7b3432d51d7416a
zbac4653e4b4818a85f70f753e8034d94de265bcaeaf15351c6f5f9361aa54df7314a4fb3aa2e90
z7c323fd8121b47ef61c5a578c0bfb2b241c531395faebb319e526b12be887ebe42bbba06a6a1cb
z6f68a8dbdb089e66b925a37ed47f839838b422845b6583a7016c34db32e8d9394f5412c5741ad3
z1bad9f365a818154232aab3878b5d251d191e15c153b6b4f06024e27bade03a52993f3a75e606c
ze36db598283428f45ac446487923fb631c4c7f7526b55470826d9104bee84da4faa404b586f79b
zb87ed0fe7a535b44ed435bd2382e142282540f1d2614112052c03065f03e9a4dabdf8b1befe559
zeb281ddaf44fff5a6f38d0220887eb3c8cd523ffff34a644b408c95b118593ac2e164ad2d441e7
ze770fe82fac2fac48ba7297395ae06f2f4a1179761681abc8b6a7c84fa9061039c20964ef9a30f
zd1a89208a4934dff7922de939f43d796e806cb82fe8f4fa27c34ac42031727a208775c9474aa84
z0df0fc53065983473d0d6aef3af938d4d221c54374570a0e73a777631718587f27ed17bc46afc6
z891a0a8cfae3f58444e9614fce2e0970e65fff0c6d1a19253ac95ed593b1050d056aaaf9928269
z8c77845078cd5c144624108b4603e4b3c40a7a5b2ddc8c3ac65246e126eb564699637839f0095e
zd4ed527b2edeeb322c18d1f29f2881f3538434c46b0c1a40fcf77d012603fc8bd219630a308a5c
z28b2f2e8d4402aaad162820fde3991833fd0c62100f5788d8d528ee9a477b5bc4b56ad8ce3f78f
zff5e287d5d8d0b51482067d63f69af28a976d666851945b9c0e4eff553832aa88f9c372af220d4
z5ce770a62930baae5e27ee349b878183aac11caf8bf8331ab974bec73785a57fbfea8a1b5d6522
z0eed6061829e3ccd24a3495190e02f1713062bb81ca4b043359d9548a3cee9a18080099a240640
z3ea204c73d3c7a54de3f41187292089583782e5f9c257e36bae55ac09c912aeb2ec9ac2e5278c1
z0f5dcd08396bc6a018f2e818a3edccab5fa3ed976c265195c743ef3ec85e13cd61f890f4ca4827
z22e5052da6b59942fd11a760359ff28c8629935f5c78dba572eeaa50688a5353e6a93250edd0f5
za273b83261065bcce604aca08d9679b8e54c86250d929c518278caab7f005a4b4597f6b10ff20e
zc77c7e99910e2a89b426c35d6bdc65fc7af9f397e14af30d011be1ff3d356389b15f87419ad15b
z3a47f5a413eafeacef2adbe205401a2e6e19d23baf3fcdc55f3724aa4c815d5dde06c2489cb7fe
z67f22914a089dafd98159b0aeecdeff585d0d7977fbcb720338d4a333243090ec6c6e9d7a6e948
z64ce917361758ab8f9c76d472d9ddb1af5b8dbecfb8f1c5a0c1f93d9798c0e9ed6e4828bc87d19
za8fc258670e8d6080ab24c0a379b0b66f382eb3138cc81b2421c5fef2c71ac69fc6bc92da46479
z9aa776ff051fa99fa7fc2d91a079d38fab6f9467712636725c9fccd0897ee930ee67f9db0780d8
z5d7505419963e4bd7b06e8c66d463de06655b140ffdcf4461bab645be56a16fff668ccc716e2fa
z14538b1a4033ba0066e57d3b8de1875b27a084bad1feea2bd5d627972b68e8da4bd1e824288b5e
z7688fb3720e8ea732c9ee7aec649da0ef829f4c03e18771299694b849dc4aa97cae967141eb485
z595a3c155961f38ce3438fade041e3a0dde2941290e3a50ef310c5a89c8001c60a3eb9aa36926b
z0a22ba6a92797e708828c4609cdd57db0b5b07204ed1b668186c36f383e527959a4dcc15045013
zbc6e634abb6c8f27398dccfefe1e3311630a739a44c11ec09bb558d40ffdf9e64270c29d59ef91
z7e80c5f18ce35ba705c91c39391c734a59845e7536ece874ec0b178adafd3300d97f0e71828f18
zeebcbebabe9e8fbc93868e9c1919b9a16ab6b3d9b91b881f47bce6f7fa32642bd5ff0e07f579f6
z108a2a49d295e05ae843779c5e19dd2ff4f938ca5a8a04db46e862e681724be683352e8848b276
zf4586dcdca0a528e2ed3ac1c20625c18589a40d63faa3593e0077d3ada2c86f3279f759c35890c
zdd5a9bc8548854f482ba373fbfa0c8ae10e420b5f46f61b1f1c9eb80474636b051cc3ce41f4210
z3c2e16d5c3ced8d9c0527e377265c88c210ab30c4dda548102d3fa2319bdbf9de00f690752e3ed
zeebf54b5cffaa8ecfb53ec98158753b5436fa449897ad2d244921d75c23008e740555964607acf
za1764c4a065d821375a39bb3804e00729adb474d0f445995e6903d2f0009c65b38fe65a16d6fcb
ze09c3ed66cd5d8c05cfd825f126fa747005e6f5c2f68dece3a87bf3bd84aa753a9d57fc105cf76
z1fda7d59e392158ec37f4bf5cbe3ab9ded28527e464499820772b0b0cb04bcca623c8faf470d01
ze3f860448204ce807c2b28c9d134a9e79d1c4a6d80d40f247c6a59b85d1003ce55c0ededbdd685
zcf71d7140749e0f26685eca51c60109cbb284b57e3a681433f1071117b58cf40cf014d81f38352
z507e8ede73ac174fc4aa10e7ef300cc087fe131636a9da0b252f9c8f50f65505a343f34ed1c5e1
zbe763293678ccce4d7dd391b5e1f0f76b726a037d1b9b48ac9faf23c0a7925d9ddd8f34f44d808
zbe96d20a20f3402d0143c1bafc0f868e6b10998fb2639d74e9152c232ca14d3eac347aa577025c
zc546344d3ab987e709aa490d024dc3093bb9c09dd1350d1fa29b874c140331e836d4ff258074e5
z21ecab70c22b1aa6e6bb7239a4eddbc1f061d776670daa6f9d2da48856a48565375f0990556a7b
z245f7327b3252ff469ff5ae139a35410673706c35a28ff45328e85b05fe0cd6386f96d2915ff84
z1a75822134fbfce892e83d6c9dad3965aff9c8a14d95373d0f10e153a278e3e6a5e21ce4b4c6a3
z8525e2d2b5b852cbcd98fcc7c383bc3334181ecb3e3cfac6254dc2972769affe708a3f7684817a
zb34ee2b284ea4bc8994bf26dfe1b08a284bad72716a173e93ed2a16239d2b56251280b37ac7ce3
ze637acca683c9c8db57c3f4a5f46f6bf60d040d4e93fb51fce1a2cc6c137ce0fc85850cec8329d
z2b5742551ace29e1720100e0fd96772afc344b75c281ea285e7293187102f38df71ed4bcf5e24a
zcd2711330d2afbf2a64cef187dd1eab8c91657a853ed04aa7042e0cc67abd47aae8df515f3ed8c
z8e8b05984429ed28c783bce6378de395a91eceff4df368fe679e0f3c63c9aee07ac93ec62f0753
z8e9ba0e934a3b0a37c0cb5bb6bc095d4d316b48394c629e7cc87bc08edea9d5700959f800e307f
z4ca37c81b4505e24db10949acddbfcf6982dd32051fd4b99e08f62af9aa9382a0a84ebabbb101e
z39e6da4346951d0b0162ef5721575ac46571da42ca112f940c1ebd2c5c3354283590a209787b20
zfaa84b7d918742bbc1ec7684d0c0adf71f05b32fa29920a9901c007b2a8e6ec58cafc261f0f006
z24b180505fd5eb2bcf218e7938d3705401cbf26bf82651d6560763bb642e261b4915dfa4481686
z9481882830bdef2bf620cec54168eab44c921fcd052f19dc90234c39fe80ad84f2fd8bae6ece15
zf6cc9c316fb37d7b5f2fe5eaf696a17933d711a6de9c5c2b022a494a81dc8757aa4fceed6f5f8b
zaaa670004af4b8135a01558a09acf07effeab85be41eee8eaa17e7d859ee1bfd752ec222987987
z43d1968134e8f8dc25f830a9cb9a17cedc09a01a9e243219309af8fb2f2e3b0a7a4c44352b81da
z3e6a9d734c868238fc6bc0ebf92dd6a0a3f589aee4d4c8fe9159eec97861864dedca15045ac0fa
zc2d32b98c9612acb525bbb2c1de11a0fb1bc931a039ebd19d7de7c92ed838fa2b624a4579a1bc6
z76dbd0175251da15030f5907a58028c2554742dc80611aebac0d368274e9ccb683f615f1da3db7
z8e620ce11e279b1d7b8c02b6cb62983cc18a056ce58542b65d38701a128c674eebae740e7f2563
zc8137360493a816e90c32370f8d583f4f27aff5efcb85ba34c45270059067ec9d1ccf3827ea181
z7ce3f6c7d46a63f371c2f964e577bb6280a1997d3b113cc939cb3b1eef922f241691e8aa7e2990
z4f1660c2f398786a50f08c483573cb79979e3ce3312938ea4e35e0091bc82748515466e9dae5f1
z3483d3586209a1add5a30ee8d3fab81b6bb483005ec0e70220bb7e736d816941278bb1738dd622
zd9e85cfd0926070f9eb9ed896f5d55dbf5f166227fa969c8e1b381523e8a2416a17b63fa03e37a
z113e30b609dbc516c32671b7cd552c933eba2366f13091c7a517f7c31a8960ce8e85475f691a0c
z0b01d0a78ef82af1f50ae834db86b928cb79529c086015a7a608f360a6cc4d1e305435130c966a
z6245671a3ee54e263f29fdb881e6fcec79db81f3de2123eb27e042a059aee9022bdbd315feea82
z8303a926765ccbfb81745318d9fd26cc62dfbff74c70354f6dbf460ad215420e08312fb8950d44
z50612a647b68b00d4b0f6b21565a212c8a367ecf97abea44da6accd1a049f8c6db343edfa5af75
zdb9a5e535ed35a3bb15a5507ef244c4d46cff20a89992df66a880d6ab5b429f3a35a46de9ee4f2
zbfdafd501323a5469ee047bd6dd6032346ad3beeda8e7e03da7114f32903dba38aa584536e6868
zfd644f993b1678468aa87c7aefec172745fb86525dc6cc620970a62ceb704520065b1a229261ce
zca4a4b3f3f0836cf4f57559a6d1c02451894bcd7476545a1222ac915a7116190e2466d5fd75b13
z5c63f2433e83703686d4c994eba5fd92d5c4b1c34d1579b100ccf4a6383670d484388145220f82
z3f8a38043df2796cd9f6e9d4ae30f22c3753e49e912c774343fa2041dae62cc8625199f478838a
z6d984fed5d1c7c2170e2f1fc40a653f7d07e1eed853ef86bc7bac3f773eb6956fdae6f6b360ee2
z44e541e039b14ab2b243b72e36f2ebc5e7486179ca2ba8d61169750a18bb6e926da1a340a3af24
z2bd7586aeebf847e3f46bc42e78fee0432f60d0826cd29c1c32ce2fa4edee4f5460bace4e687cd
zdc28d31dbf6f2a5b826d2752e79861d16d9d44b84e845e9d543418707f14d5d4f7da25ffbdf330
zbffa11a10c7c2d06b7843addc8e836421ce6c81c5226a22843a7aa410b88639e3db1f206b5913c
za8ea01c2962cb9ea4eae9ba70e4f84f3c2947e9e2001c327694cb8a1cfccd8aa12952702046612
z292758780f9d0d4cc4f799a728009313eae30d23abc5c59e85f6d8c48d4720f9cdd55fc635a2a1
zba7760e4aa03a0d86340dcff0fe982e2784a75e8dc7ca145631029ab4882313dfb1993fa3ec35c
z52d79bfb1c639ee941f0d0e33b5af7c6c8b56aac7a07683301c1daa272afe5a8d62fbb5d995459
z6dbcb437b3b894c5fe411473130d00aedf952c2fd4e389375770cb9602ef03b697fadef0cbcbcb
z10ef0684fba2ebcd2ece43492b0e46f4a93073b1c7c31ec819447eee39b227b0a52b7df02e1628
zc78196a7980b77e9dff190807f0b9b76b79218a3ad6ba47de37d1db01b776fbb0a242c1b8b05eb
z93ead5fc76b4115d084632c6086e4687cfb39b7d78d852105fdc573ab019376f980e3d38041a0a
z8cf4ae696b95425ad84e28baa83c8b9fe5d2e5f7df1a97d3338fdd2c4975cda98fda7a554b7631
z7282b58cb93cc2f0f4017cc1fc390633c9cd340498f815ec81b7c6bcadea6492b520b866852798
zc913e68ba99ea384fe30f3af4e2b549b33947b54a9b1611411f2bb49e3f09ae987096c1863cee2
z69faf31428d940904baace96b39621d091d3678b9da8122ba5676c772d34e28ecec97c795cb52b
z969fa4f7f8705557f4ea232c915e94d8d241ea880074776360633819e238e5a78d90d2c0093f56
z66347864122ee6b205b5d505a5490ee74c6addab0a32f7bf17c81f282a83793173c648c4e88e4c
ze4039c80c639e8ff15f727f0e5244a4e5a345f64ac165df09a63f9e9b27ea85899aa75e240d26f
zb71ee1f141d51c7472d31894fe3063747a9087884fac7643295098c11c306aa7b83aa7829d00c8
zd6543683e7d624c67f8e101377fd27bcd48b2630dbb31b8fbcfecdf355203d0048cdc393956eb4
zd8afeca26c92c2e18f54dadc9f3cdc908c53203e5af5bfd8deb440cf9724aebbf70cfd09a69847
z6e161b3f8f3b77f1270143257d67f6f7edfbaf08c54b43e46634450c1cc374d3938fa53318af76
z1ed3b4ad161cfadfe0d9bb6d421ea65a10beca894b8d29919593341d0ad13beaaa2a897480457f
z53a772624103e9138c9b19e2f7612c0d7a0b2cee68daf51d963b21ac41f8a8ff94d970c529530a
zf4c9ecd5f8773a7a37601c8b23c4f87faa0942c6df279cbf259e747bf99afe10824f4b9ffe3aa9
z301f101c3b42af84baf01f300fa6e8605c7882582381f2144fb257cfc650e84af411941b6a2e56
z7c37ee8357438e4c7564e3b820aafbaeafb1baf4a22c457b7cc0b3b21a17a5f7f0cbd215ee9acc
zf3da62326ed051eb89473dd1e15ddf9498dfa8e7eb2da58b5c81d674ffd3708389be554f103084
zd5f520bbb5a69c34b12734230722644300d987622d65878d4cbb0d07abdadc3b5d002f0d706922
zefb56d4b6b4a39c34727a40c69f014a498a7f176952161c7c6efd2c81db13ada784c58e27a604d
zc2ee9bae1c67a44d697480f7f212183d2676f3f8034a8d2a3af8a273ebf65f57d9f16eb47e0b56
z770783b705a2be7af1732f12ac29eba2a5ae2e80b62d1d2c3baf233341259156c88a0e9beeb225
z5b78ab3ef1be226a9fb2c2efba6bc16a6aaaba0f0a42dcd133bac58560fb84e6ed0eca767fc24a
zb8bda3cfb8ca35d57ed86ecad06b50aab8a16e3d4e76652feefeebb91889e735990200a920e867
zbbe1fa0f2f8bbf8223e950b8449bda67e0f71ec1bb1798025b72a2ba9093d36eaf4d3e21395e55
z6eb0664598ec890e38a4892e702418c805d1c9e1ea7df95375ca018665165a9f022b2832955e66
z2af6bd0bca149a8c96593f421910d7ab3672291a828cdb846c79091cd10119f18ce976bc3c7422
z97c9257efede6358fff5c188435abf3f101fa435d7dc66168423d994bd645f5c3df2b155a75ab5
z22c4dd1606afc70c9366489611d0f61ccb140fef9cec3a8cd7455bc5083b15ab803f336f973653
z83665110576a76cfa7305b9e3d33f7b9bb432d50db164a26b7b5ea20db3d725fffea06f05c298f
z6db7e0c229a4fc4189741ed5308d8ce64ca42fa6eada950bd3bde2fafde088295141b0df422fc3
zb752e374784ae8e32cb833f614e6f70345019f57e025bd5d4de8cd28af55483ca9ad35c9ce74fb
z932ef7175c05d359e8e71f5a98370c06ef6338462b2d2e28a643e00aa0e48f4022441347d425ca
z0f838b5dcd498018b2c39160e72a56cad32b55171bc5acdef4770e280472ec568336b9eb1d773c
z00e1f1c2b2614da1b68be6ef01b16d85fa910361dd2c042c90e7831b2e6f697015e8fc0635f098
z05653a2114f8a4a0794e9971ddf135f0a876b82f72a199d5aecedaf76756190da7c2bd9581416f
zd47d86f9636fca819df81261678c12e3f34ce40f99a2aa9769dd007c97b9a7adbc5a8ebf743938
z9d010297a300ba15ac0e3dbdcaa1b16c887ced2db4907b4451759061e9aca7df77528680641791
z6f3ec5dc5cfc055204e709cd168d5bd1db158d3f5895255c55bbb2e60951774dad9bfe0ba5e9b4
z43592ec5d2db39135f520eac3e0cc27a870828a885ca74be7d05675e984fef65b5123f0ad71ba4
zce9ebca7de048e1cf0ff47119e3ee0c8d504860b8466d2f4aeddbc7986861c4893da9c2fb59a61
zc1cb06e6cd4824c5113eb91f2e67f36ddbd3d8618cf4831a6863deda313544dbc76e25e88b6fe8
z0fd87a304cc7ed2c3cb0a1b702141636dfd77280a16ad27b97037cb9e3e3117998febf4e4c3a01
z89e00b88e8a81916563e027ca340840870a129e2a11885af932f781f9dafcf087eab7c7c694e7c
z21166745aeae2801c0d31b3d5ff17f4010220cea43eec285aa5df1203e5d73ca756f4ebfa7cfa4
zee322ca4f2543bcd9b096fae8f82959429e959d00c2059616d7654877c92a9cf674b85585aa026
z00aa645960acc75242940e67eeff8be4c86910024e899c30dbe6074f2bf07a1e7eda49d5be2319
z617b476ef6e77340265abf994eb8e41f8b8706355ace0e75b50f4e39617e11b49b59abea9988cd
z4785d62bfad72e12b1796be663715fedba2ccdbb5f5484d9d6916772e16e1b7e8e81a4258c035c
zdf02cd3fd40e3e34e38e2b0aee7b59dfd56fc0b9124d0824f4472d72dc696d6cca25f09fb4b090
zbdce685798c01e3f94c27a278d0cc275136e6299d8b1ec2413ffe89d0b2e74968bd8c564563971
z2d4f088ca5fc1fcf73e89633bca5a7680da00891b95a56c18bbcbebfcc814ea4d57085fd523a83
z372674cba8a74cba5173796b1505cd9276c747c9fb7a55f4191fb7110b9e09b98b91cbfedfb65d
z9dddbfb0115508bd48d333d84d041cf122278cc55f7303b3f4b58829a36d6810695d4349358eb4
zbca2cf8d4f606bd66d32b1291b4af844c9f311802feae3f2029ab5794fa438cd5fd9b378d1870c
zac933a91fe97d468dcd42701de7f2d95abb2387b95f42056c524a42a055308345bf3514fd49407
z6082236b3076d5a51e86aa08919254932ea1d1721bea091dc08243d9f9037edebaa9c09050c558
z0d146be8aef28b0aa7ce79692a537105bb61228cc0209f6f96a2512f43003f8a93501bd1a8fbf9
z66293dd250e42fcebccd9a06a7ab2e690c4d50cc14e4a9c92321cbb8707f7ebd322ff41be2bb94
z9e04a444d9a4b904c91c6c0b146acb6df153d56193e49c6fc2f39ec49f07f5a6ae0811ddc8f457
zf9e29acd8826c84f9baa4a5ebde09fbf47f528a53a69f31c154ec9484938462e492f6a319298ef
z4fff82edbccf316be103f5e27ac2ac943fad8874bf4aa373b4a710402c76f36b4f034b72e03f27
z302ef19a94d7f94579354739535024846bc963e7bf020b24b4009453736ce2790ee0f90eb9c76a
z3dd79c83500f41a6e0330a8160403b4cf51e303572a1798ff02643be0c6f34db1af55daf5e51c1
z963c0fbadd179cdb4d6c8e0b0b3003e6e147df1f85d8bf92bc2d1d4469e95e206377cc004f00b9
z043a6205b00bad4f56ed47abaf4d77380c516ab08896ac1c1f4c23ad04d355f086bf9b1b273759
z140ef7f88a78e0249f77e66ed6e79e0217f91ba82d10627a7fd40b717f9d66dde723310ce9153d
z7f1d9ff8b622c82b04a4acdabe6a9a8ea8684856ae6a42141dff9626bb3a1cc3d1e4fd9f50d71e
zed036ed16e54e0c6be2ca5a2d92b65c081051aca44b5fa284d0a34fe8449242a890c0b9bcf437b
z3beb57fd495cc5996e24d8216b6902163f7e085f991f28f77c81403e07c193663a9fc2bf89307b
z40a93e7e87372274c4ef215c3fa54aafcbaf65e4c9c8de3a5edebafbc44c27f12069db14eac73f
z5e506d6585d525df90eb7064371eca3431deb65136a2266333dff448238b1737dfd2825dbc74aa
z26bdbad7deb3de2f5d24c91e2bdb40e0a44fa4b6e2812a6267ab4524568b26e510f373da48fffb
za480030eb08c43ec7c7b79a736ea0be3438fd6842dc29c11dcc7e56d8481f054740e6eb9b7f421
zdbc8279eebb9caf226ac8c637b08fe786dff1d37c3a6f831653434b7a52ca9d2dfd09722103365
zdf90fa5c4db638b44247e7377a1b12e836a47a3b93879bea0a4f3f851b4d52601498e6149564af
z1375afb9b56b3bb02eec2449d8d20f7e9581cd0b8d3abcee91aec42acc789c73b1a8f5db098fa6
z2b3c55e118b0959dbc7eaa636e069a95258f05cb27930059c8d449ec9199132fea6a56b83dd5e8
z3b5bd8e1a893b3d9bb672618320624a0aeff6070be2d2d0a3eab07f844415ec8db8c64ce4c12c8
z8b902617b513dc3345b1a79c86e427130d24a6d412fb5db55d52e59d13b07ac354c915a9f99fb3
zeeaf57bf2e12669042383971e34efac31fbaf49b58ae3112779d57ae4a30b7c4917aba8f9c5196
z4d16bd21ad8907d0ce4417e1b74698cf4497344332074459c0ba3ce6cc9cfbb680476d9f29c902
z7dc7e792fed9af04eea66c01fc1f05469d280e62c07955060feabac36b253730ba6d58b56098eb
z90701fbd133b05509aa3f0638868c0e557b9942deb148a8736d95616cf662e697eda66d44b2dc4
z7da5b9ea7588b6f43d235de77332e46f49215d44809837dbaac58e720020e9e2381794de8654ff
z2c55474c7d9a87f15d804f250cddda7b6cb9199dd79db48215568f9da307c0028181dca9096544
z58a502976dc29b657e46708d8dc1da65d9a99d032f00cec14ef0ac9a3b63c90f50e5ffbc91250d
z25c38218aef53517bf82df2a147d076a276bd1dece86bdacb081b531c4be3f1060d5598e46e50a
zfcb921e7d7fb97e2500d6669a2b318178353ad808102457bdf0dc296ba1b89109ca0d2fca0c4e7
z7eebfeae73f1fc5588cf11b0c41281ecd89f799098cdcf39130b8af9608cc040fc9e60a0d77045
z5aec08cae46fe7df655e99ab958447118d9b7584578c4eff2940608e19b5d5e77ab862e26548cb
z13d3c66a0f1dfa3dba34fdb8a4c4d004b2d3988dbaabf50b3d8137a9df7225ee0138ea7c85c078
zc8ffe0679c132e7f1651ef73f52545fe3ba4ae00bc8b8ef9565efd208a5691fde07f398e76e241
zbf41ee3063c1b01177815a1e8af646a3ea866e489205f5072bb86469534b97fda37525965352f0
z8a86eb94864d2ecf9ca33293653c00f01f2d4982172a6f6163d322d0b76d14080d80692cff74cb
zdbce186213f442d00d63785a87bdf8f42345409f5fe7adda9ba6b60e36d8613c6177d751399303
z54f9a1670ea3ef5a72130adbc0968d6d8c54deec10f962a85f18a5b23769321bfc6db2ad90fd70
z5ea74eb60625048a4bafa6e3eb62d0c0a341f02fe283b2fe87401809e2dc5833a8baefe8850901
zd141b673737671bc943b8b0662c84867cb0bd42f76ce86c8e64532f0a27c97c6a188ba92a3f910
z8d727506e8287958b25b52e90efc74564cb909216a10032a9ca6383734ee667055233b76c4b5dd
z907569601fd7ad6907ce00c73fc2fc7712c7906fd50d2e6f363f5c7f52a16f22a5013cc4153515
zf9b3e2d92eeb0a72acba43e836bcf8b9971dee443895e98553b44949ec80993d372b6f57d9224f
z5f11ec1acc9a39dcece7623088dca55075b0743cad21ce27f2591982f34f103ecb2deb79def665
zc5857712975623308cfc06a9ebd82cc6b1aa68434e19a8234cbe10fed6b5fca28a4561ddd64867
z920ba9594a03ea6f1f2e6152c39052c7231c316a21c3e59e82b7b33ec18560a967b2246eb4e3a4
za32ff280c06c394ec0a59a9ec71c3a4f96eb362799c6c143b2aa00f693717f37178631c2c8bcc3
z5c26778f92bcfe30c19036bce415da4d0af3fd4e95ce08b004e140d2fcc10be1e71793606bf847
z540d1400f4601b392420ff15fc484384c0caedfbe933e97d4b721288250681a2ca15785b31ca55
z48407a2b57a4a619f16f07ba5508a603dd655051507019489dacb876b48691edd0b40d45274d7c
zcc38a762cbaa8b18a51920bb849f4a6a78d0e00c9e6eda3c7e08c8f9938915ca3c7e4e10eccc2f
zd65036668cab67037f99cbf590c54bc9364bf3ecdd2d28aa15ffbbbebd00472f4a64db217f7005
zdf8e9ef6649ac2f7ee53bee59eb33100a11c8442731fed62fe06048b98ffc4d5becf40aacbe52d
z36e523abb2c14de652e0ad695bfcc87e27179e576f858ff4f8f085a139821a3f456ad7571a6276
zef81f0ff14c9b6ef378cf2c2304f8ec8935f6c0f58482b3f3f58cfcaa710168f1c2525292dd714
z6ddcc20e766826b1ce84021631a04925fdc44710191a796b049a7ccd4b13c79656276a45268c60
zf6ae589a2da6ff61dbae737fae1b9f1bc24c3f8fa8761ab803ec67c95e0e6a99798dbcf51f6b5a
z922c6e359806aac944071987c2f74eb90bfee877ae828b70c51d2d5929c243cb513b6dbc7f6e1d
z471f3918b45916f40fd2a6b81b5bdd0308864ec9627fb912f9492e2120903a20a38fa7929b42d3
z109cb113be9c344a6454aee2ac86419f61f0f2a5c0f5d1b4faf7494e9c979ac088c467b67d9c83
z6aa0e77ee0706bcb52a9d674dec923f020e545cf3b3265f9c783b55c8453a446798454a45c5f09
z993c30a4415a004acee30f5bbd6b440b5d66027f5ee09d27eecbd899a6db5a4328ccc7782345db
z044277109791c9a00400dd668d1d0a239067e732a19afe4ecad3d5c550cc3b130acdcbcb6bc68d
zfb6672356d34295b4a4eea0bd6042d4ed916adec24521cbf60932122fe7ad99872b5d133d7d51f
z1adc012385227c8a23ee7ee7b5005d5b38dba065b8507f3292b8d0d3d0d3feadb549db3b178cd7
z62d673b143e75ae620c4f846353c8df665d933c986a93fcd8431f6647777d9447759d33879a92f
z0ba680fb53d6ac3ce35f0c1f2112ae41cf898c06136a60a6e9df45456e4e044323c2556df9f3de
z911e40dfd51e88756ff3dc58ea9ea6636c303d84d9be9e27402e2f263739902896688145a2acda
z534e027ff6af8b499c405d55f3d41ed2f0973f73ab159af936017e4703346b26e485fdcb63ef96
zd4a6786e39cfd9dcfaaaa5d7f2fe43cd6a867daf4e1dc84d805d3527d3a3972dea6b87583a0d0b
ze2a2230b9d4c9f7fed9cd72856a173302b5aadff06924021ed3676818eb65a2b3862c46a90c7c4
z7b5efadced2252896686710aa600864e283419ccbf7e1a8442d4a960667f13d52876415ff293b0
z2c1c0af03486c442b108dd29758d6683b7266d1c44915f0aae1cae46e1f8cdad75eeef3eb6edb3
z41251a307c375e596346d217d23e56963ef77e687c2f4be23633a688e29761dfec7372ab50fbac
z33028ffee3ec8b16c8d9e7c1adc27d3bb979720f99135be90a46e3d4a337e6cc9b22f4085c9581
z652a2dccc4669c77b38b6c8ba2c75b3296fb65c4d2889606b8a0c3be7b08588a75a55503f9578f
z38bcec91982e5b1fb7f0bd07aa9be6d0c1642aee770360569c138228b20f7ff9831841bb587e02
za78b827fb67a4e3a926dc423e0f565a2b2d09423638f37f73ed7eb5f1aa385cdd0b74f698d2ff1
z18345a151260ee22df7b8a2e9ef02c9137c03ecbce75a1c39dd0ff99202724b2864ddc7664168c
z626e4c5c9e45b4824657bb91d5551660fd1057ca556427b87f84e53ce112c1f2f4cbc690f8242e
zd0b359c402e81ecca72963a925594827bed8922298ab3a9e52bbbf69baa76566bd7b147161bea9
z27a2cb7ccb625654f7204cfd11a7ea4eff1a44135aaeee909a9d8522387bccfc654bf73b1b3bba
z5588333ac820ebd9df6716472e1c2dc97451d584dc13d471b9b89348ff8f6ecf4478e8a927de30
z7bf965d5f0bc72113c0420c3887ae22339f0a1668574b4a9557719b37c392162a0b7213f197b6c
z361a78551e73b29b7d20c207761185fac28ea246ceb7b0bde4232c2f11ee0bb4dbb62adc411fd9
z827326cc9649b4a0ff6fffe1a8c5877a52035cc79b29d81db03ada075bbd464084cb8a8fa3f86c
z8f2e028f0266afa210b3cf65472d8433c478428cc7631c0cc5f7581fd7c99ae71f81c71887b301
z16aeebdf112b0a7f08b902233743b0505695dfb2b481df29d51574354495fb1bd61a4635e9ee70
zfecf82cdce18050c171a0cbb5878058f6b750cafafc005f36c2cd648701dcd10f9360cbc148ca2
zdd93d77324153ac1e3164fa2d95dba5c21cf5d7566c2d9592a70de202e597ae295edbfcb8fd2f3
zd72a1cd344df90d3dc6e70f6ac26f1f8c08b89cc4d5e0655d05cc0ad0aa90965d7369cc744e9bd
z8285342f53e5326c0252e6a578674755717609de031aa5007f394967676b1b42cd462d4b78df72
z85077cbaa32c638c34df5be65f4d25927e363fabc7cc34720c8dfa2f2b87744bb31a69c3fc6873
z095d01f207682fcadd67da901ec64302a9c4af62642f4e3ccebc07176f1b2f45628263be9053b4
z8ca0c0a4d0435b0947e083614c1f575d0127236f2daa584e1d0f48ec5c17082a9372ce144de360
zb9874d0dd84237f630a8452a47155c642e07b49d52d63d4ce02e73fffdce8e33856c2f3ac9c824
zd4966a677725acab073eb83616fc5f61b5fd9d9681a314af82633a8215b6bcf15c24b6dbaa725b
z34ebfe4af07d51338c412defb759a139f18166c636a289f169abc9fd2a29d24d1a775c5c9b2564
z4a18c20f43d4df5f46a6f2fafac83571615520e14c6ad83beefb1f90477e7788761159957e9572
zf824c07c9dba1a71266fc1e30a43e34dcaa01b77e84a866f63183cfba4b3dac80b777d0e190e7b
zc4e42e5e8f629806cfd0075cb4bfc90c58f045943bb59f86f314fa5c8d4012244af17d72114a05
z125e3a49e833013b6ed65d23b9285995a41f18804d7336c06202867c725faf1fb80c0920c6dbd0
zabbe36aabfe33f96017fb833bb080a1483c0f40ef0a546282e4c8d0612b81d10646053e1d4fab9
z9b42ed6f07224e7181809cfb9fee10d3a05913da32e096aeb741d559fc5041359f44826bdfab89
zc46f64e5c6c81d99f2ad46ad1e773130dca06ac1ae912a007af0459c71a0c2bd341efbe703afcc
z44d84fcfbe6a8de9147b366d65fdc615d1a214a5471e9d92de5e0306019e9abf853cfd84a92141
ze461612f00d27884af2b3abf10042a2672e752e7ad5527ea2e67182a3a33eb4bc2986d650a9bde
z0228737c1030db7328463655aa33ddd2f1086b284a64e961d9e6cef4842689977de30959a6c945
ze47965eb1f0b6cfa10637755799f72145803e7af62a63491fd49fe020d1284ccff4b7bf405d9bb
zc40c3602f270a4c21bfa5c6d4d6a294648425615fc451ccc160f4e77527fbb6084d7321e73fad1
z7230ea447b655c4fccc9d49544f88c72696aba425ea4d0dc30f84de7892783afa29daff7ea1549
zc8f7c71bd226e34686445f0d8f56febb0d1e10f19f08338133c973a6b9859e42f4ef73569c6e6a
z1db49ec981c40f3f4f4f486f4de340c5472e2166246dff6524674d5eba7e316ce3f0a769af75eb
zd4d375482fd97633a2d1d03460c3e164a401b684abf6077958e36368728151babca5fd08f61ae3
z84470134535cfb7c2dba2fca1b743f1ac9c39a29301a4e63591f70df5128a30a32de11783c9f5f
zd1d4ee55e7ee8560b7a00275b9829a6221cf7cbcd7c783d3480388984f0eaa350f1a5d319dd91f
za0ce35d5cc2a2be6cca59c102ff9bc260da44ee635b89caa7370474d5a5c9316c32990361001e1
z7c1847541a4296cd9f283af444e20f1da3faa27fd298d5e0d4de66bd8e20cc63a2a6309fe20eea
zf3a034ec4b8b2a0fefc6b35da548dbaa099ccc9e3ece305e3f5f38f45c500b5ce0f7c73f2d7456
z87b68193329530d2776aa5b536aaf4bbb90a80514f2316986bfe0b300b37c70bb47513a4a718aa
z9dbec240156f2dea4a630a770cb2924dbe180014d3290b936c4a4435e317d0ec5a71ddc2f7cbda
z6f764915245e804238f9f06d7d9e2a6adb869947fdd8a8fd9856487e4d63e03991ffedb0e773ab
zac8d71b873a164edc4d7348bca75d553246248af44a1180a9c29c3149233be3b119f0885088789
z240389f8322a1239b2af3c7133ac6038d5f6928e6222c57e8f85c980738add25f50f0d8a381c85
z4889230b8202a90c24cfbdfe692eb5927198cc7c3ab7cf61de5e8b588f97d3dd8c5838d4e829f5
zf866a046ecfd740571888e5f1b724d353a6ab63927e0dbafcea622d932d9195c332589662d6189
zbb6f18cf5f20d443a8b6c10a884d8da988b842a897c80a58b17438d70a3d8abc1ff793c601828e
z23a32c0f97d58c5899d56c5579f92149cec764a904bccecf2bf1c844bc493ce2a883889e8a44c0
zf1066d8e99d83c676a7ac1c1529cfa1f18c330c90003e49e5ae801e900d7fffa51f0425541b9b1
zca01b8946a70820e66802d979765bacb2cdf461116d0310f4285855b4339fe837346f5122aeaef
zaceb5b230f698dac2f47dcc5c6919094516515b82faa751542b540d9ce9b87ee559bddfdd3c2e6
ze19b4abc5fe898dc69f233f1c65540f04b7397885484c8af75e3bcf0e8b24ff39a168350318641
z296a32fc5ea467a26ac658d8da5b5faa07a7907efd59fdeb7bf36ba3e5c781e88a3d04c0466c6f
zf74f6ea6e71ea8e2f69cf14bb7d95af52cc812cf75bee0fafd1f1c01eeec187f6139d31f3cb17b
z18114ac14ab758d659b5857dca3d62a34633b02110055c4fb4528dda1375369e58436ac2ff0470
z3ac6ea12fee1676c602e41fbcbb2ab9df51f1c30fb1f1f50ce13aef8fef07800bac4913855ab48
zce3f50d99deae0bd0f425684ee856f76dca443004a74cd853249d145d8613fc74e652303eeb507
z18ad5ed1dab4d35e7008be04c9de9de8d394c4f282f0cc0c799aaf7ceab58d1339dcc0f01ba7bb
z8e244f9863835ee1407b9438dc0ffe28d6296d0befd6518affc8bbb3d56df7f816b967f939b80b
zba4d9ddd4a72603c70c36748562c9fe1cc4594c890cb7d959cf557fe2922ccedd4f79617fb9bb1
z238e7bedb795bbe1599123a507e3ec3c241498188fb67be5f91f83d350ad666515ed4163526066
z927abda2f64ca66b804c1381502745b9f56a11fe06de338c27973b78b7fa09d713c07973228535
z4113cd17dc76120f9fb5bf2bffd63e4312d0cc0ba5348041fa2db8695c4bc095decbd1a1eb063c
z6b341ce37364281e9e6a17d4bcbb9dbc6b8c369a8938393e453383a24fd274b0c8ae11dd61d64d
za8bae27a9525e871aa9f4ff41a2193109d0d14ead281387ce42572977c55e64565cdb7d660819d
z346e676373fc4016e866ac36e37540c8a39ddaa683393c7b782733f32f38f52200899ddd942f4c
zb83c928ec08d36681ecc9aa7f65fda2e3effbfbc145221c9aa2d446ebcbca33ffb96af1afdce11
zd00846461c937ce6b0e13afcc54673cc4c636bd48dd52188d7c483a78c8b8b63dba99d64a5fae4
z4a96ad04b0e8d7bfe083843c9599c67ddbe92f30757194f726712b806227943c9e6f0a48290237
z0318487a0f2b37282875b11da7009d38b2a510518dd534c6e14211336580bee023c2ae9f6ec70a
z6650e767515967df53198b5aa0b005b84ccc49dc2a17f6025eed10136a62c73146b8bc11a39653
z44df1c7ae0626334a8addaa9971c5ed83ed10ca83a311835bacd9b95e5c7810e2d92822ecc0f15
z4a782731ca097a3e8e751b23c579885e9aa7dca77af36a8beb03bf35d16b95c3e6ec23090be9e2
zbd3f9e3c4d650d5a47b5a9f80108b7b8ee4c1468a0c1f5834ead6748bf91eb506a52f6b0dc6e76
zba923c1c68ba2f40d30bff6d574bb24413990b365aab3ad4212363062941d7dcf68fd98ce5de1c
zffeed80b24aa95b4dc30fd03a1b3c614d071db4e1b2ed57e146bc299bec8990deb379ff0d4b333
zd82937bdbd553879809400a0964d3c6775c8397830f493e0cc83ad1731d103b84b7550885888b8
z3b64eb3450f296b269e58407a82d2c28ea1c7aba89e89ae90faad6437d802a2a51c7832fdec4ac
z08bdcc262b6de5b4f4a2dd0183653662e265dadcc251dcfc82e5b3525270ffb022c8797b9bc4fc
zeb43c49fad173d0c54cbba2d6c94368ac76da743c9f7f40887ea92fdd77e36dc3cdf6a240d89f1
zec4993591d4fa249d2e0cf83239a9172135d06c2809b4683a5ebdc4aa95357ddb5cc15b9ebff2e
z34eab2773d021006fe73457b102e5177208c83d79e902819e37a93b47e5d35d11464732da789c1
z4d8276a2d472b3b37aeeb7790186cb2234626012ed46ad8a9dba97808ec020c7e4de6b76050bd1
z0218fa2acf6694b8ca211dbf9546f4d551d7c8734cdbcde60f53ad1cfd2b6c156e08690f5a49de
zfdd6a5be5ac5d97461b5aa6bcf4b9fbf7623e3a2bde5eb3d56cc9af4d1ac6cf3c338870bdf51dd
ze2999f86955cc4a49b642f8c4e08d944febe0eaff75bcd6407c34eb265323c03dcf405515e3c84
z2536c6b761c75b93ded60a552ba5090d8338bec255a63dc3181a5d551406dc99e05c90b4593dc3
zed54670180d26fc69c69dd7667ebce1173ac10405a6bb2517d235f00d758dba5bfce5f794469b8
zb855de475065aa6522077a90ea3911586a4dbd7bd511f76c47c06bace95863e2344713207e1e54
z5c16f47be5d36c22db3c9a58be17a9dc70815a18c0af14de9fa0b2fce239780cdf58ec1e84dadd
z8aac48700ef502b61485505cf733111aea3ba09ffd5882138f3e37938416dc6dd46cc347ee5919
zbbb35f6dd17eef0b2208f835e7838eed123e39b9cf5b572a4367b33eb4d65aba783ce255169253
zc349cb0445e53efa72145be58fcffd965460181b318c9401974be591e3959d22b6b054d5b5b624
z44391cf3425c06d39191ee573e9b24ba061b579ae4d762031924e8918a006d416a2a17ee81be43
z7d6686c42ccb90481e2303d21a837c207630360f9fe4280c74678d5a3bab7ca47cf58662098075
z4de8002664a0eec9b15d82661d5381660b2c567565564e56507ca2abf76db6bcf245577b8619ac
zd847941575eb3a972563aa5530566bf0f3c56655557b850eaca01bf209e2d6f5e2ae28a07cfbfd
zd9001d1198ee8c2e1fed51f480510dd86eadc17967fca20111e7cd1d582df914b5115cee958a02
zd7dfb88443d3ca547c7b7b47b4c215ed35e1f09d073b47a68c974757a12b1a7c2f900f204cb2dc
z197e81bb2ee00573f8502da0bec126d6200c606f7a0b2c9b2692ef00905c28413128c072179c75
za36924f3cb0b9e62cf6450ffc729c190c5db2d4051f139a6c97754f141973018478539bf0b49fd
z8b6bd45fa2e87f1ab52c3aa36226ee389daf36b21084333b2241c4a2a647dbd06b33b85e82a529
zc7fbeabc731f59663536302f8ae58b76f3982f8cb113b91696fb1a6378069115655127ba5d1d64
zfcab650e35de2df64b2414c908a106143105f860b79c32c765bc06584aca78ed5e60ef8599e59e
zd356971227284bb5c4998824d52e266d9a51a58f711d105f3a5e475f4dc2c5b3446815bf429a13
zf2a03eeeab97d7460b90d69400f4d00c6f21a2400f54f83a275755e591ceb5a490442fd04cbea9
z13bc87f807f9e5d77d488c4365d8ecedea50d1b8ea048e74ae351944e24e4f1b43ad31f777ea62
z62590de00132c41d1d3f43af6465debddb03ae105f544576e86a2d8a8fafdac72db417b53483cc
z532132641912d88e461ed8a129986da99b960d2a50e6dbce6b5c88399f80ef4f3a7eeae1b7a656
zc9e0af80aff0c1889912cbe5b44f8f969ad8a6bf342c223922907772071d6f26a6e8b3b29eb813
z9603db4be89465ed671313b97a879130bcdaafd8902a09c71155781fba762e3d928964d80df257
z4c88658a2474035a04185dfff653087d76274b1b6832c3b6ced4cd1e854b5fe98339a286a38567
z50d2907551826a0240c1eff58800c883b838def27b99702f5456c8496cda214ba00f20a7a85c8e
z91a4935771367437f0af92b1e6dac965e60692c808d474614babd1042ca2550b5058addc919385
zb15beb6bd1afa2c3943aa119525ee74af338c2d8c18ed709013e0e17b178a3050d91c3c6b1cbe9
zbb96a5b3eec99d9e9bd50254f0467a477583751332e042994bba02c5a35d1ca82b79bf6591ad4e
z28db19ddb3dcea079821b1a2ffde11608958e2a64c5a225244f02daadf9659aa7dbe2c1db900dd
zbbcf7246f0aa7e19490f2f99c0275e2699bd3578533ea13d0bcb606e897491117b081d4e7780ca
zf7ace88e805109e992cf6153b2b11f65b4d79f7a0840050b0159db1ab852e4d717032bf3ee1d56
z892536829733748a3112eaec0dfe5bff44ec40648a55f9746b787f4d104f20069296a78608a82d
z77cbc80fa0da94286228b7915368b7b910caf465fce428b761bc486b85a98d03e4a3cf6be4c265
zc882d9bc2d2b05bcf6afa5663e28b631d57a9d45ec4700cb24e60ac7beee38468b122a517bfa8f
z781a6c2ca05d782dfd22e9ecae8e842f9156e690591c16a0301fb93a27272c0f54a2e0c495c496
z054ae44c937f3d8be9ce016f5be44bcfa7e0a468c2005c3bd47e6beb8916b3de6cca6e21b1992b
z905bbc25e792b0adc4d95e04e1b5ba773accd538b005a1c4b510
`end_protected_0in
`else
`ifdef MODEL_TECH
`include "qvl_hamming_distance_assertions.mti.svp"
`endif // MODEL_TECH
`endif // encrypted_0in
