`ifdef encrypted_0in
`protected_0in
ze74c34e226135848fe16db9ffd31815111b6d7fb642c521a3f628cf6da949865580b22efd062a7
ze90adae0e65e66a2c36a587d0a790699161455169ed55a01f2084f11770a774ec4c588039b380f
z6de9c5084882a40b79a175f5c2114b2b6d78b070cb806e1c0aa9258297f4687ab308bc470f0040
zb0b1de382961eeeaf2e279e1462520fc31c119af8f2b214846f56c2b3cd2eadbe4099496abff18
z15cec83ec4a77b868344aa20ba7360908f5c0de2a79abf8b3534b883bb12180f68b5d4beb444cf
z3fba8f13afb0abfe8fcc4294810f75afe452434d2d0f1166236c82f76edf1e12979f04bc35693e
z32ae028996dd85737a8f5adc1ebb94f39c940246e887647b64782cd7ab429b0544c173176cede7
z01dfb26b1f73408344a52b7e1f117f12bb9c8077b34876c2e6fdc085981637012dc9754765e1a9
zc512ce062e0b8fb16a214591f5c81e1353b900a611fe1f4886b57940b41b7f2ce99a7b84b04b90
z916f717e73bd10589c81e207ed77ec660a8cbed5b487fa50acde1b055c8870bd8676023f21ddcf
z9c98cc47cfa2d654ff1365d1f45035a045a66c5dfa8279050262ac56ccafe221d4824992a69d8a
z0056c786d54cd57e5ac49b6b8aa4fb7a6065bae21c146cc6f3a280ec9ff5fb2462d875b77aa676
zd56feb8da130336fa99b29f9aa3fa434693f259df12068556affc73d44aa85cf1fb7a203020152
zcac4c3d995d7dabacd5a5289e9ff8e6297752c27d9aba4374a79f561f75d038d6d8cfab388704b
z6c0029b1d1611915e0f0ba4e03db7c818b3caad04d3b2037c9474710b5ea0fa10be160cc4b9faa
z2d8fee558f29ac7729eba39c055557d2a6a92c5225cef50bc9f069ddef5f03d285a976a0fe0eb0
z2a7ae476c8610468b47c26df2553a0ed89c87912f4a0700d4b1a6d9dc49fefa219243fa0134359
za30bdff8de0d9b9e419b496370c68f748a21dd6aa537a27cff9e12e1afa4e56200f83399bf5b53
zc72238922bb18d46eeb145da8f51dc780befcc0ba7e0e8f848aa4b9e5411b462bdbb66f024391b
z35338d1b868355345029bc60a7c8661317e0d1d017e22c95d4390e5a10026fb958056e9dd03b4c
za64a8259d0c6f9b4be87c583df386c6f0dcbcaebb97c23b2c492ebaf3051050297d8277f7e2ffe
z068192227f1b3a4d31842a51b1b98174c136f14d0b7cf98a33c9f4436d033b89f02a68c56ff27d
z6e21369c9d5edc1f9dbe2787f9125cf0824ea8e8a4ae3d907cd9ea123d2159d7d2b1b4f1cd0213
zbe591f6ff153409bc06d130ab5cf90ad6f601ee174cdcb08b80856fa7c4f397babeb6f7e894a0c
z98647e2c2f6a6574821d4c74cea50b0760711defdbdd3a2129ee367a7415ad07c5514c9261d7ef
za9a338ea8f5fbf302ff5908eb1c5401f72130e5656f0f5733bc3cb3cdf779f09f2b2eaf5303ee1
za57a4ee0fd2442a0e814eff438ad00a9bd6e0fb91486d9dd248aa33cffe2c3bc1c5c81fb0354ee
z3f1ef4d49600f42679d6c44923a5889f446f03111df964c8c830aca81874370d0dcceae01958c0
z0a9f5f7622e3e431fbb3e89c36f8cce55e07a8707cb49373105fc792d9575ccacd123e73c3dddc
z2bf5a718cce5c5e5b43311aecdd2150558c16603e16aca2fff9b87acd3275cecc3f06fd36927b1
zb842d87815b22282bcbce0b6faeaa8873effa54672b39c6029394105b5dd7478374d3646ad7280
z4dc947cfe41601b3ed529165c7110d951a1155706336ae3a1e2c93a398e2ad9e01d1cf9177b39c
zc860776da2ae06b34236606480187a3d297778b4699a82c9d9beed863881aac1fa706d62833490
z7fbf0535b1adef90e8f97851794478e1921739a92f149141f18131de034dca51087ef786c1332e
z5dfec0bbad29d61813dff220f05b4157f8897cfa0d19126755ec6d478af42c392cf2083fa011a2
z49baa10424bb49d0de90b9aaaa4ed31ba5bcabfa5fdbc5b3b8124d80c283eff32db4567c200839
z846bf0d548e242f60740b367af6076e32731c289140f950fe27c1e3cdea7f727786724ac4dcd27
zdc452970b2e85d937790913ef69cbf66881e9e57cb7084e75b4e322291956018426b1fac85e973
z40bdede2a1f61a6cd354d1ca5fd592c18ff20e18dbf1ea112ef2c068da4a0962b86f1d9fd4f683
zf426f9d25efad592a15ced31f3be41ab60a833cb9f9d07ad702d021db7224b280559680f56a0ad
z68214296faa4b448d44ce9f0ae63e47c0ac322bd692afad5e8a7009afc27996a3c40b846b2d46c
za4243a744b630fc7b746ab4bd80bcd26829d8ef3e0fa0218b40550b5c8b34405454c1fa49d51a9
z9bd229c984477c4f1de196e3e5652c18a3989668265c8303b834be673ee41527e91815708795c9
z124869c1729f64adba9aabd8482d9b9c24ec67b65568c29ab784c23c9b25276bbb91384f382c71
zed868ae724489de34db0e58819b09bb070c6968da225080d792a5381bb1b2f4d47f6df6c940fc0
z6f00e174f8adf1a1ee70fa1cf1df9d9e21343e3ec7335acd6d9a9c70528bc8b9bf7d482dfacb70
z63a02e3d03764dc7bda4758ef680ea3d4c2a0da6a52d373ab94db277933dfa21a92f23f06883b2
z318bbb785f3bdeb4d8c99f7be35f7f46320e2bf137fa2c195e53eeb50aedcec7724163e705ac8f
z592cf162f902ca316de378da06068fb7a488426f57b2a04ca139b4c1d7bec1fa8d73b4a1252bc6
z9a513da4f8684437cdc71fdf8c40f28972fb68e0ed76b3371c1697e2ee36117066c0ba752927ac
zfbece8688ceaa8a69a863427d821c1c19b2c63a4b81185daab7699bbf99ea1e6fa4e0e94a726d2
z3e84a007437f2336e109a34501166d1f51703d5885481f8e98a6ff6b92f6a81a699d4b4924f32a
za4ce562b1f07b251b39e0755a47081b42d14830a5a829dbb2ffc2276b0ddb47a44032198e0246c
z724836a5871f3ea3e9c99116be5e93873e5f289c784cab36e78766798cbfe261fa779c416ddfc8
z03594cf58e17793864852d52637af573df4cb811ebc9351b848dfe155135f26d7f2e06af2d94bd
zce6825de0257fefed0995ed6e7f0bd94a5dcadede73d8642c4d272d03852654e2cc821d0c42a61
z2b39f72ae87308a3789b051c22189d9da025cea894703e66e582a6809f4ada33a3b699b3b10697
z7878b2f1c97d36e03f57bbd0e0b8d3bf0f07fab3609d3b8aba767c2d2d2924c06cfbf7de8aadfb
z6e7572dc1160b9d688525f7d522f1e327caf2d88c4a31180fae4bd2e2342eba2fe1b5408ced569
z6db2d000305e1fc2d09be36867aa8fa6a1856f2ff5e9d94b7d79e8435dbed275370154f7e0cb86
z89dc817040cb373e7476bb68d1387b19f2f100ee4da68c9260afb2e166d138372c21902f78ae57
zc18417661b18144ce92e6c7259762d153498181991f753b2715dcc141a0ab83f7194da067f1865
za04db6977774fd1174dd260002f3f1842b19db391fa14584efc9af61da7fb27266ee6a4c3845f5
ze48a71a84c62e1358e30dd234306da8a2db3f07da9a8c9372fd1a0a28f759196a6fe7dd9758ca1
z2e03c6b2d09e760dd26cd09f87b5f3b9e155148e05464c63c8a78a9ae7f5195e4ddbc1641e1077
zde1903f8bdc9992591eaa050cee64eb0b79729d3d97c287cf88028ba12760b6e29d1ec7cdcc9c4
zcb83b9e023e9b92538bfb6cc1d0a6c0425d336e68341b8c962901abed45b9f2208fbe874bffc20
z879367696a9bdc03aa83e8c0472e5c91f314d43312c9c53065d6700903f685802240ba1c22cf57
z0a2ca874779889592774b97d83188d51bbd882151429bda1f3769819bafe22e66065e4d10d1ae9
z9fc337cb7f338c209be92a8bfd1dc4a20b8238cb37f9075087ba32a44cc71d36d8285337c2f173
zc1b1b0e3612c676fc236d99ffbc0c492a4a6ca738820bead1feffd24dfbdb915765965be1ca20c
z2bdc254c7c4924242685d4d154339989d3a48a7e65412f9a22efe025f0dbfd9e7e7b3f393840aa
za65ed5123d928c3d32d8402ea83aa3f88184aa06096fc2df1c56830b57b0c704d522840cc53817
zc371587d88ac873d5a59e8d353b81922fd47e89109a50dd0b7d8ed9e52bd61f5c00bd62cf1a556
zed0d5c9aa88f68ba984f5f76d135a2e3517e5fb9eff3ed9716227129a0c4a7b37486ba1eb32864
za837b81b90c05491540468f5330b6900b5f86748fdb83e3e151f59e93d8a3e70701fc9fb45b0e2
z88286d2fe9b4c2751172c80001cdfb89f00829ef0db9fe666969bc26360d78e3ba59750ed481bc
zd94eeaf0d6591ca344cd0c9017151986dcd5c163566f229515e01dc81895e075283817bb7d047b
ze999902cd6384f2c33eb4708088b3fd5022cbed37a66abf73461cb561dbbf55e44bcd124e56f4b
z034332a6c1beb9b5065b534aac2095feedfe61ca4c809cc2f6e9be4df2a1752108fd17309e4e23
z37caf480a54a6459f3880f5a31a482af4514e93a4ea09d61b0b2a4f9a4f7e15da00bcbd597a7ce
z3d87e9f55edaf22ac8118856a99dd525be77edaa753ba3970d84ca37fcb366871b4bb324a0209d
z3fad4e16b6622609cbe91fdacd17a0080aa0c9968206f63d7a38abf928685290289406c0a62737
z2b85729c6b1ca064fcb9dbee63f7e2ac4ecedfdd90fe9e8d4214c5daa1e400a30189800a1245c1
zf8892e0e95c085224da9f96bd222e37c0ba05c36a85423b4be6428fc90fa5bdd8a61f2cef99af7
zef32fe4ea6b88d12bc54c378543b26e76540d6eafec2591e833ea4eb9bd1b00c4e108eb2359ebb
z5983fc7b2aea6f7abd055a09e0bc93a101271362e4ba8837e62c6a9936c1d7fcc676d0a2f59036
z12b755089d0780c4a290ad1bbbc9ac9bde57ee9167b59ff6653b3eed0acab4cfb716c72c68d42d
z508f015db13ad21c3c047a923a7b1c1c7651be4f2dffca708ce9907d254540a26f78087cf023a9
zfcfb233ac67975111839cdcf534ce626dd3aebd55caa41d2909385d3151fcc8bfd26482f97a9fa
z25a0ceacb60f56fa521795a86f93b66d594334d5d04b1b9baa8a5b68597236883632376059cfcd
z0ff3c4738c8f634729ae4edf3f28884634f07901cdf9318111c130160a2ac95c8e099c03952f10
zc7f47619372a8b734d59ae3232b5fd7abcb9d056f3c98baf9219b4d36f041c564df393190dabb8
za1708cb7dc30b40460c0a0e4e7dc3c77a52f509900c35e18a4cc3e2670f34fa9f69b0abacfdfe3
z15011e02e199abb4b25d2276cd1c205fd1463c5110be6e1b44d734867c7424d30a5bbf9e04a914
zeb8f5bb5a2ef6b5911d91eb3f73a8179ddd24c47f81690a947886aa7eec608ac24d463a106b983
z8cd62473ed676f677f710b97f0e286d1c97ce106aa1ed076435193e238bd09bcfc8a13f8cdcb0e
z2c9e892993852e4237c61974be1fbf648c1fbbc3d6ce8714599690e45a69a803e1822b59472973
z62812512e84d35bd44f33269c36026f3de6ab5b49675f2ad834fcc25063c6731f421cf0cad753d
zfecf65d598c63a6ca1b028d3e6b4c35a64f5ab56fd71dc6d915313e953eb0b2856d923dbae3498
zaba951cb046c75cd6095f60c8c9cbfcf9358ac21c8453e5121a7fe16621b70c8568dcfc0a04d3b
za5806e37fdfa52d4d44331222ba0264e72b3ba28fb5747f99b7077e39f75e2f424a33ee2f0de21
zff56a85e62d478707cf38031c34db2e096459dfd479b5e31d4674c572a631708b72fef257fb292
z220449a5a57b5992c14894774475aafe03aafca17f24f3dab511219b820b550570d3d48a0e81a9
z9495fbda06508df29e085f08cc493ea22e42a833aaa91b7ee9d84948d73f00aa6cb88df9a92f4b
zf4c65b1949fa435c362b03f62c0a804f4c97cd78bc3348b8e0a8f5977cf019bf1bb9b192f922ce
zdce2d68fa4790fba53187c253f4cc041f0093dd131b9a6f9d40873f05d494947f4147f7a46217e
zc3c79b30a752d14ac4badff371b3cd116f7fc586409c1cac22195df6fc83f417a86b53134a4f2d
z583c2eb9f2a9d5735c6e88c2a0d620da4ade0c2548825e6e1c44f07495851d7ed02882d6610316
z3441673ef525b9020ad0bc3f10c581d51f58f9162d13370dd6e2d1dbef8894c8217fd0416756c2
z229811b57edb7e1d4b14fbcf33b1f048b363ae7ee251ee4e820d9ca5c7d3ec4e908e8731ad92d9
ze273e37caf4ad9859cd64356a9bdebe32b2eb8ff7bcad918b990d496377ae45d26ba14a7f70d4b
z050f2f9d50fa0085b98a232223ac28ee4fa78e05c1ab9d3765267ae34c094dcaf59c2c58464742
zdb80ad924c3c1605bd63d6e05884a034d5498b0f861a9b7c630c1cfbd5e4291564b9e7ca32e784
z85d7f3c3da02f80f3d05cf5e9f2f4d9b666cfc5fc52fc674a9f6c1d6434df80a25a5378a011a94
zcdaa0aa5375aa2362e142a30cd08b2aacce4fe7c0204ae4ea6f10be6e08a39edf40273d7a6aca5
zb0bd37f08f1c9eebe269c50001ba6a1b23a4f4f4e4900d71e29c5c7596b5df7f1495631deca0af
zc69047e6020dfda4b42000d5a062eb8b8d02af6024e9fa9ec07e131e1630bd973985960a5bc3b1
zd57784df7336baad0e05c6714e12949ca447fa458d43d34f6fcee003a798855480d16730c615c5
zb42fdf2daaa2840c6b2e7d610aa1c8aacd8c8a65036d0a2ab9a1e756fff553b9c02f2c4e92b79a
zdef646f1838d071cfa474b8189e57000b4257ad724b62f4cf349dec7d55db3b18dd49b82daf2cc
zbb79c8c5cf13c00770f24014e89d6925aa527dea07cc6804ed990781a03a4790bb467853f33be9
z305e8b08b7afd204ff8861aa9ebb7e37e90424260f2cb6c52c31181030fcdee02b487823eedc82
z0a8a79f968a93184f07de5c8f7c8880f4124f19674e706a086265a434892b84f1e12f8466424c2
z3d0ba30baa2a1f2029567a5ba5925a8832e0384e6e7cb7f0ae411113b345bf6497559057c90bfb
z4db3d54d028281ea02404bc43f8604d0409297a0ce23e7ee9876370f37fa2ff84688f9b09b5a03
zc8d0066c603271a3dddfb26f59a8429ecf4cfd70a936e8158dcbfca25e229453015d8e5e5b732d
z0b62fd74fb957fb5035b6c327052ba85db8fee766155b119020a6b79cd5b575556af297520f6aa
zc81c03118acf41c29764b1b0ac9ae84e26025290608c38242b544ab90d8c78ec6462a9bcb19145
zae5bc58be0d1f35374f179323f6c060fb432da70426ac57e53c8ad92190a70225dc28b31f8a667
z23ec3a86b8903a988adf810fd223ab4f03d9252897a153cf3032f5f549079e5a9030bcdbe7f520
z735ad48002a371a14822c4996d6283c53f28a61d8e0b6e2ae71da585718da223c46c8b41e0deb8
zf6b2c75bdc56c37cb5bcb0ca0b46b36d314fbb62e1feb3524f0d9f8582f26ef1677edd111d7516
zabad9a4173f1cbae448d17efbb8f443d3f80960b968f2adcc35b78f5e9d73df582777768f6ed3b
z42f3e6591995b84db88f34e6e59e4fc439e52fdd020fc8882ea95f5c742e62b48b3a2a21234dc8
z8027c153310f50cbfb994a5ceaf5a3563e80f45904b85baf7716909e9f829412d82ae9d254be3a
z84ecc73e7c996932bdd0d5e8e9f2c413dcdf82433b7ad0d06bc1d74e7c03f6b2e8e57f6b7b3aee
zc2c198d4d8381d63331153ac1f95b3f278d995b7abc8029e754e6cd0c538f86f0925f34ead022e
zd68a3de20d3ef6386887bfe7d5657316d84095643fb921d018404a233d4bf7124d97c5d89f2216
zeed4577ed1e6c1fd1d0cc502ca0fae76eebb5fe8609085483c8793adb581d23519c607b4b978e8
za66cd6b44495db92bdcdf9b1ef5eeae4f17e66958475bb2898faaba034ec58d492ef35929d40d9
zdaa882d86a1a2d4de9967f5f46c0894895dc75e79ad439de2a3a8f71e72d8f1a18c87dbabb2710
z7a94d790d8b82cc83925c85a2ea3d2860cd30e3f492afd88336d80d3b92083bc34617e01b23fa9
zc3ee48934e6fc19aee2001ee990e7ad01dd1307eff2551e7e62b668236125f271c686aa491322d
zfa53ef2bf5be714a9631e0470f8e6ca3becb9a33694813470b166e141ccb4ff8f482c0d3bb61aa
z9bb41eb843c852cfeed004870e5d619e321b907e65c7c9ef3e178345974f51949c8138d1c8e557
z6e02b80f6f3e012720419c8b6a04d5b86e19c9e8a8c8307f8e38ec3afa4f42506f64cd14de771c
ze266d164dcc8e374411f33c74cf8a452052b72821f57eccd30cb5327a7e5c5e56cde13d081ecb6
z6ff8917c880116f955850bd54431fcfe09c0f48a805d484a0593a5031b70e136722bc5150f9ecf
z811fa7f131ec83f46f57d6d6911f908f72e286af071c221908b75cd5774bb01c8f2fb6a69ba1b3
z532a050d08ebc205f2cb857bbaa24f1fc6af32dfbbafa56886987b44c16610cd422335524aa04b
z5d10640e0eb70ebffb4f4f8c71af06d8c6c585349034866634a6fe2089c0b562b1b7c062abc8a4
z2b4f84fbe2123053a2c6a6f9a2fe5e3dd73f35b03551ca8507b2057699f83d93ddd339e618a466
zf94f15753bcf256c6deccad325d96c9ea2a6b97aae3d02fb82ed6d3e083e4e63fb86846c5a9a73
za2b67b5d4ae29c1bcf4954d014efe34aece30305df279ddd044f536993d71a6db395ede1c9fa0c
zffd46570cb1a00d871b98a903f07864d9e8afcd6a9ebf3712b16b8bcb91cb6c44bb149d1df41d6
z684134ecc20a5d535cba3a7554d2524f43882e2df495b172d7f4138fe7e0cbe157a5c5c3229352
z86957921a546bcdd1da81282b0351aa07c5d22f3f20d8639da4c8a4bac3c3189c2a59000e9e41f
z1020f494a7270bbbbad62eb3008bd2f3baa663f27b027e58fb809530acd41536c7f3ca16699a83
z7bc5d1e825b0dff0d5bbbd1c6da52ac0cb0fb8f532e03176c544ec27a3ac0d249e5d1ddc01674f
z85a4be0cf5120e3851a4af5f18e346297d3c703f7d2447faad64f2ed6b46a7e9415240afccab64
zdd0e2595d26e547509d1386c3cfd8088301a54428bf48f491b50d582bd8e43056d7a911ce9add7
zaec7cb1a44df2220224bf3d30380fff7b86cf90ba8249b9bb82b09ea4ebad994f7b3e64ca86279
z5b15e77d6fb95587520aa52f0f6e6455e8e98bc0102d19c1afc243ec5cb62cf43226d3524179ef
z63e57c5d1b639cc4e7ceb4d9b824b4f5740eea77f2c3caaf5e5a932ceaf8c4c57350f72e79ba70
z2682c291bbdbee999c7f564249972f5c44dc84643f048fa214197e06dc7c88993c831d58506b66
z7ed1a81e4579b65f98454ee9152faf12b7fcac1d3937c7f25a311b5fe1e55a296041af58820747
z9799b2b913dee90017e300b99afb0768a25b457b181ed9e57fbffcbcac31678cb40acdce77343a
z9847dcc903565e64373d91700cf1a6f1262d3aa95930316026653935000818c94f80f8f1ec7526
z82d095d5cc789c4a20257b16c846baffb3fffef11fae7c4cac7cb09f85112453152bda6b8e3b91
z29587307c6709d571bbd37d5c56dc47032fb5f5838e3491be0e4eb2a2c979e8ac54ea6421a9be4
ze23765006a786ec2155702768da3a3cda094e8c5db145ca2b9e82332edd6e31d98c6303c93e1df
z8b1bafa3b76f5beec4ae6b25ed77aeffa7fd9521e2fb8168b9ba8a32158f1d10498b60b0707693
zff633a904248b315eaa73b79ada178c49d564dccce537c47a6336781a431464560da8abb340454
z7d83e05e288d03dd6c98c736a9adc857192fec83687ea4bad917cdba013487884d6e933a8fc4db
z355743bbd7b1bc751ef67c5f702b37aaaa4f854966b1699a55bf98a065b516f4ccf8d0a5b6b292
z73f9629d73e69a32713e7bedb930a547192cd94c8d9457da68e20d6dde301f1f464e81f05a897d
zfeefca0aa255c9339440dfa18faabffa0143f5f9f1b682f97d511f2d8eaf4dd2d6ff7d395fb991
ze920dcf19583785f73a3f18d5b15a68627f964eb9f49f2b4965fd5852fbad8ef68c4f9c1f24cd7
z31e9bef0a95937cfd77e2e96db5caab15f9c896d1a3225ec64f60d93f2641127744792d2354d3f
z6f6e995691edcb15bfdba58e8921494a20136d9fe2d1343ca67ceb083669893362d2c94bb8070c
zff4a1c367fe99d9d15746280445c405d8c308c99c7cf585ecc83530adce2724054d86817ce7b7e
z0e5f5181ea821c621b168a675d44eab5139c9d31fb7df78c84ae04727feec41682957ef88f9b38
z6d3a97e85406dab479f63e92bd3ce077cc2d9abb1dff5b94ef90debb3ca3bdad768a1f8bc3f80b
z7e316978a0823faf2183a2aab6c15056336c8a0215bbdcca21c9271399f62a3f8ef58ae52594cf
z5f42a6f0d0e6776605b8df42217f54d988708b9a2b1cfd513659ae093dab136feb11a8ef61226f
z1326f85e405c854910d6fa26435b7f8d6221533c5d79d21b54214373fd527014b3469bca9770b6
z2e2c5b2a3f357bb299c065a09a3afc14d1f99b09f5fc7970cda7d6b7410d37363829ac857d99cd
zf0b5a56d3eeff7a7f17ac9bbe5c88759b01e9b60cbea32a425d92ecbc49a62655c9b10bb2f3e24
zf388d9d99c5d32d1c9087b1c69e2d54e63bd9d036615c2ebe74beb9c47a803ccaaaf578fd0f885
z6dc645b7595d461611cd94459a91a0ee657e86423983a66c42f8be16374391a892bac97c2649ae
zdcdb744332799cd0be636f456e5d7f2c5540aabd24ada1f80be8257fd70fbb168e21a15c3dc055
zdef011197c3e882038a88b0ebd74b863f561e92dea1bc3ce43c314682bb11c8f6056742e80a6a8
z60d958d0489d9010aa8cdabb912bb001aa22ca1616f08b799cc26f31be5d2828875f2e4e8b1579
z00bbbeb78d3df3ef8fc65e0058d07e73ea4590d11c4684cd6fd07aa77b305c29520798cb406dd7
ze8fd05930aafd704d7e21586f50cbfbc6812a11ff3bdeefa17b214dd97a4df585bd3eb63a00a52
z0bb99c6bef8bbfab0d9ef5a5b6e773f5b5455bf58ae112f55513e581e2d89e88a7313d76255a3c
z8dedb0bffd441913202e6282ccbf064527b31bf0ca31203e8f7e6f5aea75b8eca5067b036d8358
z1d7c960a72fe048553a075f0a93d8ba28420823cf67fd4f75d3dfbc098c46f554234874f324dd8
zd4db21bfd856a671cf8a82c19977e33df8eb97f54cac3670011088724a18f2314c24c560fd37e8
z28e899549eb4254d53cc60103eb515974fcccadf0ded6b554c8e4c89bba3bfe29893f540e8f9b3
ze2a67b80fa4027e8a4e2dc36255659be3d99b75d086d172f5562baca63977621a900655e6b8d91
z20f3576266cf12a928eaebf64ceaffc963032fec1eca5fcbb49d61350483e781ef8e588c5b3470
zb270d39c9eca9907f20b6b1b0d5df6ecc16cabde06cfec6d5516e94a3871bc9d2f34768eb1bc18
z80fee2404b40e5ca9e23452417e390df5bbe8d72fa0367664700fca3e8d815a6e4ccd6b2dd09e9
zc7dcf7e1657fe4623bcaf1efa754582b4236ac401d556f0f9704124b9e933616702a90dfeba206
zd82d61f944c14658601613f89d9a54e256e2e85c0f81daef5f3ce92f00031bd93b0306dc73425d
zcd57f1e1d2cbfe8b7e422e859bcce67b5220cbfdcc945f28cfda0ef2c52242f7f1a8258a8a7106
zca16e857cfb81f77ea7c938aa89d1b33f915810f6a209569201f44d17ab19a8c5a3e63a4b87fe7
zb480cfece01390011ebd1279622d57abb03d12a4728939dc56e8fe25f4f79bc71434992f20b324
z5f75d1c0fbfd055788d5564c57fc8e68de640edb881b0a1ae918c7b9995d3b332508363bf57d5b
z77d5857675921071e36a326294d4f0dcaf8782459f8e17d3dbd99751b6b70a340c50a02adde21a
z413d20caf376e0f0f8b7ca93fdfb0a64325f8633bbc5218af87140e03d770399ca15680d47f394
zc981420c2d3a08fd27b801b6e28e4fe99d5b2dc9003d10775fa5f53d008ac51c83b0c81a0d6fed
z1751fdc45e1b83774d251d0d9c04cee86806bb7ba6cd1d3169b1ee7a1522cf310c655e42f92b32
z45e7dc7d8fd29d1ca3f6a042c311ce1dbb70f659468489c3906fa8cdf36b32d010fe1131e25382
z1f82b40cdfa3f2859e5b4e68f04a18a14bfe81e032d214083b406a932e577ee5a412cd4d67a05f
z1f674405d2f88e1cdab3bd2e28e2651cbf2f430fe65e760431c09df2c61f9ccd4e1e591a422132
zeb799ba0ce9f116afbc2eee912189eb15122456c6e4266ff373c3102ae5ec1fbfddddc20a468ed
zf11bc4225faa81c665b32918827381ce7dc7c6581565dc595588092c3c4e80450ddf7c5d576b99
z98dbd2b662d5a5b304e7324d399ab3a548ebfbeef4624e5c3166ad894039f74af4a294f539ea4a
z00e6e28fddeffebc2bd8e59a0cb7c2a706e3f77dc56715b931385bbd71468ea2fb587c6257369d
zfb481ad24f90f5c00ad05241a08052ff49c9e92e1e3e8b547672055e5af9cdbe89f85df350b720
z30fe6114dd12b1c6eb4b1d5b5fdac6d63044aef230f9ebf0ad6649d6c659709dc518fbafb43b40
z3f5d8b8385cba8b816bccecc0182e4b667a63414913c5caba9e552da5fbc6c22f9889afe7a55f8
z8e0cc64033b90a32300fe61e978bfe58fb16772026fd7dea65f5f36b331f55c7d4cfbab6270db8
za25142327c5c04b3a8f122159eeb75f8aa7babb8116d3d9514d5019ece82023f9a94605dcbf6bb
zf3ac33b7dc03d5b159ddcffc37c969305d5c5cc051f8cf80210c1d8c748cae9cfbdfd1128a9abd
z1618864f0f47a7387af05e83ff498bbeb1d123e00ec504e1afad0d4869ed9f28e1264d60be2621
z469f1121e97d880bc66059ad8ea972a6505cef84458498bf8e5e11cf3bd06918b20acd886b289a
z5a1bcd381dbf826f82124c4fda40ff6c8f48205ed33ebc1eb2da2f65e4f1e7d423c66540eea853
ze9cc7b3ebb60b7a8c0a7261c5bee5911e6b8afbe3b0a21b3e24c76c75a245a33dcf7693cd6c2e4
zbf177579a10cd39e64f1b37328abf374db5f4ccdd5ab8fa5181317664ae587b363cd24e12abf10
zf638bf76adc0dc2c2885d42b718d7f60466cc168864fdc03ede29160bdc92800f86f5aee4d6c74
ze3566da967a1a34411ae25d11c7ac26a601b0a05b87d8443002faac05244cb3eededbe58ab2905
zf1a9a8565a3b832dede57273f206174299465c16e4582dd0760149787d0064cab358cc0862763b
zd1b0cdb475c18ecc5216bb5030405e3e0b189639639ca4998ffa43c1785a5109338ec94826cda1
z4983b1ac6f241f5fdd5417ad234825b1cb196434cf2759a793d7375716d79d4e2130cbee921236
z6f9da23f3cb0724082524c5cb43900b8101c8ae4a9ea09ac655a27db50c452d00e1a1cd008b30d
zfcf5c91317017dac90460de4abf614ed190dbeb6faf31a274091370e558d039e86b803ee4831c1
z5f240dfc9ea984bcaaedbefd4e1a8e4500727432b8b5f15a829a1bdeb40576b6790d09d5eb185a
zb55d185006f1e02096399d2935fa99440778fe537327f81e70ca0eb2bfa550ab7b6a94e13644ab
z52ae80364e1e85673b04504b3f90bf5732336f215ae8b8510e29ca4da4c62a0a072d7eb8663962
z2b8b0b57349de1c28b5d86d54a0f07e407c0f0db97fbb43588c7851871a67fb234f47f63a40ec0
z1af17bc6b4f371dea74434dfbc532aa0336f320b7c37e6a62be90669aa7355fa2a8534f451ca9e
z44b1f24e1e61db33acc15da007fab1e00c0ae751b3dd31278cd25e8cb1c32258ca0bdc4fd089b3
za769b991d34580c6e9b52a62ccf6e362df2d9a50b4227ea897da73dbc9c41950d5931a875c6f1a
zf9e04e07346729d194a1c57cb5ca737b5729c777a4825c87b77bb83ad79e013f9820762636af88
zf176f2d9725102d94a4f8e776778366244745d1985bda5f536814bbea3241c6b468a6110ad5cbc
z9fbe9203a8556143de7a1dab477d9714873e5ac8ab3e4b3962f0488fff3862949e286cd3f4a1dc
z654ead04fdb3672b60b966e2c1d5042dcc4c0f9d92ee98c9cc6c0846220343f601cdf64a3391be
zbcdabd6fb4c33639eb7c27b465f56ecfa76c2c5856494b55e345c73378d8939ceb29ebcf2beb9a
z76817c6a3e9f90d8c7ab1bd91bf23a722b176616978a63c084d860b393dec79a5acd819ef5b291
zfb2c3755ec0d6208cc853cc74bb3e8adfca8dfc7d84207b7bb09f4d471f841b59d309713d46895
z7064036cc1797fbef4be5fe2efb951f27fc789f74f262f418c08e4d8c36b499d6fc1eab4f47c8e
z82318c2c0a5973b28c4574c62f43e1d06f6948e7e73563369307e4a25ac40f31de0db6c279fb5d
zb0facc83f4cd70a2bd348338d94075ff6dbf3308d95d08e39a96545ab27d70192192b851fb966f
zae85e0de43c26ae80c0265d4d1980aef8c23701fa90b3868507e4c802016733195cf09fb56c34f
ze6cda212376e12c77a4fbef1ef9dc8a4fb7cdf682ab80778fc8430762011c5fd260df3abf98f8f
z5ad71f5d159bf8992a945d0db51ce48ed1460a280c3adf9789fffb72074308b7aa5e9bf377f58a
z1af1874a0f02ab93432c762c16cff8b69420d66051c34158237c375d2046b9e1c4b77f39279711
z46535e646ca59a8c7b5556a6232d6b45783f2b48d86a863bb3d60192e8bf9c9dec860e7c38b287
z8de7e214121f24775ff657922a18b68b5783523d1679dc6226284569e8b13de17372cff7577872
zf21a593582b4e04869b5bdf5f85ab6cdaee571172c007ecf2639fab8272358a021c93ea7207046
z669e2bdbadf88c02977de8bff9dda9541ad135f37535364e561087311412c426ed5164fa895d3c
zf1e3172900b7310957dc6fbce94b179a2ce639a9686111a8fcf20218562dbfb670b68e037cae69
zfcece69230e0314f6d26c90fb9f55e7458fa2df099f94bf24981b016ab37b60b5c6e4ceaf43f32
z99035aa8b0c6cac93c214d5d735801f99324f79ea68aa8f2b85af429ffb61151078a01fbad9d7d
z91c223bc79a892357c80da05906825ec00234922bd6da6886e4c7acab6ff3179e455c2b807e305
zf1c9a40f24ec4c61cf69082ddfa27a1e1bbff0aadab0d39131b3dad4c72f20bd2d58939acdfbfa
zef30036fd88938e9f2495bd1832351f3978e92a7dcd969f17f47c2d78e79ecf8b37c9a5e7d672c
z30552ee1502cef50ac6f3203b93225b0d17a507a46f8a4047256495913c98e1981235e84f02818
z7c34dcaf7880c5e58a927d9281961d0b76bb63cdb14d00aad3b5ec665dc6637fe5b9ee64eb0d3b
z5d978aec4533cf781ed181c1b89dce194423668aa82898e0feee68f9a6c32b873d2cd15bcf2a58
z9e1daef0c7734392ac712b0cd28b9595835495b83231f60a497bd3f40b47484496310fa9183551
z9eb30519253f430fd2cc68d20887cc029c000eb6398eafa8aaab00fbc9945e35b5766602f8183c
z9cb30168bfaf65cb7716af9876ec7d517d878cd217458d2fbfc874cf8d8883e74d14e8a6cc2345
ze0e6014e2553eb4d0a5f1ea4d1ae2379be1b17aba2111ba93373942972d6d7c339aa26288d5108
z3b491a0cd3cba02fd8db1d739f7c9a60ba9c92c0db3e5328115d5eeabbb8ff17ee14e291234c59
zf78bc5f0dd7f79d1d3c5f385dbfa8bb61269298f85521758a2153faa7a69789c23352c317429a0
z1e94c5b13af9b63647b7765e5368f14d2656e6ab20202c002204955198a3fa5b55d7846129fd31
z4fd2be440f22b6ea9176d85a9b486d1d2c6676e14d5399d6ab48c0502734224135be6df1eaeeae
z3136bcadcabb40a94a0515d81f9dc92b92e0f9b94aa0f09ca7c06eafdf398ec312d91844385487
zb258df6d9f31ab527a12196f0343e05d5b9a9dcb168cd65f242d2988ac058456a08f244d4b745b
zb54bed943934da8cb8f5ba24ccf5242ed550693fd9ca6be7ad278899b19c0cc3f2fa473cb8b295
z2698dd385e34c9383285cb899f120bd1d6ca9911cff64ba44d7f54f59c3e7de2d911fcba5dce34
zb359a53aadd0320640ecd6bb936d4d797a14f09819b54682e04398a83182bdf6b87f7421a5a3d5
z9ed5a2e18cb0cc608055e714207e85474cf8f6cc38fc846d6d0db874f9cde9fbbcf182f6076bf1
zd4326e44b89344546e76d8a04d6b1cd6dac959bfff8b44955a438b380fbca400b74618b7de3ebb
z98b0a48e4a6dde6bf8dabd00221cc191909770a761892850444968b5fc3a3e130b65ebb2f40c4a
z3295ed73dfd26b8dcd57a43e67939b0ee547fd4d7f58d33fe8ddbf319af6b4606b7c3572f9b465
z83ac6cd15dff6417bbc8755a466647799549568d8e508d54128e69bde7e193fcf748f609d06387
z36e99b9739ceca8d455a3df71430ecf0d2d4853bcaa9dd929d29340f5c410a6f5179f24efb48fc
zfe621c2e9055dc8947f18a14917e230cea4fe7be32eea5867cb48f17ab8b12260f748975120061
ze674b1a52522c423f57a816515995e71facde8b26761b981995752888ffc9822309ab32e192e73
z5c1b12169c9fbdb1b151da1bd3c640e23495877c3a5c72fe1d912768e625ead30cdd1227b7ef91
z4b37ca72934049452f73fe8dd1cffe68f420676e94f044135cd8b1db2c50f6c7b98f3cb3dec302
z0ed1f2b59768c645cfa6a1933927fa711b2a8d613b9dd8f79670cb959b2897b8bcb4615cc782b4
z3ec1ba81229c761f06cc92d489e14286620cc15e5c5d1156db17d256b21a38b109d0c3043e1263
zf35dabb255bb8d4a603f71802f5110ab669ea7a56b46b9f881220f7e9b911c6b397a0786de4c55
z7cc82dcfebc5e80836f400235ef258f8770a51cd167617baa019ecf01783b0b2e15baba0bdcfe9
z2ab4d5b2d19945065912097f470c0a56006761d05f3eb0d874a01f99eb085a0a2ab31494041233
zfeaec4c895a4a3d7f4cd00bfead232f35435eed340c526e6abbf46f18f7495f0cf2baecc03b55b
z14b12b346e5a7b6122ebe470055061fdde795a3eeeef1f6f3babe04a2ee6a921ddf41747367303
z780a43b7ac606db41e487bff4fbd96bac377e6d5aee06343d6b7c218b19013eefb3239c518b942
z8cf6285c8071c01007d8a2b73cbf2c63e8a692b305b7e7eb09426e608c833ce4cfd3b48ee868db
z44a8ca2e520c778cd9c3e1f3fe6148e14be402f0aabd43b25051917afb333c0d5ba0c934e1490a
zdc59db389ef883846454de19cd4c108e059e2f0e290b6cbc0a0781297fa74728033027aadb61c6
z5baef6f3f56356df3c3fc4252ebf9a486956ad6485fb3ab061d4e5c6fa6742b88bcf0dfcd53f2b
z0833165bf7006f418318e44230cb53b4a05ad132989b2676d59a523cef76007ff0eccc19baf33f
z0cadc7f9c9dd9ea3d9a035f52dd1cefaeb7d3584d64c2def37918f77f616016ade2f84f524e17c
z11cfd8548a3f9c6013c30ba3fa6d56635d3580173baa3ac42712a1bb554719a2660a72c5488d05
z1402b49b94cebc12031896023000e859ea3d906d315abf18b3d18472c62ea9600076f9826360f1
zb559eb4cc4ae335c8daca828d2b6f3b098b28945cabba2a6d6bc472674f5fc9f8810ded2a9e691
z5dd7076d230348e7e97effaba2cbddec91173d9ae9778411b45a79b818526c6b89fd38eb8d5f79
z9967b8c8188d1db1d58c15ec8591edd298298084a974932244331af708f71f55426af7c7ff0a87
z2fc74bf21868b32e52373e040a89341f379e2f7263712393c4e3f3e903497e3867532eb1279c56
z7644aceae58d16c53c4dca2b247dc8d8411f79adcedac8c3560468cf14f451a0e096e4d19181c0
z58e37fe83b33f855bbf7650e486184bb342d8a35b03b67cb98283ec2aaf3e8ef60bccdf9bd2546
ze95b22a87f76d312b291545143de60a504b83e93dfec6d44fb5ad735cfd7b66ae267b813deea7b
z390b474fa218ca6114c669760c503c75e01488e1770b22b0eae25033e5ab2bf68a851b1c8c2d2c
z20adfbe2b586305c335e0f7241664f770a04b3c86d14459814f2cc8c2d807ff75b543ee68a735b
zed7c83d6f3f5b05f8df0285278317b44d54662c9ebc9c0ff06bee78166cda3d72d8851939f0032
zc634f4c8903ff2727bbfa3ba68aca2d39ac56cf0b45447f9a4e2c2c3ee2eb1ec7348f25def6d44
zf8ead0d6af5d8c944cb4a9cabe2a76fccdbe96983e7823ae9af781653011d36e687f1353ec29e7
z87a1c3db4692e99e4cc6542334ad49080d3b15e185c4544ee38e7a46449689bb7f2dd802e4ba39
z504dd7666489e821208f9b77c239e98b8595748911f0e6f015230f664d4b09a1e9403b87d55aa0
zdd2917e336886fd9b459e82267a709cc1eea9179a8e7261c21f5c76b1163a4886975d892eedf8c
zde555ea68a628ce37185d48ae886d8b88c5328026b5090856889a05f143a64109d25c40ee8f56d
z3f139172a32b1a713ae5a561b0f0d996dacaf0252177d80afc769d914e64c930d84dbce2c05430
z4fc1949280c1548aefea2aadfcc3529ea826706c1f7d2a62e7f5450069fa97b975ff4c95a2958b
z2627e02c028a7b6d85fe26be08ed541b327a6a9f7910ac910e85a3444c8948449f893b4406a812
zbbd244d21ce8d14268028271e205bb035f9e84e33519f155dee1ffb0a9d014c9474a011a881219
z26893d688592a26449c6b7136325e437fe55ad56e538e83ac737f3925465583bbf2334ec979066
zb45c5d30bc6c64222b9af641b09c62051421e4c8047e69ee3ec124eb0537a282a8694d5dc0271d
z6c30f02c593f33d341052226f61af59bcd3f1d89ea23e90b4b87df827094b996f343228b2a765a
z189d76fd06ac2d1d191a863e655eaebe7f910ed206850fd1125f5ea134c2ef7a3875a9e880d1fe
z3360876d3f89f24652a92d849d38be2a97857f3e37b794dd551ed2d28fa08734bb2598f8594795
zda56591ae8b3799d6b84a5f2d3b26967f81da3be40cbf9d4e3f196f3aa490a907a990a77239b42
z969f1d0982072199a126cfdc51f9f4ef1afa99ca9a6239055a72e4866a34a12fdca5f8dc549cf3
z4816ed2aec9e391e5f6f2d69a1b4fb36badf9760a299a7764b2837bc17636983a75a05eb4542ed
z06a7ec39b4c386ee2f6fffbc25dcfdd4afa208a7c9d1a6e33bb633727541eba7cfbd4bc21bc3ff
z7db573d77f291028a694c5ab0a97a5a3c2b66dd3f82e429a8845f9a57092f72c044a856a9ae322
zff105456b07b7ec763c669da08d4ad5cfacb8bfcd6141b01883359e30b697beb3cf4d282b63300
zfe9e9bd562be264820e25313adc4c93f61ee4756773fdc9aeb45ef531c56bd7deed87e4e737481
ze4d3fa323e40fe246752792657ca455bc35291e757cf938788d10b5f54a9d427e17ecc67b39682
zec24ee6241901a22a5cd84f2b85592f810f183e136601c91b0732d326dd0181b31aafb0a76cb07
z2ba841d3c0f5d5d5e3ddc5cab2e2d2850c6383f604b9cc1098616e163c9a89a3707d0cd51eb9ec
zb33c612514e017c2550a70c0237d3ff581b5ccba5a8dada2b3458b530fed6aa00ea57243adba46
z119a4801b58b8fab0e10cfe3dabca4389dfe77e1e398d56503d9883491aa104e93af38d15d17ac
zd92158b22b19b2958a2b3c2f8334af33f6b1acde72d9a1d52bb117a62f25851c043a538fa9e596
z4bd66fe829cd853bb641208a0eb3c2bbbbce43b2e9e92e81a96cca66cba752694b067494fcd90f
zfa88f41bde88aa0b98d58c2f107834e21b15875ef875afd631f9e390e691f051a10a8368dec330
z6da0fa0541d731cf63304d03181b213fee25260d9ed781d216b1f15ec04731b321fe553ea0a01c
z9d4bc86315f769d14df16742543f0e099ba346428c4f2ce6973c394ff904f124d82024e942b49d
z96bcd2ca4025c168d00dcd6b371c6031b8dfc82695fd0e8db177d822d6009fd4b34105ea766115
zf72d909ca67ef880c5be62c01b9591668c38f386cfb7ac5d8cc6a07ed4810b33a84b34dc977c3e
zda546a2b1d307a57519116fd604ab47321b54a470b0c9f6eab28b134d1598463b10d865d5f38ad
z8c4aa71aa3e2bc5844e2dc8a94ab2bc3de28303e91a70b2dded84e4dbd48e458c19457309b9909
zf197ad0f3ff3bda504b70107d390644d231dcce01c2ecf6929464078e75a0433c42827fc462313
z4e89fa7e22a53051e1df76e832bf905617744909c7da58e127051dc93e9593a822a6c777cdbd87
z9eee50c0a26863de246612b168fdcd9aaadff67a4389b03c0bd632812e29bf2da0e1145da0fc97
z0ab88e51fb92f59e9cf0cd41a188098621bddb2fe28c454c58b786645fc2296f3f1bce1acf2406
zb648a6e46eaa78e656f9b1b47c461474defcdfc8dfd2cbcf978e140f7f0ec363780c0397078c44
z36b5fba245b8a1e1a54848c69537281635909420b8bf6fc25d1657bfb18cc4b5dd073441c1dda0
z9f66054c9e61393ef700e4641a83b0004a57d11dbbab9b9876d745abaa11b20e8fd95223478592
z8af731f6cf21b60502cb77de428166ed52e781ba1f4859dffde65fe5e77d4ed0cd85345879e57d
z6d4c1927a7c2482b0c39f44401ed507582a0f41418759beefca05c02a36270ca4cb7bae29f2a00
z0edc0633e30b9912694f029a93b5846747ecb6ef7073107a3e3bde364a4b67b7c720e54f7300d6
zcf0e8eac58735e8d0ff56c6ac641d7c24d5336574a2dc45498ac120187a41d851129cf7dc2a39c
zd7b06a6d91c8f5795282050549f9560a2d16461b4db7f1829a92e49cfc1d967e5d47980a30548d
z4db420868d129d0710a66249b55319e9014a23b1ce3bfeae393fc109528e622e5df59cdbda48ef
zfde8d67a783ee5dfc76982f7798616b4dfdd3e53ead2d8ac6e492c73d945f9ef8596a50e208ca6
zd4c30e6e794520937088a04be1afb684777df97a23c5b59eea1c87b6f5a2d04832ac492c5054be
z0ed041b9698fb872d67c440b4a83ec2c13ce2a6c738d11c5e28d61bfa468f2822d18d8a0d8dfb7
zae9191543f5f6ad2116c0ccceb53cda2e43b1d460615dff06315dc81d985151d8e931190837945
z0d682457c4ca94f25e06f8f8c79e2fdf1d4b529827bd35b1ce07f558cdff332840dc654b3a8a1f
z6981409e40440d75a3ee80d3ddd354c82c0520d42baaddaa91def645e91d99a2916b0581ecd6e1
zd6ce5f71997345fa5cb8bbaddfc2ce462f02299fee4c913924c1351c6f72d3981080bcf6c50a8e
z1f9ff173b8b7e58ee313166b6359e2cf948d0308c891e7ce6e5d4d4c76ffdd6fa4f1905f37b8d8
z089617f3d0ad0b316bd4cf44c487db38eac8bdc7e5c32953cab732bf74cf6ae5b60dae565cca9f
z3a21e1658323a6d5adcaea215bbf9bb893f7a7ce5d8e01c6a86c44034ae60fdb1a8d50ee47062a
z52d5fed6d32ec9a777601b4a16f955eadae4b31290f90710aa492eacfcf87d8116e6b1a5f200af
zd32af45f5466e83efdfc5636dce5c479c6e50731e853007ec49b837dfbdf45777a0d96fda74b32
zbfa1d8aa50e61d1cfb5deb8f9383963d24885172ee4bae776752bdf4eed6168915cead0c716f47
z2a89709f792558b47f798bf47f35fc337261303f787c891dba962845ca1fdf7d72966577e6bf60
z4c5f21bf04c598ed3107641bfa784f37276540d308a9095dfcb7b8907844b98271f12ded9ab8d6
z08f926f8f852dbac8701eda7782b6f11c82740318dd4e4bf4545f98f8f17b10484026a11e52dc2
z3740290f19ec6f561064ced699e6f7f3e31c82dbd51340f55985b372b37c2ccaa1c4465543521c
zef2552581833f83485450c292e0da2b44b1ec9b81165735e3dabf56aa702aefebd3982a3119b8c
z48cd43358fa26ede7505d2c8450120ef2847b62b54d06fc25086565729b3d3d8551014f427f769
zfa6759f5a5ddf95bffc858b3e3bab3057a273a31e6adcbb98ce7d1db46daa0c1460e45debf34c5
ze6ed3ae3fea602194310830598d7b6d61aa0c500dfa2fc8224672f753629c6d6559d8c65a059b2
z5da0c249e27a9c651d4330fd3c0fc3c524e31114a22e2bdf44e12c63d6771033704a7b806b07da
z7b75d8b9db7fa562a64189ab49a83d0d2505ffcae10d041d2eedbc7c7216f24be4b843d6f0ec23
z5b8e03ac0c915b96e2cec90c763d10ef9af8379e38a41872c12f3b493d415e1f6a8b763475dd02
z6a92642b5c45e6f2ec045ab749658b57713eefb190661914c09f01bb4f22ca0079d96264f3e14f
z34ff86d9d94f055350a3395328a2e7c03e9d966b037ec20cd99e20fa3af9042d47bc2c25ff6af4
zc5c0d57802eb7b676f7568d5ac4cb4af5caae7c1745463fd2762f88f058cf91e9551d7bd5ea6e0
zb0e615875bb9ea41db266850815f9d534a38bac49f9288a826efaafe237e81b0558ccf642936c2
zbca1465732fbcffa373e12a967354b1adc9efaeb00fdec43d4ac23d46470b9450d39778042c52c
z8290c89ecff372bba59a255fefbdce15a0fbb609bebf38f2a1d85694e96e2a7123e5cc4077567b
z70c00f66aeee3700cdafdef0b81946f15872d74b7c9cfd584252d8c88ded77a1d2689435e2274b
zb6187d53e30641e050cc66ffdd82ab645acad82856e29a546dda25306b1ebb1b501582bbe6027b
zfa09c55fb7ab52735ce1bc5e0473ad4a74ead0f79d51113bdf8ae08d68c28b65f5d2899eed1b97
z837a262c4afaaae17c474345dad948d1a6822102ab5404bb762efc95b95bbf559e76e353b3b9d2
z68aa747c97201e1a74a13cc4e367338cfb4a874cb0c1d86f565e63f13573b16328e6e9407053ba
z0a09044d3c0e0449ee2146fde16096bf17bcc1ef0d410e8e4571dcce07e9dcb67a9418d7d03883
z2607cc14b1c93bd768610fb6a94ebb3e0e092f310051aa296f9a62f11b29db294cf523bda71522
z3201f334b0f75c86c6bfb02b7e97d8e92fab073e1af7e23202c8fbca66ac6fbf216367dd48e854
z649fe258fb5c47c915259c0788dedb76afb552b662c9f3546cfe49e498dec7e1d33d677f9247e1
z3dc6d1e378774a238b9004f0e545809977b9276706e3a2a2a478a1f8fec4f351b4a5f0121ef4e5
z425695b2994195742f9c7fad4ac948d3b1175d6b8736fa9cc51ff24575a25fb1d6218f8a0952e6
zef6061dcb73d6cb249ddda2ea53bf834a5f9cd49060acb23b69a28a1e2a2c7db3470ff3fc373c3
z10ff934efd097a2258d4c5ac54c921935da00350f3bf7872b27471d15d2b7fd2a5e7b8aad3407b
z9a23c4a504f55fee5c1d4750489be4a744245d64ddaf73295e7869fa93b0748ad86a63379917f4
z65c529333149d2ba7b459805bb429aa3d758e96af7e93f8ba2453ed6199c4891efaed8141c6bdd
zfaae185703e5f7e945cfd7056dfd2d5157a8ff5975ce50c5cdc0e31a95567d8cab131cd9b9a610
zf90910b684ff45fccae3d6b4e35b10e8d0eebe71b7625adfb456bdd98c0bdbba1621961117c8a5
z98ff045075ed989943f645aff95ec149952e1e662621b4dfe375b7c70b7147aa41babbc4f2da04
z3e455fa731cd6ec35bd10e5bb56a01f60d6366a63eb2b5c7a8fc9fa97150bdf81c92fa5b96e367
zc188c45c3c43d8e352d4e0abac53267a72905f972bd97b6920a05fc7b9a7be86f90c16036c7550
z5543208a67ca891c596e5595b29d066e961c67a11b4ed62f37c76620bc62e89ca032b926e29210
z9b86c13ee0820eeee8c17a8616cf66633c22ee5971377b42ece2a2c4570a673594568a22b38bbb
zbd324355e6d39b3a8490f7bc38c1c8831061a3f0e6598ef54c89d5d983f47c56a8b58f434abdfd
za04c37bfed857422215222fca17935b8ace958296076f5a2d94ed112502d227e80b9bc5b5039a4
zdc7a984c956705435ff8c40b2e2029f24f5f941f848500149c7cb88dec9cc57a8ba53b436b2f59
z171566232439abf1e188a3a906cab760879e13d34e901bc63432ef6d6fa056b1477a04641c5f1f
z4ccb55c750a5a2a6b509c96df154234c9459b7b04909bc6ef59d7a7795868b7f6dd8cd8df3891c
z82f4eae41aea3b3675d54e342bf25fed89fbce9fd6dc99eff83281da0248dd5af5e65d82347765
z2f1d140f007c2e4a736f6b3a6113ea693918a86ffb7397c338c42ee885a5962f71b1a22bd11560
z7b8cbe88243c5f0967493d77698edb38595f8fd5eb73bd3868c3e8b96c588ddcb8c39a27a69c86
z5189ff56f838f980cb8834b56e6dd6b3bf26437bea2692e2800dc10ed758dd3add1d65ba2a668c
zf46e1cbcd684b306ad0bec05b9aa82a3fab0c7c0518ac96887f212c4abe9f3531d2895287d78aa
za60cecf6b448ee2c1a87cf354d61798338766efd375350101f077a253747ec164ecbcd10371564
z7dcad3b55ef309ffbaea748493895f615274117261c0244369d78ebba2d73e5042390e8c3940e5
zbb3e877385b7163e8c4ed3a1971e585d6a7448eb12a51eb06a00b1d4f39b1617e242b38bc07a19
z340077f01f711e87c92b49058d97708b4ea0c76f5aef8153fd823c25b33324127e173933ed86a5
za602f8869cb2f8a5aa14acbf2f2247ce6940d32ed823f39eec92a5b9e94e5af4a1094c2e3b8280
z1cd97b10609ce8ddec68568cfecaf4edb170e6928a4b73d638193550b30ab38ffae5897688ba8c
z3f51dafecf9e94a72a5579d0f053895181a0165d85744597b00fa6a01c986e1b363e22329f3a11
z8b03c5ddbb58d913e2ae6a97294b802ec5ecd7c1e133533723241c79b1ef0007564a80e2c49bc3
z68ace515747fb08d19d132f532bc496b95165813d1ad4fd25bd3bd34af85d44109085dfc0c9232
z071da92190fda9ecc123c5e2d46b47d2e4e2f5b8c0bdb30ee12e52db84f8536d248e198ae52260
z719ea96ade56b03598ff2a51f0b156f741b9f96cdb0b7941e3ec0543c2324ffe0809cd02477f7f
zed5a847bd76d556d5bc028a4b8f4cf637bf7469cc1fad57eff3fee63d847f9002cb6a088a6c0af
z44d7c5fdadc12291a4439d873201cdf9aea99546531b9577784d45e79dfc386ec6b46c100c72dd
z307de2e647a57c82e4a0837090371c5459a7efb71d7bceec1be31a6d944f71935b4cef7972b7a7
z2194de9aa43d85813531e693dec1fa1338b4f208bfb0782abe613d2d33c27098c6fd72a963e00d
zd809da1083d824b3aa50bafb2442e2eaba4f5dbad4c14030689c0c595e27cc4c2fe3c99098d150
z27cc83983b4f7ab7d097819002f7abe2bf12f8460dd888457147f695470fc163c420a7cc7e5e49
zfbcf52f8a921b804c146bc6e682315b693711c2c7161d877e4d5ef1e122c04a9d2ba2178fc91f8
z4fc1106b69416ff92c86a5bfdae7c1e2c83b52c3495a5d4cce9e9d78cdc03ad37bf64c310bdc86
z264ebb12df5c3faa06c35fd230aa9e612228ea6f5a8e7a940e6e8196e2e1441c6074c4383012fb
zf0cb37aee38eeb6440ff596e506c71675251460b1964adcc794777bff4bb71bdab62e40c1416ad
zd28059fdc17a18a49982cd314e7ce7f1be3bbd946609aaa1abea279a18eed74f4e913cb60719f2
z72a69a570b67bc5a596e7c999293edf44b796da305e9082c5d1c6f54d14d39cfd1f75c1d25738c
zf4759107c4477402c895873ed44f5d4bab233a404886475a21329d57337f8aa9aa0dd38677118f
z8f2124ec512318d127ceca0e7fe460c467edad2f5afd776a951539a8c8ce8b92ac6f389e0c8d91
z736aed0bb46c69b14b73ecce339de11d1cbcec3a24fdf2a7004e81e950170c94cc76705a4d6665
z6bb311eb8d70a8f3b7cdd7cfff618dcd189d8f6eda097e01cb0ed72f885575580ee62d90392ce5
z14372e680ac4a29b3e2a41ab703e376b9f226ee3d6999d164a246463c45e5b05c6473815c8dd73
zc1c823f251b00895f601e3cc679e76350ea8a26c5e1de2e9122b2ab1a6ffea7d3c0c39a563d429
z683880ecf5827b3499e21c87ed459e4265708b678f6e69e5f2b8a4b9f7575f96b56d6a38b3aa92
zb0d8fa2773ef59776e67ddf4fc2e4cd7157341c9a0d6028bdb9a92c9ff21f3c931f05ceb6ff0ad
zc524d62eab24e830233145eacf8629d37f5993613bfe4714004949986d17439bb48a7710cb64b3
zfb727bed724ed9c32e083641fbd0e92269a17aafa94643dd5f05607d03221a542576201298e98f
z5187b15cc47a3e84d0d2021545bcd039967b77aac42128bebeba3449b66c089256c08268a77be7
zbe55ac3d4e1a0de67a808f28b220d4a4f7ff4056e2a3e72783232d836c63b75c05af5c29de6fba
zc89f717f081b6e66eda82e789f707e3e89f62a7295450e898b51258daa0b1168abd4574e682fa0
zd073980c4e2ac383fe59f16de55cbe8086f2138a2632315cd8815b789764a44915ffe03462f36a
zd29dad683597f6c7566745e58542d947c63e8bf58c00eb66cb360404cf198ac55d292e4af518b7
z8591145ca4c6a518db8de16a62cff0936719bf97170471f8dca3cef61edd425a522b0d6d21219d
z975c85f92fb86bae018d7c96a12f0ed520a5d4939a6bdf00afd83ce7b87ace072db5f3969b01b9
za2ac5341899f665c186e44aa358e56543bf7997847333fbdcb3e24afc14ba8c3346dd0d09a0836
zd947810a46d4097fb070fd819eeb8ec9062c21e76ad002830aaa619110e5772d1ae96ccb279a2a
z35f46bd3890f2c3132c15f9a02a01a840d492340e5a9480f5b9e4dd377f99178960b1e1c947c38
z68e13398645d793c602098c0a512e5e6913c2befce0fa14c4d6def8faeb484f1120bf9d57584c7
z6c9c13fd94822cb5dabe577247a7526d48ae5649433d19ffccc1b264e839d733cfe0a18861cd01
z170bab2b0db36719afcf9f1af187ab7b8cd1075d607df62019181726dc648550322bc83c31dbe3
zcd3f91a797583319715f5aea467a1199bc1e8bee79999f563be7df2d6c84bbce127aca943ca4c6
z39910b2db911985fd2f95b3326c9faf6284ae12ff2a0d14e405aa502e98d8bea4ea1058b372b22
za2019b9065f30a2c603b823a36815ee12d0c9f818d03a2b01c4a661bdb7664f99c660e4bf77b40
z6d557ddfdcbde9308e621d60c8676d6a38959dc40a8506ad0902a0493703758d2c1dd4e9889026
z922d81ed9c907cd70c0ce149180da5be699372af05c0bb2e0714ec32af43480e48b161af5f00c9
zc53e8a36926b7a78adf3db415f366397a618410542de0648328d113a053f1d4d7b2b9a48871c9c
zcd9519abb9856edbe72c5d57e32192a91584916dafd169f57cd6803f3fcfd0e0921457b98a6c4c
zfca19b235f00b13c96556f5c3ead50918969b80519ccfef8b454708ce7badae2c6c2b7aa8c7756
z2b53dbfcdeaf50a822e88a443b48920dbc797500108224656df7d32e481d0bdadaa53b3a19f1c4
z401d01a0ee6e829f07900f890b7f32352d52d64fafc3b882f1b83994b3b27a4ad02b12f03afb20
z7a0b0ecc717d31afdeae9d8eb60f55bbef21c2fca9204e045b66dc4259c1e3d1f63be996607791
z9e2e3921a7c462e25cb588e3351894b90b35483166b02fda08ab82b68a24685f005359eba2167a
z2ad92fe5bd818019bc286dcda2034322c8c2ddfd24941a37052b6583aa25e489ddd4efb1fd710d
z23bf75eab83db0b6dc2bf639430f20b45625b3d53175bcdcc1953ec9dea1f0030d39b539fe7796
z6817e25bcf60b5bf9651358b77f4b45e456e33af944f42ee9125e8e2b00e50077035a388323200
z59cc169960ababe6b7f1f0b8b6d19f18684591b87b7190b479f3679868ea0dcf274276cac38ffd
zad5ef26f84dfbb23b6cd7cbf2968ea73567df13b6e4de6f2257eb6cc9fed39121ae3e92a7ade40
z66280b43b0c10b3be2379f0abba99473dcdb127e5da2edc9a00c54b3f96b2ba8e739cfa6edba04
zd986dca6998d407d91aa34dbfb3061cd4f0b134883d1bdc81b0b47af0ce7a7158db58929da016e
z75dae9f569497a63526549a63ed8b54835c00c22da921478ae00679a23c60dcd1bed557a874754
ze31e1323c9ebd73c0a9153ac6aae502f7e88b7aedeb20078925652bfb6eb391c0195330c210b64
ze716ca3c35b1fce9a957b39ac9bd59cfb951dc211866cac182302e490c2c5debbc8fb6a98129a5
zbfe840a22f6aef278080c6d224d98cb274714b7e4c3a4f06b26888f2cb6db0fa6ce7a4766485e4
z6b62c427c217521058f4dc59509a8ab19ee370f6f5fc1dc9f9a28fc21751d26749c74fe23d9b11
z9e4f26a571d2c128e4cab3febe469e99a1903ce7c72ba1230871bc3ef17fba756ac05ae8d331b0
z53ef33fa3325ca78d9b8045dc9bcb1ae28bbe410174cacbf51d039eafd6c9c600030426ce7dee1
z88a73f10dd9b0a387934dc2ab525cc163de182fde3704d6ecd86c97d6346fa58e33fb716b8ed2e
zf2c97e937ddf5a3414ed1d1df0e8a1ecca2f26d7291b45830628f50e5b2bc9b55592982a300a6d
zbf731d8661e409222061845621b1bbd568af16b9659a6feb6e155cc7fea60db950c32a0c2ac2ed
z74e9f27cd020c363bf3456f05104d0dcc05869234c4dc721d1fd455930522cb96769512665259c
z5b2dc9f9f96bbee1514b3f49279a553b9ffe4cae7465667088126cb6d44c76e905b0c3ce7ebaad
z934f414a4e6fa5a9e2248c6f15f2db6414c0621d3ab6fb42de9fc29aa8c304c5eb40250d36afe6
zbacb2abaf7e0eb2ef1b1af6da7da57caa8600bbce079fddeee812936025c354ac3e0ba0eb3fd73
z405d9e1454f63a0415d890ce8bcaa0dbf8c89143a12e13f69072175199bbcdc27e48ee76e69fd7
za6e0bce683bf8a86d4f2adfd1cde4489621494789897723e2aef675a942562c0f738b1681c817c
zfa314237acbfe1170d466916dda0eea80f693c1b6c69baa10665c325d48818ee6798391aa074f1
zb46729bb04b0fcf112fd306ae48c5e9d4353b0bd4526034b9fc7fb2e5a984251286c0eb228ba37
zaa2f067d8501e51ed68d6a40884fe06785c866d54062a98134b79fe0dd30cad72aa7d3b60fbe1a
z6c81d54488451eda5900d1843e02ee6ae57fad134175eb431497b9aa904843a0acf886447337bc
z2f5163bf9b0ecfacaad062cedfb7c5ed866af9b57a6a24fe4566eac349e9dda112e0f4e6cb6641
ze2faf8c694d6a6493569811b67af38394f99a6555d4773bef97abaddd7a494058a22a7a7fecb1b
zf1b56266ebf2c4fbee59ca65fca3f16b4a22ed5ac5287a1c582117c649da5acb4a277604fd4c69
z5546acffbe623c8a7cc061a8bd4317d8376007a458a33701e396cb9a93c8fbe6b9d3c5748889b9
zed071a7c32d5a342f9ba1403e7f83924274ffd98388d20817a379f652667b391b99eab20771c3c
z6de3a177ae4778f7a27cb676d0cd5e1b3628152e812d3f1ac22b24a7ca666419103a39e74b4b96
z38dfb208139d0fbc9716eb99f305788164602d8147acfa40f313ccc596eb9b5550643d7af30371
zbfaebd7a62a839c5b345f497453e148dd85205efe1db27c274739672f21dc9ca9f2332093725e0
z0b91dc2ecc2e7c2fa276cc10c097d40f04c795025cffe68b3d05a8305d5023250a39d7bf47ff42
z43339ef99c4153e9662204b01826b3a2d75347d1a744e8f86db4fe6899f9d79ec6cf2c88c014d6
z9124cf9827467bfbba5e516c3c1603579a7c9f034ce5fa73b4e99e40fa8d159b92a1184a9308eb
z73aee554b9386c6c804144acec37222bc284c9546eebf0bda515ed2ec8436a082491b7b51ce5ae
z46b27d9e0a4000cb508667e20d185b4572b406017ef123c95b18ffa11bf4cda6efab31c2cb8731
zf26f487d0cf272aed3c6b64f628b5dfc44df62eadedfabab7cdce20c6cd8131994d26b329607c3
z54c306846e4705c56753719a71eb0dec43421509488a7d2dcca805b952523350e1eb91a8abd1e0
z2ec396a803dce7a52bc57ad73e905ddf19bca5f88bb0aace27a9f4f9642374c882433264c2f91e
z101488a7a89c3f56f2ebc0c1aaaba6932848a7a31b4d7901749ce8c1ae3236f3a389edd98bd66e
zf606e9dc1eceab35c572b310912c08ca60ebf26f01a58dd757490e1474c5a2bf7bcc280d40268a
zd1ee2a8a18a16f6d7a814ce3cdc1d4df69b7a9c43559c102f60af8dd23517dd82633a708b8741a
zf90e8cd334458850049f62ec609c25494630f8f46fc6af005a250c6f8c71f3c9486845660dab58
za06a6a48e87e9a2322666f739d3bb1476af656b9c55ecf6a2d2843d33dba84286fbab7f5a5ad9d
z81397639364aeada14d11f6c65d5cf71720e0e1ed4d70728e2dc26942c4b1fad33bdd968689f60
za0db40430bd58f93ee8eafa72be6c06be00c08844e632db0e1c34691cce213f1714cd480c64381
z2daa08f9c5243506978869dbd71e8fddb033e809ad2a3b591e1631ecdc335bb06e657881af0232
zbde2dfa6170955d93adfd225404d593f765c9fa6fbf621d9544807f1ff10f1f76eb995ac42dca5
zcb165f49abb178f4851f0cfe3bee791f2fcbb01061bed984a94a2d52959d9b89e5dfe3270b0b2f
z0b40b1e081a9bae570ed74d266529a1da9311e09977a26a6e07931dbc7abf984b630cabbcee4b2
zde5c1821e60396f2aea428ecda131c882d61be74dd76d67873f7932ba3c88c5694374d24388567
z3613edb40cae0c7375e3c84b5b4f5b42dceae98567ac36c9600d2e0cb5ebbeb28ca3f26525361a
z4d6c2de588d7652835ad7a67b840e101d72e01958249dd145807185e004f18c3ff7d3e06d4c41c
z392450b275039fad624121560170b8d772b7b6b3b67ff9c0b539ced8f6d888ade12e0c4cb9dbcb
z7bf2d1ab912b5f465082c3b99a09d0ebc178d2af747a68032e9b78d3a27be924234775d20d4de4
zf544682b6dad424c4e4adb36982556a26e996670554f99c1733563710508eead07a4cf2b16c751
z28ab66561fe9178b594a7793c0e6fdf7aa584afe422732e13ab104a60adbcdf083943e0bc9c820
z05e585b9f39307dc009ca31ba80665fdf42d2c5abe1295b95e42099a0cd0ad8db5b79bc455faa7
zc766a6f519e43cb5194b80657e111bbe4eb131d944906d6861ce214d5a3cae07951e691e9e066e
zf2557eb035a7197b8c4154da1b899d8ae69df860661c4ed0d9bf98212a9714f0c69c8bc437efb4
zbd4d85b370e73ce0fbea82db80d3bd6a96b24a1571e8e38504ba9c3e689b6b3d1be38598cc3b80
z293cc8c01a7082300a5674908575bf354d39303786a99cf4e3ad366e9bcd42b67b49dee79cff3c
z2835dd8da8dd9511742ff8456d9fe7ce00031d0a95e50e76bc523aad07cce4ed9779eb82cd8306
zf9a5f30f9b170f9f41110c63197e793736a81061659b68c08f289295bd8648f58c6d673af8e99d
z474e1f3f0214a886871a94f835bf4b9b99be91ad002146e9c4c843c29358b210ad5f2f253a8605
z1346bdfc2c5e3f31a39e54330391200a741a7161c951ebe1efaf9d1fc88e16c5af052c2ec34161
z4f6f3585fcef9cb040d1091497ac0d907be3132ade9305556f61314693efb829ef3e881f9a32c6
z7dcaa510f83bc336632c2e5ba4c5df04392e5942f469035b6ed31bda2044b15de59cc7eecd76dd
ze7e518fad80b96afcadab53c8520f233de1439f391588d6edb9b552145411a8594277fffcf242b
ze74913520becf767f5ce3d842780326bd1aa0aa8347c4d8729d97281556d707ca651f156349f9e
z46c246d364504abee694787bffaf2ecc97220c9f06ca0b493dcec247e5465cce1ab57c30fb2d12
z133cbd60acb200f0874ec0e6f24736a75e7da746c9ad180cceff786ac334a720390f74f25a87fa
z86b48b3c8c6a4850ce5268297b8b94e93bd59d803a2de62e332a5c54664165a6b2f93a043eead3
z585b7721abb93b4e56275a5f0fdb141952eb3ee0059948ff377978c19b4075bf9215667d699812
z965af5730e3a49fe2ff846839454bb69f0250d3e87a9279702bf286cbbfe7f98a3371aff5132a0
zb8b6a4ae45e775ee2ee31c3721eb1a5ff4d7e16c0dbfc8298e9f62aeb044a7eb0d54773214d3de
z5ad6e04cacea688a39f6cef5c7b54156da9fed33ad71b632b5fa7dc7fa43537cf77c45fb098913
z3c73868c72b03f40abf273fbc7d4d4855f8776cc5cfed69cca6e47ee7f7527bd1dbe8bc1f1b6d6
zdf6f807f79fe99b04f73603f85b97845bc946d209c3081302131ada5ef6d4c02b9c1b8c4503645
zef7a996dc04f031f98f423c19074e83313d387fa9f80addfbb30b889f814c0001353561f161b69
zd13eae332bcc5897add906f04aa3ad3ac0412fb45ccbcbbf104d92cd6799045cba5fc154dee25a
ze6010ee40534df8fb57dc4aed7dc8cc90aec2f607029fc4b3d9c29694ed6bb08441f21c773dd2b
za81afce0317b5e61ab2bbd55961c3e4375ed45f81c2649ec96467876c4beaccd5a804f10791ca3
z05839e4cfc6d4c66cfc903b633b78b13305a6b70d3758ecc5cae42135634d33a1822ef2fa0a6a2
z575e7050c716e3ab27202359bdce7539a803c3dc2fe5f1f56bd82a747d9306aed7475ef84a22ed
zdb7cdd24cae08d537ba44a66fc76ef4cd5f4e057d7927870153b001315a459772d0c2f0a10dff3
z2dc0d263232c1cb6847ce36acd6ea4b563e4fbbc02a5773768267363e7a61b0a9844ee98039d45
z82a7eef4800fdce3771ff5ee4a94d354e0dbe1531112f6977cee97f9de891f969d08eae8ae926c
z40e4e00b7d9867eee002b8b62956ab866b7726cca25034960e3d3f3324028507457fcbcab12917
za6207fa92c09cf450d3f72981a02e32985fe185fbf883050e7fd114ca5aeaee5df65668525b317
z13022c3960d5b6bdb780e47201103175463f06060f5cc3f76fb21ec1f5ab77a44e6c1a2191e5ea
zb819cfe866aa2993b244a112aa4cbc6cbd6ff040256a78bcb63c553545e7d5dbe3f4365499f7ef
z3d1548de663b44dc9d89db1ca8c93220a1a9d3c19a5b41420132c38c7cdcd3543a1e3eed23ca2b
zbd6971d523b749a19ce5c17aa61c8d6949b9a63d165a22035a03d56a102d711a6586b054bdf880
zcc7425184c68509f0f8d150d3bb7b21447a900a239117dba1887aa7da84e03a863c79ec798ba97
z045808866f5e99257d06ea097780f4b047c2b965b2f5f2750b6f1673b3f9ed3c00b365ea0b0d09
z7811ae152a9867c756fecc75e569dc2ce859cfe3188abc00199b8b50e40bc225fc61ba51a42b97
z1adf7ed2ad3da2fc781fe60013236d4cbd97d2d30bd7eb9e1d43e3d2ed8eb04066e09baee38e2a
za33a3bb8a30cd87f7f97480ea69a777d5acebaae3f673e76c6d6958828e4f59cfc282c37b0a651
z7540d806bfccfb51400061745c30b7f7cc2f7083674f80d8141ef468ef7e3e32c17f5a762826be
z58f8d6e8cb8b70ab5cb4cf249235104f19c8c4221565b5440567e4480323da44dfef0e78135deb
z5f88ca96b4594acbbdc1b8905c6306da430cd8b485ebd5f6f71b7d63f58835a31901161c5a130b
z6723056ece20d95edae045b9a3e2a058472d28796ed7b916f6041f75de072ab71971d805bb0ce1
z67df2fa869c717a4697fb20ec237a61d454911467a5e6e55cb618b7a0c128db757b05369005a36
z731f55197e24b59d3bad127fdedd17925f748aeedbc7668e1f1deff52f22bffd04c152b942750b
z948a0a9f9d6b3f9a5b308519eb4e18f2ed50c74ec1f3aec4f305668155f6a204ae6409af4ac4a8
zdd6588719c021dbc4987c2c5fca3d343682adcd82f232d3fba69552252f94885f94cb63ce6988c
z6babdc73d666f938687607025181bad728ef0c865b51a9f5eb9d707d583a06dcc135d6031d1661
zc90029fa78c1bf53f83329b64643d49de9fda511b87f34632db89e0e699e8f9b1f60d3d27e97a3
zedb42ee2c5667dff2053e5529ae650b9f58bfbff456720cba03cb21b9733942df94b3e55bd384c
z1163c780ac735aaf69feebf435a9ada22b4d0679678a48e2ce1cf4f9fadb9c0906fcccf86347a5
zffabd6debe8b9e7456b7c4d1e4afb218c3a5cd8820e5376663f342f7059155bbbd6c78722d75e9
z3bd92f7d0b40d57ba7cb6170eac60c0cee88bf637ee4c580f78c3918f75eca5524a09000f2514b
z194fb8ffdd1b35b468af17bb230e33694345f2d0346e8967f655371b154fa516f993606030b9d8
z2e31141d66469ad6a16db3e5372d206413c5e0106d0cf9df692864d6bfbaf432c9d643250cc642
zc89064dabd7b5c58b34a2ae2beb9574b1521b4f4bd8f2aa7e5a03aa11b2b92ec0ae7254c5e0204
z3506769bc11f11d5c93cb8bae3be8856e1fff41196c017615b914d0c4b283ce1e3d7704cbea3ea
zf69c4b9bc8fdb48b0fa7cbae24ffd744819cb35bd1d171064eebe1cdc1c01901f14e59e8a2c954
z45fee6f1696be9fc170b14f78a21e45d9458210499661326d91056c49f03c11366896a21a1e813
zf4dbca571ca9caf8e7ac429a9e8c3d755a9d306460642ed423f3d3bd2187dfa2617ad13088bf49
z3e8d7c826872b3647cec9dd77f0bc7a07ba2806854286b870dbd9508404a2430eb62de2c050f68
z0ccc9e72c57629667bd05301058bf7ae00fd3c2e8f5aacafd4d935cfa8ad73399367e0096f90de
zc112e2f1d953295a587d704365bc71585a8cd40496173c0fa090d84bd4e6a9e41fdff6803eed13
zbee3c129359129b5123088b2454c3a19a199ef214be12daae15eb6e1a9d39d9bb7714f99b1b1e7
z4056d711b182122ff74ffc3494d58048301bceba4f7c9c95acfeecacce4e4935b17cb72b0f3082
zd9be077a4ab0d15ec3b6199ddc96c2b70d50d0d140d1ae5395f280fcd7e77965ba43550534c5bf
z2de48edc3a6694aacaa90fa7160fc91dda05db1c3ca5ef017cea25f5b97d8137a2d85469e78abd
za6acb794db98b18bf69a3804ef1dd4bf9c7a694745e114289d4dd599cf007acb34cb3ffcb5f146
z8cb69f4e0decedd1e85519c23b8f880cc7cd6a875a5a6a4909e0ca7258881484509e34ba30cab6
z32392fb0e6f8d14a29475fba95eadef4241c4598f2c684408dac9e010689797137679828322666
zd04bcef3252fd4d037ac13c2fa2456d16dae5c203814aa4ed85170159b949e2e4f0bb5403f4367
zb9e0028f16a31c2ed607ba520b233efaa1e948da81937e93711e08de590314a9ac7b666ab6f7aa
z746a6371c63d1e57e593f1318ac8b439171925c9062a155edc89b18c9367ee471af78fe568ba32
za2b9ca6b1693a0293af7c4fb03baa6cf3aebace50082b64523b8fc23e566c3435369ddbbc48153
z7c4c4e2c17c463063cf220d4f30880d5bc77207beee5950ea886769173da66fa3accbaab321272
z0de62b0a115bf6e1a7c3d8ed05375fb5859cebefa64b86640af800bba12502970384d62a87c23d
z779dd65bc6b49f85b2e505c6142a49391970164d3339f6d81da342916d9f21592c7664d40c1c17
z39ff286bbec443b687697b305042824efc6f218b2cf5a25ba280e257c16dba13402b84c4af7387
za34d5742a050c0d9d3b32b994b766a3d63b3220e6743be9a3c52d1428c65b74c046c5a50fd1dc5
zba4a90df21fdc9a85fbb4106ea1a28204e3db2566d68340d3cf7ed2683f87fe908f6b95f80b290
z7cf118a8e05d99e8b83434a4012c9cf5c2d8208b8f37601551757c9fe9ce86ca2c5d87bbb0b7b3
z2ad07256a481e15865a58838cfbefd4df65fd13f45a9cfd749dd774f68e3440eedb46ed8521674
zd01b82afb7564fa818284f4e0ff0d69ce434fec96eeb2f15fd0255a73ca98bf81bdc2d65fc65b4
z4086b38e28a44469aa87315b7d55cb8a14a8de2cfd0a114fd2e107f3a3486abcb71f23618aee7d
zdefd6de9a31e1b2dfd2c4285120825930dc91174ef0eb788b55e260443c4f3b0d30ce28606e98b
zbb34fa5451ab0305ba5ed56eed6c6c4b823b854b63596163d3c687914a933306e386657dbd7165
zcb81862b465db6e7464b29154e7896f8ede3d89acba78f7f15f650bf9c8f5705c158a561ebb35b
zd730dc9539089fdc957dab48109e8b8e817325295f963e5ca330c6291b1ba96e0b57b9a81f09e8
z994c05856fdfeae295f778afcf70f301afd51f9dfb5ebb79414f49ecbb29725d5c8bdeaec9faf9
zf857e70274be4e3e198aa4e9c0a4cd5ada6339a92ef08d1a126d898c8decf6f94e35c0b5cea056
zea0c77ac2eaf8967d602155bccd732b87e06329db70bc7efa50504c3fc9e74d4cf9623defb4b92
zcad2dcf46323f0bf15786244216b6780c1a1467fede4210a83253b57fd8e8a5c290bea235c829b
z1ded341b2c650457a1b27cefc90b485414f585e7aca39ca7ce86479523a3e56a8695a12b2fd3bd
z2f6f8fb79c17211fa43e626f59d1df88d05be5d3156bc5bed431f7a72de3127df7b6cd348d416b
ze0e4c1e94b51d4a2594235ad74a6d49e927586c87f2d1a82b7f56c872b1225dcbe599dab908c23
z6ad7ab4920fcd13e3efe578baedd92ebc6dc6e455acccab35689056b0a849a3efd2d201c46e7c9
z80835e2fa335ce4fb1d2042d82bbaa9ca24755eea94fdfd6437db2d8d47f65d925ab07be1e769f
z1ca6d446995d27f3521d2644b3317cfe5bc82a11afd47300b5412cc077d08c57f01d7afc925aed
z14ee8b779c00ea3627dc098458273afd38742cafcfe13b0a3a6b138fdf2c9fddb52520cdbf2c10
zafb4b8900362ddef744bea3e6b61a92973d133b7206f78163676261d119c06482b5cdd88af4fe0
zb2409a327d34d632b8268e3a9950c62749dd562b61ad600c2fd1bdbc83cf0ce11b9c0e23364df8
z38fea200c72ce8242e7a6e9cf2157014a0a99776c3e07f4f240ce1b8999b89beb76b44f9d12da4
zfe80355c70b99b0a3559471777ad77bf5794b495d6d81499fd77e9379a0ffb742a3e71b8f8be9a
z116a5b2b2db6e0d6f6e9af6eba374c29cd343d9f026b3e6687b71847d75f4656c2aa9106d3f630
ze46511c0968c5f0b4e3b7a843c89e4940c710d4fa1703c6eb15aee55abb0a7be6dbd9117eff680
zcf22d82802af4b07ffbe70eadd3ce3ed8f27197732218eea2337fa8e8010b312343b7f3786a12c
z9db0cba9cb1976fe80a224654adf74785f7855d593d0b335d948f457385b29451c6d39e8767308
z8e25737e0f98935412ed4199e2fdd6d08391d7efa34043a1f98e77f35fcbd3be5b741787107d14
z0f01ff6ce4bce64823d2983da332133d1e8d587f47fe1e137719b6927b98822930cc90accf441e
z14346c0179908705291494567dfdf95812f1b6fe85fbe9a3572c855b0133b89349b78a274c7a4e
z625c2aa9603431c3be2e2bc1d3834c74c1d28f26431f28e0d311ec956b4004e4ad0f79a064824a
zb8327f670b25410bda499845428895a7d3fd93e7612cdae03c81001d56da52f325a27347ff4576
z90186a7b29feb65765ac1267a4ac1ce4c225ae330eb55024dfa54a94040443585b0b839f0a7972
zde058e08ee2637c272093b32b01631c2094f3004f1a57d3d53f39ca9a2983c947597ccbacafde1
z9fb55fcea9ec955333e0925ed3ebf20271489df032b84264f00b78a9613d86e71d7000a640565d
z4c8bffc0429109321385ac630058492287f9635b83a4d984629187558493228ac68bd1c5ac3a88
z49deafbf712d099f00e3064d564976be9eb2896a3d6f61aca2c9ffc099600d092a1f43b6140a63
z568537cdb9157d766b1f658f9b7fc49c846655c94b390d1f77e02e192b961213d42fe1d7a0f442
z48f49438944d0e1aee7a1d1b4b5242e4c1fc50915b8e9dc3e8b93c227b110f6b2d7b5f985a008f
zef100569c4002da21f03bbfed823343eb0932f7dd5f51d729ab0d99d9c3dd62f22aeef23d84561
z6ac3cfd8ebd20a8aeaff0b9d6382394912dc65c585f00617dbc3ec0d73053778e4f84b93d26181
z4fe9633641b98f03798350b1c7049041feaa6368373773e0a711cdbc7ff48e425e61251ac429a5
zaceff5402714d25709b18d45c4d79fc849ec21ee0d4801cba8bab3727b8543d5a159e56fd4543a
z2593af89f0792a24b36899edbb03c013f063fae84cce3b1729a4d8eb8b3d998d05ef43e2a63c38
zab1df7c59e5f9f3eb5f31312c3e127949828c6ce38a7ce51e1ff9e2540c8692a0d1d4d4053128f
z35c6ccba725594d404ea24a59b439290101c488a3040250c404386a8a96baf8b4b214f5aa5982f
zccf9dcd16db5d3d64ac579c8d9fffad1fe76508169fd8aa31a40e8f0af43fd9ad2607cb48768c0
z35c8661e6b8b7be9117310b003d9c321de6261e37bff6c092a035f651e7eadf66132bdf4fe888d
z8eaef77043c8443d30f80907373e53e3b2ef84080742f8e531be08da98af9a1e574e6c8c93e309
zd9c911a37bc91148021d140d5748f6283e67a7eca42fdc4d2b19e05ebc1ff7e39712244b7b90ee
zb44573d1319a4a40b806a0d729c8fb9a95d7de6df629e29e9811796413608d6647646bfeb03e10
z3e9f237ef726589ad483a832deb1c0a6c7de77a7f269bf1f1e4cb09d838abbf473f627ae4e784f
zab4926dffef500466b36b9089b81451ab9c9a9d3cec29becfc5c9a553ad7d93c0825a73f158cbc
z41eb7a8120e20b411416e4ea57be7dd4c86985db71ba7908ee9c022b15384c6ccd5b416cd4dbfb
z7a3697e04e2bcb09c149a0e41db2ae4ca61234f22fc2e8ebb4248873c7f0f0ba611b8f6346c8f7
zf4b680074d670bbfb3a5d7513d88f1fa9726d8f8c385abe45a1fbfc3f22c36774cb3ce7f6974bf
z6430d0633356fe43f78d351f6225b12b791c49fec6c0cef9943df582011dec7b9afc08473fb449
z413bcfe0e3782381d6b9e42fd13ad37759702862b4721ae0a8216fd4c9ba443ea21a671e5b6caa
z0c5057ebe574db651eee3e768be76b9806030c10c61efb0d2db6e865ccab2ea92fd65977eff35a
z0c87266182a04bc1680cf39c7b496869e10a4ac5a4cc9e61357fe9d80b43f41dffdba46dd6889e
ze9b046161af6c0bf722a88011b8be50ce8523a8a4acd5143f6957cc9e7c26bb14ba7fc97f685da
z152788a21e76a15af12f731967ab9cc90fac09d2348765145883ca4b447b6d0ac1c7a828191312
z09c80886eb7e0b1071375788353c050cb2c0b52adec18df364eaec05af605499135b54cfab9f93
zdc0f18dce7d7afdacd52404ba2805201d2ba8702e7bd0f0e778b31744a656d15c4f4578c5d9e8c
z8eaa735f9acc633a83a2c52957a0bc3c6322a330b00f5f62eeaf809e2288a08826a90a47c1485f
z9aa58f764c050e8b3a2cd562ce3751ca8f20bfb3fdfcfe1d35b7fe530d6d85f87dcf697947e44d
zfc86d768b8e5c0f91f3744c826634b6f8c201d4a658f305df2700312ef4d27695e0eb4b4ec19ef
zd6956ce7d420c214c2d67f4df284ac1a4cbac4243be610463e8f315405ff2b32ee0d98ee6cc998
zbdf88d59cd6c4f9b00fe451f912a749f6df74374d00e294f0a08516e1c936734fe14e69276f066
z4def1dff7855bdc598a9892c0053280f04a65f9db0c52b02c2ff806b4a1035e7ea392364001fa4
z94dc8e1547619bfe64fa6e79249ada5e5ce65d201f6be46796f7c8ee35c2cb9cb5c1f53d3bba3f
z8be60bbc0ee0975decfd0c1fef4efe29d74547f7b5d8d142c986e5020b8b461dcfdd71fafc7aad
zeba9d48b8bc87e52a4b004c8f7a03d7f405093c3410ce07355af5c93317b00341733e77273dfb1
z4f6dc7a45eacdc1dbf87d7bdf258fcb65066b1aff1ab0799ad43f6d5189df6d28a729cde6821a6
z406529faac0e9307aa545b8fb96e5a9273f9f1113d40fbb3bc3bed12604cf79eaa78b3709b3ab4
z887d3b575c7282d738031c247137436bdc02b67e1643089b57a07d6901d66d19e0cd49806f2d5d
z08f56739d41a080ed10e8700b59b720c6b010a1d1dd6fe1b7f19796ab8cc6228d8c65efbe61f54
z1c8ec3bbd33c602010852789c6e74feb69ef8b98cc998574c7c993f5e849eef2f15d6f5fbf04b6
zac1ce01ff90627f7f2fde10c372cd4dc79cb9a4fc4f2aa1827eec2ff170c32cd40aaf0f2d44936
z2b13ba1f559d32e244e2a0f833b73196ab64b12cbbe487cae025f21acacb056ea83a18d28019fa
ze0e88900c4393f807ee1fd92d2bcf5cd66ec00111606e5051e85ef8aa9125b58f40e5da40899f1
zbb0e48655909415b6f5d8f9fe2c6fe2814c81a5e14b4efb564470298418df0e3486a313640d085
z26246225d1459be008a84cd561e20c86b2509f2035c04f8069049e967b8b90dfdf8e50169e79bb
z15dc11876c8ebe63bb5af7610c4509e81436a1dbad77c8a2462beabab049000f18f9ee9d5ab4ce
z1598add070f1c719e013c9ea0b431f0229d8a29ab97c1d6ce9493f0deb68f3edea3678adacae1d
z2584366302078cb78410aa375d048da8977f70f3a533756acc58d990e9f4ebc3e0ef31ccdf9a17
zb45bc89679824b88d160a8299458ec77cdb1e40038a8b60456bd522e9026c4e9708958a4090965
z7031de33dc7cdc8937c3a433c6c15dd55d588c552b622619377191319aa80846cfcce175eecb1c
zb2c8b008fca8011458261644012fd5bca74e1047e60ed3109ba3be045c8ea72555351b16cc85ff
z2c8dbe2fa9cefaede525e7d37ccef4be2096e36d235861e74940f9c167d2fe2d043c64000bc88c
z3f6a5405fa43cca1b4ad104522962a8832f6172e36e418f5396b259eb4ea08beb0cc4c14b08e0d
z5a569a4c2a4c56042d736cb85565c8b8de51e111e9bbaacbfb628cb08748f45bc5800a627f6cf4
z3f1f01c6676a19ee376169eb10c7028bcf39b968c6f6fb97b6e88d0d44166dbc33e98e01fb25a9
z847da110e4311cfcb4b9543ae6537d303d934722f36acb14d7d8e65fd23a540aee2e4872c75b5a
z7f5c61e4cc0289838128ddec201e942e843974e7a671413c50b5d1c9f88a073a0ca6f2488f04f8
z39db753e07f1b0cfd90a437a92fe14a1e699e29445f7f56e2c011fb72ef5b9a6400c67b91d248d
z2a9d17dca08b1e539fa7c9e681e362cb7f005eba8a6d9b7e450f2fe428ecf06b69ec8847999ea3
z9dc217fe2b3e1c4cd12ac3d1e1065d8f5528feee2febd92c6c157ca41fe1eacdd704343c710622
z68339136327ad9a059cff2944255036fb4fac7c6c7290af5fa2dc0f80f8a739e109e3df10f9a93
zad4dae1670d067f8c69bda6222aeb2db41f7118b1ddbe7b6093191cbc3a9570e38860052f94bc0
zff9717ee873f6f90309add84234c70f1e959bee7b1ff613f639d4786f45b7518a3ce0b0c055510
z25fde9cae70b11c4eaf907f0fb0fa09c7a57c4fb03a347081fab0a7ee73de7c07a13916e579894
z9d64b523940c5acd606eee5d6970d8e5c043e632225c9b012473f52f6e223e5d184d019342594d
z1d317c68511edba9b8f0dcd4cf70ccbd10e8076dbcb5f70ed609d9f1ac08dc5307fc7d08bdc355
z4327049d6cee58a3edebb370e96d72255148b41bbddc00d22e55f965855a35da0ba9e20a21e91e
zdbbd43788da7aaeab3deda5e35af7ca3dace174b13ee170dbfdd454738667bd10fb0da09b6de7a
z972931cc34e5e5c77cebbbe769e49584a51ad25ff1c89a8a36b6340bd5c485d05221a0dd824221
z2e75af1f6493763baaf0078130809e9ade5b09b33079496a182e62f7e9a69e60a5a25fdf5268a0
z70ff89691358cdc3faf734add5d34020a5071e15afa0f5a42bd5f7103666532592cec5d96226a0
z8bd045d853f4ded9afd4e52dc46abee0415486d609569cb09243947ad55645ba34c28d956f61fd
zd1b2542ba5ed066f524a6856005d499dd0a31ebe34864cad1abe8b0860e4e4650fc28b82feeb26
z0f423ce5d93b050cbcef777263dbe78cba7584c946bc5e35c1fc7fc0eae2de81ff7671709a6689
za3b5df69fed3009cbe63fce47053e81ac678d1fe5948d75311e9d488516807193646b9b6c44cc7
zbf4e2e9dc53f1ce8e060cef30d904af56601bc43fdd6e630aa0a7c69b011114b6abb6bbce2b534
zec5cdaeecc05dc320a114574b2f5b361eadafef31fda6a9576799b3d4aa6514bdc239d5eff7211
z39a77d7cbfb4ae129cb1bae9689234e2f1641602b05d56628669bf0ad64915ebf998935dd32e2a
z15c48d495abef744501ddc8ecf422c0c832d58e1431193e4dd38526ea3715b9e7a56a36bf790c7
z62b39c6c803bf5904d93e1d478c01f4b6bcfe7676edefb449010b25e4d0ab3e4dd19e6461957b7
z939ac68090dff62b03fe70cf7ebb5198d9b65fef6fe7a6956c4214ed76970b91b1be5403c66617
z9faaa6d8815ee2fdf8fa203bb94048f068cf791b876557d88ced2d4fa3ad9460fab68ab9df49fb
zdc35e9eac0a95dcdf22261b14080dfb18fdd2d92be1825bfeb3a88d021d288f36381d3df275c67
zc677c0d735484fb7988577bee60843057a3c2f9575cfad4ded68ca490fbbf7e01efdff5a6b3074
z7e521343cc4fa25f6b9d9670347bc4c7fbd7fc60c7701abd9fba266699c9a20868de1eba739704
z62b25332b6ccf1d496b76a0f4aa7b2e5b959a1d66517a0ced9f930745ea60588a3786b2519af14
z0e96ccfd247ad0baf27746ad5ed7c35467236736bfb1829741b6f93a120df916258ac2925f2156
zb58449b3837b0d7eda2b60d88ceb7a8501a13078c324fe60d11c2e31f0910f90ca4435114db9ad
z4bb4b7f3d3accb301022a68a0777c7d02191563762ffecabf9eaf85765250fbb10ec1efd25500f
z309cc2fa8803a9fe45958f3873172b226a9ce6334fa23b081024738bfc5b5046aae5173d699aad
z5ea0f56b4e8736675175173ca26061958ae20156d1e7480976996f8097c69997005fab9d71d845
z1e12daa3fa7db820b2e71ecb1838e9fa90c034df9eef9552f97ee69878c88b03f25e0e63536771
z5448a33200080401646e420b745e7a246bffb00e2cb9686a559cd1d0f4f21958be1ed4573564ea
zffc493b0544f2428ff7fc58190e932d9ec0da05a73afc9f35a50c49617247e2f1e47cd0413e316
z8196403b137cdb63d5861d4dc6abffa992f030c5191043ffc20e4b926ce2891789110a5f7eca91
za822ab43f1334c5949444f4d89ffc83cf160560e7a0ffb5a8c082c2952b1395321165a9bd3c3ef
z2c0ede4708f66c53d1212af62ed8768fcde082cce15dc75a1f91746701dbce384a603ab24c39b1
z757ad490effa43dac32c674e870d4c5b1bab05549af257b86bf1fcbc1e225f95c02eeea373e9dc
zfd0bd8f51578d21a18458bd19f879c58dc873a6714ccde6f06b9f664d670751bbefa10415d56a8
za2b2379a96849a24225d7a2a92732346ea2f8eb2520315594cde9c1e264ee739309df5a681bb2f
z152a5a9f113bce724d3323db7e8180338beb598c1a949a590c5eaef1f8b9385a1b3fa7f6919e54
zdbb475b7c66b88d53103760f3fc41bf78298c57907bbe2492a32c44e205900a5b83e1029e19cd0
zf53a6e3c6a09dfb5fe5a59211c0c13e6521faa2a349966cbf1e1485d27d3d4d8d24eac9b636cd1
z8d8c5d187e1bf1e5f67414b2240d0c979739e4a2735b8dcc4193bd3df99d46a5eca3ccdd9d43e4
z8e99324a3c8fb6899dcb86fa546f4051d99508eb313434dae5d0722738550c30c27f130576ce92
za3b509cbc81305f5c2069dd8cc93a89606c0a6e00d9c4dabbba27e5ae5e0b1b9dfe101446067ee
z98dce6e6f7fe2bef7e622db4753359d737601603dad2bdbfa9987328713e4a9120d86a4497d781
z7fc6230ae0f9e7f828480cbba58522bbfae7f8f6ced72cf7f50d473c5a76cda25f0f3173786b37
z3d20cc168bcf73e97ccfd13aa0bcef16853fe1bb390ba48b95f28bbd01b8b56ec2ed8d93efa5bd
z998694f7319ea23505b332b85e857504ad2f3af4fa071fd9d1b22c0ab825b804c2677a926a3c2f
za754958646fbfa3b361ba6a7f4fcfd28c4ecac8067b9923167961564b7f420b4658c279d2a3968
z58bcb27cf548e2865282c1c2b61323a958f9a086dab996c4bb97bf2bca3a768b69c54b2291b3b5
z765b5615d5759c8207263001f8b079dac9c4b7c8d1117efb4dcac36f725f6a67b1c11582ca3f0a
z6dcf9d904685bc45ebf3c76e417289277f8e19b4d3f7455115d5f8f1e72dfe0e4d1a10ee5e6a81
zeada11662ce8e88e0bb7a80b2347e148ccf7c84c6a366a39df41f5792512198fc8e7c231ebc460
z6baaacbd13bc5129899f2948a0a3dcc1a795fa733f9e7fbbbb5b88edb830c425a2db5a7e12e76b
za0fc9a688e78973aeba2b4781c0959890115d7698d37e85ab983aacebc8861edec1d3037f29c7c
z3edb3238043eaa646d3756d9a066a678462b29a5c3b2ee07020a18e17e264e095dda8751bde85b
z63923d69c250a75fdea7da2b05fe4cc27bad4162b13d9246a537909beabfc03b58f6b4d9fe8f9c
z03425caa1104a18e36baa4852d3fe9de9a1296d017513176cc590e2ecf2937da88971efde06f0a
zbb6ad00f51b7448ed292e9045cc8b07b6906d4dd21c4d536a23d82f5061b4d39541c00ab97d6b2
z2696d74ad4ba839d95f02294efc30ea4f76ffa2111f9df3a91845b7484dbf8910661ac51f83ce9
z6a9d504e78ff65f0c9f48f469edc53b28f485d16b8a8f88d9a8d0294cd61e825f6409394a38ad0
z5747b6b47bd5c450d49eecc0b602ade97a24117794d07dd976314d2ab61fca5d3bcbc759b57b64
ze24a1fb4df3c76ef843c1bc7d434185f7956e13e08a91739f402d2fe18097fadf1da4f645b00ce
zc97f6c4c042139a4dac68652636b74b30404e4577cbd8a69ed380840e046eea43157ef61d68ebb
z0c8916241d8533d16382508a564f63d100446dc7d1ebb1d21896db4027cb7d8bd97e08358600d4
z8c4ec5d363f702322ee6528dd5c9e4fcf634f3faeb4c65dadd30c9673c64a04ae92c0a6d16f3cd
z02d0a5483c3595ff091519c8cc197dac5be8475f7fd02782742f5e1558797a09631c7895ee1299
zfc80717ebefdeb5688c68e42c23cad33cb66ecc5c034ed3655e3223c359a45b3a79f4a6901625b
z55a71237c20c21c80f11c5cb97078a119f2d66ee59e862d614d8033c5adaa07b51552c1e715a39
z7cb64afa2d8204bd3b47b76965b76f747de730ee281d8b526c1794e8a4dc43f77d0bfe8205a530
zf26fca7aff3f756a46d6a56632c39173bae5965683a56fb14c0e61f3ede5ae6276c3a85f27abdb
z7946b1f617ebd0a5756b5bfb6a3bbdb0b711e5df7576d46a225048c5ed1af382103489760a181c
z2cd401a79601cabaef34370f3a7a577b18652d76e892a1f1f65b5eeed7e12e8a3660e42d84a03b
z8d05089e92faf8f22cecec8dd25c33cd56dd053febc27db3d9b43789af69de687478125e647be6
z2dae9ea425ea36303e059ef5ee995643a16e92e83b329bd86caf3a1286f69167bad078b4f29b4a
zf783eacb80263684dc6e93c40bee465de64589c1165ef22dffabe19970db65be5d2c1b5616b9e5
zfc758017d322b39a97444dfa5ef4d0f2322994ef4506c5dc2ed68e8ec2231a31234538cda3dd10
z33235a6ab765e02de6f622914eb6d83aad48b4a44d2a063b5f9f2d95a1bd80b7d25e745015bc0b
zfb91b908fd6619ff25ad30ae46883948eb3da84d294ceeda18c4c5578e18445715c77602a5c683
z61dabd33b23bc50181f02c60b36a08efb801f67561c49386d50986a2c6ca4885cc11f977c5da22
z6d9623cf8d7ea46a780cdd4f6a7e2e284c1704a7eaa5b9d22a04d5056fc29ac0788e86aec092c3
zdf5a3914981cb6209f0744f5d14190f7ccdc5300be10a1a3903529867801125233e416ce738622
z1f991fa2711c417e63ff0db56c263f3c7f700ece2c8460ac9dd5eba926d17c0328ed888c57f9a9
z2dad0728862ed779051600503b87bd908610ec393bb74530e22e9fcc7f9cf8aafdf97e9b54c779
z7fceb62d337405cdcd310adbdc75ea8ed301dd278b3ee54940434ac16baea3daaa50b6518d0b91
z2c29b58e751a0e3555c80dfda83b7611ab3fad44d60e5b34d64229bef20822fa5db71328155c9b
z2532013609da1dc1dc1969cfd3c399aefa84a757c217e057f063a140b68c7e46ecd51f6036c05a
z57b9341746ec0ca3c895db5c814a2372a3d0124b9c627c3ea077ef9d91fbb5f90c137834deb254
z2803c210156151da6b3d733db328aa516192c9e58da2467e483052a2fbf30fc180290083202ef8
z322de04af036320e272e67dc96b0acacd2af6f2637c2c579cfb0c3bff94d4ebdada3a54600c9cf
z7bf459e065297b3aabe99f6b9cd5e593670ff971da98fc34bf35e3dcb927e0fcde15b0245de01f
z372e9f54f15ca7b15fb191afe57d7904c4afdafc1fbff1f8391ce912e176b923cda06393a374f8
z41574ceaed559984b0600c089270b2c62e84f4290ea6e8492c2d11c123e2d612cb3c83798db87b
z876fd4cf2c541b0c8971b4a18979d5126932065c49ec1c242f216c877c76d8e8ec9cc649cf6855
zace72494e4962ab4a541d486a439577c033e428ce0e6faffd67d97297d8533cd891a42698030a4
z872c9579d71a8b14a6f698d8647953f58aede231f54a4884f9fbe864faa5ee7ae76fa5f1acbbc4
z264bfd1e169ba4c291dcf55c0d3889ffe3acac69e04435b5984a5a84392b9c3ad8500c95935958
zfd36d837143503b4c1
`end_protected_0in
`else
`ifdef MODEL_TECH
`include "qvl_crc_assertions.mti.svp"
`endif // MODEL_TECH
`endif // encrypted_0in
