`ifdef encrypted_0in
`protected_0in
ze74c34e226135848fe16db9ffd31815111b6d7fb642c521a3f628cf6da949865580b22efd062a7
ze90adae0e65e66a2c36a587d0a790699161455169ed55a01f2084f11770a774ec4c588039b380f
z6de9c5084882a40b79a175f5c2114b2b6d78b070cb806e1c0aa9258297f4687ab308bc470f0040
zb0b1de382961eeeaf2e279e1462520fc31c119af8f2b214846f56c2b3cd2eadbe4099496abff18
z15cec83ec4a77b868344aa20ba7360908f5c0de2a79abf8b3534b883bb12180f68b5d4beb444cf
z3fba8f13afb0abfe8fcc4294810f75afe452434d2d0f1166236c82f76edf1e12979f04bc35693e
z32ae028996dd85737a8f5adc1ebb94f39c940246e887647b64782cd7ab429b0544c173176cede7
z01dfb26b1f73408344a52b7e1f117f12bb9c8077b34876c2e6fdc085981637012dc9754765e1a9
zc512ce062e0b8fb16a214591f5c81e1353b900a611fe1f4886b57940b41b7f2ce99a7b84b04b90
z916f717e73bd10589c81e207ed77ec660a8cbed5b487fa50acde1b055c8870bd8676023f21ddcf
z9c98cc47cfa2d654ff1365d1f45035a045a66c5dfa8279050262529d2cac9e64fd27d9c7de62a7
z731bc808811ded9016570962244887f98fe5440167bd0088f2f049df882af501358497c3b28776
zcdc5426c7f52a851c35106bb93e16fff98478405cb2c034d92a13b0536cf592c53efa2bc42b272
z5c52ed0dbb9ec35d0cee158298601da1f4ed68fddab40fec79905f12dc96a8110d8da442bed2ae
z163a3ad607d09d5a631332004ff962ee40ad88fb1ad2c6bf195702b896261672803134376ccec7
ze5247175339dacfe422e9e4fbd7d1adb9b57a18dbdcbb3bcf18f5d8846ecb4275215193ceb22e5
z8510c5b0421f0e057bed7958d14a606e5acc41a1afd241da618b04d639e2b2e5d2924ae18a186d
z74c585fff3d6af936dc334e2c0b0c48800932f6d6318b5d409771391101f44ef4d596e9216a5a5
zebceabec4799c93c3330bcd108cecf3ff9fc7c42a31c0875744f98e462b1e7eaf7c65b49328cd5
zfce1ce9ff4f40e6911c4a36bd8e414affc7016b6782119bb4f877cdb407d39402d4b2454e63108
z3254c1c30cd7d1258f48c1ce133afec518c9070d2c6d97318d498c218595b2711f473c61743a56
z9844cfc2346ba2148de1d537e3ae2b6ec18c8de44c6219b5abc7a155c111de7960b8df96f320ca
z2b826e3772bbc72eda23732d948de8cff05fab007b361b2b2d5b54d763563837db39a27cfc2a72
z7da1b187afc72a56308892508ecaa9e1eb788adc1d89c900d041bb10629d5815782e3ecb97ae38
z59b73643e3e61a76d04b000900c573a13b019cfc3f5ecb2f3a21b6658bc4cf74f81e715c21b599
zddb7790605990a082e55ab6b19e77c94bfaf4c53617f027899ea018a9bd2a02f0da64d26aee32f
z7aae4d8b97a281bd8c3c57b9feb1a1ed890c3001448c2053590497a7c442c067ecd877b247981a
zad2f9d897e55f8040c52c13250ca3b574cb065c5fcbf50d23757507dd161d72f629ec153c0d298
ze2179b1e84b39523e4841598ce0f338d7f914d82c57df5c7beb949a276aa09ac2b64e165ec1345
z0d7c792302e01c0759dfc9f16adcd0b6a251694062dd474ebf2e939296cd9d92b3de12b4eba617
z8346cac376809ac9e4fca4174788c29f2b61e59d6f23e9804a13b4fafd6654d050d5adf9432036
zffd946041e21a7d63fe04fbf6c71bd6c231ab7e69710f5a65c6bcd6c02649210cde92cd9c20d8e
z72f520099fbc9f54a8828878a8fd509feabbf6edefa4e433b1cb11deea7676639d43084f8dd45e
zd84f009abeb6da05227c5aed0f4cd087ed4182ae7763489bd4321680a4a0ae291fc2b5fdb01636
zc707ac4c9948e7aa9aeafb956ff8035bd645f2599228f275c426acc832b89e4608f53aabcef54d
z43fc583ae598dce932aeb2ddfabd12b5d9433b8cdbc460de8191055a598ca038ae77c79f44607a
zd9b5da72740cfe976cb2fca7bf9a14035d358867c93efd9140fe13529f3f18412074f2203814fc
z9f17a7ddfa55655c7b412491d231c7ae32570081b9ca43982d61903f0d070b692c2ab6fe1300cf
za2d605eccb694b29d4e83bbded3bd8521fe11c1a404e67ad456e0839971af45b9105307e8686f3
zb226e1e5b433fdd52a8221e4917ab16b88f8644cd8202fbf0964d7177ffa358a4abdfd6d7a80ea
zc0cda34530a25866dfd6e644dd19cb7482bc578cf783e3884e21c271a68103e276cf62aad15512
zdd2e17bc763365713f660f1a285db7c7215b98ec474ac6c73b54416b528e2e976050a1fafceada
zaba5f20415ad9ff5798252eb3ca49a1708bc9f7dc133980b2b5b6a30128980dd6f1689a6c57731
zbabd3e09e3d7b1e986f0570814dd2a307dbdd171ce8531dd102877ade512fff2d2a6706d87b7f1
za151d94899fa8a0a767144ae8312a25856c82b9dc7c1964c32250c3615b90d01daa8fbdc66c37b
ze5d626f523ebcf982cac0baafe60a823d02043d04648d78d93e8e656e125b5536f80e3b52e6c74
z0cede1fd0d1a9a92673f0bd07698558a2401ba0c34c25ffbc759b7070a0cb74ea996975d74b596
z2ee40512cb051404e0f02c22bc6050e12e978673b5207d2cd424f80ee5a0c4d5c1be8f1e4ec189
z4b03d5cf4a29eaea3325cc67c638c94196a409ebf92a36a2700c6dea60f7e4a017d28c7edce4a5
za59744a479a163ae449780fb373cd8199eaa4551da4097b9ee096516ddd618467d6430ae6f7799
z5bf5f2043ecc6937142b5cf8c00788444e132572917339b7d4b87620c7c2b549618bb8f2ab2d64
z90bd07474cfd09fba1a3e06d780cdb21a356e3063e622a05a43ba0c117c6fdacd0b91f82981719
z4437e93bfe342acafcea403ba3f9edc11045c0ccbc13fa2c1e9d78f766388e0b631d1a640c71f1
z7514c6e3a0e34daecc57b5c30329a09f3aa50c145114f0d1a85e4959141143205817caeda57b5b
z34694d66afcb9e0c666601b2a70debd55748a3cdb96bdc6bce0797e639aa795505b77980c590cc
zae38ecefa3b1955088e3942d3b6044fc30079a6009f5832deaedf94ccf22520a1aaadb2f1e2bc4
zf9cf09f5c2430805217354a1a889ffb2bca72ccc4ba2ff19dd2a06545c2201d2eb1fe47a8d3407
z2d0781d75d1d94757bce740a953675361d1bac15916133770eb5cc6864e5c75b79b8e7b7fed6d1
z73d41331dee33a5da7490428f9cac6563e5bd78e9c51f1a3bdd83542aa182e63ffdb23b87fd35e
z9459940f4057cc2dca1e07038f712a8c8d24d0d35900f7db82a1378e0fb3479b9efc0324250461
z87082dbfe96857de406b3e2a6491d7ee8ada077bf376cf424ff7deea84cc190841e2ce00af7f56
z115564160f88f64fb4f3a37a19c3f0e56a796ec96c041525a9133f45eb310faa05c77868843ac2
z54e6f2b2e4118bf50394c3665287a7e611ebf8c488a6d9754d5cd153c51d9daf16d054e9924f4e
z028ef83d7e404136683dda62cb3f2d99023903d01c5e8104dbff1c69112c6d1390a2f14ceb9f55
z3b21db69d6ee89bc1ba20265fe886c11aed6d78031dd8abb3c38c80723cbacd77dc85c10509f52
zafb4a9b8bd6a1c1b7efa6d39443e146b4748eb0ed70057d73095caf321be6af90b3db760d00a16
zd8b0279755f4d996b9c2d07fda48ba6d2d97dfc96cea278fc66e335e497b3e95b2885276dbc553
z619f953e6d74845a77813d02cb9f2ca6d1c73c6ad79fd59e0b7f7e0826382049661fce2181806e
zad52d91d08b7e539761ad527a37f6e4aa92f7f2a29856d4a769402bbe68b4de25ac7c4215ff44b
zb86e6e7d1649371f130d6475da7527b0b828f0838141404cbe15bc6b7cd39176bb2da4b08a342b
z2a9fb03d375ea016b29b493619e060563e8fa5d04dc670720eade4d784de3bf978398b8c4d696e
z94238237ad847fbb375cef38e1af6ab4997284df682792c323e261ac347ff26e059aa0400539ba
zb8ba8eb3a88d7d9adb51e4311509bcdef5b4caac7d4eb8e59f0547698da5c82482387ffcf63cd8
zd8f80bcbf4f16b4e5eeaaf27dc625b878f5526cd4a4a4ef77ccca134e05cfd9bf58b4321b9ff23
z4d1334567c3fbc2ec678130af8c864528829abb2273f5a62cde004aed9a70cc3be5d5cf1e4e524
zc125d4c4be9cd835af02666f29502148d8a0b2889bd71ec9479e9bbedf3f07aca751eec9a435de
z59d146af5ab980fa1a7ecc54e34fdbbb11aa99e44ac44d475ccbe41f01d24f2dda22c0f295c1b0
z82db2aa5b5212dd26862866ea3160d4525845a9e77416274f85d18a824c2cc680933b0b7bfb995
z6432b01530d5b0f90b09174afbc532f875ae20ce462b853c849f1dc4075b96d4df9c31e2b25365
z2a4b29a2a87c4e256f36647567678387afad1c8f1b5a6159957cfae38f0a52813f200a0c468799
ze72113a208fcd2f3d180636ce751d036e40753cf64f1fe5c32386a43b49f20273bd57c119fc1e2
za94f147969106a20922b011b3c3865fea9805cc136dbb94ab1242f9a20df2b083e065fd5b80f14
zc7dbccb71718d45db61b9578aaea46f51828ec6ba85ea0bd31cc30806cb656fd86db7cf1b8af4d
zd258325edf5faf0b316cac469290543c46ada1e78fc7600073940fb84a00d14b2182a459c0afd7
zdd16bcf3001ada71285a20d9b36b712ef5d347965221ed6c64625f8521cf6b257ec0660fa47b52
zf6f97de32eaf5c98ede9cb50ce12e3626e12a4ec44ff0bb348099e6ddb4579f217ab33a63d64fa
zc2fbd44635582b1c0143af96e1c337f525e874e4e797f903630325e972c69ab85d6b9c6e513ed9
z5b29f21f174cf86a14083809f6dd0abb83403ef84502f4e626816a7e9127b4f131850d907262f2
z620dae3bd752b2c5895651ab6572a82a8f72ed68de266de42caa922ea956bf984167936f644993
z95346c29ab2c50d47b14506dd943db47602768f97131f75b59da4063d1a7b21dfc8621a9c571c6
z1808696abf7a42ca34c25ea5ece8cf190faf0dc966748d4dcb60ee135b6200d2fae521a43640b6
z9866b1d5dd80d87d0ea61238b855e6809d773aa435317a70c18778abec80b99805dd20683f77f9
z5b5eebbca6d4af254af565ef2dbf56e2833851d0e25b5d71336b484d2c40d2b18e67d06fb50d36
z9bf4afa0e8690d6f7255a6f61c5314031834b90042c7a6a4168c4a709b109c1c155549b8921b2a
zd3f0bdbc49d2250a481152451c9a65600750349a96ce9c609752484ab5b5e700905f910a9553ff
z7d0723dadbc9d0fe276c8556b7215911626a01ff39424049cd32a54bc6ba115baeba4c35cc65d7
z7396990fcf03154a8b18d7fa50d765359d66c3116dfa084a9b571d2beeddc67b11b4f7f57da0ef
zb83e9f6294d13285ec3c96b7fea923ea294ddf097fb7bf820c542580852760d8697e10fc273905
zc3aa74a0c7cb185392070f84b69acbe1f35f116c624d35ebc3e84d0e453dec6330dde8c2bee79c
z2bc8117d66525b9494216120da29aae7916b1995ac48fe6a121bbc30b39eef44c214a15b41ed0a
zacb9f0de85286136638cd1ae44a602291f506de6635faeb39eb9b7d1ca577c3fd23a1bceb08011
z6fd962be06e71521a982809f7071c8d3c6a666178435ac58969c2de7e266149c5551f79f8866f8
zb0b7e2d8ba938ab7f4bf231eac03be151021e8f5048238e34abaff9a83d2d1248b4ca4e02c4bec
z23ce40b678bcb7de28faa2fc0d67d2aba5d4384344b21d66b897741fc87ce52fa2464f5fbf5dee
zeb7ebd89f66d8945500ec0f1aad50e865fb4699b6f8702c985e050fc4ef593448b301f60d2122e
zb8053db4148b0ca1170f12611032f7d83bd17023e19bec2d29f3da47a6d459a65e1bf1a6532818
zca267b572c6c143b5fcf82bc5c28d7c333e3806c3cf13fb8f1632166de954ebcc9692e17276f78
z5ba7ed15b7fbd76fcaaf36b13c0e48c908760ecaf106f5ebfbe8ac18c85fc35efcaeb62d0edfd0
z8d555dd79c16168fbb4fc71020a52c87d2649f9de71c62ee2d13590edc25b3ed4171ab50a7fb60
za42587be16acdfd91018ff4e79b556621169862bc567d875c22aa728420ae8bfba63aff3874480
zbeb8e8477c8cb2dba60b35db08b594fa8c2bef3beaef3fc757e676c3c9d6fadb238a9d840b1ccc
z7b2f208dcf30f77477e8ae0ff854909555c7b0ebb6e19cfa61ee31700cdbd3ceffc3988c51f126
z6ea895b38d6baf144c3ef07d780fde1a53c1966fc699d69ff99ab8b3b7505490a066931b9fce52
z3ad41180025b1e66d9b5da43c8555e0b1b8ebfc4a0a3d8cda596e9728971651d4abcd88197f298
z10a93c0b9994c87a1a9effc21b6a9a83f909f0f7fd9853c701bf6d2129681d4ece7a0b8473d98e
z44020d4d4b2bc73b3d7b1b72c24245e9a6458d4bae7ab7b3c64c449a48f4df8672e17b95f010a1
zc91e71fb60fad6157a21eaaf71f86b56ee2b75e7596f302a864908cd75fe5b020b829232c31ece
zc797b55e22d6e38a63000bca6e6faf123cca97fd10a0efafabc9c360f00d250bdef1d14039c103
z4c5b02bb61750ee0dc715144169fdf31a2588af763e8193e0170a34a3a5b9cf64816f5f33ead84
z47827bb422d14c7da038da817ee6aaccacb1f229658da8a5b7124c48dc3d13ac99c880255bff9c
z6e6fc46a7ecddb498ea2f92c3be3fee445d4fd4fec01734280f5d48676ddbf99dd66bc120b2861
z95ffcbc071c5c578dc79c3fb61af6c2079ea2636cfa267256978f8b4a0da709e797bd069383b8c
z7625f99bf375de1eb2966a82148b136783ba1d6fc5bed91d08fa59be6e8ab5aad17fe3e1a21ad9
z307e301cf6ab1e250fe13607252ea6457b7a146601b25868386b28ad477e37b825049cd6aa530c
zbdc525beaa3385d052e64ea1f13b15ec6d4fb40d80f2b1847f8c09ef16321c2ab4eeac3a888c2f
z7172c69f29d9646a798ed9cdf13e967239ae94b080ede569d8f1b1b79078313c98669bd51798cc
z6266029d7f5d73a68722f822b8f696fe8ed5e02fd841e30a514417fa170007da9249360863910d
zd0ddfff4b5d057a89a81ec778c7831c58f13511961f86426f5ef493f22e326e728073dad244cae
zcfb5907c891b8ffc69cbf0176403e7374b2d5dce4f72a4c08f9a9e5a5a5af0e7b00289d0850731
z329e3b045d44cf78087dee20adc73e9c1d6d5c0e47844005a5a99c743f6e74e378340da5fdbbd8
zc5ff945bd9b81ad353e0c0b169a98d4832e5c9236421d40ade2d2e850401d98966df4080229a21
z53efef3d34339614beccac0dd006b1367b9d562e3ff6e7168c7973fffaf6fb4b2902128d91677b
z6be36d371e33be6d0e3a1fce6b4d551953492a403649f4605dbeacbee5d43f5922c41ee597aa12
z827749ae00578345f1c77141f505c616d2d39ed28917efd55cbf16d5bafe8121c8c610cfdd832c
z447e81e75cc124e36de0ae3dc9d17b803c5e940d18cb84a354d2b527d437049b7be5ff825a04c2
z06a283a88177a6b5f076daa181df9401cce532f126398035b635e715396faab19a886142713563
z69d21c6c683d35c641faf9f925fda1c54f7a5bb892af68df665cc1d209be60d5eded1e093f6ba3
z887d0cd01e6ef321a12e0ca659ed0216db581d8b7608781a5462d39b2b76f6cfa0cb3f3efcd55d
z5f22ed8239ce1d99e0d9d755dfcd99f1254ea3b3cc151daba69432f17c1f3d987c8cfc7a0605d5
z3ace6512f9567d297db2be5a65e1e2db9b7a3b9ff041c6d6d8ef830ab0ff3300dd8bdee8245adb
za221a95e838d918e5637519c30c8be902e8c6afe3776451b23623a4c85116d0dc788fbd4b9fb8d
z43f64aed07ce22510dff4888d9688cd40bc6f5ec8c3811296d49dae2a89afed211edc3d279059b
z9e66def95abda96a3ecee2a4d10ba2f982751ec20c47af73c0ec1ec13bbe1e55b844b2d062e8d7
zc973f001fe0adad0270e1dbd5162497e264ba5b1098e8fc0f34de632e7b194eb99cb2fb5ec7d9c
zb318d8e839af023fc2516111015ced41ce8b7317c4337d23f50d1301ca46b79bb9b6643ea66d8f
zf6c5db9a153aa5f4ac729bd18b5f933f218ae754bc9addd2a2c69821528e748ad5baeac8082734
z362231f87bff218ba1f42a1831dd743dfa91ec9c95d7cd1e31e47582611d97f6eb7d6fd0d303a0
z04c0797e7775bf78c5220a83ba5f37b9f4d890951cff7b7350f508da00ed03ff67e4618b921185
z0ba5e843c3260b4e188e0945b355882e0ce7176959772160bfdc33e45472ade006d8fb1686974e
z51d27abe134f52eead4b4bca9ce5e7d75505b02f6c65c7cf7fdf9967297221667711d59a1adebe
zfed8e36999afc7a62569acc92dd7c3c357a7439322d205846a3bbc89e1ed7682d42c777f25e8ac
z66980297f51595bd5f21922289c5a9f1314e76704d479a90ca35b18aee764e96b8d49a853cdec0
z70d64e00969a4af6b9648efc0bbe463b4d8b2b0bdd150b9727a891134b6ac4f07e3404d5582136
zf84ed3425e3655991ab160817ffd1b1fc911c53cfd5a58efc9aa389faac9af2596522bd558be53
z01a278b3cc5cc28c15173f92a5d56581e213d75ef53386b415563b3015456003d864274f56a8f8
zfc685ae4847f191795a62d989a92a251914b0e5ec084e93908216dc117405b6ca39a9c3b6086f2
z5f387d00198309df60b3283dbb9cb4932940578041f2953467382e82b167435afe7ccec90fa4c4
z1d50377b4bd7bbb3306e553c16334a065613028a7bff393ba6813936c27af9b32f99c80896eb25
z5a7ce9a62fb814bb437b9473614a16ef329d2b0178ec2053a6bb92d7617b2c45b0680e0d9bedce
ze8768e066b4994e316af87c13e8cbddacb2560b3d14dea7c368cd298e231c31e939b537611bcfa
za721b4f22754ee053701813fd9721dcc1b03d6dc8ee0b5a8e8a66dea951c9e5dbc05e802503338
ze861a1b7de66fc5599bb2d25074923fbe5ccd4a5d639074604c0b89d2884dd6e65f0c541325418
zc976184646c95dc86c9ea646d835b7b3ff601307ad51ce113d09efbf3c611a6dc8e77878b0c582
zca3e1bb7ce45dcaad049ad6a19796e4269d46ef71b89a6d73f70a62e0dd87a1607f7192076f8e9
zd0b856dbe2e3a2b96a500facd06972bcb16d2aac8e2114cdbac6e3583311000615a2813413ffcd
zc4a2365dda061a024832afdc8a546cbd32eff470ff164f36d2be05bde3787fe6938f8e4266b31c
zfd224b681c4df25ed1895789a680d4388f9d5545c5ae91c54de1095a6493499d542d3b05338feb
z9657efcdd4953614c5fde421cc708c5c483344cc7c549d1c680ae42a43911826b49bd0f18a0884
z7589697a3e9cbc294f1de2059ac2d3b4e448f8071f7a9135882326fd456f72f0ce98e47febd631
z60d9b42556eda4951b7d9b5917a734ece7a4a5d4ec1cbec9a59993623313dc31836d55138335a2
zf7b6faa3ca12c468da7fd240ada1baed5bc9201acad428a6ace107d28b0b39a7b85cc2f2d9efea
zebaf946f3a73ffd0ba62f61c1ca3a9bab51c84aff95b60de6332e389905799273f28fd3d2fe1c7
z6132d049fcd93123e9faecccbaec6482821a86e90a8112cec9f2f825221523792f935ec7c33e3d
zc3e597493b31f06ceb0aff7ccbd66359b880b9f5637814c1a4c3b005cf14365f85ef81d0d73599
z175b4db6068051403c380a0e654f5b54c426a4427d2e899fb799e15fcdf3f64023b1cdcc9d404d
z313e7d10998a6e198325ba1fef1e0eb55d7f2aef8324952e1e57f4eec1ed5af28535e68fd074e0
z716f8777e97f2fd5c8f92e86ca8a99fa8acbfbfd590fa43efeedf3cf007397d8c5006ad0f53329
zdfd707ae3a8c7e3faf207fe867da689985df826a771a2303b1594b8daa68f3afa827d2bab2531e
ze7c045255b4d89a8a0cf1bbbe493dc09a35b7c167c6109fd92285859af2a38506a873825f0363d
z9381f507bf709c9e676ff00bb4ea5da1243fc782ccb3566d90aac8979b741f6314071cdf5bba25
ze074b4c32b2a69d4af4dca952a11b405f6335d227b3ea0b9edda7a3a5d85248440c55b1b2f1f05
z8ad4e4e3e1c77cb13f32c0eaa4cfbe84682d55b364d72097d6f5530bbbae776bb45f019449e66c
zf4448079f5a6c8f17a39c3859d9613a389eb10390c92418b4f211d8ecb121e078e8787db3b6195
z1a80b3342f040097e3acd09dfe9533ad4bd3586ac21b881c6892cd4d0c432f5b671291f2b72c47
za3be727584374df4f2401b6b7b29f014ae6e362f0aa1149fec89595c015d24d9a4272da25b433b
z66b9ef2cc755005bfc1f506b7225e3cb82803ff72196012a229634be806b55e01256e60a3f6828
zd767050b1e1a046a5a255dc104aab786286483d7ba3fd2aa454ba245f0d3097f80a91e9b33327d
z2514a9424f2d67cc41800fbe332f735754592ccc10419e3a9b7705da181fd0711509263460c994
zf87e7829e2a4168a31666d8b1845355bbee71421304376e2fef2b4e49b5e967aa40b165386c0e2
z06b08f0d0ef1b31ce5e94dc17b51ec9bf234580f2707ea0e8411d0dba3fcd3986fa286d9214085
z66da21e85e4f2dbcf136332cb0a68e4f6c8c066c94b2947f3a0ae6dd44f8eb5479044912237c79
z599fc6b1918fed104b30f569e346b3b057238b12dc516b95c36d31dc239062a7c390f8552f4301
zd86cd5722f20f0be25d530133f4abd8de9a36d3a69885710410e2df992e816ffef8f13491a2847
zd6d6a2db1ec5435cc188f2d4ce3fdc534ec41051ff74a83089aa90a14ad61a97aeb7ce2ca08ac9
z48cda0cd2bac11ce35f0939af4caa299e1d2d8d453d9c774a5cdb6d567f58fa3481c49da9f1517
zaab4a966fc37ada25296dc20028c589e6a77f6c9108a31848351644744991720254bee19e7ee15
ze1a96400b1c4fc875e157ec7603c1ead8b1fc62b91249dd068fde4d8a44f5774f177c0e350c7b4
z1fc6872f063093dd3b21d4af6ba1a009e5079773d836d9adbecaa4675b0a4026888f5dcb1b87cb
z2e09e1f4ac8dc0c707ea2e2407f7b23394f827c473655ada1297f79a0d863212c31e3fbbaf3b66
zb031a58cd75a2084ddedec12cb02cf2686d251ed806d99e3b7f026bf614eda5b5bb3c5f1e6585c
z557afdecedfa018f6ab93a0975c55a7d74b5b7ded2ceac69c001561528e1ecfcbe05ccf7d89f5f
zf7bcf49feddcc3deb17d8705d71c75b92e1a18f862c2e1ce523446bc5052da21ee1aa20c9bd973
zb6d4cdf6fda01988b612cab410cffb34a8dddd183bde400b14d5febe67938e5cee81db0af0871e
z9e9ca07df658023a4c5b4b6922a9e724bb139ede7a56bfb3b265ee84a2c401178d11872af424cb
z27fe73516b8e919e3a1b15c8132467e832774b0f054f20bf3636dc6c81758e3bdf0dbdea1e1dee
zd8b538bc3aa3bffc6513ccc3212040dc8905556e067ae2240fa6eb364428563a584a0c0769e830
zbee8f48e5e3fb37f3d0a14273a9832dc0fde4023e69b419f2b3ed8158252663cdba516a4c93113
z4ad3ed35d74da5e37d8ebb71216b87b9f29671ecf6f99f91a595d351c01eed5a098213adccc946
z10970007bb32b7fcb561b9d52821d7d1cf85fe441fa770ed30a3f16f87ebac1366c726619378d6
zf992880a484bb736fc11fe0baf99da5404b84e67d7759a6d39ccddee4a643d5fa96fd4db8d3da4
zad275ee5ff4cda32db7119d44a2d71e53c176ffde70a4101142fa48639d0465e74d3ca6c68b34a
z2e5112652526a0ffacaecbeb3b0226a2f8bcd4e892fa9bd363e4067c7a15d740cfd2287a202112
z979eb6cee12ad7de47c157d6fba80763028c9b92d0138ce9f8ed238da1e08c72b9400e22898c07
z9a06fd322ac83476cf0a9ee285c4e221df77b37f5e1864437067d883d55bd2c46c415911435ada
zf42ae82d33a892e004d0febb125e3415b4e48701940e12f3a086714518c4fd298fcdaefa6615f3
z13820461a8ca68eb6544634751119f0fce45539af56772125871341f387111c2cbbe3bfd2f3a28
ze782d55a92c8fa465c5902636f129991c9a9072f72bd56b4aafe96cae89db59d57c1fbdfc21321
zfa6a9e9537a7465d1ead78d34c8535a8075454607e21a11be91cdfa15f7c57d1b7d7073d9b819b
zbe24b2f2168ccdd8a809f89eea3a745e4a8b6e90a3c7b013826b0eb46a737d4dd62396136fc34b
zfa9d254877e8bb2c9bdccc41b781da18348235fb9f768c79cf8580caa81f91e07ab59f57f8d5e4
zc39dc831a45c4eab6a57273c8647c04e53c6bd54f24d33a2d09efb885b23dd77ce6a1d10267139
zf56f9b03041e103f3938f83c192cfc5073da581562e9126f351a284804944b8bb710cd3233ca83
zddc3326dea8721f280a2e2f023760ed9a54b34300035a6f2b3c7d8b2e6753423290ceb78d89712
z910245500259f6ab79a903544e7d76c9601127d3c8522ba943d71d0430c8303b4a04dfbe1d11ac
z25d3eb517f0d785aa5c8c0753b918495f8c7917602fe1d2e12e19236ea069b625f8183c976ac2e
zdf8bdc5d50baadf7793aa42c3bf9c9c0a871007e9edd8458b68e6cc66083f3dae0dbf57da626e4
zc2b715163cd9c16b1be72ac3cba66bf5fce2068bcdfa2f6a8d769d87c4e0c66286d4eb1a18eeed
z3afe7757f11161d8434f9177cf8309a75c751d19b88097f24e1dc7bc6d301a8dffe4ea213f1c1a
zbf5d511f53f6bd2b2ff606fb2a143d7f6e998dcd119a8d64d04853fba277982cb9b49a53513eed
zfda2d1ea44e7a43f6f8dacae66df08ef2bf0b69d06d674ab7b9d117db2638520a72ec7f42d647b
z7941a9f70414ac99e4fa5254811ad9a55167b961574e3c126866142dd6f872742d70fdd8e4c490
zc57e9543ea3b7b4fd0b903d02d94944275cc3e28bc2e527f47d5d37bfe9dafc632a5710aee1fff
zbf54de91bbb4bae41862308047309f748ca2ba3f66b057d1b6c00102ca2dbc55a38ff754aa124c
z036f11ff6e965c5ce8bedc99179e140d62f8a1522ba0b0d0777509f51750f8c3ffc253695250f5
z3fd49ea26174e5000b8940ba0b0732e6b28e5a0dcad1b1b04845e8320d241e99777146bf47fbe4
z6dd331a09642c35f24ee776ea43a5d1e2e5373e2ce2bb113d8103b0729898a0e7d90549385bb89
z9b286ea151fcdb1adec0b25e7b6c5eeda8cf822137fc61f12fbc5dee556cf93ab3fcac76e132f8
z669cedc047cb667d6a1af39d934cb3c080aeb052aa447b9d056442506fdb9d90fc8f654170bf26
z66fdeeb9ff8140ec89e6c9e89d364cc2e9a0f03a6083f23593de77b26d734666d0d5bd2a8d6ca0
z6b48ad2eea2e9b4ac60827a7d4875b41d82a0dbfc3b098a56c9df3831bd703f710d2aac699b67e
z474b7a016cf63a278f6992ad49ef773c96a29487d9581823f25d91cee780f1e03936f294d88788
z66d779b7475abb2b2ce4e130df2ecaec6b40dc06f83068086673aa3930098aeb078386a1190219
zcf0859a7b81ca38396064933add8d1946faa2962ab26c24eb74a7fc5aaac30a58169700198ac79
z9acdd8d5c1e752556fa2b189a30222ff9d08b977790d0e4e9a30378061eaba0a51bef86cbaae09
z604ee8f6119daf00acbbbff8c77ba443ab912f514d3760140fb701c4f4ebfb6aa0596ac06b4eca
z40f2ebd55be360f8baf604ba9c4daef5aef1b6bc674c348cf5302207f250ede9c8cd41a171939a
zc664ec171977aefdb2ebf4acdd27469404f3db5c43b54861695648450b6e4707b149c3a3f4822f
zb988e2d790493396271b45460df81169fc04a93479886bfdc17617a1c788e30bc803abad4f98ac
z7584e96ba16fd84d9e997da5b294f0c69dbc9f1ab9900d9364043a491cd7ff1e5eef15c4bc7f6e
zc6abf2c203a2db32851795bc6612c8f54d4ad7a1f74a08258ec898f30fce2b3f2c0ce3057ce181
za47a93698a46693195f318e8b3a930817d6855a5f5b0555fedf32c2e4f0fd945672ae38d214930
zc268bb595d5e95dd0f7624bb62c71223cbc8e7b7f7fb4d23414f8757319e281f61c39be12f36d1
zb597ed98205f6c3cfa0e27f9b5835087817b2ce3197bdd40fec5fe1546223070d488146013d380
z446702a946f007707c9709fe6f60994bbd62e4e0273b24aafcebc26a5cb380cec117408af41211
z79d2ddce9fbd4e5500829429a35971f3e1e214d81c9be100feada1fa6ad72c9ca45f4200cb57ee
zbae62e52a96cd2e0376359f0b6123cab5295b2e233eda3f84e91da82c949192ce712a36286a082
ze077a217d950e078aad3486b4f31df0cfaa88a3aad47c497805637048fbdb62bb156cbb9305efd
z700765d2c69ce947920269edeb519f5a81a1e17464f622ddfa437517d8767356fdfd441fc68ce8
zc0d21fb73051fc1fcb6d91e35a4389a119a458257189b53c4a745bbb67ab3d38a1b1fb537cfd2a
z3f72b667748b4d4d065aff33a7c183b70ecb86aa55821f7d29c29294f1699f1959bbb19c8170dd
z20f2c1cc4d1d441796749ddb0289065cc828e3631e44ac9145dcb052a44da5c53b4b02608b3b1b
z98bccd64f2e22539e1460d90fdfb021920b8385562f80dd6dbf84df076efa26a7bcd2cf3e05056
z64625bf9ec101eeffe8363eb14701daf1d8a0c249646fbb40059b07748d3d3d051cdbc1424b4ce
ze4930c9e3db8b31d9bac031cedd708ccdccabb5d205caf7f2387e17ee935c8d00e3fa7ca35c160
z1ddd616c5e9fad2d499ca7e965fe1d3f7a654c8f23ce6befed950001e985fac61c9c8429bbb6a0
z79e1c8ec3503d48423054d35b48b51851d3f187a69dec6695503042c044a616565186d1498351c
z46fc6221cc607937530d896ba9cbac682e8df7dfcabf833d040955f4cebcc56b0f848eb2f7d9d5
z87a40530dd27c82fca1f73ac8fd826d6a25580355e4dc4b30db9070b17f26591294939a8911581
z302e83ec51d7d4fed28ce77db5a2560b60ea5e345a14ecb549e3b2075b09d33096af42cb9fc710
z99f56045029c080c470ee464946a1145df043941c4d19228c700477003834e2fc58eb1ed443ecb
z220df657bb8e71422be51f04692004c89bfd48433d5e074c8ba35db81601b327b31891305d5e2d
z5be08eb9a6b409fd3188a3eee46569ecb39631978fb30815b1cc8be3c8e847e3e49518a784863a
zcb712c7f9a051b637184b9a699471ccdfe884ad9989d66de8146f08423a8bf397368cc6df58f7a
z89b7f7760ed11422fabf105910516dc832788b26d891792d60de33fb90286c4d63ddff537644e1
zf4c5866c7e930de6fbeaf55c21a937b531335942c023c6364b5a8713c2919c4d31638d5978ea21
zb1fcb38ba6540200d9a5df646bdc40ee4358d17dba0084758aa666d3c7aef55d03b68340cc12e4
zf3fc2c67bce79c7f69092701818085964cd66a97d0ee2d2679acba9763ffe82e9174be38f88f9f
z90632f02509a3a8d520c1ab967757333c351c846687a549eec09c8738267571951be6721f6ef4a
z011acd37ca995f1bfb3c2d0f2a0956f6dac432e478964407c3ff7a68cd37d2f1bb6d630b920f59
z08d3fafa725a7711d4c9baaef9c4b2c58fbfb6e523a0790df1609176aee5e95151de5a77517505
z046557af129241357a26033ca78b4083c17f80f1fc4db12126fbc255f7ee4725f0e5bb0480b141
ze4084910c30ad7b19e54f53f8b9e3f873bb8401b23443c0618c1a13ab4fcadd079fbe5592423e4
z779d5372cd7fcada87d56cae9f6fd7bebc985a4830ad3f97f448bb96c17c6353289a72c8b89092
zf16c3a59a3f8249e5ecb0982f041c4683e89d23d34002d369bb817171aa88b3ece34563df95dff
z2ba8290c7bc8fc7212a75775b67e44b41eb464f4067cf83826a22bc305d8ee55c83988ade5cafa
zd1b195a769be6c7241ff0958f169b4927c69f8b6e5bbd08d04c4a7c943168e2e2e7caed3d800fb
z9cdba455f6d3f13b72972d3b34965285a1691dafaa56cc308d4e465173f0aeb5b8a568d7ce3632
z0a7ebbd0fb92cb8ddaf3421462f4e668f780f481b14e09cfe15e8590ccdbcf7bdf7e06491b6169
ze4d8467e003c2d4d67bb6686a09ec57e16438cff2d867363f34aa1a45a9ff24340631d4d135ce2
z6954cf8f542c7b47f8c6e91ebdda041eada3734d9150cb91289af64d592a18b6327fd366a83b30
z7d7b7e6fdac99e794d24b14e907ef18833c015dac1216434de2eca55d01888d3037cc6c5a920bb
z618294e70332eaf6ec13f2c32e10d46582d14a43374a144dabb2b92e527b2ef79e50f6d57de7a3
z87d2d6d5dcc31e03d0c6c409be1fc8bd0cdc924a008f45f5f8de78192a9829e946ba193ee87248
ze96803fe54c70e49b6a6f248fd541329a8b102269e29287b68056f2ddbef3ffcddd54b601a5b33
zfc41dbd02ad8a6e1006cdb72629c9947fd3a47d8ad1dca4ad996894dc4a8a90d6452832a6fc931
z407a97b58b9471b3e7c10cbb85b967ee93e1f5d40540eac2da1aa4fd67fefe7eae62106dc3559e
z3a26a40d2454aa283720c03c16a45fd1cd9f15f68eefe644d5e9bf99e5e9449ad3efa5f06cd962
z9d76ef438a7f148a754163e90d2b63fc3ca3cdb3444cfc83927c1464690f919cafa44336919243
ze92b75ef6e91554b4ae439899e202452469ddb5972e1f8695f22c8b441155a8041603a4a4515f8
z117a1f03f79fd0fe4bf75f4083ff978f69da1796f9756de5b7b1d9f6fa45f44a21ba62f51ecc70
z87fb97c3e6f667a14a732960dcf3bb340d5aaf0860c23a00e94bc72a4f18622e23e84568e71aa5
z77fa418d9544a90b5b40dcd2eec049be73bf8e1e04aeb94fd6d5a4b65cf5857ecc362a7d5c23ec
z0a4f4c981564049150f5681561c8c8ffb9b00028a3b0a60cab0cbb422a8cc43a8762eccc001d34
z24ea667f9b888701629318c1308943435977ffc0d1916cc5b7fde0197557c6554110b12ffe62e7
zb9854828af14012471a05625abc379f51c030c42f9dd0e144ebed6017fa4dd2e80974e618be6b7
z3299fef4d6f8aed471f6c9db5b472c567073ddf903d95488e0ef57712bc25fc07cf10d9a79397d
z2f0f5b7e4905a5aa63b768f2ee4534709cf5f7cb111c10952d54f9e372ae206453f399455a60f2
z8c5627e70bf54b9f392ebacbc38d83038f73cdc0873a194f5379a1857e89b630f728f2e3e69dac
zc4db7e940ab28c85be9a026efbab454ab5ce8db82c9a02880765f9cb6a9c533299716f5f1448e2
zade1447690448e1c2be3dc5b1d1db617fcb1f17a95d97dfcf31c7391a466cb096119ad4ca32208
z40fbebeed0da1b88f362b6227c8b7dde1750276dd991a67df6140545a5dada1078c69ec3d9b362
z707949dab8e706cb45a1a7e27bea6bab166c20ca7e7faf45fcbb0195e4cc5d99504b1cd6485653
zc04bc6c89d2abb648539c8d49305bb1fcca3ad92260533f0b1f0fb435bcd15cd296eaf88b8a940
z912814968bbdc5b0a2bc348149b96d149c1b76a06762cee5443afc7e7bbffada2a335a69406dbe
z76b49d6419391a8cbfca86e96494f63d04e50f97c0947c938a517e0be87fa9234dc3e25ccd6578
z8091921bbdc8c32f8ff4cdad05875bd60e945aaaa545987b8ec1c30195931e0b6c0d7eaf7a76fd
z5ae43176782505e292af88bae77f749c6e16f41ecb1b99e174bf6d0c2dc1258ade2cad868a4f11
z837e0ddc13ce01bb0de626500eeec45ea8e390c55e9c69bd4389fe165f29aeac9285862ef30bd1
z2edc00ffc20d399a438e549986dbf4d4ae7e8c79eefe87a0f98e5994b8450ac04156ff01d21704
z4b067c0a62bbf285f60d65e0156add3829e928428902b305361b9b3fb8e893e98303e018852fd5
z3ce29e45e969a61f8a76dadf5036bb1c1a74aee08b688b53c8b1cdb03193422262a0691604a198
z825bb947a5bc5ffec99b0401d00bd46fdd00bba4eef217f5b66ce25ebad4c99d8d5c3413186573
z239645abf068ac4e1907277cc5fb8b6454b4a1da49e638ea931110f1c3c687733c5ab7db7849bf
z98864dda8351e605af791fcb8423e8915d6e19ffb414a36462b3e46aa7ce7044c5093999193a48
z9d314bdc6cd550b7b8a20583299bbaf553ae6f456a0e6fc0064c743b832f3cf1a2dddbb34551ee
z80870f39bea4426b949e9cecd56b2c8d48c3afdfbc8024e1015c01becdb2216391aa1ef67ddf3a
z80885bd3fbfcb4279985fa573113714de8694430b2cbd2d5fb4e444a1708f9eac7de1d35b7f974
z70c36b09038e1828ea6949f8b765ccaf168aa62b15b8a0cb58cd008b27ba1b6cd58fe405a7a7da
z5b6c7f9835deb400c9875694adcb72de2cab8d28a7b1806f3cc58b27a884662a7337ecc26de3a6
z75aa32fb4d496825144f2058c6c62995574f4662834754aaa4ff11782f4c64ee716ca6e319a6ca
z22f6432656b3c088a9ceaa12ffef7dc73e734a7a457f8c741dae5560b3737ac386d02afbfc8a65
z8a81d052d6436ef7d4941485465b02db1f37ac36b43d983a6748cf4211be77b7d56e8020a16a0d
z57a622bc7e54afe47937918d1b2802dfec7a58a1b72331d15705722458ef1629f535bf567fe8ad
z8458d4dea7b26113f0214556a21f88d7f051b9f71ebbabdf37fee065c1c3562cba5b666281ecd0
z51379d23c5d34c7a64320f95a88536f678250d585cbd0716c298f258e70eb482c4e9b5591abd93
z2659024c0abcaf8e2ef3dc0696e93403a5957ae510c7ba889bb4c9c01ccecf5ff079346b5a970a
z39a575743a921e87c4be489a2f08dde96853729c0fa8b18a2bc28080fc7eca018c1413800b0c5f
z9f22f024af3d69d20e393e2e9fd9162e5f9d136ec1e84e1aedb4e716e9b971d87b7ab1088c1b11
zb4903304cd04aaedf1422647684a7a49b8e0f9ccfcafd3b4b58194575454e8da803ed2d1caf2a8
z91c5a77f0b61dd0206402b652f75e15427f0aa4a58d507fe4c188d4990ac226a6a4ac65f640ac4
za27d5aa2a278ccd3be494336bf1d6320caf31f821de1c74c0247f649c56844f232266ce8e915af
z0dc7a0633b5c2cc4c7aba47692bdcfaae8d4018dc49b2d1610e47b71ae3a5439c319abc96592b6
z1962501f45a364ebb6a52d2f3493abf1ae2a9652586653349446195ec6fe0d2ff94c4ec9eabe9f
z710f457473f9b0797709540f680a17b336eff079135f3161cc10a923a7130ba202c2b376d7b483
zb1d83eb2df6b8cd4bbe1a978969823d05729f916b5d6ee2fd6f3862c980fe67dfc01cef61e584e
z5b14ee806d8d2c6add42327f12bbc86f73099edd85c157bbef83c74b59ad94b8f76a78f3057ba0
z7fe125dbbd75ea485c212f7c665ec54a9ab32854b8f2f87d361855fcf265cbf9f25f6aafd3685e
z594b3b3f985c802805f1072477f81a2df476f18ef1a728a3225b09fe880ca78615a83215a1c5b5
z5ec106e33838388bcff6530fecf37de7b73f8090845567d91a815ca63952e77399f1e2afe38330
z8c0a5c11b944e94b22c469da40cc8a4496b4265557823b25a049dde6fc33e0b6e1c4fa6bb95051
z3d67ffbf6da16b18549b480e17aa542a9116c4c5ec7127b054b9c5094a083d2119222c1d0596e8
zb5d2a843390315294d1395a30e3d7873089cd61986717f9c71726c8f7ae46b1bd4b2c40830e8d1
z083df3fcef252d50cdf954c495549c5444bb765f0d4fa0442a5cc1e63b081d203bcc71f55db45e
z04c56c2c33eaaa32daf5ace1302d41ec13c326463213215d9fbcf89857129fe4dac9185b869f4c
za1a6b8d25d5ec8c03b2ba85ad0d2849c8e0b1a7de23d1e02bb1ab0243ec124cff0c1c6284da55b
z7908f2192cd20881f154841a189d7db746a62072fcf0be0005181379258d227ca2754663420d72
zd92e45f3bde0e144ec6bb375f2a8eadb46b2dfe832a58f8bf8f6771abdadef4253fa29bb685537
z705ec38c72e7c11cd84be24053db82bf434398bab9e14f9df589b5a737bba19eca79af36d831ac
z0df43414675c9bb38dd3db4718c8235192f4ac643c9acbd079396c5e8bc7b12f1a73ef0815ff5b
z143c6125db434394456bb6f25d64e253103884d8d2d511e6d8ce4600eaa049928fd1ed1b45b257
z40585221a893b8648e68568b3f285f2a350eb0d97c8718c6c16dff521d969442040c0de181da3e
zabed18bedd361225edef5f6fc74381e87c5c7880d8e0e193adc07b4e33d0e586e8219da87f9af2
z942b3e8d2f3b2c7c4b52025180fddaeb7b776a4ec3526652c5414a32ced8c219c884be98c274aa
zf9cc5fe242a27e291d49445bccfff2a4a7abac94e6b2b691f31bf66b10fdc75a60672450452d76
zbda46ce785ad9d99fb74ae7893fe3f4554e4f61bef3e0c3b60234951bfc2375342775a12034dd7
z21f895fb8a7af21d75f64faeaa4e9a7064a3c733885fab75786c76a75ce7b059288111febf8199
z5b58ac14c18ab041ec87132103b3d1f5ae16fbaa22bfab68e784ddfe3ccc87037e43bbe5dcefbf
z2e7430ec399ec4b94a437f21cc1b1e6d1138d620fd7418abf6c37eb584bd626d20b74b3231f484
z76774c125cde8a209cdb64f4035557d0369799b60298661d710eb5d277472f7d6b1ddeca27cbb3
z8ed48d0cd682dd2e4ad7faa1639baece012c3ca4f85c3f61026ad51d1b19f4b42e0b086b1d0757
z58c38011ef79a9ac432585cd063909d134583ae3233c4a648e585f6668f0cdb019da3c0952fb34
z5e3bd666486c7d7b570d04b2197d036d122af31a562cd318a1f2d46a73c1f3e75df2c34b0b1c39
zaf5d47358142cf3a0e7b0fe12641776902a9d03c5c953b4894aed927086d1515f516ffd08f61c2
ze600df692593f9d99d455e1f197b3c77f267f55caf2b77252d88a1540619f0c5e37765c7e78022
z6c99859921266c74fcf35c91f490022b0b19ea54daee07e97b8f23477480eb211cbfab7c111ec8
zece6e5dc01a1c585e0404b8b4423115af740de172d60b1830fbec868509e1eb8e00b0526713a58
z7f971ce410c928e8c9df145e0b67245a309fd6b21ddeb16f0c3a102596bbfd78937e6141e824bc
zcfbf153f38dd369ea83a81965690cbca9e3a336f0260750a9a19c07247e7f0f67224042aac5c69
z8779c1abbfa60889ea869f7524dfc1e6725bceff13bd44069e896885f50e8f38ca1950cc8ef1fd
ze89d6d4c14feb33e4e82d5861bf6c17ecd6ea710c3126080e9eac45cd869b2050ea4f343ca1a79
zc2db1b2a45e31702d48684db5dba0b1b1fca5a7661da5f57222f9a8a7899e8b276fc3b53c9a52d
zb08f6f5f73d09b7cd2ef4937899eab09480806e5fd04258790856b578dda4c0b4bbe3a5f8e38f0
z9fee4b48691da473cb5c73163a827991418f2e797a98ab99aff82908fb4fadb8c1876419a1752e
z8138c0c11e1596d841122b37a779a7828132d9d2c233a29d248701fe8f256d6843713977b887f7
ze3f1e08eee18c6bee22a629f5d03ae4768065f26298e0ee5bc179f25ae9fdc6a2f6841a5a94590
zd99962287f54a34cf4c0d4e28a51b201133b4c5bfb0cbf3ae56e72bad13f3ac24b24cb18d0f381
ze5095352f3ed812aafde497e78c8606288eeb7d112ab69bc11239be28e8b88f67ae380ac1e9ea8
z742afa8b229a470bc8bdef5be9b8c33c0420724535db98615968f0a7d0be02b34a0aeb3e79b9fa
zc0033f635e8a8ef53ccc2de7f9bec7dc6c2ee6222f824c6bf15ebdf5c6ff8acaa7f7b15d3418ca
z89730ea32e5f004c5c3cc00705d11490277b10716c052d70a6dbd9a25c246bc0a39443f62d72ed
z63f9111e72d8fe10c4452e2d8a17382f6feefb38de28e0359e1324de44bf11d67081158987a5a5
z04bcbf88715eb2b5d00331293426a5688b79c561d5bd94b038272a3166366dabe47fd9e21ff3a1
zb95aa764b35b510c01b1da40bfe23a25e0fb0b3f8c7d442a9415d36642695510f518aef8c3d774
z649edec4258111c8a3a22a826047e818ba4e2ff617428f6f41d7cca8f8354fb812d7547752f9fa
z45b0f7c8a2523d51582b44671a809714465e021eb64ce7c41eb46b784218498ed12377b2e9cf79
zd9d78d218a2aad31e1e6470f1ffb5379afb464c4ef3358294e53a2d25a1b2e5195bdfd64e4be69
z8b823bb608a785be0e6fd3d7de07509630eb0350ef756fd3f7ad7240c2ec3644e9775ac0f58b32
z1ada6794d67f6bd38d35b41b3017bc8cf936ed9d8bd1c19cceaed789e9f8598cc13a5442a767cd
z91ca93187a2587c8e1833c486b81dce7d44098f00f716ae758d89c5c2265b3aa79e65fb70ec59e
z1bbcc7f66572bcc36febf7827b1c6c94b7de4dc0eb0c001ea79b011735dd41801ded7cf3a84c48
zfde6686aa945bd0e0ab5e57eadb02f5262f75cc972e809493e38dea464151df6c2eba1ec5847ad
z6edebfcc323ff2d11d4485fe63d69e7decf2a8bc52c00cb0a0c96a92083daee1df5b253569f858
zd6c06234968e9c9bba09e33ec1ad3ff555126456b027f47cb05e76e7edc89b8f8f5bbae7bdbc82
zbb2ad55d98eafebf1a830f72bccee759d6631a02b67b6a93e1b5f69e02037af12867d8ba725f81
zbd8ef4ae2c4ea943f98ae0146f4b15c499be61989808ba045923dcd77a1f8bf68d4318b3f39627
z45ab15847235f71df01c9c209b0cb06f2603ee6b8a7b831773211c02f1bad91043914bd05795d9
ze80404ade2c5a3665b4c4e5f207a48d90086ec91fc399c470f09bcb274d19e8ebdd1525da63a97
z16b91bb303d4092293aa69ce6233854b06c2251201b241539dd809b34a1a858954402fbb01b8a7
zb13651bd94f74990381d8e508be025d2e85c5d6fd6833d71429466515367608025ca8713e754ee
zd3555a7a4b4dbbfb45dcfa6cbb004d86eaecf0dbef0bb0326679f590692302ba28481f7b434edb
z05bfc64c9c8be3867e5337e5c0357be8914b2eb34c1223ed25b6718b5c57dad5b519624fcc2e11
zb9d51dfacf7f0d58032164e7abd6675d00974eb48536af11c3e69c0d5cebb84bbe5c2f39081979
za3cbcca02cb422b165a68dee28033e4853e800e5388a20dde14ec82ddb53c0e1c448e08a84b0b6
z1fbc50d7b9837194a19ff25013e7ece5b1146015a268159bb61f9fdb047c3d1e9c2540b436a674
zbf98baa5f7fc1726e3ef43c2eda80e8279659f1d4c29e7d8ec8611006f071ad5b49122a46fbbd8
z34ea8aee6238287e7a3560a266911a763d44974968f28e8e5e75b71446c562d5ca26013cb50793
z14959c32c3904f304b244d4e6fa0a2e2092c63cad8dde07b07133ac627564159a7bdf37cd0d68a
ze7381253725a3880beeee0504b283144d91bff8aec0e7c1fe8fefe0db672f04b268a89ab5ca5bd
zf50777cbd10e545a14585c0f64d7e2d0338420b6daf2d981e4e2c103269ecdd5513052b248e9e0
z8f992b6820bee394ef256d4499e649bd397858092b5cad3bd33c8ac38890ef211d891087aa1a71
zf49a561c59da73534f2d7e177328e0a66c6fd358c84e4d9b105b58717922383de99f3c83168113
z9855e0dc9a2bb6a5d04e64d3eb06074ed055acd1614e316a636cbfe80b9ca8d7f9b1ad513a6b23
zbdf7391fbcb663d8a6df76c30719208680ea3b1eea0bd05a11db029f6497d566163a50d920c4d0
z89cf7c93963bfce236a8300fc29f183a54716a72a1f4150409ed7497304ac5da97c706111a16e5
zd3a5d676f5fda0d56da9c98bcbaa5c334970ec55cd490e829b5e41d1c212dc7f7ad608a565a8d5
z1bac127fe57832e426cc14779f5c09cbd04cf65607dd8c015d3cb4cf60ed0d53b18a1142405865
zbb58d578828517665787f4b8e97719fd7f1e563b2b24602b0e4a299936cc7c95c77fa15b02e750
zab1974e56ac2f342fb5db28c79968b2c227b58304e0680613a03c5e5e12035dc4273481e4fe725
zabaf5d5e3887b28f60be2267c689267d5b0441231f5d3980e40719c56f049f886d810043ffaf3d
za5f7a5858fc7fbf71dde3d919c6dbff35b5fb9cf8a46b1579a98ccb99491461d1ad651aebf86ba
zec8375ca820972abbbd53aac0673fe6d1cc9012081ea29d34dd1145994b016e81174ac813f0bd3
zea2e07a68004b5613e1e0b9667933761e9d8295a7617b6637f1abdaa6aadc6fe188130e643e9b0
za8daa1a6e16eac39489016d66a9d9995b8979d983fb82cbfd8a5bb40a759b777d2ffbd52fb7784
z422ed6cf67fd59da2345d78c513329d90aa862f4767ee87e5aa299ab66beb6b4ae58221a4d7577
zb970d3f273f0b408f7255c8a012fdfd886bb8666a7074ec7298d62fe68e3292abcf76bf94766ef
zbaca9dbbd4d5b56ff38285ff602976bad65a8d1dd0c6d7795c1e939eca2c3b9e451164d99e2b07
z8f92913beaa057b1f383068a8110adea12506bb8b6d46f45d42fc73f4385729b6e85610108ed52
z441188fdd80778ad93e318282874133549c35934d74f4ad64a70991787cda420ee26cb1b7e6e29
zd30261fabb65221626f5fbd76d21ea0c7682541244f7387b3a8bc0539db445b1e9517cf27fd634
zd9dadbee81c7f88dabcd809be1c51852e4c53d02953e9c54d8d43c1894ff3e6d0da0a89c979a5a
zefd844cfeb9b7a1b0855e8ec0dec7843fd4eda28f13a35c42ba0341edfe25860c43ff1987fc109
ze4e242937bddc2a105166f2dfcb409872c4f980cee3a38f39a0f490dc73ec58de218a533b55963
ze1cdcb2d75243c4c41b46aef75fdf97680a01e36aea1c7d7c57f17db312085bafbcb02236f265f
z3564a91f365110cbc7f7a3c06b19da4b4bb0a730414f34f4e5c2fcd2d1c190b588b91392656679
zfef16caaf56d19c7f616755f6a6f21e5e297c8c323755a0d4d1e080da1dddbccc5a779fcc042ac
z84860c803860c527902798fa2050cf55c22fb2d0ec8a03904c8919a4a9f6eb530542982d178ad7
zf93f74d1904c61576dec060975ebd2a39cc89f5bc394b61fa51f249fdc3857700275e80fea715b
z6d8a7de38f02e4695d79b190291413d1de564ed4d03b6be9daf01f2400d9c2ec164720a920391d
zf5418b207dd6ed8042caed0fd6272205246624be85215d75e4c1dcf32e81a7efd3067eed4d3e78
z424ddc006d75e1d56ada92b255e5901ec3fa4cf3c53935f451d6bf180aa23fae6197db42d48dbe
z811592bd2215e59767dbd3bd51c0db04f113a78634ab2778946e1b77055679519e5335371841c8
zdee646d435a85fc1444762e042c88fcf4a012ee39b276ce7613f86f8c2691bb45fe9350d3e805b
z1b2ddad528cdbc87fa7e3ab67611842ab55a9d2625177061462e0a262e06dc3ea634d92b10c266
z7094b1fa15c7ae80a5de13e249a993074fc506581c1ed9cfaf4d2205901bd6b833a9e25059b8f8
z9b8b68304e3e16e60028400ccba954ff99d0e5596d9c16264e7d8ef87a555d744c994af833c7e1
zfe7a0f7f7867934ecd9d937192d80941cf8c7acc48f3f842c29e481639b2abef80e6fd2f29341e
zb1a7175e21f0db9c8e2f55ce3b7e97e8fc78e3e4ad4a9dc9a1c65d8bcca2e55c1fa7d38c8db944
ze1fd68824b5716141d1c1441de5e5f11526a80ef4f4abc7cc2a399e840fee1e37c4321dae9506f
zdd9b1bda2eeb58245d262e1a0326b99bf13ef0ac29f0d737f5c66c311c00b72b4dff78168b4f08
zd91664e5dbd4c1f15c8c0c4d549d6c0d0956955952ea92d74a3eafa5982b444875e110fc5ef958
zd1889e596128c919b0688d657de544d49ad4b5e0ddf922be9be70373aae03cb68fb824508b929f
z36d12d15c576385d70309a01790be001b371c60a75f44a3170d96f65dce903ccb0ced6308ef082
z6d56bf3ad150c3a558f964a7b837fb83df546dcf15abc195c4ed2e4c482a6378b250210ebe9223
z840b537550205dd9a2d6aaef1479e3e74250fa6516934d3464cf23fb204e3aea6e8dead426df29
zf40d8dcdfeccf1d4d61d47c8498a45024afb80d900c4965cef864bb83dd00d5e35e91409302ddb
zaa738331a181107fa228d320b400a67c6fe1ffde81e40f73d21d193b9f5bb35762aec8b7fa0e73
zdf838328f22adbaf6f87fdd5275b930cbc4557c5d3031f9e782017f757511ef575d974835a6f83
z8451e907779e97bde20a3001ecc5b159bf8f3c3b0498971968a6dfc668c92b279d360eddf5356d
z0ca79534c94ba06ab63653dab64ad9276f03368e71fa4e6c06c512701462e05f70a973e136a486
z18453c6175857eed3887e2142cfd8b46cee6ccab9ab7ddd7b8f478c21e94a8963069ae40a27ff8
z92a744383ab124de64e98ddc2e7843793390040526dd6ab09c47b03df8eba1d3f546decad4f6c5
z0b69b9c62cede7212e1cc0283412d0dfa395c7f8baefe77f47b24d4c69c980447e25e18c6a5a2a
z9841e63692271c875ed0f8732176afb5eb3e7fab58daffe4f239f6024fed4ff148b959a116ba4e
z522db55bee1aef931496ed299a09c27c0a1dbff3fb105cc3371dd4f3d16acd9e8d3937d1555c7f
z8b71512a0942a8269a7407fd564f1cfa7c695598079fec8739623dec34b22cc04a2be6e1021c5d
z5c6298bccf3495d149e728c802e0c67df5b2949cba8926d0d74b556b05b549ddb1aea66a0c4db0
zc1545a33925d6046ab565054d97f4d35b0de5b266aae6279401218ccc2cd26d9206b23b4e234bc
z09398872b3ffb465acf31e3123168b0120bdc51d69d63ae3906aab5b5c62151342ad36e19c7da8
zf5fc95667b1ce98f926da348606bd6dd815839c7eec470caba3c4229320fafb882d3a916075fb3
zcdf5c12fee2585c9d8cc345678f2abc7e8113d85633d84b5b053b2159c5e87a03c97b3625e0153
zdc2279c37c38be4140fa4eab2f0352ad69fb835d6001d6193755bb68318ae3b44c763c15cf5fe3
z13ff3f919273d7d2f88c0f2d2032e5f51291555d3c9876b503f0484e54c8dcaaeec59bb0b02ba0
zf52962306a22d2f47169942da3eff88a78ab870c9d32fe0a1705eb97e575fb00049089f91637ea
zd664c09a960e1da1a612921afb3b9fb81dc61c9a4d408fef2bdead9eac9b1f41edfe12f4b83212
z61617857a4efe2368dce1b904c26f2b9125d5f4c2e9075c33655f6366d308c8c2f416be5035de1
z99d2ed5d4bc6f2b7e8b35017ef29203ae5413598682560f0d55f311fe3c6cad717449bfbe15296
z1d0362c68c3d8e66c248f64c4b4b673b9200b3ba03850dc894f804473d489e9b6519a3e8cf3fc6
zb872f0bcb8c693cf40b762f72b7dbf073d25595bfb1356cd557ea54de5c53bcd7f9752c41594bd
z43405612ba894f21cad79d4102cd90a450fbaf2debafe81ee2e4ba4162cef030060be81a07cb30
zc8fd2a5f0ee99553f221c1a26812930704d3bdec0fd97cc0d32d562e9d499a41716ff6ca6cb1ac
z5c9c691af0a55ad016f83348532565223e92bb7f753a4c5c75bc1d5bcc7e1e82ee4ad83226edb8
za13e7d031ab6ab95d0c68735a8e148b0d64e9059012480056b9d06d6cd88c191f30bada2bcff48
z0109b806cc42d9346803faf59df46f6c1d1d50ffa890329999d10976bf055ae0eda3dbfbedc19d
zc76760c123e9ed224369aaec06e9c9565a6d26dd06e90e41a2e1edd458cc930f1ba67380336a33
z11f9858f95f18bc8e175ea7a46877a0cdc5458c90ede5082e03b4e4008d833a3dceb16c708c88e
z68472a9abbeadc18c058612cb0775e1e614714d3e8a111f3e11f72cd7ffd583c58c1cc9db414a6
z44bf26fac7c7fc3bc4c34d752b9cd883aac31c648bb0dee83c46f1a3f8e85094019471e2cf3367
ze63a9e35a3c1369a01f0b59f30af073847b09cd335d5a43b560e92407f9420dbc12eeda8e1a9ba
z9f4ce9ac5da51295b0a4f574c7b9b5dbfa9254c7ba41b32a17afe43a8042f1c986ed47c7080cef
z8af305ecde69caf89d5816ecef502a89518e3efb9d080a7a90f45b98a291d31fe2b92f49efb481
z2a5f1b95989490c4d6dc2e31f9808f9e85c710e556f3c758632919a92b77d46908ad1d9a4ae079
z798c4f71fca9dcfacda3cc4e48ac92807f50eb552b092ec791ea35e645256cf34414297ffaa254
ze0cc5ea10619138566595da2f21e9a3319cdd67ec776dbb85c1dcc5cba7dcccbfc8ea4f7db7935
zcf1db89a4768ec7e613ad5cf8a8ee572a950321fced4e9e549011c323d4e86d143942b3a6cb061
z496e60840fbae97f1a2b799404e4ac889a8db8ae1ab790abd5b343996e1ccf136ddf593e6f200b
zfbcfca4fae71d533a2d5f7da5bd81de00ffe7bb2a145c2fe38e58259512954194cd7dd2c319426
z66c80fc97ffba7e75ad4272288c1cbeeea6bcd78183199e86316d49ab810441a228371090ff0b1
z7214f99eecdd7b365719602282db4fb9069411b6308b5c57170be7bb769b8bb2f93f50d720df61
zf305b523cf55c3d6ace7831ee183abc0a1d69b03935c60cfcc64c28799726d97d048bbe84043c6
z356045c150be93281d6a49bd2fe966f06c583125bfd85a63cae858a2e222ff58d39bb0b41da036
zf9902a524d2d73c637d374f886f3e5e31cbd353c791cdee43f18df1eeea4baf734e19ce337e359
zad0339a279aa277dfae958c6c6b512e4b2a3e9f803e9ae99552012c970b671bba2450efe287467
z1b7151c52e4d8da2421852b33c109f812e90bb912f326700e9813046a912e36db618dad9dceaf4
z79cd3ba2133382e1501dc587da6ea81d498822e4331d298f79673632220b9ea050c22dfdc88f5c
z55eb40ad412452394658a833ad80b383ffbb7805f88c5ce73d3256cdcb43228d85b4b5847042d5
z3ff4fc323987ae72c9ee0696422e745e542500f4d8960eea2ceb9872c0cc61fcc7b19d477ee008
z4b90f8edaecdfd6fd371936c468f386052d6d6a00f3c0fc6ac65dec879fd37789d4695b904b6e9
z7e40d99c7fff1b7a03c12c371ad7a43ff4f5b7c1409007e25037f19586a2a37419c1918e663658
z30cb65eeb21b2f77cc36e5b4d2e694e9cef4d42d7e53f2b328ac5eb6f0f75a66f21c0703ef42f0
z8eb2eae2bd5c1527627b4c6c6147d97900d75ccf0ed0b8a8e50846db6d20f6e2ee39f586049f11
ze0cb77aae784f1dbf930b552207fd9fe59b49a7c94b72bd39d29836be5d90116248e5bc08dd7c1
z8ec63407024e9781d0a027d801b0889a5285e85fa9063919995695a75647abec4fbd43823b7bfa
zb892e4223d44931c935be32513f88344f90350c85ddb2f9281d43f34499d9c80a5803a40f96cb5
zd7b32e106af63dc14d99c582df9b408d0ae23cc8570a7b833a47194f723d03dcef21f994a935fa
z525017e5e901b9cadd39890ec4dd8f3c364dc27be3e301a9ada3396ffeea8f57aa6a034946ad41
zbefb38bc3d0bc385ffd15a03d60b701a85b5743b8eb845754fcd64d722c0e57ed16ed592e4eceb
z4af28b2bc4c1ab7b195038918a068cc3a0e1145377827870af1cdf2159056b08e980bd8a5cacd2
zfe73149964663d7f1bff03db2602f8cabeb4f67f4ae454467560c0c7d3cbf9c64c846898e75ecf
zd8c4545fea64bff1bf6463e93f84b8c9ec4013e757574c2f4e766a030f5577c2e81d31114fcf7b
z98ee59b96d780f0231d45f44c7fe6c3f7804cb2cf147a7ca3221bcfeffc808e351e438dc38dd99
z4ac0921f06c42a71b3404ba6a8ec0e45fea98b2f82f33b32257b7759218a80dfbb279097b4f6a2
zf43217669881db57317069c9b78a58534f02f9180a94c61656e8131b6629fc53f1f4e5990ca782
zed73c9bf666af41fac2dae253e70cd9a3bf17aae2cacf5767d1cea274ffc7566f0999be5c5e84e
zd92e0a1f5eba7b170c2f7a8f651dd42253bdf2d28f8f39222d379c99a19d3851ac1cf587ffd7e1
z57f9abf8521eec13d07ac1d37c0fd01009bd2c34400071301afe1b3afbeb30ac91602af28ee715
zfe5e8d92a03da997d3a73db68571e2d3359b2363c5b887d52bc9ee19ef2d8fe6589e1fd7ac9ef1
z2335111517e41e026bb663f730ca07829ba77914b3c80b73c8b21ca6d6f5453116ef6cc16d919e
ze994329d423096958907c83d62f82eae81527fadaaf42038e985ba64dd83555a97bddae9eb8333
zb3f79d0efdb39e58a3d29980ee34b1862e62efe31a5138e135cc6c1cd4b56149872d24b0ddc18a
zff2bd3588797b9aced012d6eaa54e94e98f6c67683538bab6202406dbb2594280e66caca9a8de9
ze47590ace726d444974311f4c88ebc1b85d1fe87efbb1b7ea8aa2cb6493fb93460ea09c6e3dfe9
zf3adfea20ba43a2465b1ec8a0aac2d3b4343f79869c9002e3f3c549c1b90ae753146908ce48d7f
zb295f0fbebd58693e3897707519470777a9d7c11f0214048d5df586ad2388b4cdc8bbcb76f7e32
za3642545e0e34da87d5c9ef69f23ca169784942bb7f923772912b257889603f1c1be40628fab22
ze44d29e2cc1b3b883b8e2ec61fbdd52b32c77ba2062b10bb608dba772a2906018d13806446d81e
z8952cab9e2f7ab317bec3af72acb6fe161c53a7a318a0bff07b3a6741db2eb56759894e23e1b27
z57ec5883eb026395e2c52730c133fc80fdfa0ad3491ca12f60c6e04917ad4b6237c98bce27a4c3
z5b3912a0ae3513e656ed5ef5af5c1770610945c07c4fa7cc869820434a98d23eab6d63aa6ae033
z7900346440d8ae8f5549a0dc275c50c6fd5d8bd03a1cc809ca677821920be1baae513bbbedb26d
z09c48d8fef6fa543b3e953f8aa0e13b039f974109a4167bd24233844e2d86380f9b0f5677d1dc0
z53132f199d8c28e4f98eba9f0376ee8c7d6c66f443c2c8d0d2cfe19be9bea96023ac1457521f8e
za925d69fb0bb7f5a5ae358ebcab0660ce170c5da2313979abcae9a5ca2e965d67af32fc39c3a3f
z4da125ea832c21315be0d2d034efb20716479a3a1c503671b195cfcb2767f5e34c625918ae13a1
z4aae48977264f553754676875cc0e9cc329121e5a9242466894f255571ef8967f6c2972fa1bfd7
zae610fcb3aa7a7db7dc8a168735145f3fc7dacb7b154811412eb0f9fe2e9fbd28658100867a5de
z115047e0214504c75180c6aa90d49318992225c9fb75393f27bafd85ab56f965bd908b63092aba
z81b8b1497a31082daa6d1ed61afcfcfffdfd1e786cbf9290c07b5b7ce5ebc72b10919a95509d35
z8b54cf7f6030bb8b2da2c0ee80f3438016364d5241e5d2ff98c0e9e19d355c31fc447509e08ddc
zf70b96aaedca4e609e682ed92265f6314b6e0d76577d09154d218936e317238be041f1f2fe8c6c
z8650cdd1210ac144b7021c8795f09e79629f3da95683fcd1ad305fb68d3ab139e5e75a18e5a98f
z0b891ce629526ba68562e09de50f1327ab11c5efef71401e61f7170624532e436ae0cbe095d451
z1e7f01b525abe25855b493161f7a33e73ca5dfcf744c69c7482028a2a325929b93972a6997ae53
z0fb600d44e65e3368591a40f398f9831c6407d5f6f471114c49e53fbe9ec201d1c1246b329a311
zde63ce3de8a6d74a555ccf4813a6eaf030d2993b3742d75901e8e317214aef77c797ba64f2f10c
z3b45768d34998746870ecbad2245c11720d3bc921c065361da314fff2a9888b66f51ffa1b03710
z1584087b2cc283f364f169816a6183dd525ac2c668165138c9b0534313a86899f50a1b16b747fc
z92b251968e268251000362a910676a08d6b64f881b1ee0c01153525ce7a69504e1e77ee3fe7c52
z8b31acceacd6905c043f09a9f9896a29a2435b459a9b7cc0ada73ad0283cf46c5e57d851f2c6f8
z1f767450c4c63546bd6159331632e15fbfe9552d290beb6c8e557d6925e23e55cf0fcfa65fdaf5
ze3f81e74cb8c2449a118643e8204cad45f4beea0236e84dca4f0781b19621889f80ffb74b297cb
z533ec7652677444c7783f3411a15ed6e3b60af38a7b6ab9dcf2915181803a3b1470f4638853f18
z3e2262c0794a699ea33de1c614b082b76b9d99c8eb7a53df5379e12b659d14f33a9d276e0af16e
z996ba425763bff3c3056b9611bfd474258f2c043c8d9a733a9b0b28c3942eec290cbe6ea43dbf3
zc50e5820b5986d319658aecec69cb675289c3e35f1135bb84e5e94d0a04c6f4155a3206cd6ff4d
z4db26f03ad94cd7c42f255a20b2f6b50d99fa43686fecd6466452bc3d8d5129e337d878aadc4f2
z63bc9a37f06551ced4f680aa55b7edb91de9bb0c29e1029ce1ab1216af3a3f2e800545dc0c3087
z8a305aba6d226dd244d9fb36e89a704b0d888681965d7e4f6c32bf42d8fc26f771967f7075865b
z46ebe52f5bd6e241e977e934f00961b008f1fcab35a673a301c6395652cb723c93a28ffb8a0d67
za7bdeebeda1e3b9d42b9333694b245b2d9aba550853ad0071270140b284afc7999c89484e8a24b
z754ad5b5dbc536c0519c2535f31ab05b1d44b0b61a5c7aea4e7f0c737ea44b9dff7d7b08c9002d
zacbc5590e79d11acf9af238b015487baea363a0f1e89844099f497930ea043cf949786f443e447
z50178cab40eb0e8947576b4c3ab5b03eaffbb9202bc8e724f3c7ada71fb49079818942a82061a8
z2ac2b0c2d0de828da411e5f804c10ef7ef02af937a31c8436b12ab5956f62bd99c2a12334a2e63
zfb24f052117bae0a2acd643799c6781104c643690805bfc2ecad3ee0171fbed222beda7ab384df
zcdf76f441b0ba986ffb7e2ac6d60d05b026a4c77b9f9b1b03886d8aa69eb27ffabd3da9187bb64
z06c70af105c98cd85c343028fb9843770bf358380c03029250f49aa4d3becf17acd0f5789ab87a
z10de664901b305bd414f1953f00e39a1a6b34942851929da46c564292174dc060649ed6343f7f5
zd99d7222090af9a2f86a8c747cb7bc62342d79cfe4e9916f2455de1ae936c28ef6e490b5ec9327
zbdf9fc04b6cfb7adfd5c7326b452dda488277dfbac635feb087418fa1614852f6df74e6c538373
zb957afa4f1c34fa21285f71368e77f3300a06320f1f13af9df3e7e68f58cca7119f421bc320c0a
z4e7bedc37437f4d2e66ab6a6b7199cc8b1c8279fdb779d5e8f1a9006b93f8626fb1e971ae06dbc
z6cb9f093857c09c84d11c850607b5e8cb7aaec570b847eaad0fb9f384e3bbf03932543483f550b
z4b4aacef7fa05cf7b0404ea085d1c074c8d753f2d94900c8291f417043de47d84303f0d430c221
z20d694563aa719dd208e930ac9621bc3ec72ad60ab907c343a512f0c37939a7a51c5e767044d95
zeb631146a1447cbb657cb379a38c484c699f7637f36f80294da99a6d0e00e710868f5c472b5f91
z6733cb5eb7e5942a49764e3bf5ebb15982244bbd5815faf4ac51c7fabf7649901d22793b692eb0
z6316beae98f0302d6627d2c1b4185cd8da62ebd8f2aab5ff69f1637e3ebe65979f3fefaa795e59
z60e0eef647cfe9d2fb503923698305e4d88ac7c94c10f25a5d7e0a8242193154e516109fe563ed
z56361dcc38bef5c8752d9a54d0b5c4219da9133080d07c4ed69046d552857ea7ac5bfa85db9f43
z6ab33cde1c09460d8886030fc2d16eda266fe93103fc8ec944adde0ced7046372e9c19eeda4fd0
zed319ee7e9874603ae0f457f02292ae53dcf809f82374e8197732fe3ac4ceb0e46a8429944a3f5
z0484d0a281663647c8accf4ec24dccc2061dfab3048c2d4dce9f944cab7f0e6cbfed8bbbcf88e5
z169b172dc9bf8c25ef40e58373ac7148fb5533352e50e88ef1b97f2850cc0fe361c5a55e077015
z6b79eb0395d9666029546c4a40f3120367f483efa74c6908f9463a77502ae23ae2285fea953205
z91eff84cdbc314a0b8111ede28e77e52b765313edfbd477b33f9ec21e540bc5f0891567bcefe5e
z80f4976fd72df25b88542959d8ff4ab8dca2944ccaf4d6f28de0888fe864319357594f5bb87cdb
zc2c915edc2ba5a3b47f25b55cded4998d9eeb5bc6ab49a50d687227263b9b15f3c68f74421d185
z7bbb27aec82404bfaf2b4550474010cd3451ec0d5c5a01d701debdff21f6db11ef881b264be67d
zbd93c9fadceec2025d249aa0ea1ea58eea6053575d7fdcdfa2bec268d5d1eac1044c512e5503f9
z3120cbdaa6b6afe5ab6addb067b01702bff97784d61c7aca250de83972d775b47a176aec766bf0
z59b5b0af41eb5b2f2892be9264dc74f704522ddfb8f6bd8823d0d87ddd0c41653929e1a8ec96d0
z6e3a3ac4f2098ffbb585a3020b80d389198ed67a64560bdee81481af9fc3a1a358fcf1760e5893
z369606f8ac6846cf1203697c9ee9985c8c4dd6f7a31856899d038528280b9287216888ca24de92
zd2eaf312ec6d20af9e6053c92a1369dcbf8a512ac0c17f01626ee41ba32c44afde24b6097bc90d
z54f25f4e7f8ccb552d92f999cff12b31be99fd68d3c7d69c15d7e34daced436bf50fa684d6c48a
z1df728dd35e0ca03fe0274b7968569d1c2e0e1d876b6d89f5b4d115d2c93adc0fb7c02ec4c9dcf
zeebdd6683c3cc30fe2ae9e5a79b4e5572095bb1d06358628b697c0981424cc0f72ae1e934b3e17
ze03204f3caaaf80360d51769c80913c42bd3f2dd950498f39af629c4d78b425fe76115a9f0d768
zfdbb5d6efe8a5e7b2a5266caa8e2a456cc260561feecdc3e804abc27fa47d0cfa77d20b0f06c58
z499d58c75de28b32a0fc59563512a3bd0d3609789c93b48d5350c7f013c4c892ac1764ea3b3dfd
z63e929adc7ff3d13c9ece007c0ee6b523160443bf6e7060ea7a2dad035e87e1dbd1f7c2d3168eb
zdf682f143faedb0367078fad585d0db899ba2d3e66aca5732c4b5d8d1cccc010a9fe9d56958218
z5bf4cf65712c370276ab5547b27f275114eb8d285a723b9f2e8a2ddf483d55589110f8b5e66aca
z3ed396b45926816b001a355509f4e77f085760663eb63d542623bee316023d41f11ecfc54edfe0
zfeb5e22be821375f6ee3fc6cf569502b1e541d8e0ad64e49c11fb3830dbbe74075431bd6593094
z7c55cacc2caa4bfc59720907349525117b4ee70df4e005807993be2608cef62ba88823c2975262
ze57d7438a667d34358311f87b920bb082bcb8a15e2f5b5c438fab5f085ea0363f0ca35bf79bce3
z874e49493807d93fe097ddd5d914d4f2c744e9191c8d8b9eaa92581cd2a41007954becc69cc7e1
z47f211576c61a29c5f0d54827b77aa155efa4ddb2008d2943f3776a9dee5b46f8d7b339902247f
zbf72e36092b517dfafb48eb6dc2c7650fde05ea2863cfaaba778a151f4631a4416ef6bc4671359
z18aa3ffe6c539057f6b3065f564773c240734c3339031cfb9e14228625c0788eab8ab0933883da
zec46513f85e4a0617b9c1762b58f9989a15e98939ea4dee4ddd505c22ce911a1125ad8e525ed58
zd6b564e2f12b7f2dc975f049b38dc01bacc39c520488a41d0b5283fa03bd6532ce8025489eca3d
zd6f4bd26d81870602355d3625842fdbc8dcec912a5067fb5bb30bc35d2c9eece57e01aadda735c
z0c7073bcf0fb487780f111ab6f06ee5731681c4a8a4decc2837a19185edde601ec8f4042a75fd0
z65ed88770303a177a5cfa59b30f5109610e38d412d419d0cc0634815dd1c9ff7de6c985793777a
z6966c53ffa25a530e8fbaa43d12a3696764a6462332932dedf9584ca83a6dc3c7c87499899bc5e
z9386909e1c9ac677fbde7c31d2d839e34332e45f2583afcf9ac76af178d67043b243606b78ec3c
z11ec02000c3fc6de6685799ea2f08039c1185340f01d18bdb3c40a48009d8b6f1a855911dcbed1
zb30d01ca062a22d343cc19a35977d66a63e97e7abcd23d3e99ddac1bc4e24cea8b558b1c02a8ea
z880b2a5f9d99b1abed988a4b57dcbc5a4b8e652d812a5d7333476252defaf222391fe910cb2f2f
zdbd27f35ef9e245945cd19ef7c9fbea459fc089dece89c87f10fa265a0260c4c108c0415aea307
z4ffe8167054147b4a64266a0547becf9f549ba0a6e2d4c95c805310e36a549c89e80794680fe13
zd7ebe513ced9fcd88d1e8f405db875fdf30d1b1b28202b8f5f626e86cfc7e8c3b4b1c77b547e77
z512ba0aece8397a67d47197ac9f488327be03469d0dd08e7cf59041a4a0349e234c5074ac874e8
zd2231c7dfc2270190e7f9bac09f5339c6c2dd5a61fc1cc924efc192e541dced33ac11bfef2b05e
z5eb801af2825fb9d0af5720bb3b2b98bba25d2c2a7539dc5c99aa612df32c02d94040a38c8b828
zbd77c02ff00cb4758151db4d7271f5a328a3f3e0c83e48052d5cbe82aa82267619c015d65c7e62
zeb63bd641ed2e1e7743cb115ca832c093faadef1ac970c8fea51b55da847f89d421c8ac320e2ea
za21235518a2175192c99cd218655fa0af1e8655f193d876011cbd30892f437a04edd72a4a6c7a1
z857944bcd570bd658a3c387e8e0c327fed93b143ae4c228e624e0096d0b7caac13df8b5b484694
zb34712bdc059b050b30352c3f17102446169ebfc34842f30aa3436b525e45d8d980bb0f98ee58e
z6bd2f63460f444bcf260d951d1cd7c3758398d0bd58d53157abb26ffd3e699969a9cf8cb981461
zb653f22708d7c85d93239cfa750889f6d2d5044402286aedf9898d5c9af705c1b50689c270b52e
z0929ee57fd0c52e5c18ca046ca1afabc7d9f3a019713217ac2efb293c3ead940b3e80e6074af16
z68725fc74218a999369c055a8b947643a957e1e0695600e9b272a349cabb883e480755add04247
z3ab20c3dc575a1a3ce08ac59c3f3bf37b25ab03134c9d284cdfda3f56f09cfc87cdc42d5f8c0df
z5e3c836ae59df8368f14e1070c1383684c008dcf74e476bdb00bddd836946bb35c21a44cb5bd48
zde5fd091def2e6063cb6e7478990aa19f068f84ab969c5597f3611afcc874d2483970c3043ca48
zfda17b4d0d667b4fc23c180cd2abdce6a36b5e06d54c62328f6f19094c804c012deaa4c170eadb
zf4548c116c6a895a4ee0d94dcae31d5b46f246f296d3f100a1a58678c4f785b208c24a7d32e171
zd21fe35c14c1c9536225185f9de88fc5d9f9656965a338d22c2f9d302d762669280473d93b0123
z95f025fb3604bfbee29e67d3a68c9570e63f021e784194876f8285280e703ba76927bc920370bc
za58ce44a01ff0e43b96805b4c0931f64b3c00a40629f7b2724e6637de9d8597b865dfd3248d9c1
ze3c01689bf4e1f45e5d724cc66204e1d25267f93df058c707519018c33afa06c5fe1675eee2c59
zbb812df62decc71d0cc3d9bf42b3639ac744ee4a9326c1fbcf8015c6153eaee16081c95f57b16c
z0ede8a8ea3ab434cc577af78018d517131a7ed344cc6c01d183b5b16586899b85378dacb8b4e33
z2b2318c9912983f6a0aace5df8a9cbfda214255f9cb7f58ad61bb8a8b4f6f171f8b14a7b251fd2
z5eef036f6c81cd63fd6754f5fcd6fc1fd07895398750f4bfe7880dc53ec2bf0b463ccdd857a1e6
z9b9dfb0e3de63f6bfcc606a05241290c4eb11c3d68ee1318ecf657237733553af003e2bc74535a
zd819fdabfa8eeca13f054f0172b339121784ac8ebc9f7f733182f3bc7f0e166b6e285d0b6a8d61
z2c9429a5bac0f67f2a1ffced7665beb8e65576b522a6fb6d785e5207c323a46253d787a9e4fad4
zd92cd50a96abc6de205bf7c6d5db1642e3cc7db16781feb3b8975fcf638d719cac9567ff9445d7
z411bb920a65c8105e9d982df8cbd7ce073e0a2f89a1f2f9c255241625eb61eb298b90ea15e967e
z670c2879865c2ca4a9c6f3053c96243c41a1c398e45bfc8592f0bb2fc6d97c324d738ffa9b8611
za92a8852d3c460bf7cf5a84344ddad8ca6b8eecf343d1d220a0816043cecea05278b7fdffb16f6
z11ac0fc4ddd051152a1298a5c1c7f1a95ca72c1c00b05ed5a8dbdb1dc23876160c90398965ea35
z228de9d644418021a93317ef636c968e09904ab9fb94cf2a9a1f21940b85708fa10e53aa4e9b7e
z4c5e590e7e97965d13b947eef3b865435d48291f698aaeb82f1222e048385baaabf2b3e6cd518a
zd0c51a5fa779746dab28ea41288069eacf4156387b73149b3c13a37c5bca36644befdff617a450
ze230094388d18ca08d3407ca8dd455a3830e34250c438b3390dafda752e1f26c2db8b7626db77b
z0e72687874ec70f44dc972868956d5424d639c9b874fa023f99090d85c16492c9a6ad0223f7495
zb52852940c9fc192e27348bb1385f6fe4ca49e98828d9e254ad653e8a98819d269f313985a08c2
z111883cb109bfec6e205f291152f5aba9fd433fa745c64dae55ea236e9f92097998a91ee1207b7
z655925f8d96cf7019a845b285cd3f873c0a8c271d459b937ed61499153e886a6aa8a491b3bd93f
zea90b67f51ddf0ab6b9f09285f9402dc895db62186994df4c2a7ae7f01b3993d840e70abab0e27
z7136bc2609a4ecf1757fbd0af067400a86098069d7f55b6db20689b0df3ad7cdc85f054da2d020
z9d8f18ffa5faaea8fa16c616bcafd5c6bb2b6cf51ac11ad1a2bb015659cf7e4e4d582f643bfc56
za4772983223015d0ce97b265662ff2c6f2f567fbc389d059912e03b24d48ed5d1722ac5903ae5f
zcca720b8c7184ca33fb238c52f2f0fdd74b1eafc3b6bf7ab920314119cba3b82c76f4796c2a620
z33d268823e8ba579a7f650aa0921607d0d43fc935c93a17c5e9d2147a4bc05437de6675d43f487
zaff4cac07921f3b13034914a6070481fe1e2c04f3c2d09894aec05471ace056a7334c178bc0768
z182275d8802aa1cd9f33839995700f6a5391ba790b423e08ae240c691a2de839eb82ec77a0ba2f
z2360a27835f34ebeefc1f80c47b884636b77fb4c3b202510e0d003428d1e1b935512a03f0d1f4e
z0d6e3b22a392dc8152508d88d3359f3598cdbf5a7d6f0f10043d4711d44b763bef9d72304fd67d
zca27ae337a91042198eea3117308858122513ea362cd0b29d53708e5508c0b65846d5ebea25079
zaff5ab21dc8dc02a9e646c27ab146093167ae97f08a996cd1bea83e701b86bc98ff43cecde60a1
z181e258b5c1b3442d4068e5f2f2ce5a8bdb8d4501e42232bbbf45a70ba0960363f1922f5f43e40
z2edbcb22c8e9e5c0dbc9f2473534b9653fd5ea2102462ddf22a12e965aa43a7306cee83ccfab54
z19a863f19770a1d9f463ceeb762d833e97d93510271fb44bb21b381bd9260ce42e8dbe21517ea8
z233089c1a630055c85c9ac3528412fb9768c81b742fd02652718742dadd55d8e7457a7176a32cc
zf6d32c11661a0a4127f4899a88000f1f93ad7adc8958a331dd259498c963bc0e07a80b02e34041
z40af4962c4341fab368c2388cdf0f02814b0692c8d63894ec784f6e6c938b3f590691ed8b54537
z0af5f040f34bdc9e772eab8bb658edd8bdea610cd0309e82443a921791aa77b4bc53a84eb6c82d
z280ece98ba16b1eb226e37821766defb35138379bdbbe6a0e207eec2b232991502ae45c635adcf
z295f01f94332e94f49c8f93b8494f132c211294aabde9d286dd9a6de2ed37f07f57a98f062b4a5
z27c4c7b7d5a730d259442a6e0666c19da312c614532535afeba260c7bc4b5bf3f0a6d11c618cf3
z5817ce4c01d319898024bf6065cbd027ff8152b3407866cfe4e9856facbb1812b31f85e9ddb8e3
z719234e9dd8032e1270930baed134ae73afc44f24658565cf261496774a53a214dc6318a64c3f6
z5c3838451c70c83926ff341d6253f3e23a65b5b4e0713934b87dd57b040a7b865aaae5c2beabf3
z88ff7786aa5c09e2bf372603db7b3d612b46fb39f0336cf95d8dbe07c119122ecf3ccc6293b5c8
z733b94c9af86f75cc0cd251e595760e6bc2e17e3ccd2b9639a4f2a9e4e598f151d31a9b0f0d9be
z3d44c276a342235413518be35708254d5405df2b7dc10e00de79ef4946059b50ee0bd588ad9570
z23efe35be7bae24e6c00fc89132cdb7abaf49121281da95d8b8999e734afb3e06966bc3e084c71
z5b2ae29e7583ccd5279c72291866b4c3f8913df27a8f3e7f62c98e6c21a869fe944a3899a96161
z1d8e173f1c7885822d3c05b23459ef53fc47f76f6eefe1c3ef622e0a03df9340b9e2b9178a53c3
z6eba48c9b97f32a7afb81f7f1786453d165cf79470885690e48f73c8eff37bc3a054027bc69841
z8381848c80b5be013d3c0e5a4bab3915bec337b6485c598bc2cc774e63d7d049322941e0fd1aed
z6a3a5bd3685f5d4b729607ff3bd2e1272f34384fef139ed4f17fb242209b846fa84ea776278dc6
z440fac575ca181f0876beb0742e9660c4f74e57969f322cb1184f7d92dd9ca12d19f1db29e3669
z26d6b7c19b36f46427741965093319a2cde1a75c6195544ebbfd654dd0e623773509cec361faea
zb5e1bdc68df82115f83b2dfd694d6ec4c5ac69f99bbb99a7861a386a3ee0a6a42bdd8d980d1ced
zbb15e901a2348b9c93b5db84520f92c1371dceebcfa91c41d242ca35c8b06e133b846b9b14a912
z7c0db8396844a3355f0b6a4848ed5b02a8fc2459d010ef4fc9eccb93cd4b69fa7d85c10d39849b
za4e081c80a0d05d8824b7310182e2e5c4316501b0d89a5cd5c73fd2d1e3bc0461a27f116fa89b5
z6694e3c69907986163e3aa681fd6acacb15048a8273147ca16177795dc9c4ce592206a819f8417
z77782f07395fecff07d92180b44a44988bbc52bd81492da163ff009a062f0795bbb870704b454d
z61bbf976d951a9192eef3516ff669ee111b9f05826560d07a5a5c94c4184eb6904455e697d7bd5
z44e6a0f702eff9b81fd517372aadaab1194732d9de47ace8b0498395b2094a09959aeaf3d5ea85
z116248785fdcae5313cf7e7413c90aeb4dbc921a7457ead2d521e90b49d073e3557ba51bc95278
zcbdedb675997d45f39a83d6260ac224cf019b50a4b5366e3508a5c9d3e0280e81b5da4a6893eec
z770a9df907a0762dff33d586c8c5da1daa3c20d45581210b2b26855f97438cfed5444a55670040
z343911233138883754422c3aa7dc57d6aeb6066455b54f3f69bf4899290e16d0bc4f19f24779ed
z777009ceec104c556715798594988f67c5154eaafd9bd0f504bbb036fc33b1807cbc854c4b0122
z81489eb0ab639fb3e44a6e09021f9b2f7ec31239ef53c9f6293edddbb4466a12c75cc9bfcf12ea
z4d204c2f79d1b99025741e30677b044012c9dc72c8571e103bc4769ce53d96c614aea985a551b9
z6aff3f5e2856a5b45a08b363b88662385c2268ffc544745b399e7e6262397c1bd3a94e29646090
z7914e4f5f9e41ccf1b9141afee9bb4121aa2758fcde43d2f0a37146b2d25bd2363b22747b1eb2e
z223cbd12b8355e892b2a283c6073d05a575bf9a0bc9701802fda14d90c6873ab761850b5671c41
z6f6da4c326c8451361125ce7f0c6c0b75369c78c1a894f423c1d44d11213b32deb170fc8d49ae2
zde07e23724d94a9b6df088e8fac860a5730b4795c06713448f15ccb47d11c7763a06e8fef6d1a6
zb3f0835278b2d05e372af04f6a9a4fd36336e9196f5eb0441bfccfd99756ff29abd8e0be3b4c56
zcfb5ef16464d5c06173b07de4b0125c4c1121fc1c62aafd9d6d3ee3a0e5c4198fff61a8995eb00
ze6dc2174d1436c47bf1fe5f44fcb8260b72e5a859cfa68d9183421d221b8c97b11ff15af847d54
z8a89897d2839ee967afee387c7b57b9b84f5be9243c6bfb571ba82cb267631af4bce1d37fc6b5c
zcc9a032ffa9053ecb996626b054d48aadb55c67c7898f963af94e00046c0b2197ef489a4a1fe2e
z7b211f12f40216523a9a4d1298bed70efe935672e14ece989bc54a62af89e50cac37c1a29c9970
za8359a1d61373821da2b173077538344323dd28490bc52ac35a0966f79559eab8c339ae03a8549
zd17ba5ecd0e6c96d73874e7b55c1217ba36ce270ed63055e16d7e4a72dc47ca57099d107cebe77
z63b260163328e75478d2941a2377ee74d5665afcdee1d0632df700580b21c06e29d67adaa2a1cb
z65cfa797601b80f0340dfd5f4e5caa51a1db47d99047c13bbb28fa6ad3a67ecc453a5a5fc88310
zc7d944a2a5aa7f18cee24182185662d27119477adbe4179d4b1ba4e8881fe94ee81bc995a5d136
z858449124f84fc36f6199f2fc9fa0a5148d95f5ab45b25c74d5707c23cd2146d1b44d85507c041
z3f186e6ae9892dd355af6b1300dbea0f3f049cf1c4921154f003f5b81687fea012f9eab5559151
z0916789b48a9012a40b68bb33bf20f34cabcb565b2fa5a1acc7849bea43a2903b28f850a30130d
ze8c4f846d35b9ae5556a40466186d276cb23040adcbdcc7ff8202bbf785bd300be1fe55d8cc3b9
z08012d24305238db1b254d849555bb9232191cf3ae971bbd9ef6823d3ac4fcc6da68872e0fa1c4
zcb223d07767826f19f86cc4d68656277a840322b9d5022fbedf7ca07c8d5ab12ee0a93cce2eb88
z457f8fa81bdba8dc7bc2e249cd442b2591360efb57c01667665e725046da69505b9e8583fdf6c3
z35dab9e34cfab13e1bf297888028f181f33dd20bed6362c08634076b95545efd4aa3e3e8553500
z0c70166b80d98c525d3a54811b7c14b8fc8ab652db871d1006648ed7427df89f11fa1cb15cb602
z5814b06d7e6ccba6036f0ca61d514db73790b906b04071e03bfd0912c49f15caef4f51ff60c1db
z276e70d0a0b36c4d945e520fa752c05833bc9ff6d34154af29698c0304a7f61713b09aea9877a0
zad9708d9cd434ff6fa34f709f9547ecb3c32aca20c9c51917051365257c27bd0712128ebf37a91
ze2df9c55485c6be3e254b02262332d81affd85188c8d1c34d3085df3b3bc6b8791104e31eb0d58
z06724e82128b8c3f1dea476aac82474638f492ff631ed451c61bddfabf6db8f009512413f8cff1
z13411fd2d84d7a838477cef581a8af6b3204922528d1e2ab1afea88b1f2c97bcd6e6c6e6f240cb
z187ca36197e613a90476729f7ed219279e2e412137dd23e59e419fe2313a12b55566d07dc622b1
z97971970e3b5a9f739e4e50f4d48bd53885e108dcfc68c2f5f6b144792b9aba2b0fbfd7cfe2c98
ze8ec1786cd9e756ab453a51eb5bf9aaa126ccfd08bc2a127ac36f9fd71648cfedb4495535bf951
z36ef4613ed805e3774c13862148d65c33498eaa013c6364fe5dfee8d37b05d241db267c9e1cac1
z9ed9899ed75a4a3c5d28169053d5b2767727fe6990edc3d891d403336faec17e7c08b3b292afac
z26be100ec64393a0728bffd8175b1bb5c934f9c1873a7c40919811da5d7312d1cd993b0ac26d82
z4f16daa5a3fc462624cc43e9ee9b1fad0bd7a5e56824c0eed9584a2b606b486779520491c80718
za0797fcb980cd3e19b72e624706d3f07e936baf355dc5a0d7c4c59b45f65e9ff32b24edcdd13c1
z1238006e23bae111a6fb406a74c76c6938b71bcc88963aeefaf8e1fb8747c12154ff8852a74293
z0001904ab53e27ba02dbab2a816d289b7ea227a466a27f7d8088c897bbd446ba6bb501509913e3
z4c66e9e831ae2f2c6b82b2377669e949910d5c25d24e21252709f0d806729695ac9a1fca002bca
z523031070e882c9b9ae39acaa189772970689cb01896a48120a87773aaf7b4e2b9c41e02fbd2bb
z81afa321b1ff4877c5ebb8e5aa54b2a08027c66aea7f4350ab4673d9e3ea56fcfa302a3eaacda8
z97f09ba7ebe6cfcf730d11e18e5952654c3db4a7b5c8875f01aa3691935b1531c03a0b1334ff43
z6cff81b8f8343ffe6e52e30cb99ebc6630cb58199be53bad4ecf107fd2ec4875b782f2f277ebb9
z47cfea0da098427db55c64d830f0dc91f4da5a180fed512aa8b75105bff8bec175027e79e87c21
z0a7fdffe9c9c8bd502dffd25d96cbf4cd36f3be4ee3a0a702877631d5732cad8f258dd35123e3b
z816eb5ee647dbb7def202b1eb9754b8b74750670c20e778578701f8d04dfa52536e0c7be0f0f50
z602ed16c23b4cf94cfdd3261a067590f0fb7a97628cf3301344e28d863bb96b1f17ab9f6587651
ze70afb79a18b3a35492aea014d20d04f71f60048b1a40f4117523af459dea1b25cbe2729cb9ded
zc6a491216a58576652ada6f936e470b26afcbc856aa923b5cd2bc88652e92f6509081df198d244
z78e01bb320c19995116e52359510cb49729c19ef61d5fcd99fbc8e9d87c25757e1c6a1a13ec1ec
z70dfc6d056160593bcefbf627172a5c9d665bcbd4010049dabf7fed207703b3c88ab8a1ae939e9
zf6a8dd2509b384c7a6d99df946dfef95f0e38c05b10a28c1922a30140f01eb6751889efc1146b0
z5ff7dd1871e17ad829f1cc07d7d6324071dabd91d59a08023fcc5bcf355f8deaa270f8082640a8
z7d4da5aaa777abe0b8366a880e48fe691e9bd334d282bf7cfdf3b57d87bf577d4e6c9fe35164b3
zef52df83237658fb04b13cab941b81179cdfa128513a2756e3660baf4bcc21cc812022b6c776c0
ze80f0686e7d6ea5ca670afc087f8ce37afef5e4facd7a7a03f23e07b49b14a217f8d5e6da5302a
zf836e2502ae766e0a65468a642253be86fe3018fe73a72d0762861b5c60aef85bdc0e2cd52fdb9
ze6f0560f04485e0f465766234b9dcf44300ec68282d481836ac07698bea7d8c6220bae04694ddb
za560abdca41903de0928c8a38339eefc6c1f17ea5e21254b289440413c18bb56993c4b6e0e32be
z7404fee84ce59fc08d22a1088ec7e79a995a6ed02905f4c73021711614bd680a76aeb653651afc
z535b0e88a1b3c340adcd867be6b2abcb742d39f9b91cedd62372e6aa392518eeb4ba101a75bb56
zc0b81c9945cb9e392fe7866f0a609e0d8d5b2cca85090a22cba7ef84df8e79cb8aff8daf092c75
za91816b31fd28ff77ce1ceeae46267e5d083e6d7c2208be8d90eb86e9cee8950d7621efc4106c4
zdd051292ff55b46ba8f550ed509a8a1a4161a9e766e4228f89d493c794ba7f5049eecb4936fde7
z15d14b807a63e3694425111cae60400b5c9debbbe4532952a0a3c6cb2a4eb833f3d9e63877e11e
z6d75de4022550fb89d15e10d4db0cae7ae4f719ead29bfe597287053891febadd8521803276fe0
zea4386a8cffc4f7a6edf70526200dc341dcd7ae4358603686973551b0f47bbc18d13a7b9a113b5
z46369db1f81b0042106f6219ac6785f694f7b7804d0fc932925418ed9320b5dd2ce61f64ce8b8a
z0709835be08054f5dddbfa04e2d470e08735b97ef2c029095ab7e0202c9115e7af447e819a387a
z039a6f4cd7ad5629fe0b8d84bf9b4b631c919052b461343ccbc583783431ff7eaee86d436203cd
z4b9592a0b06fda1230018cc9226fa21f3b4758320b8934fca347be31b6e2f4fba7d0241ab0be01
z3fcabbddff6f1ee0299e22b58a75ccabc854dc305c8af8fec9d80e256c662179a8335dfa2db65d
z8e618b56dc1c0ad6979b14d1674aff6a8438ba2b502c3e82d967856b94cb1272f7b6afd47823fd
z9db187c3479bad29b8c2c4cb89de3b0437f11cd8757ba6b501b48f63d95528849e289d267fcddb
z23cbf08d43136546b6e8e600a3be6444ca04d84d6f9421bc786b05dc96381698a0b9ea1440707e
z510d0a21c7de48032e6495e70da464107dc5ca5440b7065205b9d89a765a6dd96452f750e51dc8
z170500a76e0034fe54769a8641218d0decb9d8e33125e3d0e558f846dbef070669b753a14ff0dd
z6ae101db5cdbc45220520bd58032d7422703eeb15f6f4099e5c9d766809781473421d4ead5ef1d
z7a8cf08919676916d031e6b8daed3a0ece2080440f71dacb2ffca011347381b8fd5d66bcac1a1d
zb01474d9e18aa7a74a174789b41bab457d55a59133f78bd0433997209e967e5e1e04c2c50f95c1
z0398ff666f6841435007de800bcc76c84b62ea792d8e2a2196fc1c9ba3d12c7dc25b4c58654081
zaad25a7afe57f0b20f95fa2ba40bcfb3fc318911b3c36a66d2555042320cd8ee59eb09c657c2fb
z31bae7239a75ef5512c517ff20dfbddf2e77efdbcb7852765634948ba01a8e8a64f55a1527e264
zc458d42db51330dcfcd24fe3f0d5994baf5c23c80f6e84ad5a2ec2b1ddcfc39ae3e11e05ec0052
z65dbd8522b3fde6b33018fc6e6c520c35ae010813c12d90e235173765e6e9c29756b893bc142c3
z32d1e7ac567b711b6e6699ecb2ae71c790707598402a4bb654ca4131583dfd1bdc6c98443fe4c7
zeab7b94267515cca7e6a32f96a329a91e48ae73604a969df1ff9bb67677835fe7648083c72ba2a
z1d0bb38d27c5c57c579a79b5979b60e86cca789618091639273dcb40978a3716ec0f881ed47524
zb6e81947fe40c371e120aba69532fcb7b6bd775ad3c3b3f15fb78ca748d61cb9a698a1bee505f8
zb5e2cbdd98663fc29e7fc84cd8261755fbfab756c70268cf5170a78ae26c872f77461edd70a630
z865f4c67b874fc677f222a61bb477bf7256a8674b9100b2c63ffd2b05fd8d7ddf6e34f2b6fc977
z7b901cf4c3470947e087fe783d094834a7b9f89b1cfd628b91f5ae6822fe1c8e13645068543956
z279f75d6309ea0c02c77329569a580d1eea454f03f4a74f1eebc59378553f82f3d4f1316788e2b
za4f9413b7f3d2581def6733cf975c1023fa733f4757dd04cdd7f2701ed46d7fdcbfaf1fb71cbd0
z7ebeb978a91edf308c5a9f9ecb1021a07f1a7ddd65b6b6bc1dc8ce7cadb39e19ac85276df70a91
z7431135a8b7c8a029a2e429157551a6162b97a12cb58b0acbc35c5cc8622203c941893f3f72abb
z3e928c91a78fea1198a3f0ffb2f4e5de66cf7c74314981203551945e97d08c3676c49268269a24
zd6d7d35ec7624350fad07007ab9454a6bbae5775a19fc2c3436bc4b27cf0779ce97d321cf2e658
zbac09fc40553399289b03333a2ec3544112a905f90ab3729a30a8812844f26381a1d2dba2642c3
zf504fb6744d1f710d4417a7410d626a053a349ed021064ca9cb06cce307f0d626be69e3ade59f1
z65191b253fa88fe7d6922dcabe10fe257e46b54ef616dc3750e383c222ff43477368c9548a1652
z4666b4e66a685ff52e3da4b74ad205de9aef02cf454d8779fcc958862663eaa42beeae22eb6290
zf87b2f5b0a1cc5ebd592ac7eb98fed42af575391e7594e0be39f7e20556d162b3e4ff16b493055
zceae4be1961aac7ec559c46331277c13c916e294b1d196780faeafceaf390c6ce2e0a8f1f627dc
zadaac1fe0c68d0762f7b8185e9b7d4c5e1530576ebb0be8f8002e7af82d580a77ad282ccfaba09
z7ed45ed8bd5d8f059a40c1c4edbf64241d280fdf6ff2e5af2497139f5c6bbb45a1a144ce17c1c8
z33ff5c877e657c375311a1508afc1d86d160af924fe30e1146ed9dcb7642b8e699252ea389e89b
zc83549730a6ea5c770113f2117b17151bfcb57e62aecb4f5975bc5676907a565f48d9e8fc631b0
zff986e97ca2ee617599d236d55f855ad64da4187d805467a1465b3a2bb3f6c5caea3609762dcdd
z4616db367a55fb3b71cda4cb5f2558073a9f21bce055f48b6e805b1203a6f1ca14d7a6ac48a48b
z9f72f949bd3b0b5ee262c0a1a20fe49ca8c969b7959945198fa6fa80ff921bcefa2b5bd127a0d7
z1c1f4e97c6d5d96f6017cfc8fe77f8dc52de1012e1cdbc5a4e9631fc1003017ba9304a741e89e7
zc19d89763a44d0f9a59686a3fc50c1274d3e012a7302cd8f2b7a17ab126a6643ae256ce3535275
za63157e0613a102fd58d7d7f794e289a966d4f30888d84fe3af1ea8cab21587b7f9c7a448f8c6d
zae42bb53bb38a7aabe1436af720f50fe24e95dde738cb0dab39dc5b2e266fd4a1c80cb23c82bb6
z018800fb5f973771e877aa6970a7f460abb96c291b1122b8b5a7e606fd97a63ec022752629db9a
zfc5635fbf58ddeb6dbf9887751d3fe3113adee7c547fa411f2e87272b1af659652f4bc51d83a9e
z51502c8d59dadef0791500d327e2a8a311ff4d9f5ecfc37affb8759fa773e1cb07a540f38e1325
zbf9a8b83a4436dfd72d98a774ed18092ff005a996dd672ebaca79beed9c50630fff7e5a7512f11
za4f92cba5d78db91feb93e74f9d77619083201d634fa7929986fcad01d32e27c5ea11cacb6ebfc
zf0883f63343ab710b70f35404df58e40e25cccfe268b1e49be4ad1c9758a1d4bc6c11449ab4106
z5aa1579d7c84c3cc904cef99118dd990fd06277a6bcad3c57ccb8ece6a432c889d6af63760e50d
z8df4c64e0869eca3341629f999e90e97582f272a04eaf1aeba0808731747a11246417ebc9e25c2
z42bb130af83569580148e5002b2c0c6487c95b5a757b6d55d4e0eb03a31e25e5e29872dad1c790
z9932541152260893f70810885830e999c1992ef6cabd169670ff67ca5e03135bb31742b887423c
zf90eebb548ee93da88325b816a0225186c2acfe563bb472adaf63530991d6cc54be63b6112bb8b
z15d647ad95ecbb28f6c2409fe749df8c4e169091224de4e9330e68431ea8932dbacd9bf554eb29
z22941728aa80bc9b3e291ff32bbc1b81ac383b26c69cfad4bdc812d161ee55b6dbef5c1b3c41cf
z1a65dd7eecf2ebecd5c1e718eefff7107e51d04405757ce813c102702293383ddab0aa9a2250aa
z0399ed1907de2099e72345a0e091b12f975f4ae48966128778ddea6c3425f217326a5e74673f9e
z05f5ac4dc314650ee33ace1f0353ad68252b4d2239eebb40d9712bbfab2d45633cee7326f70b44
z75ee7f113eceb498feba51064e83f21aa7904bd0d2aa620f95e86b831e96ea1c39b880db866511
za35349928539f7c01ce7fdad613e9988314b6115f7271642fea3f198afde662290e1acad46c18e
z4921072816b0549ac41f9bc71670ef3a2675a7d1822af57d8362a395d5f6cc81617e1960999cdf
z96d2ac4a8af137fb55574043b811a2fff648f3dab58efeefabc0db5af68ad9cc48cd24ae119c05
zc0e5dd8ac60995bb16c4c075b7e11304103b955f0b8c5dac7e5dc219bf1c13917a61f20720b6d5
zb84943dd00e27d0d8c208114026b02ae483888df526bf48e5cb10ce797650138c8f4ea71d40da0
z22adf675cb3ca61697a460f22a934bb758836409f7f233895fe0e9730defb558d9f895e51621d1
z7810ce701bde536be2a8be7173514b3957658c4ef7b6301c68a3f1c3055f1017beb275ed2ecf01
ze5f4906ef6411fd45414f3566de8ec0e9f2254d5b37a1319066b400959f013644ba8ba88308d33
z323a58f6515ed012bde08fa715e25b14efb5dd22e8c9d7ef49d9f52912f61fe35d6c1933ced709
zb5e7bf506b4f5f87a97f05c97c234aca0f82efca6e168ddcc7bd80dc0706d772e9c538a17ee72a
za03c5b1a43ad16138a8d86dd15dd06e4e4b389cbd53f884052caaf35cada4e36557eade4fa0586
z51878890bd4a187505ecbb318f013134184eff31f16461e1e303fa255babc191ba27cd26872b04
z5ce8be1ef190a4ecd15aef01038ee1e2c7f008e504023ede3afa4d2df5862a33d512ee3c9fb164
z548ba79ad39145b1fe1153f309e0c6866c28f3a8c2ff7320d9a323e7e22f5778fec2ede27f167b
z6de59aef436f23a608c64e2005fa8219fa0da7f138ad69768f9f68037cfa46eecd58d619ee42a9
z538c9fd29f5534ae1b8add04e5efbe39edd701c93e846fbf4b89a964c42f35ab406b9cc860de57
ze920244f7a28515c618de9658589fcc9477d63ac2cde214a3803bf650956f4423a223f7a0d8ccf
z365577b8edef5c90e78f8aef5647b12f5f20aa7647c11a4a33b5f658aebd036fbb3274418099d7
z0cb7e2274b15abbedd56790dd9bbaacd07b3cdd138eed86dbc79e129e0859d5e447222db37f3fe
zbb34576068c95f069998e62054161e31d07f03dadc831f6e73489717141bafc12501239563b0ee
z41300bda66a7445483b5bdbe0329ff637c8895524d404074f457348706c57948937bd058400210
z525d14cda0bdb8c80c86d5ce196c4f099b12b87a3032b6b0212ae1a33f2c361a8d08e9b9442842
zab05578929292636385625ac33708d57f0e81eb0c7c3cefdebd38481e08655f47d4b0b3ba88869
zb3046b029a304af0b146db0fe3bb6eeb2b8ecfbd4deb5439832b23bfdbd923846090f96ddc3452
z8a777e057af2cbb0faa0a16b124fd79c5796bd831a133975eedd20537c3bbcb9d7da1290ee189a
z59728190928456826945839dfea252d852b414358149f8de5594362b875e5a8642badda6db273c
zf5f474e43d8fb846c3b4f2efd1e4e51f6c96dd9ac1f385e6c29863ad6b3f73c2aa31998009d7ab
zb67eaba95fbcdab01b8ea3898321419aefeaf6560d8bc7be74d11b182e425925863cb9271970ca
z9d384de55316ca585294edefecf0d362d83a6e034c73190c8df53640994f572a6b905c255946a8
zc722359c39e90d3c0cac816db0f2e76192d5ddcc3f0ce6ac00e01f1b59512b4d1ba688a7a6f4fb
z5ae3d90daf7bfb99de7b92d7975227b7d18a528029afc30e3a604de660b02e51541054f72b418c
z94910510ee82f3f430b89f79f551745943737963333c0c46c6e369fba75ac096901b29d419d8b9
z8b8a1abf516b81763a91a0964978d7a3c4464713371bcc5adebf10327934157b77bdb8f5503838
zad87761dbe4b9b27a783af5eda3945b0552f51aa151674801e3dfee5d2cc9d8329691808136451
zaed87b3d6904f8a759c20745d23a00e096efd1608f7fac75a724667fa86786e1845193da70ab02
z1de0c07a52e8b52f90b656311759f8970f2f4fd49f051e5898f6180d86aac5aad7bab0d20c9933
zccd543601a985f2836f45a4f268c7aaa429cad833cf39868efe196a026f6aaab71d2e723758d26
z0e3484b97f6c87f0a064321705bb8ab3c6066b65ad79e2a1547051a2545998c747fc4de983ab79
z3af92f158bbaa3d81d1cf7ca4d3ba9ef3cf354f2fef56d778c4810fdbfa7523d60b8c43df25ec4
z8a89cba771ca005c520245d5647870f7cc9480b5df3ae8c239633a5ea8ef1e53ee3530de4f5e93
z2d306e2927310d3940c21ea7a1911f841a267e68a280aa4b99dfc9010ea3b826debf24e9d5d931
z035f4c76860e4263694dc1de5e9be4e32734adfaedc08f3b1d0a044975b0a6a07b8cd5465688a6
zbc4bfe6e27f848b8d4952821b901c1d781431a622000ea4e871367107d71d77ad71f6fd6b8d284
z63253d9f692c80263ed68cb5dc52fc836d837082f619e1ab63130a382db5e828fa4634c2fb5233
z4716eae35a5b6b301449ab250e17a19d09faa8ab47b99b46a7fa67caa04d239c88c2634e9f26ac
z75bc444229c1012d9e66678831da9c90170255ef5e3cb609a9a67897df696d7860c208d0dca992
z3c3e4a5e18119854c49eba08ebc1fed72d7cd5dd2bf2670e054a66d762305e9990b5c3aabb22d7
z7b04fe973276a050c17455a378d248d77000df1901c5638a1ed37cbcafb499de87ba51e2be366a
z94f1457112856525e8bc8dce7c8ee44ad6e6b1378d70a553afccc9b12b98a6c3dcdc5b88736794
z033f384095130cd6acbb9f91c440419cb50f0122253158d6c9b7d018d2c1059624fcfb673ff030
z9beee0d92f721fb75ce9a37d9edf5000a8de9c712519cd6c3e16c538ca28bf42677771c096b05d
z8339973c26356fa5591530fec1728820e4d50e9fcfb2142da78aaa80219d523748dfcc5e5b7724
z859747d7a0dd3deea4d7414395cf24621f1ae80f88f2f62d6681a583c35a0dd098fb88fcd4afa3
z1a39b94cb8808daf5656688b4111d1403bcf27e21fa845d1f000c2c58132b4ce55f6b5f7706db9
z127b105e52484c20f53c9794864f2633572ea373fbdc81586021a562dbebc3673743e348c14d30
z9c26bf0bf62e1bb32cf02db88f11f536852417b2231252e668edc4a6474b24e2a860bdd08b447a
z4fe99ed411feeed24c07c8e15b48f00ced9ea42a1b7461aa2c314a72f98aa7bf1a38a1a70914bd
zf6945ed4a925b0c9dc7a81d691deccaf8beaf3e0b76f6b78d3abbabeabd530e2459d8383337761
ze5547b7a955d6b0557eb40e15ab833bb6225cdb38bcad2f77471ed8164f92e2743f11ed0d6cd05
z14d2140a0c8b9dd1d83b320a6d6698cbb9be5236a122b71d2d98d4f0ba813cf4e2d5f268947708
z1d0fe3f93d2e5ab6a5a567644fa99f500878ab620ad0e92cd6bce8c57bc384fbc0182d011eb0d5
z7feae5841b1639d7ebac563defd53a098399492d206dd5d230ce4dd2fb58d327f7a61b3c8e48d6
z0e7030452505bac3587fdb3e990fb0ef24d9626af521838b4ec3a37149e7e59991eff0556c839d
z0202118616fa4730e0e8faae8e16af2f50432dfb4d1fb5de815df0f04928d13fe778f9c5eb6f5e
zc61c710e81791967e38ba5c9babeec04a983ae4cb654c140af75f1858b83bafd7357bef451c968
z7df91d54cc9d12b0f9bd2dd61c41f97fad45bb5e9066547352b260a099b823c14f7876ff789e71
z048863dae35fbafdbe8d6f89fb6d378504ec1cc980fbe6adc5f0c147cba38ae4004bdbf851f24b
zd6e00b0ddfbfa8bad7addcd3c55091803cc0a3fdbf53e2cfa8d6276bd3ab0ed2a1a8b80eb4a89d
z8693633a4691ae024d231bf7a8196c97e151c35e6f38b7f34fd0365e2ecd85f6e671cf74e3c43e
z0bf4d8cd9919a1d1fbe03e0f7d818c8c73a290f22d3a18d065664cdb415ce5cd30dd7960fb71d1
z68a6a4a1287fe976623c24d4e2e27ddc9b1166b85746136c823f81b6aeb9fd42a661b93b43cda7
zf13ab1140f7f298196c14a9464a4a984ad9cece0e8dc2b8f65ceec43c4faddb0a627409e25a93f
z821ed43eebb5dbd8988f1f0bce1534a9094d10f94dc012dccce5c2e14d69ab6461629f145f1a35
zca9616c298775bb06591b0242c2223177604ee0b2183925fd419553a706a16e60363a710304e01
zb980516a5d58ac6435e50c07458f9c19f183422ae2683cca62787ba7ed2af75f650d915c2bc258
z718eeba4bec159fa2c260afa8f855e05d8fc2393ff6a104e6754b268ed3c2b624ee5cf2f1fcb3c
zbbcc55410d02b1579dcb4e3be550f431b81869eab52458f19add2828af00b36e45ea93dc45e899
zf9c90de0edc11c9329e9b457c07556123243987b7438994545b3d15af0a3b47102950360c9e1bf
z78c6bcbdeff15d864d6343c2d256ee74660fe9a471797dc14a537b00d32be42bdd45ed6b0ef654
zce00e24bbd897ffae84df540b0f038354d2fed6683b5357922ba3ab45b4e86cfdcbeb2adb84936
zf645802af384e17868fe66add6b270a6f269bac9e02b334ac6ea7be44e0a1cae4ec80fd924adfc
zac851c31020e11c02bdd90ddc7bcfabecbfa43eaa9d0e7ea6f159cf0aa11fdb74c6f888acb5867
z8de1887a8fa07f108d43ca71fe9cc3ac6b6fd7a43e39addb935385071d9b314111376d91e51cc7
ze3cd844265963157ca25801be99d52f625bd03faad29b6457688fe1ef5dbb86ddb5524dab42a1a
z551386a904512ccfab6a52936cc040aca196977cf5a749cfca0bdb57c395b18a60dbfd273dab69
zdf8663f4732bc2be5117304b0ad37aa96208acf0f3388eeeb40a1d98a8c661fcc9b04437f5a50c
z9f166cdb40e5ac868ec62df3d86a2e929f8593a41ee1b7710d00d8b28248b491f146ad8df18c7e
zf25f8065456edd331127df30137f812fc510cde87a4f3c833ac42a4864fe1cf4d87571d1e79b37
zf2fc6922f259103b2074774a6fcb0242842f52b657f141f469ee5f297f9d750b555692371987b9
z98faf98a45c2acf7bea5cf8609ddd7f121a387850082ed800ad1f9621e3239921aecbc8cce8697
z63df8f3c3b83b0d16396cae6fc9a9b9579fa4537b59c50ffae34de933994a3adc0f466ce5df652
zcfad5209853f2a7d6b9725fb9419a948f6d7ce9012f21ba50d646a64b1fedc26c8692a99288abc
ze1c906c5b5be40e1cb4a85a34d4a6a02aae3ff1b05e1999c5d78801ae717d1cc88d5f5f1d0c52a
z222fa2f644cc16fc028745b5f8cfabeffd98d62d9bd90d8e8002b816686247e1eca3a0b796a08e
z8ac6ddeec19832f54964037c658187096a8805d2afd8f94ea3ad99929d16e9bc2b9646bf780d54
z68e375c598864f7bf49bf00284cdb905f1c743a55b48415b0e0d01fecaf3482844359dd33161e4
z8c095c1e78c2547830ae0e064637f2bd230ecaf90b55d718266cc8e0377cf7f879443c19c5b544
z11cb3c30eeffe29375beb7c5d7cd643462ae166b983620f54236afb471a2d98841b184fb32980f
z0f9a9557009e38c087ab291f5a764051d3b6eee9637b2e85a30421ef0217daceaf9d5cf5b8ba5e
z325761e2e35ca7af91d1a31748d20f6ec4152246b8ebc773dd087f653cc386baa8a42db701b635
zcddd04d38ab4a3f9d4ae12c345ed4d582aec5c7f053adcaa9c2f2564534a50d2360543c53c66e2
z5c19916a146c0bb1d4574fbe588f7796a1442fc92ca23a1fdbf337fdf2920a77a0b7d18dc1de1a
z782324a948cff4b13edc07c761411e7e7b91fa153ee83246c038608556a84e9e28c6a6970cdcfe
z23c0c7181761453c318e00f92d84adf6e09f76ace37dc517f1d708dfd0a2b1662261d7821073e0
zac05c31caa05703c1947915bc7f0559eda800d3fdcc4d55f9d5a6b0ab4808a93c3099bb2242b61
ze2876142e54f02b32221aeca15bd46b62e0e0934c171e376116ad180395ef40c657fb4dba39615
zcb66a88e7cd33978eeb3f1fc25bb1ded42c0ae86ea20529e4ab465b360bdfd99b26191524f9018
zefca60e15188a9412ba8d118626d1e8081ab593ff33ec473451419e3ddbdfacf9a88da9d287562
z51ab469a8ee24ee90441de09f2dec38953584b6d71356e51941ca5d9d776560cc0ef5d211e376b
za6c5fb55fada2c75ce3cd4a44562ce37e90045e746225c11fbc6b97dca97dee87ad4592e9b8db3
z1b0313e9a917d6b99e8956d56e32c8e679865905ab7254e7bfc67b5b9a8b550c7f4cdff4eff01c
zab3fded7d540d80145293eb24a8737014d6c4d6ac9cab133df7bbccb363c03987f19f3ea8319dc
ze4c17dc3ffdbaffadbb97e07ed08963d0bb3287f9cd3b9b1d8e52666d6f4018a812251d5248cbc
z3df4219f119a207a55d9635a7ae2804213a4b800e40a0425c18c106e7db982b01fd3fc26cefc32
zb76c1628aad68f9d4711786f30b80649c6c6d125082d9e72f017bc416c02e18c8222f2a66c73d7
z1d12634518d3b3288dc286a8757da40c7342ec8e1e51e09a8f34f14edc353621d69b3a7eecdd45
z048f9e3a3b06f843f28563fd391a9c465f663c3c30565c625c8122bf2565ea111dd80bea070de8
z11e1790cba63cc32f4b0f221083e37b165ad0fc4852ef7923dfcdabf11bdba0d9b69906a006fd0
z941b7d806a87c3d6fa4028f52b560772c60de016aa78f36868fbf74bfdef132f7edb96b1b552d3
z03b9436c0fd82022d7dbb216a88c414a83fd42313cfcd058aaacd9fba64682e6cb300c5823d38e
zf5f342bd4b548c7de6fde47628ce4d8d036cefde001365af3d156363d4c2dfa8fa56df9ed69579
z0f7f19bf051c9f21436dd46281181a76c3b071b413eee949c285a4c65fc367c86b62675a187eaf
z17141238b29d77b49ff831de3b848f79ff20aeb26d99bb1c6cc3f1c810b86ca4f8569d4a06ddf0
z0deea7821e8edad50e589763a242ce52b48593e2ff1e53134e2b7c51ff76d6277ad722ad8a3586
zd1048db8225a48b51b17bc83829d03c4840a27b0916ecead0df007b9ae5f5c7c290df819175426
zab53bc95f5fb96609157c2cc6280b1c293273aca7b9d6d40079d83a3f301d0f0c0b4021fce09c3
z803d9e9ad28afc347f977a41c0ca0cc607dc6f301e7a99c2d34651411587b5841fcef13721972b
zd596eb1a1209ebd15dadc715f1e487fe175382de324385d00d26c0accd45438e6fd6190528e61e
z00306535c8fb979e10c23df835906d7ad78c5675c3008b70a688df4519aaddc08455aed611df3b
zf08e46b3b2f4aac5c8290442a44ae6bdf150802954a3fdc69ea6f475644f478e08056e80817a93
za253cd3beea85cb379a5619869184a7ba858b62e839ed25785e0870279ab6df7b119bf166c424e
z026855f2c9d668f080f3a90bbe54977a90274f8123a0a93671b23f47dde52411cfb4f1407ee9c7
z4df40a3f41c3650cf1e16d7a0516e53a593cdeb3a59b87b72997f72d1a8e05a8d4b54de1ada800
z706cda23b113038dd1376d700d72db2459f20542ec60c577eea0de37b6e0adaf696ede6b496608
z1406852984b5da33046851997dd158ac254e8591dc600f8b7d1d957310d0c9a984f92004437a6d
z484a9473e8f8f2a8543befab6aa9a66445ee000f52ff28d7bae6b16d12da273337e059bec22259
z132eb771882ce8345402bb2862c3f4414b71382eea95367154037f36f3e7a773b33434a12204de
ze0e19c272261af33e224695f4ff338e0f8d848cc7df75f59e68068859de2d9b117981d81850952
zb9979e78a711181139863527e03eb9cadcacadced23d0e89a44ca1ec98b45df1b68f630dfb0797
z55986553559697e95cb70965b782a546522fefba8063e5e4181b5209c3bae49e4f71bd3026ce7c
z422929a40e6162939b685a921b899d825896d6d30c9e76d01e13fd018d6d2a728aebcf1b6c03a4
zd1346e060f76a68e3ef171ed2f65fe0af85d852f101386849e5638eb1238ee8bb0766b1dd2bb99
z24bd19860942acead4128749c3bd777d2301bd90851d5ebb3e944f768245e06d3ca0df61d22e3f
zb0ee2f48bf4bb72422a59c5ea8824c616979cb394646804ae076c67a513b406aadeb8206b20f1d
z5518f02f99da84d5e601f92fca3a176db2359a35406b7c8e629b60428e4ee425ec53c2fd240581
z78d35d3af98f2747f9982716dbcd381371f4e455174ba3901dacffd837c0cf08920f3bd2e1752e
z030ec678ac7cba48d5e14925815b99d6b65b42d72c552d77453ec247ea12591b6b51bbb9a04c65
zf63def0eee1a6ebb6eccbc5337afb4b23f7ae54f48e31fe214addbac7eabe4804450e6b7c076e8
zd1af619550d7be73067e7670bd0cbc1f6f58c19f5c961811e5c822a91b939b80c208abfad1dd80
z93c5b5609fb126fab698ec0ad8859091dd36d32f710aa8301cba3b16f779c2f17af71a1ed7fec1
zf1179a81543077960c145b13bc8c12b2a258b996c5a709d03b88ff957ecfd41935cd480e880a0c
zd67fd4650c07e4140fd8dca567fde6f1a2ed123a75de196e6d714d03c075b47633a67dc4eb722d
zbe84a068526d1aaf78ab8667c383c79d476a751a3ad12342a0905dda12d885cc2e2a8923510eb4
z71f171fe261d04f9e0936652d5af520ff12e184a1a1cfe8c20a6d6dbe75dda19580513d3360943
zcfc0b5f5c467a6b78200bdb4d3c143ffb907ed78ceeadd3ce4c03a1e20638bb8e00aec10b1acb0
zeb8d24465d114f6818e30e2c0115f42e85ec816097dfae418879fdd82811edcbaf7d58ae09ff95
z3bee25dc202b0dfdf3f36946cc6f8dd59c3de8d0c29b1ba0435b4df301a5a3c19e696a1d25a5b7
ze6664a3f7e3ab0682303c3acc76e3f8321e147515ccb72fec8589c9018957963a252595420fbeb
z54778f430ae3e65cc4c6b92e8f9e4d44c9a78bfba613e106fd18d1df199f618f729bfb485acb77
z95a100a21efe173eb878be7a5ae5e3a1c23f912a2b62fff28ece32914eab10918a5cc2c438c431
zce7740fde840c0d3d8fe63082487cd47d2ebe9012a1a88ffeb9583be1b4a42363da83aa414a998
z6230606a5e517e3a9d296961907be39d42312dac24543cbe09f1c917ba8a56fb43d37486a49dbb
z109e91600f8a3b885ce7cf794231a26790d8315baf570039fc1b141e97c4810ecd676affcd9211
ze959faead912c58414a0d43fccf05d8afaa98164dde3f7fbb516e91df55ccbda4d605c8e4df830
z893a0c639bafe9c720b16419ffa8874ebcbd06a500fac03e334cf383b5a2b92e832192f71f8f6d
ze43aa4c17c2a36a4cf4dec22242cc016ded9af3066cfa955d9ba9424740ba5899aa8227c901e3b
z57e933393ce7cd0534302c63ea170f720ea1f4ee39cc0073daaf4c420971560ff1b32c927589e7
z6459e18672dec315779e38fc34bddee59d9542fca51a26d4fa5797070c0be8f9d5539a916ab912
zbd8dd2d78d39acb5d70e0c05d1b204b5410dc9bed42b8221a9a486a53b4d12f9b28ccdbc958d2c
z9bfc6af566102a12a8a6af36891dc5db554a9ff6d797229ba85d1612c41f3ced36b1a772e5cf06
zf288b4a00eed6750c4b2f21f7e181f09f923551eff40b93163c1c9b9f5c352d35098b8942fcc27
zb2db0678b3f3d2303aff44b6a5f94711603bceb97feea319c27414017257a71c6a5f5073b4e783
z82cf942064ce6baa717409684540ee53044b04b06fc135f5024044ff7a8e47a00fc05a7ffc992f
zabcca4a17df19853edaad49ea313eca9d94a68a07fc7e79e3f825990e90d3ded2f0bf41ee4fced
z82b823fade5dbfa4e0ce190d252a2c64e9d30cfdfd5933754b848d6f402fd0c79251e46621167d
z1f0c6a7d83664c4cdbc464cf5753dccf6f2a41451cd08d0594272126f4f66ae2f06d699083c370
zbd9aea48e304930f05eafd6fab98e81ff7689bba6fb48255dc93417f94936580491db9b22d36f6
zbb3b70da54b71bd509481c49c8ff28144c2b44a87b9c7f5abfe97c1b0a76a9771edd9f6e56698e
z9528814491b6b99b53b489f16a37c88c0030e680a64bbcc699ce0072427df855007022457cf57e
z43bccc45c60cbc127f200e0ddf567714dbd8aad36e7ceb03d99183920923c560509ae623f264fc
zbd2170e8b6228ce4c2ddd816990b20af2cf4a7bdbc1ee5c8692ed9728308f50be912feb75cc9d6
zfe6c56c6e94d4a82cd1d809b4db0857567d899e40181d353c5af1ed072e56ece3d00c4bcdcda88
z5116a9019621ff7b0d57c7719fe8416331a1a09c77cbce06dadbce03077fe9c3c61f90e592f2bf
zd47fdea302fb5a8fe70b471891ed56a91d45fc8e2f2cb72872940b4b1a05e535a99e537e380c0d
z29e31715caae386c3a139bd6b4fb6303ee1232f36ad20b27e32b6cad195e3c34bd2480e82bea22
z8c86131721f204fa15dabcdc8937f321998ac19aca2ae67967d045e0222dfbddb2696ee07f87e7
z795b22814e7fa90d19e1abc9e5bf264012f15af874597f65de2a421e32989eb61b3d07c0bd0269
zfdf576407c25fbdff3367b948e284f326218d24ef5de150eb61a130a99b4bba1a4e8a43770b7c9
z815578bd4da060e5e8da73f56180147767ec6dd797fae47895a10da65d4f30e0b0ab9c3bb2c924
za43c4ed93a76b71f96a995074ee29566103ec8a75871b2c9610269044c1f0be5716587a0cf35b2
zde86c12bf8cdd33bae3e3822b062a4754a605635a0b94594ecffad79601ad494e41de4f5817c6e
z22c5c0b69c35cd8961396556d9456a0866a210169b989f8e242f17c276a8dc82915e26f4f3d160
ze384d0744de1092ee6535d69c08d16e0c6ebd768878a9b2cfee212d3ae5dfa5737c603f17b724f
z6e871cb694713f15c7d4056ed7b0335e9b00ebc07f587b27a033d305b111657b8c45c31249b03c
zf46c50aba921284a7066b32a1c47b5ebbb9d4f030244eb9c96818f28676482e428c55a70bf9341
z4a2e0d0c45228f72f22220649af8d2af6c2bfd5e42aa164a186eec3598b54aed60b71dd3c890b7
z12428eaf5d1ccd7fa3e2d5e82fe6febd7cbb8ff31ef17966955d3944ca99050eccd0cbb69f2aa7
zccdad9b7702b2e2623781fd8430006a8bcad3c2f21886026f29d8a200541591b5c653cf25d5bf5
zab6b865bd30620593e4b3e60d5502c3f3c0d9be8c6a18d4ed26d2abd8336312efe3f6caa7794c7
z5c41c1bfa9b95bfd4d2d36fd919a42c53a07ce20186f6342758170c48fdd2e4dffbf308fcde6a6
z8c05a36f7779c03f0459d04a0f6365aa0cdce7af027ff056565f9be696a22ff174a236eae20800
z53ddd850e8fbbbbf30f041ccd94cc82148b35772abd7caad511be738f4bd1a4d1c2c794dec7086
zb919d3a14eec1b93ae0de86f451f157a875da8ee78610145b5f97ffb1a00fd931dcacd61bb41ca
z94043805d69b6fa8f8d62da69ed54bc52252eab030030c4d323c8c466762916a5a99c6f370f798
z0f3803d2c15b84added08191bae3f25f555694ad4b26758f0cc644a48021d59a048e00bcbe6119
zd0f4288dc720cfad62eb29ea179fd5d0c2e9f231d1d3a901917a13f7f15155b210d5a25f39c770
z0d97d47c4da2a1afe769282c69bf4c61c198b2f05ad2f73845e41ce0409b46c18c6b1b50bd732f
z8fd63704c7d77fff3a218ec369456cb8c7c93b6ba330ab02dcf7cd475e5e84f9299afdb923cbb8
z27e720f79b8d40d3e1720d05191e153f70128e35637eb783ee8ad006948ece4c7e34bb3dee0039
z362600ef2e2b156ef4c4056a620805ad9b1e27b0e03e03836f7afed25a58bea1605373e872914b
z6ec20672e8a047db0056bec2a47fa2ab0126b4923627136e7bef52c596a3686923fd29eb7c54c9
z5f94b51d5858e1efeb9e356e3cc3276da99bd9ca5238cb8cfb377b5ca8814f2087f186110d17d3
z7e4df80599431e0b7fd89a7b84d2a2aff7168c06ba0c769cb9a4fe3234b427308e2087f23fb929
zfd1b69df0a944f53f0167aea88a04575dcbf7e7c1c2d146945b69c73b21cab2e2deb3e1f70d414
z0de360eb03963aa95b16db75666ee2bd3437bc6bed7a57266ea9d741379c95324fd6a403bfcb5f
z05f59ebb2579589e226a7dc6e9bca6dd7b50bc9f0e4d4ea4a23fd71613f8b6a6ba6fcb1a0a0cf3
zc5168746bc5ecde1a3e8cae031025fe35ba7f0d8963765319f229b49a646b51ed8efa10f5dfa72
za0d142d486a2699d77fe995ef3094958a307efbb2422d5d365f66faa0cc2b800c032064d893a7e
za78b084c0ae6f8addf913a5d70781858a833785162341c2f065460eaa97ba7f288499ee6b4846c
z4cad7b446a14bbe4792bfa693eb236436a729c7ad3692d65a5845929991068885f9e09a6cdd132
z84f53dc3fcc88d60aebfe21825e1abb30cc110a71ce5e8b560e5ef2ba921db7529efac9cfd0bfb
z33f4d0eea3f1e46b0782f5b49305595157d481c2e2cef07d6a684bef7f995d5cb985add6d65a26
z4da3d4270b14039e4361660856cfec0ae557b7d31aa3fb7ef99a94c036fcb761397d116ba040a3
z36b42a72e5f58533c80f65c17eb110bd29c689d161fa1a5505a329dc0a3a9574bd43e1457c1ec5
z1f62d921fddcef4d99bc94b0b9cb32cc0335f2bc49088266901a0ba3b8adb5fc5eadd381a7764d
z99bc8003d125eeaa667e3ea49a99da0d9a45ba9d36d1b189846df768a859682133a52fbe23dd0a
z42a6ed419adf127e82fb51d29fee9982e029f99615717addef01fbff3498095f5f88e5e6ea2358
za4f619cbba4d2a5c30bd4801de2a8ce0582df88d88f49cc1c347af72d6117127a8f0847e302894
za342c8f36508c66df7451c6fb595ade8f441365aff378b2b6e2dd4203e9ff0809d52d6f195994d
z56d2f4967bfc310a813f7436f0f39bdaa7688c4af4c336dc5462495422f8c3b057db934b3219b5
z9983fc2a0cb919c2e29384b70336ba4479ec09aadef42494c0c6593e0b5345353832bffc6f9019
zac09d638aa07286826a175d7e27820c789607bfeaea097d00dc48f3e4c0461fb8a2b3f7181e236
z239c387d8dfbe60ad14e0a89599f43332a4c4f62fdbed2a36cec04d2246544119bfc5d8d56cb97
z7758f2313b9ee472451fd2ae89b50c7a019b9ed883921bfb0b2e478c69f793ee5883922cabed20
zb882054ba55b148e040cdf24908c5c52f237f62b414b4d4fae17b90918ec27e7c7347908d6d18d
z81cc90dc310e0c534b1a9aa3297b34fcd8bf3bf50e7c0e16426f2e3ea40427c3a0e61dd562687d
z07c9a23e0b349e8f4d9cf02fc8bcbb505388ba7a62e326effbfd983bbfa1d24d26b882686164c9
zd7cd0ed613c44caca73d16e9cb730f8251d4f3f8a811a82c45dd01c4134889ec2e25d5d7861456
z088c71a190234ae1cfcef02902a22ffd8874a019c42a26e6b571162fb0d88ed177f79300242343
z53a51db6d1b3cb3acc07d0cc92c241ddc9f4390dd3209b8027569c02209fad55d045b6548fea01
zf297be1ea277ea5436f371869868f9d2d094cf7b3feba30282d3b3f1bbf66e377d36c0e7491de9
zb2f396226ee7705cf8ec7e2077b771ff00f00ac6610d8a6440fefa2ec8df39177f767f996ceb42
z62fbc20b9bd6c4ce093867d1f8346c2983905d5855da11241a25b8d5ebeace3bd9cbfa074b8706
zf8fdeae256f9c3ab4be80c6e6d50e270fba724d393d53c06ee11188f6eb492a985595620d53964
z69afbb0ebf2e4979e54028c7ca89e4251b5fc493500844d0228f067ccef2f5872bce0eb587cb8f
z66a38b9bdc67f704e813090b5251e62a7436cfb2914efa33d0daf0ac0e1d9575e14f8b2b2728f1
z7e56dac9ca348a12365b846ee4ee2c48dc128c50b80fff57bfe2d565badf4dc664347dd067f397
z0329970a669b6666611fde0166833a1ffc1335afb5f33c153d923d60381892552418d841bce873
zb5095966bf5c7931ccdb81428b9e1396fb965e9a0c1dee1ad037ec6c3799b7c680fbeac4750c63
zbc7b65ceedadc4d61a0ee0b3b65dabda95e3b9539563c65276e54be1c457086217cc32c7d91af4
z7f202ff3b3e91d8334a628830774552bc7ae04f8d5d79a3fdbe004f7fab884df5de542189bff19
z317548db6094d053763e03c6f4ffa4081bcbf067e83793ee79765fd57bf9de9ddf03a0ccd018b3
zac66a9c66ba24c7506e7687d7d9d0d0dc27f2af5aea347bfe9f0f42ab7b0c1645c0d8e2941fc7c
z32c39bb2cc96b24d6bf08dadcd46e7466bfa8ef362842f7026ac4dc8b8e180714bacfacf0a063f
z1e19ccb7e9e74efc3d223694107ec67003da38c32c9c514194c199bb2eb415cac116e32b3c62d8
z2f59349464e540d0e838a8d8c180aed39e1da73d7a761a9d0ce01dd6b0a4c9702073eb9c866d55
z365af848f246563b2de812c79a7342a64cf97995c4eca06dbe65ee9ff8ce1a4af10d2edb3ff572
z4208d92dec8d329ef05fe45ac8bc0904b7d55a38942b95f0b420923699c5001c7c375c39ac55d3
z015a5701ad8bf0c8e925a6d70e687e10a986427a44f10f44c0d826ba7f5292a8719ee31fd379bc
zbea546be17e1df96b811f2077f2fd96b93c43f17f562d4e9eae5fc292a9fd620700af1021f3abc
zfb11eb0414ccb693fd4c68d2431e5e2a1f16a22ec94dfb8da41c8c06eca3eefe05e3a34b993ed1
z24103f7e1510d86ba4e8bb3abb2ab8ba3a316ea2805bd1f8bb0ad1c39489d8585521e13d8856db
z950f73f69d9e3c7ace539b5fae7983c7ad18fd21290a76ce3448edb163bf37e9d01f9e635b6c08
zaf6775cdf35030cf00ac2a5dc585361e5f714bab709f18314f1d35892fa3e5d6f8463ba76ef898
z3a5def8bd567bd047bbf0d1cba5ff38840e9ed882b41daf3c23e04a4b33863c732ed28bfc4fc71
z6406747cb38d83bd2456b84e41b19ec471147289765784e0bc71800eca3432567b547be200b93e
zdc24e07650182725f7110078980d30886a2bae8a432c5f424923f6211080dc1d3dd5d7763cb132
zbf06546e0e575e9b3f6964799f871da8446282ba0fa2836348436b04ee6690d9014c3830fb84a6
zbcef5b78555968b38b34f52dd4be66fa22a6782a2b7df6ad2e3ebfb530c6f202dce2ad508bac82
zcb2d9b96c1040e8acf29f33f8348bfb22c84485dab5fa342a71a18df130b6e79b53fa7c80e4b89
z598ef531a71376e638a5f89fc2f46d6673d8e8edd3b55f3aaa04c78a38ea4ad4f4434fadf5eee4
z0346dc980c282f46a63e388c7634b60f5d631f5248de670f371d38c422e3c5d26bc12f73f1bd9d
z7d43f33d5c56cb3734a8bcf060049533d5d0db03036b384ce6c304d5e220901e9efb7d82df571a
zf8d47d83118e15782f637f7adacd73658e57e9db63117fcff7c0fe29666cc3c4f0417a036bc196
zb31e65fb6d525b89039836be19a9acda0037a70d13fcbaeec42571ecc9c0eeabd01629ca5b3612
z1d91679244154c6e7159cdaa8ec0fba4630e091604c1bff4354120a69490dbb718f73e25a7033a
z15c2e5b8b8ca8386053c97aa10f4f6ec7217877f59ec39154c2cf78b9ac6d3e9ecff346527c490
zfaf0206de4f02fb287d33877406d92d67edfbeb77c5fa05ca02ac4ba6365766a60bdd040157c8f
zeb18389493c4395c806408f7c9e9fdcc31fca23e05d164de6564ee675ab3b923a2f11b75d3e5b6
zcd5a001a348c552af26aa4c9187c31e919ea940ac8d0c0db3937f8842bbf18b2b9430e62af1b53
zd6322cd7706ee932260d726e60d1b9f28703750502dc4d20005a79117d83db4ef3b297dd1c091d
zebb729a45114a9ffe45485c939437169d947c9279d03cbf536e2c1a6f540df91848ebeaebb03a9
za95290c1e425ce8b54a04fa5b8dbca8dbf98be233adbb5e9a7cae10b095750320ec80ba764c882
z14760dc9174833f2fa38e103fdaba5aab55ae217ad5252dfed8cb1d25959d5f66e517960c0c705
ze286b16d4c4e02722a41f4097f481fb9bf35d4bfa894998a2443dd412e9e0450ec3db545eb44db
zd6c350a98d89adf81669b86c6852025112d95f103205fd89612d0a784e0190f95f0659c5c6058d
za2f0763db5cac73454ad2fd7413b38426dbcf5214ddb8074e328b16906c5074528ba9fc75bec28
zfa2f74a7efb6a0eadeb4c1ac69336232d49b6082b067a8e4b859ee5044088cc7de0a8f27b9b8f2
z6d51631427ed77d30d26c082463ef00f9034977f4e9bc4ba1a6d324bab40138f072eea588d012a
zd962edd5b29601dfb237c059cb20c6029d6cf5a3a1ab40ada22e258c7764a0f9681718b8764e63
zc142d056e861d48a5b2da1afc2a27c9bf46761d78bd02a4b07b9d90e5033f1cb50b9e94a729411
z5e19f60c7ecb033d555de4b60207b52630370b40442998821267eed651fe8d38a2dd02ea2ac638
z0ba17a43de3e45a7e6785c08fa4e2b454fa7c7ac178fb0352c98b113c6b825bec69143344ebc71
z7720a694bf40d78e6efe208b411dbd7327ef3899403723c51ea75d4f22c95d1d8c9f644dc45c83
ze4e23612a282d1f03a2e79218901f6d384defe89eecbb046cbc790e63c298ae2591c4b2a0d439c
z6a1f54953e64139d793c7fa33fc35081e64da9b9532af2887287cd88394550f390a49826c330e4
z2bf5fb7f3ff06463d679989ebe0b5a71d863878b6ad6aa0dccbb6db389d28c48a18210d3d77261
ze341c38d09cb6aaa3a7d9005b6bf71f2dd07d33659eda0b897866adabf8818355e4effe50a3f35
z3e9144af11a3d2d0928acfd483fd2d673fdb1a23ac54b02aeba82440fc36d0e0a8b09a0f707961
z22761f93bcedefab601d309b832ba46270beca9d0dd9802da2f70b03ce2756f7204322116766dd
ze3c6f6175876106334ddba10c332a20bf5e1231a750e89365f0d712a23e1dad19b8a57e95a01fc
zd8ead9b2fd13f1af19fb44496ce31807c9754d819b104e1b1684b27300ef019cee0870f4e8e685
zf3bd6eb24f43665726f90442c1f8f0a435de58b20010765dd48bc8dcc000bfc4b5882ddf2fc1d0
z4652a601b643275a666d259814bf2d8b71776a7e5fda12be5bfe4cdc45232cc41c44fc509a65e0
z451afd7d4d695893f2e2fbd5018ef6007c8d6f1d8f7e8a738bfd50333f2549702adbf11fbda4e1
zb7a53ea8ae47610628eac4f2f4c2b4d2f92be3c5e12c5627811008151709df7a6086a56cfe6969
z4423933eb28aa54bc83c85c2606ba45aa8964c1a4340af7cc7c1c06253f1411233506cce56e808
z66f413e877f45b87d7600ecaf7047edcdb61408988b3f2257c5a588cdd419b311f8998d038d3a2
z5f69b3a6412bdd56b65f4405b75dd979b2764d3351b862a99842931f2037ce2c638eabed38ac3a
z30131aff091b6db6de65a38bf4faa2bc34abb667e546f8b04f9b9de444dc1d9627da6bdd974240
z7570f3c204fa358a2b6b39b345c33ffca0a5a4be4f1abe2e50dff128ba5822b06aabbe06c36eb5
z761008348db3335b81a66038b1d9cfbdc7b744796084ddc6aa9d71805c1de3305244603bdd4692
z3a75ec5435eb82b24d7c939f0a2477de0250c7db813567e433c5437f58e68bf77914e5ca4b1549
z3cc7ca0a57833d6c133798524d46e77ba94470db488c00eb082a1adf96e3aefd889b399950442f
z412424be816fe36c4a70158c7ed5a34e54b3d9123b6f0c9974baa844c5d496b7fd5e66109aa100
zf43ab7c650e504fbc53627361e6e57af55c626c8bbc59f9ac7c594dc0088110a8fd8bcb6f209c5
zc66fa2269219441ffa17f335b9f087ce127bfd87d3a4ca37cc265459a0949b9f096834a44a04b3
zf17cfc26ce8e58454ee0c83f96a1834f0556cc12e004492c3bfc7d103589d24a27998e42c2ba2f
z734eb8468aba7cb32f5608e0c3bba419a1cb1eb616a87f6727b2937134c59f517bef9644df39f7
zec1b06dc3ba23a5bddb5674b2fcd45b40628b373a5086a107a333da8cc363d5cf6c7f3ee07ab72
z86bf063cb2c8b6111555545344c1a1a2523440ea3bce9de901fcd3d1ef91d6ada11db55d77d9a4
zcc6b71f786c17be7a3716aeef7788448c343c1ceda17579ae6b8bbfc3c53cd313e214c2749ad33
z240c4d4fdbfb230355cd4d25a5c4e2636b6181ea1e7a8e1324664f6828ecf198c0b497781d6fa5
zabaf281cbc62529d7d990ed4fd671cc5b5b59bbf80d1a137b456fbc1be235f5fce17a540d14f82
z5034ab6fa7b1f04855c2996962746cecc18626998cd6cf2b80d3debaa145b0400f826d68c5d2f9
z93748eb29ecf5c9f3e101e6c28542edcec5c476a405cb1f9e0e691ab396f22c7b20051faa36398
z710e70d9dded585b34975c0bc80c4bc9d9d41e4d0924e2cf2c727b243a6cd8cd7a0c32ab0ccee6
zcb926360811a958fa107f1f8b9772d13d50ed8657bca24040d66adbbb96f9751a48bf99916d720
zf1854fb9c5a63a2938aa8fdf32ae471f51a5fc0554775e31eabe45b289e248a7bffa3370e11cfa
z38ae6b5c80de713380ae52228d7ec46e6af464448dcccd7a69edfb0bb424ca279f9b97909bbc75
z963c5fd3f39a4fd6c83884dfb58a037d2cf480223e796a3f941db01ed1b2dfb25e0dd7cb63a811
zf9f2bb78daa902ef02fa1f7e1e2deebb61bfd84c642436a0543ce7318c259137592765e409b3ad
z6b4d08df57d406d8ad56a8eb7d9a9f0406780934771a3fa766b52f4c4b5a5222f7e3857fb6c9a5
z45704612c397ae1f7ae885ed4af76aeecc95ed47c59a495a9511c78d419b3f7a12eeeba1b01247
zb60b3f9c59e422133a17bddcf4c6174e7b2fea4e7c131d4e0b11ec191d81ee27ec524e5fe642f3
zbe2ebaf517b7249bc00853764e0ffdf5f58f6fd0b5f9e1327a03344e0ae87bf5c2378c0e61fabf
z80fa245fde7f0ae1d44af916373b2878198872504716ca322cf0f712b087efa4e0f70cc0774496
zf771e218a584951e9bfa7be7130cf79d8303b57782695133d786211a4bd08dd4346ba30e5375c2
z8c8d7a2da3b0e6c0ecab90af89494bbde2f1e4ee0b575dfa6993a494327583f3c72b8b1b17cf20
zd2d6a686c55a41410b0208746157b85fa7b136a932b269844f451c6fcba149b3bd6ab3ff2c051e
zbffcad895ea0888d47e51e98d7d08cdcd7d9864f1d1c981f32cb97d00e197c4208c071a05fdee4
z1bf774902b047eea859f5ecb8cce198515c1120883fa624550b54f799f6177fc7f181796229352
z1f662ebeb31ea6225308b04c861f1bf031e1d1ed1e67952fd24df0811fa0421eef7e3c7ea1f1d3
zfa76663402fa9ce65ee57df7ac5aa6f8a910c747ef8f40af792ff57f519b2218e7aa6f135210b0
z93b8b946989df2ca415aa9d6439ff570fc00075455d9aec4761df4a3c11d7be5a6200f060d46c1
za7b12c10fb8556b2c513bb62485df899151dd3fd4679070d27ed06d9fa4959f831cc1ea1d20a07
z5060a9979a9e009191fdbda0323a68f4d33bdc48375be43a6e81c6ad1cd10ea819a4c10da9e130
z26491907d7f9a18448f0388a9112e2138bedd09b9327f57b8931a37b7669fb006fa018cc7fed79
z7fca21232ed921ed3dc14b76882b3011b87f36687fb4370e108b50c093ce95c2b22367c25beec7
z4e0eb60de37c573f0dc9c769973f529a1a7e256fbcce73b654c6af6fa04d34f71f5f660cdc18d1
z61aecc1c0fa9beef8468e32d51b869dc8a535629c09c5383b5e48d317d03569008361c7b4dc3d8
z72927b8bf44aee6eb7a464c25c87b68667ae22c14188a431ca888d82508c37587017a39fd2b395
zfb5c0fabfa2650ab0718b698579869511289188042138342743ec15256572d87adac4f7e338f9f
z5b331568b5310cd7692b5cca84aaa7de8bb55e0d54379b4e6f974846190c3d1c022ee1c3fb2eec
z3f0eec5400b36483df383cfdd1c3eaed1d6c145b1117d6b0ed595316c685bdb4065906ffb0f20d
zb1a2eb99541353d1813fa4ff2e23c2cbac1f357a131ddc84467a10485ce20f5865b4c55d91c2b0
zd49181bf83efe2f3b3dce61adba3333892733a1d564a0ce639da1e6c31abf2108d1e1378a82fae
z3187c9b45531f75d85e075cef16e86935f42b50d8d4583e257709205b46e89d63336350e85be87
z23b9576f611c27af330ce97fdf554edda0c0d138f92c7bbdfd3b974f4ee6578a409a29f3226b1e
z7d5d84a4dfe32f1afcae1b40443c3e3564323d335d7f37bd70327978ecc77f820bf07e0bf1a690
z62f5978e375e144be79765b707dd2e75f8f216ca2cb175f875ad48cea89d3e207b7f221a462102
z48d89fb073acfa2232f049e1aff7f8ccbf17b322ad621c966907a76b164a5c2c4697c44c98b0f3
zbf86ddea1b4317d74309d0655c317e90bea1de27575e78f9764d8df6899a00e65189d87735db57
z532bb82b867101504a0131b5b49bad659f0b739d143df67c351e2fb5609be2fa0580a15d0c251a
z9cbfb84d3b091b4fcb73529adb08cc8cb55700204fc496194320e4c14056fdadd146ee140c15a5
z6a4e99be153f5c37d6239852d9423ab6cd7d66472e4a33a3ed27e881174577adab0754f671f6a2
z42cdf8bd382f0d175693efedf8b7bd16070601c38aa903e028f4281ee926be8d58583d68b195d9
z5d99f44aa773a0cf71f83cdded7c1b3ab713378aae63d3fc11a4443dba180226c2014a178af623
zed61d0d7c4dc1831773961882bb4a2f1d383eb8c58a44bef77ce6a5eee77656fd51ca968056c22
z15dbf8e0ae7d37352435e55fe951770d7bfdd38007764ffae7fa4a971f508fe61e73da5e7202af
z08f04fe136cb90d70542a7e84f01e5b83df379a692022190c3b5c7d49cd0714333f415ca89037f
z9ab71c7cf766973d9b7dd42fca4106a72d67db8906ac73167044d36940ff08432258eafd53ac21
z69bca0eb40ad132c978d7f5a174ed4ba1acd3ab6e92919faeb584ae71388da9f528d525de5d2d2
z11c42bf6cccf68db2a4589416e1d40f430f222f59a947673ff1389580fa4ac13e787ea5c2d2fa5
z63e0e2158e76bc9a7d60fdbccbdbc8fb728e9b3efe9a74625c8eb49cfd02f6ccecfeaeaab4f77e
z24991b620daf5bb20176fbb5e0e5dc72c54b10d992a3db23231617190a4ac8fe42d1cf008101ef
z9dc02323b374a6cad7963e36d88fe84f304abfcd0a691e2ed8ff3bf52037939dc62de49917ac89
zae3891fc813ab231ea1874dea369163abe9f32e69f37010f2de3c661470e6805dfa06a24661037
z453a675a252924d97a6f54bcffb7a77ebb547635ff5a237544ef798afb958d75cc81f96aa41448
z4989c22042b88999fa1ba37a8d7923a438328349b442dab77ab185c362b4f37fbc90e745725daf
z6700012f197c84a67fdea74815782e279b6c4b5315c0327563aec045a4a95649c6e609080c9dcc
za76d4dad42c09f20bdecd3f2f94ca60ed76cf585b60b1c73fa0e54f4a04021a6cef6cf64bc3319
z73b00d8346ef665a78473ac22223d58fe7645a6cff2d2258b9648eb33ed68245131bcacd70eb38
za57417df660bde0ccb6a839e3515439281e8fc691ee7f7879a0eb681cd68313a9c05e796f9d3ad
z9ea137eb689605b4a4c194ba827307c60cf156756fe3a83a9e2950f6bdc30c761d65d919a25cb8
z1294a4e212d20a8771ec9bd3fcd34b701c186d1af78e7861335f6d65ee7d2bdc15ff8b8223d92b
z5d2c9a948f87d6f8748af9a60065184a63a17f3e58aac6f5472813e6898c16f7665ab2673588c3
z2963020965483da9b8ca49c604a3966b8e3b642bf815f47e09cc306e29554815d20ffa3f1e6356
zdd5fed34882f2055347a9171735913d1e0d0d74ba65f0721fe084a62e649480cff61fb7f28ae31
z8368803e29daa19d08e379955afe7f3c0d50ef5d3684e04d1e4fa08f6fc48a2684f786b0cee2ef
z43606465d7758ac162072cad86fed24a3654a0ed652415bdb5f43eb643e4579d7d65be9636927a
za0645b9e0b39c61c992677260670ec030981a89808cae3284baedd9cc87953e3120f058c5c7b3e
z754182c8bd7980cde4deece5156da10e83a12eb0ea4d69314b414dfb949e24d1a920674100db64
z9cd3f7b5932ead856ba8ecee743b4abcf1b78e23568561f92ea5236a8dde390ed75b40f138be12
za757143eb963e14bc0b8b221442270992fd3e3edc1681694c31685bfeda1e8c3e827b0cefdd7ce
z7f15a416f2d085fb01fb059cd484c430f2b0b79308e5d30c33aabc15eab48c15960db9ba06db61
za739c0f72b550893a444ffbfe508ef3f724b43e479bb2e8250e24ec081de5290d03bbcd508afd6
z712c2bece050168861e1a978991eff5f6f531ed1ac4e24f96a51f40cd7be16f5936da0f4d5ef74
z1267878e1dd80d6f4901891b8ee32b3fe3a557e983863497790bc30a41cfe0c1749b64a6c9e35f
zec6634efebee6f12dacbae5c64add5249bc04808d5fe01df6aa7c6bf4d6e4f0bf3a6f5547313e9
z09e8cf934f6cb417b903cdd6da5eb82dad67e28f90e99dfe3460a9ab758fd483e330e36345eeb8
z46fdf839c50ab50bb277921e1c71e62c92ad94cb5cb0947485ccc1518e8f3ac0d071da24bb38de
zd11e578a485e4387d1fe9bd3c3270c702342abe34c5d493fe623769af92c833dd02fa651e82d79
zf22d90098bd02917e29854c691cd36b16c22e8bb989ec6bc4d5fd4b200b6a5c78f616ef49c60e7
zae5109d106d31cf21a348304c89cf0a530f0533d9cafd5623330efd3aa74888b831dc000c8f4a3
z41431ae07cb41f7ca2ee79f32b2ca2c183f96c678fdfdfc7630dfc623f1502f2bdb0a64c396e0b
z79e9276c00164b62acd553bc8a3b03a4dd0b50ac18fe428ea2c59e435d1477b4ec57b8db14b5ff
zdf8bd9fff25cdab7b572890f3fbf11326562bcacdd5a5de769dedc659d816fc6890c0c9576fa97
z8b9a5b0d9cf3e883d6fb1a40f715249b30c3369e460c264e37da4e8ebbaec1df3ba54817096ce7
z3fe96432d94366a243544a9c37b5e65faed9590dbda42772a869c9163da3eb443cbb62a9e56920
z321dda584d36cb6a11ab20503f2b58ff2433444cb92b40dd8419565e3a2a0d6431bde0de4bdad7
z6751714147d4783a2b3b16a69553e5053bfa3fd27504a5826dcd3cffcd152001269f978f81f13e
z34687150b94a723729838ea1ccc618699a361b366af6190ff2a0f3ba845b8032776948f84f5294
z0ebc218104a3813af2d7ab8888491c5a7e8f9478d835001258cfecbf811660a11b91319f623617
z1814c019c10e96516e5cc3f0e667133c285f4e4fa53e0ae91286a7f532f5641f8cc4fb616fcaf2
zd7f6ca834729ad1b051275fe8d33b5b168b910be09ed6366918a5093ae16ff10d1fcdca64e066e
z6bcacab25ef893b9d87524c708b7bcfee4f75d997b49796509c84a6ff6563571de83064f3256cd
zae4492f225c077258a8a366bf16a11989979a3626b8e1b863fdf22fbcd332d16bab436d4c7d694
ze916d6fb2cd4aca63e1432b5372458e819f533d2aa1478cea77b268dd9ec6bbffc722fdc213598
z0ccbd9ee6412513730066b77d16497ebe40db65bff9236c61fb87d6e8b307a97dc02749f076244
z8bd6ec335f3ca5917be51cc1dd7c77706eaa0e2961b4d46cfc851dc9592c52bab69ed187710ac7
z5bb0edbe1027a0723ee93203b11a13db724b77c5036c758bf31bde70bf48826d80e250011eb869
z7459728e8306ef5829f3b2be5e0971d0fbf0eb15c15275873bfbd95e29b6af0e5e6bb7aac4ee2a
z8d57cb6fd3b30f6f3a674a7649bda48eef49d691e2b0ecc6bbe8e383a3cd04fccd4db313d6c052
zda2b7aa748dcbbb09b6258c5fdc8ed091f89c1f97bc89e3872319258c6dfd130a49fad822b2c69
zb54f1a5d25491083bee32f505f6885cd9919caada219b0771150e6f0f289af0d314329af135c53
z36cc2a058564a8fa9f5151038f71cdac1b1553c56148d0e5eb9b3fce4f3ca91f1f4b63321b1e7b
z2dd42a84ad5efce7c3224ce9984094b7249cad44f2c2a4f4bf98616abd45778cc77cba6946066a
z08fb3c640ab92ee462073429dd44981e554dfba2b3a8c3ce5d0a7c880dcfc2cb1489454aff2d69
z69714e744c6df92fbd0cf3c39dbafc69b1611cf247dbadebf72e08ee01b05185700a9a30caee9f
z0cf936d0b6573699303713c155ad0f2b0edff1b5472285f338997a838a5b7054243d2d65c96bfd
zf304bdb35702cd7c8317709bff8e50f7ab06321862c56c62608fd7da2fcd6f4e3600b20d99c702
z97339cc5d35db944481218594867af3cfb23896bfe2d6cf56cda66be12c5c87d6a047633b44def
z8154efce7815c9a8b4a94e1822015dd487af6e15dc8d6db8bba0fd47da7acc9910618745bc4531
z0e1510e8774886c01b225354a29d64e1153811d44a4b92694cd5a9d1093eac66f4d0925ea187ca
z81cf8ac8c00de15e7de785e1aaf7491b6c64980d9203b60ab2271d62ae6403046be0bfa6b2048d
zf4420a29d7fc2aa98bc4488b0e15e5916ca338ef2012f89034d6a28c98fa101a5ca8340a80acbb
z01ba34e6cbd23322b2547edc0dd2b29f8081c25154854eb949df49201ae324765fa1f7979809e8
z269542269c189869d86088b41a1baf8ec8c64e92cb0e2347855cf24eee583b2caba099f591b8e5
zdd95e0d785e8aa653044af68f6b50640ce782232c252a38d49c5ff1b742dc7583e1218a68ef2f8
zf6478635ea8ad28caec296b3d334a45cc628766a327313e223e19d2321f11f8bf4c84b30f555ba
z0168b099251ac7665ded47777aafac2add7c1a996a7aa1517104851e453170dccf214dae3f9034
zad2344ab0028845d133944b3acc5d15d2bf017d28053bc58f77806a946408639101103f6d27f3a
zf2c203813d28a9aaa62699810b9a1eb825e150e66b7f78db91fe146e5ec34bcf676e04c6cc5ae4
z8e7ca294798cb1b7e72a4038ae11fce3cef1373c3a22e0e3f8be10d2068c9aae482c3fa9bf9a71
z04d94ee3d6a1bfedca5a80802f070cf057144a599d733d24b9029f8c8a185f2cb8b80becae3d5b
z3470655ad79b5a274ce339b7ef59dea177df078d791355681aeec67ad1bbb224a22b1b3c422784
z3ac8b2c626e09944da2376b53ac4206432f9e9c3749e049a66fc45904370b54f732e3463bfd982
zca5a0c2f70b89a55c5f0a5c26cd9366242257e1e4ac641cff59615d2d962c6c5ed62fd3ce39b3c
z92a4f48878fd2ccbb15cdec2115d943b175413268b5f229b6241969e5287b53522ec00e6b3feec
z1010b946e2bcfd6b22910a605bbeebbdaed35863ca1ef3314a26c75d28755ca6a653945e7b18b2
z3d8466c219f62e42d4dfeaf727092b05892ee577d56bb9e7b99df64f1ce2aaa3db3a9dd3944cb6
z1dd49e24e93a8c133990d340119e42d878a18c4a650776df4cbdfd8233d1796b11716683b7d283
z379bebf671ed3275d38c0ec0197d603814c5729976d33746029aa20a10144aedfe61ce0e739efc
zfa881ef1f3b6095547f2cf37631206fea746b4232a5c37d9ed4f50aeb5be82f63fc54f438f34cb
z894dc62e2bc64bee835a417e8d1b0be186ba9e60a3cd4022b2554a20cc07c04b4b57415eab3498
zad887d6c191be1bd2908632e287faae849ac65924ea9be44863780dd69951f421e3b9df75b4b67
z9159a97a97589e1ecafa65ef6d2ebd4bbbfdcafff90a5715f5d45ef4dc82f2b74b450be6c29f1e
z2d5ef0e9206dacd9cae6d82649a4ecced5780b19bbab5788d60e9496d6b20aebbe3af11af891a6
za0a59c7e2e1be05272d2a64890167e4467defa1705e225a30ba10527ad71827592dde2181466be
zb7fde3f60fa195442425f12ad42f0bd7b89edb9bb42659e652116380c9edc95647c5a28337a6c1
zcf86673a8ecf10077d485f0a459f579c45cbeab9a84a67efe7587dc1e358049deb154777e688f7
z19f49b9e49a63aace69cf5b94f5614a59b91f8a71b8823ed1c05d5e07a20fec91eaff12b973c18
z094708530431d0f432e9929676af9a64a4fea1600edc3b7391f36c93eed9ec0e158b23be384564
z35cc7adbd0a9912af70076a5597bd0ac04195020a381d6fe5b68f7a43eb2cb2eb48201a1e67190
z434c048d51331f58ba5ae12bb5051d2904c3e6223dbb4917b0cc2e5c67ff3a840a2fee946612cb
z484cdbb7f3c01df570147f7488dbb54e376b658b492b7698d4836724bdb77c54c4c5bbe7122bba
zd7b879440169dac9f64880d804bbc2449ee18583298987a875f4a26feaeea644ae8bbcc87addc7
zdf28ee531da00009d2474c528f27910ff9b2b5c7484d6edabae279ad35501c40146b39cf4b698d
z9ee1e9fee541225bdc431b558b5ac29430e0de70135860aa5ce2938758571941124c69d20046f6
z620fbd8a9d3abae45df8c5a6a858f265c6790ac3eb2c0e9136cd5a4628c404484fc7cde89c3cdb
za5caa35860ef0dd9633fda0b481193c431830c64d67461cdfdb81e3a234338ff93ecaa80afb25f
z2430da96bc3ecd8a1af675205de545dd942268f1befa86ebe315e291bb4f8870b5d060fc599bba
z302795e75573991e0318b981047c51b01610d06e99cbe2c7cf91a51236d0c75dd8be0561cd9e15
z1904284f4dfe9de3044554d57ad3acffd94d227719feac471ee0d79b5538292f7d81171d569c08
z07186b8504ded9080a0b7fa44e1230309b18ab496003f1b950f85166f58a77e6e7e460011aa141
zcdb16bc440f16c1657905bc6249654cd1ba5d5b29cdce8718ee0fca5c823bb03361ed5628cf278
zb912ef1d7966a9e7c83ac3c5a5b4867e26ad2db8301b48f2420d531b0e1a9ea8f87f8fd793667b
zfc92d65afdad94c09f721fb45c7e6229ec0cb236624995e9223c13a01e33972a526330c03c71ac
zda3dc7800ef008b967ca239afc8b15ee51ed87c20aac7b3a1930e7a6a06332dcf4c7ae60b9733a
z53318a2bd28f50854c7d32cb0cca7b1ae99ddb008a5a4c66bafec77726592aec81f499a22f57ee
z26bb6de43ab9bf2ac9a34ca35a25f98f4c6792065fd99cc1e59304de5878ee2d4519aad970a0dc
z9ff08199d76f6988e3c9269b404cf4c55788f3a93987e3639ddde181ad0d150c0daf616dc6287e
z75e7752d01c769f1cfb232688ab1b6ad413884dbe16c0955c6045bc9bee8f15b24da5d0fa9dd13
z26e095dcb8f8d8bfe99edad75ca6bcd8dc7ae6074318660c02f5b8b7679731c6dc2acadb51bc1f
z8cd7849f9f0e3130d176925b394e33a78fbe18a7d26c4f476d61d531e946f380293b38311895bd
zecb6b050919ab577e0bd936f5173f9e08836c92f98fc86763becd9ec4af6186f059ebdc9b4b17e
zf2d14da00fc7f59a266854c39a1dbce5fb2caf2ee380c987b3faa51acdaf85790828ff985f069c
zc8097da0c0ff5653d71d1c24a339fe3e194b51a7daf76feede638e40c5bbce5f901a09e1f27bee
z1d5872f321ce3a68e485d2165205b4f6214962ff37d992b40f86963b2c4d5b59b8eca2b783800c
z65890077ef1cd0c1326994193c1cf9051046aafac7afa73541f74e52bdb1cbae2ea85122165cbe
zc05bfecc9b846dfc341b5b83c95f74e8b1ff6bcb4a58738c221f6af1e3b9120cf6b9cd35cabb42
zc766cd46bd8dcb65b1bdcc175fb3ab389d831d5cda93bee96eea42dbdfa06932bbb27d56a8fc05
z28ec93b90151f5e26a870fa17e82224bcbeb25d6ee16b7a3f7e28d1c9347af3b28172c37aa4082
ze8bb99664bd75975c39d805a21501915e3ab00e13b3c21eb0b2b5dae9a78991cd6d13fd9be4482
zd5906ef84758cdffc73c5309ecfe0723ddd3ad2b49d8409a92ee2ccbf3623a673302c0342b7144
zb9242682fc50f055b79a883c0d07089d2f09ff558e6058c3e6084de080637b64e0dcd8c911f321
z1966f3fbe636246688497a32ea2f4e1cb2d876089b5df238f0e0a5640829609aecf206f82a6b50
zef6241f21fde845b79c9405e0d5b3d372958a439edd4267ef9f516ca79a477163ccb55f8d4e567
z01accf01cbb09bf81dd0edd511c0d38d4f1fe267c8dc31ca3c907ad502173b9cf5b82c550c2921
z9087ed884df0f1c02047d18d44f20408500907d3fd7815c59696a713b4eb66a4d72c55c9a3603e
z51786b1b3f32fc3bb0d545b9da6f1c1df2ae117490e19c6b6f8b207289b11b6ec45595d05a68ce
zdd39f78d8da724fa2e5f408a3a281ddcf9a9ab881fae118197df12251dee8913136a94ca3b78a4
z2ad9d21173a98bdaeb086ceadf52a5763740df56828e855772c8891f227c872ec05acfbf7a3ece
za9aa08c3f31fa7f3c9ec3a9475a151cf489e532a0bf944dfdbaa86d6fd647ed4af810ea1d55ca2
z8094556a5017d70233ab7d388bbe81d21c49296c61647f17734f24d83d1c0a9c5bbbbffb0b0654
ze9df34849adeee4fb7310a429e3cb9d2eb7242084eb064d3f13bf381aac8648366f99407697390
z85aea2410c71e50c9c1988fca08593fbeb026b3d7a7bfde7a690302dbd328435759a0733680fd0
zcef3f78b0f69a70ca9c6d23c9ac5749c2851d14f47bf7a7eb80847d0c9583c8a8fe3a68d2808e8
z6563ce7d6b8d632a6f937f2e132bbab9102a7723e5561a014cf45c25469481bc9d2899b99bb2c0
z98acd7ec0fe54e9577a6f3b69cfda668cb9c3b7d8d836cbdcbcce4ce400cc909cc60bc011b6621
zf56db84107daa93dd2c804deba63869a0cdedaced928aa54390a956645c6c9f2abf31fdb482afe
z13659d676711176b7a792cf9fa4ae127c43094065a9f7c36065c7fb01901e5da83dec7966e4a67
zfdf8aef224035ec7e5f689c8dd7cfa3af178f6e4b9cc724c792950ba78eef5b40e2eff559c0fc8
za9b36b078f2966fb3e7e91a61f09d71989537f6a7fd0f7df5399795c12dbb918ce7c1aa7beb221
za23702c4ca7e9c70bf96437fe4dfdb234ff4b69e835ff1954b70f4833db2b887183d0bfbc10c6b
z42577fe9c89037968ae54c83bcbcc274a304418c978213f453899269dbcef33c3e96102504918c
ze7c7402b5838631398fb7b926140c432d0b7abeee5833c698cde9f21f75dea263a8b6a727c941d
z0ee4d3c860787df0fcd36cb3d26ae52f60599ca8e975f93776f975669a875b6b37416b945f8bd1
zcfad121083f9c07e7a610568049b5a07a04c01b9d8e10d6a1ed8a4f01ca64cad0f2a7bd40fb5de
zb054c2e7a1443c0b3c8b6b9e35c6828300775fa3d2276bd918b74ae42de07afe63c29ff0ce5725
z17d48b49e509f7cbf028935255d47647998c9199b9455120796dd9d2aa5ebb548575b83e76fbb4
zfab3d858f53abcbf130982a21053e3d7480db21d89bd405046d448529bca4df3d216f5c78212fd
z29b81e9b57e7e5e6c2db2696ca4fbfc04365ac648b46f8d424083617c83cb6a53f5c92e96f6c80
z834b8a944d3ac217656ce68f120497632c394cb91de50f914c031749eab2c4d9106359611b148c
zd31a4a2b187c20e505279729c102ce6c93faf79cb545c0228631b3b06130f9364dde06f008b85c
z510414a0d07d94720579f5f0e7054f20eb710da260600dba2af2bdecf5a867f4f56baa2773e76b
z11e837303c0c479b49f4b10245e8d3a8b5c05963b3698cc511537fb5c5ddaf8c54e4306f47c8f9
zc03021da3b14953c1cead6d6c4826b9666ff1755dd1b967850e05438f6d7a58516e2fa07adc07a
zece71bc5efcad8d9984a6de1f30d407598481368a030f87cdefbbd1614069b912aba76d779cab0
z29e087d6ac7da724b7939f7709bc451d2866ab3fe5a91c66e8a270bf74bd1e82c48aa263822141
z4cd18be5476ab50c78f78645ac3c89422b85821bbdf539a8a6bd1c038561e793562038dfdb722d
z5aa7ebcb54281d34520a4cefccf7ce116ed3c2415c65990670f29b5ab90d5e9d11fe1cbd973453
z4e244fb6806823044f382a7c4f40c7bfa48c653f77d6c09687461eb0c1f3720f892600d6c0be66
z7b3e76fb3b4c08ab3d156283f2143c01504dff73c619ce47e238c78181ad3c3edc753c378b4103
zf14c7f57b7cf5ba4705368d6668c3884834ffc5ffd68a294d458e28877b0eaa6bf91933f4b4d35
zae18213bec3dfbcabd667fad8aa856a4d96ff5a46b69768e3136325796643ffb3300c4e9d77100
z10bbbdff70388c6f11863129e27820c4629ad02144363d167c4d844fe52826764578eec4d30602
z5c21212eea754b141c3c86b55604c956baf686f820612b2154360c28de20d8fff67d694a9b1254
z14c0bc168e1ad1456460b203e943bf0a05edeeea35571e0c5095633f33178debb3f7d65eb697ae
z7132806e4e349035471caad54f3e8b8a6106cae61120faa3def37209a5afa823fff162a168d628
zb05da0193b6bb50750c6411127eee29bfa077a3873bb27bdb9bf4f85658137fab38b1dbddd14bc
z57e888c232ba7dcc9a0d5c83ad708822abf89bb2934355470f90111623e5e520e74886e65ae4c6
z5de06bfb125f7dc958a9cd1b43c46a5b0e96cbfe7016fb15811c549e727a37176470fc2515aa9a
z7b5a9fafabe7b10ae2488a337c43c3256cc86052ec246bd0c06cdbe8afdab4591e12c57ac1934e
zb3ffbd87fb6c994c62590eecbbcb41c035f6dd860f89ea4a0dd46a4cf417ac19cc3a368469f705
zde2b6d60034b4bfffab89be39c60c35e0e9ca9d0ec6c1532dc9c7c939a703b30225f525b1d1791
z1daecfdd9572bc578513d20c44f2d74d0ae794c293ee90db53b2dad2e5486e243a55c4fec18b97
za7cfa100f02fde06a03d12cfa2ab5ecd6d8e7f4762c01f1b8d22e25446d7ca29994303724b0fa2
z800650894ca30e36e8602515e2513415abc97bbb7179d6eeb67a2bb912a7e790c0f335969ba836
z8c151a41be5e202a5815531c8d2f4f3f3744e4c02e487f0cfe3a7f5702325b77f5fda0f86c2ba3
z6fb334fa734954867ed107b70ec7bb3ed3347a3b1540682a5fff3556d26c4cb154aa6f55891ecd
z797fede14b7c1d34640bc27701c7f8553bb476c8413174a30c328624063348ce9cd44fa2034755
zcfa08da57f27e730504b79f4a4e6b21f1a719684f6a049511817233fb8b99b136061db742fccf8
zf08e6c05e2a622eca990ddb2344bcc4a052d7949cf66ba42f0af97f8c5a4387cb8944ebd6dfaac
z99bbe49734dea52bcf967d36a4c4377707786c634fbf8cb64c2396687e0f8f6b63fe56d88661b9
z3340fe64f880e3b48225d156a7aea21db6610a94340ffa9536526f6d1f8eaa22c139c9f68fbb31
za118615d88faaac2c63e575aa2755ad56cda858f900e3a89a849a658b52253bedcf4ce12dde80b
zbbbad5611c42c8e772e165eca576d5a68495fe3e09c3ac930d25ae102aff08fec98c20e44cca5e
zbc925c5c7ad4a959782fb565f3cdb906fa0296548454ff74157196e3dac6f5919681be11c0d815
z757ad37c334baa13449751e9f8e12fd43dccf92a0291687d4842d6348abcc267a8dfabb8a92db0
z91a6db6793be8d50fdbdf6f67a73b17c123e5df00cdc864e75046e21cf8bd3e353e2b681086568
z04af1bba2d7af04eb65cde67ea9c98d10e7a0d627cdf209d5c1263cd187e5d3c5639e452091469
zcc130083cd85c3ef2a7c03ff3cbe90b1f006b95ed56874ca41045b554c8fdfb0f93be57cf595ee
zd5e91300f08fea97e8fca1d564f8b99f6f79df990f26b9fcbe3056670464230c9a6f4e9d70cbc5
za399973a290925eed8cb3b9581353aec754575c2782e8d21904d245e63356431b6b0873f7cd273
z328577c1edfe7275e9ec95e2c516ec4a0896b039b59f495d118ea7a048f3535e743a2cef9d1b55
zd74e6293269cadfff68a4f681c1e70e229ac63593ed0c99e270f80f73425b9f0c3b2a74fcb57b9
z4447512ba57370291bc29ab5f19d625a5de14f0226cd14677d9c158b90dbec262b8a54a1f5359a
z341e10cffcbe686aaf06da28d47fe74cdd57e5a61d94312622beeb969121db7ccdfcb47e04caf0
z7068486b7598a110c42c9080ee74f11523d736d01be1be52bc380169400d307d9f4c8bb1ca98d6
z689b0f7456e38c21d76617b362a7ad6e43963dc1cbb423883053cbf5cef28434400536e77e2679
zb09a7ca89f06a9ba36a57cae64602da00f8fdd9294146c4b58589ade9352ebb2bbca0c71c38368
z9bf1c3075a0a72061b28677495dd1ca76b9e50686e8194913a973b0bad44f9238bcf388603a301
z93e7879d55b6f0d66892af617905bf2e92067772139a952cd3e9554f47f2b86b2bdcfe0b6c9e97
zb082576acb3e58c1e2ebfa7db83e9db62f90bb50ed0bc05e553fb3b78b9cd74864edb873562ebe
zd092e42e27e0191effa425dd57d6a350bc3de43174439414ce4943534070de7d1b2f3fc9e458b0
z0a23505beb0b6fa79d45ea53b96c91b239886dd9ce1d82bf118b401fa390b742f77dd4790a52a5
z817d9b81980e57622324884c0c10db6ca6beb119266f0e537e26fdae9cc56f1daf49d1e423c925
z9c6a8564c4a3c816efe812b6b01972754133a07f42372d38c0370bc4a79ecc41c7113561c929ff
z48662301a17ebb09c3dad3efb47cf76651a66f97f5ff3a0a1d17c4d728d0680ecddf393e419adc
z9f52ff9371c062d12de75dd7348e2e3773b491636d1ec3073f9f8313afa355ce84ac3c6fc19073
zd97fce8572fb5db0ef8d0f1f4484b957c4d091b8b487234516828b45c38d6ca7aaf8fb690de1f8
z57033612b2a6db5fd0cb2b8bba8b3996a32ef9afa7bba4dc99774ba9f7f460eefffa94a741f6a2
zd5c0aa82241fa413709faa5909555afc30162704af9452f3912f58c12fdf43660a0e40c4658d28
z6dc70f7c10d2730068d99ff4dd8cf4707198272751912551c32d46bd35d0b98e2ed78d62caa6eb
zbbc697db6790f8095728b518fefd2a30e90ae2ab41a426ba146373785efdc11fa1bfe76d6481db
ze473b83422465c97271dfd7a3ee9a32ece8904f0d9995146c8f9b3a4ade4f0711d074d5b6aeebd
ze6f81bc51dd6a9a6952b7662abacfcd80332d4c2ce25a58ba1858dbcfd64e226fe4ce556587123
z522708a5d1b8e149a9c1c01f7009504dfede6f17374f146557ca6854386292b8dc8b189fef6cb9
z203f52a6d9c1769e9df67445a002d82801ee383424b1e08f5436ee824903006c1fb56fc097fa1e
zab57212f8fa06a5e281a52268cd63005b02aad171ad266c1abe8be0ea193f872c9f359b53b05fc
zefa8e6f47be8c230e95cff41c1cfd42e34703676b852cbb895c00621177bdf5eac431e90402ab5
z8e7342e8bc31a63e036b1941136b423ce3f4902e51addde55965952f239a2642eeaedbd9150d45
z698b7ccd0966c43118b5bfba48f9f32fd49b6c79c73c865935793c5f3d0a539008b949037e9712
zb368e1df10d17006249496a540e250cb5d34f5b0ea90520815658edccc2df1d58aa3fa0f0627b9
zaeded7f75e8010d1b30d66be904166c431177f711ef38556da3c40297695b5d1a9d5366d4e497c
z468d893b20f4d9bc882aecdc0c3dbb1d91a856f997a4583a5cbd7d3ce22f54cdc9a888a1130028
ze5b17577c6c8e52e61512b8b6aea1b3f9dec20d7c3e0923803c4507d6c3c3dadf4b6b595b43f35
za23432195be9493955b1fab4b91b948f86e0dc28f477da0e710a2fbce1747cbc8ce0c952761695
z87a7233a8b84da613c777aac743bf6313a26ed844f0c2ec3227ec2f55f18c7989d1e2641fb2dde
zef99bb78238b5b5e055ca5b6ba20c2b80a6e5e1ab4e9686057f0d31816e62b6f9130a0b0ea864d
z6a7cf76407b03e0cfd15563905c4ef4bfcde645326328c187d5618f7102d0082c118cab854a074
z26848f19a5df6778194dfaae804acb7709c88c091ac6bc9c0cd8b9d0763b0ed0559297ad847b0e
z6d8373067eb0fa054ef68b916c3a5cc0f58432068322c49c486e9e57be4ccecb98e4f85a3d0f3a
za8d35d4fa219b3012db4885108dab113e5d11e80e058eea44e9272bedbdc2e63156cffd1b46374
z833ec6e56f40d1911efc74bcde4a772de97e41c4e6ccb939c65ae1ac07b24411b17237ac6e8df6
z5b7916d74eef8e81d6a41abdec93f14eb619058f7feb7e114fe302cd179cafadf4abce3e62f88d
z4d9659283ebc91ffc648ab9cc6d059f51c6b8737f864c433e55a4ed55d91196da67a15bb51e763
ze1b5eababbf15c6b406f9bfb088b0d6030fdae0fc73ffaf601f6da7ffb6fccefae7442432c5b50
zf2e16c14c90cee5e4e86460ed7ada0f2b7abcb15c2d9e38d2805b64efab81911c030bf52a9f592
z950bf121d50d49cccdc25613e13587219decb2bc56d8910fb0a3722a145c2bb4a33ef35dc6c689
zb9f9687146c72928185f7b4977995935d97bef55588a72f5a4fdabc20cb02cb53fe4bce8c4d98e
z3f577f6a999c86697c279040569373cbfcd9e5cbf9e0785824007308fffe4341387027e1e06709
ze5ecc4a0be1bd67be2cf36e768f029fe818937a732ac7863c5736c612b0a4f0b4afbf32c55496c
ze9eed56911101d8fbf568ce3b39896e64900bfe130720a3b639bb1dd648f57247994a9baff5188
z1f83c0ebdd3dafcb39944547e3a4ca24f7fbb913bbcc2769d58b1697c874323e0eee4eed9b6867
za386dede8542427c8311f382f7700211ded7283c48bc329ac3d58853d083f38627929ed6718f42
z267cdd71c5191490c04f9c3c736cfd0f6b6fbb9428ad4e03614ec25e8ec5c7a788dade04c5c118
za3b27192cd48f51d13fa607c5fc814c48060a9b7c442fb9e3fa993ebb5c81dd4e31cca9cfe508e
zeb40ad665b6fe76a4be3945cd0450e81bc7d7f6d57d69a287a5ee7153d6f565eb3a23db567a0f5
z71601faaad87d434d2ad9a100b65ca103e2962f5b1de3e9fa921e7de00697c8db0f405625be467
zec142a0fc8d544ac369fc378c34e576941ab71db8d6ed14e24174bda794e51f4ab1dce5075e245
z52d4c9e8807613ed0b5dfc6565f07c607e024efe7b618bd5240e8fb4034d70f8b856695bd93e29
z221da570146ecdfa078c9e2d3b38db1032e1a5d20d84633c7e8ba143e360922206622e07c9f5e4
z83cf243aa5ca21588f059f6d58f393fed4e97605843171581df1de6132c9d38a7824a6b17edab5
zd2abe8b0023e366f68e919bc9b764bb79b0b9225bf761b762f1c8fc087e345a6ddb94b35416e56
z70485f040c78cda2ce1a0c91db31fcc009335345b314802e75a1ed2169e413f70c53e372f33d6c
zf4fc4088b3b6646ce178325a9613e4195adfc1e58965d1cfc80cefbb97ad53dcad59a90c90cf92
zfb52cf323e464bae3d167805b957d8bf6372ff746f23f276b75af920ae8d7f2480e04076cc2b9b
z198f8bd04bd78531537f6eba7a37e8e178faa8afa87731040b101e031e0251b0a34b6bee0c5ec8
z92e1505b85a753ab32748dc6b5721b6b411348e24bd86b81b7c01b3bb822004bfe8610b331e0b3
zba11b26fa75d10ad096bc2e0a8a0eb22c7bd52053bda7f85133de09d5b685473b3ef733ad0ef91
z26f22f96f9ded6f3ce8f9decb4eeb3e6574adf9cbe2f54c0f565c3f30f83a65784a314f170a77c
zcdab8788fe5d095e7c3bd4c2d693cdef15b79c128afd0410225110b77a4040d84fbcc88ca2243f
zf58dd670d5e03a0e01916d03ed98375dfc75e9c2bc6d817c8ef0934b0e05fe289c0928358e7ace
zc03eb1a6f4b246b037b9263ad7482e063e479ef2cd5786c4b5dab7b4da94a08aacc1d8aa05bf10
z3b80cb46321b8cebb9f913d61d303d15eff977a089ced64fbd3b8e06c68243a9051d2b5b9670be
z8ba3f887bb8541a50a35c656e4c58e42f441f8485c3f1ec0bd0514f241a8b94240f4c201c1ae34
zee8914b54ad516d7ba589c217095a8c0c9bb063892755f9aba9e6cbfae690b57024f4d2f0c3f30
z79c57b2cdaea840b652ca854cd8f380c07e494a511ebf359d7e54a53a1125bd55777ad84a70335
za6415b5e13a85e541f70dbae2536e6a01b9ae4671d76701219299e98b792cbf1c31707bf5c19cd
z62659a684679a48aa62f30477096780a25f407e61854ffb5fcebd7920ce0d34aef88fd0f9b0a36
z369e12c54c44831cb2af59c93ad9f5060d7ae8b5fe4ef22b76be3ca94d7f1bb87757a62f5386e4
zfdef37a73389c2ed8a15bbb1bdd8d5805da113b8aa87b2e122896122097a3a26f1d2990c96bc18
za0909d0d31b3bb8c40e6d9078bfc9fadec4a780bf935ddc9bd6ee0409e3ac44f48f502fea1c236
z54758fb87ae4c82b5d332a5c900a952922cba1cae878ed1987af6203869dbf5bf292a2cc6937fe
z6c1fcc1855a41619f27237c76f645f167f0caf76090ced10b2412d1076047cbffef90b55854aad
z2bb36217f0c62094f6b79c70d39fb589acd681318dbc92a1f9ff59502b2e4d22a96c975a1f99ab
z3a0e775c58fc7cacc33439cc6f57b93eb43e4ba3e58ab4c9447d5c8ccba02b4850051318d88507
z8fcc243705c343801c030933c40abec832b34ecf3446d08f455c09b2ee06984b77dfecd9d41b71
zc5adff10597e83edf0640d7b59d01b58863b46fdedcf8f62d2b68e2c4267bf179f99269c3b890a
z96b41b989d5a8abd33b5d8c062ede6b0dcf3f7e3b7755cbdd6d6dbf60f740e059f8a712c8037c3
zaf01cd7d3f930faffe25c1815cfe7206a7f522e9c8b3feca658aaeea3693c18561dbbd44215ca3
zc9332e17ea3c14e85d52cd967813e6d079e9ab26ba880414403e1f32e93a39661fbe98c094ef5d
z240b3cb7f5d4c88c6f12094e903f33a6ca92a50901bff8dacc37946c47aa71d73594a3bd67fd0f
z3366be81a00a15dc660a5d441c3de049b562cc6af6abb66a4af731f60f978b3bb1c0928f77031c
z663985fc64732c8c321769d4ee68ee8602d9e928339dfeafa6a1a6ca4992013c4f36a303e8c994
z418d714d9166d6dd6de1fec62080c590b5c8c652bef9a1be5e8911456245f93f6c0fe791115902
zf159785084763563b1896e212609fa66987976a5b80f1fa6c38131f7e248ffe04c206b3c403dcd
z19886990847c0a07fb579dff4c01150e88bebf562e4da8298ae3a00d36daa1d10a0d2fe61e8e49
z37f624242d5d7a739f1e4c97154777517b8b3130ba97e7097d6f7a3e6bc43559a1b9e58f8899d7
z2b8abfbec3a440adee4dda4ce0e91e0a831f45dd2024fedf84e4c3560d63e364409f8c6d9bcc5f
z7e3560aabc4724f5a3e5e54fad49e8b2e55a9f8d8716fb382188d4a3390784b1647e07e95da040
z1142d4e4d8227b8162c2ae110e486a3f6ee40316987b86e43c7a06b3ddad07a59a1125b845ae2b
z35e7fb1f3b4b0e36ed89d6df2b9a326ff668215c89110f2c425ecb688a61c6a899369428544701
zbdc6d14cd2f646b55cc4ce6758363b674059aad59b281d0e3d5671d486d2704eb5fd6378bbfebc
z3234f4c11fd43447ea92b5c9bbe22991b6a7fcc2d7ab0bccd6c34108fe88a2a35367e4e30c519d
zf58803dbb1b9b8f7c47160d7571d4c0b8031a3e2aa58bc92a3f63d04cb1d3cb8b9eb61a54d9b7b
za9283d458fea9960339dccbbcff5e1c8314dfce3da2752e4c8e2d4d995ce17a6b6ce3e621fe363
z8585c4eb21e6aed2548aa55671cc91466143cddb4b220bff69db0abca54e2cf6c002b2135d7cb2
z5ea5d5213cfdd3f373d39657c3022588643ec8b3a729388386e8c849e96ac8b3d894db5c66f057
za2b2366aa158118b461b67ff5d1edc9419b5d2c671727ae427336dcae0589087af6e5a6ab5bc96
z0c5de578e94fff86fb0acb1d52df4f85692a236287ac60b67b62cd176987b0c9148581761fd1aa
z8c788bc8751f77eedb29217df19ec45e66bf43d970df35a5d1780f498c481332ebe8223208d13d
z3e7aac2802c106addd0d8ab79c885788f32f9ee0df75c0e943c080c08880032d139ab557ad81b1
z0835bb45c649eff341a311af920d339c0cf8473f4296b66cfd9d2683ab449294c0eb286e843dbc
z4e8a93f7344caed0a45d19af7144f3983829b00cb2fa44eb5d8a6ba0a26b843340caddc0318180
zf0f14fe0f3c8e666068cc789c0e8dcecfab4ea7def2356a2020216359036e162ff4b8071a94113
z17cbe40163271ad81a9d6a7e72da28d5834080511bdc72284caf60b9c93689855e8525ab41ac08
zad40e6e6195668f35c04976c18ccd171080fc0b3b58ca4fbe8badf57cd7492475c2238f9f4587a
zb4f4d828e6f7fdcbeb7ea56ac74eb8229a71069a9b8b1fe2aa327b00decec8dc8d9050ea74c1b5
z92a5d31b4e5c3b619f0883d7c4e5c81781b6b069e6f39e4aed33cc011e03941726edcbb8413069
z90aa2bf757a1d0eb98010aa12640c5a5a01ccbdb8ef6e39b00ea8a93bd0f160a7273774c728d87
zfd9a7ed0ba3403d710daf43bf026800abde45eab90d8af699d8d62cad419888981f5f498e1c791
z21c3a4591c5da94ce8e58c75a5dffa1d8a7538818876b1239c28bbd09bf7255103f9155d2bcbba
zb8f97f275bdd047033702ace38c221f9c077cc82a74bb4ddf6de23f854aa3030cc302aca4aa3e8
z91f1d5214389efe45b00f2b68e631879bf91950ea842a45308eeb7599c0f004d22ac4cc7d7c40c
z4edf0f9b3bdc61f1075aae99aee5a98f628aa6a6f333f6e114b2c309effb0b5a567917228c468e
z581e07d5600fbf560c17350a6cb290c77148e9d6dc8c4f9ff91728e78e1c14bbee68e4ed7f52c4
zeb1e4b753980c202fb596dee10d097b92c3e141ad2983321bbd2d2b03183ec4d6e65e29d8f3746
z18fd11430e91aaa55e227282ea838ba449bcb60a8c4e80372fe255174483d26102ac282c045863
z1a75a6930577f7130912b5025f9be1d8c3d94a9d3c169da19003bdc083791ce18f0207af795831
zee2b7c13168dbf9b1dbc3b260db9e6c8e08df3e9fef26aafbc285a3e026c60378d5762a6b185d2
z18b3b52fa4b4aed29c4e0209e410c3bb70658d1c78aef7fe46ffd0dcac9bc69b6e3859e6f19839
za6a7bef808fc945ccb2f6ed1ed050149efb79bf1adaf1b6cf01b5b11ed145c878a58d67daa38bb
z181b9eda50c216d037baa5d08bcae9d82e6302bad67a481f8b3728f9a7d1275d0d4f5554ef129e
z7b54912242fe155d89ae9d2611ca726f6b7bee8064b19ae4045154eb0da383e8f1579cddc4eddb
ze0ed5c03ee29f914bbdda04fd3e99a865ad6994bcbcf8e36dbde037d7dbad967c72656e2cbf599
ze0f298902c60e7654df73585352abd9905def9b19067d39d77794ea167f4441c4d5a1456c58bea
z5b930be64ac5858113f18444222cdb60d6dc35efc7bbb699d96d70f04496d7589af5852acb3a6e
za9680fb11ed7eaaa482efd4e0ba2ff5694e170cba448bc02feac31e1ac8d50f7683da52e056658
zb54463f0c10b704fd9fc82079b4f530ba860541b792fb06e08fcc54e54a592e031729408718154
z13ffd3aa9fc33c5a836e07c243fe180633f3c52e337e0e32a6bf08445cba768e4ffe9ca5de625f
z8703c32014a623366d28d150fad3935e560ff19e6dbeb810b931d29b5a6318e11f12ff69bb2f50
z306d2f8210fa2ad8b2cc6310f484fd09d4983224d5f7b3dcebb284000b87e84cf0effdadf3b694
z72af458da566872236a3de4f924896c1f7ae3949010d5fd23f25282f6470392b7e0da1b57a4af8
z2b39bc0f6cc474ccb7852ba95519ea6d44cc5dc5b84fe1f8cdc5b8fe1063966475e5de90140550
z6ad39692fb304a8ffa588477ef4dfc95b2d7c4308434a5a0e896d1c008d5820caca1fcd011bf04
zc355377bad910a1299523e272d8e3f36d46c38829023ba42cb60bae62d25485b12adb250f5411c
z69bedf19ac59722837e05da638d14d3d41b0d31678f1e92df869d41a6d7ab4ec000c6e3993e3d7
zcc9c6c03731850e78986be878805976ec165bee65f254e0fcf24f754acde8c3d656b664369b504
zf67bd49d62edd45684a8c7f5628562d5ce9b05f99aa51f9264c4b543f58f4c86dd7278a26b6369
zc80af8d3b6a97f82cfbe8638067d4e19d3764600c773ac93b93f1a5934d98c6132e87fa91b85ba
z355278caa9e6de8206863b96e095b654375c1620f5a5d73137a64aa8b095b307db07a0477c7a4b
z0909e2a7afd8fbabc56fb0459aba58e1e2ee68ce6048e6dd91c75bb147dcc326f0f050e856d59c
z9bc4dc333b4b3ed5594f5231019733640fda5dded0db314fbc9fb7418f251ae182d3f8a5dddf82
z7429a9a1141b955fcae6ed4c20f7bcaa3aa1e7fa02b135170d56ef1f45fa5b99ff0dab88b10b90
ze000165e51d77fe1c12a3c58d69c4ef7cf59e3ba1fa5f7d03d5fddaccf7f47012f0b862532d350
zf36591846e8788f3dfd1c44843f4fa5aad88d01089f91c8fc45e3de4e7bfe0ea744f4a4b17f0c7
zf4271d3982d3e7d65cc65339bf343c8607b00230064254cf798d82394d108c318cd53640ad9195
z262b4d29c59b99644080fedffdeb260e751f6f1c26c6ab27134963006e21030f0485a213b2dec5
zec364c8cf64ab6d2cdb0744409ec0bf552ce38cf9349ccdab4f7cd9be05b7b9ad35e828aac72b9
zc95098d34bf0c7a2d6ba4aaaf0ae0fb7631e17f82a0e492f9017b6dc20932e0eb3ff022639dad8
z01d7bc26a55dc743983d7c48d3c49d0a7a4ffa60fffeaeb5681414e199e7a1e0a4a7ee226e7ed9
z7b492282955f6957471d62265b0168d854b4be79a933c2155a27fe4d2fd2132a739e8dcae1acda
ze7592ebb8a47d402410adbf6cdefa8ba41e01a9e365e6efbe77145d554f30b3c2c989af9579cbd
z64ee6788c223280aa0128230d4cd26066fc2e366d5ab0596ff2e93459bda41f0097984ee472c7f
zcbf8e703fff802cc8acbeb8edb1f13e342260c76ac2e404e9230178331c0e8c11020cd68d8849c
z374f660d54cf448494344667ae734cf663fda125a5710febb454ade18070862c38058237bb78cd
ze5cf62d4766713193a0b00c2b8f58ed9aeb12bc0f2d54f1460161d7a00b1e8e7c549ea877bdc7a
z7f877badc44d171d99ff5d9c2a9005af98474dd2d6ff3f279a8dd63bcb833e69199420574cf26b
z2c06094ab871a6daed9bf8ce2b897ac11d1604da5b870f8e2478d32c48649796e1bdb01ba98e3d
z1b3976b66d201c4bb27e3de288b88aff3c789285b662c80a20eb4dd5f62fb28bb2b987d41c901f
z6cae847c2dc882af128a97d05201ed4fde0aa18b61a61da5deb7b3a5c208c760e78a1f95f53149
z21b60aed28224d262d4b7690c759a1a03ebe13d25aff65f9719bef6f303ccc2f1e6d9b2e7ca89b
ze132feebcd6077713fda2bd3d7eb1832da1170c01ba605594673d9fdda10b206795f76ea975d14
z9b8374f78d52845bf5472b339e899c7acc686f70471182b087d2cc15655cf1ab20b01aec2f55cd
z8061ff68c4d29fc27f9cabe83f489c886da386e19f67cc45b48075e5f320dd72c5e74d7b9d0245
z86c83671d77e745ccc660029249a99becd6f8d70b26b44899eabf16f7095d265b05bf347d92dc9
z58350384fc68a5def6892ab10eea632fd1a4d455ac8512bccb03c80fbd834939a34254b79d5ed6
zf3f56b49988f8b28aefe4e67e49790fbd25062d7d9c84f40fe5a2894b9d92af36ea16c48e45275
z6e65c72c1b7938ff5abaf553513487f0e5f37bec6c6b6154224fef77e5be3e5c996dacadd7b808
za6ca7598fbb37137cf7ea8e060df3f178d4f45ae71ec8d59a2eb64cc1a647fbc4d2ac829e5b92c
z9417939b0e67ca78fb9c1f83acff638151671914bb3a9ab5f430508f33413815bf0f5179de46dd
z9369a2a2fa68a5a4e94a711513e56fbdfef209c4ef517282144486d8a0fc7d9564446fedf1eb33
zec66649e7f7846f67d3d666086aeef4093158d032eedaff3e1a926ae1638c14dceecf1617304cc
zf683a541fa74304c99afb60d90ac5778946aa2466b5b7b49bf7c261d168d510a19107fc35e75fa
z639cc56396340e381094d62a45aae20a0e69addcb89384a70a9cd458c02c76c94bee9bd72d8491
zc0306a15f4bf2d8bbda83a820b14519a2b3219bd7640fc28763ceb0cb34c455fb9ce6ac74dd963
z7499d2508df4383389186d773a2d9a9346f5dd1b4a2a06a29c4430dcf55faa92ea843fb9403047
za71d502dad6d76cf82d54407209203c404b9e717dbb3edba96f5d4f911146ed99adf8bdc58a4fc
z99c7c71ea51a80ec97bda4e054cde532e71627e1589115297df71a4148352e27103e540852c1db
zd0386232d59b5cd252886755824c84ec3f2ce9a73189a76c7002ca3c032933615bd627e7815374
zc1af82f7711efbceb63e722616d7d171fb6baa880586f5ce436046c458ac473aaedb5a5dff5714
z6ac9c8a71e967aadc5794929a33714169e1ee395d900ba62610c7910f19b4377b0ce0b9c30b47e
z88adfdda2b05308b2cffd482a8c8aa2c80d4f3f834184e9c6da307577da2acdd03c0eb32164934
za116d66397bc30fe02494994df2de9c12bc434d2ba1fa76c6a27c72d47c123524a1f4a572b728e
z725af6bd9c4d0db09e6cc46266b33b74db47880e49341b269fbb9e04cb1a6e2993187b06088119
z6047b2c0508014e8ec2bc2dbb4893458a257366925378335fadacb1c973d3a8e035629cf568285
z2da3c7df8f30f78a24c208dac386ee4823c8cadcb736b55f6bbc8fb023bfba788aa34e18534199
z491d66aa9115a25627274fcd929a4c14c1fd17fd0e0504cf2ccafa9fd86e44aeb70e73b09519ac
zc2f07420e905338104a8bf54e497db168e7e9ee3f20b458d1d8e55bb9d7a8fe22d25cbae9b94fd
z4dcd6d93a247af32321eb8f79aa535b47e9b7f1651fcb36a8e2706a9dc1e2e144458d2cf24e5ed
z497fd9b746db4ff596a4d56632ab6b14f835974c15169ecef80c7128434412962a3d62e41c9001
zea93a88dd25cb28cc5b09836fd6fecc18ef95f4d2d15faa425cc6d555995f88d88d5235f0bda0d
z767697a54a59841facd2fa702e369f73c1ff826ea190d2954b609ce2dfaf6efe3ff79d758626cc
z4967ae76dd77e5c01aa3e24cec3c9d08ffe02fd8ef43e83a7e7af0825a40b7d269402ca0976420
zd320d04dbdbc29d671197e84398e0da056e2d3b8adec23b445171e8793826193687fefb081beae
ze8fc8febbae12c3e16ed6ace760b7ceac2276088ed51865c6beac6c68ee1d2f84ce45f3d1e9fcb
z95d55a1f4c020b2de1b553ad3b53f96a4e18d4584dab1c390308c37a0d4cae292d423772551620
z5952e3bac1731013cabc0d761a80584ec7b7fb18f11ce9f27c72e2d1d750b676cdd910d2d945ac
z65e61f3247009c625221facf93ea63fd687e97f675ff58307e81d732075a18e4bb145d384da5e3
z1a51fc79f6671220a480e0d95dc956f170c7ee8c6254dde1ada7b451be66ab7fc47a34b4d8c41b
z6399f833686cbab0ce8bf8be9d4e43bfb7a4d4d4020eff8a3c1eb215643fe5d92e97512183e719
z13c9b835828029b0813ecb8b0f55c649731e5cf8dd38c1bf5cdd69a1abaf033b5aade8f921f2f3
zb6025e3e7aca8055b3e4e2b23266d3daa360d87703884b9f20357b87ad5f00ab185a0c3f60d4e2
z2436b09f278f7156ed2b89b63b7bdb79413b05a809e57e9c8b0a50ec336d4eaf6f0f9111e24c3b
zbe0fe7566a7aae00399c3b1d65f55666e3337e68f49e7906973401739317a6fc4a3037b3afd3b0
zdefe41ba0ed25387488e2fc8d7c7ceb2486d2bc1487f79506cfe628bad3d5339ae20e58733c273
z2f49e4ca6a7dbb589477b40ec14268900397df80753fa89c5bef1c25fb89dca00a4819bab769d1
zf2f1e01ba82bdc8fff0363afbd48d5cbb58d21e3736b07694ba821e8cef588f1e6fc86770e77ef
z34be3483107e50b776d95a84ffd08ff411d956c6619ff46c26d9bc23159f9ae220f441feee0ceb
zbd839676709e15bbff9ca1f042590a75d38d5389d841adca5f3b11f1bee3b4a6e6ca251298ef1a
z104233dffeecd7a12701825dc434aa35c704f23fd9bb56c08a835fdd6e7a4293edb18faf98de67
z52ac3772e3241861785c1bc3b21d255cca8a23424920ae0b0590721d2d554dc1ad2240b20f2ba3
z6bd94b7356a868e09e1f918c182829e87843c9807490efbfe4101aed27f99d0b80729c824f73db
z07d4e7d64d7cb5844e6e6bafd45248a86da0512439eb175cd4a31354add05dc2d41dcdab916027
z08f911933f02efddf126bfe7bbe1d2f27eac6a656a0830f2e3e95d8650cd16ca87eba6e2541ef2
z49c1319a59d40c8155577fb983f296c95e8a6eb0efa7b10e33f7eb4d57c088f66619b06a986b01
z63efacb6ab5878566922f90d735add6892ecf28d24d2e5f2c11c8e4ddd7b42ed3f496a8f655376
z88511b4de6fb72792620e04b9b7d1b35f5ef44e9513b518a22b78a26d87560d40cf23bf66ba0e6
z6ab45647138c255478b27b7eaf98a1ff30439aedf5ea3996fa961e9cd13a046e11ace4069c9b2a
z65cecfd291ea45f9a5a25b4e07a5f1520fd817032a59170f2493fd33281fc539867134c3d1c471
zf163b498922e2159d9d8890f7d6927b63a2b439a4adb9c1d6e8ba31f84a9d0b4d3d0b5d90d93bb
z939cf64385bdc090ac85284ba3286ea32f345dd0e48008daa7237d5dc990735b01d6e093ad421c
z3ac0cc59f5dc7634ddbabe2707a59d282c8a99c879712df9abe6ac1cefdeb5568aaa0df0c2f975
z0cff48cf7286af09b63a8017fbf6684585cd4f0b8fafc82d7db9ead3504ae7d76bb83450adbc43
z4aa94ca05b5ce917613056dc1c4145d1e4466b5f86b661b08e808049889f336ce8b5c9126e476c
z7dcd3d7f9f80490f1d4220e3689d3b28ae438fe7554c585d1f8e396e498c88f3e5540fd102b041
zbe8314600da2045a9ce7ed6cdfd706f776abe155c271b7e6a182961178f790ed87aa3afd76360e
zc8753591dc6e2599c09daeb0698f9f07f01b19a9acb524ae55f4f0ed9113fe5ca2b617d693c5b6
z1950c444b50c77581c2d6000f6a4416daeb46ab8fed40e542032e00bc4ebaf079d7b93e707988c
z3b88055ca5ce1b2367e6309bc4491ac845c62ef0d67b3e47dc37f245911e30e26aa48dcedf9046
z01f85a10dfb91f38fab5f64df3831e3219211de401b33bb587210d81ca2124b719173d29bc034a
z88b784da8393478fc87be9a83eabdd78e3bb9d8a3c6a726d91de0c311fbd373f12260085ace77a
z10608c04b0dbad49f9510c2a0536580f093b8dac444626e10877a5361baea562dee634a6152a8d
z397c01fc3ff8397a054bad7312c88728edeaffd5f708dfc35deaa5cf56bf192027ed357f557c28
zed636edb6595f5db3fa68847a309d6d1c7eaf83f54e6ca249ac4dabc1d3d57455e4e64ebcbc778
z42f8d4525770deebc2df7d4a16d13c2caae7ceefc8144841880f4f1a050d5e231e612474793b77
z407dbdca8c6c3e6a9add05320d928ee9794930073b79baeb4985fc1e8a23c3274f74eb76e50f5c
z8603e6b03ccefae4679f10fcf380403e4eb097c8ed83d2cf441e49a07f5fe2af35030d2f9f1a92
z9bb6ddfc61cf79ec4c58ebe64a7927950b70c8c085b52fa487e07290e9858a8be0b9d375bf8477
z1939ff51c64adc55bfaa8939f2b87dd5de124a7a2362b53bd7937f77492fe2ec4e2f250c5010d1
zfb9f69c34ca88d7e4adf07571b566171a644ac9c601356e24ac48031b96cfc39eb06ad71c7b569
zb15500ca04e19cbdd17eee56665729d28eba5f9e59ca2c3d2c85acb14616e1b43240346c296b73
zce1a5c755a20a0c87d7261282914742fcaba3c48b408032279bd0f7bf62173da62c5c1a574e042
z5c0938e133a660b05d2201c125de502d9f8af2f6431a2dfb29b4fa33ab608b4ba53fdc5c794a35
zd00c662fb78188e750301efe86e4a8958f355238daf38dbb5eac1bc1e04c01d90c1b6f458c7cc6
z40ca1feb8ebce447fbafbd762ada05e1c9211ac66b72abaaf40d06ddab353b5d9fdfa3df4153d6
z35cca7f01e9af0a64c1c587ea078e97bd051fdb7c15d1eba0963b806f47d19e9d5140ffe26ee1b
z6c052343e69cdef4cfe0669e4ece6f6e6c9d76667f793d63c24dfae22089ed11c0a5d780ab6f93
z714a38a72c34ccdde30b2bfd45d487868a5f5958b44137749f99bdfd1062ec98e8c0594d4ab9c4
z12c5cc5015047e959dd6f31351c3b1aaa9de4ab13adf2f4b2b4648b04cc7ec95e6515f77382d82
zaf6ac74faebe95d81eea2f7ef86366b0cbf395bb5b2bfb32e88a96d0e876e2e5dca966430c3d70
z54a6e1a26953bec1b39a5ec41dfef5e99493e787b2b698a30b1f8f8e45cb427eae3104fe235d6e
z3be5a7d6ba46d7dc46229607cfa3803de7ecd5a832d606af2fa1316ae1cc545995593d0796c841
z517be542b0901eaa7e0ddb253687cb584e4d192a559cd4348211a9acabbc1c989981df4942337a
z66efd084fc55cece3d873fc5fa5417ab6c9921eddcbd72b520deb3f7ece6b880ca6ef5e75d8992
zb760fc8e9d1714691caf5179e3010095303f582b65f795c12828f6baace1d38d8ceb796ef1210b
z7bbbdf49510c6e9d2b501b195671051589f9c2e848130f74abd736f9c7828c1ae8ce14ef971a3e
z898f1f4f6a322ac40b43240b043b3df1f2835492ae4309c1f3008fd413922de66cd89f961ab49a
za2188c86dc421faa1b7613e269bd7e65be4e59e8f90700e5ba129a0bf05d1535b2bf960d555111
zeb0c52a8aa2fb2e895abee1007c8ec8b6d811d07986dbc1971f92adc7dbdfeb49721426d2b97f7
z0262fda524c469fc3f66570ac71d666899e108da635841661a768edfbf855e7db15b7d816529c6
z63648a802b9392885f70bb39dd2bb45671ff5a5166cb51458e62c44aa28db6ab669d3a5dc1fcb1
z1b685adf773d057470e8dd799e2557dd6481b4881e5a547aa2fbc3540a82b36ca9687a5f436209
z1befacdb56ec77710a77891ea1053944d0ac99bdfe7a60d7222190a87a1b7af8741dc5a6c9fd40
z1a3d618cf0902f439f75696843ae1c74348f01406de495b0dd2deccd8d5173872940806f700b3d
z6fd4e3e99df0c22edaef5340ac0827e61bfb38085e1f181f096e4ebe2c90c10906aaa71fa43873
z4016d2cbb96d99dd2ff395881783149e4d1db149e3213555fa7a87dd0adae7e31d15186c5aa933
zd077628e5f66219173d15dc555abee641e03ed2f8aed04afa14e3ba518b4d81d4df0fd80ba76d7
zbc0640535083e991d32b885df49216f93175bd1bf15c6469d6853616b7f829709646434d238a27
zf6839bf9b40b310b3c08053a90aa57fb879624ff3d85f07715e550873c3913e25ffd6e77f8d0f3
z4c8002fbd1dfe84c6dc16a7a5739124c9351645758f905e004dc9d595e8f9fcd226d61c4124e8d
za76615453d2cf4be498dc0e96b1adf2fc6fd24831ad5d343dc6437ad0deffa4a8367a12354129f
zde59df17d19c6b73b9e68f08102f6ab79329bf040f28ca5d4003bda1d22d486e5709121ec6d332
z1dfc8833093658f1039562b41086da0fc555a25fc4a83594470c2ffe9deb89382b56190fe1340b
z666c9440a7df9be5a86db065274b4d40b5f5c0a6b24298c0209ef17cd5903384fa0bc5335d9059
z5e3d373739e2aa6aafc188d70878037ac83ad76cdbaaba92585d9467eae22e63da7ce1eb372c96
z2b1376e90e64eb0610221975fdfcca6f6c2d0b274591c0308dd05a423bfd892f9933f10ad21e07
z2b971d84fccbd71f191e2d52cbbeba706e35eaefa8339b39e6b642c6f655a127bfcda4c44c248a
z95ba1192c45db04ff5bc520d8be89ec6859c9be3914a910108b3258493c947856caa0f816dfa24
zef06750bf8761357093021199b1f023e251eaa1ffab2c18e4f8a69451c081d22c9c8162ba5737d
z4aac83d73b64962bd819a3ea20ecd04568fcea187ea68375bec1c7c4057d4e91453f9034eec4e4
z9b64a72a5f245f87a5ccfd0c2f37be24bd1102a19e8a0007f21a8ef4991612feb8aedecedabd91
z6e06211361d82eb6f4a677b6577365ecb239f54e769e24da3eb7f56a1f6a9923ae350534d6f5b3
z1f961dd678c6799ca64fc1253182582c875cddce9487f326353e60cf27bad4fd978b685e2112bd
z64d77b7e624d9f3305e5f43eb6ea32581bd52a7be65dcd9c5997b39a5360492d6a99763a190678
z993d6fd12b71989831a1f6204de828fab859e457019f485ab1127af4509b57570538df9f55ebba
z9d8b85c1211e2f7584d7307c7d76ffe1a26f820d9c06aa52e8774efa945caebeb23e872b2f1d35
zd325d69c0ba60a691e6a556c7b0087ccf7a4386c2b5e5d244561206f1e514b005c62255ec0c9cf
zdc14656d15d270ad695bc3506db28243b47822cd1fb60e70f74612e0a0cbae1dd1fd9eaf1f29cc
ze8a860f2d9531862a9b5c63aada9da80af6b5ce82e5fb71e6d394a9d0f623df1cc7cd0e47604b4
z3e229f49bec74d3cf59e0be99c45ca14533fa99c28e431904073adad00daed8adecb7483686d90
z12e7709a090f710a0e41a30cd0972e8613256a2d9b4e7246192cb2d35a2158a47d08d7b15e8051
z7ff63545d7e374fdc0eee3a539bed32a3c4abc8d5fc5ec2231e53cf3a0a8bec175ef13a67eb5ba
zb7b7055cc44c3d668415dd8fa4f043087e83ddd46b078943992a00ff06f53561d7a9960e63d181
zff7d8db0567456148f8553872f0e5474f1efaf2984b9005e4fb52d639c1844001314f8000e9b79
za2dadcee96fcd48c087496efc04ad21a26c338fa58c331e069b2ed9b1f86995c5b70b44523a3c5
zd8313b29cfa00f773c4e599a999b8e288266b015e2655227f5c2cc087b44ce8a1b3e6cd9f344ce
z4472e672949350df29fd7ffeaa1dd309bfdfa43ed5e38e8ad9941d32954362d68e19fcac7ed3fd
z0b8db4b8c36cca92e3baae06244e2e8aa8b8dfb6f98e09d38b22d09822fa0a9437def7126a599f
z0e34b7db317477b7f584c8bbe0090163873a6dd020c791ef56ece9e6c7c6f42568454f466f7217
z5713c0bfc7c42c26ed774e994934a1789f2a13fda0040793e85838b31fe10408fe7c785bed88bc
z5c14b53f21ba00e6c099bcfdc26f6bbb61e2de7d4154ee6fb12092988d1b760966fc04ea6ba191
z3c6214a9af9489c3ad238bfaedf5b39671bbeec410d57a85760af975274197a5bf3fbfa4d2e1a6
zda76563a4c1f0becf86f33d48a43e8eb58dea9472c2cd6028ad79f5dc1a8910817dd630cb2f0e0
z95ac645782ae2c242ccf86b1b3c1ec16abe34ab4152ecec6686cd48670608aa9a57777e32b9c75
ze9d43127639e299af56ba381b352ec5a63abeeb11045a0fda7654adb99a2e4c8ef29bb51f15b90
z46bf98c869fe55930065a742dc0dd85cec860e399d722073a681d0007963ba5f8f34eb5e70b8d1
z056348f1da3d9b03f31ba1f4b50b6e34fffda99a96ed0037868a92734053f699c88d9225401338
z2c4615313111dfcb1ff04c536826e0a967c7ae39e06228d1a6911d72ed5082de26c6096690c1e9
z3bce4aa54a1404f2caab3db1b7b47c2034b5f6c5370f49586ac95dc3c30dda349938dc6c2fdb0f
z44c3cf23a62541a15992c1f1dde896fc2c6131472c0335daa1606b5a4a47e7e102a6f1995eb3b1
za5da766a82794f17cd0449c92cda916e83b332a482fd52f2c819aa04b6b168b62df92958a16353
zf41a28bf1d4840cbca0565e90a97eb93edca681ca311358e8ba23bf231f0548e58b62f8f85aa84
zbe2612f539f74817eeb3a8566513227000d99236049de14e82a7541b5c38a55cb49720decbcd30
z9b7dd2eb6f7b287d8508865991152e8e0ae3866d284984fd294d4628d8ecdf871ac63ed67727a1
z146391451a88afbddb2549f6726ce0f3b57d63f0ac509bd5db1f29c0728e13cb9fa9f381789a76
z9f1794e0b71d01e22572b20857365f2aa88561747395737d42044b3007c0b477f3c37e6097ac35
z19b717ee9b77875fb2a440e2735f8ee52e5280771ad59bbf8629a26749bef0b9099717fe477560
z9596099ff6fd56d7496a3d2407a2e358e02203c1ac34896f329c285d2c855f15ac1d41a7e0d1e6
z99c998292fc1f0f3b53b4479138ad5304e2dc2b60d92fc2aaa3a8d2be10524df4e298bd3241b74
z7a3099e2c0d7124ae0e17ff693de2be9611cdff8ea6732e810ad949c6b6c1ec723879b1af7a762
z88999a56eaed0f6a36a7ae1027fdeb1b1e09b2979fd7671ff15c477629f34beac0f4e17af4e319
z52a028aa023376f9c0ef83c151434e8403fe222758504a1a87afbca9987476d1a4d885b227ce88
zb652e8afb7b3f4b13fe60ec3ea77c98d4bd06f31cfe97eed8c516f964104980608accd64e1a42c
za6e46e29d8c932bc711fa39f5cc9f0365714131850075b599ad03655d38334c4f3a2d18ca91b7c
zd70e98db15c67129a4eb7d5d908184c4546ec0acfc9f76d201313a23d9e03e44d1c413f6b04992
z564e8c645a1e6bd9b5d93fef365cee55cf2afbd52262014a628a05d793316e4fabf3c2d624de54
z42d0284e31961c966a0d9bd7ce9a5d6bf0bce6e99464e9721a7932050b5505d25c7e9c69f8de1a
z81ce2413d4c54f74e64021ebcb4def89f6f40f9ab812976325bbc7fec467c8f885b9596ecd1fad
z48f2d1bf0b80abafdcd2b794c4bf3cd0f7eaaea9a10e54fc83ad41299065d16d8acdba0efc7cec
z91f41e9634704c6be09c55af963e974836f998bb782778e8ff1fd5abf22daa8170b4c26739a7b2
ze70f6c7295aed9cf711cb032aad5e9eefa6b8f4efe03beedb715aa323458f5e630f8952b7d6083
z5564a9093488b048f4486ae0ad9b937cdfb81d4de2b6774a3e0a2bcd9374dd9970d663e14776bc
z09cda4e65bc1c25b140f75dca9ffd5c1501718cb7b43be5f3ed92d68133110ba0a32713d5922ff
z3ef2cf9fe8939e8f720d0424de357d856ccf34fcb878ded3069b491db1775cc4f708cdb68e3b09
z4df5cb424d0319bcdacdf8cb37ea5926c602dd9fb81b88a3ae89cf8cda9d526bfc09bb9f743431
zb2f4b4745b7b92b22c7990b67d5530c517d532bc1114a60ab0fc2d00a8952b0497996da6e6fbe5
z585dde3335da5d1c65656cc16b483fb9103a5ab0667315e730115b0ff8b194426fd7c7a6b6d1bd
za27abe1ddc1571309a900f7579a61fec50312df78e05775df0bf0f3b23c1877d71afedfe3063a5
zd7ef2fe38908dc5933ca48f69e9cbdb17e4e45a280f5ad2dba52c5c5ba56c81647e7bea7e237fd
z71b76049f8ac4788ca9c83da48b71ef6815c52089c452beee2c8d9f77b7004335383d9a97a6ddf
z49f2abe2c0cc7c02d0b5ba26c07a8f6809778539715d112e371b81fbd23d103ed8484465901e44
zf89afbbb80bce7f4a553791cd46f380f0f479b3180128f39a37d34578c77845c2ac25400a263fd
z01b3472b575cfca83073ed94e08ee6e46690e3e4818a6d180bc0eca5522e3659463aba31804b69
zd3a1b7d8b4e821d053714a0619c79cc6ddb224d136bb796b41069f9b7e56e76be1ca4ee7d70a84
ze83837244c9328f8a4c51964301b018f13a30edb73c5d9f3f732b3f16648daf0fe5b3c488a901b
zc7ce1731e715f195574d8bd9f0fef79c04d750977ad9305b42232cc9edd4604d8f7394eae0fd07
zb81264d185df6550b839340bfe1b9092bb682504a0c4be4c541a9b88ceb3cfd9d3e30542c514ff
z992ec0ddaf3b6ee5bb54b84c9d2a1aa21b957d8cf44306f84aff7fd76f7158a82781d270e0ca91
zfe2f547a883c12d47396719458b07a3084ac49bc1bdcd0de3e0141da7e8bb9343c16514c7413d8
z65a5e7f6dc42f245a628429b81b3ef3e4c1d9bf887fe5553211b63e6692ad5df47e3d14533a801
zd0c08e07cfc1ba043f67ca837fd9e41e898537d245bbf6386a146ae6a4af94db309cead5a4643c
z6b3a074d5771e2c7ffc91a9b15794abc1ccf83f12f47a0dff49b621d6ceb720190a77ce44a460b
zcca2f0b6e778edc2e887c412c933237ca60c071a55bb47f03101de42e41823efba4f661e5e6fdb
zad25f22f12fba2e04f884dbd1dc9c1baf498c65ce6dd699bae77432a21ff4b9ff27c0ffbd27edb
z33641435b809b34e1b68042b33ce87493d60d8fbd7e7940cb5439172b6440bd1f75bb21d8bc183
zba083e202ffaad6a03b68bb9942c93fc0b28ea14bd5e86ea68b6b67389f783de53669931df87c6
z34a00594e8e4a839530f0b57f567b1be884a9bfebd284223102a116c816365e1b41ce7bc9f2014
z4e54897b027eebc8b04b2aff26004ce33061540c19224351a1caa2d255899e6e8aa8754630b2f6
z4dae1a0182240b97996e4e669bdccb5aea21daffec4b640875c31fab5009b823cf68540e2860e5
z90d848bd1b5da3049e8b2b277180665d638712c5692d0938225d773752ab2720d841987256f4bf
zb4dd1dcc3add3a19170e6855592b89507727fac2cdbc764bd28175993896bd954b47b3aa7f0e8e
z6c4c13208bdca28d085eb18ffc1f13052ec96f1024dea041f382c26f9f5cb0459b3080e7e6c0dd
z25430c20ea19d526529b1d66cc18461566ccf11511bd7c1816de1c49b54201caa347b6b956634e
zc7f90e01aaa0a9c8a2e37e8ed0efa2018deea78b8bb4b3b94e5546ab84201ee6bba081737157eb
zc23a4f3e5adca637d32100e296331c118f25ef4348c6d6e96a74fdfeceac74cb97b8ecea0c994b
z561b7074dadfe571b53ba50d8eb3d9caa4f4d29e05909c98065954683ba32db8f5af145a219221
z9b0affc78499ce23918421cbf32cf4452a18130ba615d7a968c4d147fd8d7a6550ae40067848aa
zb7b6e46d158e402ec13b88a33d9cdcc38382d18939a21c8a0b4cbbdda0fbff4ab38d9f22a200b5
ze771a775475e86c08e465cda006293f402d9c64566cb08ce03b287775143edee03b005871f7b63
z1708f7cbb5afde3f604f5682cba4b7a58b99e0f0567f68519d3ff84cbc5405290383ceaeb7fc34
z73cb5f06483c887781a23cb19a925618e00e4fe50b21be32b78bf5d4ee4b129da851db1288ba10
z203cbc4feab7ecf7bce92f14747445544b9a0c0066f228b923392c4ec9edf1b79e8984e0da8162
za2258587d9fa368c5c2abb5dc2476ad48aa4032bb8ba9eb6093ffceb92cc98a6b7d60e2ce02daa
zaf76e34557f3cfdef96c3ab9abfe96b0c7caf7de84b82636da9760e8d9332f957d7399d686e50d
z47b312e68a5caf1fcd274e33d1fb7f166dc201c25ad8785533cb8375bf4fcdba4d1fe2d9ef4cd9
z46ea66c7ee281ecbd9f46fb13bf72dbbe7b3bade4ff9c0010650f6b5fe4ebf5333bd83001d09df
z5524f45fb6a78c4cea7806556630deb4b655ff5f5ef48721163b2f928f955b8477c4eab6817d37
z10ea957376f9330055bb7833d02c5d708df7428f5918381082cbde1797131139f1ec2eb4f1fcd8
z44deca249f3476562bb3f06f5531acf5436f34405842b9369dcc712f645110173427ad2f1a8297
ze35a6e940a85f61c67648ca6479803cc27cab35ecbf37b1f8ab46d59eb8d7ca596416b05098171
zc40e634ea58f5ffb98d71d983e7f230a767d3d7006a1562871afbd66e659927f21bbb477d03078
z3f857436b2358a985640e1920db9ee81d1eb3e80127ce55f090917ea3a3fcf511f68e0150b29f6
zb41e187f1bd61f8622d62c979cd5a18c8964c4d5656355e4953cd095ca786dda4665728f591eb0
z67c1c31a3268cc8003354579eba0fb8bcbe4c762eeecac501afa30444e2f12d21e6d63c021771a
z20b6c3f90405da434d802d6ba6c887fcc3ff46d79e0780fee8c3114a94a23735636fa62436d5f4
z058a26098703a672ca3124dc61bbdd8072e67e3e976cc8349bf4c4e119c472357160b350d9adb8
z278a132fabd2ab882adb0da46c98f1e075c4517f669d69e70fbc2afe9e2a41ec313985bef3abed
ze79b6de800b87a8ba7797fae94cc88d4cfaeb2f9b13553ac7478943570536f23f4d6c8fccd8f2c
ze297499dcc7e9508c5d336520ef58c288120b350a9c56a8da38db9b70fa79789b053021c1c465b
zebab6415e9b017fb583b7beb30881bf8e286bb26ed4e034aa42325dc0f0277b37f8033a32c76dc
z0541b677a4ffb2e238f322c328d1a26e04bae2ab7af3bdecfec30985870c12271fc179f3ec3d8b
zc7599b99dd616d196c2caa507f80e18a13a0c1a1c11df23822f53a9e6748b7a1445a80d283a44c
za193807308e537d1453d4a70b1c552610d98d5057ecbf8ed1364e56ca56d13fb944ea9b533b55b
z6db060c5d5381d8ed60f43bbd6a6523212da3ec28c99d8b4aa038c819569e5488277ebb81197ff
z577b536af6d749f37d01b8a44549a45a231d2c2e9a577e1f7cb14d3a449c08edf2df1bcf16ea06
zf00f6668c05c14647bfbc92582da73eaa484a235367e8b6724122b350ad456619a508057cb09a7
z2f7784e0b64c23d11057fa2b75e7d7e261513c6aeeab7332bfcc399b834f15e6eb6ae2d837d93e
zf876a1b53699d47173dfa1933eaa611f0ba1e1a19e0063dd844a6e22bb3ad2515f6ff661076a55
z6ee5aa16ad17b2efae88ea36f57c87e8418e547e0fdfab9777055ca134ca8bf480dd4d5c0cd16a
z5ac9a9e9340140336c244666174c0e1dfe445cb7afecc4f2b45ebe5f96024f7d77d025c93b13f2
zc5f0e79f972f674971cc14e89ef0aaf6256d52e9997e8a7c1b5a1c540deea03d2ed3540c4377bd
z37c706ba5c97b5a63968e50a2489b4456668f16bce17096b0e791541af342a406463b4f0ca599f
z8022376aa7c28404280b2c95c6d57064228b58ee331d551836cdc764225d5270fd124606f43a5e
z895cfe9f118eda1c0aa4c9a39d95803f304825b0ee8eeeb89ced1f7954e8b238f9f2da85aa13ee
z16bedf33c849c5a14265bd01f6332244f22ac8014ba480ed9eb457f7dd2e0f477cf8271bcb2424
z43c42c3817af5625953766fb28ea4a69df4053b902fceb3339dc66c3b922320afb977dc728cfb7
z95fc41b7278f4855882937ed5ba1cd2855d76fe6adb56dd7f12616eaa069ceb414fd22fe4a75d2
z3043d8e63e017c3a8b88a6de5072ba5bd06012d58766993bfc9da5dcf9431c72da88009bd57b2d
z835a13044b099e9f066c43f1799ab742ae1675daaadcb6f4e6e74ab87eba73684730deee7999a7
z89f94a6393e571bffd2bbb21025cc70af4ddeca88125bc2fd213ad298282927ecee0574561efd2
zab26e71ca9e4b7d1c1de747e194dc0e1d3d0ef017ab9926586fd79b27bd1d551b9aa28d095822d
z5e22a7b57546622d17bf79fda3347b1c6704751ac7334275fe20c937cd2d6e528e44d4811770f6
z2eb546fed67882242d54c8f8c47c2f9a9bdae6c8fda0057186d7d286595107cf88462f05e357ca
zcaaf83acfc79f77ee6c33a56e7a9b0a63f4cedc00db42f56d31ccad83efa82217cd27f033acaed
z201d05571ac00350140513ef7cf60863917b92db2962ee9188973734eaf1107cf29a7314230cd6
zc59556699c3946f42d3909ab1a2c28213e06791a00ea4219910c263bea8f8f2cb1ea4020f1294f
zd3617f42f80388d18cb90b88592af1b3b537b80ad67ce6bfc1305a423f185255d2f66ee3b0a896
zcb5a20f84e75addfe958c792747585bab981b4a0065de2f46c93e26d5925bf7fc0af7b32b947e0
zc0adbee0f5cb9e40d5f69a7899f01c2841903855165abf8b895172ff46cd01b7a203b11148b52c
z9ca2b4860a54022da70dd66e9dcbfffdfce8fe07a585c9f5b24b505364794797216fd2c8b45531
zc454a56e2a8bfe3d0982823e0df0a0aeff07a91466e032bbff4fc4c74f73733fb7ac110cbc48de
z88611aa0eb08f51fe1985fc3ffd8cc1e8f9071a43cc751bdc4b82aef01e496cc84d680965949d5
z24ae2594a40e75f73bde5124f34d667de692484b5351bc98b0b9de65877bf420162cc02274644d
za3fd6b97471ed4459806563b272a5eddffa221c223315ae501175f8f668d3204e1e8c1c9b6d6fb
zccacde7facc53c4dfe205b1b83683970eb01ec3f88a4af4a3ce354638c9eb61953711ddfc16059
z82c29087f27dac1f3dbadaa558202514c88e47145e58976638968263416e3286e350bf8335e13b
zeeb3d4880a66a5d9bdb71962157c02184700375426913250d8526b3c84e4d75c309f28c7c1a97a
z947794c12e99cd14396955efc4dec4db03f9dc1b030ca7fc6ef6965cc68d0c8bfec9570a89ec24
z1377a6133aa3b38c8920f6ad02fbe618c25654da502408a141c83b6a7123a23e7a74f4961a5370
zc178c949e8a385e17b34b436ce083d4c5f3194a7388695f7c0b8c357635387784b9a3bf2b6d5ba
ze935701a7e4b734e82ae7eb8b33d359c45c8624f569f8e4406c7893a6bd095ffcda54b31953c86
z7ca79b2844d7f304c540b5915465971070012fed8fedad63bc63578ab06a39eb2040da48a720cb
zba554d9a6963af25b5449c62f08a23277b44b58fdf9fe0b7f80e0ac369e0ddba5255ef3bb19052
zd8162182bddc69b2f7c8da6e2ae1f458438c13d6c3eba7066a1ab2dbd6f79e4d951d31164dac70
z37d4c1f3af961f0d3f58f016a30b76756068a3b212a2149c105bc34ce05c8ae0ff138315ea16a6
zdf74e2d55d5297fb6694c8e0791cef667f8ba69fad55d3da190ba07cb5e926c2ad48df9707d940
zb2481bfa53d16afb3cd7714dbb78e25bca493721a748a75b549c51b80def99370d8fb8f2121646
z40d81d564196fbaa97eb4c62410818d676fbf2f61f379bb00302568ffef6c0e66be897ef071de6
zb278c95737db8b7b7fa7585d212c700e9252ef9d45c6b44d95222049dd1681959a42bea7997f22
z7728dd88d2d5feeca4930c7ff33e45f3ce981ed294fbdf2e7cba0a6402fad162f4b887c081998d
z35a2d9aa86be9ffa6c6e4d83700942d051c4ffd0898dd85137ec2c50bcff883bae5699c7306ed0
z682a90ddcaba3348da15027b3050705df91c945dcfe7a7f0d6fb41e5a7779967f4e1e9f1911337
z04f37f8a1a987fe3d1af4e8e293450f355f6f6b4a0f12f51f2d26483fbb957a530845cab4ed77a
z586dff0d97820372a541ca9d2e01728cddaac996d11aa8071e201603fa8e425521a1f2c57f9529
za483bfaea702247a53027ce18d17c4fb0de7280833d49cd92755acf829f2192e5ac9ac043c5c10
ze6afbfae1363b454cf6ac914a7bd6f89623768c8a770c6dc113ff3686e53313db02caee895076d
z1389cb4fac9ef8d393e891e02e299615f0e0cb9995d59aa208ef947475e17c3908a9d080971586
z21b81da38bc010cbd8b99e98412341a6468bd5b4f791acc885ea1263d8f12658c29e975078ae5e
zfe35409bea5f413d37d6100dfe3e0cd34bb0dc31dac96c83aa7225c3f11389897c96a2903c4e9f
z786f0f61cd7ea3fa1ec4f87af3ce6a2f0db9c542ee85482ab26c5eda4648b09c86f21c1075caa5
z6c808b18758e70925076b71a160429e27980a002d68d10413777b6e885217cf6bc102f67bf19e3
z81f62be545eab132b1d8de0a838e8b5cabd011bc87449b140dd36f72cb194739d432667457a959
z5f1132cf83fdb37b8fc93b974ea930ed10009385e31ddea5c8b83d84783efab48eae1ddcf93077
z7bb1dbcdc55822baba646df44702746a094ae4a28495e116650b86ac6b4d17811209e5d5170439
z87c1e82b28d365fbb44f60cb23462d8c4c59a6c00232f030009b3e71999fb4fb7913e50987cc9e
zbdedb075fe85dbef2ac0f27b2169c2c755219c696c4af1e7ad44ab2efb399a11ece6b2a8a53274
z1c345e2ebf602bbb2c3fd61532846b14fc93a8db51b237a46bd5b9bee7f6116e43095986dfe4a9
z868aa6558423eee27373a4baacf16ef4cb17155a4bb7ac278af9bfa00073b5239fed3275721b2b
z0a00096b1bba08733c72230f64d7f1932a8589c236f1e5197a1064da137a9671db7399b9c525bf
za8d94ccd217cd63a96184a749d7b7479dfbf121ae8c719635043327788c031a0708ff3b628aa41
zb3c8c2f953e4201b20c646bc8ae69d663c960e8a9e44a9d1fe93ce169bce6416163591e91fc480
z595f80fdab09ff3f9abe6587915abefca399d53580025761fb512ca85f5ffcd11529ab71b7f472
z1e3bab06fac85435667dcaa612178c63c55a2e2e0a6ab1c9c108cef510b2f96f511c78cf9c6e57
z283e52ee5faf29093145c752547951d714b19eb77550235d38126f725b15437bf661a78a2a4e2e
z9ec5382245182c75a8f9073cf60d8571a0ef9bafbc289a568368aa4a92896a37aced8f93fc9ba4
z9558a22995cda1d2e9e62fa707e84c476e860160928d2ef1916458de697d82fd79e3c43846641a
zc075464009575a238941042f965233fbe93ccfff4f23fc2a6618afc66d8c8a73db3df92e0aecea
z22a9406025bac4fc308c4b0f2eb34ad2c1a308d0b403ffb48abd5f86e5dcd64d544086f2e96875
z0eafbbd789e9f4b959bf24a8ea461f915f64fb4acc2b0c744a30b46d42b78532254fe18a04d795
zb1176311814fb1048b055581f8b0de1b06c1511bd459e1605d6a590641dd6f5a3319439ffc9de8
z94772d84bbebc04b344c9f5959e929fbc81867165fff4ab353dd9f289669c17786ed0f59cf613d
ze1811d5bd689616a11294bca67f493bbebccef5b2bebdd97857d7501f0f0fffd4f66f202c8c30d
zfa90019343112e53837d404f437986f5ca1290308a6f481e712c6544cdccd02e6eff8311d5f130
z192286127f02ef3a388f20acf115f8f6b718975b9a61b6a7e3b47a7593d0fba02ecd4542b3b1d7
zf6b5c592b023ea7372a6f5a1983d0ead9b29b802331e7df6533844ff32320b33a5ce47311a75e0
z2568dc692d5761966e3d06015e381c55bc767815152557d9006284a6f4bc8d291e9400fd444511
zc29347e31467eb9bb9789156b75cf4c75cd9d98a2a51ceea695539efeda431c458dc29c87c749d
z0610e814fc7f2fc291493c9465568b85e619c49340b4ace58b34d41684cfbf8c03d4ff84dcc487
zc3efa4ec591cddbe9327e20476fbb00f83be17c72c6c92f632102fd5ce7a665f04a9ffce7068de
za7028663c37da45c1fbea331fd907d9b60eae84237318728874fc1ec0c0ce2741dffb2c20f3acb
z8561232dc03cbbd22a2100e801cc62ca24a08712abd6f2d1ffff6319cfbc093bfde0dc68be307d
z081b3d257c59c0787de594782e8c6d7db52c12b13443810d28269f0665fc4fd89f65a0283e3902
zdc827d0292c728db9161f39f485cd5895e72dbefb7de6ecee0b98edab5639f3fe2b2feb59d3bd6
zf5f7aa6a64468ee03463f549c1b0a265f09b268b47977a30522b5d9060c7f593e0e991f58d71c1
z1db27199980517dcd9c1688efe0fcb9fb5d7a196a0f3b316139a50fb8d430c2b9bd90ef38f3c36
z67d9db9db07f55df34092c10cd36b0b4440964b9fef29efee493154f9419a1c465e1f9fad6746e
zddd6c661a7b1f5ea22b59852539cb5b5dfbe094586d4919fd38e4b28d8a9e5a5a69e390c39f8ae
z6d6acd3120f27de6cf9c3c11112ad796a9d507ab078cf92ba245bf88361b11b932cf5e8616d0be
z7bab9971d8e5fb05a23cbc96f6922b77ddeb911e43a540bedff03d0413ceeaf6d2a0c1b7fc9efc
z92a5717f5a307bacb8dc923958eef134b4ddb53a9d1c36c3bb65cd61f83a9fa96a00c375cabbd4
zb13015f142204ebe768328e29e2d8a3147817253d4db18c4e68012dda693c552a81c7ef12c6898
z2ace5fdcd14b73edeb780f28e14d8371bacafae7e2b7a93bc0acf958669ca7143c9ff3ad6f9834
za6064b242640b8029720573afaeabd55feb08a0333f0274e6caa682c6cadf59f210c77c5770bb9
z6e2397e2d2ec16a88fdf996fb301b95eeab62e54d7171e83eaba8e5176d9412d3b61bba43fb034
zc702269619f4205258b4484ad9e132e448af654935eeb3e1c7895e986bb8e23c221660c257babe
z68fd086656c21f8791863bd3d5e13f4a25ce55d28c5a606c133af910f1e3d313c576ee35c44876
z03db8d939645192a08d6bbd44b09e1710dadfb13eadfde1083b3088fe6c13efb331c0cef8d0582
z5bd3ecce687fd2499c21ff89a56c8d9c5dc8a293c954029e4ac78ee41e6d9a9bad351dfbc944f2
z99f6a2f1cf2e40f5f55f33ef52eb36fcf393e15227e6e34ad791759cd0463724e5437fb1a47ad2
z11cad01f3b301db4e5b82ff5d75b64f0634ac1a0b3a8eaa22f0653e609595830ec0a2a1db723d3
zafe3df87e8b18f8c0bab92b520077961c3a1445f29bd4e3abae4ca525ebc65198bc90aa8d2eea7
z7b4b2e2899ed7ec69a6eddb90e2aeae95571a5ea6ea5674fb4b54821064079a43774bf6c6be2cb
z8208c4d3fa213ac7bab2c1b9cca77ff2d608d5943e8545dc457aebc5fe3236d014122f7c0bdf11
z5f17821688940c0b95249b2a55d093acdca4a4a66604160042d91b0079f1f23c9c95a962ec63b6
zc1cc1920114cff6ebdeae80cba7aac284df45b4381e989b5b6bd6f66ed3a5a6d985afe297ca542
zb60b22be1aefc2869216a24f748249411f7532e9c032d18a6832556202c8582d651af6d4ba999d
zd6d2c6c02c500f22dc4e34a09e2955bfec1c4087f5bd063bac8255ab1a2ea299918f13425e0aa4
ze20535be4af6ebae675a8a44ba5cf0694b133d51d047d9b5ca8e523a7fc25f7d2053712c8ac5ed
za0b8e09adadaedb15742dcfb62fe0002b59dcb71997279ea0bbb8c546ee76719e22eeb1ae762b2
z397f47216f743a0eeb6a27341c4e4c8398eeb97742eb3f2e8db9fc13a494cdb1e3a38e5f4cc784
z2a329c440d0b78e94d1a923aa958764559e120797251e84ae6e908714d72f467e51e762d2d7e62
zba247c56c92b13fea0c9c81cb6ab5deb86100184f0d12b9a09f72e487753c9a0b326330c8388d8
zfaf6cdd7fae45a66935a6bd49b21edf99c8ad0c74497023401fd4a495ccdc95cd1342768d6a214
z4e4d675d555ce189087b343b99d06797c0c50855136fe6d7e0ead4f765c837feab221e066503af
zc6f37b5679bdae7c14dc0945bd39b8408073676613348d21ee5ec069cfe6bd05155f7c1106cb37
z3b403a041641dca1f637746cf7c745f737631d03b8bce8c5555ca703317e614d87bd0946c5bb5c
zc18cad6de89b35aa8ae3132c9071abcc36b6f62b94a75ae904d4b73b479fa77ec9a07dac9cd6a3
z9a37a8d3c76c45fc03648b24facccdbc5dbd69cfd030e6770083f7db22a2fb1461a02d92695197
z96779c6119b277f9ba1a329882792a7ed6b3dbeab9bd1144dd60bdbc009428bc540ff4a3da513c
z40d85afe7c6397237b486fa4180b4bb928aef9fcb091a3234ca05948f178fcd452d68438426b5c
z036549a0ad48f9e0c08bd3e8b2da437f06d1b83a1a62d06d40b926bae7903afb2c499b0bf76949
zf00c5f4cd1824c33592e3a759b58071f256d3bf9f0c225c484b089fa3d325bf0da9aad43ab5413
z4902c5e65ab2d75f612056c7db8552a181f34fc6f1887796b84f9d58e7b38fcc8db90bf4f8483d
zd657947896e90293af94402c28516c3e105962f2e19d97042c0a1a03ebf144a47e0e97a56fef81
zd8fc4f41d084b33c2c1ed0d77b725186faf9143a530b2ecc0d356ef64574b096065e911e2af251
z7d53fbb7fafc16f75101fecd67000a1361ddd6f24441097a913c606860fd31ee6bb66c0f5cd1e0
z1bd38b149988546f6ed0fa1f00ad54dc6eb78ba9836e9cacbc125cfaefb9040d261294bdd64bbf
z51dbccf25636e9fb6495ed12168cfb037c787ac2e6f5e6ce43f16c9c510dcbd63c27e3b6c4b8bc
zcaa0332413529710c8c2ee6baeb2f01059c9415685c28b20a9b8aba31e9bf1c76c5a0390d1a1f9
z63a5549ade281ab4a198a950872e8bad4ea8a66eb1974d39940d5d835948fab2f9dbcafd6ba12e
z6ea25d4666d33e725e2230f355f3245785126c442a0ea3df660efbce22b94a7a807231d1acee2c
zc62e81d96a33cba1a1890ba39ea05a776ee07996b0fb8f1ae56a4ba9872109797321d8879eafb0
zfa15d33d8ad50b87690eafffc35f950f18f89fc2650ef5237b0fa7ebb7286934048ccf5e78ccd2
z34d578d35c2d6e1fb55b6ba5d24d049d546d204e6cf1c6af78554cd6be351e57a679e88b0e6cb7
z3786811b646a5db1c6429a5a251c092a5674e1359a80ff271b3e60f81c57d5be93678cd4833998
zd27a5c5d49f4c8fdad12a13e5210a507078e4d7f0f1dfb18d7cd6df89f7409c6709f99a94b784b
z49986dd02f838701f62957ffcf9f281de4d24b6a038700d2d3b85b4a63f50fc7bd3ca8d1fa9ed7
zaaaad396f2cde307354828bfc90bbff090611c7c45f08cffd3a8ef48516ceaa2715f4de9eedf6e
z1ad23bd51fcbfdd8d5bb1213bbf9a192788014b657ad67560717eaa7acbdf9544d18e4abf673ed
zcb553cd0c5ec80e7a5d3001d33c67fb24ad579738432d612c9375069af6433dca30a1f8be9faf6
z161bd58276b314daa227f6d6a5d47292a39ac81988cc72e692fb3b4c7b61fcc2869c7dd05943d8
z1f1de1dec6efc92f71754140aa923f56b48ae569938a0cd84368a2e16b9bafb28ebd343b344e46
z4e3ca8a0427c93347170ab9bda30009a243020cb6543f9157cc9558bae38b26bb436e26ebc85bd
z51a9fe621f9e2f1ce82fb6e5d17f6952e8e2c7e5f6287a107772ff7f4516588460c6684531d341
z729ecc734f334a0dc2586d38213e38293a0ca84dc3ef04e40830038d9b61493a269c7883ca8927
zc3305ef4ce32095485413e814da4c6c7166c3e27fd31b762bbaa33cd9eb3bc60a5086b1ebe963b
z9f21d169cda0a9ff3d5978ddb374c7885c0fc470c3e655dc8c16343e22c5ebfa745715769515d4
zf47b421134e20ffbb7047c3c3a53bd785c5da070a5c3456cc22e8d63cf16229fcbbdfdfe3250ff
zca586a2a182dcdd08aa0d331053392b1113c37d054f80df9ddd9f235e30f5609b8a0cdcaf34f0d
zc9098c2cb2dcfda429d3b002bf22e318298955f099243de99bfec4666c73efc13c0368f1857ff1
zc6f5652f5d52c95b0f99428619dd66fefa4c5a4c545af559f2b586fee9f31c570198194f459ac6
z07b52a1b8b1011fba67293fcd58b3a8978b4b0f40642f5d7f7801f95a44c7cbbfa46393e592409
z1145a82efbb4a026b806323003d0c949935c0d317c136933917fe01da3bde4122ee307cb948e7b
z4601d13f2f88e3aacb55f8700601f906259296d4d7a7d48bdeaef5fddfed7ab36cea0f235919e4
z05bbb1c4a60554b369aa40482db8050a7094a44153bbda1887d775f3e67d9ccc483b43671e7294
z206c5727cb9e28da7c1c3be2fe0d0346a8a02b824bcc22f35c49414fdbbf30ca9ef0de34ddac47
z4f0f753b8d01510f1356b8ee746d81a886d32dc2ad271a1164a66d45de26a80d0d91058733f04e
z30cfe1ec2af2207fe022ba29eb024bae74fe0a2d9b7b95f142f911361c10dc740e84a6032402d7
ze49a443b059b3c67fc15d274ae2138ad446612fb0c989b2fbb16bb7d07b51cc7cdd7523073bffe
z4287654501d5241850e4ffa79eba34ccf8d113b9321cae80922b4e0ee4d2c747cd247993120168
z940fe407d9327554ebad468d99f53a0dc1b3a0162034bc8fc5750ecd5211e1a93b901ce9612299
z635606234d36488288c33d60f1c75086aa111d023f1b7f11e090e0ac648b4719466f5a5b826fbb
z6b04b1c5dc70c018edb21b0f168221c223d006561bb1d3fe60fbc22df31831388ac60236c1c9aa
ze7a53d0c6fcf7355a35086407cbf40be6eb99d401443242b869900e47f575e5379ddb4d5f24d0c
z1a000edea56b2f5ff46a19088edcd92afec98f763be743fca3f1c45c0289ae787c64826b360009
zf46f64179cc300540973f0d3fc7ff253e9f70db22e911eae8a3e0b29634c56e32180ee35710bff
zaba7ab1f1614b713726642be89c7bcafcea8d51d7d188216b914f338b06dbd6d320b39d961af48
z0a81d7f879fd99cadcabb11caa662820a376275bb8ec3ff5d78c4049f7c0eeb5c5ebfcc252c12b
zbf39260327552552b276bdbe7268a8e627192b475a37153885cce5447ffb3fa8660406ac7f9c93
z83d5282523199ad788a60c640da3296ace93dbe12382e10e286a6461cb4fa8f451f1ea76a07851
z74d9531417e7f74c42317dabdacde9ebf4522e2cec12f842d4e2872e8675964d64263d08ffdb06
z6fade136a777395a19a8268a4874b498729d34dd1d7b1cd229adab1db8ac42a04a7446ff79895f
zb3517eab8fe7d4957a2394320831f12fc759fa8be0485a3016233c3065d0dc7484f6cba3583116
z2fbbd76ba14551481686f04946756db6b58c5ace561cde4fbf1dfa1069998c8b1ec9c80ce1e1ae
za63a584f458121ee743b6449789f3afd69e01a25d9d67336c84f8deab106cf42e8883c57977fa5
z6eee9b63e454adee177fad5d3e846e4b54a6a30b42f22bbb5f5d2f790e9b52c9c43c7e67113249
z318d29eb8ce5e72cd2295a698a209ace95a3497f7a36495b0560d49c9e003d407445d5ea500026
zb0e1310091d44384fac0b0c257c253a1ffad37f71bc17ee51b333f0cc0544f39edfd619f0641bb
zd44cef36ad9b5087beb7bcb95e3d1f21a2ac8cdff981980578c134477cf9f099e6f5e042f2bfdb
zbfa123374cc64762a8f83816e979e62acc8e28aa034df1efe4d0016b89f475a70d33402634401f
z9fd1aa0109dee63f13816b25afad2b31a6acbbea926175ae58d285e1966bacdd591e8a30eac355
z99f35c3904e39d8246fdb6f3c668cc35cc933e59e07c48145aacd273e52194708da81637f72b30
zbb4bcb6b7f28385b6e99cb62ea376e6fcb6dc166bdebe8904acfa04c13ddfb8737eae695203f20
zcb76881088f4e5aae0eced85b3287963ad6ce00c41c23b414692985f80a678763c446d93945843
z47b7382e4c445f09ffd4a8cccd29f6639bc724e44606ab72ac478de9fae914fe34c4d25aeb2e81
ze5af7f40e7fe0d23e9ca2d7be612157cd9157b71c887aaf2f682602c3f2a49ac93208fcbe5a3af
z49daeb5d163555405736848e3303527b77dd3770ae5d49b37c27d3a1ca5cd32174a7f9cc086731
z84b9b3d9425b7f96bcd950dd9d1e6cfd5e259a027b059b28e6b671cb6d22f428480b73c5139127
z26a1bb09fd49d1c7089f344227054d62ae6d489e40c6e3705f4504d4f0b7d2ff25b0247be3b1c7
z4a407eb8fb46bce00e3be1a137357315a077862bb59adb5636a70e8aa5524b04c29c04e95581be
z32393fe998f28862f810ecf9de7c5f391a1df71f60882e4ba73fa0c8e724ffa189b2b0721c62f6
z1eac906030dedc4bd7bd3d8a36f2a2c2eed49fe8b885a5cad520de050edca12c664aaeb17ea52c
z99a47afe38cefa7fb69c954cf35d34ef9393c4967f2a7ae1a9d573e980688c853b35b0f8b7479b
zb59bd8a091147c3046c96c9e3f339301c1206a1e90497650bf8d2a72124ea829e7f1d5698e6183
zdefdfd61d877634b9331d21d6e293ee4dfc2e447f232a411904bc11e03143f581ba22aa1324343
zfedf469c2217cef3ba21967068d85d15c1927d6c8c85b3351b8182379ab84f54611cbf5e6c51f4
z31da38545b5ec8de2b187ebc5e5eacc55425b41c3081df5d401d258d0af2f55777927a611881a0
z81c79ba5a2f94fde02865f15c8e63bc9224fe3a759fbb7bfa3c1459346e8b4e7abe311a47a264a
z7ed33e7bafa878edce40172cb0435e8e435010fba675032ed35e5005326c0f819e24da935c147c
z210711e9ca0387971ec27718ae44b70648b87b03bcdab2a7cc79c4f5231a7edc5ffbbb63c5b68b
z8fe30c1bad7ceee2ee736cf9f7b582608aa7475ac99d261bbd7a79386e20ae39a0720f3e09dd7f
zd5c234bdf14428d21cffce1f8e6c2fe720f273b2e68f339ff9c8dd8c6ce91de78e887c09dcc2b4
zafba428ae12ef855b37cd90a3e28253092f642d93f9d4314c7470737a3da21631dee1ffdd9e90f
z582a1507518de565bbad8f0a130b706ace9b2bd3252144266acf688ce83024617e57a587c16355
zf8f15613c1f96375b48b6abd0a0c84af9b8827c633fa55b9b39aa3316f55958f0196b517d21198
zd13fe41686caabb040f3a75a3506831a97eaabe667ab4add5f8aa645ece3b9740959bc01de9aa2
z1ffa865854cc68f4c7a617f2ada71f68c2aa32252b9f31237b3338b2279de0f62eabfbdd9010ce
z513fc94ea5a2dc3f91e336c8d4f84b7babae1b6871d26aeb256ed4e1d280b444567cad9b5fb723
z1c753998be3d8e0932bf93229b64f56f22673f739b2d03734dd10a6fa1cd0bb4eeb9a00bfe29b2
z25b58c24ea1685865a1d85c6e5b51bee7c5d7d8b93f21c2da38eb8b7b54444d6a429b7d53e3b36
z55cd5ef5e96181903526055e65fc52706ef7fbcbaf801f5801edd7ce3a64c2174ca74e238bc92f
z8f37cba8355d8e400dc929469d2ed9b0cc03741c68bb624f99236c8fe6e3846a694a2fd13f0c95
z5f6e1a356f718ba65348c861785165d480305d722d1cb6c94bd38f05912221d908fdd4b61ee14a
z0a4ad81134441f02cf4769888759f99197c993ec205b9c4f9cae7fc308280df4ba0cdbc54f5bfe
z0b11a1cd7606b4aa5aca2bf54d9d759c99d748741ec2ba9eb4a4306aea3147cb23ce906e36a96a
ze9d3114d06455df9bcd3cf1c2c3e694ca9b23ecfa163db6ce597c716eae8c99bc1ebf34eb8bcb1
zc34e0282cd1aaa0d50cc01079f6222625ce36005878573f5e5421ddd1f33f74afec7f3ae09281f
z56d4f135ce1e526f4616871f1a2b653c3889b17e6a77a0cb11606f385bb3467d6d7172d404e1f6
z33cca46d2397591f018960e1c4826adde4dbb253d5ce2a42ebc4e1c9cb03a7f137523cdeabcba9
z0cba1ef39b607da8fe8b4681cac8ede75e8c3aeef6f5817c795a27b90b778b4c216173decb7ba0
z1ffd6d8bdf0ce0361e3d60894b02e917aad47b973f8a04043566d7d268096ef4e9db331f8b687e
ze4c7aa36b98c1c77c0ae1d6647cd843c36ff8032d8c5d09001b937ab4be54e7a985a41d6aad267
z4c634ee60e52d4e11f19cbcdd4bd9ee4b2ccf26a7e0902e00f32667cf34b39f42ed344876ce576
z2dac18067f90c6da1b3199908f331795026197390b6fddeee9af89b9ec1100ee1dd86d3289f1bb
z70038de5c5eb7ad9fc998a1d1592c005168dcc955f4e6add562fb2607119629599b04255ec4aa1
z68ec6844ffad5e9862506625308f11ca6e0ec1d8312b59b077d5198b44aff4af32818a9f5a00c6
z4b65f580d425a8aa0cfe3f4889bfa30a896f6590fbfdd5cde967089841cd438e9d07014436a882
z0f0f4e9982fe38aea4d3c7555fb77f4557c852e7e576f795329c1ff8566c29ff6f983b3eecc7dd
z46fb7589d5ab471624e31f5b6bf5e948e3099d0c9c916e725b17d398c243eb72ab11a46576d96c
zf846e750367be09e23d295e4d12a66166a93c0bad8fe97b91705011bd1953647f33f186b81827c
z4bf98fcb70120b1dc74c88912fc38d39891b385cfc1bf6691f8812a04161367d89800febe7398b
z9c6710ca130ae2e36df7a84a76c40f277bc1753af0febf943d2026198dd3168c5c0b9b2606726e
z2a95df2d1c41254c336d6997f893dccc9700d4821eb75f983b0299e426e052b83d98eb9fbb0388
z8ddbe062ad5773723ad7f54c8a64de13d413081cf4bb7ea37e26e7f90864735a25e2c2f334d270
zd93aae516e5e3352aef2010eb4e88abe9707d3855229d89c77a1a1009872e978470995fa52e9f0
zb7f4db281c6c797c9ad1bf96af81bcf3c5d3150b120e32583c43af48ba05d16b873ac577df85c2
za5d853906867c7be59906c7bffcff7f998964bdfc7ba45747018e15b6f151aec3b1dfea6aae3d0
zdd424eeeaa8919e6a34a8a27d59909f31bf7c79dac6bcb14e0b14bf36cc2717803107a3c38f0d4
ze901e4684a74984abd3b081806769e91cd0ce77c2bdec6334a0fd199c46fb6337b59142604dd1e
z76ab25b653cf94b65a028e654cddfe90fc34489b5f179419760c02bf603404394377529d680f62
ze5500fde56de664ad3360ae89697d12770a8086203b41f9c19f40ca53d2f3b1c5b277db27f554e
zd72f25215a8d475de90036fa8eace5019f9e87f38dafcca917d6fb616b9d86fcea7bb6fa6833b3
z1bdfbeaa64edfd0b81d393e348763b5f221143cc9184fc59c9ce88afa9bcb34036d2eea7d09225
z671fed5255264d2e16997004251b94678977f82723b3f3fceabb5b1dfdf53fffb9eb7dd48c9348
z85a4718ac321222e4d1bbf5a56b60450f0cd6b2b0565dd2a40c206df6a8f55dfd2fb3e86a04899
z1dab18b13e33c747c71f8263259cb12871fc7d5736587183fedc686c864c0451e49b367479d8fb
zde9a8a158b33bbd1e4f7fa2b01faa79c0dfcfd5331294515fcc239177ac79c07f8c9c16e5d7110
z0a89012514939219c274fc5029ff927a983f0bfb93046c4e48786414becda28088f731d9f4a67e
z855f03f7d06e4ff8c6ad164fa3545c45676a90b0ff96fa83e054e7b4f087d5cdcab9e9c7552808
z0218ca74f148c202891878138d18b197cf0ca2059d617cca45fb16d70c372e44cf943e40c5bc75
z80175425b3e8f199dc5c7a919df5c840a71d1acb64a6c3dc65b3552c3e6cd735d34461eadbfdb2
zfc5b80030ae094defea2ad6b03a4fa6fbdecac3a3ed6941316d5d9f2c6d44f4e92cb73124a91de
zc6736254f0a6a10360e4987746587c81be7aa97daf7b4b504636f56ed200ff84d44589468a2a61
z260255aa177397eae49c7941fe6067b70b8577168a9e560908cf20290f0e9efd72d2829d5ae4df
za2aad4980da55e41906a1045a1d5def671d6e4116807ad85fa9de4f5a3e7a7e159c2994ea9fdf3
z602975844544fccf8653c096c8d74dca10237210831ff2d8b4197c7b8fc6fa3910dd3fe99ae93a
z100f360445a5f4b3b571fe7d66983495dba9d1e105adab7b77123be103005a5a77b98563e07e4b
z300d6174ede586dcdc57816f656d7dbdf698eb3888e9d5249296ec4931a767907018075c4fba02
z3fcbefbb9c2335b634d28e65194bf31b3011da0cddb307476709ec8acf99976491fd75f10f40f4
z499ed1c7c4c3c33842f6639d1ad8ab5a24d0519d25023a61bb3e67d019b64dabf624ce006129ea
zda9e3c98a2898b48ac8c4548cef773c9684bb30d344c539e69faa5e8514bf75e8cc52a9f125886
z073a0017a4535fd308e14da5181a99a2d63cda91c0303f3e611d8dcdf59c819a6a3dff4c36ec72
z32c4a03739366a612c10650e62f06a0cf26edd291a4daeaa9b12f1e203a1f29b25994e97423488
z3ac99dd5a7a5df470777d1049e670dac91247b51425930b20a7a1870d9bb601cf90fbb612e5324
zb6a915f23769b64a890669550e444c79b5e612978d6fd1cc972f14fcf9689bf05bc079f717a932
z5c9c95d28f392fc460a6c860ece02d2bebdc3f72e9ef3b2d447d7100a6515565e2da3254d4efa1
ze2d47cfbedcd4d19a39af92707006742fcba67358fff09b6df5e6e2c53e78b4a65b5abd0bd0763
z4fa792e079e299b6ba3831d9e54d5567b1e0e505c938cd040295b8677da21467fc7e098bb64544
z18c7b0862e448b156f88c2bfcf434874fac590859e0df2d259a845a1f8c28ad7127f1bb9d88850
zf10c3ea9613d12cb11d77f0bd40c5ebcae8c36edbbf8688fe740013dba4bd96f39831f19217a6b
zadae8ffbd0664f4a73a84fb3e14d0edaa209aed6da6adcee6600ca66ed4ddc2a198906ba47417d
z2e08c5a545f40ace46846971b01a8b1ae624bb3ec242f2b67319775344eede54ee04dca7593b14
z9425f43f9a7059166edf5e23667a3db18ac3cfb97f650ced645b6d7c5a29c736aa6b64e08b2921
z068ded182cddd02f4b404dc2f201344c4cd5999077f17be989491d5043c428d3b945dfa5709c6d
z2e4e2c6296cf395c53a2914c5a076c0d2810a09d8768ae867ca4b2a0fed6e2be6e5f088677fd65
zd39a3647839bd0ca24d2b41e63b0bc3584121f050183340f815302bc05a5b0658fa0364db5ebc9
za37e94148ebfa85538a119d3e1032472379ad0e9522985fbdfd4e53c03601f83159b83de95dc4f
zf7e045281b15ec8a6f15ef34f8fc781bdcf6ecf69d5b3799c0f5052d0533b241e44963480ef44e
z4d42a4076ae44eb5805b0c3cbbc6c496efbb4d6067c7ba385577983d49c46780d98c4e871ce6ec
z1d25c2f957bea3ad83c7d25249ef0e563eab111e673e641daf70a247115a837a70f07c048b79e1
z3d449f57f9b650e3967735762d77cabeacb6e90493fb98d5b6c6df389bf17b8d5e7ff8b30218e7
z9fc7ee973917a52dc7f82ad0971cfe3d250584764f9aa35cba59ae235cb1c7332a25da416c37e4
z798b90ef50bd3d3cafc65de892408f663f3ccfa7b1f95e7790e985cba330f3d678571d9c438261
z67e0f6208393aafb18a470c50d8420769bc8b257938e20725e0ab8a1138e8dcd5f71e4b89a85f2
zb0f7a1736ddd7817f4bd5e672a93e0d748f2e54b38f9c00fe2c110fd9f613d69fe477109e716ab
z31d10717be7557f70efd5afd861831185b2701ab13817e05bcd40dfabb7e48ae9eb988cc8d72b0
zd4c1a8e17466e28a903fa4d029b727ce0f4c148bfc3a8d4aacc3a4d35dfde4734431950ad4420f
z3f4c48ef492b94b2a925fe988463eb51aaa21a10fdd8c40313085ade7768eae68e80a815821544
z6162462df6041409cf9d365505ace0c19c2758a19fd27d2b8ce87d1721e9c1953a3a0e88f025fa
z08d8c54ec825b4a5b1a8fcd283c7144c39aa08c17d534ef6d1eddb97e113755c05397feeb1b3ee
zfabdbdbdb1b6cec50d6efca33081ec165241ad71a7003641d50745507a4591278073acf485c7c0
z77afce2329d583301eda57d68b23cbdb3a5fbe0bf8a3bf218d5eda5068cd192b9b254838f2e6bf
z5efa829359d9f7aa5e52fe9ea1783140bff3ad752c49d06f427c517a339d30ce4e9282470c7a61
zf20f446b933a050ca58270c633e302f6d1632720a77a2d16f93151abf89dcda5e4bcd43dc5fb44
z162f85c8228440f74f5b1eb8e08656c3e15a460cb6708ba832065f87891ff0652441352abd5de8
za00807a6d341d81a541018f605540a0342cf5ad0efbfc2e881a952e15eb82fcc4862762cac3e9c
z6332ba556600e0cc376a820b5ab36b1663bfcda6c6ed742ae2f86091cb91d436be5670590d1272
za690d41d9c89f921810252d0f8e27485b707ec331506637b538359bcc3af8502dff7776db0f797
zca7eeb4b9898885227a7a2e8ff7fba8b1e8a26df4ff673a4ec3fddddedd645f7e6a4c723a3695b
z915692f4c3225ea20fc5d949fed399165af9694d4719a62a5a21a5c2930af0518ff79b0eac9e63
z7412ee17029e4550913a43bce7f25c8e7b0e9b8f0972781e51bb35c6185e8dffd7ecabdcc6ad76
z7e7763c0eb78b813ea9385a9be50867d66d4c0e18dd6ff71939a043dcbd16bc7b83e4edbace520
z5b24b86c5d0b5446d520a51c6b1c3af7670d5e204b7e8f738dafe9da2d1c3d80ca3f2863b7dbda
z10296267191b3d213539d68e7029098db51c24bf66a03116dde2011b395f5433198d45d536a9cb
zd399d4c3556539f43d5c4c9522f48545b061414673c800f066ecdcf2246d2daad964bdba9c44db
z9ab0a2327259becce78cc7e480806d942a3855c4ec0dbd225d073f2727b0fab2b1d2fa42c2b6d5
z63612b587a5b2b128b82159d4723161e0fa4ad67bcc76d0135dec7915efbac46ddcbcd051a316c
z9197c6e24f224fea4a849787653555818d228a36d41684b1aa758c5acf62a199c0f9bd13fac2d6
z7263d207521390876418fad1ccac902eba6c5a6daf35e853aacdf6781d99f126538052c8b227be
z54dffed77f1cffa95db89822a8cb5c466c59850e630b4dcfe031d9ab3d04b6cee921980852e956
zc9a0297e8e2aa03a329003b90b6d7cc889585c134d71f0fd99915b21a5b464a6e70b659d8f78fe
zfd0f2b323280dbf8fb6e1306dcd617280ce40069aa2fc488eec03ae8bd8686883d4d7c16322205
zaed0ce92f8997cc998a3deca4ce522c06ae8bc1afdb9416f9aa571139965c6f988134962b5c1f2
z11f136cc9382e969af451a57449f397ec7eb557dad7bcf0dd1547daee6fe7e35cbaf3c31cc04fd
zd177a057005476fae4630297a3770cb04c0a2d6ec44982bd24face9ce4757faab1e2cfe6b43a92
za646b7f857bce61918b94ba772253b8cc0fdc1d5968a9d31d47b7d60731519966dcb6661493ecc
zd61ea502bdfad87daf9ca3adc72403986f7d6ddee8f0e5edc6829feec58ff17625b93231c80c9b
z5ebda718ab182c370818c320110f590c5def2627b3d0fcfe6f7bf03716d7e1186f2c06cd83f1de
z8361782103f23daebdfb0ee10d5675999180e939a6663c7d4312151dba83c52383b6ac247ced4b
z8dd6cf3eed3403da0cd47ed98b71fb583d24e02120aa52cf3757f5132b7fe8c553af74e7eafd9e
zba620d94a5bc73790d2508f8c6ae791a75b11813fb8e36b607a8e633ba022440a2fc374bd6e726
z613e721fa3379e1fd6deffa6d662b29f3cb42fa95a6b113ee974ae587fda20c1c24197119db8af
zd8b1d099888bb0260516c01619da92a4efd2df19a9f29643c00157611909d1d17a39326fce9f54
z8e22e8b1644a342845218ad84ca59e30ef7624138344ddedbc70058f6c16890fd3f3bab73125f1
z01a27fd037945b4849b9877d984b5e800418e1051c34d100de2e8f181ef57989ef334dd30ac048
z929d434a5914810b262242fb543c1eb0421804f83aeb89e2834dc8e5221ebb0acad29eee64a9e6
z72d3c33a0908879c01f9c6a3c89f99f14860d52b794efdce13e039b71e47e8d6846920593f63b9
z4316985b7e9f41afbea6ef935951aace5dbbc04bd3b34768e7055321db41d836d1286ee38e45ae
z8e91b3615d26a4402d3a0f25a098f092240fce463cb53a10637adb31494b0078f350d7f2abd74f
zdc825db85063e5dc1836b28b86b9c43b865e949459a677b026ee1ff337ef2ee6d7e29df0699a0d
z986669820af7a1f9b39c48299747fa6195d2ca5b5be039a337b58b4adf5f20ca318cef3cbb92c1
za0396ac9d06bbab1683cb54833f383fe43e4e22629d876599595f367719b6a4be9a1f6f21365a9
z4da686fa7fe5c2c89d41ba7648b859e3911a5fda38330c726dbddccdd22c106bcdbc41c43d359a
z708cbfea10de6ad5a863b973434f82d4e36d231dab50351a840ca31ddae56c33317a0368a7a8ad
z3aa071e003a4811e6b113c47654f2fa7ab0cb1af2a0f7dc9a35e38652cba23a4bcbab21890a8b9
za3be5793d270422ccd5722e63ed292116342dd224b78a805baaf3a87e09f2e11ad3ed4359bc855
zddb0234be19e61ef560b07ad2e58080bc93e9117c7ca0d9bd08083a70789297cb98fae80bd1a78
z37d201a143c62e4cb5dea35bf603f9ca207c6c58caf04d9e1acd6c411bab02957bc9ff2291f803
zc1d68da9909b946fa9e474993cbe41fba66b3604675f41a7d986c93d2b45dcf81688166072b586
zb634833b7ee86d8d2b5194f48249f5299132bfc73b9363eb81da35f4727d6b13375c039846f290
zad9aa77107c492fd9fc80c855623f81e64a9f46b81aaba6f730eeeb15821d0b5c7fa1086ee44db
z4dc44a00572d7cc8e8889b78b5093eda0ca6cfd4289da131145698abbf6ede037f6d1d1d87a38e
z97e60f8c2820e87edcb83bb921ed57664372c7086fcbc5e213317cbb010d6e70cb0c2844df525b
zbfd37b54fe0498a58c1c056c9205f55a05874c00e4f4c06d7a00f1cff19975be90941834c87df7
zb960e00ce0b94f5bb54e697654515b6ddbf0d10fcb3f60479a7b4fe341cf5acf01ada4336f2700
zcd9126952e08bc0a8b6cdeb8500d5c67edfa0a10dcb16ce28a51f0d1ec376c80f667c39674fa71
zddb346bb0b9c1739295be2ccde9dda8f422c5c35a695365da881b58e5e975ae7d82486d6ff03aa
z671e47c98a2f6116af7ec33b734fda5f92f3905ded52054def74d829ba68013c5b66be279f1131
zfad5a9510ca088214cd02d2fe265727cd32634de1d66d2fe2a209379c9cece2959ec75506ae640
z36b23e9b5b0e7942f9eb6bf2243797ab91e35bc1a713b7aac8c86cbb0d6dd7b3d4c03dce38179a
zffcbfb2d0bf0623a27d3d6e4229edeaefbddfed30d17695c995265b3ea3f1475da280136549773
zd442220192e4b34958aff718da93c3b64efb903e4cad77c7d35d18cb0a8251ed8db07f28c2a9f9
zc19c5d9c253f29d133407645315701052e0ea336fd75261254b2ba56cfaf64d8e1cd972a3e8148
z9c8df507288d83adef3069f17b5c59aa9f3e7554b14c8cd0afd010516ecef9b713efbf9f21a198
z2621eb02e52749cc0fc404faa20ba9321c94c9ca05e076182c82e44ffde7af268810c460934bb6
z04742e781dc73290d20bee5860f9ab375233c12c742a0121a2be9b91bbb3e5c38b7716ba2d7c60
z3eb62698a8eb15277a16e72fee74e74a1225b10a1f5920db249d61c9003074bd5c4d0b378a1e02
z93591f49a64c5fb7246647da122aa4816fb0b71eacf20659c06bc67dbae75ef81795c5463c93ad
zaf365cf884b6f11d3c3220e36ed9ef61521194953733b3913366c569f11ff87b389d969e21c61e
z3b3dc22262b6a18b5c196a47134859b7cfb6b3af3e524032a39b05122978b1383fada712af0196
zc53b09fb39ceae32d924db1476078df4c137bd012f98fc2be43f8f4420ae58ec83c8c94f329f97
zb4ada5919d200f3eb2f84bea6dfa25c6308cdb6a642ba931d8020ca1cbfe7cd2f48bc334511c8c
z25bc67ba8e1faa8ab12dc425c9068ab88a14f2039eddede99674b7365bd657df2149f2c4069457
z2b6e5211239ce82e4ee648b952115f1bf20a80b8ece4b082926195a09ed2031849d20d39ae2ccb
zc0d71896ffb19993244892aa6f3517de1c4459ae574dc8c6e8174fb42307b0bdad4848a3aace59
zb202b7c9eb04b44a03009edef5c373610ce32a917ef1806080261cf62f4e1c294d68bd6c922671
z05491398ccb0e46190f9bd57a192a01300a4d21939caede9974c62b6ccd0a23cd564d608921039
zbe17cf99a8f3a879af80dc44798ca4a335a0412f80e265ac44c073096a48f63f16f0bacf081624
zb98392a1d6ec8f9e92919079fbbcfc37e2b376decb1366d0846fb9d88ca3e5466df8258402ce44
zcef44e834cae821b42e3c7292ee8b5a8d05f16c580dd3362d9ad7fb210a816525ea782539e17e8
zdc20e4f820c52229fb4537709b7ee916e5ff69fd0b8b015ee6f0286baff97d4ca6567c4ac30f0f
z4d975ac4097377eb455ef18b80625f9a1d3f591ecd6acd8c656636c2a770d219abadb7b4685fd6
z4414ff5d8da0e9504803db47388b7c19bcba4d871615c442176770a86235662c3a813a2cc63953
z7cc8f4a111b5eea654d30ee7c385c32e13bfe043b2725307f744b7d5532d40879d6150355a9774
zc9a4645a7c8f4d82a392b4de9632113022a0f824e50b39a1619e6236908d46e0974458b8b0ffd2
zac140c811d361cd189ee64415a61c46f81f91210c0dd88a249396a57426d6237178e98d65fd31e
zcc2ea6649e683461c3e84e760224201f9d77886a2cf63bf1ed06ef6b2703d21c6ebf1d74515680
z2cd94ab5207ebb7ced3a24c466e268981af5550ed054616d97b240b5dc4d0435088844ea618f5a
z0942b542850280befc94b98557d0575ae40071d869811878d57aa14db021c57fd07ca08c471dce
z98c4379a6fe4f92a6f5cee20799b65d53f3086ab2403dd457cc407cb7ae5cf5bf160d0899d87e1
zf6bc8e2f30267a184b6a303f934b2af491e08efdb3fcb84e1de365788839bdfd164a31f5d244c7
z854fdeb25a9dff0384c06c18c4436de8d76bbbcfe9f3ede972e6a5145f9ab04c959ebb61e7cbe8
zf02298c76165c60ff35f5f50b0476543be5613845c2e063a7c7640e4802e36f69f0b8602f09aa0
z3c3715775ab9286bfa1583fcad852467fcd3755b6ca54f0a021d8defdbade9ba4317b5aeb6dc87
zc5a3e45a831e9967ba494d29a7bb10bdb6fb37b2de49de7e0a029b7103c7aa63bc8cb99ff8662c
z5a0967b417b670daf5c59f44c9c1371baac32f58385c3e3b5616bcd7cc8805dbe47b4b12d317ce
zd89f83f1a3113df4068b0a0a68ad002ddd202f4e00e3b41b820db4e2d5d9fcb33baa236fcc62ac
z22f5d39aafeeee748570401c89a00c6713027c62bd57d034a4610228e462ceba4afbaa42748b13
z60ba6b70e46bae97c67a585af65f7f89dcc3001a77547634749284c151201d9372213a70f7899a
zf2dfd4264fab585c50795a9635e0788e28ff92ee592b9893606200edf34a93d8db326ecaa8e6e5
z5c98457a3ee752a848acfceaba4711cab5ae12aa219aeb4c8129abc1d3509d19a7205a5052edf9
z63e5e0996f4348455235c032e73a4a34fb47b42bfa17d862833fac6172824b757190e8697fcfa2
z662ee02a55bd0110576b5b321e15f6756ce7e35cf437717d02fa7f26f71345e9a836c0d634e9b3
za95e553b2a91a169a2e9c6f4b56ba4d8f94db4d958279013c7a6d9c95a6c873297ade9a131cd12
z9aced73e04ada9bd922f4b73557a9d0d63f6ce10a7e836a0b46dfd3e57d09db2a96c27df901cfc
z4d01b8cbff55cd3195da98715753f008284ef8c2b731510f12c1545d9a1ceb81d85e3bc7404688
z923b6d3a821afc38af242e4fc254ef6497356f7a4c9afe73be99a9d1f5da8a6324d83ba03a0a56
z6c717997e1a12ee6eb7d610be54a737694d0549c2eb111196b305723b3fdb4f40e24495282dd2c
z1a534538342ef37ee1ceaf47d944783afa5d220e91d956d55949579d9cc07e0e42b116f2522015
z22702f52528c870e59afc6341ecd8503782737669b364a61c79c7c213ee3f1b2a20b9787121d76
z60f0d63cccab03e9a92fb9fec73a7279c07166521f6096b3043f56db8f2c3b4bdbde067b91180a
zdad66c5c901558ad6c74b2edfe615ba683ef57f744691f10579d9bf962aa6d4f8ed759c1a2d298
z1fb042b5d50fe747f1b6f8857ea7a52f7184d70cb61addc3e171ba92da16db23cdf6c8a10c6ace
zde6183a6cc12b7e3999233238116fc24e950d0fcb81d67923b87e44ae215b360a63d21e9625846
z3de9088087b45484b54b2cda7a61e0fa956bc561e5e477f712731ccee6ed934faef61aeb0c03a2
z45cb3f47167ff7a18a1d603797e28833811e92ff7333e90b9cb028ad7954aca5ff2f9c5213a380
zffa9675358a47c1490a61b56e606b73887dcfb1ed194103d1e7f59edf74c65ea9bb4c9ea47b107
z7b234ed25188b95d96738f995f8d0b798eb4675f3656038c0235c2bd92c4526b0ee898937e6d63
zbad0fe9c14d3f480dd8effa41355457e5038bf429ce9b9220f54cfbcdad145393326968e8229c3
zc41d0a8bbb7d958d55eebe71623e4c5d8a1b575129b753bb0a509ff94e88f1e3c0c9b044e96c15
z225843cb41ede22382674710a52c72e25a47929746f3916726450f8c23b4de0e6bbfb0910609bb
za321b54379f72108d96808e2edcf7f8a55ff3981ee2d52b7e91863cc4a5917809d2629a29927ff
z5eff05ba918d001ca1ccb4ff61c241140098df959abce79a99232d8a34794b07c9bc5d86ed1af1
z3cf48573f3ce235b3d4e1d6adfff8bbdd889f7efa2adcdca460e69a070f7942502671012007a88
zefcd136a4158aa51d1be4fd773b19b2876f664d0ca481f58e5189ebb95bc787e220946f7a1084f
z072950c953e79af10f614a711ada5e964c4ac0ce1feeb6bc637f6336a772a6c5aaa4353c2eed60
zc98a9f41f24da07f4b97609fb4126f1957cfe7b0974553f39b7da0276ef27180bc9b9881dde421
ze3485ef121c3a907ee7245cf257950c83c6eee905523c9c9fdf97f252dd6107e1af378bb74d7ee
zdcd86a2898929cf28c556804de591c13a06916cefc5e76b9c88854b90a2c6ae5ca85ebbb7c5638
z4ce02ecb9dab2c3315a4fb621ea476e5c5e4bbbec61bfa874e76705d3d340354c80aef5187be52
zadbc2f66ad5b17091b705824ed5c8fc13506adf974184ed889ce6a84a45bb01478dd0446df40f3
zc140b8e68dc41e3d7bcff7ace0cefea2df073f68ea063ca25837bbd44b7e35a6b36ce4fae944af
zaa6ef4b2aa966724db9437b04e195247615e513f2fa84baef13775fcf4503c9b16783515c3aa66
z1d2ebcfa5bc024adaa6ea34e7d57d6e5b1e5418e8c144a2513f5916b53a0789ebf038d70e98c32
z11e9d8dee1c0d298ad3d842b4008df96f4903a620f1aee7e965ec1fca99a3ed0a90c5568b174bc
zf6f3ee5e6f42c81fa69907fbe43e01d5bd9705946851b1804ffb44e56670255a806e628012cb53
zb840ec3063ca355cb93293107a147a773ac61031c41e0b050e8bd14c7f5cbb124e049b02d19da0
z8c6e9a24118f40f415a320a8ec285694bccc860c66b276b18c44a3bb4df837aa515f6e94e25e1f
z6bb5a3bbe8545a2b938c03443d76fd1d4d967dbe618f061e2001d8f6029fe7588652ae76366922
z79906203fcd122a87388b498f359adc2836cfe9d404c5a78100f6af30441132efba403a09b88d4
z9c87ed6fd974a1db56311a0714790ae1e3f375bfbf163dce66f0c6196bdb04d02ea490fc6351c2
z6fdc96c78bd4b5227d3c166085837d6d30a8fcabf5205462717ef34f07369cc577114022dad9da
z6c7de4a99943f1dc68cc1afcf91788327500211644c44e95227ccfedc37fc73550d8945a6bdb0b
ze4be7107af36e7219815b43a4bd5311fbb0e7702881d88dd4ffc9ce22582042951215481bf76e7
z5e9ee05dca0b13afa509af5b0b57e4bd835d36d808b6292e4e60d4379c304c3b35eda8d18c212e
zfdc264b863362a4777e75b0cfc4da68e66bb8baabe2dec5fb6d35c10dbe7fad2a1a0d91c1fc685
z18b5f8c475a3af6af6bff65602614d12a090f1ffae986219ab23d8ab2d2bad9576b016e8cc8312
z975b08755b3322491be92e5d93b1e5f69d750a56afd8cc1dbae7642903958d70476985e5f1b9df
z3cba25855c4e8cc4671c06e6389c3c244211699067e06c8383c557134a5d8fd547fcc783edab8a
z5a651f19acdeaadd748670294b6a4edfa2614627cfef8df13e9a7aadca8d15dab31ad0f23fd701
zb863fbf52191430cc7c106d41849fbca222e87a746494cd0c1cdd15396d3e2e335cced1a2e8fe2
z7963280097ba321db13e04dc29dc161c142d0d480ff0985f7e1a7ed9940963767f4917c2f38579
za59787847141c149be33622f63cfd03eac4b1e853b04ac80b417eb14d518067d6669ac2fe0b26a
zd69c3a5391c4272576ed337517a25a91faeedaaed813ed71a4be9d17c4bc6cc0a7950d02e61d98
za519e3dd8c12bdedc0027798bd09f61a2ef0f38910e58b28c2dc8250fe55644077a2b0bf984299
z6c9e819a0abfdea6ca13531b8392d2e523886e7c16ca8e527a2461550a750f5ddfb18803db1263
z6c20a625ff90380ec831815c55796f8d10679178b174742086367cf9286dff18a28933d80147b5
z7d786b50af5c0b3a7ff8baf1193e84f516c8f6bcc115b620dde3e7a30b3bdeab56aebb32363d33
z08e91e061448a1c5263b5ad368833efe4dd4533c4fe01f4b92ec7967b934367d75fc8a4dd99f42
zaf9aa751d8faaba560ee306258b80510baf0d754dca291400b618582e4aaf6428f7acfa8b8e24e
z3a802e0b3cb44df408d3cf6550a2998a0a6ad3448d3e7e858fde9fbdd3912b46f186992b2d99ad
zfd849dc66e07b2780b43d90fc54b39a6eb06d785d7a49b9d1c20af708419e7a4190fcf7dffcc46
zc83baccc96cb916132b9ac8f3de7b6216c6892e829c5222b809f4029055bb65d68fb7073b195ef
z4abd68277b412915ebe3d43aa2d098f8b200de6e31e7638636adf371dfdea709a6cf9a07fa43f3
z39da92502b2caed1581f91a6292cf62b62f568717442383dcea2c0c3dac6cdf0854564c67712f7
z462c18367538f81c347b3eced897ed90e7dd5527b2078d8090fefa8ff5915125c7e121b1d881f7
zf3ef562c5c0d3c1ebdc162a6c665d3c6a218ac3c5da37965bb0e8ea33534fbcce123a733086d4b
ze00aaae167ead7d337664e5d9c15287cce4b5b064570f71835b8f97a8fa98f500a4fb8fe509693
za9e3c76ce6409970a7f0da36f4280323323eaeded0fc316d1471ddcaec101f6fce8ec133495479
za2b9dd6f53b548ef0ab5c0f5948096a2cdc4dafe2cbfba7ca43eb9f5bb9bf1c0ad3806bd1571d1
z8c593d1a9748d50954be3a2f67d7138bfc844493f7f8575c1fca66237daf3fad527220353fb6e7
z9f8c45746701190c21268b1948f4efc8d97c1b8ece70e724d32fd5c5b79059260dc3dfb5144ed4
z8d9615e9abc173fae1a550059805f72e8ca5f8277ac612cb271ca37b9a6f7a0ea0e7999eb0fbe1
z518c37453559949d508e642768772c612a6579fc2b2f088eb9159ad12a286b9b87eec0fc5bf448
z8d65f119dc8356b4a2fde0e3b8e1c12131f937c7e7fd054252f14b9651f35f829a8a5d11e8607d
zb17bc84f3075e5d08cf7ba7d7e02501198d93ddda908e4a5090a5d88db811bae2a095c97591963
zf36ecf077b5ab2c353490fec5eabfb840eb6f486d21b0fff3ca71e854c8f5b2209853b35f5e9ac
za9676d0bf06216e5fb5f4e76fff01544ec6f4ab10ba3aa8cb014ae9709ea1c5c98cb60558887e6
zbbfdae492a6554b023db9966182a27940954bafa9b3a90ab089f0e13bd2f60acdaf00aaf79de01
zf803785b60269acc34c1ad3c3f476c61fe303284dc0cf68f4c29045df2aa1b8b58ba91bceffcc9
z59e46110384418cc670de5de3e94c0eff6b6ceb5d80cee1ea1a359b8f9469f3f631b500623fe5a
zcebbf5fe4cd09f708446b5fb9ae23fb614062f0e396fdc3a6e98b27a73cc3a30e1ab2e8e2d121c
z71bfdc201808eb8feefdcc770f6e50d90fe7d34a25fb17fc086bcb7b75321e8081c7c3c5a4ea43
zb90bbd148602c7494a6d0abb40ed2531be81e9f4409ca74ae73b8b39636d5de749c1f2d9dbd853
z008e19d7b9599afd9a24a9704c79407232655438e30c9226ff21e2d914083fdfdee265c3457ba2
zd8f27eb915fb6a7f32cee3a3fc0a5bfa3ca1e59fe33532c514bd397e86e4e6c4f770ff98eb4f74
ze2c99bb44955ef232d867eb31b535901cdcd0ad15cb202f3d1029323e4ba11499d9de078886ad5
z5d97a61c96d54bd05d08cea0c23125678cac3adc64158526b1c544a2ae0a01b70357bb32583d76
za7cf3816432063f789461091cc7aeeca019d8d061b7e92e6a9687da1d9ac9c1217a61649506bcc
z739c7975ef6177355ccf625503f72dfa42b7a2e6a01153638d84e4c30bc1f5dc128322a27ffca2
z2f147ba0ddb0170127e72154171ba0673b988159b5d3347af987a6ae5942093e8dfa3e9059000a
za8286d1814f8e7366ced86c4713a4ba674449277c4ed9501ddb559b5c5ad114a93d9bbc621e0e4
z07327bad5c47b58fd2fc904c933e6efef7eae3862eb2b2426289a6d925544b3bd236ba500bb0da
zc13a79bb5a3faec221fe78356929868c731c1ba11ab401307d398b8e996f250c60c78c3dc94e26
z64a43485a12d759fb33306574fe2a779fab88e6e67b3443c378810d5472bc8b8d8c9c0359e290e
zd00b106f3d2c90f8b00f8cccf58e3a3e94e9a1cd6f6b7adcb49177da11f73c23bd44bf55f536af
zfe0cab7ce1f0f1c854712dad293826cb75e5a94dce65bfa032252122f5983e84da55824d235d5a
z13b973e5948df8047587d0e65d13646989e26ce7f3ca074969366452d107aaf4488e773c9805da
z8644aad6449e19267d184594ec32190137e9328bc812845a273c6d311067e6d3e2469f5a4f408d
z1e3d3beb0ba478e8d4d53f15db1d3f71b4cbbd23467d52868588cc8552492966036f593d7c9205
z4f215bb3577a6ab8e12128ccb1495a953b52586bc0bcbbb5279d93cf7d80f7bfc26659331b6865
z134c9f4bc2e4b590e8cc3261bbbd6dfc7320cec297bf29cd726f00945654e7262b46074a48b303
z45c91d94867121d9f65204ba273ba8f62058696f6fa0dd64965777a7405a8ff84498d615207984
zb3559a9d76af94c460283001f24fc1d12bccda6106047d394d03ca4bac4b8b1044b971cc822226
z15bb9c6f871bc4739f52b16fdba48f02dae6d75708b05b13163f1c283b34914ca0005be970caaa
z61e6d957ded1847d364e223059fe1a6f70d144509b26d6fc6f9229fb21f2ca072a24a0ab681aef
z816fd4d175c7d03c434aa1cab6d0ac19b7d95e3696ce6e90a5c510755963e66958021bd08b089b
zd551354992476fe74dae23e1d58217178447592e1718fb3d7e9a305e28143397b5db4f55bf5df4
z35d29dff3ffb5c17fb6a0d18b0bf374fbc1220f519bb8e8776109329972ebf54626834cfcacda7
zab462005fb741d9f0e57c3ca5bfbfd53b91f46b912ef8a176f3c59a7d323034d3f6807583b80e2
z244540f13c787131ac5b824dd69aa31b2e98529a8f25745b17374cd59c8c879f8f702054a084c5
zd3bc22fb96c7ff27f8bbae9a80bc7f12df53b2075d3070ee574f7e7d39c5d444c616e4bdb30395
z411ff334b9bcde1365eb4d6d1cd8aa414a1fef34e0adfbe6f72da7e9d3374f46a8914f4d17e1d2
z2af3c4aabb5a844d6d99b64206ce706b53e0e0febb5034ef28382fa0b09f831bddcba8d5fea605
z04630bcf24b09a9d0d840bf3dc383cd462d7743b1032e143c0c55b633080bf6c5fcff09f30cd4d
z25c6bd16a795ad178ca88cb7efdaffb7ab176793aa76c9f3e64e8c799dc6dd485521e3059c45bd
z3da2282bad0587144b79fcad6e13bb14500aba96bccd7f2d1f96341ac20848e7e9a37bf588edc6
z7dbb8fc4b43580f703f28d4a58b18c31d81eabcbe6b04973a3e04c480374a5dc327c0d763f2787
ze2a2f2be1b61bd486ded1d29e55278af893f829f60540477c8bbcf3deb233b2b01c1cd3d2cb35d
ze1051fab29a1f4feb797f8b96b071cfa252287dfe06f715abf409c1595bf29312b90991ba2edad
zef9d5ec9459a29756d56f9d9a645bedae31c6096ede65114a2a8bc211aeb2937db4eeb35d653ee
z610f1bc69f1b6b97ea3fb453f44c3b1f219adc43ef7b8075a367d9dc06fff45c2b6cfcfdf91b19
z5fb5866b281c468a9d3eac60a1a07fd2dac6b1a810f83f1e72105fe2ae0da566a9bf53a899362b
z4af68757ba3bef646c8ef3d8c6c20117b820ac58ef7f12799ce43bca2be2176bae883776086a74
z16e851e941c86c53a5c879fd604d8f6ee5bc2545a236740f89defaf3621787b467eabd2c20e2ac
zb897fe9cccd3dc44a1241cef79667f824a540ce02f07f3376fd123216b77ee5a7e112afc20ec83
z8182d4ea9445d84f6546b32f60a736bca6bb06d3d3b6be947bd4226c59844f786b3eda20b2eee7
zcb1b33d8ec95d60bff25415e91828076c35f93f6560551ffd2f35b5c449c644ca2660b16d73a54
z4dc7b9c620f4ca95aa797151cde504ee186d25562402d061272eac75a3026e99c947fc9363353b
zfeb38fd88b93f7a4890300892aa07f2bdcdd47359dbd70f04c0398c6e621e75220c564438379e6
z80be2102e1ca9ce941c8cea99b1748157763c11893eec2beca17c2e17568347bb30e703e7e08bb
z5354fcc69f18919994f800140be34e44aa5f74a08fd48917da72d44b0d6574bddc8ae20a8fb869
z7058859227131b556e51bb2b22a11c4dd6d774a25bbce1ae2533493cc1879b01d4d03548c725b6
z61a8e701daed2b499e263b26fcae867b63386495eee8ab826061a6cfd327b6785c50bfeee26cca
zde9b010d9690f560f9f48aa83565736c9fdcf50c8edd4ae132687bda1a5cd11111e0fe6e156b53
z8f1afe2ef37ee71bd0d0fcdfc03f0124ba965387d9e9a382e0085d30712f927adaea3ace26f053
z4f9b74a7907cbf7e8274e525217e00c08f218d527628ec02bf8f4fa0013be80251ee193b5a07f9
z03ef09d63a9223170f4a706e525e3403550612a484a727a46a0751fe3ae6126184d6849e5266ca
zfbe8ace545c99df466a39b5aa71aabec2e7f1a8de674438792014fe77f816b9af17bc484f5677f
zfce7b4316d9bbda5bc20157f1ab2a76b107b28ce65e55aa2638636f513f65c702c302d8bf812eb
zef6322bd05046f089d198f86a595749cabd66f08ca38e30c1b1f42c85ba852034076379f54daa4
zf4d9647db2c58ca1ff88e4963d2359831ff7f1b5186bea65ed030a97ee39daf7eaa8797769cca0
zb900b4d7120d26efc473566f8a5aeb5d6f56a9729ebe78c6da3ab5542b8dad1f337fe6283f9cbc
z49057947ecea0c36196f00ef4b54bb96eec2187eccd226921374e18f010d9fa9ffe9d76e0234f9
z4df680e9956a463f6bada28f27612a3845d780f19be28e12cbb2a082efb1b7d0b1852423bc8c23
zecb917d89d282455adc2b21a3e3232cb313e881568f23452aa688853b763221044036882595683
z6d00af9ea0ab3f00be156fd4238043dc6890f2e23816498665a1df113df49b30e8c491b6ebd7b8
zff59317a3649db397e71b6d45cddfcbb9c157fec4dff4efc8673ac5ff75378db539ec447c9eed2
zb689649ffb619f5407c98587e18b1908d9eefb40940e93ce111f23745f42faf35b1a9fb9ab301d
zdb9be5af171863609e6e8e558ce587e3486067a4194c1ccae3e20dcc88738d51681f7df4e79d1e
zc4b02afdc71953494bef18beba74c16272dde35d33bbd9f5deb7233c74eb207070b06c70b9e8a2
z2a25882ae1ed9c5e03c98f88a98d7eeb7da93f783550eded4a62a25744ca8ecba659595bd0ea38
zf6ccd28a6e76bb2db0f16c4ab39d60ec7ad8b93403283e905b5b9f2ab7768565567e6e3ff87cad
z5d3c0f3a65fc1bdf515bf2bf65285e5e488b370df6ab135a0bda6b772e1a6d72e8fe0d6153c6cf
za4031c9abe0fc275dac0d13f3c9708ec74c180e54ea3b6a73c55ba5f0b7fce94d4fda5209e6631
z9c8beb701ead09f9e6d83e27b952ecbb25f36f42bcd0d60638218d5cc02e18bc5173b2ae807b4a
zbb7e5fb10aae6dbaa9ab76e54650c8eacb50635a18ec35ad1bede022d8b1b94db19913de83a5b0
z26b07e2ea04ae4307c3daa8fd164d0bbf35e681092d9a4086d92be4920f8b332a473f966fcb674
zb7ef8602a5d28113c2b9bcfa3c396e3f7408506a76e62b4de98a337367ff4721852d20fa0181f4
zb82eec0a899af1c7947eeabebfa1c4acc76f8dbcffc7713a53719ea0d5822fc40775d81a6b26f4
zb25aec8d
`end_protected_0in
`else
`ifdef MODEL_TECH
`include "qvl_pci_express_link_layer_monitor.mti.svp"
`endif // MODEL_TECH
`endif // encrypted_0in
