`ifdef encrypted_0in
`protected_0in
ze74c34e226135848fe16db9ffd31815111b6d7fb642c521a3f628cf6da949865580b22efd062a7
ze90adae0e65e66a2c36a587d0a790699161455169ed55a01f2084f11770a774ec4c588039b380f
z6de9c5084882a40b79a175f5c2114b2b6d78b070cb806e1c0aa9258297f4687ab308bc470f0040
zb0b1de382961eeeaf2e279e1462520fc31c119af8f2b214846f56c2b3cd2eadbe4099496abff18
z15cec83ec4a77b868344aa20ba7360908f5c0de2a79abf8b3534b883bb12180f68b5d4beb444cf
z3fba8f13afb0abfe8fcc4294810f75afe452434d2d0f1166236c82f76edf1e12979f04bc35693e
z32ae028996dd85737a8f5adc1ebb94f39c940246e887647b64782cd7ab429b0544c173176cede7
z01dfb26b1f73408344a52b7e1f117f12bb9c8077b34876c2e6fdc085981637012dc9754765e1a9
zc512ce062e0b8fb16a214591f5c81e1353b900a611fe1f4886b57940b41b7f2ce99a7b84b04b90
z916f717e73bd10589c81e207ed77ec660a8cbed5b487fa50acde1b055c8870bd8676023f21ddcf
z9c98cc47cfa2d654ff1365d1f45035a045a66c5dfa8279050262529d2cac9e64fd27d9c7de62a7
z731bc808811ded9016570962244887f98fe5440167bd0088f2f049df882af501358497c3b28776
zcdc5426c7f52a851c35106bb93e16fff98478405fcd4d89273452c559f93e5926bfbc31a6dc7d3
z54b24d4be133c2e8791d1a3493ef5eec5ddc7946ad0ea5c76e2a70b7a3c0c8ed8a71b6eca7e25e
z09da4537f69375b93332cc993e3bfe7a3f2eb4e2fb77f10684aae015976eac330f6e2dc4032528
zdaee88efb81edb67f8dca962dcb4f8c831f42aeccb4591b53c1e74ec19e8d7d3d27eb793c8a8c4
z99d682ef0ddb26fd7677cb8de34f0b2abfbfec21dd90aea081f28ba71668238d70bbd904e74e92
zf5c87b830220684189f6b35a94f4f206b05d404252ca15608727dd156ef384dc4cfcd5d3cfee56
zd1ca09fcbf46898229a03dd77676c37eff12e9958fe2f11882f86bbff66604da1fe6211739677e
z6631d595308687f912f58bc7035f936c1cadd726036f9bb142e5771042f0473a2897b452833754
z706408a32beb1def89869a4c488c6f81a5e95e930890fe82532abc10999f247e5144094f2e9fe7
zffc8be7a7edd161a0e0ab4caf884e334ae2700d1b9fd3037f5dcd7e6342d7a2e4324a5f2808b7c
zf3bc405ada533d9a5be4826336f1d7de493d338839c860c497719251ca3bea45cf5f8186a4b172
zdab56423c69e822de183945a63f5563f3288a1369fb04f3effe170287074a6df7676c2353e49e2
z663071c104a637ba480d15faaedfee764aacdefc5c4f018390c766b7af6934cc3ce7f8a3da854c
z2925f2893c323f9208b7211f930a0d7a2a18a35a5b4376916a1d6d2378a09fb3b5886be6af5ada
z58b226cd7ecf98fb37cd81f22a98814325610396e177ff275602d7d3dbde80ea90d4092a29028d
zfd35dd24c5db5cfc30aeec4c43fab38f1c9a5790e97624ce234ee8aea07b74ba7b158ecb8525ae
z2b2840c525c8645f7fcbad5653f8e40bc392a2c3c78dc8ff2bb7d030f845d85c46772bd24ff039
z29786c34a5b0dbe3e28b34cb88b08ff7d31c47f9d3226f7fe8e9f4428ead631b23234274f9e9a0
z099fb8e6a907009a0c06558e2865a9531b9011510e372e5d41c1e74009cbfbb4388db0d70a4a43
zbe1832160379a388269b04f81aac6efb29b5b088bcd8865c170fe0bb2009782de4355e051ab647
zef28989f9fa19d6ff39c0473da1bfbc43ab67fa8ed57c28aad5828e76ede20ebcecc016951f880
z3fdc8e0d769cf78f05ae94b16ad79cec085edbbcfc2bf52045d4c98b52589a625fb47fa8f98681
z351b2970db68c147c30145d511b20cf5e991b585210d6cdba03eed6268d41035e147c5d47a6fb9
zc849cd639f1e510a85eed56625794ce9ccc225fdf30485d411d33fae357ac52d49c812a86988ca
zf1dcf73bffc8967f31c3286721b35669b6b5c6bdfc61999f4d5494dab3262705a4bfcc90241b9b
zc75b65ff7129dae691af63443e35488c2075e264baed64bec64de38254c056dd7bb4468c7b3673
zfc70a2d4f1090d0044d1773d0dbbdce4f03a55e16e277a0d4d55da52794bc9245a6a3d14d4768d
z15d5e6f42b6d475ae72f59bbb6a827d6ce35540a895473af043c418b19570f4c62d5311c19a092
z323f53a8a478dbe1fc647b4962227c9207cc0c58906133b64940646a88abd142556631c3bec51c
z791df0ca9aec9a8b4c058bad241976b54676535dfacc77ce2f19251ee1a0f9d5dc2112090443bc
z5005b21e4662e1c521a5fb646a021a26b7c00c14f49bd9ee0931fba88512ca981cf8152ea5e804
z2b48cb2f2ed2ae30e2170905008eccd80668a6e19d0a215f5669f6534786794b852cf4b77d0b7f
z18d7ff735effdcdddf60ecfe76ca3c091ab89db36a8859f2c45d2ba7df40e6f89e62d29cd949de
z6935c0d6e08b292ce25bea306b1655622e19b9f69d50ad7cd914c234460743704b2d24e7bf328f
z452664a36fd6cd151841db08a94cbcb2f9546ce1ff8d8d6cb5691417a73860d96e36076ec2e24a
zaa740c987c98a44824c2863d5ac0e6ac788c0ed81a3cd459532d7e3da4d056750de496be102f2d
z14dbcca8fc6498d3e0620b3ad5180f8648c3600b9a0227e696ff707e9e7e9383bd0daa420ae12c
z461859e08c9fc16717b0e820cc9ff46767f9dce4f1cd1151c5c2ec117d2f2095af563d18d67f64
z370811b691ad7c92893f571c20060e8bd97650df1a381c99da92827ba9772c15036ad173055926
zd375b3aa31511b470308ba7e2185d82e53ccbad3480c9a8687fb1e423fd8d40614d7bdebdec701
z5585eb193dc2b75e4c1ae2d57480678b63a7784ce980c4824c99722fc4e54ad7b69de84573b4cd
zb16cafb1a98262e21c73baba89eb53577a119c58e29145767a179e0d2f6410f0e8e7f9f36975fa
za4ef9b854bb94625a3b3297fc8ee1ffeed6476411c282c0d1e1286d356f83dcdb0507b00f92eef
zaf6dda443cec1e8c5cab53315898025875f85a6f4137c2984449255bfc137c7229f2dcf77b38ef
z6a24780d1068753796cab2234f0c89fd995de15b1b820c8ce8d229da7c720303c05bb1054ea61a
zd89da0df64c8683524da4dc5ccd5d97501f37c50484686c559cd8dd4d1f9956d37546d2020b0c6
z478f9a255d917b44eadb1fdd5fc2d40cb49edf5bf2d059681f42238fef23a23653f21b276d5d84
z5d2a01e2c44f57484a4f0103846405de6078e4e990591e7ea4135114b063dd2cc320dd194354a4
z62610f8de83ff1cb7c80655ffe1a8bfb81f6b6361601a5337761e1fcd0bb84a67299f31e404aa2
zcc1c4704cb8b8e7c8d22ecdbdb654d01f794a4e6798e08f2f53431f700fc72429c800fcab94440
zbbc66667da0eb7c20f6c29b53c09bd22d47fa7ed0d7fcaa1273a3e6453459989102a3653f61440
z54e883b0664489cd6bde16ffc8b3341563137973cbbc8265759e755d704c044fd8289218557afc
z6bb9fada1fa9d99f20be49162538e2751e4b9034eac2631c91c81245ec7f525d6d0bb8ec302fb7
za57b7bac7a7aedbbad3751a56ba4ebac7ce4f1225df896bed2f632633eab2310b9aa1b2be8b679
z0e87c7edbe61e57b856c76dab7ef785aa8c98151ad00d11fea646c74bfd9e89b80f2b502ae192b
zee7cfe24ae5892c1067b19094e36be80e3ab7ec41d3a063633f00dca24ba814dc06dda377d661f
z22a5e3960e8a45d3ce8fd9fa579c126c1f4631cd2610df667b71f1fdfb54e015244ad6f1844b4a
z55fa2bc249b75a5bc0fa0341c38985c6ec6c3aa8ca0e7c6aedb6e2b41ecdfbddfd007c359dd1fd
z4a21f860e1424f808c3c79f40835bd44abfb2cb845d958cbf58cc4b0dd4b469e82e3ec8e26fb00
z28a111694f8fca4b6511118dcb6b1652495df2b46557d71602d88efd437fe92a7530f12a9fb569
z37dbc8a8dec96a720ed25afdc4f9d51293858d4a6838c3428485e93131c12dbd872f73edb2ed6e
z3362c91e54104dde4ca24b89c66f7c9aa0e940b507967da82a070fd4ad36cb76a4dc30338d15ed
zcbe922622d238a4045b486878b8b2f18dfd72af52d235c5be5ec945d0400c74d674ca0c13a4cab
za990743b1eff86ffcf8294b1eb83577a00208592e05425d35d381431ba78101ef5f3894b08378e
ze966d27f07c1c09b51abaf33d61d405e276f53510381d96901acf723b509210fd3e5d0f956b739
z63bb753929796da3df216f19bfbc6ff9d598f3c0dbc5b5e4c7bac125538bb4c496e9205d128751
zd42f102a7a356685bd4552af92a1964a7e3ec0d1882e4c625ccb5cc39ce1529383b9120752430c
z45dbeee9c5a7593932a1fd122853dd3e36d682e1583b6b527f849628ad528f16f328012f235313
z612fc599ba0bf451c130dc06d96d5235643ae0a2557cfb54c000a33bdbdbb1344fade91106d055
z3b920731cfc1f58bd2dd5d943c0edcfcafb86a8d2cba5fe0a15f0384531a3b5fcd9457a620d03c
z090fc9af79b3b271c8c3cdccbb8eb47ed2fe090b321daddc7347e76c8a119abd1157f3054c3ebf
zeb247aac0ce6090648936f5771d98d152b8ae37b7280392b5fcb31e4e751c30fbc2cda08c69a3e
z0b3c294aa870de942dca144b28bdc202edb8eadb3ea5add1453caf22a5ea48bb9520e9fb706b27
zc6a39d938466937aab222ff66479a4a318e7812f900c7d547f8ff0a09b2afb9b70f3968821507e
z6f9bc88187818119767d5beb70c7b6e5a70d3077b101ad340369e8109ac12649dc91ef3939dcf1
z0302d144b275438011b001728227bcadacd4ab57ea28b0400f45d4c81854c95b03a9a4174df905
z1536d2abd0740040cc42e40ad49e8dd03c5fdd4b262cf04db9943445b780a4a8373da549af68f3
zb5832d7f7e9e00f1a675cc0483a18c89cf4f911150350377fb07c69b159cd011534ee6617b6820
z842bb65169f163e83915ec77e25e61ffc9a353f35a0476666a6a1165114dfad7a6161b979cfb5d
z8e506647f3375e9db616993eebc29aa26f82f29659f669a87d92ff88c8c9aced9cda6f25f637a5
z224c9205083f0333074a6ea48a9a850312515e977ea23baa2a841f4e37e995bbdbb607fdcb7e54
z12b919721c5875823b14e2da0ac87494ebdd2614b460cb5d70f6cdd6fe0249400411c73f0acb43
zc74ed64c2d0a48e03bcf7365b47e7c599985b4a91a1cb3da50feee95738eada4a42536e461deba
z66a6f50a913cadf63ea8004b39eadead83ab4a57da3075fea6fa1e5a64d93cecc6ce71e47928c1
zfa7e7d3531c82141da60a170f81f506865533b4cb500cd52cbd22fc338a63eb1c4a139f40f3a3a
z9b1692e8ca0d2fd31d32ade2b944314ab7d96fef4057615ac939827d4ac6dcee3c9c166e53bb7a
z38d1eeb893d77b33af202e8d9729757ee82127da33e9bd478970ec99a5229ed25b648c4477952c
zd4e92f9cfc3a420d11574289709ee1fff0bd40dfb3d0599f7b3b8d4c4c0cf85129430746ca4261
zbad1725cf2a56b2decb3fb98b440781a7682a58c4ce689317a43c38aed6112b839939c9dc69a04
za3a0d7ca16c1f46d594a691b40683172f94502cf0c7e02db238b72bc1c034c2a8319cb3ea0896a
z6df7d0986f5dee4ab3423efd8fa5f806212dbe4755759e8957b5df28c701ab0a5d13c7512cea8b
z1c03431296e1c8d300cc7dff8520482639ed4a5914ebba80e22c5a31d414d4bcd27aa888920932
zfec4cf44ed712990f0c4cc3a674739b13d7a48e95e90512b115c71f9371f09593a7d1dc238bab4
zef371f36a395163713b830d68804b6cf2a239ba8f68c84724d074cefda779a93d0231c07f772a6
z1d3107262e0c9ff37a0a7c38b77985a7e4c8b413a0a446665963907b5c047412b66ef7c7301f09
z34b4a4612e5385d1bdb9616da8fe384d09f1212100ccad712c0a5bf3ea373948dc1a175bbdbe1c
z292ab73c8faaef2c0c12c25853cdae583adbda7a0396663a13351a0cd82a300e939f6ad819c55d
z92c93ee52def457e206eb8eb26eecc2ba8a8f4aaa4286f848fea597a4713eff2885f96d85d944a
z87f95fc51dc52d3aa7df9a6f10e187ea3005ba65f245cc8616f51a05bf372d0dd060dbf12f0383
z5e544d0ec36fb5adfdbbfc74408b19714003bbb3822b630364422af2d466e8f83c0d9430cc5d03
z66cc0753a896fd73b9d244da6fdb3ed4de0bb81db0b001b805094c100d596cf8d52c78dd484fb7
zcd306a63f678ea45a4493ce0dc888fa923941fd3cd0181ffefcef8d9c58884543ec9496a2d19de
z7957a991a6c71ad986d7bdfbcbfd126d8e7c401c500aafcaa29beda922e0a41fb6e6cd0b1eef9a
za1b1f1e7571f8191a15fa10f724d93f266aab5e8a1825589139e0baf23d27bb6242cef81a6e71f
z1194182852d97999fcc72dd6e0363155a455354cb7a3e6bf5aec8c44ac5c036d89bc65921ff572
z0768b5ca4c8077e985e9a27729aca2e9849ebb4d3ef56436f3c44aff1539d03bb0d467e35887b9
z6164143375cd83681ba34917fb5499cd6b7ec71917e5dfba47d5f4e6cb90d2ea458eca06e172b3
zad66a84358c0110d295129a57c4c0a715fab7f74610b33a013028349ba2829d21ef0d91f9b39f9
z503e5ba8c35220dc626697f2c4f9e9ec3b496cba3eb3e019a989f8d62fdb37cb56c72982abb0d4
z91579250edeac0ff2e2241de779d3a653c61a8c8cb5c4a07edaf821cc1c11e41e61ad34a5464d2
z5196358c17719fbb5227964a75b9ca5b59c11bbf41e190003ab3b27a08f67ccc90137c437bee85
zdabcd9f211b777e9b98a6faf54768d138508a8b62cd2168b0b4df357a9620a7d62a6816a5ed6f4
zd02ffaca070762637f5166db7838de15cfea0c826058702a8e6d926188684dbe89c3a17c0c0e9d
z911effa8dc0e98f635ea1ba6d87a1bee64682e5d9dcf8ddc6db58fbe13c439a1451d04077ab79a
zd3e3e7a5b86973137a8b8590dc8a4c818f820b5512ee5481f08b8841945adff81f6d7db763d755
z3c5752a99990c449842471c348eee9c2ca69a6b66e786efa345f6d4298f24382a62b8c7f668e3a
zbb7eb6ffb9d63f317b9621a89caf1ff582f633acd09c783abdcc05bc9d63c17d4e76ca7fd5e55b
zd423de4845c44f27aac30fc82379d77eb754f812d9a010f9e8ac42cc32843b5e4a7a5aa9416126
z33a0ac6c51a824d9af8e2bebd37161e2d75858f75d7990b28fcb3c94900ae47f34e888fe07faa3
z7c09cd6471c5ce134b14a4a6afab1d8a51ba5bc1923dba6c1e692868cabb67ba3e87f65a8a1469
z4eb05ee62b96103fbd84267f84a85470da14c0382aa5e0d8f8ef340b28aa87685a67a8df9ef474
z7f2774c95f96ed36dc0d0c68571d3e02e87c3460f9854ff6e2657962ba65e6f75f408fe88b1cb9
z22b562bdc96add831f3c3fa4adcc7f9ac3bb9af81c555826e185e6018a232f01ae179de4cd109b
zd1a983a17952a8e73f37916c498d14d19d7647c7501fa3935e8cb5d0d49163a8da9a3bf11af796
z5b192d6d3b5477b61c493b9f45ec9e3467dc46b0eeadae88c85db188311b5bb5eca7163b10bf9e
zd7dcf0ad58cac614217c9aa118279e11678074d05f9b9fb65a204ae9f65786fe58517a7f9228fa
zdc62f7f371769dbb803eaf79267f59c6cc863dc92e4ad9e0fb9e842d120f9a6090ed44aa0ae827
zc240abe3cda0eb0137385e615d740e5eaacba3b8b7de604ce7c82ea9221a4d2a533edb8c287a17
ze7b046ce8dad1a7a47d12dbda4c12684f5eaee70ca9a0a7cf2f564717420373d3103de758daa3a
zb1453937973b56a6ef384e8e3518b88571475007616c52b67134675886bbf1d09a6c0b953837a4
zc60734b8d28674957bd57590529b02d97ae49e829d486f6d758ecf31b06328f2fea4a5f6bebac6
z92f43929b2d18d105fe527c5f06d531132993ad625c7319680cde02612c6b2ef358fb4149ca436
z6909afb69d462f2844f688cbe82b45a9a72dc7ed785750aef1c07a50b7eee3e4f0baaf3ffa5bed
zb11563a326d6e379e5564ca10af61715da0c1a446210c565c785d614d4ae95562a78b3daf705fc
zd18b229f484691cadc4a3010e4122ae2c5d6d586237bddd1462db3f3eb28fe2ea8636cd37207c9
za8c53b6103fcaac4e8bad2c61db08d03c8cedcd609c8e89374623f0f3b15eac2d5e153892cf609
z513d0c36a7c4fc475d6ee6126c8040063c31cf4ff2d45d6e02fa9a4b8439066ef7612017f77f08
z33a42dfad7159a7f9faa8760aa1ee78deb1af7fd0822f52f1a0d6ce7d50df656c438d053805461
z8ab749c8effcfff4b954e58f54804188383be21c4ad81611ae7fb0dac00332e2e1a4cef0aa62ef
ze7e234242c58dda8c7b776a83e41dbb03236b0ce3dc87ff17130e1f085b4ef10547c3b5522f6a9
z803946eba4b37f067fec2e7b2fcbde5c7294db8b3444e5b0f95ef21e8e3c74124f4d7c44c637da
z5835ad7034e81ff4858927ab73cfeec341e57a37623c928eba5fd4edfa0803ec6f50984489761d
zfbc6a149a3097c0ef68042261329af19b510db6f20037b4c3a7d49a0d7e352902033c3dec1b72c
z67461ac1ad3bc627be540f680122c686f1da17a1f12c21acac34a535f368d567e61816f1687b9e
z1597ece8e9e2fe3f834d17671881235ad52804cf3eab9f0cea004562303787d23dd8a17a6ebb15
z57172ee06b9bd8ebdb7f5194913a1ec5a85bacd1515be40267c8dd76615c84574d48e87a06b149
z406a9976ab9adc060d2a4d68768bb583bfa2dbefd89a0cf6c3754aae0a6eec7fe18950d3a5492d
z9baee733e414c0bef5030a155777c585ffccee5fd25a92b0cd370b4443695475d5ff8e1b670c44
z69e26fdafa0e6ad9e2cf9cd4a588fbf2a459741cf88d961257deee8202182a874e665d287af2d2
z118ba4758251c4b000b8d2f1ece259a05929fef4562604731d534cc1307e3a4333826d250bdd02
z99083a8525aa89acc54b56215d270e8b18db8b6876edf646dee8c5b5690c36687de9935baaa17f
zb74136184bd43ea7c932140942fc1a4c7cf40d005560dcff1900d9b8933c54ff3bca2a3e7730e0
z24b2d5e80afb9ab7a8a1c5429eda407d1c6e1cec1d88116c9935e9e68de75c05d5bab0732de318
z458c11edcd34cceb08e05faf14c934181ad6c46614cfa81d68c77c9d31f5eebfb11d1a158a4570
z6ad9ee0bb17eec5089c226ef13d78c5d2069f8036a963da4b1a006fb99eccdf60bb4eb7791e990
z7dcbcc11f3ca5c56b7de935a21ac8b5d1fb3b7cdeeed08e6a1f64284f8fce42fe30872d5b2df8b
z880ad4de59ce8ce6eeea34a812639007f86b21f21193f9019d028b3917896d0a3afc3acf7c4b5f
z6cb707d749387cbeaf43345e63ff89344af33322763a3f03e34c38e989fc3f6cdabce7f240154d
zb5fbf5f769bf7216d724b599bb89163dbb40edbded4892c4e8f6400d950343c1cf143c2a6a8d19
zb59e25cff2e0ffdd681968b39b7685f983de2f9a62db36c0ad99e9706b5d8c2ebdad060d739793
zfd9061070e686cf45a11cb9d631ac6dce64d25c3f6ddab2a19a0215362fb86ce4338cc559d37b3
zd2ce47be3e06641b8911033471b630e69c11f0e60ab080123fce1d9671152e5837b5116600db01
z03124892a64c72e1b22dd36cab110909cd30f1fdf7827c6df7448c84750dab2f604e067ffa7812
z80f2b9c53e8c8a003fb29c1d2b45d2ce3d7f053834c1a05716169a2dd5b4585e6a257277db9c2e
z382fc51da72cd9d7e1f7cbeead4b743f7591bc542957ba2b7049d1b2bd543201d5f8635e914921
z8aa3d449995c672a2d52b1988a1eb2c3dc6aef13c068d36a27c8cf7234b41878acb2eeac033118
ze1d3ed1c1c6df0478c229154433009124805affe952f176714c67f6a59f8528a50dbffb41a2180
zbc184c9a345f062b4d886f704aaf9c375448c09519dcfd78f85cc8362ef1648852e388b999db12
z147d4c6e4352ff25f1f6ee0024704da5f5be07236b7468e561965e250cd849658435ab18619d7c
z34c6a172cb57880caa5f8dd5f07b2c7d2e9db7ca6e71a1c922cfa2711e6eaa450b880e2a51531a
z9d8e1b5b9fa80e618394a2c4e023ccff17801e6cf28eb2e8fb90708e03b78d6076b7473a0c3901
z2ed58220328d24d1abea0d511295caf1a16185422002bcd4d769dda7c68fb48d677b2022469c72
z380ff8f244a2e5ced9a7ae085bf1c31002f598b7fa10166d287b7af23426d6fc6d03036f310d84
z60adb916e8124ad62a6348a902e4af5044578ba5f4e11fb46bf60d82d70f7f7db5b50ad612529f
zc6716a6f7ebe77e950b65a055c0973977902eec508fc83a097027b731fbdfcea3b42b00fbc9fc0
z4b4ec7728e9f51444628326184397779339caf0c9b0596d5d423fbb77f83738bc3df86a5a32301
z0804ce92c8b1d402f6227724c80da6597b72beb901af4b064a588870ac0a417f0c4b4ef4c88c04
z5fc861a1a44530d88f2aa08fe676a9be9eb9acde184ecae70409b6c5c7baad1e2abc7c79db596e
z1391cb9604d0763b33ed3c61b72f15c489a9115a5c377f0fcdf9de7aaab3b825ebaa08a9f1bdc5
z759ec30b1c6e85af349a20fcd6e933bba324e32dda1d61637886f279270e1d73f8e3485657e930
z7eba9bb17048de0bcc2b6241f9d16a155b3737e187add1063cbaef15a6f7fb4b83ba0d506bae6e
z38fcfec822aadd79e302be14a196c36f7090b4ffa45f6e6fbb9a84b04376097d51a691925f04b5
zb62bd19df7227105427e1a080909ffa7c84b5c6790c43073cacb93e25589230ac94a812404fb12
z2287b898beb8e7405d7c574f478e6ca28472a60831ba2f39298ddb6ad64a2c83ad7c836fc5922c
z1b3c2839a933e8dbbe7b86ce3f6aea13b83bdfcf970ddc3cac23f21067cfc4aa980501f15fcd9f
z46950451043a8da2b1e945d6b2b9b07d0cbbc60bddb51694a0baf05f342241c3bcd78a6748b6ba
zac4596380b3c252c7c4e03798742792749d9319c3f2022c60c737be71951784f7df04383555cdb
z79cccad056b4bb00a7ba60765c82bd824acb2a8f9316878bf7ef393bc060649dcb1eef4129a29f
z6a94efed98b3ce031cadfd82943e038910c22a8be78298ebf9bb5f013ec070a495239d192a4e01
zcf627edddf03f341b56c497d10f07bc5858185c949a2c8c7a80af9a809e92e7a65b2315b65c4a4
z685118bbf84b5e084a10b07f345db27d698557fa6081b248a4932959c3029ace0daaa2f22e0c91
z934b021d952b6670025c0ce58e7968210856875e9f04e047f7b2d7b18163845b24cb2be7d17558
z76376ac80b7bb7690454ed323810b6b3d18e379d033a7de6dd68a428f4df8ebdda30f67d7613ec
z104c21cfe0cf6bf9584857c8dde7aaa18b79cf0dfb414524f206cfbe9c847cdf9d79c72ef208b2
z85ac83470517d0b7aa2d2a50287a2db71a704e0fe9d754dc6424f68347ef6a72cefe5d90ab2192
zf726aeb16707b14023eeb580a17a5d919460e0746f83de3b546c24d6f83e886a1264dc994eb56e
z35b7724a09d75143e64bc8f578bcdd62b31bf339539f4c8b8ac60257b6fd22fe1e5db324fbb4df
z902aeddf5b1d69ae6962f7612bbb44a0fd72ce81fd35c27d98f8fe5390b1ea3c939b6925b19b44
z084fa36a9ce57d5e7b16223980af6d71dfd0c7ef12d28aef461d9416d705fbcadc4dd04d781bbb
zc94a4ae6c20ffa276ed4035e40d044550ecf2936c3b13905262f710ed56700ffae3a0fc28545d4
zea70aa3d439dd8f376c586db20575fa07da1d0961b02e68a8d731d0dcdc36492553565ada9879f
zda8485aa00fcda9f3307bd1e66967e16ab84b0b84faf8bbec6a6063af706cd1e4d41f3c7fad63b
zfde38e6b7c99ff8e93416ac8da80a9625a7002c6e86efb6db832765a47c8730320f3a214b43794
z12f8c475c4b4ad55d594dff0ada109b1d23dd77aa1ceaa86fd336399a73ed5405dd2b8b574d8ed
z7a4348ac91f6d6d49d4c59c5724fbedf195a63c461d9c6b0813f3778fd42dd66ffae13ece5307c
zaed2a52f18a431aa8a8eb30bb48847bbe238346d591b62a51378f31851750e5e432ef287aa899a
z09af29b91aeb575d80dbec9fb707ee2202456825c8720cf26a12e84f3710ec6d7b1bcec116e263
z81c60511cfa612db738fcb23d970c97332c2c247b8e0d6f6f2fd0086669f6ef5205a3d9f5146bb
z96d638ea17da981ffa86e40807c6010164a1c96a11bee65200f3bfcb63359e6ccbd66a9583de59
zbb0a6ad22b4c820e9e3a1b035658b16814ac24c7288e7199265bf303e73539338ccdf73e21febb
z034ddc467a8d0fc3241e8725c83d7e1e4387493e72b63c7d1b32064d07e9d0c2ffbe60d189f70a
z2187b4eb7733e8e78fdaebff6218360e1afe623a2e374d1ca3fb213746267f4a7ea5c943dd70b7
z9d05e0222f8c2dad4dad8bf0d7d80303a7969e95c897b69c350b3b8c76ae79a567590182ee86a3
zf4f1ce770330a3deab453e9fe8c5c67646534314ef30f2b3cba5e7937743dda86811cfdb53bd02
zd8a1451c3d314328ea80b482b9c019d5e0e0bf818c7162bedcb620b826c88151516a7d901db90e
zbf6364ad07ce9d7056ce09b89705b6be23c70fd641341965b5e9b00561576b08a0a796e2e35e23
zfb2812a5bda232b6b1ef1d7827202c007e29281da63df1eed86385a99922f6de0bd72a4d30661f
zde96bb3d6fed6944682ccba9a1914c647b805b47a13918964fcadca52c090cc491108eee90af94
z287bbbecdb21ef3ae618e5a30a79cf15dfa9df448d65e5af08f0f4acb6d487fa498cd998c8ff6a
z3c7ae7d8fb2679ee43f77af19932cae4b94c01a8d592fea3a42cd35ffbd246cfdc640a739f429c
z64694b73880e0d3f951e169fb9969765156e31fc798fd79ee225cb6b0f6aa7d3007ff7ca6b50be
z7a466c99831cd2572b72f50580b45e7ccab260ee9118f9f29326328f1bb3f4870501bd0e6e3206
z6358ebf64df02f32046643427dd9c638427d40182c0449c27ca360043b852135e1e8da7feafd9e
zc153270af555e7c1cadcc85958c4aa545b1a9d54b260ac093d945b9a727794eec6d815d6626d94
zbc6cd57d98702509f15540aa91efb850b6da4f42d80b99ab536d660bd7829c6d29a7d0ec8a3562
z7f3887a4110981f53fc064b92810dbf63cc5c30e6829624bc4b209bfcb2e3164a3ca85f3a95acb
z45d620d76c9b8faab3c5f93ffdb540bcf985f74dfba86e0a35ca014b0d4833dc750133bc356ac9
z4ea8b8f3b0ff41a8497bcdc702bf6a243b11bc66d6a83bff59bc0c58b304a65d18c46dcf65c426
z6c96e18cea7988c384574ff2d5bafb8ca075bfced1e1eaa72dcd5ce8f9042b35249ff847ae8ca2
z9e75f8113f40b0be5dc776365d5dfe533ba89462a67f7497e157cba2c074a48bf7ffbe38dcba55
zc1b36a935edbc3ead657d584153629c4c7838a5ff6da3ceee460a34baa2a0a559c03a9699a3ae5
z793cecc5d0a0018159a149aea9fde88c3b8b704cad553ef81e6f412f0fd5f633318f06fd8fb186
zbd494ab3076e6732d6fe870a238b23fbbc851051e26f60f6de503d94a7f9cb941156818cc402db
z2caa3a773404cc1fc9827d17a39f5e8b57b97c09e74062cd35dbbb7a521080db9369d086cee94b
z599ca7cad539e73fd2b486c99f332ee0082d0a396fa5d652d362d72dece2e2aa81c4e3e3bd4dfa
z0fcd720d9550672046586ecf117f3f9ad11350a68c9d64a62f2aebc85b44c2bf0a982c8214ab8e
zc81f12e0e59aa84cccfdeb991504f2152e910bbe13321d0120b14c5461f17cbb54de4a48188219
z5bc61256301e116fcb394f0c015fa4d8b3d43d84a1aea2b6231f2928bc312e0cc729eeb2439a75
z943722eedcaddb357672c5f20249ca2001b7888221428d9e1d16e76d095b78b51b607b18fc71fd
z5229d035b7d1e9f594d3764462232f4122afd0247cfd56e2e63c485160fbf7dc251bbe9015013c
zb5a33a250ff0beb6728e1fb5ad9696d173f7f1f966640a83459ba096c40a6554742f17d70e4b0b
z6fb79ad5e1d41d1749dd9a87ae1d95bd6ea46475bb171681436a12ad3ff0f724d1f587b403975c
z2b4016e7d729f6400b11368132b5e255bd4b973ecd2ecc0c618bc8333f7813425115090b709af2
zfc829dabc9a763bbfbf392da4119a6a48a7f1e2104cc3e645917d76e235ea4973052e2cacffa1b
zb0f237d101a1ed4de03b7c529bd3d7d5a303d03df41cf2cc7883d4073d92e4764986f548e34047
z15cd3630aa9342d85844088864b101f747941f89b4c4a9a66e268922f740a232ab7fb994f6fb7a
zd59fb998f8ff61c6fbf453f8ec166b44995ea05adfba1f4de8dbe396c6daf109c3a79d778f4467
ze148a581c770189aa31b203b17c3d0c665c42e8f74717c66a26aed4641524b6cfc606c24084b53
z06831698a91c13a31b13a7a2417bb42cd85999f430bd0c3ed8f825f2e6fd7cecdececbf6840c79
z1d05302b8a162f0114a6c5d7c0eac593d3891375e3497a960149424fddbd004454687d1e1fb372
z4d9539559aa7853e0b5f83edb4c1c6b037db48085a8fbb86470245da2e95d308f429199676be02
zaa59f4773306d9649a70f4bdae0c6b0abd25edce03be42e4fca0106567a75521566ea42e3292f9
z80e8d577843d8892f9203cd69437e9dba36104ead56f59f7044871abddf4155337a3787dfec391
zc51fe8bc80c6866ffda62f95d0f5debd42f45c3b445cd45a45affe93acd7046888cc7f62c3aaae
za746cf05acd45db89647b60085741d06487480f696f6d3f4e280b90f227e2c1bdecffd448befdf
z65ec96850e0270f04b1430f81d8e444999f077f3b7f24a75ff081c1785dd07d810347f2155c1ea
zebd375e0a5ed8f62ce96dcaa90b4e7b326653316053ec325390cd499ed435e5ce7445ebb2825cd
z23fb7b24572c45c23c3c7a9532e4b242b4b61e7506276b5f2411a2c39a9039d20179fb883a03b2
z9b5a8df87615636d8646261221ac8d7fca3aef7970aaec04a3e69b1f3afa655c6f8db0d5936486
zdf3bcb1f4b2b111f33f770f2485ae37a25c79398bf5f20e57676dc02c120c5ff8056ce6ccc2ff7
zc3171c28f058881821d834ecb0153d53e81995c74db1825c36af6b5dbc539039be4fad9e7f1766
ze65bc1a1c0d133f4fa819db9f73ab1314fc9de31e8458f1fd169f67f210a2cff0433dd13c3fd7a
z07ab108fca3b3f548e2b18745083ae175ed0d84bc3b9367cf29c13ccfe6b78ac70b3e4db74ae70
zc7d53ef495730687297ee8aa0f2befd335f7312c266d66929a915ccb960c17a634e022dcfbff17
z5ad3792e2be85e3514ee24d0a14dbb9fbd4938e0d49aadc23f3750f6d5e27962d1edbf08bda3d0
zadc69bf639a5d5c2451a0f614f06bfee3087203a6b2a8f61c419c3433bcdc4a9bfa1314b610f2e
z9aaf76908ca64bad0d7ff5eeca058510f7be38864957322e197832df17b6f16cfe46bca4f0396a
z3ffff345c7230cc86441da07d07c0b808ff8a716543f8e607a92586d597c69abe3546850950330
z640cbb3075114d6d7f632adc84d6bd2640c7ae001b3431e2d283e62ecb817ceb52ebe4ac45ca6b
z01d88b0e58001190de35f964bc347df3a2bdee962efa65b804d8c773190ee3be56f0018262ff2b
z2ae4fd65cc7090826d8e153ccfb629595644284be2535e5ea2b36b4aef3097519b37d397f3b3f8
z3f9d6dafc5e35cbb6ae981efb6ef68120fbae6eaf66a38cfb96cb0308beb1d6682f96f707a87ff
z8a878c1099f1cae6515e04549f48dd038d01ffc0ce89ef73c0f11ce2b83c130cfc7512f46f4a8c
zda0ea38a5f5be9c599d4dcd3d9383e23e48c0f890cc021db9255f2dd5bcf8d1a0f7480c1fecb26
zd468f3df1d62f561910489fa4deaccabd9b8c04e730b8c2262a140d0adc77f868caaa3399b16b5
zb01246b0b7726bae2c96a473f6ef5873000927b7b069f12dc0aa6545c15e8d36d4b4503ef5dc57
za1c0823c3ebcef2329a741538557521c070e5da7e6c5188e10c5e8aaba1d1e8bf3ad75b232db63
z6a5e44555ecb166d29c64101bac0800ac5dc68fec2d048fc41ba94bd13e2f2338fc0aefd786284
zce10fe47280a893f408b216ebaa6add780337bcc67c877dfbab55b70ec8bfe783074c34bf57a99
z1319aef9d98b90adf80c23647e1fc1acf38bc47f1f100f1a614495202d41263ac27de2dbbe765e
zf35d649266b8ccbd617853a640e41e7e182e433322d21e715894a7e69fab7f5390485d9612f219
za5a92f10a2736626e00c9129c45db16f8e06d0d5191b982662b1d3bf8ad08c6afaabf74aa77369
zc63c20b5bbc26e4970a43405eef818e1768beb92e47834b278011c1e0072c0063167ea31568d9b
z7538cd1927ef90254e0f9cb8006c80a6a3001c8e98e5a9455d6003cc5412e7942fa957a2baf9a9
za125b90304ded2d102f0c736902b6ef2c09cd047f904347f4ef632893a93b419d263a1537c65dc
z9aa020b9812fc38a827e5ea2ee04fbb321cb3a5b13d36534c4b22ece089d3ec5bbbe7a6cbdec85
z3847d750107ef6162613d2906cd5f6fb9dbd264ac008f6e1dd30eeed109446951076dec1e6e174
z23f5e69caaef193e2e4660c2e77b2c8dcff41763e0b182126da497880bea9914aaa8e4b40b2c47
z33a46babd762cad72b0a0944cd2f360bce812eff0816ee356f33e425a00b74616f4ac74ababa50
z4bd0fe8adc9afb20005e19e4f3d0a089bd040f8ad0c811bb96f49492ba0f0d0d82608a0f9bdad0
z2fd18f4faaf0ed150c0a5102fe25e6340a277b09141cadd2ecfbb5308e2b4a854b812db4ddae0b
zbe518930a83115b635326049e5631b1207ed4cb0911a3f002da675b3c20fd41b7c3ace9a5f3d13
z1eb1548e9975cebe36b955da7c6fc290c8149531a3893357438dc44f5206d78d3103b1ba995be6
z3408cd7b99388cda3ba26d77c96a61b7a5194d892407ecf39bb64a15cb1738dd6044634af8ea79
zab4850431d29169b2e9ef74da5c5dcec6affaa85e408d9f2c14e24c5b9a8cfa52a73f7ebbad215
z398d7c0af11184d02cced3ca9cf19ab69959f6ca1c98872faa8e3c9edba5e72826fd63f73df558
z7964c49654e89810bdd49fc6a699c2c9538b856147f803cdc84af75e632890ce3b7fd73427e038
z8d7ed4655e2c59c6228a07c9a656725b547cf10ec4586c36cdb07adaf88b88b1a48a167af6c4f0
zca580ae348cfda5894ce77fa21be38b2f04ce517965dac36f8552171456c02ac4db7f207584eb3
z913df1efa92d7fe32fd7afc2b6d949a9f851a2af64f3225243f42e4ca8e5ba79bd2c7b7cc5e36c
z08d217f8f71d998be887dd708de187acdbc6ec05ccdba451c6c74b0388357f1fdae2d4cb05201b
z9f0249caee907a7611a7cb521aab82a5ddefe76240b77f2a48cac33cc405e1d855be8bcbd1d72b
z7fef7c4807dfbbbbef1438a15ff64781921082582a008d39c643d30a7c994f856c9155a1f0b23c
z32f7d4c02ba48176069010e83435ef14d7c6b251b848c02119a19ba0fd7072a4f5978d110b1902
zf09ddf57963112879aac745d1edb5a7d41c394058bb053014236507adc182ce2789ba2edd49a2b
zeb596d308345e5f11c4cd3399eb4cc9bad360fc44c1b43a43afd5afbfb522fb1a62be3c01d89d5
ze6c57d1b9fed0645cc9f2fe296a426bb7af6a516e4e4636c8d3ad6d4da8ccdad78b55a73fd65d7
z9e79980f1a95f6d8b7e268f9ce68bffd8e8f8c472f5c7fa8cad669689d9cdd676adc0741909964
z01edf0b93e2d393e63189779d7c4202c87582f76d28d5b9bd124d9595788f86a14d1e5762c5647
z9143373311ce37bd3be649f50408e4475b424f1d72a979f17cd76357851e14019e75ac76491ea8
z656d9827c92a366bd1819285faae92abade2c3c0bf53194e5d725aae435d4c3b1bd800dc8b5c39
z498d95affd575fd5a69e8414247b85065db69c9da04aa54fb4e69cae4f373dd9572ba3e3fae8bf
z8bedf30873a970cfe80b3d7dc6cc34cee73b9e305e316a9397d26333b44d3c8dd1d28764206854
zf2666aa4fd54a418ee503d04a2b3d8315bb29a5bdd6ee2e46f28c339bea7e60237a3ea9545164d
z8b3d635e63a9ee09f02b54d21d8d55f4458cc4c81b1aeea782c3f6a148a46f89b7d42e814602af
z8f1e81ce0d176ee262fe122c46ba558a6c44df77cca416256ef9a0460258f43e87861912e01b0a
zd8822b52b9e1cbc70a973111a4c9f29014956686bca0bf851f4ec1174f6118d6fdab2c74aea71c
z0df08fcc7bb7b9a0eb50139857ae8a81020d6257a339476cb163f32cea54895d3c3161a8fd3c76
z11d734b9d47d03d53e2631e3f9713e0c5a85a3fc3830974d89be17fe044455bc2879bb77f8c74f
zd7bf34e8ccb5323100996a9e50690b2054dd78b6e7482e15eab06884d8016e2245fb1d294d728d
zb4b9472477cf19be67c0cc218200a1ccedc911340f71eef5e7be854d890214eb77c6491cd41d98
z2d1ff541cc7395c75deb0d619aa45e61d17ac97cb02c816e587a5c2cf4f9b38347ebb14db697ed
zba4c5e2bc96ced9f5e312f618f0f322d2efe7dc253df86e9793fd78b6f9762f9331c4589251fe6
zf0463b7bd46860c1dcefab31534427f6c9287ad4b4d4d15cf0e0fbe9e2b058f6c3f1b80c672878
zce9b641bcb822b45c29e61ba3fccf5466204d5da66c291e22b35e419ebd1ed340c9918c1a98eb4
z163a54ed3e32705bcbfb45a214c1a2c07e167504d88a76231a7db0fe9f8f98909c23bd0e11a33e
z7324bdb578b8e312cda8f40d8c40fb60421af2aa9f38cc83ee53aae0829e8345d0e65bff71cb00
zd60c20220ecab6419c0262aa87de4b0b5003ced27d4505b269da778fc4ee71930f88256a134805
zaefd833e5cb127076b63e19fc76ecc4055ce680c99623731ee93dcdbdec812f269a4daaa7cd676
z59fe92276d4073af0f994af17768da16ada65ce5fa54146694082d63f547ca5ca054acb8c9542d
zb5eb8e6bafe80dd4ddea85ffb6843344d584f4d5d567c8a4f4479cb441c7172c548432add343dd
z2613e6e1c120144ca5642cca09b4bb8d33836981dbf95282abae6992b70e0e7cb0fca2be4d1319
zd753f92c8169aac230d98b95a6635af17d180ff57b90cd29aeec64cc752484df05f4fd09cbb126
z3c36f8f3e8a0f18c5ec8b03e0d740f855fd1475f02fb53bc47ff1127244a221e929cd80322b04a
zc97912b7e984dbadca5ebb8a06c18f8adf7576b8c7d1b7c827c61cab69de8ba084a0461b39e62d
zc5320240a023353dd3c5824f068adbe750602f0ee5da81450620bd896ce157dbc49c14f4301aea
z06f5bd8dfff141016395a1df4f20e7b6b692e7ca937d1c8417eccf4a6dc90fc5b704a8b8aea075
zdd73bf9d9636440c03af80741d1d629dd5a92114c4117b680504c6f157c33007e456b69be17344
z83477d96303220ae02c793346151395a01e52d9dd8685cd0623bc57d18e73a6344b7ee764cab91
zf1ee1a674813a0eb1aa490034ca6627190847d5b6d22db8e3957883fd1ce40a6943781d5c3086e
z482df9c38370b95cb1d88854e7dcff2859f899818e80a05d332a57cad6fae33629eabd421d9c4a
ze657084178f4e2493f50bc71e262a23ebfb0b43637dc9b3846495bc592bfb78b58b1fe7ef4805d
z5f40b02f5b77c1617de55b61754feca13abdf6a29399390102102474abc0e33712aff52d66b91c
zbda6fc98981685d5cbde0ea214d28909a6325b7305aa51a2d0bb2fc3afc89a9de23f15962925f0
zadd9934645dc598393e298df020d5227bee2e58329575b8616c5107e220f3f8f69d0a7f4c75930
z5d9866ddee712366cc145c9ca26ded3a6178916c8286ebb4b6cb552d1495f370fe25b80a7f4da9
z82d32213e3db5ad5cc03a9d318c89150b03e90def739be0c7201943589cad7227aeba6e4405c45
za8c4b83f50ed86f79c51d41693a1902ba33e912c78cc25f642a016a0c9287b255c4b6d8e23cfcd
z1d3e4e8ebf34d59db382acde42bd53db3b4ae1447911c57f21be63b84c235d62c8320cb5d1103f
z4d023c80c3590f88db78ab807a7bc4ea987cf5990b5903df75e66657e665396b824f6193ba12ea
z3a3b91d130f7ae86bad82bb898ef99ddfdf3f214f00de9914ace248ac2b9dc718126edf0357319
z174b0106b31ff8d1bad636859c328b16d0f6e1bcefbbb0a6cc4f883b2ed1f63d5af86e6e962078
zf8e05dd87ff8bcfbe0777747df3a1bcabf490b9cec26acd5058559a5e92533c80b884dfe34bd0a
z0468bb69c03c55ca3aa96c7b722433c65e274ce16019bd39eb235519dd7cd58a9291530f3683cd
z36b77f9a202c775d9af5d67ddbebde3a9ad8ab18438d23b1efc80911e26e9ded3491d0b4655660
z6d28670688517daab233b75ae11a27313e942487108bad79b595d1add86bf8e22e72de36454a18
zdb10e3bfbcec77e88297013c4039ebbe271be753f74a0ffe8feb42c525e9273e7d70a652209768
z813ff96574eb3cb426fb7889b8e8ac8a886a349c1b3298c5fa971977f2ee934971b36c5b3d8756
z571fde9239ad60c67a8f368b09b14691c014ee2e9d2dc497872a66a597e24fcad77e8d5e69a4df
zefb6d07acc18ec6cbf43e89822fb389cd49c0b934f0671c5349fbfacb83910e97e7b8975a0c716
z23e183fa11ba33e9371f02a402db643d1ebbcede17bdb323e7e8702a1c5f772757bf7071cadd11
zfee990374f79adec12fc674ac4982f7c83acd0ab7b1ede921292bbd1daaf9a3750b258b4c21313
z59e66df52f72dd2eaaf9c07929acce76e9a0757703dd0ecb96fb15c02e541cc8e3ea0d55453c7f
z47d1b788f37b29ecfebdaae781d70085125b6dd6b858526fb43080e16225816c5ad42f9717a74d
z76aa5c7e6c14241dd39b82fb0c09d77da1d13d703a0e86b30aeb89553609b05449a4ffc24839be
z6a4fe07c46b815f97623d6c1e958332d3dd449780c752fe4d3e760d10f3cd55d2951f83ec947eb
z80b1a37782117bf9c421cd50bebf0f54d7e15aae718eac1102da181f0557e1fd4707abe5d9cf1d
zb3270a0ab8a987eac845e3c374f983384003c3ce4daa61b582f0e8683c9fe89d5aacf5e125e8cd
zcd0c0dc3c720c962c31fb2cc5335caf489e6d58e713b789752a17fcb32c19bc2d3e8ac8775defe
z8c3474aa43c61ceca4f9dc0a8ad8e63b8272cc2bc5bf0c67c14bd42b6ed1e7f7c403f57fcf2e36
za9dbb646302cfd421e94ef75fb1be68a9b03443dad5c8912c91890ccf758a6234eef0bfcbdf097
zbb320fb5ad00ae8bd8a897a52123b0bb918f70fb384ed4aa910686d59376eb51bad90ea6d7b333
zb27e3268a959990fdd96406963f1976cc12dcc32d82acadef7d78245fefee68519d0811792b8d0
zaea9155a107d89eb274204dbb0fec369ec8efe56c5dab8d071eaf6f87e12b24e9025ffcc12e81f
z02bff668ec1f3f8edac1d0346a64378b27cb7b9e9ce6b351e0b7899a76be757bc3d03bde771be5
z86eff2b93505f130f488d1a11d6d12b2f6e683181f9db7052b2393cfffae904b73117d3be93df4
zbe232fe74702035a16f4c4b6b116cfa86bb3cbe5a65cde00879e9db3e2515866dd613107c5b8fe
zeb150321db3363e5cb194e2d5844652878469751527c7de67c52d2e30e331c703f6b2ef138187d
zbbbe9c5f1fc1ef834fa55398e509bd9fb42420063650f2cc742b416a5341656744fb9aed69f427
zd86b32e184bbedc4236247997c63831c368f9a22c603f0ed5e6601dfe7bb81429da6118823d793
z77ab8e06abd8803c5aed4674ffc559c2792ed072ddf5aaef49b9fae43949a0855ecb1fb9eb01c7
z30b2e7f2533d3d731eb6ecd2284fbbe190f34592e430fc456a3cad6d57d1c9100298b780270dfb
zc8a826d38a8aaab0c7161f4f954f8bab0c64cbfd4ffe51526160497ae8f3ccab6dd49bff521824
z1005df4106468ceb6ddb4eec73207e19b91225b33ebc4d212557b207fbeba0d047276aa996f314
zee7946ea7d98e3624a3d05a791f2f8b86b0228afdfb783acc6421602a0ed238da16ecb2c580788
z163e65188acf452a40ee3af9671501d0c56f3bd307cbdcce36d81dbba81c3816c1542f80221605
z596da2ecc36b697dfa6e9b1e8bc4ea623d1ae41384574d952f3d69109361e871b6a7b07f9755c5
z19ea0927071ffd3dacc4c4ed3a80a5469f5258af371b244477ea65bf58ecb3975fbe93148312df
z757d835892566cd703c622f126ad5fe517b858bd4eb91a84c3cf4004f55e79cc662cd180dddcfa
z4cd9ce79d5f1846c8a5261f11a391dfee8d3d7832b73b7a7a937c7671d0f506e9af74b426d159f
z35a98c66c2c047680d4068841b97978147cf0f558ed88f6dad744ec5587c721de8d978a2f7589a
z58429f194f0cecbcbba00e55bcacc6b56758806a3b99af75b0dbfdfc3b3ab666fc3a9b8bc2a5e1
z2aa62fbf6bcbc28b9659724c0ab88b7f4d6859329d8b265604b97529c46dfa5d5a209bc4857d4b
zfb670fd8e86dbb7e9f5bcfa8123dfad48f591fb98841082d492e5aad8c5cabe2def637bb3d411b
z678307f39bdab68cc37dc3d45c0f76fafc1ea8b999729992e5ac9bc86ec623956f90727b13376d
z523fd27f940787b6f82bd7f83d09d160e3f039fd4420c44d575c2b5bff6bd5a35793cf7bce0bdf
z9a03bbd7fd6617e7c79b2a20b4771ad35e1ebb07fae82d993ae7f2bdfb2715c2d8bb1085a76cc2
z1a2feb5fe9cea7f01252c26607b99d88db7371f2274ded7b0ffd64b602cd21886fb2e2cac8850e
zb1aadde845b03ac9ebcf5663719a73346a32fb3f87ce0e5d6f9cd9035d44b17ddd3fa7f660f32c
ze416b2b1d962b784e75fa32d9c2f5f89b8615aec2fd474393efcd22982588f58fa4a37beeae2c0
z145b61937818bb330c494b86ed176bdbfd9bb99a3577814302f3bd3ba9e2b3e03eba3cb843d5e7
z2f51958eb3928f6fabde7f606db931c8845ba051e573287392fe6bc754d10b50c3e83cec33d0bd
z0caafa33f82cde9db1c14c0967168d650b5c0f08247ed8f6f990699b93e8da51becaeb2c009a5f
z4bd149275f1dbdb1e31889d9aab51e1d1219022d8ac4bcc47282241516fbc897bbf785de4b7ec4
z2521fa46e389b3e2c94b8e048ed29cc12096c6eb4ce2016c02af7d937ea9d94ca114d51f000577
z3d95e66315c79e2797cd3ebb99e87e0ac5d04a335be97c0db5e40c45fc107769166a1eefa7247e
z23b48f73be667e6991d85936b7644824f4ef2c851ef54dcb521994e021b9bdea0812e82b1b04ab
za9d759fbbf3d72c36ba9bc3d1c347a14e90978da08ac315a766a4419fe8097b5e2680e36fb5615
zd346a7530bbc8097ca0d62e59da7de7b8efa217bb9ae9866634b84e628d47f2a17111be6795c6b
z851ae85cb56ec8798c85bc10590eae682a58147be9a55f217b59a1e4a91bce55c8564222d40da6
zd3058ea01ecae403a310430f8e02737f53c00db1c3a23af2b52cbb3e1c0430d348b6677dd1f20c
z09b1ff55e6a05eff6594e61094238fcba2a66576698dc0617c4254029baae08ec9c043de5b79b1
z94f9030949fa5ef6f63f584e78952a9b0c1dff5047cc884a0e883311790409a02cae35b6dc3187
zed68273c1960ef91cbb41b76569183353f886f39258d1772ddfb0c9f5aa6d242e50eadd3c23291
z9d9760d565660c2af1374ad1414a03a0a051475c2ee0db87a0d137ee7afd24ce84e12cf79c43e6
z9be666cbf744c52726974ff4dae03475268286df676cb51b0328a03631f5ffd829970e071eaf97
zc21ae5692d03645ae6c6c5f8ef39a281778d712b7ae1019f06ff6306c9b852ab1b4560f8d62c3b
zb76f44f6c02af268c8d37b289a75053e1bb19a291098cb015ee0877d6e0601546f9e7817bee135
zd885de1fa3ed47f61b410d97079cf57db5b965a0616f4983a6f3743b1e6bc4219611baed934c34
zdbe9a72869213c51e4ab33538f359f3a16c4a4e11e117723090f8ab63e7f3e62c77dc9e719c93f
z4a0d86761c1577fb5bc930547a1594fb98190530ef539d80327b639905202cf67c84c6e42df096
ze1c8fbe5bded144cad0db16f133e63c42a2c7410b4031992bdeade01bb902363f8d89b484cd65d
zf90a254e6737309e21e9d31a8b96dbe627e32ec327b77a51ea6ed243b2613beedf7f1d72bdcf27
zc8457336c36dba45ced6c29eec920fdd063e74b1f8d2673045c2abbf73a8ab808a726629ba896c
z427a39367f942a37a72024aacfbfb650b958c690df93ac370187f7d11c4ea34fd9b5acbfb695cf
z57b2663f0815f872412f5003dca9b6f5ddff50d9f174dcfe480f71de169a50c1ba8d2412b3bd3d
zeb0ddab1b7b63b50f5bcc30544888479f8c6755ee80a37004d624bbe64488166ca937f751c02f0
z72029fe3111f6ae573fe745d12c3c570649ee74b698f52f57fd15c5827e2eb67ef816d1f20aae4
z6175030fb1a53fd7bb62b9ec4364c61d026a1b4d296f303f06e521b15d366cdbb19dc53cfc5ba3
z24f896f90aa6c0073936c5880a49684a57614326027823ff3d946f4eea99afc104fbf05f6919f5
z6249574c51a6cc57f93141594944ad1f343ee0b00e66c16a31a5dda67265246e66d76060338467
zd96213c85060c9a0ec21542f9cecdca937aafcfc1d43ab60aec085da515e4473899b4e446db8c5
z7795da77b7177f43c6ff2f7151c287a81c9776ed63e7e5733e84226704c137235c2b8e276a358f
z1d5c3eb45ece33efe6584eadb00d5ebcf23ad011fd4e7003dde8f749254cee50a6c3ef3d52ae15
zc85400d960af21f4ad122b033c21c5d161d1ab4412a479dca5604aed68e593c91889d61e1bb0c7
z1f8540e3ed2909117a754fd617cc96e21894b3057663b65cd9fd8c1f803fbc59304c863a3cac46
zb73c1c49c23aef6bb409bd1178293e59ec29e3ee628eea2572bd47d10bce00de38f119b08b3a4e
z9dbf7940d1b120ba28892778e1d917d7b29dac15ade510cc602153a32e4fa54bd105b1672ade90
zcaf3965439b99404a6ebf5d9d62bff90a086f822bca251e4fdaf997515414aa70ab906b4bde0d9
z5f8f17a948863ea50321f8158c2d17a4cb93c471007278c124eab11b9fee679bf9ad419cdcbb55
zb866ef0d6c5c7661455a7d2dbeed93655100a37c294792a8f1e7ef0cad42cae424f2d2c1bd8bd9
z6a847f004bb90cb59eb85aaee49fad9f2f66548cb832e5209e559ff8abb70960f31d914ba0cf0a
zea3c59268166359fc5b457025f73c26df2bbfa76115604278972af85a58d48aaed7750b2ac675a
zd8ec9cf9fe6ad7544f290c44410beb2c8af6ade5c2e58785b13f1c53290df7db66db03fddb3417
z9d9583507291b6a25ae30f8a6776c53aa0a5ea01d8a011a3bdf908f6db7b190cd0e84fa640b223
zc3881755777c5b78e89bfc409ba95a674d211980a02fc5162ee743fcb05f55a0e2a932d4a41782
z76d10e06bffd8b56a279d24ed1240956d57f2dd45b61f04c1c82dc62ae055550a8c4e3d4426845
z73e80820cad98ddc95b14caba6c632d59fc3023c13dab0cdf757e2778647aae670d6a8957be46a
z5496e87a396ca50b2fa80d09d9c93403dd241a0ddf7900f062d99594159a63d53bdb048aae4779
zbbd1b4fb74f37f1bcf91d23f34a6213608e95de453dc2dee69fce46bc23155a05d9941a7059179
zfa969c6e18c92b487bee1de7e40abfe9f778a0ed9597744d888b253382b6355412555853e03dc4
z569d3223b68e37c11337dfccf86eaf42f7abef218afe7328d5988095623bc0c4c1e30827cf8dd6
z1d3fe7110c5ab99c7d8c35e874c8d105461f8fad708cf325e69c9209c2f7a4f659b0de38c769fb
zea9f922d5a60472e975ca1408149acfd107dc15ccf7538e4c75c203dc03c43a315b3fe33493e11
z465a4fdba415e24ee22ab335d3a79bc4cb317f9ed8b79f40f065841fc2d066301455502f5a9f08
z626c05e100f699a21735eff18d20671b1b077ee664f86a65d6cc4da803d9e51073166ca697ae71
za73477455d8c88a7de81a5381db71813056d401634d4d19c8a335bd77f60750d71baf7a1025fb4
zec2b3fcb182532c659dd328c31749cbd3c56acbd06d702b612495ba64771ad7f118ed30589d78e
z640ce8effa44bf6f4283d1172ff645612c2983d840cb4f415236fa58f5a1fb1aba6252c612772a
z99e48ee040f9a25b29f10d2e4ff2fb4e0dca219ef1ddd69337422d10a541e2fad50bda5e5292e6
z6de3986ed441f6602eb87108f9026f24867b68dd9dbde2fa5d87f2983995b969330853eec7d99b
za92e3225f1cbbda21bfd926bc9f26af827aa17f31282210f593f6d5826f2f348bf1e2e1b05362c
z8e8a5e57721d9646cdf849326ba51b5b8ef6fb140b2c88a2c681e225e0803524493ea8b14669a4
z787e3a550755e770af33adcfce9fffdcc3dda3d9b7a3ec3662ce0063f811618c8c78ac11c3db3d
ze8034fd7030cd34d2922633f3258dba9ba9bd2985ac3f8c02cb783caecf217c08af93a9d5515ba
z88b603ddd0e99d23f34aabf1dfe3c5cad88a08b5d4f2e9986ff4305676f73ebe4f2301db721bbe
ze0b5c19ced2c64a4ca7d543d0335326636fdf2a6a24cfc5fbb5c09aeac206099dafa8fbeb9e5e5
zd898807827b81deffad9da1fba4c848e0b77c24998b05ac3b7ffa0b1fd9a0bfc565e1e8f8b3694
z69c056bf4a2f4266be6d2b736eefde1b16da6a3cea914763635ba91dcfb72d9d2b6b95e3f212be
z7a137cb06a5b85f17970cae6f18214659ed6227a3e2d9c161829122f48443861f48c4f67a076a8
z00fa48941672633b95c928fd7a3c853d9da39b006acd40cc8fc54d4dcc7d2dbde60c86016f3981
z677e9081aa224234c4f5a04480c807c5559b808ce779c1d9706a6df0cea93b46b602f5f05ef4b0
z70d5d8276596682d378836da74d044f04d6a088f99aef39468be99adc1d80c5ac62d466ab7c32a
zeca465ab755ed1ff918af83cb8d49f38aec120beb182bd04e76440c46a5572d2ce367fc90f9683
z6f3bbf0294fb8584a55d98b4f9261fa486209373c369ad3c126aadb943d71af1217b91735bbc4d
zdcdf0b5af0fd0837e2d309f049dcd5200d9f9d7dcf37c9e7275faa7ed70cb6ce8fc34f2c5a4f55
za7abaa363c17ebc3199c6ca0679f3ffa84387cd8d15d32f3a1dc141f7bd02ece0901100c0cd74f
z39d109509c249d8ab73500a2acfce3451613a9f396b71a077a79ce7f48aeee9040a6fe09c189d4
zba8f5fc985cf9012a1e9c1f446fec2e19fe97cad9ece78c8bcfcfc97a809eaca86f428adc23dfd
zed079ddf69da6119833b4ea8130e72c07230a7516e5843e08ba62c0f410ff6a8e0aaaf18cab7d4
z2f1960626cbbbbf1e48232573b4c3c1d2f2bebd383547e9df442ce0455735619f0c788c23047a4
z2584d3856c98bf9f22f24867cd7d69127539d0905c94186e5cc6e5eee2f9cb59cdc745bcff00ca
z25440e53dda69dab0580f60783f18fbba2a39ec51a6d40205d44849265a9708fcd9ea181e2b80f
z527602b9e894d0fa9492ff8ca2ecda607acc5c74865fb1080e3880a945d7d2319be5f636a1e2da
z272c920d016aa11da81b0d1b42bc2f41f35385ef693334a25b855df599abe8e1a97dca9eabb7d5
zfdf80e6787daebfaec1cfe9f58c4e0109dcd6e0297a7d7839d6664b9059d4c8c4a651c6b68bc99
zfb809bdd7736da2c8bc4bdaf735b06a4bc2cecc36623797ce47911c6ba4aaaf990d0df762656dc
z70c87981cbe8c6cbbda2e0d966aed0e02fead68dd94bb6e5a784b125f5cf78c9a68cdb6a622a3c
z99312879fb4cb19504ce27ec83f1058089a4dca28c3a3c907aeef4a60dfb519868bbf195cdf099
zd2c53f403541c11ea6d9977cf6dfaa28e6926f0c27b3bbb6e3d93198d9b6cf2a0f7d8f5693be8c
z8f6de1fcd87635cb949b341500de9a9cbb419c4ac5cc3b770250dc35d341b037429e47d7b73d44
z6cd0d98488ff74ac5f2ff64a137ae3f2c08d94a15f89b86c3bbce6961bc6b49972216edb68d40e
zf9a153efeb89b50a57705947f2d52efc35059806622d0bc5350aedbc260594eb517ed807f4f141
zb07f96e1eb905ddd4253c8a41984e7819bfd20791f50e7c0772b50591db43297dabde2c2c263bd
z58d510f054113f69a5fd804b62cc99da9c35a2d1dff4e5e183ab8b2de906cbb7a7554debf318af
zeb35fad7e4435ed787fd1bb989907049e46bd44b74e50439d4c20ba87e99ab2080fedb9da302e7
z4314f0fdabf72b597bbfd1be3a3cb171991141e2d4bfce8cfa442e653c01516a307be0ce0c2579
z260272b34220803128fd7d7e0c7998164586145090ae686727bb2252debdd803693b98fb18e722
z9a27051270e05654ba66a9a80d0dc47c6db88af1e52071127acbcf9ec00bffa89d238dbef11c28
zb8760057705c86312ab1e453083d85274e836bd92fefddbd59faf723f50f914583255be49bff5d
zfbe9249acfb994b04f45eb800a0b2c09328717eb16f85e41f744f0cdf9366b83ea2751166ee110
z7a9e7b3d10dfe5cb93de6a523d413d7ce51a83b0561541a1aa375c166c25697072d053bfd14a1a
zae36ed765e80494f6751acc1b9396cc5bda511c68d5e25c99639d486bb8cc386711ea1e0d27ce7
zb76c8eae71d032fc4a7e519f4cbc0fca542860683cae3dde2fade0de69008ac1a7058b7b00a8ea
z402a14cd6fcf4311e383f408297d3df4189328e654fa9ec975efdc938f98f2e043b3d06b6379a3
zed648b88102a31b4eaddfeadd8635d64a50db0e9df10211a5d1c08fedfe120e530e4710b20e640
z8d4457b1d011ad98028470412493a37fd630bfa914116d64fec619d1403d086b7847c66441e66b
z3d78fad86debb1d700288efd9aeacbbfa35184cebcd06772119d78143182e58695c0a672975cac
z103b58cf6d2e9dfbe32e123f6178fac4da19a9fa909e647db722dbbab56bfca00d94b630dbeed0
ze878cdf621a2c7f16d8f42257bf15549cd922ce4e882ddd64b63be1bc7a06252d8bc2dcff6ce37
z8f7104368bf48f4a31144a3e20b0ff400bcd64520bdeee62132f297614c6b7fdaa16455a087c8d
z7fce515be8e3d0dc42cc2a62b74cc7242c77ee409c9318d377958ff881d6ddae56f01fbfd26e27
z3946c0ea8676d1d30d95c17c37b9b54f4f07139f6685226645bb62d3179d8b49cbf378f79355a5
z550d6580d5179659fe6b3180c6b4133154f4d65ee3020cb177b71a5052c429ded3be175bdbf062
z8ad24b1b06b5f86658ee789ae71d284fc350a8c261e8542591e279db7c4c0bd245d2aeaf964873
zc34ed7fd3a214874ce053839ab19de663fa835a211dd9ddf8eec5b24a023be93409c2909f8c185
z69450e9a47f38ac3bda77f649954071122192af0ffccebe3ac08c9620462f13f0375a6fe864105
z1fcc7abff0c1c7761edbecb2bb5228e9067ea2139c366d6b36ad2c6b39c08da3447962e032050b
z55de4dc4756a9dfaf32e5632694a94dd4640de5c9c3fd865a9dcbc7b3f283cfcf91e75d547e262
z1f2efa984e076d3b410a3e1803cb280e53ef1debe5bc8e14882adfb1e38b2ab3b9840629185eac
ze8034daacd921d3ba06a72513230c28950d6000e329e6a76f3d2d6288e5cdd63160993b658b65d
z1cb397bb240b589412884d1e098ce282a686718922c13351d78dc4655c3dfd5b7952cbeee354b3
zfc8109d24fb3c1e815cd91d24f9bf3fad0f6f440c1bae818dadbcd95155d30fad51f6ce1ca2996
z2c51a9006143b827409f1e56bb7e047e2c33019ab8c576dbd45c5943c4da06ce2ab36496d1e8a7
zb7caa824a5eca5dc9797f70197895e53376a40b91d6f076e4611812d7666f8c3b64570336c7bac
z6470403676e031434626b96165ad195ee419086a9c36373772da37929e74dac0fb73a9ae7bfc79
zf288523ff736c8ddb3e1888fc5d27f68e572bd5ef036593bcdc62bd63a9e299546501577226ec3
z2b30ff9ca545c72078101470ff2c4d1f4b1c8ce5bb51d95554005db3b1e7e38db158d143c10b0f
z15fa7f272b972847a9ada9cfdc6350f2105397d79dbdfb5a11b55bc66c0a03c817e0ac2e7a22ef
z1a23a4bb210bd4ba69bf8e467431826fa07bef8d6dd8ee22fbe17537784d52f6b520047260c6e9
z2fd7f62c9b00d5c3e39df6e41ad6544544fc3f1110a9325040de3a76afffc3b3bb6dbece367c24
zd811272b42a7f5e6ba88ba214ecd8ed2fc93a29c33c70469a9fd8bf8f19171898fa18d2da8b6bb
z2c0a7392f3acec595ab22d8e353894ffd25dcb0a411f087a4059b6699c365412cf314d1849fb18
z681e55a5bb5647c323b4593d3913e72806ffe7b5e333a8d2289b4c72cb10390607c7fe30220e1c
z2f07c874ea8a3a6bbfa6e081139773b1e3cb0eac984fd3ecf171285e6df39082d21879bc385de1
zb8b5f93c183bcbcb0d35d1b7c0de9acc7dbc7d87165cdf964ae72847e83ba384e5575e4da0dbe3
zfffaf1635f3808ec5d6325ddf039a17a0af959963b972ed8dd72ec06c87b97ea1fa395fce5b3f3
z875f6716eb866e10123265f6ca4661038700e6a5058420a1f92d0cd9f3a6b191e1278c933c464a
z83bdb4063e2b77f598d8f30997826932c5ac851ade2a7082ec300d99e41d6e5552261ad8a2aefe
z31aff6409e8a9c73a829be0088963cee8b9cec082e372a93982d1cb127c92d349400ac7325f4af
z44ac803aa81d54adee4b11af7446cc9aa479fc0b553be0063aca727ab08771cc472b31b7b0dd82
z242d8d22189cae47e721f3cc7be4e82dd7ae29c4643563b65fdb5ea3ae9fdaa919bcedf6703696
z894537b7844dea6c75312cbef674306ea1518d36e60117953619b8766590a2fe9a0bae56ed71c9
z380b4d854a6e7cd624da5049401daecc04880ae278bef3620599280726d9f076e2137f2d2997aa
z0a1b8d516ebbe81c72f62314e645a03ec12f835e9af85f9ee77e3af2288c1a32068e319b447b81
z5239590905bfb80b90d8c3c933d98891386ba6b4f5d48b688dd1162e3abdbf81945d16a62b581a
z0931e5a73167dc55f6d8d941c0151d99f1893009750e0ab90e2f1cedc772a7583fc9f11ddeaa12
zed108c94ec8d61bfe179339725840a2a1a67b28721dbcce5364741c909391f36b98fdf00688d19
z87b3e4217bd0dd73297368f64701c3ac466229e1cb862b53ff2760d4a7049bae410375f31c6f7a
ze5ef24572c9a40ba37fd8ab46955ed30bd975a639f469cbb2a87ec41ae687e3317a36c5cbb6c68
z9a1f66a367ebb72957c3ab166bad18b2916742ab33b4e517095863d029a6df30de3cca7af2a4f7
ze699470dd5f2a54780f4dd8c68ec2cf3187b0f24c1d185521a42290e3741e0636f18809b3e4cc3
z365c523009588872cb67f876f8cf6b18cd148188086a736d8776b71df77415caaa465999103678
zba540efd8d643d37795a0dd26673e3d271690151338807871fb5ea138cb5c94183a605974b05a7
ze91421c6c5a695c088282f38c350671663d7a4c61ada1b93067e5ec5195007ae9ff988b63eea33
z731e94695490816c74fa040e30d07ddb0c329d2f555abcc1583ffc292209a77032d1aabebbdc4e
zf72acb5ebdd093104d91f74565b306b4214e7ed9374633458fe7af2f23260461dd21616d397cd3
z44da36a37ae823af847aed71f8e6f350476cd228362027e65d4abef252e6107757b3ac88011ad5
za0a336af7342cc61fc1257820389992b5b95d3dad9305de28b443c85964dc52abcef2f22e5913d
zb3289f88812045b6073ae55c1a147b581c38b637b8f130b68501408adeb4b56b21f1bad7c79376
z0668080949b31b6454eaa36f93208f7077510ab565a242d6b18f066fcb88ac0f8a4ce87b277144
z93518b83f5f8a6299e8a416b5c7a5c37440a6b4f448b86ae78da633f2538230a3aa450ad93ec05
z9d31b2b1b189bcb94e6d16b954baa1f2c9cae5ae9a3f0b1e7ece747960d6f9699e13f04a592b91
z264450e19ab01d598a668b6995c714dfb8c55f0d7ffa5ec8ebdc42657642cd664c53f1ad0d5c8e
ze97ee16eca1c589dd47c7583eb757bb279fd69d54c49a69940f4fac04f39eee64ab7ff5c1bd01c
z7c4b3189e5aacadc46f1c1413b154dc7716259038f33d7226306686e3b7d24188f1f3fb57d68ed
z8912a2411729c3588ffdcd402877a76eee0c886c8b9969eca30a209f58f920ed7824e347643e1e
z06eda41770c96048bc95a73f0a3f92135cfb0c28e8c7dd6db65f0933973f0d768a4f635c21acf8
zf38d71ba6639c8634a3ed2697e1b008b0d0c6fac8a90719e9f61798cdc6a1d93fffd33781641bc
z899eadf2bcdf52b015d33d050f08a391e0012e9fd6e4660be13718077a340c29ed5dd20b3ccde1
z56950627e878cc6df143cc806b330f6b996efcb10b92256a59eda0aa25524d8baa1359fe13fda7
zd4c2fcd9e45adf3079876bc1559c7e1002775f0843064d4e3bdcd1d8280e5650ad2aa61018c98b
z08e7acaa3b37a7cc6c9d153732410125df92abb73a530a026aa81918ff49767622f0b85248f1da
zdbe52aa46c7b662bcb07ee079fcac837820c19a837c73dc6192ea8866c99450e6875c3c8af2a2e
z71d58f590acde142a0d1e617df883abebbd02532ca6798f550ffafdd6f366d85fdc0713040cd0f
z519347b0e4067fe6ce63b679053a53869d73ce9b34849b81721b4700d9a7838c88fe42b0bd82dc
z3b6b1d726a1d6b1ab69f53c49da3fc3449cd496c8ec00f36eec7dec620fafbcf09854c4d6bbcae
z174dc977e7a6fb98a02f360d974d70db51a474fe50b14e98ff5a7834e8dcde9e73e5df198268cd
z6ee22aee302373a8750cf233de98c0f3762605332504f51e4142f5d7bd29bd7c17034d7f223604
z43b91bbe7b8752b54291e46b61e53ea2d4b7f36e796ce3ea7e05cbe2b049d1f2ebcfac0c45001c
zfccc8ff780ddd1f5273bc478c86073cd4e4f37e22816fc744113498b1a83a10c8208f213d464eb
z7146c1f38a70e73903af456d89d618bc187b1119ecc71c7ff870370af2611913e2694228b924ec
zd72e85c1702139af511ba9b6c240412823dc39e7f8e3d10f0a346c498d3846bbc3f2012684d72d
zbbcade675dff6a98f6ba0c154161c9ae1ff510927059a90d7770a2a5c11ad58ffa3153f574a1e9
z5ae626389bc54a29ecff3ef2ca933127a226d7942cc99627b0a907529c95881803443b07235b68
zb966f93e540421159c7130e6564ede9bd88a0e6065abaf6681c18f841e10a28f50d10228a17be4
ze958afa3f98303900ddc458395d1cb1fe745dab7a4c37a16cb6bfba4f0d211cae6d41746c2678b
zd42d450dcc0e60a345e14142535e934d24b77c10218771872b2f6fb80ac4b6b9eb20cee88ee38b
z6338e1d3c059af6a7ad1d4681a2236723597bf7a36a20f3d5356078882f1b8f5bb2985242f7a77
z99d2628b610b34715dcda263ba89a4f8bec5b923d0ea94d0d8a6721ad298b276b38398e7ada88f
za7952243d9a8b2203f6bf5476d062eac21187dc4c76346ca5461faa7c6c4a150dd09d8ee69a467
z07efaadf10de1200742a99b0ac37eeb4d7a10ff31f929c961062473d6e4e1e5bd5ff55b6b94867
z7916bc7d48a286968dec686646177979f0d3bc5763d31962bfde81dc567b8c6dad565b0dfedfaf
zbaeba2f7702ffd60043119f26fb7513b51600beaac01885d47ec7496f5faa1761665c44b9227c3
z6631004cb92ea71ddd9ae61146af14faa54fbe779f19f5ea463fa6df787c5092ed892ff09f4946
z4e25353425f28a15725c1da09ea10b798a305cc5e2ea003eb01bdfdd5c3ca59bd363b443ad6ebf
za7d86ce4e994ec0895747ce8a07631affdc7bf414cf214090dfd5cf3726caa9d9a5e04e36db733
zc7c1b69d30acd3d4b1f48e0440babd19ddaa6b9a53a25ece190bc25c5c74fd529e2621dfb7bce5
zf0ed5cc5cf908000d2b4cd5bba10a7ef5597cfe68a501c1650ff985f665aa1a9cef4a3d3dd17f0
z698c766c8b534d57f8f9a87d518857ebf1223c94d125826c0a0c288ffca48262043a07a7f64b17
z478e29b93229ca63f48c905d5394a7c44e2f3e1ffdb80d5933ea59b883c2ab517481a0f48a5e9a
zd11340d8020d4201533d4dfd0403e50b0240493bb562a249d60cbf9a7d84e2a296ed1c1848f674
z88f61cf834adf7ebf706ab31e8132882b296e5edef6620bbd1e62cb71f7605b1390d708928e308
z20059fe27ff2acbffbbab715264679b50faae4b016cf586eb8999e30aea85a8395597909bd85b9
zec96530e901bfc92f6fa89aac35508d6e96e175e918debb41f67f2ecd8665323c7096f441fba8c
z30e6e04477086ee1f0ec50e0ad747075070bce528cde286a03971d498b5dedc08f798b07d6827d
zb3a713d1d50756a2dff154943ce85e340d94e595cc5b6fae79a2941e81cca6e8bc65c04a70a786
zead2c15bfb771261921706050b31e08bfcaad0751e0575717c13b64028e72ab18c3d007d2f2063
z082053adf2bd661963cb123c452c3c2ad5e6afb7b48c56339df40a6805c6a77935a6ac723e96be
z806bec4751baaaf8a94e13d26e9197a5f88eca8f9515e7c1993bf0613d9b418decef703a508bbb
z0b349ccaf0f7b801a218ff3cfa3d1c7e6bd83c05ab2acb623193dbda460ac249ef20e23fa230db
zdf8c82ae1a3c356cd3217cb086a4451bfbbbbbb5e210550c6a6c8938714bf41686afee8917bf33
z5f2e90f69d3afc3c6e15f5bccce5abfd3a6652deca459885c34020e612b6bfa18ce8352da1f490
z751cdf5c533a529978fb89cc63a3f0a9764d2d727d59ba32a8082e5fc93f3a2c0f65e15a656c71
z28a706772ae789981a10f05bdabf47a441ffbd33079132a7e4c50cead61e780064887d0d703012
zb85188f9a5529c9aac6514e6f6fc7905036a0c9f48544f29d421e2c6e19ff6ebba109c13e17360
z94aa732d391c98e300a4e063569b643b2f747b32cf13b022c0301bb221abe0ac402d5a37adc02f
z41368ed5b5a81107bdf20a21756aede014912c8b761a57b8cec3083527bdfa263507ce0a6213c9
z31b502d8e1bb9c015a3c39ae121722fe80b944eb90192351b2be51526617c7102b8bc98a487920
ze996322fb890be3c6bef23a664db1444dad1deb391332f1c249f13ae3172fe163bcd4ae5fd1a29
z87a018cf43d28bfb6db45ff9b2311f03f76a10802cf1d1a9a4702781e1908f8b9435c8414d4fd7
z3a6e31bda504e0baf34ecb0a4625e4137a4de89596292488bd997f659e65518e21e0114fc3fe81
z441ed46999204316268751ee18421b946e6d816a3922359d02f0571fc7c8f02a5f3534b7908c0e
zf2fd082e5ae27babd519518981838e645473c214525305b58e44f06ef2f0af688582b47c655317
z69cb472366615ceb7222944b3864a2e42be91350a9f50290f591b5fea1c3c4fd943238e09db76c
z0647770160828e26628e01cc201550cf4fd6130a4e160102a702ed329a24107b0e193c66571ecf
z0d3b0145740b48bdb5e7b8ddf019a394c3586b7b2a430f7c5574191d37af95a044181f8ef8cfb6
z24b9301f08d9a3925c775276e027fb2721360e252eb37d8d73dbe93b3253a1b7b97260004854d1
z23de23a52e234e6977576bf6b5ccca748e2057ab0f88d20ecc9885115a82c8a10f3d7bca7834d6
z6f1e137a75889e35db927c4be37bb845c650ef960758c6075953d266a45e938e3eb1c4f89e7b6e
z31a9f601f07bebce16982ed9b5061e84a501670ec6e6c6f75d8df1a31a651d7762f9b0e5902b76
z70959774ddff3d0c87be2dd104889aa3ce8c815ffd723bb5fb9cf39222bd29947e7a26ac69ae00
zb5af78e1bbe135c3b0d031c2e274edbb10293d9ba5c72871dee77515cefabc744cc4cc5ec00c2a
zb1412c3d8c8282cd2990971dd087f86651d567380f6097eeb389592743a0f2d98785393f5cd971
z6a292ba7bec7ccb834817e9599583d8739a2571aa2f8fd60bce53e2bd70640dca4f3c06fc2bfc1
z02214a05a972372abb77aa4e6ad46392c405da4ed1463984a3fdf77ba81afe7017818926e2f25a
z1b181a447f29f8652e71e405de4d0c2b098eb4b8e2c6b0fe3c457b4109bee035524f135ae3ba94
zdfeeb2572695774cb1f22f49a3ede15b56f3337c8fb04653703a2eccaa623fa8014710e52b7070
z9248c618a1cef399e6071f910bd85ab8e9e2e59061bc8ebff030150633da1ed8b217535f1d4952
z8548bfaabc0b5edf7a71819df782d5f51dc76f7ff989831bed8047863c04660da8d7350c926a01
zd84d370c6116a2bd366d25eba302a8ed415a5fc7bb72bd0a05dc951ce9616e4690011363bc848a
zec6d7f9f3a266b2e307de17a330f2c8c7c12ea5cd81f4e004a86a3800a82fa878c06d78de277db
zd1464d503f768a2a0945e7954652971a60fb1e41815bcad05076728f90e5a42eff272bc17fbd38
z392eb6e856b90064a2ee7f7b35e8a76e8d5d2a84ac72eebc429b957394c00bebb977ef0a9adef4
z9bd9d80d55da742be6d804d137095ea0c41c831c3865e627bc614047775231cbfe791754e5d859
za9a48d79a8893cd2a037bb47ccd5d9dc649d53cb4ef3201667ee9baa1541618a3a412f8aec9721
z6096005b80a2228adeea324bc4d2b200e7159029f502eb64b9b99cdfd35d35c16a61a3de9eb47b
z4a90b811f789fb80eed24e33f4a9242e3da0b8529e09c8597da8543838163df661de75c0bbfcff
zf66da8750cf9fbeebe8854fcf7876b65f3d5cdb559eda12a266a3c51b87effd20d4b56a73c187a
z7d102749d506ab1ea1feaa00fa58b2a2423deb9b1f4ba8ebc320bf3ca8e555636baf45c86c1d13
zdab4eaeae8269057cd363121ddb3c6240530372cda9329c36531771b52b4146a5847840ef62e6a
z17a16f0006067894ebb06eb4ea3f5f47e80a41e49f2d006b01a33b65fcf7d11c95e93f8bec7e52
z89a01efbfb71a175a1ccbf6aad0504bf24fe794ce877874450e24b8342fe29123d04a9217fb9b6
z2458432a260ecf19ef56b77caf5e157db938d3c0bf174c010a872b468642c6d9f547996839d7f7
zb30a8da9dc11c71d1c65b3eb65b7de50b87d52bd3f1848b2b98357781688a30fe1e2f816ff7827
z9fe41da3e56b0a92f904d63d7a8e98550d864091cf498bed13e3ecd16ba825b180a1878bea69d8
z0df5fb3540abfbe4f807d86cc71f8e761f0e22e9286e7cd150b26edc96c261e7161c500135ff31
zc3c3c070bff61d82b22fd282ec5869d13cc358df4beab1fe5d2ce87cf5f6bf2abeddd7a474654a
z607100a0a1fc3e606a9679da6c3196feb2138298aab1e4e9648bea2f7bfdc15a2dbd6e6d07d71f
zf8446ec5e59cb40a3a0e45ae07c6766d14e55b85571d8c25adff29e3159bd84d30d9d5714bb688
z0650fac4ab7105dccfa80a1bcf2aee5d6ba9d162a29a321b89374a026849f7b59610cf57bb4fd5
z607347482825d47da1e853536a5ce2dbe30a452561cb248f4d8e3c1c6806d237b330ba39db4673
za440e9212b4429ac2d7baaf96d8616c78bfb2e8580ccff0982d832b40118b6bcb46bcd468a0f62
z1e12555468b3945030e13bc84f5044f7ae3115796948cc92ef7c8f343753fb4a99ce4c2e4d65ea
zf403a9d64a975c74b0ccd3f554164ffcd15cf878b559f029d9d7fca8370a08fba3fe48dcf2fdb6
zf6431d405a3ac133fad72cfbb50743fb1fc7a1d03c7ed75a941ec66ca4f9020687e96101ed6c48
zf3931624cba90134fa5368dbfd33f816b38c0b96fcf8aba99b23ba016f1f7f096cbcf235ddaa01
z61bf11ec509aa9de5fa88173448eca965e6b262b0708349d964dc5f0d5622dd597044198eecde0
zc569aa8c985d0b66df7b5c9a8af1c3e11e2351b06676e133ee210a72064b3ed70ae58b6ae67ea8
z82104b9715c9615d34696e0a75d16a435f00086f9d53a782cf7270668b1309332879eb456de5c2
zdda7eb0686ee860338952fc5838d96c9fc1477d661cd031c2799633db689c5b6f93ec39007fa72
z0dc5de28deb4eafc1a9c4f660322c09a150112506577bd1e5ae60923e304c9b1fd59491039545c
z43913eb7b4edd0ba62aa5984f0a672174328f681f1c2ee221cadcad74f24550f31484d1f4a39bc
ze20426058eb2f3d6cc2c1a9a7c150b169436c4c699b66c93c6a988ae150ac316bf8d14687cc2cf
zc21905d011e71bd72830ef0974c6896f2d9ab564668cd9c6180320b0c7ae552e93694989e83e42
z8d273def0904bc5296fb3b125ad397cb95f7a477a480938cb3becea50d0a32c94b03c8c311c1cd
z4b9fb06cfd9e66415c6ad4ba08bf4ef05aef9abc51baf1fe6c38c5022c5e9bd2ba9f8bd533f575
z5b1bc2af9b78415d303ee59012107200e28ec9555797074f9cbe288d5f1d3ad01a80be16746c5c
zf56aac1629e476c167ca803d671414cda380466c000534f60aeaa1f361083dd11163959c305e31
zb601cd0f911589851d570ca59438951ca830e7a9b492c697702dcfa9b9ccd854c776cb2b599981
z46093c7fb5f7856e81fa91a9399741bae91b3b3c5ed43b56f05b62071ecc2448b6505dd96398c0
z54937c062bb8dc80a2e0e9120e86948e7c7ecd925166152cfae1364e6cbd2303a04e4f5570d91a
ze80135658179dc5c44ebef94e637044de48caa91410f6a93993cb1bcfd56f2f43c5df5aafacac8
z4a2b6c0933466a07da01e577cf61ff54514ca6bddf8847cc8e3352f4681075ca99cd0c8f5cd5c4
zc6455032cf65de3180ae1f08f6404613c4505866571ae779fb70a66ed5df1dfe138f6b9f3eae30
z5c28487be6d5ebd8d41cba1022e77c124fbcfd0aa0d66d29bf23f824fdbeb5565f10b55b4446be
zc49a8ee56a6957ee7968d8ab81f07fc72fb8c7f56244a47b1594f95aea4b786c8eae140223736d
zab432c67f14b29e9f8ffce50a956fb5423e1fa02b5e1cac235aa2bebb8c663319c3828fdc31888
z9394957b1e4c94eafe6693f961269aa2b642316a4bbc4f0620729b04a2d2340f903ae8708dee1a
z19972bbb08b96560164dc4efbd5d4423afe9a4c5422d953f63a91a7e996da7c12621e7f9521375
z589bd48f9437b71324421297c5b6d758403b2c4051ad6ef17b055c86b5c111e163a04d02e105a8
z07932f9347619fd3a0b4305f844ad51d0eeb230c6765e98922af4fab23296bda5e01f75909c2d6
zc34fbb87864abefb34227890cd103332e0ac45f601227e3a0f47c5fad0bb5f18a94cd7967c2166
zc2bc7efa0b535a51551fcbba029d33e1f30395e805f6cd79488b460f061dd452c21f30ecc09a9a
z27b70fda5de2c35fd46aebb332415823528d002ed4bed97bd833b342fc08c68cbfe349828bf594
zf8fefec8e0f8388d7590b43180ea9ce2a9049b7766a8756a654e01998819c516379014d7435891
z5798a85add68d452aaa704b275a9f3c5cce51e75dcb16d8a3053e8c67c66fc1a3e9cece633a4c2
zd1f5f9e42398935f86425322590f247a2cef7085b196e60966424072a8572b1e935086d90e53f4
ze7769ddd70cbcf9374acbc10d991b0ade530c70398e7ae381b596f0ee10adedcbc382e64f77e30
zde09ff4742d67132f9c05407a9de18ac3f2a164f1dadcf1cd16cb06a3fba020c2334771a026e16
zec78b987fe587acd9a34309af3b32ff124e0f351b996a758da7bbb10a5798f112f9bb17818fad9
z99deb29f4dec83666de7d6e2d06400733610040085216d3214fdbad0269bc71e2ca9e0932336df
z2ad67bc621f58ea2a34a8d573212e3de9611c022d83e91b10ce60822aa72be220e576b643d2130
z8123b7069d44dcfdb1afcf604e5cc8fda5174d630fc8b1fcd82d18b31b68180482376a58cce267
z973de1cf8178c6225d56f7f7fc198eda38778f4daaa98965365b9d07f12b572a9584ea873df60b
z82aee00b2c2e552b847b9f64fa602773ace55d4ac3a00d0d056c23a2b5f210f1646d7ceb723012
z0052f04f7c0d80d863a4df020e24ee6f6aa63f45e829a6d8cd8b41b7396635662f4fd8492d0dc6
z588cc196dc119784b5333e8f65e6a40b872009ae9130b9b64d0d692ca6529eb3f61fb1209ab8d8
ze8e13ae7714621f69e04b62bf5622277f43ca5aa20c51f22d33a11ace6d299d6408a56c0456fa5
z3638c148898959b2bb387e21cedddc25b35b73d5f537add29c7e1f71cc07080111de5b9dacb143
z6bc9b425de427922824a894aa65501ef1b0ab8f7080214f42dcc8f47bc1a230337628edefb6456
zb3e5e2c3ced067369ac21b1be169f0e0d7d26f66355d0aeb781bf4c63e9c939e617b239da82662
z26723de9a54fcdb9e2f4daf695439d890f34283aeb5f69ebc25f5422ba3bb060dca1969565876f
zb05fcf20a7bf7e88ca6159492032031bd7674411a463ae61e4343854460677d2b27f44aeeb3c0a
z512260f1d80f6fb9b417f28601063823423c84736e1f58c4b779c3768d17ecead659b0fbbbc7e9
zabd397862694c752fe1b7f54f4010597c8fbf52542780bf90c68cc1965e18011e6faab2039fb16
zccfda8c8451fd309766cdaa211e0d0bff48911ef6b8cfabdffc63b134d26593ad628890b8782d0
z4e2e5ad46d51f2d2340d8d56942d5b41812b63eeb95eb46cd2d698d4cde738db08433d92caf269
zebc88dad19624aed1c4b174325755acef53114c9db64a542d529f79fade255f0f616fe80b7d55b
z5a1c6c72f87f3a9df528cd9fa971c14ab7005ef9c7da70e1d0906ee6a1ccafb0f4814c95a76223
zeefffc6e6abf678fcbe1d6f8990a33932a8b841323bfb7454c2ef8401382c0f8718f2f7a39f221
z8ecf24ec66ad3b8182ffca0c45fec57806d2693952078e3d94674ef7d8fb558bebf6a34a516b92
z172776bade484535bbc91bd4ea8aa0b38cae38e2d47277efacbdb50dca5b60f0114a55342081ab
z05a4ae97e73028d9149721480747149dd18b9645d13e4e6621be123e6303f3c8d04e75b8684109
za3a64f91ec4cd3435e25eddc20dada31ca3ece30672b587b7114b1c20215d93f0fd97314d1649a
zfac77f33ba71580f159ea8f1d1500c8308aa6e2a0ccf8b1bb1e8b49b83246f4c2e1d1b6d791fa3
z1051263c696d143fd0cd64e8942203d67850950d2f8beaf8758daae06b4bb7af1349ffca14b9ed
z2d2689ab7cfb147ba70e12c79019f04b6820af0a0958a8c93233dd5421f13dcff512765d08e2f3
z35f1aafa961fa40cb6cc92f2d251394b47468b4d5d972e7a1efadd734b025e4781a45a27e61776
zed809de0787b584087cde7f1df8991f3718d3135db139d65bc53a7050f0efe19d7061f9ba44d84
z97b69dff4cd958f2747acd5ba69ab12da5e0bdc4abdc2964653f8bec3fa8cf6f3dafa464210e54
z860f235029aeec20f96e496d5f66082a6f742ffaf7dbeea5a807093aa1295d0ca341f66b3da563
zcf470b482598e234145c6a922634015bcc258ab232c68e473bea1151742f2799b53863c6654d3d
z14444ab38a483745f35534edd554475e5554abd9db310a64027e16ba4c207a46e489ee4871cefc
zd15ac1075fda752a3ad7abde4b2ad7bcc7f2bd33f73848982e656a36ba1ad05df817478da4badc
zbfbdd7c3d93d0806c2a2ddc9c9d9fd536ac4d289579826f2d45276ac1f4f276ef65888d386cf80
z144f0cdce6e6d502cf6ff33656ab2823f2d329cf787e2dc3bb8b49fadfe5db40e60d118030cc29
zd71a950913357119ac7c01dc68887d33d9b6930f7e348ccbd847b7c330e850cf9a03566962188d
zd281535e14ac6f7f61705351db20cd4b39156df2963dad625a3086a3378c0df22095b8dfbf6949
zb6637fc2ebde2a40011fdd8738e49d94d8598fce9f129458563d06a1ea43faa5c10745b158449f
z0b2736aa4f23f9f07bc2f6c74825b55f47cad23b1be90f21b2d490a264cd2cbd48f7899a9055c5
zc0ed742460c01fa2a6c4780bfb76d98dbf31625bfb8a7d6579f0179cfdf4889e92431cbf3a9e9a
zc49ea3ea0008faddc7629fa3c909fe128af9acb724fdf8591e8b07f32a5147f33e31162a5be23c
z6bc8cd88c7c2b03a83b6284bbc680b3e7d2eb1d54c44135772be249c64ee8fbca0645d9aa354a5
z4cab70fb2a0e8975d1790dbd6268c84b80bbb0efe2a47bea1f3e466ca954cb5bca89115d9722c4
zbb34f2107e1710598e3ae9a8cc96c9e495f0b09db014dd8425548e27e1f60a4c2beaa01960d785
zf1994cefba30e5c037a30218b2af4201967af172ba1e6ae72d2967959dc4bd2f1d1e135b3ade0c
zac35eb40c83e7083f544d18305d1aeac0d7ec0a2331481a154135cd88c989e75a7be2c50aa4146
z25fa9c7be119b517c5617415908860b26952fda6b3b5ba70785e89443dbe450a38d524f7d79845
zaf8096389cdc3d462c01b0b04de7fecd8bca0f1bc49e28615ff4044664bc45ea17bfc655ae39c7
z242f0eb9b7b6010431d920ffbb87154113ed3d3125713e7b19c22abac3460508d2443d25f713a9
z4a742cb5c79d42fc7c33f2ec3133668fa777d1c76965ba38f54fd3283135656f16946cf2c70ba8
z101a53af82d7406a5fb8a019820e0186466450abe64ed5beed5e2e72a902a725d93293d6c87f23
z54aa6fcd1baa9594a274b9e9273eeccaa08b2dfd238934a4048826c99fc5a4bc7ed6d3e078771a
z5b404b9e62b51de0729d00a9a6b6bf07c8c2c3355be9e572cbcb822b41ce55f4c240f114374b6a
zc6aedc637ba808bdf1d30b035e746cb2250a59f66608738ebffbdeb66254b71d93908e78a0f951
z679167dec85036bcec912e7925a0b73671169eb6be48effa34e519e11ba06022550073d389de0a
z630ad393659617e1020aa600eb298ada313c7100d1cc237d02ed826c134431bc0c4eafd3c9ca67
zd1b14746fb72bb62e14ca0d33a3f1330b49b2d3ea5d1977c87aa5e7a4043ba7657ae30698d17fa
zac972983ecb4d05d9bce74bfb31fe6045ea2f2112db4c0ab83265d0f811ab73e2b640e123dc6bb
z1926a9f90060b5940bee001773c64a5b79c433a00ed4cd51fc459ac21238dbb72e2d748b55b993
zefe1e16cd35ad9d460b5d039a4a689dde842544a11916368598b275f410427404a606dcb0f6fa0
zed07dab0c9d8163dda6781f6443179d9d6ec52ec1da56dadd3570f83a5f1cdf0a6b98da90beb76
z92612d7d28ea44d24ce9e15accf6804d3caaba33dd29f7a938679c4088807b226b216855d8d803
z0db5466124e88808eff0ce8da541a879047de8f28cdeb376a14fd2f76c6b1eb3b5cf608a4af22b
z63ae0d1ce0eb5eb3605b976b5f1f5b64dff486532b36638f37c3d2ecf191c40157be3dd2f8290e
zda1776f1a1eb6070ae268aae47cb7890637dbb38f7e232b1a3ee87c418f1e9aa4ed46d5b1dbd47
z2d32a937c2fe98bc3aa5d75d9adc918953380652a50ebbf418b9f566c57023b119624e802dd450
zfae4d56341f2a827fc8f4084c3dc2fd0273753be57c5a86f892e4b21ed76e058be2002a5411671
z4fc90bf25114b6b52fc9bd2fa90584bb9be6c42a165023fd553334160978f6d9dde634c3fb1320
z6befc4e143a4365f1b211a15179ea549b23287f5208ad7ac759cfe01022685f8769b0b8fcff4f9
z02b7dccbf783e47d3c8ee43997ae99eca204325f843bb6f732a66d35e15faaba952654b97bb858
z775cf8c7527411da5282af1c8c0a4630361fe70c54cc2df7aacc28c5bc8ca2c41865a0c377fcef
z317752dfe17d3a0e5ccb127d2ca72f8553db82db842334a8869b7ceec24a610b7879d363798291
z8f5a83c9d9830e311ccd570b6f5b0be980ee0e7b0fd6ebd2cb1ca0f7dc81938b93efdc2d3702e5
z8b4bd1c46cabd7d0fe6449b486d890069c35fa226e61caec742543c45a7f1deb8f02a40c237891
z27092c56df0948c5aac45afb14621385fd6c461064a039374f46cd08b09a7feae49a6648c4ea34
zbe05e6e52bf5977bfd1bc48cbc324d5d8a6e9036e98a52937b024dc1edfaa4663182d02c3b53dd
z429c2127901bf7ae814b91e9ed97ebd26cb9131914f107d3685a3581861cc12013c0f72b2211ff
zd46514c01beb64318847149b478ac8bd40b2cdfb63938f04080dbf7219ebfc6702211706fa03ce
z0bb7e45167788ecf9d143db13757ae0f56c318393efa182ab3e5b85273206de716778e9075de53
zd1483d5656b7b9ed7a011d883a6b3ed15720553156ad6033ea0ab6faebe9166c6eadbf94bf3960
z42eb9dc5e7018bd3e844505d69240a256b2898df8ebbcb87287baf0fe3f72889b83443d02efc05
zd67f25b03a56f6838aa85b7c4ceb9dcea41c98750ce7e4ee197c6a4a4c37e1e9c7a4e486e0a168
z55a140101fe3d66dc0857e3f80cd243982568aa98ef945b2ab86e0113f4b7511d12d6a6d810621
zd8f2c063b3a293af05b9abbb01c2243f3a49226b2c81ed4e36de930a4795327a2b6db70c4bb218
z41894e7ed4d6418fe1563d404480da5064465184deb30c89c0453849501ee8af2a00048bbf0569
z6ee96cfc72e3e73c907e530a0fe360f9f7593218846c4cef7b0e409899ca80bb8548df1f0f2e17
z0b0f586a645d10b28abc6bdb163bacdaccb20b092f3b8af70445a91c2291279d1b6ecf5ad6d079
z1546223a7fb6c4eceeb37b9c19b6e5ce2eb221e78d1cfb0df56cae2c6296062b570db59f2d690d
zdb0a539c4bb5e36f1dbbb77e8c1679a6ed965a3ed9384c48593bc7c2b6294ba474359129a7d015
z59c39460bbd1278f00156239076ff53b4db29fea7c708a6da9d94c1241fe800a3fb259dd57fbfa
z73d9120574d5d6b70c9412664b9ee43fa7dd73bf5bef34f0c64b6c2840c889929534eb67cec6fd
z460bbb62c05a0afb2f20fd97981392165ef1aa86868b6c4ecdae92b047d088abf0fe892965bcc5
z01cac662a3c47d3daefc823501ff9c0a4e3248378838d89921b129922e420cece2287830f14fd7
z3ba0a1ca438970a06ddfef0d10be13e44a0c8b968181f4e764bb967c4702e4039f9edcab12409c
z10a978169fd26e190776fcdff2ab9da2ca6ae3b268ed34990f2de3848d92d9a9cb7ffb54a17cc6
z7e887113e923fd4e7c96114edcb472f9919cc6bebdad43e78f18e0a49cf7acd8a7f2cb81bdf9ce
z7c1a95520796086dbe96fbeb19e26e93cbfb8773dadb839260f152c8fb47e3c30f2f9a7186a28a
z89ba298626ff3467480790e36b3d98def8c79051ce138a34ecf180c1d23242fa9ec64cc1da71fc
z46a21f58f63cd28569826b293425d225a39411e922e17ef3a5abb556cab11f6e4c06079b410eca
z98407bcdfa088110b732a5af526ef697836b6bf37c09dda179c59df94252bf0ee7d32b5917d212
zd166fad74c2fc67a034901d5809098332513244385c49677ef262a74d1958f14ff6eb121f0a217
z97d5eb9b9356e2cbae1deee2b4add88ca9e7cf343ed32c1074d051033fa0d36ccac369242d32ea
zd5cbdef87ba1b8f10ae730b2d1bb3302d01d43f14bce0d49dbd390873706dc4c9da1c3a9b9e483
z198af8c0f0f86fd5271d80c6bbd51c8af30f677bba471a9995386e07e831dfbf5d6150add791a1
z5e8972c5819835589fb73e780525f71f043bd5927f85b0e13f602917b704cb21ad43f05ef0d487
z832bb3a02ba14f90b09ba646a25d7ca705bb35d5bbf328cd1756256bcec112df89a1f097313aa6
z0b08d04ca28214af47c5b826c11c07064baa7e4e65af486c947999b0f4bda681aaf9f7353fc11d
zedd415852593cd3be2285744cd66602bf7107d140cf40cde24dca07347912d22c77e6a7444577f
z0be6e7c7152ee0094725a6387ce28152bc31d0a62e9b7b356c2cc72efd05f69f6e2ac1ac181895
z05ff6ab81e5fda294a1a788a8847759a5f0f90eb5b8be9e9f49f802aa3e2025ff8762c7ac0f255
z3dc5b7c451946e257aab0b73598e7375d67b3acd9bcb0afc56bf5cf0e663cc3b18b27b9ecc3f43
zf5bc6f40c8de3548456ca0cea72073ca2ce14620b5020436d720c7d3d7682a70908f78624ee043
z0d07badd8ee078e1ebcb67de45ea71e23871f18b77970227eea6293d8eb95821b20b6318ed93d2
z9b9179ad9bc48dd76471ed6cbc2c58a9e3d294e04fa0ab3d1124f111c21b4998fe059c477ce2b6
z2318ced7936446d79a39de87dbe32a971c65a6aec71412ef4bad16af8a13011dee01b6110c2052
zf53255a0c65642293f8750cd7d3a9dc4a6c070d247af1b2b8bd997d68bb29632ccc7d55a582acb
zd6e7c682fc43aa8b7b468204ff6ead9ffaf64cb99c5da9ae97a8ec7f098fb36c3d9ed6081044d4
zd4ce4b8d048914a77e360219d1491c5b4b2f481922578f98f3e5be63c5c629cbaf96ea1fecb21f
z7d4143707f55b6cf208aed667de0c569d39ea6a1e4d8dc9d47f910c4606c3e2eeed94032c29c06
zeb8fdb6fef943421970e4750f03a689994c071dd0c5661e4f62c537ac05c6c454be95e2f9b8f1f
z32b4bdb7f9c4f8de893ba98a5da5c8fc6181e5c8a1fe887b59edc95360938ec5cdc181d903e428
z1fa9d7eed8f2f72f2518f472de0e40c6589e327b131f464c449932812a8347237431d1d273551e
za1b93c78fb3fcf11167a0e71539406e1c93134d1110723f4e3160f3d514f4df6e2229a061468cc
ze4b108c1187d9f1dd340cf1aa8b60e3f3481fd058996cccc564b15b2688d0703b8378fc147dedf
z9a9d111122b5567236a2e2883de70d2a271f19244af9cc37cc37a89c60df255750e5d3565e7075
z1c2a035fcc63ec7fd64d793f8279538b61b9f6bc585678f1ba7fdd7c25e29d1d9a4246347f89b1
z1eeb6faee6ed56f512542f5753dd36a8fc20a6bf4b819e91d1e4ed6769ee6e81b30c656d4deef5
z030cc35cdc91d3d3c67c9a8701f9958a4abe14418663f5ab90078c3a5f7ac3b168ef67ff843a34
zada0a654bc53f75c9187e2a0f1ab89db3695df73c144e9860a3cdd1caeb41fee14eba8957ca98f
z9bb715638a9dc64298d6f55b7185c91026e383399966f2334421d110894badadf1a8e98df47098
zd50167f86683553a1898aced55cc5273b3ace5f937cfb5b95a33e5de613c623ab15eceec86c787
zaf8aabdf7a22667829216d16c6c0bfbfa1b069f3aa628a5b1a53145026f23f20a13d664cb9ce43
z12b84be184b41d8c922b378e8378ef4c9bcd3deeaf0d06183c5f680e64ca8165cb99eda82a18e4
zd7192881bbecc416bae4aa83dc530e7a6544024f41cb724f5251300000bccdb40d80f4ad334568
zd15b49304ac746778acce71158e85cdcf5a9ff6c1ca43b4dc82b3b5ea50a5056ec241567b8a29b
z37f02fc95fa7f9019c63f8f51baa8634cb93a188dd656e11f9aa5ea47d56921b03bf26c4ea0670
z2a37c3413d4fd6683299b538b08473db804fa9daf85c621324fb0b869ff98b51641722d59d1b23
z7fe6af82184de0117d4971b5004a25715159ae4361f30319e772450e232c2b4df9995faaf94237
za1dcb62e84239c144ec2361e468359405ee7520f2fa206d033e2cf97198007d268f9401fc771bc
z8304865de2f5aa347b9387c43ab16cc4fa501524c43940c6938b98ee53bb562e3ca45322a3f808
z80d775679e50e7590b89b038981bdf73d118b5fcf8e8757b0aa5fbfbbcbbaf21241b2ff1fe7482
z058bedaaea2b75bf8544c380f4f2b29c4c5fbc000eaab4a3f513e54ae51d0f52aa12c4f247d3f3
zad8e7772dce671570e5a6418f21f209b028e2d493cb96f114b95164c49ad525d6dbada51d271b2
zbdd35b8bc74dc88f3c996bf2139acef56dcd006d78ae5346bcfda7cc97d56711976b282382da18
zbf14e273a4bf0c1be6b84fdee912a4b94b196846375423ae9b0340f55b9d93f4f290740947d547
z5386065b77b86b1f87f2ea5b9c64f629630e785fda926d0388e8147a869fd1038344b926a333ae
z0fa7b8fd3e2aa0d6442fcdb8635b63d5dbb5d13bf07252b757a9de496f2c257f424429953cc9ba
z3f9a51b7f1c261c1002a368c06ca1bef407c5a55caeb19de909894cbdb8cfc35b3f578456bac06
ze70df1121e13dcc8ed0d6a404eb7f77a1a4721d51b94ff9f44d305be4310f3c7b6a4755a9bc8d0
zc0a9d041b2b95aee7defdcce187723c71628da1278cb1794c77292414c00a53873b26d2e24233e
zd91f651dfb13d94db29a54e6934994c0e1edd256a7ed8d332d2ba23accb1eb37fb95527414656b
z5c0076ef2c7c3bf39361764638c0092e060de41e32cb9b0cbf78f3acadc8ad0a766dd7ba020a8e
z261731141ca1d3a89ef2e43e1e2d6af5660451f4ea5d32ea8267f7aefb3627e0d8dc3d06bd1b91
z0675a8c17c15ff542aa18b41a4b4de705b4f2af8da5db1310507d4c66a73fd43cb20cbbdc2bb16
z799fb75634ea364b994f7f8e5ac18aa1bb013f0305e8278ce64d8fe20d84d34cc9d8140b1ee3b9
zfef463ea5228360554a8bd3d7a8f75a926aa8bc12f2ec5faa097a83bd89b477f3fab26efceca59
z0f039a77bb027e30aee56b54e57092f692a42a4328199809b6df77dfc5270bdca14b436e09fb7e
z7f491380971f16925662ba964d48b0a24113da6b55c32378c53ce5727ff3d270c43701e4ee2a39
z49b9f10f0314b5b11e60356777c02041e86c5ffd0b952439c9890108d165ff4a6098d8542dc46b
z7cf6d605f656d11c915792075ce7d62f475ccd831df2e703c01260ace6ca489510daa86e5422de
zc7f88777bf26710c010a39073833f0f2fec744ac6afa13da3b73e489259eeb035c9c0608a77bfc
zf1f7cf7305e33592e84b6b08315a4874e8f3f5be5b6aa6848f0161f58bc1c239a5737c6a986bc8
z1ba6369cde385f4605e5053434793496c095c1d00af33f1030100f9d1eb165d348bdc279df44de
z3923cc1e47753649f07f36f6d3e443633b2ac8a6b49e5512c810deb034a7b89589b9c87b094c0e
zf4ed89fc50198d0dcffc026f9562a8ac7b85e932f7931e203f002a289add60fb2f28a9a7039ecd
zea03f251156e8fc8a56b139495ae34f03daa7a8874a36396d88f20154aaff7fa398e1fd1628a68
z5687d549bd5ca262f8258bc9e386acabca620b946a2e62a29a3b9509a69ab489e25f4307e85fd3
z740ce9400f075296f9f37334dec468c9ae6e5aa4ffa50128b1274f4d6480fc1c4509cab0949160
zc603cf74e93be4557e891fa5ef2c02db8071ab4f185e727f5ed28c36997b7106cbcd2cfb329eb2
z1e5996453c5ebba797e77fd28903f34bafe4bd27e4029195fa5547f29797b25c87daa617540dcf
z32bf9467ad3aeb4e1e7dd9ab011bafa80f446aa9494891e07480e63b478ee4528fddc987302ad3
z75efbb6d5ad5e8350756aa328454854287f0c978e93a2f623a56511c73573d72a9e700be9c116b
z61d1492c81d726d5f044021e205a71e3518faeb0a0d58e2b4d0dd74047a8fe8258821e7f3bf4d0
ze278002bf0b564e5acf84b43bde4c95adc4d18fb14941cde7089d832bfa439659fc43798b8f476
z08c855445af129cdb5bc6095b44c3f8d48aa44f8fc7350aa1e79b8d00ee7c4254594bc399ff093
zc1a914092ae4a9b00e4f28546f7d57ae54deabaa32663ca619ef3fb876738887d44460adc23b5f
z70965eea3fd261cde884970df817c5258e351b67f8c7290264c616f037ef848b88a8b59c961175
z6855a34a5afb16f18e7d91e0caf19822386e90097e1cb92a9407ba0fc980c3c8effc0c04ee9beb
zea1d5ce7ec3c20a99841bf4c3bc536cc034c8fad5415c788f8914e9113451336171b329668b23f
z09b7f768fb800a58654faf2a2b4735cf853e081661ca1204484ccc8c4f2489b429231dc37d28c4
za2d6c569946a89df7b89166564166ab064342c4a165bc24c96756b462666e25266851e006f6aa1
z7a6d9d148c054a3eb910978732151166efb502b2bdf43f4c8d76390d76d96a6e442df4ff1b31b7
z8ed1bcfe21bd31ad5b08aec603c0cdb988e73e0f73937626de608d3ad0a61210f20fe06604d4ad
z922f1b8d59f989a1bda3b045d38f5f62b978c064e2b5c87fcf18761e51b182fd7fc1e4ec53c5e7
z77734359fcf4cb7acb31e87ae972a00ef2e91b62d5a6e454d5cd58e3e975874246472dfcf3f0d7
z21a724f0e8ec27f61997d364d3ef34fdb35fefcaeb9940a656f4f1a4c137537e8fb9a371090b6c
zd64107ba80abd08212d7a4f483f73ffb8a6d4973096468c15286049c6ea8e4a1571140a527fb14
z18b83b527cef5962d9156ad28ee47dea289aebccd146e8cfa2979bcdd61243eaa87fe2f11eaf78
z3eb052c66c90b69f999761b0f54811e859c57513194edc107a74eda0a4049cb08820407d06c12b
za43ad9dfb6e3a8dccf5dfd6309af238e589698833ad6a9f71d4acdbb92cf7bead620764c456624
zd6d909863ecf59aa41e29d7112c1384d2f2bd9e38e6a45dd7c484c3eb19224129f2b56413eee7d
ze3018de1d71f12048b87096fe4239fd4977c2ffad3f6757e9df7d1508ff44f8aa17bd7b9000a4d
zeb3a27fe9ea858fa309d167099b87357d6c2d7a550bd0aa4fcc91448c1b1bd0acc6708ad1c0705
z82ecd3aacc06246096b7298b1e9f9f42533dc67c32e1997a39f26267f916839951c31932da27a0
z94d39fb621994dc6d0f8d7e1c81a796bbed8045fd3b9c46e2e870fd909a2d957622f986948249c
zadea45a8f9ad26c3132bda8a0eaca39528c05f52695cf25e46b6e334bc6387ce43f495fc0fcb3f
z94bbf81fc16febcbaeb4b608c558910bd0860b4eb08f26af85c9a2c91466d733a75445de66a326
z8e72641bb2d7a6d1327e9b86d42eaade098993f2e725581b714db5e63c26a0e9d9c5758133df03
zfdcf0cd077f8bd912751154cb95e51decd165bec2ab8814b75563a232f6a7f02d21c8b24cecf2d
z2de9a19c53aeb231b330eab2fe26a29aa19193915de151f219eb6f242e2815f1310df06872bc92
ze8a02ef643c6ab52d5883e4b6afce0999ab2b0a948502ce82ce9c35e207843d201269db3a455c4
za665afb2468055b18b586c07b7736e4fba13385ed8281ff5c09a64e41314878e9c635aa779ad4d
z041ef7e1acbf46afef0b53a1f675eb55631a16e16f58b552d9731ffd2206a0273eeec918dd242d
z690f957b992bcac7cf8972bcf10f05b3d55a0e3eae2b60e0eae6be41d6a69347b2b1512e265667
z247d9430e154e33f9f507d8fae0c5da0fb8851e07cd603ae25d4ae21317d92301d140342cb42dc
z5c360dba89fb04fdf8623075e93050b75aad1e8bc4f67740dfc8684d4c567be18fb0e86db03e7c
z25b4885a54001fafe5667f82a9e3da264422ea6aee9d76332f5c5e8223ca7bc82aaf80ed8ea048
z1316bddead553ba0ef05cbaf2c22f6541287124729aba27f22af1dca5dcfa04a805d24815a0418
z73d37b2993add0e5cf01175a6736027ee4ba67d4fdcb32a64f8877eef02a880fb78f5d3549b7f0
z720bc59ab2e94619e34e178f220a806059ff1fb51754728d6b51e2273c54214f0d0ac701aa89ce
z892cb3f88de22dfdcb658dbce703a8fe129023f445af7351038c1f38dbf95de8a33c0828c735f4
z870dfbb1a6a07d7991d56316a28b6ace5358119269f2f2156dc7166aa4dccda18596c821499ff6
z82ab5d9f241fc9b0071d2cdc620470c8b76cd6ae44847ce90888f0b13e4b946570cd28b206a9e7
z7474b222bb98901c3381e8eb174d564b8ec7e8886961e9261e3c59a6d8d2b5f934e6a70385314d
z9796ced70d30d634738399bba712b6187dac3c94844ee38a80a792e1b1a8a533bbb7c553ccaccf
z6d74c0f0bee2f8b4beda3c911d181be90bda0d812071c3257e768b2b9ddd898b13660b637b08f8
z7f5af26aa9b50aeab9b8086f5d641a9347fad4cdc468cb724c121a8da6c13f018e730a1d59dd1a
z8caca6b07bf75a4f86167c2051aed9ce163e6b702c6bf53e98e404955ef145e165284180d38268
z48d3b58a029abf0f1c4650437f82e8319df6912a5a9fa51e1f741f4783b6f5dc61ed44b4e672d0
za7162af2dcae2e9ee6a4edfd57376053d378a247a110169b0fefe9c2594af29a90ce56c3c7270d
z213cc8563880004ebfcdbcfefcc86491df50c1b555b5cf6acc25541dc0b8f796465d8d2be507ea
z2389da5297cbffc450da2dbb086b1778167aa8702bdd16207119ef4c343f7d46cb3c33153e3e2f
z06abdb487b655cf64db764db045e7fe1fdef5820383ad43c918943571a39490f088158be02be4d
zf0a2883f69a6098d6711694783737d39e7f319f95ca638b6451d253d84da8672a13cfa54ffaca0
z5b115d13f0f2977a2e57c96bace5ecbf7106a1afcafe8647e3a60cffe85b19e5711d18e1a41003
z6081b54ac83da9e052d5a2872dc77b8641f4b8c9406de2bb8906aa26edffa45a9ffb332dac8411
z6f6d6daf4763005ff5b313baf1b2765449b990d09abb72676a1a7191ed4f75efa241beb2ca6839
z203c58d6172fcff597dba68370c30a7617cbf45fec247d1be01ac94683497a55b28be5640b9861
z43496e5258cf93566e650acef8c0ed3d3dda443ed0fd24d9ce0dd16b5b9b0b20d11120f0e4798f
z4f1810cb7da5f1126e48b8077c02fbdb769450b77f7922ced19d145a2e58cb5d8b5f509d813ea2
zac9c903ce62c63789eade25091f85b418b56cda30fe8ff6ed4953dc312ec042cb9e80f107b5d65
z91fdef9b6f32d510f06b58f7eee921c89d618b8f7cdf3b492c2d5234221903b394b66155628cdf
zfa6fcf3d7551f42b93f77cd8344645805c1baf44e4b8fd50da66430874c5b55b2236e47a303da0
z643c7f6aa1a1c4777e6cb2dc568190e44cde670b29b45be08b5c8a536d274219676fc0f3329f0a
z8bba93c6609ef8a946690152708d47b08e505551dd655345f4c9b22102dd1a4d46e6c9f8133af5
z93cf32961d5d59f7c7cfb7ba85c1240c53676c1cf4f7f319f1e8e4866ca84af9baabea61ad4340
z4916385779f3505697aae26492ca4d8113f4a08009df0a983cf515a8493bc55e854280372cdd48
z101bb7bb6ddb15a0ff62bf93e2922fcf65644a1aa7dd7711fdcab98b1671774aa25b3a2e758e84
zd61b042a151f5baa5a29329f14c7947d55f862fadaea37f1186281b62be5b4fb0cc45674686792
zcbd0bfd0833bc67049e38af85e60cba54a069297d9e886f2c5f4b6d77b9f557b76b72b3fe5fa59
z06b3cc978786131ef8a89fa31c9eb844639e966619301d5b8ae12e9accf1e72eaef90ca407ace7
z5262b105319911d5ff4abee43de212815f64aab9494034e5f33deec68f23a2e182aab4af531568
zeff542f2fdd641c05a03d91e275608478ab6b97dc9ed455b0a61fc2c09d35bc6bd041de9667c7f
z2807d517f246a805d544769d2b7001efee4d6b096c5fc14eba20cdc7d9b9da6566534608614a60
z15f34528a2885ed69661dff660d62744a17af91b2d1d6a6fa7e408906ebad0a1abc1963d1171f8
zd190ea7ad8de5d99af1a4cda9e1b452dcf5e3b2079fc4c1179bdd78e944d7df0eae67e08403ec6
z7b67bcf88e6845b21fbff6f9957e4a0268cbbb7afa7b8c284b627405753ee48daa65fb407f51c7
z3bf8ee84f95d402dbcb5e4056ef38bffbd9ad487a5cab31cbfa75854be3118b0e767b2e02bc10a
zfa7caaa5b97d24d699a6800b755f8e0d8f8d9ccf2ef437b8e9c3a7a3c4af898be0a8d858cc91ce
zd25a280eeafe6f273ef411f8cd12014af98d240d1380aac62513368aee1d83339bf0881570243d
za94cc1a7515dec24ce26c8c49028e078db8ecb53950018d0aded10e2de21b7ec075f71246a6a08
z34ee40e5d9674b4b021221bd6ecf6f51223e810890f9559d4a021b9c30aa5f67bf82edc29ef641
zd458c7ae0eec314890816301ef19623763e5e98e6c56c534005c830408c151cafb4a1f760f01a5
zf3df89212ed647d3723e8cb2d55ebb700893bedb720b0aefc2fc0c3f00f8a7c2e8ca4d25507517
z2bffd5e5dac8da30b454877453f4bcc6e1aae21dd3f31248698ee28385043ab27be7cb769a95b4
zbc248488829f817aa8ecb8368b96799e5d4573509c9112cfce316160656d0ae82daadb4378cda0
z6b8363e2b44549fcc9cb7d0d0752a66953b52468481455bfac759b67117aedc118ac97b9fc5184
z6c66bba05c3c7caddd3ba5c1c85405a9bcfc7219839fd62d8b1e6514f9cd1b6f58e8d5e7075838
z7fba46d1eefdc979521f4dd1cf692837306a13d275f111ba637819ca2b8cc836eb1f5e5dc74e4a
z1e0640efd3f626a51fe700e0732ac91af2a70972390c534304eb66567592a1180d7f0bf06621f5
ze63ac11f6b20819ce2d1c059a45c8896ba6e94d37ab68d80dd64331316bb90ce65250797fcd76d
z94300b1b2e0e9620cf9076999606f7aa722859c3b900a4fdaa96ec37a6b5967bceb91742815c71
z4c1b1940e9aec1eae81a60291513daf35e2897a12fabcf2f41fa5eec092992b4356d467b8af99a
z7f47c09743b202dab6a67bc3eee8480a08f40a0ee3a765c0e4f62277e3dcc7c0d4e29e2ef63bb7
z8da80ffe6e0a5c68d03fc9ce8ea07273b318d5b09e11789aaae2b57e78b425f982df94a31eb70e
z6aa7713779e00f6f7ab0d7f32c3112119c760158e4a7899ab3c43f6ae4843f0058b3a8765e583b
z8d9e9ee6f803186420bf541355de1bd286bd0e9a8983235a7bac5dc37bead3d1931bc32a5a4dc5
z3781a3224af994aaa375f7bbb8864157351fa04dc54aa1675bd4507af26408041f3cd023819314
zc4a8a04d24a71e690aa873e68d388b81ddf81e52009b834e361d4122974894b33b46c438761479
zeca8a4ff964bbf217abba332449ba8ba0047c82d13e2e4ff611264db0e3c3984d0266619cf7dbc
zfe08338720a6adc81b22173cd0d594dfea620e000d059e68713f1ece3882752c716014fc4296d0
z349eefbdea6e6c48941ec6e5a8ccf97ed8fa9202a8bf5368b8a4882df4ea8890b0b6b7184e3fd0
z27aa2112e4d794d1f3d9105107919ccebcfe7684b34c445637866df29a5e42c2664c5278998c52
zc9abbbead855ba837f79327db939f1e77e6a3cb69bdf0775abe463e6f5ad80e3ee21f919d92c00
z7a7272a7914e7a693db0b6a3e6760071d56e975efb37a667cfcda3c7fbcfe741280e76adf2f484
z7b1c57a907306e52dc6d522e8e3c849b2016ecf023bb03aa59fd0a6c1b5309971fafcfee7f3c43
zc4e4d9511823ff5393e8678feef1736f98004d99ea9093b049f1203fb49e80fa0c706bece7ebf3
za569b8b64226755c8f90d329e88e4d504054e315f52f0268a59b8a9f257211ee06daa6f4c9f971
z5a21b3e2792645112ef174be5720819aceb03acb9fe1da3ab5fd36a4d31fac5d1aae402ad4e8fe
za91d73fb3b1f49db3794dda875118a28c944f0dbcf523b799059f86dace404d1f488f00539ec5e
z41f70a81ff1e77a0dc40aba8a790d4808dc2b3c3cd4695c9e6165960dbc24b8e2328b8a8eae52b
za4834fa53530534ac8f34fbf357a1af8e8acaeb0e159ab874a8bf9eacd3ff06456b0154c929372
z9db033466f3e71d46cd539264f3c0b3545a2b4f0f7357828ec0457741f42b10552a2277e109af4
zb9b0df7e450d0ef1d1d09d275baaa59acacadc7bd9785ef0d7139ba7ccd2dbf93d621d2129a6c5
zf9492a63113b73d91d415685e353b8c49f29b52c0992b77fe3c8d03c24674ecaf36143c6ba9f0d
zffb25f84f64fd9cb7034d4fc6131028978fc70e236d7784ef1bc51623f17418f73bb6809bfa937
z43a6187b98dd2335147667eb3a11a2f18c297679744e2f97e06c459c35a1bcccd02931449b1ce9
zeeaf7a3471f0b9b058f1797f0c986f0954db49bc43b35426c979a5b0bcb315c290b10ab1b4496c
z4c19e4655a8662f3b8355a8cecc785252c22fd44eb20bcba8ae9de62d3f9beb97a023cb0df9e48
z6dd718da27a5022d049a6f7cc3eb4738b1a84f2c84a0e7f28dfe5cba899852a91065d78e8aa8f8
z6e732512188bf6d1a5ce1b12e70331f7fca6cc53ecbc58f618e311247cb119fd5fd5fb6d991c04
ze12af697b3322dffba7a063ecb0535b998392190e1cbfdd30c736ae629515b5a3bcc5f2a5b593a
z2ff427017a394f298934aff9dc5c4cf29b67b2f49befd6e4fe94d89eb5c2078bf1a531004e8894
z1a0eabc8c7cedcb01a2fbb643aee26c799f5fec876129dd18f953f8a6b6eeaf5198d78a94a5e5d
z6e909329e7ac694ba87da4d86528755ee9a7ee3c28e7b335d5948ce131009ede5bf6db34686dd1
z4755befa4d94bcee08d71165831095c3561df71273e7a433a3c5f8aa044d0967280270c65e8044
zad90db9edf17d1e7d4a0df31c673b58b4fd5873d0deb8d8e4a7853fabe8b7637192210064158be
z081dcf62e92dbf2f2fe5cccbe4acadaca5c4f27f2860a4d417842c19a887eb80ff5b9c88ad2b71
z6538697a04becb9fe08535e04d1e1e6b8e628b7dd62c0a50ad2bd3d81439d9ebe55038d41ad975
zf546319f8ed3b8d3bec82a5ece467494df2b2ff5cfdd3a19fb802c235ff47cec0c6524c047044c
zd6894cc4b5a0d5cd4b35aa59993b02c9f43fa733e5da990bfab7f9c35c8ae9f1c186cd9ba917b7
zaf8e2d1fb0e65b19e03e952926d5128b9858bb634e86e432a77dfff218e28c2ae4ad931f20a025
z06035f48a4ea4ce0aa521854d7736660bd0530ffacaf683397e63c1c9ea81193fcd4863ad89b37
z8c601352461cd5154fcd3a7d4f5788ec19d6779e8cc90b3308f0ec033e2f51715ee8b70da2b0c1
zbdf1a9fb2e0d659470a69ee11f377f0777d854144e8030000b3c3eb306f2451e9b842c9f465688
zb1903c73259b71ae97fbc299f7c3e7ece790e0ba0700f9885136c8a4a6e5edcc6eeb75d9ad4fb4
z1f29a7cc8802b686aaf1567c1a4985b4ac6a48ee4ab491ab54270fa67f7981848c98d9565aeac6
z75389c3420fa594bad0a3b7ae8030a87f13e3fe54c22c1eb2f9ff954c4bdd775e69f8ab9b5d94d
z7bb873f04132e80b57f2d1e3f85f7462323a8ad7161f79224c61a034dbdc6c1f97a3f7d03ccd9e
z80c7a2eeedd6f3dfaca6969bc5bd98023ad444a6bf9e7da404d94a43e0e45bacdaac83c1a29d92
z9d4e4b3d635b8b897b615286752ffc61c96216faf38562f66bb35b17cae90a73c2a0e2067b2e5d
zc18ee92856c254ff2e680f61b0ad90b763ac81af843597da4e14998c5704f96965739bc168636a
z797a84ee1070d17e2ed0c43f97cfacf42b90ccc06759f143f8daa8109bae00c508e7085296d609
z56351730d2b7c085a32b3ffcbd48b1461f264a39e594012b695744fbb21a2200cfb91e9f2dec70
z3a34d27cb542af2af9b7933763e60d794df0cf1655135c9565883c5ad9b6cb55cf350d9a415e6e
z0122708b9bce85bc10b6d63ff7114f94643dbfaa7e5665e395d87d3d9775adadbaefea3cdc5690
zc04674477eef4246354bd5f14ae8e4d1fa09ec2ed90e8bf85e6680846e7a8b52dffea4d4f1f87b
zdf403705eb0d390af91b1b6ae50d78d8a9f53688dc13acf7b573c0bd826d26ed744bbddc701d0f
z067aa0728fe433a0332e225401b5a8cd7b1f32e46406549c3e1809fbb45d3c229e195c28c6fb63
z2369d92047e88456c2a0e468618b224210ec9990cccb9959c20b82f122cb8994f578f5719591ca
zed16a14f85800fad933147fb372bcd2137d2936b75db183b104745fdd12e298ff61ab7980cd8e8
z0108c889cf23f89290d140190ff1a7b206de198be8685d1e46d31bd43ad158560d2df915705a43
zd98a34bcc8ddd09993b7a9813e1cef8e3f4628bbba08010d050a18cd11c9bfa896b4df0d924e46
z523d02cbaaf72aac8604c13af0c8a5d0391a9482b7191a1a56a6071beadbdfe335336c4c60c4ba
z7abd8d428cc0ce6783ba0075a525d6cc6ba870f668641034f95f5902fd68686da6e095dd59dfc6
z487a5792a71bc974be4b69b194764b556551186e42ec0c4c579ebd0808c2537b084784e0209bb9
z3bb186dde34445412e828ff9921a93ce08c3a4d613a7497954cd57f0ea7c485ceb299863ab9f1e
z2d39bed552ffd49659c67ec76dfff777314ead39599a3041a0263536a7d1ff52bf8d7451d76703
zd8dd4324e43a6601e30f8bc4874289fc579503cbc3ecca2f362609453bc5dba0ed52e6b0cbf6a2
z044a67912ffb23129e631d3b851e8f8ae70486f74c9f13598656f62080668c8538a5ad84257826
zaed47c44dfbffd733fb1acb5c58d5ce58ebf3459e53d0dc428f498102b2f426da1804f97b37679
z99b2aed6ec40b54c6421c0ab0210914df799c443eb8acd36772b8c3bf95ef9b2b59138b8e75fdd
z338a9e3eb18d11c6fae2d0cda3fcd47caac3fa22e0ea4ced702291d43680248867e02fdb6c6f75
z6edbfaf574071a4c4b9f47d4c53b18d1dedf378c58bea1fedef72e673508deb30a6485850c72a1
z1b8bc0db277c7d65bf5119906ee9586e9c3c5ecf49681b6bc3be2d021bc32e4046d17f9d879c1d
z1b5c2f8c5fbf5627e97d46ec69d8e43617b177630b58450ed030faf42af545007ec81690343a56
z2bd7e90dc34c36dd837a47bdf1b42cf8864be9e1b037c6277dda9b6e08665d392db2e35ced16a1
z6983e1237256514eec516a06cd0a63660419693c2c0679eb6b371a05ca99b580285f1bfdb4147d
z871e804ec0140db4b8811ba1e8f7f6cf855371d07a8f886a02f80d2fe52396640b84756ab1f1ee
zd1b17d7837b21ff361746693a1b4ad421e0348f3ee8805b34197558a1ea373873dd03f7bd8c8a0
z2edbc882a44841a6fe2a5c04a6488d10b6fc37a4908c7844ce39b007179a97e881b777ebcc00dc
z425563a89bd5a81233ac7a368796a50a7f5c01ef4ffcfd2a40259545f88b19f15c0ed8e8b5da00
z1e0014b4c228e8e85ccbac36ec343bb7ef58984a0337a82c6b257f8b0cfb6fe223c7d761612fb8
z7ee8c74b78841067a4d718737c9770f59eb6254bb009ba8ca02a0512455b90ee1d9101b1b3ad8e
z9baa536e4d353ff17fea6084f9bc21c70cdd4f9fdd09d182b16c0d19f37734eeddc0591d8e1798
z03b0d615280261814928f0ec441e45266df9424fc3c27c01e082a186131c07c21d63ec43e13838
z8775fb626d7d97cff2d35db305c5880838a38332e34d8488b725b1382d157de43a444731d4861d
z4d5c580b4d50b16bf7d53e38c6c7891fc4ccadf1306c70e97976ac78dde299c25cc3e942e42076
zb33a0c21f05ff23ce7cdbcfd2d6d15ee9eed6927e02de4aa65edc5c992993c2d25b295ac32b720
z3f670899464337f29b6eae0854786bd3fe088a49a5e23a54a200218454b609c8464e085f282304
z40b6086b8c313d1842db1057d0a0a35fd064eb729f7816ca551793892b46712c4421997fba6a17
z1ef5a4fb5c61bf1d7230aab9cf5ca05de3a69a54bdad85ddf28baaceb37983bace4bec2fee1e32
zec937bc5444d1a9200d8b18123d9ec484e4c37e76d22a0b2a69717f929ad63b6b004df8c2a0ea7
za0f0cf2ed304790895bb9fa30122ab98fec7a7a1d4284a873009f21fda9d20e697a23dfe71af77
zbcb69a3eb25a77a5c7349806abaf6b97be246b5c73fcc727440ec7df6da38a267823d0b41bee5a
z0d37185b61bed826664ea3bff01eab40610b0a2b5a872802678741af7b8d1dfa7f1b6a10c07969
z0fc9011394477dcf698373d0c717d6827d703a4de24adc5e8859707845409433ce1ee35651c919
z0bf6f599e4d85c5e49165c6265badc4ce459fd8a0c7a2baf898b1aa1a2eb91d22f4dd1140dba1e
z0647effa264f832b8ea4777113846d77cfdf2441385e9534c824b7c924f235237dbfdcaf6cbd79
z2d0aa3d733e83e343b0b8ac67084b952064e6e8e226460f533118116de452113a9c9f66248c8ba
z76d241017a1d5f85860e53b7e48c3043d2c120a23e7b1a477364061f02fb051ecb27e9bec9ba2c
z2f88e5b7779ee35ec27c76d837cf32d8c71e99eba2b4ddc2fb08f53f6d0e07ef53c1eb5c53cbc6
z7bac06f9f9a23544a49be23ce0df14c450012d02b4801d6a248a23aa8a9c1e3ed0a746dbd67525
z732cfa1536d2f4e5812b774529e2b766b7cc05bbee967c381c1fb8cfbc22d724bdc0affa015696
ze66f3e16e708eb28a898a52dd57d559a7d2012c2fd450e5aed1d25751b966b514907ef184d154a
z53fa4b7d9c53a4925f35fd4d79c08a54a16b4e8210afaa73fca6dfd81dd334fa23c656f123c913
z3a892fd824ad52b5dcdb1c54a7c76aa86faad1a1f34e2b7afda885ba9585bb53a2fe7d0d588816
zcea68927f04818a1f947bd882f9c0a6f9a586ba8206c2ce2cf24fd6c8c9fd861bd883d994a226b
z78a4454a171a0b3296e4663b4c618f316217c242f664c47e5f9ae4c7486d0620a2e3236425b6b9
z19fc00b51289c83c3edb7465af62fe0e298cc00d51f1eb582cd61ba7dd8724e8adc0d8752bafdc
z6a35331bc7edd20576092799094103633403e73f26a6169286ca504799c2ee34aa18f2c96cd036
z6f519225b109e6e4db5c53b17a26b70b1d84f56f65ff4a927df3c6eb05d5657d05a26d827c51dd
zafb3050841e2538639a8b6538bfd43ccb9dfd495ddf0f64dcddd53ef16a02866303bcf628e8bf6
z6efaebb5d59daadbf914cba8b31a14b0ad52de2bf3200937085a13f3d5882344fd36396d70aa64
z2fdae26e0a813a7e022d826bd9f1a8f78d46b252f5d1129a118a168a4028b216e648a59fa46a7b
za1ee59408c1e9c25a8f66c1ae132fad68681c4f6cc19bd3c884185c9e9741affa7be2fd16a6ebf
z050fdf8f8f4dcf4dc5f0ca28b82c8107e4ceba705ea00917553eeb3e3c55997de66f4a66fd9ee9
z61409da7f1e8195b5575d7da2d8f3126ed518dabf960804df955b25f3f011a6cb33e9fd3713bcb
z8cba07d488a7ff07d942410f4acca59b1c92d47c674f6ba2b81e96465911448e64b8100bbde9a7
z8bc3e12698cf8b27eb40ed790ca898a2cd11facc957842c9bc02ea25dd38524931fe90148cc3a4
z61041d93c7ef79d50761f54613fb1262af140c56b55bdd68ed9357ec713a9a391a7a81a528d91d
z5a98627ffb263c87520fae0e4f49b68e2fab0baf9a2cfad58b599a8262748851020a4cd60ad642
zaefb9405ec5740870d113a207fdb58b4d8b26c4c3e0657fcf873dee28f32d43f18042559d0c2de
z83862e7faca385294567e5c57dd0d3ead11a1e19ac68099f9fac3ed1e96d6183ba04c9958efd74
zc1745d2142db0899718e7f08f4f9f58e17a95624965a5f8f798829e358aecf192bd3c8b8e858a8
z69947074c261770795e9f8f0ebd4454108b66bc6beda394ed045094788251e9a9db3054c7fce47
z372a3d37eeea25a92aaaf4d0d0142c6d7e46715afdfb2029e2277ea98175d9af79d8d208fc9854
z3ddfae1794faf587ec6c61a7c92e9f8399f57912388b30087cb5d32b5ae1361515e3a7a2ca3618
ze33b9c66e2149c450a93e27d2a52c13be445aacc4276c16eb5105ff56feaa586dfcbc236ffe4a4
z4bfaced76b8fae22e9e39298d1766d8ec7af1a13d251ebf0968bc68141d42c35017967d399e884
z4f3c11966b072beb1dcf1b5b7fe693602a433529daa79a49d6c915ed72b646d949941ef5ca7d1a
zb3284a90bfe19eb0d38716629b7800a3cefe4cbd20927d78c4fdad91b36afb086ef54d0844d14a
z6da60b2058677ca5a6ddd71b3bbb056e1c1d471f2b0a4ad3681c322af74a30984cd0e0829560c5
z6546afae8a2226cb50b9d157031b411fbcb7650d01cdabcaa13769f0667aa94ebe63493928d5b8
zdcae73ad0d09ae570c7ddda87a9d6600ed55706b9eb811944b833e24b4140efa0f11be9b2feecd
z2bb6ffdc001b25b1f20a079eb7faa1c90f34033d44abff21b62f022b6ad64124cc66ecc4fed7fd
z84cf7cf977839e374f47da1cf4ee33f81aeaf31b4b94503b015ff01f40423ffe75684cdd391007
z69352f53a467247f0ef91b3d9b3888ef27a2f3f990d4dbd04283cba58611652a98a99748effbf5
z526e2614d76d9f8367c3d6bea1a650aabd0079acb602e302d06facefc71b8490afadc48a4c8533
z1e3c924fb7296c4bcd95219acf50f817365a07975aa1c38e673aac33498ac345f49f0aa017354c
zf7486e3943a3e61e55d9cb870a848bcf05c1879ed0339ff45f8853c2c881ffc714faa4449cc9d1
zbb255b1e18e100a76eeee9f4b5ba924ab42b5f5e4b0989e0abdcfbae7fe10395c98e0bf4fc696f
z2d946b22cba05678b359f423259edc62a0053436c04499ea522b2b8746f8768a7a4313c488ab2e
z5bbd2c13fa6f84b4c215905e1f52ca59d2e654362a47066fbec93554cbcdd5074057809cf4ec4f
z27e81a26e680b3d3d6f5de0782f38e96da829325ef39c3057c9bf807da6ea55f5e54033db9f004
z6bff25ee9cf35c2d84c36b2c5785a74934de89648959ac2c6bd17f363848cd9534cc3f57d23bc6
z3235035d4554d753bdae8c9f9aa18f3180e4be41f73738a9648491041592b6ea0cb4bd7878c4de
zb32e3591189d30f03253585a75959988e4fbcca7aa99eb79a611f8768e9a4ac45dc0eaaceb56fa
z7b91a3f117b2356e3bca95ab6f8116417b7dfb38ed0a38748a92538da15a010aac86d7687c6da2
z204e9a3945baae43b0ac4dcf7f39780356c5eb11badb995339f91ac68a915a5cac8053aa81a03a
z356ed5ca31aa09317f52afbdb3b380c528fcd2ece7d45c46058d559684c3bba6666894863472ac
za4f9497e28e915736f0155645f487dad193bd257df1ece80ac8abdefb43b7d1fbba47e061cd5e4
z3e6fa68bebee38550acbbbdc40f0c1b79f6ec4c3520b45059aaa4be658147dcc65ff8031fa3b2c
z927e9cc56a26e65a5b652e383f9ecb132b3c02e4b3264d6d48d2e32c36082096401e4bc903b18b
z9412ad5e90483e346cff838afe917666f5fd8b571212a8231f3422251bc4c1530971fc364ebc58
z82a9cda67048d517d2e774d4abaa9e006ec7a7023a3fac4e8eed553b1399082bedfe643ec886b8
zd538a973fb8aedd4da66c19edb805b1162f92e0c7fd51b691140e02bec64e3da44623d0d1a61cf
zf8381e7362731167370d889816563095d6382c46855f4475da9e4c70aee726fa72ec1dc61b8ce9
z7b65fcebea7b02b4ddd852e2837ad09628703fe9f062b5b437e2e3aad5e59239670dc285fc9cc3
z9bf0ec0da7c8ffffd06eb017cd11308d45c405b29cfc20ea513c57ce6cf394b4f20f391935937a
z115913dd0da20b2e443062372a57f6bc88cfdbacaf1c0e0b77049c1b0b3cae8d7d2c012918ea5f
za5347061c09f81da59e318b6a984a6cd20621ee36c2d4505da4b846a2e79db83b94bfca988d560
ze3e024cc0f4431c9960b037cb884bbdf5497d927e9c31629a7795de38903e92a5353215f40ce4f
zec27d974179e0d2070d700b120b936f6ab4502373973f99f25c0e20e122249b9e4c6ccf4ea717b
z256785a633a00b6109f5565380c23a9128de613bd49dda1be7947dac0ded4eabb181fe7237ef70
zca6e777db6fee73f9f2b902a4376926c04b337d4aa79f774a9c0978beae106d52e784e5ef67ead
zb3f1598784a699ab64ae80ad4ee793332cd30a3ec0e144fe6b88a0033d63422133c488861a4b7a
ze1ed32b45d879830ca5da3fd7e8a9723a63f556721378284b16a59a72a33523290534e73df0781
z23d0ae4e9dc70d30218a96244635a0b41eb6f28133f5ecf2797a727726208cedf35cf05bd1ffa3
z499851e4ef34a3b810064a9b63e358ebd87efb01ab4f172e063ce5936e3e5389285e4c22a0827b
z7e57a6c5fb60450dbddbdff56c4e25bf65f20cf2217d75a7d0e3e566942c16a5538ffde9486248
z5c3419103065e0d3859af985802099802c51a31989404ca22d267c510d2dda01ac09cf6aefdbc7
z6335bfe964247fc3f6fafbe509ac698edc086947a2c5c5643493190889511a183e7a2b59e2e91d
za332d700d69cba235e0fe9ba95867538571af6c06b0f52f0230fa46498e57af084b8db1104a1ae
zd2d9087da8a2daa7815a12f0ed7994aab230e71844959eea10bf5808551235b31d051c7d4579f9
zffcaab1c09321b250a490afaae74047359eb0dcf223767dc056980d48272f68d8c42e5f87cc9d9
z6329ac6e1b491bcd537a77d9c96cc18a2caf35d12867ae1bd7799c641d61fc9f9820c609e9a3f1
z7e6d8c57ea090b739e53cd83c876eda040710371f4f503da996778df5383cb38d03cc1a8263df6
ze436bec83e6b131bf53cf315e6dddf41046744ea2dd9081aeb267444971a63c7e7bcefb0775f7f
ze815b21d372e05db28b65bbd7ffb05228a25d0d683020c42042220aa46a50849a810ce8ac0a6cd
z909fb4382beda8d005c6d540ded90afe9fe1e0f3ebe8ff53a22e81b1b35d9b79338c8e5edc7186
za745d0e2c57ece52a52422fd223ab0dcffa4482662f4301a9c393e64821ef1b3fbaa250ed2b130
z7e5b0e583db6afc24789c6cba185793b75468fcdd743c41db47650ebc3f8f9fee3c079d7970359
z5aed5c245587335ec35dcafb35e21550f890b88ea3cfe753ebaf49ef1c5aba3a4bf64de3b27fd9
z02c535b825aae74e3580627358aec4bd642548ad97df395b881de7554b18c719a38cde7806ecce
ze135d09242d1f945aaae6f5eec7e58c0baee304d70f3549ef3a108be7506a22d5173a84adbd79d
z7338b736e11e8f210874aab4dadb87703edf1348409eb8be47a635a1cebcea3a4d06938e0abed6
zc7458727b6f93aee0302abc83e64dd7ea601cf105348d127eee3e4b88d0b3e2aabf21d8812f33d
z37cd004df05bcac6c0e3d68b637301fffd313406d066cbc4f0119e3d0ee3de77a46741caed337e
zf2a41e85866a77f5488818565c44101689db7d64ee6e15e03887b1dcbd99ce5814fff7e59a3417
zdadbaf9ff48f351208f93d4077d5b3f518c92b8b4ed67faa5ba88e8367ccc3bf6fbf7b120cb845
z9c5777200e50ee3c82324a34704f68bc4c7b6b85a74fa211888d0a27be5173dbe474df7aa10d25
z0c0dfb5f4857aa997e56909d3a4716512e1a1c28c3d52649ba176eed15de4ad3c9944b70ad4e09
z7c34560a5c440a1dd5ed060bb496c58f37f14a11b1cffd32a167dec1d725fb001cd0ce904ad831
z74038e97621ee158642eb2d2add430b680c20b5696d96c1e4291264ccf102b599aa09c3848263d
z1c79df391ca7cf8592fa783989ec975ca7e280133fb858897688973fb0e7d2eb40a6ea90ff6f1f
z237f5424d333ebea45d038510b58698e1407c3c3945fdbee850568ae7659731fbe010ee98c4d2d
zafe5c8111d218e0bf183ba1a9d86da95de7c49fb5f05d030cd8ebcca38b5ad8fab82b8772caae4
z8ebc5e2c77755568bfa5c7c5a18ccba316f1b21f7d19ae1e2769a3e7309ab1fdbd1e2e994f3372
z2bd8ce257a8db93967775322dbbf10222b651722e14b826235e16b7f34c4c84dfe8a4a0af76c4e
z7d5e2156af59cb8b2e7378898a236d2548e4bf18054aa7b4604d61143e508d531ffa97150f6432
z7cf9118b8c0d877e7d2a321fc6fd79e3dc09ff2b0b1638e8a79d6b648c721c720aabbd549957f7
z392a26b1bb2d898c6ace76bfa91a806451e209ce89cc08744b82c78be54df3b3f7a86d2ed99a6d
z8b1db1653ecf853156455de7298c8c35fba243558b105a429a1d014a1c4c2dfd5dbb56d373fbde
z8f6931b331b08b1fdf59919133d290736dce71f68c4a1e2a1b6be5d8463d59137c65c185776523
zc57d54ce1b5de1c989e626d271e79b267149a35db54a3670ed01c4d4d4c41214eb9fe1b60a57c3
z77096f90b9959bc35e5bd8cafa6f9b1feb8b2f6840788989f7807e4aeff0390ff34220465b8529
z6ff7ab5c1f360fdaf8438d2228ed3c5a716c0ac3cb31193cda82760fcd023cb07c44c231ab1e51
z6e2ee75e795a95ea2763e516c43011729d861513d5ca6dfe7c4d1e249c3153bf28b7af25386496
z5c01d3304473da2ef34661a213a0c5542092ba9011388187a23f0b264518d1b0fd0e95726ea6c3
zc20e30678186f63d9d3f5e32613334ec2fb4f10699d0efda3445ea5abd0c2cadfe5b19e26e4592
zb65c1699f9dcfe50b1234dc1a0971b5d8cc178819a45cb5cbed4e1eac3133f73f377f0f1487f97
zaa6abad91b922c8000dd2d1cd3f3415d8bb3d27d9f22f756323c8505dd827519f9d0384baa5e17
zac6440869340cde9a005cd3c278686f41814f6c21ffa0cc8b2ac83639bc6cd3d8168893631fd0d
zf7ba6779d996fee6e7c3f8c123cc8ce36ca3d5a35e030fbdf8dc887b12f511a2f672c6c4907d7c
z79e2bee39cd1006bc775bdecd449686c2dd196955314e2b003d19bd143aabdf30ba811841ddd08
z0add0e1617a97a2537187351bea50a885d2b9d08b64470da8ffbe72f664f4164666cadfb22c95f
z3e088b0fc277bc504aaafb0d0fe842a2b0aa137ca7b3651887faa858161184ff21a306aaddf368
z572eaba59b2496f2445e283eb26da187d4d006701501b854600d0edc4f792fb4b5ea55495ba070
z226151066420a310bc5b4821906d010a45bb9494c2536a283b00c8c363e7e3d6d3a82f6abcc4dd
z4f62852a7638d43433e185cb57f1b8c3c9300205069f38d8a930266d43fa72efd3a971df11df36
z1307d6eac4fcc0323e9dd5ab1502545b2d6bf9636a4e152821bfea762017f4e4ea50c13027187b
ze3356dea126f43f0001bf1c6dc70cb6e6ca423c47fad70d975189b46e03b34eae06ef0c234c02e
z14e3d56f9a1b930808560699ae7bcf094c257b62e838c535c171b75c7e6871502f413de8660995
zf15bbfcb76dc8026b95ba19adfaa2314351fa387eea4a3721582a8ceff95dd4f897a39937767cd
z90effcb413a39f37ae20608820e32541402bdc55cfa2cbdebde87134919c420de4f1093a96b766
zcc495d3c16e739f82dd247e764b556dcbb71d429b548705c0b906c217ecff84875b001becede39
z4122555d6dc3051a93fb621992df8dd5a6336d813a8c23c64e0b2f8a1c08cfb074bd0bf0dc7b59
za308bc2911bf272c964efaa05d45d80e4a5f373e6b24eea1af07098516fcba91b0cd3aa86cfda8
z2117bb53f0188dbeaa9191bec1037a1d732dd82ed6d5f7dbe9a118d96421062de1331d2e568e7f
za5651c53c6edee9caf6080c0a26f4b82fbd1367c7b59e9f44261305318b094cb2bde0873436c43
zdc7d3bb8b450114b242a5f7246f9049539b8b5bec0f8a8f9aec278d916d3458073f80524797be6
z5dd002208ca7333bdf124e956abe65eb934bf0afb3d3f133e3e47ddb472ecfc6f1ac0170238d54
ze977c606f08a8228d66f12dab527ea14418096b9fbbb3d87d4d79db6ac127110f2ae1906278393
z0aa53639dfba9a2fb2799dcf71e5638f489968b499e690e6d167326eda8521a44dec27d9e6ab86
zfd04ee00dba7034c628396346d7000945f1072c54c6a3f48fa509c3487a2d518ebdeb692355b49
zdc2c98e678ffd9e79c5266357c600fa35474ccd61bd30ed625898704a302c1e19fc9c5c4322305
z1b399487ef0bf379854c4ebd0e9278ea56df065271ca1f10bc9f4d82237d2a3dc0fc72e1202173
z386ce0554de5bf7d13db1e86745ea709daea40aa329f1cc255547313c6aca3fca90741a21711eb
ze23dee07de465d6b4acbcd49d115eeb4b1d0158467b1993e7efc04eb3a12e42e246509f0ac6159
z13f32acb89935eb98b3f57dbca54f04bcdfef0007065a438635dd2a024630319a6f87606daed7f
z2ca61d153db1ab993add0f1ed877768789132eaf1d939c8aaba4da3cd785ed0acab0b382de31a1
z8f50c4c5ffd421a1657cb38c7bee6a420c4187637f2139c227f9e18846f90ae0eaacc1e229a2dd
z961cb4824c2bb0dda407af4fa4dac41cf86910d14dacd6484b51fc41fd79e38fa413d949fa8d2b
z41185d8a684b471f41749afd448b499d88980880ca514ef5b7db0e8161dbb312212637cf93fb48
z485b4fe7dce6f5ad1b2ceb225e75946b7d0c4d416ea743762ad409a8939e0a5137254f1b4e48ac
z31a5e89d46247fd1d5300b0753b71bceb29e75870c3579de2628acea57b4814cfbd62b1d2fea8b
zec0d9046e06e0bb1bd9fc86b4d4911845fc1e3ac2aa88c086c2f3a45c8702a9eb1999b8436fb89
z5ca43a8957187642720fe71f938f71ac089b56e546ddec4bbe996730c5b7d53921bcaa4598241c
z0886465e41ee14b8b72010405bf21ec7af1b7e6e4d9d06b3c8a447e592f1ba9943a96d98f07378
ze516258ec6c53653724493bb4a48610ee1e27796051830f13369ee20a8b070a5d623c01df24267
zf01d8224469065633c1562375e5d4c014f09fd4ec6f566be0e57c7cfa2bc828ba3c1545ed5542a
z45c86f94b26a0c9764cac43c7585ead945d982f2d2c84216f1f94bd625541b4ec51418facb784b
z128c77bceebfdde8e72467980e549c7980b3c12fc3e678c4921653536d23d46369d843924a3ba7
z1ccb5efcba544f53822c79513cb395de55cfb139831be5d274c7ac48d89a776c837e4d9dd8656b
z0c50173125b1f49f929539f0fbe95e27e3c9c79c123a5f05331a358d1662412caf995d0666b8de
zd82c013bb595d537b42ae23edf33f6b0b9bd2885d0a5109d994fd73e7bd673864080c8f28e3f9d
z178d74d13367bd08ad899ebbbcb01ae6de3ce85bf350a096c54a2aef5f7ea94f6b44036d82d295
z45e94a9c4ce09759a6366991b3dcbc5a53cebc8387189c4dc6902960f5bc31a6e83b3b0ae45021
z3515d3ed9a3d95ffcd1fc78399e45ca5b2c8450ab71fa8638c0667840a3f9a4470dfc4784e50ae
z806b7c518ff43432344cb96a0495496f3cac36d6e91dda88231ccd1fd059cf1505373ae1938e1e
z944ea01a05a3573d3da2756c35edecc72a79ffdfd0d65a7114d2fd5e9cb5579372617b0ad15c5e
za89234747b718064f9c2dd379561447446a880731d05cc2eb36264dc5c8a40c8d501dca9e6424a
z71779de9a02b8474f064fc02218db29ff34c21e362197ddf52f24785e93d8c0f95389e38411753
zb3f38df787563fc02b02d849d357652e07976479b4289fe7d4cc9c96ecf2db7f944e1d1e998637
z680c03a4d0cfde05065265035cb5df02c45972b44ec7a9cf96972704e7c2d0a4af1cea0911e4b4
zee7d78f28cb8d78401d10f0551ed638445c47c5fb4d41436b7407cd1683f39c05c09e50c175e53
z7eea92412ffef1706823235d407e321596355f3e6616b165ee3bd58fd2f752148095fdae86c25a
z80beeafb7986f2cc9194a9b1bf7048b3d17086066ecb83e0b9493755ae480d4a0759efaf70653f
z2833008748555952f8d604855d05b6425e732c189bdbfc5b3bfa919497fe76235b80ce6e34b3e7
zeb844e4d7fa18e4b9c4f83c2b1441404527d3e98b551a6c11b333298d0fb8dd9c0200be549f6ed
zd9b9c4b42ca4d1e293b8350270266aa03ffe5f067fcf7ec2cf387cdab746fac54a34ad04a35311
z66f15fc9477ba8d3f099b815a886a15f8c931e9368a61ee6c3b0b2bdc19e0b696829ecd1d13b8d
z4c1a0271ef98a03e40c3f418cbaff3062975ca00a0c048d67e407db2b470023ad5171a26fc2f08
z040549b94ae48c48632f8b7fa44d04902a23418e8385a19b0e80ff011c17d283077ffea2f69fe3
z3b1a52ce4df60f78a52fad863ac70ba8003fb7e78f698bd2c0502a6826d590a733eace1f956f0c
z6500b9f45624624175c30c8db88fd66fa858e709ec568c7b61ffc9869324bb0a1e50d5529bded2
z1aa43e0ffb23b523c6e8bf4f4ee4fa2060efa6707d4d1161e0a9babaa3be2812c36cc1c16fde18
z67a56e0f54513dac78aff44c0fe68dbd14d41f18da8ff0cf3e611aef85b8f7e60676fcc38a1dfa
z7b93204993caa90479df92bc85ae05a47e68860968a57116f3cd300198ea0454a52085621f5041
z501ca433dfdde209201839b63d0bf5e9853af55e70f535efa5e0c29a3a062c4b93a86c1ccc7b5a
zd70f3ec38720f879dafcb93bec9f65de58508d0aba584bba9cee722bbadb4575c786c7d54afe40
zd85840e26aa55b416c34e098217173af6122e837421b5e1809552884351e7de6894f812591cbd1
ze7f4bc30c3f8f21028ad9d1b6f654f3bedabf3d0841bbf8421063a4f700ac66b3f6cccb5c0a343
zd05d9f6b4882369cc4b676795ba040c50fb2fb956ac46e0b027e3b5947b38938c6d37d39a6e3cc
z0e2c49d321e7d84d336f5ae9939358caeb9441ef85fde31a25d5086741fbf52281d0055fe037a1
zaf010cead1ab51515e840bc6b17ad3b2a4a801f15342302316eac84749ec86253d24a133f20613
z299c98680b33f83e2110295ea61597f366291846677442bc19b08d3f9ee37b29be63e8aab71722
zce5fe853cb5e37648f7640fc0989c9949a2282c997aec428a0bc344402d4ecc15820b5e80fe970
z96ae62fdedf1f7b77c2a449721ac7acfa629032c145c7f550aab02d0a0559a32f65d2377f85171
zc00e3dea7b443bf57e77dad0aae30d36658543f33b6f63b7d78b764a5be807196fb0e9a1fb73ba
z82ea850c3a405901d04172ab439cc85173c99bff2871b759fae6cf59e88d1d2d4885bb7df4cd08
z6572555f20a506576b4b1546beed5e71aa9aa689afcac13e4b12e468fd1147edb756c8db8232c4
zf6b6960cb394d24d0361f3e531ae9de1309ddfdb30ff5e51ddaaa86206d69e8ff74210a1eb96e1
z951eb2ea1889d6ef76144e33f977aede5ed806020277e305ef8f0729d7e618a06ff0a7688693a3
zdb80c8e9d759503fb419f9b281938ec25ed95bd9b2ba05ac9f43fcf7c052c43cba7b68be086271
z6ded89d48c55685ddd1d31fb2bc10f7382a23e9a96f254b95270f7f0ac060601ae59524a5c001d
z5a4ff2f3a2669779edaa64b4b15bc5fff7fdf0419e2b8dca0a4da60114e29b99d57a79cba27844
z33f407dbfe3e5c141b949fbeaa1c1e58cccf934b1d1f749edbae27b73c30fa98f78ba66fb6a91d
ze5b40f523fe73b6f7af91ddf95be5072baa9e23987978afab0b7d0d6358ab03f20d60274f5afb0
zb8eee06fb71f671be4466ca5c930692261e5b1aba168b718ba08100200e63f5af75bd9be67e8a1
z50db6491e5e0466629d2e1095cc9ca2ccf1baf932a32e6bacf97b7f4bea223baebcad6b3b2dcfe
za5723b8a7e182d3d14d5f752e7b566b506c9082b63bacbdf346ecdd3c7af54e69da3d37633a558
zf8477ce03f74137ad6d66585132dcad7992b4274d17881e902a9c07bebf77e77bfb56ea9589f93
z5627ad34e1da3a5de26bcea99f4de1032284199994a0336e5c625c5444dd39692ffb9343a008a1
z91b34c86d60f19417198b23f26514b0e2ebf162372171bc422787979205ab72008b68ac0b04640
z8f9ae07dd8bc3e0f7e3a4d4500025c058f36bdd540a25b6e089c001ee0a0d77a4f7f72981b2534
z1f6fd90a6abf1e2f31a9f50a9bd66ffa5ec18bcf9a50b6ba495b0a1aca1fe82e9c59a3e2ad7d46
z50370ee73c0b33bfff7eb01e56bad5b4d57cdaeafa1cf563db1b0bb887e06796d0fddb3af91a9a
zf063108c7e31c9eb821c58b90fdc5c2526d52463b1134b04ed9a9b0b92657005c5cc0f228c25d5
z06ae4cdcb505f600254fc6cfcdc4d58a472acfbb93b8d6b6bc6c4bea7c35cf5c7ea28f2942b0d9
zf63eabd7bc49721aa6fa461dfb4750a106e2a5e1319302e5816a4854028dc928aa0f5ce6ccc955
z9edac949969259e94f2025d58afa994dcb088d584c159b83b0a58c622b6f517ca15309b26f0b02
z46d4c7756e06eb767c8440bbd13d56d11a64ecf8a7cdc23a5726833a552a43e6ef008af3c30202
z08c5584576ce4bdb3d1d5f4d04410c4287fe8e55a204b17b416d7c2706b115baf7c907063dfe85
z0bdb9bdc5dcd723bf77e5b3ba00823797c660c0307bc9656ab108986996d0246972335879175a3
z00e18db0d8688b0116611a3f8ea99a7204e57b995c3c5383a957bfbe94f0956db74dc3516a6388
z9f2aa531ccfe14d829a4ffc08406e335d520e9abe7c98d0fa298b9bec7ff36aa154d5328895c82
z8c5673535afecbc97286959e05f7f42a3225aa121abc4ae45d570fe247782dca43d83ca3cb0a93
z3532113996f814a5e86c0fbac6d407501fd19cc6403058a3f9317ec84802d1481882f9ca22546f
z3c68d13007f7c957f55bcbffcbc903daef40dad16e1cb9b7228fe8f522a4a117ba2b1b9eb17f77
za8b031f92ee2e0c801d773130570aace0c6c53564c5f9b0864696896c64a2c6b7f28b0d850d510
z4d5c0173cda5cbad1acc12fcc72f65fc51deb8810522ba03331d1114af42be2f6a456b10745b53
z6dd7e8adb1e0fb08507cdb2e91f31becf498a803397ce16a0e81349971474e9131b18c84c25d08
z7a09c194e0eabfc6444b9e6fd894264f6963b8283e31c5951eff2e7dd8cbd412aad916169ee38b
zb32f6d71c3a69c2c02604499d04ae34b1715b3c7b067ca19f137db823f9e5b984773c0d44cc8fe
z120de6f54d6fc4904104e51a159d4ba35b74562930ab97ae3b3cfa40f173a79d0c5bde4ea8592a
zf440f19a0c91cca13f2980d634402188d644b30ff1f7e16b3c43bf740e308f9a8b19e22822a79f
z2b6a22408771883b95f6af542c241a24be9f0cacd138b8f2ef397188c9d8c14dc42c4e68f41b14
z60be39fce1c898ca655dd87a019afe78fabf59f3f1b6417a916b409f7ff0869bbfae11e9a638ed
zcf0104e4b9737b756acc3cec7f123785d4620b83a1b4d0874e7487f8606b513351c9d960f010f8
z2b13ae28a353f0ae6475c99366dec5cc8eb7aa5fe6d6ed522dd193bb90058812495e1d39240cea
zc837c9187ebdee2a73c1f13434b4fd7e8b391431de9f0a88bef6dcac8051277f35476b3c87dabb
zd515f50f1de18ffc6aec5049078caffb3783754b1749865a4c4a11f8ce1b10570edb048db978b4
z2f0eaaae08adfffa03f1f230615f5ef1699f1fb784e12c5ce43f805ded7ee1bcf366839fb6b35d
z5528910e8c599ec7633122709d922fe24226b96b49ab9220fa5b7ccd47676ff8e4a5ae9c66c8ba
z11017126cbaefae3d6c4354bedd631a0e029510ba475ef7c32b97585e277a16013ce05fda8bc6a
zdbc56c7c1548d9420358933f278d4be8bfd05ece3ffb0b9dafd1cdcded85374ae16ac71dcc6f34
z21947a9db1ac0fec99b5777858ff01dcb1656fcb68af406a4f3c602d82c7eab9faf3b9207c82c6
zf4c93652e8e1ea299ce7d1811aa8c39ea5daf9bc091eef83f68a2c9ccfc78c9ec09295649acc07
zb7134c8f31868fe0a676cd7efa632810113c2e00325038f9d542c1b3d6db475baf661f3fa1a08c
z44ca85dcf99b38b883cd4318803ed51e78323a9b50a894aa6d117704a85e6f534ef54d1292833c
zb3b14ff98dfbb35235b16c5901ca82029a875a9d451eb93b84846fe971952093e6d46f65ceeb87
z17dc7532b4994448bc03a99e8b36a2710e5c33829de9b02d40d1e24237ae15d9087a582765206c
z71afa863d923ac63891a7445eef8296c27778181d93b553433f5b44c29ffd2bd08091d54cc546b
z61c6a5d9b8e9ab919d4004a1a85ef6c33f18a9a25768f2f516ced92a6757a456b54fe26bd2dd85
z2adf982cc367cad7570034f4d5001108d155437516e93c00511913d119e6aa3ac6025451d7ad91
z06ad55b4bfab3280a99a91ef78a4015a43552960a14c058efbcad083ead8e518c6c8a0c1c8fdc6
z20133dcd3fab49bb3901ece2d807b01b7526d1f295aa770ab9dd8c6a581e09e5890da8c1f0fbcb
zb404217f3aebbb879351f5e059f366bb230164991fdabe29cc0165131627ccf133c194dd430efc
z11671e61fa25028e06e6d85384b380780bbd08ce7891b797a7fbf6d4366571f94a7355caee369b
z2da68e5ad7dfe6ef8e76126eec2b9a01b7085d9089cb265b070c0da238b50c464eeea8a7286b63
zc2b9dd41aa89204bec5f2682b3299af47da8f71dbe5f29db0e58e612609f560307b3b8b2601cad
zfccbfec951ab36d6d3dcfa5d50b6a694aceaf3e77aa0279ef2f1395bcb0accc4755fa48c67a7bc
z64b081b1e73c03946d8b76be724aaef825b927f99b71f0bc25501779c129655b7935f1c16b8d87
z56315ff680a19ae22db720087f30c93a9c353b4813efc11b7f43f6f5c96f7c65c0d6aa20818ca8
z94539b44928ee1f6352ccf7d877bd215fbef6d494d717f05747839407feecb2a1a33486f4a2957
z690d1c5c2826836544be86957089a087087b507bf9cde7470cb16ac35ef667fdf540962f276a8c
z0ed488ee062683a4c76dc5dad20e2ee13728a9673d57d7377d4926f7663a322961d01455b7ed2d
zbf652bd2b526746b7ffdd7de1afd36ba3f37a565a9b1bf1c7824f09a081d9a3c090f7916330911
z25ee26da1d73e19b8384885b56ef5effe8d2bd66352365cb7267ef3a7b78fb0813f7395a66b8e9
z63dae49c0b6e34ae5ef882189cbf22c6ce1ababe7f390350b12bece58d56c0ab4c7948bbfff51c
zedc5f81c20a160d36bf3dfde743889bb187600c71a24172245f8028a7ee2f3a9514709082b41e4
zdbe4ebe5b75c6950063dedb530d0430838f65684f292dd1cdc8d707c06a1b51d2f6d8f0689bfc7
z7eb91a403de39d4bb7daa53fc5e19e5fe5341daa0ca9b198084aa10dc467097630caa30fafdbc1
zc1cf54d9f8bae55226c030302acbde25616cab5b69967d77f097be65b8a96cf1dc1194ba8c6f73
zcfb2c53dc807cdb8e94f0fbd8d25021cae802a5790c623185c5b69c9cfe2e522d6b840c4931b2a
zf02831088d20827ba8730af4dcddf9cd39fe66f0ebeb72aba5f4814c4d11f8bd44e2befbff516d
z1e10f175c9daa912851e1613dc380e6e2d493fcb7c6da6eba319d5be4986c831ebb054f519425f
z895622dc2fcc5329fe4b689cd98ef8e4671d9218507336dd6149a6e73147e2af5810d4ede6f546
z8c24a3b3a1cf54de4eb86d4861ffca9b87f3db3b95f8cff57c3f2d3497911e66a3645f1f47f5aa
z811b57931e1462baa77aee896470ed197b3658f44921e296006c2fe416aef42ee0192bb1b3b85d
zbd7ab50e2f5c2bc3938ac2105eb3ac90f4c7eee1555c9a5d33d1d146d4e6310fa21fc1970f1c2f
z7ac17ddfe9a1722131d927876e2e247b6b490b8734cb54d9fc7bc40329f74c834c0f6380e30bb1
z831c242e66107dce8cec83ac93f12ae2b92ce1af36e27a0e8a4f9a8fd869db29b0eb38ece8788b
z1867a6973fb87148660d8efd43ed8bf34a85a8eb710e762a63f8c98acfe250a66ecebc6bc1a531
zcdda480c7c9e7050c904a9cecbfed169fd11904d194cdbe8df862b16842a07d23c99d99b1d2f83
ze91f2b388afda2a8257b807a41eb8a47cd076e823a77acf75b6a0319460bac2b97a64f518d44bc
za453946b5e1368975486ec592b54e82827220b304cdaf77622a5b44cc60b4ff9b76254c438b180
zdc31ce7b7776ce1e83a67a42cc0d7ca82686720e959115ed188b6b3dda3f0d88b36b4bc859df3f
z9ad2e2963b5ceb04314918df985bf0614a161a3838e1493a7898b2c111dfba83dcbd2bd41dd20c
z445fcbdae020a4a1d4fb59e923d56b5588afbd7567761a3dcfbbed602f47faa0f9ee372f2d74f4
z1094b667ae8e791a752a88ed9f69f70e3cde26c41ccdc5e8912143500976a68778a9e69137e5d5
za52ad1e62a7fbb50035b51732c1eb7340d165e06b593609e7aac56708edaa63010aca5bb5d8d01
z3882a4efb6009b47d430e2201393d65350961ab0414c067c3f63505f0e036fa59d789d72790e0e
z79d4dfe76fda784eb76e1d5eebb6683a0707bd13460e39189f98f537d6f3c2673229c75784e8b8
z5b3508101eed95e042ed84dbb1440d026b48dec2d153714cd6c7ddcd5377f1cccf90462d75f5dd
zbcae1950141fcd399d1b0aaa4947c990bb5033f33492a59fbfc196941f63d63b4844b5d586d5bf
z281e98ee0905a0a60d71617b62adacdc12173f345f7bd69174fa159d6ec8ea260b0576ec0e69b2
zd959a19fdae94ce99e2cb5e5d0754cba0976be03bd8cd8f4a18353d50e7cef66d79b54253080f4
z2dfeacfc8b0a46ee76d079f95a6cae68d2963d517bdd9bd5d338570dbe5dd95239be5cdd7313f5
z38fa76d4c476dcf4f177cfaa73632e1db19a33d31ccd8c332181bd431405555b22063c2f6191b2
z050e9e289a9bb25f4ed22838f59f7e3dae3dc63992920caaa81da72db9e7c9d9ed88b9c4c837dd
ze056f4c14751c87e1d18689bf16181b20e932d3ed1dcef03faa12a2453f2428bfb2c1e98c675c0
z734ed1363eae87c7e916fead1a79f0c1d40b5a7f156416fe05dc03b97886b6a869d0f3d31b6e08
z94b4ed91e8f9ec3271fddb8cc38a36724a52a007ccabe15e1047f8397f1c728ae552fec91cfcfb
zcd8d36c0e31c0e4b242ffafc4dda1d17dff4d538b14f26997face965dbfc7b74e3a1003d81712d
z67eb9c5ec15ffd13b8e92fca15e0cd3f1c0a18a668e9a55789ba383c6073140c99523495511e0e
z6c9b1c8a81b5663b971eadac3b94a6cf30f745a93341bb39ae89867936c8cb60812b99857832f7
za393defdb4315e8e4d605bcb33a09d5757ce817d37f739c5d0e699aaae2c5aca7221e27b191fef
z546b0bf6dcbce1ecc9bbafa226ba2e3383b47168df6b5b72f51cda5db0703243dc51bb087979dc
z194cefd5981d351e6f563da8bf2b796d77db6fc4c64f61c1b8ee0db9e5a18b9c422bc65ae2a042
z9d132cfa71d4a5958f4ea00eab589c9925c79148332c5536543be964f9904a41e7feea20a9e5f9
z2afb802639aeba43708e10da18c690acc41d5f89670730e53fc26837b893fa695c76cc98629ad9
z32fcbc8d3646fcdd5fa498b4e67b196f5cd48da4777dedd3c3ace9c6c4d6ce691a9abeb50b32c0
z9c920aacadc1e5377cd6926d0fffeb66a861368dc93dd5288540216e7e0e1c301444e013e7fd8f
zc13a561b2618deee2b7ba623c00352f149905a0fa154ee30b681fef68dae86b1bdb645fc77af18
z89762e4710276ae885c19ac0b02b40d748b64b6e66637d421dd5f69f03446f686af7e3e0e0b49f
z28c0c065da160f25684a0c217f98f7f211c6c24b956e2ccd4b563d19871f767ee9778f425c9557
z45fa0dd3a9eb11c0c1849a0e628dd65c9ee9b8cb28cbd8d219df11e292f05964e6049cf0353a82
ze30d15d7340fe953b19a39d6483c40ec6e5b790d2c1a6d795fe113075eead7259426ce3ae4d943
zc5d1b6bdac8609a4f41dd00ab05fb398713193fa50d307d305fb689ea572bd8c3fa1e99ff3c579
z4913d44ef49caef3678bb69edacb54324babb691291634f0b69c53aefcb35950e6840baf6c8557
z5fec7eaa651f1408a6c00dc1cb5f91ab6094e2a4b21c5be436a559ca6e5e5268cf6c21bbc10696
ze60f0780a1525294e8f57f195f96d6a76a7afb47a69c71abc78e9417c6232759a180961065032d
zf49d26b31b37f30c82c9597ba94cae0594c70f5dfdf962108f5386631ba7f911b2d8ff21c3b189
z858ac1838a42215e4d3956379e6b5d6bc4ce12a213396897c5bc646339f286c2c8ef13a68d4631
z8158bec366101fb6bc3c2a82e912d7676a3756829267edc13b10ff6a0512b2ef6d745648363ce7
z6ccfdce163c80f5f75d98f400e4f481b67c888b623015e1ad6b3e2a3ac98fc5a5086700648a0df
zb6aa01f25f0b9450d68e1e21804dbc5d6867cff9cac313efc59f494a7a48eef3ed460b0bf91a76
z812fedfd18d54399518144e8fd3a11d76c90df4ea1ce7e2b7b4228f4f917134efd62cc12d29665
z935c888146d0a635441bdf15e636124219b7b814f22c15b87d4637e04d5c35fb5ffa8853c87a67
z5f321b1e98279febdfd63e620b21ef38799fcb999bae4ff36182b955aea2742dcef713b06d631f
zda80408f423ae52a799591f9e68b52739445dd49c9cb5b6de5db07f170a253f425a7cfead7ec9a
z73ab17c55741b033608e04cc2ee50d3fb832b7b877fe130ccfce75a90020fa825c80bd8582bfb7
z7a35ad31c8cf3b3deda1ec61808a2e9d27e2ecd5697d1f94da43c029638a5f08492a052a3c2bc4
zc1a703498fcf251e7d153219cf41e825ab7f57e48f904540b8de9921da555ee6287506124d8e39
zfe05773ad551e78d2bf338eee09cd2eae448c0ece08918a9376e20d58b45e633bead98e4368218
zf4dea0e93a2030ad421482a574233a0ef5ecc2b6bc97e7969e64f3da2a6a86cffe1f841d443e2c
z845b017f4dd1959f5d4b21e4d10bcede26d9be98f59d37b2f0e19b57fcc865a17e472fa33731a9
z3449e500c257044c29e906f8363c97999713a4456c0caee97153c651e28e81753a29e95589d934
za46236c80d2e7eba73acee6ccf17958b7f2505b86f15752a82d9267d5f6b537a7b48e05817dbf8
zd50f3531c967c35321d9f0504eaf969ead09df5375d1b3bc190e1001cdef05288cd92d8366a4b0
z345ad49d54971073ad57e144566fe4dd74e275fbda0827cd1e863630f86db8854a7b0a6b172410
z936abe310fe58a310d1d55118815c47e94e6e8f8164cd172d9724d251eafdf3765b6d031d4f14e
z613a3107a9887b53c6fb74033ee048d1c150ac47953e3b1cb90ebe1a9763989c030f2c2dc25922
z571086dbe3c12bb5dd7ef8ee8ee012195e3e76123a78cc09c3b7eeb8ede7b509dac7c2cb364b8d
z67233da904b4a85696ee7097a32d990736431f40ae88d49a7b86b0fecfc35dfc5ce0325ac24543
z7f58dfee4e554d2b93952f6982046a3eeec4c67f825aac4dadac18d4f790dc1985b183e054da5a
zf6ea904cdcab2809ad279b74bcd08bf94ca1f51c4dc5351bf540a0da6c6ed80f455981e274bb92
zb8bb973edf87a3adb77a2de48cfb445f28093fc457b8775ff47be8b001ae69090709b50a879cc8
z9409cdfe42ca92c50f091808631266000bd8f4ddfcb99f956e76a1266f06f736c36dec45af97dd
z248aa662900b075b9c0f4172f9e6c0c7f3bb63b64603b8915797d8a2539bced94ce5547efb6445
z1e5ec7ca9068b7f6947390638e2a287cb96a3ee98d9114b8d5962b141a006c238e0989daf8cdaf
z25e9db95fb9144d7559a2666e4c436aa5054727704cc31e6f50cbf838ff019a6f832a1d8fc3440
z140e99de3121b30b54309ed3fe2861fc7c5cae7b8341387c63774e9461745c34eef14bde0d3a71
z77228305585e94640fb66ddc3ca5d8cee934d18c0a619db964d41226e908568ef7155692628d10
z6e88ad1ac29b27e7e82c89ad0a6247cf9670b4efd97c87db69c7c1c5f3bb2aba6ee2c346dd6c33
zcb60534e1abbf6249a688f4eb006a569d8dca0945d4db6bddc6d7fa9b7077134a3efb452e7cdc3
z23735ad476d96b98bb4cdf984295ebffdea564e7b6ac8c57d45344844a7bc2f506954894cb9940
zd5abaf29d1e1fe580291bdd3dd925a5410abb88237ac6db752c123902db8b9742887ca38b6c6b8
z3aaa069ac920d1192c49fe77d59309e9f9521e8942cbb60e6f6a8cc8d7a14f38180463122d9d5f
z3141f0a8ac39b1c5f017b068f688a7867a4028a1c6988ecb4501cda0e6cf9cbc5bc5cca48809cb
z634762114fecff5c669119dfdebfa8669343df08ea3508434426f5a3c7b7bbfe3c15f32e15f377
zeef7b7ab2677a42526408285361053b5c4faa2c180d71354bbd24db402de85fcf0b7aa8334ebd8
zf59ef8037d35beecaecfff7c1be45c0f6da3fed189911229f39b38b0b4fbe30b987afecb7efb24
zd1d330e34e9e9489a0a69760a98c463738e57f6fe8cc37517f6d125d5b4a89cb5848a82e5fb9a1
ze8efb83c850439e7660adb117f312090ed91814589dbd9b702abc44b7e7e36580e43a8b98ed047
z61eb1026fd996a7d5688f084d7bcc0d724178bb1cf8ac82d98cadddd7e700bef754ff1dd33ff32
z4786e6345b60aa8906e132f44c18a423cca70b8639b6995b8ff52e6a87a9804ea9786775f102f0
z51d79e210192b44e5123f44822f25158813fe5c426b0d73e72ffbf00526a7ac521bc2e415f16b1
z63cecb40e5569178aa512768abde769aea9fbfca1aa1e831b424b00f27ac65ca97a2a29c16447e
zdd876c34a347b1d3697740c476b260974ead0a22b26be13e7d0ee65bc12e1c9553d1f397713885
z2fcc2a7cd2c638cb965f81770335517b046819d67ef4b4ce455c4099202c0d0e2c11cc0b4b5bc8
z6b892f90b5b084cb5ffa27300b347d6fca9e0461003d77d27bb55668a4b9cc91e40708a37c4ec2
z56b765651aa0e6415c3605ada78a3db223dcdbd8058d024090857a3dba53e650c70d6e9d349132
z11e19fa600d453d60e062c00a2e12aced818e0ca7cf0acf143b0b3c66de555a3afafedb9f0d2e8
z5866b9cea52b4e2b588f99f4dffa2f8b0b0273d64597dceda78e1cac8ea25c96060e442ae65d5a
za5c5042dd539ddb3638d0fd4f22fc878b303fae646c26f636b109ce0db413bc66b402a87b4c6a3
zcfbbd56c0afac8f8571c9c32ac79d61e13d4bc229f53e18df4b30113ee38352c407908bc983a1c
z02e29aec1342060d516e3cffea688a4f6a2fc613a63d18511bc3e75692dd889540820a963eb18d
z0c942aa61491aafafdceaecc5037cfafb5a193f328bbf7c2f587a871aacb33679462d0d75831e3
zc6a328b78213474a8d916796adfc0444331fbf210436d15961d75f3b09d3643984d4f123ab7cfa
zff84a86c9dac9132710fe1e2f4e497987a74ebef9ce86441c477a62fefb1b7968b2621d6710717
zcec781a82a017ea8800ee5eb9a907300ce7f5a4c5af92db727ab920e54576823e3be2412c63fef
z3b666971e7320ec53de417ccabe990def55053fb3907c7f7da86257f80390468a51e38c7345869
z5bdc18d45db96242a7db67aced1d2178f45d1ebd2eeaca89957d4ddf2239cba67fc3f8465cd546
zffa0b6b017b473b3703066608afc206b0e4183c7e3e8330caa3fea34378115d3cf939306386c81
z5e83dab46aafca6feebd0377b285127587d44dca7532dedb9bb622cbb95e6b55fade87e2a8de53
z0d786da90d87730748b79ad5cbb2f6336755411cf6e7ced6a60fc4741e1af64e3fc74ac84d3653
zbe45c6a5a99f40e1634bf224a3cbf4f9a949e4c991d83c1fdc75bcc202e0a4b09f273c3e4189cc
z190e7f6f2df22c3ec2e57d9a9b3a99d5633c1cf3ea514542b3a3dba836f09bac5f10670a85a2a7
zbda886520f18378bc798126b332c255dd2f7bbd6d5329e91e3dd8522189d721c9ab9cf3502cb1b
z303aae72705977176dbdd626c452e14bb4ea095c27af2f24725ab8096d00929cfa7986ba34f612
za681492d8f9ff04caa0a857ffe050d5744efdaa5251e094d34df148ebaa2f832830919f4c41f9d
z2061256411a499cb0b3a3635932859e6a2d74ccf232e426c77b2f4bfec8262962c46fa0e1df385
zd2d821e58baacdf3e62c27e9cc2c83df4b92d843043664c41c46de492080fe0ce8f86d79d9b0ff
z145b47dad7cf83c96947165bdfb95a95aaf2a52e585a8c7e7ec971eb0d3fec0db7dcc1b9176e8a
zaec7d2d0883b6b223a7f0dd48c23e480d2f58526f3c9afcdf7bc24bd013b1101512fdeafa8256e
z451fc07c63f3886a4494c42682f0ad3650cb0c8b42e1e47dd47897e2dbb6b6ccc0e484f624b72b
zd62d0c201d57c5a45cee07fa6c87701e90774e54f58b065796b40d069c2f601f4e96175a9bcf9a
z43a362bcdbc83df71092e7046b5208c01c46eea3c2f78ba9fcdac5a2a9f63857309709541b3c1b
z4df1c3e871efddd97a7f500144422008b67c2abd2961ee6c80afc652fa50a4067a898c9ddb5222
za3d7e51a851c3bc57d07b21b05b75a49f0e1bb4880c10dd5dcb7c6f2480c6e4edbf887d574d0d6
zf81d239a044786314d86015d75f094a5557f09f7be984df78b765e6becb290248f0e7f65976f20
z0168bc66f7b4964e14975bd300f3e95bc5ffc6a03cc3469f2480994467472bccfb8a29e8195e14
z5b11d33b34f26898c36643bdb98690c8d8dfa5389cfcf016e078bbb59fe4284fcb634593a884d9
z3349f559700312e029c692de7ceacc27499f15dedd9ce3a8dff8d4172482a605e1cc2305293591
z6298c528b6e6da80c120093a94d603a6cfbcea2a7b497fd16eb3e663dfb1818ff17a4dc6911815
z2577b2718a4ce4554065e001115be918a61a4f8c2ab219e275d54235eb4ba1714fc5ccb5f39441
z685b286808bf344e1976d5a81faef6582ef4896c2bfb0b60be0f40f88d86d5de26ce3cc932b8e4
z493bf16a5ff063f23c60bdaa6d9e94e10fb3f7a4cb28aff5cb9bb34ff7f8fbb3bc7e2dbc50c314
z34ddb0c8e97920611b02a22acac0d341e7b81049dd31900acbb35866b73ffacb295484d16645c6
z00d2a37c0362ef1ba9deb4da61447569324979930509b6d728e9f9bd8f4bf8b7d7a62626155e0c
z1b3b5c58f10a93939122a5e41415735eb0924e47d2d78c5ffcde53aed95a7d7b45ead5c534bf1e
zf524ccba185263eee8eddd4fbd489b1c969dfbdf155e72786de49d0462a1b793f320759c5760be
z3d2fd023a6e6cd61cd1cbbccbc01bef594771f694e2f97ee5ea55e9a3cf0a8df1bef89e2960aef
za4f21c71a38510f6dde227ace03edf986bd9134ac4bbede359b55ee808c2ab08ff0166a46fe01b
z36052ceb575d4b6a435560bdddcec01d6c1dc4a5cf24970e6ffe2b8157f026edffd148e9468904
zac07ec061343553987daf59e8cb37d7c765e2d0b6f13cb9a768955cb8d02291f8d46444796ac70
z1e915857db5d2c425ce13f8341d2f411b749b04184225358838b83cab4dd46ac0d8d5a94763ce6
z7e46b6a01a2463153bd34667c68677a1acca8b392d1e1a4ef37e34fcbe85b79602ca5712ad5100
z5e4fa3d24f6eca1bbe467e50099a3dea879b57b8c8837a93c6fd12b0ab806ab6b670419d955f96
z941cbfc17232d05c2ccc0512a1e88561e082c6360e360f4e25d69161f1455c4722ccc9ca66d4e5
z5c60ade62ce0f996a7b3f5f9ddd6ed1cf03af29fe685bfaf267115a2090c5aa1b55ddfd4ce74c6
zd651ab9f6a378716f553d85d1448d4b222f4e76021c83b96413e57510a0482070d634e5bc19738
zfecfa08173091be26af616e23ea89a00b9f092522c9f03f3ab3ccbcb6bf9fbdb4d509c792a2c72
zd163620d493e1b66a379ccd74be84c8b01f524fcc425472f1876f71c798f93722f62ee46d33837
zf25bfaecee349bfe7a7934955e8093ced3a920894492f7771448ca3cee1c953dc129af4bb01fac
z34b75da9579ba7157f6826a4f4e992f4cc297f31716ac0753fa58ac9addda389b6580ff1e87c2f
zeba98ab39c8f1121b811996c516adb1fe506af92aa3a0147ba506be2a81b1ddf2b52dbbd5a8739
z6bbdc6e15aeb555b3aca5cba6c3e23cfffdd9415df95a76960d3ea910eec107127626ced0e2df2
zc72d30adb341e8d8c30fc34d9746238f003f178b5fc98574433a28814fbdceb20007a4f3821efe
z71895da8e424c7a335e936f6f2e2fcb28cf69d8174f66d05c27122fdf04b85cca51a367a7c8454
z98d90236f2ec89c6acd2dad486abbd00a5faff477ec2130cd5f2cd3f2991be19462dabec8281e4
z56b613c232571d6342b9e6996956b502e6ed7b0aadbe1cd1993d8b737191b6a6c0e2e083ae864c
z6e192a926c1c9d9ddf93d4df316fe0751930b3d4390dcd2687623db75b0d15956de48f3af512f0
z0ec2e775da6615c211d5991385e654c7de7dbd372275515873e917e777e779683b927f80751b66
z3f3bc70bb1cdcf2fb705faa07ef08d88dcb3535e5e71df27397cdb02c9f0f52eaa59548320dc05
z58d96d8a7121f350fecdbf148aa5509808c198ab8e9c8cd668d0b88cf81d40e5c549b470e6044f
zda87fb74f3aac29eeecb62699c54acf7b31b23a629286882c98317788669acf655671dfb8f29e5
z87306331c90e22164bdefcc57a29bb813249ba19e6ea840d76d09e5db15bca2fd7cdc26903bf16
zd6cde1fa2e51f5583678975ca5deed2b0ab962017be8079af0e6097482012be60cac0efb197e53
ze93f4f95a10362ee5e020cf9be987b4f2a0d701eaaf52bb1a447edd0ded7179cea62fa4dfea7e8
z7f9021fef6d553edc01c97e52ad5840c7e88fb959814a6ef9c79611adc36631b48cf55771e09a7
z1829c19d60644221e0214dd0c26c92e8fa026ed91311b23e08e86cac0c5b9eb26021081b1fae66
z8d9094ee2b5dd3a23b83385d1effa84323a0b24183298f22bfc1bd5fb5ecbe4736b8eef30358d9
za836c2b103088412335056f78f77d0d02acc1daafb29cbf1f4f166e09b484b7784797085c414db
z417068649f92d33d268d3f5b84f0f106580deb7abb27f8eaf5d34dc4d3f44b9206b55d5789b298
zd2d098e17132e55ba908e00465093c51606b2e9c034e913c50eb11b07338cacb436be9c313e49b
zd929417b97f8a5bd5bad1f56645327a4b1888103bfb55f66967b5a47644936a900fd9e06162f88
z9d72508be352fb6b789cecafd4cf411668215a61e235db87a43c5dc6a8b39d674a579612d2ae01
z1ed9932579dc1920fe96a090b70f068dd54d402fcb9436d002fe121c2224ab7e3a43c56bd3167d
zbc7fc4b73cf79514075014c7f551d3eb8d49f5bc19a03a5b55b6ed67b08c79f400728c7993d437
zdd5fa3e59b28d70a5c3f5d6ab3086fed8110ea90884373a4b13d38d85c9d76cb3e364ce2a5eadc
z589a7cb8efb0b790b91dea4af453a883086dc8ae7d0036e5b56caf4cdbba1bbf7947ac8d6528c8
z0739ddd49f2544abcb33504c4745face7261b84279770d50640f6eecaf1bd4f419b7d50a7a3f22
ze741acfd0424493856fe1c4ab8a773b2560e819930ef08988189c40daa4a0cf22ab4de95da33ca
z618ab596e9ec524d5d33706bf26e443917ac4f927d43602a4e0973a5e3812278053132633e843f
zc1d4c2c7be58b6f22689544f34c6a194ca6fff4ee116e7a7634300e7e9349dedbe44d282e2ea18
z36350c26af33ef2dde22630f475f6bac720f64b15dcf4e28c7894ee11714af2147dac25bd814e1
zb23578951d17b2028d54af8b2da950f1bcd43414f8d17f4c1920d98bbaa8d733cda5076770d593
z5b4fbc7272fdf7919fbe671a7e2485c404af6df340545daeeafe75de7347910be5b2faecc3c581
z390992e7eb5192ba10b859f94f6bf2ace7a819bcfbbd77428067d191b0f3b9cba46986845f5a0c
ze7a7015c807128b2100584c8f422860a0fa9a55aff8a9a1dfa47803e7997211e1e0426a57b20a0
z2be1ff6162beb9314e5606f8cd9739487c7ade5b39954c3268f1530ee119c157e8063426cc8777
z785fccfe17f4d0128923e47511a363695d9b71d3ba6ab91e11acf976de663bf15aee935c75cc26
z4f8e6fbc711e5001e9b252009012cf502f8c610ce7c98c29e905ba63a271a29f8d20ed05db58c1
zdb2033ef42ca7c7624e41770554abd4dbe308adc61309ed37b131b0db00d674bedd56721803bfd
zfa94227b2c3a98010acfeda6130174e80d9133d4e772bab36c687730ba95ad521ffe5a03e8a6a8
zff19b71076fa2aacce350ab416f5e0de02422e61103b8cd57bf7da3a415588f3651c83590d8c54
z042f78472cca820f0560b72e155e572e653a931db4c0d40b9af56dca7174f99a265b2140b7dfd3
ze55a827e6778b5c396e185ca816a3542ffdd48b54a5cc87a48d8cc5b2e8ecc341a4f1fb702b28d
z0564f43f9fbaf45b25ebefa3e56d62ef0742f2eacfa0a824d554d9cf54f72537c74d2b5e315fdb
z507bc441629c3a35ce7f47ff0b6aa8559c226228b1e0f60cae63917f12de0ca4f10f9d644ae4ea
z682457965afe7f485ce2bb673daf3b3867f55a3566cf1ee367c481e582811d373de954f5ffd18e
zc0d130246ef351307df76947f07869d7ce3ef9a9afac663b52f68338207570a17e053f367bf068
zafc575f3825560679d8b69e6bf84a8c2db07b26515f0cf46022ba645b9b304e5f0b2b825e1cc0a
z05de1babc07ecedfdc14c6708820d2e35ba9a6c1291cf941419cf35a31fb1e09f7879166f6b12d
zcffbb705eb1f171681249972c6a70c80892c799c7669ad20afaa17169195faedea44fb1fe0583f
z1f8e4614d91b826c6f9b6d77ac76dd7272df4fe4072e48a611418b193f98fe5f5979618f486525
zd08c2d5a3d685d426d688b1c591e6e60711c5d6d81d218f3c9e96548e8b13cf2138100202d1edd
zf7d185352eefbb5f759987d698b645f2bb8f7046a1d2b4878651111112b45075eaca837de8cf7e
z8d3006174668940d16acdb719f73be47c52d81ddf21b12cea60af64e35d75cbeed0ba26a04a22d
z40676e270eaf91b2bd07d1e7127af21c482eea14daced4b40b10f749d05bab31888444ba2fdbd0
z3d7b4ae4b73d3ed20627ee87a4a403048a9cf6a53afe6172e03cf8ad7cbf93d685b18316d8b03b
z1ce39675acd28e6079fdda2fcf7b9d72467a1f10d939b40bff2ebe3eda0e1fa5a621290e490006
z41e9088637acd5d684eebdf177da9627ff5a6a2c5b0bbed7078c70e587285f20ab7c1ff2aa1070
z81be5798f3879d9a1c313e357570b70debe1a4040c94b2a77c5a642b7068c2920a3e7e58faef0c
z5b46078e8f39023e3f084a191cf8c0c97952322ada4ba91ec5a8ad94d41206ffd6dd17d6a6f0d1
zf7d73f44c3774fa8a1490e8ead72c5e226210157e8f8306cbfa5520f8b8fa01ffb2c62e1386ea5
zed8253cfe8fe93cba4d939c4faf2270aeba1d352a9eab80397d7f0869dae94aefd4ee115753a5f
z1209dc595c5b3ce6d823a136b74f84dd02b3283c63fc79c1a5448bec768c436da846e18bdc0461
z23a5cc4a7b63d924debd455a321c3aa306714fbf202b28c204a8d4898d7e09dd3b0ce850de6d27
zfd2e163ef0a638661cecfd90155395ac09e727073a119ef3f1b06d7ce8f096857c4f8b7927b7bc
z9ef5f89e97c4402b15734faf2520d9bd78da00024b8b1f1c3c44abc51cfbd8bb2d8e0e1cb2e176
z3cd5aeef87179b40343d848461c499e83c129d6a49bddaf5de9e06e33dbac539424b647f85634e
z63970b5129258db7d33e78d0c280961b1fe188b3dcf96cc428a2ce8c55bcdbe15efbf846107406
z2423794246fa8140a81a881a4450732bbe62b6df398dfbfc0591c7359c338d73fe7a5d5618f96c
zdbc4add76fdefe832f72645f90ab1f7d22fc3db0e4005feefde208d38b5174e8212398a9f6ace9
z41f8d08720076bbc1371be45a0e176726eb00b6ca3de2e94f92b4a691b76ea9e9be50e450b7f32
zd5fe97252fe79a46e5999670820b6f70a6fdc21f9a6805adf80c3bf88730ce4374bf4a649bd9ed
zcc397c2c0480594a66501b2da68c39a33863a526791d4c6fb906f78657fe0382cacad958d72b36
zec9d33aad5eccab2181eb4100e4e05edf9a55806aa25bb2c1c7888e47620925ca7b3e4850f8038
z62f79bd7bde7c60a7e63fc397f1b04cd421cc16e22094cffd1684fbf68f8bcb6fa3a806db92407
z3ad61abd6dc9944f75d9adfc256855633a600ec247fb8dc7a4d8ff511a9068c544c5400a342022
z082feb4357c4d95a71b0eafb6b8dd9b7d34b50ce11ad78e4406a53f53f6d0714288a17929aa63d
z7bf22cb61926bd446b677d45dd706bd0819c150bf23453750acb542fd7b7dafed12db3b998a92d
zc7e46920b5e48eb8fe70c6d6700805a48bba13fc9134d71c64f6e50b72898cd0985bf8ed53ad73
z93e80ff54b75d49d54412e84ebc24bd4b559c39a1079c8c1689dbfe712df801477153fc28e6343
zc7fac25031a27e5df22d561bb88ccc61623a83848bf603faddf2f45d329ef4c281a0891f026b07
z33487a4639cf98df7b31b8860efe06f00fc6c7c75d89c5b5675b37b9fa68a0b22032a938739475
z6680070e4dec0caaeae2336d990fd66e0c8f583dcc0afd4134d3d5d0bcfcb190d06d16549e8ffa
zaba4f178e65d32539a88f98afe13042eab071e3d22e3df0ae8e5e12edf62b3fda21c4a91fac4d5
za1a8280f20275f3a970a589267a6660f8cec3b325a9edb2ce29a0e61279d3915f069fdcc4ae592
z62a10b3a461e38bda0609c31197dcc30d199a8257f124bc21f03990f7d15b7fc84574c65be850b
zfd4201f10737083fa504d7a8310613275d82332c1c3375d0e6de3c21152dc17248f512273a9a24
z8717b97debc85e0a01ac4a077c69413c683b6d54f977e3718f972af6352105fbf875abaf1c5fc2
z94dfd584ce2f3c1a6ac1174b59415999e864e850f94005418f982c48daff2f03743fbc5ed7e22b
z6c5f43fe8ceae811c642e59a8ec9980a1430064ae35a5ba597f533a76e656be65a6858fde137b1
zbf51b324816fa5be34ca3b12fb2e13f8c5c36be6b9f72c84cb878f0f70547633d1ac86a37be519
ze5cb05529d20fa76454eff05bae23481c38011c26427f7dbe9b80b2c9e586f3bcca448076239f3
z7c81ed3302138d868b88f466e5e44d27fbe70c37444dbc7e87a8367ed35db73e43e96ccbce25ec
za9f89aedf5d7a88366d0a1006c70bf79d91b6ac0841db466b7e200f4d6313c50f73a34682e4e07
z6657867278827655a93aa0e7dccec4a6a68b16b26313a23d2f53cf5869dd3e84a0f4062add96c0
zb1a83f4d9d2101080eb547b151944ea49755f1d329ab15ac696d20b7b01aa7da0bd27fb19ddf85
z821331e2644c2e865b4059136e7e784d94579368f580240bdffc25afbd01ab4461ce5e1a591e96
z6fed820b1f205cd959ebedb5172d4934f9ef700c94133675feb682ac1d3d8b685b0ea71c90625f
z5872173d684a782a5f4751dc1c39860bd0b58501ea20f420432bca626b9a92120a62691f5bdcae
z19abc98f8bd20a2044d758d7f27c39e74822609fe43781b69daf307ac459a1cbea9102aefde3db
z8784442e7723a669d1e03c793e84ce09d9b7fe51f3660399bbb0cf4d875b66e66d1d5ee439e6f4
zb1ec96e7c19f09237ca46c549eb70f2952179586b82f22812df0775ada5e8b953c97fc94d4b901
zdd4c511a3c96f9417fa89d0b1981c3e602dfc80240bbd16c5967086431c0c7b113b7b7806c98cb
z21979d3616f8f0b949e63e973ee65669bb790843081ef45a61b1d9ae65d7e0241f3990ba63bc6a
z8680ecc1a2eeba7b767c782f7a5b1562ed46ddb2d8157213a1b3598c800f4a78fe4301be950bde
ze885b4890c2fae3aec9a9c1f8bf6744f82807c1175fd5ea34a56a1ac0619814bf9e931ee38a375
z68ed428e5294c8edad9c5befa9e761c2a4d74f4fcba655820b1ee953ed68808d06032938e69261
z49dfffb30b513eba22c4345a8a8867d97638ae86c3d72edc72cb1f2b872ca0d2d3c03ee65962a4
zfaa59452389983043b752acab863b8e451fa44e1a82d856970c4b013ad35b159c2a6db341def24
z73e61034f9bba29f41d0159a684f05c57829701ff7b7afb13c90c4c499886ca63b6df33b6d4542
z2e2b2eb7c0ec0e767198f5393524244cabc826e22fba9113e6c322c171c7caa11216d3f84f9af7
z9df006717dbf2ae0662d0aa695ac7fd20bd5e9bae2c1c9a9d5030ace144b263ed8915436adb692
zde8e6a76dfdc70c55dca52896422fe6374fbc358e48d5835d8c5dd5c7b9107dbc4f0855ef257ac
z2025964107e8120a57091ec322612cbb500cd53fde2f226d5013caec9d24668f2502fe96043b17
z5447497336d2f23a695e668ad4fe456ccf5ab9e75e0238066a19871bd48b08972753fcefef4547
z3e88c0f18cb5d46f5e654a66e7706ac192a01d767f1957c79ee3053a9677b190974965c294650b
z95c704167227166fd700bbab47083fb94cddf096172872df5f2902a3e5cffdad78c725aca3317e
zf85dfa8ebd930c2d00799cead88e4e7545e1fcbd176adf0efcc4a3419c0fabee5ce18572f9184f
z155defb3ddf3535907177985e075efb361efcdc9cbb5e35eb56a0c1e1ffe0d83f8176caa7455ec
z94970d57e9b79f1bcfb0c8d58fbbdfea3bf108817a1b65f9c8870b24d462f07228fbee30bffac7
zc49ae504a9797a999f1a3d145c4934d7d192ae7bad3994fbd36e9e4c75a4a451d69021b07b850a
z50ef73ce0cad5217ec3020ed6644d4b4a1a4ec161afde3d9229f24399c024dd436aef8e3a7e2a5
z0ea11db5aa0af7ba30fb02385e47e755bb545bd6de4c021b0bcdaac292fe49d01f243a4a227eec
z4517e166b97fea7e2087938002131c8adef01bb11a2a59554ca35344df6b60944467cce6515584
z0cd116ff67db5967496c5024e8de58c5724dda3d18dbf779d65fcddbbf10f77fbb083e311bd111
zd7d38aa7c28b183f64e3407aebce5233aebe1a4790be5c8c992b73d3812c82d378117821dca9a6
ze94d0e92dae5ed63c811f67e0c4dd5a1ab5ba2ed60a4d7ce215e0b995e23a791265293be44cd9c
zeb4f2fab2d26e5d6495ccc65e768904722710b539b834331ebdd49fb5fe97ad41481dacdf8f25b
z7c97af387d4e70d5357efbfd22f9fd33567bbd547daddbc9f69f673618a6776f375baae9b1f4a8
z2a8a5fc7785a275d55b87087bca9193386c635b26b595ced5ff74a5bc081ba3ac6e0c763741b10
zbf197f842f1e92fddebf245ddcc75fd05e6a0f7bdb7733f17b307b024150d4e8edc47695a54ee3
zdfa690dc3d746963401a182dca76b0e40d0704871d0602cffb90dd30501f373d280027e32a8b0d
zd6c5d185e35519bfe8a2df4cdad62ebba50f6b9989090b4597b53fb5297d9eecb294fab3d51adb
z91ea8b796062e487e3d9bd265901c7e20e7f56001f83a6420212e2fb406c946bc97c86a61b04eb
zede168f3c14ed98d7a72da67e788f003099c12d15b25428904729d329ecd7757684642419282a7
ze9f17684b0f5fa09341073689286b09adc7656814fafd1b51446641568bb75c2ad7baa7e2199f1
z058b871391fd0e5c0467c8197e1359755e3f3067236bd179e935761eb8e0ada48f2ed2079ab91a
z4c4a61b93f090d9f36f54a1e28a7014a9974581027cbde2a20e62d346e6a6ec60f97147d9683ce
z519b8fee7dc7d10d61f3aca29d1e4fc1929335af91811fb93d60a057d4d568128c796931968e09
zbe87a908d6773f6b9cf74f00fbc5e733fcdbc98da09ab69034dc5740e806636d23c15b5bf5bce4
z55c4193af72a27b3aeca5dcb2a8af8c905d61f60737d3929791347bd2782447ecb80ed713d7bc1
z761bc5a5909e8b344a817654dddd52ecbd8f06ceefdc6ef586e271b69cd2cb3bded7ae17f8772c
z746fa342b0434808456722984f1de4186ffde44165f8e96993a0ec0b9ccff90c2a820eb4843e6f
zb35be44e9aff0ee53ee74f7a6ddce2ba5332f4d872b1ceaa0d8632bdb908ba72758fbb3c9bc80d
zda61152bddb6f0ddb2c5db06e2b761388509480b61673f0599e51ce8599da8fd913ed2338dc77b
z206b8fc80e4a585978c0c93769f7ae4b86cd12d7811ccd946d3f1f66ed9afb1a0d8fca174b1b5b
z388c118f00067feda0febc449e73ed571a6ad91b3c84fb2959f7811252205cd88f60b72fe2a9a6
zd0dd2d56ad2c128ee522345180c13451c80c24135062a75abacb74a239aa81a023382cbb3e3b57
z31618589a4e73f256408bba81310e2509157adf05605d7048372f322f04453ef873c9f6759b862
z89d17cf023acc0ef96fdfaeb9626f1ca21b3740c710f27316b008d1e99c5150d704ec0b4ca45e0
zf822d061409c51c468c19eab4d18e9711019e30fb4a21cc9e3374d9a24f6622f74126b0fe731ed
zd43041e6baff40e0bc858654784c3c6410d659748d507fd9c495dd4bc85566c43c384b13fdccb1
z1b416d30db495af22f4c440aa0ff30852a885037fd393bcc2e6cf333284e98df75d136abc4771e
z91f1e273e813a59abd22542b9a230a4620fb0f2e9125a84ab20a7d46865dac8e905e80f0174977
zd03ca09ea7a4f19647e7c067269fa1cb0352b79bcf27092dd2eea4324d86dd25438afe6ecda517
zb7788b3e2423b743012b18bd06f59f3fb87effdddd939758358383c4882afad137ccdabbaa535b
z2475be7c3b3a99e2f5698696fa5d07accf8abf4f3f2b90fd14b434e1f46b4f04b406c57d6a00ab
z2af9e4225b4c626be5029bbc9b221a8e78e213b957274064acd058f72e6fbd85e75423741a3b89
z758ae266d444512fbfbdc0ae8b1b42cacaa6632ec98536a2f5e0a4468fb6b1179e8d44a01fab14
z03e7e3997a0bdd3ba8a7d33e5c7b0d9f9b31281436097ae5b663d147c7f1d79f48561c6af96fe3
zd3b40c4b23216553b7ab3933ca71d285aacf60f06303947d54a03e6eec4348c8bee89e8305f238
zbc8b5d580da509ba0af1159a21455f6ceabe516ad8b300bbe00498748adbbab6900e272d88c19a
z8b7c952199187a9f39e22748cdfb3a0c60939080854dd9f61c640f6f08b5fce20d70c6ad0c0f22
zed1e199e7d69f4b3c4afcb86fd5d189ac4c432838bd6fef8f10be7602c0004bf58d727acea24bd
zc5596212e7e36bfbc476575caea3627dd787e15266d7650a2c85afab7968e025530f34feb9fd44
z8b4519bb67c6cdbbe4b1eda885b09936e5b60f926d8196538ba3f97c02175f2b71920b27f0af1c
z934172b841657c966025df0fb315cf48d6e2f740b35bef0c96a16e6e9f8370b9868d11557e2af8
z90f6cbf4f82b98d414738a72f4e867202d705c81234b15e15cb0f0f570e15166e8160490be1899
z943a8766510b510d93b17ffa3fdfb61caa297a1a1cfb01886be777f3687ad794059654e336a320
zd331eb83d7209b1d6a49fa34cb24fbb0e56729deccf9b640ea0aea9201ccd24163847f67d10506
z3dcec96d137e71cd2d818585758dbe92d34484a69b17e64255116a1c73f158d0116b67f9ceabe9
z41b5aec6669e54d92100195fbbc9f98665d7fdfcba9f44f275c01a7d84237bc1254af58cdbb96d
z370f24da085ec45ec1744b04eec01fcace1b429b1cd42fc70e9f528b3c316f0437d26b59ce11e0
zc212edbf965765dcb8ebaa92766b9e13e3c7cf206b54fcc8c7d3f9b6b6a1dfc7a9614ba12b1a9b
z3788fbc04adb697c6e1d7bb024faef5b9cb966a30c0d02a4d27ef8678285c0675fb674a7210c06
z9f8140ad24e2a20cc2d2a527748f619eae556784c609bf3dd5e215e96e613a48e7e2561979f618
zb24f021c31742dc5e39b3d2c79743e81ae23d44093d784cbe944b40748f9a56802af566951bd11
z05739eb6fc52ead7b3c4639dcba5e69d87320a7758f809c3e9b127866833d8a4b7c33f6afc125b
z2ed6ebdc7c4f78bbb2e2cab43ef70731d625307a96eb0d0302003fe63a79a8174a0aefc965181f
z481f5cce746f4fdfbcc975123fdfe4a7aa59a2acbd6e6f36b9723b8e1452dd4476117d7fd93a6b
z9db85410a81f899acc9737fc5400bc3109e76c74f062f0009050d3dcc7ba0d2129bb627c3287d3
z10dbe87ce14e5813d92c1273630676b2a791992b31fbc5b9df17a66dee4ce1c4bfc1d5b1ebed64
z8523877599927de1557fc1c52b9af950b1ca477b49b153d821e98bd9de05ea6d64b4880e6652b1
z716a8a3a59b435d8e1600ecdcc44c6611fbfbf7ce0cc9671b69c7b410ba1baefa7ef2970393d37
z380626cc4260d2fd13440ad0b5b8c5afc9acdb30b8f5a4b3407453166fa813e38af070a06adfba
z2f60887334f903469c0a8a40e5c56d0bfe28a6d5656d40fd8c7a159d4495125575a006dc0886f1
zdceddcaac465a390771359e4191c4cd80703ca9b5d1e6691ab20100837e70d868ff87327249447
zdf82e38b04f2c9cbf9f6ddcbae3abd4c4dabd81f74b794371885f432519ec5f8a52134bd16a98b
za1cbc5bc0728af861c54f734e861b8f644eff2e263eea03e2def747163e63eae5f47095a2353a8
z4cc8fafbc3d20f38a61d17f609b2d581f3b0915b73ae18bcd25cb8fde545749e096054a5514816
z0085430d6d9ff9c53ea1ebd43c47481c38e3f4421368980534fef6c524ac5b27987d0ca2b72d3a
z653ae5c720d0ae0edb02f4ee3605b99a8697f311c5e17eeca6664938a664311fa6a2d8d143f55b
z6a6bc90d2d4030057da28c4336ee4a1de6b3e3a9403557d046938507579d357ff73bffa6cf4408
z5092aa55eb1d74b2326effdb7e6a05cb1c432e9620c50c4112b578f23b047d73a340d46339562a
zc9fa32711fcd6c7555798f35f50f71b3cc3b057625ec982039739ba0d0df765832e48eb40ee3e7
z4ec8fe9e658d79c6ad155b16f54df00c8a83150fd4a74d97db432ce4bda584f01a0d59c4bf4f82
zb0ef622411dc8690451d1e81e1e270694e2574dbf25faba07cf4869e576eb8186e6cca1ec3ff89
z4fe6566a07bf8e02f7c8e27a8489cceb4ff4b052754d0c756ef01552173f3e43000493c70bef29
zbdd117064b711872f20229a21ec67273631c0a824b7ac5047355e30314b2f79aac73886aacded6
z69a574da578a28d23159704555131f9c2fe29ad05ba149209340cd52b063c3219e51a8c4bdc764
zacc84df8d77dc03e8c96183e1aa47b403ebeb761a53adc4447b687fa9628e9a9392b2f40c6b58f
z347fca3b4018e6c6087cca1ad0d064233e052e2bb42555fb7290001b8aec439e99b08dfaba4343
zc12063b6d793ab74fb475065cef61594ca75c6bef925b15feb03a779134da72e7e4ab585cb740b
zca9dbb82c7c348a6204b99dc64346df2b12ef4533c590318abee20461a9376207fd0132ea7c6f6
zf8bdd807f89b0ba62d4ce1236aa326c50bcd100ff361b1484fd87d54764cbc88463790a134b4db
zb8e4b808ceca43ff96cd07f7d27ec76670354365ced3bd4ad4555e7dbcba1f05e4023510f86faf
z6effc458f296989ae499b6aacd47afa82ec1804e47ddd857d3e4a421ff3e06dc4d43c288938e4b
z600c036f4c40313be84bb1ce9329eca24fbe9bc19f9b9526c0722d316ed2df1da3526ad4c7135e
z9cb56b10791ef73ad368254767204c1561541b8660e8defd8a6e5780fce4281e5d4bad706c6ed3
zc60a239cf6848e10c04e4bd69cea1277cb7056f45fb452e695ba5ea1254b132aa34435916a828f
z4cf58cc8fb33be6929eb9116c7d63a24729c2b58c7b17c41fa69d29118a75a70ee4ae85e6b2a1c
zf60310d65c034411a851385ecb2296deb8443296bdea75c691f783199f4588989908b6126771d3
z0aca4a6f544f98f559f36f3c6a80da4b1883ad69b00d3c5b7d61b9e0e61300aec6095ad2ebfc72
z768f501750713033cdc6b9a199edee27011d090ef8bfa9a42c382b72e6ef7adc20bd1cf633cf50
zb40d17b043cb172e8ada9ea0aa71ab1cb32c7b7530b9e0949eb16a674f0a3052c069a3f8d9d0d4
z04b24e0c8dd7120c330538a3448dc58c4728a764c7b0f217ad8dbc1f6f4357259464e41ff2f6c2
z3a2e9b07c814ea4a487945443e03d54c9028f1a99eeaac2fdd333056668179eabe3250da18228e
zd332674cd762f2725a2117b66adf89ae9009bbc1cf078a1b64e2ad55a604a25792a81b0c882d41
z1a46c81f1b565f488010b0dc55217ad85e9e38e9ad46028daf7e56cbf514eb597b3906de596b2e
z1859febb9cdf457b0a5461bbde740e8a44c3c3acee431e0a46361fc853f2933dcd0f3dbe64efb5
z0eee1648dec009837205478780788ddf481623ff7d26bd0996cadbce26df4ec510f147f296bb51
z30c67009955cdb1f597f3f7c769237833cfe7dddf30af907629a5e44b783fdec37feb91419b5ae
zc61d921f0625353862fa66fcec24b68baf4152dbe3fe70f42fecb2aeabc5921651acb14300d21e
z459fbfdfff34df9dcf7df98ad9ea9a9e89c74b14ffd2dfa139d8ab97b6c56c01bb4f007a9ce379
zab62a4f3825d13cc876731b1169d596152b363f72f5e5dc551dcf4876da299ddc5fde4d38cc916
ze8aed6af35da74d4c112fbdaa8ddc052cf7014f281ae72f8ca4e0a8333f0d399d0411a8d301785
zbcbf08987b0b9c630de01e575c861d5b6ae13c3c0afa6b931796a122ae87ee0ee6aeb8e0c737c2
z04e6818b058e8f209846044f4ddaf49ed0b2b4f1054e20ef7bd9fa756cb1cca473cfa81fadf976
z3094ceee8229e21666a92df118b99217567362e3de99feac6a286f577da2a53a3b0452db218f09
zcf9a182776156bc7fb6460bb6e8b36420aa62b860112f22462d4ebe341ba232ffe11d7ad1c371f
zd5c8454bfded2f60b846492a5651bf9fdd3d10b39b9ad840ef6c5142ed280ba1132cd9552f679e
z81ca7cc5484479d7705cd038ca7c57b08b59488b5781f7829428e4a1b7eb7097e4b4d435ad1e68
z3f4eb0df33764a0636c21e0cf889f15d32954d143b2ae85b19d21ecf5642ae5c91841dd8b3f25b
zb5b9eff3fa6c7987ed50022d625b8519fd37fb6b4b72cecb77725fffc9cb128f0a4c9a8a2724c7
zb4efc5ff3961fb839d2de215028214bc2d9299d042d9386de0318ed75e51eed8756650dd72a9ac
z7c8571ea4ad74c2c1ffe51de2be18e731cc130e65532cdec65ec8a8896872c04a6b80d4c90c630
z04bbfbd2b4ffc558253ac35c0387da72a2657b8baa4c04255d1594f2d03a8f26f64ce7deaf45fc
z164a6340b645c93d46e898f3098b3087b1df50976561f86758b7eafcf69e471a985949f6ab972f
z9a982323889e4b5ac5c2872004074ff2fde9f01953327f98fd6a7f68a111b3f628a77ba81ab0be
zf23cd3daee823db795a61738b3f02e6a1c5fd7eef5ef856a1a8645e55b0d884ffbe048354838fd
zbdc30dbdc6ceca9297e13d4bd27a6b638eb7502544c3c446d77a0dce27146cd6bfd64c1610475c
z17e8c3eceaeef849654d34afd5f4eec20ffac620de9f86409ed9a969ca2f23ef60715be4ef4102
zf53d4cd80558c623726003ccdbd8b458e082a83baec1066f2965dd362e76eaaf3b581f992f4678
z2d1445183321339b2d7afd42004ac224482621ce1dd6fe13e09a1b059a4d0d31f03992b869edcc
zc2ceeb545b1daab4921a390216696f536d370767507de2acc3f75153b3b2c32241b0efd72a4759
z87f873f7d24352611bb06861c2e5935fb6972227b453d41750ed1926ecd98599ff076c51378546
z78a5eaa4d8a2c5fa534bfae0dc107223942a2dfde404ca4fa72d3694420808de9628eae8cd87fb
z9cfa63149853764827871fcad244d0fe579e67e03988d2d05529470d5685ecb96b851c3e364d7a
z6468a8a4412cd335204100567371166e2cb3f5fee05bd99f551f8edea86aec5b34e6c6c23a8128
zb00ce3f110072a9d9d9bd3dd678c20b60844eda87f6bc480b4ed8f834f1a19802bc8776311e145
zc660a089ceaf9426a25a19346c68507cc1d52aa4c301b8564ca174c02c35430016ea3e33c47e7f
zb607fe0145d7a58efafb432276528492c046fd39968d7fc0ca0b7c43ff6ebf8503158fc72fe9b3
za8f5ab9b91998e969385f907926bfd24e9e5d496fd43940aa2aa309b9cb34ab1ef862f2802cd8f
zd9769d30961986018fee5693618d114a623b816d05a4b44ce3c6eb63a81bf1fb776bceae02ecbf
z784994d9933269da8a7a312bddfd1aefadb1d3e4d8f8b43bed07392708e19d13bd5d89c900448d
za51a653376cff930a0a73076e03dbb020aec58721be66db006a1ec436634b93439552c7c2316ec
zadf96571cb00e3cf6dff6f290f6722a5dd6a2e8885b7c9d5532e4ecd95e585a3c76b62154f6633
z23cd9fdf453879c0c32a9c6dc085b977981220a96a90b35fb6ca0b8c8247d0b2dfb20768c08133
ze692c5d3a8dfa59029943c90a3f075b0941e2ffeb52034ece389260d45c58c0b22bb0dcb6e6560
z78777fd7a5ff9f8f534b1573e1ea4c635b17a5e68c4e6fee7e566f3f8b07090ef161ad739452e8
z2fdb7d9394808a5bb7aec93f0aaabdf87247f63d807d2a1f49e485ae89dcdbaaaaf81ce2307358
ze9b31dccdaf1a5cfc6463a53e6d4c698d895ad5294d345c3a4dbee3aeaceca7ac962ab20806c1d
za3c1177a23b4a1fd7a046a1ed77ca276c686384aef5367c94000c8e615352372b153250368e830
zcd4afa37e86b915491518078273dbc62166e81f12c8cb92b2737d58240217f15d0f9ebb678a673
z2a2a2b3fc3721ffa9749e45f28f22aae272da8db114fe21d4aaf10067862a450fac16971a23b9d
z2501c46cf56f2a52233c38a3bee056f0a01cdee5baa4b466d77d2dea834826e873c63834b26e77
z8d6467726be5511f5b2e39ef24ed65f84a9c86aa1221721d7eb00171c2b81936472e3eba89d9a4
z816c8cbea0d651265b16bc8650f133494a71d32192c32b1858043d2c2b50465e3c41f04c476941
za15d684d2716f678c8fd6975bf088126e4cd04d6fb7313b48129d6c2b915d0b2a7a85ff6890fd8
z581c5cc526d9591d7467783cd0054ccd2f0d6a744783e1d89ff31f3c74237cce80865c89ffbd19
z6725f5d360b21ba9557857dfa1441cab4d3683c16ae76e3e6832a8c86de1147df1db77d4616499
z270299fac9a66435b2dbb516b7f1f0a2cc9cf5841114d0df3dee43dc3ffe17c7706536d6c6fc95
z2b7e2f37035eb0a64d0955193418532df33d2f200b02b6e79fa24a995ff1ffda34a7c7b3784e16
zcc6e9280fbfaa69171b8a0690d7f786de19d01e69c152fe48cb5c567f9f8aec007da32054a3bef
z0990978cec9a074693a6e70864c5aec7d0287b3fb376b20f0a602f163e763cb5c3aac3fad701ed
zc4540aeb3379a8249d397ffcdc2fc40d5e47bc17808e52600583d4ce8ad7b3bf06583c9c394be3
zc7eb49d3e5840e87ec181a19012d3e4e2d18d0169fcb7987c18749899c75ecbfb15dbc2317c60f
zece87197b7994cfdfc90b96e91d74674923e4035a09652d4f5d7fd793013bed4253933eda64339
zec50e4731215162aa3e7405c196e2c55359e911c8647fcb7391676605327469fad9b34393f1cd2
z81fa725172695e8d26bf75674d622e8e30529da27ba8321d2a80605b3a9adb97f0fd339cfd080e
z2acf4b55e50f5ddabd4d3a79882aa9cb18bd382fcfda6a6bd5e7069906152ee8aa9f8461fb67b9
z52ed9f545a2d15d793ccdab7848460e124c71fd2cb22dfcc4ed7cc28b1fe17cfc3dcf9046da8f4
z8c28a76b2332fa92d6c51b97b368e8f30b6d1a2e672470c4547c88751a3d4f97b9abd1eaa9eaa1
z26de6b536e5b4ad4a8d5b7ff6d248eb146a2810ef4dc0a1507bfa402c26e3fc32cb85838774404
z42ae1910a6e0b77c006fc39fbba8a19297aeedcfb7d94568ab91ce7e719fef632dbe563a8c7a21
zda7292870acbcd598028b548f8f281543d1c46340ef8525e16ce7d8445a1f0f12dd11051acc738
z4cd2e3f40f3966934e0a4ae05193ebc0050fa16bd1e0adaa2120025fa82e793efb756d82969e42
zdff205daa337287c5eeb2ef9eb5d1642d13ff4abb9721a3dacf60aad3ebcc9f1f9a835c60ad9cd
z421ef1be454b7e98aad406e001824bb0966a3fb7893418cea1be01d30e15f1406cab5141b7969b
z100e86adabba3ede7f5b48a8ed4344663332fec094d3f7f26a746b739693bac87e64ff2f104a8c
z10052d3e8cc8e5a3946806776a3a3958e2e26aac1fa6519f3f360b5be0dfad49474407cb4aaef1
zb0e82f7a1621ff352a757578fa0da8fe0fcdc71a7c2b66e7b011e27ee9e0203bcd5a6895677284
z2e261b2bf808c976926a8d2d2969a73ef58bf02e1c582caed7bda664d774df9b8dbc4f82f0a8fb
z64b42478cde83e4008d5729dff44f96b1e2ec934809f5d5f1c9b2a6b4d497babe135a704364ab1
z7e222e6c1645941809a1dbecf85d38b0249d3e22690a1109c7ec6f305a2cce09f71dc1767e8629
z4f5fa3025f849837d05329107f91370c581e147d92713d2841296ddf8dc59cd70b34b223129334
z86eb370dfa8fa1f38a71740e287d2be49647501546ddd80feee75314a6c7529d98d1d62e4b9d12
zcf823aa84966819bad76893d5b261f1abdcbbf351e82e92896efb2eea82762a07fa0088dc8c3b4
z70e97e1d85ac221a6bda98be8a6da3e0b3bd5a4ac7268327eb5a8c4313b6dd828b9f46f2c98b26
ze9f3d0aa7c94cda8c0fe185ffff0270d52c74130d866acfd94f3d0ab2594be7dc04995b9e64cf9
z957a8d86bf42c53e12af4984426054fc0e263421140d35a71c90f0999c726efce8f71924bdcfba
zd0af5d105dcc53508e5518cac9f1df8ede92a3cde175f4b4b27d8d1fb272cfb8114e61ba7229b8
zae632b4cadba3c12c6c2b1eb8439105514a4a272ba62aa490f4c4f2d7f7736a7c07ffd80b99930
z34c6296953ec2edbb5f5e199390f2e1f33d89efad160cd3fda42bf460a20e973243bc174a4a02b
z64fa59f89e22180ec02027ac397ea0bf3494f4125551c555db9f181a193958c95b0d55fa321280
z5bff8886938845e889796cbcae2b53d02c565cda21959d4bffc203aef7c92cd85286780d8f0878
z64ab0296cd3907f3aa7b365201b78ca0d0ee55a0bd162556a530efceb8901f2a4d1911c501dcd2
z96c0dbb34dafc12d0eada40cd04ff85b3a22c720ecd8e628bc64b56928d77b38de68db4d508075
z5b53cec32d1ba881d787e896abcdc306cff97460f1498c640fc836201428c73507e79dd61c0709
z9fe6935dab5c70c87600f32e653079683b2e696e1cf8638cc6d278322b5f57a1004fd2eeec8905
z1daa1ca0a280f74b8fdd0a5f413e8cdef1e7f0f74c4582372c9cc3ea744411c01d0d7580ec8448
z989186cc4b88def7a1312ff3df81a8c0839505bcea477aabfc223fd429b849a980b8ffa6993127
zde55d3852fda9e5bc38b72252ab45324679e510af1cbedb4c136dc842cd3cc236244679b253c3c
z9c524c6dd7870ccecc39faf04521ace214f5726dc43187ddfbfd8ac0743834accb71c731f30d63
zcb2cd83fb37943313285249a84de16f74a3c121b455277941a308a8de90015e788378e1c1edb37
z12b2afcac67f2f9cb06bc021a65ba093464b4c754d52f3f5c7398fda887580b3032383e0f60d04
z0936e461f3362d250c557f22b6a54584699002e1c5c575508575e8561418dfc4f3a0237cfc71a3
z5877d31a517a75a772f209e6cf28916f1b88c0617899cde75957d05762088bd4d9c5182e03b712
zfd72507ce661506e1df5300ab395d51694c74cb1ad0b1d0117ed4b92e44cc74918405601d2d3dc
z09e296e1f84367c1f87eded11f0f390e15ea66bedf4cee16ded4b834a0c2775a88a1aa3662c215
z36400bdee7506ae1326e6da90799672195df2bf49a29a4d83bb70e9390c4cc749967fefaa8a08e
zcb387e961c9158430c4d180b8dff582c240805504088ec8d7d8375c1669bbe461f01ba2edf9283
zc223bd311079c4fa9d8d458866aea37291158e8973a26bba0a093fc53efd5160c946a1f19c4653
z2fbaf2d6169f6c04a92fd4ca0ce8b224e5756ce98990384f41d5e9e69b4efb930087d74487d0b6
z16feb55a546fa8e8c8ef9d08b2a54e6836e85f48c8d4d5a650b877edbee9999e48a194563ecb11
z8047fcc0338e04602c05d9791197b618e7d9ad96b1ae4d2918605f2a8e5ec1b9e08a9e6cbd4b95
z7a6f48ddbec54c5c012dd667d780308d777b624504942a110235319c1e241f92e1e8fa5e1bd6cc
z418c09cd568d0b6b79f6251377ecf177e843a6777ae19a8f058d65007e00a68f21b3c68ab79e93
z9ee6abeccc1096024e37e5bb2e1848d0079a2e6d1a2ad1c5a2638b622d41d31eadf6b96bb63a5b
zc27174f49731c14338e75c47cf37a50a5ab88e270811a2426067425afafc77ac0aa3e52c993464
zd4ca7cd118ef084004bff3bc02717c874df2641c1a9bccecb2c6634dc34ad65b7a096e2745c0f7
zc5971c1a62bc425946dedfada3d1b2c864ce4a49648270ac056376933280a6867dc294340f7784
z28d710387e52043fb655ed70ddefbd416919f4a6663fbbbc4dc9a35b53fd8c2ec7892467fa43ac
z7b2ead90fbdf406885c68a28eb330456628c2b7a4fd8e0f2d9583010bb5499998b39af6917b638
z13caa54acf08b9250c44eab539c6d29aacb9ae4aeb50894c3a4e2c22702ce8081f324393ae907d
z7013d7607b04dc305c234e11f741f5bb87931a2da9d391ad27e915af41ffa23d211d1c34d8cc08
z4913252cd1fefd76da449ab81984df2efdeb57a6287cca195688704714faae5b8865af4f3a0478
z9fd67dfefc90be555a3bc103be15f49ac345adbc26abcb5f96a9188776fadeabe34c999e2f97bb
z6b7aaa8ae34b45f5751f7d894f9feeebd32dd53602100922533c5c02bedc2ef2b31f12ec8a9709
z4a99560b7d49446efff995f4006a91f3c85eb0313c2ca99911637e58326967574eec0ab3b89069
z128582048d242df70053bcc36e2a26fb32103416a7ec6c0c77015e72d7e49cedee78c7993492c2
z193b27d6721eaf6c746befebaf84301b31d07c4dd0968520984606d73812537b28f2049b549216
z75d5534456020a0afd6fed2d205fcb87a113625ed28e6729b4878ac982aaf09d251f0768921002
z9caf4f43fff2de226af6fbaf2296cbdaf7ce2cf6d708d98b4a3ec2ad285c379d814b4c6d816965
z018ab7952853f47ed856cbbeeceb091597393c2b6fe1373a58dd291b6dce593dec35fce09fd516
z331443cffd1574460ea00fc67096d530d70cc89c637f6c676e735c6807b29b2de30ae8b9ff3ddf
z686041fd1c424f1d3e68ce9737088fe35acc7a5cfa43021e6e165374f9dc11ec00ede53bd2def7
zbe4ca48f933a0a294bdf1d8dd81c356ae8108d3f73b69c39edb942f355a2d9dea9afe79f0265d2
z0f04371278a4347b7e6a75e3c3d2c12dd0f6444e8d72119dcfbf98fce8f733e7e754f6a74c5fc5
zf10f27f6c21cafb2dd94c96c399e98a58264c1e5c88ae5652fae31d1e012e241701c371be8da39
z2f868611f48aa3c334212bae22075a7d09eaaec90ae4ac1f42e98c3efaaa7ec2e66202bd275b86
zd3e7e52dee44285dcd3e383b1fa0bb8c2697dd910c931d26562075b23fe932437e5e94a25f2b2b
zba9fda2ac390453ab33738985183db2fec30a1de9784d13bfc18a2afbd330005bf62fcfbdeb502
z57df0dc3423f401b0d8482394d7d6096d782fdb30cbb65874b54b2ba1ca5f38d44fc05d0a5e392
z15085b5c178eb3595f316d65227961b2c8209f4339b51d9433e6937d89f5d64bb0c9138fa133d5
z7036283393d5477082e0a3849b9e4857df5d0cad564c02c5e04bd850919d0463efb0d00754366c
zd7fef91a424d01abd7721fb8683283d614a96388b6ce19d5b8eb7f6e2b705e32cd20d992ab429f
z6c8c8e1dbc9e3b88066b6033fc8085bf7ac6e923db2a92b1b1804223063692e02f1261450ac27f
z1b8419cddac29567c83791589502c75edd9d92be5d47704cb933d9d04604c0d01f70123515dbdf
z0b55a6ffee58ec002e7d1ade89b7c420e7c69672d66bbf267ff4cac3521786f1342edb1ecbc9c0
z367dfb15d1daf22425ade826a302534add1ab920ce19360cbe2eecca87ab8a079349a164c8e2fc
z840313a6b7f7c0256b6f9013fe77c4a05253cb71f7709428c6b301840cd6cb6f4388d6efdc2293
z371d721dab48d5fd4d7f467f9129e85f539822270402a3560c8538b9d8a8340f2d283a8b426108
z81f11c22ee97416341a1a786c5c0a5683995ab6ea4b8527a28b7f90f6af2e654264f3d7db06d95
z4b3d6354dd3d4e994884aadd484d93a32e55e1680b0b12eb9da87f8920658690a736664df26df5
zcaa7c76481c6e4f26f980f1fa731ce9305128d50a4d8b87dce891bc67e5b9ffce7699e53cb9347
zdc1a18f463affe226bbb1949c63ea6de46078ea86c665586da5514fbb7ac83e17734036a16edfc
zab470157291f062a21267cd8e4efe0b7cd131b3e6eae0cff867bedd3cb963981ebdfb53d9acb22
zdc452a8435ffc9983c8c97b6314a5fe9c9484703900b683449338d185c38e2e5b1876dcb968494
z7ea7e86cf9d1eeacbb74480d4dca6ba27df359965676ba1772bada468cb7cc05f535e4d5614ecb
zd81ecb965504896190bbebfdeb4811ec2bc38cce3267cf7518de86a96e2e06e74ab378e9e2ae3c
z1a1a0d41adbecacb073dbf696afdf85bbee45e187581c14ae927a48e4573edb73d984138d1f2da
z60f26bbcc2fef36e29e84132128862ff902050e55b56f02127f1ccb7e453d2444d3ff4782ce780
z90875dee731044d8f0fc37fc950516b21bdf95a2188e0e2bd839d3bb62e6f13cebcfbdb2379e85
z35fb1a07a999551088548ec06412c383d0386660e85727fb805e018632d3718cd430aaa7586c7c
zcc84425429877cb96f6c2c1eefd845d13729bf98e2b8cd06b6cc3e29afe93399bba7607f13682e
zf7b0e59ba8c5e94178ab3471584fc6fe5d015bf7305f3ad7eef1ecd830c76936a01dd23977c13d
zc3894fed444d45a5ae42edc4baf9f9e44007164cb208492c0d44998f9aef62c8ab0c9678aa0d74
z9b12634791af2dd9c818065a96893530957b4e7c34a307a972691556f10f1f54ff81ebecb5167a
za6af4fe86d1e64a0048a4cf878ff9441359578823dde830d8fb7bc9b628851d9808e32b1d7d4dc
zef1833debd3da793461721d4f598ce7c0e17d93da8c98cc88268547393828a55c7ec958e666e75
zc0a70bd487ed2690428c05ed036d0695ad5e1ed8e74a9f540acedc0686adc2e2943abcfcaf82fd
z5de3607ed717f1ea72a650541d6a408cb54415112567f063d1b542fa8505786606b964cd740c45
zbed82154897c076266f23cb351023137ffa48c865f9f731aafc46ab163b4a1b28733b5eb0ea91c
z31ab27cd6a48af742815ce39c2cf8b5a4a5224156d027f516a9f4f38fe7cec3bed497323e90536
z5d6cc5ee1e1acb3d8a97e34f733318e09765217735d49cbeebab930845162bd1b0316095dcfc6a
z470a11f46c81caf0495f9111f2fa11a510f17141915fa83809cd8b956234f487e303db9fbd17eb
z67ec8d1b49eed99b545d59e896b74b2761daf78d252107b366068012a87e1ba9fe7b387eeff76e
z6334bb59ae3ea8e8ee4ec8dc74fa1ba21b779dc46cbacc8b598bf765c43d1509c20318b6644400
z1757c1108133cbac88245f66e59a20e1257d2809ef8fcc0d9b1331985a88cd9f1be2ece7e20e70
zcde7c6d553bc5bb55bc0ae40e3668d2eacbeb60595e75b2137e89716aedf254a6f29fb9a19cbb1
z7f49ffd8a5a4e172532e0f95d2a6cefd5e57855c8f928131c04100851a951d875672cb5b314d3d
zf5890dcd52aed7c2f3d683e6f22a8f1ab8a8686f4faf98106eee19fd232402bcbeaa8f947f6620
zcce7e41e5f3e7223dbceda967360a852e6d7e8a84b1235f132908d79ec87fbae4f3926ee1b25b0
zbeec4ae934f7f34a6a809f86088b15379cbb44e457b208c8f62cf09590e115c5f892090877a52a
zc4f5c7cd2c2345038c13031e8baa1cbdf36362845b1e5cfe25cb2239205d301e3b6a81aa962726
z505c3d825bbf925d255d9b45c1e00b9bb56e672da9fe7eed213b046854fb6ca6a4cf41ed62fdee
ze5265de0e75651f284f1ffcb3fa60b5dd0e0c22cd94bf8479a580574d1dd9d83796c3533c3a8b4
z2c4326f77313fa2b48e90da0bdbb6664ffeb22762ab1dc2aaf066810f81ed80fbeb46d3755f60d
ze0bd038176b2d41e3a32ad6c0bc42511a3f2a1fb882cc52137ef2ea049967d6ec32c295572cc6c
z57b1e62fcb2134b8f2b2ea82705c153017c808ff70374c307bdad11e396c5d02c76ca67849667a
zead84e857c9dca8e37bf262e6e26a776fb5d5080d0ae9dbb96e38b2517cf9aeab8ad54fb27478f
z458625ee15599b27b5040986e255432567effd06c6ba5c7f9e1375c67b075a0d0898c81acee72f
z0e1ae209d4e73dbdab8f81174898e8044390ba720053c3970eed8eeca8ca73bff1a305d54962b1
zb38b7a6f4319ed8bf7cfeb09e0fc721be4a20b77557c915ee44b8d3fe0c06069a79661cc8edad6
zba762a84d4bf4794394d124af74a9e1618d993a88bdbcc42d404cf0b01a8211a6153f86f492fa7
zc41fc85e1edb5685065ab89f92287dc9e06ff0d6fc5bf927c0343f55cb42d8971ac43c83a797e0
z4840b4580c4e2b3c63c696669d90f3120d8d3a35d4b81f9eb3c0460372c3c3f00f9cc813ec7122
z9fea7f7e58c1676f47c2441b979bbc89c5134b7de66d43f6faa74524ecd69b32ae4531e09315d0
z19943c0230f12cff46426ff17f6ca8832f5805197b351d2395216217b3ac4e7662d2829fef83f2
z08c19d850d453e3e37a86f6d3bdeb5b92d0964ea7991aaf0b7ee40cb1e409ff0de34fbe8811df4
zdbf8aa0a06a10c66837e36c024c2fcae81ddaad3158fdc2c914fb83cc2cb765c82b5ac4137af5c
z34f9aa5f61ae4bf5e4c9fa8a19d84dd3b17b6ebd29dc2ddb98a8541bb0fc228dbe25b672e71e10
zb609bedec4a967f06c7c296032c949031e8024429dca441108e872ede8a63d85e94a5d40435abe
z8a54c26a3863b67087c428529b5fb132c17c160ace056f17256fab9d831757cc5991e7ac3cf62e
zceeec56712f0ae6a5aaabeba48aa01d23bd680f0b2d7208dcd884387ff98451da62c8758ff2965
za2e37abe61df8cf6686f3225c9511658b4210ec3a3227a7414a01818b40288205d9fdb7f3eee93
z754788c7aba79d5f6dc646341078ca35d7e5410bd1f30bfddf1ad2299f2462e852b6519e58b1c9
zf42f2d035b8ab3c19c68659f3b4ef0e1121e68c371a76de3c51c03b98c0124bc6849e0eee8f660
z6e70f8618c9e2ea01789b5faa40de6b2eb24a738215bb6488fe658a5d3ebf958b6f9fb04aa0c28
z816ba0af7fcec37621bc1b6db51d8f7f0b3bac12bd9a7e5581366ef2c37e277ea6ede7e89fc7da
z8775009e521aec1d9e2ffd7d45d51b6963e5dc17b2cba9116309f904601078f7c052a1d19e115e
zfd5c6436664773f37d980e0259eff412339917a416d187211756c318feefbff8596198b6de3058
z501b8037eab249953134be205dc014691d4442ac82a5bf8163e389265d6f3b90aced0569cc0c2f
z373ed691f25883d5e8aae9029aa70592408ff09b4023d85af6d0cd4d528897ebd156a939602415
zd73e20bc37891e2af304c6ef36c80660cd601de99c76f51b709ed5d414e7807040edcd56b6edb3
zd2e534ce8071adde1da7565a2411c5e9f94b78a13235d40041cd968fb3fdfab325c7e2dfaeb3a0
z33d06653ad50b2fb66a81ffdedca8a9777b3fe1420f77a59e6cb9ccbb0ac140c22d3f28b11c728
zf2f8fad9131c7105301c1315657ddf914e1deedc9594339dde7f98aa77aa66c0a92843779ea82b
z0c0d5f3fb1d8dd16db936d50f3b56f51e4220fd0e5bfe5dc4f29032eb38d17d5431e26b3f208c2
z0a04af245b10db391a12c19c6f1bf4930539c2cc14f4733a57c2d956033eeb8d4df29312dc19fb
z5ff4470ba930d131d43e092879a1ad7a8ff7dd74f132b0b48e5bfc28eb42be77fc22a34ebd16a1
z00e39d6f0ba176d444844739cc93afaf74122141f6de81fad564894128e9e72448f253bfdb6b6e
z31109ac7f43dc5223a9da69fe18d93a6bc96e0fe53639d0c5e513af4f248de074391fc279bbc2c
z2b57eb5fab699b4e29c40c2a0aad00e3667f6051456a94e88cb084d21925b9eb89c1ab7b6c85c6
zb628342f05914eaee46a8239da5e3772cb232e35b8fd36ea2361f5f9d4618c37fce2bcd58a42f5
zee1bebcce1d6cb9f7a30b168c81ae2f96e82a409bb0a0fafbfaed637204f8388e9501b72b7b13b
z0b0b039602fe4f080e741ba7fd741b5904c6c58e9c4a5ae15318a2698cc9f916dd3595f3be2227
z256d8663c9ed51c501836de25dcf0ad18537478e99e38fd0f535a2182cfa52c4e176a647b23a8f
z1e4916cb0edb5a5b5d7815c12927f5f3dbc549654db7feb99b044d9bed0de1af4113cdae50ac8e
zd77a426ab810842bbb261667936a4cd5f70863dd81bf79af30cc3106f6cadd8c8b50ed1b563e48
z700026cee948d4ad49f25744c3af393bd3e9cb01edc2ba4d8bcde485386844fa6fbbbd05025157
z1e42a3b3589d67fc369d56a14311f7bd8736dad63bc5d7e9e688b753b7e86bee9c0d9f63a5da87
z3b3a3b54cba4b59774d1bacf755d483f1f7b1b72b0e3439410cb367e21a817d62a0d69de41a622
z92ede19b7b1a5d5dcea900e253f1b333098e68ef7ffafe7ec204229a7dafd485096302fe8a9d64
zdbdbc8cb46cf58d2b62e626865e054dd44b32fc7165a80d5be35f27322527f83b73a0e46234d49
zc11fbe594f2c24a00ef0fcc8d265d66c7b6f3335bc322df638cb1abea492042acac431cb695ea8
ze459710928db62f1a21265c97f05ad346243a4f87f7d8ecd113bd916bf68dc23537394ead386ea
z5dee350a85e03c2cf52066946124a32ca52dca1cf180a321c22ea798e8164f03e30875bc7a2399
z4c2561809253a58431bee31b60ed3ba40aa36324255e8d461a4f7f6cacfd21656f06e0a6ff5acf
z2df60bda4c3b6d4d3de63fc173bc4eab3d342742976a310062127a919b3d6f320a2b50ef78af1d
z150387e92acc82090816453e009b8602d6eabef3aad5fca6bc827f50536b9b7da1d262bbe0e5d3
z783dac8825193f57059cb2b182f560080601830e226b58060a4acdc131b3ae4f488460611fcb7c
za35a8f06ecdc25add09834177cddcda6bdba8b2d1c5dba74df308ad4fb003fef30da7c0f95f555
z58ec69f5daf593b6575ab39db8af61ddd6ad367d72a993b12e1619c8103750c6d92f91e96a56b7
z65175ecb44fdf153bd781e0a6d7c40662750ff6c16eda8245c32491a9c62e68ff8f3289e467abc
z0ea2eb5e79cadb969e696b73b57d33a847bddedd5fb8ffcf0fe092fefb1e8657a3e5a0ae43c538
z4a025a1ff2afe4c4e06e735d4657034f8db944af3e6cb5b997a399ff31649658718297c799acee
z5f29f1de72f9b78f0025e781fb86cec4225e7bf2e667655caae389cab9bf15b82ca54add51056f
zea118065693e2c91b4c0ff04243c7ebb9f6a365eb94e13139fad1e5eb018c71978ba393f715e83
z4090de8954ec065c21f4522ce0cbf6cbfe22b42692f3e7ec8260d42461f204069d57acb0f3fee1
zef92dce60620ba97a9fdfe82405922ff694bf5cdf4897e4045b39dc2a6145383bdf2f9f10abcaf
z773040fa67d8b2dc65381771b099ecf92a80368720a0e58557fe5eb41d7eef6a8230d57f3262c7
z8e2cd54723aa7073d3edada215d70c887b788404683e3dfe4d221828a9e11a37e7e07d870ef468
zb7773e61fefbd2b1e4d25268734a66b5d5ed5ad5fe358f9919424422732b7f64c5699a03b727fd
z50f89075336a9fd537234005ee0a5c6b9b546f85ba687d594666af40007673911e19ca1ad50eaa
z23e1686a89ded82fc5284f3a382097499424ee02b990f8921c50c95b15c71e69d1c2f39525b0ba
ze2a83a4bee31b7d93654010a67e5bade760cbabb8e14d082e05ad3faad1d6c8bab9d39befa0c00
zfab8464649e54b122a6c57f71f40faf7142183780af4f977e498ad552da7eeaca47f4d02f9d3c8
z929873e31cdf190d5d8b8c5996ab46d908af17cb6c45420ff07ee7966dab80a3706b4a6c10ea5c
z2f74f2d3f6b7857f0fbd94ece08c4523d78d28a9eb5d28fd181a812a334a343a6f5bdd57a779b2
z5c6e8e215bf5d7bbe74646de3945c3bd830e493c1447dfeb7cb37ddc4406735bb23efae4e76561
z898cc98520e3de7dd300ad07e574e94c34a8dff63d6b2c295cf6f5285b4b0d235f0c90de6ce232
zae78802b19d030c8470a51ac898561602c3e1044890c4834479d18ce970e87c40f3e7b6a84bd78
zb5b80bf148fa99fb8c3205540b9680948ca0898fa9f53d0feb46cd2cf5ca8e4ffb8a81cff25a49
z16e7c45c36f8fda9684f2d62ca8af7243c41ccc2b44e63d86d365d0d611b163016a173b95889ea
z71933030ebdf4bf1c57995aaad0f926a11e97cdf9b5da1142fc6ebaf95013af282a89d4b4b2100
zfec24c9d7b193ef4cfd2002cd072040168b94ac5b76aac337492b662f1b6dca9ec57b6f2e6f81b
z35e07caf6e549c823cf9d62fce75a7c24718d5b50babf6b4c8c9d541da65741eb02cf349992dc5
z7e04c7a97d2d404f1bb9215224970e9268355cb5472f634a35732b2ad5c40fd018ce586f174b9e
z31a124e957c38c21c6fccd3067b25316db3c11367e7c3d2e9e1d09c41f34f139e2f0da2149c5bc
zbed22d37978e88267422d02728577edf2715697cf5044049efd9766721ff4d5fd64f4a0bb2ee38
z4e667f6f220b98e0a2a43e7d424715f2912c2b6baed8138ab5b85d9902a573c9b690cef881de2e
z81944041c8671ff7751e09302de98a0755ca530c75769e0501b43d99f5237786fc3bc357338f23
zbe60a2e11e0348387b12e20f2f955fa15bbc599855cfaac057f92f659258e139ac0f98cb1c4ec6
z4f6d6297df85b0aa4e1c520fe59fd0f291fc6bb9ee415940c703e8a9db092f0c5e6fdb4409aa97
zc9b1c6bfd77132df9f6bad12c588b8a0adc2ddb9530dde82eeaf58b45e6530c7c49e9f1c1a2857
zf5478525a81d5aec2876159089b6a224299087d0bcac77597539ae30154a3415c78ae9129d22a6
z9c609c05e9722b8cbe5b7f83a09c43348bd4984194b0ff1ad0e8afee141887d4fb13bffcf8e2a0
zf63078b1409a3e29c4de25fc129dbfe5d12e3ca0316365425bb062eb1abad30e5748553361cf2b
z3b46fe19bbdb576c048f6e85c30ba05293c9fcf44a7860a0227dddc9e1b9fc569defc0ce97cec1
z0f6ca6135b19477933d5a1f5e1a958e3c14785edbd9e4048157468f28b11d2729863ce3953721a
zc9fdefa451d339793eb5eaaca01f58f4594425fa8de4022657e824820b36963d04ce69d16a8d56
z8546124aff12cea68090621978fc8f6617ae822e5da1f78230566edf23c9624b3f7d2f54e09e8e
z9ac550f0d396798fd11ca5a3993df840958150a74985be988d55fe0971a8d934fda4134c6b6436
zde728efc4630f4386f3845c8690c8e43523f3d758f0d9b1c21af5a1733ba7d528a6806e6b020ed
z176a2193be1af5a2656deacf8151cca3d72eefa39c00ccf531b5a3cc0d8e2fd1d4394ce5161f2f
z940ced47b363d480699111d30dfe0baa40252dceda46d4d7099873dec360034a8dfc59fe173951
zbeaa0bc7fb76cfc354ba71f5d03b0e147f2e50f5f336170f951e6e21a03c4050fe89f2be911bf7
z9dc5313b464cbd73b62850e5699a519829913dff500de23037bd81f9d0d32cae7c3a8a74cb1d74
z677a7431433de6ae3835b99ef11cf91d259dca366f4df7a50c9219c2f76496171cb9ad30b53edd
z156b39896282f7afc0ef89e181a49e764bc00607cef34d7f1a40e0d8c070b24821b9d9879ff0bb
z403b085110a3e9e118145ff0ab9f379bf1f94774f6bdd220427b7587118ea5333e2c1d1d968952
z6c1642e2a74e5de8cd0f8105e356fd9599320632feda462be405bef455447bb740d5ad83a45f34
zd36cd74a15b4907ba718a2e254e424e0d57633412109112abb4e72202e79a0c5a6bb49bda11360
z18571cb9f928176d90976a7479d7776969ba39cac815e653cc4ec5b16fb54c3679ec8bf3e37a37
z08dbe86672c5f6efbcdda5772ef1be6340e1f63f97164cf144803eb5ed6c86424ffb817bfd1829
z41fc0379c026637105acab53deee5f5be7cd809f7486b47e690501eb41a334230dab370fef01be
z5554a8772c12487d4faf000dbf9fed3c450be1595cbf28d92d3ebb22c4ca2d524ad50d34d6887d
z11775206d80467c9c36d9d2135d21f401d85b7f825fc42eaed4420c4bf201adca0d4156b883863
z59a95cd0cd9adc0be64e9ac917cf9ad844b6834eca0c1c53b763040ed178b10ef19c4cd2241c50
zaba0e6fc4986deaf75d663aa5cd0edae94ec3c2ba2505e4cdcd98f13c38110374cb47b22f5f8cf
zb72b62768c894eb5e1c2e0a578952b3065e2a70882309373b0443b2513b6207f0d4738d89688e2
z13e2c3219d76bf0bb7a749451e4b849fa3dc27508e0152398d45912672a2899f6a43fe91f652fd
z4fe5fb01954e7db391f62208bef826a42b037a43fa62440f2bc3b5c99fe4ee18be904e23e9f10c
z3ef589248af3406739841686ffb8a1ad1bbd9936619bf1cf914d463032f7a487891a1392a22944
ze47922f71cb2c65bd4a53fd48b66e6ebefd7f495be5df279af0842bb1a48f3da75cbb67cafaf09
z2db80cdbf6831e7067ca01294335c0a6f425117e29e233c51d55f7c701264d0fa5cb4470d170bf
z36bb871e
`end_protected_0in
`else
`ifdef MODEL_TECH
`include "qvl_lpc_logic.mti.svp"
`endif // MODEL_TECH
`endif // encrypted_0in
