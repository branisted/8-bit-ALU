`ifdef encrypted_0in
`protected_0in
ze74c34e226135848fe16db9ffd31815111b6d7fb642c521a3f628cf6da949865580b22efd062a7
ze90adae0e65e66a2c36a587d0a790699161455169ed55a01f2084f11770a774ec4c588039b380f
z6de9c5084882a40b79a175f5c2114b2b6d78b070cb806e1c0aa9258297f4687ab308bc470f0040
zb0b1de382961eeeaf2e279e1462520fc31c119af8f2b214846f56c2b3cd2eadbe4099496abff18
z15cec83ec4a77b868344aa20ba7360908f5c0de2a79abf8b3534b883bb12180f68b5d4beb444cf
z3fba8f13afb0abfe8fcc4294810f75afe452434d2d0f1166236c82f76edf1e12979f04bc35693e
z32ae028996dd85737a8f5adc1ebb94f39c940246e887647b64782cd7ab429b0544c173176cede7
z01dfb26b1f73408344a52b7e1f117f12bb9c8077b34876c2e6fdc085981637012dc9754765e1a9
zc512ce062e0b8fb16a214591f5c81e1353b900a611fe1f4886b57940b41b7f2ce99a7b84b04b90
z916f717e73bd10589c81e207ed77ec660a8cbed5b487fa50acde1b055c8870bd8676023f21ddcf
z9c98cc47cfa2d654ff1365d1f45035a045a66c5dfa82790502623b57a3af03bf0f0c0d35b51558
zb8b5f2d29acf03737a9ca2a053b7a8f06800d50b465c41b30eb585f62f3d0c2c5a43bc3904db24
zc5b00403728d562fcce00b0c730547daeef59c218114a3913acea226708dea665d2e9758f03559
z97123e13813eafa16b03e0b48be3dbf74bbb91f056fb1f204f4bd836417d735769a98952c6a322
z1adbe2f827224fff25030d8b004f4d66cd871b76d4aa4d46f7de2cf2a22174412ac5aa94bc2374
ze88e33f3d76eaf46f8a8b0c87b981745d7639e697d92db7593091aae53c9c7bc9922271652bd7f
zf9985f2ff4d8f1652ce9e2a6813fe94247cafe1e3a4eebce975106c64b8d53beda58d020e94b65
zeab0e49056a1f411d9dc7e488cfbf7ec55a0fec8a1b804330ac939070ef575f2755beff660bdfb
z0d91dc74397b5ead1cd7bf564c422095147a5172a34762a5bedd70cb938c2fa73ebf83d150bd0c
za6c31db5993f290177c81c736931d4f19a51b11f0b30167498a0a5f6cd7cec7f7e5360365a2651
zb9e34d7c52779021dbafec3eceb4105c2adb199337796a06b53959d6b5683d915eb2389c185db8
zcc94b359271f32f7198737351062728d13e1f8713238e83eb4e00f029f51073d86ebdf779e035b
z256c49e92c1e58cddd3c6f6305a24d5dff1110f67a845085bf550cc02083d5702dcf216274cb9f
zc61044e8bfe11b0248052d1dcab3f3a056fd95c28cc3c5b2b4f7a60cde4750b8ea0a4a808b80ec
zeabe61923307a001478d163f158729bd1542ef56c294aa89c79464a5f45376bcca812b4a163aea
z81ad0638c11f1347ee2b61ee28ed03357776df80cd60bbeb83af06eb4790a9494777084a6a899f
z8b2713e2dbf680df482461df38d195522277b610f5ecc4f068f45bd6c31e9e1b77b8635def391f
zdd3f479ee56cbc2a90af2ac39f646e03af8c237d4554a13112837832f352fa456df2836f10b7f0
z5c01b8cfc32e443c52d17ba942a05c53709b947ba5da76f3eb3dbd8188fee9b139af4bbc2a05ce
z48dd270c383559b2c4f5effafb7db6cedd47f7b1152394c6039818c91765b75a5c234eb3b14dbd
zc6f7a8c3ad97cd54e94c623be09aaa837c61474341c77a5802540bc5ab09aff71b31c48d3b1fad
zd90fcc9a197ca8097be8bddc490942251bc0941f60e997a124047e6cd676cf65d97ee70b44a068
z09242ee397114b8db2a4aac5bbcb001e5550592bc87f045cb9167959271d6af892c6610ec3cfdb
z70bbfbab4200d06f8e8f029e87471b17fee448a98d796a1d45cf907a78663009b1380bc189d0eb
zc5fa4ee014ce3a0d71e5a29a3ea0e6e3e6ff04696be79d3d2c50fc4655aa88e3b2d1b0642a1cf2
z126d39a22ac2fd3025b630b15ae94cc339a6de6554863644588fbec8e6e3b1ea696d798306f861
z42568f318c9f6fcf7251ce98f35aa9ee873aa68e99a4abeaa2321f796bb0ada53aebaea5ea98ee
zce97248f557a5ac352ca8ddea60ee68792596b4688fd6b007fddfc7c1f4d62ace6f033805a8d35
zd55a5aef64d9db0c34b58478f019020c317b690e7d0f6d424741e9cae9714552e247cc6d232d2e
z735ec4f861d9e6e9deb14f3fe4dd1aceb59650f8d6affb2ed37a7ab8fdbc832bffc0692bc0704f
z4e82cf692255571a92793800f9bf1fb80fc06ef6b51b50fbc18bf6ca7f6feb7c519bb4c0ec0f69
zf10e9aa5035290f5ae587768ff65df74551a4aa6c70e2f9a05b42a54e12845e8f8b7e90bf5c774
z390b8fa25a390116c43f9d21193c59c0b6e0f6df080d5dc56a3db7e837ced17d700f0846eb2b86
z55be6818b0af09b64124c3830ca6252134066dd8d7730d2607e5941c6823c3c56dea35c45a3d1d
z7d33c387e899e75a94682eb8ca4d68bc8f71e200c209036db58a4960a4f788d21b924faab37d9c
zefd79250b4e2012b648d6aef32ea638da4be5295303f7312eee611f87ead728760b25a0172b81b
zc801c53b03c1b81030fc7adf6b17833b4a52ba783424a490c55a5f97478e87c85270233f154226
z4894e908382e3f638d2281522899fcd48eae9ce074d5b487421fbfdee5d7da7c9436db35d9aaa9
zce29b0c33d31d144324ac3f58dfa625e2ef9cff3bd0aa0d6ebfd258777e6dcb65fab49b3a522d6
zfdb81f714c2733e94397c0879cce826f7654921be53c14e167f8c80f532dfa3c5d04713621ba3c
z5ef8b7f92fb142c23e51ae977ca342d51c5b4577883338856034eb225b1cb3a83543b209ed8591
z05a4a27bb15ab633269aae5d272334ac56e08907d150666a156c7c453cac6417c57f6d394c44b5
za66611b17882d9fc8909ad3673d212751e28ad2595e052bc9283b206a9e9f004c1cb1b2e8e7ee8
z4749bb2bdce12fe58ef3d166645dc72629c1da08fc12109b84469e0e6d7621ad382113109e7288
zf584e757d962c598d2006061c909f025768227fb5bd85aadebb47845f5fe11af731c8effe0b5b9
z8e0cbb9bcc4a5da44f838762a2cc73caa1634117e5999ce190133719072e8085e3499ee438cc40
z739780c608aa39078ee160377edb42a512c8fb50904e64dd720f0c6dbdbccfe9f44b7408cea4fa
ze370925f804cccead6331cc9a5a62c7bea77f858ff0820a335430087e8e0637236e608e9da216a
z1f5a324a3ef93d83464a0f23ccdafbdb84fcf561ad48d6c4455b18800aeda661711ce27c7df34d
zd824d415f1ac7c6adbc5962a2bbd3459a2d4005f8a86ee5b46e39d1f4279908b6310b48bdbcc66
zfd8e5858d2115b4b10400d40fb4256b96b3bcfcf0eb40625fe9c3a566243b767912194c39a753d
z18345c305e77a8e60d35152ae692765f733db094ee47ed1b17ed9ca922d7d1615856fedf1a28af
z1428ccd48d32d12fbc1cacb9745b5d54264d2ee66d8667cef0fbd6f0fbd55224c2abcb8b00c0d6
z72ba8f3373d1bd3b0d42890e4717dda01e685973c142787402c25ce88dfe7b83c11e54308472a6
z66c063f29c1ce901a78ef061d9ef77b2cafb4f224d82f39bc416a12a9366e2be4c04a77d3ce163
z9c0fbb292d8db829e5a736d1e89729b180335e72d1380a288fe688a73f69a3e6a1c9d252194812
zd49dfe6f8ef8b3b10a124881a12bfd697e05ec4aa2fc212fd9e00bb7c5d663fbe10bd5e7564468
z4fe495a7f5b046de38c684f26c33586252ece4a11d91d6d20d5be1059aa6ce2eec8e1bd52bc3cd
z188be00c5dcde22af304418e1542c241cedef253be87a1aebbfa5682ef8df27bdc6f55e0ae5dc5
z84937a173b087db8496dde9155ba23947b11d76a8f3ed41e0e8ae5b28cc116aa8c45fcff622d7e
zf38ab4929b01986b4cdb127223d735185ab891b44b5fc32bc8761650043aba84f81cdef005f711
zf349a993bdde1ad9a173248dbb2513f8138aef1b1c870c85d2c58d9dbe1571ada66f056ff17971
z87feb209e4f05dbb1f2795bd9613bbc22a88e0a02f74711fdaf75c40f47f76b2162e30e33d23f3
zf9ac85ecfac251ed61919397c9140233ea710eb0f51fa1d4466e5aac65a1e356ccab54c289b985
z8dbcee657421ab23a7077106192f545e084ee2af7d4097e948bd5f0d48b739e96fa75fdae03d4c
z3091feb25da5cd4644547cc2a4808950533378767eccfbde14505d66040b0053bd3c6c4a5817f6
zbacbf1d4193f809ee9be149aea1e7568e121097542b219ad0317fdf59dbd6149fb9168f46af147
ze1b5611647774b4ea9b534cbf0dd242f3befd22efa01877ce0837c078b1cd94396fb9401365464
zf3e945c9d8a83be46a6e226ca42ccf453f844f8b424ba6d31408814ebbe6752721fbbc3b55dc2d
z9eac342972055d01ebf6098e70b97ee14f9921f4c20939c6c8a106b4504a943cb8506ac995020d
z64996d8ae0b6b1827aff514e910851654c294e8bca63dd2ffa25c357faa1092b3500bd00a77406
zef05b5ba2c2efb8ce9caf4183a747312788d8e4655f8b245e8ef9bcd24846fbd760f921e256ac9
z118b66aa5ad7a6707533ece8ce5c572a85382db494601f9f1fdeb255a3adf20fddd19ce10ad426
z0a9dcbc367d84240a73e9f974e7c7058a3500600f8454c906ac8f79d831bb73ddb7ae169a0f427
zba94ddbb93ff8de6bc873844f09543c77f08af897b3b107fc0b1eb78f76e17eab34a0843127f7f
zbe34a10963b3e028f154b84b1bb1ca02b8a0f5ea9b145459771fc2df6f38d22be1f5167e352e49
z960497dcfec17f43eab7162292cf3924cef360f93c3b6712efa8b4ed5ab6ee6cdb2fe6bf9f0249
z31550566e2564aabec41448e071f7685d6a0a586659bc94a6624d088b44cf520064376e5683c97
ze0e20a70b0a844dbdeb28d16b2e59599e5a1bbc4359931b3d16dc77b1de4b8f239f101d8e91fa6
z8471ea7fb118a615b69ca0e30377a2b475d4acb722e63821507736ff8e5dd1687d174d624edc7a
zbd096ae2aab88ed7299fb56b0ac890292955bff929cbc3a86b56534f1ce4c8a3dba7b89f526db7
z0a01dcaa2584ded3ffa5aab679d3c7f5114c89d0733c2a1ff0e01521092fbc559217dd588968ab
zb27455b540c2d5e945de84e09044dd2f7975aad5fba9536c31e784c67c5abeec20c57a3c35ea9b
z8caaad3a486a9819caf6803192098c7aa593c3833051112305fc79b00854beb12d8a30ce2eb570
z5cdf3afc28c6901504826e8dd5988d705b0ee5b5d7d6223e61dd4e31f4b8c5874886ba307bddd6
za5e214dd569b199cc6b7cad8fabb70741f8d89dd5f7fa7aaa4a521e2f636d51a26d12b0c99f69e
zf6fe01608be07126aec0a807718c27b81cb05e7580c8d802552677d40926017cf6eb7d67afd42a
zddb76b283a316fa06a9383f9cbfadd33e116b2a5b4800b84148e3bf0e82c3b66296e7cded710ae
z663059af4702e592b95c38b3e3b6fe92e6c90823b226ed18b799368372d7b24598a0762f23cd20
zc64ec523a393e1d713086e869b7993e24feb42c3232adedfc9147d992f0404521dcb040e43e19f
z3990fb6c63f6e94076463ff078e96a23b0a5ce419fd135e095a01a516bdb55f85f41697a82fa0b
z4f743c31b551764f4f11bcbb49775f412e2ddc88604f4fde92f87d8fe011a38389e4a4f925776e
ze021fd6d75d4040c563b2801c28ead7c4a15a7b74e35def9c5cf5de04b12ce4e1a7063b3cd8031
z91ba5a3cec5031f847cc7f0effc6d75c2dcc274fb63d57442c69219ef00048f2ec3da7651e9b0c
z22cdd1545fbd28991916f3e3f3a479ef9c80a9280155a89b497d4cbd3f20cc5aaa8abe6fd6328d
z337d5e61a1ea25421c17dc23edaafcbe26783780731c3baafe6662f052a678cd60af2dc3f87d49
z39c40b21389e0c1d98752c0dbafe8c515f7c0fb8f992ef6378c41519db21e551d7125ac3d74f4c
zff5e4fe6ce2b022138a6c6f6dc0e739fee7211c60666795eae7df68318cf87b69c09c8ad7ba6f8
z2a726b6a8af043a5b3dedbed0bbeb0b26acc0ecde9e6751952efed8b5161562aaca7a973ed88d4
zc03e8a9cb45853a543107f334a235a0fcd471b657ed6b46b17e05bd6ce1cc25e64528fd021cf06
z62c996564056516c75579cfab117c18207bd527a5a42f0bf1a2002586fa63af71918b6c318badb
zf403f18434c2fd73b25e6c983f42754e5b01daa7d60500e847c4f4fd586b3ec8c828fb5d055ae4
zc886d09f96bda5f1040620269c2de8be9feda6730bf84cfd21084d1457932a15d423d4e590d422
z9808baeae3dd3bc7a76ae4a7692121430f3640ff76663cb59ec7aca2b3d08c93b144a5aad80125
z9f347b7107e0ec5ca489251f0e09be9f1d20b3f727a41139f7070afd0cfe70a91744bc9f5d6970
z494ff6ff9c3e2e5ec5f3f8d7994b8eb298141faed896db62ba7ec7702f0d5faabf35d6669e7c6b
zbef9d9d4550431ca0b94bab897dc9a4d6468be1122610630136136e28422b600c386659b4a607a
z30b966fd02488dbd2836fc5125c63f251674e14b25a23d4bcf75d6b0290aafdb30f10528c1e673
z6e8ee776e17bbb0a312ee441d36df056db949099439d89a7d64b815d1205dee5ed2b83fa3c09f6
z0ce4ddd661396d814ccf9a4c67ed4e7e5ca0e3336c103e80fc4f0b1d172d7e42c6f414b6ea6632
z7e0f605da99008de8f046d128a6e60b6a3b3c619e7ad8f82e87e6704881969d749627aea0ed4e2
z131eeba2c9f8541dadd298fef22ab6a3d23cd4c6cb96e30e0a3056a8d16baa6cc0c89bc1be6f03
z64de08f95ddcba068e6b6028d1e5e756dccaa8f6f3eb0dbad78c2bf45e8306a9ecb6c042569b07
z72f7c5d2114b4929425487bd8e9440f8ac60423df542908a078ede125d551c91d913ed29f1dc1f
z022107a757ae87d699fff026beba1fa3ea4750c924ed74a98ed6d93a8a569be06d7fb057270a38
zfeec28e48e6b22f1b4d681c274198b00e5d8e6d298247388696169906ae88917ced29a4a34d64e
za42ddef5f62d33b2e39d52c871854950676d33b576ef9c3462f18453776ae4776604604ad6e01c
z23f08f434863e724e25ca7f395626c0826cb6d96395a317470d0f2ceebef7555ce96ca98de1b92
z8d92f4f53d68c98d7bf47754656a6f682298d8cdb35532bd2fda91e934104eadbf4188765ba30a
zbe21ab07d641dcf7280c3d1cef0b0dbfde14731b75b22e539265f88971a21368995dd340601476
z7de33a3ec5b7171ab680a493691b491430f0f288fbc2d9314458cdb60a37275ee2fdd4d43a60ef
z042234c8bc65632229ecb86c5e4f6d1877ce74d4e5899eb9ad9170af1bdc9212178fef99056f6d
z7983193c30f3497d80b14110ddca4b4867428b523e6b5f027371eafee60dc57b4485f2d75ef8a7
z3ba1d9cf5980f9febb014e1b9e2e9025b2b131badbbcac7166bee4cc2950121e9e6e96b2a57a3a
z8297b33349e230bc2f741506174d4c5db8a2eed99bdbc034624594c38c3d67bb37586848411e48
zd4354c5f66da8cd3b09881e897b1406cb270397c69cdd86f4826c26bad4c3124eadb951eaa223a
ze17e89f8e166a69d425d2fa322ed741f36aeaef958efda919777592ec0167189650c2cbde6542c
z291e831c627a73d95d88127b488fdfcb2f43b82fdb52523b37518aa39bdb580f8c6c1366194a03
z7f35c2ab047424911c25d06d4137534653e69ea9869aea755c5c6a7000a69e88aae02e59d8a146
z84c6c311d45b27d8dc68fead5beb26cb9a6146ccc7728e6cef4c187b4a1803dc5b675713eb3704
zfe76a6576635b3988f7503e10c744b35243976188922a511e8e370735a3787e23b060255161b6f
z812546d270b7352fef0b638ebe87d17bdb5c1e44e8d416ed49bc575df25310e310afcdfbe65ffa
z90d970a129507080c4c648d00c21d4c565da446072864c8ff567800ca6eec72a30c1081bb3255f
z1be90843ece5a4a879ada2f929fff179e4c0d66e72d70aaf0acde279ef1838f256aa59d47d8166
z9aa29347c4f21f50f3abf2b55c17847c1c54639647bd94849be5f7e1cf645f8a12890ffcef3496
z93cae3a2e5142d58e3bffac70786ef87d1299ff4679d311e2833e7e9b1f872376e100ca93c053f
z323fa6d6dbf28c3708a0cd286d17a60a1611a9cc54febc7a8710356501e82d37ab5d9a99c1d09f
z25764a0b4604d645d5cef4f3e5fef3a44fdf863163fba297b9307de6c4aba7733e3757d3795344
z0bf7641554f71054d13fbbe7f5fdf343b5fe4b8f1ddab23c03b58fe131dc9647456438b0fe8551
zf8dd244eb20a83eea59ccd0c51102246baf75a293b4a1c0125d68ed81ec15ff1fb89a53084670a
ze3113f2e93bf5ff155c012e51ec049d4ea6bc760ad0f2ce82be34b92705c27a17b9eeb1b660da9
z9f72645947d451b21f381dd82dd21962261704bd7ae85c1aac0c7c644a0b391017fce5017146b6
zfd5b85734648e8c2bb3a5f359bcaf390621f5fc12331310a20500929cc22781908c2b09ea0ff34
z23f4ff85b269429227908f8c271004619fa14f3602037c089b1a4d7ffcbb3e9a3b25a5f62702ee
z1eb2be85a45076f129c3b87b72f0857e031806993d10f04ad74b8918d151c88756efa3ee74cf20
zc7698d3e0d283f8bfa6a814e080e61fef1c76864bd8fd1c7749b12703aabe79209ccd7ea733cf7
z1de5902087f02d35e99ccd4e93652636271965b7f0811bc504991190a9f7967aa959f8e7f4ce21
z664ed0f9858e0fa42839c229c641cd4f2c383be067bb8de2bbb5c916d24f781f69c243d761bbfb
z3e64825d0ac9afb644c3ae92c159325c5304bdab997b83aa7bd8a8683cbb6128b6cb5b4fa81375
z67dff2ffd1a7ea129dc66cb3627aa255a81afb1ad214fb2da338213a623508969c30476eb051c9
z1c72fdb6b2b7bd9dc40fe9c0c1730e8c19d4246ceba1a223d404e2be7a4ec5f2f1fc2f7e8e1c88
zfe6864d97c440c3cf6a52b382b4506dad0ed490beb0564ba326456ef17f636d547d827dea8bbf6
zb0bc32fd371db9eb8d12ed9453e656eb432712bdf1967c10d6a5548e115f7a5bcb2552ea618cb8
zbc67d590d67f35a4a304050ce0043b3badbff44712833ed733ea9cd41fad0fc34ecbcf512a75dc
zeba592e06d8e9c48f27af516855b6177124c12c8cb97d580fe1f9ffc9ef37d61bf8e945feaaf61
z0591062b97ff65f37688158daa272821194e75adf1eaeb540c06e1df2e44a78091cfca93a85d57
zfe19081ba28bbae3e265ccaa288c9bfdef55e3841f631b5ec8a304f485d26c5ad2080b095a07e6
z7befa24675b6eee4496f102f677dbe684b0ba61ca7545eabba0f89b24b5094f3454426dad82f6e
zc1cd2be93a09acc1a0e4e333ecd6e4a879b43e88116ac5691e84164903b8c400c098a2498e1a64
zc8d68a453935fc6aeffc49a7d7ec53e78b36fe2fe57bbb46d9beaa7d6b91148cb6cbdf765edd47
z6234463a7b32e7eb5e3143370087583a896ae8589b2444ca0ac195980e92491112740e6f6c6b4f
z5c54e2bb5374c682f2575fa9d066b747a3886ea81b48515fb897e10c3f50bc5fbb6c8462e3659b
z1caa54fdd8ffab381cca85e7ecc2943dbe92bb92bf3fb7d0650c72abd773ae23db7d571cbe7c9e
zfa3aa9b91934a632f180a4a62306ee7a888a60e1e70397f120dbcbee171dba3b433e0fa81353d1
z1b1b824354fe102abe60121e4055c5c59b6d0e648e5f1ff0f7532661c178b8a7863af0af769a57
z34f14ebed4d3881b9624c87ec933a14f1fd6c562dc26485c0e8fdcf46ea5119486e72729fb06f7
ze508ea8f98e181108f0b49dc69f6596937580f14c1986c2250060944ea1fc1ece631e2970261ec
ze9142c63cd55ce18e252dcc90010ecf6b6d11324e856c51edff7f5971488f3f230008ddd1d0c09
z42a2e2f9f9b9396b4c4bc5004b3ba0503271ff2a57d55d3853d9eb9f93770947b683e05c419a61
zaf13b9729f27b7c243e9fc7f2826948c1847eeab38126e3c735eba05341b47d2fa785e946da916
zbe06a9baef3f056921032c0c572103ea96f5a016030cd7bde61f6712bf586b221cbda303ae6a92
z4f725c2f7811fa45be8f0b42473541da7fb639307f154d0ff7539951a29473c143b9b35b5300b1
zf727f61f4dbd50de1dc0a7176892195e0358b0a97e28665c605a3956854dea9cd434a71e9d5905
z6bef4223e916e4909a5329c4104f06c271c76b0548913eadabc66b156ec29c34bf30f939522e54
z0516f1671f22c7ecf1f8eee86412abc790f09077678768aa203da4b0690e7c114d63475c705bde
z9e5e6a19365cd144a2b03321e35fcbf60a78d897d643c2a8a58a83482d37abd4711c8ef8095f72
z2225b733176d0647d39c416061826cab2a75bb9e6a01b742a2a801c0095584b25d4bff968484e3
z59ca49bedd354c74c6fc5342b34ca74788181c79510cfb3d8a9b6fdd74f301e44db13206f3f180
z4d8cb20e0ffcc093c0aee1e14f0bfef41446380040d2312273a6be474d57ebdb43f5dffc94b8f6
z8cef94912db41dc44376eb1e7c7bce015cbd1126754bbea1b45a7af0f98b9f93d859abdadde8c0
z2546bdd66743cd09a8e69c98df4c5e8be9597e91fc85f61973f176648b4fd7ba6e5083db32591c
zb68fa36a6f6e847b8e391516c00907c21996306a7d31955fe9774721cc0e3d22056c81da88fe04
zd49dce9dbec37148b05e3adcc5ff42ad928f609f0ff9bb74f47c336791634369a7c4c0adef2422
zce5d36427bfed1eedc5b869564895a47a7157e77f869cc22b2bc0dbb15ad8917dd30b4354f31cb
z5d378dfa53149dd148f7b99cd9c939246c7591cf9d41ff87a84ae83274a8fe05ac8698916f868f
z3b574412f3fc17004339a830511f261bd97b78ea3fbcac2d14cd5307be1c960dcedc76fa699400
z20099e489f59247fd8f3e7d977d145ed229b65d9936ccc126d423faf3e58c5c81b34906289fb57
z16645d3fb438c05c95eef9591e02a18a6da86bce85fc0e1dd960d75a1fe82a7c341390d35cf307
z85ec25fa51b567b0118fa53391b17b0d79d46911b83b16f0ea7af9a2a603c8983298cdb16000a2
z04b3952d873f35fb5ebda5f7ca18874093ce569b67aa350048136b89af53359bfff739abba0aa9
zc71a1323a6ae53fcdcee1f002d0dd7e9a50913901ef567f41babf276ef76791acb4948d09b123d
z9b676fb5b9dbc6ceebede4dfb4af63f4db460616d6839d3ab39504bb19c93f96dd5a18ef2958fe
z2c772f5d54cf366168283b8344417945bfac41637b6f3349518ffcbc30bae1f6e84ed3c0835f9e
z889cb92d06fca8f04245045eb6bdf715c8c382e5778234c898d5a0d25c7d39fc3566f984b7be94
z7f561b1a6d716f1dd1c1adccbc00968c426dd0e9228ae3731ff039d75738b91a122218138f3725
z93d90ee8b0a8a967aa323ba8b7457deafb406f4479e28506fbf152bb59426454bf387c2dbb724c
z8856517fa3a9461f2ec79f6c9e8d8d55e8152c12796fe93c571ff7539ddfe27b3c36c03644a877
zb370cfa33d11e57ccaf5d7ccb8fee0e76b0c85187ffa80276353900b18cfbdfdef138855474854
z63ee18b43c5b8bf0b93d3f57a2d1b5ed7e695734e3232126079e2adcd5049a52ff7c90ae38385b
zf9811ab606efc62118bb13ea1c93db24d0c809a6698a53f3264ea3a81b0d962ecc4388214811c0
za2f0ec7ed5f360a85b44542e76002f0e744471798a614a070f375acd45a17746743170b0a8190c
zff6e4c4b30666c6b6aaae357b32f9af0b0549ae6d7c9d6e491d10a1bfbc6d4d9491716aa90489f
z4ee999ac2f9fbac9f14dd39159bcf9b70ebad37579e26cbdf643c6c1d9b832e5edfb95a0e67925
z3e5c0584a422cd11761a989a5ebe1399a59c041ce2a6ca0c84ffcbf638affa54710e694a3e1c9f
z28164f79b617303b7a0e2b18e17f10de18bc87d9430c043136da3577cdce833a84a43d79a8ed7a
z28c49d98d9423cb4f6c9afb47a02add656de6ecce7285a5e0633529e9a66de2b36577547f2b011
zd889dd9ee73f9a3985a465d1447977cd9982cacbecbd1e6897d60a01e634dc943db2db171233de
ze0a97fd552bc2c30d232fb2bbbcef469ecb962c6f1e5382ff066972774ad0e5b2e2f51522665e0
zd71800edf74ab0a4c79e8b6fd3a9f0f438dc4658b5685c409c7db09c25812a56bb092699fe99e8
z2eb89b948b36ae71df9e46ef69a9dd60b0d90a55c84240c2524c11476a9065fed2abc8bb9140bf
z798ec7efeb7a3472deba10c97a3594f8aa6d3487749ece4e01ee1503cecaa96e4f3d79123209be
zec4aad83ecb266199107dcaec8e81f3e0009fdb3b7a46b3e181c84899dece3bbb8816034683275
z0b73bb89adb114c4a73b665f18c9b74208651e54bebffdc4c439c757eebc09be37064085bc7e03
zbf4bffd6f8af441e4b8ee46c1e5383dc01366bfd46c0f07f9dcb16688d47abb4bf8ed80c675d81
z499d302da4376136cb124615be457f5d8e61298bc36cd7f64aa58f8905b89d007ecc6a62f54c69
zfc83f47ac4f4baf6d6d92d5b039feca75ef7b38bd20f2bdadb403dfa4c297b11dcc4b48e000db1
ze2f59f0e3aa31442353fc79487e0e8aea934bb13d3d8748689c1024b473fc7a7cf3ca4d0b738c2
zf1662848ff283391f7aab46e121c4aea7c8fd4a6e5bd5f13961dd208b5feb7bae8f22225c20ef0
z022cd0208ef2302fe96f6b236e24785f423f9dd0e308a26676d942af134610de3da88504f73e7b
z6e08bbdfc5e84a33eee921ce62150a838798c7a42ecddea0f8adf4bfaf8fcfa66fcef5100fe0f3
zdea34ade5d5fa047405ce21b259f75da839be08c0b7e309b97278833ec9e64d8e943a9e1c5d92f
z4aacebe6a11de0d4e4a014535564827b0fb99a4d3cee45af669b2b359135ec24f57269a60bdfb5
z160dcfb594fc4d191ea7bac13560a450f9a8bf9b649fd22616baec9379187b30c84d7c935d50e8
z599b64017f88c3f226dfc0a5aff1fc1e252a0c96b8f410decb1e6ec3b97feac45c97f4b503a515
z698b8ba6e3fb3d6bc2704fed93762177c761caeaa2b7c3437a10dd835f86d26f80c716c2c143c1
z7daf130b8672110be7fe23c6ab30d537ab17e60ea0151de64d22418718825f4c7ff237c1572f3f
zb18c25ae6b593fd6653042bcab68dc076fd049651cd0e94d9d53def8b7eff7471183f2604b8f2b
zab1d0ddb7cc6591cb09301fce14aaf74b059945462aef95ee9ee5a366ffb34038155069633b4f2
z46c4c86d3c7da531aefc89fe686b8d9e722d8dc082819fd7ade5fdf116070e92bfd248f51fa784
zd7c42abc1ea82aa89185b850556d5cd685528230d1cc239fe371d2cf62bd79117cc92e47258b6f
z5b7ae5f989fedb92ed32efcc114f678bb95eccf9a184c0350a043e39dc4d5dc7e032b3faf66da8
zf4fc88786381bd2212bf350ff5912fffef546aae7b927d34deaa223b6809ea024c029e7b0280ee
z0f82a030bc9085b6bda4c832084caac6d30374ad0ee7d8fd1dc88ac77354eadc44c1f0754c6d13
zdf5af595538a634ab8778801a7d2add27bb26cd0cea1b2d8fe7cee4e2a35fe95eeae04a82caf82
zf040678c4bd0082ef5e57245916ebef3bd33a33112ed2731d19e01f6a3c4cd790b8caac3c8b4b4
ze7b3f9a58a3a5ded2623f572ed147b1bcaca96c5f989b35ab4124b7860aff0327555155fa33879
z6b044283c8d90e668dcfdb2ba0e30b1d0603e86227a57977060087730a8b6e1f2fc4a6f44a898f
ze4b4faa916b5f44ac319dc1f9a243531b67200466f7dcdfd3daf0dc6a416f281f35d2a9b3709bb
ze42caac78c4c7a36b8aa15abb0444e54468ccf21ac85118fe217f9fc23e796db7dbdfca42f2321
za2545d3bbcf617b014ff3638f69f48d275b6571bb5ab0f3c6bce14e727339e90ad01e079a5fe76
z5615e1067aa8dfc272940904fcc459ca81508e0203d5b1bde5a905844ed9d20690b6553d715cd4
zef330850545bed8cbadb5e799b0bc25a4538e9f82bbcb9d53c5871cdce5f90ac347e0014c3e5eb
z8bbd78e553380352afa09df834791535d20b101d2b0cbd1d052123999e470e940b4367dd2399d0
z5027cd058748639f4795c101d07a49aef762d8b4049a2f04fbdb9844d6663574716c64920c33d8
z35e91d6ab4abdfb23d9d39d7e2016aeb01d5a18d74e446d8ac7006b18f95c3377bd059fc06e936
z7017656a3e767518a29796f0e420cc2074bde98e84841b561d9989458f203be66f4895994e62c2
z14bc8b862026884f73f23d78df973e1b3221557ee48f007a12ca68df1d41cde0a37bb1e3fc699b
z59b7035cba59f8889e588e4bc7e30e269835eee31d5c13d1916c09b315b09fde4c534ef13b3e76
z7c96620442d6cff5e04c3da3d1244ba97f34bb1804f432bd688155dae936d2236db36484a162bf
z3cafad7354dd7230993a663241c7e121adf2ecfb3d9490f0f63b968f8fab111b69ad1213e25317
z5909d81271dee54cf28625cb0adad0690bebba454893bfd87aeda8938a72a79098f448d7d19b3b
z9905856b8227856608de6d2679b716f11cf498b86db4644c8a7cd927ac8c6d98afc33dcbc9a17f
z2a76b5790ad5902ce3681b0c0d3c8bd990d443f5443906fc3768b8a8e76c90ebac1e11a7ec3244
zdb6f01d639de6b4d08360fb4ad6df25f2accedf12a9e1de42325c511d1fb9bc1bda0b412895b58
zdd05fb543f76e9d1da297271bb39216ed38d5666437cfe269b4692bd273ed7a67701e5f7342e32
z70270b3ca6364e6462696eef85c43409e8698aafd06c4026b638e26abed078ba5b260103c78755
zf8448348b1aa8eb4eca38c464a6b72d4f3a347195d8b5a8d6401a0ec853bef74f4f713379225ef
z52e12e89d88afa49896cbb8563d62f18f37b20979d6c9cb360a7e88504a21518b98b5605b7f4d6
z1762e832001a5fe2a1a563f9e517881847c44533137e5e52814ee05372249e64eb696aec956d8e
z24c246083fa634d8f08cc260e8f1f6b12bfa46396557f6ceb4b8c01de045d80e5a3591d2b3f457
z0a8a558ea28d7f5bad2f35814a57203d3a66a659a8007961750325f5d6897ee2a84f73923f5b48
z32d8054577829d57b5cdc69666106aa4971b1f6b32b26c5f55653b08989c984f7853e98f258891
z2cac9e7fa00597347488284963cf8fe54585e3127e387406e27b64b770b15d90e3e8298c5712b8
z631a62c73b1f1c91e52ee2b0c4bc5dd17305ed400f06b938eb090a572eee125f997f9449108d02
zf73ed6eb0c1179c8c5ff96ff71ac55c56b1ebcf1ecb1a2cb6025ea2cc688bc46699c72e8a283d4
zec0fbf1693da5a57c20ecaf54d98d122de119f7fb19af75a63573cf72045799842e572b291c6be
zaf85344918a3f3aa64ec177f075c8f319302aaa8a095a923fe91d028085a230bc014e2f5f23dc3
z94c2ac43a1aa2770468e04b99699e33c7f3e60684ccc8b6177421c8ba050d1cb133377bd9f7861
z9ac1fbe1633d5fde744b39fe5b36a3874550a71a8f389eae0dce6bf9d85d8271ce677f9b899a90
ze861cb463fc551fd264b42a4e78c0a6a3cd2791da7996df166d3a54d0468a7a33aa1f597ba6b14
zc0f19e0b33c2fdb6bcef9c521c59aaeb587992281d33ee466e62477e58e2678301029ae1c54045
z089e25c755b9b05f9d8e2482e4dd81dd18c5b360971f6a0421cdf2825104d524096fa1fd43fdc6
z940c9de64071a4bc47b7168b62ef68aae649e4cbb60b1d9c0434c43afc1d6b359fcf43289217e6
z73e6fd6bfa0694efee4862d37945b3b47114702657cf5fadffcc9f8d6ead961b0a5f0e93af4af6
zc26b233704329e7ddb41c13fbba2b99ab71dc34ea01b27a915cab6a8eff322bfc5ed2ab85d1f0b
za79a4d6a55ea85f1c2e48500b81e238e2fd3dcaceb2d9fb452fb11ba0593ac8b35e91a09a25079
zfb5bef36480e9946ccdcf97ea33e01b8a71d7bebd63b962d588219a14b59f05ee3229ebbd5b853
z7b6e55570cd936d373e8229961e0bd96790dd3d5a07a5aa8981ccbc44ead2cc98c55b4c770d444
z3bc53bc08ed10cc9a851937917b8dc9d00552d1d309742ae932cbdf07f58851ee9dd30c1bc52e9
z82adf66be3cc3b8b1ef398857635bd79409dd5139f6606d5094cb7b722589319de28471cf3581c
z92fc20117a56d72929185da4cb9719fcda081d2f68cae2ec671e5c345c8da0ce3a3168e73644b1
z45d6338f057ad1b76df09018577c72687ecb6e64291b08f78e98d62c9bd2bc9f78b20ba0c4de5d
zb3f59c397e1053ab009b068ac5809aeb132d243e2cb05c921498f4a6c4324fa1e3810e234a41ca
z84717f76715ccc4773415bfec2e075f2d47f0fe4f39487e6231c0978bf6a991257784c7e176fa9
z5e56c519e7b3e2edd66ad8074f3fa2cc32a646b3ee1a2efc125e5a1fad3b5f44f2ecf52b4e90af
z86d51fcaa5cc6c134ec76a5f830a4029da0df9ff5ef1809ca60891547ebfbd1d6cffc341e847de
z2e7fcd1c3cb58c2f2d04db1704a4e12d18fb1ef3f849aec2a8235b3c9fb456c72d1f75565052e3
z2eb9b680ece6625cc949286d3e2e06b1ea69d8b21699fcd4608f39dc8d5305955320a0c7d94e79
z7f37fdbef6d933d774273f4d78788272456bcd72970ce766faa330c697bc84737bac187fccf0ab
z5bbd98439d41d12780c93bfa96036b7f952f44d0ae8f8d970387d39679b3e089b9934ccbe73bf1
zaf32786645cd43d7002465129b88aa799f15859d141f31ccab5a50e77502e6346ccb17f1891ee6
zc95df4fa360121b3c96bda10443464e37602c4cdf3917e76efecf86277b32d04dc3f51ad258af1
zf22b88d4c3b8eb2fe88b9d74b2478488745569bd2f06edbbd45c2c740f9934bd4b2fa762673304
z6e9375e20e540ae4a7898252ee0893d2d087ee6429a131beb2badb8c3dc69a1cabdc9fa5778ce4
zf8657f651e00ae0e85a236b63f5569327a4dfe987a8163b8817ceb70967f597a9f46710bfe8cdc
zf8f0c05b9c60a56cc6a8d2d5ffec7b896b8dde0ad880fb6ef0c1b510a3fac44693953fcbed5d68
zdc1b2ba7db67eaaae259c06b9e04d59cc83a0567360e28c6b4f8bcd0640869f3c51023f24c8257
z84ce50da396ef479a10ba38c2e27de13b8d08accf4332e2361734ab572fc8b7b5d5900d35215f7
z5a3f20eaa52be39551e62b9dd40719419880e8343b61b45e3f298c5998cd1def1e2121793aca96
ze96c6e8ec52d4300df6d7794a2b501cec0b600f7782813f76ffe193407cd7c831cfc23a9b10bf0
z87c0e0147737824a3965dad82d386f84033af36782aa886d739db87271ac6bf82313682023c808
zf86adecd4864cf6cb93a5a2afb0c3b313a89c24674e4f2fb09ef8ad1adcfbed7ee740a3dfc5611
z625e8de83651e274c05390ec5ab5bc600108e8d1cb3ca0a8792ddb02d79d9194d81320f5096e13
zb93c9cf8b33d75957481b4961d64f4b5ec8052af281fcf5512e21845fad8c1b27d06f61d150ecc
zb005afe1df388762911a160d3a30b6fb6d9b7e462661e70974d052a907603abbf8d97c95b34d8f
z823852d307356bda0ac245b88e2a9bbfb7f3e504c38517231452d244b7f016864e6a227839638f
zdbb0c567d3cc719c8da268c85d21914570ed34e7770104d4b0e624b25b1b39f83c7ba1e424771c
z19e10e994066f5baf374ed4d8a9492489788deb5d8114e6d848d6dbd7f03ee9439896a0efe7117
z42351f9bc690b94cc747df531613e1e18c069285be55d91c064489fddc8197e50d02379672d5ee
z67f9a1be73ea5204d0ae2b0c4c6afbba3a838fad2aa4a70c5996c856a10678378ef4ce6c93d03e
z223ab0518a951aeb491e15a13150919e2eafd73ae84d9210eabfeac6538f51fb75d2464ffa5579
z118d56b3ed282e59fdf71930a5ceec6fd169b989d77059dba592cf9930b596e7fb49eb3c66e773
z505e9aed7bbcfd737c28831b4e10204b3df289dd93dd1f4977c3253841e8d6377d0fa1378c3a06
z3b67782e116fee4629e04ced86bdaa4f9f12aaec2b4fc5e8b2d4696031802388061c60d87c9224
zcab9840fcab6b2579060c52547429b2114211459b7869c26932e679d53b741c8bd45c13120cacd
z1ad51af61b54c8371fceca1c2526b14f535e09521450bf854f186923c3638062c1c0fe857567b8
zb7a38765afe0b5491619002c37467af44cedb47d30c090b99ad882aafd4e3c27cde771498861f8
z4e5c395ad359864832b21fe4d51dcf7ec862ed4c9f713291a5da742c0bfc4b694546398024e39c
z9b15dd79bd04cc649f8e042cc6d5c9d4f8bbcfcd9ad065f9535117007e297fd088db22abe818fa
z1e7f7478f46efed07c0f60c55404d6c7bb3a26f41ad6081d438e197eec45a24ce0780690cc9e98
z4b216836c1ef20d2ba5f7b98ee464e16cc09a243601d01bd991c3cb3a8798709b8eed084f3efe1
z15ea4c50da2572dd62028f6246e14f1e0e29459b373c3c5e690837c8e6adb4841accde964e287f
zccb49edeeeda403b5770d48ca36f3bb9d944c7cc7b3b80d9f4b41d2b7c03e83fcc9a6c28d1f407
z8274fc1b5b6af47dd84b6874b151886feeab925ed52b2e81a40743d096f3c58012b6519ac0ba37
zd8bc17c73b3f5720bbcdb79e08d0952a4ed26b109ffca5b7ce8a5d5214c88e937788efbf17702e
z154c100796d915bd41875fd0b237257225a7fac6803cb5d24da63351d758417d1a76609f472faa
z9a9d921e7ba4d62829c9a8d4a5e8945190fe6774be25c6e533ec32fcd2062eec666391dc4500f5
za75018cee778bb84a001c156d5bc07da2a5e4403a878c6277be124eb37b793252b2ba8c63cfa08
zee5d5ec8835234e31aef75f60caae1a0dc4f5d15de5663b8c126bfcdf77cb64f542a58441406a4
z42a46a2fefc15935a43fc12e6bf536452f2dc4db29067e801c26b1ef66ad048044a6f6b8607395
zf323cf752ae922ccc0e073e807c34dc3708d1cc0935eae3b7b5e0c943e469f28f44dab49b297f5
za4d690eb369573cb5fe9c9c8363dd1b6511dfbb38d3de963ca70711534b068fc3a1dc5408c5500
z12987e41c4ae8ca685aa12f226b038b4213cb46af437bf6961e803e7bfc30a12fc982251f7ef74
z6ffd96de505029be9b3de1c56cea7c4c42cb75ce6e51407d0b726cfa5251a6d0aa931f390f8378
z34094c960c4efc22a6cc0e72ba53f0f7f02f2c3e028edeb6a9ee585263503585a99ab2975fffec
z9d4fa9addb241982521fcee1a20150a71c5c314171193bc070858d48d47af5cb48dd1e4f5ce38c
z37d498cc7f98d92171407213001b05c4fc3e1008cae4f1a0f3f1cea489241353be639ba64a46d0
z3f79ed0e21469fb05f1bf729a9632021217eeb6876791b02ea49ab02f534a93e93f02e774e45b3
z5b8397cc292882ccae943912d6dc6b2513a2981dbabde70b11b265601d7c1ec684c9529d316c78
zd7e40615003a13c53333bbd96e8b7e4fee1ee53cedcbfa615a5084f1f735a99df04ed83f1c24a6
z1a6c1309ce6fc940fe75d225cf895a508c96b9b11fcdb41d2b3882306bd37d5f9f9ee69ec6b86f
zaa8bc55a858920813455f51a56525b666084298c85faf6675e019a2b63d35a63585eb4f80d3e42
z59a3e5467863840d05cfe9543d80835c349fa92c61a0d4cbb9c4133a761532a3f22acdfc34857b
z550ac1f648458c106c66cc557a6b2f13c72d37ac26c254094135e8314a6ef61f97f227d61b1a09
z4a0608be034f3bce0f68fb687e911ffb7f7ecb6838185549fb3c2cced1ed5c4cb5579ee772e7b3
z6f81eceae492c44227c06d9a2d6959b0c73edce8413204ef03c337fc5991586470a019a34d9875
z45fccea5e4aba6f612731faca0c8ac44ab3afea6941601389ec70277723b35a824309a6206b598
zbf02291c811e6d04b63d75cce4cf6480f124a5143986bf07615480bd735b115f5579875c701787
z9a800785d79082b0d3b9ea9df90758a2f4a8df59eab841358ddb9c1646f45f86cb628ba1711634
z6aa14f121a71c19e543ce51c0d3bddbdca5ddd66209c3362edb7d15ec239fbf8bfe02c9414cc43
z54a2c5920202cd7192dc5d8949ba13608ba55450e042c8c7673df6675fbee94825980a2e0c31ea
zb35cacdba6d83bc7e1fc06eae09ed98c5009fc9ec3c6f18217722bdb6a7eb06ad96fa554f80583
z642fe966db557c366d29ba651a0759b6ee9a0c24dc8507106d5cc0909a3851bbd92be12302fa24
zd51a549d360567684c46cd5b2dd51041b950b41491312eebbd4c193dfb217c60cd277cd10696b4
ze9ea3592e1fc6097d10bebd890a785a003b34bff198bdb41b41812983a35a447374bea5b887ed3
z67cad487fc5ef9769f3ce6c6eadbe508a8b76f265d7566dda13530c83be5930bc2ce5208ec1881
z409293e8f161eefa28d4c77a541e57338984b18cd3238552c6b22502d33305ff515207ac7a7a42
zddbfcecd520026e15cc3d7818cc39cb09a1e62a46e0ba35ffa92cf58cae8b37b6cf55ffc257c5a
z22e8f93f4f8370ee489c86acaa9d556da2e22ac952998283eb29cad7cae5c09c74e67e7d8c11e3
zf7d5f8aab796697ef7f1f9e69a6fbba3cff17575706de1ff6f928547282fddefaa7b419a9850cd
z46a08a173e9e03e385524f62541f778e9725b1e0ee1ebf6324e76c908c2bd0aaf0e3ba3a72d812
z4f8743853fc84bd066059bee041aa436c39a63ae707b491c9e89a10f2f0a09283e94be488a295f
z4609a69ac9cff500d8d04efffcac71712cb80c90719613ff97ba7e84be25b0f9c7963508d7040a
z9cd6747c807b0ed4a494240ad4fcbf59d267925919c52bd5af7a84adf15c4a6c76caf196b87895
zb7a738ad0e88d067ed29a5f4b1e726a9950cc1337d52efbda2fb133239c1e844ce73b2c94b642d
z9a3ef5bf78acbd38b6fc2b35a092afee8ac7b265c1e5cffd5fdffdccabc6c4451a2e4e672831f4
zd92f73eeb75aab1017c1299f075fc6011af52e608836271c6e0fc981692830923b14bd55bdbc65
z2cf7cfc77a26226f5680b9374746a286699bb47e7445fca048dbab0f0b4164879c1a7d49438e45
z4f791f008c9e8ebb8f3731f213f3a2408ae9f51be5f3c0d10a02ca69918008e45db20514532505
z4d02ef87ffc96b5ef8c72579b39e449e4813cd16ee2547e28a3f3a6802409ed168e10eb137f486
z723a03f6a2145b734f61466954287b6c062a630e9ac7ccd31a6ca37dfe4bbf2218deb3392e6287
z3fd204ba71a6e3876dff9b4cff13dc7e31d2a356464250c5cb63ec4c713fb4fac20149512edbd6
z46fcc0005761f03328cc27940de1d26072c1d296dc6913920d44e01cbb0ef68ae11d0656ca4245
zd1b4446d8fece1e6a44f357473b83e1024e43286656612a0bed2406e6b49568c437ac14d7f5cea
ze6090d356b6a7ad400c0f2d6b49031595dc0a5b65604f0b5e7f73efc7c4a6a8086f64ca53897e0
ze6d1731be8cf69ca60d100bc470d43c3c3804b0c53ba7987489f6d7740610bae360a106770b500
zd883396b861038d4532fe55639813dedf7e0943935b2381e0da7e045f49b5d4e283f6d4326090a
za3966476b393aeb1843d44f18706fb054f4a99b41e5541c7eda9579fb92f659a1e31eb9de6d736
zfb6a9f87a7505b38a39e2eddf20586c5052e5c6402b2ce32ad6281ae03c0e8224d856b26203cc5
zaff84a327e5c7cb20785ed646405d5f35161e984f2046f80037395618bb56a9e183e0b6b6f4bf0
z06a41f323fa9672d8ef5683b12bc67160c88f9b05c69890261295cd5ebe38e2862ed060493a091
z7a662bab5372b9a02fb017955ea4b981cc522903b9265e8c064e823d0821b6ca9fdd1069ce1f84
z834c13e88289981324d692634e9a7952b413ea9c43462b54659ad67770ba269c53c83dda0ff3f9
z0162c800afa3d51e70353cd1e20051f30824708bf7e1b1b4feac0f15ca09b32fcffb81cf7d0c81
z24addce27da8458e0e603e67bfe3bed4c87ecbeb897591ff718405f9421687d81663afadde3271
z862d378d89eedc878b059109b034e8463795668a742d95512b93bde163d572c95e4d7a25d9646d
z7618f92be759bf10dcc86fdc7018ce8180871f9493280a437836eabb664bebade328404c21c7e9
za9969023dc3dfab9dd1ab07a213f39525779722180749014a12d2f40dcfee95d21702023413805
zc2eac64a7a3f0f5c3baaec1e398843f6cd55d414bb0e3d3ab8853ad34ee999f7ccd5c4cd016c29
zbb1e7308f9c8a693d793737bf39a2e00e332cd1e4a7e6d779b7137e3a706630c2c1a4974e8288e
z58281b359261277630d682401d80a52396f4b81f7ba81f45f28d7a5f197f479918c0444eac8844
zf2d342ad0578dac86753d3f567f9a5739373132ea43f8b57589f1596184d442b129c9fa197f5af
za8d754d2e53964ec64f53bde998be3ecd357ed63afe086cf93d82ca9498f508f770029f8218133
zb48032819eb9bb9e29b6dbc31026b7502e9061859b9f8f087c3590c2aff7359561d7717bc74451
zcf61c613da4d784d22e47e7a8b8b8a02059ea5b11749ed0a2a177c58cd2712bc3007799f7ebe17
zc2d7b723df0fa1556ae20cca488c07ff496ad6f9801c9fdc28f2c376b063b2b37b3bd3cf33f75c
zcb30a48063488d7c54dbd3011e6f15314c78e287c9fb2b9b7e2427d6229ca9d69268047eafab55
z22aa32031de17ec6572dd97b51d093ffc88aca5cee81a115ff205efeacc757438234b61bc20147
z1ed540f96e3442a381f5533e2414a2dc950f11de52fd50efafbec532481fc9bffb379969b7ad57
zbf3f7ce46e90e3fc5cfdb8e17caa052b752521e01fcf7d99999ae43b1e7fc787506b3cc41a0448
z923ac25b6032a9e2b52fb9829a42fcc9c07d4931ecc2aeff58d82889204830f32d448239af5ead
zc9a491cf3b7a9eb13508349817f494c062de6321487c25b866879fb2480ca086344c11c7d5886c
z5b7d02796f21d09047aac6191c62999f49505b6b954dcf2a534ce9125b4c4634e8317361bab398
zceb0b88b40d2a832afcf4dcd42bf2671fe6190af18896d972e6774a2ccc72ad08b399718bcf5dc
z6d1439b85b781eb90c09250952a4b87e52a3cce5b52528a5adce3422c7114c5daf9763c40639f9
zc3aec3a172e4cfb133aac8f440d79cd4e3e9f2fa5b6e46ad6dcc55bf570f37e86a2053efddec08
z87b684881dec2a2112c5710b9cf55583fe2e1e7589bb913e9c25c72a263ed66af381abec881c70
z6a7f6b3327743e887254777d66f50ce7fa9812bea142e53b55855f9948af208fbd2cd2a849c749
z66b0b1e5f7c6f037b3aae25099f3a8ddb34200813d1bd76825e20fa6b4ee3c17c7a17794bc1615
z23345c273cd31cd6472f0a8fdfa900162b76d8129e529af36b091c98a4fe11a432c83cfb68c73d
z74a477a9b0cf1e299356f1e54268fea1c4d410cf7d8abd9d6873d9ad073cedf46159ebd5d44ee6
z5e6f89ec082ec17e34c116d2d3ddf0c5481ba59bfc94f2e9e2bc885d30ebec6857331f7f18886c
zc21eae74a54991784b45d81979b37f8765661e0f1600620c37c60e931dfee74d2362ee5250edf3
z77c429232f603dfaec226810a72cc3cd80c9037c87f28f7c43ca8c6ed6bb6c9df3732dbc7893fa
zf571f1a3bbcc230648bb9ebf08755fea337271b13e33751c826ea587c285f14aae5af55ea59f81
z3cca5b1c245967f73936a86dd84124411aadfb98b58911de2a6378c722e082b7dd823d189123f9
zc4528001adfa92a6e8dd7aadbce3612efb5ef82cc92da253bf3fbd25361741f04cc3af8724094e
z8532479c2d6d01295ab3145f648057c8d3084e89d35faf2b8cb0b17e9bbb650166a090c42cd9aa
za01f092cf058d6f13d8a8b63c026b8e3c6e1eed27d544bca68fb5f8ab73ff667220154f4e5e0f4
z17dc93bad166713f5b5edc0e57c2534756d3e8eff4554ee8bec8abdc2c7b668598139160257702
z7a54b57e443f3e256011e8ac467d03a916e6a2f02319a8e3b3a437cf1d4415036c463dd829e8fd
z62e1732a82297665b44000680f0d1d520783977a5682feb60c6a6097b399526faccec140a06cde
zd670ef27669a0699f9fa186cb9f03afbba8f665cc6b6d6e14c88bb71a118b43a5d011f21aca359
z4c8fe1706264e23b2a6c6a375e69572dc58640baec7c600af4750130ee5fbf6e4ab452959d9039
z90576cbe42c07f1bb9a69e631874ddfe97bce5565166614abf2ba8b881c4d0e41226c97434581d
zf5b2d990a95cd1a47320464754bbc47a097375a24e1d87d5b48ff6e960339269bdf4a2b800cc72
z126de3def75947bb720ee32dd62d07d6a418d378a1d6c8f3edea9564a415358acba4362de6d1ca
za4ade6604b0a70c0dbdf54c99650aa41a71a5ee21a064b0bb6b78f9df2354f4a6d412ece10f538
z28254abed3f194fb036ef53bfc04ee4ad70b4976e320f957dc55e14b333fe8103d0dc170aafeb4
zf1c8c8cd2a1c65b36be32e1d8327f3d23fd361b7361ac62806c2547ae130068a6e7bfaebdd5439
z447f779d4ac511e5deae0833d175cf223649fb44005dc21aea84dc3f91d4ea8ffff802ecee8989
z330a6812b51f8f1da965a126ba00ef732a7622f718633ee65478d1d28656de6cfb528bbdfbb861
zc819f93c9a6b7957a20b34f261604dd480d8be7e715e323fc43aa833da1abe53bef3a0e03034c4
zba2870eab09ad06a17264ebb3fb087cbf3db0129e5768ff58ae736867203738ff9c1256a4b1155
z544895b00d798def92ba90eba028af4218dfbfa8f883620f903a5412340bab68b9224be3507041
z3f45dd4603b4c40e4a8a0a5f36a43476275d0ca50cd8f8896e76fdc56a3c36c3e184acd54c9206
z914297c96f44440c517a1cb7c9344cc79fda93da19a31a4aeb252d12c6b5d23ab935801dbd049d
zdd38e6fde4531b7edeb8420bb20fba8f7817ab0d77fef0d363d7b883024bf48fd6a99003f2a0c7
zc33fb0adaf63de619f5ae53c2ef7737d8687f07708fcca6b571396a82f74bab667bd3b898d87f6
zf29f3997686a59f8e80177fb44d33ac3960318c22b1f58783cc25f470d52632ab001bafb396f72
zd4d1e14cd6d8eb3a94f7ac587207a4e1609e4f63a2971907cf389cf081ec6f4e719f17dba29b7e
z25a5247e8ae3a43f2a2c09f0fefbc349fc2922f9f7b4dfac657453b6f7625f3082e93bff290b2c
zfc486012c01bf81a1f293b38909218d480a33a00144247328ea76ecb875799504b25e55bca55bd
zf6e16f1855d2baeb95ce09a1d93a071ae6131479f2063f4b921a0913089cc3bd7a318f4d6c940b
zb47223d694d447327545f0e6014ca15b09a17e68749d67a0cbcc7cbd10a791d583f2d454c92b4c
z79bdfcd469efd1228969a32be9ebea376f8010c1366dfeb9bfb39638659c931d2d233d2c7cb604
z3245500434696820486270fb909bdde1a12e097ce104e7d5cfda425c998ac9de103bc22e4246d1
z00011390bdae9f2de5f15d492723fe1a0fdd2a67a78fcfd6ae0e01515e971afa5074710248b5a9
z6733d2863821d841d33323f0b2089b30e7d6f274968c58a9c424bfcb796714ebb7f0a52a6d3bf8
z9749e13e1bcfbeca44860fd9502968a6ebee3c9d3c00e8588d192af14b9549b0e23a017702b012
z5630a5192e85b9b7ebb90d5a7c2fe328183bee0581e410220c6f13d80a49c6adaa3c9a636ee0a2
zd139497065d3008826902d04c98fdbc2a18707245605bae899295026ee18b232017a45bc401330
z4a075edef0e0dba046dc16cb263969b292106f197d518a27f270e7cfb1d14192587dc784ba9d76
zd1d92ff7206bb396613c57cbcaef4852c2cdac850c1050ff370acba29f2acfd0067dc62974a2e0
zecf3074c5173a71ac8c893563559354090801b8eeb18097648007043ef1ec04332b65d4b0e7faa
z02b870c2ce34213d22004f94fa9e9adfccd25117d198dfc34bc164951f7510f14f88a0571d6fe1
ze70f58b907444bccd816c0ef573d474e5506338b623f7fe420ba992b2d8e9f8d512631c8f7d7dc
zf35258c439295b32b8f951c1a804cc28acc85fc2bac2e25d6a78a6b1b6a65a87b4b1db9aaeb8d3
za796fdbe69bd435d5270fb8cfe93d3bb3350259c894229b337d94b936dcfbfcaeb3ccba088aa6b
z64a158d6f862052f5f2d1b20de11fbdac85f42c5cedfe8fedfbdef271533e9f4e7877ed7d75fbb
z93c6f3421e966ee26f5f6b31e037d272f12bf3655bd7f3262491122d566aff874e7e339a2b77d1
zeb39ecb065f9354be6fb5790ca76f5b287c76dc0439a850f8d2b5ba80a6e676b9dfe8e8d7b207c
z2894a04fc40c59efbaeade54ea2548631125b4697001c7811371293d275b274164c10525d2003d
z66226ec783eabf5868b5a4c0ecb9645fa731cfe20f58373ed845bea34d25b0bf1a2593d374c40a
zbc863999318cadd34ed2de298fb155b8307bdf36bb7704120d66b360aaae352cbb69a638bf915f
zade87d445f09ad98a0703dee4b7ce6e7213cc9779c47a384fd0fd9d3f581aa13db1fa861c8b964
z7064d962bf456490bc13ebc59383635b1e92203babe810ceb0b477c8672e05fb539c5f0f76bd5e
z749a550cd0a5c8e14b40e64b62060b35676ec7208e2fe2cc386ca92c2f9bccee20d5d74070b579
zb698715e89c59d4bdf762572878eb71dc2c24fb8e42cfce7fa6172af7e48f3e45260bfc3eee231
z7a87a96be8dffa87f6dc7023398050b241786d6a0c40593335ca13eadc4ba2568a7761ee085eb6
z5b76d666da2f873998cd7a1098c4ff7ba519770210bca4bd30e92e366cf6cb6c9a26f0108f03dc
zd98134e7587431089a2b99ec9cac237410e71e3232003280100a320e5541b980f75212e5eb6fc2
z23665db6a8deff0ffdfdf5ecd81594928cc756c23565b2350fb0313d2a82f85f4e13925560dbb9
zfe4dc134560391c1dbfd40f246273a93ffc89f324d37c0d8e35380c51ab25d8fd4c6ba3ff217dd
za788f164c234c2affd31afca474928939e77a905797e239f5b813c3cb296c86a54fde7f512d59a
z2619f362698c4478c6c2b88f1358e409192709a1461053bd221c9837a5d49949c0fd90fe19e98e
z7407ac86128f190e932eb194b3b045ae9eeff7e0a11ec6914075cfdb33bdc6a36d82ee90164eee
za47b44f8e0cb0053eb212dad6d49664aa5185cb4792b6e80bbab3fb99e755b20c2b7a728c68667
zc01f015fd26ed4dc21f3189b92ae54634cc33e19c91b66f7cea907438e3b6932cbc52e829ff656
z29b4517f53447a2222e1076e40ad0dea1a87c258e857fddae27bcbaba1caaac97eae9ce6e116a2
z28520447e908ee54e0f35fecda5202c932be0ccf72aee53ef5b3fcbc8b4207a4fda0354d34eebe
zf19d64f6a1f3a90c672e0c06d4fff96667504b7b8a54445375ce48eaf3017face015c7ac4e3226
zeff5a6f233b51641bc463087376668ea598f0189e3ce6133d26c5a45192aa52cab3c50b6822ac9
zffd882d4a8cec2d8167ac1b6073f85e748d9731a59134d6ceae6797c8fb1df7521c5e53c5eb068
z027003a28f04fb48630108ef6a79e6ce1da3c763694f97532c0e68dbe350614f6bb0df2e5aabea
zf9416e5deb3b3add4d9c69d40eeae0b7dbf3a095b8bc5ff5ed30560a973f43133f8377c2fe4373
z5f5879cd8ccbb0ea6da8a74fb196668be0b132da85701bb22f28a1ccc204147dd218c2da526251
zee7a68e87db767858e1d23f539d9a1e2882646842a995d83370868908479bfd4248c41782179db
z34ff129a43b4f8749bebfbf4536f3c247ea2ee781fc068633653a99d16a6a7e9051f3cdfe9bc7a
zad4b26f74a8852a4a5c130b7685eca21e8386d5acfb7e6c9612324b24316ee20a4fec6f4449c47
z5f8fbdda01c3be153763f2df52ef88e7db623ab4bf5867e73c6f985e89720c2e595e4e5b3cf862
z944fa8e17a3fdcb3b270a95271c5aa3402bf637cb302930ec88f35069795cb096fed3c60e31113
z6f7eb78d30a280062ff3418513321ac7738ac225e1a768595c8bba7bc0e1c6f015821844ca9aab
z2650a845ae84b84cc54a3685107af518ee8d0b1f89ef70ac1cec11f9c778b9a84478af5f65bee8
z88fbde561498a12f092b3bb73cf5c4d972b379a11621eb4bd3dacf609a773973977e27037aa377
z5681e20cfe999cf66ff564e4aaa1c21eb60155898e2e4b1ac0de1f47c4b2df232962614e4d92a9
zd957d22a787d578446ff2196ba4330d55173333f221ea98e179ad0105d510d504a26fd37ed4440
z8b38e967ff810ea6556dfcb178345ed17ffbf6ed4c16d0d8e23c3485bececc089c73128f59b889
ze9ad5b9c0534b3ebeb69b3f333946f50ff8d6ae9c3af93138d1ed5acec90c83551a65d343d3371
za85478d53c37d45cc53a54aa55e8cba7f9d55cc112d3bbf57915744bef614320aea13547494d18
z4a742106e0ab27517690c15f84f5c4699be59bbd7b2b9255de3ec8c530d484094e800745077277
za52a2af45162a1da3ebfefc50fb8850217e11984836277c45d70ca63c91f89a51afab938262e24
z900247a6120601efc1b2f6a533c9b79a160bcb0e3c3dbca3de4baa75b24e9c00cf3ac2b8ce0b7f
z4111f4d600bde05cdda7e331508e706e7053d83d8dae989b66489c1c0a2e65fd7e18cd9c233f8c
z27d4dcec5ec62b91390757dc17d6f4e5322c01184479326c55e086e86193a38479b65f058556d9
z997512112eff7a7a99900a5c48a41087519647a1513cbe09db53410713f0cfa3acbccb6bc57057
zcb1c41cd8a95ca23ce07d3f61839f5a35804eca0245a033aabf761cd7aab3c2b9879d66fdfcfe2
z297bb2707fa492ff6f2a9096532a258ffd4ba0c812e3dd223c1ca855b9e06d31bac3a602489568
zb2c7b635d73a159645cf8c516fcd70912cb333f203708a02cf6e83ceb0fb12a32df0e093eafd12
zfb4963974f5f8a38e141785ca9054358cefe81e5ed06bd4303fba04d53e72613319a35a8f19515
z0399c33eb5a4271b375b071f74bd1d0be65b3dfafa18d8946a3b217e43bc47227f0bfd1f9a9afc
zac0fde9636029932af61d31159937d8a7f4adc4b0d0318d8e47ce8c9ab32107c06eea2172b798e
z813cb465ca47549007166550fff5c186c00593238dbf762aa9afee77a96c81fa0d808d987ff772
z04930c20f70b91970780bf9255e907314fff0ce02dcd5a53f4eb30940cfe9cbd5e2fd4ef539adf
z5d7a541588db4227b2e1e3146b21f768dd57533baaed75b5b8956da92f7c0b6bc28e2692f9fb54
z189191005f17ca933649670cff7b2772f92b999eec4f4b891a0b414b25dcde18adf62365da12b8
z97459ff555970a4e9bfaecaecc17f7aaec3d0fa5b48788e04288bc66ad86e142fee31b37358b22
zeb75f1d944f67f541b34fc197596994078884ce7ff02500b9f10920e0d66f39ecddaeee4bf1ac3
z63315f89b9bfd0f8b470d500e66c845a57ac41069aed70bf56cd4fcc5b64112d360d2c566854e9
zc3ced34dee0d56a486042f8641d05ed0d0c58781dcde2a7b6a19d0d17ca312b67edd33304e1eac
z5280616267804f77c1d0d571b6594546170beab9b29c10d9421c8ddfffc847db0ee5149319bb9d
zfbf64ae3688cc558e858b370ffd8094ffe55a5b41568661ae66ac0ef6d738faea9741b7b2eb51a
zd6e7fe36e7452f5c9416f61e8add75d1395e4700d0019cc69b0c5c9c2aa7410f7aa91e8c6b3839
zf9ccd96904175d9b49bde06de6bc89fc67200d82a68532b752884b16627d2281f20eddac5aa5a6
zbb3051bc768d35b44e399d9836553fe64a13f2d6986fb4a81f21b58dc5e42309f71acf39a41b8c
z51cf9d44662da2c422fc63ee2e34db4a75d3cb410ae9a9aa1b4dce79a952d2962d6631141757b0
zbb12d67cc1db39d6842621086b61c25d554275f7c763014585d5929c89a50bb61495ed4d168df8
z537e83fc01e96897474e6779ff598bf509c5fcc38765f1b297f4cfdbb0a8edde34e2a53c5a5c37
zd07aa4e0fd2f5c618be6dc37a62926f772b3eafde844a6ca16fdfcb8b489fe7bfffff7b6931544
z3f7c2ceab7d1aed53ed031583138d0f04a7c62a78304850744d4a4a0d3b9da5aabb79534a03afb
zac06074181ef66b6b9b82b4b349f9fec3fb968e01201e473b5bfbf412ad779616efdd9a22f061b
za3914d7ea64351bba6f2362200d6bf077184422ecd8abbda1a4861245d59130e1550fa88cce9f6
z165e3e2a35cdda60c88e498dfa676a37c8f8caaf17524de66550aa5c6b6a33ee4ae54f7673e1f0
z545dac46af638ed9147cbd051326b5189427e04b2c96b04c9014e21f8c9586cc9fb2b30012764b
zc9bfdafbf4742413d75add6699b59ccd8399885f935e46e7ef11299bd6f07c768ac6a8b930d502
z23654b791ec7b19eefa7d0b7c0ece01355f46abf779660f42a897e49ed1951b6d945730d028b44
z3e858b1256833a710b2ab40d8bb9e4166eccf97b9988ade768635a2e8d068a3558f31156c66aa1
z9a0f3aebe392609361432aee1c832cce7929e6d4d7809d313df2df7970a3d7a8d193f63b9fe741
z5a9cebfcbd43ee3ebeea38ba836c156c422f55d806e51a8b1de25609c729d759f321c20d2d1c65
z0a8f84565263c7f388064bca4ac5a1f3b5158be1f7b31cc5541c770699cc3c5cc5ea689f244dc6
z31d0af54ef13435707c57120ccc2110f82db5ea53ba5777bee6f0a1315c7e0951b1abc4454e206
zd271cc28e4f6a6c7cbf08e64f348a84fe1a3d48c07d97cbea1aebd6de33548cadfcc211160e2b3
z2325d791ed5b47b64aa0a2d379a8e19f9b953d4d8bed790b301f3ea2d7835c8b6448e5237e5f22
zc06905653bb69332695ae804358750c57142f9304ffb6a056f06ee05ce101e397841c58d7339e9
z1bb7e81034352fadd15ef0cf320adfcea37dfd968cbdbf33830c37f94aa7d88c3b647154b9c751
zdd1a6919e9edb05975ac5d968da98634098067c7d1888e524f7ad9354a8666a949c56a6d2e39d2
z8fb62219336a0fbd02cd29e7641f0968bba52cc040dcc3b62ec0d9a4fd9c2bb15e3729805532bf
z9ab32c0349d696c0d56a1e8e48cd6836a5f4b858f0fd17212966f493eef0a8662787e7a2382405
zb44173d0a47d52a9e772a8216136e8f2adf0b29e30e35d9aa0959d54a8740ef5d697feeda7ead5
z98d378657ec986a57e968d24f1fa0936cf8cf2988b68497c534ff8a9cfa00c5377fe9a700e43db
zce485df201f0b15cdfe86613bb5d44326a9b77f4624055a96c6ef0a43a5651b5071cac536ad556
zbe7cb680c887b6b88bc66f4f898a72cc0cdcc1e6a07e2584df50d19d8197caead05d4995e9b24c
z9b616e5f0df327f6484b05e937b3b9cbc341d8226e2b98190f3703c6eca89825084bd865214582
ze6760dca680e114992246b0ce05429b875eb7b8ed789d67725a1e66844a16ea1834192d1836dc5
z2e84f2dfd16572e6f1511894f8ea524b3c4301c20ab83424f298bf1da298e7cf4b57ff17280287
zf3887191f7705c17b12bd9e08e4886822c756ea164385ab0f53f827d2a7e10ba5d273021a1d0c4
zaee26841b87bf81f230da515cc20ee3ca460cba964658896eba0650b5fc78d5f9ccdcd595c84b8
zf9c5b6ec38dea273edeeec3078937c0d4dd7b312899691ecbd15e7f86cb5258c9b7a6c066f7740
z2f0447e8b9032ab3cc57e130c452b46b744a0d65450d63100558ba96acf0f153174eca5696886f
z129caed2c8e7c4280bc7b847930f6d2a0f1f01f37e1a12d703bde84cde8c58193ecc35defd2a11
z83cbe5705368bb5683a4c816564c5fd7639ce545b8e1998e7d5c4d8300c3b08395ddbcbace0c84
z8634581db3e08a84f4801eb5a9cbe11af92cb26bf1b4ebe7d57677ff4211ad912ceb22ab354165
zb46b95c1719c09551b70e83c8608f12e11f7cc892aa00e1beceba6b21a6ec0bd529da270716748
za064a7d04d16480936df2eed6393b6a533e74ceb3ca1d12a5792248945a8cd2cd1c990f36c097f
z7ae8f5004cc2afd72ce364475a4361d57713571c6b4d4681b1893c2492fe5e1a1d6c6858d1e641
ze3bebe3fee8d007bdf6631f388e657cabf87a3e750b8f3966460e106687049922bd55f87af4008
za654cf3e025a24a21686fe83a86a7e3ca4284f89627101f5a911a5fa73067843b67c611c92ec50
z63171b2148f69eb60c950cb1c8b5be2b2ab11401ebf0d52313faa37c42d5c9e5de1a1f1ecde2b3
z742e8c81d25caa34974bf2dd9ad7907efab6d1a4a168c5a001d29cbe48380050fab518a1a0997c
zc1f2f961906747671961a2ccb6f93f54c457efdd54ef7e1574ca603c2938f2c621acf93ac83131
z647b43961f4ce40f7a4f4ee2bae8699c44fb96bc2c69d9a92fc96845460b502aeb55acb1c3e5b5
ze4c48e81cac174c28ac510b89e2e4f78d2dbc54dff04059f482f83dbf263a6d685388d211fa152
z3d4777e08f1d7f76a79d1f6c5724413e14abfb92b67dea42563d7f8a28fe9a8a8bf58c4fe82fa0
z6610424ac438aad2f4ee9450dfbfaecce2cadddcd7fd6d876d060aa53fa167f8c81eb9abaf5d0c
z61c0920bbcb5d52a1e94dc8c4f094a82aa9f829786a29e324e59430f2d92bf1c358b959bf4dad1
z1f637587448421faa4625694cef10b5c8d41f26e237e39132d4e5ae27c29b37a78d5d464735c4f
zbfecf212f400b0dbd4767be838a87bfecf4592b28c561dcb072f4fc650168d84fb89ceeb641425
zbb9f02d0302e8478c742baead9262988faeee069f6068951777015682e9c468836a7dd2b4cb74e
z9f20ed425e6964a778adf8e653e2c6948110b47102081e34cf596e82294059c92d46a0a3d300ef
z77636e4cb1588cc4eb340179982c9423526b64ef09389de21620642ec575eadff70fcc2e8615fd
z4ecbdbca40576878b052342f97c980699cd142f6af7548394eea390a88e6d7da62bb695379122a
z4a8c891833fffbdfeab1e7140c8eff5870e2207e1c98d06335b66a91f256f2bd644b1063aa31db
zf21292a1848b952e8494b3f8c289ecab16e0df9e4e5e233965c9c107f0cc15c6023f1cf0b4dd60
z8368943e4f8563b678dfdea2040c55831f5fbfdea85fd832ee328afb8afd652fc3b88f8599da52
zc6ac6c70550fd3a43043c354560b35f33aa12baeba3dd12c83b5ecd9cd38ffa008aa37bccc5fc9
z81059261c1907628dce9d0e84e65cadbc30eb43cbfbd9b6616f5dbdd4f58e381ffefac5eae570c
zee7bb0eaa6d7dd9882143aa2381a81791d08932397378511a5cd8a9c580e177a13ff916f5f5939
z8e619624833cc923cd13941743c89edb80e74a4aea344ee099475a4b1c6ce125b418fb96b0773a
zf20e02c0a747bca7ed628b628ec681f1935e4e694b729e4e398abb627063af7667cf27cef56f3d
zbf9bab9d3c8d589cb1a33ee1442082a62b5ddb35ccb0833259cf6e6937cb595cf5286e55162630
zcbd8cae9d630987880f58bd7055e802dbe1de6c380b3665d6cb7d4e90c8904edca87d1efe5daef
za21dd8140536c0576bb9cf8d4b6195adbc29c80a371fc12945e4126f3c44ca9a8636a2b166f1de
zdef33bcf141a914f53754d2286bf73ca12986c4876f6c1f33495706d129d5fb469fd4073dfc5ac
z04349162ba2bff4bf203e5a1fe6ee434801e475cedc8c0bb6f23b9c48315fa63719ea6ff1974bc
z936c597f1143c92b50fe1814fbe3e7d023c36fa3f5c72e3e7c4dfc760ffd93b110027c07be0b22
z10ad1b4ec8f68f2351cd7b57073c48226e11f1c010ef997a9610490abb7138dde1c94373eb257f
z233b24dc4d9765710a0dc5b204b99cbace5eec0809737642b0fd30091bbb1b9a90204ff96d5d16
za9c14aba1946e1b49c2e3790b8810346b4c942d76b16421e1e3e412469fe2abc0a0a0817f73c34
zc9ed92d343c2371a587f398efc6134d3fe3b239882d4ba3a41bbde8aba621657ad087f3476eb99
z4e90ac49e42da16f69a5da2fd29b19b44f94485ccf23f4592bc349fc31a6cd7ddd688c14cd77a2
zea01857baba6c6c154754d8ddaa68edab12902d9b3ee143ec0c3b54da34f66ada909f7b39bee56
z9d1e18b78842f973a8b7d6059574328f9420ddd8b72c781468a6904f8cc2aa62e2b3b04ea7724e
z11448ad96035c7be9a5d2cb1c746bb80c65114f940169b7586f5a13f1479d85f6add1f1803c232
zc31f1ecc01d829069d9c12191640ab3b9728ad913eb14905bb062d9b4b126c5beab83189b8a386
zb3141c89240ed8e2199250f8e17c3edc16f93d10d69663e76e5f2623335a0bb6b130b577948de2
za6f295dd05c63dd8e4dbacedd35420cb250f2947dc08a21af4cb6cae85c543fe6ee0bdeebaa4c1
zd056f2f44a9aae6844221b66970d8b155c65a1ffb0df1132925627248e48c2b25130e64b63e392
za46dab56a8083051a93fc37ef5a63fc7e6968121fcfc889a995ad47cee1c0269c99a4eab83d068
z05fe11fa39277dfce10550d410f46754876149b66288db669509806dc4f475694c23056c07fd3e
z12e2a968ad41458bf48dbed330e5df442e48e67f50a731725d9fbb87c9f4102e90775f8bd03274
zbc3fa230f0dac448083e2b702cd9549c9fd6b55157ed50746453fb09ca63a7155882770d58cd19
za964de8606a4d3b715a79c831075a34b11db008fee6ff753e126fc044d9b3e107aadebf4f40c5d
z167827a70c6a208a5309a519bf1799b82ef846f5cdd893248a78c703c3f5cffed1e36beb7a31cf
z1cea06e24e2e52ad838cc6ad7328b4b49e6b062de37a1b7ea611c048218a63acf52143f73c6224
z67fcc857c9af7f225807ae6de86c01f99f2183b16fd6ccb4340a0a3c28ea1ffbec8573e89c0bbb
zdbb0881cf3c3afc415b3ee8a332051817ff636b290e20b04be168c9cadc2ddf79d5b8feb26f71a
zcea43cac30b443240177e8aff80ba2d902ffc72ca5c628ce5ec60ffb2f2edde5b3f241a2fdb36c
zffc71120efdade13fb891ba9249c1901fe6a5d3f216ff185fb19fd329f009dd5efe2e21644c3e9
z168bb47299cffec111942a2e2f87d28d16f3b6e42f5f9eb6a5596daff430afb14a0c509b432e62
z5ab7c786d638caad9cefc5259ea2b0bda025ebe8c06fe86fc8fa257ab33152381964030731cc24
z892d2cffdd8cd9b54c8f138f733cce148d4665f8ecfde5753424ded65332e4680070b43cec3e72
z3724b8521c59282423121842a25cbebdb25dd6578f4175ffff75e371dd92a1e45d2440427db6c6
z5f244cc5686032852222308e9855877a5e718c5331310af1a682bf1a21ec4c662960de63eeee1f
z9242e1339ae974d07de9dd440da417325e6c253115c9760a694778a5e97ad25a168f6d43320954
zf00ca27fbe73f1e79d89ad4605a32bbd609da397d85f9296264fde665db162ac9dba0b79f2d5c0
za8f0341cde23c7d4a10eebf53b07641b6c4dec3c3ee1ee4ad3d1f33bb4f6b22831d1dfc5c9c275
zb789408b0d61e1b01b175793f8b28d4f1b3461e12c2021914eee9bda1e07e880042794be1f4c13
z3d0fc6fa7ed67e68843fee10506ff0cd973b11e1bdace4426fc6b4e9856a7bdf59867a52d883df
zbaa09d2d2155e3c3b62adeb1f1ef2db59fe3f93e6f0ab50535cf492161120f2cfffdb61ee18a10
z086aa1817635f9ba9cc11f4ea9a4cc224f4caea5a8e98adc01af5e066ee2da01fc3a9bf54eb700
zd8e7f1660036471f452966413f0b15186ea5884a2a82d3becc1b8747be81011a4572a716e4150f
zfb05b1086c6a4a76a4a1e773633ed1aa67eab51e6ba704fea4ecd92bc693d2abae75997602778d
ze70a2644290cdeb6d1fadb3f66d4edec2703cb3828d736862aa651a4df7f9539140fda0bc27230
zb280544f1500d01b4eeb1ed7aabed91f034b3afb37cd81ad9d9529c3acdca6f37b61fe2ec9f3ab
z423da66c39f1eb521a96350ee8bece27d0f269faa6875925b56b99b34d249e633d7f270f781323
z88bfa7cf6ec7fff2ef9589de57e14c04d05ee9437d0ef0f0c0004dfd036c4d7b4ed39a808776ea
z4c59b1f42be29a4d439595111751d3c23aa3ccc6c56ba8aa2f0d224d41f66c96f8303c0b3c5c30
zc1d681e9f2acd80f4f628344c456c63ef4c0cf1f8cb5ceda877ed8d41b8c4e9eaba8b951894989
z503a5337c78faefacf6c5d905367bb3ae7551b8681a51d0343cd49be4a993b29ebd3b748009c32
zf5c541f5c3c3430af76e0e586686434bc441d5fb1ec75bd7cda7cb26a7f061a5c8616953bb4e78
z8fd8bc8a56e033ea63108066b0ac09f4044f14de4458c37f4f863db400e89c5c8009211c770d1b
z444b51122fabc256f8b8c0d014faf347edeadde8d309e5b6815e175f1ad8479d90735967c2de85
za14b9446536e2d961b48d3fb2c12e7e4f22c70ffa3ad7354d4ad76e4c7bce404f0745ef92983dd
z145f61ad652a3543f70a7b1e1798bb9fc827ce8e1a8810ed03dd6ddc2abe5513bed2dbd15c6fa5
z7c23e1eda5e2f231e587e316062ffaf626a3cae77a1f0f028e5d3e98c28c59e1dacd74ac7b2384
z656b169edd714c31f816dc7dbd0a930c62ee4abf19581b8c3488ed07874d7e2313e4ca52259806
z54d32c28ede6f0faa4fceb48577a0ccbf26e934e38ffc31e649b211bf6c102c9cb5bdc183c7250
z99cf8eca895eb8790dd5a820db8a94cf76be8e13d45e03b725f43b3ee7c0944db03ee0f00de28f
z4f1a64fce2359b5db71471322ce87e7b5fe144c25018ecb2dc9b06493c6b4638fa57b30b5665a2
zce15dcb7b71eb3a0ae08f9dd0083279363fa58412459eca803d15d6eb7fa6a21f903b87432ec1d
zeca43482df53fb55245552b2dd9cdea02d14d1af2d5884a21e39b509e3ae26d986b1ffd24542f3
z54de9d931946c0ef186820972964a9e5fce506859bbde690e7128aff97346219bdd09c15292187
z936bf0b4215b95260e5c00a8e49bd18894f86d70b1a18ee7022feec964b1a2d692936549513b78
z786b7130928d9dffec5cb28f0882d131e5e8a2d61dc8c46cd0d60d9d2f7a5e1e22f39d1d690d48
z536b92144ff098bd76b72b71399cebb68d370c70c08e7e9777733ba237dc5b8423b784dc9c2cc7
z6d29022a08332857b8960a8691324147739da9ad4ff6a95fbee7e7ddcbb8efe9f421c82a82d04e
zbc8296793ede22363a6676d1b7e357d8ba5d449363c92494537789e7ca078f571b0538b563ee85
z4bbd1624adc9b4cefe7a794c85c1253e450eb1ba9805d687843668b766d0fe906351daf275f210
z39c71605b39d78d883b7ee6bbf4ca23c54872cde1f1a5e1dee5b7cdec204d6138a6daabb234b78
z24786f5850c4428c6c8bd34c82004dda8ec50f5d01f7514ec21272ee5a49fa788a0cb9e50f8f7b
z4866e728c5eead74ef362f4e5c6a42e6603ff5c447b231d74c131efce21086134ae0d0b3227f8d
z5208c2e36f11c5f89e5f0277b148c3365cd04af43ad6dbfbeaf234bac85e9b1a39fff032aa077f
z805fe731ba2225642f4124d0e18712e9013bb42dada86e83f2e7ec807629f878710898585ec3c4
z8670bfdf6c9cac6e9b785f2ca96f282447fa66bd095cfef4d48858b53cd1830a512bc5ed48b0fb
z40c21e1bb5b5cf9ec7940c5a24903664f1edd541e2dfaa136e0a364962a51cbde3222a82c97b6a
za4d3661527c9edfad08f76c8f5257d34f0e265689da8b526fc5e9b16f891e3728845b537d3fae7
z275c8ba584bcaa51633050a8c1c0dda61c3b2c90e61ccf7e98bfbc43d623b622b3d47d74935a2e
zbe9523db9d4d555c5f6ec2380afebd46050d3984d40d6e93124010aa5bbe5c3dfa6592bd63f1d5
za31db750131fa1e01ada3425df7c6f7c793d5157624478e54d219dfe3ab84dbfacb1d47b1729b6
z8b4285e39f6d5d9a5729f071a8248f3de7cc16a62d22a536de81102d3b1830842b61d47558f3bc
z39b0ec80238ac5b3a64a9654b6a4907240efceb7705bf4764ff3878313430bb6c426d133dfca93
zf30733da13c6bbebab655337224550af7222d36de1ca0ca584327d158efc0cdc4941dab00d53f2
z2adfc91f38d00c5921e624b7ed3556e583cdd3f29be56c1ddaab5eb3983f9c0ec9be6f1ebdedfb
z3e22b9feb2d884e4a5245927f776aeba363b9497840cccd7e7f17cec9ce20ba9227d0d48d9abcc
z5cd6fa5194056a91437133f2e41f1b623ee3d698266e54a28de8a74fb4b3b1d19e0e7fa4c90bd7
z2796ad79a8e60f2297c83fabc1fe9a0ee3d798d027bda91f953d6670e736dda5c83c15b50d6b05
zfd8e58f36c147a98a6d7e63b7fb860e7cdba82f4c0fe97c301ae08aa3be5bea1c498fc6b882a88
ze1660cb3ce0c8d7c8913647dda8c78245f91ab3059c50cf6274b040ddd4bddd49b241f93a8ded2
z674b6690a2905986646a58d5b1ab7247c76be9f27b77c2c0fe3589dc422bee60d09104249c3176
z2528da42106fc5f69346a0b5d4f7eff7ec2f4333d36925a957eb3e9a84f8847cf53119ec9842ed
z646eb27ef1d4abd74afe8dcd4bd57f8685a5e1d82721eec3f1a43bb136805a7b76c79a43d92f59
z95bf76f0c08ab3bdb424a46925668d34bc4d9534154add1b2d8074acd649f7253713332bec5713
zf098496c713c8525b55254b975832bc0fc3fad1a65068d79f5bd703794e4bf671d694b69d5eea7
z95e93b82ef6966340c14dbd8c4804649d322e46aa1af35978b54e001ce7cfc47aee73327517026
ze86c1bd6218f473f0772f512d0210e55789dd7ee66f6bf35be68c1def0c1974fb011983069a2de
z3296c79dbc4c6451fac9a0b614bc08cae12654f7166c103bc9b163147b213f3ea053647ab676c4
zdcb56f279a5087f072ba3701047bdaebc1c42386f62ef7e84ca833de0861bf29cae89c57b39899
zda2e9f913f5a22bd07f62b540e5200a76ee25e837b1882e8f07f3c412e71e0554c4036a25b8f02
z22816b14240d31fb5a24ce37993511c61c0ac7434595bfe8f89c6da8fb25c10894d2d8a0e5d851
z825b1b81f040281dfe206317b56a0899826ce0873bf5edb0e1decc17c14691e61d6ca5599b45e9
z833112bb9ed35b68307c1a0e9e27b5d77d389361fd9ba3025b575f1fd8463090a13af3ce51ab7b
z075310c26722aa8eb0897f002978543241ae01c865acc2cc081c52de784abf271a3fdfa96097c7
z3bb8f4e566b98b3cf587a771f1430eab973e110af13a22dfee73e3210463afa1ef8d3cbb50f3d4
zeec65264b6770c07e8ed91352f63850b05171abee4d646810153de2a30778c6c983a11228ba467
zfd0d6bb66196718a7ef991081937937f42aa98540e31596f456c276ad31b4813a3c4103a0cd8a8
z555d39dbd824b8233489003fc7e2c2bc36035672af3aae9c52a55065499f7bf63cc1aa8f90ceb2
ze39cf4c1edac752c6daab8f170f90f45e547b836df55a6937c5cfd774318db1a8c6a3cd9303074
zad9f4a1e4cb216fe8b688af1cb4ce8e7dc1b13e866ffefe0b19838273875d99cc323a092fdbb25
z70a93750de6496217981fa66fe72d6d1644a9306fe7d46fb071d418a1bf660dc2c1230c8aa0e1d
zdce4a740b6e5d37f3bbd315b91c35e702083fe817bd2d2d316cee27f7d09161227d5e519ea05f8
z015bc790ac88a1e3c690b16cf8d1de18ecb0a964e56be2ed1d87cbdce969e4f85b9d0470fbcb01
z2ceb30193bd6ff03ad2f9414aa01ff3605d86f942947190f6b4f8721e9c03baf11fb75363ab387
z5b47827f3b089b3c57a7b35d4a78df70042ccc4813b1c3d488689a3b5cbe79fab58f0569f51f05
z5aa4a8119bed4676514461dd56929cfecc7c056405bddea0b278020998af63dad0601fb08cc65e
zd74006c6a93e9c26a7b8b631f5d190e1e49d8a61c8bd4db6cd0772575f6fd81276936adb5b1099
z29789f8fa10a8d381f380efceb360142b5e8cce2dfc2f3d2f75f2a048a1dc2abb3709fb2fddf6b
zb371841b0addfe040c16694b6e137489305d0063e5d515ff2e988333f3254d54cfa74e03462fe8
ze394d5ca3a387015a64eb46f671788d45a2fb95807739871bca45f30c594787c721cb210fa7593
z1fed059fffd1b063c7863f542dc228c30a542db77dedb81f519a1ada0662b3936913c7a3a09805
zd192a53b3020f88f6afb7e10cbbc2fef8005dd15cc88ccfc1ca908a2450a08a2719ee45ef8039c
z5c2f3055a2f73481279afa8f323a73f2571656b29cc81d069ce0365b3caffccf6a7e95caa9c174
zeb67c0126fa11df2e6b1876c7abb7325fe86ed4113593d5dee48c8c7f5c762b81796394061fb02
z8739e502091f74093381835a4f9422e19c0588ab5833a8c012d857966b7156ac7ec3122d881df6
z2b092c3b57b2c6c5057e7361a4c167544fd485b15423e58d0bc091eb4ac17ad1aab687c937379e
zd4695cb9bb355999f2060146f278a8b703675e599043b3c3fe0423bb16050796d114fa13bffc53
z93a7a1128aea6056e5dabcfbcc068a690ae8096d1c7005ac649fc9ff67fe5e1522068f5edb5d63
z07d20b9008da783292070c6c1499c863c17b7d407121829263b91d12cea17912a9abe68dc6b64b
z7bdc7e3b59a3172eba7ec51f9be5f2b976862697316100b8776a261cac25637868d3bbf37d29fc
z111eaa9d9de5d15ffe0e5ced84a942c3a89bb36d7c94c726255dd7faf85780d86e097e4125a98d
zc1be0b5effda64aa7209b845e879b37ec911453935748b194f53d686ac86dbead233710c81b37e
z90b00865f62d292a633bfa73f35a21f30fa363c217a9c19819bf03891023184c0534e2fa3dd358
zec17b0b5552610b075d466725bbca18196bed1a055dfaba375f6eaba182c0d33cd8e09165e47a6
zb60cb5af540e3e93155dd0061d953c07a828e2c04d7d23dbe7c69c4f3070ed74fb22fdd7f133bc
zb4ddef8a318ca548bd681aac48c94ebbf9b9b4f9231b78f747d4bc36e012ba44b4f8bfdd35e2ff
zf7757b7894c614a2ab28c13368a3379b5f00573e5887d9dbef3c8a299183ae12af13f9c26ecea6
z517b06d86b4fddb4c760d272d702f5d940506162e71b692a9e34a29dd7d49cec0cc75ab16c2791
ze20379ad231e3e533d0aa251d9648f116525655dad12837a83a50ab61a6ec2e22941399ae473a6
z64a430b71532776edfb28369f8d8a1d893079432dc18732b8828b8baec7939179726dd369701ce
z8e9c81f99c0783c6e65101dbc114d2ecf624ff6e4ab11d031a7013b990f1fbd38c0c19502944fb
za35cac9e63cae62dc52d7edf780f3e4e4c52376ecfe842e12907a2db0e38f1ce08c437f8a60b1a
z11b95a881763f6c93a684a551e8fa059de279aafc34b7767fdd98e032b44276d98314397f8f426
z7543e86c79515ac975bb4d9cfc54602c464f1e967902170caa09f6190d2ee807a96b2c14ad8af3
z4f4b57b537508c753a9ff19f20eae21295437738bf25666c8e5ef78b37f256b381020e71bee135
z8604002280d044d14b5d7d1825d1425c6c9d3c4938e62a33f0eb7cffecd2ed363934640a4b5775
z9f3e10d1c4b1456820f11b368800cb53235fb8bc192f4e517bdb344e185128dfa842808aba5c3f
z3dc9b4cd072160be8102a3dde2978ac282efe33d7c4b1cc25b0abacce2e4d1be0ada377897bbd7
zbf7b81f689b5b58c72cf5a3fdc03e51b1cab2b6db95b667d1823c761ebdb0818d2173c3c1d9938
z8ca7836bafcb676884a32b34204ab622348bb81142f6ce799fc62e75c6b877bd95df3662d3e3c9
z6ff38ad9074271d08143a377352a339e72bc19f385c63d67207796e35531327f8e2e4139ee1d5b
zb9b34ee9546676486686de91365200bdcb13e728d77a2edb48614b3bef4209117ffa437865e0d6
z6490d9adc784d99d49191e9d4dfd413f11c13f0e08992bfe1ad1e31c21fd492aef28448fd92afc
zb6eb4bfaeacc277a629f479735f948de975440cb70152235a3dc7a8dde755b1a4dbfe2168ca6cf
z93991ab730cfd7ada6eb2a488ec48651ec0fbdb1391fa88be43333021c161e926c4b7e5838c6bf
zde8fba2977d27481a28199eca04485d9197fcd20a8546925066d1d1bd3601a1b248504ea54a16c
z517c4b6b4f5ee01efdaf3295f2cc0aeeb73f914b8d076e52ad2200ba44ab96f30390dff1fb52ca
zea41cd75d0cb1a38773e4a347817b0974b72807d1d582a3269b90bc517cf28cfc7633ee0b912d9
z47bddfa4a9f10d42f13866be67159de7d5e70183e8d5920a94a9190340ded5077e4e83dd92c61e
ze5793a40d340a8c935fa45a54bd3c898d1823fb086203358be6f770b9982cf4f222a747928e26b
ze0d20ef942b93def9112858b61ce119431af3e304d807da6755fecc1909fa95e145096e4937636
z46559953883e85fc4e863e0cd6d1430f26459e687a970db55673a3360bef9b154d3f0bea06b72e
z9b3d928a19fbb069e0335617a54e958f9259b46c2597628d9db1200eb58ab63522fb4863aa8104
zba18941ed8dea0014e763624f285b8e54d9b15dbca0ce0ed53743fdf263a80e6d8e8dd129d688e
z4eaf5543dcc2e609018e52cf765aee56d9d86d7cef29c00a6677f61cf3799092ef9c942e43ca3e
zf0c4a51fd54b0c85be6fff3bc75054dbf53be2c7511ad714523b56903328cb12c5bd07c3395bbe
zb1c5b921cccaf23c5d49c4719eb01ae13d1e80286fe87364fe451edea761ad317f1198b3697393
zf90c376f238347dc94bc09dd5637f9dd96157bb91c125c706d4abc0a18045d0a9f055a79f67de6
z0a8c380e32dde6f155745a20d82bcac2d60822f00e9b8b81b86bf35f8fb68c1d76d69012cccdaa
z7689376e953ec9043f1e908f598663f5ae1083f4e828f5a5e104d7374970d3eeb0fc97680fdbd6
z60508d80d24e784d71dacd4df54a366843f60c3dffc23b6a179e77be5ad4d24e63aedaf8955b04
ze8c434f2db75f52741f0d282dc15182e6c2f1c2c886677fe76cf421da312a2541bfba0b9dc5f6e
zc4238975b2d89a100df8b13a9cd118b8086a88493e762b593d3f0c5c41be25a1fced8b1a80de58
zf2badf16d562043f83196b36aff62060e7f0e328dff977f1bd08cd40ed0e9d44fdab7bd3b8f530
z0cdee626b5af586346de5268be46f7cfb9eb78b4ca9da162bc0f20ab6058a24574f519e225aa97
ze02d59e72698f366bfb4bd807b26b0a0fcefc25295b77ca1a085119769f0c99773692c566a9230
z83547ef35e0bad794a254b9c9083f63e1bf47a37bb07d3b6dccddd435ac103ae9ec04f4c82fc2e
zcee7d6945c126d8adcea774da0361fd4d158358631806442c9da0149607d685aad0ee06ec2d5c9
z0036aba3a6f7a2f69060929ad81ba7fb4946c0c95d2318d4955e6605b0c7fc54bddff99add7b7b
z0b0a32d176e24cc322f654e9bd4cdf32bc4d35bdf63c4bec1e46da5f4e5ec5c852592a6385f867
z592b5703566f115c160a707e0c4e8637cb485e3145aa355f9740e7a9986a0cced352c7ae7a8cd0
z514d33565e666df8aa9589685185f2ee10738fe028fc86db1ea00deb8d0890726cd91b4fddf9a7
z249915e452505f31bda7c3828b9c848f04498d0cb9ea0b9eafec22bfa736be1cab858319b53cc3
z5c2880d7b5ad51fbde73d69daddcd27f17c08d8e7f4d58c7d0d38ffcac1321d491f9f03577b820
z1b22cc26b33e5541fcf07274ddb56131ea7d37d6a03edf7b9039e470642726403643ce28e872ef
z3fddaa90ed6189cd4838a66ba001b403d02712d8a468a75532f6ff09350af8dc24455038698284
z07cb665ae161644dcac27570413718672a5895130931d3c32c402b3d4991ff46da277ef3b0d7c8
z0a142c291494ba4e3d5af4a44e7665ead49333f86da9b359cc523d7de4c5b7bd86aa626501c6f4
ze2023852e1df130f06b1892cd4ee90b8fcd14ebe1edd8657d834671f3c773da239f6083061e7a4
z992d812fe6bbc8bb5843545fe1086ecd7d27c7d57a971ccfc1fc60c34db3da58a3876c8ef06e55
z7f4a5792902c99bf03e653d9302a22de9d7fbab1fb1f6ab7015079c7e31a275efb37e1f21abcdd
zfc02a5a123c51597867eb891e04320062d645a71007fbc7d66e927ad30a87fef24de67695a34a7
z646398c389b39948b00f62dc827b029bc12a2830da1357036393a011533f995a5792ae948b35fd
z70c5e6176f1e0a3c81461137e3da1ec2b14d8201a2c90fa89b44a5228ee11e585b3cc4706d4dc7
zd2c6f83482881982f462ca3a289e55604b1fa9f0aa16dd75e2df2b7846c35f1f0c9231593f75ac
zda807b4c8c96f68a193cd73ac81bce646b2feb755ca61b9cfc8565f18493166b37500a2c9e8862
zb180aca53ab0f33d725599fe4a732b9ea4a8f43f37b5c6f0bd80d7f4238fe83e42f708a2d5fd6e
zbdef7499bfac94a7e3b8aa22d88762049b89f6afea6b8f8aa6264dfe07da091d84e911bae1533d
z0a85ce6e38b69fc7943fc39b75be5296493505383262b9bd2b05cb7f774f239d46cfbe384bd22f
z5beac66b594ae6bfb51347b3daafeedf818caa98024b3438dcfa5b29aabda88fed5767b773b433
zd311590ce48716e4b83c875c28952fc084dbe9ddca7f31a3c5ead07da182b731a142b19d2c7e60
z8061c1bfe1759e291d425cbce3efab8bf831347e569678e343887ca34e6a7d2e6172d7c04303a2
z7c3b033966033a21cb7c8c7321357ed70cd0f1321d2f1131f89855cba5ef4c1ec397fc810d7dea
ze9d7b7bea09eecf84029681a08afcdcfae834c4b8d9d21ee9a4bc75d2de17ef3fd3b5122700a1e
z2c49db8c3babbacc0baf180287a02f56b80f80451bf353e0aa951a5a0c9370eeb30a7868cebbd4
z3208614893b351204773fc0ae6d89d26932fb5cdd696bd763f57e14591d786d92730981b411bd0
za1d178049155dfee525dcd5e2c71eca364f38faf8158fcb99ff9f5529501269fba0bdfc86a7ac2
zafb31126ed01954b4cb365571d86af6c14e61d592e2a89e54b943c6c4e0e80640aa6bea1dbb501
zb6ce4ee79efe7253fa4e34400437367fc2ea093fd2aedcb2a1d7f1b0577bbb2f493ff72430a559
z4098e19f73bea84bb95d594ca883c88e5777a131d8777ed395b8f46bf7cae9c6d048705dca8baa
zdc794d3c43331b5d4fe86ebb904fce7d6af08cf639e45327aa90265d36073b13fcf5d3b41e2b0c
za02f3d3d94306b7edab74ad6ac9e074aa70eafbeb7bff8ca22caf22cac7f1e78be7b38c9e4cd5c
zf1faed2f86236747c505c48a0d5aa92d1714568843006a3d9ac70e7aba710482648729c7bc8f45
z37643734309f70b0e9c16433e57ac5a7004f7714fb6f194000510149d4577065b1475fe124b6c1
zd53e66e996af32621fe3508b3ea8aa3d74ed0a93af11822259b7f0bcfa8eff4a30e68034dd5f57
z663249380021e81cff3f940acfdb7d0e16422b2c61a57cdd6da6bdbb31cf4ccf61ca9ac79cde9c
zf090efc7aff06358f6ac274a3c6c56d7754cfc85ced8e0dc1525a402ac0fbabd09291cde31a7df
zf7e0bc1264936ec8a2c33ea17dcaaad39fa01b7b751bb31baf4fa0b2dc1da5a6f66cb1817daa8b
z4aecf6c7a5228aec9ab8324f328171b8ad08fba50dfaf12cf57393388cee4b7a42bc73363731da
zcf8b86b045a1bb1394ec50a3b31593f93f37133e03afe4587d89f6e260320c5827409f65fcfdee
z7d83d3d3348423f718cd0b4ada625cccabebba27e507a31bea616e6270f8fee4a77d0a2c822184
zaffa0bb463e73d0cda86c3e5d865aa84a56bb2ef3b4087cd01b8153eb6bf93f3353c0d11d23588
z80bce0401f95bd5b880ef9f684d2efebd41389723acb7721158edb348d5d8ba4756b125f74aa9a
zd1cbe1741d2d4454ca829059b952196b8c06c0f7d658dd8377688acfcf089a0f9ab34091e7b1b7
zc1f77cd60a30df1388ebfa7ceec3ef5bd77e4ec8168ab20f2a31b821278aff0065493246349bb3
z247c8d910f8c069f1e3612e67c1c664517014465c7fffd393552bdf22a6daaff2ca89b68537173
z1eadc5a1464e9090f913f33b887b47b794b93ca43f319917cc796e260f41fbb129f471d7cbed90
z216622637dfa538340486c74e778e26f9e672a7f1588d710d4ee12c0617aaaf7fb582a890e68e7
z266b5c6bbffbf7d04b39e6942ab4da9b55550815fcc9b5e4da482d761db54e992615c624b9d971
z4c9e82763ab75c10d9fe364a5ce5f0d25571f62058cdde42cd75958cfe923043924dc8ef689a86
z040a46a01cf4fbbd435be86dce3e2d1defbe2705031ff204a902884393a504721b5388df66cb94
za596861154bdd751451da724cbae17cab71e8eec8709994945d986811b171d2cd6f09c716c19f5
z4beadadb7c7f062c6f5fdb55000939f93a116b67a1b850e6e7f4d1fe9a503d280e65afa0cc0d66
z8458c84ec56106e35c85aa21e32ef981be2ea25b276316f1655bf8806b8c18b48dd4cd082b96a3
za341afb062d58b0728f3689df6dd157ef046eb7a975e98ff19380a08ef14715078815b32645cd8
z2e5b3f4cae06fc2b50864eb5e39fbecd6fea0cb0e5134985072a3977ea3115091013c2ea36fccb
z69871053c517f2f54139ed487b2a1127ae71c8a47ad921422f651988099b1df4935d6fe6f2763b
z7d11de0f7f99b83edf47cc736f1022ec7fdb91a75865e90a06ea9a8edcd3054ae2bfda8a836898
za4d3cdb2ee37d552e0fff8c4f46e2fcb74098fda013108cdedd306169a4d8291f3035d000fec81
z2ccf0ae65d8b81267bb2af28de949a1b94629fce93734fcc3aa3995d04225f52954f128116add1
z01358cccb525063c1f0b603f44b3f2740e18cc8504126c3a59026511db99cae720c6885516c216
z70ed8a301d90893df6a0a742786ba78c572de71023e9f9d61d07bd606917d395737596bfb682ba
z362c9c23f56d978a19d1eefe877ce75f4103c439577aea9a398f5e96d060466d49117e418da6e0
z5c5e59a9fda993c06e7142ee0bafe720c0bbf26d6d7098473ed0e964648f52a83a1fb92a2e7171
z86c0da0c0f06bc68941f99ed08691b13a47b1d59c5a52451e54ec9b961f0fb2b9afae64aaf2c4d
zb90ff8e872cfd549e4d8c1b3cc6de5229d4712d234785770b4c97fc38255da917f4d4e8e6aa9d5
z6183b44abce0df2bbb11901fb0269878678b4bdeffa6b4eb749aa917dbb45ddc363ba0d244d15b
z7df8d224e53c7b1ddb293c902b51dfc86c0fea51da0f099618d75dae4ea02dfad7edbc6f9ed72e
z3a45ae76262e53c2f32c1ac297ddfee31700d750180a0f08257394e9712649c1293ead5278986d
zc0a95b0e82bf8ec8775f567fddc3e1aaa5343e31888acf4ad914946c08deef0dc14f061951c431
z4b67d36f72d613c6aa3cd96d3ea644e3a85013de02749edb1e9ae8bd885f3f8d3f4ff07ee5ccb9
zeecdaa1244cdbfe38f83f407c887e76ad5e6b5e0044fee45839c708939a04c4c343ab7f05b4f1f
zeaf4ebe72057e9e11934ba5d1e3408a0bb0e450914bd23634a12a9171b320c348876932668b156
zc4556760d3007fee04bf6dbd20188254e2f0a6fdcc68d5469856a8834494b22a66158a4102c603
z341d8c7baff8fb69574cab91400764d7905f2be342bcd650643a4b965958a0838bc4c1d64d8024
za308ead60dc47880fe340e4fa61e7965aad4cd7264ef257a5a860b00ecbf650dc4790907beadec
z959b9d470cbc3b9b181d8c25f85fa7bce66e822e05d54ae620b124304de699ad3168c9233ff32a
z3ba72a4117a999df3be35a18f4c8ccdf974c867b2fb26a2527d530ebff819110020e9f52887c05
z241cd93c19d8fe1cdf5a64129c2a1b5f46c28725d9a66c7c531131a2d4717cd8e5c0828bf39b7e
z1bdd7f9515f90aa5c8e2b622437216f5ae793b19d6abad054a5767d01e40938ff072d7a076567a
zf986be751dee28cf124aa5ad0e28433d28c66105ac62709033ecdd972155634e591e3d82af99b4
zcdd597de3526a22f8b455964850f2018cd64e35f0c409503d3ab5c43fcc3b73eca8e28b9d3c4b6
zfe541f6a12071e44a33fa9e9ca4fa64e45403a3a53abbbb1a3e6b8e430ecb88f9041396a93626a
zac4fcff30ce2253008425dc1f1e40dbba019fc1fa12bfa889e967f5115c338827437f156e53f4d
z72eab0a1e0b10aa4f9ee070f524fba33939f993e15484b27acea12ad625a6652bbffc6be939120
z182a26ac0115d9ba64fdbb916824a9e250db11874bf91bfb0d0851e3eac59b5680fe72ec95d8e3
z65bed2649862f310c8a387f3e529c3d8f0ed2c1afe07dc5b32c16123b67c7cc3ece39bc9ada4a2
zde7054cccf9ac7307403b90a4c1bae21236a47f39c5eea24a1ef61cfd41a1078133799ef20adec
z6865dbdad94b781a3f62455b2d712eb5223187536b84a8e69440464596b2d941e8924e52d85c95
z25b9080091393ae3a15014eb3b1cd932c169517764cc98147c59a90307587e4a63ff2d7a4b853c
z3ff15e36acb44537bc4b803e039c26fb317e596e18239fa66db2c8ec1f1c74332cee5449f78584
z7ae859b40dc598228edc8ee1da0f1b2b2912c9e6c59aff0b88db38db4b544ff08157f8ead353c7
zd1166f863cc604586b594b2604d137784e6875e3867de084591e4aebc6a464bfcec50d95ff0850
z0a91b9cada45cbc74a953f8388f25da04d59e074d640a11da807c92d689be6a431a602260f59f5
z4c9146f183f45f56953e00e420b7b281ab14fa07bec4908e5236621f56298241c99af975a1938b
zc2f9096d3376b78bc907739de34b61e17beaa13c7c43128133e3bcb50e57c650ad224253edc42e
z01502f658c8aeb535f543f107927444b235e7acc7922eaae8897e2fef1b9de68ebe7733a83b8d6
zfff1904abcd6321d41e959dc9899614820fdcfa629ad245e9d080b37c3f49e752f33d857a7a836
z39c5cce45f9d192b3233047aa51ee00fbea9e4d6557a73ebc3eb4322895c783c77cb25fd51f1be
z66406f1bb455e8ffe66030fd5b58bc62ad0540d0575000f6917e67b6b1d6b4ffdae0a82451b7bf
zf9441b0ae311f7f4e616dd8f92bd215eb72ea1941733c12a8bfc50d709c64551ecbb30442b8a45
zf875f108781c132d5e592de10dd271cf952d5d0df8c9c085ae6ec362cbb279892dc402e865df45
zbac0cdcc67df49831014178423468b784008eae2b027cae2433ebdb21008eeb379098d93170fab
z5eca0855a4a6cc639e748fdcf9840e32729f44227e815793394a8606a077733ecd6d910dc8e28e
z391619d09dda5704608334469cefcfdbec90c1efe7bc61f0326bc4181f8994b12928ddea1193c2
z12d9cf75089b637415f9cd2db4b4044f1e7e7c6309986d82605f0f2925426a4b0b8e21e8934fca
zcaf5c0b9b95dc2b836364d4917cedb471530c5223d452c066d949b6f1f57124469080e77097391
ze6caf42c39365fa2df74dfca6c90cd241e493138135e4908c0aca322bd273ccf9ec4d6f844f9ee
z7e7e6f5661ff1f6a4b0cb3d382061024106718561998bde75fc47ebab7c6d7afb5b0c0f24b9fd8
z59453798d3fb7beea9af1c6b5eebcc64e7ff71a1a403be2ab6d1b45d86ec36a603647f7739c800
z8636203646b9213528a744ab7f33cd6cbc09114c96a77a59571722f28aacc3a8b7a52d934fa91c
z51ee8ce0d599a2e7b17611cbea8dbb4b5865946564d1287ad2fb84644b2f41cddca624efa8df26
zeb6116283df295fc1bae7ed32abee92299aa60156427801dabc006ab6cafa7dba88ebaedf21312
z95252fceb78c469d4eb7a822aba6a0c7e0c2253aa017f844c1de60377bf9dfccc207e33a9cc737
z19fdda777dc3930e149d17a95bb39b521adacd7f3dd0753972912a0fba4ea5c31e17a710fb91a0
z6fdcedf5287ee23f112b14bdf00897b4e6e9a63847fda6b1f8d17ddd3f19624fd4a48d005b9a12
zaba375a6dcce5e954b3bf985f12bf1fdbcbb32f23f123b9553ca745c388e0409e8ad9276c460cc
z7f84244a57ae7f604e3a03564d6a2489b104bf06143032482b612a074fe05eec14a5b4f87de99e
z581978397ce1e3e32546471b084b4bdd56c612fd27bf84b38d37e6613068b0aa7e291bf1f322d2
z93b58fa06d933ed48b980841db6f9e9c9e02722913082ae6e72d4e10dd010dca3ff5abd0a8c08d
z54c4546b9b51588a523d85828f5a63840741d3c1757481a12506fc3915e11bf7354648fb2ec1b4
z2b66948920878ca05be985cc58dfc87e13453a9cd151fdf3bca2c71c57304c94c476c1454cb68b
zc3fd7cc07ade25af3eab17f27e8beeede98627814f36c74fbca51e1066fdea511ea8d01e93f87d
z4d86a219408bfd4096582fbb8136c4ed7df181bb5db83702601db8517c180812cc85bcb871c5b0
z1b5523ac79437e27b419a6a43f4d40e21092157edd881b4a04787c4c7cef00a8277021ede9749f
ze9aa97e28e7efd148c7261cd3ca5fb1acc98b6756b6a35b1b039d6a7707e3a5ece4f746f7d3b69
z6affea0213402b948c284e6ee50822972cbba9b54100b2f48fcfe14a7d7a4b8ad29d8bcd01ce7b
z6b2dce55c13b48f85137c390efe21f0c1983bae67b7be0cfc24a969abcb6821b156996a63886cd
z5fea27d4716d8c4797c6bd56a53e42e3329fa6b6be0e6e4124fb7344f62dbd909643481f3ef4f5
z41ce4edeb1293043aade329f38a675e1f488aefce4fbcb873dc285ce170139f4360b54e23b0268
za0fac961cfe800dcd592af7249c6e8e0a59daeecaa6808c263244ffd09157789c3c643d3ac4c80
z6337835718dca1b785691e506fdd022e342237262422a8125c54a41168de5c5509778f35f4f933
z8399b9ddde70bd2a3ef909658480cb1585d07fb8f23425520238d0b1639000a1216f7aedab2e3e
z9087026c5285e37809eb821c5f386b525e34c027b388182290e72276ba3b9164f7a943ce18d20e
z398579f558fccce80626103c092ec4abb63f93a3a612befbd45e628e9bfec2450d19dfdca33664
zff6eccd6e13bd8bdad9e61bf6400452770952eb40cb39a430efbfd1f496591ec97241b2f45428d
ze6e629618010de7641154255ea3b7273b56032f61fbf078be1590095bd3a643d8debb3cb5024dd
z7142d1d9ee1b908123028b5c0bad111bee76638a5b1146bae7778b457b33a6b3a4eeea8726efcc
z3cba01bb1870e23ecf6e283ca82f2a814042682c45f9c5562a6b46d4c2760b317933f5bfb1d813
z05b61dc2edeaeebe618ab2c3cda65a057319f92cf5d01f0ad8db8ca9cda1f7d5b85a84990657e4
z7933f4bf059b4222efbb7d0212e8521a42143fbd66eb250ffca1ed24964ed88900c4fd11a5ead2
z7aede747b4edc24a7687d82f51da9d4ec5e9864b6a3503912b8e63c4a248697eb1f14ed8a3be24
z34d1e2c6d98d57604c60b917fad614887f156b007c64a216e19f76c827afd19449b79332f5c81d
z4ea60b553e9398d7eb2e2736212c1d494ff3b9cfff4cf48bf64f1afc302c1aea89bcc045ece18f
z744a9b2addefaa316a080d58badf394ab15f02b1c9cbd3bb481d37e88adaeba6b2e0216808b286
zb908efb37d8d8e4bde33a685f26576b00ba3ca642854aab7421bd1f04cf52243fd9f640f9f47b8
zaa46fc792219976a345db380f65b4c79fde522a9896ea9442fe7133958efdb8f88414224806333
zeaf174c24ffe4aa498d8d372ad985487701170e412a46bf4cda78359a9bedac918473af82521f6
z0247845d4e6be5cecf2f0ffe72197c3e9692ebbcca9f795f865c095dd2f13ce89df9a3c80bdbb9
z80df1c257836469e645a0c7b2ae5ae122dfd060389983a3d595eb124b786dae385bf53229890f7
z616860c8c4d55ff94d301e82fa4953f1e909610a4498329c824fd67fd9dc70f115dba31ab6fda8
zc2308853608c88ff82d026ccd672ef6ed0ab19f9ef508c54b5a89a0989ea8d0247d395ad15cccd
z79046b90e955c8ccf46443dc04dae36517542179a181b2d671f80448cdd90b4107a4189cf39480
z029aa0a056f11844e9eb3fa24b3f77b6197cc574892b026b764d620bc662640448eb997e697910
z398e3bb2263510cb2c4ac2a114898f9ab8678d8aea2878b1f76f184b404c3287ac8394cb0ff450
za18ace339990a6c411a7ff2674eabfff5e5771e6cbf1618b5719aaf0d164c1915fbd2e71b3af43
z645761cd08398e75741a8a0976d6a1d41a4b296987425b89bc46700d7dcc3e6797f6cc1576c1a6
z3e98b58418d84e9c5eb45fd94fb6f42ad32eb85d6f2a5b0f92938aebf06ad98145153c28eb4371
za29c564c5cbe368bfed96deb9fcde76d57828442493181bda08fbe08b5d2d242fbc1eb81b3b5de
zc54557f53b0fcfbd234be06023e7cac665cfc005bf89f8c8c9d6f0b262dfe9ea4aa617ea6e7073
z17923ecb00ba58fc1196acfe65f196bcaca854774722e53205868c26c4ad63d32311f9d1ac99e7
za6fe72aff3b32e9552dcca57bb787c00869155702ff753d2c54e2b9a379d59ebbffeb0593777e9
zaa8216d15b3c6e1a5f4d4d2e9e454da349cd91e1729367cc537d623e1473a97904340e1620afab
z5617cdfecb18058cf9366937416e3bb29f3edde5a987e7787c6977ed6690a50e894a3ea4e0297b
z77624c21382e29e5b494e949638f8723fa1c3fd345841176642cf9076a58cd1b96bb1d3dc5689a
z3390c2fa50f35f2b8ff538ad2f6430c7aafe5fa43f429c2074c2fd2635f3062530a11fc9f1d0ee
zcb4175b2cd8c7d1055ed4dce2bc967ed173fe79bd19632dc72c691c748d934bab0010e10637f62
z220fcc8af472c2404bd22c068a70945da322be839fa8114330cdf3e9717611039c15403575d580
z14d3870b6a6bb6d2a57847de58480c15a612c7305e995d7f0405e421f1ed36034b20f3ea10f05a
zb5e7b1b13c0cac3b85589e80fc91889318d83095b0ae16455ee5722098cb9c7b555733aefecc74
z2a32deebaac151c56ca78ce14bd0906b9a2a39b80b735616d1b26feaa90de338f506582d5a5ba7
z57315e69167dc8eced9c57a8be7c914f68978f04d8ae52d3cbe20d6aaf42bbf54f42b79bed2f9c
z9e6076957fb33f76a68010850a7a12746bcd646f9e45098b298089519c01139786140ebe27cb15
zedc6e2da3112266cb7e273bfb85cfda5c39f939407997ca16aa2da4c629baaec491105900d8eb8
zf1499fa376188de6279fd7b5d0f9ab32500f93760a54bb11acdacbc5f4dedb3adac71960ddec28
z47c8f2f062a1d4b6eba0b3465d0e20f3db1af91752005f81a66c505b17cc01b4bb764654675bd8
z87e16cc47d30ed9c4d5ed96eb515f233cd5b772b4f3702341500050fcc4089a3c03721235b0689
zdb8540dfb917f59c633148d87b9d3fa8922763cf082f24d49925d0397e00347759b05fef18c83b
z0cc7e9d706d96f5d04757f8cce7d90da82df36c7e8fe0dfaad33bf832bcb4b2e0e8e67d0bea0e2
z984f1ff20d1b10b0c63a2a7ba4385b5fa9f20858f2949606d13563accc6f191422fcdd9a441a1a
z82f589753003ce8a0805a4557d711c3aca007cee82fa1c11fb758b670a811cff65b59433ee2333
zb5e5bc29a75e81b4b393d3cef7b2a141f196cc91d3fb6a667c5347edd47c7f5cbfad5fb5dc2974
zcb9f3ee0935c74de75ecf57d81f9b85ba9c52a49bc8fd3d1e3c12b8da3cd12f659f528eb70dcba
z0e98fb69ca720ab1ba469284e79f6e9273eacceabf31e5e6686cce34790048b48dc4cf313ed676
zd47419a1b258d4c1dacce51c15165b6b899db0baba67ba504d41a9b6b7fecb2b57663ef4ca4418
z987fa8a74fb3faabf1530d4719d4768959f9b4f88911462b6b939cdb2ce18a9fe58d1cd450c68e
z665b4f62945295c8621d5ee5273d5e709c8583469bf02ee19eb7d89e53cc6d9f02a7c994ffe14d
z3d42baa1d7bc7041bd64c959f28dccf53756d953091fba7c2033562e19def239bf7ac5fca0c7a6
z99fde148973797a259aefb9252785d44aa5b65518ba8dca7e7ef826272358e8d63996a6a5f5a6f
zcdbdaaec53b287a052a6c09332edfa1f5c3f769e16ac1bde83bbb69925f3bad32019334ecd242c
z3c12d912c11773ce3e0d0bd76c661c774dc783a9fe0f6cd501a328c737782dfcdfceb39f37317b
zf6569a84415dc3b52f6550ac3fd31f27ffbc2e7e3a101b9e2c5ff0fe7998f6379808ce9d3a54e8
z808e3db29ba348ccf99db41e098fe239fd0ed26acbdea7ab39fe2d91996934032f2eae61d56c29
zec4d41120f9bb4c8fe51d4e554f63820643cc3c35c3acda8cd6c85558bbd6412e1015d25d8a736
z7ec942c9e74e373f203042444f7a447e7f9ba0c44451326d06088928a39d3f69be995c750dde1f
z94f84bf8aa48f9c9424534d188288207c829e91777b7dccf605894f49a9637d3b7ed97fca7d147
z0c34e0c47ae52f0a7480f96ae44a966fe5f1e890c052a39361437b765d022f6784ed7f257c511a
zb45100281614479ba4b273e1cc5c8da8c83b02a6a3842f7786b4f2d34be5c576ea7536dce34a34
z9edbfcfa1233038afd818dfa610c93852ab394670c3f5c8305a8abd0e42b67f872dfac97477ed7
z71123103d966fc434e79e2c5aefddb77a50cf7aab2aca6e4a5751b220ce6965d1870449a4ea4fa
zb6939c661e4000caca87b7daba50949a074b91234071fdfd6f38565831f2891d50db933135982a
ze5a3c4d5bd6c337595c104eebb050a6115bc119be3678d850cae0fc16422e7c88016a7306a85f4
z3700517f164a9f5a6bd4a49d3e44f370e8eb5cd113e6d56819404fee1ed19db8292207c621cfce
z54d9b3aef26183395af315dce1ce34b3be54978ef8852da452ee9eeddaf4a7122279a0be7f9b68
zef6e7170ea7c3a352839d626f9421018c8dbe21962062dc57444b7ade6600eed95b96471490e70
zb343e9236081e644b5790e570f5e20af46c82367f80c8ccf78793817b3d130efeedf659343a602
z90d6058face31eecb2b184f4c17e0cac5ef190b80c151c6d8fb941068833207cc883c358dac35d
z17106f9d89aa761ad2020e1d0b8e6dbf3d0e390bae58d0d93abc7238ee9a53e12cc351a497b53e
z3d44a7309f55685ddea0e31c5f92f846f80d1756408a39433bdd6227335143f19a89cdf298fdd5
zab64c6b93f47573c55483c3648cf7e7240e47bfabf342e4f3f75ab2679a5cfbe46493e51c1f653
z935a0502d5545506333074a982a911ae88f6bd6222c4ede517ff0bcbbdb066fc4ede5f9aef20af
z33bf83d75b996cfda135f0f0b02b25b52d01ad94c1cb5298ecb70ebda1a63432b4201d7c702f18
ze05c564613a10bcd2432422fe44cb953aa487fdb920834ca9b66eab5e95f93a6a4fd19c006088b
za35c02ccf45f98692934d5aa5a6681ace6e88d0d7e88f40772d215612170b6048af0aeab452387
z8792928cf2fbc2207c444a8b286894a29b4dd05da41f6c9cad9419801e304f7770151a9fdb719b
zfed45e8d3111a7c29abca855e7c7c72eb80c0f15f147c6ff2fd87e1e969307e45a92172c0f157d
z35577c34036432c60102f899aff563f582b4697bfac323417ca12b7e862a0a3a3b17f805d9aada
zbce2e85238b7d1d1bf31ce5b995ebd48f9c0c64729ad8339bc2d0a38d2b46d92bc402ea4cf9fb3
zcf6a3fa725aaa2579999a86281e7713feec479638cd62c8e11cac7b4d0c7b1f7c73924d9576c41
zc8070996570939dd2cefe810139278a6af9abb3a7d1a11784acf5d963c71556c5bbf1ff24fb197
zf4f2fbc4bc18cf1f86891bcd6aa3d5157928e9df92b129ef0c0a9d5c408cc2480dca4595865a2b
z3dce96cd57747f6c8cbcb0a3f127d4d386d55ff4fd118341020b2ce4a35ee4814085fa541acd23
z4cc69faf8e5a6c3103c5fb60a74991d9c2264154224d22ba405e04eb7d51559b2d04713269732f
z8119aae471431be0ecd7e0387437c6610878d4e030aabb32153e645f16f23abc1d1e927cab8ffe
z31f6a399eda9718b1d2b0ba1eefc8addf26e7d50e637c326652ba73bd819b3e863b395cebf6ed6
z564489eccea4d8ee58e14c346efafd988d79597a8331fa34758f9fca14d49152bd0f239ae4fae8
z67dcaf134f3e2d49465ab2a6a7efc3017b1955f9ecae78aba98ff29c0297e8cc9c52348e440805
z292c62949153b8d511ed4e5a5b7a9f68ecc7f146317f44fdc5e64f998f824c27184f304de0f5ef
z382e0e59053f0801e6ff092dac56910ef40cd12d4b4eccfd33e0cc919e13a3af8c61edfca25add
z628d45899a529b63fcccae601064fe89a41864232d3614eb6425762de9f6ace5bd4c887ca7d282
zd61e4c3a0554649c681c55333074788c880de13f7d1e75926a56ab6ad9ad0a1c35ddbcf58f452a
zc8f3f19bfa726e411df3b8cb345fd0f697fa2c1b4a22dbd9cbc249e1289f19c702b5c226a60964
z3acb6f0966bcbc518f1da4baf1b288f27eef05cc7454fa221ccaa86cb661310d74f7da95e275c6
z602724303aee3b916f5f2dfb7d85bfd2c760fc85436fdab72a0b21613f41d2b5318a2247d0e822
z77f7ba73266015640a83f30490f734688b36a773173ed717cd0411ec66cd0ed8cff368e4a41724
z8fa08737974fbfd0f26cf090d07da7ed80cf5b19e267d7a2a6e51c0e90d458b74aa2e1b5597f21
z1b5c66be750a8510b05454231a0d33223db58b4461082a24a9cb20792d3d255bc0ff130b6fcbe8
z4590b925463bb9a882c5e3f69feb1ef5f6eed58df7d43d61ce60e699d0b692d9f69dbffadb27a9
z4007f439e926efce6f6276f9154830c554b93d9b9e63bcb2f1878c0bf48d329fe0d2ca83364c57
z4ed8d993f10b1ab464980dca1d2ff9ede97695ff75c94e4e1f5505bc3afc78cdc8218c45f614a5
z2b0f546ea1f58dd469cbfc186d560c6079984ead4059a6db9d5a00b30b83afa718a15bf18f37fc
z44c826f2d13f2c2885c7e1549a4127fb34a235167e0a0e92898c2ad7e25a286a8b44bc49c05684
zd266b25348affd4d9d6877f0c40ca9acb1a73408f4bee98b240e42ba7581e27e9d040b793ae16c
z4527e7e7598fc1b4b9f3b72afa28de4b04dbdc673cfb068a43ff0225e8434e58f5d5bdcc80e13b
z755548287eedbc212bb9c6a27e34feb5b81111b1b48afcebd230b33b43bd3358d6a88bf5954249
zd3ee4235fe129f0196fce3ffb36856df69bbff6c5a12cc2be746ced6a3fcf2bdfd0a633155dcc5
z7224810277c88dd3abd192946a8f7ed216435e3ea309f9253b7a97af844f6497e449febbb1739c
zcd6f8956aa62716aa084afe0795ba3e75e34db33dad6409910d8c455ee9ab2237e585ca2042928
zc33247c2d925355663470c2badfcd9aa4da8470efce1dddaeae5f29098e3e9db4777b4c7094f98
z771f5bcd633aa4a323a155d772b2b484553ab3594956d4a591079ce15b0c79b590243e8cd6d38c
zf7ea3eb235608357a1fe27a3aff08e04fa8376143c8b09efdc5a4fd7f79ed5eae52214f41acdd5
ze9d7d4ad2e201ffe32d71598603d4781fb6d226bb5ae048a77f58fb98d1036bb90be964c422867
za831094241d342c9d74e8da5f10fa8ffed06fe5127f629e233ef4e98d2a6943a77ce43f7291a4b
z92ae79e1ab6f12bfe92216c5ef1345decc962443f80e82177143b28cb1fc88f87f9f41f9d9d9ba
z25db06ee5446e9bc6420bbb3634576a0adb5357ff66f8cfa1562b0f51f2c3d351e3e75d9932790
z2572f7663d0f6118fe70a9bb7f437fb28ba2dfcea9576719fe76cb684bfdbc09a3284cfcffd2f4
z70e35599a56c419660b362ea7bc22de4ea49280917b351cff0fb1be4403e2b657c26ef7c4bb866
z8af60d6537015da38684e8f02ccd25126a28d6339dd95fe65d9f57eee4aeb5f359e3e15c0fb642
za519f14e08455b63b023374094f4be34eed22f1e7d507fb9aec2d816b50647ae3ada2a9ce46610
z6bfa1401efcad1049aaf80898ff68100884e1d23743e3742b7f6c9f00e213e053d2ee67dd0588d
z1fcc261af0b255770162952ae1cdca49e948c7754f6805961186d84062954352a03ab78d4ec0c2
z6eb58b77f2e96f9b032f2c3adac15a1cf9c0f03af95874fd3d98df4be9d284d8a5c9ac10af0dba
z4ff3ede9ea533bd56e37d6f597c684fd21b226f06293fd672cd60a825d5c20f41ec9edb8871e74
z70ec033cd81a7ee3e0272eb0f3f7e3f82fc414847f25bf3577c642ee37062f34530726188ee076
z6da92c54d0289d68c51b6e2e57938993093fdce177d70b49eecb1fbef345ad8c5163816626abf2
ze814bf87f93206bfa8220e0a94ef3bf9e109eb9715a95dd50638c92bb3c38b3d973c814d36cbaf
zdd91fa61def742cb84175ef3cfdff3b183735190b24379cfc3dc07bf57c537f91dbe730497e27e
z4a886f872d635a2aefea582b4d07a0c48eb88e0848e19553195eddc434133024bcdd804f5f4623
z7b2453b4ceeb31125a378e33973071cb6dd974b397ae9021ccf93ff222b4ddf9d6bbc426e233f4
z037f121e1164221e249a00be5ba84fbc8f272968cb128782569f842dbb5cf4044b630688e9e377
z2093acdb5eceb318c2d0a0a5f61a646dd7486cca44a65a5815d6e56d09f4405de6c2ecd6c1580b
zb60aa15f890905da82f5827cfe3bd1cc928acda2325d7190bcc2321d5dc94f9465e166e6c86716
z1eb16415f75bb1ac50768528332a30013dbf427dff5f64dc52659b8f18f647e66f0caeec615645
z4d0fff23c4ed2683e629316b6a307c28ab3a02f0f773b147c5ad9b39304a62905b6599fcf95bf8
z1085d0a94352328206fa56e037d1bbef3a1b1d540686992bb5576890912a32686180c3929e62c6
z8cd59d85cc8b7b7676294876c623d1a45cc822f14fd970c8e2f2a877e15e7b3ab121dd640cf58c
z58d167ace65aea9ab72dbcb65f7bdad58c62df1b5f67bbb37f3ed7dd14c6b1e417ca9b84cbb77b
z92781ee8cb4c923c7875b0e83af0f23159072cafdee46623d63b7aacff632323723dcf2375c9d3
zbb7bbc9d4021b473a3fbb0004c70adb11672d2295de68beb7f4eb360e4771d7168540c76c66539
z7735751eaf1b79502379c2c44154698ec4cca9eaf5ce7696bdba4122b433351403a31a93208541
z80f1f7943d5311377c4f3f1143d9776f24c5162ccc4cd5f76e529c42554ee3425babdd374d4707
z859e360f1ee69e681040030c117bb4313d1fb272261ddfea0dab4fd9e6ab7e411d5a1748f6fb53
ze59ae972058b3a5b10f9c36d92c8a3ba50352ecfaf3552cf6f23b7c1f8c0db7ed39a11882322c5
zc7cd698e702216a958a4bfa8272d234ae6df48f010fde94f9cbfa9815aad60a3034d025dc1
`end_protected_0in
`else
`ifdef MODEL_TECH
`include "qvl_multi_clock_fifo_assertions.mti.svp"
`endif // MODEL_TECH
`endif // encrypted_0in
