`ifdef encrypted_0in
`protected_0in
ze74c34e226135848fe16db9ffd31815111b6d7fb642c521a3f628cf6da949865580b22efd062a7
ze90adae0e65e66a2c36a587d0a790699161455169ed55a01f2084f11770a774ec4c588039b380f
z6de9c5084882a40b79a175f5c2114b2b6d78b070cb806e1c0aa9258297f4687ab308bc470f0040
zb0b1de382961eeeaf2e279e1462520fc31c119af8f2b214846f56c2b3cd2eadbe4099496abff18
z15cec83ec4a77b868344aa20ba7360908f5c0de2a79abf8b3534b883bb12180f68b5d4beb444cf
z3fba8f13afb0abfe8fcc4294810f75afe452434d2d0f1166236c82f76edf1e12979f04bc35693e
z32ae028996dd85737a8f5adc1ebb94f39c940246e887647b64782cd7ab429b0544c173176cede7
z01dfb26b1f73408344a52b7e1f117f12bb9c8077b34876c2e6fdc085981637012dc9754765e1a9
zc512ce062e0b8fb16a214591f5c81e1353b900a611fe1f4886b57940b41b7f2ce99a7b84b04b90
z916f717e73bd10589c81e207ed77ec660a8cbed5b487fa50acde1b055c8870bd8676023f21ddcf
z9c98cc47cfa2d654ff1365d1f45035a045a66c5dfa8279050262529d2cac9e64fd27d9c7de62a7
z731bc808811ded9016570962244887f98fe5440167bd0088f2f049df882af501358497c3b28776
zcdc5426c7f52a851c35106bb93e16fff98478405fcd4d89273452c559f93e5926bfbc31ac074a0
z0eb509dc25747123e8481c4f7728976370d53c0acc5b7a10882d5b25ac1c2eb5b8866d0c37cae9
z9de4d2abd2fa8c576bb458474de01f84b89f9c86362ffc56bac062e009289adc34add479dd2395
z1d5b66a61b1927c73dcc2d92451f6f0018939499d867efdcfa4f8946d333f9af49c73898f14ff3
ze6b170f9065a89e725796d3a1ad9792052fd6d520015953a681463d1987de3f592a9cf054f5df5
z7ce96d4867a7e9d802a4bc81b4244e666483e6937ed1483bc07dfb43ccdad1555389f7a385762b
z5e9d31b1f07c53841ed2f610b0f8f4d06671a1c8f56b46d46cfe73bec086b93bac97b354796098
zeb462ee3ed698949008aa8cb0ea3cc494aa276e87466c26de178ecc8afa7fcfeb445d3fdc889e7
z1c1ce85db92f203aa6544ec67262c856e78ee51879ed533a899e547b9289e71c06b719f81a8f8c
z813aea69438e3c15f6893d16469529f728363d642a79cb70f3972622fb75e0ac263a90c9d37215
z50c75a34f0934b01ad5934398e3e812e6a881df530d488496b65579c44670fd0ca2cbba647b099
z460d8c2315408a2b3edfb5dabf1232e0245dfae4fc34e1070958e7dbcd13e2b4c93c2da608d50c
za4e476aced9e61a96e70f2ea894ee218e03b1b1daf6d6d63b822ab74f460a01e729a78650cfb55
z0c065a896d1087e4763d2a8f22ad6d1a72a9c1d60a890395483f24a8b4733a8237c345ce2df426
z85df0dfaedb34f8c1de6159f3fa40ca43fc0df520f29f1c9d7ab28e721364b8e20f9b59328874c
z63a0aa540d679086ad5736cd5d5aa7af2daefcf1612f3dd9f54cd6cbd2a8bd64d5572a706a96a5
z7b3595a0887cd1e0fab4e24d8422cbbaa53a2d4393f3533ad6df0a0050f0704e8c28386123a00b
z8893f3c4593f27d500675dde7d4f8773fd871ffb51ca9215c46c5a3ff096d256750fe15743a601
zb7476fb1cf9c2de6bf983c20461c9469d113f4a906e96adb035f8242066245cdd248fc08b01da5
z9464955235dc66eb6c99ca2cf1f6e64523176b45683c3b2b72e3d0b6d83b119d08a883e3c65e44
z964b41b023533006fcd5610df5ba4c31ecbba5037117e62c6bc9b417f05377b12cdf9ad8c6d303
z7439d9e035e59718f47e2d87050334dfeb5d3678db8d2f7790dde7a6c7a55f5fb5794afffe67a2
zfaaee6f373477d281e7254667dfbc3e1242a01e84b7166e542b6fb14ba17fcd333226259a40172
z734a57455f723a5f93dc01a5611fe370fb074e888b762c4e3f69fe6e72718fd35dfd74f9ae9bc5
z0363b738863bc9a65db9a243187395aa22c49f420a7bb69f9f14a7f0dc36fe4b229e51e03bfeaf
zdb2c5b98dc9a5e90f8e4649577eb59573cc3095ca0736f75e8738c0d50c254bd4fc4a652343267
z5aa28f8469e58d19a648788228280f4924d82cf00977b4914cd0857c802f524094df1cc6b67967
zb62ff041483cbfc3c5862ca2ac923ec3e2fa2193d8e4d5da6ebb81e1c65d6a2e27ef74b8a9f11d
z294b98ee7b9fdc61c67dad530e46e3038cbb62f7f2c7925ef3bb624db3cf3f45c1b374d20bf81f
z9d52958dad65377241f258c34d50849f06d8b14705f3628769e8d3b0d9c375d3a022d6da41536b
z088fc77db81b042c03b567fca61cc9d9c966049278dd77edb33d437dda2e96c144876cb53b5186
zda130a7b09fa9a300eea4cb004349927fc366aae4b1f4067d9ce20e6ad28d7473e08208fa60bdb
z9b5c855dc398a815bf7c709a0791109a684398fd82c579a8a3a5fec2229323a1a194a794e7d2b7
z60bf7e1dc588f66dbaa3756e425c577d0bb67103bd50f5716dea50533abad85d00d1a2a63c888f
zc4efd3b768ed569cfba51a46fedb1ec5309573bf1f5df31c73d3bb71fa8a71ac5a853a2dbe8c1d
z3678d0e1e85d839ba70093a1617bb9806ba7033b02e780997478e996a9165bbb792edb359f777c
za8da0af8280675fc971b4c41162df872cde50c4ba5841502933774779e7404b23d7e4da093f84d
zb8f6d5d73b90773e272a81590d48394732b9e966b2441ef5d86883b845db1272e1cc577a5fc72e
z2b847ac6b639ec2588f7cffc2f12e665de185a3d32ec48602d837aef06fe7067160e1a40642ca5
z40b866514246e7455dd9ff1285e20c6841638159a0fba98b6f47ba0a20a9677f9036a73c0e8133
z16c44d4b94fbec4156d83f88655364876d089c9f76dec35b9c166d5f6599a922225362f2d77b53
z8ccb3fa12a38092e30d4522f7dcf2595be75032156b2b31b2e0aea73de8ff03596b8e6ede05d91
za19ae90632506047f92fc5ffc35a89e9b3fb3d599483faa14d7da70ad6d139541c992c7667e6d7
z0f3bff1cd38e6513acf6d9ea5d4b0bffb99ea2c76fb8086f827a9be0be23853453ba9fa0d74943
zed71750589e477f0aa10631612b91155e61a14f860f34af04c47c820911d43ee49bca903f0f880
zff1c526f232f97b07d3bdf07e63e220badfd0876e204340516be01a5e840542b6e397c3ae60a6f
zc88610993446c1953210cfdfe1b1de7454d5a90fdeaddc088c5dd86b2365b2def2021fe6b5d712
zeaaf09ea5ff35eeba5856a9ded9421365e84e0b753b0061ba3355438a014a2a61aa3b733670d14
zc41fcdcdcf12a3a639e54a3e6282fa1d440204c3602bcba80bf080b0aa329fe19116458d0c1262
z3f5a4a45d3fa1072e6a17af80d1a8f45199a5f99781d7e6a001689af3bb408f7b78e96df8a5be6
z7951d048981b3ed1006a9649ab8f9a918f0e84cf506cc2d009cb2dd9331e5e3225645e09bd775a
z6e6f90c3155ab107c8bf1b2dc8759d88e436fdb8caa65a97e3e70a940ff9305ce8e2a3371ec737
z4eb97bb9e8a40be26cf267043feed2ba1a0449d36cc9ceb99ff1058b3111118baa0c54f60abd3d
zc48573370c5eae4cafa52d8f38d79a43e6297668aaddccc54d1e5222f8c0c26a47f30a53d1aef1
z568bf03a2a3b2fed29f146ad7cd2ea389e11612a7c483305837fc610512fbcc1e4c042268080bb
z0f155057791d1c669c21ede299718415d50f88130baf982cba2600282ef8d337ad0d7863317db5
z01d863100162e2ae2f57dcfaa233a98d9cef8cb819f29b21848b8374b4b3574df68eefb9321614
zbdfd939f853eb23ef2b74326b798d2899eb24bfef2f384f3cea48a3f6ca02844d93c7211bd41b0
zab78d8bec4bca1d7cda3889d82890e3ce457d7f40086861a273caea28785726b108d07110f21c8
z0511b7c89d78b80f1578ba33e0a624720c66669a8a4b4d1fc4f6ad14fdcaff5d0bd1ecd51d646e
zc23708f8011c5b3ee3f709f3a2555411bc323640b16aaedf77d4bb204ee6c430827885b81cc865
z35404f9051be9ca48f5996bb636a75761083beb4ba5e03584fd0330ab53f5c80ce30b1368de52b
zcc2fd4c6451bb65d2e968be637af7cf6441da8394725703ba47ad9b713e156d9996fd3e06e484e
z09046bf338875c1d1845c9c2edb27842c7d7ea5ccd6e73737c7d76dc77c53a0694d73b025099ac
zeab201010797547c8bd71f956f661cb000afa33cd67dd2b35df9c738b6ff3042e2aa75648db09d
zeba3d14116d788d9889b80610bd94f29a138b0acbab7b0a4cae33dc9815d689d6c559ec0b2740d
z96227e99efdd3ede4cf21606ceae58340e3fdc6f5c91615fe0a5e0d2bf729fe85390e658a9c432
z8dfa5e9fefc465d4357309c084a4c6eadd161ebaa370d3a24e16d9d4e796a54490faaa47a641e1
z5cda25f7f65c25999c99673884cdc169ec0372f17d91226097e915acdd425ec74cb7219d970a3a
z79b14ef5c3faec818853e2e9c61d9fa9bdf27080e98d521fc9bf9279281a74d07bb05e2caf8cf7
z92aa8309aba9bcd4dec9efb41ad67f7ce5f1fb11c726d8acf34ec149720b913f476934f67b6d50
z5a92f1cb4534f8cef6f67a2176baf14d9c23e8b57bf484a43cfd9eaf3560dcdb0dc354d4c91c82
zdd8584e64d32f61b9bd2cfa4961194016ad0ae9d1f6c2edc21dedb13ddba67f6304efbd0e37219
z5b02152aa1740e65ee6a7e75d0bb84675651e45058e66a385a0235bdf909b60f605cd616079a73
za39d773a22c540a3574f1e47e4f61c527fa66ac2d5bc0357189ef44887f2a4fa31f5b70833af95
z6708353760f2bdcac599218e9b2de6c1fe94511a45b010bd9fd0905bf3727847541c03917c036e
z33982d67729d4f720f58fd698d8ccbae10cfe08300dfb5d31e593c8678de976317a6473bb35595
z95cbaf3893253473865e2d8ed6c77d475c29f10036ad1eb166d8bd3dfd3b99ece60fd79511a2e0
zfbc9e4eb2edb42a2524800201d17e45f5ff2603b1638af7828aac5e2d3f232264e92cb89b33241
z8c0db4bcf00e147f43a3edf5867c0309d5834569be1d02ba66a83e28b418cc303f45f66e1c8f49
z23d73c3b81e2647cecc466ebcb0fa0b9e6a9b65eee2845fe2d2b51c660f63d95b78fa509ec2b93
zb6f91d051c7241b0b50a738e312becf17ed1e08131a392e5d229081c558ec7dfe5a9a3b9b8df6e
zd080a0badd806d017ff85b4985519d7562eb514ddf5b8e0c0faf6a9b2719e3b476543485f1df43
z52cba3acd9517ad485557857fc6b436eccccf42fb7950ee5c99dd1a069a8ab138f8997afcda8ee
zc64d40c0569cb1efbed3d5202c1f6500fdb7f182ed4b8734ffd73be8b3bf2f4d2334c9890067b5
zd8c102475031d4f34a4678a4635bcccbb989d438b9ff3d22b41daa34468cf76be7e926300feecf
z538fcebe7f974060e9ff7b99a5041b3a9058141dcca2e52ef133378de6b27a2915f9e7c191643b
z47a83bae92a397537820e5e4a3febc3940318fa0f221ffe3b4106bbfdd058ddd072a38f3242e62
z6d3cc13d8535017bbd541af42744cea597675be5fccbdd81f556a29c679e24a18b884e35179a68
z9c2d228aba1b7b7e71a40cf03b3fdfb8da8abb22ea26ac2fbb77f4e0c8eacb586557564bfa7c19
zd5479b8a21dc706ac372d4e479c712a1d432a6e83cd04e9f807434ca96b340d904c585c326882f
z891ffb1e3d56c26448d1c0900698a1ad3573a8dce8107cf3d00756c356cc3711a907af184d9f48
z7e247b94ac21315798b95920978b440ca9fe9eacaa2057781451755669c90b17f89002bf711f27
zcddfa1c4031d3d18acf8b6df752022753d1373d9639866efb0d62c25225dad403dd7c3a7509707
z3224d1dcbd9757d76c6bd7c4e275b26657d01855036bf8469c5002c7cf2d115c1bfeda74259df4
z8281cab44eb9c1696e96aaa0117db82d8e47640a0397312cb97a8d2fc9de884656b9a4281bce1c
z12ebfeeb04c7494693a8d580497ac0489fc4f5e5728fab0cc4dd269a7ac743d6f1a264a314abe6
z6f918705bdf8de5df66ef7dd20285c0dce3d08657f232c1c6ddf0439a05ef1b959340877841e57
z4080fde2cdf511cb8b72d8659791909fae5dda407c6135b4a9e870437bbba5399bc6fdf3c11173
z83aeaecbfe4c85e93e6bc343185e982cf4e193e0bd0c4617ad2b4944fef71384b9b80601e6540f
z1821f407ad546312e41a490dcc363d4e970595bce8b57509a0bd70c00effb3bda2080149088f10
z99937a4f8131b15de583fc0a3d29c5d362a733b340cc64f80f29e65bee746f93e788a7c514d9de
zb9e88269ae60de23f3a53ece70e0367ecaeafd4262165bfae515226bbe8422faf788c03bbdfe81
zaea6ccff03f94dd166e61ca6b90bd405508d895a33ccbbb367f992eb5ddb99e34c8d4f83bce23b
zc15f29998bb63fa9459541550bdbd6aaf7aeca178f4c0b2e9c714c8f5a46fb2a5739354f45ca3c
z6e7d39b7a3af5c2d589102c9dd475ef0d3b56bb80d3a0dacbd49fa256654dbc7b2711b0bd21c42
z6685af975ff11daf5d1c0a6d2f0033dd79740d96c4f5cbb3a94b0ca40d886b6277e0660b4b39df
zd4a7178776a62ebdea283d1e6206a973c6256c64a8f6b1feb03880152158333329253a3ce0ec20
zedb49f521f63c312e68c4a50322fc38f3f3d6f47e92891299d73c1b6aecd794bfa5dcca7d12369
zff194c19a577c97e0cc93fd9e93fe2a4e5a1adede0940c1e97029e4b76ebc95017639b7f038b4b
z00cb424259cf93c8dec42c0ff45dfb1ccf6dc85b242c98ff7de9ce6dff040e4739eae621716905
z28fc47b94ad4d147071d30115aee08ab5530c3612567c2d5497f1d75aeb7fb5f6578a11bc685be
z87fc237b9e0c419d3ff9c1dc38b0f4265b9891ae319f38749b24472c00dc4faacb4d993a4c8939
zafa8182785e21e8d0e80ac2645034203e7161f93dbb7f4a968af92c1d3e23a073bb3d1a47d0701
z096e44ae769c8b0658a2893507dc49e8a5517b58acdb9529aea311cccd4b975aaa0e286fb0f0da
zf01dc933ebabaa3a4c3191987ccb255d191fc67d4500c4a6354f0140190a4269a2dd1921c5d0a9
z0b1ae6736be8268b01b095b4d2897c21026dd7a47ebd4027e17016e36d781474d6594e2099a72c
zf568a8865e9515f0ce16fe4d475a05fcf92274b09be086a03c378d067015715f17830f923bc475
z9c846a2341ecc1bcf1d11dcca6c2389f441ae6d297fa458751e6ab1267d3ea4b49a850d2a46b76
zae6449cc3eaeb1cd199494ad548bc34d961cdf1f074aa98cb0179a59774eb4c8ec3219d6f3ccc1
zae9d928284ba997c59474376d3158bea49fda86df8a8f6ba676e0eb447c1473e370e351d417044
z45a579207a344480cb0f428c77eab0717acace13f2dd52c060141d340f69f8bd03ace0495c1c50
zc23e688b5763c8f04843c2e9aa719936ab025885765495ce7b38e1984ddcf80954fd3dd7f97ed8
z0bc783e2139f3ff1ea20ea39112664517351056b1179797bb77b2a4c2e529ebfa6b9ff224975a2
z1fe9d659f0c5289071f938519b3bdc5e0292f2aea5e2a997d5acbdfd870d87bbbfadfe1fd7aa22
zd4a392510f5d6541ec6804fd0a111523da7744502e0fcde950eda6e0c2aad40723c5d124026162
ze2a4c2ae702ec42ff1f08efa98471b2049aee78168cb035ba968382acd6e05a8e4196214e6684a
zc1c916cef8e1aaccd32f194ea91762a6d65833658fdcbdeb93179b0caed4c8c682fa04b8ef9954
zd081ba5ddf46c103cd3f7386b487ec35b1b8fe8ba04e4645a13b7ed41366a6ce8624cc8cc5d2ef
zfdfe762a9b932203e49850e953b6baaf6b475c8e43f304fab91d54172478e6e655b96426e9d6b5
z778c843f62a5a5a5536a7afbdac4ad6f6c99719e0cb000b3608f94003f9400c54f3f4dd24fb1e1
z9b8b844006ea481e4edfdb6fc1f7d3f9eeef6a07fd627e883aab6bf7443943134057862cdb3a20
zd6d9f5ff4615571b9c08caac000b1293a338e0d321c3bb1a7995539a8d13da380aa6fe94007615
zb552ba62e21a6572c0fdcef1c8bc7cf057c55324dffe243f9f60b9ee8ef057bb42e345f341e494
za167e9f7c26f98fdcf4bd636df90350e2300e155f991106a21138f3d0de828010c7388d026c642
zc19bc5f29cfa0e3e86991729c23b25a44eae6e8cf769667e18b3d6ae0ec6b49b432ffd8f13d249
z4efe515c104683168cb64f4d0738a8453aabcf766b67cea7d3cfc6f07e33a0460a0b5e4b89f8ea
z8212eead0a7b3b4e5a8e8bd62865f5383cc78b586c199065a54996be45c399c2caaab497b958f7
z2b2657906b5e24b33c54ef0a23b1c529e9901962974fed4844fee167340bf1494ccb9d42f9ee26
z5c75cdb3baf6b27c0d4f20fb4d04c61964035e1d10ff071ef98b11050aa20fdfe7c5b221691a8d
zb14de560fe22fb43a4be1747e2e55f14a7df842b97c763da01b054f267b8a1c43d567a75b49c58
z2732f50e5495af3ab545c174f9ba1b66764b2398ca0136d1dd2adb0e07062ab9456b1caaf2485d
z930fa3c3bd5169d0e9ff9825730d4bbc744d2088b760448c4aaf498d6c93626bee9a3649088b6b
z90493cb1e6a3b574da82bf72b471f2a2b61cf054d905fb411fae64dc4f1f282ca3bed58ce89db5
zec10a81c93191f50f4754a2d1d841e6623b9f2d6e8a57c902389075ac1138cfd83129557407956
z3977a9a7c87bd1e71e8ef7d4f17ee8c23e97ddcfc61a6dad6f4191019cf19a95c634acf3156116
z5478faa542c30de3446e3ce04552d1cecb1920b6d45b1a080d54c8b7691d762f5bbd7fa0f96d9b
z5eca6c4965b4862b68f40035c16c65eef2f6c4fc031b61f5ce58cc7069febdf6d187724e31dfcd
z8145743eb17ec54597bd593e418ed3cee143f1a913daac79bdc2911f4b811236a43ec84c020c9a
za5ca7e1a95d7ad3d3e4d6b346afc09700d7c34b3784533f166a7a6306e5467454526ba21fe2f7a
zeb813e258780b77e13a7fff1b277dee3c4cb90442f063d8b8b4476d78b02c24a1d5a75a0c5ed82
z2c94bc8cf72ae917f5b02ecfb2a707d99acc84d006fe1a856988562e447c6bf896d0daa372bd15
z4e79c00607d96399d24abbb04610e4cc70e373e33f7214be82f5254c9ce6801b1a0bbdd9ee6dd0
z258670f8d432b9ca8975b0b449d26867f3e584fae16a5c80f12968bbc7925d7e0d2f49047dff70
ze7c8b49e667d3d8e265cf62830efa7c18a0b235fed716889d1ad3fd1b44988461ab1cc60007867
z3b761f6254f5ea0352052013585a65327467286f5deec6961ea134e0369e4d5a9f485b91af453d
z5309d8ec28778f8952f828d9b20de129f824abba8e41705494c2916dca3d423574ae21205f71e9
zcb723028c3b44d6ba46c9d13098f829a27de4611843edd8dfa973e2514fa8a14c8abdbee1a2337
zc6ac0195b2ca024ab09ca73e592a439b963747f647853991b7cac874d8b1bc34aa38aeb07c23db
z030886a98cce1d986241a956f71813f3fd5aa31b6b136bf9eaf7a65a71344e67aa2bcfc0ebf87f
z162b2dbc639a88c451836986b2046d154336228b6b7fb675c4feff32d9281992d3c2282621c43a
z8f4d0c71fbc311b0315dad11596cca1534286a9c9b35282c4524081917d79c8afbce5e9ba75605
za80e9252fa8ff48e0da25d090c4f3a2333be2372e82d090bd596355225c324e1c742b03be8865c
z5ee0601da109a7164eb5f5349262c87cddfdc8b913f98e5c33b2280bd3d38d0542f837a2d7f35f
z2d7d16c28a620248c4ceefb231ea8abef634aa18fe680ee1ff50e50b1b2ac779a40a00808aedc9
z387521342ddf5384422ee687206c706a747e85f12fe049283f5c416cfd49a02d418e7eb892037e
z9311d37b82bc2f04177afe08113f688f72f96049922d15f9df3173eb5aa49b9599c17a8d3e4d57
zf7a2267b5a3461e5a6038e29be55889077e9a41a9373ac30d3ca92e137f9e2d4fe6e405f4f89e8
z32cf66690c114b6f54c00dab822fd2f5c6d8b127e78ba322960a085138c3f9851f13783b99d5a2
zc0033a65bbc564d7252e516db3e74fe4d36a2bce9f1ecc9ece31af31fcb7be9b406d3b6aff0bf0
zec84754391e51ba882653e92460769e1239301731a4ffe0a34fedbae83c0dc80b2d49b1ba12b97
z1b74562af0d64198aee653d072ea5f2f45b133bab8e70017b3ae0c19da92a7059e317afd3b9697
zfb86d30ed5471c7619298084562cea1e8f94fa05f04ccee184eec4ae9e5ceb1ab32bec86483a07
z53708a7da4c1b91a0f55e68d05d578a7fb339c2becfd6a0a7870a47cc39d73637c32c84ae1b7ca
zb6fd6175c9d5bf6cc0a4487b54725e85fa06ef3bf47fcb61e21d306933d461b9526c4b22d18c5b
z25d4fe09be6f75ed3ba8ebdbf765dba6784f8e7e1d74c3ee9153485937382297614f4c6ddf6831
z2db56769313023d3efe79ef4cbf34168f4337568463631f16f8bce756a56d951b220a098fecdc0
z42c57893132fbf87dce1238fe454c3e908c6650aa0c292d5005b4cc2d74a4fb17f00a63fc9c6e4
zd9b7c5023c7b4194296989b04bb1791c9549a31f365646ec87a4bf1ce31e8bf84efa52e9500d85
z30200aad80f0e39195efeb95b0b5bc72ee72ac500046a0243a2dc8fa436dc93b6c1c6576bb3d47
z441d8361269b787de57cfe364cedea0962c95994ecd4819478ac7e07062c7e0990e18a1dadf899
ze164ce7da23d11a8363532a6c0a607c6d8b10970def64fcee854f4539f933a9147c4d3f84322b8
z3392c98160667891e620b705c9eb42ee4a606e54b1bc12733532a4e1f8ecf28893bb7cebae928a
z9dce9efd49ef702cdac53b0fa746dfc72ad5df840a04e778e88c948c7bba7cbe880a4a653e38ec
z969a99a04389cab7181394a2997080ba574df0743615eae21ba8501e236f3dd94db484f08cd34c
z715ae55accf3134ddb591c52a68895cfc00bb1de25f3f36a1bb6d980e5c689fb5e4cb95402a211
z08e39c0fb63065690aeff5f5227fb4b1e4bf0cc30e6fdade9ce1715ae6c2ce59e87da5f1c1a259
z8db24e2830726bc6b56500b1db3aee41650f00da2a3fab8a7b2044617be3b32831c14096afccb2
zc8b4399a0830f992dcee85bc454b895e983b5a06f7d2eda93d5efea1c1b75ee5ad31d4e129928e
zbee6026608bf023ece2bcbb4ba89d17e3d0e5072b26f98b1032d5aa258002d01c59c0ca912c8f4
zac61c6fd33540d98bf78f7d6475055b4cf87a15381efc520607c3838a645a360d39f26fab60d6c
zab7b5ee2043d49c0d49ba1be40c31ee3ca18c00f7cf26e105fb61b5d0cac4e6105ba9887941721
z1d74b0250e3d7b5da9759ce59de48512a9b123ec71fe04c4a6165d3da7f3cc41100e429e5ca7a7
zbf85a6cc49fab49ee8a4b8de47cbfa9ed3ee43bb3e9f727ead684fec70d0f157fcfdb6db87db91
z47c682f5b97dc92baef54a76182ada769f41d226234a31a7724dd1a565ca2339a569403bd5ebf1
z6b22830f8abf0df9459534a51127a8a4c0a41a58d0f978a5acb15ebdc6fdfc2d61222a09b2669d
z70e9b62777872925a808666e86498892202e8bdba28ca8fe4487e952265653a2035e273d85afab
zddcbfb77c6505678c44c683e9baf8af7e6b82a0e4cf03bb6d0b5bac2c024f28d4cd95438076526
z81ec35709761d54151386d3f0bb8ba7f59ee2dafd0109411477b47833b7ae91a7ee836d0b5bc5d
z01fc7809e51a37e0b019b5f59e6510f109348b3dd99d60645333c90422b45dd7071a068e2fbd5b
z403f4cc4768b0dfc098ce2f5cdbf4e61aa4063760d5eec36f649db0c5070ea597c7158508658e6
zbb4eada1432e9ff4a2f158d4f80a4d10bc9171490ce7f15bff7e9502c877b99b6e1dc5e7d6836f
zcd814e9ce70463ecade6a4c0b08543dc6c87b28d142b44a311a6df05ca3776bf8385b00a95c74e
z88571434d1f0e290c9d6183bd638e4cd8f0c448b2af0bc2a4b4adc6bdedbccbb0f396ae8f48916
z41286b0fa6d8d6bdd3107d63cfd6e188cf89b3ca019789ee03cd7dfdd04863060837def9ed0d01
ze84814c04026d0ee90e469ec7c9765cbe7d87e5bf5840702cb99ea95b243fccfeecde7a537d4a0
zc09424b81fd5f792affedcb6fde94bff16d81c32eaf2a61264e0128011f83d646e4b4cbdc4631c
z19b525b0f9aa6e33b6bdcad06ded663a2ec23e43e7760afeb34f41be4629adc8d033f709df358c
z2fcb619a7d5acaa6eb299d23a33b95c5cf5f0a83dd6267b75f67ea3d58e53811bd1c12287b1a56
z1b7f622cb67259b98cce05c89c19ee95a70832be93efac65ba7c90246ffdc5ccdea8b6b3cd3eee
zf2344e7369f66884ec933a3ccffc05ab9ea2b7ad81755048c9765b3f898b9981f3c7153ce00769
z9b935fb1ac89f74449940bdaa998e88e97d75aaf118296b4676df4a1ce3ab858c4ebb3b3aa473e
z3b9faa2688f58f66395ea83766b48d3ba7ed1135eec1300e6a346e7a35281a54f4bd1244505c42
z9878b037cbb3c46ff468cf6b083c78deaa0eba279f3a2855dbc7d684f44d6562878c5a00fd6189
zf09f194317f97813c75e6df739cbc8d63b31d8a79f7f54f6ae700c7fb3e0dd5ed4b6e026acfef9
z4fbe2da2fcc219406d697359e1f0b375cbd583687cda05c04e85e6993f2bd6466dddafd883899f
z35201bf85626fc286a75c188ea0cc39e7e4b0a704ebfc1e795e0b8113ed81354df80b9d3a71439
z90ad07abf2cfab94e78dac7450ac6fd4bfb8eac0b3d2ea18c43f3ba4e20fc9983d048a1c3ee5e1
z56388f81e309b484a1759b7829e4e2333d70ce7af8ddd23c1d49e238b7cbc11b6318741f37d773
z857ec93ed40cab7301ec0f2db262a84f318f08661392e0a5f408ec5b7b37db79a0181775f6c26a
z47b1471cfd65afb9c9510a6016dbbf8cf35018b7fbc44346ab703310d7946030eabe2d2c19344d
z81542795f95c04fa91c8474b21a5b4149d6a701bda177b961dc13b366a506ccdfa84637229f701
zfd905c9a77ce3f1df69b3447b9426e8b5f55bfc3e8962bcbadfd9d0c98cd0f7b36d503519ce694
z55275bc6a7b5ff36b4834114f2e9e5a63504c136657b7e0d2f07c9d1f026545207328ea8641b3f
zb667e06d1d100a06d4bf3d9f089da88e8da5384da95f583f341225b12008a3f727304d4e68f0f4
z51249108b12aed6c75cc1cff3d0abf1adbd3486f73c27fc4c3845e11489849ff0719e7c392c5c1
z6906752a346f8a997b33b00e9eee78cbec88a189fe36209796688277ea7a82b376871d985fb826
z1c7c7a928aaba522f8428bde0f26660b69e175aecfe4011228f177818227ac3f30b982bdf47e94
zcda100ca7a4ec48674587e28cccc183df3f27fc0c8db7b40a27f8a29e0a86bc99a1b985fa5cd50
za22fa382f245f2b104a3a28548e37a5a8677a158209fe9d78b902ef05d48dc4edfa0efaafa5c5c
z2e90764ed2e276505b8621ee9c5bc5f885744a5bf3a51d495c4fa7d7a21fb52386712da3e6c306
z66884b5c037378e6fe46463f2948d7c3b496ec33f1c4c77a86228c515fc764d360f09850d8ee63
z1eb4d2af6b15710532eeea7d6328cdde7a1ac6178095370c44bd393819b98bdae95899937fe869
zebde0262735f485c50e6e51867bb7ee65013d0c94dba80436aa02672c97be79fead6d42e6d4122
z12798b26259d7133a7824c4ac9a6aa945a024be538281c1bad0bfd53574a1ab4af1f73cfecd695
za63620a789c32f20f1a1484323bb9e99539f7961fa54e27487f90a940d4cd6b952f96eb37531f6
z550311f357a4b193213297f2ab528c93eee16d68c73599176a63fca592fa861472e5bfd64349df
z7f4a0b1aab6c9d4202c59e85a6e626b2fe4b349ba3ec789c5e7510db95d0858c74ea731c4cf8d6
zf1ea275957e5e7098d5bbc4ca007552898b00f33a51556b40c73256d2a9769aa4068a4a898af30
zb63de516f52ee175a716f2f54de3949f029376b8a9cf1fec30075a476a5cbaf6b33daab1b67a13
z66da4e0b2a6f8bf85e911d43373db7df29fa8376f679e37009512f7cab12cd131dc0ee8a325a35
z8fc52d8df918f7d265b88f0a4914639166f4d121278c813f1763178e6307ce1d13fe84cf7d8450
z1294d72b40b4054dcb4cd0413b84e5a6b06271d30b942a65586ba29101f05660b025fb812ef7d4
z51c10848bdeba5f98f379280d817267dd6bf8d84c6c07111862e7239f74665d6763a0346719dd9
z3d80455dfcb68430e1cc9bb58508004af08991a6e65ff97e4ee846453209304a9e523633bbaa67
z6a401386ff1e7b7b211295f1037362b30a83492c10e1ac4b7e0ae7235320ab17a1922cc4428ccd
z8c8c916b57e3b3aa2c1bb32d9a156220e4050a60a5c5b8a46811c4113f6771a4b58fb6d7c27121
z976e05783516c9bb3a2268452e4698cc30b78746728fa24d2b693ab477fe77d3bfa512eb5ba1d9
z13f8963033d270c7fd84a18b4c9c72c0469bf333323aca4eff3dabcc6e5beb359f8dcb0cc39767
z008a86d6605089a27b3004908e7891c9fce9d4bdff7836e501bd53afcebea3ef97737d74ab796e
z8b97bb1a27245188d8dd6e55d99edfb1538ba293e6053110201756e8dc7d11a10ed40812d15adb
zb874011f7eccde224f732df2e08c9ea4897f8a383fabe95acdf0ca542db7ce8afe87c6b28f2bca
z20dbafc2569fbba84453de3f901225de3d59ee54ec80ecc601bafd10983643b967b1bd3a714b77
z059c98fdefe2ae674566137b1dabd8e84ea7013102e41c2e264ac48dd8f71f5cd261f6a2eba63d
zf391eb98ba64ea100b48dd06b71a90cfe826202215ab7a7a8394d8ddf3a31f4558728be6dad41f
z94e42c3f7c6bf1f8ca080240c1cf7457d6616dd795a5fe65f80b1c14f8706f5f21c324b9f3c7a1
z293c02547c5e83a925ac072ac3c44cbb360d4d69852cfa5a3ed9f3480e3fc8c0639ae8a33fdc9a
zeb1ff7705d2d26fcc3259ba1268e89e01d5c7881a13339bf93c9262856cd99f2b88dafb29d70ca
z92d2bcab8df3273b758c9f543df9cc8c4ac078f9de253c62758c7db76c1402e3d97e41e91e16de
z1c1a7b4dbdb1e8018150e2c4da9e8b1fb93f54235a0ee1aaaddc482c18d68755b64a0a4438e864
z8ac35324e66f9756009cc5cc0684e2228f081a59583d158329f24c17082571e2cef9302e1c39c7
z50af8d589c19c11249d8b3e2f5424da681a4527cb5fefdfb486d92045e2ab0250b861ff31afd1a
ze9dee1099018be88883acb3794ab6b0432445a5f0c620f2af8a7021527ae7a3da75945aa2bb6fe
z1a38c1fa5c65326ad54ef319126c04bee7fc93aceb2e0af5060d80881335fca85a7f80e2b46ba2
zaf35264b466d783038d3c3b3146a92d54c6212af9cbf6b8ef7aa9ac9651130107bc8412e7652ce
zd60bbfff70d48ddb520c981b5c36e09d45b94b5521dea91485b7218e80652568ead3c3f0d6b596
zafc66e66f23e488dbec65f5d17988476f464ef50a44bee2e112c421d0dcbcb4616b804da1ab5b7
z3bf659ab44f36eb968fb4ee6bc97b977f40984abe435c325a951b13c726db32d0ee20ad3bd06a0
z17765eacedaeb1457216b34513e090a39758c6b38d2a80b1a475e7180453cc6471d73d79e720ad
zb8deff3f34759667d2063c382569f15451a19b7364fc2ae08031f0df03637d0fae0500b28d50cc
zb77fa8921780c6c21adac8c65466f2ac09b47e28d7839be6f7602a7dd0ff112b86a7a0ccc2a30e
zc5cceec89869f5406f606f058b875dff90999ca35217c6d20768a680d3bf1e5059a822def257b6
z11f413bebd97095ddac4ab29a685ba30ba945fd0999ad6de4d8ba8003f73487254818a7f8d4b79
za93508bed6a222a9e5fe82e8a2075ac662de91e9185876a932243399331f824d27d3c30040b40a
zd7aae2ca880974d496f8069ed704e0a49cfebc63ed9fdf498849a655e080d13c2048fd343a1b3c
z7b2be51c3308fadc8e810d63890d92e8730a95d66f8f3ee847375e37808bdc2a701626f7204d9d
z82899b1679b58933587b82041e226612e45760b4e5f7ed065fb775986b82e72da1a4cb5fff6a24
z3607733bab9b722373fb0a8a8731452d9871717da08c6308de7ea4339a56c87dc4ba0778fd0ab0
z7729b60742a5260858177102310ecb10b5738aeb6a52189c6455439686d79ecbae6330f17ce07b
z307879d460271e9ca4bef5b04edc00d408820335a23ce8ea0545e13fc844d57932665c9fafedc8
z13801fa23718126dfb1bbc22e40824d5ed5b75d877a3da741fba087d3cb9217159f4ec067b32cd
z0b95cbbb66e48df202cdfd7b8c512bc8771946083a155f44787a1286c7df9cb84ae7c8b17ad4d5
z37b935e2fdaa63286c399ad4c460dc8f8e8d8d848597525527fb504caa61ab0833fb4f81d401ea
z99e99adfc97942ffaf9865a138e48b4e80391019e580765fe69e99dd6af6378b0d9b0f62d5e25e
zeb58a3e10d3db22c52475e0cd35dbe25ceb17b9b2bff48b442f4d5c66b7c91bc94965ff3981a36
z134dbdddff3e36b36a3b9f1a38a308505ccc7b01b75447cc94b93c29b561d863f6c5429d6117b3
z667016960aec58e88960f961eeea2f7b8fdf2981160d40e5fe572a9216ba7cdbee68c7a4812f21
z6780c1d24c09c506d3f5bffa8bfb307488de2d8f3fc6c096aa3ea2387240a451b1a567bc5a78cf
z12b5e6a59fd09d6b3eec44550f7ee969490421ca75ff8f6f73ab71f479c15580dc86716c524d00
zb209e198cba67be1345746ad1ed359af300b0596bd363388dbda717dd59ed3f5ba0d24bb21add6
z7eeee4750fdb9c7f3e95cc2b479320985367d36e32ee80f0028a3a543619031afd48a3dc468c21
zcb019cae0cc62300164d7d44359a7ccfa0d49dbe1b0d90b5be502c8890e5637af09bfac5245b00
z8b43295a5160d27bb3008ecd5cefac5eaf58b29b32b199f71c5d126d40654419f31177b9fb3c6f
zcfcb97ab1983c86e026f147dce7999fa4b22a869d3325fc8f118e06ba6409c3f6784aee9b38da2
z568504fa999f6969f5a4ab0fc0b1e56c0c269166aa6be9078055b7c790d5de17494fb029200dba
z9f20ca4cc3b0a933a8116f7cd668955f69c78163af74a801c0614980954b363d3001705cc4bcd7
zf387bbbc68a5790cb535b18615983843607d31fa91a25d8d9fe6e2ea036282ed4a887d068ffe81
zad3750c981c5daefea85ccae3fb191542c342b56805d8522cab70b15ac6e9f17740dc2c8e71551
za1e0e29f8ec2df996df702a175ebbb1e6d7a244a5dc4e1b3fae589e8621bdb9b56358c57d2d8e1
z95ed7b2b54c94f8e22f8285eca65d5eba472763836f5cbb613cc49320b585a8a9d84ce3f9e189a
z3ac3f1633b537c33af542f1599e283b884b8fa4f2698f24f77e279c6369e354ff8432affb988ed
ze8394fcdc3f9a5cfbb5fa67c96df5689f6d1a3748aee8cd15e0c27c766806d712329c04a98a345
zdaf513d77f4b9be817b7772fd35de730929f68824183f9b01c88a42b628979ef5fd21047b848ab
z4725826c1b95307fa0efd37d716f3fc4f180ac1bac2fbf4fa249b0eba2bd8dd488a8477aa25ea7
z8ffb3bb69b0116493c403d9d02aa0a0d9307a2e4ea953c83b83ccdb0d7e48937b166807accc467
zce909a1497b9612069e583272d27e1089856cc16a1de5e532280e0c5b85e8487ef7f30e28ab143
z237f3477aa746361543e74c3ea55ea69c11e20cabd8b7b8345f96f66095075544ed36ef8574861
zcca73667c0ebfb840dd5943d9766ee2314fa1f6bc2e753bbdc63562eb3e33ec227ca0e53690fbd
z49e59e32b59d13cfd94b5523ece11b71ff7dd443ef85f32d7165cbc818857d6037eedd5013e374
zc5eaa0f40995200cbebd43be0082887cd19d061add439ac212934e8eb604bbad7be872404688b3
z845cd06d85e73ad19fed7ca7ed4108be5744a8e48582c91a5e51b5fe403d2ed8b1dbae80a5e587
z775a83da5aae1d884cd9f6e0349ddb19eb3cc2c8ab5d86936fd0d3c121a8ce6a7db13eed3ca879
zdc4dcc1296fa2362ae7bfd46affcef543cca874e8f69684c23c9bf25546b07ea86de3953a53038
z2552df617c54a6307905481aec2a30eb5e2a23a35145522843d6ec64e1cb6361b0225dea1369cf
z52f3b3d70486909d7152d5862b0bbec9682e691b65a5b0f52dc4db8b4906c6fc95fcf63836b8a6
z23bc75bf18eefca945af0133503e916fd529b3ad529cbbbf829f01b23bbd93da86d4708366645a
z5af3e770618568ac41c99fa1c506574e53f7cb1506d54810e4499c6a936466ea975b7e520ae73b
z5b6422e3a96fdf2a8510c794c25d029f996885233b350eb1d92c61670ff955bb369893c1108305
z6725c903598dfeaa9276c24a48e0c25b006d31258784bc5975e8cde25c3f94d46d6278be2030a1
zc7ea668ed5852edceae8f62054ce78c6df2b45c0c4c63ed5ea9a30e41e40d193bbdb63c8eeda88
z50feb36f68d2830f8b70c961962200cdb4a083dc193daa0a88ad19f8226371e1de273b4803672e
z9b426100693023d442befefb927adb44d5accdc0b27b92815fb5f95fadeb13451960011f433e27
zbcdad65cb3111b67b012fcf5c2b92718ada17b42caf444b7ed1422816db395dc523069fa88216c
zabdc50f2fdb75b1a73d24bea193d940a90f727f48a7c8cf5fab9b60ab92f44baa1c1da05276a8b
zc4303538b4cffa2e3fa9773e0bcf952fe014e50e9c9d03a69717ccb4153b6be983dd53fa300811
z920850e74703122691396188dad18805d6b27c143f6322b9297b0fb35dd433a3a29f0a43699ef8
ze1de5a4d51686be168a8ddc83530e67430a042a4957075d51127603e0a988fa6bdb40c7c4cb093
z8296ef806580df70dd179a51b3989f87c551754477e0981b064e315fbf22e4e1db8b68a6ffb58a
z8e4be51a482f15b0ee02a06bee16b09a664213791ca73ecaf3be8906f5001cd07045d06347f954
zc30ef74914b066877fef6134fcabe05a810461ed605f6f0f2fd519f1eed1e8417403522aa2ece2
z628631bae0a574882d287a4f539bf8fe0cf20d1cc2520cb714ab82156ba2521383b9917ba33fb1
z2ac6b056220f5d7cc60759b9eedbad1606927a87ede97adbad98461eb86e1b06f820da1d3c329e
zc052680f77a775099165dc7701c7d64206192b7755d492197e58c58bebb08f760e1b2c6e7c8cc8
ze5255365b7990a6df0801fe9278d0fac1703853e08edd0a20e3d3b9dd555b620844cafc531c595
zf756fdddc5fb7165bb3decd177b633bffe3126db6ce017f9b1442787cdbad07fc7bafc39ae41ae
z419b1c80810435a7aeff34b2e564c9340a47ba52ed9fa79f018e9eb5ffd6714dd41f7ee03672a0
z2b0286ee56be8f35dd1acb086c8df16fdd2bb6c2f9cbd3e67b2d6f3888e688ab60852d4b319bd4
ze4930038a397932915c8cee2a549b16902d1473b5637f118b4f477c8a13835d34c40c48f7478f3
ze0d4451a0c5491a43a6928912c6d6533703e0c16d1c840b20918ec2ccb848a081bdf5a07f76b2a
zc5533969794224f3ae4bd176656dcb3dcb6a87cbfe209fdc01ed10a521a9c4a5ccde11d76bce11
z9ace9d682a6f391174d05cb8eaf6916f5f7c435033ec46ab3f62e82fba4c4411d8c0163ccfcc74
zb5964b8c4fe9eaf9ce07007dd27786b2c10a0165c0b2763ce7053039d709dd98a34041e99b4986
zc17b9d4dae944ca15179430a8465dddb81ab1e86515a3300151b65b7cdc770da862bd20b11dd71
ze01f417504b1dab316585945507f2a09c32d2c0ad16ee20b1e833bf683bf94ee9e68cd30547dc0
zb7a8098cc9f1e298c4d0ac7cb1e0866dec3a334ee927c7ab144c91e53458b12d927ddd3f15f28d
z11ed63008de69417d460429bd49d3e2cae5e11410b345825ebf9847585711176883590916fffc4
z34d1bd193dcf1f0f94e1892bda2fdfe4993bdc0a8600e374c7dfd701d922b653e4831ba51b1b48
z4ca3db4e8e5da207f3865251fb1d439e439afa7a4f25c2866535cf223eab4d8e3fe2920282f787
z24a7bc73e684d76f700cf2279155c05d761f0a2a2c4cbe88aad86a575d51ba89f322e5dbcbd2d8
z971a4bd66d2049a7b5a515adae836ed3a214872c7434f33343272b8f3be36f262f4da67ba6b3b3
z6568931db3a76cab7bc1cf4bfd86872071075c3e6cb574397af547ccfe2dc7752f32ea9b04e33a
z26fadb010e824bfdc4bf12d572505ea67486a96608ff0a4a78acac1518dc0bd849b8236bc51099
z9b00c1351f5c42f327ced4ace86bbff4ed90acc727fab792fb1bd972a60d9a0db39b2f96b10be2
z0b7487a4dd011d40a55e62f4a5a3cb13f8d7c9c5a554d1a3d0d840dfb0f159b30eaca44998308f
z16c07e57a2b79f9892d598dab6ef7053f6aac339001a891d0c20cc3d22df0f5fa094705350a103
z680b145feeb13e1f88e3d4eff0bce6fdf426538fae3712da109cea583d5deeb061803aff6033bc
z700457bd1115b755ce63a292e0efe5d78724358c7bd61cdfb5cf771793b5a9a1cd809e65093f9a
z4ec0128a00ad63ce89a4ab6ee6607b4b3f9378c5e980e69528f3dc65b000dbe24fa3b818ffca14
z532e2ba5b16665236fd549655b318f68a25740682b9abb7830dd64bbe2ab9f95477a4fde28da6c
z3312ec373ae19f96342a88a72285bd2cdf7125a07b4e0aeb50a89d01f583d26c88ec25cead7590
ze26b35944bee373b76ac4603b23f1d70088e8a0469a5c7e4c045eb9f098743e11f49a0f4e6057d
zd60c779dbfb7eb846c08ff84affc6921ad47c3da9017ba91ab12dbcfedd69b0c1a3458115b2c48
z0cb6af03864f454e3aad9d755e672ffe15e2b8f54ccc4c1775faba7361142f78d6839d8d42f8ab
zb6a4bb7da16d9c7a7e463f0ca7385ffe63394ebc3f6f122e77d60e71a9ac99585500d47d2887c9
zf678e906448a7815798b55550d809ec0ed7bcd4a728dd83c1048a2a321f68e9b3e2ef5932c17c2
z380bb225e842191a02230f6a7a846a1e3f3cfa63c9b4276afc4751734d85a11c45a38f12e5b8a6
z74d56c8714735c6a82cf5e6eb5f138275b6034a157ff89bea2697a06a4ff2faa841ce951dd9c53
z55a07b27a94d114a5284c3afddb4e3319a7cd71ec7c8087385f97e1e67eee4a9a687b8e9b137c3
z43ad70b7f2e03e14fc74ca8563016ae0b7769c85749a9020f95f5f07b28ca953438eac5680f014
z5ba9a93244f8eb062187ceaee4d4cbb2ac74e93794d735f5c382e343dac61b9091a3e3d3fab94b
za47be8a8f6548d32a13a9e4f39dedac7118d34801d07355e80044397b264a80dca7b91e1da56ee
zbc435e88f92fe9b0d0dad46bd90ed97b6d804262298581abf9619e5ff8a6cf18fd2b48503f2a63
z3cc47692babe074f40142eec1b6a72080d9a2649e956f6906540945f750daab28e773d9f5b186c
zd3e82ca404b77051c30d8250d201405193fe9850d8b744335e900596dcf92e9ae18b464d19344d
z8a3d1114cbd42d860ba90940b3420594c2e0171df72e0f8f82e365b8e04e26c496eb5300850e5e
ze8fbaf421b9a1d5ab4332845408165376291d78b505096afa794e521cb28cdd1d41c96524669da
z64f4ed60973082e6c8888342882d9591383ba1a11a3eba313ae4462858d01925d8cd47b76c05b9
z3eb23751127437951d06b9004358453081697f0f792d7766e4ba4e4a8315ab603787694efeac62
zbb1d8e993c82252ebd865adea24a12e9878aba2b8a36bf131876c8befc86959b56672f6b46a369
z1f37f0aa9d9e7b3e4f7a29d6878f178076c209b0d62ed901d3cd7497863b9094753599b6d5881b
z8d6b15bafc89cfc4d25d55fe27b380376b1e3cbecab3edeec1c0682e5c9f18af251c109d6e0f18
zd4213d3fc9e2b2c97e7adf8cc6a7d6927caef4ba01a46b014944d635f6fc5bc76cd286905eeb18
z6bc743a5ac66d9bc24895d70fb06ad764696ef088cb43f2ac1cfd57e01ae6da6754cb0d6f36e77
z8f750bc31d1f673319f75c1e6d83bd8d99c88ad8658d35b7feaf0689a10d891cca3cd4dfedbc05
z84a738defbbb48352fc3c9ca0c0a39c9f7cfda9e8adc3e683d496b30b965d77c51764916abed1f
zcaa0eeb72461aeb9b6e723caa9936b4c5ad1cd93c6587a19c9c6b720579cce0e39fa6900c3b23c
zcb091d6e6f16b7e2f0bfbb577e10dc304944fbb9c383cc92c4a17f829fb7dc15bc305f1719efc9
z3e4f5a885069c02489155d4f86a8a9b4595d5a1bd9c83ff1b556a74c28eca928b8ee58ed554d17
z48f93e36a5218b96a99fea763b202ca78f46b9335d8b79c2ffc2d1f1c787ea23edf2e63376bee3
z3a6d7176df0cb0408feda070cd4b5f1ab5ab0e17980cd76bc3f975990389e9e13452479d53e7ac
z320123663085d2b3d2adc05c233204f10d95163a08da5f3d83fc57fbfa7a9d50dbf8907a070775
zbb10acce0b39bfec5cdfcc92aaa73ff1ea80c86c693d1e3b1271a4289519310502d430fa0e68a4
z6dacfbd598ec9c0d5694bcb9435e04d16db42f8da1c41a47d5c0b30147a1b80a036f99d8a6c52f
zed21f1f5754c286a195a0b9e17031060deda4c84832a631b4048b26337c57f8321cd4557e624ba
zd0de0564c117bf486e2b614d34eb7c044440eda4765d27f3f459398c0f6873ee425341618924e4
z6217f2b8622122269be559f8bd4b1118eb4865ea0ad89a9487e08a896d828db175dce764e570fc
zd3ad6d78d2d4ca2ec5d2473d518905bc3ec34460c14ed55dd66388ca7dfdd76ad30ccff3ee78b9
za17b63327943e22029f60131fcbf0c0f765f3c8e7df6db782e312c047950705b7c8a131215fcc5
zde214882bb92579df09fb71dad08f8b414731fb1a3c68583fc8cb276fd0d882c0f47c1d1bfa70a
z7f7f77bf57487c058747a6d2971900204a4e2f00668984caaadeb37f17dd30155725abf5895c84
z33e5de0da101320757cdc3bd1428e490076fb2f900880244f01b451619a104fbb7e8bf90033d8f
z12dc54fe1f2e120e8ba40cc700e32c4fdc4c6e52eafc1af2ebe618d8eb14d0f65a6697ee47ecf3
z088b92b4e2debfa53b7bab028bbcad8225b4f713f9c6e07469edc3a1a33271009e58723ef465e8
z3ddcabae1fb08759855fc71d7117f9830d6259be9759113fd2130935803458b05c7197ca340762
z50ecbd1b4b4210a99ea9897544141d4570d34bcac2efe12cceceade29b865a864365e965c7a353
z5973129fb80c55f8195574a7df0540310bd72b328526042483b095bc5beb178af74ae9e7942e3e
zc646fbe4ceb1b9ef6d19e761262c7775b29a17c459dfbcf6c6beebb1a91ab006d856b3df249c40
zfc0b43ddd8079f762d51c599f3ef270988233f9365581d53076acb2380eb5741e2a619846e4ff9
z265f067bf1098d00f6da11dd4cf2a009586fb272138451c56734f4299e09c81b24eddaecd264c9
z2470a320e42f8121f3ae3534f1c70b5f074f54851673fd819912b300be146eef1b9236eb2ca36a
z6a0226f92f9727767613c705d984d4a2cc42439fbd015ab4de22cbfbdbc54b8cddd6609e20060c
z4fecaeb1a823bb58f9d323a0ce8984f5be4a826d6553d19dca47abd30ce154cdc90c4bfe7e0370
z591a44ea0b21f47eb7407b6c3a8b4eab4f284938e58dfcf380c6f247330cfa72c1ecae0ce40819
zba76693f82214f122bf3a5a4734f04f7e379d54a5b0fbe292898cf8ca432f08c473a93748be23c
zbebc8a9d39511e761e8df902fa370f5c8ecf219d58428daf9498b41ca529c9d3ebe2ca7736f81c
zd28901edb22128776e48b05b771899c6e132c1cb5db34352f2358d32a93ec147a9ffa0cc147d6d
z1909607f07b05b1d7c6017d3aa4e7f5a70b9cc80249da9fb7288c87d8df4eabff4d6a8a3c56c3b
z43356aefb4017c890b48fd37d30251757d28ab17ab7af3c627a19041a530a7c070042a711461c9
z6a47b70260f226e18fd7b60bb21bc74405f743ade101b67598ae41c1dc436bc14ad9ab9dc9134c
zde054dd335632f71db052135725c9134c5e6c0d6d8eaf78c5d674c52ab240dffd5b6e3991b42be
z6e13b5aee745e87b1189963d676a0c8713d77f406e70a8fb3d00a1ded617a156d6b5ef9b5cbd96
zc201c6fc7b5461f1561a16cd7fc9e1d00a557367226fdea71c6d4e196e19c34ead524650f5b9f3
zf628ee85f488d9690a00bab05ead7cac3e5dce6b4fe190d612d3dee088ede363b66c70caf90c64
z045936808912af745924686dc8a01076cb25104007e2235880b9945a17ff01510d6c1932dcc6b1
ze806e6972e05fea0b02fd5035344446bb0191279ce3f5953eeb948f0733606f95d3af3e1e167c7
zde38d4bf2e2e147d5edb57202bab237637f57699efda4c07c9fda019dce71a6c200ad17b897d06
zdcfa73b41d5c01fc558678312d24ba21956d1ef333c240f67c5b9a2466a8025cb5968c5ed891ba
z0e56f1e83105593a57eebc0d765a65e03412ff36be0bd36664ea2c11d08f0536b973e552e4d9a5
zc84c23394a6bdf9f2a83f53e1696682f19310681016534a8be17ae9fef03052960a68d5eb5db73
z456bc70e53388c297712871077c7c879d97ddaf3edd977630e74628788cd2098029acec663b18d
z1be28349734491c752807fe4afd023e316fa586ac1ce1cac707c7dee752557e6225925e883ec4d
z38f0247d53b7db3ca80f18fc1dac11efad64f07c252b9e453c53a354c246139e59293da930f075
zfb004c7d75f4b37f9d03deb1fcab61d2e3e20ea6a15ca01f57a41fdfd7dcc622ee3442cadcac08
z1fb50fcad4256452d7dd69ecd7c03780c9e5916975b6a8b39af2c35d1b57e17238f44982006dd4
zbaaf86990330dcc242b97c1f11df46f5021ac69a5dbc15ad7db95f9dcef58862d975713136c0a2
za1b5b40d667b75f6c2c08665e625ce4b9fa868e9d8043e19d6e0ad974df907b47975b7db2acc69
z50bfe7a74333675110959ef54c7b7fd029b46fc8d729c5331825d912be7fd959f9c9120c96729a
z1f841378e5aa3946b2c1ef9eb0b5261ef8a966616362cb969284b7900a2f906e617b2e4244b11b
z27887b081601bd06fc413205f64056efa357e507dce4f7f332709f82f9b82c21667eabb063a19e
z1acd4d16cc8c2503207a3106f70b89aec69e3861dc64b161c5339699650461fd4235f12d7e507e
ze529bd5189e1b311c330604ee16f4dda0e7fa77eec75bc3d95817ee99ce88c3f157da69cd7124e
zbfd94cc63f8c185df837355f542f16a61d84fb4934f9445a272562ab02f5715106257315b0475a
ze0f5ae0ef0147ae3191a01385b47c9352f0af0567a87f44493812ae5d94ec6d4d8e25cb9b6feb5
zb83c543e228e6e4189fc4d29eaabcb3b28e0736e464267d26cd38f88195c25418cbf3674e60c63
za22c2d1154f4efadacf424f3247a2e3effcfb985db8c4148cdda86684e9fee549f9dcdb12c90b4
zf882c6bc28e8de0e4ea2efb0a0e73c05637d037be620651e3d4a798c5baea78411ea2762e22e9a
z4985288511ed9b012ce06339bcf43b23acadef20a529b649d0e786c0009099308a89af857dbe9e
zd6c753f38bbf1fb8e198fe8c275412d3407201a295af4be397d90d4d5ef8a1142e4efbab0029a0
zeaf03313beef2b3bca4e370d3cc076f8577e3b40f871aa3e6ab58dee09cb75f6de1a32d1ea48ef
z2cdcd315e38c55a718561f15984704068752c8cffc009ea62e99043e61f4072a908344c5a25b91
z932ee8bd72d4e4c00cb5e687cf5bfbf7dfc020ba83b240733be05dcee2dc52816b6ef1f22cfe8e
z0ca3cc9d4ba1c160692752d45975ff16ff0641e0bde0e08928435b2e01c9b89427d21a47031ff5
z999223027fe60f25cc525780232fec2ec126db1cc105a601c530bbefafa3ba7e4f75f960bfee78
z3a19f317bc74cda56317047807385a06c6d2db4e7ad03f8c39a8c5266222f328c8e6327d90b7fc
z6f83d7e8a45c97e2dbdbac4454b20cf41940cd8d19d47ebf384fb98ab5fe332fcba081609e0161
z43bd6f43e3baf5f1a6b22e4fc619dc755948e26408a46b467c16048192ecb7e7b2afb50cf11f86
zc7a7104b8e86d235db44055fd44537e8bf79fbffa03573f4a38ce907dd2e690b7f4f91269173ae
z53ad21b64d9df76221b9909baac60b83344b1cda1e232f4526f0485d721a37d194850f5f82f180
za9a061b879a82fa24168d68d47a7b888661ed46842b92da5fd802b951809603310355521238fe6
z010fc36382b8247498d21af6b228a492842d4df6e0cf6b6e65a57e1e0b3369418487120564f2ee
z979cf14d84ed2e955cb85b31810f8972c5815cffec33dfceb48d16fb66a3b7496a74fc24f1de6c
zaf2cb9567e7533615c727125c0ef3fa8b62e8e9583b5fe922ae857d62d405d1cf579a76ea8f771
z1a406c4cd088715d0a9fb1dd9a73c49aa23b17bcb81ded3d2663abda410c3ce4af0f3738e4b8e9
z224a13034c33a5203c03dfc5396a513761866384e53a8ae9b49cce442dd2d6e814b3b24ce61415
z195d4402bdf679cd1f6ac7b7c3c6ab35f09d156e66ab953576c6e12556c005ffe413f4b527a5c6
z98873c95cbb4630ba4529974330a2931c8bfb6106df6092ad91cd9c9e6cbbcd366cb88c0b1c178
ze1a59cd2c8aeebdc814a228b36702782b268e6af3121994d4433f9f6fe1b4acb8bd1bf8bb686bc
z74949d6de26c4130bbeb573c6ba3162350386b2ecf1e1c16237a32e2230c5fe2a3a40d5668e032
z78238f7e0cc6157b473408474cc2dec71b534dcabc277f9225c1957493f452487cedcec0d9711b
za9704c490af85b048b18a4bf3dd0fccf131530fa48730bb3ca0cc0e8be75abb645355e4546c28a
z4f6cc46de4962df08fa9612594226ebf1bc3025ebc3bdbb96c269fc124039e5ab769660c718efc
z62a5a07899f9c6b4b7a5f8ba19eeae030f64cd4c3de9942acbf32cbd8e3a6293812b3ad0f0015a
zf17eae95dfe0c84fea656f3bd97a98749d42798239fda5b727fc6bb2a88c030cc5945525d52a8b
z0569493c8e6bc2059c71ae56805945412c3eb616da288b25d215158092d85772fed8386184bf70
zb182c0d3f55a45183b32d6cf45dd1110a0c212fdb317147691456a10521700d8f44a0f535d64f1
z477b71b41725f7f96a08bbd6cbca654daa52b5cea8e36dd1be5000bd3d10569151ed2e134c8b96
z1f4d9527737fe6ddf7833e9dde6bdf9f3bc8ec5eda4d15fc37ee08863f5bf55e638c307de602ac
z7a37d58cb42e2d6c1ccecc37c6b56883f1e1d7e171766544681435969ef9ccc15e6f9807333dd5
z04cce216af9aeff359e9fcef9c24ba9965ac11ec98117d9842c04ea54095c69e0a7ce7e5fb7ebf
z7d5209cfb0c317547047a96bf601afa4e3900a1dcab6749cf05dc7d4ac807b86b0b35b53a3ff93
z6344c79350cff3bcc9f507d37ae2b91077b081f2486758d3c75d6188798eb9089c162a24c2fc79
zd8bbb750ef74954b2952c9c65df4eb4b781428b227cb9170d99f6c239e2a2af135c1295e78b046
z5cd011000d91dddc320dde7104a64000ba94ca36802c586d2013219be542aff5a0f983633cf1c2
zf88ea338433440cd5e5b18a10e07e00c69d4284b52d1597eaa13baace5844f6fc96b7e68aa9d40
zd7f63767a412cd9c8449b59cf65fd3c500fc521f2e741149bf8f70625ada0d1495762f0a650772
z99f85eb9bc0c37424e9ca381b74160b03a33e642b078b9fb94a42b5124765c3f54630ef471d33c
z4a84a91a014e904c963c88755428a697d7cd4803007bb34fd9b95fcf82f45da97ecf08524b2351
z06f640ce610d0d99278ade35bfd5caa6199092e00cde99cd3a8c6799bcd10ae3c750606f8f88f9
z1af7989893e525102e422a54ac623479e75e0d6b95f7be26ab784d2d61359ddf3db769d9167f72
zb1d3778ef71e8dc8accbff80aba2658c69e4736c3ac8bdbe90b3921ada9b08fd433c8ca3aa58df
z71aa4487a562e0038bb958c28a01a14b5b44e528e533f5e6fea1674c7d71ad7c0a88e80d766fab
z00a09f7d81d118fa074c5025874b5faef76f2b249b98ff2f58de805133f14d8d9fa7ab5cbde8a9
z455296ee8c989cff9df457ba24f842cb0d00ea6d19720af41d03cf25be41786ef199ef40dc8873
z8eba493d9829f5725205c1e8bf7f09d7f2fc0d0b1db3c6bb150784afc7b398931d081fbea08a69
zeed5aa05fa08d8cc5cab19eb1b3df78f2f53e0e8aaef2dcafdc758dd90e3000150ee073ae9c97e
zfc2a6fca0cc1fc94ee6b819076320e5103bb31c7223c24623a6c769e4bdd883a6aac99aed04e34
z9e0641d9737000236b739a0b2324c8ef5ab5bbe0fbd25222df045ee94c6de993f7c7745e2209f6
zdcf3587d52e4870b497d099b9a84d9ad63c6e871b4761f850ac636469a55da82cef275d95e08e0
zbcee737168582c611ddc6cb02b9c78664672e067b114bdff3a4ad2fc1c3e3d1c5e25183b119c48
z4970278cb965f928d66a1e97c0492b6e68c74f4a00f2e8f9b685d062b3377bcb8e8959c6c57a2a
zefdfcf5b3412d1494b3193b50758b43569f4e5f5dde104275db3833d281570b31a32cde9cd8177
z3d13775d0bc8eb8ec88fb042b3944db8d433b8f8a497f8678f88487fed841c70870ab4d7e719b9
zf45ad8a085822047291b6e59daab931e341c06fc45f9b56b6be7cf562ef5fbbed299072ab33072
z47361d6c73144fc8d069ca79e755b146fbfdeb9f1fb6f050353e1f3d15e5ae240cb99291980ff6
z9ef7ff14f827cb454a8e4744c92547d7025733031043b76e34de6510ef3a44ae94a9b8b79db20c
zb7a4265df7677011eca198a6161e49f56a10f953ef46ad50118c3b9cd532522ace3e53e50564ed
z3317df547107d1f9d20b8187869012edefa321d16c993fd65865fda32d4313ecaa3ddcd2763f32
za8b7eefe3723dad16e3bbe0a8f608883ac277b9223cb06152d62fc0448af544e73e22ddf6ae55f
za1a515cb3dc0c54d2c1d917512bbec3c3946865f92c9aadd81a2c0cdaf308d0f019bbadc2b2e13
z38835fe0bda354a1cb26931df0c6f61a98f1d39efff5f3a70b191df08f88384ee556e564f0acf1
za28ed052b566b473156728dc421298e8cf913f6c95817b485698655fbcbb73a08cd63170b005ab
za6b7d4c4783bf60033ad60f0376287fa8af639a11e91169869985671475eb694d0691e5f47db03
z79a95987ec7a5fafbef60bfefa3699cca5519c1302e02e6c2dcd6116aef7dc13d6c894e068a33e
z253fc6314e26634c7d081e36f0405706a007cbf2ca2a5fb8865ee1c7067114055d80bd4e8297bc
z1eb350dd527f3b2623edb960a7da4d520861e1da84c4e0aa46ea05825414098329c1245b4b7647
z7a4bb0b2c299496432e0b9b87b5dc50d62e80dff7c1071bc83e1e6b8faa724a75d68a0d1111503
zf5878be59a51401bca8d8bab8485de48655b9f8751fbf436f191ca8bc598af87d359cf3065a07d
za4a20f50cc741797f392be4e8ae56c7f075e23b3bd77fe02c89c5dd9a158f3b6c95802be126fa4
zb0a2ae38869f6c9cbe944ec4fd365b7a26136d1dda43f08a0628c520ae07061ec9ba4e673b85a0
z8dc4f7930d76c2fe5576c4b6a3e95434e42e1083b9fa6ea08e44d9b62f8c54801e11efa1616fb2
zf754aeb2e62ec965b6733559bd8bc1d346bb5d30f1b664efd7ee957bd0f37843c688f0a98dccba
z86d9492a64583487ef620bb5e29165749655aaf7d33538b2389981c8cb5457357ef174db3e9e63
z146f3f2db4e9f526d823e139844a8696c5af65fdd743dd1116e5ef27d8f3ad12d2ef2f29872a00
zdccc8fef2131c660ef8d73c3933fd9823a7dd1454b0f1f0cdd459c12f2bfa49742d8088a6297b9
z2d8c98556519f914b16554f3b5bc8cd130595c73e5f36fbb6c2299c23a47e350e12c22ac2cc59d
zb8757b531b8b9b589804f4d15f7467b3c57b7c110d2a92e6ea790a2c307480e3b3f5411e3830c9
za78f7b4cdb4914c93e956b63b764b2b87b5980049b607bada46ec707463508bdb2fe4fc70dddbb
z4bbd722a4e45d66d528a80111116398f4aacb938794ac14a3dec9c3e1ad9a29af5d4941146f48b
z2ac2d12f870b18e16eab7a02471b33ecfa777600c07c71d9c13167b40f312d494181eaf893ec3a
zeca22c9d0493f3eb94684e5ad592dd716f7e7d019c6101e8259e81ac112b1bba9c1536e0122062
zac13c42aca6c972eedbf72f5b9520b7fd21e4b169269c203b1331e92feb76e00690f52d644dcb8
za1258250092bb300f04243d909b9fad97e90a20e7aa2da4ea31817cf9436cd53074a16ddff1202
z8df0f6bb8a81af2043138945ee93689a3aaa3b4e75b9342476ec50c56f6d7d082239f51a3c650f
zd15c3d6f3de6ddb58a1471dfbb98cb9ee85692a9157015b83bfc53f8c9fcf746b9c261c2744060
zb0e641b7216f214806593202dc2820c882e893cae9345645b454e0c1672950c16f9f47620241a8
z5a0d8e1756df374a23f4f589b7e9cc0a0dd5c696ea87ded7b31b117c5c90239505ce5bfdf071c9
zf3a4a5ad439b396aa598b260388206359e80d634bfdaca140aa210bc18cc9a9713d814dc9a9ffa
z746f915ab96af34279681ece4a9dbecefccd1da719886979c6c0ee19a292828886bf6894d3180e
z0d82018c24b4ebd08a2293605465d2cd87fadda3eff89b7e53ea5a3109745e70baf6c51a6a3041
zbe14ccc4975f419c6b4f68dcf91f23e0f035b597484c75d764a3efbae670175b5be735732f8099
z69675ea66accf7be953097ab8b5fa001b006d63cc9e63cc7edc89b9b47f27bea15a92ce0869c2f
z62773030612a5d13f5145260c3f186cad7123835a9f3b4cc8aaefc2a7d2aecde5cf9e8815c65a7
z6c3c8ad849169787a0f01ebf3a5ddc770a77297826f718dfd99c6506c458a964a0fbbe7c5d15b8
z007d244dd41cf0b005c9fe7f8f45c50ab81155bd982001972c8ea57a37c40cf5c5e0226bd86570
z1901f6ec7cddb5236a58ad706a2d70c639650bdd35bfc7bf4f0b2fa347c1a6af0876193e2ce47a
zf595bb9b5d83a3eb01d87a08979dfd223efae47848c648c415108ba7262eebe94d9afc6660a376
za05739f3e42cf91f34c3224ed97c61c09aec10e0d1438118b5f4b84f44f17027f4c9524ec9d6ca
z19222293cfdf30a8c000f2c8b741dd7ac75332d8e3b3ca317ec5a3e9c665008c3555e0587b21ed
zf75909e335aeb6b293313ee3b69a2354988f73fac323c490e742ef2c03f36dc7212a1742828c1a
z2642c9e8912debf3a147532a7c7eca0ab7407615ec62eea3caeef0654e3fafce03d247b3b76389
z441af68c0a11fdd91f6e8f07583dd4bfefaaa141a94edd27ffe6ef281995a87b528fdc1a6299c8
zc794cc898b545ee2a90e6f600fca403477c29cc455a67b229ea864e453f53197384ba68fd8451d
z0a417ff4730dec87b276f65981a05f67359530ec0d9d4cb2d52929c25cd91e36e03da64f4112cb
z1420f246102fa0b807246c959749d08f1a3d9efe7cf652ac955af2cb0739b0b4f50078f703a1f5
zfb79da258b124eab8745dd2200d8d81e4690ccc47d8a26dc4441fcb2423ac4591f1828621a91c3
z351244f233be9e0d7621aa58a893a158020029b9250f5626da7e2021812ecf5690a16ab5756a01
z0c404d82e7b38557e59ea48dc23416c1c0941d994bff7e2b981018d686f7b17f48a29257660317
z9ec1c00e09759353b50860539321c326ca283ae407318c2d38b858561c8cf2c466f698047816df
zedc4579cec1f4084b895fc564bc545abc5667e93e8275ad7727228a95685ce98cda2f5883ae4b4
z0c30cc73ab2ede769e8b0b60b5ee295e11d50d381e4c2b810d1fec93baf60af56fcae7772ad7ba
z34bf0e367a073622c0e11b02db83954f69662823ae653c26007e2f53adf9c582e44ba734962871
zd3aaec2801b1068c1471e9773ff378587660392740981f8a2042a1f0b157c07d9babfdfb390383
z982e8ff61555b28dd49d57b1d916d8130409cfd150d7b4dc723a809da0736ba0bb618e445ca58c
z168d35d08233ad46128153803ff9385df10d3495671055ddbd3cfdba0ac5aff39c9ef23a7794db
zdfbbfc49cc18d3d6f9ff2a4a68e4499d333f2475275bd8f890a73079396eff75a1ea79f9369c06
zed653be511ac9a7f1e7cd0ecd846dfc95db57cc2568daec077e69f12c1c291290d599150598fc4
ze7e4cba9274a19b440e7162803c8e5d41175ae457375595624b1d0a095e5011aa6555d32ee21a9
zb6871c58e9bb5d64860e94f3c3cf45681a2a8031bff8da2038ca0fff6ab2490357621a99fde27c
z9d991b7eb99ac4326ad4344d2d24546d186d8e6b17e05eb1cb15aa4a033ff718c2a530d1983c23
z0f04dffc82e34ba4720be7eec834e819eed2d6aa4a02dd8dbfcf53dde143f76046d0cbc0f58274
z1b7dd3e36bea7dba6f078b0aab748f89a412e26e712824d4a9c407f2cbfb6d8675e229e921a6a6
zbd4ef2f4f82221dbd96d1700d374435408d72742ab8281069fe007feab8a7683525f66dcadc907
z940a7f012fbc350b403531233da3c72377a9f363d720bf9422fd94a2c251d881293c125c7ba207
z86f23cb637ccfd885e58ac755da4c84dec61970fcca43c6bba3ab2fa3b8f089752113b61b2544a
zeac61c68aebd90897184917d1df54edc2640ddf4a152505ecf2ddae58b5dd8cd3615b5bbb6bc0a
zdf8387b50380c88b8ebda54f07efc4f72b921ea7bc3d961f9deb09aa31935ca00ef0c689432138
ze944eeb75432a703b7e90cfb587066bee42035399de590a6f3ab5cda5774405c344b8cf6adc482
zfc378007a3be2a282b40333342dbed445955ad9f47b109121318eeaf617eec3b27f21ef9672501
z456ed7f31ffa4306d09746eaa2c3a8695cfe975caa974e43c591df8a48d8e8df8db05b8a9b6f08
z4c6c9af3366dbcfef89de0514c720fa8ee7ccacba1776a64bdea305ba968b36f8a40aaf5f4e356
z20477d1d95ad420747ffea311d5a876332a8650921952663cceff03c33e02c48989096a6cc939d
z2a0754d4d6f41c523d276f2c0bcd1518cafde3a74b1da948a97dfd56cd88ae4b6ed0422f783e57
zd97ea570b3ab5d92672e812e3315cc530192f63e613a5127f432536b4ef2453e9a2860a7d9b3dc
z592a2c676ac035104bd2aed4b34a747ea809703101c8c2e4b2efa61c04f11453e73d2786d5a398
zde5d5ef840f4e8c5e62842fa21efcfe1829026519fdfe6f3dce14b78a46a411469d5d6148ca67d
z1b982cf558ac834239356bf1510304fba31d1805a02273970d040f34f345104b8517105f29db72
z0492155cabe2592068f561892ea75121cfd12cccb166ad1e9b0f1859402618cbd8813828888791
zb83a13937e396fb812fd1361459a6e5b263182b864d690bb520983f7a8443033a2fdd7a45cea5b
z6ebe85e51bb5844719a8dc52d1bbef18d7b86652bfccfe28049820e29b697a5b1945564ee3e2dc
zfe923c76b9d91bd12318716abb7ad274afb3028da4036d7923e867c40125e714deb666fd40d7ad
z5055c7ff39dd941da7136f183cd0ead10d23d3ba87d10d0284a2936d1e5ebf3298c7d98e8b5b11
ze43d82829b9ab66159981660347880d8d40529379cb40a1cb1d0097f0352a757366ea97cc74353
zcfc919b5b4cb961d0ff51ed364b895c92a30479c052fdbd23ea23536d6d5d94da6689bcb0da790
z74ee56a85611c5daf4e7d85a843165689a2b9ced27a31c377f4040424d4250d3a8c87b41cd71fc
z68346cc07221ad0df4c3933e3093c2eb79d806a40065dc70c564c2dd511ddc5eec9bd618c9622c
z91e7644883475cbc1c88d41179d70183f733759bdacd0e88dfb4334b198addf6c971c5c33d0b69
zf4c42d72a7a0e3cc7618e1f7a169689fa5ff81d1ed145c048536b566679a6d4bb2dff79febcfdc
z056b139f52d05095af77a92babfd8922dfafac8c73f331c6e5959e54c61bcaf48fd37b9d1d3eef
z358fab15e96768faf88ddfde345eca7352b39201616d5c1643325e8adc3359cd4035d0198f38bd
zbb9b19e5f7c41731f0b359e03c597304e75d9fb7b5e675cd85151008f8dbb902f62b3ae629dd81
z4d9738113175fd3b188b23eb03eb25129ef6d296f82802270d0777b9109a8c8e54cf77c8de597a
z0f7fbdb0b1917112a2b9d910edbba95a4d25902f224897c45b929e5e56a2819210250dcf460a47
zd1bf05702848175deee31db88f2238377524cf967b2a04eb58eccafa6f706aa6512f9e6142fa5f
ze6033b3872ef44f5a4d7815f649a4148854d9e78a576469a24163a8b61b50205a303dee1b897ea
z42b1f99ee2c193890833437f139a46927404a3f6d17cb2d1f03ffee0a5086ebf497ddd20d29987
z561cc31b08379a05b883a29b8e210ba1da6eac389aa883ff6f84598febe4bbe660f6adb1ac6a58
zc72ca385ffc632daceef0c7fd367a02df9cfee21ee32dbd89fa0c6366203c66fe6c90cd0c5dde5
z9a89820c478937bda5791e8c2b2eb0ebd6af980fe10ce39b1097bdec9a926b9f1580cde16fef23
z60042415fbd59ac538dcad2e97fed47a6a11d558e9eb7c9e36f6058619b0a5f27643b1fd4817d0
z7e4823871d5ed49c45865e0c8b7bb72b42e78d7ad88ee5a607c2fc77274f1b19e63da36a297766
z00784602451571c52b11791d2553fcbb9785d58b2b6652093cf60f7b88a6b25c11c3638a309c1b
zcf0ca913c7da20a348d7cd52634bda053e9098b79770037943b63de0abcf171f0b98d18cec03c6
z02547ef5a01edf1757576200cef3109b69679028b14b60a29502603a790a65153cc3f287845f71
z5618603aa8f24c25da3c130e3c11d478dcca571674b7470e03be29df37585396ea19d13f8b4015
z96ac50be6546d7ec34e20f1159648ff805dab156d42c45a6ca4b23ed189fafb537c0b1091f18d3
z303998ac97ffe3d577e1c745ef536780c4aca45cfcdef8bef8473d13c21e19746ed8ab6a38fa8c
z2fda91efd10dba2e93901a2e8d6c4fd05e2c59d8d99e665e8327e287ea8747977ad0b15d644a02
z5b9de9acef7eb707d42c0c204ef9f2d5f60e8ad3e76b4571ed99d05657c039910e0a0bcd735a3f
z52f9afd849a8255c137820a697a11631bce5eaa53d7a609af0c215b26d1b4f03c357102c627798
z0ff850d1f7397ec642332250fa55a09591f3bf00fca72556f508d0d196334835e79a232d841a71
ze2900df3885814e705a85991a38ecceec182ebf611db7c37e4658da0f793b9f7dc7d20df140aa5
ze547a9f3358b800cb4603626b16f215e85c31dc179ce1f1e5dbed78f5c5f5f0094eed93a532ff3
z59931b60b7cca86a5ad43e52ec7ca50e745323eda77f98b7c16c12a5123cec487360e4df790ec4
z68e4fdaad625a4c49236f9164db7f254c4c0f4d0280fda7a670a211755b6a52cf412a62ec60221
z65aa46dcbe38949ec74e2ac53efa466e1aef47db917ab7bdcdc669974e18afadfedee768ece261
za00ec99ee49ae4981be5b1a7c92883dc0daae823c301556ac1783ba4f1cfeaf0760d6bafbebb59
z8cf14919fc4dfa1aa0ff64f14ffef4c22e61f8a0badc1fbfe96f6004921c9a897432434db0a36d
zfcd132990e4d50a8d126bd38ffa9ef7d54a1aa5502ada1edddf6e7f1898269a3948b426077e2b5
z227159e7295b799e9ab426c2230b4a343210f6ac5a6610cc9df9353a9c94bb1b4426324accfe5b
zd3e50c37e022f739b4854aa03659fbbacc409a74a12da31e3bd2452b44a5e7b27bd02271881478
z5f9e9e47a773d27c3402a6c22cbb460a4b6cfbdd9e0cc72dab97e42dd1b8b963f24d25dfc8ed0c
z97ff8d8bfc9d1c0e69de70442957b886b1fa96d20b64b2b91d14b383de5afcf750eee1f9bbd29d
zcccb3497e0cd905295cdd4b7965248a66c71f6c3080fbacf3c80e0b5507c96265bbb53ac49b7ce
zfd66c6d381a69a5502cdb02050fbc241ed4afa790685968554d23e0f132d5da10c0c88daa302ed
z08cbe12e29c21554f93de0afcb736e964265dcc3d348e0e7060d3f18050311f27a99510c03f51c
z0a89f25f2fdc4dcd2888f45d18f10d5a3e89b3d88b5c90326219ec0939f0b6c9105917392f3645
z93f9201b3d80af4e18a8200264219f1a7a62f379dbcee3ecb09a15d65c62354fd9e8fe5796f781
za1b8042f50e8290d02aa7c184cd6026bb3048184b2c0d2a87868e656874b1cece877eb16bfe390
z5d1dae5879fb6d8051165005ea53f96f068791a60e936733860a71f2bff3c84604dc2ab41a7675
zd8d942de06ce20ed9e0f2cbacf4629d43e29332d9abf8451dd577b9c4c769a939a1c50f1fe2386
z83bda4ae1de682dc88b5c6573fd025a341fa043300c2102f6e1c2c3a060af472977f3722b33b79
z84ca814570b77758524e259121bc4739cd2b1776382dac5de4e089dc3cf6bc34889ac2f1f99c24
zac64e3b4db635edeb4ec53c7fd88825b91f0fdb58f2b786a87254ddaba71aa72e6a080b6eca8ea
z207c09e43227108181bb2a782291533c92d0781d7e7944e6ec92081cf63489e2d70f5e5772ba4b
z9b6139e0a281e263e51cd9d9c0b5168ce93336ce77237b53823637c4bfef797880f2b68aabcf04
zadd16d6c900b49f8f3e9a01af2fa4024bb8d85a8acf2d6a669b0812bd0ecda17899a278530ccd3
z6198e0932ca7120ef331b5a0101e0029cac122b3749890db77c276c154de19fd8644f463c968e0
z69ed9be8e566e93e2d5f484677278c1ee4330336608ae27eb9f7ea02575828ffdbef5b6a3ea409
zc49c35ac1cd80e8af0ca8c057f758082166b07382f45902795a6ab4eb61fafeee22557acdb7793
z02c98a61efc19f335f975f5e90d73f903e571f86460487c0e4d655e98e31973131837dfbe1a181
z2e5991076c870b0743a466f5aeb497053ff4c32232125498d192b18c7a97a0e63244cbfa4a6bf4
za7d8b27560e532d8e2ecc78bc9aae02c0704f396317bbd6893ef6b03cc66a5c42e655caff57b73
z38726d44725c1f9de09ecf3bddeccb443eabd307262f2e298475e40c41966db14ecbc2cdfddf94
z4bc98f42941ebe0a0b9a80a65c14e390a89175af4a069aa19f773a41922d4870319e469c430286
zdf70df79d98e7c83bcc642e479f94b86867a993803bd5a8a1314b6717ef397496b723bd5b4ae41
zaf0c827ef9bbc1dcb3163a9b2989651b6e86ccd7e7ae1bdb5718ef0dc525c6ef90206944e68c46
zd7f8ee4875ca13539b83f088ba9310a6baa14e4808194f9d553b94f24207ddf4c7fca83ee3917f
z71852b9fe48938388d9e361b64445213794f21291ed031be902bc6d71c3c508d399170c1f2f53c
z9f4007e33f193730677ea3061d5a0944d34df2b144e45916c80f017439746433fdb88d7c451e03
ze416682cde8790b63db82da2172b13747c5713afe8eff066403f399cae65b7dbbd2099fa15f28c
zfeefcaf6b71f1ced94947c56113378caa90b76a7010fc95cb219b180a8efa7f1c80965cd984d8c
zf72dc5dfbdfb91a4660728cd7bf030647378befecb2e9f98447baf4a61149361e12364406fddf8
zd7da4e0abfec86861e435b2eac16d3ed4d1692fac6fc98e4f4e34935bcc5f53aed7b92b6b01b2f
z871c849a3923918f0733a1b83908ced6fea94a4da1c3cff251e31c4fbd1dc97a15e32328569799
z7ecfd7d3a334ac3164c6ba0b9911fbb4d4c8995ca66bfe99f08cb3871451928da0824877b1baf9
ze03f3eeb3d3223e7c17078de30d6faef918f72293e46e717fa7fb32e2c903e711fe8cbadafa04e
z917193889b873df43d95b0a755c68395ac595609159839f2d095d4ded5f7abdb4f17088070d292
zb8379a46ef08779c628453e14e9b53cba6117454a912959c1f0d0788d21fe589b832c4885c9a54
z2a1cdcf39c844a7ec5e4c4b09d8e44099c8801e0265971fe5436fb76c929d7af82e5f0498a7a6e
z368d2bfcb38e04eafd1082bc4aebb29582f8dd9e828858852cd168c0fc283a49f71c78ed4d8b1f
z9b22176209b3a542ea2aca6c6da2b4983c5653cd0054c2e59a46b1aac6bdd383a6c6197fffe2c9
z95cb8afaa13af4ed9a28c7df7ef8153c85bfbd0ca6d91421a563f834db5950002d87aa1163c18a
zc8460fd0737b666475b8dbea8147600922524cf0e7b576f0e4b55d04cafce2372e453604f1e36c
zeb287b9956480421234944c9a246c9fa9b237afee29e12a8f6b3b241689dfd2c1fa6e8c121d9c6
z08dbbe2f3fa5ca527d0aaacd2fa9f48351d54bba6ff7b4e5b73428a28dcbb4eecf6f29fbe6e3c6
z3d7bdb3e50bd8d509b6710532ad06b501af2ea01116454ab293763561bc93ba6dbb9c41b7bb351
z3437a800a146ee539749d15fe34862b90f11e31f61e29d0e0c24706cd1d2284dca4abe889a81ba
z5e138efe59dda01dcb56d06f86464ce42bce9d095579a0cbdd03d93c916a23bd2a6d7d0bc3ca72
z78a780d7d098d6abc2d81a2ccddf39e959f651fddba84e1bf8849b963e0a261e36478c81665910
z84650be2fa3916c09ff1b156862a698abd9edd9f4696553735ebdf0b3eee049579a018394b7d89
za0e95635671665f2b007e4e218fc1cb0d3d57d1d4da1b830cc394bb20c021a435106804eaee283
zcba232fec5d37d041a95addb12b26cb98f021bcd687c5143cf62fc9f87c6358a7298f9d3fabb15
z2f59e89e9b8daf452c5f29371eabaab9d17b0128027efe879a8357f8ef94c2f2c68698deedf565
zaa46417b8427d6c4cfcfebd3a6d81302d2ae765c06ddefc3f192eada976a7b3b6c79369cc579c5
zd127cf21c13c98808f5008b83b437ff9c10c55e1746211029d1a437a7e698125659daa14983e97
z9445cef2882abe33be4983af52744e215bfbcb2dc70ac9a3e5a9263194fd23052f8cdb61da1bd1
z82cd54f00b7e45203512e7b2e461ae2ad177d225f63faf8f0257a48b61a4a39eec9db6ee0108d2
z3617e1f5be69a1f51d6590368f02b690f1afdb77243f414799b79953a5c4373c526a2b3bde957c
z03a21300ceab995f729b45020e716fbec8a3e5ad613636b491db4d93f7114985c6f1548dee3727
zfa1ec0a6b679abc2a2c8232d3dae435936f00cee72863ccfa1402e611a55c2605511e1e0b7fc08
z2a34896176ff56a99ef2d0e99ddfd4e7f01dccb293c8b09cb0710285b0b4334d2fdfe616b43510
z6740ad1f57374876e0cf66506bb4776d9653a3f862c448eb42ad13d2c953e2fb40cc11750d1301
z7209830b9cadd99dbfb6a4a08125b386892075f4b2998b1f35e6b0888105b7fd9b8e9f8120266a
z19362d7e31083f253d9c5d908a5c8f58ae45e6f78d4d700618c28d43ed5af329a4e2c603615c24
zd04ce7af071e609357975401b621e93a833af00660969cdcf584d6a9d01681ea726f555767f0da
z6cda0a56188caf569265e0a8b6db96bc56ea1e52b2c794b2532e8e4f222ea0cbbb67e1613b6ee9
z411c51c90803bd2857e75282918770922ffa576de4de19c6eb722312eef0c08ea2dedc680b7e49
z1bd2ec2ef65755169d42d21658c57ace35b49e38fe781421fb0334e8e6b2692569d4b0b0b4a34f
z16babeb3da261f9698c35d4224cd56c9a6fa601e0ac7ca7167547f9645d97ea735fa6320151ac1
zc0b08092daf2b580cfa420c2032e1e0a4486f97a2879c5ad0aaf1d99812a2ee6553b3b9530d4cf
z05c29f044eadcb53bb221189a9904f4a7e07292bd4286f7d74e466c0caf13d83c10c307483e7ce
zb48781b280606a695f6eaf711bcf94aa2f19bf1c8c875f9b4658e737218f2877c7fb85316b3a59
zb2e22e181ebb1788f675fdd2611f92a75adad826b8160e2bd46e88c2932a3b1a69767c3815e9b9
ze955d6100bf690739803ad65584437af69e5490e3b7e5c86e091b3c75163f91d4209f52bdcb43a
z61316b7f6ae2e0674e71405e042fd20c3b1a7e6016a330b2016cf02ad1ca746fa21504dc98a2ec
z6f4bd60325ad2f9ca857ff43845f26b3609a7ab371ea3dacd863583e90dca3643c71712c3872b2
z7e722365e13e7f4cfbad79f3a8041c7be91730dd056406991501fb9818c44b5794f9aad93f849f
z15e4359cbacabbf4b03e4c54fd04dec31e78180e78b2e8d6b19ec8a3bedcff172bf4f8684764aa
zb43ab0d1bacc89217eea5413eda2dcb96f52425f18b0d753595bd6db1f4db48e150a8d43804ead
z41fe6ab1c975b1e5230ef21b69f082f68f197b1a9389baea922e724109b172a7d7f5448bb9e378
zf4f2d085de155de6bece3d730ff0e4d89f413aa9af14585cc0dcfc784d7a5df63b0104f98124f1
z7c4786b9b1beb87f186b58f1cc862abfc2691a72655a2f0389796a8979ae7fb85815794d04c1ed
z83a6438d70480112352ae32f68744dd6537093529bc5debc6280ec1b30e9805d7ed0d85831c118
z3f8977354598347802c0602cc37bda089d15346d9ed35a7b6dd7eba943f39fe4a822d8414db5b6
z8e0717e069a935f90cdc599571675cc96d5cf214eb59b66d8f0c606f8c02a83f279e6cc154b4b3
z27779621006ce92e1c8711f99cc8e897186f5d50940368cdf6c1df6367e125673b804b2b2b856e
zefcda6b4799aa8cadba68f35510bb532129c483571ab9c2ca87d80fa66bc9c449770f3e9f15196
z52e2dc76fc74e4fe587f8fbce8244bbed7acc5f36dab05bc230c70b809213470872bbeffe4b737
zdcf0a4b4cd24d8b9b166bacd5d2cd6e63a96908153038ffed955c569936e38a6020cfa343325f4
z72d4528e60eddc597f869d7ca1e0437f2e1adcb2623196ab099e105b44a1933576e41988873907
zbb6579c94276cd6fd384be9fbef51118e6f5fee5321e7e601b5f2eb6f17b2496e9364d92204cb7
zee79b9e3436b892fd63661962348abee478faa9a24721ce3389dddb4b1e04a4a4c61333c194ec4
z78b454513fb34f60945d5be512ffa2b1d3e73dc20c49265eed9a3bc5068360315944ca06b32932
zaa85f492841af7af08d0c27a6122d51112c6f4538b4df5add49460b96bd6d84866a9b1e417bc38
z68ffa22c6f9e196a84fcfee76c6cbc36093d6be3b4011be7fcad1e05bf534ff53a34eebab99383
ze6b2fa7d8a16807960887fcb867d36ab1e12fedf7d25599425bd45a7343ab9f88a3315dad96234
z6da9869c1e7398ac875d037ac6f49492a78749cb82fc2cfbb828365191145af417580acf606a6d
zf900ba47399ab753d851e0d696f74cbc2776d66e82f703c2b7204e70c10ed07b303765bd1be0ee
ze1bc1f73ae0045e3f91de6f76d952f126c0fb63cebea0cffc7bb76c1f9f28703e16ba2815f1dfa
z6d3ad4740940a7a89ba38a93272e24bffecaa6f16572d0ca68a970ceb8ac3a99bcc5cac2d6f8fe
zee42bd0927c151f24fd5723d2094692d97328ce7df8cfd8d62a52c39a379d49e4d05ac57bf724c
z60e710eae3b1b19902e211f8b8f24112e2c54e7de79532322ed0553d0e73987298e89df9d7fbdc
zb83eb9c2ad07f876ebc7319152dde9d0b7990eec3adb1f30e2f467796d9dd0cd627658869af6f5
z0fd1192d19b0ab8a824030bdbd21122f7c8d087f869d34bdf366d14fbf63a2adf04854e141fa58
z02ffc896640ae53d235976d43786e14f4cb1693feb4147a3dc7ed048048c5b2b42be0f3da7d8b9
ze9492abbf9ee156fc5f17ce97f01d8b3769381872232b21d51327ea3bcf8232cf4af308730d8b1
zae9e8f2ba2d66f1cc9068090d5298e9dc22c010e541aa0cbf6be53058e2afc0e06df2ea345b03b
z9078799e71c64fda6e4ecc70dac2085a62523dfe093c2a4a2fcef8da46376c25271e8ab46e327a
z505def7d202275a116d006525f303e0dfc21b8c1c769fdc8ba101970f9d619320d5d6c4e6e9afd
z172516b0424cb36d77b49b15603bb2629e4cc36ad04e9737f473ae72a4adcfa94895766d13e15e
zb832737d31eb30adaae67b3e030a66276db265b1e6e341325d9610c7258f6bf8fb4117b268cde1
z322daf065761459e76e863914b4ccf19dbbfe0af370e2c85e8f48f2c061ca3cd30f2217b757754
zdc44470750279b5c399e94e68f55a1aee58133720df87e0b2ea4cb8aab49a02a2f36738f75c135
z54142ac9ae75e92d8f06dadffaab83a1a630c77d112616d24ff17a2788950daeca32df75b9790d
z06387b04fd492dbebfab129dd29488ed317e1c6c2325bc8dd429c5ce01c88c648b067ab5c95fa9
zacb68cda1c401aa36a7b847a86405c3abf3061b07079b03963bb4c7cb0d258ec44570b6685d4c8
zbbf2f7c3cfa9991fe54f067f2d6548bbfc3523c45198e43804020e09cbbc76d5ee2cfdb4f374e8
z1f25c2eb892af5acc188706569f5dcd25bdfd500136da53889fff3ed816b06d6b1dc0e9b3ce8d4
z007cd7beb829a9852e8876136ca95af014fa6c2edcd860f77639c2d09e53c0284ae2542c10ef06
z984384f85690be5118c1731668197c51155d346102390f2c694fc3d85326ec5a13cfaa0f7742a7
z3c39af561408e16f89f3d5add4259e872ab3ec8ce78cf0078f7e668e7f796cb3fc4c8a36c1c5ee
z44b1a18dfec2dd74903f8eba0fff80e7f41fb7c72c2c0b0acc62949a61d6728e6cfeda58f5fab3
z289d35d085b0d0fcd1a3d77638e3eb600dbca76885469d40e9fe2bc723e4b5ae8a98ae64e250e8
ze6321e08bb2a46c9f68b4cd2e019672d20b3b9e0e44598b6bb6b5170000a8cc50d04b7efcd6380
z47a36bf13c703042bede995c1a766b77ac57a85d544b156a294b1c3b96a908568a42846883ce90
z75e98a132145eab1217e5790dcd7ee8f3c859711590101958575b677ba123057b2c1004dbf84a7
zdb062928ee42030fc18b5f2ee7e2bf4fc9571a6b546d12ee2f7835d06a50384e983ce6a857f078
zd08138227665fa8f0e02cf11b203e17e945a1365292ee2a67b20f29f0f590a81cd2813dd76a498
z1e0cfa50726520fec1445a12495098b1b6760c7fbf5fbbceb5f8449d5be4fd20a3c57b9f64dab0
z81dfe128e3fe018f543b6a8946ad2a7ff43a1a2b86d19d97d75cfb15b908247c6d531fbce4eda3
zfc4cad2a6dc648384db056992410fbfcc0868a0067713426527e07ed2c467eee66693c44547822
zf99fce3583d2f3606ca7ee890bd0aa31803ba4193d08d109b86877815ef5ae1bf4b6a777f8898b
zffbcfbbaca16c6e5e1cca35dd93836670e3b1a013ee95ede2569a8bf9ce3bd710615d096d24592
z56f9126cd16ba6efdfea477ac9da98228813c05319f0bdecc34adc12503d5b10f94f0f65fe214b
zcd8a66d312a76293a0448f3aee456bc035e05f3c13409459a0a8e8af4930d2170b272948b5fca2
z85a199eacf0db1f7daf6529d2178f00f5273306c8a055868dc253b0cafd558ae304442b4563449
z18c75eaaf52d17e40578db4547579b58ce5058624e9d9b7fa342fb17b4d1b6802f60bc1beadfb9
z17dfca3178de4e16832ca890fd83450eabaae06c62bdacfb150039c9836bd01bc61a925a7d19cd
z29c3a0d87cc763734f6b942078dbad9256368fa3c356f0950f98ad8551553ad757857c89c81b1e
zae7bac51572ccabcf3bc8ca9fb610f98b5a3f688b4af1951b4b120d27d8d7796b7aa72a5c7bb45
zbbe4a97eaad150d62a4d278fd687db670c4ca09d12233e25e8811d082295658e42889b961634d0
zedb0e3e1cb532f3069d3cfc85bf8d649a6fae4797f338580a73c659665b4071fff3c24f91b5b20
zb2a6c86c161f26a498ce46201f46dd1cdd95a1b513491e0059989a924de7dac1da28676acaeb40
zed9aacfb8e7c3dc102e6297d7ba5f6b3bbd9b9d9379f83a5ad8bfdcfd78d35c7d55a68914552f3
zafbffaf5078c9c11193f64be19753dac25398c1c67298a771196978cf47a05270e34821fedab4e
z20558a3e05719634289e0b2554403ffabe34426700a9ecb145f12a1e0f68280863f708afdb20a3
z2571934e6a39f4633879f7b3cdc3c51ce4b8a1192c3f0aacb76ec2ce61a6841b0d44f401fec294
z78ac6895c6c7ae5c9b84b5f743f7c8968e5ae0bb39cf811c3cb524f8e3cfc58307bb1b43f15f71
z8861bbbc01656c987b99bdee7f041c9931eff3b6866b8f45df0e8c20c8af4302c05c8350677c65
z65abaf166eff482430f4d20688ec1256027840924268773b7282c2937f71b2db7162c313b435f3
zfe1d627a0f61c88c645b1b15fb4186464ad2fce0a2056b6932e2edcbdfe809f68814604c37f154
zf2ec0f0b261eeec4c2c4fc605bd1b1634a98b863b7b12ab33aa6c0206c98ba4be2feda45ffda8f
zaba450e19d1cda639fe711c0e25f2a6c58878ad0c5ee8548f65128f35e103ddad0bebab3af89a3
zda585558de7478e85f7ed4ab126886a3203447a69e3e84e025d1d42a3c471c11935d97940bb0de
z787a128bdea2a7bf1eed5fa9a7021fe3d461855d7e9264451fb0d68f87f19191a451d60013b26f
ze9dfcd6725dd49a058a00bd1da7b2b3977bdf64d07ca7e8cfaf603c87b7439b821f4691404eaf0
z77ae187b5950e0b9739e6099b0f99fa7dc98887dc507a7eed507ebb851a7ea2f9048b5f450e8ec
z1cc49f918d4697fe661e5b89e5501866eeddad2fe3c14ddf5699918f1c47ceca7e019ff8a1ac03
z26d9c01fe92538de769fc0bd84239a6e43324c50fe16ddc30ecaa20fc53d925f220e56d6869a90
z3c4077bb05c3184ca8cc0ab4e002550164cfc690f2c080ed33039c7b2ace4985372d4fcafd30ef
z62d0bb516ca60002a74610ca366ec3cc4453a2f6fdf95e76be0952e27034659c2b7926e5b7e97d
z2f56cc18f5643d2190dbe926537fcc6afed23bc0f022ad52ef59e876ad7f859b3f3bea18f7e804
ze707a3d80bb12b6e9a9bb7f010af1e962840df58a70c02b829f1953cd095686054e15b56c57036
za10210ce0f77a8b779ead2591226e47f9c366de1a914fa78fca2cc1e90e20543c1d75c22636506
z0fde2e58450d42c65f1ab7ff87016d9d89f8557e0c135d28b162ec72ae4e6bc066014be969f5d3
z8c7dac9edd5c9f614928692fd80e2b1e97599233fae2df4ed6440204ef085be2e9d598d0e40623
z8dc0d0bd1e25afbcab38d137567bbd4cb0fa91bd97a1ba50f42cf4c2b8d34aed1a44c82ec93975
zadee24f7054c15ce7ba84dac9458ec127ba1522c5da36192dcc6c5d8fe118a518d85f70a8674e0
zf1618c3301dd367c98eee312c9c98f54ad5b34ce1d54a875841d16e2731d43c8dcf98cc9c970c1
z22ad50b1f49b42c91393351ae5e9fea809f148be4944d746700e1845fe1722461bc0630d7f8b34
zf6c0cbdfcac95fe965e1fb5ed6850fda5120258b9a13a9d33921c1e714682711632ac067d8ec5e
z309f34382b4cdf296889a2179e67db8d0ad8fecb2b67b3bdbc83d527b916979d1e5074fa7cc200
z665088586f1da59dda5d91c2310f253c8622d668441c307e74f266add31ab29c2a6acc85794780
z2f6410abc128883f7ee3b55534421a96bee08dc49cba806ce29871d32b211820569d0d1f91bbe1
z53e2cb4c4276843f034b7524d8806b99dfbeb957ecc8cf2ef01b6ff7d8a86c854d45752ff3b835
zfb21fc04833d87939faecff79c7c3f0f81585089a918d3c64cbdc42525b89477ee5f288b5b4581
zd0871495d3fc1a9e50e1b624c984355d56a9fc456a78e63f932969fca75b91e0b650a376100442
z34762c3b94e405339dc4176f30fc235745376b5292dd181d97f5ce7c2ae8431ea5383c42637905
zacd1414bc44d8f2ef375a85fb95a94f0d880330f358fec23e3fe5a6e0515be5d266218c3270089
z53af84b6f43db4b540f5f8c78d04c3ce8aaf876f36d323526f8ec71878c923fd37ed75dd7e8eb3
zee930c113950be380c47d722b49241292b24ca79b3b4cf71d163d0986ad7cd856f998d6a1b6b8a
z789e9e708d4ad5948cffa9c27e3b46cb8df8cb95095cbd2fdf39d3ab689a60388a8f1ff351f93c
z73bcf0dae1544a245e936d01b310a4a38178baaed507dfb9d7822f1fdf0a5cbc16fe0370f7866b
zecd11750760553c85f22e59c844865ef6757007e05c6fe5c446f539113b5704619b1bd9cf97f43
z94b03009a3300ed4ea0392d0afe22783421cbedc57cf84aa8793efb645a56f37b463b12efd8079
zc6fa547db34c0070c8c15b8995016bdeb15485e4ac5f1beb424e6bcff628fe2b33240f9b63549f
zedaf6e95ae5e306418ed4952e2630a01f2815fc904e03e766ae4d8ec41cf4813fce9cdb6afd5c6
z85291677dc0e687e7bfe4d1912f57ac9a7519fa75612256bb09e78a23051a57d9f0921f055871e
z0ea205992d67c58e8fcfd7ea5fa4ce3f5bbb64dd0eaf8b84167ef57e8ea7c108523912e46139c4
zf4fb515f4f14e6687a12cbf461199606ab18735388964d14a513095bbd3848dd186d5aae440417
zd62c2a8e7b24bbd06aeba8f0dba09bfe0cd3083c5cf436387a944144e09f7feb85115890f8ac8d
zc92b450a4959add72a3d92e308dfed7399d9f4c64af723b355c9b56b711a52aa6ad62fa65a5c19
z1ae663d9c25a0b1269db85bd03a215d6bdfc05c9e240610df29e2ec7e0491bb2bfa78a786834eb
z492407c698c6c6e62fd5bf08c9a90155a2d0223a4b704bb4270d4d10e9ac1221fefbd6aa9e2b14
z79df5b68165e66cdcad2c9b010a0d16e354f409ece240e07ca77a799002343438a1f4e5fd4ac15
zae99a704fcec71bfdcbfa4f29843f39b48fe02562e1861381cfef95c36c9dcda02396317d00daa
z8f7034a5f03daed8bc28c6cf9ab05ec09a4dcfd2a555ee437acca683e90c5df062f8f2fa6332bf
zb052ed0210c3991175cc536706f9c48c175cb6bf3bfb38ca1dc5ab550db45caf8bbaace4e0d429
z983f116324cdd990cf643e58f8ea368861392f9b76060954e235c3af141d0e5a5c871962dda175
z204d8d4ef1c08d1d9784fda6c51b96a7a90f629bcbdbf916eaa82156178e2ee5cefa02c5be3bbd
zdec0713dd041bdb51cc55918a7660325d105bcb0de54372bd4fe97d09d39f480310ad4a6844f6c
z2dd32366fc91a1c05292cbd61ce8bb1ac0560a8e7f3f8657ee5fcf184fea4942fc2d39489de7a3
z9881829ce773b903229e32b65f27a1f8ba1e34399bdafa3a3274c573d12cd58fa54cdb49627798
z7786f15edfce6ea2f0bfbf9916157715b16515b81611301386eb91e7280abfe09686bbc578a5ee
zd1a51d3122eb24a383ade3e9fc9589c890f1e0dc4a380da283526e12d6707fe6d195a3c2705d75
zef7f67485b13ce1d61b3bf246f8eb245e48b8310e08c472b10a8bca4974f2cc23490d579754c3e
zc320b6635baeb1e2ba422aaa2f1fe3cf28e8858b9cb242a512b4ca4e92abc8a69d0ffcafd290a4
z0e75595e757e5c153dffb03ff87df92812fc11ae061417491c886d2764436d4de9d37bf59a9bdb
ze054c1c291ad83efddeb0a67893cba4476c2cc4933c820e6eec454c5b918e9ab8c2c87f8ada979
z62d1c99817a8b1c0cea66fd8bf93152e9014810446f255d5fae5171ee124da36e01a345e0bdbc8
zf9a2810690681d61a194e400e8c59e76b7a7d6fcd11b5f572e4f593029ae3893b5ac58f2dc79af
z37b725dcfe736fa9f3121b67a636853a68b56c9c6bb22c94786b98ccbae9991b1f7bc11698d0ef
z9165dd48f52b1838a3442c68fd47479ea9485cd80011908b23254044588323dbdd566e8937ef10
z7d0c66feba4ed03c7479b4deab21dac5210af53b05daaa8e1562764b006b1ced2315e4d36b49e3
z870a401a9506e524fe43f64c9da1e55598e0e0cb852bf159fc98c73a78f6948602855c4270c4fc
z3453267a09c62bfd135f14561293ffcdae57e711e02c701f9bf7602cf58e19c7b3660d7c9680b4
z1eb26d2a55e9f856f2f6b0ec181a4b5000eaad762a1a79838e546dc240fcc27cec91226e403fa0
zff3a955e7a054984e163d97c6398b735aebb2e912f4f7b651a46f6a5cb190c540bf16addd8fa23
z9aeb689e8704a90f1eb9060099d238b2425ce454ccbb5db86755a79d7d6693c73604614f931f6e
z9fd0a70730a2351bf909bddef9364a95a31662fd0ad69281408245a7c3a01e0dc57739bb806fca
z36e3dc754db2aafd24de01c67033460a6b89cf1118a08aa8bcc7f7a49594fb7226c3fa8abbc2c4
ze6f7b17779ff53b1e796777d7e6bcc2c47983b17bbe8ebca53c3a1873a61721f362a7e23eccc11
zb1bcb74e27951580e51fca6cc984819a75733e39d91f4f9e1e4dd90c94d87231f3a3181c7a2c52
ze18acd491d789811b65dc96528de62c816556aa46e7a4d1483a88fb1f44fb5b21d5290a83d03b9
za5856890baccb0a9f9bc6ad72cbc579b15bd092f9ceb4abd39040153f0fa65d7c7fcd18db2829c
z8f6f6e2019925361163bf74bd1dd264fdeacc61bc30dc0ae67fe9e3f305904bb820d569e7f5ade
z3c698fd9c9465af10a034893240a0199ceb6a98adda8bfb2f174ce35e5d6d049c07815d7de34f7
zadf5b378299d30e658593310224f06700860075a7cfe6b500f5cdaffaf3cbe923fcc8ff0d99128
z1087b25c782f31a06a7a6efb332d8fe03f40929d124d64ad238e08daf7e2691670b172aeee8f64
z244aaf0d706885f9769db6fa9c11b1d8dd6d9b869b064e16edacd57d0455fe80902da4a1c9ad64
z1fd9acaed8d087363af9e8c09faae61143b7e4ed91fb8194e31654c873b60e93baa510d2b888c0
zff72864b800e681a93c8e53fdf1287672e16a498b0d91dc0db80f962d4c82c948fadf0dbb7c504
za4e1a566d724907c70f14fc530acb4c4e729f73fc04e562fdf005094ef50cbf41f3ea5681b51cd
zc7c59ccca0ad7fc66059db41fbe9ce43e53ec4c79d4544ad48236759f239bdea016d6783e638c0
zaac50c00b83ef6923ce5a98dedddb2bd480d40d930ad0a2accae8e820d7be8a746833bf38617fa
z5b404e100c2206cc62d365973844808bbe87c6f64dc271db6ca4c80f2d8e3ce4cb8328b8100ac6
z5fd310ae29e3003878a6ae072402926d9a551f6f226c1a663e54a4bfe582a1f44e9f928d9e96d1
zaca6ff3cd8960dd91166567ec7c8e7b176bdc711844a93c914d66385491c7dc255f98719b95877
z8e8fe88944837efe1c12b1b1294bd8cdb3dc512b4b295327742d796b7efc4caff560f6a12b6e38
z1361e01b0fccc3700e6bd0c3c026b90ea6a7b6897426dca446ad10d79ef1fe650e7a04fac1337e
z3908ce695372c1161d0e353ae4a0b6db7083582370d44f047c7835eb20a18882e46f61f88f6239
z16fdc93b8a55adcac1b7e6c1d7d04897da7734df271f72433b4b971c6c58209fa13a6f11f1d6a4
z8e3d074b381936b8813c7b3c94cb59f56bc388af4420af738d752f9e499c577bdd8e721a18def7
z52e539f42a64f46dd5e0a25b5ea6b54e8db0c8ba910f87d44db779f8197c1ad8bfb134b06c42e1
z707a0b0a481a3ab50ab6ecf2b14d5ef9c4c1e81343765e2d9765b5a61c9e250f1d233c55400e87
z039e1e25d7b8ef78c34c211b13453dba763472895710071a985327352962840a384bae0b1fa015
z7ac9f327fcad028a91ed1b8478044e856d9031c6275617fa82fe97ffaf5ff05b7643e74a03c440
z0460c649e8d95ae16f4cabe05a6e30009e6798fe11a6967d2e10698354882807adc9753bd19fae
z5106b71bd7f38e223b604bdb8610871d84f8ecf2c9baec95f5df2032a7bd1e97f1c1b068cd3254
zffc6271a67340251f1d5225d2395916fa2cb09e907b1a1b010cc9d6a0154ed446f148c772a0f19
z9d72908098fa0191e932814909970ee1389a4062f4d9159a7db9e1cbcae84d9aab95b66d5497f7
z92078152573de951b23a622d2321ea35a7887af4a6ba6cf346522515dec87b34721ad3b3c05052
za8b94708bfccb3f9a1224cdaab1d4246362853c004c6ba4a3c6e2a1c5c148dd2e7ab9691e6d6ea
zbcdd365d29cd4ca52cca02221cfa87b211c2ad83ad12cb09edde2d93995532c52e5197bd677e2e
z2d31c63371eef0176d4fc50a301fccf534cc3b47b0a0c6e67c0a385481667165a9f51246be713d
zcbc0abc4dd2aa8156ffad7efaaa5024abc32b9e0074f1507bcac8e603e4462be4ed852c78aa186
z64746ad4946a8dcfb4dc0d53db6009103498da5ae16a9bfaf826a99164b5147328ccefeb38d7a8
z3477436b0696fda0e1af5d2b95ac914021e7a9f59680671451a2eac5e94a07a3fb2ad62c49b243
z3c9033554d71a122fdfdd6940acd475ab0d7729fc4533bd3bc32ca65b2e7663e58fe2588f69717
z162f436f99bb5444a1ae4764291ac9dedbd1e5b2f49bb34d8017561328ec2163f29c412c844da3
z8dbb9aa1e9f28512d581f3ec2d57754b915cd810e06031596d6714d3a4e2be69dba38b6f58af68
zc2efc851d282d144480284606f126f19d85e8c4211be33b2dbe9c2d9e1140b784357534aabdb04
z23be9e5e5ee5767978c989f965754d36e3a63dab3480a583c783d5eef0d979f918a251aa82bca9
zb98a2f52163defe0bd8065282bf4560c957e8edf78e596187d10c39e10271595fef2d2c613ba96
zfbe658a5ff3c110230c2730b8f210ded179cfc71367f624b2f0c683e9ecc9073d65e81fbd15e55
ze8aaf70a6ebc20a67e570557b794254791a57cefe3b44cb59ce50d2a01831aabec6d653cea81e8
z0ccee149164e27aaa2f4ee303cd8c87fd1a04fb487177d39f1937dd9464f5e15d5f25c5cc057b2
z3578ad9401d8f89e8fa0e667ef7149205b02968ae31e5a4af04e445662fcc686f3b97af220c38b
zce0651f626e9e61ef43c26e4907818b75fc93a8f82badb42e18351e87339595fea8df1b224b9eb
z9a144b4ed67079ec01e499369cebf95573c832549113904216490e47c07786e17cdbc7698fab79
za9cf3623a8eba4e8b2b2d274924a327c304c60cc58ccc01138018ef78d65dc22772399a193eef0
z6777ddac06fbae3134804329075ae1ca0211b1f51cb02923526f76ff8a475e0a0f8559dc5a1676
zcd4de81db84e377a947fd0979cd8cc92ae4ba8cd8660bbdc6c817f75aee2d6e6a0b834810f2350
z94bf7fbd0fe7743a6f3e052f41f4f698022946169ba7f5240c9d972233b34aca3f33dd020bdae2
z806149257003ea3e56bc524716f09f83449b2d72d62e72dd8b52912c4b78bc417617172ef7d971
z217fc6865203529a75bfd8b053190f2db667b5f886dcf660ccc50a9cb44e393fb61294c7127820
ze4b67082b6480303625224968166ccd6f01e4aa80601894d884cee59c06a99bbd0c6bc9e443cc3
z7cd48ebddd6a3928d6a4cfd48633925696dedb46f17a22fadd1b4427b5f94513ddd8f6f6cc8bd5
z0dd85259bb04e24e7d4e036249568379a5c5c7bd0136a87549b6be5879881f0fb4d14f77003827
z9e6cc66e0f9f365e1f2a284e6d28d1bd5d00e99ae61677097e0da2d0aa8588e901886ae97bbfd2
zff1159fdc141ed1dd352205c73ba5c4b37b9ff52ae8a95ca239beaa4b8ff89aa1ac89394a714d5
z6ddf61b252ca17b8545bd94b2794d4393deda5714b2172470f531cbd43015c1305c616a1f6c1fb
z8eb800bc0c498e6a27a442480cd3aa510b85699d3bde79305af2b72867477247a90154a0bc85c7
z107181c473e621896e29c0926b544fe51982869fbdd7fae95f78236eade62383b1422320d5faea
zd4af710967f66b0f3d1ab2a63382fdcf72f46b00473b0148ed7b88623e585961ecdcd5a1f4f242
z971c95008764d151ece01ca6dd9749dd30877ca53ef5b0ec37e73f26e8e08c1aae66363336ceb2
z9216de4f392da3f104145fd861bb69e9386fb8b9f5b47459bb168a102d57edf3b259725646e2fc
zae9a22c61ddec7643af0e5949d2561451451bf878ce2d23c9fba7763092f0c2d3ba80f33cc0138
z026a9aa2c975f6f2de5d64996d4cd8412f5d823850712322dbc3dc0b6593972f028df09feef31b
z0b7e3394368685e8328ff96071aba2b01ac917bf3be95c92b63595fbb5c44ec3dd86fb2cb5e4bf
z83b1013d7e848fb4adcf8bb8c0a2da80590f7efaf7c47b5a4e5f087413909a8ed0eeb9f0011672
z6337def92154f7593e5f6b3942331f95e2bef4146ba5a1cc5aadabc22ccb34d4716d2d3080658d
z1ef2b24511cd38f0d02beb27e7c23cd9ddc0f97248c08d1201090fceec4fbe29a1b3992047b54c
zcc898500ec8473fb68ed8f24a20329a9ee9eed6ca7cca4a19a164641673ad1fe90ef1595c9083c
z400323af6b365f26c13a341bd9af9442fdc670e6d1fafbd3cee7deafadfb30040c432ebab533b3
zd77be81002489d35658448a98ea323df9810d96c4f0debc43232889ea9eefb0b10800f4203cbac
z4dea77c4f19d465205a678e1ec398a7a9c0a55c649fe8ed975f810317c4f61bf69b8ce6a33ed3e
z5ff1b67fdb13b692555677f989c6a6d9e6839a3aea52e10e2591c4bf94f265b9a586fe8cc4def3
za1efa95db4f3570461782268b94bce8b60cdb245867abac5d1e4d3d72c0a7ce385389eb28f3db8
z868b9db7a92dace5b1ac20252627f5d761b882dd2e7121f0bcb19382040a718dfe6403c72babe7
z1ac6685cc6f45c7b12f7fcb1cbbb95001915d5d1c0a0ebb244a0c2834a357058b12cf8d645ed67
z294293980c2063c0e13d87df3098c215d439b786f7e915927d1b110ecb3390e6b16a2c8cd44d33
zc61725a3075c48699f3602112afb0143d88cf2d2a2d3f514d108fa5a847574659b96210e61229b
z88c0cbf5474ed6e9e53ca69e2ab60264abb96ebb054486977b20b799a7f062a30dba09e5dce1d1
z0dee00aa794d9b0a6270223a2abfd2d6a5fbdd665c51ffc4738a80bfd36968c8780a23b0415e3e
z9a3334c5737d321cb1f0594c60422e18e12860572df517942140896ec9f2a272675f18200dc822
z8fe4156e739b99be3ee172a9ef7cc0cc296dd309f8d776ab84245c6525255f7fa89d54bac7b81a
z9bf90ee69352f05b10236fe880eedfcd2cb235fee5583813ce514f979ddae8b78543718b22fc26
z1c66080ace9a62b4ef93ecc8c966e571c6e211bb1dac8dc4041931fe650ef3a2e15754b069965c
zd6e7834a81a94f88fa52c9f102be38a3b30653fe2b2d625f926c3e3aff6e9d0f54dbc45606822d
z9b31ca65d4b9cb52d1eb09a300a0c87bed37846ded1170699d1646ce06559097373dd9de2c4a05
z1b21b0b51e75b6c24d0dcc8453df6b309c71fba1675fa8a51e2c5779dcd9c135e3398706da07ef
zefde2205b7a9745dcab611a425bbb5409dc45ff514f168fc3877c8dd2d504475778bc63be6a9b2
zc7d093d36d7845a9f5303def9a3175ad830e979426151136ade8341b78b0358164ca94ce98321e
z0fd02081a1ff727cdd422bb3fb5e419104d3c7d6ddcce1f4f52f895cb88d5977b8f36eaf534dd9
z050d5d3cc5de3d280fafe937c6e711484a623935f9308bf47b2d32649eaa52794cee847dbc5714
z1d320e505f458b32289d221a2d6f3fb8b86a24c15ce9829ce32b5088dd27e2e4092e0a79da6bfc
z4efe6fb2d86fd5c4ac024e45a75e4131a338b733b790b3db0617c36e8cebd70f15c68e120125f8
z80ff786067891e0c178e5e1a1e65942e19bfcdd0c85f3ad77dc69796c550128b20f471d0d6a91e
z98f0aed980ccd4e7470d38daf8a261a727e6c9c3796355daac93a83c6c20b3b3540ffd0a76c25d
zaf626bcd7e11ef5251980f791fb2d773b8863da24637d7566ddfeb3eb322edf34b33e056d969ae
zc4b98e9a16c1651f24e3d77adc3a973bfd6553f717512c1ab4030cae924dd3dd9db178e60dfc6c
zf6be97b0cfc3e26c882e2589ba1438c5c4c1da658c57e64e2520dffd4a96e1bc5731adf91b84c5
z9f3e57a03642140dfce019f3fe157b50180827e07ced63beed3dbae309c947831c09d1044cf7f3
z41dc51a3459d86b222136a029275f679de1724a5dbfac3c2eadf2e745717048688630207afbce4
za7fb980a151db820467a0255ea8a9228c5fa391f01b4dbec8597a3d0d163da35940c1b070c8ee2
zd64672c0bb18ca41d6cf54342aace0233e7cee90321354886a29f5268f4dd80e4514a9c6b825da
z7248d71763de70d983fab8866d0d23f9a1b4522f54d226585dc340a2643db4328758a613359778
z5e13fd1c1670d3c119848d93c589ce42f754d817e813f4ce9fe2c1bac3c8cb577b580491970d0f
z2157a44548a6f94e5cb5640d9a95f3cc2d6830dd8d1d9067417e6051a8d3607376f9dc3a8c07de
za025bd9e149220237d51de25547a95d2506c7cf01a1b763fac2a4f14fe80f52971e0bc7707b7b7
z9e7c934afe61777e26105740803366375d300ef3099a874d62b583b77338a2fe7f4675131994b1
zc01f4b5e9b955b6e82cd8a9b8dafec11fcb1a4bad2f6079a785f450d78c6271107a250bdb1b143
z47fd9745575cea498922a82ef04f6cd10c472508b5ed741705155e6595219f088d87f47cf682f3
zcca6c93addaeae619d713f05af9afda0b32301220861915cf3dce490e46a331ef45f6fd8dce9b7
zcf78680cea8a5bb435130bbf5f533c6cbf1e29717ef9c55e51fd69a2758d5a4d52b14fa4476e0f
zb697d39f6bc4f042b0d88a4a13330f128ba281ef8226064deb9069a6b913929bde120c2fb87755
z5522094e0663aaad72b9c5b7365466b98e0f5f493ed5dc41b232912c8c8b758378afc8505ea968
z763db0d62023a1de5f6206dfcf882d8db4af21f1795a00c8fe5b220b264d53f62d6153204ddefa
z7a2bc9c3ca83a63800c0b15d31f2dff919d0b0ad757db06508f7ad97bdb2e97de397a766a19011
zd31ce7476d1df65ae1075967b0f2d2b3025b2698e19bedbaecf9d9ac44fbf734b12d8ca91fb9b0
z014acb39a316762dee4a2ff1057c5aa5517c6d05290cc7cc215e58f9203cabb408c5a59d2a0cb7
zf55d3866b4a039a6eb450a442eab8f9e50c50fcb20aacba7e1c0c4ebc54cc6f7626a091f7e9625
za76570e288d84c468adbce271827557e9efb56cbb7c2009bdd7164643a3fdea825028948818fe0
zae606d0950dbbaee7e833a68cf93bfa3a090faa9e20e36d718e8f7608b75260b597a979d41272d
zdebe197e672b629bc9beacb126e229e461952199f11b6289778d44eec9abcc050ea10f73ae113b
z2e102475a08653e4ff268501a62f988567b56bdb89dda609914cf524f61b69967a8840a053ba18
z083c2da5f2c4f83cfeb76e06f2a172ecc8696e261d3aaf8351389764cc052e4ca80a2882a5d0da
z0973ebac9bc1376f70ebec6e6f4e019a05a90d4e965f4bc45844634164bac6a5bb06f91f3e0911
z9817b86004f73ac5a5cc3280ad1aea8adae537aae140b799421b7728d211d3ad17f4d3bcab467f
z97941d94bbb6a9e84746d0b2866cf5dcc61cb3c53d44a23144ec3a7976b0b845c20684d4c8f2fa
z450af352a1bf7ca2e4311f4f55187506f33f0abf7c08c2c3514427d92a5dea0e1c5ea698f41897
ze8dfaa50c70de04a5db53726db899f2a952df70330ddd0bca59c0445f0ae8f2a234ec42ac95f0b
z5d6c046261fe838ed5bcca2a8700f4215d6d6cd65924b51c8b003e782de010882ea61e2ec1f24d
zfc25c3f9d80d90765a6ef1aad0b6279b774f0958f9a0589d84fa52570859f68703ce036cf6e2ab
z099cb6580751969941890c83dfb1be65538ae188da842a931d3fdd6561a27a0a6b064945ebe5c8
ze414ffdb11086f59ed15048a201a53fc7d5998748275e8cfedac6d8853d8a0ee6c0b0d386f177f
z725a54057cbf74e109d6ba0efe98c698180f914c75f102c3d2dab967dc92eed37644cc635aeacf
z9428d85a519c5946549c5b372853bd2a7513225e5a7904fa33ddb1d28da626023f625f1923ea6c
z0e7e24ba7fdefb1b8c1c7979361d3ca242417697901a6aacb43138e0b82a1fc0049492f49501b4
z8e5ddd76de5ffff6e444f9d5cae77d2a49f3110c91613377d3e9988aceecfac5b63101319e404e
z53e21b811ed3386f731be620804bb4c85fefccef494a8f6f66c0cf39cae0bceba33adfbab68d3c
z6eb65b5d753892d1a50f34fcd3b87707dbef57a775195f0ec191eded3ae834a532ac397b50ea70
z99daaf28b9688c744fc2991da117c09774eff3f94e8bdf9f8bb94e09c58455bf302f24366ae285
z8b08322dc045ebf9ae03595144188cbeb9df78c3cfd685c458f2394252392d6599f47ba1d9e280
z8653829c53faac713b832a3494ab60a7c66dad749781b0c38891e07be9c814f53c43b3ab1f1dbc
zaea65fcefc1d2fe3ca965893695b739f6745efd5c7f4b92704c323f08754165628c0ed42e688fc
z66b6dc642282e75a8966a1746045ae7243dda1f94efbd746ffa428b76abe27da6d6d2a386eeacb
z2d7ad49a6ba8d4e296540c152b38b3945d502977f3c87a0fa80f2f4ffbbf67ffde6bf8e021f3a5
za0706ef09c8ca1a9835b2c24f0e846df537010b68c705d7876d03cea7434ad976ccad1262ac8b0
ze1b8c7626b53dbb9a5c0ee7ad17228b75c5cb92ca1e31b6b72f63167d44565a23e8a75ed9627f1
z4b161fe5e7da8c43a45bc39997f48bd452fbf1b53889693c193436f4a9eae44501c998ce7c1cc7
zf055c9fb9e6173b7ec694345fc0b1a7424ce28a9021995e2072cec76ef789ea6a10857a7db5dfe
z365e7f2524e0c62df27cf03d16add82d9eedb153634ed8c03eb74947533e48283a29b18f006410
zf5f205712caeb228d7f57ea99ef4df44dcfedd177f0208a324691d4668aa48dc4bff8cd0ab95fa
z618da8269a6b621cba745058aeb92b33542833a5b8f4ae748351907a02f65de282872438c67c19
za6c915359e500cd6ce616aa370aadff1d4d8a60a8ed5bde7e946005e86eaa2b98b0cc8c6b58eba
z9b61f094333022233f5002e2c9f359932b626fd724cae8cad29fe2169001474df1d4e331817844
z9ecdf8059a450fcd3e60020fdb8af883fac83d2da1669520124c9ac73c23db3a27fbb61e1f7297
z851cb681c10270ef51a876288716c51d6c04b3fcd2f0d37ccaf6eacad72029fee5582a62480491
z9c228a4b5825ed28ad7b20f05a62693ef43b40d64f7355f84918a08a83503aae4005c1afd9b298
z3e4bfa0e51f5e141950ef7f18332f6442613238743c4fe5e344592d0cd276cb375d07c55e87f17
z6f07a7dcf4a75ab6266ee0c8144ecfed45413dfb9371b77e5bb6965ff7920ce18dbd3216113c3b
z86a91530df361cd4f125983b494f08aec3e9b2df0d134c25b9a19b31063b39434eef5949b89fb8
z9839149f6f33a10db8c2e8c2a450eaad0c2806724906b7b4f48929c621013b8e2d3a4583f28312
zec526e360c28c6039608dea3d6cb46fa931a1f19be39a780c8da6a9ce2eee357ab8df7d3690bd2
z9be0cecf8d071915994a32658b7780880246c2e6e55437f11abc8b366a46d4c79a55cc61fc41c0
z1496d429d885454604e00c1aaf0cd645e770809412c953eefa0a6ca4ec11ef3311123fdb7e86c8
z12299726c2ad05e8b5aa9c9a751cc88078980efb03590e7a3cae0af803a8377fa4931c9dd60364
ze824188d2c917d0a1d7db0decee04e785962b8f1d10159b50b4092ab3df606d1f5fa579d37be56
zd2fa7c77cec71f374c957cc2d787752c61b864bcd537aa395ee99ee200a10912df89ee7aafe2de
z0ef565412032bfc7201a202e440e91d5de8d3421ad14c40b4961689de0cfe0f9f28a0e0c0465bd
ze1f199ebe5b4f2beca26af55be3f87dc0ab41e065807b9115c91baf5f52d302fa614f68be491c5
z16ff5843b6795b1d6fd355bdc04f7b8bf57bdada4b36cf0fab37d795b2708287869a57cc245ec2
z1d07dffc7f20994f833979e2c419871a048a33ea477b99fd3e7bcb9b0259866c79f8c39843f931
z843adaf88c7d448c4858f363db861f86ed1e75af1027f9790e34cb64cf4e962e1ade5c549c230b
z3a5688d3d4b39cb182243db350528403362f1cd7d40b55e0fa798c6ab21c40aad0e379c5427505
z11ca8e212374aeaf441828117b9635ecb593ace62270c220e4baaf45741975c528826cc9619121
zdd1248cb62628f7323d75dd0cfc48b905d9076788bb9fd282d69d924e1c209ea9184d6dd82b5a5
ze2d247545ac1fd176e09c0ad818e475cbe93275a3520c1e6428dc543948e2940d46e6924b7f7f3
z50477e6fccaf87623338f018f29f53fbad58d2560b7b1871d21b81fe531c8ec2b5a374f692842d
z25c43cc557e91be0c255e6dcd49ef66a97bbb31f0afa9908492d5d5f8e375b5bedff2e2f3ceed1
z13ce767df3326925408c80e9456099cb18c06770c8cd624e20cd21101ace1aea8af0bf7f52c41c
z686a871354efeb27a4d48293b73bf94f483e8b4afc55a7f422381e88ec43d48d4b5c0b881efb4b
z780cd458351591b9d733884840b20d064cc10a56ca66ffb8c45f17ecdcca40d9c66a2a9b54a2fe
za70841bb6dced9a65ae01fd17406b4db2472bd29472ca62ec8bc08fd066936a71f7c0f1a7485c1
zd575e87f1c180b47e2cd8b1386a8752ef6a648395ab307b8694cbfe7e5123d2fa32c850e144a1a
z8dee89370e3620c56db87bb17c986e0a11f3a013a2fe69f3bcef2b90393fa50ef81e96d94999e5
z489e9c54fbf5a495132cf49e693d4bd42c09b54d5fd353d707ca24834a0b2640919aa8356ff0f0
z946f4d7bfc61270684b6e707e68bb6703de48783775e76c773c347ff32e2a4ed2d33b00377f057
z2cd5491a10c7f036ce23abe79677733de43741178f192c0ea477c9d26d020ca501fc950d35a832
zd328a56ef50e206976aa2bbe2791b015a13534aa336c2f32e3eb49a49aada9d144534664f87d2d
zdb43cf55d6314c7e4327127a950d95c16109fa854b8a9ad9ed76e7cdb7dccfd6b2d1d955ac7b10
z862915c7c0fd549748a3e483993ff43a934535f57294f62c6b51a0e17d4910b757f02ad62fba60
z1b67c38d64b03cf0b32fa73c581d8326a2ce2a2b9f0011e6c2afd1ef3274313cd278fd19987c20
za6f3b91409417ef88b28fda2608127dcb3c3278d1ee88a3b8c4d431529835b37c18d9437b1ad2d
zd79fd3e75c1b4e577cba3d57996946a00347b6c36fa67956535c5cd744c9af8c52b84e71eddbd2
z8cb1a569c848e0f5cfa472072a37f11699220b3e0bc822888d1a428416c8c08daa759f3a7cc648
z0f2bc62226fb21290aa1dfb6194977d35bed49ebc9d409014eacf63377db5042b683d1b1f35dc3
z059bc0e0d3fcb7378f8406f76cd58c8c817f6354230f4f9dfbf460f0a2234f75f46a367e3de8bf
z0e0aea15bd9f0f2d67e33846e47b1be9e4024d41fe8503953faa0c7f49672b95822a810e5f44e9
zc8f47e890d3bb8daab4c53f01dff3fc14841c73bf1129af64773c933043746a00b933e4c408f8f
z6b28e019f60fcc1b42e9f67c476514beaf9cf5bae613e41347da551365043f734950ce484bccca
z0e3445cc1dff4b6ed9c9c81e3101921f7d92b7685f8f66a19c7809192b8542d09d93aba653646d
za3d5b456cac6417247efb4431f1e9fe2a683905230a56f5bb180e4f520c8a89f9d1403fa60e0e2
z50a3761ac601dc1269fdfa04a7c0fd61addcccd80ee6f7b4c1eb7441e14fb774bcace12fff3311
z418c9017b5a0fc86cd65236f80aafdc539d00704720f076b8e15647298df97149807da441b479f
z0a5234ee84b71a7c904b9588bb0e2b2712edd69c7af9e54384e5b09956104b57b826366f1376af
ze3a6b1b6eb183fdad15fb46a3f589940c102f6ce068a1f27ad7c0ceae77eb47d6d99378ade1b11
z544d9b0a07cd602545005300db8df0a1a63543f517df9f43cfc7e09cc33b5768149f63bbc5bb9e
z479b96f2629926fd75e707c9a9f57f846ee1b271c8227f3eddc71aa48ae3c1cbf21e7021a6f219
z2de59dcf13b70086dfc0f24b181b718fcf5e5b2a8f16a010b15ac564965332903308801de1e8cf
zdf9451a8b6b428d9c581dc9e1d75f25b4f58f3f067074288f87f75625d609e7be7c323fbc0e051
z997872b56432de27e9422daf11a9830a099a8a4dabba03a7947398191e05398e2e6abcb479390f
z7b89af3a1684c2bfdd9dbc7a897c8f34c3e701f0a3655afbe74c544b9ba71c26f95f52ccbc855c
z6ad41f8da1494645943b6e5f768800bf0a3180be9a322c52a3d1e790d44f088142d3c1c7152acb
zeb0454d0da01263b24ba6513ae0ff88d1ed99a8c35fe304647fef3a6fec3341157a581f6a28e2c
z63e748c3c30d743a5bc6e62a506894be1449b89b5dca2f574685809fad27cfa8ac85e824ead38b
z9234b3e72ef2cc424c652d1c3ae7206deb9e37d541adab3497b0faebe7926cb1437bca5faefdb9
z528613f643cb0605bd3aa303e1dac1995606acbc86c396fda6f2fa59530feb0843a89458bdbca7
z60b1989964e35a37b10fee66c0e010868db67dccd20aee615571d1b300ebb900881215e90e417e
z94badd85353ca3615e348da757b516cfbb9522ff0b027ce2445d614d36d3ab2fab5974965f795a
z40b094585d0429bf07e57adb9ed21771df135e6d4585e8a1b3422529e3a1381703d971618e743e
z88f5cb690990c5bbbfd283581ba5aff4ab4115a4a13b588511a27276e93bdde36cdef7edd8eac0
zac4fa42020a2f092c2798364ddd8cebc7a1c81dd47279a42e95fa114b8636ad34d89c849a0fb2c
z97064c8fafdab2bb7f3534dee2168021fe8d5eccc3140337b54b18c7a575053a643b2b9868d7ce
z67506b7bef06491e135ec6344352bd7c4ecc597e05cfbb91c43eedc661dd277ca83d2b4d70458c
zb1cd81ab6572194501defcb3e8c98bb7f27f0d848c8f46167f541c46de176af2da0b8430e0fd2d
z7ddbabd68420932de9b78ea4a48e17c55d988f2dc37903ac08a07c8d2dab8726518965061b9e2a
z0630389574b98f1db3badff1fed86072de76350c12cd17ffa44f70338594e82b7830dfdc592004
z32a59acbe2eed9ebfaf089399c3034e0c2b3b6f4662b914606e6af065d8e54b7c91764f9e650d0
za4d844a1c626a5c5828bf2b1ed6f27180d0f8b39d2cdbe072d4aa5bbad4a3df67a2083fa70a08a
zd624396f5362e8e0c3c220b242104ef7147199797f86538b6a586f1b5c0ee593d424453b2bfc53
ze77da61b41d8035289fdd2d46347aa7d7fc0d1750d573df9b24eda1741e793166eb06744a5517e
z5b514f2b780576181b5213b72e1115859e59bd3ff76bab09e6c3156723345036fdffc96f2d7af7
z927437b17bb6cd262a3da57f4142dd8578c9a585bda2ffbbdc89509c902dd617f2bc0464dbf6d9
z13b54f50e92ba44a545bff3c6656a7e6370c6a4ad641979b073d690ea8b48fc751dc0c400bf214
zb72d415390913720f8d2cdd394df4ffaaa5c4f6e392ea15d420aeb1445bdd75451fb3b1c047139
zc43e5a7a0cd216fc85ba4ab8b5c01d550ff5df50198208d7984f988c3288ba0ac696419783c6f7
zbfc74d599d966868ca400dd9da27b7eca1053949004dac70ce4bea019059b123b56d997e1d3b70
z00b34d0120a0fef4b4f87e66e5636a06cd597171a7783b0259bdbfd21810f22de45957f3fde263
z3ece86a3beb76c5fbb7a6d0d49a2b7e5af4971aa1efc67fc2f1187846371a5c676529ecdad724e
z0f0c6c04a0166bf6f19ac800cb8f1c983a0c5c8ad325a673bdac19752a3d8cfc7cdd694329cb2a
z24d84ae926f096240b197f5fd5d4f2c1b4b2d29ff4b169e18d83cedc5a3f064221c59b8cadafa2
z3ec807246f48af8d70888341813bfefbce93fb25ab6cccfa2e3ab6a6ba20a3004d9c467c2929cf
zf9a6252315c312497f9a51bc3f40bcd86207ce3d3241e36f44a8a76d69f02be6a008c1b1afe979
z5718d8205b2e54cbc504f32e8125d195197b38db836062725c380235ad2a857750c26f23429477
z0721aa4ccc100896b14ec728b57f1f482d1983aff7d62f20c8245d9495e5b7aa097a4f41519acb
zf9a853543fa338532627d09e5f8771d7216fc44e18f8ea07fe7a242b49e3ceab3dbdc6148b9087
zc3f757c890ab831942745ade74d5ff7601de916f9f60686b1357af2039db71741cffabc1f87c07
z2cf047a95da21492f61e7d06277c054cfd1978999dedb52b4c0c5620c441927967c03c99b0dbb7
z713587a044fd443ee2d2eae6f42e2c0a3a5178ebff6549e935e5d3d6d0629bf088f12fd3f8e541
z5f6985b565d00b967a392130476e1aec958e38f32552d04d33996b6a129507009de42abfe08f28
z6c3cedd0874da960f2d2f51084e42519fe80e625c420c141c4177eb61107374c93e60225718d6c
z5072081483381b75ebe96f9612ba2cf91cc42fc6d6c3c548ca51f9be5ef1cb95aa45fcd1fa889a
z4e10417016179ab251512a342c0040dff8bd27fac9279eaa46c8a46a6796da5c5cb4c16688c8e7
z0e6f2fa684a30d0afabe39391ba14f534f09f46fc5df7e0641af7380d3e734548cf46be75a929b
z27ece48bd23176892f738e3a69255ca93dd66bde667654c5dd6f11fdb1ee003256a4120d28c376
z05d023e78660c96d040cf22d1c3b23ed4fa2d531b9756343b679ee3be5dd72b1bf170177278046
zd329fff42fd9df4ada1ef893764ddcc7c56793949d25c0c9665672a1122727138e43844240508f
zcd820326155daadb4038cd2803e0fd2c82f9641e8d3a5b31ff34e16325d098d0443615d7c3e381
zc0e9874bc3a2ea7f82b273cbd8454be866edac867cb403ef94857f32eb0281952cb7f06e24f8af
zfc1003ba602aca1fbfb7a2d3b77c33234bf25fbbc919552704597ee3dbb684391dcfa7a5271d89
zeb6830387d330b62d8f5794086791edda99339acb66ce6c98dbf6e9d6416bb4b6c967ef31c0c36
z8d405bdf845d5e2eb29375d4ff6aea83d657e5955767ae8b98c711d56160b36e671aa55e4eb925
z4803c03e3cbd7f4d506ae6288d4dcdd62be066228d92a1b824298f3de59f551f7420886f0a192a
z8376423e7387deb664c9e3c807f9718636e61739f4b817053a8b3222e382c45a564506fbe6514c
zfa67ec211a7a14005877a0daa3875733ff853b45d27f3b8857c711b18cf0822c8d46a9889b2d07
zb0f1078fcbe91ea9a67c768acbd6f918a5aea6794dd003bde4507edfe0b73def1595b6ff166e2a
z44faf23e8298c84bcdd24230b6121b5d2aa01edde00d72aa809ee6c8ef5dda818eaf27e50a90e2
zb9b74598f4dde27aa388198ec654dcd1e3b3187f2e2c8688766bfb4bc8e04b88474412850c12bc
z27f01d0a64f353af99710e65a3551b9f7f60e5a92b48d0f766d9a0c6a217fad7850c167c80af2c
z882111d60bc44b1e6decbe54c37bf9b9bf1ad1c75aae180da056bc2738f9c8a45c15617380c1bf
z90171a0bc21f0d07e2fddf941beb258833fdeb7907d6186c12a0af149149ce38750351fecd6b06
z0a930f9805d0f5c3d8a7d6ae9c4dce07cc559afa3a5607e10e09ed215c6d72e3944a5389bcde61
zaafdc1127cc2c8abc2ad2d106eba79e46edfc567e4fde36148e5db9676f5d49ebde80b838abcde
zbae0bf945c6f2509d2d2231cda0ddf218f5e1db0b2d746ad6a1c2105b513e1cca7eef3de1642da
z8d286ce32cf50c26b1ef449f996741e783f61f727491d28e1e5ecb360da06c065341d4c06dcd5a
zc9fe51a6af96d25da3a292cfdc172eefac1958e0c5e434858d95cc036439368bf526f2f5f41a8f
zca5c07fc14f78bca303b1ed3367a61de53d367aa1308dd3d4ad1c75797266497938c98be59d027
z0c4bdf54d86aeea686cbdceee0169aaf6525a8110b498103ccfea2eb17438a8503f192baa5797b
zaef3d7a17def86d452fa60953ae178f3dda2def515c31d328fda8d6bb5a5c2633a4944bbb0bc8b
z734b10eddb544e95312d2298839b5d38d77061c3c3d22b37c0a427e0d65a37590748d11d0deb05
z1b971db7402d5479bc46fef3dd74a41b68a46463832ba3ecb08232c2e3a62c5bcd27014f3be778
z02b552736cfba417c73c979fa0fc07db533425a64246696c631145f0c0267b9e209e0dd1d25ece
z86418ccf174b685f447530092f3d78bab22c1e51ae12e007402be60003eb4feec25578f923d0af
z7a05052e286e043cad2a3230a3aedb4edd5fe13e9bd9471d95020bb9a3249f467d853898bd2956
ze4dc27a62eb3647ae1f6ab83776c57ad40340319add752a61821aab064c29def78adb1169f2556
zd9e383d2c1450f4d6aa77da81fb3ebe8d669d719c25d9c7739c9cf3e8a88e8851080aec9fd578e
zca1fa2fa9bb90eadb51a8c60195ca9b9f4c4e92c53c9836af6aa2b66cc689408ce5ce45b560faf
zf855ded8cab0d5eb66c9c1a2dd587a630fe94416a3c3dbc0808f8e45c60aab3dc4a5b20a878d30
zb8b9c5d7d363c7e35e86824f096ec492bdbcfeb55335d0381d6c3aee46b4d797b31421bed84653
z2bcad68beb987da2445f2b887c003cdc85ed2f5dd1083726a57fb5ca6106034b042a5ce74a0406
z456d4909ff18d8fe9498fda26a682f97e337255d0ea68b07dc4364b8aa3673ce5ff443b6145732
zd6f676c6c3d24ef6db2f56a29ebff3dc8ef82178e27f314360b123e4b664fa663b40197936428f
z52218f8cd4b7a08a5fe920af194a9d5b37d155301c9b11c1b6b818f7d3457f693d66b9b9869d61
z414b9c5a780f551a5bd1a6bdd45ba45f0670552c3172a86ffce2fc049d4e19b8ea07fd52452e00
zaca5540a2632d1ad86db1473172de5571b1312200a6ae4678546a7b8e0147a53b87c291c41e4f5
z2b8f3683d39666f6b1fb7998cf7ac6584c5465800ff831dd28fe135738650f50ac5afa395860ec
z394bc6ac02531910a13c94ec00f85e8ecaa62ba4c20fec86825da5cbd0e0a2a2d2c0e18092fcd9
zbfb851d05924e1fd8b1046ace863f6b4195dd8fc02d5a632276190ae8cae51ed1b8a9c99964892
z7eb6e8f7c16905a24974796952c4f8a3090821036c0e99b3bdfb51abca67e8a8acfb9d81043fc4
z5beab61e80494ba6991c8f6c9efeba146348e228f3ec277bcd45bbf1945182b9acaf1347312f75
z478d0711c6affb486c3d5e4aec60a06113f4ed63cf7d9ccf0d06e7485a7b85f0d02e8c26838532
zbb42f19f18bfe438d74dac72f8b7fc85d03fb8e94155fcddd5b68e2938f87b9670c407db8a2306
zeab7001ea821c7941f9540227444bc00fd6760463f6a6f1dabc99ff8fc4a720b515ba9f7f890cb
z9db5ad2c2523a987833107669fae990d24806ec5badbff76caedac93d9be568a703d0b4543f004
zf6971036dbb9d39212664c8d3b24d7ac9b430a3aa5a25a2b5ae62a778e1c11edbc578e211c7628
zbe735f984585a08919808389c774cbd517d7662bd56a1b638ec9f4533b51b62ebe5b9774281ad2
ze1056b285eb4fb36fad3a2d6af6b9c4c3fcaf3cf6e9e5937e81262bd69b3915e2c96c103ef8237
z7d3c55c162a41670925e9373a475bcd4537a0b25567b6ac443041ce8197f910ef61aa99bd7aef5
ze1818ccaa0f484b96536b3b468d95b35bd4bc9169a330e042697a131fcc825b0254f4c2a9d8da8
z70ea16f7a64505c0e2df9abe544c4f8fe7d582d916205375cb6c97a3b0151ef63e6f0d4a32db6f
z24a6de304ed4bf376d069a28501f2d915592b7a88b932f59ebf73ca400999be902ea253e0ed795
z6c8c72a889a93ac6c6d3935c3dc07bc64c8cbd22f927707f15695372f3bf7d5453e8fd3d612cc3
zcda9abc4b3b5c1796d3054fd8d8f8acd8f77f1bb632b85a9e2a2123aa040af399549fd1f6de0b0
z5fea6bd946f379f3335202e2a5258c2a178f1e85f42ad46b328af97c92cd9ccfd96573cb4dc5e3
z810a50722a50ab3d6753d75cb8be5a77de66b20b7e1a64db0ce6d8ebee90a0c5e919cf41de9d86
zdcb45e12817e364cb93f318237142c4cf3aaa59382c0e6cd5a286110f46020c41a4c4e08adc397
z2b342e6e9046ce6e5426fb69849628a0dc0121a8b09f897a8a2ce3e7319441401cade0f399a3b7
zbe2b02bcb0fcbcc0090068ec4ca455549aeec7cba0c5d2adcbc7dfd8b58f2911a7cce48c5a3c13
zbbf0bbcff0c7a7a8b175ebd86cdc6858bd10de8fc65b168dfdb3fb1b80cd4d3462a56a2d8168a0
zc31f44a73fbdf414eebdf439081f4a8438e8793cc8fcd08fedd333926247a4d5a466a1e1fe2221
z781d457d20f1f5a7be6f6f9dcb29272ad7684a01fb9da33d70594305cdcba43b2de3bd36c0c3a0
z86edef513cae12e61ce73430994d82b715aa099e497a3f81621e857213e21b59bafc1013bb0ac6
z092cc98c05afd602495dbfac679649b9d3e3ef935819e094b0e0fbb214ce6103d29a60fcd22fb5
z86e9566cb4c11e058fdb7b8ab6aa18338065b0de3b6aff39d2ab8b114264c1263684596e653b8d
z056a243816f4329d6b27ca7032402871f5200b1d077ab4a2702ea9d905a80105b55debc93f81e4
ze409c1c45c6ff43721fe5a4e374a76608134afe73c720c7323ac5900ca3bc1b1071cda6f923b00
z1b19895ced96937747e7abbe43dee0b80358aa45a0a57ee181e259e4aba4adc3fafc564bb842a4
z4d2c1da5e7dd3dc56fbc8b332434f93e6f9fcb5c045cc31d4e179108d46de6c3c3739382324991
z4c5ef0ebe09fa9ab8fbe148b40e05608c456212f0aa0203e39c3349f973b604f798472f0a24a0e
zaff9aa3ab9ca273f99ea8a72794dae12dc086f2a828840576718e7231cf029a252e9290076cfa8
zab24dd821aefb1dad7d3d1724bda3f5f8f9fd66dd561ba68173a61582bcdc3f0f5f4eca977177a
zefb367b24738b34f371d2bdfd3e02b1266755cbe99f71c2a6d37476d8096e2b4c374814e1f041b
zb7eab9f6bbb5eb4b102da32d1562fe678cdb437c5ebea57aae8ea34e588106ac4008af48b941f1
zc3794639debe578a1c67ecd2eddde29c6d7400dc74f5afc96ea4db0808cb5c6ef7122512d5d1a5
zf5375e1bcb7fd880f39d79c7f8499d0ade23487e36d86bb3fdc233305ec589d1e1dfea9a4ea586
za73630f9e00330d12725394507801dc719ee540a192ee0da8a2cdfa4621834a6e8f7b12a7c536e
z3dd68f27e1a4e71121e9cb375c1f68c65916067346f86c69520210422f91727dcf229a5c8ccd31
zb2ac1d2fd445282a0586c16bc057300993aa2201ee0b377e884db1e00db1f9f9cc2871b5b7a300
z3aea598462dbe7a88571bcd8e3c81cafafc31ccb41169929638defaa2c3a3ce42c9b1a2a2cf9c9
zd062cabb76e0f111bfc1aea8533e852c9f7e0eb9a42c089a814b03499bf960fbd52168dd8e49a2
zd4fb1246e84767f42f814cc6d963daa95da9d5f86cd6092ad1c1b7eedce125919c281fa7a8e013
zcc7d75cab92e3ba8b8224e962b98307020341c1eea1ec22ecf36d5d2c075eff2d2522e359c22bd
z4cbfaa5983aa577232f1292e2175af073da04742124b06fe8265425eec13e168238462b78f0a6f
zcb9a28bf07ffc7cb29e8fd781226eb911209f45014ca601b1de31a6cee02b7f359803fbec0c85f
z7c549fcec61d58e268026b5195fa65d7023eb5ae34e0575e37e1a18235856feedc81da6a15c431
ze4b55fcdac0774b31e12e8fe8e34e13805eea82255142d9077f128611d158b09550094baf13d58
z51cbb98760662a77518256714bf291105e92989abdf9140c3a4c59034eb79833fc6bc390b7be76
z53dcda63e18271d21a423db4007ef3080e756acb49e3d385439f86630070a55e1c0377af9c01db
ze18da64e7fc2bb54a337e1d2bc1060137e741ac5565ffdeb597c9821fe29eb21a4e4936002f72f
zc0be8acc1fd8621ac14f1640b3dfb37084e64a6798fdf54e1009ed63ace1a596e6405ba4971012
z6dd185e1498c86fd30866eb2d08220d19d89e66759264dd3cd20e73a001d519e280e156d78ec9b
zcff3f91d0e0f4a88115def790f41305e80786663946dbea1940d72974cf209ae0772ac4e5beba1
ze932c17e9a0f7f7483ac544ff4bfe97bcbd840b949145b1697be0a07e1c2dfe57f15b1f242b4e5
zf4dbceebbb11884f908ee6cbdd5fb187c675c1c53e7f8b85db14c52aa10a138500e4b5af7bcd1b
z7c3226a3faa2665741014dd2134538334004605c73d5c6cca85c33d374690875c3f102bbaddcc7
z427b9dcafd086c47708fea1af7fcbe9d6cc8adbcba59024c33f5b8ccb06a2bc2a05eabba0756ee
z668a5fa9eefd3874039d48bcd1f6e2381ae68a3b27f28a3df34f17ce26919949118fb9b4e31c5c
z2f63f5457688ee2727d2f73cc05ff9a913cfb91c6fd07c77278748f0d04c606b89f5e25b1cc3b3
z3ab5a6a18fe9c75adaf113f227d47b122e8963211c8236d582f2c4fe4b4d25e70dba2a902b1a5e
z345267b89dfe7b268a6d5c3c62343fdc72e6544706709134f467278aa031dc23dfa930b4c04336
z898c86c75ee4a6a25fd7dab86e50cac8ca0ace84c9a630217d7efafe2976716eadca993b4320c6
z82e168e04162d36d4ba5b4627d10c7838a88100e8ca5e15fca255485497a8e47344315ae3bfea6
zebf8b254374884f70597ece40b71f00cf0e120a8868f0837ab13160f94b53ca6a9bf0e458f2e66
z1ad7cb9d7c6b356d0bdbaf8088809b40961f8b1926a404ea6da417fb15a53496ab6bf412b528b9
zbd4fe50a13d3b4370a1e5de4c1d24c30aa2b7c0515e281b41be0c082ab3c1b3d83481dfb7f66bd
z65665be82f54a8e55571f3c87a197cee4ccd1f02e591c2013ef8faf5437d5f4eaf0d317066623c
z484e85f868d1da9b7bed844eb25c896394ac26cad569388ef35e479992b2ad2fc39aa56814a08b
zffab4f00b485e7f1802563b3d0da41b32cbf659574c107f774891a5493ac42875913367f9849df
z9718972c979d30d79c5f1ef54f31b69cc972dc51d944d714ab55f906177787f6461770ff61fe9e
z428d121f630ecff05e19cebd0eb23803a1397bfbcf6365bf6e7fb6803df7d9f1c341193c521651
z4f1de091a7022d2df4589ef313d210a2e5e9fd7ad09a895e950b1511cb620ad7fef2c8b0c66f8c
zd37b8a8a59e0f8036357a3a78d0f8d66d268f479b41a35978aa635547b42deaa68a3b8c3695c36
zbd85fd4e68bf9e7f2c8c981d5f7ca32421be455868fa0c80ed3caa2a50663645903d4106aa6688
zc15723da1aa45e92e6c4c4b50979f037be6fc6c09e23d13fdc38a8a5bb51df52367dd190312cd2
z7baffe4399bf462aba7403cf8668d1810172e4337acff1e24f5731c8db062b3fe129b3462f7f8f
zed2b6ee48de37aa46317c41969012a6b16aa2d540357f6ec4bcfb66c79816115cdd4a6cf3ef47c
z2273feec856922876e3056ec96832e29917c825320f064ba15c7a1803f648f9a5b4db7a5d55931
z2438924bb0e0e726c8206c5cd8d4df19b747121adde574f13e40dab1be042bb46ec62ee919be89
z650bb88795a76b8f3f1f7e1d1b04e0418610ece63ad55decf3fd860079b5708106efb23d1304aa
z420aed054d931f2eb201ef029ed3a5ff7431524c69586e80ff35e4f205b662dda8c9fc0e0f6ed6
z82a809f9319bfbc1c75bb6d557885931d93a72ab907f9fa54b17c484834d152bf2cad76d745bf6
z2a3082da93edebcc40c02482ad721003eb80782523555b5c967fa40463ce9ac657f0980bef9495
z18a574f19d5c920b05a16e1f17ff16fa0f1285b712d25fa253f87a92e9036c2554d3e15b83eb74
zdc25c8e52470aeddf3d1517dcd808a05d2d68c05dc443fc5434c2baf63919ba3932ecb60a86823
z53adace176b709ea70a5657e375d406afff5621a1ff92f7594cb5720f7dd7f06e090066814d23e
zedb971e59557abc8b2b43dee4a4b66999fc5d7ac0739683d524a79cc51db5370231c959cb59671
z9f80079562d53188758721f41d76d1922b5a856c90b5886d9dd029fe8c86a521be1c15aedc840e
ze0462b1bd7e7b8e7a43cde05db1ff66d01a653cbad387b5def7fabac87fcede12a42c59c78d2da
zb5f231425c58c7d2e1d56d1ff5922944eec310a5bb5e34a90a550a9a0ca2efdd845310d45a6672
ze82890edd46c457e6f4dd813b16618644e8d783928a593a619248ca0e9eda68421a14dee399ce2
z54376cdec3359e5bb5b09c25af65f162e74686a1ac3dc0f62a67a16272618e18d9e5ae735ffc6c
z708d7aa679c3e9ce273df2851fa61e49e52eb7e1d97c41715cc00ef22c4fd0cb7159aec1ad0275
z02e0d3876e8c568ed66099d3da7d6dbddbb0d439c00d63bbd68aba6769c00312c150f013936e79
z59c7cb66b114e9a2cafd85047eaa40fdcfdfce12bf09563d995529158bbc9c7c7f3f954d7d4f68
z24be6218bf48d5c45eb13bd7036c79877bad8a0e3c1b8a1822a11a8a1a857ec24e0cc4e902dc35
z9bfef97e963d711c3572ed34c508abce74d1ab005871f624b12c18eda30c95de8859ab697cd127
zdef0c9a0525bf36cf840407886351fa3b61762ca2e89f8db33a2aa945171601ea11410de16d7c2
z403b3565e551d501a69297c10c7df3077596810e759a57f81b6ee1d01715f55c026457a10550ca
z6b3b40113e332cae503d038f40acdf3ca595712c94233e710a2567c9c54e962c88092264ac76e7
za7e588d2581ac8a9ae8e34f88ce55ff844be8b3411f79e4645966d43f8f301826a519523ed0f83
z1ecf0a1564c888c0b55fc7d69c29313ad155933b2e294d13a892bfd3c4f876da59c62455617e28
zee3f3e76c3d3f5e4528bda43da1351fa16be47ec82804f2e6580d9bbf80aa367683c758e6f95ff
z5c6e2bf16f20a071eb50d0f9b910facb9e665220aff26b65fb08788a6a368e89c94f3a1de9b2a0
z8b2e1a17ef0c1af99f3f43d2d14b0654baf834315462d19ebfa1d6115cb8e50ddc69e44901dce8
z6d73af62690513ce4e7abac119f93b5dcb6e7b26d278d72e5673eae6a8f0f320e949c11b620410
z5c85280170160d259e3e681ca0be5c6d7766dff27617afbf876bf069d2557b60dfe9327c2665ac
zd36a88889c77e10aa71fcf1e58ace85a781b0035842db8feef4c6eb62ee5763696dc477124f837
ze58b0e102c9a3fadc99d7c504a4caf55c512781dc989a6233812de6d4ce6d6377461e1e248bbc2
zab03461c73c67c06c0e19d52944ac9cf0c81c1484fb45adfc64bace96712c14569274fb8493057
ze8b61749961607f992d6c7efda55ee5cad3f9c6278abff60fd15c725a9a779f73d40c95260f74d
zb88ad72842f22554af52d1705477425d7def548d79dbd3aa6f9bda9c7bc177af3ab92c8d95a7d0
za7b981b2517b2a2923d121be6e0f581eea2e7f4a0da2b0ff70eb500cd691452d579a80834a7c00
zda311a9a603c567c73e74316ffbaa1b0434a757b7a7b64f1a1aeb4584f8b305e625ced99de1f62
z2d7550ebed170fa4a55028718fd2e35663ffb24cb927a62c0b046549b5827381f58e2ed536c353
zd8ccaf0fed8b79af821ff84003de6075480304855cee1d2c3dfbc0035ef13718e9f8505c480e82
zdc706f717c5d867c51a81b4140ee6486cc8b2dade63c9f021560c6c5d74acb3d06f8e0ad9ed9de
z26bd0cb897c66c6ab8620549141e875e49339a7c194a583fc6f46b276125871a78a6eecc7d4afe
z52ddb877354cdc2dd38060b3da4e7b7e6dc6f1577efea849f9f1ce7c58310eb42ea3534e29c1cd
zaf5b0fa923c85ffe342bc8520bc83967aa72c7c5514b5cc08931d590f413170e053c2fb02cbb5b
zfbd66f61e424f6500d81e7d70c82c46bc562e091963754c63823b4710f4943943a0bcee48e6d94
z6c3e74014179d2b8fb1d81dc7a0f0698d8572227ef31a4155254fdc754d2913e590f6151c5c9bc
z8a91dbe08077aa8ed032f007fcfe2677251bac73e7c6b08a2254f7ae75b4d10106eb34aefd2d3e
z303949786052c7efdb89eb3f13665955b5b750afc7793636d15c5ac6bc2eb45dae9489cd76e1b3
z9cfef9ad7262ea8694bd75c0a1b7928ab30a3ca466649795a610f5aeef4e8a4f6bc8acacf1f1ac
zee4c1c5ce7f6935fc0df55d95aa43e9f25d49ec153a3b14388a5954ee8cb611e9c402184a85f84
z29caddf76ad5f42092bed805e3fe75f1b4506b3c0c65b15db2d9237d73774f1514e33d95356ee3
zb34bc3ac30e65d9d2eb25f24573d5b75eb85f61186faa4fbbd5465b4feb3d42a14acd2f176f3ed
zf3c882af3eb12b757be0da20d2a11d771b6b5cf5c125bb5813f58c781e404f0919b3b3d9a9ff5b
z6d7ada3e6b0369fe9895aa636f701c3cf4a20dff7d45ce816210dbf355581229ee6da9e324c208
z466e5e706bf278a0f0b6fca42846c007c2b7c506fb4a41f84db24367c5a62929ca23f171b8114e
z74c339b65fd607fc3a5021e1b7dcd4ca6c7d1b315bf5fb5417d42296b9aab7d24435c49ff0564e
zda72edaeb691289b7db3f509ab335b4f62c9970f5fddf904c952b0db9873715ff1886a472238a7
zfe6b01730c74bc26c909e000a8d849649de6d0aecdad081ddfcf9fb659328e9597dcae4b0cf552
zda0a68bbbf1520335a4f5193be62051ba3ae3045dc87beafb324d89632ec83049aa081d8521465
z9d2dad722b046b964b43981c83d7e6d4c44eeb35cf90f8b157a3cd47a039eb2bc47c80ab4ef773
za6ff8d4e4327447dccf07a49bbc7f6eea590bd588af70dc617579fe7c342ac260cac84b6fc371a
zee348f1bcb617e32edfd938e66d93f1c3016fee32a0d12b1be171f7dde51104d548fedc6d04685
za193844327c000a5fa34aff5b35decd417caff1f87fd9e7f6e3921980cb8a95a6d8f0fa2fac2d6
z7ac48418536a9fed1b1970a407ee38a3b07e50bc5e83523e2aa485c338092ab7681004f0e57425
z8d4ac47bcd4bae609a875cb75058439243676a97c29766830e97acb58e6acc8c14f2f1db63ff04
z1f5ed2b88dfdab7d7b7c769e2a1797c2edbc582f804e6defe99e0c8f0d1d28b7882253cd2ed15f
z62304bfd8d0e4041880d9af3f14f8886dfbb8802baac0ee27db37a559e8fd29e7ecb480e37f7a6
z277d1bbec2c840e5301dc91284429102fd447700bac9f213a67a115cfcb0495c58425024065d1a
zf2024b1b6bef33dce1f7be70cfbeca702b568344d58fe208bace551dab229cd97085c5a05afa67
zb4771a895852604c466cd8571881bd8b60d82facbe22927b9371eeb80f190446e36efb4d2baa71
z2388a3c5a79b780e22355ff0c35ca2252c305f4b834e287b4b718990d0fe5fa50f45bdcd65809b
z15a26c9a22540da5181702e4392c6b9d0f4ae4325c39c9bd06c9d77305f6a1cbec6c1cc701f107
z57d8a3f93ffa9ff1325e927efc1ff083e61f23f73d5384d35b97d9f2c0d7a70cf467dc2eccdfe9
z9f0811403d7948855dab8b73cfd4d87bde151d0eb4f62046b98b61aff0dfd439964d36fd6ebaed
z54445be6b0ba34db79ffca8df9a9936ebca9f441e46d6f32db491c4fd0dceb85f69701303f7417
z447b366fabc46d9fc7af172eabb0514e2eeeb69de8355baa4eadf93963b103cbf7d4d9c03b7171
zbd0b7aedcad8bd1005b6825ced347578fe348e1ef1cdd02d9f0cec7a5c44c9e8190d2eb6ba33a2
z6cd362bc0d43462b3f9ee616811cd210f02755bdca06aed7fa9a072ba5402b1f053cb9bd38ab20
zeedbffeb6289a26a1722060298ce536f8e3e8faf433982f18bf406a5e7d2c55c0def178773f11e
z644d3f1af694e54ab287604c35c6cc7edfd995746b698f99932a1db7803c95a47f765767cabf15
ze786544481d874006cd0c366e7c5ecf933cd85b146c49d63588e74d78dde14a0558cea2864e82e
z2506b6dd8053552816f4fb69e8147d4c596dd4a3136f91d20785986e0a7c43e4a34f59347a87a4
z7f1d9a88e1fbfd6200f08de4014d6539f533aabf3338d66f439d5ffd97977ee42088bd7d9c2862
zbf0511ce75b994e4f437a2b8fa119ee76e77eed58ea0a32ca57cfbc93d8f2ef7f6a178f38e76a9
z716bc75019a4f8f0948268fdb73d427a49546c89b64a2de4c88c4ff08fda1b4843a266b94cb0eb
z54e4aa0cc1d3a8e6ad40c63ef5669822c7b08f06741deb29fb3914d65b2e86773662254cee8d57
z97c30a6faecff119cdaec382e3902b7d12c32a3b7b473c3adfdd6350d4449dd8e28073d6db1ad6
zaeae70a5c459bc48672f7c84cc2ae3a93e4fa6469651f917103fbb775f1e9da58d4183d1991f93
z967f93c5bcdfc1856ca23419b0dc4bff49f34efbf023bff25377cff1507a7a2f2086fb60bfae7a
z05c9885013986084edf5fa11d3a4cb972dd6fcb109a3c74630d335f9637d84544d696adc81362d
ze6b5a4f1a68649ae7e1d58435704acd6c3538d7bdbfe1d2b9fa47ec98048b1914b721adeece9a2
zd3da8a6ec113c200357d47e99af3bbfff1305975810f11c245ff2e9ed031a301d4d7bae2a3ddfa
zc5db4f528de880d85a201fec97fc53281c7e74fd7114fecc537f471d0587cf0de0e6ccb18978a8
zbcea1dffc57ed504eb725471bac1282bf03efb03909d462401b783f2ff6bb6a60ce6a428ba43a3
zfdf7547b2e1e4c4a1afa018f4c8defe3dfb8cb10533847e404403c80c05970b6c436cc7051297d
z6045de8718e085474208932ccd06c618798e2544e88e7873b6905d79192a495943d1707387fb90
zfd2a9255f83fbeca90fa9922799218d4878cb6f6248a02d34e90cf50f961fca6fa2a3718302798
z08f021001e022ff8f0b9ea89cfb19beaecdcc458bd4a4a9e0fd3acc69764f338b5fae4e42e57e1
za46cca4f438bbe08cf9f4f48c9dde1d41f5595b2132c9a01f41fa45245e1b3418350ef7d721448
z1a2f20d2326cf988e83be6b07fe9b20b18d37b5317445229aa07ddfbb575aaba931c85aec6180c
z73cab01d83ccd831c922b70684e605c3d5e5a3405f1de63e8501970c1f9978bb044797d25706ba
z9bf7ecccbf49946d1031b89ddc83cbff55c7f6684fc53df8ff0abf8ab15c102b1b740f7e237d14
zb15ec955348361ef3987f79206fe6bdcbb2afe8383faf1ac2186d9c9cb6433411de5414c190e4f
z4da1c76c17272ef026cd192c3979a3cb2043a2b076e8063f14b1484438a076718197ecfc28b65d
z1ee35ac60c1eb65d64c073c4e9acd45dfec10fb6c513f3cdb413d89eb1b1295a4f11d43f147978
z22c186d1f8f940a8a74147b7815173d9044b000f437ce1b81f72b8b02fef93b7b87018348c7e26
zc5ebbad42fe95239da442e243cca4542e85c59fd4e6fe5d0bd427d56cd602092105cc360d4a46e
zae610735ba0308b8ec467c45f0d80c4ac309b1e31355980397d5718fe0a369260998dfd87018f8
zc0393158cdb0335474d23a91ba1eadfefc2ccd29ef7cada96fb7f067fddc940d8500a62dc50f50
z4db390081890a7bb794b62ec0271407631e5799bcd48da426ae874b5092dac75445cf59e5d2442
z833b31691bbc8d08b906787db075b0403aaf4557f258c78ae9aceeb47c9eacb30aa2cf77002fbc
z8890f58661492b56da7f8e9a359527264998eed1b17e17e5a9134be04a41f4aaf92339dec24062
z96ebe3a6a7936b43833e67105595085d8ad59aa55b1d8515f41f012fbfd217f1bddf6331260a91
z1eda1649b76d97c1d2de7c4bc23e839225e414e4fa04c3ce128136abeed4d04467554af18f0c39
zdc86b1622995e223b53a08f788a02316136cfcdb451aaa874fa88d8913bd52dafe21aad8fe44ad
z4c365917094a08ba5fc17fa1865ffeb174effd5e72394b8c8ea830c69ed230b2895bc71f64d70e
z7a53db69b8169eaf03376aa99015a940052c087820c8abee8aff026989d96a3d5e1f67333d1add
z0754bd09bc2aec1b90e2ea9086022ec8df10c19bbd199d6fc91dc650cdc38e7a31ca8f45775bf6
z4673bebf0ee272f6d5bc4208a0ca075f976fe18a28fbaed7321eefbd608f1e38bbae43dc235fae
zad2f651332357fe043c97f9f3ad2c99aebc2e98c170baaf5ab9c2375c05fa8fb6475d4fab493b7
z878465a3cdf31b3762ac7009e0e7c7df6203401f14870ba44ea7fc25d9c354c0eebf2c06ce4d47
zd2d688749398f5e63b0f88a7f213a4031c2e2dc5be539401b9073a64117196132aae71e3ac452f
zae27617cd20a859d43f944c27aa21e9c4553d81fffb12fdf9b44ae631e43ddc71a395603e215c6
z69382780d29ba7075508fd099a6b6622a768c8c98868eb9345a670cab7f2c269d4939e4b4681d9
z0cde656121497dfcd39111ae30a38900bdf73066c310cd82306e9559263410a6370fb61f4c61d9
za7a5c68f8f81977f58bc256be53c19cbc1061e58aecfd3f70c296bda64401d33b64dd882d4fde9
zc1a8a8e3fef2c0e9cb2c87e65c91e927c159d29819acbcb705a234a5798e9c478715ff2decab1c
zf26a32b30cecc8168ac373ae67bebb587b077ec1a62247faba772e54858ee7f438fc69ff18062d
z00a5b2c744ebbda8ee8977ecc3ab5f0d14894b1bb9623bb4b7e15a1945bc47e68e1630ef04a2f8
z7dc1f8fb3dda12721b9acf84bdf80b4bc2ab923886573efc64aa7844dcdc7177ad391bcd06198c
z84c22431ddaa95d036143f7ff9b2bc45ce67991cbc0db5c0ff6e75a610c9eae7338f1211180769
z3d4f76c91d3f0da9b61c45e5244aa6292efe1bbfe6d1709bfecf65194098dfc13e5903bbbc6660
z2c29370e85b2d8f4fc4ff80f43629e9c8d81062ed7e3c3435e42336370a830e6fde61964226b7f
z4f1bac1bf835b775ee7c889f4abe73c48be4ef0722dd9f9c9db5273ed237aa09ac9951cb2d9b57
z269f4eb86e897046648bd0a012d28aa80ac1cbbff43e2414958f7e32c1fd4044de8b17bee3db59
z5881eea358967d52943984f409909330acce38388e8eaef504512cef4b82eae88e836822724d4b
z3970d6eed99cd5f664c708256799fa8d5c6531fd80bbfae5cad81ca196f8e2f597eeb3cde4c9bc
zf814d3af302b46461fae885b0a7e8f26a5aaed0fc646fedd63961f9302efeef30067027f5c741a
z07e9691ad75d7a6d2e19f6607a4605b6987f5b4aeb04e16da004ba5dba05ac4de4375a52470a35
z6468e4066f40d2ca99d722646a84b59df1a11735aa44b656f97d065f71c29c03a626f77e6103e6
zb7c9b96d7fe7d52b5ffee79ef43144238e2b63f71b05343aaeed6ca41693b6c744929d62ad5cbc
z978025f6eb7e449b0ed7c6f3183e00f537dc3659fc0928b7ca189e7b9b1714fe9864df74c82d3e
z60272f54fb5cbf68fcbdb6de014c70ba3d407105de7e2a67a561feb7d702b7dde905f62108d6cd
zf93d00e7a2c6496372b8826eff827657c3e642623d45082f08ba90852a4350bf3dafc4ae02fbde
zfd6b826d28a6064b8ef08b3426e463d7881a67769673134ab1ba16f89180de3f0d337e82139ae3
zed29103697acd6e93bcee3055c37870919fbfe3ca2987ee6ebbe1f305293c7f6e83944963673a4
ze0c8b72166d99710a9d168246ecd77a074b0bf4aa4cc9a9000609bec1eecac967589e4a431c64a
z02973580d0c57745cc13a494fa68491781535f81df965a72aafac3130a713fb66d7e8ec3fc8f2c
zbff3897674b188900198d31c27505a02c83e8fe9167db56111d0deec62d366da5505a85afdc9d3
z42bec8f9f2bdc434620d250a01d460620d76e67109f14a3c0f39f27cb7b0a47353efaa9e308216
z0b9c2cf7a38f2bd8fe6ae463ae5e851fb12d268e73672841f82c3c35818666ce45ab864f2c0d59
z723840726c7cbd4abd59538dd296f9f8874670ad865a543c8abcea974a7eeb3d3cc7d04b7373c2
z150afe7b94ad47ccc06527128dd12fe23e2c9aa80c6a37343685da9bcfc400b2629c8d975462f5
z0e6812e0fe8bb2d7248b0cb5bded08d5e53932a76bc64b0007520fa9bcc2abe710d456f84bbced
zb63c43a5e8ca2c9581ea7a50312ab492d3304dd06b7cf4c6f769cb7c2c7b6aa81652bb1d382e3b
z50829dda3156fdb64f29a88c4aabdb5186176a10f8d333628faf9c64fb77b9fba9c0d476bbc552
z07956f482eba27245f0878ab6946b94b9ca577585f5def33ce02029611e36974bb980c742435e1
zd1732b8e1b49377bd7f168861414a2fbac841a29496da60e7f68ebb5736bbd436f2b71f0a780c2
z09f8354e90902a2f424b29e91d9d19b99e07f278016c8b210381169f2f5ba878599d14d6c76434
zf12207fac9b6502dcbf7be42a29c5bfb50f132a04175ab85b07aa61152ac68a30b8b7bcf6a9d6f
z11021b993dce64d21f86dbf5cdcfc842029de27db1c8eb23f13a700c917fbc4fa165f988a6c2f2
z0a55580c3b35c5f976a2a7f55a63700f1bf6fb01db93a4635f620eb9adda78a80cee85b95f911e
z4f7f47f30a22a8561fd6d2575fcc364c4df465b2fec0b13b554d24734cb17dc07378524ff31fa5
z3c6c4ffcb280a531bb4b59d98ff23a45f3498f77400d534df5f2ee0c1f19891ba1e00d2fe88943
z8159871b5321e7a86daa304118baa0c764c43bcf689ed91fff7ce6bce4f14e4b428c61a85db0c8
z023b6be9a5cabeb3e30d31de51783ec947a51f08a2cc4ecb98a6b837967674d6a870d0fc5c785f
z9f7e0a969dc98a39fc62dbdc41e182e2505fd1ecd78fc107f915fd1395a55af020aa9da45d8a37
zc67257525d26282db94d80341bf99df03ebf6886ba0d9c652bea11ebd40f53c436080075e8dfe2
z58cdc81cca3fc0cb26e24aed7e07319f5af582e465450690299c6840e4bcc601426c6a14964319
z44b72c9951f73836883ebd96d1792b472b132cf982b9f6730bba8f5c30a0bf9ee6e10198a3d1ae
zaeb106cc9925bbab942cc5fd0806711f3534b666f1ed9dcbe32d2767421c7cad6c07a5a55f9989
z3b74aba5572b40692f7d4c7f723b67a3b02f4891aa38b1252090305b330faa2d8490c578eef17c
z29f2f9412db0bbd46c907b7ccd3e6bd235eff136d6c3dce884a34001e374797ee1aaf8e6bd5876
z9199d426eba91283adc2d562ae9ee9674c2ccd9062fc7d1a8d0aedb7d6f361e970f6f3866289d3
z386f2498d520391c4e6e6f8d56d186766f6be8159717178b42a114be266a005c9988819c7bf521
zd8623c2e4d8d91bcc78ad58cad9e7b476e8e32e70435b06d2a23e3bb2691eee10135c46a478af7
zeffa126773e1380cb679db09d4105c1e8c401d7676c09d11d57321fe664dae6c6097915570e8c0
z9e39227bda7f42c2b2c6b96aa9801857e1d31982258dda89f984104ac977ae66cccbe40374d7be
zaef585e17366aaaa082a605611855fa4acd6a0b6a803492884cbbe6aec60ec0dc8c5f8b943b84e
z42f8b3009d687e444fa42eac7b0a771c5d5c25c94e7ac053fae62afa75e9cd45aaab1932e13988
z94a33a9d71fd91711c497209e50579d83defd5d9ee538df288a0448bf350322677c0cf4dece999
z69189c9601077282efad8144a6a3566bba4be6309e7c3eef37891e09a22c28fa637066648342fe
z06b03b3fd7107f37f74f892377e7442ecbd9a31e6a987ce2a4d4d73d5b7608031181576c0f944c
z34d8174474bd64b4ad75856f55a69ca8622ab838ea11f2d8654c4aa84ba63d51b299b519f90fda
z3df5237fee0f408472726d6ec252cf2280c7b84359bd4b11ca070b5304a1de5daa07cb045e1802
zb1c3d5e61de1f51f81f3c3eea10cb9dafc3d3134b1751d4583ed0b4586f14910c547da0aef08a9
z1a689d4f1d8091a21fea12126cd80dc73c1c51aa6e3bc4c9f0d73882ed01161d67db11a86cd44f
z89d56b3591c0a3aa659905cb3dd1de2baebac3a7945e05323de6e7e0da2893ff7270990b0ece7e
zbcbe97807bc924de66ec8cc6990c9b547dfbf59c437ddf44ce0aed8691ec93b60a75e2f703defe
z822ed858fdecfedf80af5a2b364eced5014860ed4e2f90bcafece3302a236d69489a77bfad474a
zf11682366410217f3bdf8efe767c906aa434945d18b7562c1963a56791d482f91e7bebe3cc1412
z40d642085ffb0dc43741be3666643dc4c46449f020a1fa68df8e5658406b8a5566a4fc066906d0
z173a6d2b66967ee7b4176447ba772d799926d359aae2a2698087b4222427a8c24f2c9e35e57b97
z3a773f352d2f10e27f1c3c09ea2afb42c18bb290ed03c63e10329c571756e5d62ecc27f091951a
ze7dc403740f7181f6abe0c2021db94143c514b29ea8be00efd7efceaaba465ed8089349227c198
zc51e1d6918afe5558525f31322219eb36800d836f20baed5201c8703bcadfcf7db33a57080687d
z97eec67bffe9933fef647fe011128c2009d5882f45833e6d76400789da55d4697e02300f22356b
ze9387ac4b615f9bdd0a320a288d5409b48905cad1528651157ecb3db8515e8d40441d87f745849
z90501c53f7a944c9cac837c25696740a9f37b57ab10200c761eabec3de00b88a75af208ab776cc
z75e5bfd906ae77d43de79eb8dce04716be53b17f6d7485bb7c95edfbaf1a20a34613b0801f2e3e
z3495b8032ea6438a5387fca67d1506fe6cfc08ceb4b77015fc541b897acaedbfd6e48eab7e5076
zd98ec8fdd27eaed2332e0ca359685e476e369822a2855b940b37fe0b33e60cb8ab71a28db6d2a0
zbc07e9b4dfcb654ccb859e1a69c477d0763c44e3327b48ec2b96bc4c1174500ef60094e630f29f
z00dfad9c790d2360417b130c7770bc333c7ffa601cc0a818f2e9ba65859440a58e6cff59af6cf7
z5c74f845fb4db4667f6916ee82ccf9525e3f8736936e2fb489bac6d3284a01fa1638ddf4bca6a2
z521e6e9c010abb3613a60568c1746f4b4ef6dcf556a9ad56d551e20459b02130a35f21a0acb13e
z920a8a738496011b1e4019f25cb564226ffe941482bf9123f3a80eb31a127f0bc3125046016819
z3ef44d532e1baf2bf2eccc6b53dc0d9f2e178845b7f8618008bb505a2c2ba12956ad1a794b50dd
zfaafdcd4516b1bc253e1ceb6ac3e6d5b616c4da4d0c55210a203a23f4f9e2b4605e90552235b1f
z1441e3b3207cd84da9f8b12562b74879b222baf069b1220e2348ba64827669c51b5366eb63945b
z7d9cdef98c387159d856b0dfb4c9ef6e3bdedd7edfc4c29dd5e9b964294bde782332235a6f633a
z39c29a1bae8645f832eb2dc9a78e15959a3cc064ccc2e9e168678777121d55b369b5f26311d878
zc28af1697f1ea65a85ec81f8d523aaa3fcbbd29a44190700b7dbef9073c7263ddde1dfe0197195
z7cda6f6aa696a5bf071b6d64830423494ece5ca312f1a86606f4cd40d3db3b8442f19a28a52559
z5558eebec7deb818fbafa6d77d1a56868bd56c20686063931f3c81165cb2df1e4a99ca1b11c3de
z56c5b93f593d3ce442e0119b35c23e54eb419d7000e7551a038e0fa715e5bfa1e089cad511ffc0
zc8d9008fa2742182efb751217881a1d9798a03cd78891f36c2a9e3cf97800737b7aa6a05aee937
z3e09ca63b73dc638b841147b3c63274166a314bccf0057f0d2a8a4e12b5a7dd3d80b9f593476f8
z8ed7e77cf16e9053cc51bdca7af061f9e5dff2d9762b50b649ad996675d65cb472f96bab5ed4bc
zaa1fc3ac99a77bd47ba4260d8b46ab196cba1b3aaa19480a45d29dc64c9a8e5ad50ee6acb9e57e
z4039363b040ce1f96b14a1eb6dba419ca97e0de3be81f63d59b2a89842a1069789a57902861322
z839852b3bada66f56b808067febf19ec3b4f9b829f021d4c5a7025969032742892ceb52cca03f4
zc793bf8016a0f2e6aac99eb04f551fdfced06d3d3e0c7c494127bae3904a63ab45431d0994534c
z3a86c793183d53b36c14c8d36bb793a3b9f5e72c875a3965d84f6ba7f88c043b3ba0a7a037093b
z32afe857527dfdebf249beb06e93dd8d1ca2a38d8a765314b4f51bbb6fa35c4c5ba8077afee1f8
zd1115f93787113b5dd4b8c1a0669c46f979b60f6dcfb6cfb9fa85e1be482d869e6034b6e2ee3c4
z50d0964808a3a938303f1b5975efe2c73a5ec524d00bc507ef1282f0ca22c62fdc3987e0b43e12
zd828827f6ed5c04d6bf6fc3f46e20077eb1cedcb6c2b08533de5a342e63c5148db8a93b7189322
z44a88a06f85193828a5f26a43a29ca64184802bad47b5a4831f1179c2c78dd8b13e52759e30d9e
zdc99aef5390247096346a4adbf046719f6b958c370ac51a7e01c6ab63bdb53dc233cf0783258c6
z7b0fd272c345fa91000fa9ba01e53f99aaa67367407b65e7cc55a7c7e1db51aee06956d716fedc
z5ade67d8eb42b7bce33eb4be695ba8f3c5e3c903e7287514a04a7f2ce0ed897f92ed40bf5498b7
zb9cd652426b1dfa2d0fb3931a97330e95316f3b4810779484398436605c45430cc44f65938420e
z54eb4867aff80f229379dd9e3c74ed2ef6b3a811d445fef2a71723f09a33ebe92a7a07ed787dac
z8b77c184d31c2e0c05fb53076c93e0561d7618b6a541f660a17aa1fb195d988b2d5f54ed266e4b
z0348f26fc76cc868b827fddc19b4993b116debda9c39263d0a8871ea8e5ebd73070aa0efb4d419
z1cc64aab244aa3de8794c60408e6ac25c393cd336256bc6345e3d7acbfc009e3b120a1f8348150
ze694aa046b38c79fbbbf4b3654c1fd7fadc0912da29843dcae49e8009c3c29c489675b3b3e0853
z98b0da0f2b8b5031f69b08f140bc2367b0fa07e42eb375fad03a49dbc50aa6aa25c14d666aa155
zfb926b8d58faa25acca4b394960dbc643dc9f28865051efbe0421ef09c3c232243a65911021c8b
z0c04ebe0594bd036d2aa213bb5498f80afe68e0558806ba0892d43395b589a28241b8556ab871b
z6c52dd651b23502af14bf6868711e82f2e6dee31696e2d3fee1301d64c1eb638e7735b18d9e8bf
z064070fddf19fa3eef71627e2f4fb32342ed1e7d140e4bf5f802be1e494ee098a54e01222b1ff5
zf8fa175b8b01495bb6a15cad5ba7032a80fe0e7c248d2d76c1533f7bf300518ecda60766586bab
z91bece8bb3661749546ad632d11385a09e4a7b51ebb4f3e23a0023690a2d0e1cca9976a98dc376
z1e07c557b2968acf19abf93230db2648d09f7f0f48b96fa9f087898c7ea017c00019d361d1a35c
z2ceeee626daca375f83ae619a55b2186fb090efd47c3ffe7bae34ae3ced866fe6b09aaa1481bca
z9e094292c928a83760b6e36249d709e9694bc7b5ca8dea9b0a0331f8f5bd327ef565c95eb61d0f
z05065834cb12c17693960e95ab301aea7ab9d8f49f95f87259ea5644de5bb4b794d14430ce937c
z71c81602cd6741e15ef29ac301facad242532eef29eb0a3798fa8058a00782faf3df0b17fec277
z26a4dd1f8ef17c9be3fc023bd7290f6db22fe88caa076b3085b4257cefb5df6e88262ca75df645
zdb176d60669d9c5bd429767a00b55c3f58021fa168e3ebef761fdd3f2cb3eceafddc1289299970
z9083f2b003f926288f4f463ec56fae42631a612120ac7912e287da019a8c2095485f4e60082abd
zee3397d2c24051dc6220b6c6d135f5ce44fc12da3cdfc58b08f194d336bb1f36f7a0cd5398aa99
zaf5d1bb0ee470a9cd4184f1cc3c2498a1066476c88bea35449de204851646c9532915f4462747e
z23c8abd3265d244271831b465bf1a5f7d9ed117f2188d0a5ce8fa6cdfe45153a7fb1a91c679eb6
zb2bc1d55b1ec41e5161dc8776d669112cbe99a90de9435d79d99e45db7d953a509b0c129c5a1a3
z496f4bf2ad8e973749d379acdb45ea785109867fc488753eda2b06ab77a66d457cf0d52b34bf41
z8ab89ef11925a265181f6dd8a4de3f44286c311e80038f6255c77e7c34f31de6b9a68320da1453
z5a3b583629b52ce72303a87c0bf5caea9a0ffb6c89d6086922b043ed25381393797c36ecbea0ce
z057ae7788b802984916aa8b93836042609faf686e8e11796e50324303740cf7f5d9690f576ee0f
z8a75f3e4c0f0bd95b74e56aac084035ac18425c475fb7737ede8d5a6b330643a60050a984157b2
z57e5f2790c35ffb874720a77787324537c8ff0a1a4747ef30c335761f3610dc8d2c357a375764d
ze8765d167ebb9c54d97847634c14a58e858d5f15aa743849b42316ead11ccb64f21260a432b7c9
z8481bf643f7543b2b77c73d70d3f0de2bc56d0135341d30cc12b7ead2e37aec895fe63ac5d58d2
z3e86beb31f57c92de0bb6d27cb38b322833b0e74db77aef5293df359dfc67d3a50606405bf5ee2
z19ac29056560ab2fd5a715b913ed2b87702ce30bd6d8b0806b217189f0920552c29180bdb48f8f
ze0d0e70eac4c20c72c95bad5432347d966f85f366a848b6fed6540e263ef6a2c64d6d9d721f115
za62f19f45c1596ac82b74ffa92fe55c210faddaa87e75e9d127e862223f1a38a8a94c34637efc0
z9639f478b13fea01c29bdabfafa3a6cdeccd7eae72119d6c4701f73486ebc084e2a712a09865a7
zf15a5bcf9a69bfcd13601f8c720682a52ff12d75359bddceed36484d93ec7fd0ed16bce35c62f4
z4500b8d5e525ff73fdd08e0d76976c399a445fede5bc2d0ab1f3374a313f65a2b75e8e11af83cc
z4f6664866060b9868606254daa72019800f8e028165cce003978d48ccfa17b67b4fdebf3162638
z809c132758faca6d1307cacf766cc8b2d7eefc6107b95c519a0d5ee810b31ca1836e45e93a7e0e
z965e11e345deccdddb58eb31f97706cebc60da48178f2d7f3a277b507e7976d0dc2d6de68b572e
zbfaec01f383e2c50545bcbdc59d505bb08c939f5e1b9f20561f17628275d4445027c766ce6490c
z25e719458d979950f7bbe0f3a9f360beab96ab26e28723a99275f77d2320c6e565c5b8a779aa19
z559349a49b2ae84024794ad1fda79e28e2edbb431c603795966b307b8af23dbdfcd2d414000ea2
z1f969283aa256e0a9703f821e3e5e211b2eaff14016ff438e12aaf13c178423009f02f0e89c430
z0e02fc55d4f01f0918756a9ad14fb8295266dafb2881a7e79488ece20b79f602983dec5493c14d
zd7a0b680ca2bf0a0f028c3013aab4ee6817ae88882ca592c39f06ab0ad74faf0f9d786622a5b5f
z3ca6a9e54b7e0bced6d51bf7336e9383f1d592a52b22622257e72f52cbdc5b60587f150148d4e1
zac43069a4f78462b1dcfbf82d56fe4f6392338fcd37d3c7b1b5f01dc14eb66432f2c58506ab8ce
zbb6fa14bb2abeffff1a7194fcff2ab54eba8e8aba163ef6a69cae2c3db8cc5a887a653c8e9a5e6
z049125bb3d6301a2755503b22463f79855261214a92dcf449a6f7a70a204e82ffa7693c788e199
zbabf72a2ab55c4451dcd8f54699d1804f281767fdb2a365cebac36ae9357afa50e952be0a20e5e
z6117afbf33afb4bfe0d6b2eb7796bba380cbb81e0fcce6fbb34d26cde346b8c950c174c0ecfce3
z610177000a9fbe1ea51f0611b1f3aea24b78ddb36e3037f599a248a40c09d70c4450c75a692cfa
z005fd0d739da8fdbc93372658c62c9d986b9da1fd0ac455bf38dee6c9b4bdfeacda97e1d0894f0
zf80d1281bee2ac1752dd461560dea369152e640a4b9ac806fa2f90126ab63214c886ed5ce3734c
zb2f84ba917929b0889415204c5997b535879e879d341e5fdd7a966960f2037aae1c0da597c70eb
z383efd923f98b4202b133ea3c22f2708afb6958e98ea4723e6972bdec51a645c2b5e1a9b140f43
z44abaf51488e9e9e828e6590d4df8041b4480427eebf8375527e0bd7ed987795dd79c220e1023d
zcba90526ee98cbc96ce65ab375f9f4d2df946a52fd8514fc18f0bd2f04d9d8c6ee35dd5ef237ef
zfc4c39a4c6e00a1272bbc8d4499b1109586b5e5ce9d73e0899f4e74c234ff1bd68dc18d3d3f323
zdd6b3f5d64099e206f09946f9409f5b5f024ea9602525825ab90d951cba06ae2c5f48ac9f54f2d
z8dfb60007ce883680644d283e47995949c2a636b1e162159e4fb49e4d7a5e6317ed5ff5caca8a4
z05eb8a5e5bfce3aa407f2f54839519364dc092e2608d508f6377ea71ab9194f1a89dae5ce02f63
zeef4d415131247739e24d590170d85519337ccebc25be709c72a8f00c889f2b203d1a153ef53ea
z5cc2f44f272db0b58d3a61583920982a248aedddfb1609f0edb9cbfb6a5af25315f5572da48cd5
z1884373a4c12dd7f62fb404f9fd7fd2001974692b2cf7c89d29efbe1cc630ad71de3864795ef1e
zb09b3195222495d0820b769d3cfcdb879e49d68e6a52021375cdd4b05ee2a6f6bca0a0346db2a1
z93dc619b9c9b79ddb48bd980efcf4b12476b0f6ebd9be865f0dea7ddeb63bc5443958d9c7eb093
z028a956e48571b047aa7831a9ef7f71f2a47911c695184d750860248ed9b1f94895e84c5c8f4fb
z93521d47c8571b6b99166a9905c013738e462e2f81825b310814e89eb7dc45e49a853f51df50c2
zc82c3f625565f177c8296a675924c333dadf710d02bd19b5249c38dbec9680859b3e1bf75648c2
zb851372128f5f3af95860471b944cd6d2e0e4cf4012f0ce661086931b7690a5bd5274df3ca8d49
z917996543edd264640153e03b38a2fd28a705ac1bda853a15e7ee5d86c25d06f0aa99cb4751a33
za88c69f8e19ae2758ea2dab24c3c1dba1a53a0a94475f432d4fd34d9ed0098c77b647671f2f424
z5bb8dc47f57539ea03ee72ba5d31a0deeb338b7673056dbfd20b29b62c87216ec9f464d5dc2db9
z34e81202cd841b9a1232d5f4a8d11aba9fa7a2e00b1a52389c3f68ade14cd143250a97ded6806a
zb93a6bde21d4895e49a1ff0e2c074ce7d2e47f64abff6ba29914688b7268d55017bdb81408cfaf
zb64bcaab6d768cbee31d27be44c3435d7aa2884aa71b7e09e09e6282f842069b92ea9e5f544606
zc07ce53f7bacb06295e7b7a8994ecd666c4520ecffa61eea2d146f64a15d4161b6b08e15674e10
z2cd151cbe9c98e7acf4f15a3bb2dc98ba2ee94cffadda2c69048ec5d62984b19b62d345cb59c29
z03ca0d92eea56bbe4e3fa428d8824609e05921eff96fd1ffef19349fe9580064d6035dcc15eb10
z2aa8a43a8673a01dd92662ce5e4921f0589fced4efb57c4d27635d672243e67ddd9ede3b349ff2
z99d2b684d3eba0083b629161ddd450cf3a5aea2876f258f12c1e12cd9549df82ba6b83b5e8015a
zda57e2d92735c8100af6bc55f9056df4d4a74f87ae8d12213eb8eb933bc1d17fe9e5399ac22d5a
zbaede660052693631e22b9026644315b31e6536d701d0f0e31f74780864a9d5a1a8a0887ad566f
zb46e81abecb7dc578dd0d13554cfba08bb9ab677c2ee6891683cae019a3490f853258cc7e1f264
z307ac85fbaef3622bc5acedc0bc744ed39c4fd8cd33f8dfdcd4931461bd454fab8b6fba6375256
z26417bac85f9be1abe812e8599861573e66331f3ea7d6845b6a6655b321b837e4c0025604c70aa
z07a4dce935f20643c92c51de5148732f6133730d07187dbee0966774fc09d7bbe303562a816d0b
z2531c811f5c4689e2a83a487d1e47bc2a371d338c0c634634d61b3461ed382748c298c1c320ba8
zc5a169efa72afd502856588cc4d9f9606458e7fd78aa2eac405da1b40ad1379475af0e2d38c711
z52ed3905214eaa70e30cb2bf98122b5bda38766da713375d1357810f076158020eacf3261cba53
z5e9b76ff7855e62a38ed48407c0bb1e2d77853afcfc756d8381b24a68e86ec6d5430208ea1ebd9
z02bdaf28a6e220a7c225f2c10eb41bd7ee1056f27ad2af08627e9d77b1b3a286fda927f4851f12
z5c75b5647c226399ede876997e60d2f1854377c77dc80fab29d606e3c5f2c18e5af2d27268553e
za8989c0291baeb4bad00016a3cfb496ea5964c4874019f3093bd127c60891c9e5a683f5e40d8eb
z1224132213dfb752c73519d80c4baebfa54244cac439ce646a94cc00ceaff1e146762b22f9ec8d
z7f66f4fddde9bf93556f4873a3bd0e02cba803c06d205d0073f1c0ac297e7848589925f26f9b92
z48e4827def344790edce5a16a73d83000fad693d06fefdffd0f2751458a64bd6e806c34796fc5f
z6d515e023ab7e8e01ec9d955e70c213760a5fad2e199d802aee5af1e80757b969282c18f743c86
zc1f3a3e23f4a625521c1e3aba9795efd25c1970023881a5b40c1b789987d13cfebdd58b51e0bfa
zb43bfa247edf15d78d4230c0b2ad36c415c6dca6bbf390b10c42e92d3da61555b1e24dbd2995c7
z29efdcada39ccff5bf82e8ca90268935eb55468efddd0c807dc91b726bda237843af5a27b1a156
z338d0aeef929bf02746f963783169b2012b80107ee64a373c7fe67487bd2540364bc1ec24a2bb5
z3cb94f062a1406f42c6e3f7861177fba3e518559700ead1b13c8eb815bb6485266b6d1f416c82a
z9eee287b77945939c404ec36d8b6f596e16bd2861de4651e529aa2fd18a26e66e590440f2d288c
z14691cc3e881f5b917ae31e6aa52f4e13e2d2e876b7c9a56f2167e8dde97058ed45b74bd29382a
ze3321f7cc2c8b87ce01757dba4a8a7980b7ecca21c0ab01e9f0634dab04a2591b5b7876c694b73
z35ff2897eb354a2a1073d70390eceac434549098a1f51b2925d86f212cae906021700bd105464a
z910cb56ff621ac38589187474d19dc056ce1d058b34d974683c0433e4af5a4328ef4876a1f63a2
zdfae262a77771521544794d31f8d16120e14a9bee8ffc3ff45f6eee04a2cd4a4a75aa6086d197d
ze05a096b5abe98d4d305a1f930457b4169cd6b7896f85210805ba93a65ab93a7c9a5c61b92f0c0
z13e3ef2c7ec9496f60055a4a7ee76bba5ed9a7f103da500afe01e67776d1755b166d1297528766
z589a8627909158f080c907dd2ad1af92e72748488f0aeaf885ef4ab2b596627ffa61504261fabe
zb750a125531d28fa2864b61ff16fafa2aa40971a9b18f880688e05a83078b40e51499d2dc9c7ae
z2f616168f70ec0c7855e9bbfd9fc3f4313bdf5b26704c809993e69339c9eb3e8bf5b6e0073a4ea
z3204e7dbbed54ac53fdf5c7491b5395dea0d568cb9b6902ef90d326789706b7725e628335ad557
zbc4e44ce2f34c6a510e8817692fa4cac6c58c67e1f9da33da5ec8d46416077aaf913046221874e
zcbb5b13571be18d4447cb4257131063b19df58739f8bad7fcd7878320fac14480d7e113c6f3c18
z3ec757e25719bf90af3f437add8ffe277d765d2d1c8e8ad39a053ce9d1511ea15a036666d08af8
ze88b689644f3486e8ff16ac286e98b10f9e2503e1889fbd4b988c9ef52d55440aca9147f72fd9d
z629e5eff5128c092c0df29afcfc460a2b2d4a8e006a1bcdf5861f723b687d11f7b00d2ee4d5d40
zcf787a8d14b88ec332049613b3abb9e6fd985395dc804f6ac7d8d4a71739acbcfbe829a032037c
z885be20ef646540f4b081a1b63d7a0597dabf58ccab412d9a0ca58a93d9123f32e5c538ecd8956
z2b1a9ad5d8c70a6fa9fc88f78770b528b766a92624855f219273a65c5f35d04fab26847eb3e7b1
z471fae70836b338a8aa6d3fd4e206fd348cfce2085e4c1fd23785dac3ae91fe7467b7212e166a5
zdbb273b2a73db122a4562f3a5a0c5cb9e33c8d266abb573d85f631dcd9411ed44b3c4369a5fb41
z1394d26e3b487aa15f9a55d900c551fb04d26829c2fa08e4a887c8079408062e6afdf33dd3d566
zce8a54a6bcf526d507f3c9e62f3445d7386fcfe47a146e8fc0598f05a0f7615244a5d5440b8940
z56abcfaab275554f8a161eca70819350a13b26a9ed58e1b41c2bfd3cf4e090da33f61a935e267d
z28840c346cafedd42458e1b958e66b18049227e0ada706215ac3ebcdb4af7ecb7d91369164fa3b
z260f5921f02aabf387024b61b822c0251eb4f891c8f3d37f2b192dfaf2841e75843d63caf8e253
za1f4f94c74e33b17bc60c69c847ac90c06fe61d18c36c9ad7281b8810450d0392243f10b580295
zcd442bcea68532c91b117391229cb66ed6a266bf7399335431951177e8ebe13012934b4fc0598d
z9c5cfd40ab0d3f5ae39ea4b521062d631179f200f068dd0ca330e8184b7c69b93d590782dd528f
z1ca8bfebb0e3bd395deceae0273502450528c8bab9643851b7146b35b7de7eb2cb176be036bdd1
z06b527c937e3c0a3c83e786cac95d1906d6f023962be9da8538872cfeee6aa62d51d1ee2b6951d
zdcc6cfe25a53c3a175dc777a72b315b802203499b1e8d686386e1e0942ce049f21a2e6e099a67a
z3c8830da315a941d9a038708aa0e50e163c2629d284e3f1b31b9b84c2fe7d642443ce0a7a1ee07
zf84f29d7f3e08f52180695a8a95ef6d3e527eb006fa0f7e20af1f397a8efc45737e318f767ed60
z7caf1f9f64bd6a86cfa8b30ad1d864013c39cbd4384e90e11c55bce97d6966b32ee014276ddafa
z0059f737688adfa2bf1184ce1353227e42b39c931e082a53ff8b10cf97c7676464e458818cd352
z9692ba4f43e88f5e9770af138ac104fec2798dc83a22a07fb6dd8bbf6aef8359effbb90c89f21f
zc0db913e2936ae2ce33690458d54b2ad5c664ff39d00adf7ed995652ded84a6404ca8314612d91
zf594c85562d1f8b7a4e89cc7ae647a8ddcaaae243346b2786bd4181045b5e4991e696152f058f1
zab97ef944e51271d6b6ff2277683b97330f6dc38a8700f5df74517bd43bfe2da0bf75d4b6df3b3
z7e6d341cff60e3b440165edcb54ee8ad8f1095e1a5865d010eddee7d9eaa2e0c746db18bcab507
z411344ee780041a02763fbef78d17789d892a13b715b1feea738ae531048746f34cc31155d7d4f
z6592bb3cba99ecba09f5590b4fb7eeda07932d82ba3de427a9dc81d159f96c31d471cda74a7527
z7d2bdac34703b38631522433b04d148be76d4c5390258a34798c47bed50efc2895c7c37a364309
z96589736c35778a0d88d4d3b2b6bbf1031794d03d94e7eac227ee7f1c2d125da3214a42c27f6ac
zf3fd6cc723d2f65cbb8abafac104bd140c4fadfed1cc1e8bf13363a7e5c93354d1acc32834a962
z6709d3c475f12f9250fd1744d5894ee4036d0e0e283253defe49b1b273ff77c056d5a41f9ac8bd
z6c901b86bc1fd7db347274c6b8637176ab26cd0b1e41339a712d3cb3a173139fd1f46f3dd8164b
z08f3bd6a2a952dbaee927d516f5f55e1415d2c5ff2e36524df7859bb24b548d144264929d1e0a1
zffe90455cfdb4045d4a4075ce108ca4c04e3155120308b9ba4d72d3fe1f2c94251f8a0a77e2527
z19a2c76baa38e412b837234e4887b6bbf5dc8e6bb4c0a97ee3c73e2ac367947807be768543bede
zeb5194b393f29ddfe9f2fcdee9ebe936dc3dcd96a6edbfdb9b5c2282b117797a5ccc31ee78dc71
z1f0715ce45e2e582c08a0bf0b7f637ba6cb23dd72dbda35eb334661511e22ed7245b6fb60f694d
zd6fdcff85d94eb36832c03444e09aeb9b13cbd2bc3f75249e93053b859464246e16401d8decc76
za6eaab481e0ae4b44fd6c9d1882515d2feaa84d97ab7a94eb7f0ba5df37f997a7bd433b38fc587
z0ee2d3f0635ef69ade4351ce3ba1a972795dadd0a8b6c6325d8551a385b8f64bd88066e9789775
z91a4585c4b06afddeb2164c2d748f6f9fb04f72554f4ec291b86f2d533f400ec930524ea8ebb38
z33fe221ee4f381226a5d126a9ae515c0870293d76e9fefbf07065ce44de172bc4d349457779867
z95bff0aea4dcb6bd720140e748e5a47a603d4eb184eabd468ec8d3ecdfaef470e656093acc706c
z4ded9436cc89352b8a92c975fa3f2830201ac355b55bc7283a644839ed1b5f6172e76c5be14204
z85af1f77a948eaa6a491275b947ed4009ef135f6b05408de00934e8c173623abe964aee5946433
z07a9bb6d7e1b7b2a0b1e46251c7afe9eadee426586960cb81659b2af8dbfb49a2a9a61a86f9e17
ze90bf2d3fc2580623e9b53445a15cc801ed1913506375dd0b460072cba42b9999034b5e6a91f4a
zd1ec3aa3fbec035390f2a7d7756a5c30b67e2676afcb11b5e8ae155219dc19fc7a4b946fbfe477
z5102b8e8d86b5638956b050cdc895ad92948247605ec95d76d09deb5e4787db9a045622581e20a
ze89e012052a0cb3323b938725c0e181020b4828fc8bf29ea0abc068bcd7d9d98d3ab25469b03a1
z89664e0d1f6d1e9b7268fe9649031141c137902df7a2d9d7c5a85a4477fd5d9a0369c5abad2d5d
z3efb70bf86733c5c808cc5ea771c27e05d4a0f1a57fc2824af273aee30df00add47acaded0ee35
z5707e44b161966c2eab678316af95022dfe66e14a8ba9730f81510636c1be8cf458ecf899ecd67
zed6a52af0380b19cd24a36763b751f34408639836a4f1418ac263e06fb29de43afc5a1dc4de8ea
z871d43bc996b44db5ba2f151cd0ad0a422968dbab1286ad5ed586f682b5d8c880d90193d5a9b30
z7dbc9f73c5da3c45cbdd80b28b3b8c824e54396d3d4d1c0d26cdca14d587dd40dd21ee0d1564aa
z87d5c82f4feccf8a45ce3a073bbcbf3ed159d5009927b168749759d74ecadca8a37d4c0f9bb560
z26f5332943036e440f58cf2e4b9109e6d1003367bf289173a2c8ea080a1d91c87370271780d5d3
z820b55ccfdeeef001f1cabea02177201f0ced632ef118e7f9a6f39b54033ac07d47657bd909f72
ze3f3d48e23d8137c22ff022e0aa9c28d68b5a84555c72bd6018e313ce3ed913fced251a2eaf97c
z0d50aec1419d4ea9c3735940cfc2a9511ee7bbd67a3f7d1ae85ef95131a1be309e6c5c25ed520c
z1da2652e213b19d2cbebe1262b713d5cf7d222a3af756657318b1d5e6f0b44d49a23ce6488b76c
ze6d68c07ee8679ee509d0e2158da5d360702e69d6cb3fd56ddd7de71410e8d2a276cd538933fc4
za822260ccef4dbd85257723392630b1f83a6745608316670c81177eb2f75369b94dd9f7b524c9d
zda31ac74b85e0a65d8a9b795d94dc255e05824c30e536a922769a918e6028da9fc4718e7e111bc
zd3065fbdd7062dca9ae88e3be33d32f65575aacc9365208e6ca3cfab24b8dc3238353442bffa1f
z32a5ae4597db2f5393078d98e559daffbafd011fea64616b80caebd34af45db4a95d1c8f8dd0c3
z234028b6c5b76677d6cc121c054377033f261dd033f927aa079b58aef989dd387036d19e0b6607
zf60586f4d5aaeca959dc9feddd17396db8ee402be80e6fb4656c99acf2e5f683045f64263b1533
z9c3db9161a0b9f263905c527a1e4686b3a8223e68e42d2c9b1d635fdb884f8f35e16e1359eda73
zb306294bcdd051d3b7e0729bf45cf24533971c689638cd79d25f333d83531287176371c7c75ad9
z9043f946e64aefb303de687c54b781671b5adeb5531d85a8ba3977e5cab4f852810091a974ef70
zf2cfdbcaa6a5d39dacfb03fd4a9c0a371d0d606a4e13c1f2b611c0841dc524636582a8a91e1f06
zbb7bbfef4925437787e8bd011b2e4264e60a46d92bb0f8e10ee2fb370dab37329cf3e77a4f9c76
z7797f59f8626d858a7a746dec53508d1e635367b3409bdb4072ae9c651ec9ffcc47ccd99d97183
z123c40a02ee24fe4a379cb4c55e4ea92b6640c132d06fc06f7e8c7076c7ad7b1c2425820aa1a2c
z1a1599be9176e4fca8ce92f4d259f83b32bd363fb17fb495a99723d1de365cd7806716b6a431c1
zd1eb04e25417bf13ab9d2660a885d522aa5f6c055b5f0e63084f5599fa2e846b4cb17001a79308
z94336c37c3f09353d4d05889d6594b67d00937df87700f819f6f63b2c024d88704f8c0d55ff2b8
z4615e70aca175954fb68209dd28747d094f65b22a01225e6597b1de998c727a6fee6e8ad7c9197
z9f1af31dbb4744a060110df409b1da5e5dc6c08460bf21e9dc0d024d88e818d82f3eb27832d798
zd349c20ab43731d1da43a29cfe1a21064c53a40a3c646fa344b4e2768021f4f1252aadfacd1f08
zf1733811604734663df299d9445befc9261321d8435081eaee6accb9d78efad71542beab1f3dfe
za2ceaae85241a35ae9c21254b988b5d9913d0291194fe61c2aa670b9087c12c03f6cf7bb53ad2d
z45e907509bacf68b9c302e1db94a492efab6f28e28253686a6022ad351e6d503062b6111dbbc04
z54d7d221059bf99a8a2652e688bf39e178166ee0bf30b40b326d11c3507148b3d595033ec1c0bc
z7eb69b786f5bf5d68371d902b9e0123f3d21334bb737e6cf9b403ae00c314288e18de40ec4714a
z23b8da95ebc8fa7b2c55a2a74190f0398a45a2a1a9ac7b41d4e9ed949a6225531a08664139df8b
zdf0d7fc8a177295d9fe8267e146b568d5b94038e2ab172e147b44031f5397fc77a9eac7dd763ca
z7bd38382e053a2f6310ed544a5f74042dbc1b9b3c70ac849010f2b5899fc0bcae7ef4cd5110c52
z98bd5cbc143e16177ed7a9e2ab178b26bef053d934b37004c44dd735bd9dfc62985aef4a331e1f
z9276074bc7480ed18eaa2e100171afeb306540cf3610552a01e5aece82c3664c807638f72ce6f8
z3a98cace53781e71ec691e8b1f03373ac60a281001c406f0607c32ea983e509dec3a04d06d74d2
z976abab37ea599bfba6749fcacfede538500d9a4a0bb598478a17179684d31ef77ae66fab1df60
z95860c4cb7777009b1cceee14acf22291432609ba4ef5050a550cb44d61f7a7144de74a4b500e6
z886fc56e1c0082914a962adc40c8a7ee0aad06f57681906ed2f3c752ec6fef6ccf892322f9f103
z816d3390ac88c5c3d4522ab5c8c09b802392a07336358fbfbffda95a6500cbc63ab777cf63deaf
z65643f62cf167b80cdb88426030fc4e53280fe576cd45e3d51e538152e2b997d8d7f42ff6b8f5d
zdc5802750cc29a27659fd985f99d22a0442aabdafa0030e580a3e4a018d88fd3f3081de7794cd2
ze6a2f32b8df7d94d6cb1696ac9bc39a22eb5d773961de8178e1bb1f92915792c3fff1a997a2f10
zf59254aa5b2e271dffceb47f6100553fd2fd3bf77b651530a0c692eec41cc50da87149ca87f8f1
zec59075dc47235b8c1b4a67d1437ed11e508273421a36adb303da298da58dc2b9e0feadcdcdad9
z6c3243199de56cee85651712263279d52f3b87811cc747f667df11fbebbc949cab396af98fe9fb
z74f0fb329a81de7f455f09d808903dea3ccf9039e19c6a791cbb7c76e427c7976036ef7709740a
z74416d2f9be631d452ed10d6cd3e78927883c823efd8b4700e659f32a203e1b47aaf06ce2b5a5a
z9d75894f40fd19b4839737f67421dd64f91aff2d13a5a0caed73d6a55a6a92091290fbe021c1d7
zd96b31002959374f81a078cae9d672dc6771d6546d10ad65e3821c5589b3ae0739e4325f782228
za1f2a6712bdb547d2833a6110598a3a17581c9ceee3c92134c5d0c4d87a2c1ff667afcfc05a7e4
ze55a2640d9f89b7d81827d210cec78f88edabc3adb132c7586bdfbd774b267b90f30b822bc3f1a
z048f5d36d2bc85712e30e91fe6e6462b344b0c23f16a43ffc4557520fc64a1fac900c8ca23f287
z3626425823093c0c1ae6dda2d607c534c2ef61deed97795b471971c0eba8a891db31c0c6ef64ba
z6014c68961cb6dda7cca46eeca3aec284a95f5efb76d2544ad5165da1d9367589c5baa953e8083
z5c97ba87ba4e422ddc20cae2807396b8fe46449fa98f984083e358efd6dda61d5adfac9d497f67
z180e966b43fcf7229f9120f43064891baa4b3caa9e424494b6ce5c91e1ba8c596e4cd31a25ff14
z54732831385317d8028c8a2a7d1a95655a712073a002739f36664378bd88c682a553dcc9f403c4
z39e44a70af6e35fe941eb688ac0ba5fddbe4cbc63a5a7a35dac7cd5a2c78792a9d11db962d88ce
z1d9b72d65679e7306fbf46f746d51d5a3ee68f4059e3fa9e122f87eb01fd264bec06317e124d15
z84f26fef1cd4d1a921d4d3065168974809011f4b692c3eb5cb3a702166e37d56380d74826ca073
z2e01bd072113a6d7068cbf0dcd381dfdd38f09263648fee987a01cd401aac94994853833e585c6
z6dc02ff54a1d49438b75657844525156e367d29415cacd52b321641cb528a81d304da2bd38a153
z342b2c76ed7565cb9c80cfee002908914c17dda376c54c582e2bc8348092bbb04815f206507f77
z3468ea5655cea1a4421b94d67e0986e40118f3892859da88b5f0da73198787051b035a0ee91e3b
z4d5950656f4f99f9ab93b3f1d6793acd6c74f8b6291d9e89f98131711cdd6162b0e4c44107f229
ze5dfdddc9f1b6cbe2c5bc54c381267fb6bed68973ba0dc78c86347a5d467862fb8a82849007b5e
z528229bc1ae2525c19385bb7201c4d896d25b97c7e2baf554a6f38771cd4c4a23fe3a181a22a49
zb1791c86399b01190b9d9408d9419a303698a9c948ec66acbc306718ed5c288ba66f92088427c6
zd972fcb9cc86bcc6ccf937a675e87adc81b30f8c5db78e4d833fdd8b3218461c0bac2a53dc1b87
ze97039d79beff40875467b9b62534de7cb1e49b6c909ae6db2f2c2937f1580936d23b4cdc72af4
zb3b92a28f445fc6535576d56059152371fb5197a95a26c22821db0fb49fde0006653a83414c35f
z3adc11d6fdb25ccf7ab901708f4d1813f4f1e87cf6c70c660ea59969377fcd2bd88bbd61954545
z22a4f42b14536b28ca1ba296acab932c3a4ab9df1216d4f91bd56dfe55428445bc710ca70f71c1
za8bbe351d709142815bcc059eaef23cc631b98cc0e31b2533310bee0e1ee73692edb4723fe81de
z4fe36681e432f8bf4d85e31edcd8b3fd1b6b742b074ac3de85564d4ca7304732144c8adb4d3531
z73afcaf79de40defe0b73b1ba010f8a2c731b87a9264f2c50adbecf6ca2ed153b35cd36262d1df
z0ca00132b32f23b6972d9a31679b1dd8c0d4974b7a9d15c3dca5894d91b283ce71ad507e728db0
zab443c2e54fbccf70bb1a28eb16b4a51014efb0fe12c7702ecf23f75782a233fe20443937cb977
z48c5224720f180a2680fb25951e057d2ce52f46ae1f4480705d167ce09f6901638dea3d41e4199
ze2737ef149d67f8d4d5779d8e9e4f18261e31e7f171eedf55bc1079d9ed24b1dda1929a3a81586
z115db69a74aff192900fc0380aa139c0ed0c6f5ee09f4f90075571519cef0185f7a53711953c80
zc325b8fa6d711d84118160ff67af3f7060f0517c94ddec7c9bb16f22804915cf31d332075e8d42
ze7d947d9a49bf77084eb30473a121933dbcc3a02f0ab0b6a99a6868861f15ed19c8d0049621d1a
z409b8d8b24ec7f10cd99eb20dfbd0eb58c16bdd3b2fc1e20f446c167727976bb590a343cbe9a88
zc6d89bb409270d5f66326c46d86024cd190342e821a77cc9a8c4eda94334175ea75c1461d76ca1
z8e8777d2ea6e951e40ba33c5b15c5f3b83c6987e74d9a0764aa7039270e395aa483c16f673ceb1
z99a9ba5c1d40624fb3f94c4ba17aad795f8c21d33cf539d17304f697f19cec0ea125747ee93108
ze8c915d46a8a58732e7ac49fff40e49c079a3b7ec384060f33f805f22b369cc12fb257b66a2348
zbd72b431f262f2ec964ab66472ed349892ec19dbbb64b356c2a1829e4fe9cdaf6e04b89298774c
z7258635ae94565fe12c42f4085962e81281f856cb3adab9406039a69de2654eb48921a0142eaf3
ze0e6a70ad06cdbcfd540633d9c852df29ea6c47290a49513b66cde112aaa63966489463917a1aa
ze023e23c7197c18bf48e031ad6ca50b30f28b8889ce8bfe84a15930bb97bbfa4b2c30532a4c6d8
z4038ba4dd62ad7bd2ce1384d29cb43a30bc52bdf88f901a0fcbb0d1d16d3f9437650d9994d88b7
zf2a917c41117a8e0d0b00bf845c2271c94141c68def6fbe38284192156bbae49521fa27602d8e2
zbd3accb8cb10986fad7d9d68b8516adb08eff4c93683b45a6571c4bc71de795d085771c527218d
zceacdb0900b96139f402ee538a6137218af34732f822c063c63cf5e0b3eca794581978f8976224
z2ed7c9a6ec051d9b5dfde2d77386b21e98e32f0aacea033b0500a2ad2696b1a846ac973606416b
z42f5a7ec47ee832f2ca7cbf1665f81cbc220a54c6af00f4df7c75093cd7557498e3b91395ce188
zd154d9d81759cbe4279eb0b7923d84fb68a1f0a57b1f35fb3ab832595f5c8319e2c42a856ade2e
z7294723601a269d014ae231e89e5c264a3084427f1ad59c7aeb21d3741406cb6480a8095f4840b
zd31b2fa5b8bcfad3ce527f55ef37d5167fc4b5437c02157aff3274080f09e62f9a77ca48289954
z6719a30f9a0686135b71abc8c1c1b3f74950ad5f02b96142359ebd9f5ee70774261159b7632204
z017c42e7119db02d1f88e9598a4b1af077dfb5c1465273c4d85da4bf07af2fc100dd7a97bab31d
z02175e29585bfe0dd2b1ea138721380f1e93058e245432c7bd3445b60884e878bba3dadec637ec
z699b4663de0d97620a42207ff171155504437d882383d94862a7e23f8e3ae5595e1ac36f3acd4f
zd1e5507ebcc10f8b5a082e4727d64f1257a9a78b8f387a0b92b39cf242bed37e75e7595a0823d9
z6ec59ebc44b1d0ce324b204356ec4fd51c7e3474e4fe2e062879a6e8c1a84259d6355ba6560afc
z14da270584753a4041a8aee197e4d2623a2116cf0dec5c96306369b72a341968b2040ac1530e07
ze7444908bb722536b646d93c23262fda845de1fc503121a53e8fda759c7a7fb0b5dc4e865ccb5d
zeaaf872ffc32229b42ca005b989fbb77b34454ffed0c05d0587a78681018bdc84520e55546d615
zb3a489642fc51cdc30207ff1c035772200ede814cc81407ba2a38dd6445fb9024c0cb4b670951f
z58fca07f2ff245d03096fdb83466db9e32dc31cb3568fd5cec51eebae05053ad8314445d30f964
zd7d373c0bc543f37ecb96b7c198ce6207ddcc85c2e2bda9d69d6cf40b42c3d3a4639abb342cb27
z2468fca05730b4233ca85babdda90f67f6139a85956172f8674d9d482314e61fc152efa4666d8b
z91396a87be5a5cff66e5b0d863915dbf7057283976e1f0e21a210a102caa1df9afe732623012ea
z8f8f4b8ffdaae01735a53da074186cc21075710408d28fa77a8688ba667e58f25d7d58833a50a2
z7a043f62ccf3a08ae6d946a76b5c9fe2db5bacc64a9efaaba0fe31792d388b7428b78a7442e028
z2af2e57b73453aab46f717908faa304fb515bf3ba6b15a5d23da795bd3287af4841650b6111b88
zd8556781cc033ba46ac8cde5124d2fcded9aa2833a34948f2a959df557e2a609cce7e2a8f9b1aa
z5f46feda0fff06b9ce98530967736c8f3037a2f01303792f3bd3b1da5dda8cbf7c5f1c2d4f0c98
zed3d0a3aff4d4a1c5a30171ed63139976d4dd91c78fb69ee5ebf2172af0cdc8cfb4c3d265144a1
z316b9d2f20c07779b802950e660bb48263c90315c8ee23f948513614807cc5ed4e37361795ca50
zee5ab5b349570d6d05b2797b83c7de1f2aff8ca9ed16e786863520bb7815c70ceb7cddad83dbcb
z8de7d1e0bb2e07c78525f647f2194f6950ffcd8ea28425b8eeaf41136d3da1555f9b69bee37869
z570e30bea0b5748dfd13120795c1a22619a901bad9dc29c8f36ce0443ac51af0bbdf0b410b8a77
z1ab8e5149e53db100df19edfdad2d2d2c5f897f929f544e077a678c1addb0406517a37b7a8654c
z6ae5ab6c1a434f1babb05c15552c433111652f705fa58fd7c0f87f11597c95e88bb07c19cb9a1e
z2d17975b4b906b4d8df114be67d077f9c35f438385df40202367d65b7b4a807fab729aa6f61104
z0e15e38760712f2d8acbb333df777a8913228f8e52a6d5dd28dedffa60f979e4d1711377125203
z906e1d28db94ac099b969f30e39cba1a90a1edf321f1e0a20ad6695f046f203c51a3d23a0229a7
zb3445e94065ef23f7b52f2c87a0a05a398a517b0fd96f8080efdee4aec0de41402f3e7253d3166
zd0c08c96cbf1e7abcc7625007ef11a5e6ad41ed27526463b22f3865e486aaeca59e675003f405a
z1077023b8c2a9fee3a06578e345c2259cb24d9517c1a4e1b4ccfd40d19b5ce07edae675d27d70c
z649c7ef14c92f2adadcfa27301ff3ad836428e030e41b3968fdba8a57d87f75b9230a53e14dfd0
z9b7ed0f633c1a7a656a37dc1ef5716d59d25047af52d2eb58cc2678e4e9646256b1da5b9be6572
z42dd59ca822e3ad8c201d4e7d135360b5ef71f3d70411515448bc23e21ae19291070bc90087729
z25df5a9c4f6efec62ed66525f11728b0195f14c6be5644872ea616bb1b961b471610cd36501f63
z227b28a3dfb4f82238c1dd5799377629888bf4bf65485968960f6a79019c6490865942a87313a2
z8aad04d927b19949e4c0e78265f7f43a3860a036c5f569c75cf6498de2c2aa1ead97a5266bc784
za3ee0536f60f02eca3247626389de7f9121063c060d45deb4235bb8b41bd90f4f4f93070a847f5
zc45e7c1b654bc32356d88df669aafed806885af57cfb90ea53b066bdff196ea060afbeb51adaf6
z5f8e3861c7494d161b1d8672f77b5289347942c9e045f910be62e49c06d0e1707052e1e26703b9
zc1a6ad224d4170b52786e780de4b5731e671b83afdfbf3569cfb3d9aadc06a698772e657b6d523
zd65eb44234bbea5bb316093e33491132dbdf3748905b8ae7e9da4a6f20712f1e65c4166d515a62
z8b82e3474c2c4e1e1ec34ff0dd60db8bc969d1b724686f3ac659602b5020dd53ce1b750e59bc34
z06365ee3c41404181404acd0c290cb72bb5124fa4870c7f448b6d23e3c3ac8a32670d355a50c53
zbf0b94f4c23d5e9cd36852b43c7e302bcacdd5a460ec6ba0d57cfd479b069e4dddbb8adbd80a97
z1ad91e392728f98b049052a653129a417ff8f65bf6709a42065ff39dfedda6dc32a92a5164c7f0
zea28286ff8dd83283cf1873cf1b159d21d1d85e05bf7bce9c649d59e340f1ff0c04e384f215c0c
zb3f14fc45ea8ab46f16dbdf3bff32e429bd21b273f9c62985b52253ba48ddd9a33ab998b340dd8
z479cbe07b651c025d638baaa543a0f19c40921354fe44c30cbe45efa52889f39c5fa4c779ca1e1
zf9d2ad53bcf5cf8cfdb682c419fa919ebc0020e9a48f1a082c31834f703d837f14f73dbde325f5
zfb0c0e57351b756792bf7c3e6714649a5bdddb4f5666af86e3494380623f619dcf08fefb333dba
z0eb1214638887e19e6dca02e9cc9ceca1c54c9eb1f96e923a0e02a5b04d7bc9f13d8fe5b0ffdcf
z8c027b6154408542ff1c1570b3316a965d1614ad6d231ac240f6e6516c7b1ceb616bb7594f1843
z466adeb2d0ce8e2ee5a5c11c7c642905bf733d254913b5828259ea46e09b4c841a0281e5f1c92e
zf289d0817e7fb7eb7a17eea545bed15e011f365740d0647b2918e0bf0adac08c74d3ab2ef6cba8
zf0e1219610d9ff4843cd8bde6d89fcf74b23f28cf44776352a187789eaf65d4a63ba48f126c260
z1c7c3ba3849ed8635c8bcb675b1bdf10307befdb88763354bdf3a81be107ec8487008fcd6b2ab9
z9d92744af95177075357c3a77cb6efb60559afea9a4e4e1b92e78d50bedae01ed050b10781c88e
z0f997965caa2b3b5d4c526ec29ed24b916073ef917e01fd91b07030170cb7725d9ede3e494f0ea
z9db23c1d98802f71d3cba9ebfebdcdf69e48c3ddb2173c88088cedc54f4cb5703982bafe2a84b9
z125fceb944d1ed08a6b0b6fbbad74f2ad4b30a9c8791b41e9353c98e649a25e381c48d8a0bb379
zb06fef65e30b6e466582ee2dbf4106a6ef4958794e8c88c03a4bec047edfe8a01c04d2420dd087
zb627af218ae792327a288be922cde4fcf27539606eca3c6f2c8506a6b5582edc2ba4d026370516
z58225f23fa7f013a58c8c4057019be40710b35642a0b896b38a667c775256a7ea1896ee103d5b9
z84777e884feb09d9fb3ee60098148c9ce1810fadd4bb877e2ae9a7786dc8f85faec57fef196824
za8c4e794532f996f4dd6c359f355a131966582d3d07ef7f2ab973ee83b4c1a94c194949a442778
z14ca16cebcc2e9ab50d191d813b4b51981f06eab9286b9906ef7891581d60117d0eee5d5f41edf
z6bbdc9e36a84e802f5d839fc840baca97ad9754f1a41329b7b83b9cafda79be5ec32f4c14bb0b4
z93f29e9dd67f395e88d6a302ce3c777507d48053ad733028885f85369116d4e0f156a45fa73687
zfe12b04abad9aec9c21b64347f7bda2f59fe611f4d414577b5b33c8455f90ee89ea68f6ab9430a
z3e9501d4b603304f429f2583dadfc1b2256c48b2c72e14efad18df3bb940444b2f4d55d094a8b3
zc7bb739d6f32493ab659067296a014b3d347dbd462c48dcd94e6445a2aa16894aded3d0101409d
z166174deb0baf9aba4b762eafb311384caa387eec105644be2d50da0d90b84e27aa776b3ffe1f6
za1f49c46dd32345b028b5f068acf66bf6387db945080833ce3718ec26f7aff20eccc2dd556a1c5
zee1e42eccceb0e41a21f5d256484fedbc306ef9a84b086321e6550a8d19c30791d93a5e515ea60
z15530f673850ee1d18ace54af773a3823f1093fd9a9b6238a2279f953cc4536498276ede67c836
z8942b41318ec92f19148874dd44a0fe8e543985c35cd7d5a82d1bf97d1fc4df449fba2bd015310
z180363fcf5201c969bd60264449266eb71933913fb7c3a53bc9d62a43e9542ccd8c3d368d37af1
z5ca219fd8718f5d7c22d71832e6b2cae561a04eb4bfe146eae8cd73bba8e104f98ad8e2710660b
z21b458328c44b928d94c1a3def2d9238f5181d280845a0503620b5eeaa720de7504f2028230cd9
z007f40a55962510816076456da7eb6911062d7dda667663de0f5a91d7df6b3489841245dbb40e2
z63ddbf024a5ed38006ba7643a8bf80b4bc6d0450df7e6ce2b627e10ef67c48cb695651529e5958
zdf6181107554f20aeb1898fe9da5bc723854937470c457978e179d35bc023379a6ead3f3591088
zfa1fccfdbc9e48f5573cd88a6236b338e5fbfcca96a1aa2495863a0f5adcf6079a4ae32901b642
z67e98744192fda744dac2b7d4acb42cc796019084959c5f58fb043836db6f6a5509b6da3df7377
zb44ee81e5db5a230f862efa89bf5a7afa2edaa8fd75f0ee70843a9936c0efee1a81f5067c1f433
zea38c2987e27bb78696d86d857bc8ea7eed480c11d50b2dffe433cbeb65d9e4bdbddac1f97424d
z1d909fce08cce7d02d80ea580650aa06f1ade608076a746e0b9368a191fd6548c325fc408a2f06
z649124867f08c9ef9cd82b8b09af383ab736aee4d4111a006afdda245362200bc50195f7458dd1
z53d77cb07c0be34cc7f830e1ffd3273179773dea17084fb69721b062ce15395a1e571fbf04c750
zb77213bd1304fe634b3d1a41f3d44ac907468595cb749343133a1f1422020bb35d8d8a308b4e78
ze927e820c5540590c66bd5f072b1b33218430f8a50431f79853c9f158503f3e3c910b946836507
z7899a1c23cd5812edf3da62d4ff67e4989df72dd44c32ba65d106fcfdd9c2772613d97a361e8a5
zfcf41fd7142eb87e797a11902bce3cac6653a094e98455801e04a033b31b189c821e3ea7696fc4
z1e468afc189dd6a31d02775ca7d2bcf326eee28966c678e32e4cc5c9c4436f8315c3d59e62fad2
z2f4124717bae7faa8a2d4b9d317b9b3a0d01f47b7e45574ebcc38ec9f9811eff1fe2df98742c1e
z7ed383264dab3a98aa5a913b22672dd77e5698086b0337a56cb5ee7c2c75d6d46a9e73c43fc307
z09426096d55a79a8b4c22ad52b33152f64883cb41f161ff0b7057216638140fa0747099e16a10c
zcce5e384f1a9b68fa592f69e862c366a8c180564debe97160500d9353ca2a246f39993e1cb7264
z1adb792b5763080443ed1577767b9bd87b344dbb35bd45e4c9d5ba26d1d6aaa8bd7868e464254e
zb73f5a4c9c438477e841b6514c00fc04bca7491cbe19e30c8ad895c82acb1dabf6b3777fe2b878
zf9f094ea6ef21a41f598431648786fd1396b6c38db20c8cac6bab7a7575f3011ab216c9b0b72b1
z12c94d370aa409c89f50cee3e8c46afca5da773b804e969d47338d98eab7df3e7681aa6f50f7dd
z9d90d9581d183c0dbf44720c645adffe95337a52
`end_protected_0in
`else
`ifdef MODEL_TECH
`include "qvl_ahb_master_logic.mti.svp"
`endif // MODEL_TECH
`endif // encrypted_0in
