library verilog;
use verilog.vl_types.all;
entity tb_multiplier is
end tb_multiplier;
