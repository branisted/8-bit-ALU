`ifdef encrypted_0in
`protected_0in
ze74c34e226135848fe16db9ffd31815111b6d7fb642c521a3f628cf6da949865580b22efd062a7
ze90adae0e65e66a2c36a587d0a790699161455169ed55a01f2084f11770a774ec4c588039b380f
z6de9c5084882a40b79a175f5c2114b2b6d78b070cb806e1c0aa9258297f4687ab308bc470f0040
zb0b1de382961eeeaf2e279e1462520fc31c119af8f2b214846f56c2b3cd2eadbe4099496abff18
z15cec83ec4a77b868344aa20ba7360908f5c0de2a79abf8b3534b883bb12180f68b5d4beb444cf
z3fba8f13afb0abfe8fcc4294810f75afe452434d2d0f1166236c82f76edf1e12979f04bc35693e
z32ae028996dd85737a8f5adc1ebb94f39c940246e887647b64782cd7ab429b0544c173176cede7
z01dfb26b1f73408344a52b7e1f117f12bb9c8077b34876c2e6fdc085981637012dc9754765e1a9
zc512ce062e0b8fb16a214591f5c81e1353b900a611fe1f4886b57940b41b7f2ce99a7b84b04b90
z916f717e73bd10589c81e207ed77ec660a8cbed5b487fa50acde1b055c8870bd8676023f21ddcf
z9c98cc47cfa2d654ff1365d1f45035a045a66c5dfa827905026201628cee5aae21fb892db766c4
zb5b1406e11aebfd6dfacc9da5ec03b70c276807a3eb15e28ec7ab1dddec42388b9424ea285623a
z248195c9f894b36317ca6e59c86f11031163f5f5bfdba36b10b435d3cff56a90d9a15f1244c71c
z9a4cc6c4a91a43573938f48e276eb68a35116c6f2a5641cfccf667f074f36c3d65ab81e0e96800
z60ab106795c065140465a1ec216ad1eeb32cc32159964d3f9c49e0642ee676d7e60343979f26ce
z92c77b9b0ff0e99a07efb0f2f9376cb9c0049a695e104845ffd4a5b6b459c3e256168a74d8ff2e
zd7845dc66131c3874fe76c65a208eb9b003a1a0475d4906c7d2a39d1eed852b974267d4012bae4
za2b0842c00695dabf7681e458cddd4cc489583011a454e9d923e21f38502c7b28892e5817c5e0c
zc408538c5067e2a54c8f698308634752adb675ffc692f71bba8719b0c7135e9e3cf27217b52d04
zc6cf6abcf2d977ac40d1ff981dc8534e3f3513366d6328038df8ff0effbbcf9bd5c7adb10b9bff
za427f22effc874b200498576c0c17e97db17459602a89695507c527b087f9608a82b8855cbf3f9
z6bca95919005741959d6d489f2d7afb9346a1f1563c7112170ad382c658b7ff0ceb2b9b3077f56
zcfd8c5131db99a69b9952383f312bf178c975e8db8e6f021de3ddc11a7e86922a6577092cfe8cf
zb58ec5a55b61430f36b327f788743cc75d0d55cef672d8cc910899bc25cc13dde850e222c1f2b6
zd0d1cf8e45e58ea74a3e6bf9e18fa0287ad16eaeb76e146af24f6a22a671ba71ce85a50ad024a5
z97210bc2cf39bd4a1e7f1c410dbcdb92c73b005a4d396c751a17f61e9230b917395e929d75c893
z745d944b7f1ef16a86396789bda901eba5a232d550ad7e24f9af02f035f3d1a95b555a78f94b6a
z771b76be9614f3fd78514f1f13013b261918ebfb8bd8fb4a3d5aeeeb3b5cbe1d10c1c00f5e219c
z4d0486935406f1c99bbf096500cb3b68061a324b2c18284650d7bb501a898a1d0d4a7a2e41abd5
z4a70812765adf155e8e32ef80ee53cbab3bc6a7c0f00580da1ee2cca803b65c7965e5b229c55b5
zd29ec108ae44a8e3c9d44e29b2e8dbc3dd88b0a9cdf3ecdc86847e9a0aeb0760a31d2293d9279e
z2035bf950db756834a216c701ab0052b6aa9d29e4cc5ba07a4c3f0efbcf2d4092111faa9c24419
z67a3bd581f036ebcd53fef938a8a30163661c107735a08daaa8c33f65f366f1cb2e2fc670a4b98
z0024ae33a624c60916831c71b6f55c04bcd02a0128d46f56cce1aba380530d4e9e27f635c26916
z57dcff731e382aa591f19bb620b86c2b531052d74865a3b97b21dfb6917c3d8462fe25888dfd34
z7e4f28b278e664d29586bcdc2a467f2481a5a84b9aceaff5ed6ca769a3d480088ca3f44a981497
zc5d6d36b37aa9c9bc2dbe593e2aad1035414c80f7f9307d7f392452d3ad7f75d70407277206d34
zc7afb3018dc8d9323d275f578d9970dbd0e8b1760289c657a13b28b23f62ff8098e602fcad6b98
zb455d4409de513dc01ec31ee122ecd4408dfdc48f547fb236044de594f29dc1e4bacedbabf2d74
z7a446375294934a13b9c5fc6e3a075ad18ce7babcbf06d99b6cc70ea1ec7f65fa1dd42c4aaf925
zb548ba5b793864aa9e85d080b42e8fdc831d2ccb6c44dc8578b629e5f0f007e54ec586050d9d0f
zbf6a1c4b192bdd0a9fcc537f08665783f6b1ac332c4b017bef2d762bc3c317563f95ae74530036
z203b63040128db029b55de3905171de74b9745409994a2015c3e542c5221d48ff8ba463809868f
zc3e416c5263ec9cea3b4cf023d701c439fcfd66ce33f4778d1d5cd69e44ec0492360aad37d4905
z6a3db6dadc16391f1e5e519e3f316bb051e91db631563683300b448d77f5261a7aac3023896355
z0063ca021b53a694b4b8133b13bbdb4cff97a7ba26133aa5e8bdfc999f057327d637a5aae4be97
z2451bf99e1b18596b6b5737a5a72ceb64581010a0294de3319bbe8e5c4a05a703dbcaea89d48cc
z25905aefbbb4ede6bb014b8613bf1c56c4efad1917f3eb095347b4a26b06d1237ae6d17e63c1ae
zd39dc2df52d78029329ff72660142f66f9741bb5c50b0987b6900a51a6fe80bf75161e9f831285
z970664eeffb1da9ec1e6526e1794e59c0a8c87562d4a4d0ce5362e2904ea95a3328a9688635a5f
z4ac3bba5e9b4e8bdd7c29ef28a4bb78a858d32d8d6afe1f470ef460b4ef01c50f1e6e639f10688
ze9a7c49cbb75b6b5dfd4fdf577f437af1a2e75b605e088ecc5dece4712bdf2117e1db59eba11ff
z11a4d2de559c5d13925334d917a82fe6b4ef5a27f9f82afd8c8499295cdc7d422f1e96f075eb56
z2f0af3d347f4be6757c0e9e4cf3a51a4b004ca0ac7757aba1fe449f96bfe7969dfc0563ec29505
z1e8dfb3c5d29ef83186d0137d232f0a30e8a79f09bdc7e12c229e737b5caecb792bf411f18c5e0
zb79b2884befca4a65968c3bcfe9c842bb16f360128bc30a59516b228cffd40017ca391d09d1a89
z812e2af8c5fa9b4335cd4a0775f42193df9526e0332f83e8532c49979353bf6def0e577615274f
zf6f589b805e43cdf4b31c4196426c31a2a82525eacf53218c9f06dd3bb521949c9a0b1914aff0f
zb92e15d3a45b7e5a206cbcc84ab5a77a40d62e021243712e5165c5a44017ec28ae830595071537
z21f2a4adbbc164093a791aa0d40794784eafc24d823e5d4dcfcf1f51ecdea371e98588ff8070af
zdc4a750f537e91d0ae71f6840c202c3390594439701de658c7dc3dbb31c2d71948a59826542904
z772c9ae6343bb4d50d5caf4072c05a14455f9bd8a261202d42548a52f2e8fed84e253e302bd54f
z96d38e429715f843fb27b2d642df1669b5df9719dd974cca6475690a0204a2773102edc2edf4de
zc4f0b4fefd9079e91f286f659235ef333cd01a3af505a7a4803da401b6800058597962464e0034
za6be022cb8666d990f10b76ee4b93802347e9812d5b48edc282dd051173d74266d24b87198bef6
z085cb1ed0d462b46f04a263f66e1e9468a660c610a9d4a318e3bf013e750a0193503530681fded
z78fc10c9ad56e52b7de204756ffbd77c773cb5a0a1b1c4d2c0615b52ef9daa430dded32da697d6
z9832dcbdcd1855d3ae951f6c9ccfeedebaeb619527e53eacb5548cc9f7c9edc5d997085d7bd76e
z5433b7bcaaee17ba069c0fad25141dd532f6e33712a58da7f058c4936d1eee94a3d514c27cb444
z74b311a4b915f95e6fb14221b23b748c1b8e87872f5160e9a9a2cde2c9aa1be9cc4ccb8324dd4e
z4897b2aaa9c0c39359c66690ffbc43f90be0e2f2712bcc8b628f97934ccfc81d53079699bbadb3
zda98ecfbfd95a23b34b2f5505559d76aa6f2a8ca51452fdb2c54c6b441e51054c56e0dba4e8aa3
z1b4df70185cbc0ccbdbd4d264780b1bce0726cb27a00bbdf15239391932fcc4a1b85799a9b2085
zd36cd3559876deb1d34e0313028bca097c8f2b6a30f25b8202077516df914f2d388f01dcdcf67d
z083c0863ad6eeb63accf3ed5ca5ff092d37ec536fe98e345958bd74cd72f5cb547e517d22278b5
za203b0ca72923dbeabe8183aae7a2a4db72c59b2d9053a061fbb51bc016b32b8d51b7541f54488
z4c28509833f450eea9d8d8c12e943545c9d5487057890a4dd289ee43951016caeb91a93c671d66
zf1af3b40b16cdcfea99067c2753c5582db8af571662a16fb247c7f67305ed5d7b2a6277ea46a68
z982f4a10e5fe5e2c65f357037351d5bf03ad3f742711751e3c56ffec84e7948288fed627d1813e
z98b0d101b8279eec59b6f12dd6b371c1ee702873133f1b1f21522dd3421663d479be7536c40827
z873efb7684768175c526873118bdf0a9212d7d6b205e19993b9de6eb54e2e68a29053e0f7c47c0
zefe9f89b16515a469d6631f8036ad79542a7e940fe396d64569638c715ffd7e191a98d4ab805a1
za20ce45769ce9e151f0b015e4e8b37209c2f3bbe8979199bc57e1a14c545e44024ab6e24900fa2
z711f1ac89ddab8adceb00febb098a7c12af74b9f02d39e80d973ab76836bf638e2b2718feec209
zc76dbaecd6b7bd7229b3012b3162f0ab62f6f88df0abafe0cb5d83f713053a1d0f33c2529491a8
z28e2ee588f69e3ec939dbf4bffd5c1cad142ce91b01ad6139d3f82706df8667ae765d9ad7bc358
zfc5bf57751259e139976f2fe5c2c90a1065425c615e12c604e6dd5ff008f9f25498bfa61fb4230
z0312019f7fcbfb51d481995ae8b4abe356addf858d9085d08b61e3246143e33bc1a6c6c3065a00
zd27187ab2c412bad67f01ffdd0a82d593a86628a54ab546a6847d31ef9bdaf8e51a534f268bafd
z0893df92007da9a273f63a7e5f9e07b6f593e8f559cb21592561710a103aa81f81ba382964249a
z655045d6d0fc8e52a3e00e2325d16c8b50a19d5bbe59cce6cf8f16039d73be45ece1e944b9d173
zf5a42de8959af49ce983f07be9179282766d2f5d909cc31332c2c060a0e3c1324ab544abba484e
z61df638b56af4dd6e6288fdbd982045e29dfc7347dc50a3cde35b76c084c8621a2876a54275416
za5e80a56c1ec313c75616a2575bb3bb2572d07010048ef83c9ab2105d83e9b456f8f77f847b1a3
z264f63c53b0733d2722a2272681bba6946d026250c831737d473fac5515d6facca1263008a8069
z83e5e1e323d298d82fffc6974c20b18abb6f8ff80a7b2ecca525fe84ba96c24a1313f340936095
zc42271894c65c12284de4d3794161758a44128017d6eaf9bfeb7fdcf21b05a2c233ab1437a66d2
z168f0d275411c0081e02140b7336e3fec001da92e1843992b035dce77c0ed94543fdae77f752d7
z5cf9eec98254fc080fd170340591c5a262815b74c5ba5a62b25d1952ab01d35e5076c8281b46c8
zb5af788ebb537cee158b6392f4268dda6db747669332a1bf2c9ff77d1413754b26e0c252080a61
z9e388902e3ad8e8ffbb33e25dfb6ce910d9174b65ae0f8aca81de62cd702508cfca579913e4fda
z6f1bd2c90c377e9a4c591e68e1b46239b0eaf541f4b13eb4af1938395715ba34b0678a08f66e8f
zc69658de119faa688365f7363bba354daa22a13c7823378a88a07f4d2f114040d102c094b65392
z637c50ab7327dd236faf97bd65ed2732f03f8ae43541e69d5a1fd83e83120b5e436f75fbe15557
z751253371d972f258dd431b5112ff66b5e7fafa90888a837e72842496687c9b4ce144911c62865
z0ff4fb3aa5a41620ff44e84378ec76205c84548d505d4dd1a7b2ac24b3a85d5debc06915b2b3c6
zf0859fd280c27740cd6108ac30f674c87af16c18d1d80493476ca2ed6df3a72c517cd8d8fabc15
z3217f23091ebbf11bbf45e5cd5540ea5b693417a6ec00d9f8c035124003800261ee2b8a9cf1608
zc1ea464eff60bbd20ac257d9f436b4bd76ec443528a3b3dc55902ce4b0fc34558886c59a7baa63
z39f063551fcaa69bd195aa060831bc6d71d7f3ac604b7edfd85cdedc27e4686340e94a4a787426
z90e6132ee37fe58e5cf321dd3c5bb4346675b672e78c92749154e5309821db0eba03ea25c836bc
zdb070ebfd64a48c08e4dbcba898218685ed2b3a9f1458607dd72cb1b1f99434dd80c305ed9c290
z4aa0bb05921da75020266db4df3b990ac8e8fc09abf3af0fd6e961fffd68e654b8d4f13b8a7564
z9afe0a360f82cf591782b3a22d7734339a4f15a632da4dc6bf1fb5f79b4fdf135664eb465a6ddc
z62510ce7e6e51af05506c12efed3c96ce7865d9914670e55809ee2d71b3bd5532ee7558c1c30c9
z2d5d7c5548aec15d463c4c4ad5926a503d7e845e9aca63f8273a17ec416276a4fb076b1427aeb9
z697c6d59801965780fb69b1ca0ee05f365689070a2b6feecd3b3a83e3b0e54390a3d35b9a87fd7
z92b67d526403c89ff106e653eae0b854d581502d749875b91fafab7544a923ae597fde53f378f1
z1c2e82bc93628d9f20889883fe77d12142083fe9f7e33d36de04d225026ca2f00910fdac993b34
zb2d8999a809bda538a562ff8bfe457827bbccad9ce1f807c471fe559876253778a47a68bc3f583
z62aafc732708107274b6d3839d075c2de587d3c390cf3c9f5846e14ecf7cd614e6d6bedfea9167
z761be3ee429bed7156adb35e74aea9c7853cfda13e070ba452a068f73eba8ac872459c16b52ecd
zd81f225e7817190731c3e0278cfd8ced63e7edf77fc4ada7998c95318f1604408a303fb02fa189
z1019d5b6c07a854f424148884f34c8a0bb6db362f18170a5414152026936db6b9cd1eeab9b3c2e
zc5c2c1cb1d5019981fc3f3318d1b3513a1acaab0c450040eabbf9b45bdd222482b16eaa1a52076
z86abb141c78eace8f876451399ba597e09da3c1e4e4817a5cb53d7cdde187ae9ffa40bce3cabf8
z49b434fd176c1883effe6a1238746031e17626eba0cce81cbf4cb6c8ffb4f14b945f60ccb18783
zf376313bb727309ce235ef885667d7500fc6abd9a0999a46c6bd7c4feb12878245003b4fcf67b9
z91b2f52c4c3656bb03e3d0c16e17e4377a749be0cdf48dda86882d709667ac73765d32d2f0e801
zf4019de7931a9c596b5a8ebc253e128883b19877af2602475a20e0a43b60345b6a1bcd0209bf5f
z573ad272e464875c93b32cdb7a5718ad9b1e7b513a9b1abe71369c7fb62144b917a4bbb3f4abec
z290eef217a7ddcfa4215beb2ec35ef11bb9b5b36faa6fcfc59e112af19c9cb12d5c479c9996cdb
z2b9352d058e87e170c6bdfd735f848341090be3dd6dc0d31b55288d4b150ec3101b826dd38a6dd
zbc16b41de5571927643908f654fb4c274b6ec1b4a0f883e1d81a68a838607683b3494a855cf585
zb171cc3fd41030851a93f7ca20c9449169fb2023938310aa3e815762a3b06798ccaf84c665a742
z5b4a32b032537227a37b73c4f85d28d89f54ea62faebd78c4fbe18e7189e8af21af533ab47b2b2
z7722dbf1d5b7d07e1c85cd5877b458b965262260624e44791ba801f02a52514f7fb32575d8f605
z66e2edc4f34b693ffd7b9c1308f7ab8458fa8f83134948e976c14696b08d81da93d0ebc9648877
z1f4239cf84d35e301f1570cb94424be89ca083f01410b24744cb06e3ccf90c5022ee1597adc43b
zf35c297881f95d0d6ec04bbf023516de73e54a87dbd455e9e9728802db3c2094fae1deb7b04a3e
zb415d456805ed4bfd29c8d500c2e3b8b4e2bdd3298f80bfa0fa58f57e4c8856b8d1ee4cba8cb04
z27a38fd39c2f961a2ac978dbd380590e24ad4b1492c0d87e4d275fe0fa636b453de51d62612176
z42817adf0ca8ba9d03f0b70ecec6ddc91d48243f6923fe9fb0175f61d3745c8e5584f8717920a1
z1f918e8ee894751d4729e8da28cf2f2bf4a4f460f37d58a818bddc666ee23dbc2cb21db9c5b723
z02443edf3507b00c4810dbd58806b51b0a24ae46b5819fa91dc3c0f967ba583317b6fd34abefe5
zff52aa44107b9dcfa40ae9dfdbd29d272d79d0a0249b71a56ec01d8ad33ddc69ae0a1a5c9ee54b
ze1e6c8dfc577f2ee1b3a60163e7f97dbd014160456bad6df6b2b3eee01911e7be5b65e4d86c907
ze5105c4fab68dabba54e502834519489dc3eee1826e74339f9f764fc9cd739c5131439ea2b1041
z800982eeff76a193abc7e44bb69f8087f203a73b6070da6e268d908bd27be38eb389b6cf32d218
zde3e945bb05098b44f9d26d38d1f21efcdf91b15700645c63e62259f30268cc13b95f522465ec2
z874e9cc7d68d621563114896322d094cbaf33b9a73d5f20c7f6ff695ddf487e6f96e067d6463e6
z37d7166570add49dd96bc037943e1ab492007aa6719a840456c3b20b5ff6a6a34c1df60b061224
zbe1e201eeeb8b78a59bf64ccfbff487995fe5e7000a95b4d8c4a18e6703571a5aa022c10b5aa6a
zcbbd636c2ef7406c97e97b5fb4ae98b8d9a15ba0e526bae86aea1362708b851c00464ba9c2a4bc
z562fb15c70636d9e8c300e3cef86e30f376b2bf1837c9ef5692facd28daad95157c30f88c41c17
z92ccbe387752809e23841f6e3bbf0cfff723310e9f8a14de5b88ee0c3e699dfe27cbff65af14f9
z0ca1f7943eeee92d930ea975d3ff549d08dba91bcadbf9b318dbc5acf1045c80b1fbde8e067525
za168cce1c4
`end_protected_0in
`else
`ifdef MODEL_TECH
`include "qvl_clock_recovery.mti.svp"
`endif // MODEL_TECH
`endif // encrypted_0in
