`ifdef encrypted_0in
`protected_0in
ze74c34e226135848fe16db9ffd31815111b6d7fb642c521a3f628cf6da949865580b22efd062a7
ze90adae0e65e66a2c36a587d0a790699161455169ed55a01f2084f11770a774ec4c588039b380f
z6de9c5084882a40b79a175f5c2114b2b6d78b070cb806e1c0aa9258297f4687ab308bc470f0040
zb0b1de382961eeeaf2e279e1462520fc31c119af8f2b214846f56c2b3cd2eadbe4099496abff18
z15cec83ec4a77b868344aa20ba7360908f5c0de2a79abf8b3534b883bb12180f68b5d4beb444cf
z3fba8f13afb0abfe8fcc4294810f75afe452434d2d0f1166236c82f76edf1e12979f04bc35693e
z32ae028996dd85737a8f5adc1ebb94f39c940246e887647b64782cd7ab429b0544c173176cede7
z01dfb26b1f73408344a52b7e1f117f12bb9c8077b34876c2e6fdc085981637012dc9754765e1a9
zc512ce062e0b8fb16a214591f5c81e1353b900a611fe1f4886b57940b41b7f2ce99a7b84b04b90
z916f717e73bd10589c81e207ed77ec660a8cbed5b487fa50acde1b055c8870bd8676023f21ddcf
z9c98cc47cfa2d654ff1365d1f45035a045a66c5dfa8279050262ac56ccafe221d4824992a69d8a
z0056c786d54cd57e5ac49b6b8aa4fb7a6065bae21c146cc6f3a280ec9ff5fb2462d875a56f9ad4
z3de8931eaf8f3cfd310a65b585f2289e7418087419e699c1832e85936e09e6739133dd3d7604d3
z97061f8b9c90afed7ce1433542064890d559573596efbd13dbe29aeedfaa8de76ee2e259f0e48a
z879a310c03c4072e61157a32d8a17565a3ff7022e8cf19ed589f99531f4974684a962e8211ebf1
z1a180fa2f9cbfb0772f1d3e3cee8acb202b2ff875767c1109dc6eac271187d7b7df5cfd94b188d
ze021486c9e420d3c31017147d2ad6f8203b641aa0d1013bfcbe3afcd95eb51efd18dee75bc280d
z0a2fea72994d4d9b34cafc1016b66f8a0de1104a3a62e23141c294bfe80a8ad4dc7a5afc1af0c0
z03043bcf586f4d173e39e87a9768b359796af05f0d13d4be0c2a4fe2b208a9899e47c8bb2eab75
z7519af13ede30bbb2504cccb78a9df45eec66360a0690f69601993ea6c2a16501117ea45c21c77
z74d1125217fb10a580f7a45724ff1921cd67d9c1164cfcac1ca2eb25b6bd0fc988192740c3a1d0
zd03b9e8d53070c4f0c8f004a526ed67a887ba6f039d7208916b78073b93ecc4582916c73357916
z950c36132f042b2a638b0591ce2cc2d9f714e600fe58cd3aa30721249daa08739511fbad98a67c
zd34e8f38624966b0768e9ff1bb67f774dac41a18a562cbb2aa4442132afaf274f6211e32da1857
z28847a6e6b4e7c0e6d972022cf7f4768881931de786c80940506ebb710d372f4200d5c34d14734
zf574859e61279fa6f67590f76ba69cf5b097a1c8ff7516ce30e62eaaeaa371452ddf17d13e4e2b
z3eae3d019cf3ab079f38a95e66f9988e5785466934a93ec6ddd59d742bf06b8e58c3981491d6a0
zac792aa3fa9adbd1e12364535e5b5f8b97752ded2b217879221481eeb2b29194539070957516df
z889d29f894f27200aec9fbd112f32808e9999522940c694b2d9b52fc04b770f83c7e0d1a0152b9
z3ab822cfc3f0250032d5c30395adc97d0fda33133b2097b7a6702825dbbc169c4362d6bc88f0d3
zcc01f760acdd3240b5f86feecfcb14a3f7b9c8b5cf1f729c5e90fe97548d7af3ba187497987f97
zdee8aaa02d47777a79cb612ac35cd10ad185a470ec31f86f6ef904c09746c831aad7d6f630462b
z3a3947bdd55047ba8af47e750695526aa553427e76ab6213b3668d7c0d76012e4b2c3a16cc6e35
ze199e56650cb3eb78148eaa4014f6c13c1fb15d7912f3953846eb0cf2a43ba1f4ae52cd5c18807
z759065bc19777c8633d8711934c2f5f7e05df467bcda3a6745089e24472fe44e2aff2a7c78b502
z98db52b14c45abe92d0e2f2884b3fdd5c52530cd25e5ef6b3d1a39709ff54e29e331d947cbd858
z4e42fd8cc0a2fa311d2e314206d405bd0ec9c6f806dadd70274ac92fa3f18aa9980eb63c225550
zfb031584c7c0b57cc3800b3728f4f26c8faaae753344388d0fdb6dfdb0dc1399371bbe2f083a3c
zc8ad0e292937fae358af1e694b226b7a52c6dfa2b2fb7957ae8e848fdb5655d973a157c2ade175
zabac8592270f31dcb30bf354325cb7994cccc171df7aed9a312929e2059e1f7d5541c5dd73363f
zdfe41ca62e4376b64ae7df7ab39c37fe9c0567fd244ce6afd937b3bf392e1c1e18df4c2f15dc1f
z9a524cc2004a1eebd72c8612bf385c01cbe70838bc4a84861446b4660bbe65e2a161866d683610
z4d4cb6430c86d348f49af9a1b75bc3d7064be800300dd500b97592e742c400ba53a06b6b4acf1d
zbbedca25167f93e70d49b6c2ddf9a87016f1e42b0cf312d5b9b2ea969f50e9bcbfe95caa81c9d5
z5d2319cb8e536760fa2f3b6c519d9eafa73a1f2d56b844d35944b9c69b7fdd921210e6d1c2475b
z028e2311c3e138b6dee5dc308ec4cf246964206a0eba7ba74da3753701342d1a411b388b6e16a1
z0c75637e09b49db120da04f0ba7aed03d4ef0ed4fadd0cceb3fb042a4b00a96aa64c4740babb0e
zdd570788c0bd218a181a11b744425479d7015fa4b375828c51190ae4e3b09334f640e001a13dcb
zc76be0971a940b931aa43262b20225ccb9f7fefd16aec3bb7e013833cd931def6a4dc62163cdd0
za9a1d4d43e2fbc9d0c4d1031819adeab80dae5a69791461726668dc531ace9f47abcaad9ae24a8
zfa58e979adaabb4d7b5170ffcf09507df33d16bd00e078c6ce1a95b78defc9a7b70b3a54e529bc
zba786c22acfdab43f22ee55c09e58ce8093bc23c3fcdcc3389283eb3df5cf780cd60e4664cbc48
z9c30d771335b811fc1fe16e98cec222ef9c05569c94f381dfa9553314a45bf4814237d50908a65
z30f9f0fa8732d4810567bfad82d202650219eddd756563c594caf3c2cdee10a9bb8aaeaa28ee24
z513d266f38140b0af2bb89e56f4765d5cb2349551aa296739e934b6a08f8e20769e1f05c4d4740
z9cc5060ab2fb721756c4db612c21333c47044db7321ca0890b382cbfd9ea73c39f9a3c0fce514c
z0a0ca4342005495a0fc5916f1f985df5417b10503a6493020abbf78da550dc5bfe978475254deb
z57e4d69084429850298ad6014bdee546b54778cde7651fc676823e551c358ffc1f23e678e2468b
zbc013f20716d8ed92cec291e2110ac2b3ab960e0f5a9c2dfc889a32bfe60510437004baedcd28d
z7f5ceedbfa4a69a4fdbd7395296a3d9599c1ea52c24f36f4d2ea7897e56f7bd739a6a27f55ad80
z160b4952861f7010b013622fdbbed8e9841cc6652cfca3fba7d5e2ab402d83cd6f602b84f9859f
zc428db5b4f5dd42297b5d957bd421260686f0e2c9e3e017270735b1d8a9634bd137812e14ef841
z540c4643c1545d04fc99028ca81607d5502db1452254e9acf4bc44ee9ccc5bbc2936fef705b21c
z24033ced259f537da7d3cec7f215ead4805da493ca3acaf79c5feeda768f78f61d0587e26a1eae
zec1c021313fde2b0d0dd5d6ab6756fa6ca2039bc991854febaff5ddc63d25cc1a0413ebc5f1c51
zd462d0327a2d99d8a9d6d1f7d4ef3dd3fc78ea9add4569371dafcf0dbda9c5d8a050d98f2ad714
z3d5c3446ab4675cc1034281c3460a73d10475f6e99cb1946c04e64e47a5c309d19ddb54299673d
za3b64de9ea52dd62aa6fb5a402c820890c47c8f1a1a16d762d37cc98f6d95af03c6e1c5db5e8e0
zdd1dcdf9fe3660f4d8f31dc39be29bc768c90963bed20ba90b39b7978c816302dbba155c933741
za175b808d1fc5a5529d7a4e814af390371f3640a2a2cde1d5b3f91d9d320b9bfdbfba06402d2da
z2af7ad18c347f4031a689de37b8c061f6cc09f9fd9cc991b2590e7390bcde5605d7dc114eacccb
z618715d588f7f200309049de34b9642041737423dc10c0d6335b4e113d7fd8e51d78753ba1e7be
z7ca72f6ee4af02d2fd0ba99a64bdfe94d828407a97570688f08e38c647e874af62acd8fdc8aa18
zafd2da3b974462670cd922e75a3a906ffe8f921f0601ed2d0adecadefe8887b95ff56915945aae
z61f687a7257ed34a277041e0ea3af494e70ab60ac7f17be85ba3ccae25b9cb7ea86c6617243502
z23146abf332aeb51cbc650e9c0bca2d38a691039e89b0e72ecb06d2e2c6e59c6ebbc8e71b4dbec
z2e8e8bef13e3f2fdfbc98dfd59f37846636ef035d415a2ee95038c0a954ca6ccacb8406c9dd1d9
ze0ba9e05857d68728698b91e35e731c7b044fb7af162d5a36c482e1c29436f69bdff5dccfbdb17
z964d21815e76d478e73c804ac4a0e45475d6269e18bf03ebef79e01b8aa95e94bca40d15f46c16
z88c02e55c0e4ba228ae5918fefa23a8468f03cf6752dddb39e1ae773af5cddae6953200879cd74
z6cf4d834a3fb0c67ee42bbfc669a85b77185d2621b98776ac52ffbed642672e7b252ba6dcbd5a9
z1fd32470bada5ffc4f3a470c032965263a05bf3aad3ed330d0c9de832c59915f12885e717cbd8d
z94a66b16e63c1c20ad539a932095f7b72f379f61521f8cec5d2faeb15a81e260a74e9bbc19cc97
z1d6e5b00390db96470738b733d3404afb68f4e7c3247b3b33ab56d5ff265c229e04865a9a987cd
z32ee0f0e0b57c7a761e8ab78c8bae68dc0e6d7f99d65c70205248a5754b8012206dc836bbf4131
zb91e61f43c10141e96f236b563e91cf62eeecf976ab851130cb97ac9fc58f2e0f5909e5b0406ac
za39ad529c2dba877da97dba726985d821062753f14e7b8f36e8270c4be3232667aed921e146165
z825c9b11a619f29bacd824b48aab6cd22e7ffe93419955138b5e16acad975285c4bcdc66c5fcf2
z31b4d1cd3183f867fb192922b91966f6eb5d67d472adf92bb47bac67fc7cc4c11fce2868ccef52
z97c834423e23bb8e7304b38fcb1904979a619cee48391acfda7d8036d2d0e3020a77b3a2721f9b
z81ecc4cbaeb4f1b98ee7d83ae4bfb15cbdc37733c4dd3db570b55eeac833bde82446cf800b6222
z5dce93b7bc7ea238a518cc1bd59aac2e20a3415b7660f1206aa6127c6bb6e13ad7d2e86b7ffe1f
z07751b756f1cb901c2e9cee1057a248692fa21d1c6ed6523d455dc81188378902036358e243238
z71868a0a69ad9b760f1c8a8ff137527f76276a4c6cdd1fa93669b7979fb73973acb3ca88997ca2
z587f80fffb4316b4bc5ce30c795b1d7e6657e08c37d4446298770a1c2451e83c5de9f8fca6dab1
z779ff4c48e0660dc733143a9e8d09b1ad9ee5eb802f9083f9b0066cd86e73e402090648cfcaa0d
zb25929fee2b926a09bba8acb107008ef8e7949e8696c04e0305e73b9f90ae21aedfe1060241595
zf85dc6bdda9a1a1fd9bf6af8d438111c4679b7a35415b0ea3331127ff775239f369f7ff4bb6da2
zedaaf992396fc0c4ffb2b5b9a71cab24bfd117754ec57b16093452a5ab7943955e705abe7124ab
zc7049374174c1d6ccd3d0e6b903b7fc62e3450fb49e5d3ac66c56f76da140574a9d8cc36026d9a
z6efbd648a6071e9689e68ec648fd66bf6e2693e757d813bfeccf7c704106fe718b7e58cb1af7e8
zb6528bfff49dfb3075042b36ce5217d6a6c2e07e364f0691b1e9a52a67c4ae2152d8cb2fe65b11
zd8c17fd7231efc4823484a9963068eb2baefaf2792190364401ef4c685c6c167dd72edba3e717e
z82d6b10458f12253cf6471c6a9f51658af70d624d97b17b3f8405a90b3eeb1a699621733022138
z1ffb2e4fbe530b18eb56aa5014b90086349a6ec71d3aebd96cdc72cb42c04d14726e2a4e93ae11
za60f35ed0d5e1a2ffd75c7c6150f755f575bad0fd0dc2b94655d02739770522ed7ef2d84ede665
z6499df38b27a11d1c7cbd19367765455331b85d430a76c4f65645a2ddda5ebef86131e311f7413
z7cd87dfe7eafec87e674a895073c770142be09d540cbd8a49a893bd83c6e6b09e0780800cea4f7
z49646e3bbacab6842e31c109468d5780b1f525d3cf34b519d049c27e3f8f2b54c610793cdb84e5
z81d83fd6fbb2e23b298f8ba518c574f1913c44d3ddacac77657756a79e28c4689c75b3de1a8830
z1170a8b5a7f7bc80c4e75949a2e0649cde78c5285af45de897cda86e8f9de0aae5e0bfc352132e
z6bc1ac9bc0122bae748b3f06af11a217786c150d07506a4fdc4763f6ddd27a84234b4b0e1694a9
z0e4e1a4f18598779ed4e745cb24904445a37e60286e548ada9b9e1758df8fa26748880a723f09e
zfe23897000cc38ee6b8e05a601c115d0adc57f5ea17ffc486812e50a896187fb0690dbcacd1bcf
z003b8919357afb4d64024b01f83eafc57dd7a600d6ce8c71eacd08c106383f455f219d9b11c6a2
z9bbd762ab3b1956947286be28d6cefe0d71bf5a716952e36595de69f4e1dba8336e8bb3cf96501
ze127a52bb28793cc7459b1958b79152dfc392bbb883ccead89e14f963ebe31f6b9c73efabce21f
z727d6298bb5e5efcbf5d9f8f28da951d7eba780afc1f2f58dde2ebc5c278d11d41197d0e57487a
za02ee58e1a0acad782b19f00ac5f0382a60e0819d864393e6f4a36076cc74c166468587d763e10
z6057ac9253cdb763a869aafb8aec6e44c3be41875a1680b6a93cb5098c07bab85df8247377af09
z631d051f2f0c8bda25e4db54dc7cce4fa3dceeb6b3c1690872d37825d85f96ba22ec4c7e802588
z56cc3301d733ae2ed51223165f2d5668cd4bfb7ec3829e42cca6716dba4c6e8593d898d697ec5c
z8ef7734c3e9567b91bcfb58a76bf9d725b6c1694541d7a22c01d67f01c9badfe364029a8adae28
z202d917820e5a1c0b44fa1aa69d503e0c6056cdc0d18541df671ecc87aaff7a1beb167d5297cf3
z7968883938969bce33ad0415d593b7e239a8d97861652bdd4411a57baf365c9e766daafb088e09
zc4ae0d79db9a22fd6ec7b642e2f812f10643a9a456178482790f9c2648f9f8bb3e95a5d95d773a
z10ad83705205d196a22aa33cb4ea0a08b7df76630ddda1982edc3c6114941ba5e93620fd9fe997
z3c6b48061e8869e28e78b12f162aa97abcfd68a52816b97a7cc05c43bb64017a2f298f99ca1974
zf5277dd777b2fa1e654c18ad38f8ebb39521f47747aa020c3cc53b1e8a1301122ccb32b67aa57f
z2d88895b8336a260b792338211914686928b377c227bd5471de4ad83565c81734dbe1c3af0031f
z66011409f7e082f2aad29b91030dda85ad84bbb1e042105ff48d46a6cc114d453aae7627a20a1e
z21d6110889eb94d6b7979b0e7c5f8d875580220c45021626b708d8e1c478f98e25e7e2936d10a4
z6a4eaeed1426638f744dbc7b99cef4b382b4e11d9e956125b838f97735c388b5230ff683dec5ff
z5d47bd5e9fed68ffbd2e1a35836f8168a7f2564c320d27fde945a5a3852704ce586f16fb4e3beb
z969d51945c1b30f2a2a2cf5515fd1072362da73a0b3eb2d4aeec290dc0ee05633197d48231b455
zc09bb141654292fad270a06537734e1e7fa2f9c01e8bfc909e2cf0908912458f747947efc4ff41
zd83169668a5bc3811655a94fa7b9c4a2d73972c98f55ce8dbc8ca5af888232c92dcb5213fabcda
ze5d6cc01dd98b2e793c1c7b444fe4b84ccd71f418c3bb16560b8dc5baf54719e6c65d0c816b0e3
z5607013ceefa5b5f661c001d4e0c04e51985a8c47913fbbb7fcaa659d27a7aa653c05cb96d0521
zba652d17cb22ce648097d73331e8c65343da1c18b68309f89ae350497873c8c61213c18515931a
zca783e2d877b06da7d5aa9e18e9271e80e71ea0f232f56ac1da2b46cc22199483070d83e658448
zafe4f0df8604d12c13b83e23a9b462f1c5a273dab97a2c5f5d5a1ee91fc3c99ebd08972e329202
z98c110bbf1e16e376ffad79a8a2702c57df108c0db5f175fd707279668a80728d6bed09dc8a3be
z7d44a7ee977cf34f7db81607d1d179866baf2ee67165d1fbb9863f2cee11ad929925e9889c2127
zc31ed678436327b1c7c7eb8b298712be3a7b2e710fb444824de2d1e01611bd98c62fc9eca5ad65
z428b40b3c6ff4db67ce009a3cbe177cc4ade1146b9a50beb15b3098e3caee86a0b2fb5153f2d08
zd6e8b44087ef7df9ef53deb4efcab0f9585268d68b5a39d40e756c822f6503662c8990a059ea44
zd3ee0135c1fbc8241406ee30d7ff6ec728e350dd2ef613d25b2f911b7ae9d3005263675efce609
z1e32dc3b6b55749cc4791f5351737bc7aae6a2c10ba94a9314a0c65b525980f02c45ad12d9341a
z7ffbbcdbea78c03352e0cf6f85234d265e634112bbb176fde7f1ab419236c4d1f18782a66cd02f
z922ecdc95689ba35875b5d46c18c18bf8c6df7a495a143fa25564c6df7d095f82e397205933455
zbf8e20ae7ca4193984fedd203d36f8b27e75480c4f86ea96d20ac7bb2f97b8be11245d50480554
z15116c28471a2d4c580a1c8da85d2e754933638fe35387205f34ecb8fd1ea176e3e28832964f06
z4dd696270cb2426e0601b1d401b2744e8214e7efc4fa079bc9d9e84dc2e62ae590ccbb7741ef08
z416e1dcfac2d7202a09d8ea87f63a873050b973621c3be199c0f09cc1194f67e4d8fce5c7e96dd
z00d475828bf3d3fa3256c2d537b9514d73aef12c07dcb9b0366a22cf841562bf6700113cb5b937
z1ad639984ecb61296ec51144d5ac9928fde02112c50b8e30a465bfdbc2e18017025d75d6863ab1
z823bc9edc88a5aa26986b52136f7fcb4ab0ef7cf80812cf7a417b6ca9bdb1dfe2dcf2aa5f7a531
zbfd1f160750c5c952bee24a0d654cc110a72b888be044bd7d7b64cd3b1655df7d9629f5e108661
z4e8fb759142f08046d76d77db3e2223973cdf7be483a9a03cdb08a7fe0233129d1decc5dea836c
z51744f14835c1213237cf76b736ff3190d7060fdcaa3ff67
`end_protected_0in
`else
`ifdef MODEL_TECH
`include "qvl_constant_assertions.mti.svp"
`endif // MODEL_TECH
`endif // encrypted_0in
