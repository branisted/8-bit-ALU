`ifdef encrypted_0in
`protected_0in
ze74c34e226135848fe16db9ffd31815111b6d7fb642c521a3f628cf6da949865580b22efd062a7
ze90adae0e65e66a2c36a587d0a790699161455169ed55a01f2084f11770a774ec4c588039b380f
z6de9c5084882a40b79a175f5c2114b2b6d78b070cb806e1c0aa9258297f4687ab308bc470f0040
zb0b1de382961eeeaf2e279e1462520fc31c119af8f2b214846f56c2b3cd2eadbe4099496abff18
z15cec83ec4a77b868344aa20ba7360908f5c0de2a79abf8b3534b883bb12180f68b5d4beb444cf
z3fba8f13afb0abfe8fcc4294810f75afe452434d2d0f1166236c82f76edf1e12979f04bc35693e
z32ae028996dd85737a8f5adc1ebb94f39c940246e887647b64782cd7ab429b0544c173176cede7
z01dfb26b1f73408344a52b7e1f117f12bb9c8077b34876c2e6fdc085981637012dc9754765e1a9
zc512ce062e0b8fb16a214591f5c81e1353b900a611fe1f4886b57940b41b7f2ce99a7b84b04b90
z916f717e73bd10589c81e207ed77ec660a8cbed5b487fa50acde1b055c8870bd8676023f21ddcf
z9c98cc47cfa2d654ff1365d1f45035a045a66c5dfa8279050262529d2cac9e64fd27d9c7de62a7
z731bc808811ded9016570962244887f98fe5440167bd0088f2f049df882af501358497c3b28776
zcdc5426c7f52a851c35106bb93e16fff984784050fc808fad15da330f6f0607eda2d0e0e4b1215
z2ac5b11453f6b6c5c6b428261a64553d70b4ab9f1bf3f153bd631387c118a296ca10cbf0349426
zcf2ea5eb241fa84c8ecbbf7180f10eb9ddd4966d421e6ca571b198ed195474578ea51160ffbd6b
z0f73216703aef2bba31d04f6d0877540c760cd2535de4136d5bd4771107747c34c07fab3aaf6bd
z67c5eab3938266c996e67839bfd448cabe88dac2c17438997a3ee0a0543dc656070eb3dfe7c0a1
z57e24e01799b1ae1652a0133882b63649084f8bfaa3118d2448218b5c4119ef2134dee0d7a292d
z80c07e69250e6cb0856a07c01efe3f869b070b26474ff619f1ee9676ce10b0179ed9855d8e02bd
z3e17bd42a654e974019a7ca7de85bfb3ac5c169726f832c6b918eae789fa38ca70f5115a2ee7c1
zfb52b503ce6ce35b7dc5989bd64a1623ecf327040db427ea1518177d8423992586c82ca8ef5783
z63913b3bff1336b6e3685dbd63eb482c1694cc8e7bb0121103cb3f779f1afdb33a5dc4caad3fca
z3ad61f9e6798c7fdebf82270990759ec1a4107e22a744a216da0132a2888c982add83dedd55b92
z473c98e970f0292cb4fd1c6ac764bf3440c9b1318f8d50bc16bd1ece42ab2031f5f07b6b7ed034
z152d8af907ce476029716b8636a467a9c888befa1aad211cc2ca016bdda818d13849dd75a5839f
z6756c38996bf1fd29a8013133e827e128411df96c03f2d4dd330b986fb25411092dd6139c75755
zae52747bb133b5e191beff769d22d214ca12f5ea628bf4350ad100745bb8418051923afa248ffc
zb61c3a9d6421e116363ee723e50d4973bd4e31f429ae9a31099b059a7218d05a2309b6684661bd
z80481131eeead0db9cbc172c18256c04e6f854909427b806aa0e0ee45ad69e377208dc83a693d2
zc5ed51129cea272b74e9a010dc83dcc178dd00167ec5e7e5f6dd890ae4f1dee78cc49cb3a7d51e
z0d40624f1fe20ee0476fc20fb125f8cafa0e4c9168de2907249fc3abaa5ecac9b47411c2faf2b7
z1f13df756c63fbfc408c498e1b4396217c17c4aa56c80d379aeab6541df49e1402e596345a81e1
z264386c800647d62069c86a3dea531ff717cefa70c101dbe2932bec2d510f674217f108df23142
z410dc139440b2c0beb7c083e845035fb9a40eddaf0626828824c795409d5f93663425225f31dfe
za37643bd06c48ab6bfbbeb4a558b79a05eefddec0052f5893d504a969822f8503fe3fb4115069a
z76ce7cc6839a7c2889d111e55a83970f76ee2c0f39e34e59dc46841b1c34d12faf4ebe3f901f92
z8dd1bf5177c98874f81b204af4fa8c7cb00df097a75db15b83f72d46511f6448b2fb5b196ca583
zf8234bedfc25e8211a1fb586dae3d7cf0385401d4fda3b37a780e2aa2037af3929736399fd8875
za8c779727c15e851390118a886a847482cb6a0102cfdb2dad0d48e5c0d099174cd5bb2be3e2b5c
z119fad7b3619acf84d96b68ef5af92f5f9d0ff3584383ffa24486ae41f5eebe6ac371e9fa65279
z9eda50dd97ef1bd952e8005f9de9fea7a2c7991547a2c64ce364e5d29e50885007ae7b93db4e3e
z156be804358116f37c63c18b171b7a6b571434ebaaca71e1a7e5f01b70a82d92ee7a693f4e8253
zf41a0776faf54b4cf823df2fc074909a3b0e2899ad3835848249631040cafed6d01154b585da31
z57a5b95d8d56ddb66918b6a5f30c6b209c45339cb52ab02f6e169dad91c934603fcf0b17395797
zc456f44ce617110457185996e715ef67869366231a1f2fd55ecd7ffcb7eef5cc1378b93514e041
z42f37b8ba620d5574f3c4757533f61196c1cdce70f2f2bacbd9d4aa02e7b7559f97201b796d1a5
zff3386575d149d14125c815e4f5e6457c7f003706612bd33c68ef113673ed54ecad10fe172b076
z9a01cc2a3e8228e8bc3fd73e9cfc0dab58f0984d62168afdf1da4564b3ba4968ea6bf4f2aefd71
z4294103ab7a21505204592b50cec94b1ba731905627c8fc14d8356833be1d0550b4e6d88b2cea4
zd4289bee0b820d6cd2c87ab5f877c78782049d5b9127897895293b93f18d5f5e30219eac9c713c
zb9c3159c36932fcd77a90872c0cd9d142462700edd6ad3acd816b1102dbcc6147e789708f44c4a
z71b9271317b2e5a8f6db4f09936d47f2500f8a4283b2d5b119611684e0a6956f5f8e2542074acf
z0bd779f429d550028facbd4c91fc34bec7c0f242697b42d2d0693eecb49b627bbf6a8b7eca7f34
z165874073a609e37b11c05d0a83995bf0f5706aa82d7f0a92e956f40afae2be3ea9fa1380d0a35
z451bf3c1f1d6e9c3230afa53db4449ce2246b319eee9273ff49b8c00cc89eddd1bad7989aa0292
zc304096aa0a0e82e85b7e797318b57c4cf8d989bebf0e28f194af27608087a2e770e78d2239d8f
zff2f3b88fee9b56d368b08405f41c40d7aff14664d372145d740abe38f256115d0635ae9ff6a15
zb75c4c9af5390707172461580d383ac56eef80ff7fe41c4f1d72e6f77e805ecc6cfe4344391ed0
z0ccc668dc445477284e4f87a4849dc68d974254f242a390f88f9d77c4b915c6770f51273f2c8fd
zb54c6b2db3bbb196967856068bb259e0789ddfb9f90143561c154311f02753622b204eccdb6e26
z0fa6b29a78c1b419ef3d8255b0d8301f069b1a5ebe8e2e57b89fbfed11aea5686e6ee6d8794b68
zb6ea7d978f9b27740fda65bf63414a4c6efc4ba8b301f7b6b8fe29bcf1ed4921aa4b4b845b1ff7
zcb905f8d8f7bb5b61260ae7aa9e4d952677ca591e7bc7ed916c84862675669c7d2109f0bec82af
z61b6eb4b4a2eac8879cd3cc1a6204869f02951a753cb0a43112d326415a656ac9ac40e13a6ca27
z9d9b8894eb5a429a7c85b291b977fa40171e17352e3e1bd6198fa01532e63de18760c618b30695
zfd978d14a243847042b2fc0849a94f78df5d1274fa49b6f36dbba8d9003f0d9f4a14520f0a04b6
z7057bea75a66068794a11e8a78e165ecd1535be3cc3407cc3a49cb6d8aa18ecafc7d455f991b98
zb38258f2ced903bea62a7c97526a552b41b44b8bfd550c9ee80a31993ae70ee98bf1be0362a099
zde87b1f53fe2746642de29d19e6336a193cb794aa6872b6bba8b36fdd2aaab1d22829b222a2814
za27850e24c0f70805715c26e5dd9c4febc7e61fc30538ce3144caa78b8f55a8bf5960a682ac9c1
zcca9c2f28d3d29fc18bd4b15592d97164e04e0520afeb7e46bb44f4e56972d26f7c31b94e96a23
z7d750fffb27a4065cd5feb9d6a0dc382a30a073a794988d212beaa31b697de4524e86cc1f8dd7b
zf3ecf0884c03d220ae467fa3490086f0207888e090077f557c5db65a6e40df72c84c0a8fb9a082
zde877f7b83c2ea81dab9f64fc9f5dc56b69246ccd368c744ba14ca1635c37d2d18ac2c2018c49f
z569689734216bb347cbad1b43d6fc039dea0b5d16a8d33de1d2cecc1b46dcc9471a9b2faf9f9ef
z55a5a5af197bfce38fdf35a401d26dc671e7ea19cec44401d165f4b9f54fba3ee767d10b1832c9
z9cd9b07afad817ca2dfb81d528bd33de39cd5855927ae1acef773e5ff0d8b46257752db799957c
zc4fbb4f8d3e234e765758345ef79a4392ba91bba66a396f0079a0f139af057a656702160fc4e7d
z9a76af0ca1eb7fefd5f358081294ce8e59d0961f7be0d1553d1a6df908be63a6c15b2908ce6d95
z5f2c942aa52dc0cf00900169b9dcc317ec090527587432ad59d4848a1e0aba12e86f0f18a25197
za13b206c8872f74d0c27468288d91bb43d3fc409e5dfacaaba58f4c943007c03ce1885a4c24cfb
ze75cba0259b24231663bf6fdc3227fd715ca5e5916408587fabcfe03d779042a220f8138f410b3
zbf2d0e7760358dd2e85512fe0567409fb17f4f7d4925945ee24ae2ded5dbcbf11d64cd3ba526b8
zf28c0be1738c5cd5fc14c7ce3c555f9d669f99234c86215b2caaa76333da38173ff0bc77b65d3e
z89442db510f6bc4c0e47afaf4f6a5352d9de6b18491ec0c7fe2739f2cd69dd1b938b341a2b2109
zb2c26bd0b9d94440a787afa56913adc828984b14b3afd9329007a35dac948e28c024923a6de1fd
zc239403ff6eb627b55a860122bc0fcc66a5f4e45dfb2f3e24d719bfa794e311574306f0907f8cc
za0cddf81b1f2f60b937633f8ebbb32df04e9acb300065de07dc08f32d34c758284d6aa3d68af39
z75f2d446461062348fd328f03ea77d4973b1ee3978149049496b503c5e4c1523da1258fff36bb2
z49d2ac0e3f2b817675dbd9c0cf437e4096cbb661025e3cff99ee1000f578828239724d6820cc4a
z5e695f2d7f5c8d66f6743512c1e8cfd6f06a6f3834582d39d490ee4d62394e0397cf221f4f9c8d
za62637602a4f08670baa99b5741eb7947e55588caa0cc6b86cde6f34243d7e15c396bf64d0794b
z4b7fd361b3c4143ab1a4411627445f478c306f98e399df017ce999fe66bdd5473a0cf7fca1955c
z3530c8ec972d470fc33b97d701d439dccf50cb09088716f39f7a49377b5be8fbe164abd32a2aab
zbb8e2795be01f1182d5ed0ed0c2214e175bf29dcc15cc8b2e8992b6e90e5684b93b199b522a96a
ze3fa0a844cc842dfec7fee2ebf2fab4ee67cc9b85083c919ab6b6112acc09d2b9bde3efc848dda
z6734cd65cd815a7b49fc29f7cf93442005f273826eebb78b297581b288da99954166a81e58abba
za493ae1677e3c52ce4e878dee6b550be728e3d33d2edd79c56ec0096371112790f082bde75a145
zd5a9650a227b5704404c1860e601a0ee26dfc1602202fe996e3cdf14c7c2eb062e224d7d19c7ff
z4b5f2b1f37c40812ab7c732c42b1ff540f2002c5ecf963a30c71f033e2eba2b013a52ea607bb24
z2ef5d38f87f5086550999c4428f94b0db666e6e62a4bb080f94c1ab7d04668679943e0037bf723
z415057d6ec4b3af6e1a8cd145555df48a62c63d7dafdcacd0bed86989985c529454b6d51f5faa5
z85830ff0a1b1f9862860a1ca50f641ec3fb0ca889e6b894094584a5ab4f3b4d6593c14e380ac5a
z4ac53d6fc015120957c1fbd4e48cded646e7ce4683a6e47387d5aaf30076128946622321778bce
zbf6e456648cef107b94651fd592f666c9f2cbc904fe2a1b03c5175f4169d3ea03a52dd08eae653
z2450bbcab4af2181e414f2238d670cc3509ff0a584d93ac70d6b52bac7d88c030934d584cc19e2
z581699736d44520ee558f1ae2dd5b1fc8523bfdbe6946b8c04b72c509ba45ef09ea5bc5620daa7
z6f767b443d2e675c40f02bd602b4226229b22cf70511f7ae2471f199327b3e36f07a143a962286
zb26fb06ba6aecd687bdea1b8180e91e9c43951a740f687c9ce642db7197d5136ef53b4c89a3482
zbec23f3d2eb73f6625a549fac16d0007953eb162564c1a7729bcfe5b37fc83814e1f92c3041f3b
za679ff180c59a821ebe22beb3e8e18fa2adee743bf3936fac2964f7b5c7edcfe8714795b83217a
ze878cfb33efb0e2e09d0846ff46ea9d488a7eeb643e973f1864e87efcfefe91d7f0eb654082d01
z84717fb53713baad8f03c8b46cbf5120e7ebba01c8d399ca1f64cda753d2c368dab69207512077
z18d9c7f58d8f2113587a949fee5484578f6a39f26e0d0d5fd92f91700589abc7c937eba6c5c88a
z503e03a5ca5fe6ad9d9d4d04c0f9502f4c9ea89badff55cc7279f647742a164de47be176ec8cb3
z90d15a003681fb6f023b872913a83e193a7ea9c2b096e2104b2fcc17a1a1452226670c5680015e
zfac3d068c7f853e207acba8b32d8379743af07ca86094c9b3e9d24005f203f1ee3f80962046896
zd874b2068cfb01acae33c121ef1b2504c3761de4710b612d5ee4806b1f0e45f8e8ae511109c313
z21783d2c699639d3e8fa874c70f83f9a7a2bf6cf7ca0b18db796721a0e0e9e75f8b4e871750550
z2bc01f44ffb7fc85b8aa2803b932542ca64fc2a0943671bcd06f48947bd06f1580167cc72c7c0c
z9c787480084e131df46d0067f9b8d944ff57f53c60ba848f5414cf3438010d02bc66e4d3674915
z748aea5900d31377b1e9f099e9e3cc38e163d6f6acd14eae3eca946a89bd2f761b339092f1b4ae
zafe8a1e67c4ae6f90020f56eeb843c64b68efab897499369fb48b10d8e74142bdc5973de845f37
z15f3b34662a2adcaa693627e1a87abb979ab68d7b25cfbb80fbce8e6c48929d4f7a018f0ff46bb
zf7016fc6af737fd41394001284af93568bee6302e42656602e801592d17636b053fb18ddcf6a38
z5d1d9e9041a26d3e12eca39b35e89ea075da22e0be6282b211b089e3280d37d904a493482a9f4f
z8e6f4be8997de33c297b19fe62f46cf65138635ba07ba6b8fe0786ecff050813e820c33b171d19
z3379e6c323bfcb523197cde0bff6c9a3f1a4db0cfd804c1d8de12fae37aa8536a6b99ab5dda907
z95623334c8848c51088691ae45308bcc464f89efa0f283ab434ed400a4f2e060845e6659d500de
z9f78bcbca5181ccfeb287ae39d2ae2d6be27238df8ec2447a67bfdaedb7cc5966881cb214949a2
z964437775da12ec4ed52c78c285d5ada1d854cc7cfa8c6fa74c3a42a4d7d4fc3def5212164a507
ze6fd9354de777baf59461a72fc6f6d490892323edea430c71cb56af1cedd7daa922cabea083c73
z9f2e08d9bfe35a2579d9ec3918ccf77757d6eb316645a67f31bee123370a96e5b2c4a3c76154e1
z39cf2995c1279051ec0cb37ae4d468edfff0924cba9b4cb9e74ff75cf01440230bf08ca4cda1c5
z685a8db54d46a9e0490d5ba0eb16036a0e8bd0dd0f1be65dd0ba46ed7bb1ee784044ba14c11996
z65fdcc13fc041b48fc29c9df78296af95675a0a875937cac1a261e790258bf5542f8e3cbc0b87c
z1253fdfab79f516cea7b7bd712a9b6d0446859ef25f6b4925f61c3e47ca27d0193174c10458b1f
z6697954268fcd79ef70449d28d378ca7dc81eae301b5ada5627cab34a76c90a55c6a6d582e585e
z41cbfda066ca2e415d4ce36177a00332ec71fa103adc0ed2d2906b625a4fff443112de8f1c06f6
z88e6eabb2aa95413815dedc691608da2c6877ba772a7c753dc51bf2e1bf712148fa4e5896feba9
z36423b4ee406d8276be4beb8db5f09e14afb2cc6efae0e1146142b9441c511b59c66a62e7cf0bc
z22dba6c454b7bd13a3fd1bb7a9c3dde6741581ac333bb11b53f85dabc7e1610a63c74416a3a7bd
zeadb254288fb90de48a9712d65430c75da80afe25f48d4c4bafdb270fe04b71d762d5e10b12d28
zc462d3497f47349fd31c9503f3e3ec65f056168a10a6c9b1cb8d79c5ece58305d0cfd7cd7942ff
z4d51aab9a24ef9448824ff4113973e0b572e422a0d2bc0d77d2fd71b7afde32feda122eed6e2ba
zd6c3417e9c98647cec429eb6b4e83be90412d0580f746b034624b96bd875dbbf7767d6bce3cf53
z8f11b70e7a970a208fd7c6ee00549754a8e44b1beb54ba5df7e8965ad5921ca3d2603fd07b6e72
zfd070e4ae8caf4d44634a9fea9cad256c224142bf549c1fcaf0cddbec93fcd95eafcc795ab43d1
z8a1d69e04b38d4a9d28fa1da983cd2d20b5307d4f122570c056a7b231a727b9c5fb244372a94e5
zcfb5f994f047c7b1ec131768073f797120b69becfae79fe5b88b7c0dfb3d8833ac1ad4b31194cd
z314450ea361488cffe21e5795db82729c20968f0be9dfd0371d45862863cd1c7626f965f98c3c5
z8b1c3b2c77131dc80ab47eefbc2b580418d9113c33b44511f4392fd0cf5e99458715ba57256876
zbd2bd44d75214449f40aa89be6636d735aa588c75446c5e60b0aa058802cdc1e106b2293bd0740
zbc6823242f3463c2e7385557a40649de48380af0f5301a95e88b0a5a904d69febdf0a90a3d5147
z6f1f8790067f59a962643df29b7d91c2a8c341f07927e52a0859d11043d4d95ee0c32fea907af9
zf1f600a1f7ba0fb264515534701f683a19b015829ecd0c2cc3c8324cde043ea3c7a755146c38a3
z40cf69d8bdef05848502c4c50cb7030b5ca994a70b198b9c798a3d4fe9c0eb44dc935dfb67cf58
za1492a4a7b9df88725690bfbdf69f29fc588d1ae889aa48894fd1ca786776e072cfad89d028993
z260616c98ca5faa0cc150c3b2644410a3023dd39c005ae04e5df1304740aa3d0e80f7a23780264
z84cac1d546edc1dc976427e142c09c1e647d7fd3838ed852ea501e4bf3caa88013ba6b0f594c05
zcd34e9bd1c465c9fa55b0cddc4923351e2a9aa8c0e45581b90762581422080eaec303511653cfd
z865b4217e2f763a7faf80822acf7f37a0aa04e0f66921986e61be23e46b74925a76f2ce52df35d
z2574d517f73fb706374f7bbfdc1a0728d4ada433dd4df839bf8e35a4552f30d56f216d93f1c663
z9e52186f56465d7af0f9db916f3bd0e8df6f2e0b2da25d831b8c6699a67c642a9042f5183b8d95
z6b4d8d6defa9183fb39c5d7ca07df1449c53115d35f28ab045342c1318769629bb2a77bb8550eb
z05c46376a9c552de7bdb7b4cdfa28fa6a3408fe29118a6ace18ee83f1db0fa546f9b7f99686c9d
z29c219f8a5d2f908fd6eabf1a5bcc4de91fd0423d4262180f8179250589eec7f9dc3f85d758b95
z088b98f542fd9c32cbed5520619bfc8ff51917c99fac0e4375e7cbc5f05d401a89b9e2dbf60660
zeba3c30f642ac3114b668c3d55d62a43635fa031b1c2f844e1eedaebe0c0aa2442b9573002503f
z54cd33f641fa2a505f63013c6538dc2c223a0ff3bc2bd26274f7ad1e2eaf7c21c769dfac463606
zf5425f87ebfcd8f6b1276dc1eafcbbe4b63e5f032f5e3634fb37f5936730bc6b4295aa2b653a01
z375e74366b0de978b895e5d0893405721d8ddff68dd16a40d996ad2a75c5ca5463a97beceea43b
z4daa3d7050938e74545cc5230d4f4c03856fae5af1cb60b979da73816d291ed1f807caf64162d1
zfced5466eb454465fc74a8fb761a85e28f147212f6bdf1d7c4db9e0405cf4a3fee51aa9d6a1d10
z63b2f51d6db747886dc74485d75dbf6cba965a12a2413f78cca034603ad37d8e1de975da2e9b9a
zfd543201ca3c244467bc6c05eebdd8c639edbf0e1575daa413d4b9b56e6265b0042fe28b89cde6
z05cdf65ff9805512a4625c8e07edddc149afaa9c1bfbd74d2db93e07fd26a8123d71bc44ef83a8
z66d1b8a6f3f20219cd52aafdd8bc2065086cc163fef764d5fe73e485bda53946a75338e1879c8c
z6514b7f37cbe1d0c30ab3278e039d7f46c4d0e8874bb444bf213d5e4508cd15f22eb72805856f8
z63d768324f5ef71730304e295959715ca9d1cb6d1435a2ffb59c51eeefc514cf99c156bbb57fcd
z257cc8eb5b411f0e4f161196022ddeafa70f947c0eb57951c7766d40b4047896ec71000b5d8e3e
za655322eb6d94a8c501bb6a183a5dc45b7956a33034257154db00d38196e8774683be96151f214
zfe4052d44bc5890cc876ab3c09029dac29048fcd6ee7509c4f9758fad75dc2962e456652c1b22f
z89a69de274c0f20791d29a276d4018999111268820fa289cfe06a39812b71bd28ff7806df427e9
za85822319b294caf90cc25f3d53a20a3250178670dbcafb9ed5c4bd52af81a1cffb7322bcc2091
zb19c48e4d898baf773a388c9a941711a570ddacc83eb8ac9d45294e29b5ec51006d9aa0d79917f
zf90fba9090c413effc252fab9735e042e3ceaea52777a35060ef394bcbfdf8325ed23b9ca19167
z6d29790ab1565e5872d342b039768700d1ad9ea7d547ee952a8a38fbeb29b7130c0262e3a16549
z66216dd56b5d9b5772099262171fb5289aa87227888157651b3ddff2ef406d77c4ddbb8ec6c7f4
za8ca321590ae41db0cfab1c73d9e0077ef11d065d9879bd35c9786d59add4369329cdd92896789
ze21b6ff7be0e4715dcdc8d1f21022b70a94f81e1e40ca9eb75de9851403f17a42010f6a8e15ff4
zed1e5caeb934c564b426917dfd08fa6106b8f4961601b98f7c7e43b4f2f4a59f6a163efc6b2780
z3fd860b6749e5a4f74f02ba7bc5c01febbd3bc4cfe438a94a074869aaf547a7132008322df7809
z9a52239de9f466ccdf5f50a7a3ba84d834e015b874ae96af7151014e497f36fbd1979a4d29e836
z63e82849c742c80e59ae029a3ec04bdbe1d5723a2922458c69f1e0ca2f936d968121191f8b9a4c
z04c3b2753226d699b56a35e8be1ffdfc65821ab2e51cd3aec352cbb1f159fdd22957810de049c0
z2257c72c910048e545f8a48280530e01b1c8f8eab3b0678f6dfa1430011c11db781069c65712df
zc4b39427c7299d807be16bb3bd8d040cf9e1960e13b81ce30571355e605a5ed996f092282be950
zb34821f2d86517e11a6ccea778874bf72aad3b91fb1f986c94454fdb941a474cbd33b066b46830
z1a39de2baef874949e2786273cc8567d2dcf3bacc0449fdc6924d8d047c623da4e20b563659152
zae45176db8d555ccf2d0d24d2e96bd8edfb21d6a8cfbf791708fe5600d2c022175a13bf1a37a26
z31f6fcf3613c9c45a7a03ae6a1fadfd23c120cc931aea10e92a3392044be716e730c04e270d9ca
z07b5e3e8101d637f9f04cd7468f6c74d2fdcdbc73d135efc2d90abd8c9d984990329b1b86f80c2
z9b35fa3d4091508363d2d7ff32554e0ad402628af7d56d8f389cb23b3d952e9d1ae3a253fa5be9
za817ad45940824c95fc95d83c3252c576b7106c98f31cfb7245a97c8434efe882ff8250fc9343b
zbf46b4639ca7d823982b4984f96f5e3607e617a510906756c4de69b5fb4e0c54c142b9cf935016
z5403dc7589f0a8ea703435dc461e91414c81ceb7d678c5080196a2b382087bf83af9dde982c11b
z416c2f081e3c399fb080078a1756dbe6d462d4baf02cb7483f28d45a127fe3e30f334948380dd5
zd3a06048f418d993147639726b1c510ab5855f2fb52a6c8acaeb50c35c6e9f063e563e55752889
zd444e917f9a6b94d7fffb6be50752a7aceb30b44bffccb45b29e336be98827c83b3cf54474b017
zbf0cb437af010a92ef52d769a24b96e47af7f05c4c65597542ae66204a3aa3a754a6c2fff6119a
zda2cc1b3c2eaa7cede4bcb30bf13eb2ad51c41cd88826d69e03bfa5b24a93c23d2c33401a27608
zf9eb8a11b22fce67e9b2d8ae62b76ca1caf3637894c447402d7dca47a53d778bb56e162e3f7f8d
z31c83813e34e6acf4d47508e5797827d169c21e99be49eac40865e3e33f94a09b172b45b69fd54
z47592d04c7051188edc426594e4e0d74caa2ad103a225f817a48cecb7065df95f7dacaa1cfa332
z46b2693f89724ad120b7669f261e08f75ea468c1e97a2ab2232a64135e1120b47afb6ae505a143
z392027475a4f83d95c5dac0d7a7b1621efbca80cb8d69c7b9255b0ab10593dd3bb31a224029a7e
z7e945c1e3e54c1a0852a80f525af9af501b4aad13838110070eb623aa0db79eee30f1703bb753f
z32ccc8962761ceb36adfc6457db4fb4c3b9ece86e6114b164877bdc0b5fb1a02e1ed8118425b15
z8e7bc27a35ae855999102317d6ce42bef1f2b698ec5371f363d84fe33b8ddaf176ffc444a9a21e
z8451ac7695203777f0e7fc0f13bda637a3d00ae093ad62de012f577a6c2ecd293bdb166133082a
z8eab31d40fdd6e948b34486247e26f2c9a6784497d69d3686997f7fd3035721bfa467763a2eb5b
z372f6cd59832ae3f5703c148bd878d90a246438c8695eedf3f107c4e146c10122b791201ae5a83
z0cda6ec2d37ff8ef66c4a50a0ccb54e75a6bca24c777f718e95a0eede8336cee2957ea2ab58a0a
zbbb172d189248f2d94a6a7e899b2c233b34e25ff22673955a4b736c4d26d7cfdd22bc343b4e496
z570490692de329981c11df95d5d78a6aa27f7512362c267c7a6d651f2cc2f8eca0e85a60b62bd7
z29d3512b5d9f902df5665763dabfbdafc9921a2d467109f575687490aeada9f17f461cbf5b55d7
zd2841e274dd88798533d64b087ac7164bfe8496c3713bc1becf2545e3eabc98086298a3a9d09c9
z642dab0225fddb20d7ead4bff1bcff6871d301637f5dab862e6d937be297b7d9a99448d5c7513c
z9973e640ae787d017abe157a8950f4a2fcadd17c1653838fe7228446b6509b4a22d805999b2879
zcd754435f4c3f2896b1f9edb665ee3c7fe4a0d203fc055766c5fa0cb4f33f56cbbbd5c52a5d42f
zd2515276f93e4f521e790b85a2894758f97d3ad33e8fdc9d61a2e8f4f33a7c3216f55c110577a2
z720be3182debe97ac24df1cec55d934ac91dfc61d5bd3ac0ebed928b1750b58208b5a255e68fd4
z94a7f2be879e6ce4380b793399455c9d96a15b3d2d48494026a75af3a88bcba7e6f5a96550e2e3
zd00a0e1d4916579f32269eef6cc0eba513a5bd1eb0ce9d932c6ca189a9dbccc81b2f0966c4dca5
z2dd4b1637af5ba5e682ebc98a00103ee06ae93aa5877718e50b66921fbbf581d13ab74f768a105
z71594921e89de320f430520225faf3f68414166f9e0a9c46732e008ec15dc48010f64603b1d173
z8867a5bffd4fcc51a2ab328e3330f234d9a892db3f67ac0813deb9db239b41c4342e2f1de11a3e
z9f9364f843d6fde5f2b921b145399d8e6affaac12205357eac87a916afef25b41fd283c16d77f1
z121ed4c8bbc1d596ab878ac58b43bb8d87b57194fd7ccd21dbcdd6635ab06508f9a7e7a6f18873
zf308539fea595f823066a37ee6fffe2fb332d2710af07f8bc01b00216c1c6963a678ab8e62ac24
zedafa40a488d2f004269fecaf28a70d2f4590a44e58dceb69b71473668f562a18a3940b658af7b
z6b0fa95f1246bc08e9ed7d307ea874d3b7517f046a671c7fa74159b621364a504d075d71b3dcd1
z12be3640ebe9dd67825cea3d42b7a54e021ad0cc30194fee9b47435714afec9d75c8333fd5e318
z4a7d923dd10b10912b1b08ec80d83b7dd00054aae8118d58332570d31adf2fc0365fd56f050b40
z9fed7fbc8bd693d2077009e8ec0c86611abaaed3e8f086f0900dac2a1c3a6593547776a97f79ff
zd72a66c90e7fba2ec7d2f6826259fcb169232aa984abbe6e15f74f3b14bc5eafb511807fe5d406
z57dc7f217383ee6e0433661346ca2020ecd129880292520bbd8c091677557d515ca3c7e9729175
z71955ec44fc0a7040f5fde6ee8370485070aab5b3b07d8c677275c33213633baf749e8c85f7128
z4edb3af79e04c6bfc141cc78d24f273fa27c7a9c4d4d2361ba3f81a21e3bf62730cef0781882f2
za196c260ee2877e35060658c7ddad8c5d3e82b7ade8c51a79971d4dec3c7fad72220ae1894c793
z7139d6193c2e5fd3ef5122ed9eb29afeea8f140b14f958b2b65bbe02d24caf83d514b2ab4f6603
z600178c1fe60aca44cb230b2cac93a3711d96a6f3f4b25157400caf1ae3bdc949d8920a1ba100c
zb323e7796ef22f5c179705e333522b78f51471d6646c81d3c3a2c2257b73ce656fb1c819210199
ze3efece633a18f2f5b426f96bbe653f2c30c38de425bc8dd2a4309ec2c35c657cf024dcac0ad2d
z654811f07ece3916a1b5946e63794602e54ecab105d2812bd53c6dbf248e907eebf9083200349f
z9a69543890799a156ba3ff1f6f3b14c730e39e48508ac149a3602f94d233f5d4c79354f30d0ade
z7bfe74adeefa84271754e0b32433c34fa055e23572d83ce134666f9601b42fd38466aba51530bc
zc806500fabe258ca4b438fe0d0a7f84743f9039313a93e85414d0ee7fe06b1af8289a023e92869
z58f74ee514048528752eb575697f6d0eef069564dfb821fb759b4b7f0b440d2d7de3ad0802d036
z3f0c7b581a74e27f2d7df2134d7336705eee9f42c8dd7026cf2243452761b97b8324056e5f7939
z198af6b217711ce91310d224a8c9cf8d4620586ee7abed884094328c80858802b585e77c6d6188
z866d52b085bae74c0135b1fa7407f1f914784e118f5b8c26c25090c26ad0abaf742c519dd8161c
zacfc2238d3588de47c5f2f143ddc72b21f35bf361ec56ff6300d2486990288809061283935b7e1
ze9e11fd2a5c77981102fb909e590441ede84cbccd5397b7beba8dc9760aefeda70bfe26111904e
z976b5a240fb523555e49584937e2d66cf40a0ff22ab4195b3a249cb9525eb80a81d04059a0cb27
zdb8f3556defb37f9d344694dbedb5a738a81c548de1850039f1390c50a9662a5ea4e6538f97c62
z8640306c8ae3da3d98592f23560f8bd4fed1afeeb40e38cd40728d459736dd7fc63c31fde7dcf3
z701629a5b7788aab2adf774d15f31a290474cb88c52642ad17ea0addb3908ebc6fc754f3d3a6b5
zb5989f7dd02372330b62b67cc4e6e54c97fd4e79d336ecc776c15e9c994314bfcd4e16ac61aeee
z8f9f79949bb025a8ed9723dcefe95a61b8ca0c1bbd44b147ccdf22cffa8aa9ef40e22f6422f4c9
z6a9f29b6304a26c1c6a27234685517d80d695274f655b93c9662a94ec9ffc614a42ec90e287675
z9c496819026bc88cbc5cf538a983fa6715f600288a9a030823a706ba9ee1864fb5f2e8999ecc38
zcbe566353402b347d4e6315451e40e8c11235ebd754d68b88308ad89186bd1804c8865014eae90
z82bbb547a0ea05ab09da6e871ae08267ac5e8ebfeb1b73cd6917658e08ae307b6c97d7f05fe140
zc7465814db4af1a8b04dc5f642e38284b7030008fd7122a5b74b8ee3428bb9e9d98ef04bd054b0
za7cf7fb35a7fc04186427bfec0fecf41067608dd6ece53c90b0ca2083e89573f9a14fb73d24fd6
za26008fb4027d6a2beaf2bbed3aef7e5f02ed095a1b8620691019938c5d76527e9866f98de6473
z15bcfbb4b0cd3382371e0dfff0f9c376648599a604ad879a70b330394de241c0fb76dab072e77f
z26a160213b6565688a4f0c6566a7555bdfc7b10c4dac79dfff63166a6eeed2b3a52d185b04032f
z4bcc7a7fd90299d2867b5ac83ff8dc96879f523a03649c89e2c0e8d3d1c8bb01735142ab1a21ee
z0517928ab62e1df5bea226b2608db1241572586df2faeb4138204b904b837c2549d135e8323647
z69748caf766cc2aaff96d237bcf8e5131c3fce1926eb26113453854dc346307b0abcc3cdaf2d14
z19ef5ebaa4738ccf97a9809fed403cec1d6075ccea4a8b17d3a5f49a192c3d686c3589bbcfceef
z0ac0def029de58751fb2d397f4eff4f3024c0bf4e35fe2a0110d41b443c5de7576a5ac743126d5
z74678631309c3e0035e46efcc01080bd4c0550321168228f6dabc7f65f364a55c6fc64c2bc3599
zde8974893c885d3d681d6440c80fe1d19b1cbc2f49161b7907657684ee44e1a435d39b6e654d55
za13cf528dcebfbb62047decf9705692b6b7e649c84e905d4e8c39dd85aa554f9f8cc6003701654
z6ac3db3880240e2a7439d9e2c2daaecf1c40719dde007b9c8ec6415d6311a58acb25c455c38d84
z69755d7f4dc5004ef19d73f5a556c55629223d55c7119fbedb2e8f872a5cfd801635b230ea416f
zb72dd9ad471cd0999d6d5826d794c80534f099b5adbd291a043c40d0ec38030933138b7b42e763
z6371b3c91b7c434595a7eb940414b51d731ed95db3c4dabaa730a7b1d7d47e1a02f1a04f0ab503
z4fd470708512024d788d858c24f0ab57a58b74963babc32c53468011cce629d62c168c2877c5eb
z152bc2191e0f91c288e7dc0d497299eeacdd2956a4829fba9648844a42e24d6793d55549c53445
z2472278d22574edf069f93f1fa9296cd8a2e6421c0e1ac30a39018b6cb3d22dfb2622f8510ad13
z82a6721c09f031a584213fb2c3d0ae492d48de3c5fd2ac1c01dd470ec962bf72309a2f85f9c92e
zcdc9ba406412f6ea2329cfa4000e94a732a5345957c29c2073cea947e9c3a3db4a9a14141ec29b
z706951293508e81e5389c8deebf1d05bc10b125c328333c09411c54cc85679ff66381057cebcb6
z14c5e9be65d3d5728dbbfd188824ea3b61882c968a1840f0d05a765c8b2d4327c4cf25b92e8a51
z4eda012656f4e3f0eb6b9c844ce4dfa222d32a645a98484e6af900da6fa4e6c380f3fa6082d6a9
zce022c2cd99636d08f58b0820680690e5267ad0751b790e25fed26f7daddfb712d599c5a69be9f
z819502552aaae00150f05b1d51dfc3d188fa851f68ca32f5ed23627456075085031582ffa9df50
z9d5f3f00699a4c858d6cb47467fe681bac2230cd770307656d7645d775efa282e05d1151437b94
z03816cf1ed64fda02fa68d00c177240b81dd3dc2c5ea65e46498ebc9a3ab3aecf9548255161759
z832ced49311e421ca53d47f199a917c6699737ebefc629d184c81ebf2f0f6957d7f48a6684095f
zabff382f3716345df4b5b1c178dcb0b6653a9fb81e15efc7e0242c5664a6021d1c7ccfb1b54d4c
z9897d2d70d9584623278e7807e9bd97bb6029003d0a87511d0287d990a9d5c79d2825860ed8993
zb07605f62ab8e806bb6e6b8234b54e761f94e3a34c9aec98f39e18698b784b7f17c000e539c690
z294904f821d775ec0ab36b3ef00e1263699ade83cffea086ea5560c4239b9f74159c93a2eec741
z933cf755494a6f5fac21a73153469c757a4a155a5435d31a8cb820a0bad87bd1c6f834925581a8
zeaaa106ff48c78c80506189468fa283ba9614b23f88aa7f8bbdb75ff6e9b54bd09a7ac63ffb6a2
z5d102522f54ab77e7de2be42a002734deb4753197e28e0f7a88995e84f41deac658153de6d337a
zd64ef7ce78364190a424926755de009e9c773e9d55ca484396176c5472d37c6b00cfb4f7f3dac3
zcda1bacadb52fdd826db148c0e60bc1ba0d78c87a0b5c01866fdfaad1cc73269b8ec9c584eb7ce
zb853647d5aa879df3d0857c03e2204ea69be10519dc40d0716255afd5c64c83e826edc7e906679
z1abb6093c054c1fa442e8c44dbfe80f0ee477b5ee90b4652cd2bb0292e7bf066bca0aeb9f67b36
zabe95b585ef4d3fddf07a0ab06afc72e813c62e92dd97beeff156ad1ef86a1fa7fefcb9a53ccfa
z6f3fdfa8990fbb78ebc55ca43881583508962f8b920031f5be41024caeaaf2897ca20c3e85cb9c
z140e116fe0abbc9b2ba5c4c5fdb5c5516ab142c6a818bcd82e4918f60a8c85a2bd22de974e5778
z374cfa7eb985ad32fedb1dfc16569b80307cc96bfc7da1a10062136d5141390c089dd3ba070f25
z09d000b542eedd7e7db8a83a7844c144ffdb162459a548c1e637a6ef29c41040c30a01fc1464f0
zd308fb7ca85260a36019dfa48588c7f0c37dea4cefcafcab1d9bb96a81bdb506991ab9dc8df892
z75e297d416cf16f69940e4ec528977ff78a4b3478500c88380ff8f7bfd82e6fde8dd248bebc9d7
z7ec573d1cdf6a80d177010d488c0eef4be433cb579207981c351948497e62df27383fcd48c32a2
z4f7baf463a3b19e2903f58f75d1fabc2dd32583d7fb25675bf29a508954bd622e3ee843f4e54f2
z0d9b6c6aa004e647d6b9b8404a6176d655be4eb87658fcd9df45bfd1c329a25f6ad20fdd2eed42
z2c496a6340b1418e9dcebd3e3339c32ac2e2f63600d2014213edf6ae683f65bbfd369a498d0c5a
z008b002fca083d4f7c775ba50f30cee2a937a5f1dfb4f44a8a1aa89a1c4e30eeda0b324b509c5c
zed45e4ba3f3a59dc5eee85321fa0e4022654b13fe1bb2e702f655a7a3b88103e0e8fb5aa363064
z037da532a22565af1f4d404f1e4d899ce185f2a1a1dbff1f0ed4dce8cdd8fd0b4dd057e18981a8
z30ea8144bf45fb7857d8a9340e61f53bbd3524949bc49c66c5e68e0d81eeb60f88000def33861c
zece15042fca1bcf4a7f6ff92eb95f4dbd387db6092d69cadba8c0c4d97fd238e27e7f92f818a71
zd69efb695a4e0f403227c25552ca5a87f1f8699edd06a5b3576f455be38bb7c3308792c5663e27
z11dd3b7af86f858dcf0025d2ceef5e9b5c7973e76eebd06b1e737c8b8f7ba901ac590052377835
zdc6ee5c53d881b73e85b6a82886c5a9928f9894f796a84943ab45527ca02510e88498494f82080
zac59eae006900a3d85f6646bd3d8c9a130cd74fcfd92b2c3352ce7f4b388ca3caf3b2fb567d1ce
z21e7b50e8f9dd7e9fb0860db29899f68a9db18675f411aa9466015f8ec5b7fa29d783a4e0adbca
ze29d2a97b9ff8cc64339e7030cbc10fa0edb0afeeb756533116d4e1959de9e94e5dfe8deba1f5d
z63082453d06d510a0a07cb7fd055283fb931e5c26ef509c79c4b6b09e07d5b63a6f957ef19a117
z63bf1df3cf4f9ab565e96912910e774dd7be25798e84103459354707560855867dc74c19dce26b
z7752be3b3226697c013b641887f17e0504aeb82810b575c0e06e456e182e726952fd31100c2978
z1004bbadc871f7999efdee06b181b75b7d1ef46096095cb47ec98fc7fed523ae522be8f258dc32
z479eec0f7dc739533cd7f5e80978d195233e4656259d02b7a7536ba0da7f12e520f116b6dbc47f
z0a49aaf849e2598b45b5067e532268c7ec236ae8e962fcd9c410e4908ee6f3bf1a16eefa1d53b9
z5cbac422333e9747770f45e7c2fae056c10cb43174f1d04b1a24439acdb017d9dd2e791226aaa0
z7e55ae04d93dcd867525528ccce21a1462eed7268a0223c4f1b0cfdfde514b9ccb0723310398ee
zf7abe49a512b992a467a956ca97fc8af010066c6cef3d63d24f2b5b823868ff5ded2d34526c6bd
zea24bef8254e780d7218441212a3bb04a8a8d5523365340d2a8e1cf081cee13bc082a3b68c3818
z89338e59b7c61ca8b9921b8dcf18c534ed8dcce4df8ee49080562c30951b55bca67db76017444d
zdf4af7978b711a42ea0f0ef592e399864c9e2f7f0106d45362dffba460734d03cfc078a7953cf3
z194d8328776cd37c7d9762eec6570eb057317cfc192e24681661f7507ca028beb07f8ca9c3deaa
z620c75ec7c42dadedb5ac2e57c4b5b096aaf3b48a23053f05a1f4e1bd931908e727abb1043e3e5
zcd1dbccbc6c5a8ecae02425f051102db51c4f98f579da10b85460e35ed936c9f55fc75e7a1026c
z2a41257efca8d232b3db18352206e33c6dd5a9a4975f05f83b1826d0320ead536365255cc2c2db
zd88ef5df5e7869d3b4a0d630d7e456828a2a3db22da069a60ee59954c9902a18e415687b3eefc0
z7648ede54427ad8bbab1bbbb6f8ac3094ac7e0e93616bf79ee9a4516a1caa3d553523a67d6f0d4
z44d2e3f6772a29742bb479187a8db566a8db308e19162ecffd04b234cae0b3f4ed8e5b5d15dc48
z444190a64bc035384ed82a53ddabebd86141bba6aa42c6eeb30db145935d878fed685d8e824135
zd738269cee94a796dffa5fcd6c66b2146154790b9d11890b663acbd54e5503917b0e681be0c18a
z30aedba40f57a67083d308e7d5cd06a5ac64220116139b1061e97c299f1d5ed9c7528741c30d22
z949e6ae43bbabf5f3b94a62cdf91372867a6bf0ff7b1c0f2734c8f02bf2570b6a414eeacf35b24
z6647ce61b5c870b0bd2e362153dc7c5e45f34e77e8fb9cc27cb74acd642787c0e119f108d3d885
zc54cc9b65f9c3b5319790b4ee047efac9235e60b1893bd5291eaa188b47a9e6517661ccf040676
z514961a7f52618fea27705f02188eef6b92bce72076f794ded0fee6b41e14e61641fee5ce632e7
z14f98143deeb586bc146f23d8fd872431eb783ead926fc2c7debb626204565a830dec2408b3ddc
zfcda6598f26102839262cfb75b221762004866889801f8287514942c7a3af9dda9f2acce1bdc73
z3107825edbaa6103f3fc3149c1a6774fb4cbedc817d668b4147aa35cc455f724bd1ee3b98fc8b9
z462a4872465786545fe79cc0707369cbac630bb64aa3ef021959ad51eb6b2bc080f53826636956
z40b76279e0bbe168fd48aad006f5a9f851820ef55cd0539e567a9ee92051e367c55a853f86fbbf
z5c799750f8513f7b793788033aef6d4fe2fcd1874deb30e2d2c9471fe086804afbd6b58612a081
z5086f10fa76f656a670b436e1913135aa388a4ed4b8c01209ce5c7f6b2173c8ce1863cb86a6448
z970e789c47d0fec341c1606064f96503d8386f21083f0a06f21f6edd53b3a4e5b4c48c9304d8a7
z718f213b086fce9e0b668d5c4bae3a818b080d7e97d933b9cac6de3a2e6a091f82f1af289d67fa
z691a3acb4c5188fe0ca89ec59e0bac349d49c967bf1dd1004d01565572017aaacfefd7e27d571e
zc2d14c2e89fe2dbd2546a1e9ab053be97b83d560d6820de5a6892b8473df918cc95d6e11a72977
z81c7ea78036eacf5533c2242382dc86fb742a5d98d1211e7fb5b39a5c24bce3d75eca989a37826
z357a2027f6a169bc3cf85f8d24019857a97e32fd096b05af6b3dca6e4c733e68d15672f64894dd
z571162594d25a8cd1fc44130057c5285f71c494cb1f652649dfe75cc4ac6da38e7450701f4057c
z2e85d55a1d82b4db28ea01396608fb637290b2ef1ef1fa64eeebfe288e3fdfa178faa7b9a310bb
z75f2c6803da8eda84dd034075ba65575f50a4aff940acfd4d91c7afa1756adb135c1130540312a
zd9b73a6db76ae6257ffea52c31ca2501ebe364392f3e5a591946474222208a68a2f8534d59cea7
z7f15ce5dadd8757c77a565ce219405f5ac06f6e0dffdd2f993fc88365c684b0a96beadd8bf9f28
z81b7e9ffa9eac13fb6f614b884175bbf72f162807e5098ba31f1679bf4698e83dd1570c208a990
zd24e44ac54db3bf64b49def447808b7f6574f035d87baf733e1c0e7642e81ec397d2ad7f7aa35c
zf8c52a43a6ca7ffad46249869553428b3c95a37c0a866127b198df45474e3fd6489829f9301cb6
za88f87bc2e611595d75c5a613782599dfa94b48c78ff03cf39f4a919f7562a154890b44923c5b7
z30e51b29c8eaa951c3691c079b2a89aaebf6f4e182ea5d1416309b3867a7c9d04bf7f93f8b4989
ze365a632e96b233299acc64f39c762c00a5d6c20f193094255ad58f1fc8bb17031db02a91f1cf7
za7f2f062bfc672a7fb9c2396c2758653fa0d718d880db96b06232a09d9fa9cae2486402813c98b
zcdea30d40fa191964890d5527acbfa4c25f5adaf33ec821dfd55164c078bf1eca30996236cb451
zd706308fb96eb4e0e164ceb9682f3887943a63a08fa175141965589639af1ccbcf06978f302c51
zb9fd65a145fd63efe900cdf2c9e9551a11c56fd01f07945dcd173ebf847725daddeded10c95c15
z39b781502926c27e0d940d5843d6fe7e0d54d929005480077ad737a8ba9a95a4b95d50415de316
zfd2abc70ba3c6e42c05a3a03597fab8050fc61b41f8e032e45f0bd13258913f63b55836747f487
z36f78f9b335d4227cd131f9c5b1ba98240da939e0026ce1b0ffac1a06164624dab902c39887130
z373391d1e2cb098b4d3c4cf677bbcb299421ec93baa29334531196749eb1acd23a1e20c311b8cc
za306c21927e8a60900f191e041ecc89bceaa7cbe19005d8e25c109feade3c6f8f6db88a745f4af
z9c3b34133a72844d47e378e4fc1326115e6f36bed330d10e74a8bc7e0b8945d1d0a554b236bcfe
z9be2817947d7ba18b4ec8f310c053b2c2a2a1d3da004cc464db75907b2cabce12e2206100d80cf
z8035e9105d9338e2a90d2583b7797430ed9623c14f69404f9e98db645f3bed02759faee70fa400
z458b234107af7bd9127c3d75fec7cda8df00497956bbb35b0c68519e088c0b3c265263a2fb5fa6
z534e75062d2b7dbd3200af6dbc3b2b28b59fc28ad90265c014af16baba73a5832d6a01336cda39
z327af851f18d937c34ad7532b47b0aead01da320af564c523f42dea2b4717623129e06914261d7
za443c72c3e884e01007307468349f741cc922147ca453e72d3eb93717ce3da6c53e418c4c9ff05
z29b43af49be1f9843668e07a2f1637fd5a1f6951c78439288d8fa237caf196953c121d2eebcd56
ze26fd676fa21032c371e2064245cbb2612a38dae91949ad289621d0eb60618f96b2b69bf33d849
z95805dccf7434e45de726795f88b7773ef75b9f69db9e0d57caa4f2810b0cf8496a841afa5ffdb
z29de621828a103a9c643795c46c39015f5d764cddd601da7f893bdf7f915f5c85821e5e97d1d48
z2c429a9a19f2c87c8dbf6618e204317e00e7878b5db7e99e0c86e9db74839710b8e3dd8c0e81ef
zf4642b74ab91e30eb861db766ec3fb9c652bdcdabcceff76151af4f17f7fadc572d0ac9969ec5b
z8fb13a3308d631abe8c8f0cd8192dcc20e6ce0fb665ce2090862a196809a34fe2bfd8804004d6a
z194b07c88754ca3ba421486d7350bea4412645377c1995edb577d01a454b40058df2b8c014c60e
z78dd606f5e07bfb6b40bbb8dbe46837a379ceb98e10ca78842eacb9b6309ae2ea61c01b6a4cc36
zaf879ebcefb849575b3c14292fdc829b891db4960ef3a71b56dc1e96ed989b5bacf5a243d17dc2
z8e5cd4107c5d57b474f92ffe9ad652e0409433d366125864037405659c3f48d1df9e26a6ac08e3
z283ebebd9df1ac052f0642b30e2abc34a7f8b89ff0f069bd1830ea66f9c61e8d72d7f31d4d5a60
z982129d8d55c0cbd689c78d9fca743f6da7415e4cc078078c49f4d4bfef642357f1242d8f29dd6
zdabf937344f8a043d097b8e715afa4e4b6f69f766bf5424c6eaa5e3ac05f8abe32edabdd45c05c
z564cb76e72fc3013e8c8aeadd6ad500b29ec637ced8841e3afca01a634dd2a3c61cfbee309c14f
z986f0e2ac7148a6772297610b6114302afeadab7042220d049193f7348d3ba2ab6b2cbbc490fc9
zd8099c87f7a289f4495e8465048b1ea2b8e4bb5c9d0b9142de4f9525f4cae62f9260a435454337
z056130664c837e623f75300f0d89fa162b3880f8e5aafc3d3dc9d9ac9bd83302e20db33e7b4023
z38b82784f5f40fd54d28ddc84238af197a0f7df4d6905e6505bad8861153fe3e819cff943c3b14
z55521da68fc4f24ea4907c3739dd0dad806e95c0eff590f1072a9e6c4bfb1fbf41433b4f4a0fb0
zbc12d18e6f7a8d2966cf88c32a14438d77d39a79c33167ea48328df6ef01dcb8c64fc7c4e6f3d5
z8725ce6df334471c580ff29e0c1b6c2845256c2c1c62aa8196bae1d0e3d469829efb6971860586
z6d542d59e039f993989dc96850d3c17051bb82b68ad135f35a62e2d14610beb406d9661f37e941
z9c43c1f7ab3a49f4e28ee65663b0b332b728900fbcedbceb16026a3f3fdbfcb79e1833816fcb44
z48cc86175fec5e7fb2738c050d896b21c7fcd84192947d477148bd19ebbfdceaaca69950735182
z5b6373cac9b1efb0f321cdfc1361214389aba5a592da17aae6ab285f45c2b826cec5504cbf963c
z8f02cecc6fb8827c6519d74e4d0066bcc7f3e235bde0a5866e24b148371f96511643a7ef35880c
z43e63fdabeec2014f7d7962aadc63e445f4a91a14cbabd5c284ecd1a9e90e5fde54d2cf6944abc
z45cda2c8ef3316a147eae4489114915911c85a74bfd30e43c43e6d44b304443cac53b37cf87e18
zaf94e5542427485048980068e0474cf99268434e6e318835e57658e7892ea6a1454c730d1b2861
zd1672fbe9784c402c4f14b341658cd93c4f4c84dee1607ef29e4d8786fbd09a48fe4a14f500d8b
z7287ac1cf274e35d74e70f2f878721f61461e32c838b3f14231a91bb7c8da10c2da611250803f1
zacec19ff0ce2421ca194f780c7b395384429a3b33f8d4c8eb80add90185ceb18d3b8cab187ef20
zd15c05d93e8115cce5e5a046db5c1922126f6a6b4e791d8b9446a210271bdf1068a9afa61736dc
z431588090688a24b0b19b89ad504eea43a5abd9309013b87c664411d84ad13c5e17f336d954031
z8494e8481fdd77247f726f511df05242a3c4ef75748c0ef8be19b299dce565765ffe31365e88a0
z479d9885dfe228e1cace8f89daf2128789da028bb0ba2016f937c6eeb4b81d779c49075cf59c27
z1afaed9170804e2c5de4183eaff26aec081b75e6f2e40bbb7287e3962b48123ba8987a44ce14d1
z17ffe108faa2a497d0b70178e01b672c9b3a75ea4b4620ed0a961cba05fc9d9ee61af49f0c540f
z90abacbc36d9b459cceb0e2821afd71454b4391c8d16bdf3944ab72fbbac40092c17c65e317b8d
ze6be4184417f93838ee78dd7243ab352419898f8ead8123aa04f002af021dba02efdb2a1505550
z23e706f0a18cc5dddc10d99457149eb1537ba1eb1780450f034d18fb6aeab1d57a36ba4cce00a3
z844e136832f9c382addddc2e2ca3cbe584fb1f7af5afa0aa9899b544a6688cf9f667e598e59420
z46f3f27b2bfa93c55694cf3d4b4e04ce70ee61869e01cf50302f66ccdc21e9d076fba35372b0ac
z711f0006543e8d43152b36f6db9ec93bb0f0c4b814ab80968f6563526190c9d6a4be121465663f
z4d8cbead87fdabbf0a1854f8c06bb005ca30dc3ca3c28d8eb043b5d27ed7818eca3d66c3fefe89
z975fab6c0601435211f07d080dd2620a8fa132bf2cb650b1e0aad03b3293f15e81c65f72183f4e
z651afbd3808aea0bc49fb16725bd592c5054209b2f381880babaf35e7d3b85a6fd8e97b914d9a7
z578a80bd8e495103aaffd256aecc5eb3a7700e67ab94f55dbcb5c63636a724979f8ff969bea2a2
z9499c8402e8585daf0863053d04c6997d9be239a5a096f82733a7bc74eeb1d2093106fde79284a
z4cd85d2d6b6e1819d7df824cc37a3489ed524a7ccae753f856ea5c45037dd02a8058155163419e
zc4fb5558cf30bae2224ad6256a967798d24c528220f862a77b940bdf7fdd39950c5199ee755028
zc2c024b37e9f5653ef83c822ac06c4e9777e98f72e4bac9df0e31d147799f9c1a1dc2a3632a23b
zb49d00a56daf49c02f2d97057ddec13aeb79e256bd2d45bc3dd15d02ca176503733483d52b72d6
z5e7e29d5dd3d52da39c341c800bd3723f5c2dff4078040f4d2afdde3ff0b53506f51dfd0b1e35b
z4b3a4472b3efc1eed1cfba2ceb0a8fd1214c93d9d908b9bdfe9961884513916fe3a35dd2abefa4
zccd814415949d0447b3113965c52725d98b63e7d5addd529080345d357f46b530f9196b498a409
z50898d4c362e89ef5c3d065de7c3a2f378c39b2623a3c9b9246e986c828bfe97f5f6846537842f
zfab9f86b7de09d33f6f4708993ba8844f76a4baf820e0f7c6c3ea3025266c891d2c2f33a90a913
z0253e24e07548df4c78c594c22d6f59d424f510ef8d92f387a30a64b57c921113ffeb2881618b5
z3da8497cc06bd17b594f72714f3902203d8e9f00cae5d5ec464312c0adec0056e1cb02d316ae04
z56593ec1f9bf66a6644798becfee48113439adebc6286ab05f235bc4d8813a624b45ee3aea4388
z7c7b2ff650b8d4dee5608b05e33df1078dba07c5082dcdbbe83560858f1b784853fa5f943af9f5
zf12630abb4e8bd7a7e500139e7189ebc7a1bc34c164a19cde4b8e306d7dd0ed0219421e759c0a3
za6ca6256171685f4594472a8c36cba41e67761f4f052ff87db2e3072f7bca4a53728a5b35b8cec
z76db45feb00aaccd50d0c42e15897c852b13a1a876639faa581ca09947524315f111c74d39b89d
z27e45913b407b1d5e1adf61687a3cc0104b6fbd72f5febc8f821b58559427f846c0fb556ced8dd
zdd0d3921a992254a42fcad01a674c76f9760806053385ed3932a8dd27ec5376af6aa8242381aa2
z79be121dcff0e93748c118e12a29319bc0efc5ba176053da86f46b1c606066eeebf959d5a21bd4
zb168f5550c1e84f25c98c96c7fcd2bc9077f27744103a078090b24e76cc23af35122b407399189
z2f5654cbe6846a67ec6b851f8dbc8e93a76a4ef067fe3c55abc47f2ccf37fe89350c6df4ad87f8
zec0dd6b523fd27b51810d1d0a19d8e69f09ad1a6398c58da871cddc3838ea11afd74c4676bc937
z2ed8ab4de87202f9128f01c9914689989b4c59f3d1dcf2b0acbd9f39658a91e877098f8c2801c4
z2f7822023e445a8a24ce0196a2eeb045ec48ff7077f855faa34751f7906e84f1a928586c14216a
z0ce7cbeb48c3c0bce6212de31913269af633b2ad6b64a044190e826638df45a39c93d819dadaa6
z26e2c063d39966f6673c6676b61bb6abf62a290f5c13a987d00bd7657747e60e96fb1ed6a55ecc
ze975f0c278f0c7e3286920d875233cc1149078629bddaf7fb75e5742be1dec23f3b4438d0336a7
z2d04cbfd562c8a722f0a34b20ee1858f65f1a5eb4508ff2ec85b400762a26f6ddf899dec3e3f7f
zce030bbbebc1030593e692cb71f079b345d749829918d67d720825eaecdfdcebbbb31ce681392b
zd410758bb37b536247ba13cbc11d940ef1d61dd1c7d4097b846498a401cfcb8b2ce56351356575
zee9a1071e5cad5536fae79cfa52890bad3b2305ef7c8aa5fdd51f9243d0e1ca75250ae9a2856ed
za872406934395475bc6efe06ba01a6603ca25ad7a9ec6939d807143e582f37c9ff8ee136f02569
z28c37e066a1f12f10ce8424aeaf89e11c1e190642f34ed054b2cbde6f31fcb82082aa6501c42a4
zb010643ddaf5482405828f8dfa38d8945278b83199473db010a87f1e020fe727c930cef8e97e69
zed7bce347d1889ef2abc1f88a022cd2f91770e8903a557c04c2ed37809e754a80a59b57b2a553e
z8e6c7c5891d1fb4bd1a1df1922c89eda7782fa237697de9ef377760c161188c6d463354375400e
z74ae18e7331217dfac8e355c0aacd0e4e327c0a7779e87119ad92c5b4ab1807fa91a4e8e99d0e4
z6d65740750eaf84bbdabc22ee4873d43f948dc31a7332b466b761b311f091f8c2153d29fafb30e
z898bf02f1d4b422fce38854b6282ec499cca66bc49fb0839bb94de93f7f91b0da464d6c3e474a0
ze7130f688f60917f882da002170903feadde7fb842870a11be338c76a353cc138ea0568ae6718f
zd7c6b57e92c8818e87dc9c9718645403de40324db87f825144b436ff3b36a8d2394062ce5b597e
z5f21b92f8bb130144412b4ea0dd642a9c8b4a1067017887e97382da0b0d7036fd185c7a5fdab1e
za57ed23d5fce3424880da8b7119af3fbfe8d7443abab86a6c78efaa2810d51ad8f950a20c14bae
za377b403534478cd0081df32bc9aeb07473777170255e6dd635ee3e0d3a6767cc4aecadb411b20
z12ea50d023312e6b30468259eb688c4c2e4a3d613abb6778bacc51ce31f9faee4c613fc148a1cb
z018cfc24205b14c66e55145c919b418c4ff8801fc0104fde0a81fb357dac6947489ba09bbc7528
zf4855a7e3d46b8473e42b10ffcaff2c5d72218c2bc321dd4eb18315e27fa325ee898b5938d05a7
z06141bfd58e7884517b979c265076564900c09cf40abfa45c25d9d34d5537c35874c7cb2378fb3
z7413b90e30a6493f5037f0b450e190583f768f13b1e59c3ceed3bd4e991d2a44f41bf82c6e05a1
zdbef972a2fdd2401093b3bbaa11e5131f3f9111dd41e1de2d5ce321f2f7be5ad369aa4ca75bc78
z6f4530ff0063fd609049f8a8fb57c31b8fca9d22fd8fc5e0dd6f58133d1656a0ce5ba303414e83
za2ea8eb900a54cc789b606d82f77a63f9916bc2c6afb510a40be3af77f708a73b2626d6516e651
z387f12e5f5e3e07cc296fc88266ea46c24c2a053f43d971b5c0e429c07b07f509620ad6970e908
z5fb9913da551b7b576424be8ff2c50f9bd3cff6b997a4becd6cfdb4e60f7138ff644b4ff57d853
z6fb1bec82723497f2d7beb88ce96e9dfd02170f1b73e0b504cec86dc53b24bccd372d6a7e5a9d1
z9f2457afb77bf0abeb8a67ddff38125c3c5994e0aef9e341e9ad0afad69435eb5732b40a3b03ea
zde21eb407db72fc637f25e769f96969f313c83cb18f5d2434c0061bcbcbb4096eef234f196f92d
z38e1214b9810d1303eb8b547c82d973139f9c7c8eeb81b8ca916533cb39bea9a18f68bb01205a2
z1bea3df0a94b1ba214e5c548b47775cc777e81fecf92607a19dd3cbd97c45ce4555fe21812df7d
zf09be5ddfdfc363e16733cc771ee57f8fe9e103f6b30055c0d1b4afee91c0ed17f217ddc6bfbd7
z40826a047044cb360bb2282810718dadf21b33b2af0c97b18b4de3f60459888452a5bd72b8f36e
z08a87fd5703879f0c22b1058c2d171715fb2886e6394c041e18f8650425349a5dcd7aba782b09e
z04b59cf5dad0a5fab1add97309a271798d8828f248f46fac9acbfc93be005f6eedb2bf0aeea3db
za50d2becf582263c290669b3917f056b73d89a1186cbc1eeb892677629c62cab6e5c90defa38e6
za7da5c2f231c8332c776e41383d3142c8524a07196aee6b07cc5373cdb5adcba2029e48a569be0
zd88674c68a380c595ac6af01d0b8c4ebc44d3829303c0a3fc43a3e374f106a445fa129e24b27fd
zc622a95c082c49aabdc1b70e03ba7c0f55dfcf9ea2f9be992fa56ae6e58a5af812107530a2ced4
z705bb93e90cd8c4b06e480358e3079162057da57c25c00a7aeffbdfc347d7496610ed11dc903ea
za9717907cf0e793c111ca1a86d6eeff1e4410419f5eac096b06ada1e29e2083563520510714011
z82408b08a0feaa61693e551e871bbe5bee330f6d73b1ca35024abe4f7d3be760dcbd6b843484d3
zd6bb26590ca9fcf9a050dc95969dad70e11655e99f933ac79b87eabe042b4c75cedad30c5bc73c
z40ec79a980bbab779c9c8afc655ef34b961613dc798a0d99b986d60d5b0774ab2c9685ca15be5b
z46dcaee2406bd5aece0167d93dc14c41a1c15652f9c35ec446417154648d2d0b5e561025a7dff4
z65fcf9b5032bd07a641586786f2570feee17ef15c2ecb528f91a46680721952a7cbf944764ca31
z312ac5e417d9468d94a65e3150b9b0a895f1f06a13821978850cc76feadef4726dc4213ae88553
zb4c517bc0a68c95139420750e93be7966d0b147eb451caace4f163ff9e6145df351e9fe251bc72
z5ddf215a46ede208d1a594a3e044ce49e0da59fb91f7b59d9a8e83c5cb0439fd6dfcbac5d29e8c
z4804ce8c40d6a83850041f07030c0d66427249778031a6dec7b7cd7f881f42cb7266160cd90ada
z6687641fb90b7351fe880cb04ec2571e23301c414c7dab30c146812f6505a0dd2d2b05d70c3778
zfb9379f5712bf537fdb73658db65db93ef8c3992414196ea6d2890b93c5f4b08c38f28744c66e4
z00488d53e5bd99a26c099ceaa0d9d3d9207702b1b0e755d3f23a6be8f37a5ebecfed36ddf45933
z613d80319aa3c64fd43b67d39bd8621762db23a3da0e65e3a0a7528264d493bff7e106d37a740e
zc6c87716765b1c6367df1c77e22f3e4a06ec5c41ee638c92d5e1aa5612ec4f0b5be83aa546e107
z51b26d37d8ebc0e6e441d20afc649cf78ba3189dd22b9332f6fbb0183f95209f9f90707b1d5001
z39a395dfc61f48d38dc18a03b89829e42cca61cf79545611e42bc3df758c405608a6fe54e55153
zee3ceb03313189d242fc38ad0fcadea361e2e7ed1c916e945e2dbfbabada128972c5555da1bd0f
z22b419db1b65158695b5b0c3238e6ed73702c554e726bbbb06e12e93836d6b00b17b25d4008713
z77cb674e469991603bef698b5fd357c3fc8829175d80a1857a4198562881abe2acf0015cc189eb
z425dafbefaa82f868cf7c8dfdf59fcad40893dddf4a9d3222bc4a6271b1eda06ee95c4da0f5b36
z901efa52b8673f1233d96ea4510d6225122ef62b5fa1c834e0b71cf17a72e11d0887f016df426b
z669954a5ae1e94a647d634607ece0a36afe515c5c4c6cc92e7bc4a0e84f1457c72926f4a13bd1f
z70ffa3cea3e11ba65e670e384750cb79244f0ff886a9174793526dc0eb04292670b09a8da0e75e
zf836707c2b4b3a759d50ce28b6b690288293580e10af942bf35dd41ecf0b532e389d935438018e
z4570a7d15ddd6f68d5ea7982e3303941b598120a6ce71a7300306e3278efb1c0a2efbe3bcd848b
ze3fcb9041aff75dfe9879727f29780a1411b24e621dbe5186b12e37511a55c41b2c22e89d81f9e
zbe2f54385a3f07197ec428c175834f5ea57569457865ec53ecd97899277cea807324d81285b11a
z968d9ea80306b389a75b4f0018ac8e01f859b4f922779c2bffb635c3cf3e1bd1dc58007695aaf0
z0917ad2e0692384f741ad84805e57ea08e3d2b0685bf9c629008ecb4888ecd71f757879ada1dfe
z5d1177a93d1ae32f2b05ed1c136230b55171e0883f98a874f75a94f08344bc2f64638d6a92948a
z0a36ca8f5ea5e683ab35ca3c940514af654dd4f540225d55d3c9888a956287e6b3d4276ef8d983
z2762642a4cbd4143057efa92acf22f9ddecf8f2e890858c39d24daf530413ef8e4db33d57f8aaa
z8929549a568f5efe0f43311bfd50856afb400eaaefa31601fa6734fa17ae5ffc5e58b18cd68352
zd6aabb5143eec5a5f4a11ff21dc8c11c72d4124da7198605dde8d242751978bd1cca8c92e30105
zaa0cc5943853bbb253905f95f6e4b0caca3375bf6e7ac61778bdb0b0f302b407ce725f125bab40
z69cc3cb805c6c83bf447770be4118b2f72b34fe283a98b2a5c286533dddd01eb5453970ea0991f
zb2e2eade52214c62be76153db341297851da1121d101b8391f2e5d8fa73e07d000e3045357b432
zbbe7fe55df8ee0555f4fb646e1055bdd209a90b898e88c57ff8bc6a7271c0dde48cb87dc379682
zd2bc04e2b7d3904aee672a126cd66158ec784c6568c0277b17dbe076f6b33be8907e76916e0a0c
z123241585f7e216e8768c27da8e9b9614b63bad17b84c7d283a395c90044e608452898568c39b8
z03e1f1aab22902868c1eb6657ae1d66926143d11d260a5157dac5fd85c16e0db2e13f2b0ce4ba4
z073b280d2b2a8acd39e6dae0e7a774c9c7f3f5154b4d72542232ebdaa5127d6b7f2ef1a258925f
zc7f777ac147c7bb7580bb06fe5c19b048264d17f8ff2ce683273dcb3c7c8a7284f16c88df7d075
z18f8c827a97bd84d74e1c645166e91dd39a1e8ae8ad448499537d48218057ec5135d73eb8b1705
zbeba5c4d13fd47869de255c1d0a4e11b54fc56f8ba3d3ab28bc24f6763a03ae1a449ecdc3ce6e9
z26bfb10cb59323e946cf5c289952fd9a2c202d149ca5b75349cbc5dbcd6aa363ae599662536907
zdb98297e1884a02f5aa6a3720321ca0cae0bc55d5dae672ed0ce621cd9c9d8bd59d50dc42db63e
zbd6943d285245cd0bc3af217dde39c07954cfc2f06d72d4bc77b0748f8785e051930571e9b1c29
z09c4d60fb20a48dd61459dbe64ecce26e9964d235692f1b678e36110a69b737bd762e1a55ba5c7
zfa2e0d43dc0604755f8ca2db2acc49b3a6772b395427df36b1507108b058cbf4cb929cc6157dd9
za92b2b62582ef782b3ccc0cbdde4b2bd8af835217cd369017af8743901f3c7db4e45fde82ae791
z481b410a6c4cfba13a9f94332bc237ceca9f995cc08d2c6a1b280c4beb69f8839644429961e637
z8c9de4544459d0b3b0c97b2fd58479172b9d25b5c9d243c30cc3e295bbed66885974292439cfb4
zfdf7d0783cb5d35089f4cf453fefc70c20e18374654fdf6222ed574327271a18ae2bbe76eaa259
z72a961eac18b40cd313229986212d288d9bb78143ef18b402c63f52f3d34fe5f16037b395ecfa6
z3e13477ae1e83ac054e787175db0df641ac6caba0ce19a2a556a185a6651b913584d4a5b62f19b
z74585992672c1b46689c174619a70161dc192114263b053b93c714217bfa8f91ce86b87061951d
za126c04ffe1c673fa60747e3e1f1d2145386ba90251545b82fddeabaa3e11f994448d2951628a8
zc6e3e466f0f229f681a3a6b1b3c38f6019bc033a3e272373b9e4b2c709953f8f71e503bdccc963
z2e1ccaa9ac71cd53419a3a65e60f4d7d4731477afaae0282cc1ceafc909a7e816a4af6047a74c7
z2c95f6c1d14dad9419634f0ae82a60cfcfa9564075e2f8e2850dc815960946795ebc7c0bee9cd5
zc4325f6992699c7e52adbfc5eab8838ab51fb192fa69ef4ebbddda9d612f3284e4305b5b125495
z5f959f92bd37dd9068ca713a27250ee3e3690a930fb9dc5f6ff22342ef50c0d428553b9b46f5d0
ze5f97b4371969f9119bdad46cc2bea6881afc0c6a46e33dcad57897a35be22f1e51f11030b634f
ze1887984db8d02a20761c0149b42e33de318a4f33d991516898f64ffa06b611bffeba063319731
zf28e61581efca31b7be86b58b1907cd74e53a77859922bfada7a1b37530913f04d51f5f3cf0392
z6a3ef37fc2c38bd2506f0304e276f0650b83c25e4e605e21f570a17f0e531019c867135d1f3779
zd818a5f7c827188f17026ddc31264423c12c596b362deafd82478903d505752c9feceb56f85711
zd90d560b08f6f861b2e85c02093c0185ca8e92a308117e1d35773d39829872d52b3bf735722281
ze92b79f49b071257f1badc667598fc938c4113f482035d63fcb4dd7c864107972362700a3142f1
zf2523426c89a818ecf2be8fc3c72348fb47ad24ff35a479584fb94f49fb3a40ea689a7abcaaa5a
ze8057e42626a82ed8f554d4d56c96ac7c2a9da9043c25848bd70ab4ddb5c3792079a94a342f050
z1f6fc1fade8625f7ef972b55536ef48b944895176e67804875cb7f590e81c8594f01025e833ce7
zd8b70b803dd335374509034dd1f887d82a2c6125c1fde5d06c2e235af242ea8b1b187d28fa8660
zd884c2590909262ecf9399b307a25311a4471cb0822dfcaad5553e3569331f7cef0bf16a414367
z9e174b7f650cc626a6ae114bb0f369406649828dfc7f9c3fe9e22ad4da41dbaa5e061d482258b8
za2082163a5a1293b8b600cc2c66dcd91a8f47e7d4898c3e4c11c31be2b35e608824638bcd89f98
za5ba278d944d7e88cb1c5836071f57f276cd8baf95b4cfd5d06f8119bd5d838d1a902f6ddae16d
z0f56759ec697cabda73c2b7cdc6517293586a19a37080d6ced68c7faf08ad10cdff677be1528ff
zb3bdb8fdf87a49acdc111939771ba34e3ad3d36f5cf294be3683184b7433e6c9d26189e7c4edb6
zec2d9b757b299a585e28960859b88c2f7c1e40b6614aee9b25a910b68044bc3c801d76f5bbfad7
z74308409883b3e1203f40cf800303257aeed01e60aa3a59194a687d12b56f5a1161d903feaaab0
zef581a966d0e2ed15ac24e13bf91032dd9c8241203a7c5a1d8f8cd0e339d1af74a4aed8c631d83
zb27b0cdf108a6550d4a65c27fbc0f7189d0fb45ac24da0c1f5e271645089f45800e6aa956b992b
zf1b4f13ef60f712f2ea22c000fe844df45b2753f1c3c79b4451327a072aa6dad9ffa5c683da2c0
z193798a1a6a508fce1397f20d1ce37ee775eb3b7f8dbff24c394e77ad96ee2170ed595bc7705d3
z97898fca46198d42836dff87115e09518c0f528b29bdfe16640586e47ed045aa1b62d6a42b48c4
z870b81fa34a09b5436e7f184ac16ae936344ea3798c7dddb576a3178e16ce9981db027e3cf9efa
z5e6443c7a9b10596cb48ebf342f3f3fa199e90e5883211acb2e251444947fe7e04b46505600bee
zf6b52c70d5dc690f1beb57afe5a127facc79a841fa8d610b8da89a7ccaa6d2fb37636da517e757
z61acfd4e6464198d2dd3ab4befb239c00e4e4c31fc616b58ce13c5059a0d706fd6dc21037a07a8
zf27307bbee8ba591944c20f25d43ab547550e7bbb8f7bad19748cda86ed7ca16e1d7da0fca7f1a
z7b7fd757948a4031864d58da2f17672e425cc7d2c05020461891ce3f90370877b7756dbeb56437
ze4dc1a7bbca1fd06120e31c1104c2f1936497b9447ca4d397bfdad996c49572bf192ffbf0bc6b2
z6c7d56caf74c5c7d72f862bbad602d919d522973b4d5d317a34a11384e1cef737d251be9991f50
zb00ad79baf0e0dee1fca1fba9616693da74f8b106e729e9d28802e6daa3cdea8b8ecb740287a42
zf326b8a2c4dc8a090240f0a7af604d522b3bf5ad47548c43adec5e2eb8ad10f1da9272c521d8c7
z1d6dcff58bfb2b6ef07f4e57445a6223f51ff3cc192fefea0688cd16965d401fb3aa7be85052f9
zf58e50eba90091662c0ae6e380356ef9da70129233091e6d4d351b0a81bfd8055ea7a4542f50c4
z0e2d7a44d4cd2bfe4cd2448f8f0684bc24005c48ccd72988186e9ed1d18e2769a741c6e39da6f7
z3e852eeeee1b1ebfc213645c78fe60ce2a0b7a732a1867fc96af5aa51fba9bc19e60d6c82c6d8d
z323d28a42a3c52893391609876918d276d59c41ebd6e4c0e2ddc025a428cd2948f9b17c65d3892
z63f1d1d3df10e833138c9083dc8f572bc44e6b55e0dd4afab585c3ba768ea591c95f17ff925115
z1d4058079615931d9eec6898afb6f7014a02cedb7fb27182856e4ffc7849dbc746233df3605d64
z8252fafbb9f0d288027e57960d9a099d8d017d127b3e90258b911244a61de1bb7af23a909807c1
z3ee4645bc12227b6a938897218acfd781661a41f8170a01d0274d52080e68bec4b7de2df24afef
zf5056eac1303f6eae17d06cb5efc97b6d881ac86ea83f4fd35d47f6434c35bddb412bb47ceaab5
z60cd24849c5706f1a05d3585e97daba8918ff139c00a8f341ee509c00b1691e76b27f78fe6cf10
z13d1cc132a32bf75f0c74c1de75ebe80c9835614e6961d1a4b1aac0882c245d81fd6ef32bc00db
zba8c14d46ba9e47c5a831ff7738e39b064ad8fe751703377318ffd346ca680d5fbc8298e445825
z047c68f23fbab6901b776f84dfc564f37a16c9da699c59596fe6c378e123329db9bf13da929dcf
z5abec1de66f2bd51ae0b193d198d48c1fb9a908c3cc29586026ba42404c0065372fd06d92525c1
z53c17788db216ca488915c38b34d8e9922c070717f31047666123f1485aaca24c5e67d0c1d5bf8
z903c48f94d05206536949058b06727558043f545167cbc5c16c7abf60a6e6becada337ba876480
za50c3d9d7bd5462735d4da500f02588aedb40276231db60190071dd879be7595875698a37211f0
zb5ec868b8d58002ab0b90e9da476ab22ca74368759f369e37fa063140cf4791dccd7c70d1cc555
z6731e1fa67c69b1dc481e67c2815e4c06c98809a7abdc30279c5344d51269e7d18a9255516d41c
zd503681cc584da179c296248f49303114c941d4b827cedd56fa32b34cbc3694fbc246bfaa3acc8
z2eebe079ad4d40d3b972f8c879a8dcccf1af6cca5795b16c5db7f415a0bb840622bdeccdfc5218
zadbacd36cb435faf1b32e8abc76f57f997626b922b5b395a34968ae35d29e9f10939245d04cd72
za87c9f4d1fbe842a39907983d87a3eb8087d18645a600cd79536d3afe66f8b730554de13e3f8bb
zff09c215b4d701bb74a28dba1ba7b004b949f435655a523568fa75081a8892ac98efe61e162ada
zc9c6ea476576f41477bef85f955b1eb33660f9e9af08befc86cfd518ae1042a85a70cbfc3e9caf
za8d27a29894aa0c21a94fa34a4145f72a2aca7945a77d6d344e89f24688076eaff286bf69a562b
z23b0a88d4fd6e28ada3bdd1b7949d147772adc7af68bd5ae8422ec739368998b5a5aeafc406a1c
z9ea19fc99e51a2e21cc4b11fbb2e81ce1bac39ae73a531874356062476965da6230ff141de172d
z9363b3d47d87c15b6a53a9a675b085483c23b8b6bcd31d96a82f4d3c9a66329c84962b737a58e3
z224ebf5e01fdc2c8f9579dfd86d10841415cec9f3ea356515c169a115bbf83faafe0af846a647c
zaf3fe60a80796a4c962be935071616c25e70b79620416ce14deb7d47122badf17876b75242cca5
z6e10e06aaf0e03aabb925d2f8d655150bbb0524a5c85cc247f8da0237d82eb183fd4aaffcae99d
zebb9e993a92c4f345eee765db384fdafdb488d0d5776cf0d58a142e14c5571b74c020cd9ff0408
z77754ce04140e6152ff0d10f4531029c19da92ffae08e47f8154ae1553f2e417211364ec9539a6
z9ce42780fdbaa400ac09e49417d0e1f46fc3e18fc0bd335031191bb8eee293a5826b386a451677
zdbfbfb8af8ac1b8ab48f4d76f69c73abd135909f126c73fa5c715e6d5e893dc4ff526cd7814f47
z51995dd07ca4daa3f224502fdaf37cb779cec3b2dcdbe3b48b42ed64db9b603257345e357c3759
z9306db4a90bc84dd8836b2ed30264c43112d5a029f42a7076e6930b289a4bbfe6843a3e04c488a
z463b6571a7f1b551572adb5f0e6da9e1a3ae8659c1611c45bfa18f22c05736a74ed429db799897
zcbebe3ca7df2f572910237336ad1b596de814644c1ab35e570e4c7647245e3f6fc0225276dacc4
z25037df60b37fc4464354a66aea33ec8b251ec4a4659aa49ef2f521d419a1054e3ef5be6f17ec5
zae55b4f18bc1608bc86e83f5dec7c09a576dab409c84287e6b990a96dfc21d823dea30ff57c7f2
zd09b8a5d699411c6e8a5ca89da572035a3fa95bec742f00ad91497150c464424e71be08322db99
z8552831d849a60f9648222fe81da577d246aa2e18be439dbadaade0c3fc976b1e68432504e19fe
zfcd0a8e44567c2abb1effceb122bd1a3e6c5b3e01ec339869965c58622b2c2b11d3095d48a2538
z64e30709ddea95b1f0e42c1550b7625ed8a2111cc2d7fd0040e59a086f4741ac12f5d287260dc4
z28a84f3894fa5afa92a2dc4a08547a153eb45e23560c2347d9531b3ce995802a4766393f09b938
zfdaf3b87a29371e69839e2b4a1fd1c2ee807e0d0dbbd84d6a56ecb4bba0e7f3c16ca7079da76e6
z0a0f06e8ac57093024cce16496d22fb622b3a0c434f1ba9bc26e82134740b25d1d88fe2e55250f
zecee341111e5fe50df26e153ab8620ca1165b3754e39ac4dbaf49b2f44d895b9d32bd7a135a647
z24138841bf331d958829162bd7e26fa58d967fcc168bb7c97305a81ba8d4e78349f6d4f1abef5f
zced777d47506437bf0d22f45baaeb1c9fb23740d95c9d72db50bc805cfa932db76833cf573c750
z7512a737543a61bfe96bca8be225969c342da3f81cef391ac2d6f76e3d64622840e9e33f042306
z8149bd6d50e3bd0726978197cb4a38b3205b3d31ef322993edff4b86be418af3891864e3e4f360
z6a48ab4a9203dc55f8c950728b25a010549a216b1e342499f9832adc89060ece5f1d6995a4651e
z5f85c15048cd5dcc6ae98ab362b21521ca483aed63745101434757c690cdb3fc15fcf9db18a912
z94be89383d33217a7d3e2a4c4819f983eff20d4f3df239b650344506df447386cd33c8d06b948f
z781f1bcca133dc0f13a307288dea85964f4e7b851a520418b41cff58419bf1b3f0e7a6cf89d286
zaca397d0a656968a12cfc8cac8a30a37ccd4c5f6aa863636172e992ab74e5ce56af1ab4542d719
z20f644e8604fc305c0bd540a624e79faec0e95266dd5bd964f36547685bdb20d035acadb9f2dfe
zd479a17cd5a5816e0eecebb8d6624608451cc38ca302f1fa08e5193fc92be2020e236a9cd416da
z68e0ddd3c98d745c50af396105bcc8d0555c05e4b2e633d7c36c9c3aa3dfe51c6fe55e63a57fdc
z979a0026f0afe714d116fff8be5d3969e960f7ce41756af837265f49dea8774992c9275ae994e3
z8af312b0205770d2a19d224c88dd0481fc34eb4fb261d2f7e99f52beb05efda60b82f2f66426ca
zfe91da8c79f55af19ff4e7f542cb88b5c4281ddd02f9bc814f9eb22870e8c3756e3bb6c1fca1e3
zc622f98117d867522fbfa593856b6a702a22b4ddf552510dfa56043ddaeadcda762d1ddb220ddf
zca7d8bb85abd9a032bff9422f5dd6472f192f2ac3cb5912f1ba9f11d953f5aab04762c89ac9981
zed3dab56c34c2257421dd63acff77e0982412d686fb8738c7c4abb6a52c368fa5791e32c53cbdc
z36ab68327f3852b58c4d96818f6150df904055413aad95bfcac6b3c00534410a5013158a2977d2
z2ca803c0ea30a3eea23e2ad4ab87eec0a33ab58c9d2bddf4c95de6cdfe4daafaa3b41c3676f7a4
zc4bcccec1b787803bb79fccdf9d6e744f5daeb74cbeda6670bb4550b0510d65b61f20f4b456726
z15b9126f5abcb814c0c42bedab558bfa0668a2f542ee50d2c862ad8b5e871618ebceff20779823
za14d7ff0836739437d550078394948e0745522d17bfc161fa16ba93755388e0f988da7a85a12eb
z46a41f150ee1194de424cd3c728f9f4361a3e9b3f582bb18a8e641f89ad2ea1055fd36ec77b6f0
z81e3e5d03de1b961aefe437454695baf383593f1ae615227c8bca563d9e4cfdecea9ed17e99400
z4c074adecbd16c219335674da3e384dbb6695ea9e18de895df724d97f48fe5674da5028a46448a
zb2f75b879bb1d19fa8ea41fbbf9fa36b775efe3087ddfd185aa3c18461bf4ab69f2e9060eb4e8d
za1b9d8b7899ddca57a183bdae186512065b0a83c8e5573afda40f512b90c1ac39efec034ef2232
z79441675cf04bc1733bef4e52b150ccff464b5759f5d0f9aacf159466528a0a059877cead66527
zc20dcaa6c054a2e7ba88d4e2752db66e08b8f09d591f2987fb2ec534a8b999c789deaac32b75cb
zc9eaaa6cd5672bb890c0f86fdf95341f96991d3ebf426c70579effa5af6f3df00411fa4bcd9d77
z84eaa9c49af629bc013e91f3d53809bde495eee343e206d0dbdbdfc1477156d4e3c2eb4d762c54
za83670fdd7393c695dbd0956d0b1a73bc020c5ca95577490b960ea4308b44f2aa1bffbf2fee50f
z64d5094f51d2eb105d08909677fa41e57c5ef7a887f1edf1ef14ac44c8a52602e5d5e6055be479
zf1358176eb0c67613439f86d2d7f19fb6c772c4e9c4eb8636d310ae87c15c8d37dc16fade6a0d7
z933d5964255406d236cc4230dbc560d78633c9809b5a3fd0087a3e27877294a61beb69c0c45fd3
z559a4825f9f78ade1aa8ae749926f68d6a91b6f1da925e774a53baa275f256eb2eb7c6dc53faa6
z64ee18650f9d06d0fbbe414dbfe521570e7d8029cbbd7fc0b4e758cac30f21dfcbba91034a6f6c
z2144df96dfabe51d26b81d9124653660c5ed1ef421364f3110a4f10b4117c841b5131284abad28
z7d3380bf3957dba9b6f5a22b403d6c15e0a5a4d4d371509a2ebe9d7eb49989b7b12daab962b89d
ze9d70b404fb6e59d2efcf280d81f5aa008585bce19760fa0cbc92a5dc45d8ff5f5b8dc33ec2443
ze99f870d5564bde14a61e8040e21bffd384258a1d0c733b8f169eb20d6f98cd02e07a4889ea8c6
z8b4b694356eccd7da690d173a9890e35143a83566c8fec7b1e59416f9016abb03fc040b06730cd
z5edb3b78fbf741046eb356a5045e15399e0b8b0b60dbf4bac98c4e6ce7e994fd7022ac1403002e
z378aaea955fe96366637b9d04739f51bd60070bc99d31fc1aa71d636aa14077aadbf0e39b0b15b
z7d7ad34524127f3c249a1027b7fa4d6ab2e96cdc3f6d80dd44c54b5aa4c07f315d6edbfdd02810
zb5919c89ac7d9dc834731dd2a9f4ef945b36e811750f97f2fde47fed4a2dcb65782c61b4aa0d58
z9173035fc627c0fb29b109b115160a6c87094ae7d8e787d7bb92ee59ad0241558ac1e0f9ecb325
zecc47a4460b31c774ac9444a9f1954238bc9b6e5a09d30dab02e1b3155473f7ef766d2b11475db
z85e7aec31383caecc7998eb027ae715a85956b2f30c5725466a5013287cfe1f906485395b117d6
zd24614290fa6a0bd41fa8bd06919630986b0604b4d0a21ca608553fa340a581288cbaaa95e9709
z9d227266d8660a80a0c21e237f08f6c7ca1f142af22a4c1a8bbd11f1ceee1c96ffd7d035f8cfc3
za30938bb9463e9d87f59f1a416b56625ad1434243862f9fb108e9eec15e21b3256ac7c3da68813
zcd0d4a9c1c0ea3628e8ed1a0ba4556fa4f52001fb73633a444430dd41f2a3ffdc70a62cc7cfb4d
z8f53082e84dc69e13c51c0a4d38019cbc50ffbd26125ad0a14a2e2879c93f66b3d4ca9f406e70c
ze0b00bffaf41620bb41d9eb618a285145446385747a848bfe115259e0fb79c59811673b7c4a10c
z48cc83a5cb2e836e92926ed163c0f17019d642c4cdcd1ff376efa50b8b3ecd7578a3ddae5d0e59
zd676732c57738500dac8ade64abc0fe9018ccf4b64403326d68a280402d4a5809c37ab26d35fce
zd05d1daf984ed1ac1cd1dc0ae29375b17e411fb9d594cd8b3f7e04e66896e719331d476702f11c
zb396bbb9051436aff80aadcc0f51e883435ab660b3967b1ba286f4b8e1da3ab90bcd2f78e474bd
z2d1a05ee95ac2167d72a3981f79fde629c81da3121c7e9f5a586245fc68099b3d20afac6222de0
zcaf40825a2877371b8525876d8a937f8fbfb01a98d9b12f8bf085fe09d7388588fe746c4da8d05
za533721b69f3106ec3227058c973370ee9cddef09d6cd8bb2be9999282d82afe7a58c58a915194
zf9843bcd5da2e21fd8fb5add249e176219e674be6a31b891f616adbd9b6449f1ab942da4f1cea2
zba35f542cfefd2d5c8a666ff3f31c660e6891bc4e6e3dd4a6927c1b2f904992535280f8de43f5c
z35679338e5af6a1835a0ae8f01c5b66e6e5c52f8a60b3d876dd75db6ced213c1e8755000130490
z5783ecb823a1b5e8b80ae68aa0874759d57bf1b9efcb2b439ecc4dbfc0a08104b9d0d44e227c93
z2ab90ae9efea679b4645783fee35f294a1d1db5b0b5d0aaf9b9492903241c8bb8cdfaebb40a66a
z78057a365262e505b797476e499140417575751dae8bdcfcd8b19e0ec21ee969a1ce84a71abdef
z77961424bd0e350ebf70c264e2391ccd15af6e718937b24ccd7cdcedfa5b06a50cf7699cf48ba6
z5672f55aec8447dffd70f5a9a23dcb8d72a49315bcaf9489d606fc5d578fa4219f3c239140c45f
za1690f0470d7598cc098dcceeef99e0b71ddfb5bf7c82bab0f55b10c1407c89bdd4dd6ba0f5edd
zc447eb46d3c95549ad73e9a3914b1debaaec52574db8255440504b85a9664df147f928dce5dfb7
z7fa56b96c5613276fb510042bb2985bdd9d968e54d1fae75d683300f80c3b0a5629f16e3709648
z79c86b12ff905d7aaed2a527df0697ddae6e5d95136c91e5b7637e89c2c6d0799f4a217fc4e145
z3710991f9a882cf00bc3308127c5a1908bff6d5ee6bd4cf972f985fc5ec8d3c097bc1947002797
zcd5182c1950a9a1a7f103e4aa751102ec6911eb716ce75602ad7799e1d65bc6ef457b911f61c91
z302ee252537b1d5aab93cf11e372016319d35d5c26461d7c2c2f00d3dfa8d5a0e289522f0b5909
z9128fc1b4b2a3a13a4f3ab24a6748190a080cec98d37fc01b0aacec9cfec070dfa7263f08c74a5
z3d263480123a9fc2dbecd0f59f59eec6925c1d4303e7cd8d989989f00ee1265d892b5ec0be526d
z34051578222bec498dc0aa3c723e747b21a431e18f5141b064dff36ca39e36f82577c65859e904
zb22e7d6c7f48b53575e4dfcafb12b00a28f20b4dd5487129608431c442eb733fe270fb76688f88
z0263997dba227934db0d349ef9d83e841f776b34f93442f1199450a5e1c2bd5031e6662d549dc4
zd3bf726b47ba057402ad91c0708aedb4963eac4acd775c4aa6ec25bd1c4f822f75c49da21253a0
z9c88db8f7c5621aa8c7f4875f20ae17076287faa4bb7e95c0fe84a08ffea1c0576eeace62e6d96
z9da6449e65482118cc641d79fe2aacda8e19c9095ab66cd3c4254ad3a81ed09ec58fa68487b3cf
z76989e65ab8c54ca9645b23ed7a4b757ab11a65f0905861862cf7b1eb96834e9ac9e5914286b9c
za9b867182f92e5da2e104ef7f2965cd5c06c8653eb8435108796a289369c7549b12af5c681ccbd
z063b57ad68237d9960e996b371a405232134c49a44845fed886fffac7dddfd6d24c103c7e3fb14
zdc41e1938989c0ca1cadbcc98a788cc1da941b8902bd6bf67fb05231a78b9b395e08c42f53b3ad
z6493cd2714f9376c69976201e2e90d1ed65c9f59064fade12503ec8cccbd12773a93c1318991b2
zce3bb750f8970ad7546edb37b8d805cb31f1392a579e52c7b94df33103870b3a99c5c744bdcf6f
z6b8650bf750354b19405891156a945c1f821a03d145be79130c14f91f1a2a81cdd98a088486f86
zb0fb9f253556f6e318e01f11f2a023d37e6bce7b9f6d5f61119e71eb81edd646ed24c7a73ce06a
zfbbc4f5119f3cc83d7d7c41b06fc737b41bbc4f1602dd9d164cd6f2435da0736194ec524abcee2
zfa77b53aa277ffc08e28862d6555cd927824445fd531407f972faddcdd8081c90e9735f798a65f
z4338363c8fab307cfd2d121c39fec35414df036f551dde0fca9033b56c2adb8364374e8654afe2
z7f778776898d0b697f22c03c341087e42498037c7c17ca95c65c9e27c7c2dc2f7844eae5c1d960
z66ac7270cfa208b5e1bb6a2a3671173cf51df63a2b3ecc4c7e1f80ae0e09d5eb09e701bc4ed384
z3046fa850fccbc69629b3b5ed7fbd0eb7031bb97e65aaf44af0fc80fa59729d930be26b67809dc
z6d3839e107077334263f1a7a64bf688a3ee4ea698d3086c8b83fb501695a1dcfea82a7d3655fbf
zb99cee960cc1b1a4c6fd7fb2be160db48de2e7e76577bbd813ff71c793740e8e550dc5e8bfbe6c
z600a8117f61d0a00892eb5fcd0c8b457a064375555828a9cb9e0dbd6dde6f5b8a42b04fed01c60
z8f7c5d9876b8f12a8c06a0a443cf078c370662c0599b6c2af9653152289a82aa3236343c259eec
zadf6b78e4db8744df49551b411f14734f7a537c1837f56fafc08d814d78b57b132fee25f96e792
z962e6aabfc623a065092b4bc2dcbda6f37a95eb4e9862154c901561721f2e8605736efc64fc5a6
ze819624c7c1284787ea32a833e49ca20863003d3ab172a83d171b89197c7e43bfc6d96e4d5ddb5
z420a86ecd1e617ac2676fc5d224829f0652086766e68a886322ddf8734503403a5b3a2b81295f0
z90bb61ae77e21b531c8077f2517519ed941a951923f0c58715c3146c4e79c2d918636ef7b6e47f
z9c43f477b47fb8faffb87a01944bb49a0643abe3de9d885b9ad09fcf1677e3870e7223fecacf4a
zd2090cbec8ea88e121110112edf80818e9b2d026c8d4eae6254f25e7e330c1e505898ff46afc69
zff0a34dd6229ae7520c883cbd74de407e777165fafb9a582b3b49bec22b6a43bad4fb33ba1e49f
z6161c762e988ce691be462ab19bfbe881b6477160349a79386507e152875f2a0e183bbb9eed39f
z26e3ded672c2005078cc3f26878a496bfad1efa60d4294e163d9c48fde8c849cbae9a97ab6ea78
zfa9c6db92630c43189a821fa54d12989f61e28db4303c4776a54c850a857e724b43c7bd60deceb
z4235b163f5c6ff440ad58f21f4e1e332b4c1e5c3b9c8dd26b66f7068e628d692e8b14938a828c3
za35459b5963e78183d08486442c17d4590d61b54c1a0eb67fb992b9fc15609316dd31d0f9980ef
z8f147c4e29ab66ea361c288b9a01b5be7bc34bb72736d56903aff4a834c953e335f96d92fe90d2
z45e75c38a4aec2486721992799009e044bb89c03d22252596cce28ea36631d25970252dea5475c
zdf3a4a6aa36779adee289ae2cd3d90d05bd6ef7d3d14f48b13da5cd33f251bbb13886c23f0e4aa
z00bf0f8ffbbf26e1f5d66388f3d0703f40d43933741e1d40312cf5253affd1428246b85df695d1
z54979c5f2ec2be5b664ee0cd9ac6786fa86295fc0e988de8f0917d57ea1b820f2813aab209c04d
z7d4126aa33323e2cfaadaaa7589b7701768f5235228e907cc2a8c779578118cdeb2d0cb6f34fb0
zd50fd30b8fb7ded9dd1cfeda4734dc55d4c7d684c2de2aca3c5677a7db85339d86b85f8a3d6b0e
z2fb78711a246537c361c15c96b5133c74178ec3c4612d060b3e51e0064c42b1315020d44214cfc
z1b5c7f4fbdb78e35d0dc48a9a89dc7155218a9b427ede3822e57c222704044f7094eaf8e9b6315
z22062a19f1f8c20fb06fc81dba3e09b0cc17b77bd21857eeaf7dc2c254eef805486d23f1787534
z3419b2f672ca3e1fe62c0f466285ba3ee02418c06c1ffe7bbb5c779d43755f6d7a88d36c2c0d32
z53c40e647b606e41850b45a51f57e78de1f0b06a07c20a14fdfccb49e519590e462bbd2faaeecd
zfefa5577b88bf3d34581ef61841b525bbd117acc4cdb60e20fc1cde9303d8a91ab6d536602d224
zbcc1f17744fc2d40c5d0ddc062a959aeab4e22a36a35b37c74e5118ffdbcdbdb7eb6042bd42f07
ze55aeb09836294c12d35e4cff44d81cc445e4544802f8fe1263eb41ab4d343fb1af55a42d7c2da
z4ed8f58a61a99b356f02d6f89df94226788f9b80eb92ea788a4bd910a3b25e62c063254fc9d555
z8b21ac90429bf2e289a785b3f8609742bd3ca2bff12a317116e78da1ef6f708cc43b622bc3608d
zd5358a40a9bdd7b492dbdbdefab5c14df29e6eeb250ccf98ea9338176e9a842de62009252a4b83
z72d4e7e690216edcd854d6093e391e8aee42dc15fd36d355de78cae1e513ad7ae4642f93f83442
z9edae45d2dbf86cb5c6915144a677afcd08e41f48bf44e6ce675743466db955fd0c864eed11372
z1957f0213fea666fa4c1182c8804359b62d88c0cad772b990a61dce26fe1c9aebe2ccffe75aeac
z9fd17795d68550dd30f973b6ede5608e0403f06ab5d7117c8b5b7f0a2697064049e200eeccfed7
z50ebba17ca3861160950630496e5fa0762000a343f92e354ce4148d952138e3f36a10552bd5caf
zb333af2a4040b3073f252a2f9b2afe6af1e20a4686fde5a755b9c411e6ac91a1f05c7726353b44
ze1c6ed69df7866f96641c06012ec97a98a96ab36b62095617888a4c129cd0edfe7e45c973ac645
zc731d6001c583fef29d21a7ca1576bfa97fe39f81c6b19cd674d351dcffe362d7d1d00b056dc4a
zbdb3fe8bd5b4ef4f0037e124c2076fd304f2d679c1109d8041f01066c6fa2c42b69c96be97c8c0
z155bcea4160e6efc56ebf8454888083185c3f934854e411be065fd13324684126bd3ab0200bbf1
z36e3a517b0344cb23ebd656556f41c6a20d3e8a76d4831127047b4c8ea94ebd1300bac896cab33
z2f513bcc8b13441d5c563bf19b85eb94b27a93fd811fa1bd5359b10f1337a464336ad834541f19
z30611a446fbbe5324797331078d19350cbb5782e2c2360dd64b431025d3852fa9094c2b6397f9f
z16efb7d14faae09d80d4eec9001868e5da92b044a1099950dc5b7c9c8f43f0fa8dce44cb995a7e
zb78a88c0cd561b7ca7f64d003480689cac7e3b34ea8bd46ddc5ddc0e05c6d04ed592f6735067b3
z29fc319eaa238c7013539ebe13bc11133a7411c3c7373131e73b8f051eef469f1f8fa5f56e2e16
zfecf2b014e4a0890d75b6c8e9dc0900009c23aa9f194a9f31ee91e33c3ee403f9e54f2db4a1668
z8c28a9114f2395070c4d1493cfb3e455f75c8a731011010d33e176692234476990536f206444ac
z46a31876310b3a8cc1254c047d0fedd8ada6179da84ede6c30b46f90163b5e51c48ffabf1d21ef
z0d6cc2505933dd83a0dc736def938ccef4f22fb6e861c96ba1b504b0dba97cfa75ddf0cd66c6f5
z0f737ba8cf754b60d96d316c1e44ea59291bba8be0221bc09d0ff04b5eb40c897e404cc2c7134c
z2164f64495ef4191e89e3e7874f970d7c3c20f77c13a2557984364e72d0b877e93247bf0aff85c
z74c89ee5c4299ad34b0cd04e266ae79a19d1d40891debd7d9e1ee85d46f742fbad7d8c2f6030c3
z54c874a6262541688e4027cf16101aa073bc65dee619a9a5ff539446365bcb02500085ffd821bf
zc62a6238cdeff8a0f27f8337bcb05927e3959e238fc226e4b5760b92a78ec3423b6a7ac42e2543
z8019a321afe3c748f469b544101c58077bb2826a783b8e05f3c05406fa48e922a4267319a016ac
za0068a55b6e277d3bfa8353e61f430d808c2651cf777a2e47110fc8fcc3b152300969d257fa83e
zf281036cfb5c038674f99747c175c37e7e73bcbd9f96a8b0900108480c3e5655e8be26e435c7e2
zaf59c5a067492fc2363a78d3ab087b5462338ee00423a5d2214e78c49bd885760726bbe0969738
zd5cdfbb03559eec162fa16eb46d0d03e8f3f5445911ed51ea436a16707eeff6705cd01e30dddb0
z999b98df850419eb81b7b9d86a6c1f4e1c5fc52effbb0951d56c3d38cde23b2bde5cfafa9469ea
z82d1f0f64ead25e3ddcdb5733b4065f8d2d5deb5906f3a05bf42ba7c6d02f9ba989ce099a4deae
zce31a8e8b85742733801228120154f11b581249c2075739e45d21b083f0d3672847ef4f704a675
z797a8bb8f4976e0a16f3bed65d1c212580a3ed627984ef85d6cd59b9e2df6e02f07353be74a097
z6d360f7e4b1d3b50ef4c19a44f8b12942c05f64091d3c491c7a08dd586a4dcc725689833c2052a
z0ae3569ac93b0772683ce71cd5068e28aa2a95eb2c2546c85af9fb958d97f390682145ad13ccfc
zf193c5acbb3460da2aae6b4299506faedea00203e402f6c56aaddd0ef5d90744786f3b0b890c64
za0e0e0cb54a86f1b49e2015234a56dcacdebd87473d9661765f791149c1d7e427531109eea539d
z58ba41f76f6685c0edc758e726e3732e89f17cd546b25283fc942f41cea1409286197fae57586d
z6b0c9903453b06061370e126b5ab01a45fcc063e58d3b14a02a709a321a671283caa8da8c0d3b9
z5e08c0c3e57a19c1461b30acefbd0974c1b58aa19a27581980d16e284b2730d377c10d50996f05
zf960c25fe3061e0474175c66d44dadc5d4e4a6b3c7df21d55c72a1f37666e47dc76fe8f0d48be5
z8fccf55784fd4e4c2c5451cf5c8fffc8054398d9a4ac439e3ea9e76348897da9cff4708ba9a4b2
z5d7e0009f2d0082710d5cd8cf16552c060338ccf7a2bd4725ea09a9b9246212a69a5866252d56d
z53b6587b1616edfb915a5ecd39da2a66b603ff67d989f844ba6dd7cdde150af24ae698d8148dcf
z54762567558b71c605085e61b9efb9b7c9badcca77d8cc0687b1c852965755a14a6183e7c7b592
zfdaa4cfce8d0c7baf7867807223cc05e1241283f9db2ae47e730a153380faabfac0058255eee45
z2f5cfcd30788601a5d5c9b1a4f2f7d78e8bbaafbca533b6a7ce6b7f3bfd5a3f48b6b3b2d4ec70d
z003b828283300ac4c8285b1e51ccca97dee1890488ca9b4820c591fe9ad2587bfd1fcd0378c172
zf68bb91765838eee01fef06be9cebf054d4270e9a2dc69061cfa24970cc42798eff22292e9e0bc
z3c0aba4eb0ef0dec5a70e0edf22395eb963e473347275a4bc6a6729248d57631ef3c22f25dca64
z46bd042b0805703b67a0c15d6e4bd09254a1ea763cbe22557ef459ae3822a3d89f44e97e24741e
z70b745afe2ccd25381d946758063a1bfccf54497b2d8e7c72e04911181c976916512565e179a3f
z3e13a0d86fb28ceb87a8c23708185fd94d5daaf84abbc2754a43830e82cde2b3aef2d7e89869b5
z1b28463dc004e87b53696e667052054cd31f9527c08572b09c71a30972cd1009d9ce3d47d06799
zda620ab6a17fe17b2ebfc5f83e603d4591e3bf31e55e86d49a4652ed8418a330ec74b9b1157abf
za74d360c197ba90adccb858ce552d6b54b7c6e67521de2396a3385f7b34de3b174a03ce204b718
z307a44311dd7f09a2fad163fdbcebda3f362c6e2dd88709ac8fa3ebb5fd6e97b43a89c6f858c2d
z77dd631c45309abfe587ff1090dbfc583eb22a865d22c239701c63dd7f674b565112e69df022a7
z1d3be65395216eacf164715089d8667cbd487852491f2a856f6119883a872c1addb9c1229844d3
z0b86d4cdb164e4df720cfed81718489cdd80509f515bc5c20fad5635eda3c7789b73a65c032a76
z17530cea618634b24e94e2c68aa6833ff1c62dff943a491f6318c72d3a64ce35cb2433f130be5b
ze1b52b8e07387c4d7c45450aa7fe105ad737202764619e49c2bd9cee55eec49f78a6f70742206d
zc9c074eec0048dbe39509807d5206a4758b0ee1ea81f6b8b312c5233bcb65ae1e8d82b7a8aa25b
zf7bb862c64d450456cf0339e4805cec9a51952b5e99f3efcaafb526fbdc4207ba00b2f12f87b0c
z1d78ec5ecf0834334d1348ed0fa434aca3970edff877c411e71dec6a3a7133bd1f939f53c9c3f5
z27272f49bbae7b1c234cedc4a54c55d02f20d2573418c2d82a11f684ce50850060a8301b00921c
ze6292c0d2dee9c490f5fe79d7e406294714e5ac8808951ee3933d94a7e518ebf321a371e57c19e
z939f1d59152bba031ad21fa0c1b9d65390e588dc050f3f3145760c960c9644f5a4941f892067df
z483e46ce13dbd3928823aca404f63f9f13938134dd6a999b537855d43058d9ae3d62d8a5f1834c
zd115cb34b528a71967bf482fc18e041967907451e95c9af5697c54088e4e9c01bd1c4e236830da
z1ab823a5f420be981cbf463694672e9374b550174a596332c6181623fc786208b88ab05504124e
z319deb0c61a4f4abd3537ddd90d13db36efcdd0e15e6a215cc724e8768475101f10e6e42227a61
z0ea7e24cbd3b9648fb4b3e20dda03501758ca375c596645d6d377da8a36f2f3406aca7e0037479
z8533c55ede00fbdf5551bb6ae65fad10747906667466d53f8131dac8f7b88067a67e2a22af33a4
z0424755384231a83ee0b38284e973fd18ac0c55f9e2ee56572a27fcb7fa4fa1f5a91e89b96f0df
zbfd8154c57dd945d802f4be41eb406d740e3ca09575f79bfd52eb11d20406a73f2f962eb36c3e8
z33cc36a8294c1d06ef71acae69d55b3b3d40a7c5ba6da1ee26f935872680e5a294370f94864eff
z158a1ef59588e1986b5d978f8b16af478a509ead220da6cd78ed9ecb5684ae67e6345c828f1691
z4b896bcd833a7a25cda76c7fe4b96aa98972c078e72c5c1efe54ba2da19518ce9f48965dd3dfbc
za8bb9cf2f472c3a8a7559c372ba7f2ecfecdebadc75bbd1eef9b2065ed593f86e1148662c3a95c
zc301141cb000532cc0b0ddf5e7ccf5c20e521174a0a560c5d789aa4974e350b86828a07fe58d33
zec6cae313a46a7b7e05b797eb641f1f27fc45c3457a6a503670bbc58665793a54696174786312f
z620433c193e9c141bdfe35a80533892c7a6e1ac00e8f302d475baa1e5fd7c51a64a9a1f598a9cb
z98b8d7009bb18102860984ff615f772405638d37d80897ce48250b29fe298d8d5c2ffe672f8c4e
za29ff369e28dbcee0a5e10bdaaaccd361078dc229d018fc50be7f5a50f8473c945640576f48ddd
za28f4c3849be9819dd390363730529081312389eba193928574099a872a6a97f097588b930ee66
z60a251d6be540eff368f0f6fa05b0bd854fb4195f11fa9546d1106518b2fe4138f14ff5482c80d
z65ef9a7987fc237c8f932c7a63068baa1fdfb68fb0c4eb8102fbe4a5ce6f2a2a27ab6b69c5b4cf
zf5b55a59bba6ca4bfb0095daaadd86aed33e87b8ddc3d1e721d304344470a7130b91b2e11beda6
z236cc9bf6bd814d721042ab87a9e197f15e1238e2ec3e999d552b7a3524fdc6be268896c8acd66
z2d70a4dec3cd9d813df00d84574d2fbd4a3a3319dad3da81871b9fcefd865182d778cd555a57c5
z45252032d612b87f70161f1cb8f79c1d81b74bd19714243b0c4672440c66d1fcbe2f59d617edb3
zfd4fa8ddcba2bf4a135a116260e2f1df7f85dd2bd4efc36830b0349624f89f933c81f3da3e909c
z224b8c3cd891623fdb48c4d783d3647aedd139d607294c86f6922d14fcdf38b0c5f90a739f99d8
z05263dc9c24be1919e16887d930e0127ea6110e4d4d751a64157c5c9667a8e68d937655cd6dfda
z1f882940482ac4427a0472d437ffaff51e1c0e24af2c09f826f35f9d4b73f0718d00d41d92ed44
z73bdd3b7f42242e30db6b22f75905fe63426f4ef37178619c0d378bb61bd5363431cf200d92413
z877a68c1d529a270ec37ff78c265aadaaf920321a1ccee596e0ed16915549c432e8ed66c0c0b5d
z62995cc97c83f07ca5fad06218d28cd23f21413a33325f593567df8c337a3258b71f3453dbee18
zc0d859c40f7ff5e99a2a99d1ededb8d2661c9869b2ecae6098d5472d800f3acfd2a610d077a6ba
zad351b4fe2d56735d3dee3d04ccc6af2c21a956f06fac5a59291554874ddc0565c79e8425ce2fb
zbed6b4cd641ed3c535688139cb67f54d7d6999d06da11ad1ec1339a57ad595b2053542cd2094e9
zddad419e59cee62dc60144fab58075cbebd7a845b3e873ed181898ad45ffce6ba791fe405695ea
z17f1828da2d53abfe9cfe576a42c247adf7aa37c2597d140ccdfb6dd976140f42d88527f338c41
zcf71250fbed7a6daf260b8b986dd4889fc6656aa5d8f2e70c35dbebf592825f1dfc69b9fd4abd6
z0c33db493476e47e3e6765adf1eec75d77e5ca9e4d6d0ebe154cc200f1a6c77d1149b1ae99b3dc
z6253a65e80a6987825e6aae8c523336c892502b0b0138db1b64856d813094250e698d13af76e06
z75bd46b4c1df242487088a0b69d4a95066ed3b58bc4c6fbde55d7d1e7425e0bf5fb70ca429b049
z4951c3710d6215a4734a8c3cf7ad8a522635826a5f35b2d894b5eb9a0b970a24ff84521a3cafe5
z6214369dfb8ebfea6fa86d432233f4acd129c7cedb35a00fca2e8a46c7ad3aa0569d1271250464
z5123005b0227ecddcd906a8c7ea939e193615ab8f3e7cc2af0126db60e1ea34bd73df285321e96
z3436871353e521ef30a27820fdd854d1f03c6c8e5006c181098d9a73c29388ec36dde50b0dc433
z76f7c2b93bf28d1742a2c38263e094d378c5305738a9bc16f4bb8d0d55cb8c8f33fa32853428db
zc5c3b81a98df73a43cbf7b819427ec2d0ae259732335de7a8159facdff79ad94db7268600cc571
zd85420c0fca56c2580a64703313e338d11b21a3aafa5a51778d9ed95b15dd5233edce364795d94
z9a400284fd2e11c7fd48f45ecc927c2512b0cb8329aa231b794b6e466938ec7fca1276dd679369
z18775c650fb72a7e353673cb388b13a36d6d4589fc177e9700122a3b7f9cb8c9f7770428d32059
zdf135748c83e55e23c7762bab421e9f836050d9a7aa5f5e005ad1e55ee4cffe3321f23387088b9
z7eac18374f76faf197c2a472fc1f5225927fe4d52c69e31349b2c354edc6ed931d31d2fba7a38e
z2ecdf45caa92f97e0257bdaeb7327474a7deccd1e4f7c1f4ab2d35c46a539df9e4d7c83cbe1202
zf67b268386928f2c0283a939640f9c5adf4b21eccafd233450173d71a195b05d93f70ab1a2b37d
z02f710737a050fdfac71c2cc9a73f78b7a62fab514ec8cbe49c0aeb8c6465d25fd8c941bff2431
zb8c66fbe610eed1ab9420a03cf7cf13a343bff1be7822f3b0cb01cb8c606b77579ff288e79886a
z15862d887d1d7eb83095bb6d704c1ea985714bc41c67ae9166b4d21dd2e75b8d4a5d692311ca07
z9e2e6e1a7c071e28b4050e8815fb944e71e30459638be29f402f8fa14ee52b4764a1b9f0e937bc
zeaed6b84022f3452a0b5119d3f723e397cb6cfee59fb0b058d5cb4cc0ffbd6b21e172d74599e96
zfd8836ff70344bbbc7ac75b0c51f228addf515b0fc9b4b81910e321c0565e533d0b4c6c16384f1
z25bce065f8ed14e387f4908a9da34fdd533e63b53e16667ea19273cf1bae62dca5cc5eee1a26f8
z5871b1c2d8494dbd5fa1cef44df48727c038f367c2a31d877b431f4895b5cac5f5dac7ea520067
zcd4f5d8b6e436fd30c2ad269685bc3e43d7a434d335daeb968ddf64545c4f9dc824311d80b2b4d
z23543e4d4fb393caa24e19a0e90442adc3437f53c94cc810388095d8cd7a53e2d85183a4df8361
zc36409b252edfe0ccbf84689a780c3e67fb54f71aa6ee12af6e8b9d63bec34d143fc47b8985e8a
zb2aa66c1bd4587e31af966ecfd48fe90155134f359b93065ec319a3eeaa516e1ad284b7dcb76eb
zd2f0315ed4b6b6c5aaaba5d97301cc78fa02021353aa8a886d2bb54d81fb75a271b9c858e21d60
zd8b288ff863e69c492eddd01d2d4ae54c5e97a19352b0b276d0fd3eddc13a222454f7d46c421f2
z5320ca1e851371983a9bb8066541e0a656c4eff988db491f2dd9cd5457ce7425b28f6aa3ed7b3d
z8919eda7a8a764d3d07c4bec5a58860b3c0603e4e474070b0a8f0d0164e658edb762b6a82f6d9a
z77502776e34419ed566b8ceeed9f5f7b71d47f35ab3ea155dfe8075d2267e8c2838c8380a46f5a
zec3e24de4e70f10ad0bf46946c429399a06870e107e09a2dba351bb9c4b2f35ca0fcf4ba496703
z59c88717ff3970f2110d0f5aeab93fdd6716bab6c827c32f6b4f6e96e6705dd69cc0a1bedc8aac
z7621835a847e9a908638af79e688f475e5b7658d935e2671ee24f999d9b4b4a91c28de2766002e
z558266729d70bab4612f46720217670f560b27e0757ad6ec47e69db4c857fea02285459267f620
zae04a8e2997f13959e01112c644f9c8c244244bc1cdfef222b8fcb9b8e85a1e8781ce3575e2ce9
z57cef2c95f926f8d914230193ab005d7e1426814253f36eec1ae142df0880fce69be018eba3e27
z88bba09c598cca84de3acf566a6e960b8fa9b9df67f4f85fa677dcd7889fc16476140f29815d3b
zb4ab843118ed902fffb8f1573a8acf88aeb822e5e9a4d707ad36b8cfa571cfc5e9a25bd5d48cac
z3b5f4a60a86d27662bc0e4820635134d64dfa14ca099efc0dadd3c7676200034c1a3fc5e5e3088
zbdcb6ac31a4b88e31d29cf2aeb341e1b7b3b3f3ae5a1591500df6a968bac3529de850367d90765
zb8ef8cda2c454ec26a87c7b8581b039298c61e99b3e3fe0c4c86e0c7d4125bd9331fb00f4180e5
z9edd3459b03d79d67d90be48c9d74a43c1ccc4bb4aa8aea5c5a7be16fb9f85cd21f35f96428cba
z6190638cfd52f717a468b64806d4c7daa06a8717a2e6f0445990f3195a016395538f349751f0a1
z16bbb2506e17ae3fd53b784e90e95ec1ff60baaf44a6c3349f7704854d82417fa08f95a0ce0306
z1c5e275a2a339be2b7056fd81282c35f80685d937cbd5dd2680d1d4099e3f51cf01fd36b603bfb
z54ac94510fd86ac6c5b9a8eb3083a4f868c6abc027a5cade14c3fa3112862e61bf3f8198b17a18
z4587c2374827fc55e11c7385a92f63bedb1285365e286ead31b799763a4c825990ea7565884022
z4d4fa6b334fa07243798cddbeec01eee41b29df74404b53178053af14d57467e04460136be1ca9
z435eedf907116d57209cf75c42034e529dea3a068c7f2c34e299066605db027a7a7c0870ac5001
zd550a96a5f485cf796b01152c27c6753ad6dea6967bb6da5ba86e06bd56de8c8835a528dd99d94
z026933b4cd3d66802d15190de0fc61bc1d77910b9e2594591b0f32e437ec57cb8b7a217da4daad
z9e7032dd825c013b7fe0e3cea81694b984b7a558cd1021b173fe3b7c37f2ffa47349158287233b
za383ba933e1d8ceafd8159efcdb128afa854c505899dbe38e7e9ec61ffd93f24298a834c3407ec
z72033ea8181e799cf5f677769a9e7bb2a3b9b246ecd2268709cd3f2544da3c61c9222439dca9d7
zc12aae4566bd36cadeca1b4c670ae09835019371d208a3ce7f52ed84573e9d5e4cda8e42acedbc
zdf9b01cfa526c545ff5ef37570de92a7e5b74cbc71c990955bc818b4a51fe5d8415803e7e91b6c
z1dd8279725c3d303851f6d2e46c2f968d4c1e799078673b632f82207cc5034ec97fe9996dee9d2
zd28ff406b338092c61e13a6bf11fac46ceef6ebf99e71836800f1c05171e0be84d64cca8198c78
z02a413382fe5d35c3b44ad7bb9c61e91f2a0277603ee1874886f277f97dfc90d0edd42bf5b571b
zb0f4d446369e9164e8b248bdcc99bc8bbed2f3d50617b25250e401f6004249201c2dc986975ae6
z41dcc2d23e5e53581c4d1a5421068650b279bf379729a365a61c618a1d039dc12a76b253abba29
z92b679822b3f1e663849e369652a8f39e96e657ae066bf311d62af235d9f2a8ffe83f1d460e79d
z4527b6571adc6d3596f6d8aaad631ea9a27dab06e1fe1f434dd2e14ddaee9574543a2ffde66c04
zca87da8a4f516a476cd09d4e4970272454c0061f39662b3e26f09db620bfe7a8725f9e5b262e3e
z7a71b5f4a799972a9e2bc91bcaed95b5853c96ed9122443cdc12aa7c5522637ad4a27f2639810e
z7b877b58c8aca82c02e4ee8fd58c13eb82b5bc3e7e274d9a66586016494610e3c69ef006662f61
z4844f8fb734116416f980780f6a1037f55a5c6c3b8d020727333c8cb10c9ae7d546695dedc32d6
z66eec7dce35792972e7c06831c7701ad41df986001f2413cd8a33f8fe77ca2d26fed3f7dc0bbd1
z304ab7954fcf5aae4a861123d24101ddfbeca8a78145212108e89b7a4e350b798f38a7f9afcd9d
z18eff9b4d0871d4bf674e9960be0d6347b5bad08d729c1c3de46a5b348c6ddc228a137521ffc90
z6d345756be7fa16688968d9fd24002b1e187bd9c393e3224714df016944380bf36ada715089bb5
z763c2e5206c56aacce833baef0bcf7c041f75408ae98b09de555388e51a1f54afca1c365ceab79
z16a26dcd09a465a8f2a2e561a6caced79e3a7cc4eb5764f3320050a73cd7ca0b9b47e1a32f8871
zad920dd673738679b098d3523a81a6631911a4761d6fff0cc13f3c17cc9a2898c7fb85eacd3e82
z2aa0f2834b0a73f8146a9cbc6e2bfa18f38ce8551684e2e4839b22c7b65d88caa4c17bfe8292fe
z9dce8adcadff964e602341727eeab45e9da58d621d5af66062e443683cd17f852885a2e32f8e87
zb1b92cd86f82292ef2fcbd4bef09162f7c2af05bce03cade91eb0724ff968e63f1c0773a009fd7
zd70aa5742da61163db1c20d48bbc2ce544914ac164771a33255763107c83d04eb3567abca6bfbf
zfbd44655c642f514dc7a6f674e88fd33c9473742c8e24bc8cfd679d9142524fa86ff6811f7ca8c
z2b44cb3fd6cecee4ccb79eefc80fa0e1d9bc3bc734b01c19cde5ae9bc6b066e1f3cd2ea03ee64c
z4913323d7bf859892151c45679d347736fa3c7efc2f631eb4a38328c620370884f0f8172877d23
zf5fdfc6953a0c21ff2241aba0d152d62d4bc9c396125bf1b8c8728ec0df15a176e4b2ca27bc220
zfdcc452694596ef1e9698d16c53cf670757443cf8702456dcfb038be4d28a4e4b2f95a1259e437
zaf90d5ebe2f3dd073d1d3a68bedeeff9e227fc65ccf79ffd07ab01e4f734c40532e3a3da6bc6eb
zad503481db6aabded310955b16e6cd0ce6100adeccf815f10734d78ced77814826fe924520837c
zb81dc2661a2c464b4507f77a99d5825a5b3fd3f6ed94e67a71aa55afdf05a0d07a7c72b7ca4cc6
zc6deeabb7f6896ffea436cf1ca93d0d87c525b8b750d948be1ce8e7ec29a63cc7b0dc46a2e85d9
z46e9c368652881c061020324893aef2a6f22990373554fa3b3ab68091f29e5d5d8f95a85d1a042
z6b5bbcfa94d3aa44d659abbf5d25390bd223406d88cbe465a21c8881443ec974e0e5d50331a6ff
z7dfc92a21274269851d6428cfd9ea623dc589ed7d02cce43c0036622173bfc14c3b45cdd5c0172
zae8875489bf069246bb2f27137b8b69cb062ff56c5fb040de88a1f27917cee7e25969dfcb959c1
z4460f2e482e6f56f4b8999d03e6f4c56297ac08ceb2ce3c8a82b4f67f58a1cb2ed286bf7f8dc31
ze3a78366acac6219fc39ba7f24820e8669245ff6a9ab95937aa1cf5375d4243a908c081ace2ddd
z0b6afb2fd99daee44a662f8ff997db3118bc789b4eefeb0b71208eb64b6acde2ea2946839a6366
zb32645d1a64593f55625ec7a4421ffd782cea44c1231805a96f98acb0dd61b88dc29059fb8d604
z647bc0420ee40af99ac15d05368c75234e691e8f7852eef381f6b9da93a2819e7f9d515a67c1ab
z841a1364d23a35fe03f9110ee6426602acfdb73f42f5bde0fce7ac86ad569220fe7ab40ef13ccc
zc8738ddfa546fdd32f9bd34166e17fbcea78a879ba76fb67e5f9a2d7744a0d0bd10c7f64ccca11
z9dedd70b43dbb7c826932865e2c185f58e73469e97c37691949a1899eda405a8bcea7751b84f3b
z3b84e60b90f29f1bb806782cc62ea2f8eebc1674be3c991a1bc2f573219b35da7fd7f4a4c90ed6
z77ad0608f6483747f356d2a77b48ac4db5d23e91246c1087b6338bb762665c377c6b0c36ca9b27
zb0c7a13a959ced124142b46d48c0896c36adbf7eff4b6c851386a6433687b112d0ee56a8a07bed
zc696e2f9a61198dbbbf4b63989f333d02e7ac71c8a5912a96ec269feaef602ff6a49834998b5ec
za7d07d5518acf2b515314a901465b3cd6b31f4563c387704321f2114b60d42a73d5dc112c4c424
z90098ce8c763ce18fd72c00327a563c31290ed72197e3d967d274c9c91972e37a87f40bdabcdb4
z1ec13d9d2a0d67cd4658a5a3d251d7ada4bc86026ddf900cf36d97a267324e4771d1bbe25cf6cf
zea08ea331ff133a96f6396fe029ce05d1024ae4987a14b73d342b978f4736c6c638cd7d8f11d27
z6f242b91f709e6f71cc3a0073676a44766f4521e766bf1629c5297c94373f80030ad478b3a9e34
z1f0c822f084a8d8afcd6a383750fd62c2ca7d0100c97da112ed004d4cdaf62d23868bbf2b12e6d
zf417e3b223008af26ce3ff2c2ee02c8bb946685e35f1ac006f8f4d27b5809e9288401d2de2ede7
z6d9d044d9874dd3ace615019ca4c9173e155eacf523b49dc30bd4b3b25c1417a23919ead48260f
z376627c70e3819cedff6c47d979653d6981d316fb1cf2b372092d4bd1c637d2b9d5eabb46e7ec2
z90e67cf2cfe4cb457cdc19c527082cc0e6908d2690cba714c982cd999376eb678ac72397780d25
z4401d501b50e85bd0db8f85198cac14257188a51f65348f2751a7d308ddf751c9dd26e8ca1c862
z9079267046f99b3212ef158d85f7b37f23e61576832b9357d0ce9908f500fe6d5a8a6e2c2e941b
z8e025f41643315153a65c74dd92d0ee2d4e14ef8d83a2eb8ab7b0ead26675adf395158f79a4f76
zdbddcc11822ec96929c688ef7962d2e25703056361281620c8eb517ab4170658fae841abc89499
zc970bac3a7d4b4232ba43a178a21a8bae34a5edb2c1e296ca83cf55e0d6ab6cd161755ec02b104
zace4022ee90760bd65712b1565dc02f4068fb1b0f36a5a8ebdce710fa52d1b6d628527f6dbf476
z4aad6b186846ef17be288879028777ab22edefe3e2a941c9a4d29c12e277baa741be07a61f7503
zb042d1b1d8ac358db1a25cf79bb303a324183533651678c431221a4ecae2858a7991d3bec70555
z4b60d0d29b751c46133fce9bf4065efde0776c32b2c344d53e69bb87ae3690302d30abd4a903dc
ze694ef09c8095eb1042fb6e170398fa2535e5faa40e50c127b1aeb1725c3db282ae1e0cf49eb5b
zd05bba21ed76374d971e034a4b2db1025d1e0d31a3674421d6be08776bfba2c27b5862a4f8b62e
z902b8d0142929108a2735bda9f207a7081be43626b1ee770d93e6c77f184546ac76997fc46ef42
z746509ac81a0d5da755a5430509d290c0b48f6f6760c99d1ac3b57b9102f9363ef7baeb08d9bcd
zc825bfafd5686d678f7660293f6f19e2ef9f6a07b265368eab11c17cf751fc5242e6988934e7fe
z979dd7b173ce0c4891e8d3776cbd689efdb0f9184700906e59fdc01bbfd9c28166544cafd1951e
z71dd972e5c1e3110514efd75b44ec093fd761379230cb49761234857ab813ee3347fa18095e2f3
z3262b60f1f6fb7c8d1d394c99a7dec1475810c2eb6a775e3bd1b95ac7fe09c260b2e4db1bda323
zf325c2015a43ea2c32dc96ee2959188de6cfc9c5f54ef29a18b7a5a77ee8ba4e87823f6e135a6a
z0f3991817812792536a1f47897b8ff1d51d34fdabb836f70ed146ded58182ceb29735d8ff3696c
zaaa7a03fab75ab84a3f5c560c9d67e13858f4f9c6de20cc517ef0863a2cb407fc343f7a1f879f2
z5496dcb5807580988adf3f3f5dfcd26c6d9ff0060e83519728299e279ec5d497f5669228c47b76
zd32572871ba0fd196039b22adb761cb9be791a208e4db777676554377eaf4276b43ca073886dbb
zd3cb4cf1f07bab0cf08d96c27c457c80131923db122d98f16a55f0be7727ab3c4e8736e560524c
z905e51d2afb913ad2cca342fdf3af194b4dd6d91a4104afff8d928fee9c1a67afddf08bb0e3449
z0a52f6a8a7a24c0968961bcccd1c6c93fd68454cd0cdc52e3e9dac6a49002b6b8152ef5842de93
z3c69a606595ef274d7d639731a506bca1d4642ac343d5d9a8f259d53a4eef78243fe67aadcfef9
zfe96730ed51d8565b34953dc395fa1f904472586344e91242dbb456e41d489ee1867ff95929013
z6a2cb3e869f92d9ca57eeb7568d64ba279ef179834d58a8c2671a5f14d680d9e561f4a126dff75
za26c88e5ffabf4f5c58c8d689b4476ec1c64aa8d25ff2f2ff49edc2afc372c07ac0d88179c275e
zd11d0057ffda7816c5f719efd02b8aa52dcaaf9aab3086e38fc670af2ff4dd59fe997265aeec40
z615ea183860d5c476f1f26e20b88ea0dcb9fcb346d26c4666a7e05fd253afcc45fdc9bfe1a3231
za5cf15736dc68e630418d33574e4ffbe093474082bf2aa989932c2e326934363a1ec395459ca92
za74e838b8dc03ca13ce5262bb630a96d08108a447da0cd2bf5a011ef8de6654a396f7a56de173c
zc603a2ab93bc4ecea516b46031d9735ad88e7a547c183dc2a29dd7981b88ceef7f486abebb8bca
z7595c7090894300dda6f06c3b3dc02ddc67e0f4383e8c3cda9578460756d26bc8600b58e62b815
zcb4317549fb7d7122d9ac22b28d0c7b11467c6d1dc77e10494ac8cf91863eab45e0bb2e65f656a
z8dccad7d8e8514179a041b40a69a018687d26e6555dcafbd40d478a59694811e95138540160828
z30ad47af8f7a566c80b67caf7912eaeb38879e3c364fabc03428bfc17ab78721df170e0f222cac
z0d5f4735e0c8248bfec322db8aaae92c5f5f95a336194388af856a0546d096724bd2c3d799488f
zb82e8b1f690c0166ab90005695e12f8965b505a4de8ba712c95c14ba433ba8b2bba61ac1097a07
z5fc0485ecbec33da74c0a717ba60c3a5111230573cf1909abfd6e036671a762198440fca23ad8a
zccba18fc3b6e8bb269e8162088d3c75c91373e1a454ffec3d5f1ac382bf4071c1878d1996ca79b
z33d46a564d765422f18cfa6751d8c4932fe16e4a3cc38e2858d57a77e3abfc37329f9749e2e06c
zf69b50e1adf1eeef8959a543e00ea2ea6de252e2f70635522370a1e8094785f5e0cc22fd213212
z27bbc42bf450ae21e23671cf12112941d00df97c1b799203ba88ac7f1661b33c4c6c8354908dd6
zbe23db7c651f83bb1d3af5c6bac98766359a9a0c644732b3c435c487fad938ad289dd59789a504
ze2dac61f2413db5bfc3736d50644be31c227134923f3f2b5df9896ff71643232db77e31a13cb02
z2b18927629a4130bb85eb3ef35da0b95e59075b911751f64d0535c35d5a351abdffc813d630cd6
zdc5196ef34575dcbd9fbfeb3093c8a07c7ff74bf228c2d4a9ee1c603b93079816ebe494f4ee5bf
z8b710e0ecb56ef730934134c98c94e09ee468833b139b449c3e6b9dd4826884961545dbe0d5341
z4d9fa0dec872ae62fdd209f1e6e451624de93fdb52a6b0e228a49cce60102f8f9402900f37b816
z090913028bd3764f7f7e1b215204000548ab2cf29ce564854f603342d559be534fea7c516764e9
z5b4b168e4b01e9f9d25aa9a19e9c911cf8a269c9ecae3e80ce9c5c9d4e7250e3335393adffa72f
z3aa59d7ed64c3c10d27f6a39c926060d5c9ed9dcc219eee3886826254ed766a1cc82a82df8595b
z55d5b7ae36283247c08d424e4a527e286b485328ca52a149061b55baa398ed6c3d6b1341101638
zd658941f3ffd14e310002e6a12a4fe58fcfe766c05c243bf3a5d3bbecad68417833c71d127fee8
z82ac8e1a77b87e3270d5d0937afbb10b9212a616e3f302d2c064d1b4635de428fde9490939f1c3
zc1f33324df24611fbafa192775f10d3e7bd7cc3f63d5065cb1d49b91f1a1f0985f0bfaaad65a32
z5fe014d136fa4d4594d5a9bd7e9d72213d82763e613f605298cbe127af8513536de1ed16374c4e
zc05e9caeb3679ea895e5e38190b38b1501d962f5baa880743ef9b22a7fba9726d87060f7064d0c
z5680fe8c48a8ba0e17e09739d2c9da41f8e6ad5bc212362287dfdcd95c473430f9b8cd2dd0ffab
z3bcadfe7fd8f88b5afe7b083227f2089680610e52590a44812d558e429ea73f699198e18663cc9
zc18ca04fd20b4b90a7db6dae7309c701354ef3d63b02db200bfa2795ac201100f1ad20419d832b
zcdadcad3328d400d018e21513db7044451037218bada7f1634ef3a98cff93f59abc763c38539be
zb71318b41069f649a63268f3bf7adf44dbf2ec26adba0cb83447b7fb32b34179e49a70d5a61744
z7195db6e1c9ea4b00595326e38874754177021cb888aec6dae9ab42b5d92cba772b52e4e9cbbbe
z23ee9b1b395eabf0d7d5f18c0a2d97a9031610e830384b6ba33511bd74250686ef1d331deffe7d
zb9bd02aa674184d7b56c4bf0448684aa7e7395aadec8e4ab30b291b775ed657f6da1fe8596fade
za705803ad4c85c0b4fcde85cfa597f027354c34b4b9cf084e1509f7e3ba8803ce618712b226278
za10d30fdc2704d3befc602fdc28697b7c3b415eaf533f5b3b2a46334a901c3758700f103c52525
z5bc6e12f87a3bfe427f4bf968a48b8cf9143dfed094c0a6156dd17201a751b0d3ba2ddeecf2e86
z423536b58d1482ad7c1aa3bb5236ab5cb70a32d04d986532d31ff54f49984125c71fa2ab22de02
z9ec754e5d15a1ae75ab4c64023de1b08875b51c0fbcbb59663a8dc5f7c61b5bd5acad3230f604a
ze2c408105b8e58b2ec213fa8abc0136f66135988a4805b96bac8d14e74cd955c11d07eff095d78
z67f4613d838295d60aa8d94437b0182a86a9d46acb3a3376da945d91b1ed3eeb305e090e9245c0
z265888e7d5de648e81591d52a7ed1ee79a48ad844eb3d0eb62628ad7de4dff000b05f5edfd9a6f
z346dfd86de56397671df971ec3dd16d29ffd945537ac577aadfb52ffd0294bd968b77393a3b113
z910c5d0bb1d08dc0eb2bfe3048a6ed44b626851ae8e023e323d0024bce1d8cfab0839637d2202a
zc9e0be3942e636f6a14db9e0241004d1a886258e17eb0de5ae77ed28cccbe63d4627031e6db47c
ze72eb776853b31daecdb11a60561a1ae81406f81af8e3692d00b32d84e9f87b41e4fc13966bc04
z235eb94a7da7d52bda8475c3809851c6638236a710f144009273fc7dca8a07c10d11e3d97a4c99
z9761d6096cf69f05369410a4e28b05f0f79183975dd53b60af6698ff0646eb3ae7fd1c622147bc
z1e34c6d0d2c68fd4440fa16b40dbb3085336993a57f0697b1af43e3b250e79ab24bf4917b63c07
z10bc0cb7a359769ca02ae2885b7bf2480fd50e46460ac92de0fea010da73fcfd858eb88eba56e0
z32c36b826a849dfbe2ddab381d06a963e5007b0b5b8367a2c94977ec08515c19a9aa8b18f62165
z9457c07cfd20bef2e526612d55f4ae287e6ebed160e23577143a6cfa05178a86062ae3fa14eb64
zd6b8fb608b492123453ab9f60ab537b8bddb1a112dc9002f041fdd529713bf42daade5cf2439da
z2d25e4b4e17c014fbe7027df8463c183ccd969b19db19ddf843fa2d36c89c2dbd773107b9a071c
z713823b75d90346b90b4be14ebff3b190666da91b29cf14af0d50f2680cf20a21f94e7582a9152
z255a7d6d180d7d1f3639615d1893219605f045398a13542a96fd0d1f4dd08a8eb0017ad2259d1d
ze542a94edf2ab54055446f3bb5e2dbd65182f7a5409c19623958a057932b0de22f8cd55e451ff6
z9c865b493cfae699cd3f734aa4c4553c35ffdc70c7a0902132373afd1001a5c84f4771b8c947d8
zaacb70925a84c64005028fbacc0af9c7ade7cc021f021b26416eeeae33bf03d27df62e97dbcccf
z703de7162633be0f9a894d30f817c5ac623ed4bf8b264856b3aa843db33be462a0458a3dda36e0
zd92b29053920c62bf832379e8be76120f7e62a26a5d29aba4dca19194fc1a2ac72925b2afc8805
z787967a2086353ce3fffa994220add28141209cba2a988073deabe5ca9f7468f1338f5d1462ae7
zd1c794b98c0cdd304f9a4b3261d25cfc215cadc68993a4ddda3fb99dc9be35a47608008701dcd5
zfcab74360f440bbd205e11692f27a13468a44bf0acc02a2be47f3a524b7cb57dc0deacdb6b7fa0
z3dd42efdc170a1a31945da177a16a51932a45e6785785021f788949af91b9745e005f8c77d083b
z75b38bef746720b1ba6d82095277203132d349875210284dc4384027f2b8eb6f993ada74e2dc7d
z96030eed5e8aea012f23ddc8566a5fc2d95494cbd31cec65c381589b159344c425e517a209b6de
z5ae6b49a7ff1444fc633b00de6e6908719def2045e5c72988fce88d91adc17831c5763e6d51d57
z3764071226408f68468ac9e41d9a723ec0da84e8a8287826758f915f431755b490035f6c5658c3
zfcb6d6d340e0bb67ac40f3e0592744e665e2d1445cb06b2c493a51210526dc195417cd70e929eb
z2e6a80a752ab3ef9a7fa6e02d4657824f2e08448fd5568d0ff81c73e0cffaa9fac3789b6a2ea20
zc9c83ed94276ce967290d39ad91885196c4338d84041ef843af38c3e1a431c2d5323952bd965be
za730502d2435b3283db4c4ecba7881b51e1db4779cf677ddd264441d65ce0570532dfb82c45beb
z716317161b5311fea10c8da173ef5b738a926ed64d274b690eb0c0a3d6c780f72ae59ebb013bb9
zd94a83c75e8814d56f601adb2e18ec201bdfe6788b0537d847e069b5f2253e1f1600ee60e5bc66
z082b7f7318efb19c739872ca0746391c3e83dfb807aefac31881ed2ca1819362055bcc69e6a6b8
za8b922b85b8c8b3c0f228bd77d8aba008a621e3d1aa61cd830facf58445a3f51ff9c3a0483c65e
zd76dfca20cbaa91945112fceef3c9a486c5fe120c5501c29af80e866056ea6467db34555c6179c
zd855e199d4ca35e85492bd417a3c4d10b620e1f14648937f9c7b5d7a1bf16a6076f4edbc0ea91a
z5aa451c41b5899686dfa9eafe10573a61c7d69d9e8c74dedd1b9eebd888b16328f3e13feb53a1f
z95cdb377f2d5a211564a636a9005a1c7d52530734d1ee0adb8cd541677092a149856a6fd54dc6a
z7acedc7825e1d40e668fa2069d68899cc89a97caf6b283f74d66618c0852d9516f4cba0511c770
z502a67aac7f03e3fa1442d17fb100875d6246dd9f1125de12a5b9c2241b5b2f35d691d6eba4668
zc488530cb0ef8fbbf7e3716fde6c45713bee32161445f101f5395fbd1df1fd5a1958de06b7f23e
ze2915606f28648cd9a2969b20cbeb80b16d0755359e838b681da911f3b90eb9494629b0e2f3e9e
z25b512d6678ee824620e68670fe47e53c76cad226b8ce80aa807a4771a317c2074bf280658e2bd
z3b0b2c51034025af97562e30b845529246d634bc53aa5624d97397eb7984c6d7b94763812fb829
zc40b1ea4797729da3f8c76a919870f60e553f3ba7795d5fb978caf93e01686cf858e52a81be945
z930c392237b0463d9717de31d5530b357e3682a84e7eb709f320d62827fa064ae58c93fe399ab3
z128453444630c928bbdf75e2679e18e16f425cfa3c6a7d8e42ef20daa58a07b31b531c204c2a7d
zc6178f93bdae8c1eb8bd11ed6741521660f8b9bae3e49dec0945b710cd872f56088d40f20774bf
z069eeafa5543acb660053eb8200122695ebd0ed692b4451b776bcbda7207f03b847cde7e0cec2a
z8bb2d2eabded93a2ddf462ebf1fd6975b4edbf0509b8495d229fe1499907892176b3c082f90755
zf0bef46ef4beaa3a2e20626105a9d6af8629804d63d00b6052310582d33cb8cff7b9107d709b9a
z2589876ed2a67e57393cdc24f18e616880e871b9399cc98100bb1a4e71d3083ea1415af29a7d92
z9f6f48e6a3ed7c4c600cd51ae0e06249c855016cf29ad3429ca8c1bf817270633e197dc4c55ac1
z436d2ae4fee7fe858c14d6bdc21bc0da5d4827e1edb68917f1793ca23aa1e375ca1c41bf9fe655
z02868b31f04aa1128e455cf4bb2a16192467fd205b11408d01fe2bafa9a3f8e36c853db5f5f002
z27721167508b16de301993931dea5d3b5c947fabb67c4b45496e7ee1225bbd252c2307d17f8a0c
zf6888d3806231b35f1d11981ab2c175650c4163d3bfc7e9ec74b7f2290a44ce9242f76dcd04b75
z83d9d07a632fa38feca9b1557b6b0e3d591d2ec8170b9264588ae0dc98db24d7a3a14b1bfc6a2e
zf2c559f647427bc61e3285cf69d8bb7646fd0bfb5e0fd05b18092e61f1fddc3bc6887d30b0e9f1
zb1fcce0a6352c9f837147c5b3b1251ad80f85e520761ebba609bcc5cb78a7d6c8fe5ea555d861b
z083b7948cb39b52cea399cbea144332bf60858e42470c382822148a078195942bf9a3374fe5c83
z5ae21f07b0f87e62a05aca38642afc119b5c12da9ddca0ba433a295f71bf662000b33471d2a048
z66eb9d2c191dd255da12e367386bfd8856dc3b091ba051189c4b76de17b51c9ab2df4ce71f66ef
z4a76abe38b774de42802c4c35fc655c8d4c2523db683094881d1931c17eec2f9f42aa23285697a
zb41d538aa8ffbf2637958c63359d01161ea885fb0e75268075949f6c0902217eb03893829a06e9
z546536b467eea18c5461618b7f2aca28e3c727c66cf55376b3a72dd0d4ed30c10ff2d11615f58f
zb8970ec3354a981aba8b221cb6007251e427ccff580d5faa14beadb65cca00d097ba9de3108576
z12492184d25501916b594a443f2c4af15badddc7c405ea2c19ddbda11e817bea43168d439e96f2
z7dca6e91196bfe543f4fab0fc4d054d480917674ffa04ab49157104efd21a0a3450af64168aaa9
zb336379bd17987c7b57494143049f294669677e51ccf4c189efaa59bfc2a144d04aa10f2748231
zd84264f3bb0522b5c9ac859c6927cebba65887b4faa7e12bf86f3625060f20096cca52eed4be3e
z7a266ea4dd233b9e7f86b6d85df9400d90360c84e28da4b4900d2e832f04365ffc8dfa7c851280
z9d88e4b553fed859d63bfc888c15ced6024a6b1e2e2a105a19659e9c7aa24426e6880f2816c7e9
zdb5f94275ff4a52e4a2261a6b6b9af80d7b7a838834cf771109b2170217c7fd4ccc729ca8bd0bb
zcdcbf633e08e24b8bb2c6755556ff548a5980802a236d45fd47b8854a4b76feb154aa5c5247db4
zc753e3b7ccc76eed5918a380f461f8d347ecf7b9a7aeb58075b7a3ad04fcffe73ef4f0ff346ffb
z821fd406abb92d3099d3f713fc07f52abf7de5a4e1a09ab3609ab6ed495381bb4b2f5aadd7b7bf
z187d815c0e58bda1ecdce2edf4fff9dcc72594274cb354ca56888e12ea0b3c00c286d4245d6cc3
z0c2bb0dd5150dd8ec24b6c883d45eacda857512fd11e4a04a85532b470c4f9c1758379f3d5499b
z2d6945009a1f15e6b2f65f7f18ba44996e2abd2fb6b273a140b8d90f693a781f325987b6d846f5
zad0b5a8268d849eac0c1836c72996f79fb04a7603959b4d0c1d7bb22626d89de38dcbf5e78a2d3
z3c6ad682c447ff532392474509b11d2664e71d36f257c4f0bbfe28be573f648aebd93e8ad35551
z894d3dd88dc3a68d6e63286808ccb3b6d6a39b3fddced2020c3d1e1495f07a177ea4a1f63378e7
z55b9b5e8aafac99298809b3ab6a5624fbe87a51ed86c166ab9eba943bd3ce5635fbbc86aa2f9ef
z1ae8093cbd9105ea21d042fea4ca6e5a2a001a621b909c62eee91df22e2322312c7d4635f8e298
z71807ddbb954c055b17384247da781a8c53551c2f407e65063a0fb1d3db48ef48367bb310b57ad
z6002ba6873c4b2bced10f24934a6e9da65b3639ad06916c50dbcb1e5e33fb30100fcc13f15ca89
z5bb46c202bacfbaf6ea06c3d1b1e098850b2af4b835e7cc79cad0deb9e81590307e3cecfa80348
z77052d7eba1a4c0b06b3de58864a718abf9bc5b9f0b3199550889ba12296ac063a31305fa6e717
zdb1a1b65cf8a2fdc31324f44ffcc4a64be923ef4aacbf391ed33efeee4a507eae421404d515f9f
ze6a1a13fb992c272ddca289bb96aecbd1f0c1e14834774f82de0e89fbf33a6609f9d7661b7989f
zc73d7371b5671bee62cbda3ccbfeb8cb2dd0f43bedfd996c8d05268191ff2c3f1a90ed216fc4b4
z93e518762223d6af17ba80fdf44bf760021c6bbbf26774ba84c0fb6dffe21c8bc3d2ebe3abad3a
ze4fadac51de85eacf21eea7ffa78b908114e782788a1a932bf87dbd0215a4dda410afeaf6c65da
z5c228b27bd241684b90f52ea8097d10bdadfd2f661ae55a7cc90f5c5a884fc1c54e99166417f29
z3aced7ee2b79fad4412501acb0ba3b0eb020f51d51920d6c40bb3c19155b697e0b7241e21eb930
z03632b16d1935edec73f653ffe1491f8ca58bf0879eeb6769c20d09accb56c94a6150457a56249
zae7090e27111b87ba58dcca1b6920a0003d8a4ad6019f149f5c7223009c7edafc500e586411b8a
zc20f5950fd6c62acd804eb16d600d8ccc9f5544d89e96e599c94ae783da0c76e5286a1f06d6a32
z7ed368d868060885b3a0ccfd2747cd0ec857143bd232928f070fa5c864548ddec0f79470d1c9f4
ze103923516c57b73475c09bb2055e52886ec18899814f19529cb90e18819a78b9663640445b261
zdd635d0720ce1cbb46f08a645aed4c42804eed31312346f6e5bf9bf299aa77817cb34e2e55905a
z63a5dbeac7d7716ca57d6195478410d146d6749c13d6411a5c4031588fa6b859ed40de34642654
zf4389d8295ff997044c30561259b7dbdc2e91450aad45c4745236e6810bff0423a5da5f6bc44cd
z9fa526d54b63f1fe08c2b989c55133ed3575304a19419dffb6a7a9302270177feaec9baa1f0113
ze78da26c3598ba7aefbccdfafca42dc23a89ebc0bfdaf8902c633429d489e157073cbfc5e97824
z57a8fe9f1f7f41db25e6816d609b2f96998cc3629633467892471c8a693c6f1609d20c735d9634
za7ca8daf214575a4f3d2ef1a0c0569ccf158c6a9a8285aa04e02e7a5d543b3a8983c7504151080
zb2adac785755aa55497d510fe99cbd993baa705791aefb554007c394363a3b4a0181a093cadb1a
zd09c1e08b63831300618cb6fdec3ae9d9a288def7851fb6caada68fb816c971dd96a40c8138e49
ze92f39ddae0eb4ec0b2f1e7b2c2f826dd29d91d6f0caafe3257dcea3d8caef33ed75b1b992e807
z9716b26fc2f58a7ce6c9481efa6764e926ffcbfcba3a6c3aa61bd85866369d914ccf772b8f7670
z06d1f213593760e36245e3924b1769dbc7ba6fa0a01e8dbd2ea884366644acefcfe7e13868f9e7
zc0a088a417acf741d8f1be25a9f87e00b492d715558dd1905ee3c41a2285c447d9efb4fbe71882
ze19ebb4adba141268ec324815914b2d6c8053fcb23026f7d70248da3d5ec2d676c3ad77432e783
zdd6e66da1f88e3ca08230ca33dc4b8bd37342e6f7c7dc040c7a68e0c53e33653ad8d3dbad7ae18
z450dbf8fd084f14274f8cafe5b05052f30a612a10ad4d38da058c279474730157d29264afcdbdc
z06ad1ccb2bcbca5689b479373a8500097d2192f01c7b9b0502427c7e88bfc820c4b0fb628b37d2
z06c61df9687fd7a106d6140006a0a0fe411cff7f87a2f7cfd95743e02fa6623b6659482747ea28
z15df582a902139ae7d8436e353dee37f42b7a41d6d6241b22fa6decca217d3747ab543e619aa73
z51df32b562395c4f610927b3da0445c5c8d5c055891f5f1bb843c24c7c5dd1daede1d8a201e7ec
z26b88dff33fc467a4151b0bc55db9c22e78c3b6667d30fa32efc34cc301c40205e16f0efd0c2b9
zf61997b95e9c9b2277f12b835f3fbf185d03fad2f74553cb0f3ccb46beb531ca0f73bdf8a5de95
zed658e171dc847ed93929ff2eff484b10745bd3770e585eb244bc25d5fb4fd3d37eeef9e8b7a59
z233ef929b1cbcf115c262ae29dd274b4dc7097f4763edf45884e553ac63c9175103ff46a42e70d
z9a9722c21e49898eb15d98130571455129b780b59218e0c4feaacc06dafbb6c89a85ecc26ef80f
za1f79a04172b1cb27a1eebebd2a2311d133cb2aaa3d12d254862fdce243af17eb9a35279002276
z738dc826c9fe1a2ec786a16bf94f20970ee087981787828908ed7a850151586d68be78cea6cd41
zd0716a03cbb70a35733e7c2919e3d965214a281f66ec9270b45621cfeca775a278e1a541f94d24
z21b72cc5ee7b768700901a196498e52b697bd8675a3dff0c4ae4264e7e8cb3897367c9decb926c
z512fa4dec12854a9e37c82bbb308badcceeb5b5aaa41c97d7b3b16b6ce2bc6f8384bc096d17b5e
z3136cf837638d231ebe1ebdc3e08053c8ed21ee09657f36e1719af06444870e49c88b6b2bab3a6
z47ee408becb4e21721b51787c941b474355d1fbe569ce1310a9ab61c2a8342d95d6f6b833a1f7a
z10633c89a1118e24e6b1ef17b00ca31425c356812677797be17cd359357d926cf01fd78be5ea3f
z1e34743f0c3380c678b0401d0256e1096f6b042bd622f1818042007a46b2239c085b1cd8fae5c3
za2908e8560983176419c3406113f2486aced7b9127c58ebf03ec6e85f5b6d94aeaf5daadcf8d27
zb21c63855269d56f9f73cc971e610c35bfbae53a21a195a4aec90e5a9d746db65846daf8a4d69a
z7968ecafa1ffd23c50e9472b979a05dd4d9ba8f2fecac9aaf35fc6efcf359d1378646f0dd9449b
z2e1b1583cd87fd32c309277ae30ba82623a0d1175b40579dc23ffc971e1c675b53ef9b013dc0de
zb9bc24b0a7d69c1196c0e2796447da8746a767c2c89e134b834237e03ba706a79b2afc5bdfca5b
za4eda9f396b45ef0c3a54c922688f6b12c01be75956f0a1fd1e61acd1e07da7c1ba98da1db155a
zdde47ce9513608dc87529626afc5921455b6063b90a463ab758464aa17facf95ac06a810c43194
zd6ec8e77aae22da8cd0c9b5db108fa9cebc718fa91f7e8c443525384b3ad99ea4bb2d822cb93d9
z9c1095469f733092a1a9ddc7ad649a9c71487fdb682655a77b301916d545ccb4663590c9ebd998
z2cae2caa8c6a514dcf7f9397dee0af18a0a6bbbd9412ff5dcda65344616f5f61df01d53db6e989
z1f51dd3d3f4aa7fd3761e703f01d09ab70bf9106ae96862b3b717d096c252d108f6361a444b88f
z69b50e92295169bb83b4b79aafc9ff6c9b1d2b269c79c6494e52508eadcb576b1156b176ff8450
za638638e1927c8a8f842e60c4c3ef06a694569e5568d97d500aeb35b7eef05639da9330f5d24f7
za13cf76f753ce1563812b502e4607f2183b8a563af8eed9a5b4e549d2f9f06a9c42d6b010a4dbf
zd1fcb935ee591d1d740be1dd62cfff53c022edb0b14df1b247fad3c5eb1062b7cc33b2eef41ea6
zcc396bc68780fa0805d00336ab2f03f5bc1b51c53783403f45b14a4611d8994fb08b52219278e8
zbb2d55e57c4bb63251a4ec7532b6ce681ee14f69d9af8fdb2f49cf9cb76ddc7710dcb229162759
zf281b4be7afc276e99b79585adf6ea6e896c12cc1e57918b9b4b412248a9f6fda67d1da7f5d00b
z0644e6c9f5e248647472a11451c9fdd8f5bb98c3ff946858e89af1f4fbc1d6ca88b1bbe8e32135
z9d7280f7356c9e6140b98659734536bfd9b00923c3aec51986d7631f0c82ba5fbdf8e841121eac
z2d93a017dd4530f057dbf49ea7fe9a02a6f541eaa671bd4bbcf3a5465f953aeb2c642566b2e156
z3e9536e1db0b7c9d4d2733014ab534289a1d1aa60bdb9de4e8933ec149b776118f0ae8f7f1b67e
zb8d428b5194bbf74de52904f179fbea565453d7a13c8a6aebd011c4a609633809defad857c6bc4
z9e025b247bdfc642598d5476d22f7395fe143baa1a1bf34dafb7741d2dc6f8a642470b5fa4891f
z599d57bd762b24bfbb4fe8d7a4668526ec92cc59eb11a7a92f4a4f1fc18d1bab38650b12c3be22
z981698cc7e3d781d5a32e91c5622f26d34be46ed89288d6806ea68fd3d73bbaaf1f515e9997257
zc885782b65f25204db3c449966898fff23555a51f362928d6779a25be61b10d684f470f95ee654
z52f6506e5c2bbc6ff293a26d5dd7bfa8f85275a30e919e5391653d05e6862c799cbcd9e26ec67a
z06d6f699253b3f787ea4856c5de5208dfebe07a1366ce4790a653b5bbc2d758af7fa97ce7bc5e2
z7b91c1f06adf5c25ac4052ef915fbca02db3ef37dc5c5fe32c5d760f3c4793a32acabf22e1b971
z285e8174d2621f1b1612cc0176aba39a31bc375c6d78a42ca397f5520acb7b23481655de1489ee
z5104f9e273372c781256fc28345bdace4d56ff531e095f76fad62fedeb57b8824abd3de1508765
z83be40242bd5ee9204d4d05f1c771ff584a4e9c6a0851ae7d43646fe4b44dbc01b05f9697135be
z55f3def9f0f328c98c44e950163144d7396f73130b9ea1ba1d44b21c60e9883473252077f2aa68
zf0db3725b064503fd2f6650e4d58176b0ad62d31c4734cf0635841780b7f30d7d5625e3ebe6d5a
zf4eca62edf26f4011b4a9425b8d874910e7dc8912d709a48ebd6e26e46701a16697527c3dd0c37
z55a110d50c3108165cc2fc98da02635cccd8ec62e102db313d5912c35b709fbacbecc2f6245f29
zd15a14e4c28f5b26cee685b070ed30edf7384ac86add9f20596c66b5723c30e8ce6f8048147513
zfa31ef2bb6fd188734957fb77d6bbd2bab75ba196fb2fe10b99831f439d201128f10c9f9397c7d
z167a837e43d3c8c0482ae6a9f5c87f0721145cc705af3b7c97513f1ab917504fda33f94998d022
zfb0a06f3d2eef7124d432511260cdfc63af3397f79390fa9a5dd52a0176351955ac82a9751a630
zf821a7a5541ccb9688469e0004406069e569293e9269dfe36901e92ed3c95767a2ac39f5831856
z32d282cd52d6f168a1599bfcfb244f9c25521bc4a9ee76a0d554fb6a6e732afe8b0333ce3e9093
zf85f381ef396f9d41e69f059ff11e34de9c6364814477129c017dccf2ba6421fd7c5c2f28b3a6d
z41a0910659d02720b66ac3b9d21dfe6392a047bdfdad23d4166f6fc3379d173ed7e40ebdcfeaad
z26e2801e7a68c8bcc7cb5275953dfed0da670746c2733d47fa296d46a83db23b0957666c864053
z9a6986242f35ac0fa38c3f06708c26fa66a53d992d4cac86ed162be23d4e4ba4ba955ed8e078e9
z330562e55999442b096d44e6b50a1fe59c00d541040d2df4ec8f02d5289566c5beb732d1cceac3
z2a52ecd4f73e1ee7048b4c06696f1e5906cd21f9be24e19bfea1a1906da41e900a80700579b53b
z796b5b19a4b301f1cbff61110d2bc13e1e457f978cd186a8e61b16f4fcd9ce4cd0d6cc5db9817f
z1ce83827489ff470242573f4390b9f933d3439dfdd7e01d0481aa965e3c10b80375991c6eb25e0
z1a0af1b7f757e4efefd35bd0b4c7620b7ed9a7e882f8bd189842b872729cf45409dd884ffd5b8d
ze554c645dbc2c8e59a1669bb98e9c6e3f94170b582ce5444058d586b6b3a54a91faf7ac786059c
zb99c6562ac7f2c0638ba91190e8f451a7eecd1ff69863a40c4a80c534705834454ab51d344f11c
z51d7df9da0e6119b74af5917f26b50a1393b7879b867ca1d7600311a7549c705c0f8c7ecf249a5
zf1412eb5af261177e8b55292155e7fa308f34e27bb6abe6dad6672db310f5c2c0648d1fb50a5bc
z6538b771b86ffa6b9a703f2cdaadf3e88e3f7ad26aebf6983fd96d94a4879a331fbe91b47eb4a8
z2807ad9a2d035a4c199a1a17a2813aa53519694f29bda711942b24ff017043c7aacd69116903dc
zaf571fe50e172cd72ee848824167241e7b16c7528668dbf71f22a3ef9cc99311ad31dd538e9806
ze165778f687dc7d42d51f23d360649aae647698326b4af6e8f9dda02e44bd03896d728b22eeb65
zd3a2f5e647f9bc0879144257efdc30d8fbf0074b191f25172576e3bf25517606ad08738890ab19
za10e047872d59aea6776343ae0ca6b0802245d1f136025d90544dc826e6d4c0687348791ced99b
zb638467a45d8a57857b682ae5e9d8f8e9d98600d77f08caa94de5f2d263b15ec3f64c2e8d702c8
z101c2826d91eeaa1e0b49a015dc9c47934e49852991018a372949ae8974a87eaf5513089d829af
z7d0e0a8522d8ccaba195deea7d9d2d5b96a3c895d375c9789bde096804d4910c57a3e02d3f79ce
zfe9e5fe5e3f96a6a4aa09bae65ba33db30a5f063d0f35176f2c86deaaa7d45cb94f9f3fcecc8e9
z3fe595bc8c520ec6ea7787f3a59c154a1e3dbe2859fb183a4fa31ae06c7c5b90d807c1ca573e09
zaad47c87b6dd8d3dfe748496539dd245eb979c62510f430ae01d8e9778e0ac61bdabef40eb1e0c
z2491605594d166b9107e3ef0a6a5e71ff540ad8c6ef28c4d11e2115af8575bf775e6e58763e736
z5c45ef5c3d8d716c01c2270f7d762e4f4bf39d376880f01eb87caf839800054ee2cf2bd85726d7
z2c79b0168373b9dfd609a1c283a07e38b49802ac6274358d513b673dc247e78f122729269311c1
zfaa98f25e9c791f4835ccd87443ad749c0ca0b37f903e4b2ed91d99da6995a8ec9e322239610e6
z1d89d449c8c219328392844e723b993ee246943165a9b037556836dda303ac233f89d539d30d77
z8e5d26df3634dd79d9f8b66774083bf0fe8a18d516d05db0e7ce9b4c9cee18324c2f7838903fa8
z57321e64f804fed008e4b35bfdc9e47e60dc04d6cce4e83c45f76481ea5c16e151f6ea3bff57f9
z586b014fb46e38e4ff5690c5a2d9f25b63d90a593e5c46adc78546a193ae52bc2285aaf0c2cdc3
z2a8e7c2ad6d9f073975141b6ff1bb5fb1069207d3ab56aea46dc0112a18922a3361fc549b334d2
zdab488106162b7d42a7cce58eba55564a1a5983b5752df5036e63a291a8d6bb388ef2976b959ac
z634d6ec82df4ff94b9031daea1e156645aa58714783afc60b06f9161b66fa63a5467c8c4a68e4a
z73cd37ed82d339c84737541fa86e54d0b1908a3543242548c0517d3a399b6b628b9d14167677ae
z915d95da7ebdf7fbee7ad2f050d29165130f6c9b910ee680c30d59cb1cb67dfa8d7ac6d6ed1597
z754fca72c9d9c03dcbcfd633c22978b4647090be690609829dccc8bed56bf50aa10e4736ce4eb2
z3024484721352eb83db5b0b84d181a805a882ccfc0ae016c0f59b61b31799033e8e259cf0857aa
zdb4efb1e3be46773c1d61d2bb34ed3805d0fbbc3157fb0907fb234a34de2e444247ad1ae6c4574
zfca38060f4af99234b7c3f8a8ae3a700ad1f508da2bcdf34c2865708df08d102a9fc913e7d2bd9
z3d536a9601e57c4f308bb260f2e72475f15e046398f944f7598fb88c482d7b38aa22b6a6e22fb7
ze3ea99eeec95f972758ca17d839c7fb7e50517e5e2232a6abe868b91cc3328f9cc0ec95f4b6092
zdc4201ce8dd07ef6bf356758fab9a0d9ad07b697a4f20daa26f4551d55f9ac98e89c279b1f9816
zda105c83ceb4e4517cc8db8e5527f46ec2ae6faf3a412c4eb5d1bab1e95e147b7cb081f3d89e4f
z79104353bb2d3ebc42547ea0e7b74c5567b0f99a464b6db0a7928f4d0b4de0b697309b23967214
z208a9031da6aff32a556df16ba37dee4dbd32277525d5138cc41781e2b3282bf04e116f705a436
z4b52822651fb1852bd2974d7799abd1c495231ce31379b21cb4c00e7f12c727c7bcdbc3916d396
z94c2903cdeebc7c82b9768c0471f00eeec703911d535c7093be755a6b31397beeb16e085fb0599
zf279ebe364b0ce8eef059be387271e674f8297f0d552020d50020e5b09b7741a8a17bd36fb147a
z46ad574b88223272a05220997e3764acc483dcf3fd7e38f11935309aadec5e4babd32bd147276b
ze14ff15a6646a2f9ba155208aff3c722253da14662655f74f01eafd8f38c7c05f90b5504f7f6d7
z4666980fcc06a68091f387cfe820d2f33a6ec03d095caf0ba8a926d8ad73289d53c5ed229f7b2a
zce129778b2fdf61a6ea7cbcaa2c181acd8f7072e2796c54124452c2c61034b87a8b610e1bfdf8d
z512c1567dc8cd0518e1c2f52cedf92a320f13bae05c76190d49881fcd3e073e6d05d00214ed2e4
ze2257753bc3fc0385a2e8a110985ea85ded01b29bb6368ad73833c1f9510cb3e9d5391804db004
z9981ec1ee02d1a40445ecf67015313ea4b014e395c646198dffd20ba37c2f28febb6489c122886
z23e34ac96d034d94855864e7d2765f56382c66f926a2e9f1a466ce81b52db4b72800e2aa0bfafa
ze570964fa5086ad3a73c8638a762a4cd4cdee1da7536776aa65c2cb020e40f187c31e238a8d3c9
z2d2f32408b6e5e9f4f7dfb52e69839eef8954c131aa4ed7440c36b920d352872303c14e45ba631
zeb3fa92d5aae61f868c10999baa24adb205433f09e13fbb76899e642fb49cfd283358b8cd8278b
zced48e1823e5f3f1ec6d116f887636830222183211a3c5bf3781a3ff24660de8529c2371fbb4a5
z5727a9ff77a6a449639e4ba9ed0b9a6cfb0b9a5ae5dbb9c78501fa71e601b2912c12673a9f9858
zd5311e902fc95545c83a61470eb7174f12a1a5f5615c00c12f770fb36c4288c16701f9006c4511
z18f508cbc29d4f6580709b6d0c1fc5ecb7d1d163b3acb56c49846c3438143ea55bc16c2817beaf
z44502394da05fefc3397722ad7ac71d359e0fc2dcb326a052d55b5afc56013e45f916d25e3b1ee
z2fea76a1eadb1a7d405930cd263cd8adc0e608d29eb6bea7b2beeda6778b461882c3917e6903e1
zcaa60f0271eb822874ee2eca0fe20f4c7746183b6b30d9b2811a941e8a754de7836c55413d3175
z0ad4313f942620659beecc0964ef3be754d264ae49350355e206d651c6735354103c4d3e4260eb
z8173f319ad4067937797654db203ae521a3977ea4850f92153118d609d6cbfa3386e2194ce6bbe
z11e0886a98ca0634996dc5b0f267f4f7b65d634b614856187e8a2a93170b6f1346cc3cc397309d
zc53ff600b8ba3e2c8560cfbcf5bede66d0a546d45e0463fdce705d5bb7925ffeb0b1731f834cac
z6d6cb6a41ab396ed5b7ee8a79a0f7eb39561d3a009e7cd75b023eb0e835829beeb31d0ea9070d4
zcc56f490dd0c3d71242179cc4dbc14d6e7aa8efc0cc394f558fe198f9abe2ca20bcc674526be22
z22cbb07ae17b561b40e9af8b859f4cf1091ba36e335472f3e85ba9672535fde45a9707a29e142a
za838f792b948880bd32b057d90a6fe7fbd189205dc137391eefcebb31949ca611296116e728754
z95b6c2853c7939361a3d8e840a708d41c54e9c01dfacbeaaa1f0b77a8a6e16df4b6c5e1908fdcf
zde1b669b24c02cf4dab19eff7baa95272b8d80141ef513f8fff602ae42e9b55bbc645f5aeaa44e
zce960c086420c7ccf08a73e98605c960125893a4fcef06a5422bd4f7079871a34d66fda3e1db65
zd00e5433164b3f25f996efec5beec514ebeb7135dc3abf7deffb40e35807677365d0c29709f42b
z9ac85602b2c996c9c5401dc94e0d191b22b06180ce0e1317239dd20fc546e53352163ca4e7cc35
z50aa9e47c6a5b90ecd7041e0eec6bb0c0aa66bb603422f280d29ef5854cccf035397564d822145
ze9002be5d25e94523515767a731b1d752fdc07410ff63c9f00e3feef9c42a1087a18626a6fb31b
zad5484f7dae365be8a85459ec9c52af747c624099d9216e6604fb0a52fb3a1890a7aab04a4a057
z17e35873c5b385db98b391e5ddcb63a32ebc2a396d0f33f15e2d32da7f49cdd4fb65c92f32ee79
z5b39798c9b0911ceb599ddd0c5abebb398f9f0223c3724ba460024489bf3c4077b56d2bb20bebd
z8309a092a4f910a2319cbb7e3bd3864179100c7c169f7300016950c00a1a811509337eee2a8fe9
z73016ac4e5249872b43777720ef585afaa7e40a1697a5606ec96766fd81955c5022da0edb557a9
zde3b192c0d06d9627809f60dc89a26d52cfd0d73d60ff8ab9a8c7921e1389667c6a610d7c9f9b6
zce25e3f21be3a78d2e56fcaf85673c819a11c17049e8f70ad5ba26ff2938dc647bbd597620962b
z514d76813d6481045830dc57f2cfe8617a8f7c4413a57234a65659364fc67f0657b42fc067a9bf
z0d220983bd96c3ef29d5dc87df13ce7c572277167d1413676e57d2039b37ddc09909fe60711e45
zaaef852d1696dbdb245c05b0c20c53131b0062d3f76d85b601011043ba030e4e98ca899ac1c8a8
z20a02cec01f6b107f4bfc23c6108b09f75b8414de40df263eb9dd234f72081bd17ecb3502c5837
z956fdbb64c8066d1cbe3d82e754187c95368bfd571b80bc9b4fe65b989b12b064a5206c616e31b
zd67a67bee30a41838b0ad026cb69536f51c96f1519b84312e626d7e7ddc1ee453b56c68afb81cc
za611c965daba43d999719a625d3c013c8343e11f242282dd4aaff13341db9d255f2acbff022a72
z291829b8d1f9f099e59c51c8c95cda48b2f67b2782d2041b921abc1ea1e6a1b96e47a469958481
zc418976da104bd235774c30fef6eb77284f15a553790e4d7202ae94d48a9c7537937d1686dd850
z631799545dec2d8611168d0d76193d7761a5c6bcfdd6770466f5ddf159108947f6959dc4cdd4c1
zcd9f6ab3a793e078757866857bcf8de715c6c8f4acb6ad5168486874d77e7456d64f50f4ecf07f
z70b5067deac3be701bb2ea254de8c4c4f23613a97813829d62d8f79147600170ed2cb3cca996aa
z5254db00404290603ea07c8360f1041dc098aad78bd32683f116f1932ea7f651f53c30440f49a8
z68a3a477611ef14af5f432a5a246071c8c3f0e7a5cc4f8a8d9d06b728bc480552e417660214965
zcf9510db4cf412594af39ddbc3963f7f9e6926c192931bb8e336a9120cf41c0c015e9b3c9e11cf
z56a38ca6a84c5eef7b3963dab87795c84714fd8d3cec9f5b71e2a094483c546a591c93ac42668b
zeabc32f72317b47239f5656ef01f084e2a1faed20e03a862b74562936dc37f7ca8e523003c36c3
z9d00324c90cb73df41bcec6f291a19f0bfc43d18d54694753137b4603fde5f40f2ec7b6595ad59
zee5ec04db2daf86a4e0d39c03d0c1834b3b0837c9c8ed557f6c6609478d20f47d65c2c3396984a
z8d43cd64dd9664736dcb5c30a04a42d1b061dfd7910dad7fdbbb3858cf9e6b676ce54e3124b74f
z0fb5beb63e7310cc0be73db8ed8873d90698125fdc38e2633dd7a3fa73e37ba191993021862483
zed36d6826c98d51169a16700925af0cb2783d72b1cecf85289a329eb9af9a3219b67de5432a6c8
z8b7a16ef6dd57768a82f772d5d6638f867cc43324ef8ffc9ddb9de9231b47bb306be46513cd467
z35def325399e7fa7abf77f2309bb7f59eb72520621fc714df76bf6ff059465c82980b056179489
zde5d6b802746069667444d6009f640498c960314d888da8a2a0d3fa7e9a9e46603b37ca56f9040
zf4acff1e306c64a527166721396200d2812d6778640d7bf77da83a4942fc8e2f88955c90f960a7
z0d525d4a8895508adcfff2b5c08467fa9918cd7f0bbc65ec7f2ba3a81bff23155cef237f20f25c
zca50c47d28df3e818206f45f3ebb8549312829a34deda3e646b8dd2032d29aa669000304a6b1c9
z970e21126291f710f5c5c6ff234ad1d575ca11739ea93d8337edcfb0071e3b482e6ea22b08a25c
zf041248c0fbc074d1daa267f1b56a52733063ec118c1ff754ce74960aa09ed2f0a9d960b04ece8
z7e71657a47be64f2efc1a50c9153155f8beeda290b9095cbe375d237e041c3d1ac9d3f976649f8
z4536f14ecc33d12580e2bcae040c3bb48392c6405089d61049862acb1ada900dd81b4210aee066
z2d638c5a0ba8c0cb6934e2e222a55b98e777b05cf15fd4a2e665f38ada9069ab72fe5095048e68
zc300eaff0d806ec7a449ea61af688640313e0afdeef8e04250783d22fa8399f1851549bd72c6ad
za69a626648c3574702cef17db9565b409954ff0f2e4b4e6dad5bbfaa01820e911ccf404d0eb709
z8e365267d9c94d690be16bb4ead2130580500940734468793d9eb67525a30c690a2666a662d5bf
zfff285716b06a962164483f10082741b9cf839820d11f1ea0cff972b75a920bfd60d57af996f6c
z5f7a7817ed011f01e0e3908c27437ded0e5b327ac85793df38571c826319668698d9c04c2bc609
z406b2e4397fe990efbc7b874a7274de4b96f273289d11dd1006c3ee93ef5982a4c5d3ed7bec737
z9733a5ecaf2ac2b02ff9b0a3e336caf023732dfcf5680a97992a463443e8d44efbed17e432ca32
z3949e67200e92420e2624d480c7af983aff7f2dd50f19d532ba82965d4dca507069da660975edb
zf0acf503ab458ff753b1f6a53c9303f7ca6b612e22a1bd228c5d2f166920163a91b3d9d0fce9ad
z9445ee2efc1ccb3e2ac2f58215c3eecfbea8c7edd05592e7178a8a05b2e43d74337b0fc1b4028d
z17f5f7c949669645df4c345e793b0991f0db7641b98337c622d5541b051e6f2c9d180f534c1bd5
zc9db9f7b3222b47e70932b403ce92b33bb9480af6b10387492d9ab86991d267acfa9ecf6e27789
zd059ef351988a42d4559f5cd3d24d6cea868defae598b70614222b29bf9f26c1905aead4ca3e28
zdd514d07eb8ce6f3f795a4af5037563232500f63b82bd8718cc7a03ebd5a600f394d85fb0219dd
z79e7fc91c1a415bd3198a88d680baa9a528e221c8dc50870679db507ed51bbc1af7eda71ecf060
zb827d918094633dde2ac7f8ea46692b25280731e1b96663bd658f62ab36afb612e37614f2ca7b5
z4663004416a5669f5864c33947f66ee4b09e6aeb8eb48562f30cc95fd94acb464124807ee61f14
za837e2f010faab89273d477fcc33750f175e160a4bbf532a56ccf717ccc6a4535e12702743dbc5
z10cdd4ee160511eb8e359a205e6241c6cde3f208d8e908c5e5fb8019fb6cddb7a7108d642ce818
z5db2016cf5c0b0b61e06f1e482e4be16608bc8012294109383e37b027b54ff3eff7cb456f29364
z869d372d179314ab0718d31773357e116bafcb228fd1ec7128525fdb4a6474a8504bb86ea6163b
zb84ee553b10940326f19284f8885c55f9fa071693e8d6d6f46ede843e38b2e8cdfc50fa4b52b9a
zb05c807f97d0648d5a560866ccecdd8f62dc441a9ea9cdcc3d636a47a3144608e3923921f799d6
z5bec7924512e2da5f160b111ca39fb1fb8737a000bb747dda7bb1fe07462eb0799060184b0881e
z0d09715ec2cd21643f62f66bcd8e2080263d01a7c71f6eacbcc0a775d2ab476a8805a72071db35
z6572d42659a1bc2e42573987b0da062f5ebecc23926a2923c516508d63d692fafcf2304f8a7862
zd8b9164a0e05f77e47df2cafcc7bd600d05b02e0a70356662cc60e4805059c31a19ee882e3380c
zfb38867eb4f89737069e09f5fbda50b502c469a3ab7b8b340375223aaf893725e7eb167d6a1784
z10140065ea6abf75857cdb69afa07ba2abbaee8a2de9d22cf74b5d39a79e63feb5b128090d08c6
zba51459e36fe7f78319bdd66c3ff17a80b7e3f307d0764820789a7d654d748bc67709fc295ede9
zef78ae0895d1febd175849dc8efd0d9d77521dee756d408667f90b6505258eacf2a44783774ef7
za9bd3542478c581dce136344d5ec335c2e2ea9a89697b52dd5b32ae1b506a634f0c44ff431f8ee
z7f6b454e87502cb2e7db08edfc5ea04af72e72706f270d163437fa258ae6ca1f72c5af09825b22
z19e726c840e6542ca59f8b27449dc4f93842c2a486c5a782fcb7c5e115c62614e36e278a87909c
zbf079d86937709bfea25c0a9ad8d4cf9ab53f57379073ab6c3c68eb667a044c734ee92b0304167
z7135370db6cbd9eed74bff3c91c4f0b28bcd9c45fa4502861a232530b3534014e0f93903aca9ca
zec151ed2d572f98a8d407ff9bb6b7e8391945dedfd1611b3bb1a1ec3475ddba81f721296fa0a8d
z59ef99fcf060a7622093e8f34f46df5b77fdac9afae7a2d0e5de96e9d66664414309690a9521f3
z5a349695eb814b454d25d5aabaf72dd510d953fddbf5bc5ece7d284f11eebd2c5d50f4781b9b60
z55326e668923377389acb711c77984915dd8de84272325b30a78d4afb2e428828ed23eaffda607
zff2a1e3f53ab52b58d3be1e534a6d909e4328d3e4d1897e54bd777edb8bc6e083171d61111be9f
zf683db116337a7a02fe01de199a4aede0727183733152f606fb10a0bac47e6c8dc7916b759816c
z8db49d611b1934114bca40751f0b884b220050f45b02b00cbb9c5271b882051612a7d96ecba7dc
z6d5b02b65449b5c063849ec551346692d4f7ef53365d5d9ba2a3d75c92790cc12c4c61875dc3c8
zc5cf13ec9e472b4476457f17c2d828c2d34d675f300468a22de8baaa0011a5a9ff3621052df6df
zd680d18a7966fd11cbeb62dc9b07c45fbf4949ed76bcbdc3606ed28d47d3111bb675b9af8f0df3
z6f0892ac1724f0d55d6354bc0f2e3eedac829647a9b6fd3b8fe9a8e454ff2c3ecd890f63a0fbe8
ze5a7c83876c69f3944ff7187b67b333ced2d15dd81dab2a4ecb8170fd37e7e52a9b4cc725733fb
z09136ac22877309d3f0754351d7147765267d704fa6330c6214c9941d2bb9e4324864fceb6677f
z46f846674668917c316460b06a08688d96c69696715cfb9e666a85254e4b0c12d461f3977e8563
zd2d3bda397e7860098a0ba0ab24ce23d3c7139b3930d94c997bb6f566d05677254fdd96f6855ec
z0b6b8b4b2d0c42c9791ec68ca6a79ddc083f1aacfcfd6b932ad5efc33c06f9f1daa704aab16044
zaa061a577b585d23c715152f3e1d5031920b7ac5fb28eef0049f3b388a148554f5ade8712b5845
z7f47ec01f75449914c0a74ff0873db509da2504a706cbcec9ac7de2bd2116b2d2c13e7aa206225
z7e379d0ac5bc9a62e89b8cc9dece56656dc4b71b664c816ae601d89433a77eb4a60f8af059dab6
z74074998604e1e09673a2e53bf67a8b8258b76fa314a864f84941f5c95ca25f74a156af281fc21
zd6d00b7716626d3d2abb18cee53fb8e4a9a1f32f7a4fa1f442dd827a60062fed197e6134a84fe5
z164f1ed1f35706b8646e05946140fa29d98ae979631c426803fcbdd012b2167719e35ece328013
z64b444e85e2ad72122e05942c33a97547bbb80bdc53b67eec5f82bb840710ac1a4a499e73c17cd
z34030893b51de5653f1fc90afe7d66420a6a38ff9d43c44143e73a30f7e0b4c1cd5a2a6e05ad8e
z1b86163ceb98f4da58a683094cd8bc52f304b096b7450a90f8f1a98f274ac321e2a81e1897dbbb
z1919b232ed529aff29a5adca813d5ad2b772ec05571d01102e39c241e4290049395c04af05a5f4
z2abec887ab2fbfcb1e47284dd7833073b53e12cbeec801fb53b40e8d150aaf7c7416e93b3d26c1
z2a819e2badda41b94c9608f30b75c9b47e79c5ecb05cbbe516762c78c7c0fb9c932db551437d09
z8a1f039fbfbd2a57546328650dd1c53a71a7b37edc6e0b0071347fe027ba2273b07177e5d7189a
z831dc7394ae77896d051a7902bff564c726c1c1719bd192175891487f0947b7453ebbd84b48d8e
zadc4bcd21513e9b5eb53b00d962b5d59a77d92ea3d337ec98a402de8b3242465f1155abacfcaa3
z8f341eeede9082616941e68e1bfae25b6ef8fbeb62d4cd2c6a0632a5ad5d8299e3d0983c724ac1
z4626b66d822ddf85538dac666642927359d9d152b9f3e22e7ce56328a15287a1cc7176733571d4
z636ff23ec63a9e16f090cac80315bcffc9d076064d0264b80f511ec1afe3d3325638ca5ad8bc3c
zd3c260620fb15eee927e7f983d82b7c2401161c49b60f698b92452e6a00225b194711dc8b3d0c4
za9ab4baa6c8422fd6e71ffc5ed2eec4ab4f4a3789d8c59c894d919d10707fb7464be2b62f20ee2
z99e419b3be60fa0cf650ee1d42b5fb9b6cf347fb9fb25543aa4d312ef5388d8f26fb8f6efeae19
z44d984abdb76836de7ec56c87d36eefa4acd4341a5774c88afa9909d2382ea77a5930c9ca4d463
z9fce5e67d223f9a4b7d2178b158c39390f14f4093d12dcb3fde096a7966f7e1637dc435ad9876f
zb36ad0873878f9544bc1e96a2fda8e86ef5fa858392f753582a699797559f71a555fb87d98f1ee
zdd45cc77a1c5ff2f7ec22b62951f1c113492d23afbc5be24e5fb29e8e59366d0d101234802714c
zfaa5d53b801e79f9526dcc8e504161e9227751f0aee76c20bb48fb033e8f0f121818b82c2cbd0a
zbc1ab1a500f207093a70bbe788a1353f9899d0092ef1ab59114c10540bfae074411da989c4ca3c
z9d24ab072876fac74b970d61dd68a36c8fd4181ef43f649a75c95da11fc7b056ecc52c85f863fd
ze7c735495555b83c47247796c413435f5d6237e844d54392829b3311700028c4e9cfb6c66f34c5
z69aa90c2ae16b5a0678f3b06a8029aa7caf8e9aa66c0304658dc6840bf297343789663659a2d07
zcaac48dce2fbd3d605864cae9efc7a2006527921aecf4a8dfe91864995e6d0cf45db190a71dda1
z8683a8fe63cf7130e2a00c6f650e9afa32f662704b39223022dfff44b433ff4ffdc6a51b638251
zb48efc53bcefaf344462e4b3abb4dd1352819336f7f7ed6d360f5154efcce6f2b0627fc8b410b9
z830af6f05a41253fb91c56943948ecf7909ed4f55ca29f518c41afb1daf1987fbe203730d865d3
ze7364acafc1bdb82f3ed5b105a9d2832a5d24dc04be6478ae5a2881eb30fdfe9f69793623b3587
z1d4e51dcc286e8f3e809036cfcbe74c9ae90b60eee893ab9eed4937df84ab70f67b04b44973357
zb41f6e1be9b2f9e1205994673c8ac1fede4108ff8ab43418f7ac2a176f269cf2a5211d7c8b7bb1
zf17ffac32548b2964b6a49c9cdcf40a6e401b5b82d7cbf448ccfdf553bd0a9114b43769a9f8457
z39d380db3bff6a8143583a603a3fd0d242e661b24911c718464ec8c9bde8d03f4684e54069e125
z297c7c31d8e3685bad837d3ece8f9788a2a57e87f2e7227fb1ac53bc258dd870f87aa745441982
zfb242b2f94735307f32fb6e7c2413d876b120f9a349c47e64a1e32c9422a52c8430db7835b041c
z8bc90d86f699f0be78eb663dc14e0ac22a80cdd8960f3cb03e5cd1ccbedb35c00432c97b1553c6
z2a06fbfd39301413ea14752605cc5ffe516a33ebee34a7f57594e4acbd85b84f22297d35573d67
z5e064ac8978a73b670c59bd5bf6ba318d1e5a8996822f29eb2485c40832c38b7d7955aacbd5e54
za96fa59c56fb9ae5345c9cfb619c43d0517140d53e7ed30272a7041c18ad3b19e8209ed534a35a
z769fd0f52dff3dea9547382c1ae8880d37340585170c6f54bacfd45ed577b9b53a971e58fa34fd
z76f9356a9403798f26bbc1801015a7beeb9843b9ec53ec686f8f86c27d9cf688649a02b90484e0
z70dcce7a29bcd7292eb9aa00265a180238864a7e70b45c6df5c32204627bfbacfb0d7bc2d73f95
ze6348cc8800dab0a19b637be4f8341a0ea7d98510685e812eaaea5ca2b44eeeb2d525ca3f4bcab
z03e28065ccb1afa8a47495ddc6225bebebe6cb5b973cc1a495ace77dc9f083ee43d6f5d24a7466
zdaf58b2cb2d447df232b73955fc49b8c0dc491000c10fc7aedcf16bf8800ee83f273d50e4bad97
z2412e493f9136a047b724c061ac859afb58d5979ceaaf3c5e000b578dd20b1c05e7e89be2895d7
z51d1a3478b54d2518c7b6341686012f42bb7e3b575f4a0596054808f77d7cbc5a043f98ba0a46f
z11e394490961715142a6614f9486fd0dcb0344be429535e9aed82d1c500b453bba4a41197d062e
z2c879feff9f8dedb949634c629c20747fe71205dc52206fb015e01830e0c8ae48d3a2e21bcee24
z78ad8269445e683dff2bc2d4c9d06a36f54ab1ee6d1da3b43053765c1b56e1859d48062933c382
zaa042e601fe8865ea4e6021838cb3dcccdce7dbb16989da35c3fef4c499f5b922adce5ba624a43
z41393e9cf907066c13a7b4a4afac8bc41610b2b958ea35189127ca23ba2f8366170a904df80d93
z80ed057524960a94952597e4c72a6a700518411d0b8bcd1720972b57f838b95602ecda6710917c
zbc667e0c3ebc73627ecb2e433850ea9f0b3e2175e71b683b7f1f6f075cbf1f3d089b81e70917b8
zd7c0ebe6581916e97982d12ae4fd7b9f765f2c3b62ef5cab986626ec4c9812a185d4c9e3c204f3
z69fe5851eb18b2dbac2aeca788fcd9d7490002b6067a8e19d473468239869204851d81b0b43515
zdcaec6c5bd9b1e04924ee48e6dc4f923b207e3dcb5505065c3fcd6df008d8c157dddb6ffc8f1a2
z0e07eae3f43b9ff954fb161360c807f10f4499919edc8c0d6f5241951671bdba83a4e3377740b0
z307eaa43e9d80c8a22fd7368cb997f50a6fd58e5b8b9e4e4a0b7b220ad73dbf4ed8caab5277676
z630a13c2d566803fa29b1c77a3d757569f4f66ed72a4201d2155740f292b1db123d0f0a083d02f
z713a61e5447c9ef0576dfccad9369f4921e02c2088c3b1beeaa9cb011a5770b57da54509700a90
z25260038a467ab07d2499a5d77aa87253d8d61d647efa1c126475a58670e03918a23b013fc4374
zbde0b6f253adea07144124ca44dae3a4c1fbb78518f7d5c82d7d39c3256eee9e1291b4edace7df
z1547e9054db87f21c135e9ed9aa8fc9614aa77607b2857082ce68312c409730ca1946debd866a5
z26471e7917cda0602d68ced3e16f041d49da19c17df6b2515e31e94da30ff544549bcd44ba1922
z6d53a274058ac6d1c1ace72197f24d2c9768a4692a91e7deac6edb5b09f203b723860ed521647a
zd71c11c20e7e37e054c9e26447543bee6d971375b97ed5168d3889ac68a515b2145f4db9d16bd7
zc5a5ca56ccc8bb0a23bb61e082f678dd29421b888e58338e3c53a853b1217da49c58dec21ecf21
z888fbd17fde74b94223bbdaa349efb3075b1d1e289549c1ac207afd9471580b1ba38a1c00aa1c7
z463dc9b809c993a6ea47390c256e39fc9049d043888d419e50f029aa82393ad83070e0a1a44648
z5478663f2a349be6eb49b66835187eee8d6f91a6a3677458c82b364c4026d552ecfd2cba2f8e03
z26a2307b760701658e326991727f7f7dabf5614331e247f7b1c90592a400300baf206b2606d3a6
ze0660fb139b8a6628fd53c4de088358d5efe079f1ae58cb76aecabacda7864ba077647f18a4eab
za9a7aa0eb266ae68bd742c6790cf4c06b3a26bbf07cfdc0d557e1bdef847b7e9a61deec5a11a89
z8955fd4d46ddcef2d2b43e4c31771fcdd3b2a68cb8bf44e24783f75f904b0385eb74deaf2bb492
zeb190caf88359fc9400356c5007a0e105c457c595270f128cfc2a5cc9cd7b559073a5c4940da67
z0d8893d91d0d6881fd075e570c66c65b07637e948aaeddee00aff3ca5bd21c105af771549ea911
z37405bdd3cf928d52c021a15b6e7959a4d133854481445a09c7c066ce12b12442d6971b3590fc7
zef5f7fd3b734538d8d0a2036a984ea25a05ca8003ba549f5a1067d30f3a70070dbfc23f899978f
zb6ea6d60ad338478fcb680e5bc7ca4b448a78ab4f1154c1c36ec63514bac002414f9240619a7ce
za7cbd2f74444d618884956b455acc897922ee6b1eabf378205df17c230e425c7246b404fb0957f
z5fd16684e7e5c23f764f3fe2dca06f632c94c7caa08a04a5c7c936c592563500e84b0761d5c0ab
ze296d2a74f120aa5c89a071638d6a356aa73762b97ec9e7a813c456d1829d5706de55d1dff9df1
zd7b86e308f66a08ccee3f523cfab7331cdc7d2f36b455a61c7d78675323828fac529ce28b0ec58
z45d12b63f42313b44c094b765142477b90dfa763c649d49d68a878c5546bd292dc24ac5307743e
zaf92ba9996e9118b9aac744482d974caedfa905e70c53b224456ddf48b58f285cef267c0f30119
z5fd3ceb50022c50caee3d433ff62aaf9efa949adba6cdf23bed1451f74607a5241959784319ef7
z7663d2622841c44442dff6f17a706ec39475c9af3fb375c264338a3670d25252a1eafe1d5f9220
z775c295e9bf52788a9547146cdc834c78717f5edde5363b3f3d117bef59319d9f063c45c49098b
z0cf62294480737c26f1b04db0b902ef388a4d5d69ca650d42b1ccd014a4e7bcccc675f2600f54c
zec173efa598f09f926406a7d24b3263f29e05de0690b52ed6c14f859a3c7779e542983c41b327f
z969d78e997eae84419e62554a09f9555d2c1bc01c1dd7300567248c6ae2b23699fafa5a0449100
z6e0f5548408639bafce3b5bf47d959e43e674f27f9c902c80c03a9312ede54d83cb1119c45c0b9
zc6934c34aaf545fa274b6ac4ec587745d0fa68a9682fa1dc9722b51f64349b61961d80a4d6abf4
z3ada48b8a28833b41f5c725986947f98b13c2c2a227b6b05640a9da8bfa1256d4fbb54f7387e4c
zb898c5f61bdcfb3dd1db1d8ee0efa8fb20b34cba68dc47df0ba906ac4772173d179cf2470280c0
zf3240b927b6efab13be5a61d21e07e074a0ffb61f7b0f72c4d9a10a8562e0e4efdebf8bf6f19cd
zf635c9081ecd95bf3228c73cf5c896e77413fbc885307abc56cc9d85b62be8ea850344041006c1
za01ceb767591a12ebe6c564189b9bbb4d284d346c57aa885e601dbfd74f28dc94de41f5c58f6fd
zd695299f66e7b55b6e45facd08448e68763d58761183a61c4d05c0f741cbbdcd13c550ab5f917c
z2fd32e4b99c9abbda3c3e25ef052b1f01d5a6b69fadc1c45e4b057b653e9f1c7d91bfc6e3677ea
z3c6ecaec90bc4c5b3022f1edb986ab343bc3c1316c461c6da6c7c10be2cdac3dc61154af16e961
z3643abd194cba6f317e5ccf51914ee34f99e11bfce94924f7805631484c789c5141b9cfafe3bb1
z908cfcdda8fc72787921ccde5056669d5b0fa6de9ec07407106ae9cdc9259bb97cb466aa030a70
z78dd53545bba586d205c24b8f71b9d344562e771b4a7759b1e1bfc0587c4f345ae3f1b0e60f4ef
z026d79e5d026ce70d90c6f4561c831a7131b1c473c596466f6018225c55bae3bc226aeb39be9b9
z818c6a3edf789aa1bd34ccda7814eccbb9360db66264f7328e49d8557ddfe807148f5845cb1fc3
zcdfeeb156f866abade5ce6eb20381043ca16f79a6cf5955fce6abb901a80090db1db4ae76685c1
z1abf6d5597492137ccdd9614217548a344d3a2a8e5ef756078d100cffcaa6ea99b97b97b73720d
z6cf6d653898d3b8a1ed3836de69a544fb7eda3fa7c2e7257dc07b151b4346af4f99220a10c42b6
z34c1665c5cf4dd59d0b0a88d30d10b44202af5935a36ce75ef6fa6658657855c89af3e38f96393
z7ecab7079cd901e6d4bad759301773b6edcda345793b0c8f1dcc114c30129b2fb90ba4705803e3
zb2cca89f1031ffe2a7788451bca0077c514b20721dd090981a702f16681ef2ab4c06eb917e5637
z14f9aca006f4edef20a36e6c57727c532a5ca9420f553547d0cafa3a2185e30551fb4fe76db272
z28e26aafef47ce80a5b91435895b334696ccc0290fb72cbf6d1aced15f3b6e72e000e04a5b9f9c
z232df69bbb03737e792480798c657494ec2a79fda37eb1acdaad195d166ed5b605230ced3476bd
z19efbb80baaa2841776f3f163dc723213a1f6caaf583d4f26a7fc51a7af53b2be14eeb6d7f1cd1
z73bcf424153e8c5fcead26903a28b02d2961ad285d5c5805f0562582e756fdbc5f800069920a8e
z4a56e1905326d1e6c7ea5e48ffd9224867e0e1ac7f0a315eec9cffa814d6fe979b1b9f7e93e65e
z5ec00ebeaffe14fab143ce2981eaf21f0641c6c6a31229fc174a48c612d2984a16e38525aacd1c
z9df5b202b562c772d312a64c47ebff195b6eb3fafb1db750be32688361711048986574ca39321a
z6abcdde5f427a1e02cfbdff4e1ab23d1b213915141e32d457a43d03832f29369621d48a6804ca6
z42ed6dfe4b098eb0f8ed1992603c32871be0c4d3027b56fb0a015769f5502814535b3953791397
z7c691524dd38a2ec05c0eed5b45e31c55d8ef28391e030d4587b7bfd12e3afcea3cf068007d3ad
z2e526174eb200059ff4ab4457f26d0c8a1980ee1d3f4b097db9401f667e6b687125d999480adce
ze481ca99e6aefcaaf2cf1021f6965806510226f4509b9cd1bfc5dce51e983d1c3be1254a8afec4
zdc3a649929a096a9b6b92efaedd2b2174447022d9005d804bbf5177f98f9c142950d575d240786
z359685dd5efe5dcaa1c82501fb911516b3830a16520a3ef7cc067630a886cbb9befeb1720b622b
z8c68362b9f24112d7299963b788e989c2b4389c1650b657bc108a7b3f0867f1d44fa92145819db
z342bd578849df2f70f3a4c97e9b1eb271f71bf0e8cdaaf2fdbb3232c248857fc9f28d9538d5095
z4e9cce4c3f9c919e32678a2a7ff0227ca0102bfd35a570b52552c7458c12faa1b75f4f1a476d60
z9c43fa44ae8201ef533ad9c10f9218e3c32889dab4a98729cd417bddeda26f82347f40334dddd4
z3fd02ed90605aede49de744897c3461fdbc08def8f8657ca552ff410be41a65d637a1e727339a6
z8904a2d59c44535a80460a897cf59c9d435d1f4daa222ae84c0597b306f622cef9e607a343af9f
z38e239b7d5da0a49a703673e754dde5b85dde5ccda3c3741763da0da845b12e4661de8fe77b68b
z3a577d9f1a7e30c755d29e0cd81f109f810fe0d9536b57f60908a886d49bd833e672bf1d0126c8
zdc159ff74552d908e06dbdb991642b17f7f4a70a8b27a9f53ee78bfa952b3cb35408daceecbdc0
zf5c1960f709c8af94eebd6ddb4a1a98d6e5c8516e0c626bf1ce19724f61930d0587c79af7ffd31
zdddf4eb4df7533e7de9efac72ef8a8d5bb6c0a4b5b7c9e30113c784d16df9bae621a617202b1f4
z2f0875473a24c94b1599e8fb9b33ab1929b8c7cfff54b6ddb526083c8121280124548c55d4faa5
z0cdd927d46b369d36942679e795b4dfc51e6d970fc19c70f82469440253ffc76c62742c71a1fb7
z1a72f0385949e29e43eeeb147cc95c4ae4c2fe6e8955ddd946e5f7eaf148dc6a3129d4794d1c86
z3a35e4a9eac17b5660ebe426a65ce1b692b73b28ddcc865b1505b7b85d4a74732c11f0c61c093a
z0ea645857f22e6ae2af81fbf7e229313331c809f22436999a5442ff916a1cf783b550c2ff42d2f
z2fcebcca4913118129d04d577af3e7e2e3e4b0bf1c49da0ded3d9d31513e9231e00f46891bbd00
z2b7948a97e6af118dda0d17ee79ee844adf926d0eb335c651c33f626020d8ca096b2f4979d5c05
zb1359adb2be12c28ea129ac8bf19c054a3caac0d89823c1f827628908a40239282ff1f51c7db70
z932a1cea6c4486b798e9be37347185479206753929c06cb30202940141d969aed6b7f2948ccb5d
z347dd4e55bfb2cf095a13883e63727cf6ac9bde8bbb9cc56d75f4b0293c58713d1696ac5c427d8
zd7e750450a9f496fd7f261ddb5f479ebf88092102dd1b2966d97320ba056405404cb8d3a4af827
z86e4f560885c69cca469b3f3833f033347e6ec10954909e52e4a4c1c88a0d18681a7edff08bca3
z6a210b6313a3a9b6cc826dcd06cdf1a55cdf47084f3ace97d45391ad72f8e0198ca595e1583ab7
z86cff84f02da5c541cbadf7a7cebe746d9bd5b295652bf1b5f0ebb6db88b9d53ef279a07cf70fb
zfb1768e0c274a7ec1bfa1855991b255bc33c61d2eb1528f0de7ac3b969cec4ea1632b7210e8863
z6d0c92d5ea79848d708189d55755e43576ad23b1e7ed79da5a9ec6052b4ff8f07134956afb781e
z67b08813c8fe5fa97a4f89333fd6ad6fbf36b3e42f3d6de907171b1e0bb6ed81b60745489217bc
z914710f09940ad85729b4044f1ef2196adc22af1476c4ed3a3263d15d08fd309cf6abde368c54b
ze8c459bf64cf863a785c417dcf8bbaf8bd9c3dc539639228b3837657918dbdf3aff5690a3d22ad
z48b17d9027e09193983eccbbf269f3f613c5e6b077d5b82186943d64e8825f6eca4fdc64f5d692
z85b9db78d245fc25f60c13764ec5cf272a77b83b3b439b1dc434eeb6602693a207349cdbaa61f5
z25189b172f14dcc46ce4b0d780089b947f244ba1f073bf0d2a9b9baf82d961e6821a448b1ba864
z69ea805f7ad2c340191394f90e7592cfc4f0e30ce572e62e8eb7bd0f17222ba6459943bf7420a9
zb9aeb18445770f33e06ef84fdd37f0334433fcc307c48c20818b67e1930e2d6e69d464d7c5ec07
z54b34fabd9700780f8e47565f6f4455b494e88aa82d3ab4b43fb212451b69f4a90402a49dd409c
zf46d30dca863f146a54bd45955de0ab3d6a31cf7d8d9dad7b523babdb4ce5bfcdf7bf6a54f4522
z46c6c38f06e779f4a580693a30ec062dfb59d1f02e8e0a5dff7c331b026365d7a78cc2d780db98
zb309e5ab25543bb49680babac8967b1ecc616863e30cd2265b31e274218ad1567015b7960327e9
z1606ce2428611dab541aa0676c6aa662b991a7375699ea9d7bf81864aba01499361dc9f9dca971
zbf34f51a1692161ab47cd85a5fe14af2576ac5304a32e3c89ab62665fa1aeab78b2a228e9f1357
z2dbc1437a818374f402aebccb8c7294c9432a85f85d910125dbe2a93e1b270fcd178e3e3bb4cbf
zda6bccaef25892e11706e13f1c0338620fd1ed499dabc97951ef870e27fdc746eff3ce54f974d3
zfa353d8f0ef022be5387d2612d97adc591b5a908aebb286e3175a431a919f3245508d8c62ce023
z62b36330b6ddd340982e5e4c5821fd0303ac998c70b6598324e1fe94008bee0da7fa38b166151a
z5f6dd9a84ffb4c8a87e89d6acfb337c4c67f4123c139b1fb285faab0b8f45e1b72ddd648827c0f
z6f08e4fd86a4d93578a26e12cc64b40551ffcfd5bc7be96f3afcabcdf885b3738cd318af887a39
z4fb159b53682ff66393bc7e51a0d46832aed48005f01b23ec2b597b7e5da1f56583334192995f0
zb2d80caa9e090d3b03a95943dada2e17636b2bc899d087bdb0bd312111c9f84dcdb593c66d54e5
z9557fa4bde37b1f35b53f304fcbae9dd58330ad4589c31a36be2f22abbc8b7bc1ce83e240607e0
ze2d6dcbaaa4848615daab4f2df5591a2fd6359f8e2d3da7b8cbe0099867381773f035343ac4d9b
z5ea7fced5642f951daff6f3305a9ee3c2fb600b0c7a192c5f68089b2738374def58e7fbadb9fc1
z1bca8d76e3e697039481ff0d44e0672a7ae0f1b37994842adeee92850a181268070d4ac854e66f
zae25efb1d3b72f57bcfa1c1f9867676947394ef704beafced373615e67f7d7a70639b42aeeaa9a
z6ef6fac3d055f8e38cfe0865ad7bfbcbb38ec39e7f6052f564c3e403162f7f059ca31d872aa212
z78e4ca683f4e414a8d5d88e6c5c14b2b4efdeca47dbedc4ef1ca7376f1fbf66f29681d53856860
zaef5de7edddea0bee0a1b53457a44ecb76303d8828a99ccb3fe03d03e86c901222ac8783d4ab1f
z4a5247ff2067c22e08ca846a14668278ddf05e0ba8365fef62d023d705c479d2228ba7950c4d9d
za247cf02d2bb9b6a2ce3a810beaefcb135d72029e3b90ceae1fd2c34f999a0577146721ec635e3
z67b6c422fdaf490b10c5b09db441abc6d3cebf741cf8d533bf09a1c7faa083e28ceec665d3dd48
z7e332e6526617aefd6e87a9be12a84466d6565c638dd4d83431b6df855366c6d40a165375484a8
z62d0c2b16d831731ecdc1dab975f9af89c575c6c5f12b0b21f249ba45a6b49358a2f835ce5e765
z9de66ab222d620dcab6ac674555e1dbfdb7e2b41142f2372caef5f76c1cfef5454be4df5026e44
z2ca79cc04551e2891645395a4ff87e5dea1debbdd17588a4b0751e2676f91a6a61b03f28088ade
z1eb3f39f799cf61e771b954864c9112ae5ce16694488e45ff46ed60ce52e76ce6e229681c63101
zf3cf270c8efbb4ef6eafe053f75be0ab1705515244c2652e4bf2120d48f5198eec405c25408c73
zdcb315a90fd6771cd7d7d5968260d2331a8b8b50783ff0f6f783b74cb163e7b01e52f708783f35
zc541decf2b48e35d7683e17437fc755dfe3d0c0d173aa6949a2e8f77ca85cd2a9f5db776261d10
zef250280f582640bfd6b182dc17394bdf88d73c903e58b37571227989ec379f700881b7abebba4
ze41d12797d0f7cf782347ddf42de6a5cdeee8db5ff6521a31f0830bd10ccf00b9b1080cabad10b
z2c7b31a29bcc2243dab14a1ef0f47974ec188eb053bea9854ffee4fab69fb44670f55a78f44dfa
zc14f67d7e1e1fc8df30b3ad14affa77d97f00e6d4efb2c6b78120ee52e98483eb40cda34d212ad
zbe5831cd8c3bb8ca837555ee0df84c7664c77372e8e936e52aee61d19358b6407951b12e112c38
z1563b5159de984eb6a2ec38058d49871b5f03d6dc9f0c4f517fd57e72ace6db38239be6ca7b48b
zc8976baf111b76d9001119a82c43e696ad4a21eebe13b4e9cbc7d013d2df29793c83b33bccec76
zbc19c377bbe94a47c398f55bd9d6cb9cb601eee71bfbfbea357eb27d05f82242d4cbb146edb31c
zce663a191cacca2816c4c54aab3b0ad23ceb96c9871f74901581eb71157300e37b1a905e03a5b1
ze04a447f952e1c70d66a3bfb6c7491afe90c406865858309e5f47d7967e7d96b28e373115b65b2
z0a44fdd62417fa83ed8b97b05af5690eef106a4555b7130f4978edf8eed58776f9eab9782ec5b7
z9aecdd3d345fe9bb13e9e2bccbcba1db90ddd6b759992be13f9702b5c38175bd754d68191f1fb3
za010284bb5d038f7d534044b2e59d083e202a0bd050b8ca9ce13e2782a37f5a0cfab7a1c462936
zfc3d02968deccc905e4acfdbb41bfc8fd2c333aa4339aeefbd2104874630a5ff3ee7d8f7fba91d
zb4b70bc50ae84e72447373b5b057c52e467bc3318c50a7d03ea380f9d51828f908cc4e8575f9eb
z803666a5522bfab1308eea069c4b022153bb664254f7bb0f98b619ae77408fc4505ca92b9b78c8
zfe852f07cd87781630c22f00ecb3f86e4ebfa6b10cb8ab4243f57f0b92d2186a862ae1444e38a1
z8cbebd65322977a2a9b61dd2d1388566e125f0a45f6b378a9e5e296725c27e8cb4390585ab5972
z9824b8494cc168e478a8d3a1f4b0a683e4ee6741179aa6887a5a10fb24f540af69359bbbc1a228
z7a22f80df93029a0e971381012ef3e4b4edd5f17a08dff7dfdf33d3d5d57f5900016ba5aa3e881
z32f242eb293c253d3176348dd07dd024e32b340746bc2a283bb2ea1bdaddf4a37be07bb01f4d9e
z7fe5f2fc8761e5485b593bf03bbf2f997e834a675396313beae50d3f9197a81ae6bd8d541cdffc
z2902d95f8c73d46397f231a3e8d30864e59d7abe9ec1953fc7a6001a2c1d3ca9d375309212afc7
z47ff74d0527031d9cbd3f33848e84d4e54c01098a3e477ae04b6c5846d0c87ea2e4c8171420988
z4b0a1e78a182b7ec90da5668cb5a545d2c244b54592b90d4bedac6242e78e3778cec7db073a36b
z9647a36e09ab58c0ffe97fab4c2d9f97467c372421fba86f2c6479c464e3ce4a2e423d47bbe72a
z5ee4993de54a9e7579cc02eeeb4e9b40cb081fd6e4d59ef4ad1946524a4150cb317f4e975b7a40
zf5c8b12fb7d4b8e0283d752ae4d7d18317ef5c995a0582f85131f377c4bded7e81677266d4cdb1
z1c04e14345b451ec9c139479094ac5f138e780ed70d6e857560fb01ff9b1d2887b90ecac0b7f11
z40c7882bc7602d15241f261e03bd6493c880c90cbe3a7ec794bb633142095b6d83d46ccda2c1ab
z6ad2a018b4d0cb13448b86c5a819cd90b735c772de2ed3d679f451363a8ab84b3d976398d946c6
za0fbbd9f8b35a97ed79a059262daf72f5a7590fa85f92eb91674fed865416f7439c315cb7e4490
z155ca764fb19f1fe71fa4628219c14bb0d1734e76bad297fa9ded0edd1b761cf9afe48832f30a0
zc73ab50ca0ddcde8afea15e6ed60cc375c6974d0bcf11a52f810db3346c86b80632718a38f5459
z0612e18e38a9089834a3dfc6e155d9118aeb1ff4fe9137c506eab7e770271179237a5bf38db186
za6a6fc91d57b49517feae7bd7889b629d523c0e8250f8bf1fdcee5a155a93d3af68c88e1d21e93
z9ec7af5e51e1a961a51b17adb9a38b3a11e0c62375dd1d8799429b8d7532bb840c610ca1855be7
zdd4c6d684327b275aabcca0b5a53ec0f1f2e3cdc91fe43757926dfb08cbfc4e863b9e6fba2c261
z3e9e573558e0e9c53b530b6b3140917e92aa5bb82647cd48b263eab4b3de38d4cb5a8dfaabc812
z6b87f624f055ddc01f43170d1c3a0742ef2ed036eaf48eb60dd6a29a56f75cf0043fc8803c23c1
z1ab08492757c4cc559230790441b54f8759e6476c76b78c7df6c2cbd9c12ffc234ac47647c4600
z4e3df32b6738b08e2460d4d984a6cc2418db6f83a0890eb39d32a9e66f628978c6b0d612b73dc1
z9829c4a2ef4a33cce9daf464977ec3c8725ed2312636054ab408e65c0955b190eb0f422ff752fe
zd0d5657c87c9c661dc32025dfe5cc9787a13b05bb4107edd341774907fa58bc0847bb85f79a436
z3da8fc0d190adcebdc6a0037ddfe6dc99e2add9d5f84b12c6c5a71c7b21a6e984f3067692dbf51
ze96d1bf239d94a99cf638f6dfa40e2d8e1768c1e9b90008ca7d4515e8ff7514f16e3033b660b61
zb8d197446c826ec6021b201a8322effe2372ca1946465eb144b10f293da3c28dc3a5110be86cda
z4b4a504dbb89ecdb1653a7bb572011e7f99b8f1873ad28d852f3c0a01e91aaca87542de47d7e92
z582327d7065053bf5213cb60fb8c8038595173bfb98ae36144910de9500e459af3255139c830ed
zac095d7dceac9c6bd8cf097005bb1fb0a820f685cb3d8bad26a51853c7d2b93a2752a4843d029f
zdfa1b7054a7123ef8eb48e40e15cc594eb521f7596f6d606a948c2d3fe87a2a4f798c7180268a3
zb5528cee81773a4c42675cc7b55964186c1548062cde1c5ccda6bbd46758a2645bab3870d791ef
ze6cced379577a5920ba6142bccb1c2dccd3293f696dcf173b00452b51135578703ce9501da26f4
zce487b55623db4144b252081ce209f48975c10b519afd9d1d109371eb4bde8132fa51817e05f00
ze3bdb1d5d28351fecd12cc33f6a4a1793cfe4c54e98e6194d25817e12cbfa9ad984d57b1527732
z1fef9a7d2dbdf4909f751aead235fee6b34dd15c5cd1ad490cb9702f6f71c746b22b13525c7ca1
zed2ac2d11958d5669d5920faceef96d5dc249179ba85f9864e241e6659d92774eae63c405ea88f
z9e772e7b83eaeae04acb71123d336cd418dcdb56e3bf59c32f11f41dd4a8144dc45ba66f9cbbd7
z3534b34de7c640be0173142f2b17f3e1e18c13e506edc70e8a45d66e18c474c7c8c00f89ce8a0a
z180981ff62aff16a4aa6061d7f4b6e4c7baf693d4d17671eabf2bd5d44d7eca8f6e184bfd6dbd3
z6096aba049ff0e4078195d7aa3c3507c6fc2b40fc4f6d5a91b5a6187a9fcfff61d5fce80cd77a5
z9f59873f61362d1875f9a0f14f0775a2092d979225271c7d344f97e3356ce0104903280ba7b05e
z3e8840a709439ba64d49e3e97fda1095bebf2d40eff76ac9eb5d91f7306a82b8a06c7531ab75a9
z68f68dbeeca73a7bcb8c6dce2deac1808185b42a33a7fcffe629886c8c425884f03a7c8a451a04
z7c877f5d45065c3ef849b256e738ab6a715d142a69e80c3c297b261e48cf9ff8c176a1818025fe
zc2aed360c1d0083b7f1bd5c45aaf3e08f2d98a0392520765f732b65c859b391372c1a807704cd5
z4b6a1726630ddbd016674e19192d24904f80026e59d96cd0cbbcd07fbeeca5b1b83aecadcf3c8a
z8d6dbbaa8bdf4dc044af4370056e528c26bbbfa68f77a00dfa865a76ca706ff12ad56c1769e632
z2b11bb93a45adb8d22c61491df3b2c4630fd8d2bf6e0d709ac3491380b1c8d5f1fb605eb76f717
zf729d5d9cab03c3b4fe52deed32f4fa4ff351103161634369ca00429c72a153139079fa6d6e4fb
z173e853acc2defe399e122bda4ecf926d6d6aae931774333f5b5517c4b672bf1e02508b5b4ed8c
ze4d6ef1a34f03926973c327ccbbbb5c0b5fc081bd42c47491d8a7d6736ded11ac27bca2813c965
z5231fb319f475cdd44dc24a0010143315ab15878bf5b26c8ae30a911ffcf325c401a422716f6ea
z327720a3648826fad8d74f675ef6cc64035b7743822e1b3c58c143a079cec53fb07128c8e3c076
zecf2e00ccd11cdcd9915181370a19fbfa109927150cd2c557061b8598dad43d25d9ecc023302da
z0c038c401a2b6e1cbbd94e050045aa81701218fa6a7b0e4a4f8e421a88675c713fb713a198059e
z6abdaedbb48a28d17ea025c712f37d593f7dd6ebbbd6bba659b28a15a6259cd394662324df7e9d
z885e0886caeb9f51f31519acf0f1a86eaaca0b6a640e90f6788c93c8b8264b0102cedb05308aa3
z0fa693213164779877244e3a09913b50d91aff42a0a5b61ab89dbe47cf512161d53f7038384098
zd265d98081153bab4d267c6be713cd26db1df35db83a4a675e13f62b7be8e13f04c40357f13e94
z1468ee484c3c2c5145b3ad1567ce302469b0eee0898bf287b2698caa527fb9db61acf92d19b7b4
z9f42567a32a19e74ff053d00bb74dce2a5c57a6f850254a63265eb6440b7b3fd1d799b88f23880
z9288e9c2843a44836f62c0a4bd7c150a23a0519ea9eaa95223ac49aaeefe5bce48925405766a62
zc9005ed2fcf9e503d7354cb2205cfb31b132f3a96fbf81add9e434254ca6e377d8112685cccde9
zadf6813c999b913647e524d3af2ff7cc6004b86323ecb7712ca81469a10e39790e95826819bb76
zcc4b28d45d987a3c75ae571d28b2a764b96743ea358373d6b363f01fa91927978e53578e4aceaf
z0ec60505977d812ace19a594325e8d3f1048a10f6cf1f4ca0af803d6f7743c31acabc6f42c9005
z57e77b2b5c9a6d6f14f249f3c27a096776f642f84ba72ddc50d1fca54da2eb7d817bb07c21221a
z65fcebd8845b0a03891d082321c0b1206263ce71403e35f29409d5bce2e865308567f5bef60d48
z2f707181e005866faf496123ceb426f0decea2213471b28c87cadc02543c5d4cdfc0fb5679c306
zbecbdae9033de3cb06e90f198294a3daf64ac5c5335d81941ada1f2df9c8da19a8181d77a28cae
z54a2ade6b5799fb4825afa9473f5f1f82375804af0b295eb37820c62ee16922164ef530ae8e346
z9c35f9514a8f1e5e29f5ee89a6f0e21ae840304a7939e785a501818160aa95b1c48a819d5f5436
zf78c86701ce8d7eee067aafbed716a258268ddac4a4bc8be5232e608f88bd5773351ce44a8e5f7
z8d5587717017c37bdc80af62447be7146387279cbc9b0853f68faa10c360c6a2dd385eab9806b5
z5bb07f1817a4c73bfce57de30275013bcea425c433b5566251d39052dab7f88eccea35e6b29590
zc65129cd1268f614bbe2587b536cd384253fb5ee668703db8f163f6947ec72009d29e0f8cd9fc7
zd13f02d66a36ed0fbf335b393182ac55aca64ee55c650d60c01848ed428c11ec56ffe9f1b69c10
z1b325b512815dd256a1c510117519d845cc761dc7ed09a500eddaa331543db074cf1de04279be8
zbb85b6333e13c72058a9730cfbe13b5be3a97db7379f663fd58d3f4d0ed1c06c1b44fd29e6a385
z236b710b9a8bffd50c76ec17b23414832bc1bc9858a29a9b60fa9429f4a7545e619aec7c631394
zf98c7b3eb99722948ca1e04cacbaff14f83b95253c11746fb88ca885be1e1b8e37ce8a3173575d
zd0f2bebf1be55ab3387224929db4c302cd36cd4dc3980142224c4b86f1de4317c6a04dd36a37ef
z143acbfa2c220fa69c9c9c8068af5421bdf45fb75351f7016e439f78640147098380a408ecfbe4
za69edf7b32d72869b4609a753ad181d4b63f43010c0d500848b3f1adc68b0a08204b8c990e00ae
zbf799ea96aa06c7219e0571bb70bd62a08a82f740aa86b06c98cf67853acfe8141100ea25474df
zaecbe0979a6bdccf4d7f58f8c0376bf79c21ae764573d03ad7e11b0ca1aa2711508304b8e94bb9
zbf65d4535f78f967905a738f9cf22cadc3168e27981684ce842620b58154dbccee980aa9e2501d
zafd2920020d5d70c53323fc7444af0cb938ca050e052d1053e52b9e87e212f6114ebcc46ef51db
zaf7c59beed24ca92b2274afec26d3261a9a11c16a0f9a36511e48b843c1d95b89a6c531c0b4de0
zccda7d4668af3680753d41dc95c80c1104f90631fc6c07cd498a1b9c43422cd40b4f4ae53262d2
zcac3bcf626c87a0ff8f27b224a03ea7ff9aff3b911fa234562fe579385b56cd001119db2c9276d
z42962f08e077dc73726a57c2318cb133121b43353eda3e76ba14ca783b4538c53898bcd388724f
z8b2963faa003ccee68383c0ae75ad85b01cd25a1d382aae41918217c3cb6a9dddb59a8039759c6
zd7b3e67d6d8dc7f4042ecdc700aa9d7f8bbb026c044faf05c8350920ad62d56f046b63265168e1
z9bcb9a4b1dda4cddb93c2097a7c269003ae9b172b339584a10a981dff35ac92df559db6156ffdf
z59258818b72a999c3f5d7770f09f7859481acf641bf334fda7351f5640aa171662e1f1bad04ec8
z426b04a0c6a7806af839a21bd7ac3d11320289f7363a4382822f07f8d0eaeee83f425d8dde8b5c
z0c13878c39674ce12e2649d1e96537783dde685cd6ace5ec6e5fc1ac898db69c409a0d80d91418
zaf3d3f1bb8422e2e487eb321692789317228fcb80062d161495f75a82191032f22034acbf6e4e8
ze6d5b0e0434ed27f6a40f3e610f728fef9ed13078fade92c5e8867a1656633336cb1e581e71b6f
zce52bc25ecea0ca810c75397a07caa7e83cdee7c469eb6c176eab78648ec06c6688f2884319901
z4b1c090fd10bdbae9d8ff8f2413e70fd2ad86ab58ffaafc46125061c14d06d4b24e190aea614e1
z4c395b98c8b624d2373083fd3bcf4251446d5d118bbacf968bd18c05e1bce1248597aff5819180
zaa8b621b898864126ba5575b490bb6edf4d0939ad224f37a4a459615cb35a2600565d1ac4204ff
z95b6dda5c2158916c7a74d016e3c5fb0bd22720f42c6e54d8073594fac7feb1ccca70b302c54e5
z4d3fab3a15fa673bfa0d986618f17dfe1a90d7ef16d4da1f8df66a094521badbdab225007872ea
z97e494a7f0298bf26ad8540aed67c42be7d7a5990cd69466dc8f9d84f588fa01921fcd803fbc08
z94cbf268e17f88ea80271eee0a64eb0fa110afce33f293d7d8116db878b8b0b1c678ad5f95a501
z94b5c6a5e00f7e67fbb17b3029eba987dd440f9a56414d19872ddb94e32d2340f3906bc10269f5
zd2f84f2191cd175d2ff77f1826c2631ccfb4f0e49a7a91430ee90e4d2644533bba6875803735d2
z75b66dfe92930d52b91b0d0a8128d9312478cfbc9181299083839704a55ab2480591ba0e1ccde2
zc8d253615f9f32478cb7fa9e61f84e9892e153ea356ebc2f0cd4d91812a111ee04d750ded29ffa
zc11b91d38eda020dec4515c58e7b1fab7678e3c1e17b05cf2fe37d4317782a926d7ffdd3a2f425
z67cfbe9fa6473b90692e945d5d6191aab7de1acd14adc334913688a2aa4c5bf576b02c1775cf5f
z6b4c98b54b93ea4ab6d18956bbe9cbd735885a47ec7b3ffa138f36f271312184cad06b9b1aaa56
z9b809ccb8322d92c33c75b1c1a77a7942c0c1e8cbd25e43527c98aae95cc15c2a6a7b6e9a420f1
z9fe9df9de37b7e06d6f93901726ae93981d1746f1097a9b1376bd2297a03f7a07a8026fb3dea14
z79267856d94cefad7f1666f4e43e66070f35e771b30c2cfa046045160ff5e8af5c3483eb57cd68
ze605e0e9d7a27f56b45efded73d4e3cbe1a16cdd601aa0789d3008370ea612a5778236b11507a3
z5b5dea3ce76b7e865d802d992e90a57783e386d7d8bd45e839e47a3b1b385790255beefcd13819
z94dee2eeb97712a31a5ad360882961cfe4934295dee4085fe1291dfca267e78dd6c7be7728a54e
z47242e95cb3f334a115b02987f7f55dc3a44d9e1876e80e11b42599016f498790d8a4eed3dd8c4
zbfae4cffcee16166495da691d32fc8ca30f92df9d52b88be4d90e406d230765a089947f3c9f855
zfd8c1744af406cc0de4db421223a3f04c5f1f16a16a390e68395233148cb5ae80ee8333622798a
zc6350c62ec72d91e253e17ad9c3d80634288ec7ff33f0c9266d21eef8982938db49a1cd95359a5
zd040f972e4ef51703fcfa8145cdacc2d347c8ae8bef44431d130eb6192f97bc19587d2a69b385d
z7e0b65237beea2830321ff46abd54b39960ca718154f6f442bef25c2452af54f7344f2b5a85bbd
z4d203b4d5503e50882d7c3dab215e7a5297424f103629af2879bcca8ac25ebc8024bdaef06f5f8
zb8804b8a4fd30869a9c505bf867ff07da0997355b8c40ad1b15b47cd58bc02215addedca9363b8
zedf1ad28cd5346f5cdcf79f782372ab826826869f7305ff3bda1f740aa75c111a813662cc253c4
z22fb22e04723d7c1c8a4c150a3606db91f41d4335379ee6853af1119d9c7251a8539779de00e53
z0920b03fd90328e8d64d31358b22c6374e5a0a8b8b9bfaae2837659a5b489073c86904eb067307
z82e464578f83376501daec7bba9e0653e55c0aa2269da7ec14bc866eb62cdfe2cf02cd0d1070df
za90fb4572262a525ffba818abf7a7a7f4f3a18a6a562e6907331c8c2ccb9279e17f30a71cea197
zb5b2d817c7e17a933aa6aa5cb644b450633ab26c4800581ff88bf25302dc23a3d3b34a41053b06
z61ecd9517b088b7132deddbebcff180c055d0c4f7f7f0f2be553ca2614128052f143e75644f646
z5868441c36e70c534445aa9189b5c45293170a7db14bef6cd9dd295c7beaf996cc73ea1f4abf83
zed9e2573e893cfc986c90deb4c780dc79ee969b259f579dfce7100cc41385f2aa5b450b84da16a
zb06a87f2880485f10f85da34540b53914e3ea14c9373446328db7ffb3ae1f81d88af28aded7235
zb2057ef3ef4f354381507eaec6c88a15bfaaa55c593194020e303b79d63adfe39e66f3124b2a04
zf55432261ebc1cc1ccb842a0c518d0365add5b676676dae22cb6337dff2cbc0b7f368b3794c1c4
z70d470529ee2ea201e2e5f1135a7fcfbe44fd9bc7c6134efa48aed26cc4bc3d5d76623d3b25d95
z0bf919117c77400ca8f33370160f37b173c1dcd71805308f3412b036ee4299121c99e7b852363e
z5c2077470e0d42da48dc999b6df6773e38685ceb321d667afe58d310a713531eb48ac6569217e3
z2aa542cac35aefb4f35b51551a7abc0b54756d92fb4a8ecd3a3eba2a5a233c10f81faf8bbf68ef
z6fb7ee751e31036a451c7fa72b4fc85fb3c43021d6bddcbccddb961b4e426c00bd44218ff7cd09
za3d91272720119b5d9b21f1dc47e4087bcc836ba302318886464c3a830c4310804e4fb4203b977
z7e67c2dd3a6f74a7a2fb82b3414085601b71bb6e21c2ba27d04ebb21ef9b85f9bcf2eebc93b559
z99de49390c6b6fdf1c446a76b47f43c6b95188ee7d7de2f255e5fbb838ebe337364e8091d98e50
zb2bd79408240641e60ce773d7554ed5651a8e9f48921cb5f1240e7021c3f92b4692d93756293c4
z98bb41c991c904442a1254303523a78436194e208b7a9150af4bcc0e9a70197ff2a8ccd0c5fbf3
z9ca40ea7162ab7fd2f6eb1a65a419f73c8aca9e131deaed4162de9dc0d2dd460bf6ffad5bcc0e6
ze30adfc5cd9cf8f75e15442f2fb39128d289ab5960970ec0fa437a3e0f66932eb78067111256ab
z173152d65f446c6ff956c32e53fb0a4bff3e3c0a1b0118a66113d9430204721f8961c0ce325095
z5dae050eabf9660eb8ba3d84f73d08a004e8d7ddfe4dd21f46e2fff47912960dc88dbbbbc4ccf3
zcb1c3f87136b7a392cef11cabd8790ad60ec57cd39e1ccd71630e2f6589787eb1111ba65653070
z4ffd408cdeea6c49d69a71e0f865963ca1db6dd513575f862ff77cdb43d89b9600a72a29768e80
z9e8c681c3c605e55e51fb7e43499669d6815844f8e88cecb5884ff0acaa5fec838f63f2a2778ff
zda39c9d8ace1d0982022fc265ff5553d92fcf1b3c10080b61b7e813ef88c8990d3da51d3e80e52
z26e4ff44a22a51bbce44eb096368cd1b570f282f545083b8fe4998fdac78b1b9762adf13a40b7c
z6f7fa7c2a2c83fbe7039ed8e62e882f184414b6ac95f8bea26de7ba93c9126bc45400d8f7cb037
z7d0202835b5dddc2687f5b950ce0fc711f61f43a552ae36ab7804de3dafca20f33a008afc49025
z9d5711047220d887874cd479f5eb46a2c0ea523518a3299cb7261e85e54ad2fda100ab3fa32c89
z42bc0be5117d34907a46bfd8caddd50cecfb06e3459bc3577dddec1bf20487f2c288f9a16c456b
zbb26d89d4ed91d7726d2a7eea2ee0e37be2c46c3a66c0ad95022ed8e58e4a3f7baabb4d271711d
za7ccef36d20069f7e2ce6d3dca6f5ef61929d37f25162d6a7fe7d7abacbc955a37476ceb94982d
zc908367329f519051d0fed4ec8383b683870ec4251ef5764d41d62b8f8df9e083065d539dca876
z5b6cd3e0e8cbf7265100562c2270409960aee193efa45846e88de46dba5f919746843d3c00139d
z1937cf9a237638775122ed126a3b23ccc6de3a4e8a5222836dff35c77013f5618c1e0da6aba14f
z65a2f2ac0c31200c67d7eeb5b9b12cbc8b8c1d277e7a89e748a26c78d2acd52552061de964824d
z478beea2b5c5a2e01337f18aba6dba279c9467e40f26a6ece8ced0f8e25bcdad0cf78805783ca7
zc41ca70b68a0f7cddb8cd4b8e709731a252a7d36d3d3617d6e5206738b995c5da3d09010d310f0
za49985724df6b0aa5c718b10a260ce6ea1f6566db1634cf1eb1407dd53684dc2c4d2c86e412278
zbfaeece18eec11e4f8bdf1bfa9865d9e29cb18c4d7343f9b23a89d5d09bf4967ce54ffbde2125f
z74fd7929c164a16a477dc89aa822ff83141141734de0b2201973a445c89bde5cc80a1d2ea5f27d
z33156541cc71cbbd32f67fa005fe783e629a63e6eb5073535f52badd9ef78c818aba7a2af9b92e
zd0c9bd694e410a9777352316141587ce56a64f65e752cc456f585c18eac685184af25628444f73
zbe01ee1ba5cd28f2e260e8bb7a89347638b6d78f3a66e7e04ce6c2d95c4bd2cbaee69cac6abf1e
zecf3b69e907c20bf44eb21ac0013dc833dae2b145426ddd1221f0488cc37ca35a6107e149bae6f
z3b3136896be267f1bfd553c710fc66f61872ddf569786d8d18e8662428e4ffff5d45d6169faee3
z282d270c42da9e34703a0eee8bfe41fdbd7639fc355dbc14aef8aaf2d953c617b77de81a21f876
z6f8d1e802d409bea7d7f85a85c5722934ae2114bb8eeea11087536fe09eacc332a775ee0f5ac23
zd89f40bc84b508d579b6936e1472b8c48535ebbe3d69b74320aa511642ecf935c48e44e319be4b
z699b709db0ee77cd4761a26885ac5b8a11a1dd0723e493cdb57d4e4fec1a3bb6d04c7a2a946b4f
zfda4f7abdcb21ade0634f96994690a879610cc272cbf001b89ddc8e46851c4b64d245c22fb09c8
zcf0938d1ed74ea0fef062d8004116bddbc79db0aa1cbc75f8170e566fa2cecae663b4b0f30d4a1
z23629cf4d67d96d5f973318b699084a2f1295969b565ef9462d69f866262007371e0735c912e17
zb81cbd41c22a22b938bb1b31a037f1d9caed405a101c5e26d5ceabbf09e26a098f1dc0ed274254
zfcb1ee5877466d74471a54662f2bed6f112583bd94719bd748345cf9b8701513c51803fd07f503
zacf83e8ec0c678be1e58e47295d432915f03dd8d8f41a28b8284c10b237c3fa70f2ab5a1c642c7
zb38bfc80ed9fcbbf4e0a729de45d70a97eceaa30fbfac54655f292ba50892d2b57689405d8ea3c
z74b991dba349ae1f3313ec57f82c9cf0dc892ffa17a3c30f8d4e9e8fec071873a0cd1f0b628557
z9b51b70c5c086f7546b1a44768239d79aaecd7deec7235f88f70921da84f754e602ad867fd8741
z54fb479ebd05f30b1724600d5a3e95999a3fe6d3e1c32c2477c5ed84dc44c72d6dd3ffa545edd9
z9a913170575925202780041c3e027ecf1236ebd4b7bee7e6845a31b9c0ebda651086702678b1b5
z9d06b1f700bd0eb7558b3b0ef802e6277c73f0d7e46f16e44343b2187c52f3367d7ae5e1512333
zf73cfbe0f529b212059c95413627babaae577215053bd8649b081cfc60d550ad916f80622584f5
z80678f464f0b0c6b5b62b527bcd508815e68ec8822189845d7c20212006bffe6294964925386c3
z00b73cf8fa9eaea02a26c798c6dcf904b34ade5900805f287706c20816ac19987f829f530987c1
ze116c929b0ce12c414f1a77a853d2ac4fce770e49212d8b02ebf7fecbc4deaf6bcc576653d99af
z8db3c915e96ef94ac692e7b7c2a7273e13a22aae4ae3343981a75f3901593c9ea750e40890c7c2
z71da9d178d559650d68b05ff89694f7d082291f87eaefff3f9f98488d4673f0c249bffb7e7ba3a
z4069aae493fddfc2d499289e23b5adafdfeacb222b493127269dd2af11df58dd291f5a65303416
z49d97f643be33d39f3465d0cb1bb65b9115eb476c57c90a709e1473ea0854eef14f5163437ebef
z4b5d86be26fc68beafcf718b18d039ba7ccc22b731c7ef6a281072a27376fccaaf8bb3ba46e1c4
z340d52964dde20d56354dfac68916909268e8f010e45d9abac067745eea4b70a503109b097332f
z995c355f351f3f0977a1df02be803bb49e1757c3817deb0343b00e1693718b183b34b50b647f8a
z8c4879d5002430d8c0be96d80eb359402bd713a815c5a45bb522a5d1a6296ee1eed0b513bd7cf5
zb28cb6063e1f5cbf83b2ca23324a37cdb2d3a38b78e60216119a6e4b6d2b227118d3650de07ebe
z4e0430388f1aebba0637ab2ef5c4d70a877c86a741280a1627a34270b30a0ff099cc3522044352
z9151bbf3e3a030b5c2e2c0c9df257f070776ddbf83a5f5e8f45348e50e4dfc39b648b9a6103873
z6d24dcc7c7b61a078b46d4a38ab5436f8ec8df96a98e374dd7c8a94838d0fc1692609d52d152b1
zeead703a2aa169c41e393c34a842ade6b1296d677c9f195cbc6fbb792efde5f0fe9e4e649dcf77
z6fc012f3b6b6d0f80c6ad2daec80fe73a6e50ab01ffa344bfa52266c65bff4fb2c82293d9ac30d
z27a646c9a32fdd015fdc121c7bde802aaf1d0d74c77cc33f0650c9df732979dffce287f0b97db0
z74cf7911fba5b879bceddb92b4435252e48ca0433ba257ddd2a4cc7e9a4d786a028f01748b5f30
z17fde968bbec067256f8a8fa3341154cbd29ea73e54098d501db4ab5e19c0ec7c811b5534b2b2d
ze02907cee230c370b0097bc393179e301e900d3305809b31cc10f258311827435154e7cf9f243b
zc73d1fcfc2345ad09027f03841bf4de8e238bade63f9fd4d5081cb1cf08c057c8bfaaf583d787f
z682cdc2271b3e2d9ae5ac89fe3992860f9a4aaba797bb64437ebe2e6a716838d0b5d21eccb7e28
z6eb9dab492fb743766905b4964b08c5d438e7dba1d5e34a9f020b7caea380bb38ece8d40c824c6
z0537e5fcec494496ac9f2136042db3030247a95dde2695e554ad298a47f8a23005e74751fdb769
z565102d8719af273b3b66167e331d27d5d35b49796bf23e94052e2c3bbb9ad2e9a05ab82c861c6
zca8356034e875467c731cd6c05bc54e29ab83fa4f9038a94288302d889e9ea14c2477a05e09442
z1810b4bc31bc6e6abe08192cf601575dd0cd9bde72fec66abe2d640b3c5f1a4c051db04b08cee3
z5560884d9c25d721b17df3e89c4b1b513b1d8e9c6420924b2b95949b98cda5396ff914226e6296
z771518ad1bbbf1334c7c63bac7df3a1f429cedf50f15920d865b3be13277432247730b8f483493
z296b0b8339e8d5c57c0f289ffb65071e1dd392cd7dc111cda2978f7a7d19cf810a7a97ccae8340
z5a27c7023b07cc2b0e44b1c3f4a662f730d9a0c360aa2ce1df7baa996e7d7ca7f86f8d7af5a3b5
z61a2b228d7cb8ee769b1562e77aa01e3408f1ee723d94cbce21e40f27253dc82b5955ee7dfeaa8
z3b9b3b956308a8cc1897f78ef2160d8460a2322936fdec30a491ef9d9eb8c02fec4d60cdf88a0d
za520208eb89fd6dc11ea3ec400b6b444528eafa2321085fc8a10fcdd03e1faab679df103946aea
za8aaf35006d5269a6865aba7d8f61757618d7a0ab873291107c924080267cb934575858384fb96
zc7170a72e2e03b7c7356e1e22890b802bb23241fe02e9e7e92d0735e3aaaeb0dd5b0e95f982b76
z750918ba56d9ecca02ad059e04469ee0604a96fa846dbdaa4faa4be74b7656e667238b8c5387ba
zd8c953c4323074596f16288f84075d78d5ec9cb182f8212f76d7fe4b15df10742893fbc0d96a6e
zf83f6351e4872fcc899bfdd0289f425b0002d873a9488d7ee6fb72e631dfb0aea43ee599099d4f
z523fb60cce1a5b480f822d06f800a303405c28e969377e970c4b563a579b989ead1006e1b07fbe
z4a6ff4ebd50bbfda9a5774d82c6a5d4022b7ebf7c27a33b7ecff1759a8f6b0490e56ea5dd376c2
zd528b83cd30a304c6dd7949e72d7a6f9a5678c59ab922d6d3e7ba6c6df3d4e022731f43fb467d4
z0f38c8ee353b4dc5bf41002c111c44e6ee57e238daf8661dfe7b96abaad29bf64c3b020b747d16
z455c53964c10d71de884a34427795fdcad80630839504e1ce22a4effdc8c23338b7e9a8bd5e3af
z6749548b1ab60550de4d75e5cf3461af8ad62a13bbb00f00275153995b7ba511507c8a0f76ac5d
z5f650c60d1826ff735c55f7fc72551f62166d26e4622bbab920daa9b609b6c39fc6ff52ff5fc47
zb4199ded11cdc6743553ee2a789506081268d48d1a6cb822f7a31beac7350c24ad5e1063526f24
z408a97f20cc7cc87377b17ac90cd992e804933ade0d1302e3006845e994b6381f50d0856a37f78
z4ce20bb709328133c0bdd58ca80ff765c33411da47b7aa225fbd9ef5ea600ce601e4ca6b3ad906
z09d9fd329bbf393f5e93c9a21e653ed8788c0c071534d62b10154a8d7fc94e0fac6f160c060d21
zcdc07effeef4a08eac75f285b5565468a0bfa18a3f3238e8e14ee72b7c05fb8bc3f66280567361
z843386663e0a5823b8fefa962df638e2e49fe18ec7a94725c8a95f6f07b571914d2071b67881df
z8a97a5216145940f24eea9281050af07a356c88035df1f2ac4ea71a7dfc4f0f9707cfd3eadaf9e
z5fee8ed3570bb0439561eb4896f1e53573de48333ea21c35e8152d203b98e00d2b7f6fc7d79383
z103a164024d32e3840005deda9d9bf57e0f7810bd039897b1f4da47bb0263f1574fbd2487a6605
z0c6b15381731fa1fe7ab2ad88b6791c8f9661ffc6d49a0b16a76974f6c64362a9cc0c76d0748d9
za5bb930135edee59f107a278801d3c07370bcf60eb70639d6538bcb744b70b2949c382ead3efbc
z2fc36805a713a49007fc8569e6e6ffa258f01931404ebff1f3103206e6287da3f29792de17746f
z8f954387496bc49fb3877d8df49a2637b8e62c6857421590adaae0e699851c8d8913cf2ae60a27
za28a22f4d2f1958bcaaf58166f65ae7a83f30eb2fde2a6d59d125dce1fce115b26b2a7a2753217
za71025d2248c30002d34435a60a4dcb384baf8aeb1162019018e44019b9efd53703c846d26fb6f
z463aab9f8a91acb8e4b31cbdd1e2755435a18c129a583953f1211403b531c9a28cc8a418b68a01
z183a443bb389130ae1bdf10ca7944db983448b286202d2c9fc1b6ba7a6361473fb4c9ee8d7e575
z2f2852fad1f990f215d32ce69efdd5f8d22290fc03926d98f5f8194a21a754212f1046e215d2aa
z821eb28f42ecf284af3210feb91be935d66ffc19f78f66104192d35c7006a633cac8e51277b44b
z754f82bfd8b064415bceace788f2b7f6fcee873a2a795cb622780aa34e8942dc4a637941825f52
z4045edf33551a21a19a4bb49b7800d80cde2784f142e11f1e010d0980d3eb5330171e936c1ac75
z6a4a252c915b0ebb9d4fe41ef000e35d0c591b38e7419b9e94b6e59435dac03bd2cb8bb4b63818
za8848e4a325c5f4c53b4145a1e9354fe8d42fbef203c5070c60eb5d1ed241bb25df1b23ac245a1
z421689a207e79978598c2d30ccb7a0ad281e2dc4a57663a117ff8bebfa0486897a0bd05abe1f31
z62f21509453b0bcc3dfdf23ba899b7bdd9bfbe001c2acdd435853cc1913ed98b8b62da8da04954
zafdda037c7d0607679ece66010fd34f5cf94e70c8d423c52bf65af03d1f43f62720402962497f4
za44f085487235f74f2cdf7ce42d78e987073b43f0031ae0bf2244cf643532b052347ac0fc5bfbc
z948428310fadf04cdf390e44da2caddbcc072de1fb68f3cb62d3543646ff173072d23354b50dac
z59b3cb90a088227a22c73291f2c6bff97e11a6c02f12fbee15f1fc1b470c39cdc8de2308c2954e
z77e91971dfc532daea7be71a889a497b4cff8c897750bd453169cb0aa68cd88ea1633c20ac8190
z446ed6d187bf9ed8b93232175d6dbbda308a2226d89a89d444f15d5ea1550c00f15550193672b2
zb22f46fb1da76227a3dbcf66e73d2d8396f58c24e97b4ce6cf5d818fd8171b968ce1eecb6327f0
zfc68082de06b860ca6ab1c18973f74b1c467be81796729108a57795e60eda98adfcc5c5f0ef551
z5d518356e2a43efc26e80efc493c368d6ddf6564daf4cc1c2010fa651945bfc8904890f0a1f766
z68e413cbf58de2fbe97ca0b1fe24cdfaa86866d09d65e8e3aadd6653ae2adbdbfef8bb7a63a5a6
z4a060bae9bd5ef1da274de5371e44f4adebde142819ad12eb9c7e77e205072b284fa01f52fa43f
z8b1dbd7aa9df249132cdc69ef906a9975e08d575a5a88e4c5e813fa653062d3cb5755281444e33
zeab80d6f885040e17863ae19722cd40ceea8b9c398f88f96a2c2861d00e70174e19efe31069e77
z1e251bfd747f8f2336adabb9e18442da9dfd7a69aec75df7f1937afe73116d1656b3d4ec5df5bc
z8de4b3003f9c7243c3dd43ee2202ddc062282cd10cf9ba6208880262b21516afdbc33c3528964d
z18c9ebfb12ff494ab4cfc18d7c9095d19ae52ea0ce991cfbeb24063b3cd9c6d09ac03def4c40e8
z91679f95cb6ddea3beb3508c39882d69bb70950594f4a003c28d81746f3681fa2c42b1a15d7a1e
zc260d518cdbbe7a001e508757ea07a9d7c9bc5d5c9aaec45a77d66faf2efbb28cf49781388c179
z4f3694df2840bf97f78099d0039eb9864e9b1a104eba184b0c9a7584b35e6fc544f5f3f50466f7
ze6c241d2c68f6b52a9348909beaffaede100ba639bb9fe499bdaa368b38a3ddee04d75f77c5bf1
z2471f206a87a58d8358e5307e51e822b04123ff1f8af8ad1d1f1ccc52eb42f5d732901b629472f
z863d876028ad6e7b0cfdeaa0d60e02e0a125b69e1442e345fad5cdda08e2a60c5aa534bfed1176
zec7c67ea0a141c0082770f3a6acb22f6435be60a514d7e18e878feda4ca72ea5f306e2563f0a77
z0b150e74bf7620443f66e8e054f4dc303985df84c779c0a394ac06998a069032a0f8e8a06277ea
z9e1a90f0cd9b3a49b0132802b99c96c7bdf25682bf3db838b8314141227a90fa41a41cd3a19a16
zddeaf3ac446b8a3197958b373bdf2b10e1d33e3e2dca999c81b9052e6bdc34e04fd572e9724fe5
z947187dceebc1c2b4c276f526f15b7e851db988710d348acb6398be805d1780136cd26f94deb9d
z8d20f8d1ab61a946f561997d3122f619553afd2d6d1184e7c245f38e805bbdce059464daf90c09
z19f89ea8afa120ddf68a974f81a7b1472352867d4e98aad6e65503d3a09546a98b6889dcc3f5c7
z9da5e76040c434675292ee44442d68a17e39900235011192b55bcfb6e96d06bfb3916843a3f8e0
zcf6b7a481e9882dd02db7703b7a8a0d96fddf0d63d675b41e727c33b42d7b3f8678f3c2ddffa37
z5c3b22ca44097b8b45883a4481813dfd15e65b969b4e9df4899c3e6cbc43b5f54fadd164efc55b
za00388b7e6124985fe356573d6caac3794aa6a712381fe0538276c2870203767e68d4bcc0cbb76
z7832a475adcad8318f4d1601e8262efffa47d8e8e0a19d731a0daac58691286110f9d83a4ccd3b
zcd54b714a07fc426ada9cdeb8e3a8f3e5180429dbda92cfe4dadbf90683bc16ff5396f0f402eed
za59b4873e208dd6da6fe703dcad26fe605c03d38ed5d622f074fdd6f5a9fde7659d0f437498a72
z5ed25554faeed866336de9b80d6ea4747639ace838207d372595e409eac5fbcd2a8f7bda25d3f4
ze94e1e9ae1ba87500739081623001429c9b7a58b2c37a6a1cba05fe743b1d5bd89e90c679cd8a1
zb9467a7ded241dcd0f217c1fc05a087f47b015951746f31ef883a0f7e0f45e48b0442476f1fad9
z7e2ad186494b54342928e998b68e4fb0db113e198c060b48eea666aeca20df8116c7b1acd3e6bd
z91de3946918dd55eb4bc2e3635b12bf52111e0680005f102f271908e39a10d9770d23ba3c78eb1
z22c17b87163798b331d56878b3c5a2695dc412978515642f72066cd218b411139fe8ba0d220d42
zc30fd592a55af2f7a42a2fb0e82b52e704b888dca04a08ba05ebad8a9ac3c964a56411de1df8ac
z9b0e520d6828d91d41591d5a7e298089752b97c003c673e145a4a99af8a14226a16f78a5c115a5
za10f365eed8d97163e37964301eca94e8b24e28f178f650ba6f835e614e06c37a464901273ca14
z6d82498256208ff1dafdc1ffec09f62b7adbdd3c26431822288d18e7d7640bbff122aa86841feb
z42265552476f006c0970405add0063065382ea40cbc8530f621ffc972bd214b55993ce8365da08
z3e09e239ee0c16dfdca8a527822c44cc5686f7fe748822839ff69470a9be77a7dd0655cc962c62
z9670cc93f6099e1f444fa6189b8667baeeafc14239f788bbc5b665dbf372b5e9a6fe40ea8e1aab
za62d2bb4bb33afadf484365af3da88aadb191afb894cfcf4c530f0ec3f2d7c45ed757feae03671
z9a5c6d04b56a5de38bbec57f5d7b6c8a13e491c8035e83517bb21f34dacd59ccc21e47f7c7ad2f
zad750735e484d82dc03ce5955833cbfedbef0a6460ecb6f67b5e1fb7082ea114326df497b302ed
z2928e24d3d051bd72d3996486f6f70c65d8a40ead3c8199d3ce43a6b1ce611e41fa0d8e44b1834
z439da7385102ee65332ef1e1fe83ff5fd7a8ec7db051f519910d15f5372392db2e47a9cb1c0483
za734fd8a861cea9bf48c348787085c15c63a6d7c876a5e22fd544944e37ba5164ec6ad19bf77a2
z5abb2ed631c99078b8bd97f5cebc8505cd806097d6bc4738c029902fc3dd749f0c1daa606702b2
z429c459a57e838e581611ad8371d9e0491b513f6c337cb21a1ed1daa0288145ee05381cc34436d
zcc2ab751f3722a882c1af733e60a3656cebe0e49fd7d02592ff8cc66d7f44353c50f296a3cf989
z5ff41cf7b7ffc572dbcfb765031b3e13efd71f255de1b17e97b977e00a6e69680f4082445da20f
z119f863392f6e3c4ac3418618c88c2fe8be31bfbabba721c2b57b3b2b57d8b352d69473bcc45ff
z41673f0db0d85d6662511df3aea3c062d1a99d868df1cb7b75eaa3b2598053fd780a897d329369
z8a8aaf8f3b7fcb3c24a0ab62afd3a30c78759dd1c38ec37ba3ebae846c82cf093b665560822b53
z251d6ad8dff524dd1a9ce66ad4ec9e0baf37ff4e5d7317677aec257cd7c9b16d46b86ff4841555
z9bfb1e18415d8bc741d8674f358acdf013941350c19cf8dd64d0078d993cd44aec734274d49743
z7b3e0578c47801cc9be788c8870e1364f070176e44a9d24bfee401d73ae46a6e0e0d896a70c102
z661736ca09e314b98eb7ce1b009f0bc17b35b5e9b080313587a6e88f11e7e29e0689a122aabc0a
zabab2fdb986584dfa982b814b8b45c6e496415b5e0c76ff16b0c7341dfc99b5a93232fc7ce8922
zf0b8a3402513f2edcad162160c2acad946cef795030e9642db9e2213fc0f8f7b762a3afd2aa1ca
zb9bc2194a1bf0b949a4d6f983f0c0d3a6ae5379fb0bde62d7fcfbef79e4b20c47aa29d6185928e
z32a65d2bdb0a0d9cbd583eeb60cdfac5d84a830f56f16da20159db61d6c7eda772b540c86bf4af
z68a4174e5457edfda31d91dfc1e4269ddd3be19bfd49bce92621aaf5d8e87ec51212876e2522a9
zda60993114dabad605cb742b54f4a8fad5e417ff09cb738f2754b5dded135ea87390d9e5c5079d
ze30471360bab3f18eb586c8de73f18e457474f8fc23bb3175254d92405793f90adeccb5b5796c3
z6490571fdbfec9c1f77b0a2d0f1cd4d7c7e8c2e5edcffbe52538050139f55656e0da90df53802e
z27d8448cc3ccd1e6b2f59392b0b02e71403238b8ccd62e76de0605091984b1391dd1e7f738e94b
z0b7631477bf5a4a338a28f5b0243736f3c9227f83d10b0070b6241c6c7a1d66e4af0052f936ab8
z610bf50afef61d19365e6cb176930e354d727e98cb928c85058f5ac9a5ee5701ad7debc1187eb9
z5130e363205ece6c78317b72fc8ee9cedc9629073802ad8bca1dd083997c6618cd6f2aeffbb238
z71fe5052e161497f41b12df35d42b0d7bb544c3c1bbe3342752f37f4d40f6f35a9ed0adcae2f9d
z571d2087df002e40032b5514ed14c1424ab572bba55e50cd860716aa720dcb755ee8536b4b42bf
z3d5a38e2f61bf5f9d9d9761c1a908798560ec2e12df926bf69a36084a27724e499a273ebce05ec
z21d89961391774ebdd30b42e89be654951e13813e11247e1e288c7d8fcc6f3194a11c030016b1e
z9a35cc4232bf0c1dda14e3249f3e6d71d891e50be9c7e40ff76a7a7d03474275bc43553ab399c4
z2ec7800995f77d623b0b52cef50fdd643d39e370116ce9aef0b593e12fb67c3cbddd1884a2b2c7
z36f43d7c7e9d7882a58c067dda0614ab2933d238b3062046853c3f793068f6e35e29d18bbdf872
z0580ac2e51fa898ae7b1b4ffa876b5fa4da9da04ed4cb01e158b40b96288087c2ef97d2f7f1803
zefd897cad8c234192a66ac3d67833fb9deda3cbc890130b87bb7250daf2d7a8cff78b9f2b75ad0
zf2f95f9b17c78de311971297be62a98dee27f508a8b825cc52ebbd76f85fa69bc5ae0cb8e0e4ab
z5c67f39c3a69c17dc5d5171dd1cb167119de610d30a653cae9295b8fdce8febcbea275adb47f2e
z793ee36eb265fa69a8329b87017614d11a74f2d7efe2b5ecb9614ec856dfb5f770d5b7b7635846
z9a936aa74800106a65016377cb43e6c3bf26bac77ea62f24816e9629854008361f4418b69ea693
zaabe0d8cce1f2c5a4738e4367e50efe0df7071407e3a9917326094ff7e0b2bf3abef9b3506d296
z4d6253662b867347fe6b0d7703a94193ce57c6d37c5e86717ffc5648c7a47f53d5d5faf269e0af
z745eaff544522fb7ca9b73c8943be1cb193ad1113f56afc35124672b0a16e7b05ea0e22d192411
z6ea2941c9a8872bf8f778f1db584fe29d3228ccaf75e6de7f8fe69b957b3cbeefddd6c23c5c841
z1375686e5880a39332f06b25e02e2eb94e000fee3b80da545d8b77d53bf51b9795027c76e77cbd
z22772e00d5d3f2e50f822b6ac40f4007357a97b3535ff473e609f378056ad4c31c9102ced072d3
zde4e3f48a8de16bf78dcf5745bb33539cee40f4541be77f3a4ce55adf8c52ea66e0f08cbd49e0a
zb52e7031680fe6e102867ab96efaeac0543ce051f7523fac0c9381fe3922b2061822ab082c09c9
zfd7b17808d91cf9e6ff3113798658fb8646414e0088d1b058287c0c76120f1d73c69d02ee28623
zc2437457c77903a3cb3d6f961c38bfb586406e140e2eff815889b2963c513d94bd2c0f0954d8a8
z8381d219b044d29aee6fd6c5dc7d1266349afe526f982016c0a5e3890d70d37babca3197bea7fc
z4050b5868aaaec1cf3c1633e42081655d66d7ee774a66f4e51d92811da86fadda01da11682d54e
zb4b93015e558c271ea16528f3df688622b3d9456e85896073eb2809121d4b3c0a9caaaba1437f5
z49995d6d96c78c895acc2765f59c90d99b08863ccaf4cbaf94ed7aa2c744d1b22be394abc6577d
z64f65adb16bb4e46e282c2529cdd04de4743483df8c7000d4728337dd0d43d1233a7a1642d77e4
z9951c8d6f2e040e03559596681fc6b95b8e08f68b482d682b8694277102591b8809f67da9f6d22
z83d65c79d26b60a5e66d470a7d0cb9f6ca33807b4977b9b059e0fb1a44f58f9f6a815674d9d781
zacea878ab06f4b26b68d342d410d4a22098d5db804046aa1f26551b7fbb2d7d3f358a9c6eb9dcb
zc5577f4ae7c3f0f2a23039008994ec048e86461627170285afb8be7d6471fbb4a9c997bbc980d8
z3ed7e97ce1da51b5831e1b26d5e9583f56316f5cfc9ae1e4ca379f185bba8a62441ac16349d900
zf7cbbc4824a8a9c097819239b2a4050b63a2b98d78be62f9cb314d2d079de320f90fb511c688f8
z6225ab6bce379a3565f54f6e7b48794bf2544daa0308be1327712cd2d40e74578438bd10d5e6d3
z7658e9713864ed50a4d51c8f74bd1627dab2e70ba9c9e5603160d368a7ca8b3d5d1ed47a4a4785
zce9be9c5103192e8d92b5e8357a072a0e6259f3e8894452e13203b6ca6daef0b12be4c85516873
z3e03e36b7fc48d51db16f731103676a7ffde6a6a56e65951f375e29ccfea68706d3c8a0aa057ab
z9bcd4ab816c55b4562015ac5c2680a9fa67eef8b459220363a6daac32f918c52a001a84a402cb2
z6888ac5b424a08db9aec556cfaa10e30aa3425e9dd061a23dc687c07a6bbafbc8b133371a83357
ze2e8437f16e7806f7e684a0236c80c52cbdd505631af330c1579ae37e1c0e94efbf56839ec9c55
z39e902638e8b92b999cf9156c801ad1a462ecc478266ea6b569826c51925f69783db1866cd5ec5
ze717ca6f3bc529771c08741cc90e5b4baf122675a8f7645c5d3af43622713a9a39100d6cc0ecbe
zbb7817802ec2c40e44936bc13d97cbc1d40da891daee92cd6647d81ddf8ccae74ad7ca6f23c663
z4d5973c86c8411a0595fe482b8ea797364b0b757f264a180b82aec3ef4f0791b54c32b9aafbbda
za95761e0b3b77c9997b0f2033647bb049146f0333dc0aaeacd716dbffda5323a8a19f77a3d914a
za132157690ec83e2f780d63e3f9932f612a86c05ad2db476a75ea2ca58defdc48ee8f5d9798dff
zb76208c2a0b48ee9a3a9aec25c002c8c99d4b4237c5dc8110cb6b9c7f7ea1bf98b71b5ae7d50e0
zbd39fbdaf5f28dd2df1afdbb70ab7c8e6d9529ea3b1c5e10d74fb38005593b5d2451809c513aa1
za0f93714fd89f75941f2ffb0fd6d560cae10bb17ff7ddb5b0acae05f6af112e20c70a8f731da75
z42ddd5990fe45f38b7cabae1999d64878f2f0d74a8c197c2b50ba6c3eb4a9e5a8956fd00ed582b
z34d2d88c6d006adf1b0cfe39f8455b9fca35aad8b39cff24316567dc34499dbbf255e973306c8b
zf31bb2e851671b2259aebcb64da6e12067ba98a6e9b58749e61e58adc4e6b4b6803a6424008bf7
zf9e1bd50f9858be7887ef8e2a4a0f7b2f0ffe15bcbdf9740759c18fc95aeef8b5df1959994be89
z0ca789ad24fbcc99fed2ddfd881042124f28525563ade484b7ad707c7656bb557eaa5f3af4ec60
zd0a809ad5f0a77428da24cd799a8f30475342372f4def5bd0e43f2775f98299c224f5054d80a4b
za135c8264c06a554592fd027a8366acb30289fc949ba1b2c4a0ea5ff3cb9aba1f85dd4624b5403
z3864ae2031d653f9ecba64fb9a1f6260e023a30c035902e2f4e412cfeaa21ede2f22f2757e7723
z28c4b9e19f28b4b218a97b7d03f55fcc0c954c0f60db4323720145c6171d362e4be5ad60df7c57
z21d09449b489797bb7c0f1cbfb671876d352f4b829e8cbcadda3df3dd21fb80f61a795c648a28a
z4fa6531702842dce89f7661541e21dc632f5e5a06f316821209230ee8ffbac9fc2cffb2d9d53ef
z272228c5bd923512214bb07bc6b22c439dc9182f377129ce21e5aee8f2a84104193006b83fdd1f
z08f4e7fc79484972cfda45121c0d4273b8553d76e7cc09c942422569b2e2b09086324d4360eebf
z8f2e9597c8a23bcd3ea344eb2ee3ccb798ce876d4dba9f4ce69396884ee9437b475c1d1b651652
ze3578d2c87d974718d875eb14d2ab9b26d564c90b16dfd62b1fc5acc2bae51e16fb65211085bdf
zf4c92862525ec32251758977efdd7d07053453153532950047f3e3c6588e7d9433122b080582a7
z65b0b27b3ba677b0ab34b15a68ebd1012adfa51b27f279deb5cc7eefb9e99670eddd2cad0e5896
z0c50800b9e770aefc0d91d687827fa5bbed186efbc800365426099c0fd8129d3148c7ace9f2b1e
z50207020a53ee697ff1de7dbdbcecb4566e5103f14d03c441e97f1fbc8949010aa02f9f1f7184c
z73e96b5af176a25032569869c89ea0274b88de9988ceb5d0af6120a2b1a0cd384044a408458e31
z75ad4fde69bc2ea8749740c1082f9800c75a0ac6e3b7d43cf19d9e658a197442c5e704e9fea11f
z7bb0522a728f94e0aadce93378a5871a230313a462d89d9d62717a0a5e4f626d69e0dcdc1ffe9a
zb7a50d1b6a9dcd74f7853c085568990265e1c4bd852134982e5659580dfc176a3ca8a5449d21fe
z9368232ee805ae72c327b4a6073977fef56cd55ab3288024d62ad944ac88a756c4a22f1eaa17de
z59deae5e6de21a88aa7fc73f0e388762162d5c04a54aad95386a8fca5df1e6914fab619502fbba
z888a3963af754cc4f2c53acaa887b78663aaefb9118284266e7f9410b0b25f70aee1c7a2080738
z05b6c601280ff58bb046f1a2d1c5dd956cd68696a79659497fca19cdbd74040af8ff232c1b3671
z6ee051aeb0c2477ccac84abb393a83db89cd83c599db9b2fe30395a0ff5e04d9c32f6bcb219098
z5ee8012c78b6ec77cb36c9283ece2dec023ce18465f848d281edbba3f1ffa13d5e4002cbc6ce7d
zd9ee23d41e5d7a0eb811a7391b22b7a7424c52b2f1c310f8e60e99e851c8a371bf81d84d3e937f
z47fb6c8773f66b98f111e782d81ab78576cc21d09917ee66f410c35fed0b5673b2b01d86113265
z80a3a59c27c1ea74375c5cf2f0e8d9e10e9fe7dfaaab6a359e3bce66c7af716d92d78fb9a3711b
ze53e2e98035e1ba18331c482517e603060e4fd9e44f9f107b6b9ca94a1d09bbf54b2bf7cef5d89
z81b6a4e6440bb637acd48236ff4f88fe63e5c745d41ca96da2b2ee58cf907d8e6bb86f4d618669
z67f15070ca3602c7a2da4ea08e96981b2f43307639224219478f7fcbf31e2a3d0bcb5a629eaa50
z0d4c810786db3d6ed84a506ee9a6b05230aa26da7c5d545ece978e5d9d6803f170076352d183bf
zb829a67b7982393692cf2dd7f2ca018afd834c6b484b41488f9dc6b7aaaf21a972890ae9622f2b
z04aeb704e09000d3906d354eeff00610338b694a0ec8a02864e6a8a7c5d71c82a03fc74d29f2e6
z214fafa6fcc24d02e228889166ff5370a2f6b2d9566cfa4ea61f803733482a544110b5de3a06a1
z4ed6997d1781fb4e30af8a4e7ed4e6874109be15887016c902c1634b61bc3e2f5fc402deb3d5f0
zeaafddab9ba678d8559c2371cb7afc21b12938b3e7f2494328398e65a19fd2e454711ccd0cd9c4
zd5b646b14969fb35e95c6ef44504eb8c4c75109302a0f28d12cfebdc1eda71d5c41fe637c22c44
zbd8f9d7e6defb06857c7c96c639bfad850e73927173c57a7fdc426d6b3361939485d9f7312c1d2
zbd90241d33a36e4eada1a6ea3294cf836574ca0c0fd8145038c9a3a22f58fbbf00dcd093802dd2
z1fa65f784ea4f04aa643cded5f04cce62247d5c1a857f28727640adedfcdbebf509d4b5c82f9a1
zabcb2fa591d35e546c2bb6db8aec82af40c730b08e4c49ce044fc70bc04bffe087070d0d2cc243
za846bab0534ffdda3308f91770121251f10d5cd34bf3a1b067d64112f62497b72468b49268399f
z0b886c0a5f9490081c2d96c2aae29602ffd450915b7c16c4301b731f0b35f2a3117676971ebaf5
z511ccc3f5524de423605975f8256434bc11beec2ae7282871ad6fbf1366fdac2c187269fe160f9
z0a603eb2c90815ef29bba544e45b02856c7866c88c49946e3dc4a998c8d25c664c898427497d9f
z18542cd2887b5c3f898c77c32cee42446ccdcc01b5bed619d7a315066945d13036337b948c9010
zac791ab72246e9d9df673c4aa412706554b43154f0afcabb3bd4f8fed801e44a4a71fc00c448d9
zbfe881dc4479966b4fdf229bbd880c8f359082b16deda5ab273c7134e2e415209b18de1d0e9138
zb761f7cf9488088ac545a709c231469c169d930cb8054f0638b4a3b48e2af5db8601136608b948
z20ba5ca70c46e7db867bc7f133945e85f4c7dc5e66bcffc75eee7edff3621e55c0aac13bdd0c71
zba0c1da9a5d5d623df026fff1780ba0ef0395bacf6326dcab349def2473ff16bf639ed6dfb5a64
z07ca5490bcebd67f10cbebaefbd918714b05886e8a022005004fb7173e22655d740c95411b05a9
zdaebc0d400dbe4153f4a64ef574364cb4345a163bafd2b9a1d1193dc3a8f1ee0e3d865c7e7b0bc
z4fc4c7b69e299b02958ae7e2e08ef97a34db3b688ee0151b5820f7e19357d8b22527c56c67951b
z2fefb95684ce7f6654f54f4680cb1e53975b6e7b1f99201926a600f4a9468d9a7dd44620d53a4d
z8fe1406dd7b80d6db39159d9e558f6dae26785ee9b5c05921adb64a42de6327838dd53af67298f
zf5f6917c7b833e7c6c264f4f39069f66ea2c9c92105ba0226dc53a416fa0b42ac824bcaa4eaa07
z95695e385203fc4dd14faca67a2b6e04f86bf685ad1a0136e1ad445da8f316b3de8e81b9b3ec68
z026506c21635ec84c62d4780101f55f4a8aa9601c655208d97433d00e20570e2e39d0724a15112
z35d2399d537e6f3ad192783cb23ae241a4dbe2ed8f07df9a682c4200abbd902bd00a2ecafd21a3
z933e509b6d781ea0a74a0fdf5c5bd2472e43aae5d74a1c8a4a79eaf87f876838ff7022763f3dd7
zae67ac537815e17bc525131b7faf4c43a6348a7cb38d9638d520ccc2cbca8177db000dfee5e4bd
z1f733960b7ed3f9bddb1c7c35adaf5565104f74050ff571502139e605e84dfd06e2636ef8e0af3
z6e674c5b9fdd0e1b9c45a1cc4dd0580ffbffe05c86e6f47f07130e9f6e26da6691642a03678634
z3c1a744ebeb7b748fb1bcf5b9bced6dfee264e1cdba77c5699f7432355adf8cb10734222369b07
z459e7b80d0789c7c8a503baa0c2533a4892cee03c86475f2c31534293a1d511c0479f2d5041ee3
ze57bb817c9aa7bcafb82370f9d658f6f3631ab949caef7f8e0cbb5944ffc8285d5115be0a5b5db
z4eb3a3e4ba28cbeed9515957d6d0cbaaec32edaa87817e36ba7b8eeded8750185bc2f790abfd6d
za583f44e387cc6f23ba83ba77768f32bf8e70897a19be336eee5ef4113925b1655b4b0be6491c4
z273b9d3e3e080b5028c9a844513db3b3370490b58f6a16f1ea003470f1be3d8f90ba347329fbae
z8b901ce7bed0158ef8e4d51e180e3bb17e9945ef67b7f44db75de6fca8cab4153f20b6759409aa
z3c0033a7dd1e7bf33efc8fc990850a45d86d15fc2f81821c016aea20d8ea2828a1f759bab2fcc2
z57148154bb46a505c687318645266396c5010d3ef286201b0715bbf8b142ecfe419115ee9ddb93
z27db702c3ffd252b88471d58a4101c30a4bd3360e45aa7d7f4e8504f9ff37be6974824c7f667cc
za36da8280f5dfe393ac5ebccdf08de94066770d939df8a7d587349368f680f14029f87f58cbf4c
z295ad92a447622a5682050cdcc61ac332047561611c1c471e3f4c8d289b667ccbd5be1a6624aec
zb684446b4907a397a1a6fff42e35359634310d7fb099da3c51f1c09f4d2f43364636ea884d8b6a
zed5972151b5553204b5733c0c8b93d2dc74ce2f5cfe6b206d5a9edfe2bb1a711ed688a57c77dac
z37600c29c79eaef4da39ab7e895e1c731921369f414cf91027ed110c20f5492fa73fd448ddac64
z8a0a82c2af4a0529e130a3ca43406391c3b15cd66bc142bc4741f4ce48d75eb6eb3adee787e9d1
ze979767137b4a78b27f90abe24b5b6fd3860593f0b46b70727d3994ede52afcf4bedf1dbb717d9
z8a59d61944201a7c2b27b3a0bcc5976745913ad78922af0ccba147f77deb520b9bfc55226b333d
zbd34cdcddc4b678ee4a808d33b764cc04d8b106840d3b99572bebb0a4f65aebff149ea0e06aeb0
z6e27d250c11ab3445241d7fc49dd798f4bdd486901d318e9dac7277c2a026b04b0dbc607cb4ed8
zd53a19fcae11fdb622cab90b814d742cf140229bc5ded509b88d505925ede13d17205a489e825a
z97d3e4146587e607ddb8747473a0fae1962849cd7a5422e38df891fd040f91fd1d4fdc3e268625
zbbf2f30d02799aae6027a34dc5bfeae88fb5308f764e201ae97b8ed233eb88bb5b66dbcb8d8e79
zd08324033831c6752f3fe70b52a65ebfd88ed70336dd6c5076828c483e9bf2bbf7feda2a6eb2b5
z49a13e00d30a3ab63ef947ad8a17b19a7e0028394a0d13e519f0bb66ea1727a92160c688fd6341
zfbd831a020c5dcfcb443c3758f2ca9d662765e22bb7c394e520642bfe980bece99d6530fb8f191
z193fd1cd4a7f85ac94138a0dacf0740bff2fdeee25203c4920ad07551ebac15c53a9df71141169
z091ae529cbc4b4c00618752b9bc25332800086262518d6741800f9ce0cd80262ebfd494e680138
z601dfa1d05715b08e8f30db19655bf22817c7b36a3e964997c7a5395903caf931f562f0a695b74
z6be5a72c51eeebc10d9c55a60f3edd1e8743386e351b88e24daa430573eb8c3d05e1598e5f10db
z477b808c74fa363a7f383cdda193b21b743d67c9f5a8f635c19a71e1725dbed08f2c0b0718bf47
zd86bf4977b34d9969334bd6da16b1f6ef7c75c888e5e0477c7db354d4ca5d480d0473a2bc230f0
z3d325dc7dd89b3226e4ed96be8fd64ad8cf1af376b874f5a020145d55659c9846faabd7bd97de2
z59284a5760c915f90a62896f38a0857bc0f83a65f28f95f91b32035e4c35145472f85b74071ff5
zff93014b81e94c6b980173d50002c88e52bad7da5a7a766338d06b9d8c36bb97d67dfc391573af
za94ee04fcd70b9562de36293fb8d561aed272c9dd81d0e46bd3f95fdcbd31a5f5c991d893d6ee6
zeaa84bd8959f16c25651d09024599a5e5738cc2b5fca61dcaa987b5ce141a5a241b89df9f4dd2e
zac2430e4a900f894d397cab0d75aa6477135659c534a8e7b8adb30ed770686b3ec2502045d6286
zcca80454100ad98714f72f64a76198bf3c93256e48017aaf39747044f146f4da49c0005f923acc
z446b5174a33bf5850235150be891434c83d7947dd317674e9941615a1013001e109f0684b9bdf6
z68abe70d643b43a3127191b77efc874e096967a2902c8ba51f2819f220c0c218b31b68210da5df
zeed0d5dd879e2e3420e2802ebac03b58386e4943ab346a7158b0876e4491a7aa48f54d45826eb0
zf28e47f60360f8708770f479fa45f864aabf021b8d7b76b22e5b710c4233f06310e4456b5ad76e
zc2298bbb127f865947ed2ce01755e032f90413b5407d3678a2b1b6f6d4bc43752e0ea6824145f9
zfaac73112d2d0f927531399707dffa4fdb59ba601e50386205ba5b8bdd6925934fda154694d0bf
zfbf6704b9c5e9cdccc4e3551ec3ab3880de9f34ee355cf80ef9aa2f896140450a4ecee8111bd52
z1340fdf2361aa9c21337f6cdb48b3b8adaa000109265b57de3d233ad2c03136afaa1c78dc97a43
zcc2650e40fad765c30ac3c2935d3fc9216b9fbef83d9d7fb95b2552af257d0698d3df34ccea206
zce37bea0276aaac455fd8667ffba79a7881919186cac7fc25da9ae058a9bbde77a3b800768e3b0
z332cdaa9853a2ce8a2883d77ac8377edf59a7cd453459aa11d8cb8f1476651c352dc963a2c0475
z8160b5e99053b1afbff811802d9ab9fbd314eea3e4876ca62b628fb9665a581008d8eb14a26879
zdf20a621996c7e9e4e63d503eb5803603db1a98910d18bdcc6d308c45c8c2305a59486ebf8ce7a
z41327217b1462265ae3f7dd58737e901a4eb59cc890acb07f4de96a6edbe879a509ed01efd4775
z8290fe547baa3f0231c73e23fbbd2bfdaf86bdaed5c029eb7f04e0b6a2e82ddf2e4f9c17d0f2c5
z67d8bc261e442d425620a0ee5c1749cba2efc7885f1ca2a66d43da61e7af0fc597b09a5b9839f3
z64e8b3eaa78423134fe2468ec8e3ff3e45734f1c0cfadf9c6eef6d9974c309db07d5d05448b297
zcb1070fb0c153eb15957953314be75c590f88808c5e71125a6510b3b129ab091102be7d62e0a7a
zf4f8a52ae6eec666bb9a86cb54c27685dd901c82e6deb6f39260b1873a24fccf465b5056355929
z81982e49068c1120c3498a2c8fbe51652e573cb9c7917ab2caff7e1950db56ef64d2d7bf5a0350
zd1b5eec3e1c8f16672d9b7d71131dca7ae1a8dc2667847f03f7fbdb9845d2a4b646610264575e6
z3497960e7db9fdde2b8b112a9a1297ad1c74f9b27635be30905095e835c461d105fce2447bed51
zba5d26a18fa5d2de2d72a6f0ce5ed7a9331ac2f260ec07971b8f92b96285567c8c60ef4e172bcc
z2ecd1774c04183b8e116d36217f9478143b377b7455ddc12cc26a77ba68ad63910cae262600d34
z0467db7950c4a951d910b52e56d0e7cacbab586ec942adbbb8b9bf88bde74b4a868d9ee1ee3483
zd6eb88fa65f9f2a8184510d8d7d8a7c7284a8ae31674e1751107afbd67df3b291377b3ecd515d2
z6293973ad2a7161d2b3c03f04627b3197c5ff4dbaa0f6aca4d6f2fd3cb93658205c2a1884b2b5f
z04be2d250318423c4f59c166100d3b81d37a925de01992dd76cc0fd527601987984dafb9a21d71
zb33f53c44f620c02e54f3c91cb767bdd84f5f7a6ac1fa5427e9ec40373f90ee3f139b130eab930
zd18df6d0f6448450caa6352aa5fbee2d2a4b2ad53f7e5e41444e1348c1bd5490d0aa1bde93aea6
z47fad5dd7bff2f2c0fcf6fc4822bfebfa3ccf826b18d275618fc62587679491da5ced2f7c04f73
zd5943dd5f4a19079458ea3c8b1f2b2eb44b694f0b5f739cf442661254baa7a6ea01111ab5d4483
z9de8e22110e64cd85cb4c9a45f39ce4b8e39b6e6a02132c1676ceed778446fa5e78bcf2511229c
z6c12d0c1d9aa1b3b5bee1fc823646020aa7bf20b857d24b555d680015235ced4bd59a2df8460c8
za5ab0f21c070ff06bcd92f02b5c354c6030ad40d975e88be809577639ef62fd3fdf4f7e748d13c
zda94fc104511676601436802c710562b3559601999c03e1a9b40a29ff248a5c7acd5d937e8f16b
z7564d4c6c56aad620174ee89d07e5005a195f34bbb3b0dc1bd0f62ea3174bb0ce144c7b41ccf64
z7470c2946da204868a9c41072e4fb2961b936cb7edeb2e9a7cbfc48df49fc91446f3cfafe16e5d
za7255e0a3569d60516d2510f134bdf579da54f9a19f74e0074283a113801fea19b4e75db53872b
zd4eb1fb53e3ff402572b3f21e59d0f43636dcfc74ef3f01202f3064bde0a712e68222d514bc223
za7619779901f952a6f5217a2111adc895baa30f861773ad0f5a3244bf345ffbe584133bd2c69e1
zb6108d80a23bf18436980f81854d04d33da5193e37c285a998d567af872f83abd4fcaedff38ef9
z5f61d71ade2499fbb9d90eef04a8efdf0e9338898b3f6ea6c36308ea8ab99006de92fb432e9bcb
zbf4b8fb0ad8a772e654723d31c7ddebb5fbd9c6775ed82816c872147585713dafa05b8f33b499d
z2f6d9d13a057d58da8e3afd6428abd5d98c366369cf20e0d67154e00d07248a1bd43c67f2dcf26
zd0c4ecdfe945031429ec139f15460a9a9161db54e83941bd9a76da412c12db9d4e9afe6197ab94
z8e2c295a421a7622f15e6aa4b3d4c97284d551bdcc5dc537cfe506185e6d2ce8b910d8fb919fc1
za50a75785d74ac8b2a203d80b87c871e824f82b5c814fb67c10993012a367623d33a56cd8481b9
z1f2d6b19ab9da057fbd92e560c201fb60d0407507be72493103c41d98ece5dff0bf39a99aa0c88
z7e7181e4293e1fab1a5ec85059b2352dc26100dc05642579448cf9d35beeff5e51dc6ac6a646fd
z7c87b2bbfcc0472c163e71a9ffca6bc1a6f79c84521b2d70af6944168d310672d8f3ef80d80baf
z9d35a95f59e5b014afd6708d6a4e5ae5b876a4667eabdc698888066c1e7d641bb4168bfb78a7b6
z2ecda28e2505726182697e59a7f7858a34b69df9e7374cf3373808f58240879fdaa96166857e79
z3dd118b1741536d5ed5b24542eb8524d0950f89ca370d05459b62eaff95e97c28befa78ae022a0
z469b14edf5159351e023cf49e9dd15a059e3e97339986d3396e42c2671cec84340c0aa2fc0e575
zd051104b7f5b6d1f8fbb22630c3c561cf2f6a1348cf438cb760f0b6473b1629d0371bfcbe3c1af
zcb82fd21d9447e8b35cc48172d4e4aa749846ec02e34dd93d20089ddd1336815b65a204bd970b7
z16c9598c27656dd9616ac52af031f5579f7094d93b5b2d9678d7f9a6c6ec3e31d35d48b765f27e
z3be9aa2e0e3cca22e617b174a12b9eb67dc8056f9914d1f4b89a6b7bb23fe768811c51e6c46aa1
zd54fdba2c17f12058b8dbff4fae2314a23f93d4cdce0c1fdb919c32e12683f73733c1500d8744b
zf296f0fbfc7cd832c5070aee3f85e1d09aab2091fb7bcb22bd8a9d9fb4a8fb01d87f0b936b769b
z1ab1e69dc2bbfeadbc52046253a9a1b036a9a67523e63d4896824e71914d05a741413844254409
z10747a0cf1b0a05b0da8132fdb2861d4bda988a40cd3472dde7ff61295274ed37ad32639ecbe29
z6ba713e3c2795427883157cc074d9b35eea9f99cdb95921ab7ec79fbc9599033a8cd152add2fe2
z3099556a3ea43912e51b367c377d59f6d91e221a19858b925ed0a5e39e95177815dc640f31e332
ze2e53014379bf93384342a9a58bc56cd016e5732f1cb3cee50b75d441c3c03469da06d969087d3
zdf6eb6d9f8aa046da3780959e2df11958135015352b95bc4b67095e140fb9aa33b12c7921f5e28
z5d93ec6eb4eeb390daff921a5f3d1660deaa5e5e0ac5204e04394ecc2629e935a51bf9fcbc8580
z730431a8586fed58731ab7fcf29bb96f3671ee645394c7cddc8ec2248dfc02d86d475c8b97f0c3
zd3feb1f1c333c3385670598fa85578bb3464ec04c153ff58451315e83688306555bec09022dae8
z56b71854e5dca0a93b399e11bddda8bf88e86597ff26fb048a60cdf76bffa25766d9caa8c4aaef
z6b401ce542b76b176cfb9532d18ec61cac5bd43eebc792a5df97792ba59a0fe9230bf830eac63b
z0ae9b54b66420bf231af3a6c6e8faab41c7b2e8717bc8ea2dd0609254a9f50b1da3e3b10b6c694
z06bb5edcd858df4e26d40374f88fc2eba97b7dfbed2fec274bdfa8c668a03fe9633743ed4f069f
z3ba11f0a0341314b802ef314807f27b1d793dfa0bc171689cd5efc5c51cf8df895b538dd070650
z5bca21bc2f13dcb68697eea128a8e2db6401081ae6a9adfcf3af1844dd7ae800a7ac654a82fc06
zf325ccc964837fb0e01a01c6b3212a8129d00c49dfd45feb508b781471e01c0082be69538afea7
z662eafb92a2686beb0816fc1a19bd626d5a9730f43fc1b11184b63cca0c78003f6a287e264ab6a
zc806f820afd9390c9c8c227969bf31b07b7aa1c6b71d4336c9cded895d1b659f29c63b5fa86b15
z7f501b9378f2571785916c04db8bb7ac9ed607beaeca307aac9bf5858efec50947c32b6f8e92a2
z19b2c8f9c0cd79f5d93b88b73886f74df8d65bf5300f00fec08bab9a601118a4db362e28437fc3
z70f6b331e18656bdb10212c17d92610d4cc3bc938e3c3b0583ebfbf3674df1c1eaed82a043e6d4
z663a74247635dfaceaa9da73708fedc67699c52b364e0dc3277d93041e892b9f22e57bad235010
z5cc8e669d62dd71e2a2d80a3c3fca7b7c5914a1fa53a57e3fa2850a4d7c4303f15780d325121fd
z3caff67f32cc1de80f1349d561da8e547d4d4765fa6397fcbdd3b243581bce7c016050a9c8368f
z6d8b40d288434f58d6c06ee708ece7b48c46c9049ac30d34484cdb7e95ac646fdfba8df2b60468
z3974e84a40c9e1d200a818d64319638a84e0914d1c5ec451afe308ef1082319d55ac329edb2953
zcccb8741bd8d1ca3b77459ad7a4ad14c626544afe676f0e2963e0d1c68bcdc55cfb6dcc2d673bf
ze299ff0278cd54fa3e183be4077dab4bd2e3f319b0bb15387010e268bee0ce529d9c5978296608
z899dccb84bd5f7d466aa08a5023f54f77d4a2a6d0d6abbb410a03be5b4c4ac0cf39848bede933d
z9e79335b568e38bfe0bfc7ddc0ddd55e2d3f2decf43cd8d718d9c522c60645065b065529e94ba9
z582ff06ab9d84eba2525c5142af53404418a3103c5aae6b0eb526516ba66faf99604dfd07bea24
z48b050d39bf776d51bf2d716ba568ddf93b354fa5ee37ad1483299291668309e0e18a018f8d7d6
z1b34335d03a1fbe631149dfd3bbcb160509facab73418ae5ae8d5b552e714455d04edd33f55cce
zfe1cc1e5e374ba04e95fb7684235a61bf6763cf4a1a55ba13f9eb426718681c82b32ebf08c741d
ze073c015492ce8fa2887a0200527d52bf86668a36b70091e94b3304f21d263c767c0693b860ede
zc3c55034e1523432790e24467e0db9575678e121ad8d5947dc0e583ae1832142c85c9b768fd12b
z0be3c967d01e9931a9b4604c1330adcb109f695363c0f856addda1a7d15b8e1827b8acdab02633
z8d8aca3e06c68351cb27733b37e04ec6ab5bf101888cc0b84b4fd4b798ac16ffb74826b240c323
zce24dbea5e1a2c4c45b0a20b8cd1ed5823cc7ba9d2ae0f86431402f4820ec268b84896d595ba6c
z5c5d12975b83d3ecb7cf9362b007a43b3f4d2686f2b43f0ad69037fa2f244355915bf7b4a52707
zab4c4dce97184e61659f4b62bc1eb91bc5e6eda352dfb7e0d80eedd6845c9d7fccf94d0ce653f6
z62193b5d5a435bf281883e450668b273ff99b5d225cb435ecb7e1bd610c9205ac0c3d495c7b299
ze09212f69a9c3770068ca88510c8474159fee14da7d9e62a1c0275ea6b558dcb7499a16233c800
zdc9931bde635959b3d30c25c1dafcf00342699415104d6f98068be062d075f94843657d9880372
z4e65308788d06e402c9ce07b4fa25f6a9a6a45d9774d3a61201c53ea3a6e146f466112511a8cef
ze6c041739b9764147c2901b49857a3d69cb6cd74e6ed9e36521ae5e3ebf7d68fc025ececfadee8
zf57ec22fd01e0461761fc17139df7924b1336aab38715f382d84136d2f161541f9d33a88c93099
z372c09fad42c46b76a99348fc2972d6ce5233973c649f6c00a4ac138d1ec8e1cfc0fbfdb98da1d
z7cba3fdb20f2e8abe6b24a0ff4bf2fee4a6fec08f515ddd3d83d2d61af2d873f4cb10a73eaea1d
za868744a7bf1bca0774249d7dd997f8088d96b7446a901c82ea3e142f385c79bb014e9e1d55419
z2e863277aeda98b36476cfad462826ec5e7a08a8e90fecdd8dc32f4dfcb93c172c460a2cf1bc16
z8080cf3977c82a110656319bb93a72804f68d6e15c24557c62ed7cf6c79a8486dc99eec2b2f6a8
zb10566f35d3ec05b0d755b65f697628aa81537ff3da72ad7e79ee29ed686da79eb27ef23052965
z1d461e732e9f96e1c87d2651de96b31bd675bd586bcf3c62f5ec52d0ebaea1065639b3a9a46055
z6fb0ccc5ee312506cc882576aef0af5f33b08d62198a9ea2991270a4f66cc996d4c843b0aebad6
z9a8442b7000654ebe4b67e8cf5a577a369df4de988eeec50ad269f076897fe38d0b70bc127dd60
zd88ecb0a2170cc8c3648082695e763e20280b7349e66c55a73ad26b3712ed349df35d23cab6aaa
z107533b42b5bd620a68f6ee324eb544a5c99b4af3faaa36e3fbe712ac283d197336d524104a83f
z5b9dd33c43adeb4de796ba846c8297c9a55f691f64ce8a45fbb99958ceb27b3762af6228486919
zdf8d68137f47a6acc6a386023790c96977ed86dd3e57f291b602cc3ec39e5933d773bb7f1a82b8
zc267bfbaf8ca648a119047f5a4a8028bf0b669c8472ce960f87464fddaf00a9eb1f40a1321d86e
z2e2678c1cd5b0895b4598cba6792b27ce242de5e6464e3f5845aa9ef5f042ecbcfdffafa0b019e
zc50e91d8045fdd315d3ab4aa1869598ea2dbf70e16e0442d570a088d4a16117491340e22a4116a
ze1caae7c36c01697de41569e9210cc7dfa19d038ba19f2d3fd7a6368d617e68799c38ac94faa62
ze3ef98d814842d6b851eaac346b012641f388440005d962ddaa30f9724a90f57cf96ecb2985deb
z675fd4eecec7e6abcfc011cc5d84a549897a815a3878f3497a0c9d628884f203fc82f2bd2f3be4
zd17a9914c0895ec01305a284a54a87bfa17fe72b3a6e2998b54acb366ab185b8d48726e7ab3edf
z125103492a9677327d34eff6857372ffe6a63c5fbb6adbd71a9a4b811c4e86e820c22ad65773e3
z9a7793abf4eefb2070173ce99c922d787ac226ec9aee7946f9c0adec636025c876d6731f3f0022
z83c5fc77e7e1dd54da145b456746117b19b84e7596738a49fc0d18d37e20be7ddc538a17590256
z823331d94400d713144f504eaf9185afd4d963039dc614130b1afec61e0e936d1645b64433a493
zddb8aeab34a0db4c39f02a5687d2961a323e963f305275c7b90ca24dbe49e179ae5a202b9efe65
z83e6dc0ed3c0b952495e2583522ca9588a48819f7ec52588c9750bfa85bad885ca70f211f03a5f
za6a388f631b397aa28099e2b780d3c204d3ddadb38805036c878e96e3087e7c2a4e5948b2acd9a
z43eca437d8206b5e6a7eb67f38bd21274caa3d4a849c8d6ffa6187e866c2572eb9ae4effe978ee
z397ede280a0ad73889e2d605061f7e0cbf9a3db238176f13d6648c396fb7ed601e25c3ffcaec87
z2d30207f4af709787f406a1084672ba6d1d62771bb2c6720276c6393d205a9f76d234525c72f40
z77bcd5a8789ca659de06063a03258d66763b118cf58ad4d5a2fc485997271de51788f78fa9b4b4
zfb285b5123154bd70c4dbea556282348e02f06c7cb7540791b896d46c9963a1526ec0c45351d33
z3b9f88c85aa5e13fe2d62170c5d7571e4de48a4866d1e76de59c52bb82554c7a9e0ccb8fd4f152
z700ff5999ba727e07b2b9663b803d08c98b9a84fbee7d490a9553aa087bf24d44a1d93ad71c034
z85bceac627f453ac99fecf6b78d014224f5610891debebd298a7242c1326e038ea3f69a2bd095f
ze4c60234ee8a9dc856ab1aa604cd775e93e52a7a1afb4648036031a181ddfe524c3b545e354170
z00a5e832783412a1742d5497f38aa9f9b566dcb15b6af3fb6d408c57360eada02654e135b19789
z50eac7c2e9b9d33456bb87cc6d55a8980a34e04513a28de97e220bfb78fa05667906ef730ce420
z7bebd839656fbed17694ddfd6b216c8b27cdb1a02d7da8958d26f19a1d6a8dd382a2377840e09f
z268520bfbac60c25b872a8829c94ca7d85f99b7ee123077a6142f450b5f9244149c6303f511cbc
z3963bed181c418514a11d98b3ecb0e179e4a5b5f7706800c17a04452252e00bf1f40fe2b9b10bc
zd142bc5970880fb43b32305472cf7a50bd8853e4a5d5010aa2a06d9bc87a161111509cd47be4da
z2e30bd3542f873a1c454daef46a5fa56ba2701581ebbd27ba0b5644123e33c486042876bff06d1
zf3f8dcd927330130c754e3f593227624bca6625a5e568f911fcc4ca7a1efd03dc929a02257c04d
zf187ffe941c58d0d37427b8334f8ecd1a639429ca64f31a8ffe89afdac7f62ee7ec505f8699738
z795a2561ff28ed8e9ae9bb9e72954af26461777077681069c7cedcbf8089504dbf8c359941656e
z11c9a7d7da2c4f70107e3e339d7dbe63a67155581598b4a92e057297808ef1e3653a3fd0cb0d7a
z59bceaf30e91f904fbec81768b4cb54a8dfe1091cf9dbdffe11efc790a2dae16c71812f8c1b8c2
z7ee6959dec52cff060fc25c3aa923a9432732885046d64e49bfc26638952901e01a2c5c8038203
za613b2e4b79deffc4630faa31a9795fa07d54e83a0557d7515bbf8f5fb17d779aac5708e538891
zcdc02e0a9aba063857eae2de96c8731bb6a24fb904689fa42e5cf4f658bd974176d29ab31dedee
z94ee3630a7168c2625c2f5ce79b9ff2df9f9c8cba8d23131f7677139b95f67eb75f6147a821dcc
z03303ba175cc039b282d4eda934d851749df0129002832b590b69eb29f6d0c55394096b8d4543d
z25b8767e9520f0256b175dd19ded81030be8ac40a9edc66001ffde75b1f203b2742e13b845f57b
z8b06f96c54e9c12be210c0da8672640bd84be1248e2420c3c20658dc99d1271213e5db28309d5a
z5b7b28acc7fde2b7a2b39457480e8d97035d18936ef073198075363033fb6b9296aef3acba1ce9
zdcba273c9354b610c27d07af70893239a5f053d5b237aaad56a3a4002d92a92c02ebfc665b3484
zed8f306025c5654ecc9c0518b1131f063936ead719ef1e60a6e39d5085f3eae58241aadada5417
z1ba17507d1fbda3f75b4414de46c411aac405c9d402289fdb830997abd4b4ba5b40b0738bb0f96
zae9f7c4df764181b5d847462ed6ba8408e9dc84347202aa0e9c05f2a11ba98e187d67cb697b580
za59336c8d5df840f1d269d10450dfff4bd5b0dbadbc70d07e819f5c93d3eba7f1e5332c7cdd9ad
z67c47e773bbd02279acaf78588c4da1d0b034813008d90c3d243d75210af175a3c58d4beee9314
z6d7aace5f158078bb4d151159f36b55e9503128453419862a01285d1cf3e0a8c9f7b06b417497d
z3fb5e31012ddbe7f70f57640764d00d99dc455519b03cc275fbd91d526d989ec543dc8075f0197
z312a578ac1d43b149e24264402bf63acb6ff044b2c1bf790f9d185866de15364b2a7fa52a9c12b
za2695ef02adc6f8973d81771e39d536ba0c0831604e90f9e37ddcc043e72f106d7975043474712
z0eca707865946f21fa482f46b168229d7b1fbb83cb009c68fca0ee31d8fee2a7b7a1ffab5fcb96
za02e157a13084629abf55eca938317204df01e62c853d7f4edc2a1a97f2be976200f57beb9198a
zc97bb817a9c7240fddff0e5e624820bee3949b7fec40e5c17bbff90f9b1d1df6e3212419bb730e
z799f01354f3f6491adee238438f3af61a225d0489204e65a03565ea4e226a20cf7b43659e07cd6
za9155578cc88cf2b7aac1a1e6c11620ab33956d1af7cae8b2abad80b6892dc7fadb043f71acd2a
z53d2e3f0412b661f1ef76cf4e3918cf7c7b35bd999cfbae8b61cbee6d40a9839c8033920c6d0db
zb32e0c554ad7f956a486d3ab210de39ef99ea84b121b8382485e6fd39f018286d5eb767f4ce9ef
z8ffbbc7f325f1f3104e1234948f777be0ff3b029bc2ecaa9f54517d72f4555dcd6795582c84c29
z4595b7444ccce108bafde7018ae97b3925ed3f9c754d292e755eeea10f228067252621f351cbfc
z21fa8b3ad8424dd229c42da5434a9a19b5505a8719c26517c2cdbafc3b56adf5790ce08e465217
ze8f279e3d22f2b7ef6ed529efbe42010c256371ad4c027b608adda8fe2e04de36941107c9b1611
z153631fd813c14aff3bead7cafb30df1e57b52544345f416755f36a4854bc4ea5b5c24ae88c63b
zddcd6a50026d59d1347397d053e6728bf478435424cf7141e11e05f11b196520688b86e56a48cf
z09758381275503c5b6afd02205152ccbc1dccba62ff7a68d49ecc715b9e50a25a8de8a403e0c08
z8adad0d7faa96b632685d35ddee52a755b565f12fe75a369ec1e83684c79063376eb3849873038
z3515919e8016e646f4b691b90808f2f81ab2409e417649fd3402c3e788fea49e68f68134eed585
ze2d5a9b5d18673490ffb5d55f0e833abe1db4572d578cc929b4946e02f119b8016c8fb823e3cdc
z5db6ee6774ffed9754ec91057b3be800af60f3e4a2d1df8693deba930cd59ab8d7c10d36391f6e
zc8398eb40b53e8803b8d0b207e50347f0917be5dcfb6da17b5bc8853ed9636e81bc99702ad3dbe
z5a65b4a8600cd84bd905646c02dc57b72ec20fcd45b021e05fc37d27c98d2e0333ed30f57a31ed
ze8f82f88deec10dbce5788d440f47e22464cc91b6750a1076174b7c0125bcf15a2b2726b902085
z4235148ceca1a259b8cad1b3163b2f82a2a25140a3e93e4e70cc2723b0c1c26a546f1067d110bc
zc9c9b59eb027995ea23fc220edfde2aeb21a935583b17f162ac758485573b4cae29ecac5e1943c
z30914ce0368fa2eff4f01c0e6eeb7f599aa6557d266e2bb11c7774b88b51be3dec292ca8cec695
zc13b030603e6101a43a28451713753e115cbb7ae9fa0340c1213f8dc947744d162e655e77b4c24
z84b4231439bd5a97c40b0fb59544b9a362c597c398a5b348f001f6c0103805471d78b9ccdcafbf
zc21f1ed9ba25ea161734a1b2479d298759f311a528e4adbb06e254e5d03207a536d8c494e032bf
zd7ee480707f66c6361040b77f923f4daee4b699c12d01c1a6f6e69aa6c514cc4a66d6e05e4cb3d
z9f910686507f8f2f4ce1e6126b281e1a0280f20465aca82e61b12d09d8d7ee1a6525c13d1f71cb
z6a715c2592baa2e09b35883a4945a14dd8db60c26d43fdc417e3ed3fd6154fa268647b3ae8c85b
zbc128041dd7d09ef4058e9d6d3b62d251b9e8ef13b0cbf14ce656196f4b178499c5b87dc4a2f56
z79225681b90c954fb6b9a7ad5f70f9bbc8bcec3be0b11810692071eadd1102f1790e096f9a01b7
z723fad8552e6cd8d8b89cc0502693f6e6fa6a7f6052c45709b2af21c73523da537c04ce3d8fcfe
z639eb9d03889ca5aa18043e338713d93f1aa89b882eec6105be838fa369f206f42e7bc7f4cbcd9
zf9ff8205ec063e30cff2d9a118e8cd8b4f886ab90ec0984eaa91356b6feb6bb4f0cf135d30957a
z2ce571e26431be293ebf2a12bdd1628ce0a8f317bd11b45272747f2d61f98fa654af8aa5502aba
zdc57ca973e0c4af61c20900ad7bd085ea6846be6f110c4faa7f0a02586d39eeeff306df2684535
za3f822457b6e3870b5f22b030a9ecb6055c2d46c46c0fdaa1085f253a2f7908e42a8000f749f48
z9e0e95c6c04d7b02d838da4ff0522d903cfccfe58c1d3cb8c016dc7a63ba5cdc2cc3fb00167952
zacb59d13c8ad7f1f969583624811735a3f83f3a3fe1dcc39f09f1f30fa8f199c6c1779b8d8ae0c
z1087b19e42140c4f9f9f07fd9dfe3e88ae6b101d69bba89cb84fe6bcdbe1c5f671a5ebfc4f0fb9
zff007ff80c1bf461cfbad7002f08095fdf23b01c8978f63963a5366ee0dc6700a757d067cc41fe
z87c15af922f7597a4fde713ec59a927a3ea938785b31e2145c73bca291d7d56216103d5504c7f8
zd0a386c6419e24a3a1b9578ee37f291ccca436f94449f37c51bb18e60d860d4e830e3916a97bf6
zbcec490daa731801eac859ed7aa7f33dcab7cea0c69e44dd45235d201e71c60440475e2453f1b3
z470fd00af46382591719e4ed1984974099eb8bdfab2fa1e807f4e514f79242d4603a8361844188
z9ef4b0f0dcc611ad6b1c6adc2a87aecec2d6d064b29daacc1fa15aeefc1e1026b33dddcb5c7e3e
z18b8f1158d5012d15fc8fbf6738ca4682d17a020dcf4a3536f36466718d0af7082eef0bb34a408
z196a744c9b187983cf056af7851fb6ae5c381847166189a99fa574a4afa3866d4f2257b8d1ed24
z56b1ee28548a9d5ae4bfb64e536a10ba85eac0f82b1ded7035c65a48a07b34f51e2047ba6c9f0a
zae2748f8ca7a077961a013c0aa563832a0c201fec2c72728a6fffea67cf5c6f3209e1c30cff37f
zf3134a26dc4e7301a88c3fd61199cf5c29057a284a8d70981f7e779d413480dd9231ab3c1bf9e2
zf8014ec2612a5ab688ad4b884700615821eb38917da5d9aca0e9dbfc2a4a5b12cb2199269deec3
z82cc7cd6c31139777fc01bd3608479159d360801976ea583638b9659a2eb08b7e22c766cfc89f1
z82481bf4cde88164df0974db7dbd5f469411295dd499749c64d8e68aa3366caf1d4da8e4560844
z30e6b1244ba0256a5b5ff42d7fbae2a75f3841b5cb45e0c0a1c15d3cc8deb5ba1c7f36008dc81b
zea7e4b6479ca3d0d967192e489d5784f9db965483158a9afd63f3ae3d2262c0b4f913d91815543
z3801ebdc0592593eebf0d795e2b0f03fbeaad9bdc3fad45a5e1e306dfaa679894fd13b07bc062c
z8c0416850bc4601241a9439ab568794a1923c5e92e98726ae5d22447f4fac245df8884d16c4143
z50864466530cd02703b154e31e7729504c3596fc7ed113de89004b1b67a9cbdb3f02ea5b65d702
zc14bdb1259c0ca494d8aca0013549cbe958e47c6d05bd6dcedc3eb4351ff49ae7192de5dd48f1e
zd189e6abd34d6795a69132c8be879828517451504973ade0d9f6e2469612af06b63eba0ee03e9b
z5ee56fce76a81a0b1de58c3e1c1d3d75460732bc440977ed1a1b650e8930cf09128d7958d11bfe
z5eb26aa44598ddb7b254f80aee9e0eb4c0f161f62e79dcf8007ca358705feaced2604423b64999
z9db57c6d414591e59e60c16354f992f10ac023d108e55b7acee29ad90b1ea9c03dcd529af300bd
z1de707edc76de22f5e07eb812ee196301cdf77f552932ad5935a58a9a8ce08fa8bb9633fd4b470
z4f4336e2f399bf52184b6fac658f6ae552d00d02c1e9c4ea6910862517e1867ad8b1c73969f5de
z5b223e21aa550086df3bc14b345f5d375ca055d2a37ae6dcc3f13f656fba85facbfd20640e0eeb
ze8322042f7a85250e02456fd37dfcca85e9ce42eab6960c1f4233c681fed33dac70b3148455989
zed3c6b65e94bac8a7070a4eb48e519994465d9a3abb170923954bd7786a0ef8a2af2e87e58fe3a
zaf5800162d0d81c25d4c425b1130ce86554080ce93ef9954a2d5bb5e8fe15b594c7dda0ec73712
zb1efcf96ae9a7b9a4b2c86c46d3f28e2ca8428ca9d0aa868a51c57e56568a076ded2b868072d3b
z499ff536506dceca047fdfe65bcbeee0a693bd2a1aa72b23e7d3d12d62cbb68247b320b15511df
z3f74be8e6068ce86ebf6af4bc03b9182ac4ebd500bc0b7aa436d8ef08d54a9a826410274b65ba8
zf7eef8932297963e25fda853d7889be8602b25447835191a19920c2a4e776aee07f2be59a7f992
zac2252922b910d4070a55973d5cced0fa73bbfe6035bb06c56ad293e7817cccf0422a83ade921d
z2e0a7f8b58fb080abfa1e87133f56063d74ed3979dce4a83cee3cb464cbe205a9d3e2fbe96fdd5
zca872e0ec41a7dfcec911ff972df6abed69530c365c19983d10064f49416009b7ff746131b176f
zd6620e42102371efcf9f3c6b0044f4a990f28240c88621efb1d2f74093ac1133074ab5a530e1ed
zc964c8ec3630051ec544c4f0644c4ba8edc16a3e4d711ac0173e4269508e2370e205c55d348ea3
z6cd739f56d055a4ad8ec0c25c332915fb40afefa240f7caf42d4e4d228f94a405a1956907a54a2
z37e254639b0fc2353a2ccf586c146e2f1361005e51df19fe0cb4d5ffd307c6a1450ec1e87fef98
z00d2d8f22fabc3d036c0ed890365b3a763ab9d5ddc3380e3229c2d4100a445583ab371d2f9b3a4
zd3dfc9cb138a893280181be7410c2389618f10f71a7b1f42ce0936ee99b0d9ae99cdd73e28ac00
z4f3ef56e13866b7b068d269235c039cac5c04dd8812e4663c9886db0ff468e800c19a8067a288a
z3e93ac505f956076afd96f945f67ae2c99bcb0b46eb691a79cf6b0de4d46833b872b6b9973731d
z3ca34e6f7e7a211e3ed565245a8071648c6d80a6139212396e7fb714190aad39206a6829f2bb7d
z8af6d0875d1def035a56d6924277d0dce71a0af9377bb944b1ac80bbf1ac50d5da16001c0bc180
z58ccda1f7a1d12127699b9e17abc0d1335dba1d2be56c9e91a631af9ea81bb1159e9ab37c678af
z198b6f6e6e281a409cb4a26e78b399c579222bdc33523e30b8dce6e66693dfed194d14eec61df1
z61329d4e6ad009bee808a5a8e16abb29225f17057e212ba4bb1be471d8b02ef7668eadcb2d4fab
z6380c6715e77adf09a0a3ad6f8a2e992d1da55b06d66fa009ff7c051b408309d6acee74c6dee46
z3844229db2753ef73116d1a8227ce4eb6c4c742b36da0636803044dcf664b3f72213b8ad5b083f
za94f49dc9080034bbdc4c1134e96907e73dcf53ac67ee9fdc08b3229973355f07345dddae97675
z53b1cf753568ec61a32dc3a99addc8ca7d38f103877bc847a69cbc612f55c610a04d877e032fbb
z07bb3871e126aab37d54635362db9974008c27b1e90bb3f212e87ed3a7b3c65462616961f144a0
z819e44070db7a849d8cd90ee2842d7d9c6cce51140eb8fc8af16340d6299f2ce82135476443af1
z40b0b3f733bedd3ad1fd3d6e4f756b76e1262ebba12eaddba052f8c45779db2c341bbfadb89403
z047416b268c510a1aa33c8811329e87bfd0cf94a865c0f186dff11297bee46e062bdd21f9125db
z3c3ed3af4a03968db8a303c27b00da017f2c181d05067071128abfe3278244f2a754db08fde811
z4a01599c3303aa384703bb863aba31a5ffb79987da8b8d252480fa8d21e3e431442cdea2db6ace
z608721b938a0ec05e85cb08c08c4b0dcc0b3cf1652e3356bc34db91003f2d6aa8802e3b32889d6
z3974025bb5c6f329e1a492098a6561932cadbd041de4e6e57628ba0a80f7bc3024d4c1d04b7b74
ze4f41a88898d06199878eced017fe06149f9784159c128e405ef152bd6ba0cde5fc6f911276f98
ze69c9e1437bea9c07de34bac35e05612d92f8cc4a445cda4cd0c4780d3d1f2cf199818538e0337
z5c3499c0c74a0b2e2a5889e2d6f542822287ae5e2d4d454960a904778d0eccd6f565fbe63fb8df
z2b4a79b9c3c04deaa5a152af97e6716dc56d727ce60cd3adc7384a2a719510276935386d62b4d6
zc6152a5a99fd2a4a8143afd98b91da1ba609798425ce9989573c8fc7a167ac2cb85b30953b7f83
zca9d71b6ff693dc23218bd019b1a27dfc7f4fa7557f6e0582230bdb070cc757d7a7cb3e9eaf394
z1917fabc0cda3cc4e861ffafc3896cac23ab4213230ad6e8283e88d48d9950cef90c972a769f50
zb2cc6c6c67227f32acd35247032cab809790538ba1b48910622f7c57bbffee81204c96239ef1f1
z5fa1732116530356d9d4f45633f83c97171909108c4b25957ab935b809379d07d3e2b14c3f2ca3
z5662991fddc9a7e94a44327844bb2ccfcebb6ff6754675bf2ce16f628da806f7161378939836da
z67814495f6293de1ab53ce7ee377aa4b7d634caea20cb0cb0ce873314ef6e861cc7d3269e40d41
z9658af393d91dc1c108ae99c7792753c1936b4fca79b00f799cc1c432d49832089d3800fb86d3b
zd93c974b661a30753c775b022b5113f4bbbee158319c1b0d5175dafd7fe49fbafc9c4aa24a2115
ze0f70f9f6058ea6d7855b9442a9c9d0b4c0a9a96b45ac5acdb40411df76f70377a27008ef74b12
ze2f89f6322e18e3ebb316aa43505b76ac3ab09fb8b5f6c013fbde4f36254704aaa3fb012156428
ze6ceb3f811523a7b710eeb48f327f7dc4fca676eaebc881c6f1b34dac8f3c932184182062753c8
zbf7d723885dc7d382826b8502247aabfafdb53789a8ae42362b2ea60eeeef8435b12a50cb4c0cd
za7c96f1d0b79bbef12fbda8cdf1f1664c7ab0ab24f77d10844b4f905d7443734f9912b32f2495b
z985b3a3a9e69de83d4c834396733255b6cb314bbb012db6d46be73cea28aa6bc04e17ecfca63cc
zc2aed669473a3a2489d473e55784a571705badb88d27154ca8d2272eb70722a050402824194b32
z4187e377a2a13985d57232077b69e83398376e08f23f632d2483f3db16562d9c08c4a635a4170d
zfce09dec265ef2c33af0514f6643e4ae254c5e914a7c457487d8ce3e411b452d567be010de3b1e
z71e14b75bf5f56645eff6c4a4b489afaa0883ce76fd3b947b229226f9276a48953d263b5a80647
ze21cb825f40cf4f4291ac2c6a56dc47cb6378f9ee201c2b8c607227629e13108b2dfae0b5e9e6e
zf7fcbe21a525b254cd7fb26f637e2b4a17fa31f75bad234ef2f164e5df86d31545ffabf676b6e1
zf42fdb135e75940af54eef6e819a6b5b7c0323594b715f3a235241faa6b3ccc9bdf576401341a5
z1d502a4ec32161eb5a51a852cf669c50d8e186c915726bdaf80f2aec221d6625a949366e9ef17d
zc9a148188898a213812dcd7f452038948a295043cebd69ec476fd33e3dbac2797ef7a3f377baa5
z55447a7804b3526f3befc7c8359a71de7d6ecd164d262dff63f46bd248c3522e0417c55d90361a
zc4c6f1b6517543fcb82cc406fb88220fb996f0dfa1c979fb807941fa2d88b9b689b33f848290f6
z235eb0ba2ded1db12f8f2896f569bcb4247e01bf3b0c02773f7ca375c0445e59ef726f6278c514
z6d82ffe2902bf08cd6d8b18d31e35cdc80be69b563b6466075c9fddbde0f1e8c72c12515e6b9b0
z093a35046ced41fcad0c637b95a930705cb0d000cbe73e4322ecb73539dbc503e7a54e27a0649d
z8a0932ccc3af8ac5eb88c4edcc2cb2fdba5e42cee208ed13aea2d4ddd73d4cff7e9cd9f31b7774
zb67d1ee5b7055d70ca54af8c37c6872b2b000fbd8a2b450958211094633ec6588978b954498b8b
zc5d03b40022a1817137eee851c06333aac946a8e185b755afc2c82c45b87c1d1dc8944e93d41b8
z491c03e6749e0db18b4d6db3d844abac24c26a920940aab22a84f2f7811b549f12278094f40662
z68fa5e4a560331fc142d31e710072d64f4af74d52cf7d7c535ea7a8e0f3ea13dd0b451fd618075
z655c68f1d29765dd5c392b37ad6753d076adb00a045c922a2b31a84c109267c919e7bdb5b869d0
z686e41f6d2dec757a67bf58b2dd0296bd9508902690886aa1f7212b54f127516fa37a299b2240a
z7ba62b8be05864999c22e856bea6835831476ce7acaa29659090ab9f7492ba69ae3bbd77133599
z157fe0aac8ba012a12cc544f7a381caddbdab97dc960764ddf6ddf4feee138f3e80df7ba72ecee
z18d8ef808fd7633084fffe0bd708d53198623e80d9430fd10a54649f197938f81c55805bc46902
za04175b630e073a69a3282d19c7a2a8e1b8470042a5fa5da8c1be69f58b0b996e8a328422eafd9
zc28b028d4a2be81dbc2314435c4649709624ecc596d295612cf2f3a64beb43c8dada26f94a27ad
zcf9cf58fb942fd6dbf4d20fb7d96db8512d7c54734decbca471ff14604ec353ca4c0711edd78f1
z900d195238db30afcf9127c5700bcc6585df96ec2ad6d98cc0cb0a20b4188b9cc2dde6c372cc2c
z8f39be6b871d289dea788f2703ca7c26ed7798e786ee8829e046ad4bd7059e9b6cffad8de01e1f
z1a683f4141517e75ab3e5a7f6f3fa10f56f2209635c99f6498779ed6447c5d3a34540065e38c96
z383c77f2f34216bb21f1fd8f43144a01020b60739fac77b94232efb128603e847c6b5136607391
ze48a4c14f99cff99399371c0d81fc4a060f76e83df63f2cb46b49a19e736baa4e49390952a24de
z778a7e2dc6e7f2197df9ef0dbe6cb9fe75617cbe1daf1dcae8eeadf34c1431e87ee8d17eed87bf
z0427132a3df12d39800f0743af548f92adb4f67c371953d922fb4fe353a91d2f6626e30e83875d
z1b1c2d1f151f3c562a646b7bc9d0aa81c4ba06c6c2445eee035f4d6017da56d7eea3471814be65
z20336ef381ab6e806edcd8fabe02ab6b67ab2223e958d39f2e28dd3b947fbb361bed1f6ca5a359
ze24a177d7db74ec89cef99a63124b800e00602b25ea22d2da85d9b5693665b6ad48eae44e0b5d1
zda55f3cbe0b421cf39ea4a63897148e5cfc6c63a3df00f4a5545c616450ba28ec2a9d6f0ec337a
zeeff9e6d0a907a375f0cc68ab9bb95ada690ce3dd4e4647e16b8bce81aaee6546bdef55d35591e
z5d23ab13caf21fd7c591428f18965b0f744e75ba66b0427da2364cfc4944cf1fcddc1e515c2cee
z8093b2d646028887a4fb77012ba2593fbf05336cadb165ad233adf06fb86ac9e46f4b766e4553a
z9c765ee93fef8ee5653537e7c7fa9ef66995283071b5eac610e34ffd8c998987715ae3bfe0bd24
zfec2934a3770d2fedd7fe26549ad2567d9033eb981dd28bba503da001473d559edb02c7a16c8c5
zd43aeb1f4ef2b6e87008af2552e85c26adcc1ef54127bd6e17bd470ec0b8b7e9587d43e5f0f465
z7d32b3c11a0d87d998b82669043399bc2e387bc3b45caf5784016272c98905f2580615c93ae1e7
z67ee1503158222e00793da91f2a6878bf1b60fabf8862992c075d96f34bf887673bfb51bd53550
z4da865cfe374b49e860d14e2b3095173190da0bb62ae08319d30cb45cddd5b1025535fc4a65da1
zec970132d39cee4814f276b660d7933bb6e38e0da913396525dee70b3814daf8379ac83b109eff
zaa5cb5100a12e2d999ad86901d1acea9cccf32673e36f3a8b58228a69aad02068b87043d3dae29
z59b010dacf1532b914d9b5e5cdf19ccb349ce5e47eff8da927983b27eba0a941ffd953e0c7bd04
zc6cd468972a1ed74768224a19f7ddc90c5664778e8a7ef2148aed4b5a36f0818047f224a6a8c27
z4c4232a4bc9e4bc9d0307353fa86d8a5a491c9ce736b81bc2d6e55ddde639dc70b0153584737fa
z6e91a4e6cb3e13703df89090f5836072fbb3ea80f823e2d5280c01603ea3ac6c3b067f8939ec8b
z2b20e812e0d3583862d2b920cec823c3fc98851e8e11208af98d5d94cd597c6afdddf503e49a63
zf647020da8e3575e7ad51d2bfcc543740dd2422db85a492b9591672edaa990ac720d5b3f203e59
z30555184bacebb9dfa78087231dfb976673ee2f2275098fe1df4343f52c51190914ab7e64058bf
z41f34cbeaab7da8d6643318962152a1be5b0ab761748ff2d67080e5032831d44d77dbc310e1c08
z8cc036d6c989033362e871de3d607c55ddc9d898bd4f2381f93dbbd415970fe05afc514b0981ae
zab78c6360e7e106dde537df59ff17325e0ab5a1c3087f5e3bf5e382c65b3ea7a0200f1e8d49f90
z1a381f80c9adf9d16d92737bfc00a8db4ae6017ec3f544eb43b53c8bcc09a8214df1d82bf70626
z4cecfaa8c38703ddaacc28bc96c2c81ca90e6a8b1e8d5b6431773bdcfc6b82a32a61c1522bd64c
z17de98823936257839b0da6c7382be755e0b83efa92ea646b20413d1fe64a99b711d7be6a63d70
z1e2d913dcfeef8ec6e15081e6523e0ad9761dc1bf25eb07401e2514877929a60022885244b3efd
zf8c5f22846133c5724237b1f8634dde250cf2636f8020b4f1f9a8f97ae997350d8093647330e97
z5ec839be1a2519e65b733c54a692d21de4229d8ae0aac0217c1002af7b07731a1132c9276ce26f
z86fcaddfaa52d203b1589dfaa04fe33a60d13a91bd7cdf2c24c2ddd7142e527d8f5be36d0eaf55
za596dbbfa98b2734e5beb932b636d2f0943f2b1d7fbbcee565e0f563c880be595678c717b62a03
za40381cb8ae8f1bf5cc030db3aa4a40c11d120cbee76d388ebcf8ce3705fbea610506b48e51fd9
z00bb56ef14905cb39eb189310a7be6957cd8af9f3b86dd54f3a9509c9781297c2f7aa20b2e44f5
zdec49c99a0e6cf2dcb841eb171510f5b08a0b3d63127fc79d04f95dd0aa4a47976be0053b8b9de
zaba1ba3cd35bf2d171a3bf1f69a85f9c06a21814c27a8a1b1091f243c9037f77a8b99c3833cc9d
zbcea284a27222169d1a203e4e75131f05e764ab549b11960ffcac27586de8f5a238ec5aae76589
z0d34ebdaab56ecb8f8b5fc8908727d678dbd431fc963453ab75325b1fd2e5eb8f08679ed4a9792
zf6b9d57e769f1034123517de27df9c5fe6bc9f141bae3344074e2edb27498df577ce04fc91bc1f
z162abfcd0247f2a68c6c611c171de7966e24ceb4f3875d3e692af2f72511ecf0253065b780d7a2
z2a12f3f1c64424645ba12a49d93b7f651a4461391a276db7c9cb498e576f319457f4a0bdf46864
z100caa3a0c011ce98090175a14167960f186d456bf861069ea327d416b3fb36679edad1d57bd51
za6ca14ce4f7e9b072b5345549a7d4742d9ecb25aad7759c314a28982e74a6456d2f9910ced7f1f
zd0382c89b29a71c31c9965625dd1a5cd23d0f52f20dbc09f366a648eafb5b33a27c0524d340eac
zf9f698ba5e7a1dae1b8c36ef90383bb4c858326618b9f2bdc1369dfab005e3ab0f523c50205314
zb12a1e7371e1fc69fdc5c287cb4257c41d6509e71de704ae7c15c8f01f2df3639b2ece7043c716
zf1a343f997de0f27e2d25ca0c6f8ab57599ce7adeccd8ee1d915233d327c004e58f58b610958b6
z682eac8492bb635dca366dc20dda0bbedbd528f07be26889fde29c96f6c26bef467c94badffc8b
zd21ab6e11fd1978cbe35478289fb855fafd8fd2807a034f08daa213160cfb74c790ab79353ccdc
z749773c907b01773957a1284e353a1e033145c30b440b75aad1e7f0acab365a34bc5833a8ee478
z9024c28bf63ee351ad235b117a36e7160ea8c982c2701b571afa49b35c2b071bef75771547ab4b
z8f2e72339ba161c0fe2d6c1931ed7be2add3ed14cad9b68a82d3aad3557104f28d2df5076b0caa
z5cf8a7cb225539d380a89d802b72034c3317369bff41f8816067f52d2f94301457aa61533ab747
z098e2cf4a5af205261ac11d927ac4d2220aeb0b1378a3e5deb512654e60178f563d1507b9dfdbe
z28ec5b08af94718fce4e62dc5f87bca276f25655f31e2195b4a453b5de5ce2630f9f2b27b2487e
z4c8606702598a28d169159159088900d5955534fd388e9317fbd38cc58b90e0d8ce4311aff2b82
z39ab6677f297b691f43fbd81876118a16c62f8ff0791ca8bbac25e813447ca289013a742c8f338
zb3e44024863e18ad15e369aed56e082ccef7c87377d5c05e2580b0dcc45ccb88f532a1fd069eb0
z9ea37cfa8acd43bee4520aab8cffb4af4c1f9e3851d0f4530d62c726548f9a18f99e578a763af9
zbe9f68eca1a60aa2101b4b1fb65c36b428482a0a61ff1f75864a8b8b7531b32055fa5a8537d98b
z1d9b2f84e17a473a5f764812e70a699e3400eef6c8706a93ca809511567b6f31ad3a023385008f
zb7b1fd799e9329f9553196964d97a2ea57f049c4d90efb2eacc50059b79f7f256f9e4fe55a71ac
zfed885518bddc49c38ff52f265ebf91c624aaeba45e143aa7a2bf50077e041e6c5389c9364b8cf
zfd7145f5b2b839279cf85e9326ec1f2d4ae14288b1d2b9c1cdce92f165063475ebf7ebe97725a1
z0f0bb26fcd977856fb4ed6829f720d0682c22de019bcd17c43aa5d887f582df5e55740871db086
z366e4af2929535de6a35cc77598226e86562c1d3a84f041661a87a8e2c8dcb55d41ad2afdbe160
z0f2abffbc44bb1745ea8c58bdee9dcf3a582a7bbaee6f1899c3822e9ede6216aebcf8e13bd4ad0
zd6d8dcd0a4995dcd77b12b2d3d01ac75d448e965117dac397c04bfdd08c8b041ac427b7342ee96
z7bc3c7d842d05db89457ba2ff3e9502a3613cbc961e93ac25b90efc88c012d785c8cee739da599
z2bb8bcf386238a485cf3511f2b1e7e0b5fc359f3d99375af8d0e289b6701f81306342e6f1b0973
z11d61bd1d8f872a3bd8febaf3e73c8841db54c06bd11addbe3c470a5caa0c7e1aab19423cba6fd
z7b897ffe405c688eed983d1ed506d422b6103fce40290b54c4d669064b580bba90ac20465542f1
zf6b8a7eeb325f0ea46c98ad17b7996d585b53661074f290b2eea2b0eb972c9dcac7f452ed38ef9
zb3b479aa1d5dabda5d83963e2b20435e8d4f86a9004a53008338a6eeee6ad106d0eca2e05db56b
z9b70a242f68f005f5589fdaf01569fca4bddb8df9f8a9c20402c55ee8d16ee2c41cc01158f6ee4
z887bb35c59deedc30ee66baa07d73a976f4cb5643b0c02f780af0425d030fa9e9b753ab169206b
za2a4b95cfda7d0b43a6cdba2e60885565c1330bcc6d08ad461af6d404f8ff2117710dba745c15b
zd81fb9b0948dc419ee95e2dd92f08dd3e49d55e265466260392d1a567b01ea4c10f9e7b4e3ffc5
z834df6e38edb0c83ec0a9c1314d7e4d01a52af8b1192b09d79e3423858584f9c5616205e25d407
z9e6896f46d787e5eada532094c7f24ed238b4ca6d733e9f95f412d6e2d1f7bdcfa16e85606fc6e
zdaba0f07be2a3591f3b01ae3010a975bc1bd24324ec84f9c693692d2cd303cbc2c4a3235fc2fe3
z390c77ff5fec5f18b2b6c9952abc1bff499d881c7dd8784ce11de521a642f958a8e57c125180c2
za5217414545927b1134de2eec8b4e88f05a9a23f9ea9d3e603c2c9e342a1e133ad984e4cb55116
zbb459f68f49ef433f08a15c9e6764fc1c411122c6150028ea57d31540a3ba2e26756d7cf240a72
z1d191ebae0a9dc2db3cd2eacab598c9e1bc65cc25f8b4a18d26dd5ed48d945e0fda2b1d20c9e8f
zae4bacbe388f2bdd21e4fab08d0e3361c230d392b6f9d4d037a415e46c82e55e8e1127b4bc2c58
z4da94fd3af4db0f996e0b27e416dadd4a1f054cae1f6c5c18ca222abe6f26b76a3acff36310573
z5a3c5f1cf75c9217c2851dce4278e30364e9332103aeafeab50bab68499275249eb298d247f7f4
z8db337b293d502a07c11d043b21742f386a32597da67da5f24b07cb4ccbece9b6691ec2dda13d0
z735615f7ce38cee82f6754592db38207fc7d08e07a1df5fe900d345c60d1b12a7d8664d4fa0b3c
zfc674a16575672ce03d7f6f20461db9df4be78c72583aec5990887e2b8bab50de11ea378d8eeb6
z1191e80d630787be8bc82124567c70f481b3d796fc4c4239da13dad7821b31d7dc2fb885d5cdd2
z692ed5bb62c5e2c6c23a6bcd38c53aa54395d91783303ba76fce0692fb3e1eea9f28937f9deb90
z9d7fa49df90246e3ba1891bc94d28d6b08e51cb3a5c9ea5ab96db839c8c3eae0e21a75be76ffeb
z8c101292ad794ae1f498d9920b4378cbb731e381fd3eb1dd0900d2f3238cccf1439945aefc7240
z2e2aaee82c65ab50b915631d42037d9d3ae4b060d2c62cb57fbf0f0b50dd46c1efd498c62c3e1f
zad73e4ecdd4074d10700edfd277d2c5a75cf53d510a6af7ffb99bbb442bd8ce8fd0ad88a8f85cb
z1baf4f20bc0ba268fce55bd6942d6a5ea0ef3e53cdc167c474b0ec4f64cc94828f9fbff86ffe36
z249565a9b9b0da3c7a6fb0568c243b1a64402da0ce8b08838fac0b7bafc21284c42e4c9e65ad08
zd07bcf0a9cf09591cbd5bd2d0c11ce972824e1ef86313eb3f2eb718caea3e3e49b890759fd5732
z7409dd39f69dbcf4f75ca0c68591c4486813dfab8d72d8839279fb6b2f59069c2bb86bf4d91dcb
z34b80bb90a95210fe146cb8e99ed040df271223cd166bdf0a421fef656b75fd0b12f775c049a01
z7cdc5ec1851bbcffd42867f9af15be519af054f664150d825fe1e2c0b463e4b41031a03bc0030e
z66dbfca55de85e79cd3a799b9bcc445c6023b7a5444b0fde1a46a26471cde6b7f017c2a3628e18
zf740739d376a661972f105ab47576c3e5eae5b4a0e2b0a6225d672f699c5325cacc3f70228966a
zce55fde1f95854bf200c12981be08ae3d7827aa6ac5493d317bd6bdce6745efe6edaa2f182031b
zb2c7307fbb5310df23011abde7f2e44ca19c86b8f27191b347c4ef86fd87beeb8dabfe71534b09
zabb8a2004f986c14d01f80074cfae06f193987ebf9aceb53ec92180ef6bf59d3fe96d0b937fe65
z29d1f74c96fc2ca49c3c73c7b58a512ea3d6f2220ee3c7f37c6df3512c54ed765e652460c9111e
z15a80da4e435af5c943f7d970002b1d25e839fa1d0537e28a35c3e8df599144e10de9180422b85
zed7ccd68e283a56eebf664ca4bbdd745fe7c2e7be5f299d4aae964914070001f17d4aa1f1e6c65
z5db03c9d1325d58bdd6abdedc9e334209e92da1cd164fb6779e4230be4b4564107cb57463b18c0
z46bbfb6a82c13d03ae0548b73e5017e796eadbf9b53560da56b90d4dc83a9c5aba3c566eba178d
zb517c2ce91ecff811813bd533447bd25e9b9bfd120777f0c571adddc40cf4630c3fc9e00615c73
z4908f3243f66215b71f46a41630f350599499dc644ed12a1f8a0512e3159eed80637ce26942d71
z0f34df6e565e80a659ac9c8ad353256ef18b56b163b25cc9396ab6168e1ecf17b8b6c08f23e002
zd762db6686b3e143b87022c243a3d77ef281ec496551570e3db2d2f6ece0f1ee51c3c29149fc32
zc6c749feede202cfbc294ce6c45b8951997a1e2d695bb2a6bd6d3f5a7f090ab848bed33000211a
z5eb045e88679bc8dc68091706afdef32a8c4a524be7677c1e06dacefe8b7dc16ac8e659e1b9bee
zb95a6cb22132115c6b1245f6a25a95d97bc0fd01f2b5f87475015f170c4be417098277e63e2657
z54c3447ac55817d6520050cb170da412b7a880731cccdc9aa1af576c9c32650892a60521bf2066
zccc7095021eb33b57f315e18ab594b8960d40e00f56f2d79d3ccde3326c00597d2649b273f8290
zec3c585ef67a7d656a50405d4456d7c5fa1640b72179393783ddeeb75f792546d3ea2c56a7055e
zc7d98a6a3e72d5c076129c1ec13f967b49acd1254a9b128c81c7f962673910416904317befe129
z973359b17f8e58e58ce5ce99c0b74175582be03ceb82bf50b76caaa1af595b76eb76b9516bf9b1
z82010f95e7e83d024b4bdd9b6934ab114db00a58ab130919f1baff03035c798f46fc8c2b975c3e
zde440167664d0e05877a8706ef4db7ec3367f574a0aa89d939f1a9bd4d00eac01f7b58bb455f71
z78f330d888a3290e9080e648af62b141998305a4da5c41277470a2d9c10262fa89957c0e7cd32f
zdbcb102451e570ee4590b436bc06e84c06b9ee9f9ada8c34d5f4c2f15da1a4ebf8567c3c08e154
z4dccc85f2d713c76d3477e7e5f8b7e8301522c687b5b6353e06a38c5514619ae1af2517ecaff85
z8341995b4054bac967101ebbc56d535c71f92ef6b3d5b8109b07dfa3095733dc0990b01f203c15
zbae3f7219f335c878fb74dcc0c89e98572a11112236300e2b3611a6bf0d4ad1ccec01e666d6049
z0f290fdf46578e02979589219e1ecaadee322876e7d61a89b4f96de5c6d741b7589ec4e9c2ccbf
zb87d64beb6b1c0fb905e9bb285698bc1895d160567c0aa20f34acd063d01c9e1fae4ef35f2ab1b
zd030d0dd1335d2eb6e54097f9618e5c26359e573d517e8fed2e9faa6d6da3fc384ca465b76f03a
ze7c9f4916af59d17e4d487e7cae75957f71dc8671dc87957a2bda6831e2a558c0d5ad949348fab
z21896ca00d62f843d5e9e254674bc4ca956175d3c5e3646817e7f1abd88e3c765a0e8feaa8affa
z7b2c704e9643e841bf1335422fce9153af31b8ab32f4015775a3056d5b18907d2ebdff62ac152f
z52866b09e0d99501f54d7573ed7b1830c30f333a540bc20a5fc6e7fb1525d91c10e94f3439f024
z6818c75814c7225c6ff87d376a74b7e0914dd5f49c9a8fd07f29afa4baa509ddc192754dcaa9c1
z635aabfce3a672fe7f2439b8d1bd635928c87c6a16e8a60e15fe5e6c80ebe85cb35bbe9d1a8d78
z8b8049a6b5d57e64649803add979236a4141cb45dfd6b006130f4b844fb954759841a31b9da544
z9e0076fc1d6b261d9a99d20586a5cf459cef40a386d713f7aeb21b02acc9e40b9a44484116dd06
z42f9fe5d15f2840307f7acf9e0a35e2da13a1fa02c1674df241f50ecaf55316ce41ed6af8ee453
z51b4e9faf66603ad4d2fda856b396a1c14122097e2544ef0ce2da7ee2fc619ba565c97236415c1
z22f319ab114c3168edd1061825d4df37f4d762fc04c9061cbbb68a0fa5692f99d67eeb80cc4fa0
zf932ae717543279fe486d059f6476b525bbae54916fffbf8183e34030261ab618a5c86669ba931
zc264fccdd8b84333be7e1db1eadd3fe7088b657d2ba4b848052a3ec1918ceaf2811b2674a92692
zecbfc41525721d4fb1cb4b06f125676bf4dc74255d78a666b2235b56fbecb4523827e8b0492d4a
z526571a00929231af2a52a8dedb999c9b3cca428ded77e5700c4b9d7072ce8da0f73b1398c7d08
z976a60b30d41bc850fa52438594864c6529df58f9d91c2795d0a02c22be720892a74aa0198888c
z9d77d54e47deff64ef192c213e695d57b24cc657c8e32beef3d76846fd5c21c66ceb2ac269aa8c
z7855fc325954804e6252a6f4279bf34dce3663fdeb56e30c09653dbde98f41d06c6f2e5d550ad1
zfb044b79e908438a111cc47b99a73b43fe464afdbd34bdcf21951761812e2d982a819d14d3c06d
zc1ca8b2d864f382f4dfb1a724266e039175c40db7ec26394b5f456d547015ba29952e13ffef778
z3b18261f4926b64e5bea43065907ef869b7e83690e1f082ae1ce7f7140c46090a9a758421066bc
z7cdc3d2db4a29e9f4db0c899214b8a9a13e4f9bf7fea8eec55194fedef1e8b325eddb7d613e704
z9746329d55310a29d7e7f9c8c41ba9a2b1c212912de9701642db9b6007b92fdfe82945c2e262f5
z60750858712c5fd7d100e2f5f9c0e651b3c749d382a036641b9d88dabdbdacda08bca40c08baa0
z2672a192fd22e01cca8e640a8c4eb5f1a286b7a57aea89084a992e7aad44d714a20e05ca5221c3
z8f9524b7222d27817fd7d3684997ff7ea46b7a5c02e83cd520309ee0a57a407abdc4ecbbeac711
z35b910056811100718b268c851e7139a277f8c953d54078538b1fe53bf9d1ee2465028e5bdef83
z4de2c721fb56ebcb6f98989cf853ff3f7827034f9511db4c523ba5ca0ff84de7fc58c26c3d1ee6
z715361ebd35caf963817ae699753c35064312a1f316f7fff57702cb5f398b6f6c32e4c8337ecac
z5fc6c3f1c3ca0d01c0c8f2da68e698ed9c079d7f6c3df4e979e351f09ca67123917e083a587c0e
z178780e3a292b2f4a7bc4db54df05bb82151e8d993d09b72b41db31675f4c5d8a61bdcc529d35e
zc382303f05884fabf750be9e79543288783d8d9f8089073a2665214a1e51436126ef7ad4577175
z8df83bb04497b98da3b4f457d5cc4acf57ad14b61e97a074f17b6f7e8364c172868cbb8763b0db
z87349df24e04ca731fa7956dd09231e8c64adb81dc5889a9a37bff8cddcd632e272ab90a8d8fa9
z84ee5a8db5073749c7254f466b3d6294965bcbf1758b9ad3b8acf6400ccef17a9243608ce60cc8
z1e9fc92c1d000740c0f1f0678e52e9a8274133607511ffbf5c3813443f52f2b615438e873dcda1
z6d9fb3290047a2878d602514e8d4a39229e56c06f741e081517017b02be8090620781c85f96939
z5741921d840d2ec1584c16b8181bccd106b85a74480d4ae0e9444a43dac1a913c8f46333f632e8
z8eb4ca9880ff74e394e8c97e165e59c14b4078bfa939343d2848e855f46713f84ec6deb8109a13
zd640e016ce20fb7b19bc1e44734c71859b3115e43439dba1c97f21b49b76b6b65cceb612a38b5d
z3e05039255952844450a9b15cdd6c3f6c4682789d4751ed17de7ea00093ee9b6f5ac4ff5ead8ba
z7a062b31ed80a1c9d755f51da747ec6d71081d3e596ab3613d31eec7be0e3ae2128252d81f4462
zad673d26d8a8b1c4b18a47c25708329405af6373e2af33b3889f4321989311056911f0cae8eec4
zf974eca41270c23cc0704133b5dc734f59c890b265da5277c1aac57bb3e5cf045af2c6aedb9e54
z60f08f115cb15383c5f7de89951d70c559914b33c47f98c380067b316eaac18694e9a6567ed47a
z0e8e7837cb30daf7002943932e0d6122cb7a80c8b14488c60e50979657b9e43198c7da66e7feb0
z2f41488b3f207128d5b3c60e39005ab0e46f471c7275c9e7b51ba61f5ea7c680941285c6915b4a
zb0ecdacb35770e59dde01cffc0fdcfdba11b0ab85f4b54dde36ea8a6e0664f0b6046af9d36f4c5
za39133b15293033bec5485bcc7fe09ea5b8b7678e75f0d611d82acb14628e5916e29b9f57b9d21
z8c22941e8df9b4efd614cd29868adddc619f46b91a885899bee9f43aeef1440edcd0ca59113efb
zfc777ae556be79336180f1497199e3b3e1a4508848629795642cfef52ccbbd3e8527fdc4171750
zabce16ec7347d25f57b16b2abf538650e2dd086b629d3801808661979ada59f040024de456098a
z83039f5c1b9ebc9337389f79d993420aaaecc51153f52ce8b430b2c86ad9a9ee7921bd26b9c5cf
zc56eafdf681fc15bf94ea4cb4b36f894f25b4fa8308383ad24c72bfde348565f3e2342194b6905
z3a16646d10a13533a66bfbae1144c281db3a3ef49a0c3ffa49d2504928aefbc7207633cd7381e0
z61bb52ea1447f2119e53362c882673dbedc25b122588485afa98b4a585cd7a936d12d841821d6b
zb383321c5eef15cd7bfa7ac6a2ad8a6048ca9ebc68fce12a69d9d10e29847508ae33eb85eb4d1b
zc6bb547dea7fd4684b6cf0fb2effa5c863c1fa22c1466d9e34edd08d5bdc84a12afdcb1b76dc8c
z062139cd9a26c1b8ff9df57cb5c49ae197919cb403751fa6736064346306779e9108a9aa30d143
ze8d92593153f0ac7dbf22633988e1fc1201b3cc6fd8b88fdbb1581be3c45fa829d5f7ae6fc1b91
z33d6201c3989e066df8da377d5edffce935096bbead6cf651f08f31c22a49112337b9d3abbcee8
zf5e80a2a6b323d3602627aff6e73c6fd0914b109e6e3f732eadbd6d855b98d617e6544e31cd52a
zd0ded8bce6fbc23ee0e3ae31639ecafb83694d1e4ae396f9b9b0be085599844044f014883fef23
z2ec3a47be48ab2845377997e6c9ebefb3ca154ca41c0c3e3fbca334141aa665fe94c9915057e04
z896cd90ef06f5e0944265b98a09aaec5c9cba53ab99b32304b1ca96b96a9e6b458342bdee54027
z7d8107636de601cd0c762eb68618465c2d0b8af5c657a0f92d77caeca6c8ca9cd3dc1bbc4ceb1d
z750aef8d793a13a6b854fcccfd6f4b83cacfdbb7eed3486975519b878ff18465a77e513bbc8beb
z0a5195fc6a74f47f8a57903d747aa6324e3f8f8412e7644592e68b7f0992775f27b532048f1f2b
z85314ce1426f0426d10a10f1e32c6375f2fe442625ad627ccd0dbbf54a23a5e66340033abe56ac
z5c5dcbab02279e7286c5a1aa72e2b231baadc356fdea256bcf71f32046b8a3979ebd4d86775d78
za236ea02c5ffe1dca7ffdda52e19daeffbccf286b2503ed93147405927ecc30cf37681505edb3d
zac1f49c2ed4d210cf2b73433c7eb6e4b0aa8c4ac2ff73349f1ae1e2b269ac4562848cc0e161d96
z05d1825d34c590c5e59f9b637f6ab031e0148fb88b44c106ec7a71dc396588edd9b4a339c634fd
z9e9a32a517ddd1bb80f24eaca100d68dbca751674685b47ed74f63d0fed4c472b533b1469563e5
zde32a3ef6971d5cced91c369175f14ad91c5048d40dbe3810581f8b0f4cc9399c38d4ebc00c70d
zf09584550fd9bdc216522250f975f359bbfa81334e17c66845779b09521d89fd137c9469f5e86e
z07fb14acd81efa79e238a706085c62d2e0380f2f7821833ae335d4e1b6ef575ea029156413402c
z9b2c9eea2aee245aa3d89d25fd38cb731663e61910a65feabc48c2dacda416020d5bf6465d115c
z4da1c5f13c66a0ed811b447aa26eb211d7efd76ed415aae66a5beea1a240d60e0170f3bfb81f96
z86703135fcc43d2fdd75bab3b949d6f3f5393957ebc46c20512cae1dae06a5ae702d541ec11702
z0e5b11d38487334bbbf1ab65bb665def85474f101290001979715c8df138e3856ced78e2c19889
zd5b31bae3acf786c0139d4055d4d959f716caff9ef93f499368638b85a0812fde9aeb48f5c721e
z4c9e8475cc5cd5afb7b645a724f4b0b2961e7bedc5d3733380945b42f2aeabf840cb2284bb3a08
z3190af6d4d6ae90f933caf95f9645ad4a23a0787bf11ced68bd841c690aea1b3580ee5da10e54b
z9565394c36f5a80e11607a7615d6125ac0b658c970d74e781696e2e3d3606cd7ab5cc7b231f0ab
z2afc517ff41ae4cb0c4b0389e2703b7698740168aa233e9146d337da5c2bffe6d75c672c6c5814
za52b85b04b6c751d9a830e7ff29b0e49134c6312c62e12697122b444b3aea759d6de08a6c89920
z87e770afa8984bb1a7942b1bc3c16a8a9aacd6148b55af10c1479db57a940e9a3fc68f114c7822
z4312569520c6b37328cc2dfae64202673069b82345a81ac09587e0879579ab2cfdaa58c3c58132
z2d3fa462b0c27ed85cd3244057540e95547060471afa42558a43bdb95508b292479ddc6f9f9ced
z2bffebc7efc1305e7e74c46a142dd28cbbe0cbdea7383833a386f16de6363af7495e79f9260813
zb3ff9bb76b2134b42c75657dc2b4b9035855340753c5448c8a2626e25e4280fd67d63d7e007926
zfc1d44ed59865f95910d81042491a438ad6b65283ceb4d8d4fd07a19739a2e34d8c080ed3110a6
zb8e1c43a840ea90670fe5b4e281fa8a743d198ad96f99811d3c19c3d1858f8124efae1e5d25941
zd219b4a05533fad1d204fbbada1793fc1fb188963f17c7caa6eb35c792ebf5e99715240a8eb2ca
z920dd3ac5d74baf1b50be0c3e7add3e731e51cd33ebdc9d6d63bd56442b93b3a9072e0eff32fa6
ze2261e09b0b8524d25b20ac21a00dddbbb8166304b3d8794ed740ecec64c1cd91e3681255a6d67
z725e42f20430b89e464d3ef879486cace4aee6648f045cf673d6716bae5325743f23f25c3d79a9
zb18525527a179fbca4776886dfaa196f5ed8e4cc2c8bf2212676420b21dbd8109ab2b57f31413a
z0337f1c70d6c2fc6a16b6bc809d9944e7b246732a1e6c71d30c37725293ca3dfbddf33d5b98de7
za03bea0e9da153e6a16399820453cc66a2bbf330d10e9470ed8dd1d4cc6b5664a1ce6730f10bf1
zd846d2cdc5c63524e8bb08423693b6caa52e91b0805b554ab9561857b0284b0593dcdb3178e9db
z1dd8f95e6450cad841f4fd6e1aae84d7668ec913342fa69247010933770e2af5683eb9806d41de
zde7530a9332cbe2576632438e79d06a5791bdaf54c5b631f23f2a6efeec4e750e3bf7340d04c29
zcd60a9c5d5f79a05af716eaeff7d2d9f7ce6e38d3ef483f3868d8f7d666de23b6c1a257485edaf
z84872040727f036a4e5843740eee18f6530bce7db11be5a64e821b530cbc53dbb9ab51669659e2
z8b7e1aa5c92e22f348e8eae541a81dfde4525c9c8eee9e1911a514c2b89b7000ed8e5b714b86e9
z58299b055d1013cec183a137ec2bcdb126281766249e71bb719fd94b02576e684173d196a42c61
z691fe77bf5751131839602de36cf1790cc5a304f638a5c8e65bcc519a50b7a15d96dd40f5058a1
zbf036583d8f0c5d49cf86f779f6942f42bacc5bbd5b2958a0a9f51e813cdb4d065c1becc39f887
z1c356edc4d5d7f801f14d92324ac82128ac26b9daf8dd1a8b2c3ba9ca0a5ca9f11a4a966c4cc4e
z5c1cb56ef80f81e7142f0138ba80f7adecfa51405ab572d9042047f647703154004ad460aeca09
z50cd9d43818861eb0f1584ffe01e1a041e95990dbf151d6081ede3bd4cd9f505397ac4b17a6c19
zbc4eea31a4b7e278022a5fd4bf4bd26dda9077bde3409aae0ef8ea2af4b3938a517aae2df281df
z395049334d4404cb4c376043512894c7b525b0531aa789122dd47503ea6547ecbb76b1d5750005
zf66035d55c3b06efa63da738403d91feed8ae2aab942ed66792bfc9803856b00ae5f7794e71d83
z00df28267baf159f2c45761aa63c4bf4ea8af774630e2af11c8502a632f0a4112f0eb987bb8300
z7f7ea37ad6f5ae64931ec2bacac98b808ca5c3b80a813ccc42c4270894c2a2a4426e79787012f2
zf81ba476e99d7b5c2ca66dac807e122a936b59b8946ab3393030cb88350096217a5b649572811d
ze2de2ff43e1065b0a03644df449d7a8e6665965541cac04ad60dc66323bd977e6865782414879f
z21745cb4dc7f2d29282ef406ab6405e557b6b63357eba437477b8db427a0f519423edb6545f68d
zd51c4957a08cd8cdd15975920e89764eb6edf1a9d1986574110d0949c55eda6dafd22b7a0a4f59
zfba1429808f131ea0929ee75a001eb1193b6fc034c575f0884f4effd4b9d416c9f26fc1d6ac9d1
z6dcad93bb4b0ea75204d7507bd7f930466f05241777cc41f0d09eec7bf75ea9abb7948c4a4599d
z360fdc34f89f715f20f8d482e8a47db34c5840d042148bccd27614d552ada221a8b675d7f2bef2
zce0d1dbed7b21f2bf683f976185e2db6051e6606a05a3956e722c6537bda5b5cfde98ff3af8fe8
z67ddd0e8d9c945a73f9d14a11bd33f475063384be340c76828d5d5369abaf1929d0332a8e0bc65
z6e4983b175bfc3fd4d410fe9b38f0b10c56fcf2b92615e2af60b92431b4831e9ed8a642910a6b8
z4f1d279f9afa0b255a13332f2726a63fc1b7540a3158ab60bda327fea35da8c3666e5a4544ce95
z7931c15fc08641ac60a019bf7952411a21c8ddc465aff148eaefc538dc49cc2c20b19d56168518
z0cf3dbeab10a5bcc39050a97e05d17fafb77d682e720e3ed9b8cfb5790c2c50998c203d4c785b3
z33bf42cfb01206c9f4a3f3b64706993af5ad4d6ace9630ff25297105178f524e8c0a1be2c00e6a
z8651b79f7bcebc2e62c883174454662d028704d0900024a942a35ce17285565e52fa9c2d83f80a
zc03b459add8acda0e0cf00c5da9267991cd1becd5a35e3b2ca9df8257889fbe3b65688561dfb92
zfd153bd17e70f7f3d77dc2a7585e94efd6429d87b3380b7b6b28bf44d22ef32cfbbb609a2361b2
z5dff67a5fd7fb644676edb6692252d730be8dd25090b8ee5749dd41a05b990f87afe4712b9e652
z126663d1b0243ca7f2359f237043b3df78543687384cab9b99d9094c92968de46e61654486f754
z61fb6414a034474b5a66ff66eded9439510827cc16a76ff1189ba546cf3ae1383793d29e467665
z45fb7562c2618ef2f037adc5e333711ede0802dcf74db9a354303991816037df4d6200a6a0ba98
z5fae136939ca7ad13f1a71f378992f95ce48e0fa9f7aa151d04823f0c09e16a637a2e2f999b721
z0e0004994785880ed55ef8e5d194fd04da2ff0b3e061266a93ce0a66bd0b668f07a1558a1b87b7
z1b6382c28ec862a192fd26699e841a3f01229f62445cef2708f3b7f92b0e132256583e783acdfe
z162a8419b82196f93746b0ca626f6d3694d2fa3a8736eda59a64dabb8dea01b792783446c7ec62
z4741c9ee48de90793fb6bc53f3b1746ae64e7687eb74f4a3eaa71fc3c17a2ddb2fc9233176b72d
z655130b7024365e48d16a307a800fafc5444d49d4751cbb22bb6eee6e1189952486990d90ade90
z16d8602346375e1d329f909bfbd841dee6ee5c201415b298fffaa0b8adc7bdf519be8676d7f5f4
z93344ab127fe8fc52026982604dd81108d4cfa34e06a7c5666ec8ed15276fee317e2fd391e8f1b
za044a27d996653804011aa512a3764e496ec98ca5897dd3f2f526b2a213a93e4347eacfe3d76a1
zfb94eb0ad93c819669108494c002ef4be8cf62888f8775a47e7fb69aa823794adb3e1fb5894984
ze89c4ed49354223c08a3158df5515f6c07dc4f811733cdfd632c8ade008c0c8e40ec3077525644
zcce301bd37525a137f744eabd02f242759e3307c5c9054a3a5de5d539a9fdc2367296729414212
za8d8605af40552b0ad33bb4d7ae09fdc6242f587ac6d9bc2e32c1b5a18df13e5949f341d7f05ba
zfe1251f0ecec1a7662901bdd2bb72e3a031a73ff639bf3caee076a8f6082d70ae6b3374f98fc77
z2f5e3b93c44e15da948e7d18595748c497f18db7d3f68eae399deddc8eb83f6821ba8302008ab2
ze5631137e189aa08f29c94a1dc72e21e6539d8c807f90ed478c9d403b0ec43a1c09fc200dc5cab
z16a3534c9115431626f19a4e86cc265842e72cbd50a6eaa094e9f71dba23049ccbe5da47a518e7
zeed0582303ca2d6bb94c765e102a7e1c51be6d8cb953926eef0fe463bd236ee461d163507e7921
z667da0ffcceda5e4c06a40fd4468723dad9ed37da4aa326d1906a37dfa3c838a72851c2fa3a82f
z3922606163abd16211a18ae7a8310ae95e7a2d22adebb7b4f1e2392b9842f46c196cf3611b1360
zefbfc19bc72cc55cce3afb7d58ca37e1848e490434573e888f0d38cf47ab736e2f8f3fd47b890c
z7bfa8a7a157b419230ecfa5dae645e2c85d2c778f20cd2084fa2429304c257c1195d1b5ea436a1
z76d59f198ce935ee1249c58aba7bb53ca5b7c097d64e5196f627e5dddc805a82d1d45a3f7b6eac
z532ac940150718c2a8de656a4a844883288efd66e3028c9f26ef1a02dd7d66e6664b0f44e3e154
z475e7926ec70a9cdab6f348a4769b130cc8abf93ba3988cb275cdbfaa8c30e888a4c04a4278a31
zb7508dc3c384b9346d1aa2c8ec1afab1681eddbcc7e54a0b3c66f341e9a53bd4096614bc1531bf
zbe53d695cf0b16a54191b06cc373cd7b42506a7fa23b95d4bd0d9beee5a5613bb2964dd1216fe9
zef81e2f86923f90080eaf911d11d95cfd111ff0ccaec1725c814104f16c4560c93e0c7498e09b9
z56dc1b785a0d7ef2e897add4b3099c3642c10fcad5d0350147c32bae864bb0d6afa815a110807e
z4571b2d4e964d0d7b0df59d948bd2d8d4d651fb0639161abad9b0362a05df2b3b97acd8375c52c
z2c9d03f429a9796987ea82899f6d105265347f8b036014647c06365764877f4bb80b89398bf887
zc4c714fcfc45ee5eeec0be0b6c899cbfceeaf3d1e9f4ccaccd02e8a05d827e9666bc9e5d1f9999
zb43b4de1b4bc9293e77d4984ce508bbca340b749d072e2da1d03e12a9bd09c2a0b2fa5ab9a9cfc
z189944a3041fe510572950c85e1dfef61c32eac3d0a58cb2e619c9cb7b23633ea6350835e57e30
zfccefcddff656b8cb0a33f34ea4d1e661449297e9cd49cd5b64b2b886c9f72fd3e8528c526eb08
z1632efae2b02b3176392d6e037a2cbba998e5771b2408afdd1d89d044922d5c9325883faf3a744
z677fe08ebbb749e0f2db2af49e79f0c426af29cd10b0e7bc58abf190b8f09189e5abfc14832790
zba5ef6a0ecebb3089578b821e28fcc360ccc3de86901c11f80f83b2284da12810bd325db5677c9
z22c0c9b8b0231f975c89da04661352ace6525428adc121d7d8524712e3f39c6b3d34ac31c91b83
z23ed18c28e2e77d27f258ef463c95c8e820c8ee53b0c8e1cf59b657e5b4336af6591955587f843
z5505eeab19a2fce8843f7114d518172fc5d63d3ec21e10c230787addc2990f4d92118e8d8c8d4b
z1564a60e9a827f2d312499a1b887c17471d95fd65e7416cd3a2b37bc7048e66852ccc04d8581c9
z326b220613bd761d1fd57c96abcc5720d23140670818781a8d5a4cb17cdc2639463eb5543add5b
z47f20fa539aa1cadc9a2c4062454eb7a1528e89635925f9a6a911854eaa1f581ee1819127b80a9
za037f5cd5264f98457d89da01e60bfc1fd9b24f26fd82090d595844cb912af93033090edb76bd0
zdad44ba494ef2eca1073be3feed888efb8f3c667f1708c6a0ccb2b3f0b4d712b94a1d10be3ee58
z79c3f89a55cb54e66ae38bbfc9caf2e574cb785d4542ebb91f133e422c7a2dc4bac5677d923645
za54ab68e8274efd41e281b87d58df0e5721c006c369a749710d70444fdcb69d74d03548fea2b10
zb7238278c748c40f1bbdeb9d3b8b0936627f430ad4887413756d251a8c0e95a1f1ffb70ab2c5d8
z4693b400d6b90d17466f5b7652724823a43d8e2e05c59f140ab8af23f25b1716670de8a6ac4f8a
zb4135ded659d7939695e79ab57bb4ec36df5d5b594e5471a79553887e8b24da73dbc849cfe3a1b
zcd1f8beedb0492189a58e4e7f32ed08907c65d0cb051a740e63d9faf01a01b77973407d4df3cba
z2cd055b6dcc87efc1175960c568726fb8a4e3e648758b77c0f0cff82315be6267d2925681448d2
z32d02cff9de50b23f822d53fb3e05b5cc4c05237c2303779f0298496b1a56d5b6f535c4ba7ca0f
zae9ed83a1b7d49a38fa4c5939f7d2029f26a7a15918c7764dd1da8026f65d07949c7782e1d72ee
zbad0db51edc8209a5e8e7b77fdd7df81d6d25a624bd3792420c6fae2a6e8cee4e1fd99dfd47eab
z33ed0311602ef246924a1b815e5cfde88585582a75a2396a51152cae386b3eaad3e0a7af050fa9
zcfb433fd1edd9151e3953c5fdbcc17c64fa2286525493e3baaf4c60e29cdc08715187c78ed4258
zeabd6b2ec24b209875de77af882105d45d70b71e0d4dc3ad2499d4b25df0b0f7b64b433123c156
z67c33a8f8c7f3830262bf0e360ce906e4c6730e85c0bd198e653cae1ba04cb9a8a2e2f5ceff46a
z6cf407e3303b4eb8ba39f756a1119fc460bcd57043f1d272df0352cc2a69ea436de517e87c384a
z120231d02bc875c5c763710c820ec06d9882bcbe45abafecade5769cbafc18148f92027c8cb062
z79c381bc838f980aaa9096c4988348c9c8a94d24e34580c379080663e2a282d0f900020de72488
z997e1c6aef7437274433970a9a9eca6567e5ad56fbaf8f84c76b5ded33f31fa3c2cd324e23720f
zd704e68bcf3c1f9ee3cbe86fc929c34ebd6e38cccf383477f8bbadd312ed58606a378969ad8352
zf28fda34b77dfddb528fdfadfd201ead9700aa8e408faae0b0436601d5b283ed8b804b5882e17d
z0ac624fa4abd7fc5a33ce5a8381fb8e4a287f66a8973c2a5618759cc6e16b03b8f1f3d84ccdd3c
z0601439fa2d1b9686295c5f3666160a59109485b4658bab905e1425953844b2fc31deb4c1456ac
zc5b20fe52f2694da55c14c5fc7da5b1ff4a2a9ca62bdfc2302a54ab0dfb62b5e67506276204464
z7b7d6a433021e35a44a2bd2803acb8647c2291885d5702ca11bd483b02a81bc2e484537572ce5a
zf7e6064cf4ae2573136d6004e32fb4622b86dfbe3b39dfa3cfd77788a0fd784da3fcd86dbd32d5
z088269b9746930acc45640bdf542381229b8cda1e5571e09da1f00d0c08bf76e06dac3ff19cbd1
z42ccd3fe0f288f13827083cd59bf9d629f38c519fc0f95987d452610e3a1125d69bc77e12e797e
z8f754452b984b6ad3b1b71f93e14dc01103a159fe473d10cae5c9b484ecc3a69431d1ee155c0f5
z98a98893e656f599ae16e9af1e8a5bc6286d837c0bd1b98878a2f2b5719fc22f497668591f9da7
z90916a7ad8d07dd45826c29fa14d6af33745211e672c637c48fd6f2217075b5ca6bc3410881828
z0680771b215b999133992fc2c66a66ab5053cde4f002024518589bfe9123fb2907ed3d233d2dc5
z6b7bf8129b355eb11d91bf1e3ccd731ada3472318bbd6000ff4be3cdf4435f12bc75a95543568e
z42f4da57d267e500ed1850bfdcee3d5a1ddc841595401fdbb1b3ab402bd5c7db44c5166b0749a6
zded1c16ee7c3bfd13fe5c911791197494b8370d6f48570bfd75869fae56d367c512cd54c2d997f
z79df059796ce978de9687a9154d2fc5c28e9c75c00077119c697fe12509c2e214aa076cb1f6aae
z5a80728aa0911da60d2dd0e01b8e11dd6d036e44e818e387e03bca5b20c510214a329429c84092
zb4aea96e0c144d1e9ef4ad414a8ea4d7d2816d8a227cca55e766df30213e1912f78fbc8fdf6f2b
z97223f620546bcb456483cf27271cc6039a300fc5c939f71cba71c4a30453974f223d9fddd8de1
zbc9bcf657cbaeb8a826053123ae6872d9366d55a27746869a30a2ceaba60e3af5888a3aa92a8b7
z33f1920bd3fa82156b59ed9784dca2cbd071f885a7916d9d49ea8e1ecd116d71f9c81745f67e02
z45ccb4990abc1b76f056e907efb2d7e428d0455461f03fbf6deba9d508e29769a73517fb706982
zc3eca3ae0d5420b6c12f87c6a879d800bebe6f8d99699814448993798f1fe540f0063f59f515e7
zb07d90e20a1478cb82791dbb786664855f676e9203a8631c59d98b41cc983c0fba1cdd72d95647
z8acd45338112f187f8a890b8821a53946223f0edc1ee270fb06b42611200580908544eaef41ce0
z5d34b182e220a458b1eef51cbb42642ecce3874d38d16a209c52bda4706a532cf38d585a7d6094
z904d3b1d9d42d596922ec5a5c727cc1047b7e7d4acab18889e4cffdb1374c3d50dc717c8f079a1
z3d852232a031e8baa1273fecb3523ac77f17d75e7f44ff9bc7f5e8040b117ad56fef70147181c2
z3d0a56ecfd1078a5b6418194f65f9f7317110e65bf77fc6c4753178d6d43c25d4bfc716157fe03
z68221ed3013e7d3a7a8dc20d64882ef0650b884f9f21aaf7d8c09d097829904ea862e7c3167b3f
z944ca0fa7c5799a5a7e7e1f23d56931ebaa6bc54b263f267a63e309bb63e5d6633d87a45ac89ec
z0995684d3255be06edc0522d70aafe994cab25a43e9a9b169a6743b41f4b5aaad120d4a1a903b7
zab3b8771e7cc973857f784da78f937663991870b713b224d69642f73a70b543a57bccab376593a
z39cd9e6a61abf7fcf8c00e5d21a948d4380314e6281537d38c081e8555ef7d118160b2fbcc5c8c
zac25b212cd60ea25e164d6f7a67ee1b17edc36f5291885eb8c0b1276b445dca722fc3029105359
zd261abf490f0b074a7431ada54cbe5881a277cb365127e0ac89100a048297a97a092637881c790
z821b685aa51c8e92ca176e84af430f437c854991f8f1d2ad91caece9b1bcd0cf57aa2f7a5b7d2b
z24f92ea17e25b181010ad006c364cb079c4dc15673ca43e5bdeea6396b50035c2ae3c84edb5cd2
z7bb1d59b5a41f038b2a24abebdaca490017211ff91601d91c0b065f7c6c578dd9eed8bd2da0670
z79a7569b7f7c6d3d14547bba6a87e0427fe4b8523a3e3d3a8b42167f3279d0779b7c2ed5033c24
z595a83d8dadd11de9062e3ae50e2213f81045dffd2db228c2184f45e8adf328e80086521a18212
z78c5c2cc4e65d9d91510de4e2bc739b4abd8ae8fd78f39eadae60543c1ec8efd4ea1f693ba08db
z7d55f6bdcf4e0027d7154fb07fa198169bb86dc8a07637e69095ac4deb445a48bcaff2e4a746d4
z4a7e94115ba5ba22b64cc6600d49fc1b50e7703e3c7bd8c80edc49901a37389efbd189d08d544d
zc0625cacdc3d3b504f1e60e87ada9abfa7c673fb4aafc20c47e940909a937408bcea81109b4c06
z1c0be88ca638bad942b96bb51c535c881b0e5d71a541b0ee978c54c337a0299b4d5ad51a57059a
zb09c0b186ce9eef812dca3e8b6b03924e13ea764cfb32f0f5d94f0db383ffed317efca34a690fa
z33a3b528d9756ae0563c5fa571d1e5689db94215fc1e28ac9c57e80b952a1db881162130aa45ea
z6da8633ef161a42fd96f94200083281df32fdc315abbe63cf3a5cf7da376b2bbdbf3b89dda0e85
z64878fcaddb977c19c5e0b577dd51211e6f58cae59fa1983b3563b240245a264b3d601939388ae
z1a054f185f1280f6e78d4e4acca9707a955b4f62aea44989e61e7dd041a4239e3b5a65049672e9
z1c18eabcddf099da4f088dedfec9f1dda6177761cf311ff0828454a7ecd0b5f19894f69b28c9c3
zefdcd45aaf1bdee524ee4c51fe818fcfe8d9457d84b6c7266a858337dfc677ded9cecfc7d745e2
zf46be2b594fa43165ec06f70bdc94cf5b4a5e0867889137531bf93077e481a78802de54de4cb6d
zd59810b97ef867943527c3cf92cac5d077783c719b7ebcdbdd5200bb144430b7ce86bd8a6d8140
z4ca3892fa79892bc35fc82ed818a1295ed4052e0ff947c90b2163f2814ada5c5bb50603e89084e
zece36b81df44be5d5d53a3b226259fd0574e9952bc5e05a61b3b632b6d0d420fc90c0bdc568c5e
z727a618432010f29f590249f48b9f265ba71b3bc8927f742d59b614658d57db471f66d6bc4262d
z6dbc8788c1f1f7dfc82023fecd8f4524842bbb80dd609511b8e86515935ca984ae7fc9d8625e77
zc63d15f9b9aa58a2c8b0747dcc67a3b2eeb38ccb2b00e2164e6055b8db0dee2534996fd8002608
ze12de555f1a725b7476e476d461d174e9b2044e361ded16c741ace6296f641936d873dda0458a5
z82d4e7df50949655ccbe1ca1119582634a298822a8d77d9d45d07449158be2413a53f8fbe58f1c
z8523fed8e3357a68d73c9e19b0e96ca97b7083cba37f621fc8b0c380f8a05d71b2b4c2d8642156
zf5e13f80bc359c231fab8c0e2f9cec70c5b65f33c662ae822097484f25abf618babbc69e6f5268
ze5e96dc4b06919fa6afaadfbcdc49f2693d5bf2652316f8004e27ebcc8e26c0c712e8954218a72
z36e570a8c1e98ffec820ddeea9b30628c2d6d4f40b78f16aa6055360c7c19b2e262c6bcd7c66e2
zf8df5d74f615bee35719e12810646100d75188dc73c6930109f1656f77170b531ffba100435fa7
z79347a030e74daa2d735a24205db4d587d7148464bc0eccb8535a410aa6ade7f97b545dad22d1b
za2d638cf046c60cee866c215a093b032ede42975ae3bf53961ac7242105a2531cc7031057ca42e
z2e81cf3e5726b92ed4a8cb3fc8c894ff6f601181d137f0df3392c68eb1e1e62fc5357a17004d43
z7836e50d189aa5a238e860bef4d2646cd74ad5ba94649f12b9a9da1e421f0562ff20a63475d11e
z52f9429bd6e500ad1d10a4d86fb5acf64050119c4ae322f950d89c4557986bd8f34e9458838a3d
z6bcbaed6c058b873b2ef48af6cae0b4af0aa68b27e9843c5c61925af3f4e5d9f81e013e4cdf7e8
z945d2f061df79df5b789a366c69deff1e0afc68e19c348ac659e648e1ea06af6ee4fc21a9d84cc
z9cd858485ba97ab4700bba020ba97d7344364cb2036784a1225b9db3506e03b47eea621ed8d84f
z3847279191dbc33aaed11556aff814f5c99af9273d382f5e650eefddd1b031a14bc9e3012ae1ec
z68529872c05cfda1566b4a77d16ffc6d4d9b8d03d411c15bb2dca85d27a63c00ffd663318cfc37
zc445c30cf861f00378da606ef8d16241d97112432414f8dee9a39bb3a8f404e678f3e88709ea70
z904e092fdd812895ffa0c77c32d6c5b7afa8d309fe5972758f8730ea65a25923b1e72275410610
z3fbf1def685776ff75394fabdbfe85e2fc018cbec6fef60f1f0da86df6d7bccc9352c1b3548a3b
z85d9bb9dc9c3d199e5757cfbbbbb2d53ac722186254b8dfaefc0e5bb80ba518e6e4287b3ded3ae
zeb4c5fcd7a6dd202611216752a0ed2298ace0cff178ed927420bcf0e11aeea74e3307d0d1aa339
z2db3afa7943e6ab7ac2e2ce921afe49ee0dbc25e3978a26c5364afbfea4bcad7b4138fd92e5aa1
z3b688e58077c4e72c7f88ba710ac2f7bd038efb5edf538e739e20629250262f932aa45f795987b
z1fe3796f52ce50ab2f61b4d4006bf359db59f1a3e2619cd051c26b6d30cd2461f011d26cb0822b
z5bc95f834db829348e6bf38dc21abe06be92fe434599273fafea70b7f10b014f975004a6536bdf
zc5b4452e35e18e3cc5c2a74289f4e57c4f12cdbbf0a2274e86dcdc7eeab313d69aa9eddb095cbb
z7bcae349d0a49f4f31c1061a7a0cf9ca60f47c81052841e8e94d55918a54aa963fc56347d94508
ze53aa1a786b4f65aa831a25c5330edeaef44c2f3e7e99b2b273770af37d42c1b088c58b835c765
zae0427d4e69701dee6de70e12c2b4c06682b47412e88913adcbdb8f077e991a13a297bb4265d6c
zbf27633b9d3dfcc52ef1fff459b1856be0be797a6efa730acde705487081ed067a81a766c1bc86
z433ffb5793fdf3c93c6206a36ee63746ad0702ec6cea4de3824ecb465843e4851d73620abe40af
z61b3637cba372e65b8046296da2819417457db8c042b4d8a0be024b09b27558e0394121ebe3989
z2a321c376899d3cecad6ba0a79e5808eae15ef04cd9ae7164444b5fd2bf06c2d19c8804e89a9fe
z85578e5d268904a34f44c1e20d9c48d433d9204a0f906eb93a7cf8b40d3d4229d80d7f92e9f8ca
z0b5f85a5b29c25a99001fd8b1a03fd212681741ed373a9223db6e5ee16557e8d476f71feceaf5a
z6ec2edd19219282a961ed2cb266cd1c61dad7c75740352c4f7e84010357be441b022a63f97d45a
zcb459ed747db89b2905426cdd20fc1e1a0435216f6a63202e412d5fbca1e48364c549df5322be0
z40b189693e49f9db6b2c4fc45b17c2d810edd8ca967f5a3fd9bdc269f078f2e5e2b248ec54c2e4
z0e2d5e22f83430f8115fbe14d99b252bfed06811bd876cfb4f72a56448bd71ade935f99a1a4121
z2dade97ad72973e98d29529273ed72b2ddf1cff736f6c8826469b831ad374493ebd73024726054
ze17d30904135a8afab9df5ebdd69275aa1d75e8cc370b4b8e06b836cf055b5302ab92a3d1dcf72
z45e912ee4013da06ee9ddb1f0dcff4682584435ccb25d381d88c62ba0b4c36b3a18e76d0e6096e
z0caa10b37f49b506f078987a4bddb9446f2829a11c6a97106166e1460e24ad050c297482d43215
zc0e55653421f61e651e17c02c2dfd396b5f1ef2f2386395e7ae56d3d034008418fe4987fcc8909
z9f35ba0b0e63b921d838f5804ad5d8bafc5646606b431ca1379bbfea717f6819b964295c87ff4b
zc19fda8a296f7fc4514079ea81fe77e8717c3441f1cbca55e2618c0e86ee69b8962f5632979025
zb9f6d2cb27d431d67f8e24165f82f9baaeed0779f7097d51de007587c19c73c90b1d9624f52ce9
zbd5f24cb512cf8691e3a3fa98142e7d37f25035e2e4e0f4c7f8f9e2867af1c23419e217b953267
z684e44f057faae71d4d7ac079088e6744d9be114661b924a5ea0c88af262b47c46d8cc3cc12565
za7bb2d5c7b83a3af36c8b2ea06775f16456afb8eaded21eb4abb52291d8ea65ba733397ba05487
zd01d9935c57136abd239241ffb96dffd9aba80bf65cd3ada93bc8eb281c7c7c0102cfcd9f0ea67
zfbbd258f618ae3b6e59681b0138164d92a56bfd076d6edbc55b63e2cd2d999ff44dacae9195669
za9a6d30d510492973fb19a44c313eb4563fc9f1137cc9a5c666029d6121a1e57c8803209a6b47f
z710e0c3812111825e982353c1a3909515616856a646ca9ca253ec8f9ab8bb73454b0565fe97e93
zfa128fc873080af2825a357cf27cea83ba2a0fd399eec6b11bbd18f191836de4b45af778ec07f8
zdadcce377f0f30ed9eff700cdba68a150ba0bb88fecd3d41052b2bb27df7928840612fad56a8bb
z53968cac71223463251bea2bf3980032b220f3cbea3edb3d0843ef957b58d937aa445fbed85c86
ze6be94472691ab0013a870ac3df1007f9243641e69ca5302047fcaefce387de6af44187e3901d7
z583bfee700f42f0385fe7d5e814d3020d2d20d68b87a56479aa165f68b9f8b38b375e8d8cac3cb
zc2802fefbb4271528e50fd5140d8265a086b0972c9dffd10a4fb164c11e57863bfbf37c7ab4442
z1018f6fb3d12ff1702c0f801d3d24502eab538f60bb9da8b19f8dfcf0b13d0ad4e519967dc0104
zf54f9ad8c3e64cd614200aec1d904b37924d0a17d682afe73045a2cb0e340734819c1f0224ab65
zb23543e685b926a20afab41732e3b7be3c7f6c6e7effdc6b44293e5e0cb2ec595677a60956f995
z6863b9fc9b74053d667aea7d824a3cd1f97484835d3aa3e5e7b13fba8d3d8b073e4c2fe5358071
z04532b6a5ff3037bb183b34edc9bf37dea6031627f4962ea1ae97612609693caf9dad3aa1e5ace
za1fe4ef2da2b04227a4ee5c19a7d0212b448f55683be1620a3e3fd3a6c6c4aa13d4fcf9976816c
z8d8159ad179f98155ef393715e82c779c929dfbcfddf7311469210656feec3debc2fcb4749bde7
z017cc4ac701a8c0a62b3badbda6ef075f831d39b17a52c1faefeaaec937b32727e203da125a345
zf636a6b465a42508bdc2e1bf771cb63ff8bf3eb1117117950110670b4f46cf5802527991c18f2e
z1af5951808937bf311be5b088436a6fc476e152af402095c649bf4c5ed6983937d530ae9cb2cf7
zcd513ac2faf48cded5e2deab74ebf6c5a362989738aa2d0392f8ae59fe0206b53d5a17db7813d1
z7625b3693c1a3c490b3a030f7d3087b79f401eeed38a5ab993a76cb6fa94acef48dbb564f9b904
z18a0680183ae01831690a19d3322d33afecf9b01b6289f5d41de2085429f0f3f1703d3e0a27f6a
zdb9522afd60758f270e19b58f4630c2f8370f009aa995c240195d4ecad34532cb1bf79cc0442fa
za868624f8456a27a488b4d6f3ba3c817b49bf4296592921a1f16db9490cab7d9b280bcd7cd5fcf
z50d6d3707b842d8b74781e338cc21c6be815eed10493507553adedd093af287a0b452c431217cd
zb60e986dc7dd769caf9877382e630013db8da442e2276ee7a3442a7676d0ebba4add10ad23f534
za40e7523e82d1d3baaf81e2aed1da0332734ec268f8401dd8394486428a7c1146143129105a49c
z170618b4b683b09e8d859b45bd10cad36c2c5586c90e2fb830ad19f0c5ff4cc322671f1f770f99
z92d9e918279447ab268d4108b2b8ae1400645ae0ef3f9c1ae752540659432f419673dfc9254000
z0f2148b0a90cf25d7d5d72ab9cac9bb59da10895a9313a4fb55089df2ecdad26831bdb3f7cab3c
za1917d991be6e43e2417ad0bd5a2b3aa1c503511d17ba20717b3c0ce75fbab3d684a7bc7acf806
z33edd5c62fafcaa00760c81a53953b957fb1caa973d9cca8d65e46bb8ba5886e020a079f0a7fa0
z7e9a584ad210b9589cc3893ea2bdf6a445127136538bd381548dfb23b3158044e68ed602a815bd
ze78923089d94189e33ecbd53d3c93fa3128606b92f9e9a505a6d918ee9e8b9f415c981d1a8cfe1
ze9779624ffa7a52abc382f7a5b4d78be1e3ec4c20806ab4a02ab0f86cb0607df67592ec8ee2e7c
z47fb6c84915cedf4224a62e16f81d1885cb2d085e7b3a4792ff2262b055849d2c391f1486d5a21
z07b00f8cd7de41ab76b2e7f313774bc9053984336d9b04f6393d6709d7236be28ca60e7f369282
z5a6d9bc6dc7f73505701e4e3014f87fd7a18919dae07a4b7dc65466f5b373cc809e39e70cb7e07
za5624c764b894a9b548fd2fc4f3728997d503595d1b77c35b6d8e31ed00b363925bdaddbecd63c
zf3a046d1435d89065370f1900ac10de49ccc73d57cebbc48435bcc34a86724a98d36b7f68161d7
z2010c70d39903199df96fc1923deb7a0726d8882c2964c45ee55c38b368e5b5f96562cf7d7f644
z7965a1ec218cf6e384d2abc2840b2781ce837f99320fb126ef88fda9b39eb859fd646ded2994ec
z7e79f59385f169c373246bebcf998f98167c270291202971b94768236bea6aaa2e07017dd5b941
zcc97d7242da2d5995dafeedfae1c695b343c0e543d7cd4a6c910c767275b5d29c01a76519e4798
z0f4e7d8dd589d6e25f2a0afc81f1de7b9ff48a3893f477d5e7e54dd15910bc5b134755f5b3a344
zf9085941f19666dd57b9daedda401e78640ea66dbc6dd87d34fb79949a93a41f6502ba0d0803b8
zeb1e698e116fe30afbc6255416332a8792ff4c616006cb9951b8a13c25aa9ae4af31c03d9198f3
z06743cc644db9f7fbac384818ff38cfe0a61415be965161f654aeefac74b16bff76d5a840b9627
z16d15dd015314f4a8fffd1077a467cc7b380e19669d3deb899dbf7a9788783087bd6b7b30b8f0c
zc28655d9a3476be7ac1752c3388edcc3ce9026e4d1504225d4c9d01826bbe436f0927af4a03b8a
z381d5af76064809b08472ca250f6dca1c3e56ae6fe332b229fc1d8d901958c638ec59089e8b538
z936922c6d9bcacb55f840c800563ed55d94c587f9b434d64cf17b639c776fc3b0bb28b9cbe75ac
z2afb1ba5cebebb76a0669229c6026d874df968b4b61192cd674be020af11315c4565b54a5bb0ed
z54b324ad0c5f2fa3078933cc2eccec3c8d4ebe36753774f3aa2822b18d4b28b8e8b359e70fd6a9
zeb230ac72ea9d1b3f98f20ce7318510e785a0f236992375c57dcf7ce1739c14b9e59e1f571c73e
zcc8c5f90a68cdeb82a8aff7912f5f6e58497c9d1d972400eb37f60af67c8b6f4f732912bc3f341
zdadaa67f3b88c817cc4cfa467a772b32ecfae128db2db8bbe28f8879beedc73eff5f667c955f81
z79381887e41bc57dc17c2a91bf62e8055dc307845ca581bdcbb3bf7267fa6088417be55a4527b0
z8cfd681ba4585181c59c2e03688f1785286721e46b4d6c3ab20e5ffa6b3382d23650c14a51fa4d
z95561a9081bd5238724f9b9f102cf709be2084515c4f10bf9d34040e32a205bf045fbe9f05a99b
z917e359b2478c99a2b03dc1d3d83245250f0c020e844e2e7a3b47e4c4ae343246b3b2c855104a6
zd295ec8953c283c54c7c9232920116785d30948bfe445043f7ffa0bd82224c2f5c3be384478857
z61ccc84780e952a9b28ececc59bf8862a07b9ce3c0ace743e3521141f4fe8a09e51cb423a86fd8
z5e791481ac7808b00eee3afaa57eade21d973cb5b6b4a40b07048c44c54c277d3691f7e889320b
z7d7e6ed0265857edd7b3c30e0f7df6e8547c554f3b2caa1114275d64e65cb1812dbf9d29bef46c
z2ac1ba7507d9d37d06522b4a8435598fe5a907978181138a21d1b75d5f0503328720f800f7ea32
z183f982bae5921dae0382157089cbefb0e4a87a755f1ef3434f0f7990729f8af7f64212e1a5e40
z712f598be3ab83eb15ba0715c08d36be90c5fa2c3a12af54be0af9b3935578317ff8b041a91e39
zc1afcf2a2d947a3354c7f37eb8b49cdd9a181d079284b7bbe85638d3aa8020b961072892279a5c
z66ec139be6645e5869ad3caa77cfba2fbe995e0dcf95911e3528b8f09e55a80764540a7347b520
z22b9146bdac50d26d7f03f8fd4ee23b24980f715c160395d47b620660aa5aed0b283fc6c86c68f
z9d477086ba62c24b340af58618d91809e4880bc11eadf0b8615ef5d78fc44a41e4652ae7e5ce25
z533dbd38d2cdde56d46671dac71296b17b8fd5882915a64db8fce1037cb4240cbb8ffee663555a
z53a7f80a657e5267029e05f110cc7fdaf045ac88fb77677d17909034a90f5870aeccfdbf9cf853
z33076a7bfd7add4e7383fe75284e87b181025e894227c091b5ceff60d0ee5c6f6f00171c25c1a3
z47aa579038f31b7a0feac996d7e317c8edc1a80e6fa0792f40b31baf05b9d6fe0985e8dcbeddf5
zc9c64c90c84b3187510f5fa516576e33dd89f35f2b17fc92b14913b35eb3b13e087e7aca8a6a3a
z6154e9120a1539350a3b497eaba5468e85ab89d1ab1a0543f17f9431ed8ae1e667fd7dd0763a44
ze3b6fb5a24ccb4c2b0e047568763d497ddcdd1e161d5492d78b33b7fab0d24a5445dd67310e660
z24c04e9c2277be411b5550fe5e9dfcf55fa2c68aa5518715d41642eda7e59bd6ba9a3b6b9dc05c
z46aad8f5356e8cbb735377c55b8fb74a64e126108299d712ea35f2e52ac73d669d24541d819e67
z04b5c5e8af24648390a98889ff5deca2b35cd21ee0d1d1a054d77d15f4026e1d52a05b4cf84d41
z9fa2a61cb8879d914b1384e33cd0a64da2c914fc77d5e39f81d6c855b26ba8d51b94c5e7490232
z4d034d5270ee4a5f4096fffa6df348072e8f22546f4761209f6bbf50a8531eedbfbf531cd5d782
z4d0b0b3b70e1bc5ba6eb168f1978b01c460d05b7dd25900438f0fbff2fe7aa4fffb2002279b4da
z8506776ccaa30649bb801a2e5f70bfc5474a570e69350377c9148d6d586ab60bfa09cdf4986ea5
z414a3677af9c7e12bfbe6daf9fead0c432c08565869d1dc22e653287404782697adcbab9c40657
zddecd31332cac246250aa4e2ebca0f214be52bca555a40caf5c5464afe4cfbf84846fa26acc319
z84fe4c9bbb4fc368de16124281783c1fe4fa113cfb1b2a2531c7b610b6eff8073dc38becc22be2
z2ad825fe6f6d2b6338eb442f11cb90daa8b2b83039da75974a437a29288d9ece55b2d8d3f6afff
zac3d5f98b3cee01c2b7d233d50bd35ec8ec1e7d5956dd1d3c6ff49892cab368407247b9215486e
zcd01aecc85dcff2fd335f9512c88e71c05cba22e4cc16bc8309f09abeec1a961173ab5a8fcc93c
z92ab9d91087ac6c62af9dfe751ce829f90db6c24093bf1f07c07342050046ae86adb93ef048055
z476b235247e8ae11a5da01c02ad8d282e38cd50371a7965c1b9e46c1d6c78dc377dd49addb8b25
z647213d71d98ddc4f058602baf5f2a75b9036792ac67909238608b58cf2e0f8e351db3daa15450
zff49c02edd4274d311fa1e0a9dd7b82fa9775c083ff868c0bc66b5774106ddb361ae094665bf05
z20185d3ae4deb787dc967ce9fa8f7f6fad36052155f15f8379859db3ef348f5f6b5d1fa6eabde2
z78b5d884fa34abe61daf56ae2dc3352d3fd517319f5623f126b977063a0e4daa3dc59ced9c9956
ze903d232d4f0c0cbe3904a02b550a1e30f645f2bc74a80887a7a2e49ca5e32e46431c461731b43
zbb6774bbe85f443cd90f43f634e18f2f6255a2f68761e68f5e7433fadaf8e37ac8d9efc8032bec
zaead978825259112bb69bf8cdd51157f7c7fc870ce34c972ee252f82aa5ce2fdf59b6f66561ec5
za090e1c5f6a10bb28e387294f2f9a7d9c163bfea319bdf4226089353b35d0a1a19bb995201759e
z0750916b151df4a9e208e006a8dcdcd951cf16d3944c887996fd26d0dcfd6a0d38d6c4c02ddd69
z7fbbf0e4d6fd9edd605a8b5c7efed2f21cb3d04946681c4c343816ccd7c6ad3c1a01c7cc2ceb72
z7612cc02538c49facc8b8d8520838ae026723ff3c2a2362b91936430a5adcff636ec63f19678ee
z62366405f3b094853e8ec198cc67934cd72b27903a09448220c57f5176f60c0390fd723d2f18a4
z6e266df685e2304e78126411154a8d62bc884add4aa94fda60bced239440bffd50d4b33c86918d
z41552ec3465b9f6991e43381ea44300f1ce8c5c27fe16ee174824d6c57de49693df4a430b68ec4
z3e4f43d296b66c4496db0c56b500a16806b22e11db25bc3f5386eaa017389810fbb237e875bcc0
z437cd48f109294f925982e876aece11a9a8a136ee98fae3a8235dfc3eecfccff7cc8c80821c612
zf59b10c4692eea6dd09a5660205274d08fcaaee49abf652088803b4ebab1078af5be1f1a4fa8d0
z714b42c4140cf2abca7ecbf28d28ceba43184a8f1b0c68ed95c30a3966a500588d7529e6fed8e6
zd8ef83ef72e75eb9afcad8d99183bd6392f00d4525a4347a350d3ee4f4d85162beeb14c48de142
z6d3505bffda81b6574412c32fefe3a25d911a3d20ac1db73c97bf7d12ac30227094c7a914f357e
z98f04ff7e4e8a0a6d5bd6b8fb0ee55a224956c3736c8e097a935984b51d68e40c64d04598fc6b9
z4f23c38699185da368e967ee44e6a2c40bc5f3e0427643cc8e4fffbbd9af4115f56dfc7273d579
zf5f13b441ceeeaaac13a390df6e34c1fcb8ea82289d6aeeffc1138be22c2f58d48b2d07eb2787f
z46fdad357f69e74a910a9a00bbdca3e3117a87b3cbc3e18ac5205918579a6423bfe3e2315469b4
zcc89cb3944a2e7f546846743dd46d53526c197dcfca38173ad441e2e1e757a0ba6380031890700
za207328a33c538ef09f179b6518d7797caa45f76f23ce63f6e0daaba0082c6018d280e1ccdaf94
z5dbbd00f753b7903324c6418bc02fdfc41446b1f97019399ca92362c13cb105bccc73ebfe43e08
zf4d3264da5a0463bedcaac2e4e737d79780868dd98d0aa42bff5414447a5b08e97924e6431f52a
z695a48a21095c7f8e8bdc3176b3992dbe4051122a2db52cbce9f5e2bbb6e1cb77b1b627e44abf4
z4c230a0bae0b2375b41368f8a1e355e19876f1e5605527efeafccb41a394d19271a0062cd71ddb
zd0862d26cfcb7223a04c5fb8bd6f0e6dfbbc4caf4bf89fead8d9e8bf1295d8c500883ea849554a
zb5c85d3098a6cca87b94602f27710ed33af729e85547679b05d923d40b79403daf1d674b41ee97
zc6d160392f2ddd1ddf427bf25d2a7be96024cdceb47b1f25cb941ef5443ad28720c5c185c67dac
z6604bb640c8ca186b3a252006b4b3a7f2eff1e6de8329bac410c926a8f160f88cdfffaec101df9
z5a57633a1b21254909be62e4888f49589917276c9c7dba3f13585ef2c6a247a141e50c9f5f8190
z114aa708f66a67bc81a4f695cc30e823f00d1ad1b8a753ea7ff4eed4f7582e6d1230bd080b9f17
z413e7b37a61d3cbf8d7a2ce0fb088cdda84ade0c2047db9659919eb8817bb42f1511b68ee71f5c
z66374f43ad901d27c476c036c94e7866ea878a628d9f2cad431a070f14bc6fe0fc27044c6bb2ee
z87a3f6ca7d62d72a1cf8fe0835e2a296ab1a9c8cdbaf7e0c123d0ae1ca7fa0183a544f50127e7b
z3956c8ed8d54c8a1c651a2c3082fb169e6f51304666c7c6d96c18cc9412f3e2aee400aca1d3fa2
zf8e2dd51d5584fd14c157d04f17de09a6e760315af26f7fd1a77dd3a33a39df0caf9e59d68a0ed
z78c11a93fa1fb60c8ec17663b2c7351d4406a71cadd9b0dcc704968121d3a4a38075ff2b366c76
z5bf439fad3f0375951c08b40de6d00737405fa794b888862fe51697e10bbfb3fe47545d209e534
z1affa0234230d5f1327382b6602ab5b51482d7d4bc1b4ced897ff795d8adae17614956b611303c
zc3101212dfcae21df17e601419890f31c35e531314d35e293cfe98177fa0f79d2f30a286093b58
zb2d0fb2ccc48e9118d2e3b3e0524156cdc1e6b5e00baf5a4767ab8eb99b468dfbaf79ca9bb874e
z4c1f758d66b7f400fb72ac70dbf0e7ecd5f00a42584465b7054cb7c63d533972505593bb371b20
zc02dc88a12a84ad1367e7a3a99d8a44b374e43f5f9173c54d3c854da9dd4f3bd595de2329c01a2
z0de87ec36a7359e27ea95bba3a02d663fe6fbc2629d16e66cc9f7128b87d5bf7622ca75e55bad1
z77843d60abe11e04169d59f179dc638ab2c6733120da420cff474028373f724450fd879b03b3c8
ze821909e43a268c414f9da2bcf5af05827e8a107981b31845139494f6e75be3442b02045a0f70e
zae9030d03f3aa3a94ca7884b9e00847cdad5945e7fd13194db1eea792a11de9b9bbf0ae360080c
z315e2c5f277c45a89c71272d6d079722d5f84f6bbc50fc69a0cfe851d0495d0ce2cf32cfa6ab5d
z7478f41d93b6ce122ee10dc4f4f0eca836495e0ea625898144aef352d0949ff3f610e1c0afd2f5
z53439e68c2d53dc0b8de8283bfe0bdef6e579c0060d08fbc017ffee9feed1e1f79d94a595de7f2
z811a62d2536abdcc5f9d2ccce8a64936fabe38ec656ed2c37b0dba3a101f1d55a6335578b71fc7
zc4e650cc82e834bb2cb319ec0bc7a0e74b2ec87011a123c1015a1350eae34335ab2e727f436e1a
z374ffc09cea3faa418e60b33012d3c95ec2fda91242ffd3c3be3e5e2e30125d4d17b9f83fae7ab
za51538eb333c9f22823d285224172b6ac09e4b1365634cebb64c9f5c3558fb6310657fe672385e
zcbc2b1f3bccb06160865e13783737179df6e58af0f4817e9c2e83e0b0e88e223cc21c2a954f7d8
z8ab33dc00cadc0b13cb923ab89bc58e4f6f258f24fc9b441978e0160f83af08b55409b3e576595
z57aa78d2d3d906c36c20f2a6bd50351865951fd9fe28eb0d44cf3f20a49e7fe95a1735c2c32f1e
z41c87d9dceb2907cd16ed94446f60867eb584648283381a31394d5c58c89c665dad5f846b8f781
zb5b8ce3637bc688e55bc5817c5be724cceaf9a8375eeeb9c0a24d5400e8c3696aef6e0a6f38698
zcad6a7e639d11b0f0c2b51eee43b04a7145aee98aa1127c5138b0e6cd62698a0a4823caba44c07
z3beac4ed6a9f59d3b020e1114dc4537484ded96007c2a2cf34fff11290a7b0e8d3805079e1327a
z8f2e4aa4fa636750ab34e436c734b19495c8bb0c371871fee5ebfbfe641b6c9da6ab59ab1ee80f
z29565d7d56b0e5989766d3b31f0ff6e3c9637eae5bc973b3476eace7a48414e8557ebb353d978a
z13afc818c1fe84b90cc5d99e030d77441adffb0870ed6a652415394cf73e1f5d9f47a7853d7f64
z6e13b79247623b15ef5c54cae8ccbcfd08373bc35f1f3bdb0b75e65c801145284e740ed0d91069
zae7781879a4996af6c89537828b8009377acea8abfff29c888d99bd186e6f1af054aa0653e6451
z5aaa459ee53788d7fe14e4c340134cad826cd64c9b12b72cbbce1d32c42f7083c8fa17b17c7fda
zfde33b214e90311e59364ea7813de85dc015eca57dd5dd694f23d07d37c5fef7b4a8797cbf4ed2
zf29b8fd64d94bda4bf9c810751a91ae21ff00ba8e6fe7d0e64aee18d774f53cc7c64e573a9f09b
zb92839b91889c4644836b776b28c34fe46439dd2ffe9bfd6bec8e970515f6cf21b314acd04f217
z6f3ecf4587e4e39d6082bd80e6fed11b458905ed9e2b2de7eb3e854bbf17c8895dac0fe16d633f
z58f71d760da9ac2fba85a6789a55b7e78156e12ef29ee419af847e5dff9d578564b34f3e93caf4
z032f1e98372b63ed0ab6007133c9addde0d7b7876a6dd67b69fa8ed7057f21865756f6cab9b78b
z33c14b5c2d3cbb8a74e86555659c01794217b5b4ae845757c79048beba93ae10f0c0f57b921721
zdbe94dd22b291167ba89425452de91c6c2d8718de2c527e0eaff6639151e05fe918e9e89337485
zeeb26450de26b4170c59de3220917d71705659963a01cd3e3840f4998e5bba0e188950a4706770
z0995c5e6fa31de24f94c6371d3e2ea3f0a3be8bb08e5854db281fa2a9b76cc2b816fe9fb990d81
z30d7f955bcccc7e9fc4b45ef8a72931b1c336b6469040893fa69053cac8c227e621606d00e61c6
z9f2ba106ba4aca35b1c7ae3dd8728d02a88a6bb08c0626521c63d4c60cbc5a8f6cf215faeb1374
ze484b2e3d404b3414ebd1d78278555743453b8ee90d4850c333ae3ed8116e7ce60c3c79de15aa5
z81b50197b16c16598d86374ef51fd91604f759d13a22396cd30cd34eb515445bcd9b3a41e9e0ba
z962c4d1d5d6ccaa1d197347d769b9ba18e43f377c16ed1cd6793f922b2c84e23f23a6262c4e17d
ze33ca68999fbc88c2e61a9c8e2febfbbceacb95aed5557ab107a99534c538132c0bdcd65546182
z7bb647e67caeb33c922120f321884cb76af89bbfac9eb58406781cc4e3b98f594ff0117a0c1dbe
zb403674de52b7d5f02dfcc5ed2fcb98c8f9c59cefc5cfe93605fba9a67ead8d822dc25719eb144
z5db547e6b2157cd02d8fd8e4e1fbc15d00dfe00232ada95e64b6106c7c740b33a9b1112e0f9269
z6a0fd50bfcd52176de6231e0450439cc0a3256e352b1186efe59da2ae212c9dc80483f736c9c87
zb86b09ccc64da049c7ffd0388f3d30ad41ca6ad6d246e74952fc78aadbc320b4125bdf9ede6acd
z6ac6b5adc2c445351d34cb5f305dd5ad52108349127d6dc88588a7125d27075a4cc2d5b068f7a7
z82fae4f6b99ef77ed77e330c2b72a8ccfebce9e0d96530daae06913b22091d536e189aaf3d332c
zda64d5f07f089979c1a5e45f1a103ae7722b75f150eb0297f4033d082e42ea6f9b78f17267ac6f
z22cb93fec2013b0e2f5be3ec0c5c92e0dcfaf648ec0fe0b8760b7060e25213569ed93f241d01fc
zdd6d94bfe7c1ed5cc40d023679bd2ae139d3b0fd3310060cf63aac7b7d4267a31dd074deead4f3
zc98091310be05653a73d846c8ed6f5ca62694015da1e2096294cdb389a06a570dfdaae4245e37f
z10630bc0f1af73d0314764059d802fb989465bd8ab5d4c1a67328d38d244cc446d0206c6a0ffd6
z763a37429bba9ab0ddb9be75ca3bb7f25b80f29affbe3dd8f75d99c106a40c505a2600021f8432
z3b0aad10c2e3e3ab267be813a5116e560a8a0cbdb3757b4f061213c35e6a2bb61b653d9a9f7ed6
z4d7afdc126c3da7bff737e050f08aa501fcba24825fa6f7058df60d119b42f83ef3dab10dd2613
z5d2baade6f2435f28b140d64def06687782d1a965ac2e7e6592c17ee05d22fdfc86df141755341
z1464e5b409d5601c5b5ede0ebcae3bc999564b057133a23270c8acd3ea960cecd6bffa5ea3daad
z12fb91511e12d173cc0b74014fe8e11e469ca0584f0eea789d65ab160c171473bf0ab6a5161cc7
z51ea1a74f75438f563f51768ad05c7aba3747c288fa550ac75389510c15a6d5a624c3337c2c5f6
zc8cc0627d4c48795c7668025b4fffb6c3ffe72322239fc03e3f1182f19c7dba40bdd7fc7883fe7
zefad63133872e05c49d1a3bcd3bd191d21208d47da9855cde0bb80545fff7c7cbf3809489d7da5
zc84b0e1ec9642f2dfd2dd29dcc360210f9bd9c7cca8a90b33e8a8efb5a8a20deacf0f7406cc8ac
z5a60b665585b100b8d01e0360b789de21ac4e6cbaeb7976fb4d9944e349841d92bc826d6d78e9b
z84f66aa85010ea02d95fa501fc97ce51f235225928b369bea7017da38135950d64f4422d45560b
zd81af676e5922256439770ac72faa84f7f47d5c32fe858f699a5b0fb5d2813cfc5fff733340279
z5436253dee71e6d6329bfdee26ff53434e30a40f2aad019f25e03796a3e608cd7b0373ebd5cd6b
z9ef126f8fc134476e68f405bca0e1b2e5f0df3fb8b0c961e7e92db2e23f75b6768063ddf1c3cb9
z294ef44b07cb715db762ff226b42e21efc47ded323350a509b4b5ffb0b16f94c93fbcaddb0b4d5
z60c6ad9008d7a64f637ccfaa50b6ebdefa716eea23b9239441f28236d885740881bce3a486af60
ze7b7c6b21ad83fd884716081b2395ee30f5016fa6313cc7b93e43fad46727a86a419ff5af35083
z57d1b04a289533ae1e32e30246d4510b8913bc5fc093f33c2b13c96b46b5d1882badd0e979e777
zf3ecce4238abff76a88826fafcda82cf09bea958b25f9b0eee650718d220f1d09554fa8a9a09af
z90cb5ea357cb44a470543ca6bf7eee7440e1df30b81b9c5d050ff0c6ddb324ebf457e3a1d238e9
zd0801529c60e8b123a768d0ecbe1193dd626c4ca06a23468f6e3a6d3a14a52c71edfe2e8b4da9a
z7d77400a3439ab212e9588ad2dc9a2658339724fc7aeb0e13411cc4237e18159e75823205d99fd
z7d3fa3fe48c34a727cf3ee6859b4ecfdb793fe75c4a39aac8420326e1248ebcdbbbbdfe0e23c2f
z19285a425bf2b24b6257f1e2132b5229fb2b1adce34e6d76b242f78a706e4d9f232fd228caf356
z5dcc9229222ea3d231398584182d2f9345d4d8756f4b74aa5cd4be44917b627ce6ba0babcc7132
zb8b70198063639b955d4ee2d6582a47925b1abc2e3040f1ec5433098df8dc4b3a79a6f694c6e28
z46fa6acadd7652c8c0d6cf90ab1587e1f04b3f9a977ddb548e2cf25c1693d27f9e80975c8c98fa
z3e6188b899fa572d5835e2f8216df3f9e2376da0d3eed533d885e4aa10e3cdb2b22b156cb5f8bb
zd806557cfdd65d49d4538792d3774b350b8d5d5ade4291317b739b09de2df420b49354e99c06b4
zd1f921b0a0950c6812e6034cf28380dc0267571274fc56c8406c7b0d1ac50bb4f63fe323d0e521
z34f5299cfb5b8207866e766fa65ce4a27bae9330b7937ea7d5cbd81144e867cba40e166ecb9740
zeaf545c9ef06385b79d69ea5eb7855e2b78160ce3eedd8e41f49a393d0b17382debcb6ff61d45f
z12d1a063991f593948c32db15d64156dfd193cb46f536e52f268120052b26a646b1d53d0ad6341
z0073388b1345a96d3643523f339299c0273cb9571ae71901a3a5d93841a1e77803469f7a7ebe28
ze13c52b2bc9e3bad3d022b4e3594273eb285d100bd37e1383557de7871a9f558ecbde9ebad8925
z4bf13c26df1accb15200cad5999359ab60b6a7ad85b853f3106545cdbd2c8f199f9e29f7b44dfe
z94c94ac4c9b2ea9ea40c3045e2fc604391b91a4a1755aebd6a0ac34a247aa7f4ed8fc3fa114efe
z93dcec6eba4a6b7e95bada1b395b86d8745c6e80fbc0787e7808a978df089a92a185dad994bbbd
zdc24b94c7e5ee49c78c7b12545a4624b9d6101f72d5a8ada76a7a58d5e3e31de1d405fc408e9b3
z7a992cd46ca5dade527a13ee08443d7209c41844c5fa83195d86ad4b93a35c95f5deb6b9b25554
z8aee3e772c5f3768f9b7a4da207f25b663bbe3da827617f5859b6502b94400c0906c0f30107d1f
z2360ab4855d4100e40d932fc4cf4ec0275f228c577adf5f834bc6d4e1e69f775e2fd4e7cb70105
z34d2f9344c311d8cde8e251f4fa6f690b563a8511fa7f425bed138298bd11378288bc47fbb4553
z1ad242ff29777531498db9aa23706fefc03ba6395862f3a84b4c005dd78ab46aed336cfd71cedb
zfd97d3238c109af0d465a77e3557827a611dbb6483a05588aad8277264a56fb3f38a81c7af89b7
z6e23bdfe4b0bb717e8435b2781bc8a6630e336fb561562481fddee0604a650b8c388db28795ea2
ze2fd8f9f67079c98b6bde2d8ea45ff0feac013c3c2f6878e66a6dd546fc7465bc7cc77a9974a1a
zb1c5fd42cd4eebb669caa6391a53d68d7602cc17e35194c09fa6f4369c1aa084f90054fb2ef1a0
z49824732ead16f3a1be5c1d89170d8047a65b2c8a255330ea1ee86aa7b9e250c73f7ee0110ede6
z629567f957a037f37d12622c8faa432ec71723496703276b7d7fb2e5effcb13c9f39462890d31e
z83287672a79a4b5fc84d9b122314b95ace9038e8c5aa92ee9be02512ddde7cb16cf37ee72e3cb5
z5ba1259040f414743569bde8e17c6d67359472a59227a99e2ba5c7303519d9e4aa2ed01d59e10c
z0d452ad5d749a7a1b18676d694027a87d018c09c34e0f3438a285bfeb7c20721478754b04f6932
z80ab8dea666e38c7bef7fb20cfc8b3fdbe2c2a2dccfb1ef11ad8aa3cf14e7a0489c9347de559ca
z517537b6e54f5c622b2df6148c990d3aec0545dc434fbf62e10fd048597c9875634a78a4061878
z215a0d6405cece5039378efd0ad1f97d06be5e230736bb5cc00a8a739d55abf8cb7a9bec39ff98
zc582106edcdc5e636b578fcdf3b67c34062880be2c3294ddbcc7893d969c340f5fa13545a2de5d
z7efae6bbe029369e174eec0dcd6acb51da8a9daafe16da9a873200591fc01cafd8aac8524e9978
z3a4b39507bf8a46144486c529e53c539a1119e426177a66e44af5e2f4552b31bbb3f1f9fde6144
zd0061c528e7ccce73033434da06a4181abb66cc261ae0b782aef845b88e7fa740c6b8141714b45
zb6eb665e6c4115fa3fc6e9c5014053cf0928846d0282e45f8afbd61ac9c6e17f022583a48eca2b
ze6cbf59dc59be595fd06cd2d65923fba82b02bbdddfd7f2c172e42fbf9cb2670e5902113e4f335
z4743e30de4dd66f9fa78490bd953c17343f7b6ab21b70cf2b17926a07e08b699ebc0aaee05b6b5
zfe782480f37acc4151e5c0c18f0fde9bd34f44bb363d71e5fcefdd9ec3fc5ab67bda4ab96d435d
z159763c970270ed72a638a8981b03f6215cebb647cb354de75c65209463e28f656c49377d11321
z067b415d78ae4dffcebb9fd0fdf55c5ac9a6d6fcec21e5f03209b3c3d6522e25325dfc14d6f72b
z53d85f121d228b4e7faed5399ad0ffea9caec6ad2230e7ecfb20c17553623a0046ace9088d93de
z940e4dcca3d5cf67f70d0b2da46c7285f260047a47793c2190dcc55c53c2e9f16af635bcd3a7da
z708b6b4929fc1ae104ba6804661f64ecd203eb67b4a5b802d3de1008e1e1575038df709a6ac692
z0848f1a3a4f6cc9d2f9cdd22b496e732410aaf0e91c1ad814534ecaf86105509ac3dabfec31df1
zbc4c1c7376ff809dd04381f6666aa1e36b7d322cb169991b1340c6be75c350dbc3b578340b4dd2
zabd8071247359a6cda4d2eeb54ad85158f54039d3d5aa26b31ee0cb1a8d9b533398c3f951865ed
z802040371c87268b7917bf2d028901f2652d4fc61f9ee5bed1a5c5255655325e1934562f173573
z1e39ae15740c671a422b34879067a75d4e4254c9cc6d2e432863b50d683dea4b6c80d648046398
z67140045a0eeec6696376f736bb65e5c55ad49533b564f738b94e97031f32a497bd0f52a67a919
z1745cadc1a5f38283d771be122212a489ac6217fc404f24183ace9ec0cf38fa50c4f98cf8a1722
za1471874d8658a6de52c196b27c81fdbe0f747ad7e472b5a47ae54a0578ff349b3c34552cb10de
z0df60320f68f5d281de973b27c0ed3796a220f366443b8506b4fa5b4b584bdbcbd46c362ce517a
ze724480cd32645cafcb88171a7b341473e013fad4f0dcea4da13c2bd2e3482a46d62abda160f50
zef85646c322d0f10127d6d6cf2026c4469b7b367dd9d29f6b2954146532f8b7a0c02bac1788e90
z727be9b6f8cae1ada989c4fc9a4939cb31e22f80566c4a8a003f651e8d3f0065b330e7b6f32d93
zd272d1581a165815c8af975f66365a5b3e0718b3665e15fb48dec6a8256b3d74f0bf5f3f86fce2
zd616dfd6d7d60af28ad381a0804b418945e2480fae0443444c5344818f6cfb035a015d25ff0cc3
z21eec8e9846192701b9097e624c5cf37bbab2140787601b1c9e7c246edd0ded45a572d47c81bcb
z98420ec9479f546560d01cd2373e2eff6d2c3b0a2b87cb0087ae03c88155ee8709d96e636421b9
zd1954ef17c5840f2022fa1e5d0cca278f84ad52d3c5a57139d3041f5055fff3fe32c0e7f7e948f
z3a01c81c3ec99d63cc12efa6aa839e7ebe5063e1180894f0e0c7dea37ff61b157fa0a59de72338
z7f9645cbafc5abef2b24357794b90d7b35a4e2356f4779bd38abb6ed9464c92ad724ac348426d7
z13254836893142926375fa4bf3843c9a7853510cd44390f0b91f86204caabbcf2b2b57e3945e5d
zbc6806f25445449040d77a5ed73de739607164ffa947b5a08105ba303dd7075381b4ce010e7aa8
z0957ddda38d6e25c1c830b393ac81db1bf10397bb3ed02406c6a056c0088a26a4d505c77beec97
z8de331432d4569fe6cefaf78d472734733d048da7c7f3dc10f5e1ec591c418c5d433ced590e9ed
z65aa4e238de432bb419493b7260830f6d435278d83454a26ba6942db568fef2d4e814cb5b9a0a7
zb75ce5b67db306620afcb2ca7602ab4d15d6f68dd2ada698883f4a60b742301082027377b038f9
z3d469654e260b48abf00666eeebbb3e327fc825c09d3308131ae90f9595f4de293ab75296bf3e3
zd9e4d7dfa757894db971a442927f045422612ae7f3b201e305c99b80578980657096ab8c970949
z7a36a09319833a2a350cc852c834520bf3be0b69871ef056fc17956720fda4248b78cd5a219211
z9cdd87c96165d1285c717a572f4fb59557105043ac7925ab3b925e4a4d21188569277a8ccd0cb4
zd4498461555719b3dcd17f9fb07093aebae84ef33fde4578b340db335db8ac9d33cfa6b00f534a
z32e9fa3cb673e0cefe1bce8e5b2cb5e9b60d63372ea6f0feb91bb45759e25f162b618324f046bd
zeca5c3f361107555f5928cb79cc0479952b125babdceb7d851a7bf3f7fd21a895d1b66c336790a
zf0dd0832584d6c105414df5b3b46a4aec9f108df46ea37b785ab1c244b9daded5038faa378577e
zccb71ab633f9259220e0beca58241f6a921cb951a288e37631bff8958b6465deb582ae6eeea14a
zca22ce01ae9c88cf5e948b3f50c20d553add59e76ea7095bc45bfd5946349d5e193f5a08babcb2
z7f276abb4d56c8844800036da72f9c304680fa93d3613ac0188175cd18075bca1c5698559607ce
z5ed2203a93d0d120d70e61dc7944fd091629c8164a7df62eaa50b2abb0cd33bcd78ad4c22f26ac
z0850e17f71921dd64bfd9ac7c44807a81b01170209bf72836eeeefe04a63a18729820bd0f7e79b
z62b99c6140c85df60f877ab90a3602a060e0bb629f15b98944b2c9b7c70d8287933ff801bf2d6b
z01e1524f392e04c23cf6ec30cce9075641cbe7011e1e63a4905709a3313c043c44bc7789bfa367
zc2324696ae2e608aaaed9a94af66d76b07a0f69720d45d27cc97247992f0345f09b2ae978691b4
z211d9576150775e798c22024c91a7ff69c5cb8d3d1c7a002fb6d801d92761259992f617b3c4dd5
z582da38370580ca2959116656d698a6ea299d7c72ab1276030b055ab752177f63aa2547effcbb6
z247dac0612d45ee7c8688c9a21560d2e0fb9bfc3cd317b314bf841320fac41ce9e2f699c8cff77
z09ee28991e9f04ddb7bc0af298a2f4a93b01a94614109c9951233dea0c37fb6d6bebbf7407b78f
zab3f82ffbe3f35e287f91135acaacb4ffabd1f1f6eafff6a3b0ad309c4bc2408ed7167dad6dfaf
zcd3594aef2786c6db5f5a559a91b56f44ea012c411b27583d48aa8e60501ab56cf9b61b6b052d1
z7c33e5f763e92e9cc358ed79828169e0da72cebdd9b77cf904b31880caf758579ba07b66ee07d2
z13f37e247287cc1de2ce6ff5f6090adab323de4a22ff591bc9ff2b2a7abe74a36733ddef19672f
zfdbb86d022b084a60b4a5c75584a0e634b0990394267f0cdd005160818ddea337aee391ae53cb1
z751562384baf0853be5737948ee49f81ceb1741266e27054afd8acd0eff287204a08e8047fffd7
za9a2b02b28927a4973d06964060b8e69971e6f2aa2d8c61325e5680c1f4af64fb2c13b754ee78e
z5f374d193afb0b1668c9e3091bd1831405d2a9c2d65f2dfa7c797bc31f4088520f334197042a94
z984d35d056b3d7f83ff2c10282b71e6a9446e5a993f20b64fe8913743242d018f3241f202714d7
za6eb9536c4733e31545a26c26f0535eb82a2fb37f91ed137f55359317595ed2115326c815f1c8a
z74f244862969ed25c78c7f54e8bdf2ea2d5654b783d527618824c14c64a9de07d3b40fa2cefe57
zfb828fb6517cf86ec6c0930d14da1a70445f2c1a8e10f901b9b13329138389094f552de18c051c
z25e91a00d6000b99c5d35a6597afc0b161bba2aaa8688d3130717c093a911bfb1bb096277c9bf5
zcb9b16a2a31be1d5a254b4fae21b2eed74d4669e6f17c33add46e4a11fdfc5e235c1bd502dec94
z73649ad0d58b412cddcbf45814680c695b56efad18a9fac9b4cbbfe90b56d204ff6012240d76e0
z6a5792b33af95b0decb8567dcbfb2ff482b9fceaa86939199b1d5b07007b9cdf455fc9f483d743
zbadbc13c43988febb267c892f7ccf857e5c01c902a2bdb87f81c27379814a287dd9ec4b2fb6b63
z5a897a7cc3bc47d6e65496098135bcba761096aea6cda3a005c01dcc3cf5444a5348fa74d728aa
z46cf63b87f9633f7a9ff9b0ab7164411c1903c4c730cd36945f33533a188692f9841b2fc7ea489
z79c1abe93fddc74af2a16b9a6906b271f7a7f4c471c90418b801df81d1b7b5a7f01985b930909b
zfcfc1baf216e7559ddfbe4586f715e87fb3daefde65d11726e05bcc99660ee1b4847e451c32748
z2dc85718719cc283a1085083b8bd950698a674e52b26aa90337d77eece91a1cd2723f1549a6ee1
z0b98bbbece9839d17e067dc24424de6f0be749890e4b5dd701e301b02847ca6687822be91f1f66
zb8872a75b5c3b5d981eff7c0cad6a408c13046bcd75d09ef9c01475f4db839e45b175865b4ffb6
zc2a97da73acc9b8e0452cf86eccf38dc365ca3658b8f99c4fc7c0e0c6479b69a3c1b01d9d55d79
zd100b5bc04d5fc3eab555ee75d2a0f25182a4ff9ab7123193a2846ff5bf2a0ae649928aa5149d5
z16cbe97023881343f98715c2f6488c11ca665abf5eba160909538ac2c076db251287ee6102503b
z24d9a87c743d35ee6c30f906ecd36f078192e29666d46852f78e140f58566a161a9d04fd2a19b5
zae9ee0333415b7a68c7590f3ca67ddf52c17a84050abbb29add980ce8a94836c94b6ea35df444e
z58e474629d748e7919cb8a97070ab13c7c7763519fd02163f2cedd38a296a075441c5d1d694188
z4fa6021d714988d77df96baac46639e75783169f2ab2237b0f8d01aef8ed3fce1c5f7a373754e7
ze94ef90850e2dda9268bf9a3a956a01e0c5069fbb600cf8e5cd18c1b02516bbac752840e444275
z2bc69a35260ec85cfe4cc0e67942cf08d8084c2125cb5708430cb13d352b91d8e82009490a5d3e
z5b5c6b5ad230cb7facac4523e2d87e0e869a1ae2755dc0b4d2b26e495aa6b476d9ebe80f7213ac
z555313616124ea1326817fd974fc2b071940253ebcefee61545066d396da79d88237f26a830b1d
z11d0be4c557965b86755cecb17e265288abae0d8d665206406bef01c8c65bc41c4304137552444
z5a36a87adde3d16d1ffb5fdefbacc4d4168e857536bafc10b44ebe8484a9c845e0852c0a8313e7
z8d186795e50fbd2be33c2ce73729f4d12a0c3fbe8e291c3915193b8336f4536a1dd7197e5a1c21
zbec9012848a190b3e07266f7ac8150abc5a8eb9d00e42c638ebebb4e174a7637b7022f1ad5bfb6
z186066e4dda833601ca0ad393fabd000d0c54cc34be5c3292b84b57e9bfc17e517542cf9ca11a7
z8e7b66d46679320ad5858e9f143470839a0b5b11f73915f650da715e2ee4e3eb65b5ada3d24912
z386408016fea2827e57c55703f87b5c69c6a9fe321edda1697731219d39de36ca11bb16f5752fd
z016f7e90b0ca90816e838d2e4825badbed4295c9934acfec8f7a583b71a9cf51f8ef381f760d6d
z6ea5c68a9d4aa9acf1c4fbaa7fc55e4b400a8ca1313f25c55d704368ad0e2959fd395e5b278f8e
z78b9f78d591494257fa974741fb9fcbfb7c0551f44d532bd2ea93d0aef72308f8b9e9f2757ef04
z4236f1da65fe2f4c0d6817985590abd4155c378e65324e8609866d4301f24d7dd44449ebefe389
z9657fa1e732f362ae84c6bc86561536fd60879edf42227ca733ee6bfda406a0cf30341f09240d0
ze90ab3121b71d2b697cc6c15aab407fdf8828a422bb49c6717acde1ca3476c9c27a94d105cf8c1
z5e6de1572d82f5642c1032e217ae0ada45e350191f222e3ef3f4ad0193dc565cff396e3993de73
z0f96f806b33143786020b51d64341db2982ad948e41f6111b7d4d3c150f4c1c2260af84b557dd4
z34dc474779a3698acaa57484c82561dd064f390f184f8af9995bddca924d05ac76e47a48bffc56
z6b79168618e03c40f6c9c30c676f52db88553a3b958a405eaa1386985bbd6f3f06a9461ee42527
z54af00a56a906d2e8a78ba4485e9e139ccbe4128530cc494aa45b302765ab67318ff703b5de26d
zc6d02e8b3695b6332413d79b2b2bafdae606d0407ea13fa1a8a34485630d35d2f767848db7ab98
z1c5a173829c085b8b942f787fde3846c2bf3018583850c1202857a020dbee923571b5cd343a4f0
z8746d4411152dd63df888dbd26d83dbaecc2bdd808d3178ba97e27bf4a21fd98a4d1e51cecb29f
z83cb477156dbf59b52f9e6285b593c18f065475d3422a7c07383f5b0ee952ff0b816dfafde1067
z9b1783f3a0e6442852aa63eee4968118141bec28e3cf945cc7328468d18953a7e7f898237ed3f3
z52c8cfdaa148a825f9a44becbc2a4a2f529ffad772dc5c14eda348f545a946481e21995b2300e6
zcae3f6f483cd85c196294c57009d5db2b555ba0d7c536b36399d07772fb6b47d7c5e668ad9be5a
z454d839151e0de5a3506e0e73215494541a9155060801b456e6a16a32fbcf517a1efc5c12718a6
z46fce4e34b32967dd528b0b42050f59b5ed915c3f33ba50b1bd376a1b29eec747e26e375cd85d5
z263c29083ef44eb840beeaa1a988f9500a867ae572d1955c213623e66bcbed587ebf05a08b6c0d
z3a83219e72c0191f96cde93e82d3dd0de995271674f8d8402ef82c61894ad97ddf51ec8c5d894c
z7205b47e9c84e10af6c055eceaa6abf1182401c9e468ab671e4eb3c07236c0b952ba534faba178
ze4ef91613a0d24a7a0964caa5d5271f00eb266879130044e429af99c08142832261dd14e3da655
zbaea607d2153d8f184772ac3a864a2a0cfac7fdfc744249761e1b2e685a82734c81f73b5d0408a
z167a8b7556cc05676486c021d24884df622ca3ffbdb35dcb52ec0a31fb4d19a208665e6207043b
zfeca2e7171c5d502d8ace5faa02631bfa63ba7c174dc370bcc5795458e22e6d831d48d037487cd
z379d1d03c821f383b52be31d3a0152eefd67b86224bf8e3ca60f7af2e6f05f53d7421baadbe848
ze30bc6f2ee665dc118e1a01393ed3cd32f2f355abf812e287baa9611282fbb51c0e6c9e041a5f0
zc9a61976d42570189ebcfdf759df74a36b68aa6fc0cc0256b0e85ddf92ffa6dc49a02c4d9a6d60
z12234a8b3387c3dba54fe12943b885234a0bc22601f2db94a106b582860fb711cf474d18313301
z951b29f3c2b8f4e2b060fd26b03ab0a080060baa6923c6f176032c5316fadbee1a925bdd759de6
zc88727f7ca826b7a71f1c62635508d5f1ae67f9d16fc3f5d96ac12c1b73265854b9688d660ccda
z96d407bdd97167ed6519c59243446ce70b593910e7702a4d975fe5928c9045d43e2ca83d35d249
zdb4d6dd30333eefccef8807b76cf5b160c5075ffde403b22e73bbf0bba515ce9196ecef6ea345c
z36f25b5d48d6041594521c5d2922bb1e9e14536104080dc2b9a730e1caa1fe0c431b3becf4aae8
z5d0e0a25e6098276b7690c74d2d81f702e800dc574be9bf28c5d971222f19c2aa12f7c638f9ef9
zde2287cdb330bdd37210350f54475cc9e21bec8a51f5760e61de21f25f2a0dd4b4e7ef6b50ca86
zad9243b86b53470c49d376c12195aecd3ab3a489fff0cf04d4d01cb231cf7bb890455da57bb442
z9c9ed18a806bc74e09368566f7891ff2e4f757f3096327aa71a1022c413fb7f2ee0fb22c5f9ed8
zf3a8183df979e61051ab63bc7a1a845c8a48061fb82daa787ba9718a504573e5236897e0783816
zf133322c58d11adfcd52cafe24e9a405647e9c01da408fcbb6caa743b019b77f3d184fe64876b3
zbd8450b9d2b8ea82eddb22e45d4718b8ea7e2898e92d44214f184801c7d403da1087f60fb65cc4
zde73f9d1a324cdcbdd9a490f7c86dc5f02f70f8b1407376c0b2f4568952d7ba20385cee898c064
z41dd534245628682765a9862c241e36bfeb163c15c4be5cdd4343789553d93e11146c6b0e3634d
z4fd21affa956426aac6145acc04df636698be5e85055872fce4ee6be66cdb017aa1d2351856443
z12b0d2eb7273bfb5f59c2d9874a69e3daa108e07e3c817fad8c5ff637b9eeb368da502e58ebc34
z79d9a5b25d65ff9a049cfe32a5566eda671da231c4a3ef9ff6f8ef00c426552e036d5e8bb27ccf
zc77485dfd0ad7c095b6f68d6380439398aa1f440e9ec83a3e42820ce04224176a094ca4d655320
zb0d4bad678304f2119edf04eb816bd342174d605950e24592e37bc73cca81d60b04b5381e3556b
zcca6e805151f9cc730114c1c440a088cee872f50772cf8db14ff959d46171616692cedc96d7e9b
z6352d9e9acc416b0390a82284dfbc9a3831e645caaac22c3297ac923c78c0c2d3ac337c520793f
z875f5c6547fd1611d5f77248bf835fa2462f279647814f1042e350c3e5331ddc1bfee63dc25de0
zaacba1cf74fc4962b859a946f163b2206b0337dbfff79c7408b13b05c8289705bd2d27cc828b58
z6fbe43db4da8f314f708ee5115f1f2cd3becf8cd844db3f2957eb462b68a2ff2f90605b0a9073b
z24b9b831bf819cefe6f135aa7cc330a22943d7c3c076bd998ec17b943f3c9996d94705fd1e6a7b
zc2ebcf011cdd6cb4edd8253e097385b31e58befaa24e06b0cc380cfc1d7ac024ce91ed678e165e
zcdbe8210852786937ffbe8a339be7a6f5048cbcf8a4c619e79711a1a04881fd2c362def3a3a456
z9090dffdc7c28df1912aae6d7e250bdccab9e01d2915ad5c853c58a58cfb444492081013cdccfa
za40a6ca7631616b04fc4b2d01aa374532f4dc3063d2389bbf79826f476b477ca350ff21c612a26
z9f447661f806a5e583a097e9027ba38add4fc651c3c8f909209fd7a60234cb2c45a060983c26d1
z79e93dc4fd5ba7025d5ed596e5b241b6b69f16a558878125f799bff18bcdabe84394af4bd49595
z5a2ef5f967b27a96961bc6216913e7b5301cc5035fc9387eb7e56d427a2048a2ef1f99e558482d
zb6b400aef98cc9d80afbf9c439efce8f42de3482d7974ecb16e9adec14f4a83d92382b04b0f86c
z4d82ba66c0f81c9dce6bdb2da29971c803bd86d17409c831c4fa3d6c3eb65b60013bf5cc25ad4f
z675ae19d6e478154eb73fd8d38a5db05872c91764bab0d520214e246f22fec661e1c36400538a6
z98fe3e0c3cdc78434528e3def6a87a5122885d7ada50067dd2fbb04c838b6af750bff3ca10e657
zea0b1d4eb7a87e775ab871d13d250c052752dfedc749bbfdc10325e8f6226d0e12007969a05098
zba6fbe2deeb3c8943715c20757666c969bc874ca38f07ea0b0be8cae3afc6a1fef421aef926832
z37119e6779aeec5e840053c012a3b127b7bc94bfeb20e57a9980c958f1b02c9ea126d20e9ca8dc
z6a760e18c87cef7a73a5f4508cc13b3db1c05f1af8ef986d0f18c4415a75dd34abaac1c977855b
z2490da7e4b93f9f9f041671feba1012335dcd62dee83aa92229527cb6265f40e5f5c0da9dd38a7
z4362ba282c4c3be19546453f0a6c78d1d21232416676b68fc5e16d47fca8d57fcb58253cdf2133
ze9db9a24f878017bd4de0abdf7eaaac4303519d0c8d02aff8d6563e75a0ef04ab6d77862ee8d73
z5a3d9f0fb373620cb053efcbf8910635a6691fe24a3013b7ee9308cd2a8bbbc37f9a95a5066303
zf00d3b9bbde148218fcf6bbccf2032078de4c4a452b1f9efe507ce8a8c93bb6963a6c7ba76a7c1
zc07b047d98a76a0e5a46e2024bc15640318bb481b23c570ede8827139381c13964c2f138155b9f
za63cd193d00582f283cb3452f5f8088438f9389cf26b7016cc4a25b8415a8a17c1b1822594e521
z62cd9532f05b37e8a6072ee04fc207cc35f6e66a6550cbc92485dbdb121aeb06ece96e26be63dc
z9e429738cbeb951a42296d021847128914e2876d6d0a05255cea2e4c78b4f838876aa952f90e3c
z2a932ea78d3c624f5bbfd53a9de2480e135c52d1b5ad5a39fba97e9450a4a7d304f73e62f44fa4
z271ce1a79a9026e24d5346dccc41d3fb8a030061b8d903f94694f447614c0d2cc27c73a799b71d
zde3f1977c77e8579948319e52ecd95daf2a629676eef0fe40590e6b209c5c617927d0e46abf9a4
z17605aedcf0ca03754ce99d6d59ae0aa9e79b888a0b5c953b566d4ec39ba77af67cf1f68bb5a91
z9c13eecbaca81d58f65fec54d7bb8aecbfbaea3dc7cd8ef6b06b3669e1484badb75ab979ed20ed
z056b39ddd4fd55c288cd7894f93df48868adcd0991d3f798783560e944d28286bafc97198b54d9
z9326543f60f3a857d626d16b738a829912d5e50f7b804fb64c2e359ea18cc09d8b9b1da070f706
ze0d39e9071b3f3792681c0c9fc101ea2e5f6681a80089ee784f95d3ff52f0d8888a015614bfcb8
z8248a126d7ca8a641bd02dd7af10fba67e9d24bc50c83490f5295a25dbafaa743001658db53250
z82ecd2439787381f5f3311d7c9b01f8c5b04ebb8f3f20a581b9e82f96391dc2221a0ce16a93b19
z28db7796243ecf8d3b5421b328b412a339cf85444b9547bc663c8ab17c971ec70c7f449e50269f
zb92c12970fa18cca06244e44b6d5d8af6e96edea8ca72f6dc766a89f88f9f6a6ec0999b4f62ad7
zd916d2bdb3acfb168c874916f8a12ec1385df5b40dd2623f77a0f1544902dc4977cca423ebb30e
z06fb7e29d1d92c0c8746d1bbb954c66ea375f7ceaaf0b2f37610d95f65e1a9ab146c19a7a5131d
z412ebac309cc423b9fb2e127ad20a44ba86c8ca4f890a7f68bd10aa2e8b161a47bcee0b33f2cf6
za9580bcbe52c63e94695581029dc1cdfced58a255699d8739a46a1aa8297a1e21689e0bbc581f3
z6740a17cb8213ce2dfb37b756240aef627478329dd979151859263637b3fba195b16083805244d
ze26ce234133705c033f43e61a5b769f9e811c9b472293b3c00bd64674d9ccd413ca0630bf1dc20
zcd493b30d398d59c573b9f0fac4df6bf0972e700cd4c8403ab909c7a25d8ded24307240b996706
z93376710dcb91453002c483d188498a8ab10dc9e061345db99d6003ddc5ad886ed069d97e65135
zc762c0c834ab0539440b3fb8a38b9c2d91e60580ed6fbf5e26925795a3d3b36e09a7b235a77d10
z216fb3a5a46fde004d64402e9f909d2a5025b3c0274d83312da6d8bee32430c3672b7208d81fa2
z87fae7857d8c063f7454b478a40081582621517115fbc2c9038a5273218de66f85abe5f92f13fc
zf59d02c35b598fe6a7539cecec93e2a4fe663025d4b1479680715d22fc0523545a4e3714d855f7
z93455737a206dbb551995e5cde1ad47068d779a47479922a6ca1aa00bbce6248c6b3e36a8ccdf5
zdf66baf778ca1772c0710bb5c776c43a4c9326ba3ac22d613750aa3f3328964d237c9f286d54c7
zd6177e33959188032fe88dbad09c8371e2d8ac5ca5745bd75d12bf2d760d5e4c16e850f32cc723
zaaca1602a27448106c3442c5cfdb43aeb50990542669b97a33fd7d1091a00b240073f9ff416788
z109ee593fd27b0b4cc2837fc6aea7f7caf0e16fa587fc5c65d19d2ff8c6b176dd0fe4744a6aea8
z1b34e65bbb764560659783d463cb727c3c9302786aaf0e204cbc66a21cf6a16083d67bb6b48bce
z394efce5c2f7e8ca99d6381c50c2a15be4e9dc7c6dc6d68ecd9af492afa20756405030f624195a
zc784077d8d65785960d85f5281e3d154cc5ca8d333a8d6bada170ca5d96ba84bc5fe731f767fd5
z4b5f011133ce31fc4867d0c0fd14f9137490ae1246b5e6680561fe3b1515b37257f87461fb3c0d
z033bc850253c3757e21b72d277e61a7796bf0bae40ff51ca79278a1e3e59c104d7ab8277913f1b
z6a07307a48581d1841d226c263569f58a1cda777cf7e99e9723096b446d9410ca646712b264e14
z77a3973249a66726a920a6794e9875060b42957750a0869691bc0f45b68542cd0a96abe85fc66f
z0fdab3cc66d85cfd4ae05e52c4d15382ee4540033d0570a5724ccff6109b131a4bf71f19e8ccce
z9d57f6780dfdb46651e2f5d237aa5dc1969e1def0c228fd3f42f314f2d99388366886680d9c56d
za09b3ed006e22318792092fabf7d249e030f6562716fed3a10b8b645f0905b505a90938235fe4f
ze00e88cb48a8bce3f064582ba680f3cfaef9a8096b8ae7c0f1170b605195b1ee89bf80289ceee0
z97d5557b75594496a0a2b0e7a25f9a98f40cdf7cedefe1b2bd32a8bf7e02cee4d7d4bbbce5e759
z4afa337ae315962c3a7d1533fe4fabd5a4f282dce4191e87ab6b61e57d8048dfb680adba60b801
z9add7f0c4e08642cc233c0ef93efd5b242f299ee73d54756965088a48cd2083cdbce2d48ccee3f
z9f76fadb644124c85708c466ce16d096b28553e753bae71ae668522a89f6687812fbaa41d66687
zf8cd7170c6005b7fe7ce839bf0a79d97197e18b41d21aed933f27a8f5e17ccf463c530c692a0ba
z41a7053974c8e21fc27dcc5ab5cb74e486cc880c66ddcd9a03b3f1c7b4180cc54da425ea5fda56
z6afaa4339f2bc976e9d774cfba866aa5d9b2c759374582a43f00a96a14cd4814d8445d0440c9ce
ze6c3f4fe40252b346f10b406585d5e20be27b20a283a451534020c8dd04ae930f29ac7ca9caa89
z258dfed6784691c98aeb0376ecc6e61d322b9abeebb0a680fe6096119d89d1ebfa49ab7a70478e
z75e7b337b55f042dabf37b144f1696843df72cb90e9a6bd804bb57a44ec16e0e09162643ec2472
za1ccf7bdadd840fbadff9f872d59b2952fe2e29c1254b43e21458057d08e6c7d51f3c6fa399b10
z8c0d435fc7964dbf0b5a84daa59a6c3ef06c9c6471b61dae668a9dfd01919f5c94c971c3260a7d
zdb23c94517917150f5adc68b13e56ea27a9f98834824566e1c8ccd0683cff7220afbf132073da2
z9803bc61a1a04cb1223d3bd2674b16b77c917ef32326097a6f18122ce9f8d6c7b6bb2128f7dd53
z279609aa9282c0773eba86e75c536f371b86d42ce3f9e3e4fcb05da23ecabba44ec941d30fa389
z245cddfdfcc0b50179ecfe78a3d34604f3249fc376507f88b6d92478fdb2b1dc6f7d422c5654ec
zab86c94a35770b3d1db4a8a17f2b932ecc85e27fa2c0678d09ea428dc76d28841a188bf6d84bfb
zdca7aebc416d1c2df525235a3e5672121a83b1752c96df5aad8c3bae310e7dd124ff9f33afd099
zce3161b1c2a2e04a8c2d42d6a8a0ffc475f81a1c2994772c61f4bb35b81d029f1b3fdd91fd7ab1
z7177722022fd23b7eade63d0ee29ae9ff9a3ab3df650c4a61f950fe0f357081dcf5300532ead18
zd9e0957d6b71fb07f6458bf872094171e9890e258924b72751ab3ab196371311b79d042deddefc
ze7e1d09ef947d7afd3517a45f4814bdbee0e584d2fe12d13c3dc4ce8f24dbf1f61cdf2927680f3
z1d64017403358024a1caa5d275cecae0e2f12be496f3920615b37e629400952fb1a77d3e389d88
zd516f5f61dfa7a90cb6ad600724a1eea565af77c5a0fee7dca5bf87fde09a5b8f2425de325609d
zfc6db3ca80b07412ae1b3d86549f272b3cc8d3a7df67e9274f2b7533641d39b3908a55aa2c5482
z909bbb122dbcc74d2a1bcd244d88bab80042f8a6e6ffc2facc9ff8ac4aba3b29007df93498e141
zcbbd3c16de53aa60eefc3d30747f54444daf085c51d0c336009f9c813c59427ff515d9b5223896
z2f3ae6c50f4adde68e4a6391acdddbe17c222b7ca9d71af8cbd24726063b1a45c96b7051294c59
zd57935c582e8895886b672ea5a651731f6beb5da1878ec893eb10bf2fc50ff5a198143e8bb15ea
z508aeee1909e72c8213a0e01cc0b6486c3d123cb033f768ba2e96b21d65d480d3eb087ee12c922
z995f5402195ad40db1f58a7b9962a9ef4316bc06e610efc6c2c3a54443b7ab82fa62d1eae8dfc3
zeb70bf44ad3d50063248366e6be7081ff1addd4c3a0850ddf9c74b9e7a8c54b1888c8516b2eaa1
zd449a6215a0db51da908eb7332e00791e27de64f489ada1d7134a8cc0e40e36a8359568f64ad76
z1c76b2e3f4387829bdfc53f3475f81c16511b29f2fc8fd18f8c5124c7acb36e68e399fe2586624
z2dc33ed9b3248b9f05413ae102fa48f7fce6fb346376db3dad4b7b0b6b789c70cdeaddb6fa89ad
z5425f07147d1a7b7a5147ba9ca94a49b1d22b6f8084b63e7ab49fa519ffed2f7f79d35e879d510
z774308c4973a0ba1870223e401849d3c1945b05cb7d143997ac290497f713b00a3e93227a75944
zfb66aae3548d9f30a3cdd23cc88b93b1318b0965a72f959c315033948a7a1062ff80776a035cad
zc7bc230afd9169214724cfac0dd97fc3f424b58ea047e7698732799243be212691f0a9c864e332
z03db41770e482eeb0ece82d8f84a52aaee7aa47816ded0b2e34444071fb53ec6c7346b312624bf
z72106ffdc7dbe2bd88ca34557207ddbad35613a29c142b1857d574c70ec5e7afd3bf98cb25ea86
zc8925d91a60fd48405d8f91c5a44aca6319ab4c4bc886ceecd52404d308662a8ec69a250d3b5b1
z1c679cf57ce234e30682b68c20cecd57a6c3f4f760f38e886d162ce6148cb433074ced8e48fb3a
z393323b35af4a0f3ad38a0c99313495d1e236806ee8db735e039643dcd30eead8ca0b560a0200b
z8c9189cfb14acc4263f2ae54b8e709f525078d059bcfd8ad872638cd40addf06a830c7b3411c2d
z39dd33311d9bb75b5b5500ca42337799d736be539c95f4fef48efbe72e7d451c32ac842dcd61fd
z2a4356e0145c00a6b998cedcbc789945d6f878e1e68058e1a578e4c0e374099cd9ddb077b5486b
za08cc1621ba85697e5d2f4b090581f3a6836fbb7096c772d50d182df603ed46e71233599f6f7ee
z0eb3b2bfabdb945ae2d425a94f46f2c1c22c1da671a6fd9b261a87c56ad4037e3df52b2291594d
z586f8b3d37bb2e30969c1e20ac54c389c9a9a626be0b0e11c41c90608c89662c17f8cc8c019c5a
zd237e249d9934bce927c8d5aab3f7e85e32e9d7af9146b36b7e26a531c5dcedae622e487d803e7
zba271bf8bdc0ecd818d6cb24e4c660b5392e8c90182e9238dd763fa823a97af6e3d4042e5e8009
za3ebce5a7d86f28cd4767b6b2b9e5ae6e8ac0102359700cce3ee990102acb52b0328be4a5182e6
z0eafdae3ddeeeec0baeaf1b88619604035a2a4fa6445eee9cc5ac5d37ff2c5365dc2d8fbf3eb3c
z78833c0d715958aac382d119cbbc76ea5092c2ff0b2e991e2b1cfd8b84b03c2e8f891765abcf4f
z0ebf43d09c045f926db140374c6753af2fbcdcf66cfb0a36227238e741df016d7335f45de40a0b
z4ad60c94523f8864a2e6d853412193f9101104293193e7e87260e6a17ed87ba293364a1ad2dfdd
z054909ed2c500dd59a6e0120ae1a2a23f6be4a3f8d2894621484ec6fae64a61a448e7d24e06d7e
z8b9d2e1f0822a1bbee0b603949fd382d9b34aa7b0beccec9b9502204337470e1f7d6e71fc97b53
zbfa0fcdb6d59bdcae9c2d37de2bead7f5718466b238a8aababeeca301dbf9d3d78ea802678955c
z0196967498d64f1a5d0df175888079ab369764e53839db66e522d4c1e2a7f51fb05ffcb2bef2ca
z348e3c565127c50d1d9b82645acd83232d62a5e7cd43c87246ef6a91e6ebbdc9188a980ae2dcd8
z603fc4c81fed02077b6f4b5277a92e5b6ad9617e1005fd029f202cbcf01c56c66b769415516cad
zad24a0aaae93574860f57889ca96ffc6719b5b317e84a7f50f5937d0a05af8978c9285f8755ba8
zddab4bbcc87f5c1126907849d16970608c52eade6105808db4e2557edb963d7c12228a4eefa9de
z30837e76383936e17074d37dffd4b0d2b4c9195c53b7b2783eba922da6fc9ddc2aa745468b54e5
z5bc8a82347e84e634b519e2648cdbcbe17ec4d33552764dac77deaf06ad68fd535d48b2cf35492
z5469782d079c470210ecd202fac3d457b4c24ab7d25aef1391b120f4260c818e933a548736223e
z0e18a78ac4708a5c9002891886045d164bb69ba227606da3a2926cdc4716159fa1897e52361109
z827a0ebabdf5b0980936e4544a4ceb7c4b2872598e766b22a42e8fea96bba38ff806d0af6f8157
z8fb948ff6d82caf37f572a03a3c1b785b3eff52266fe58a90d4bfd94aa55c3ad63a2de8523f730
z924695fd0444010a9db55bb82363528cd7213fddcbde9a91ac7b8b8e9b5fc85ce3a56ba3c081bb
zb4e82f2278dbcc76ab979f536af93bdbbb12c3ed646e4cf46a8dad686ff75e65e968beffa178ce
zef87fc8cc9257824daab6f5bdc6fde58f776cbbfaa583aca122a908c012d639d0693be5e398eb8
zc785d15350f639df6dbd45a357f136a45c5686d08fa7a653003915d3c9a1559636f529227f1aeb
z22a993f0190241cb889002c2bc2357b408719a3c5be542b29a4ab32d61c61ea7ae2ee03e607169
zb8aa2c7ca054f9625afdfd136b13dfed621bbbe0a3ac18376f63f0cd71081ae15c9bfb5183edb1
zcaa61b3309a79e32536f74a6cf4729b58c6c512eca25166bb51ba502f092f4ecd71caf8801b6c7
z797a982a4261b34d0fad715de7678b25b2297b503c4e15e02d14b1adc010ea4584be004453c290
z49d68121401a35e750c896d867969fe2eef44a98e860384451b44366a76d56dc966beaf5e9919f
z139c68e3e24272ac81375c8774f2145d2d2f4135e27305bdbb5baaba072b1398d9e88bea074054
zc29f01a43df5897ffa450c6cfcbaef2bb1e09547e01a859a59192b4b734270f8eac88fb0a88310
zfb0372bee85e0e3bcac992f30cb46fa091ca56507ba2a4ce2c551386901828d329f3a3365b66b0
z9ccedb88bdd32447ed774fc52f1070a0f137db1f87c9e4058c48419a7570fab12a52b863ff2add
z84e58ca1cb7f1c09683fc72aeaca756679daca7fe79d497da8c86f5f7cadd6d3928b8c2512c323
zbaa216f3e05d32e6212cd6da394da45857074ab661348bc50f9b34700dca5c43ce1049b96118cf
zf7e8b48542b89154ded643b3bc2464ecf1f22bf9551807fd196515f980592d3d7fc9450dd79d1c
z810c797a19cd62e44baf1896c97e8f70ade646a65f6bbbb6a34eb853986364d70c51ae524eb125
z7c0c2a14395673044ea2e8899b37a82f64aa3a1a12ca31077e8ab57c11591265c325ff08b54cbf
z1ab5215c0537c4c811317cc967bdda0934609be1126c7d0c848a3ab3b31b90159a365627632e06
z7221800be3737538977834f39b9cc886c63feff5797f77e5203b062687bd7e393df91e6886fff2
z847fb681b0551cf0c77ca8bee13e4c0ce29b77d9d9d854c2247281c4117cdc178830c7f42d67b4
zf2833f9453b3aa02fab6ec35a5e3d94269c93d42c83b06fe730cace2b0406e127eccc1cb01197e
z9068b4381c4535e9575a0076dfbf283d97b99d393f560982f48f594e15436ff4a5fec72d975e19
z61dd579fedc1470835a6227ac46f309de28bd7a6472e8aa10b36fbb15061310387de2ca1ae82bc
z44d5d9bc1540c78e87a1a70bd341cb1cde8abfdffb859ed3ee3562902edf23313bf0a9f3c87c80
zee7da8a01063be80f52be6081d3ea33aebee699c506eec29ab303072817a1e4fd74fd8f541e13c
zfcb02eee41f9b5acd0678f12108c8c9cdec28db11af480f340ed8914c21d22b35b14b2a4c2afa6
za977c763d5e0160af47e66634fea98ccc03745880b2c81f710721d1cc7658770e06021b2340092
z55a7ea9361601f44cfca4dcd37bc432bfc94f340273ed302c187919cf65135380f30f778f1f299
z02e6003497b9f476835ea6b12f21a6464b77ce6f524847527c8a72aa96754c0b60107a0968b19f
ze9490c48df183d45c701995e3d8a706187282cd1d4e542bc41539d8ec16b9bea6f9dd3dd2201b8
z501252917c38643bba98cb534969470a87d34a3487174eb29d96842394ac66b35edfc9fc479f49
ze71fdb5b8159310c94d95f027b3e3abf84a0133cb089d0ffe1bd36e272b0501c9a13c76c1946ca
z139a106fe2a08c3eac70adb104e44dce99bd04c4677a2fcd9af43ee9a383c4d506b46697110346
z07426d573345946d55e7022389106947241db42dfa240753cef33df139c74deca36aafc66afb12
z0dbdb2342ad46677fc6779f33f4e3ac6c810dcd6fdb9756f8269fc5c6f82385c2cca1af6233062
zbc435ca7449207ff1c4b9efe402f27dd427a54844d6c65045c1e2770dd5a8d0f1d83016ec8209e
za6ab249f6c1434ba9976e0b9bf0818a9180eef2c3e4996447212a83c5ce705623740a16f17a0a9
z3ae2007ef85be8a34690b22a3109f3638f3198771020a1a19d52d03f4f134033304083a4c79144
z771ab93e88258819c34d4eaf8ff55b464ffa328f5021c2cc3e43258aecb02f9288f386ae371c18
z18a83b81c569a44d458ce61535402c11bf612669ed9a551f3d9086eee0ea99c296614ff73938c3
zf52524c05940e057573b1259e76b8dcfd1fc44f53f51cc3ed67194948903b94234f150b10a2bad
z7a70e4dbc00250b7efac86fd4cd3cd976cd7467a3f848492f693873422352cc716866b9649eed5
z90a5cff7409d5dbf897a0775bca8c71f9b7090b7d58d0e9c0af3a3d28c4b10ba501f100daab433
zd053cdc8c679b4a3a30c0cfcbeb0d12e6735eb8737119af11c4dd629618a9068a71fb861086ee5
z62da2b8577fb70b96ebdfaebdcd95095c0bd7deade0d451f592ceedbadfa59cf143c83f4c86bf9
z213f4fc32941e1e57afa58b000209f05890b27eaae9eba3a88bf8d4aab4a6a9cd5d3de10bb3419
z839c4a6a8d7d13ddd77444f2a9fb0301ab5ebb6700a78c755ce27e9671cfca1f0ec19424a2d8a9
ze77f1952dc154fc914f435cbfd7a0dc3376b3a1894ab60477bd73ffdf352383ef3404af734e58b
z7d945fbb4dbbb03a5215c95bb680e475f4a1be75e5423aa5d8e15d1b8adfe6b44f73f0e87e04cb
zcec5b33522cdf1ead5c42477421fff29b56d415650aa9957f466c2e345d54186e21207897ed47f
zbe11c828d17fe13e1907d3426cdae0658c6ce9be333d213bf09a88e348aab27138557204c3df9e
ze598c4cd22d5baa16da63db7dbd583aa80271e46a0b918b38080e4959768bc84e189b71a19b108
z9ddb5728b1fc1d323973a257042e7699822f1b3979f1ccfff4a20947924d64d7c030e14e99a717
z123251f240d26099f9191ed5e8de7b89f1868e2234f4c22719d70babe3dfc8c25cef2a41cd04f7
zad58a996b8d297d8772fafb42378bd4a68c0351450124ec18b454bcf11f1f88abcb99fc4336371
z39108e1384c7e11d36d740e3d1e3a30e612799c1251757f2626ea6a8acffe4888841c27b862540
z49b52cee4b1a443823fef24004499ea00bfafb10acddc2c8a649ae4fc6be18e68c699f47451a9b
z5ca487f6fbc9ee32f53f60282e0438a26be21d424ffe7c0ff42afa2f0c9e035d3cfb24257b7654
zd79770d6d0762c6a0271756873f5ab66ccd2f268857b6f2d8304578562262127611b91d723d831
za838e1b1b5240c362ee2f738527be18319c36f08787392d5b457dcafca6be6ace2df7677ed2c86
z0bc5ad98349c336fb713304650c96a90401160d61508340f6091ac887f52ca8f533c8f40366a17
z824a3d7547c45038e8abe8606849adacbc46bac42d7de752e12f491520c43eddef387e2661f84b
z9455ee241e6fc70604d8b3ea20feae71edfc56d18573b60538552ee07df7696cac334a09c30793
zabce1784cce67c283ecff3cb3062fbd0350ac1764a707b4d687eff29f2a574dde8be364573769f
z6a55df49be92e6761b03032a09fb9177d8eeea9d8af03fcf6a7f558be7a6ac70be72bca82ccc0b
z3a9db0e1f3733b20b1c818f577ad8fe5d4b15fb87c2f17a24d7e911d789d1b35826a0b8113b5bd
z63c479ddaa8517cbf864c07ad512db1c83885b8c863fde2edcb3ab0604dea99507d5500ecf2da8
z72885a816ff9ca0b67cb568bac711869f8c075700631edc748ae12a6a2c7384fa3ec0726c83252
z6cb3c3c52651ceee7595baed11ab26d84d47699b84d206cdcb03a68a9a02230b97b2eb96459d5c
z9eb101bc237f8185ad85625e42d1d3c0dc8a3d1b6cf5fe0b3f963906790a5837e6d4be56a871e5
z9f6c54e6d09cd49380758f12587ea092141d5dd0ff25124b7bbebddb91d1981baab20bac1ed316
zc5ac86c5543cd80bb0d84d3a0d5ea0ac417a0a122fa70b6cc2b2abf215f4679385347031faaef5
zcee033c2f0711101821b95c4a5de614d8241ab6330500ced1b8cd0a13fb73bd225a131c8626d32
z7c5a28ffe928eea84db34bd3570138e341fa63d5ee44324d9aafa462cb3890b87b6a6628b87459
z2e6666a95ff770dac77a58bf59dc1abe5a38156455cced218a8235d409548002fadc16e8ec9b99
zd4d7aeb4050e87945b8e7e992ae4efe94dfa6342bb820f8708977f70b900ca6c7c3c4511eab7f6
z5ee36722522066c4a044e9b02a17b445b97d238343533f1c25d24fa404dc9da9d20879251f36d9
zff4e34efc1249f7c8f462023b4f231497c6a0cd4c0f7723a9ef9d473bb0cc81736369bd32d1061
z43ddf0f69310330f6cafe2ff13edb74756550b04c6faf59311de66455a56c157595c2836c2c91c
z73ba8899b09bd2ca384db5c5cf0a1e504974f4c1b15b8c9947511e3c076a4dcd5e163c5ae3860a
z86e64499399ffc15bb270635284b0e853f2b4ccb3f9d9a8cc675aaeb3ef3bb8bfd5d261e94f4cb
z807c9fe0ddde5bc8ffa40e91398e5e3732eae17ca770714b7f2ea0618ffb801566b3b1deb65921
ze43afab4cdf2c9f094366d2ea977e3873792e166207412de4436c3e0a304f9cd2b9523686be2a0
z82821aaa199d13b680d8776ff3e48700a9e0909c8be5dc045a26371e4bb5a4df0478bf5fc4b350
z4d74dd124ce29fc7738c29568aaa52ebf3d41f4807ed583bf5dffb9638e1841d4f990e24dacf0d
z35a169fa328c9f72b0781012cabae9be5ee5c8cd9ee6e1ce6a420b4c7b536bb1c5b16e11e90fbe
z62ebe9e0463b0b56bf7cf7733e0cef4e650495bb3408f7ea25727b5169b68b50e2033150e81843
z01250ee32be25aa7e9204ceb7acf2bcc1fe50a704202b9ae8f653ba535d8861545d230d0a46a7e
zbcee66fb7649bda6392e2787f538599cc955e925fa8311295f1b52028ffdf90ea74fe400125b06
z228bdf6303f489be4b0099bca9a253cf16e34cde2b216ca532fb61de094a05843018d2a408617d
z580ea2a9f2be1700bbcb267f8e8e25b146f0287d17657a0a41d12d561e8ee5b14fd6f55fadce70
zdfbf77fe69d17c262709314ccb8c3df54d3f3b6e74d72bc8091f4b3dfeb87a341b5a1d093902b2
zbb9927e1a594e462b8d8102eca195d7aabf3dce6fe52cd2132f1f036176f3cca799e80b5e404e4
za316392d7de2c004449f6c0a1492b3c766217a1d76cf1afe7bef16fc537017af60627fc2c6483e
z4398a4e95a3809f790a4a051bd37c914a15c0d4a41813f3a377d206ad43fc64b5ff278ae39b55b
z6db1196ebaacb7319c4fd3a0382b93f46e0445f56984dc5b012026c5bf7d43298f06bc81f46a8e
z62af0befef34931026d200be4e3992da0b53a2f9cecace141adfefefc6042c8cce466019dc5317
zb82b3849137176965f335dab34b951a9e5c4bd6601ecea3463f1818c34d365e95d11951f585025
z6e8b36c2aa3e9dfb25241a55c9518bc1c36d41a0edf0d9e456418daf3d7f6ad4939ca2da455043
zc5e07d174c8c27e3965b2132cf15d552187dbed341b638115de67f1163a5861f08f9138dd16ed0
z8cc5ba553886df24f55166b702ee5f88e903c306f98211ae9bf2bc4145e40a74b97b1eb2983755
z88cfb51c0fbfb50f33dca7a1ca0a316a27d711e312ed141a29ce67321ab668683a9c01b94c456d
zc7a3cc685555cef8e8b7d15b1c1b10f9e2c6998ddc569fccd87cc2bc9b8c427fc65b23626e9063
z83fd4a40e28dc5d7f103b4e6f893dc43bb79bae1c2f031eb88fd38b61fa7bd8eb2a3bbec1f4b0c
z5194e255417782825b9669f5d310823524bb24da6387ce0e38f1fffbb5094b55fba05e4d6d6f5e
z13b045c0ed5cbcce7e4a6410f61847976db74b35fb2de943452fce13e16f9e3897a0baf057c878
z0ec7a2731080c15342ea52030367faeed166e29a506da290c69bc050a2c4262518ae5bed268ca1
z0b2dab051564d527b1ee507918b7eacf330796258887563c3dc867635a52f4441bae656826e5c0
z8befd875607ddea475df197c1100e92e511f0e6aa601a6cd7a5a5dd589c6c1c22143e9c6df3aeb
z427b67ebaf107f4b222cbe50d566f801e0da909330ffc49de6e0bcb2d4006e048e0bdabc3e9516
zc2128cd07d1745fb6308bdc07ba630c14a4c91a243ef2d28e6673cda333bb4cd068cb5e00e4ff0
z58695c36ab958b3a7aff1f18690d7f263b26850cfbcaf80387c7ce036143fa1c106424f839df87
z80ebffbc189623abea7d05956f22533307d48b4901487bca008b2fbd0c25c2796b19b14faf89bd
za340c55fb81f467ff52a497a6dcec54e0b40a92e049531c1b0aedf7938ecc64eb376ed13f21c89
z843bd85c70e96bd13607597a4b65baed343d9cf7a3de95d8292c12d7ca0ebdf8dd334e2fcfa955
z0f91c12a7ba3351504d0f18483873c424b4c7131bc33d4b92af27e16c84d049adb2dcdbe06492f
zca4f14542eddab0bf6ccd1268b6fe1f66f892b7d6b10d41cc081709a8a96cd5d7a339b203a7b60
zc654d2def007116a3a498c12a189b684f9c83b74a4dffed629298ce3c06a47ffa1e36f284d03fd
z566fbeaa6f2d70c7d1e7de6d12e28a848d5ca7d089e1a3e12b80dd5359b1562227084432949b46
z0b25c42f33112156a707f25f5e040035e26ff70ab7b3d8ce9e4c138d72ec0cc16ed059edb5429d
z844ab21f64108b37e7a8c3e8c089c4f657296077d8ca7dfcb682f28912fe336b7d452607d6bd7f
z0b8fdf9b277767ef1105aeb277d0ef046baf060c368027198fd6f32e08da2cd012794345953728
z7a7a6050b0758b9439bb430061a15a8d2bc905f7f5a4ce4e0fe82f0d72b2106a7ec96885ba2f25
z6f02b92c8dbc1635ff42810f1faedab84185a4b5320967e9fd4ab8c5b18af631bfe540ffe75f28
za68befd9eead7edb4c48ac42857bdc2baa9dc2f36a248239ce83044a3c6f6d62f51c955b3cd474
zf6825db5fe48bc6ca505c1c7599d439de7b6c315e62f89bce80de019abcc6d6895b67d55fb25db
z8e6d9105d1b06be813b597e0daeea446d32235de5b0e45235bd7c40e8c670be071221ee0d96ecf
ze49a3c027864ef8f87b098759ab46a7d6680a86eaa6daa97d7b4f0eb6535e97094003ffc35c61d
zde258153a31aef7dff42f8c919a16715cf8b01be7126691812d36664b1a670322b28fd0f65d5bf
zd3a32a267f63bc457b3bf22832d369ea38582bd9c8ad2d3a830ccc58213f4d1eb495805c630a94
z0d2ef49152922311d117f4e9babe7988c5abe66a227a47f83faa2af675b142bb97ede20a84f666
z59dd77bb1d116ab4209d22564f144e524e4e076364d901e56f884e0c8f7eab2031751b7c7d7a76
z467dfa27de5226f6c42d7a7ac1c5dcf8988db90ca5480ce17990ea9c23a1fafcc3a2757e92dda6
z1fa8fd3dec2092a75aa6d9ee39d69cda0ebfcaf43a1108ca3c439420e3f32f228d2033074a3f88
zc9418214db68ca3ab91e39dd52f589deb1a8a8d430a4ad8b989b50da94d562f26db1061c943449
z95f901c4bf51ff9922936a9615a6bf494df7b39636b085fe3bc02760562c10dd4676a1904a8477
za29e1dcbbbc2679da001dee74ce0377ee8bb45d5ed4104750d8bb0547004a46b465cd92c2734ad
z1ff63f1483f21db65f287c3c2b6a4ad8d9f18d6a0d087d92c11c3e63f894a75c335399ca8b2286
zfe9b9c06679b2ee76fae756e305a403c9104613d55a31be7786a14adc4e3279d3aa64d34f1ac59
z5bdf7765f4a64a22029642da29398a94952a2fc516049eec93423f7186978f473072ecb6aa4b70
z28d3db46e8af49d0e1e72100a7822a17f8f57d136d818fde79266cf7b52725d31eccbf9ccf4eb5
z4d623f11ddcefe8a8fb71319d8901dc12e2394ed5ed8ac42e39047fd072a43e52f61202c252fe0
z4c615eaa9da0df69a4db13564b2e9d28c0e625e5e999d4adcf77b17a8baaba46979e4fb2598b84
ze78c9e809328293523e5dc9f0dfbdad3ce5a0f3f1dbffdb9f8ab4c2504eb9d24bc1378970c36e4
z3b950af020905b3e419aebd2cc0f31511e0fb806701d91c7363310df2c35f65fd33d3e7a4fc6db
zf1cc05f059a49af01ce673f1a4c5d8df5856fc85291af34e5c94bae2be6d84d2dbd2828f3390a5
zffc41782a9e7606ed232da671c3e541a5c460ac71ae49c3983f4e3f957542cb2134a87e27c786b
z529e3c72b3252511725b7eb2d34490ee91efd590474ff02be61cee6fd5089a5963cf9a32a6c3ea
z289cbb461c4b5c162538a7eff9c4f62faf1593f4cecf6d6eb14d146c96a46f1b88a60d84799867
zede144c66c17f84435f800da1331e76424c94511693906322b09f2efe0219a1881187992992a24
ze8c434bd7f5ddda3bf4eb9d9ab1862e4bf9078545b5a95c605c495b988ee558989f3d9c893ceb9
z33057a26dd7c2352f5eb21a10e4f7a93ef1d15754a6cd9fd260303664ec4b66d5bbf40c624ca55
z8183c63868c8ca6f54c464d5d7200c826d75f33d0b565917e6865de14eb14a4be7c2ea250e07de
z2e28d6477a593f3094ec9e4edfa367871ed640abc85fdc84522ed8128336f3fc83964035c767f4
za34f0dca539d729a6c5ad898cc6025edb607410c989958b26332e481988e46bad4cf45e0dca125
z259f26beee4cdbf983c7336f62e162e60a59dca5476168746058c4fa084e80c868b8c8bafa9a13
z72a4353a853b24e1236a260efd6d9e626a807d34d7d73f34ab80e548310827347c0567071bbaa6
z2baa273c65e528d1662b9637984a16d4caf0f8d16b5ee818e120c78ece8fc4ac560ba9214409d1
z889a82a8f646c37f2e6cbd0b0d4274bd99fc65ad5995662fe5947fe117d5d2b27eb1ccf8e4ad8e
z321cac7c2b44d120daaba52917242676df97c201de9ed8e9bb9e4b78e1c95ed60c164cda0a0aa0
z7a87b2581d942da456ea141d08f5c20e8cf35275aebd92ccc80c17c5df9c10471ec1209f2a62ed
z16a3d9d684fdae39fe2051504f39b750884268f3affdad9eed8b3dbc972f046fb9c3e9553494aa
zb9da2cb1028e3352358293cd86b301f3e2bf049d75cd4adcecea1d2dc0e4a81699c1d643aa529a
z662d4fdb881754e1fc53bb8122e202ec852c5cd4530e7eb92042b7a8a85a3e0ad80965f9dbe303
zf62d6c6dd8ff8dda22ab019d95faaf7dd7e129100351c59b5efb93cef010e2c84f8900b9fa1e93
z27a9b4686f5577e53a1e956459873c82aee240694b67a192fe03c3b5c7726b312f6176153b79c5
z9ae297de169b3ec73cb2882858c87b938a35c12afc99c034967c1fbea042c39ced1db0388d5c69
zdfda2d93ecd925cd25a9ff8d7d9d7a6fa971f216bb8880dd495ec6d329154b619ae8a9d1db8276
z282d51cd9fee62fe417a9a92bfba4efe7f89140e3e50cc0de1ca7057f7c13ec1d45534621d733d
z328476604fd493d33bfe9e1b332284280ce66ece798f88a18b9139d86c1d7d7ac0f8023c9cae1c
z9901098fd7eb1257f6680e047765ba898c14608c9c93d4c4378cc606e7db74a3555357db7e4f89
ze509cfbd148ffc34bd1542463e4606f9fdca91f3acb16222fdfd2baaefc883f0649fdcdc90f11a
zb47d092d94a3fd066f93da03d028f005817f8499a89011db2f8bbf855de8d3b8f777952ff260b1
z04e6551d63d29319f61f2d3a0b7261c2ea6754e9b20b154978cc1df7febe1b2a8beb1e855591f0
zceee58d4174923f693a2ca655c46c62f5467660f99c73172fb06b098271e82bea803574211538e
za4a76dcf15a602df633b8026b36e7c6aed1813352a4b1c5d8b65acf7d61064eef3f69c1036087a
z507dc20357c784c40dea6ad377712013dab8bab8bb46d3c2cb329f20eb16e0476b500ef3f49308
ze1cc4f04de3d100ee20c96708f4d296bfa30b620a5b61143ef2e30b0b0eed923a373668ed1b360
z7b3f283d02d550b6973ed747881d645985cc9226c5b5a7f34b268ad9095fec9afef039e5af9891
zd62b6b40bf9e3d47b0a81a03fd7d936f70f448b10872b91f988367423b4b900c1b6cd7b537aa54
zdc4c8a68834c94db47c55054b55202e9961774ecc29b63de820efcb7c02c4b19511015df7a0f80
zcddef7f3659f26a324f9487a01d1d1825ac31380323ba0291f9f2b0899d48f3addd6968cf29d0b
z6b6cdb35a0922c9f740a0c047631423984c22230b2c5075b2da0590f614967ef16db3bd6e78957
zb1479c919e4e39a2d2679b03018951e35448882886fbadcfefcee31df7136cd8139bea89c2a05b
z8c2696a744869b384fbb096570daba7977b1a4b8c7f8438158d277888819bbd1a3cba93ef34f91
zb738cfefd0c30fb0ce1f1e790706967e6355bb5a2a43d38300b0a8cd29483412ec2b862ceff13c
z9db1d2d563e3845e4661e1eb53189a82fcecf208673a57ebd7a32c27eabe3702a5a7722d966fd9
z17b58c46efdb66dcbd90d754b6e23947c613ef1cc0f677184bed178b7afb76190ec0f5efb5d6d4
z49a382d86d289efb0f3d6884576474b86f55cebda65f95da20c2141bee43f490a53d77d361d1bd
z37a7c013b0f7f08546da23401d3912b3692d1c9d8933127e13b1682c15e4e7e0c131fbf53b5f36
zac9336bc6759851eb66fbc160df71123107e47ac8ad679eab9c2efbc17602118950a4e69ba2c0c
z9a59ec1b2d21d0129c27a7b8350f3b32c951236e3c9394804e97dcd3af3075d6b4368bb5202d36
z6868131d2c57e31d07a6ac0e766dff901f688033b6b69adf711bd2833eb5bacabaa8dba0878e84
za8eab1caecb0cc7688cef5774a09bd11d3582fdbb4762ecacfe256b74d406eef69394f0fd6f3cc
zade0b4fb1b61eeab2ae9b268fdf4688301dea2d8f903b277c08835bda7954b66600036f4ad2213
z123b9a0318f234056de014c3a8fc355da8c6e3674a07bc12a88926f3cc15d4fe5e281ece292bfb
z17400b19844c077f9f727d2cb621dbe17d36710161b6a06ddc0601dd56959db2a825a807404681
zf3da0469e41497d3bf7b869751995b6d9e3fc4b64104ef8a02bf852a98e827f47f101be5a9b23c
z6502e30161e153c75cfcbde301207c308c8b1233d506861c090b1e154a3b730a2a3f6b8c5612e3
z5ecdc5596f3b33d2315d17b81463fb645a57b3db510181ac16da3553cca8ebd01bffb16a0188ed
z2519ece371588a28a538894f27f34d4f4de495109d6752f41e8a3b5652e591f22cc9db3e4c471b
zb9d4c8fcf6b0c265fac61f58c95414a8705c490342eadf50cc98fb9a9dc5fb94a6a0e1ae794740
z67a22bc7292f930803f5290985798aecfc5df91484b511cde988712393ca701cec04d644eeb508
z1f72879e430970ee9ebc14a864f0da94777d7c59a6ad0f3bda976e9c867c308feef50c90c5fed8
zf40f3f9ee35c76fb69f3d623300975f9aa8fb338ec2e4c3345b2969b646c66831c2f60ceb9ef44
z05e0b5e718c7230d7dac11bd8d113faa385d0b8f13ec3c5e99ff7f2e3324f93eb141ea7bd20299
ze94cb23de15570286c2bff980dce59cf705342588bc4cc1f46884b25f8413705cc9f0848569f8c
z13296373a611d6e1e1cc0a2c99b1eefb08bf0deaba2f0f47e025c271aa57b89450fb9323f9331c
z95196fbe8bd8d7ac910239090f8ec2b41713a7c981634185d6ad9595696e9f2a455708484fed0d
z96b01f30d53868082965aafd974d69195ee4e8e52c90896dc8b405e8df02583505875724086a62
zf75fd9c8fb634042a37a910f2bea9132f09fc346032508ab59e56b69a9ef64e7a9eca0978b0ee5
zeed01b7b24c50d79023368a5919d41b010d87157b3fa3bae26606146f1288efd1d2eab1237b065
zb65ac1ea03e39ace33fcbbd893d057dd16bd3906886ed8e87880a5cc7952d0d044aa601dc9c86b
z96a2999121bf0aaec0f440fc67ba3248303efa2d678f0de133a2ed558c4e7f11679e7294601f0c
z8cc12a88c727762919c4d3408b48d43f343f6b67253daa99666ab28d64a58d2b3d981964b31f31
z969691bf5d5696305b0645e5e3a44079b689f08f27d7332247bd7400000167e8c79a5e12a83456
z3198e88744620c92bd383995829f408289432fd9ea4d5200b4ba246a4075f54f338a807d057050
za591f4c9eaf134bdd4a78d5f792150ee7f2fcb4686022582830bad67b7daa051f7883a484224fa
z3d33916c9b7d8c5c040383819fb322e9b750a6fe586efbc17f215b7d1403e2b9fd22b089ed9faf
z02d96e74000d2133de26e3eecd65704eafe01f4604918f1de82a513ebd82499719438cf3a9e7ea
z68b32ce944a161ce99b302f9a84bfebfd3f4c7f186cf399c542768c4d47e925442830bbb65839c
zfc06a1c26f9a3ad053c9aaa082c3ac1a9c5ffd063c69b7f166e954f55edfdef53e72661671412e
z11a821981f516d506540cc5308dea089393d48e5ec3c3a8a81aec9167e4b643cb0575f99ad447f
za6b39172d558e0ae3a48fd72af02bca124a3310721763d4453f47f99fcf2f7eba220dfd86a5e7e
z38b8d32194fe9119748247731ce559d0edcfea0f5f70763eb0f85ef22a6bbaeec57ef0e88c6a04
zdbf80adde937e181dd250a808dc5ef0a52ef10fdfaca8872c9175b4cb828957212230477a3c3c8
z6197c28bdcfed0f1cda40679c82bf35b8c337f87a6cafae7828c29f39358f5411935890fa20cef
z2e3f6249349d09c2f5b48d26dc4888ed521a9f0def7d05140340934bed0259fbafdec440ce32b4
z4c96fc1a8c976ce3c93b35fb87828982f8826c9f70bf006e3d3e000c50baebd61dad69d3871b0b
zaa4047cd12a10ef06a3c26e8b17fedb21cd832590339489b5a166d9cc55ee06a12409475c55b07
z04f16b869944529a6a2e94dc61bb6f9de480065efe02425a2823eefd8c4d8c8149d1676b7c14eb
z4ac60e248a494465ebbb2f118cd1d1ea84add3e9ad8797b69fe0136f9a2b20c047bcfa38a2212b
z83d41be543d7a377ccc2203bac7b0b652c49e4d8f53489f0013239942c45c60a0196b3774cae35
zdffdc699fae07212d156115a7c4e76e020e84340a19de1efb563cf3c2bb013d6dcf19e3fb4d182
za52a7dbf0fc278d850dafec07763e83af5e9e36a46bcabb34e0df7ce6ef960550102e6e289659e
z5775663ca0aae14c53cd3c115df3239773bf46bdf4ef063230b76d88a09b345848601fd659b60f
zcb9a5963d3445319bf3ae2e9e85a0dc6a43753480b54c48659e1cce54bab029baf80fcf544c509
z6d9eb84298a56d80742d781b088be897c125d026969f3b963eb4ca1bacdb93b7c26b6a12192caa
z275f4ff7c98ce0b079c67b68ebd4094e27fba3d240831ff4fff4f19fd116e6eb83033286f263c1
z6f7ab3c25d267f29106115ec2b6906c758048ce9a046a59dfab6216f978a7dc16080f9aed91c92
z39dff1cdaa5bc8b0fad030aaf65b0fd316b1924a739a185c161e766e592bc920cc0973de34e043
z5c0bd94d3756331915da3dca0fad2f4de7f0417fb7ef109ddef04bffa541d022951e7b208fa344
z8b796ca7e5929d41367b01c8734f633612c24dcc2b1e964d2c8f4e213c3eb9bea5da5e7fe68d02
z41328f0cc345a6cd5cc24c125742c8e56e0b559e763cf3b3065b212a1dba2057cb824aef6f1839
z708536d2398895c8afa55c7ca7cf8400613553c09587d5c7d18d5b1ad821dc11c884a1adfe8e6e
z50bb6a4064509e5c60d073b54708f49dd948a30416cd961533544739cd7cd50f66d05185c68c07
za808e17d4ef2b6365f9ace04c7853bbe80d24b462967aeac9395a3d779ef77a94f39312bbc2345
z89811644061416f951d23e6484b18bc6071e14738c1422a132b63d36110ca9fd1c42dec4a84932
z1514f1e3b800c6f33768add582f1ed2f2af0710162a87e3452e5543a3a4ea1d2f923599aeddbc1
ze53e472d0edc2c38960badd8460bce6b6ca035cb6f9bd4fd66f32d9a248a8162b4e48d0cc9e94a
z54fa266209c39ba050ce9d0e052067806f9db3df29fe7135ee259dad906cc7d6aa98e3fff549a5
zff550030d81bf81e715d1856aa008155b1300c39928fa968978d196f52d85aff847ecb5c6b5531
z4b3eeb148b671f681a679e42a3c71f0b1f9c44f50ca3797284d9d18df43cd47346f7af443ec8f2
z9bd7f3098f92265c23ebbb568dcadbd42c10d119bed9d86e5f00dd2b3b9aa6a950b79230793b38
zb0ded1a01ea2f85b4fd41657a486f654de8f7a2162fa8cedebde142e4934ccb8687840075fb2a4
z860277bb511a96298d4b2b45ba344f45379fcd9c965a8684da071de86174abf88065d0b758b4a1
z6571e9e64b07510294e784e516813fcf7aa96a1440cf674ec8380116935de4ae61a57756609079
z6416d30ebc9a8e2e78de80d410401c9b5e3ea4f75430a88bc9b2763554a60731770d7e21fa8685
z17b8f4d97199617531a4d08ed86a65b10ef82054abca57c2ed73417c2ad2f5b44fec65c7009404
z4fd755e0b25842885992a03ddce36f7702b298aff69c1da2dbbf8235a5e3883042ece1a4e8973d
z3915f940f963afde26c92810025310029f44a26c5412ff7f8868913abbb7dca613eecc52fc457a
z068e1ba44a7da708869573b236717a78fdb31e23e0522aa95d67771191206e1bd71fe43454334f
zfa73edfb8a62b8ae5ceadc63b151c4e8aac29fe1942567b77e24a811824b0d0f1793e004a3ca54
zb6f19b276a3bf0a94a6d586243c59d545e3406bb6cbf16ad8ce4f507f0555a489c6b753f8420ec
zd92f2321d45a50c987140df3b065b2c8b6c0f6ddc6466fa2477fe8c0e548a6aa020aa53ac9aa33
z3ddb7361e5c7d3e63be8062a7290a2001059e8aae17247c5cae31bf140a36bafea1c6a8cb6e450
za92d3bfea3ddb6c76bb30f07adb5f7f0dc256d357608ec732c7a35c02e78fd00d0012f7701da8d
z5ea79d76df0cd94ee25f5d7868dd7b17d4f75efe848bc99bee6f0ecae64d9e75fe8b88abab508b
zd3710ac7d2202980f3333bc4382a99e370a54a6111489554ed9c83eea25f74c360e34519f1f521
z17a376766fe1a48f679f768a2e79e45f08b956e1abc9150805d05389c28680b07a3bbe491d3d35
z0a9311669e98a0125c1fa65ace3fa1ad9a992b758a593448b95b86952bbdea925d001235fa94f2
zcdb676eb964dad13e26bc266fb344568efb344946c38b68e4f911cbcffc873c109e119cf73a574
z99ca95564a185610af634d1193b9098d45c991f478c53ae13a626fe8ba82d6254be9a2c29f16a2
zf2c195b883d0d0583309acd0d5c6bd30d5883c39704b38668c7681d175ec9a4a965c5496d45b74
zc97d5ceb431c785cd055a6bc0f3bdf087704a200ece5061e829168b7748cd234d8ca14b0a0601e
z0512d559e1a571decc6ed460ae8c249f91a472fdb2d955f2246d81fb3ad472eec75f6d23bd4784
zf587ef0d4886484d917485f46b58275759424f06537babf523164ede084cf1a25bc3accbd97c9a
z7d6d8f44d7c7f37c0e30cae32cff2bceb1d92f6438e41122c89868f55987b654bd6656df935c3c
z4dac4054005545223ba474d0bbffe3757f8fb324de4c55fe894b66171ca0032777368da658cfcf
zda75635a686bc71c94b4fc4693be4cbd07c07e8da54445682c380bbe97c133b4199d360e4443a6
zc338ee0b644aa39a442e884e0e054cf0ceac2aeedfa6e7c8077e77f1cd9c9d6f75ca2c33030fee
z162d472ebee26408691091fbfb6054304d8ee2e77b3f14bd51f2eb494f05d54ba25b1de24087ce
z949f0a74f9d8123dea6715e96fe3cb829fea72dd1cb158d7424cfcbe9887d0af104f7e89a6984f
z87561472a8773d8e57b90d377a7656e1ea22e8e230be1bd981d55fa25b8343c3474db33273a433
z6d79a1bfac330a1ada1bbda22b95ba5028797ab056a1da69f0656bb30e346ec0863761bf42231f
z02366772ae926fdfbe421353209edfdfc4b3075f237b678ffa3f498c76b211f395a3f7aa9c7f71
zf4df604422c39abf04b1e167038d82941021eba46136256a614a5aaca1569d554e2e258b0d140b
z135f46ba14a3fb51a8776e4475dc18a5fa11bea9b7f381b2549249a150e99adc3a7106551544c7
z5e3019e186066dac0ff78038ec40414e37cee845e62ded5ebdaf8972b95598420dea3cbba4359a
za8881d947ce599348db569e52be10452aa24dc157710f2d4878f1ceadd06db0855d9abf290584a
z2155ba40200d0fca9586505636c3f048427ea98ea9b7fb208a59ec3905c290cd326866030143b1
z9ee52923c7dcaf4f3f18d4e34a2d220c552090946d9e51d284b9e56fe1604779713498d6f1c197
zb72accbbaa91ad9d7a3315cced1f6a3ba4b297df518bd966c3519714bde45b50988b672ee182be
z168321fc207af798a7bcf19c7cb999ab21a37fbd5b437ef41d7f2444c16ae2a48849e840ea753d
z008f0e2fd65ad4d615f0331ca8fd88584b8bc906377b92b7b8a5e37d9b0f5b68e8ddfd12e542a4
zed5f0048157d9edf442f1f8958d4ee328632f07e3cd633442c16f4a167ca159026a578bd7b28fb
zbe1c8421e1f8392ce57002d4e6fccbfe3faeb6d03f9f2a4285d86313e9465f7f0dc123e7897283
z7aeb3fc514ab48dc856632bb200c22881e2bb985d6b36770a864b95647a9036e35c77003c118e0
z709cbf2861e137700a081efb6eba82fd925ac33cb7f7004ad45067cf3a34b405182cefeeba75cb
zb5ae5057f2fade7f2920ec9557cd6eed17d25858e7dd213564e94168b2f53d31a8910702e589be
z704b3dd275484d49980280759b2b3934c413f05755a6c7fb396fab8655821fd9d094b5c60ac0c7
z9200a88e6ab1d1f98df193c707bbb23c0321ca67b13ed6f1e5a7d4f64f4b11418dfd2bc3eda076
z1db26e051add73e754cfc189100980bdb78f01e2aae04f7da08d5239c9b328f5d7eb882bed00ee
z30e8285e286f47095ccc497600ce9725b3b2146ac8da38ffff9dd782f95db7548a85cf4df0d9ea
zda8fa7e26fd444f14e6ecb55a796bd995c9890d7029dd913584e0c81b759dd305402c87776ce28
z1d4ee9f7a2aad274bc7fff09675221127f0d21da80cdaf369cca4407c5f4e9534d2264e0f6156f
z1fdc28907b15aa16d8180652f5d114ac997f2848d73b20a704b83c992ae2936cbef3f14fd92fe9
z6c351fbc4f66eb548ab6c3c826e2323fe9d9f92ccf7787e01f9b7a9bd644deeed9467cdaff6e42
z940bedc0d2a9bd8130e3eded189c06433c562e54c999c1413dd9f01bc5c0adc5949b6a697c95c0
z6484403485cc9def34fdccdaf0630c142200cde9d9deaf30a9222caa8233b9beae790e3747dcfb
zf4837ee09ca820ef4b9f2b6614c7e580a85ea6e225186718c67dc03174f7c905edc7a23bbaab23
za09eee4900eafaea417329af17be229e52f1fb0b25c9cdede3ca775030b0d8c5a67ce4ea1e99d5
z250745de00ede75bfec2aac6003bf64d0cd6604b1986167ee94e8df616f3c304722424630b2127
z98bb91a3759a3f2a0cf250519e9385fee6fdb852972eec26e0d90e1a7aee229d945ff893b35999
z29caddc3bdef2b40e46160a72bc79d33a56eb7292966c41450fef710ab6e762df3df2a7d179221
z3fdad3f7d439441b448c24181792d6cc7d1a6548117c51c8ec70610caa3d566d2be4584e2c3783
z8b72dacb2c2a737f811a6bfa9dcaa48a1bc04caa04ac865927725b792f49719dbf15deb596236f
zd3096f5cd620ec22647c365c8b6d23a038a6b87785673435b0dfd5f82b7f36e7e64e2e93dae72f
z939555fb3f5ee383a379bb65e453ea6262535625e5f21bec8b88e5a6b0ae6d6e2c8865517e95e5
z845717f645ec914943fc4fed42b22c43d2ec057ee22d4fb1fdd9f83b7b011082b0d38f71ac58fa
z76eaf3e4f400774c3e7e9a61ce0fdd49d411272467b3fe7c428ed5f008b024e87a1ceead553346
z309fd664ba4a0db8b25a0ed5d450a5e7101c2fc71eed43faa82fe5aefa6a4a8d1595adf15da42f
z2f25bf074092a576545033f61f01f39ee12aa005700d15355f1ef847ccd3fff16ba4a155806d7b
ze68546bb87ea82e55328f98eeeb5c2a5f135a7fc2556ac3cbe20aaf04e5b294ebc991a8bc2114f
z18ca6171983a32233f136533074439736b5346d915c34d5607452d7d817b36d05acfe7d427a52b
za4ee3e8164b0c05ceb03ca5a01b35664b98bbed463d38092291eae87853c012118e373871bf9c1
zc82f0964dfba5913e34403cf301b6ac3105d18c65fd947fe7ea02028a9261247582f7e22209756
z6c8bdafbb81d7223c68509c658784a8883aaed70762b5e29282efebefc129f5a16283a2f72de58
z0083248848cdce308be855f1a2f7ebcdb3cc73faf13c3e9e49a35145151e1e1eac72a3ef0bd7e4
zc6183f76b00ea12f1831c1545a64016ed6378c83ac45827b0fc57063f43e4cc4dad7b2a2cd6ebc
z563671c6661e0dd997b014477b1f16a3c1dc8d06ff039572936e2c5de21bc61da0eab71b1bd51e
z7b27c4608ffccd4d136f94bfcf07d83b920cf963f54c177704ec3874b53ec71205c1d2eca7c2a8
zba403155ec598ff74e8e1fd8da29d9779464838729d74c1c81f7e05d5f970452001e8f5e4bb6f2
z8ad644b2fa18f16551a7b960b976fdcbce8d9d1612d8b8f6b56fe2482550171cbcf6c9e6d70047
zd7adfade6d1e541007a332d3a403124a279a08ab5e4f69655ac33b512ca8a3f9853b36b28f8f13
ze5d0b4a9963b8d80826cd7f89ddbbf1cc3a87f5bb53507da613cd1af487b83d61e189382c8738a
z5cb957f37bef1dfa8d3bfee94bddde4fdee382eb68ed1d797443da31a5a870152357f68bcb00d4
zfbe931ec86549407a54edbe0554b7df79e1fb957ba25daa7160b78d1c02acb70d3369f81af5498
zbdff7c8444cd4f8c0505a0cae2cdd409af57f36feecda2057b9e02b4dfd9af5e3e628a83d533ab
z91793e4077f14c1393fdf52cdc5401762d1281abbc4fb77b3d31611f2bc28735d50634e7c8d91c
z09fc725fbda9f96ad32de4f2889fcf24a6bc0d7b637ff8cab03a7095aa76cf0044ddfe84ded9af
za937acd90c5004406644166589d37e8cebe2839a82750af4289a0f53199082ced4b447494fce7a
z6cb571bbdc07e047a9c104e450d40d1f99552f09433748964aaa8b93273612a57934c5b9503924
zdb8e28e13f9ab9bdf48b6c6f3dcd65bdab84ff3bca7b32433d539b4c26818f5918933a4faa1e94
zc807aa004362286f43e56a6ebd131910a17f1c33dd37ac84640b8095b7f8f718191d426f0182a8
z0d672e125ff0cce2a0109e80f8961c4e8b8a3da34d5cab7a28698c3386ae05986c52eee4882f1d
z69e37b253ddf0f5c5bc30196983af168616ac53e98f64509ce635201f6b3e488058df6dbc6c446
ze8b7e8cecefed3b62bf713dcf9902c094c50973432e76552f3e85d1c8c99d45bd8ddb726d005c2
z590ae6e8051df453d1b02f8bf523cdeb2079a6f84a99e1c55b4bf6852c40141d3a635a8923171a
zcdba6c3e295d5030694f35396c9c15ac3db516816bc978f2790edaec6f22bd85c3bbf4482615e2
z82e34ea0dc40a6830feca42acaae56072f89c88a25668c8d19c78d26a47edaa821a6f134562214
zf936390a3d1e2c664b9759f2d4018bf3bb4237db94f4663e1c5190f08dd578df80f23592654e35
z8c54c25940f280729ab965597ab7de2f35c3b0df777ee0fe7b77f7a885b25f13b2600dc4f78d40
z2c565474fbe1071dfc323e0a4304baa6cb7329efedb3320cbf00363bd95b6bca8cc3db4f2ad0e4
z5f679cd08452b1fefde1bc4d62c6ab1d85babea9c7e8ef68bda2c5050733fe26b36303deeadddd
zca9d9972ea0609009d14841e056ae8018ec9a648f21e8f2d3a9a6b8e28306f094c56502f515928
z2dfbf91899a76f12d457e5ed599cc5bef5fa7a6508a484c7dfa0a89e81492d905f665dc972bc84
z1acf70447b174623128a999d2c5113fea37ced5899e5ed333b8f4dec0168d1cea7bddacc5fba49
z1bbbcbaade5b7317eda2bdc9a3cc350a2c4da7122b36928eed2603a9c64c185a653466516aae3d
z96acd56561b349b2ed332ddc47f04a0dce3889a8c24eb292858cebf9d83bc813074558f32f513f
z83fb2824df06fd7e979cb0f3e888f9bb006ae4dbb38fdf6cbf3b57f145866ca3538e16c1b2107d
za9c8f81931e65c87ecda0f0e0008a749f5339760eecf1b799726dc1debd31574e87ed52338ee22
z62a8d15ffe92480c1954ac04982f2736c6bf49209fef2f8c0c1e4293567468c45211ca695ed5b1
z2bc25c8fd29994f7a86c45f0ea7a69718409291d2306213965250be5ccd72f65349fa08510ae9e
z2da5d06dc7899d485097cc0f12ceafb03fed29f5342d1d3248b451e35092b47accd326fff5c9a3
zc372f324ba5430066c5a813ecc0c65bc433aa6c4d97f485152d763b49b3b00ce4a0b28dc408542
zf1d9487b1aacea4635999b0f80723bfd2acb5acdaa291512989feee76cb7dece1b73a91d09f9a8
z8cce01dbe2efe937b93e8cc6a76ac675c06a1b5aaff30da555c7cfebb2bf8a2566cf21249e11cf
zb2c06f9e71b2a9debed959034a93a36c2add7a2d61c9b6ef3dd7dbec9ddef6a98b49000593ba6b
ze74ef0ef2b272ed9135b8c80cc7dc5f6ae04cd67ff34a44a1249551b3a1794f7978cb9c0ef5ea2
zd73137c75a9fca264334cb1ee1966d07b45d3552b175f41c135eb8a75ab5e1b41a6af947cf2636
zed230b372968708df9fbd1628a70d4c7108943c6c1e4a4d90e5ef2079b5d8ec1ef4422cd865f30
z14261a2c47e75e73c43dda4a9f460fded5c3525d715fc939ee63871290548c806ea6780047faf9
zc3b99f7f6aa4bd10cbcc93bbd4939b2fd61360cad2ded971f224e271ca660d94ec4ec604fcb943
z04adc60a85057e8fdbdcbf723b2db52ea36fc145f30af8482b37c58707e8e62d59eeb15be27d98
z26b0c9b9b08c7144e48ba9bbe236d19c7cb94c66b5c504141c0d4b9c93dfa3fb1f6d4061f116e7
z89d080de4d6501941d53b9044bdabce13c88b3d8d39d17ae6aeb192767a33b0fec9a190d630b92
z18f7d82020193d4139bea0afe526385a40c64bd1b769c5b61bd56137faadb7c1b78279866757d3
z2af262c9000bfd7a7852a93546bd00798271652ae66d50160d50ea37567cdc464b3665e71977c3
z14851031237c1933fb5c0241d79747bda418a94c538072d44a44df69a5aa10259ffaccc77abab8
z1cd3ed9cc3239fccd19d69da657c26c47894c165b47521691871e44747f9eabeaab8e9581a766e
z074a90034d470fd685c15e0cbdab80960b54f65e2fc2d47929f114f2e599cdacf3554288f375b9
zef3d56ac6b3ffcad90bf83d1fff12873977f7d6c9cc8313fa62461abc85e936d0b1907f4e4ba6c
zed83c06d2642a98ac5bde9953c0e4de7316f13ae0fa8fae01734eabb3074d2cc19165554fe801e
z1561115429e3e72d177ccca5a44a5dc4e4af99f37b0a6ba87a95a6a3127454da7a17d2d3425cad
zc26326c7105d7796b7cc4ff980fa304bd1dcb4cc1c720e0891c4bdf6f5de69e93e47dd935ca5f2
z147c7cff001bd7d2ae460e93a759fa78c782475ef3ed8eea9b41e74b12346e85b8584884a66814
z7bad1265a2268ec17906d7a0db0bae828060d87549ae75ff2ab4d5ccf876401715214734a09ee5
z8e0a77ee60f59080926af4f314814ad82106efe063e0abfe94f791a044f9fe63f64b15d443722e
zde6083a72cecd98f98824e13af1bb91937a8390a54df73bcb1e13f6f476241a8791ea774bbad58
z47bbf92ca56b595903382fb24bdc4eb9909995e9e90ca4ffe40b65c17e53d4f40670ee41b092bc
z550c512c4e1c1cb4295e48da382ecee9f44295f9bd0bb09f5f150eca0c4b5c24d102c450a805c9
zde6de974ba84e88ac3d66eb69fd3769d321e5740d896bdf0cb738a43105e5a0afc8497019e7711
z89c55f26321e19c758a134711d902492f5c26241d29ffbbe3dbdfddeea12cfe483de6403820045
z37a9d29d788718f0bdbc8e7ae046b10ca301e644fbc8ff642b318cbe4f1dcdab4fc47bc4c7cc6a
z0fe6a5959f8b916cc5d0039d60d2fb09137f59dd63c35c2c75e82e5decdc520baa1a9294a41af4
zf8a9e17285af999f0723fcb76c39c36e199bd942e50be230aedf602cb0ab14bc10a740a7f65d60
zed807f2ca131d303b4bad357a968952c3b714f2ad1ab9a9669790464177c6c355c4148de47ea09
z0520e4c7d776c2eed9fcb2af3cc545618ea958d00898bfaad11650af44c07b72e5efc0fffa0f58
z1fed93c9e508e85c09950d8c9c69933c2d287cff94ddd10ee88416a3f0baf2764362edc7fe141b
z863c69d87b111f0100cc5d11da80fbe787d8e8029ca9297c5cba93938e6b83b4ac49e71e05a578
z18929afb18732cd77839886b5e902a83d29f3b08d1a72087e94b16b2b8b68b3dde755979693412
z6e03218b80ac07709e0a2a20d61534be9cfa3bd4ae1186fbe860dbb2e0cc3acec468f0fb77de91
ze8f6a651958df41b4de9f4d901e5000d0d61f703c658856ce3be4c128182bb5eee407273842731
z56da6130239b19660035c276eaaf0a5a3084435352be7ea033942a219e6fa46adb5b72c3b11a3f
z069950cde5e60c566f69bd8eb084f2c37ee5699eac5db12e84a6c2d46e3c8ead92e4922fd65c84
z63068fba7c7834d489b1e301d30aaf69f585f6a93dbffd8106a62c0edc9871104de7d0696092a5
z25043eb4a3646b64bfaf4ddc0efe8e795857ebb6762f243a9a32e88a4df951bf1baf4f522e4ea0
z7cebfd991f35bbf32969ef1ea882efb98960f1dcf7d0a9a5deabd01aceca2e69d8e73fd529659b
za1964e15f6be7c99dbe67d71cf2a07fc0a2bddf6d91f87d7ccbeaf5cfe9d46fee780e2213a6251
z60ed364ff0c7f87e93c88fada3229a4f2304399bb99d6928122ac46a2c5f60137c7f9954ef2152
z350083582b148e9301127a7e8d677378a1d39a893c01b62d545414ac92000e21fe62559b584503
zdbb2440217c0a93e179404c627b6bfe2ae9dc5709d53520c1d6dacfbf0e5441df49dc4b6141b8e
zb152bf7866ef30f483d17e8efc963407d200506e3e344d387fd227ae0c67734d6964c9c87429e4
z665c6291383609fa0a4b7bff0103f2c145810fad99e48235455c466822982768f1a4cb73ca475c
zb178df725494b085d452c8af0be2134c0b99df5df7773fd9311377b02a44eca0920125858deea5
z967b8bf2088e33c1ac10e7315cc16af5535e8b3734548495d52988d7b9b0482494c9abca5af3cd
zdbbbc862da016a457c37299b7b71088ec20cbe7d1975e33ae0bb395bfdc32052a487fafa1988c5
zc3510d231bb1e7c3b814ff38fa6e0a941a8da8391dbabe636aa5b66c82f4bb70d8ac2dfb7064b1
z279a606cf39f4ed4dec3362c53915f7439a64d6cb56c93d138189c0d8a46f9f50d7ac12bcba3f7
zc44968254e2c208fccad727231d813254fb589f73198dedec4aeb178e78807aed2e5d402989965
zb557e0403b8d0f2e90a9514cba114ac32c709187f00ac69149d64e4c535fdcfba220823d1301d6
zc7177aca99cff118b7242b01f21a19817896658f6d0a0e31b5f3be2f99e4f6aae17925f348699c
z9772e442da0dbeaa38086c90d215bcb3067065c45b5cf8f1ce5d37b64aed2af2612a696a0275df
zea3dd706816ce302679592d16b83291652c3b2d7df3fc8de0af6191b7c56f6f117c274d5808289
z9b503ab6c613cee47bf5b77a218306c092a3b44d852c052c228222de222d9b52bcd7513e83a6c6
z5cf92a4f5a69a5b3889d668093d57eeba986ce7243388a69804345949dc0cf7945adbcfcb2265d
zbcc632628228eec3893e18c99034472ad7a85f80c69cd602d5b912458d834fdd5a1404b14fa713
z91f7d6ee93ebd42371307ea87c88f91d1aa4547a58ae180f980bdd582fa6f720662c4b84f57bda
z30fa81617a6d05d2946ddeb4a766c51d6847eb0aa2d92040c1ec92e43e272401be811f5673153d
zdadbe4a8e5bdaa82d117f52706414ceb8f0f35a04b2434cabe53c5c6e41429da0b81dfabaa69ec
zdcf7f1a4ac1b00e2baf1035d387a8f99e0526025eb17c2556837526ca065ee6656b8af8b33b9d0
zbff741298d97742b35d20aaf20e02eb1d7b6d60218a2e9a056886de65163ccc17bade6b201bb04
z9f11b9fb798f2e8955b23b263f0c3023fb7e58bc47a4460d2347cb35de1cd455b29af6adf4af92
z8f9a5ff9241f376de4bc4c46c23ebc777e71ecf0e5fb17102788109db8dca2f6d8db8e34ab78a8
ze58cf40dc5a40457a6b473b8c2cb0386b2d1e9dc55c3d319a654236956aa8fc0358fd5864c92e1
ze8128535bb7a9e577cd5f492ca327c88e93ad93f1a52a80446a8c50e13f7e167ea338d8cbc33a6
zc584cd0180162a4d93434b51c06c5ae1ed3a854f4969e691fc4866464409b5a3dc78f2f8766da7
z8039bd1ad6f0f662fcad32dc89a5b0bf418cd4dedec18da6bb75fcba4684343a755ef1a3978f20
zccf297e27d749da9d4e97eb2edc67565a520e68e9e20101e43d2c04075b8481e8e46aa96e08d8c
zecc7029e3ab650e02df1065ad30f8a305fe499c0f8ac9510369f78be19e261beba3f057f658a7e
z3ac12bf297ea6546a8a9b80b25ff211373bb6abef6029ca1cf69b6c194085f42591f46a3af1048
z81583acfa96d55b47d5e3afdd7cfea0583a9d536d219e0d1e62bb6b468fa6e4b6391066e5c3ac9
ze7217e8045e0be5ddf3046446724043105fa1ba75c1a33564f4ba8f09ef449bd2f8483057ad551
zafd9ee1dea17bc7ec9e2dba9f81ad4b3a0aef0d88ec46cdb365d0ad4bf8078cb63c160de974a39
z995e5e36851571a62cc1fdb96624acc6fb23b2eb71be3179db68956f04c276bbce7830b36f346c
z54d6e3e5c7a73b5dbfb0fe82484ed60c1f2761604fac686bcd88ec55d62691db6f01ee829ae215
z900c7b1db18e60f228d78782743be395768fb2a8c082d95f07873a36d233ead7801a6b29ab0be2
zd1953d0e5fb7127734d4300e9bff60426649520a1f4f177f549acfe43cfc91b744e7bcf159fe61
zb6b2eda84a7c3f2174d3a17ee73bbe6e995a3bd37d41a9325c447aa4dbade7924abd4619d370aa
zc561ad7bbc27c66e899aff5fe495d8b07095a41ffad1d30c0c8e2681ad812fdcb8c3c68add302e
z858b0038996ea0d50e63948d79dfeece9263284160021f51ae08025b4d33861cd45a8ce6f95574
z1b7a801ab79bd7a1a3d54d7abdec4f88495edbd24efed3d2cd364144c1bd3a5323f8accb2651b8
ze0e21ffc3168c5e77aa8d28e9063167c5bff09a572eb1bc538172a4a57b73f724ff11cab75585b
zc98e96d118261b2dc63da50e3ae5dbfc73128fe7f98e6e4ab5ebc074c690d74b521f464b8c35dd
zd7d9b3e82d99122fc25b8bf649e8f0d9d42354093ae1cb96081862ef59779912a5bca25bdede50
zd6050d3298619d01c152e5da0aa42fa7e17c741fc82a80576d06b5ab1cd9735906eace3d008cd3
z0b47f90e7b00c7bb3bd719f1a9b1fd4e198595f4743a17d56b0ae6a39d1ed820ece2ebc10467b3
z6337b599bf75c92d58e28f6ed3860c968039284dfa1b15987d206a5dba89ace56324462f36b64b
z267da1c9341e59fa334f68219550bc6012c7eb131e3097bb6376755fff70b7716f89f6653453cd
z5a0ffa55bed1113c20d8dc5f402d21f9c81dfe43a1d5685fa46fbfb16fba9383e4099d104a37f4
z670e653d7a78da2d7ff871a172768eef327fa830e2d7e520d54317f0743a44c0b21388b95d9c76
zb495597a1f681d4cc0af255e58f1781774204ee69c7a21f64bf4185f518861784015f894d911f8
z49950ec229084749e7670b161ccdc27fc560cd25a08fb48ee10832eeaccf06a1fb02ffd1d11a31
ze61eea345d9624f5bdd8725b6a6d3eb47c8c1c14338f9f1943fc2f72fc972d714bd8122ea5abb1
zcabda7eb68745d2e26eaa34a3c910bcc9f07fc45b832c2ba050ff89e857f9510946cbb2a74f8ed
z73c0f25cf7129faef671599a2896555f9eb140988d9bc1dd4e8b3a061a480edbf45fbcd034ba97
z6bd81be61540c718ef428f80db8592fbde43b484908573eec79504b790a9ae3fa0652845e0f487
zc75315a88bd85771f8038927a0af6b3c1e70ad52d10f4226fbddd49481e4d647f3724362e4ed99
z672747b0221fe6ae09a8d1a075a0e7683396a8fe90e37661d5f2d700b234d7a3cfd37308ca249c
zc23ffeeea927b0e46f0f7da28871ee9f43bafb639c17c91af7174385d280ac9504fc3d8b902a73
zdd87e5d7bf23b3c53d1dd7636a89c43f8d6da1f5320398012ae10b6f545086b6e6d05e89e38096
z79d2102f9c0451f97061d31758eae9824efcd6ddf54c887f4d878851a41c9bf3d3b03a8feac04a
zf8b27b7dbb743731a5a7862d2eb60732843eeb0c65309aeb5b1ca9cc28b946494aa84055cef9f6
ze40d4c44734013acaf5bf56a192bf0a4303ecff50b2e5a648e21d1cc2082e79f9ec1638564884a
z88183d0a77f8ed43ef659c9ce9542cd528e47f0d84c6aabaec7a31b944e5377af022942e14c333
zb28445492c94f8db060f625e9222b48efcac33397e26b2313e8a66ef673cf4b7b8938ec2a5d939
z2d99fe756da5d28d9874804d0bee922ceb9b8ef85c34772ebdeb8b149c2e5666d4a872878b38a9
zb68c65cf67ab163be068167881bca447827258a4b1540532abe3a341b9fd84ca49238d1fa0ffdb
zc5263a782372c576ad1f405b93a9691be868a6c7f100d3ed71b031da965d4f7d83ef09adc99298
z8c4a475cb4fd7e142b3260255260fed1e395a34b379a12a2fec3371097200925e4dfa1937ba112
z32596d2f9238501e5248a63d88915d1cee12f71bbf2a5c830d52fff2e4772757feb5659bb52f53
zaefb89ae6bb51f188415f2041562ec1c0f7929f216e141b7722d61e0fcba1230a38ccfd777ec4c
z7fa4e80d3d43fc748d5a83cafa5c131a491fde36cb659fcf98bb8e3a62918adf1c7a7e66018eaa
z9243a8c220f43bb61ca50cc4b089218ae1b496cb93fd0cfcf5f9fbb3fbba9f12d87ddd7a4b05b8
z958f17b908b069f9d1bf3e8c125a5f1aa0c16b8594711b1c16000801f5edb9a85a467f630dd231
z10aad562c440e3f3ef607a6fb948d1ffe752f49f596a8e07ce82ce3f2281ac79782880a6fe968b
zeaea66b41cc899e4f7a2136fa38db5cda6bee61eef4c486f4430f668f3ac0b0175391d4bd8c442
z4ac63003ffdb9ac307ad0a78e0596546cfd6a0932272779b5be4d3befafb7b9ad49910b3572531
zaa599405d031d5a5513a54cb79f5a333800bf0f9031c2930e2e2b15d63e47c77eae97ae8fc1f6c
za8224bf010505ce7aef6748fd1c795edb9335961e958cb3e81eaed505af252b5a4acd3f784bfa7
zaf4bfb14206d012b365f6d2665c75de50c3a30c7d99080de53dcc3ae1b5821d133aeee126bc7b1
z833bf56b18b9252f6b592d521e53d59fec2b81deed8d70539ef1b0b85999e304395bcee6196b5a
z8beaee42a0076fca13518498d5125643e6a185968dc6cf6f327c8700f93dbffa842f342aeeaacd
z0a4abcad35ad868aa420e3e85716d609312dd0a9cfa6b8565c4007d24b4f0886088d5c8f46806c
z82d1223ca32b42832d78f7278c2c5d58802467e6ccbd16654fe7febd491e1c1889e94d360f058b
z2ccfe0281934482af90ffb696edf54a5c838f747dd2508c2ba0e023dbcb5dcf4f469fce4ae3d13
zba6c76f724acc73d9043d5413efa022ae7c03601a0f4ba1a743cf3f2c4047de4b865ab31e0d243
zb18c888cb966330fc74d93dea4b04dd2ed56f444856a339086b0dffe0261407ec3b0ca34c3742d
z39a49cb49aee48a42bfba5a65736254733eff4ea1fa7f02c1209bbf660067da7e07a10b049bf85
zaedd1f8cae76a5dbe7c98be547e872aa4f84a666adc6324965e47f5e9e26244d277def191a1f5f
z668830be14f19dd39a27c7bfbc5f26206ac45ddb7974752719ab3a3e78dd481b76b055900a84a7
zd36efe7fe4b420895474789172f37af2a6e30c039fe7c9a41b88601989172950d12b09ab0d450d
zf20075506f1496720e43911c859fcaa945838b3b6b9ccc52ab2a562c6dfe33e088432b2460f32c
z63a8cfafb64edc1235bbd7481ee9601cf9e93d18d97452490b6640f6296e5bad702e2800b85426
z09cd5f878c0328cf217a2c168b592e39ff889f30b837f959bb01524bdd6fe0a8c9f68eca7012b4
z45db3e3563c03abaee4abda63d85c385a8583b439be0c238d0ef15a73e78ba2b90cbc3c30c1869
zdfb35be72cf328761be45f6a213a71eddf24bc74dc3779c37f239efc07485b3da8316e33ea211f
z3d62c288557f998b55048a413f873474ed907f96a2449e20a92a58083e0741d2a96515bd88dc00
zfe2d35e62b88cb5d10bda6d5ad454586b4c3e6c1967da4196686c73151a7977c0756966a8ff10f
z1e97bc3db2a69ba4260df5ec22cdffe1c4267674484573a8dda4857aaa7ec49e3114c24523c57b
z1374fe612b81e8965180c077f88aaf479a7eed91eacbaa93bd742ad52100ed36b9949cbeb14a9c
z4312333fea870d72d9a19c416c5c620d6de6676f1dc32f2667ff9cb946ddfeda536fd2044b1f63
zb6b6716b4cd28b3ece58a493d38992c149f0508468ec6d04c70bd331d8f2a148917692d822c71e
zf4f5450307bce746e227b6b9aa1adeaaa85f174a251676bde87900b4b2d42b6d9d3cbdd6f0d3c5
ze3e73b9c8d076cd48f494116f4f2202471e4ea03fe730c92ad1ba278041843973a37a012c79537
z8a705413f619dc09c02f189ec60477daeb2ad915735ec580e2e40391ba869199834b559df78973
zd612a4df4bda48c1bdc37c83d10047dc706201a68d36ec154299b53d130351d1164ea8bd70235f
z93db88e76effec346e1543ccae3ea1991ddf7d9cf8847db4ea608886b9c056ae15553c13a12b8f
zf7a867c01dc6a32d13f216ab3d5d5857d529d7b5984cecc7695248790048c41d69edd2fff666c0
z350d91ecb1d94ca5f560977588a0674ddacfb985d31daa9dbd08248e1e46c33ddaeaa28d451f6b
zcef87ca5f744da3b9394a5e5697b5b6cb9afe9730363bbc8bddc909538428b3079fba7a3283c3a
z783469e283ea4aa3aa5fd99723df262db84d05b8acc7dcd20aa862d9b59d3d47cdb5791d3c74f6
z7b7875f49c118b689b64237ff7fe15117cd9c8c817c90b904901ed6159c704a5911ac85fee3937
zcea59233cee8a5c7d64403d8848ff09c5c9fb8b1644af9332ba6e32a6f90af78afbc82768f93d5
z0a599dd77dd4e2b702f2f31f968248462f4750caf9f78cc0b3d70d2702432b1477fb315071d4ed
z0b0c84c92d3cc8c3dbf9fbd5799c1c3f730b21ec690a4754ffaf1f8a64015c9e62b3676b95f944
zab546f5ae7edf0594ec30a0556ac2006f92bf2012a17027d0f7fcfabf0eb0af4af4942f9100db0
z3633ff94178e6db42f4d6e4ee43cf226bde2c7c1b73e9b7177f48f42638dafb983c56f7d0144a6
zb701062f7fe0a565b84cfcd31c243b4f3854dffbfb7696642fd735a119b3dfcefc84d8ebe20109
zd65abe8fd8a4af6009eda0fbcf788ea861592f168079cc1a95d2fef38a88a2ed03b8d2a4819703
zcd3effec0e1f7d79f22d635f2a4381f732ecfae762207deefc2810311e47ab72932c87591653b1
zd4a507210afbec814010a107ad73e7d4a4c777a664715ee2945fbda21a839d66aa849388c5a212
z49fec8b06e8fafed1c9c126f2edd6652a50f1f6f3926a6e5098d24b47ab318edccb1b6fbdfc8e1
ze8fe22b45dd1d0a71f05242eab10de76eb7d5e7275274124de8ebd3818f9775460658f639123d1
z3320885c7a3e7d69cf588cc0254c74478dfa6cf019240c90292770e927fc417a1eee7f45005ea9
zeacd320c2e8b726bf4871ecdeba0b8bc6c758e3f5583805b44c66a6e2e89adbeeabf194c096b86
z6adcb221e6dd08b35c258e111c087a84e39cbd27ebeef01abb9ab1d48c672cad1848a7cc6e9e48
z6ed9ca2da347ef94eaaaefdf7aec408796d8a6d0b492f0e67eae927aed9cef85a4bfd49950c224
z246a59de3176f3c9e3e94076d809819e7f0cccab7f206bfd30964ac18ca4c051f0a8154849c905
z581e4dc4f68e3a6370a371fcadbb9d0006133d9293b8a02b91f14bd8103d9d1ab42de9ab492563
z4622e0334d4a38c49925391c77722021143f918f175c869bc9b9946f7e2d050bae8e151cb9a87d
z764bd033973284c04a1b580327e78deb8dc42fa4cf41b2b25404f314ce97a174aa0387777de879
zf9fe34fe1955798e2cbaa286e741101fdfe29eee103b6c1c044df7ee71447e46060fa22ca37087
zc44372715f196c7307507b345b1c9c0bdbfd8fa9fa22f1f778ffa1f713fac2a0dffcd69723bfe0
zc0520d1fd2ee7eceddae9e75d3313d44501f045bd039a934c1012cc4200b19a62dc8620a624dd0
zc96b5f691d7f54a0283ec67da99cd58a81fbca53b45c39c7ee0f749d138561efa5c6d8f6087c8d
za7fee6cece8f72b4a00c38789c97708a39d0845e245ace122a158a132140f832ff63f930480fa5
z21e9dabed43b0b4a1f95e9ca826e66071cc4a7e56ec5894d65fef19de40e4d48151752f620f64c
z1d4ef3041f8062273f8569a9f86dcd5459d49129a44ec42d783715adfbe877c553d3dd5af25502
z2fb51e06747028722bb3beba6e14f971baaef3446c7205226e8930b8e34f66d7e3f1d09c14f1e1
zece5dd2de2662e37439e14fecd742b29394790d145ccc34c3730140f1256cb5d6889b25e20595d
z8b4477efde3aba9c25c32c22f3a9fc91f9ba4e2aed6dc7a216f820c807e3040c2fb1313938f7db
z54f7fc0da4d1706151136e318c07d4a86cb191a16f7fc8261e139a0fd7c2abf10100ec410786bd
z174c7f5fc0eab8ae848887f2773427a67ca6dcb0d08d04de577c699e112164a4c2aa17ce5a02db
z84b1ecb6665429158af554af6bdbca120aba2eb43e74dcdf2423a568b0ba0737c9b22a04c2670b
za9c78bcfa961cb1333d58e7447ba76818b73344bde9830702c8c908d83a1afd9e28272370d5b0f
zca4ef34b3e2ce0a306e6b3a831ac40a700d711ca29ac2f54e89d07724241dc8251755e424a0e80
z1934bb2f225309ed634fcad0497cd5a2c5740717aa2b6053b19646d1876626d7cb1295c5a62931
z15f1202a1530152018fa44dbc42e50d9c27ec8c1b371e46cfff20a4aa203debf2c5b9d99d7ed90
z92a0f64c1c0cdf8484fe2407da3e73e9a6d96f0f44f2dd9737dab52fb2f7dc47aa716be7be9fc7
ze2e01e2be169118b1a69293bc0ed45185cf799969b3850c194258195f276acd4fe6778ec4149ce
zba933c3e2542c853f1beee4c6c910c43ba63066031f6f176163adc15478da70a4c6bb870de4c7c
zf1eebd2057ed3a0255a60902eb59d706b8c243e7921749b1618dfbd751f1f3d76b329790fe0cb4
zd3a07bc1b991a7088281c449b09e98a879ff4e971e8eb8494290dafff34abc20ee97ab17d9e79b
zfd3a7146a25b7fdaa7f1dd1f013df9b68e41912cf10ba812b17732ed18e843900a8ebc015d2659
z47d6cda27072b98f06d4d4c5d1b3bbeabf4e471620b05220649941bebcbe8554ee14bed25d433b
z2f662a90a00d1b59a6e9009c7dd9d1cab014f7f772dd011523d523a2716e3e2c375e5c86674f55
z893dfbb7d80c1794fa800a751c172e371044bb6812ecb3f5ef4ef9fb1247e53c68be71b0601966
zf2f5007b4f74915fd73d3c9775a8b9b742f3dfd9df1aec25c92b3dff61f456751f85e072b970d1
zb0f6cbd36a509d05fbdce3353b35f49a499107c4f7ecda2a3e5e1e5583d42240c48e93648f3002
z7f4ee3a9fa803ddaede1afe87093cc8a1ff389e8d1825b12a6e0f390f3de6f7de2043303c6f85c
zc16341b8017082f068e2d526e8aaf9dad8c237d3141910b78d7e765df572d5528fcfdb1756809a
zc577994679f04a97004d984784a20d0b4c76053a6031fd4c5f2304dd174883c2e98ba175b9d836
zb9ee468959d8b2ff326c2ff57a49aa0bf3e36aa808fcae65335c2e681f4842d8b53d8090600714
z09ee6634df0e94d30e579d0f8876c6b65b5e65537238d5a2bc567be3c8e8a9cb43892fb8b695f6
z4c14ffeba775fff5741f0ab714ca44901b7e9fc671ad60ee987e106c22c79b895fcf6cae23fe5f
z586f759f803c003218942a484cebc5288d75cbf259f1bb0cfeb8c747de3b78dac96d69600ec8fa
zc79e78040cc1fcf9666d60b93afafcc1b120205d12da85163e928f059b651ff7b93f4a35b3b4f4
zbe441b5820fe11a600eadb1c67a8f61c9fa948b761db006a4713cdd18b52e7ab5b620021d441c7
zb1e5b58303b4405e91196b3511bcab072ea36d5cc28122c82650a72dd46241bdd3100110d155ed
zc74eea9ba4d145eee944c46fae9a620cd2dab835a2a6adeed4d8d7ffac8533b1c0096d63071396
zd2ad0e42a9d5ac0ee429df3a38ee73e0428891c87b187e9525fe9b4d418794d127fd33790840ae
z0e8552f38fc74490147cf80b39fcb9348699f56872c9be239ab16943bdc90e1035d51e218cde70
za7f71f8e5a92c75f0026c8481bf0d312dd034edc8997a5e64f53b436b2d04f1a86f1cbe4dfecc4
z9f994d712a631a5345a9df86d72b8967f7550b5f8f88d573d5613c8a31b9b8af8959952abece27
z620c4e3faa8f836315c2492b3af37ae3c384e43ff9380dd7a44a2e7e716aa01749e0eae32e9b54
z802c624a44244f02e46338b61b58a157395676997be1dfa2a94ce81a4ab6a8977f417e603db1a6
z0fef691c0c9584e9e17b76aec2ff01c85508d2bb5fee42ff50c10f4e976e3b97fd6ce69cf353a0
zcf803b12e6671c2076b20585acd2cddb9b8c6b412d4873ff7a0702dc57df7c314957eadc55878b
z189d6546b3a5e171a7e4634fd3c84aea81daaaa3eab19b0a0b97a9306e693bee20cb324d47c25b
ze0f1b1c8cf52c78200cfe515e1eb13373bdb6096dee8b6a10b5041069992dd7d481ff9778d5fd2
za1b28134ff8dcc50b4ce1268c158d5d8aa54b9cdfa85aa95f4161132076a7dfd421ac7d8fe7397
z7f6bd79e7cd11416a3a56a3b768a39164e289096aacd365cc97a6a34c0371742b32fd8fbc9ff55
z7162c4fcddab352126540186b13dbee93328b118935976ac1e6fdc7d186c30e27c0d6d4be321fb
z45f7116b28762f0171f188c4dedde8fff76d4d7a7dba11f02053c796e30edb70e522f6e48e3944
z713d641fe6b6fb3174d8ab7f6ae9876ced5be90cbff37ce41c0645ea28655ed8d7d1adf81a714e
z4a948bbc09b18abc51e19d095a4a9a457fd97197c70b9525758809d9b5efdba4dd1d0f9ae32c64
z87d14fd07091fb6d026662394b82d05f523151e5e52248f121820a11d18836a814485fcf97ed39
z919ef7da0b4a01c429ff3b7c813b4c35f6c82ab3daff7974c6422b183c7e361b3320cd820cfc2e
z742015345337a354c56d51b591e86b917f04edb088c9d621905b0842ec0f912c827592af79dd0e
zbf13089da231d264fe0d8f4129ac1755ff8639f48986be32f8db67e2a58f049500afa92cf70832
z8b5195b9c7aa5a634ae82fa3a16ceae63053a99fd5a41089273bc3fdb8423e7217361ae6f87cf9
z41a14e216a850b106d0835414fba6233d8dc13178378850d64938ed65e444b64928cc42a54c73f
z893fd5423d9bbb11e707d686de673baf58e98c3668d6724b07dac1f6fcc266b72c275eae283f0d
z121100ec06c73df52be13d89a2525a0b914a334c7081a4140f625a5e92e1db29aa790914fd3457
z935e43a5b3f4b2ab5f8e63456b2bfad575f092b5ab0d25e6212af0d8aa11ae135252b183bcb178
z5f6a7582130879a233f1855b471d41dafdc8826876d5feae630cf8b4734fe53621a5123769b96d
z01f35fb9c1d4c1c9d94e215cb180b88732ccd85242208bc8844d27110499ab40fdc97de99aa309
z820d3d4591797678c7e2a4270cfce0e50a6e9a1240bb7bef72733c3b242e61f9a7ab59644220dc
z37b4ffad55941c46d991abeeaa1acd2af56529b76917820334f66666310bef4f88ca5547748feb
zdb0e863e21390559c570c5e9ef878019c49ad2123da1045aa442421dcb2cd77361d85216e12cd6
zb7d9c897b2d39e6c6f39d047d3de0b0209599178c5b3ced93110b46f66b05bca6130334ed72e16
z93a243e42ccf4f89b1a1caecd90b8a0584c4d5fc16312d51befd5e7c58a9a31fa7528ef8cdaa3b
z20124638d6baab3a22dea3b8b23ec9e8066230c581dc554c388c6cf84678679d110890f3312912
zc45cc0358178207d93f1b31e6235c574f55970fcddbd0b610f835e7ddfb92598ee9d10adc12a7d
z91f61ca01476c2ab417833f122fd7bad9535b36b813f338f0799d8142073a09dc3b2934cccca1f
za66732bc191b07d75de1dca208d131312f9f7338db7e6da9382e413537810917c143123c7e5f61
za6c4c004cf7a1e8c0fc27675d854c5fdbfdebc479e590444a4a8fcd390b2578ce8bf82ee22e3c7
z48b615908d7101d406a86e16d22e8daf78977850201ae25023e34ecd2c46374bbb0cda35bf4605
z43d7e9320793501a94fb8e1dcddd13af721e96d38a0c96b87cb99e0b3989e22d4f244c2ff4123b
z5c6cc18c020fe8ae0b25d53cb24ba317d50b912037f91be80f167c7cc197208b4695476f994be4
zea9402c7811b3d92e53f861c54b9ee94fe93f7dbb2ea84929aa06d346d9908f222e331f68521e1
z2b9e5eb4543ae118a15d8536071fff0c61feb8f1d665b5baf3d07ce1887d500c470df032a2c36c
zd67d61cebbd20f94a7b70dd67c3e1ad63a68d33604516b4b1f9c2fbe20c290300cd1b054b933f9
zf50771c1261e40ef9cd294dedbdf75fd85cad80ab3577147a2a81d45e076b65acbc9ef50b9d88b
z8d51ce12e79a570c8cd52d9f9489f5aee0ac889c822cfd6858b8ad544978432ae3b17b28562922
z032495fa0241957d7d7f7abec49a5ff65f3567461eaaa072d317a2356b0620669e7e716121e1b6
z94d7baba5a5cfba932304030060491dc017478170c24ecdc98c75ed1f6eeb15eef869980ef0337
z532d677cc7bed0621b134d53f39b42126483356f1af40d01b746f6bfa19eef2c1ed6ceeac88fb3
za138f2b98c8e0c059a3cf5fa86f183bf390de957436a6a2ffbcc3bfff97d8dd33f9389ee400ea4
z0d8fcc926cf4546dafff23208e093417ad98c8163957f323fee81fc7ca5d644bde59f02743c141
zd80487c4b39cf8bc03748ab70e7c13a535099789fee851af52ab617be019262f1fc15ee9445493
zbab6ac03ae78155abf3bb98da9d9f1d06eda587ccc68b69b5b01ec981d9af2fb9033875e389a95
z24668e5d94020de5a108692d270536919c93f63b34a37e494223f647396f437028c3890e6ba590
za268bd925d460a43912e1f6a3e6162839379efbbd37a962988defb06f227a48b95522b2bb14afd
z136732b956b30026d043ff13ce3795afb5547e511e68f2e18cca157075d5431821855f20b798bb
z76b4c46abe26dc314716b08465a0affe6771d4222313938ef87a04295366a607d62f108564fe98
zb51b513cc0e1c4dbccb3eaec163c7d1c55d3d9aa8a17198b3b0aaa33771527da2d119a31971d3b
z788d3ffcf617b247879468c81aa2832330d63ccc4d222f665d2e7a6ef2a384c3bf0a1d8642803d
z97c4bf655c4ae5d92b47bcd049976737cfa8ccfc67d791a45e40761a1797ccc4922001262cea5f
zffdfe10692f605f26c82f9a275a524b2a450c86a2296303e1f2197d89104c88beb73becf6838f0
z9224e2b309d973ed7cd51bc4d3b90717ec8bdef64cdb604e966d54793483fbc17a0b24852bb347
zeb082aab4631b57c41fab52df076a7d2d0618ed37970ac0186fc35c6f74a669e18b3ab03d8861d
zb00c1d4b1163d6555643363d2c2a24b68d374ab0af544753b72ada65a166943c30eaccb25314c4
zdc40f120291861d5c1d653058e03c4ce76c0a33a015f6ef859528b9a169860d4531cf15e37223e
zf06fa9eb1c7ed9d30034a72071d15983123c39c96a41047e3b696dbcf392e64682e511ec9b8697
z05a821d32cf61053296e03b2d4df980b2571c98b5cfd4a260a6872c4806d3febee180af862debc
z2dac46857f1b1eab084c3a4ea846cf22c032c561652d3f9464c58b4ea29a01c7964abfd0a80263
z1b2d0db6fd49851bb65488221b486ca5bb2492527016b6114a9f5ce4db83476179da14e9c4cdd7
z4b5f0b4a521fc21677da650825668679ef2353eae9a4667bd3f7d4cd087ebd657fd10f2fe4a1a6
z471202a148aff5576b949c3ec2f242bbb1de2103c734d8faa2dc15763baebcb4ce4ef047c075c7
z4a290f90b2568d3d2583bbb29426010389d4268359c1e00aa1c8fcb46a46b938f426540abc97ea
z5188c1ed42f0a6520292d221245945bf6631fd849f27ac89b01ae3eeef8d0f0ac874a0926c28d6
z859470bd0380720853340f5bf827ed12c0cbc91db026ee7df3a869a04a5df99d75e48406d9c0d5
zc3464504116dc689e9b4de1e36ada0628b9d1e27d33808e5c3fde68a67b6bd542953362f0485dd
z211f7c570da84d349cfdb0a87a2f6e61b2c221b3de240748cd50d2b212a0120441fb3a9bc7663f
z44dac7cd86aba307cc4d9432400a8288e9daacea6459e33fc338e42354b7d3fa39ef0287dac24e
zf0bc9ebd4d4e43548d302f21db6438d95c8063c71cb09345e18b1caef9732f80a89dd9c8ea2a04
z7871efeb90d3d7cb9ded994d9f7a5de334be93412c5a46955219a550608384e61a4b4d4960396a
ze1d7ac1b894d81a32973cd94464030202f81f5aadba2730c6043ee6dc9019e8d717affded31f1e
zbbd64bfddd291988d87c14912728c83ba7de8501349833b5305185e787a90182bee98a27f445dc
z005cab733ddc7ec782afced55e95a60bf65ac1056436056d3962e7c24298b8bae0ddcfd1879197
z0b8c58f0c2bc186d6522012d156032707969ceb14013ed06d230ebbbfdac5b94e48b7cd9dbfa43
z4e2db61bb026eba13faec31faa0fd15fe9676b5aa90a585c26910cff42c5952b7d534c09dbbc37
z4cf4dd53bf83e10b7b72ffdd95e496913a98d4136c466ceb55f3bb2c0b52dc43ed1b41585b032c
za97c413257310ecf419eb3e307a8228b7b9bd5d34c4e9afedae353801436f6f4e6404d433981d9
z74f5e3ea834856353a267c70f984b0339e3e4d955231eb9dd4d83c6cbd31e2ebcdea22b8b970a2
z4eaabaceb11c3163c180dc16ebd90cbf893134a023f18a44d83c0ea1e6fba717e1f245b580daa0
z86cc5901c717a21ccff4ef5e831dd19c23ce54d4c18b1b577ce609e44cb6b3aba51b41d9f2cafb
ze455d0748dfd991287954135de194e53e837fed2f0ee0aa49116ffae07c68e765a90bbf6b95916
z00bde93d48d24194fcd90fb71c5b1e839a140f7f1003c201496ea3ac5412a19c11268a9423e250
z9ea6ba94ed9bbeb6b9b4b5cfff5d6f25a8f39f2f0c8a336965862900e81a0740fc48cf072ab6b7
z2b058f2e10e0ea483cf74a68f19be12e6eef02cf190923b6fdf7da8c6ed781cd8147f0b6cd8324
z326f44beffd1ed0f9d332cc7dc850573f7500678e873aee55c571196893c1703ee44bedb503036
z54644f18e3807fafcf0714591b0b5fce44a1da3b6260698b236dec4ef02d122d4696d2d1ef6498
z08510a7a34d95c7f8f278bebeb7c57b7337114a1baa7433c012e365c3577ddd3a93ca2813764ff
z9d57a03f7243467d2602ac26ca7e78e3527f84ad20080a85b00f0fd1cd2c30f1813c4694b45e0f
zb1e60c7747a72aaa0c30091ab48198b0cf45b3a3234108203b68f20482ee89971305b10d77f3a3
zad9258d1cc7ea5802cecd26d247b855de3bbcb7700e2a659b19c3f3eb1ab6258411ef038c959be
zd423a07a61b0a9a4e8d4132c01042143b87b8b7002f722fb97e61b3923e878ff58f9fad455aebb
z993da79b90e8a9b65ffcf37846fb4d8635b54cb89656909e1a8f3ee706c8433ead0e6ee5ce9663
zc3178150a8896242c604367e6906587c7c403a02cc5c8e4b29a02c052df8a3d72f425433f8a171
z2c2bbc1c98dd2f82b313fd0e20ad7d5c3d5d3fe481ee884cd2882fe8fbb7435bd691b0ae3834dc
zddf005c6a93d3287e376491a2394fedadf7d71e2a28f7d5b84b4216c431280e5e00dc22921fb69
z777c0e6fc6e80b752fd6c419eb0dba12c6c837fdb081e97a413d6cbbc29e4a6bb7af226de33a89
zfb8fdf76d65daf29092aa8d29cfb73ac9271d3ec670b8012e9f84f095d2f4153483698459ba7b3
zbb107c8dab93ca7f3ea85bd657c223d590c1367ea6c737cbdc5756670a02de7c3f51617b2fee32
z3904b0d3082dfd0aaf15be7dc3f21901c7ad3b098b91722b599608a5f052e5cdb09a819cbfded7
zcbcdd14ce5a5ae7c51402b02580d7f04d0d1629554fdaa05769bd8c25bc040c05b70b13f6640af
zffefe35c9a45e89db313ac7ca81db5f90db55ffdb6df3e50fabad95f1b3af906d16ad45a0d0b16
z3012a841128ac6e97166652dd6b522ede10fd1d4f47de61973b3dae2f1ef7abb88cfabc16eab67
z0260c9ef49e02780fe2cc4b8f44d00a4324f69ba92edc09eb3a3c8bccbe1f713df0836c3ec5c12
z9997df2516328b67fd6be9f6492facb1c60aee7624e5fa4876b740e9db8941e2b58552d3635bed
z64b9c4bab82b3ea736b9ea3de9d1edea1edf372fdd357238147a2a3abb90ba783e32bdb9351729
z6131e023bc40bfa80289fda5454eb422d333851310c6d73550f64ce8f756a7de6ff047c3bf0cd1
zae26e0f23d4e1d1f0387f41bbc5fda6b6871ce2474d3269089621b949431c50f7c9a5d15660886
zf7f2bcfc5ced927b25a3ac494ede33e4c99750e0e8fe9070038e47cb070c04dacf122105b334d8
z5d122fca5a771428abb23331371990bfd909e05750179787c800f586688124848cbce9419ab70b
z515c0f71c6f20ea0ff333074b7aae73caa52f99948f9f249bf58a848384bc331f10889346a4956
zbf015d02fd08e024a5399e1dfeed0dca4217e91d7b4625d4b836e477cc235e9b13c45d1b27aeba
zb8451c73613c407267340d625f6da7216c539b72b38afaf6b81adffd515ce1821bdd567df39d98
z598e235570efad3a34fe37f9685c5b4083bc088e90eb634a1ebf37b977c3ed92662e9fa38d34f4
z9981c9939a3fa56b679e635d4d145c304b419359c075822409d9bff88aba83c7f967cf67a3b7c2
z84ab59124c28ef54cc1c5b79537f22e13079a050a25473bee362079d8bbf30887e87c8d9cf21be
zb0017164d1604bac4766b97500e25b052f78b67560c629a1628d816d67e1ee116079eb563f929b
zdf4093e59b2c09626e474cdf0dae1c0564836927f16bdbb588ab09c31f419590fa97d9fdde8f7f
z1ae73355f72379cb748a98fa442ff8bdfe3ae6170a0893ab7624eab7ff19cf1b91b264d86b7ba3
zca998257ed695727d7ad1cde69eebf2b551bfcf2ab12cbee3db0941087735b59b01ad03998ffbd
z3ded92b74ca1f2d0cec768e970dc6c5b89519fe1f9636c69b4b481efba7735be705fd1329c5c92
zea0886f9332ecde2d898091293a9161dc4340b585eecd7a58c258edc906811e4394dc183660162
za786d571deee3bfb8edba040e11191d3f0dad64f91f5cb40835328bbf0d213eff76a2e49d632fc
zd3bd5947c5ee99c2b9f1646a1398369d8882443f8e7029cecdc3404665ca998e24fa83aa7c7fba
z2ebfea476a6ce49a32a7227d2fe6f6f868531214bfc7eb90d391f49f34b78ec7094089e147c514
ze3400fa617313cd6af8d92899927abe01437efe137dca16865b92865fe5b338236d452abeeb861
z150d0339755da71a94e31185c036c26a19cfd7b333e3e19bf5c5d654f3117150bfbb5ebfa0c1e2
z2f7c40bf0ea22916ccc9a69a52507428de3e8cf5d54650d0fbcfeae93f98e9ca67ea8b49bae1e9
z90ed2741d872510b2ef4a0d7fe4e73d78ee1dff8e51a263b58ddc40b8386c7048b51fc6c9baed8
z6caead927f220c33b66df0ca8dd9d37974185282262cf5785ac5fd1dd2ac85534c6782f909116b
z03cce446f33ecca59daf9d445aa6bffef10083cb33dd05b14df6165617568b5debb76c593b1534
z1564ae2d1af088e85f3442272b2e59d82a76c8359512fd22e3c061f25c1c8116b4cd28ebecaec1
z02c36f99303a0e52a1629d67451747674e54d3600d016e8ca2884280eb5c6e1f2b199203fd1bfb
zadc93286480d9fe00a68440a052c96cd6ffb36469922e3f7b8d0cc1a5b13c660816eb9994443c3
zd6fed953e6cf3d580b2a8ee2ad833ba63bdca50d9326a0385daea7a205ca5845d6192292c2fbfc
z58c6f57b33ff0c99119bf56329926fab912ad6d06ed0831e5f1108437d112348ac654de3e0e101
z77e497819d1eaf9fb442f6f14b0fc5000db1b779be9a8cca2f367a8b7dd26bc2c1dd591726b977
ze5f5605559ec53553f544c93acb7fba3fdc98952f719070ba2e5872f4457043a2610edeadc3613
zaa2c7b64e5fe3d69432bb230db0c0741f90cb3e56abc87122dabe02fe2e871e5415e869c0956f3
zcd793b524dccae945a7c1d94829d3e068113f4d907227433f26f77e91b5eddf5b2e7dfc868137e
z62855b3303910e514710bf377b2dcd9da5733aec6c50b96a48ad83a8c3ed01010c348fba151840
z79316aa30d8239c9c6ddf0f4088cef384c6bf978ba7907ac55528f49e9710a066361264af24826
z5cb031f07d4db5f44b4fa68bf96cb476ae3dd70cf6aa19e0133e69b5c1bfc5f4059bf4f0525c5c
z1b815979194dc7d38e6b7921251d4c063d054c44893fc207ba18e608c4cd821984dfcfd961a120
z39c471cc0f412228c992cbaa84df872d3d01d4967812dcfd80ad7745db603f1d32b1da23eff76d
zc84aa6c2d193551265b56b53e8ad9b963221f0a4714e20832a932011a0748e34631bd3d4ff2386
z670d386f6d601accbc266555898801260e7648548a1ff7b790025ee67fbea02b6e6a46709a0f3a
zf4e833ff14f02e58bd90728deb88d156b6ce0df6b1585a420d48ad82373cce475aa0673610303f
za047cc9578ddc8916b99e303e5fbb043a94fbe3031ed7364026fd6be2e9a2811707174001ba79e
z8a3b37906a39188b130d4fcda4a67beaa1d72135c89a54d4ea99b5ceb1049a630539c9ea7d7049
z7f502b87454f15fe1c1e2f45a0386d64a7e922e746ab103be2488b862e439dbab5aebdde318b93
z2fa1e2c4130458adfed3576b441424b318b4084fcc4319617f060ebe1e835237411f410e37eb00
z1139dc4bac2fb75c8c2a00d1b5cb65ad0f9c8b4bae18f10483edf4e1dcad5077718a308148f960
z8c2bbbaf379d030aea611d9b3e1bd8c696c983a2b6e5b203d399b004a8a102b96b1f17c339f646
z7c00cb13542a0bc60deaec2eebb7ad220d736b73368466232af11433fd3e6c65d557a5a4327a04
zec6e6a758bd9d3bbeedc75a3befc10d23151de560513fcb764fd771259896bec7678d4ec5ab7dd
z8441adc6c98b0c431dcc235db20153b77011a2250ac617baaeda2d1e2a69a6c845c37a899bf83c
z67cea8eb9747723d7e8734ad86bfca7a8c743fe16e081bbcf490db5e794916a64473b703b84158
z143603f7e3e7bbbb92597fa6bc4a1cc0a3dce7cce226c88c3799ff09aaa131d39e6f77ad72f533
z271b9ea1c152ef6645420714c288d5018eb8edc382f47eb98dcc6833943c2a131d0cc357581e37
za4fec62e422dcbc3613dc3fbc77298930b037ddf39b337640c50a399f4069c405ee90a26165270
z93105a1c0a0a62ffce2c10edbfd7bf14c4f9b2ce53c819735b270992a8d0c3ca307324712d25f9
zab4eb2667eac6e2aaa9801b0044ff116a59990efdb6fbf1fd095575e3b0c578e131671a4f1ab71
z546e44c3117194632a85d025d4a15d12ddcf3d97f494221f5bf0740c7f18c6d175df63fe7d2bfc
zccfcc09c7e96b669feb014c45e1584e02c9b04f67a67c8b2bc4e5c4f8e28b6a93fb869a6a0d0ed
z93fef08569c94fd5573a73e7258c16851eccc0f476fb86dd475d1af7c4f8f425817f2d49d76cdb
z31584e519bda9c167ae4da66ebad41b651271dfa216cd27083a96b7483201e81427984e4cd69d5
zeedb09313f051d75c9e10e5ec220383feb1bcf0811d64c38a41747113132518aaa1bd92efb011d
ze408db88739cc53b3222b3f04085959d80d848a4038c752af08907b9bdbf0b7fa450c8f5e8959c
z2dfe8ce30d8ccdb41aa7447296f13034fbdd28c47f3b29827d3173cfd3fe4c79d1d0114ab53a9b
zd014dee94b2c8304db712bba9081c4d9b096578b65a1dd84f4381adeb81f27971b9b66268cfa34
zd75511d03412b5046ddd2ce825ddce770945c5b6ff872dd29cea6796186789607439fb104877a5
z78aca81c1b946f898578239219c7ee794388b2ad5bf99d1c75dcbd72279b289a12f63aa29c1bcd
zccd606412bdd6a6b968feb4c9165ccbb75af507affddf304a3b3b585ea0c48ff9b6318b0d1b8fb
z8b13979717c0adf66a2c615a8b43ccbeaafa556e1c9410aefbbdd135bbbb50f73a34ee0a5d2bd0
z4f23cc4b694d7ad01f18d1f2806918fc05dd0f23d234ca22476120847e81952b053fe51e9a84db
zbe431f2b3fadd35d27565dd500690e62994c6c26581711c22b43737e0d63725bad937ee1a84b50
z8510e18dbfa02277532285571104195ebabd53125b497a1459474f79fe76fadb9150c90ca85872
z12c2e3da1ad36539655dc19681837beed5dd06d0ca7b601d1cdc04c15fb6183b8a48d84d3d4900
zcdb8824079c98bd3ef4f8f4817f978c6b3f61bba4ff8e6122cbe7010f92e5e2221d11e5a1fe08e
z8c89222bd2c29e05ff0ebfab4760afc23908e3a21053a86255a29e4711d1e50eb36d74cb415728
zbe94e6b5a1491252a7c4ec7363728ac56817381ab9a639ec21c4187a18c22439c21ae88ef7ee27
zdae8050ba27a9e1beae2bc9ac869ef35ecea23dc5f2ffbcb10ea1379f3672a154d9e3e6b6fcd1d
z4ce7a48897dc343e23392c0f14609219e976f6789ea9ea1cf39376fd1136da724c2c56399aec70
zf3ddb8babcd19937cb5da8ad195723a99f62af95cd4bea78149c0fe82de050bfaba74c1d3fa5b4
z7340510f157d36b3c22e07d59a74c7d7a1cd444ab7d087a77ffcc7fac6e870733ae9a0cb7511e3
z9ed12c00892a547cd57628017df4ec4dc88959e4428a09f7dcff1574d3a78bb767b0d65b16aec8
z428d257cb925b3a742365ba39017287967c0e98c4011113bc06170eaf94ba4ddce6e62eabcb0b0
zbf38c3cad61d7a959886c3c7704a6b18c9a11e0f3ad07d34c3d1f3e15937bf49b76f2a38de4455
zdf2ce48d5fe4c19212c468246fe2c5dad3c93a2ddc47f4aaa32aa650a5f8e4875760d23490d7de
zcc1de31bca2378bdf9c101bc2fb49385fafe65c78715415c117a16a3fddfff39b6312fea465340
zdc77ed1f238e4c7331a85d3b3383e67f77e5f94f693e5e950ffc4e6fa9a1854d05a2edc5279a0d
z2f54e340bfb62a4f210df990098aa512bf08e52f864272f701231173732e683e1100ab85089d08
z2e6eb9fee2698b72a601e66bed2eb4692c55196c0b179257b9e23e9a426f951d0e905c8b6305c4
zf6c9d2b8b0f6cfa4e00487d433b74657f31f86d255204bb3184d7113ae2753b85a2e6ed2a34286
z550c7ed620c32e34233dd51f2ff075d3cd82f2d4cef8bc537a14f6f1b7e8f86e13acbf1b6bac3c
z98e5707fa84d561ee764549c9cf3ca961950d3b8ca41841631cd4f3b8a803a7feb26cd9ac228c5
zfa9212a50102b7b4e917e93ae3cead915b8d45e9a7bbf59a5d086d07e4bd724ee1f7a43eb1e682
z828989af297493dc6d41005f14b93487fe3c717828dccc77e3147eef55b37eee26a44f5ce3dc12
z491519f14d0670b66b4854ceedc11c8e6639dd3762de0e1c69fb180272a39301850839975ec60d
zebba4c793367de518accb48244b149cd8c2cafc6a121e79bf05b8970248ff92d5c50c94e337d11
z7baaee7c7d602676a168f2672310dd0534c09e2f8034302a3aad507cabc0e5a285f6a17b256637
zfd9addc139d4b3bce004d45088aee5277d3fdc715faa53931d5e04d1fbc4e10a9ad6f4a83aae3f
zee3fca2e57642e836452ca76aad678a334600d5dad361a3fcfab65e611bba9bfd0870ce7fe9e99
za09a291b02e03fe2880310169de799566d278b0046531e922dcf2d76335944583cbdabe844e1fa
zeaee30ef287aaf54fb09b8309bf0b738743a0829854c2efddead106aae9a916da05ee399b938a0
z50af4c26e1a834edfc667cb6ab30dd399ffa5f27695f970b0c8da1d1f4c1ec7a9b9a334228d5e5
z26c251a6cc7a1f8dcdb365140a9daca47c708bb017402c053efd348236316829ddd77470925388
z0be149d376198ea79b3e09bd1719164bc18e20617a90cba9e2cb9e46a94061afb533897ca14efd
zd039c68681e1057dab0217d67558cf7f27600d2bbd5c7bc431d808dbbcb0c1b1ecb6d7cd0aa1d4
zffd6260c1bcc8f396096e84a59ca2460a13c5ebf5fbc86e4183501887707c19259ff500cfc69ba
z8f59a3a90483bd9fea65ce42943c90e98e81f4082e270720ec8e5984324480de67580089443b76
z6464c90a97df613c7b8d382ddf8f2d42fe2e9078b4e960a834541721a41ec41aa3dba1eaa2e54c
z7275b4a24db0ad7fb6b7c6b24fc6625ad51dd2fbc6533f764b99aa16c28f72e3661469779457e1
z591ac66ae0a1df5f74ef31c4ca34ef5f5d561e5ef5509a64cab332dd259b1a34e20916e5f14aba
za129c170a6e6047d48d2106ea77e350f074b3e769de654b1d59a1c8c64995746e1e4d29f265bd8
zfcbd8ecf4b0e8521acc0849337cb542d8bd9315718d316cdb465b4d48e788d5f19e945d000d81c
z99c122e0ae2d25dead42db6a831a5ad56b173f37b2417646380d61dc35a3169bc120842dffb079
z7fda3c2620649ec0135321425e2d004cdd232203fa7eceecaab8540b35e17fbe5f521f432a5296
zd32dc075723484052dd5e4d9e6592560b46c646812d007437fbcb91b4f8656736a571d0e2d2179
z4e924bf26d0945f392ec44263937e25d9d9cdfac242f9af655fff514143239cd5ac112e488beef
z9139bb3479e374e526fcf096a4a03653151c39ea53405d537a86cac0fee3822df37c798b3b567b
z72680735191c2402cea3dd3e68bf22b909e784e3bbea58948b92bf406f3056085421eae081f4df
zd32a5dcffe8e5385b46a093a1628558c4a063a2aabdbfec9a10e7bef2a48fbecf0fcbc47bd8b77
z011e3f63cd1d7a433affab27e0cb827914f589937cb2167285ba608df31316a43e67a736ba3548
ze81f9a6c37b1dab29c4614690329110a57508a7b5116ce65128ab2a997a4f96469f146b4784764
z402b09bdb28ec93a6c93eb63ef1ba3e58ccbe7c89beab7f35fb7054600f497394c05e9d7445cfa
z2d6331a4edc79cce0a34ffb98f9c8a94fd8775ededbae9597b1b04334811b84cfa61caaad76ccf
z57c5f1546b75c19ba86345e466dc05a244de5cc25897e051c43695d4aa88c5f0408f711f412284
z413e33ca78c2c95860eec1445d00e3a711977bade8cd89fc57991c2288424672e36ab3f60d5eab
z72f0549b07dc415b896e8d0c0cb426a81e9c3005bd8c70688f32292c781b0f37dfaf93851c9457
zeda93e30f270d82559024b4c5f50b9d825b53d6c05a2bfb4fa47a21011aa69e3c0fdb74b5b5daf
z9fad4a7ed73073ebfeb79719116f7d1cfaf75eed32caee51c0bfbf44aca61e47ade8f715339780
z8d0e7ac8a1d9b1aadb2657b933e96097f5826caa54ae7ce76c4469cbd7f95619da6621e329c3c4
zb0845adebb0aab973cd9901fc23a77e00823ac7c9c014750206f53b78a498b212ada5d18907217
zd243f6486be65c1fee8fc067b3752841c327419ef1f21824662da9633af442090c8fb938786096
zba75a3a85a13b9cd31b62e38449fdb3cf664e1de94443693a2cf35707503e6cad48d8057a67e7f
z452d0d09dfc6bc119d0c5142eea1289fbb4d981321e99450106b2e4621ab4491b3328f2808b89d
z423f81a9d006cf35cfdb345352b45f4b36aec989223adf962dd11cc18a4d220b1328157474a3ed
z53bc5be0c6b6583c63a6f1ac1e4b1201ba2cf38e16581cff92c4ab69cd2ec800328b12ed1a17c0
z157136c0e62e128cf95c1915266224934c8905c8695897720c137c1ee7717f719f9e2e5e2e5abf
z6117fc2f9db7973e4a58007a4df8cd636dcf9169ffd9ae4b0304384ceac4658d4e7da377f10e1d
z768a1ecab635c269bce1570622410b178956427a0a5cfe74c64a21cb011f90361e02f56ea09948
zec33321a52d56de7fd2e15c2d7d6d7aa2532b810182b35a99b545c09395fb9861eb12abe8e403c
z727210ab0acb77aced31e21c2130c1eb69334f085fa0b8598efbc117351a108c38fbe5795f36fb
z81c53d9b011fd44b9246f34744fbfb5eaaad42e36d14016138ca1d364bf8f83ba0e1458031e645
z700aab60699e718a6527b70735f24436c675feb81eb5ef83a112850ea4e8bf6128fbde3ac9f722
z522a392b23d5eed848f5796ef36d98b06e4e72923cea8830c8fc4e8604c3d661b84dc3a694cf2e
z238affe296c6a0c346cf4c105d4cc32a3f90debfa70d3566a3b503df7594785c9bd8b092173e21
z9995f24707630101bcd5eb5c86078016f144f2cc9d792971e9922f0c7ff0d69e7f05cdbce4b184
z67700fc48a0074cfe4494142765cedb593b6304edcf8b565b88b987370dc2f594deece94b9209d
zd327778f24d6c1c268b80ff05a938c1dad153491bd1f974941a28d63dac7538b20c76cb9043c30
zd64ce6f5e6c141c9e23f60ba696806338e635023fd23f669e60984e26db73d646084e1ee2b8799
zae3816ad8b5655e09f665d150f60cfcca368aa85e001c5dc380794571d02f45f1e619ecbb1e411
z2be9e5a50e28b427cc09161bfaff1c14d25f6fa79ef6dcbc52bf52771d5fc28ff4149e33000af3
z5d55b9907005f0c6255829310984d6f2002c786f31a7fd5ca69de8e3da33db9702bc75bb180d14
z1578e4493839c0cc371b9fc33da2728f617b0f3573c6b827b62cb704fa0203a2164eb108f46fb6
z57e662bd72e61001361ec390c13086856081c0ac4ed3be03c884846ab6195283789b55e0f7d58b
zbd4a31b741eca50f955dbf12793271f07cedb420780f2d034d71a630d6440dc1f9aa02ec8dd6b6
z8f079432b0483ad65f6a7bd5d01d87bef36b9fbe48a63784934274e22565f2bb4c766746e78591
z5e235731568bbb0f3068efc0f1b7b6a99dbe478a94890684ff494d6d0504ba4785fcad24402713
zcd818aceab59bba124493df406cdacad5bf8ad292889dabc4a9a8a4ab2c172d564383147db48a6
z1f662d7559258befbd2c321b171344ed51fabbac7e936617a92767d8138a7e12709e61d5d202fe
ze7412fac42d5e77793c32c0caba230573100c4c7b3dc5b735b7cee724d88aeb42ee67d3a28d59c
zf7cb23a96dda598dbc6d732c882d738423c03e376b81a469b3a94717340225b7b68895d8f6a57f
z3d96c9cfaabf408bfca40b0b345892106b8f8a97466032a3baa8d7e0147374b17760bd8fba4091
z9cdeb2e6d49c7f1cd1c221c7ec1c322358697a7e3c2a88bb65c2262e8c43bfe006e7475fe9fe02
z646eccb2ca19145fc07bc1bb5ff7a1aaaf731fd5100bd7ee5ab18918f717ffad3aa92ccf10a320
z57a9d6459bfc292c2efbf0e4743be160109df0dada11889de4f0b18418c701fca5315af806553c
z57765b30d167e3e5c1ac4d590db84adf597b21b5ddd5e73a21757f252eca5e671b4c09bb4f8785
z5bf6aa11f53b4e74c55810a1fdbb9582fd66d4041df945575f315c5d4abfe32e34640a7ab5cb85
z516c71acc9741f5ac5352c4a4536ed76eb5acd7df6499a0366577f962cbd59d5849bab4376fd1c
z50b9bd17e1950d918dd4424609a259f4388d3e1a1c10fa89ed94d611f592fa1b2df3b1807093fa
zf679aa8fcc8db7558f3783f626712c56dc75f02b67cf30174a5b861609dff5a446af335b7864d5
z936b9cf7274423d2813695cc7ae24c53aa18bf7fe8a3682d75c31e0aacc771476abe792e35971d
z164fa0b79db4bf91b6e43aaad8cf6f94168a7c1a1289f30dfc419570cb98e69f30f80ed8fd843f
z8f8537f432d5d7c995898a75462a02c526b61ceb41570211ffd2fafbbf094fb7b02e77a368fdee
z1a344d8891dc55c720ba06ce62125140fad1ea3f288f3c91811c9c10b81311d94611dc197757e3
z0abc9b3ae1ae2f3992926fe788ca21957a2856f850b6321062c9e57c7074d5767a20bf92061026
z69a9aee412e6d65f3cff0c15c1907e1b647c2643bda937d48bceea9c1839fecffdafa1b7f1188d
z032b454bd1289726afd3024fe33c93a085b967ea3bfccdb9d1b684528ec8893df81be77c2eb261
z531543e029c6e649fe34770896170518a2a98ef1e21556fff50b2e2b0eff0e1962560f0ade0fe1
zde37ce1a1adac7e4cad3b5887e157d13fd794c2459cd622ea663a2eafc6bdbc60bdea00db7069e
z5cdbc42fdbbdfb646a2ce0965fd4fd5f1aa032253b3af44fcb9bd0728d2a083432b12d1d895937
z4fdc904e5ef0815e2f97fcec0ad8309e9aafaef7be8fab0813dda3c9adfd0907b949ca665c43d4
z4d827534d07ab69728cdb6a3e5b2ad5917c745210398baac17530340b96e9456fe42fefcc1e634
z7cd38c7ae531771ae7734535353cb8df197d3326ccbef540a77433536c89971840fd355df6afcb
zf377aaec5f4311e4f95eeef2f5698e34f3e24a831dff755053ab4fcdc542e1ec72f0b8df65e9f3
z507d11115d021a5eac7012e7987d7beb4d049cfe87ac67d5c0ed2bef08167ff5597597f468cf3e
z8f80f91760ba007695bf4c1e89d511e9b08b185b542c208a7b1761da12f770f9390b77c3710fb9
z7d3e910575b31feb6bbaed7e14f43ed6e87b486f093cd33c99ea51e77ee01d21f4c7cbe69180d6
z17af15325df15bbf5a5c98ee63c8e9eb924ebf05abcd918dbf3af986da11755944e16abf16ed3c
z1d99add6628cb762319522df5c241c5808ab3677c2b1f9f989cb606e129c3f413aebe6d57f6640
zf1b71e7d755d56f47d6c0ce680e3f9c9d31234fd08932d1742fbfa9bb6662603d1317746310e39
z55699a5fe823360be426902cdb1e1e53267c3e4af1d3e15dec5c29157fd37213983d376596a13c
zc4d9c345b33bd564b8a2168f2bb185bb0c018d1890d888140f76341c5b18f0da93d8c99356e32d
zab4401610decb6fcf03cc41691fba1537d6b8dc19c7a1a7e4deea612e16d1c4f23cd98050384c6
z6e304f0b51114cd3cfc8ecceefa71b592fe6793ed23c8ec1f9a4890b09fa9b11b63b612c2d1eff
z457960212b446a8cf45bdbe16d5018cb15be2d646311678ab052c5c9ba75a1dc4ce73c7e96d904
z74558c1d96526dddf2f20d0ebb14a82258c021525d698fa2201070db1e46e051ae0ce298701626
ze6e2fe9ee740650ccc11d7119b72bc25d08507aaaa47fbb92aa002c5ae83c91b3ad7ffbb744908
z295473574173abcae02aa75b12b220bbbf1a1ef6ffe07c6456bbd07499959b44ccf623b833e0f1
z2d1db30c36c6345b3f902cb3bc1cd90bf5dd41a3ffbc58f83bdc8030690c81d2921fa4dee89fb3
z3b861c44bdaa136f2be89b60ceab3b803ef1d70f51492f04b4da2bd7ca4df0c5644dbfe433d57e
z1045b4a0099f095081a1938c8f17eea202f038f671d45579d0c70650c59f8d91c63ba836c72871
z464135c7a8fe5c4275d5a5b0710e89c4dd98d13af0f5c59b40e06248767215997b886e6d0ba356
zfc2db6d9898d12a2344dbab1da5b4502031851e2754ce0f4197601a4b5ca04e091da81c33a9a0e
z8d74b38549c9c2c46ae0c0771ae16e2eff6c3716ab4af0dbdd4b12e7b6aa5878076cd51eb2492b
za37bbcdec0cb0ff1aef0cd680abcbda40cd201c898b6c70c7a0c8c2fc76b5c8f05b43daa5a65eb
z170c7b408caa8759d61ea29e44306b0228bc1e3b906e7b7a9f0d5e65460ecb7fc40c8702eee893
zfc19b5a0e01ad3501a372484ab5abc08b4fe7f0f12975068c5cecf9e86cf1479386d121c975faa
ze8c6c80e6a9dbd161435291d9388fd442565728910cc1be7639f815413459679010cee0d7cda3b
za3e5dbf4719e48447ac44b7e993ccd14df8cd7946393d4acdb399a1c1b266a2e4c8814001242fd
z9b438f5d4cf7950ae8bfeec670dcb03a454915f46b987c397ae920d4d3d13f87e0c75c487cc883
z76d74070aa789a00d78f368814abc1e5745713090b82e3ac35c9799b91b4d1989015038a988753
z9430064eeacfd58184cf5260e72b2889276c02a9fbee2afec090a68e3e064f280017cb9177a038
zebd2043a058cf9b27dfd148aae5b4c1106d614ed79450961d98fc97f73c62501dcaf04454266cb
z63fb0b790c1bd9b9756a96a0cbf6f3df7cdd01989201e6c25a9d11e72b6a19f9825a4b56c82ba1
zf4e81d93ef2fa73d41125de2f08380abe8e2b691a57d4ad8885e6dcb6178066035dc7af816cb7a
zd6a3953a45a7f2cc7d5e020d38fe1d716f2bc02c4827a7d1dc82c1de156c3585c002095880ee02
z909c9e77489f723cf6fabb92b2a1f2b1988b88d042f1ccafea1fcbaea99da5c41178e83eff38eb
ze0c6fe08c54e4005521d2f55a1fb0e9fd5febbce930a16f1275ea591029be682b5cfd2603acddf
z3c938c7421e4cee41a11016f7e0ee5deee1b2e36ae184cbc1f05d32e24aa2e123cd05036a4d172
zc27d1014388c15e4877554a59d4d42dd7d383a72396c2270003f38f14c145edd3947fa597548e8
zbdbe860512e4608278181f7ae6ec02613e2bba15cee2715eaf454ecfeb73efd1a90961e3b0ffde
z1527c3498f3fbeff471b8f5d42a907ba04535ac4d8ca1eaa7a618efc111514d7667c6624a301e1
zf03fa345c5aecf1b880df4f3ecd64201f72449d45692bcbb91a3d5ea29ff8d198683fa03a49517
z6890f94f0ac34c8a02e8035adad582149418f1fe3cbe772c7476f54779d035831c6f83f2a07cf5
z06a3ef6a3d4037e86ae9512152a2fe52cfb370fb50d7007834101063547c471408a69f304e8740
z7d240667d87e011938e9a5993127c0cdb62dc08009eabee626c85ab4ad6aa2818290a189f8ec2f
ze9f7e80e4c302988d7df9b0ae9487bf533059e82fdcff10d46295e885b81fcc88ba82b1a5dda22
z4698a366562c9ac29ee889ad88f78c705fefdb8484158c3df8e279b9c17c9c73a71338d6f52ae7
zcc1fe3271b3afa3c3c8f3828c7670f047286b261168ad447bd5ab091a2644563928a36429f662b
z694f1f28925589ee3384c1487005e098dbb5f8806a3c7d5b25bf66bdedb3d01b108dd45f29b912
zd09f28d7404e8092d7f4e2bb019016e4a67d1e7ef25e88f890ef1ea2699666371a173974d2442f
z3510ba1430b7ddc922d25a44fbe41899512b4cf2dcf96da1b261cd5b1f7e4e4a93066496d73e5d
z694654fc56f94a7e0b0f71dfadae0c5ad81fe7c3c5102735d1c5fd350c0094d6049dc8c47d64b1
z2e12fa9793f4f712e7cc81d56d2220c317119213a3543a2ef69ea043fd5f8e7e5e94acbae30e88
zf4a5c480452fab360fefe324075fbdb6e240ba15e3829311074db076acd99ce377952a1b96ef3b
z90cc8247e685643c04189e07ea133723cc26c03826a23f75c734303150ed8adf5e20e0effe351d
z16880b3b1752132b59f760d3735bcaa37c1141c637956cf87677efdf10ff38725952216ff510a4
z959b52faa39803884daade20b346b4c721ea08ead1907726adeda287e6b4b09ee88c68bb5f1f24
z1c37bf18aa5b1487f29289fc62dc1728a9eea2434fd4cffd0948740443b7bfa03850e306139ec6
zdd173e8562e887effa7edc37f25a1a349363fcf2d8695600491c1bc7bae675434cae403b9c66f2
zc02e4dfde14f91fcaefdd928349456352818de6a4e202f350dd98a3b53c27f60df751689870a2d
zf027ca459249408200bbcddff1518109909a4e9fa35e178bec128ca555f29c57a2f7b0f291ce2d
z49346ed11a48a73359af4e8da3c535976f2a6e723d7096a469e4052e3c1dcb5da263ecb1998b52
zcb95cd34b8ed62d41a0034f78d119f0a297d3a3396f4c522ab1463e66111419c46bdcedbc0ba3f
z33106a50e3939e9bdbdeaf14d8e1b8d69df9440099d7f2dcf3cac4962090e1bbf31f6653841125
z65dce0231cfd78bb58b3da6064959c4eb6b2659b589a556e623f6c90d9a285d5f281351b316573
z892bba9824326ee119f8d1f78be0c46952e2b4b92a152d9959650a021aaf2a30bd5d96cdb0bc3d
z1a5aa4b09454a748a380270dda7e986f29c8f255c81b199c50473dd86f715d946f3639e4725b9d
z0f1b637efa0fe382dce1e156cd33b0599fb0773c58c803fa535d681d0dd8b08b523d53ab7e4724
zca4d2b17eb0b3ba2bbefa56786f0587ab717e7a4fc1d333be187c0fb41d1f325c0629f4b637d11
z59186361c9d7cb003250553f946c9fa778cede256c4570f5b2fb38dee04b216afdfc39fc68ce47
zfe9fd509cf326f022aff8814ac4ac27e2b9cffa6f300f8f35d95220c8a6c3d18405f7d065b9baa
z96b7645c6f37c21114783c42f209b323167b5e6cf85e6d88d0c430aedd86023b272b49934c82d0
z5da7a2fc57306e3abc7bd0c28eb92673359e67fd2730a6a8c74d5fb96635e7214bc5a2682cb6bd
zcdf6b0da0e35b39b434f48d9683ca9db281db881b981111a4327fc20f34d420618acdbd3838ae9
z963d6876637003a7370e56f231d415bcc95234ce1e07c60a989ab50940690ab0a6fce15a607302
z6a96349a008a74fc9f969d1a943e8499d327242df0938e4f0790362a12e9e5a8645b364d7695c5
z0a7fb987b1541aafd8ee63a5e79ba6c74451cd5e9140fe1ac78be5adb0b72dcc2cf8b2ac9360a7
z00c58323389592bd44de55cf1c7f490cb1d6f4c5b14e1170374b86b72738ea78e0a7dec274b7bf
zf7623c85863268687ef9f30ce0aaa850d38d26365d08deb0284393e2d095f450c23a02750fd045
zba4961cf788898fc07a4a2100a6608ddaae09f2d72604c8a0abb5fec09c32068a73f6b35831ad0
zecf6ea615006d00954dc9ee51d1f41e622ae259f3b0daadb2da6bb98fe4a3c768a8f3eebeaeec5
z9bf109e800e79ee5981889d2e242a3800ba77b57f0962727abf150dea710b549a89d918f5c7e59
zf5f2c1304d3235c1c7812087dd9780df11a0b36875f39def7b7a4f982742a9ded342c1dcb91ead
z7f79082f6d6f898833eace0e2df3d678d516415e9892699ead601fe85bd412de32f8b0a25421f4
z87e95b9c6dcac73fb914f4886df7b829705ef1b8805938c6a0e1eb4c643021a1a4084b5a1b0ad9
zcbf3c285dad01cf5ff736b79f2044e6d1a48740a8ffc8d6305d71fa9c39fb51977c82831ef040e
z8ceb4e662a3fd938e533d22f36c2a87aef8fdc088c54dbc71979546e778779139526cc1ae70262
z3039d08f8eaafe391e270aa466292f927fe7f469e428dc1ce5c34165cb78896053ee3727eba51c
z97b146f5270c9a1d58686ae30e54b5cb7a69da63719215bfd3cfbfa24c160cd094cf8d802ba4ce
zb2be085a9ef6153c8f94024d00d22b160660f740cae3532a7ebdd993077369654998df8b7c57f3
z429cc0dabc66d7120eaedfaeeb7f207a8c9eb07b21bfc4bebbe4d03bab168bef1e9e6ab59f1b64
zb26caa273fc44aff944cb14bf9ef3b9b9a97a45c1d40fd5f87edc39e835caed8af16e9b6115072
z10eb23117fe32a9df8a1c41e3350192002babdb3b7a23278f46e1a43e3d0154112a9e4fb5632ee
zdc016e055085176a9cc1a60d8ebca51aeef6595e302c832f734588d041448158cd00ed078e6f2a
ze2c005b54771df08b2cc7493ebb12e75813536bbb0f209b4fa6015160bebb14d3548b808afe43d
zc620506427330c797c357c185df077fa719e08f0e85c0ad4f755251539f78b803a28f921882859
z58c3b796fcba5f7385438a57baf1a58bb9a557a0baa63d4943b6ddc2a16e083f8abfe7f86d34bb
zfb46960ec59c560bcfc467f8470528417975704e15a8b341256fd30f07ef2e744abb344c8f205b
z0daaad7e7ff5d3f5380e1a9701e5097f6627484c1d671496f24ed9b9830d254af34839458ef5be
z2aeeabbd19004666239cb8ee523eff7aff8d8eeced10568d37d67476bd2c5a9d860f30a91917d3
zeabc22a5a6e71d605997356127312e10ba3a219df5127d3cfd0c134584414b4ffdb9071c9bf5ff
z54fabee966e6c8eae104581c6777618f8907d2c394889055c3fddad0bcdcbd9c401eff064f6b29
z97a4f25e96d907262e08b0e4171371d6d40381bfa08bdde01ca7a4efb63f04afbe900997602717
z94701eee499b42a99125883225d15c836fdcaf65258f942ef69dd9029e4757583af0ef93fb30d5
zaa1edbd6616c2baf9217aef0f402ff6de4c9f4c9b10bce7f260a923488850e3c90beae6df95bb0
z460c1c489881ee49e1b5b0512bdc3211cfc50adbf8dcf9563a89fa4322d9f0ba3dec0524c7f155
z4408d401ce7faa370657f89b6189a84c7a90056a127c9a0e442ae7f4a8ad2e9481ee9fcc015f6e
z22dab6d4c4213d13dcd0dd1f82fe3ec3cf4f993e6370f3a777e00971ee40fed383e2a2f6a17eba
z72196ca3845a3539e516f29d4b6912fe6f44f9c14622de82cf77f06ebfcd7ae5a0c2ad43f7decf
z436c0a93c922b46078ced4d9d9ac7740748ecfa524710be4f988d9f900a17ca769ec71869a38b1
z19e4c4049452127cea53f66d49d7ba94bb43c013ea53ee0d542f0f180fdf3218641f82f0273f6d
zfc2f00baa28f8885c3d7e723ad389382575b12b825b0b8beb1b952996c829741b9dab39e1a2765
z3f5a61e002b42dc87b6e8b2c329fdcef1e012ce4d653f9ab1e047458c8cffdf0275a2f112b22b9
z01dbbc0aa3c31ca6030751d925b4525231932842aea9c9b32bde7a20213a88ef370477033800b7
z3e6b5fa66cd124209747bc901698b9ac5ef2f1c5beedee71cf33c80dd18ece65015d36f60b2da1
z3ba970fc020e5f4c3319649da92231e957c8591633a99da2b75926bc27b3dc6447c6c261d7d504
z938e12782979feed18039ae6a678993fd18b9e1db0d1f2aeefc8ddfb72f6d836ceb12ddbb2ed8a
zb5bc52f17500f302514075708773b41eee08420608d4578f9b5a6cd535d9d6095296606b5380e8
z5dd34184e789482f19f14c2e23c5fe94a353e0627115eb8f67ee9f2a7dced9b8b434605fc254a0
z065ccff5aa84cfd95641fcb58739d4ec84d6bbcb70c7b6ef5524d4f7761d73f6748078d561b11f
z5b27613472eefd3e16b0923dbc8703e86426813792d64aaa4ab66dbe7f1ba19ec3ceaf613e225c
ze5be25a6d085f70faf99a5f393e1f0b8de1fa98222d280e393ca96dab609e17cd45bce18bdc356
z851c8d17e408ed554a68416c993ec3470b40dcd94f5255e5adb07e7105da70ca3f3fb2184851d3
z3e4003a2648672d70129e6e092ea9af1d9a2acef3454ef8041d0881d6980b518df2a2ea80059c4
zce311d8b5e96817731ebd7fbd053948e357694c204a5c4fa203b975974d0ab69a37226eac074d3
zc370c79847edf433b021d5cd599332872cb3c4868e31b9d555a52f1d4db0a3945a21f5388701dc
z0a9391bfa0ff4a451b01af9698e04465111a43a05ed2a9ef0e7acbf12f809cdbdb814052e81000
z7d7dcb7b34fddefa1143593ff3b87924723da78c05939cbc64ecccc3665d446f449b881ddce66b
zb6b5f0b2af9d026b89cc17395a306409a77d24c4e47217be979001f0c95e7b316ad399f5a08bfc
zf4cbf71a7854ea22ebabb751d313b4731bad9c0e5f9b45d37309b7d186e69ed854b4058208269b
z13fda0baa1a291b41bdb2403f92fdc79b1306765b60c40138d2d46f464205c14ac8265e3ae39a1
z0f956173449717c406ed0dd9dd27f80601b17c1f9a9a1192aaa6c3e9a429d8f631a962ec0720a3
zb29465772d42dc041a9c051341fe01d19f04cbb144238d0ab6c1db6c376969431af3bda598affd
z15870d019cf04ef334620970d150d3b76d0a961c917bf745d90040b38be7460e44701e067f677f
z484df757b22437b9bf12ea7e1b8cf5f0b6a0aa4561b1b03ed30fe7a9889387c9a4e1ba4c752d37
z2f8a180d650331249296f9d0209b609c865e7a4b49b310f3344f4574b3d61ce43aa88ad71d5dc0
z8bb957cd3d3181d2158d54c4e0ea60b06e9b03052b7fe8e13c51759e0d0a50eba65624ccfd2d8d
z2a1e08c1abe34e054c261958da8f7c6ac5f81e72cfe85a5d1c4a145a4b4b62547b4d31381b6906
zb8cff1eaa2bb1d286462262ab168a9feca8cde9c04d39a1173c40cb4682ee8ca3fff210045aaac
z95c822c943b210304e66ffdde8cda134e32f6c8d5180c200d63041019ca54b4774a662c57a3628
za8029956808bee67b83b7e846b93353f161ac8a0b1de111b23e2298e85eeef73dd2721a1fa0f4a
z66ac8622989a67d0dae85a6588651f047ce7134e963644b9a4cb0e68ea94ed6b15b01aec12a63e
ze109abcc39acd783f9ef0bf3b52b94f8b62becb57aa1c731eb8f0ad409ba682a54d6946c240098
zeefcf4323084c49174150db7e48bca6fc266479341a1cbfe97eed9442a52e563812624f71d396b
zf817e67ccb56108a6abc2aea244d094413228b2ec9b600e7a0d5e798aedb3cdf72695d33cd1467
zb599e6c053bd54a93608ca84b1ce57d39490f56438599e3731e29ca8f704958b4c9d28ef6460a5
zf19d656ff23887952a5a780834a7b09b1e9654915bc1d1b7d28361066cd889aaac0ac868166c80
z05b84aadca8a736f65a04af899d98a6a26def23ebdc0a582cfeab3d78ba94ff6fe34200d0fc13d
z54c0160e78c80922a761306f70be4ef323c214133ae75a971d9d098a87ad826835bdfb32b2ceab
z7f7975b65d351165d04ac5fe84779d740ce3ed29b1d79feee47c4ad5bc441f1089d794564c3cb3
z2a4be5dea03451322e2155f7ba98847301ec2a3c64ca13c85f9c9a65b100c613765813c50f2c51
zaaf10322e4b37fa2f1f29f37568553e437988f5ed9f9224374dca11a7c9c6b027dc878265be2cd
za3135a6edae344525d4e070f345724bbe2a3fbef6ced85e2fdcef3406c2ee65abfcd228d1ec7bb
z622598c457706c6bc32cfa999d30a76a2312e4548808ea3a5b76fcd3e928240aad8a996bccd744
z0c594f155717889bf5f5d14f3a06f7349a4fc428981fcfb38be69997e68d74cbd602f34e3df0d0
z041ed334c7c3a8579a5ee47f66e9fdbbe82c99fe3611cef6bc5dcf7bcd5b90c5f17181b51c67df
z949833763ae6f57ff304f9c5dceceec48a4e1d6dec26cc5463eb63fed708c471dec736561c93c7
ze3f528a281f8ddb709b94242c2ddff73f6bc007743196b637ae3e5a37e205d1eae2d68d3c78cfa
z99ce29cec11499293843147431e795f8dcc04c4886ada2273f7dbf0f3b00aaf1cf1894c62fee92
z03904b6c119ec46fbc1d0cdcc5dbb5cc4639842fb4d3ee5739cca54d15c215fa0a1795bba4bffe
z814207423193a5eef8ff0092fc946e1abb0020b71336893a2919e8c5c6e3036948fe0857cde4be
z3ea3f37fca1d0ba1378b29db4c4286a2fc71a3a2700947039ae88686d105aeba6492e6ac393679
z3ad82d8157611da9e00613c198bc52e30fe6eba73346bc1e2a78eb3e89f74d1444a345469fb67b
zdb3129f68c9b19d7621d7b89343456a1ed919ae244abefc65bc2c40a31dd1397350589555411e6
z904f5ecdcfa0d4df4b8239b23eae8c0fd8cbfd918033300936e9c1fc04a63906cf5805fde02dde
zd1bb1b41fd854c0023f55e825ae193debcf916abed2c751077278e522cca82f9fd188e5e177431
z4ec56081ad7fab999afc27872867d78564f0a5c0632e55b4817cebb6c68a596335e0bfa9fae264
za2a018e02d8e9f57c4eb40ab287a78eee60982a3ba70ce71ef53422b815ff5ba40966a45ba5e44
zb4867d1b4aafc9c04eca510a9383467f7c1b51a810ef56094b84891480cbc8020cf128fb382aec
ze1ced4efccbdcde4a2a13e5491fbd5cbbd75fb1afa67cca4c6256fc200bf6695fd79367130a942
za07b11ae019dc4b60f136888f81aa001bb755a0357681e7b785afcd825e4960717746324d8d66f
za54ee72fa4ea072daacc3ba70055d447b41bb15898fbbcf0e8e32da3402cad78ddc6f3c6fcfa91
z9a4820ca090c289045a1cfa8c9a03589a2f86f1d25d377d0a1aacd0765a55739dfae76123e652c
z7be6bc6a26275748a9c80d5f4138506c53ba00588643b75e7a9a243ca722ba93e715d385805b20
z04512fa828da670b44c2eaa3cdcf7a63f9e32ad1478c00aee26c15864d1eb5ef6e87791eea5d29
zc0f75c5cb43f0c7a6a3699ca512113cfd86df5511a26b84ba2101d95d5b7f584024369249a140b
z5e7cb9aaac3d791995b72491a36209692b50db46f5a37b06a716fd3ba9773c1cc4106fe64842dc
z1a7f70f3c6100c7d0ef2c090e627ba737cc8b802ebd64b215a0b09fe482bd545699b52f29d672e
zaf52b6367594a5edbc6e615fab8d2c3ead28807a4b3d8d1a24ce2820ea11593db0403e4c67b3ff
z81d4df63f838b1e9ed83d7e53f01c0d19174b2834f0a877d25c35f9bd6add1cfcc4beb901a8dfe
z2a0aeda211fb282e47a23e44ba54afbd20644c92f9b736b9256fa8a351263fc432e4cec339dc48
z9488090d8be69860f300cc4be4639fdef39e814d12cc61159a1f84763d69620eb6faf4eff8c334
zee8cd565983ef51d69fff267be8a10a52b79ff35d0f6e917832a9d02d652ea90b17a4321b7b87c
z26f2cff83dd02efae31a1872a0ece72f64d728a58a882e083621709301c6e4c79063dab956cbd4
z6a407435402aee97f8c358682cb3a6bc6f82015e1d84b6311d49105d8935ee0438ca54a0437efa
zceeeaf323efa92aca28afdcbc68abeff294c6a149c3918193365a994a09fcb38e0f5bd9529901f
z96072c88e28ea838796d1b549899a31feb2516e63c33e764be83622d68a7ed9b356523706b8ef7
z618b76c65d6c1fa9d0923cc6f2a04608f510d93f7ff055cb08518ac639cf38a927e8fe0ae7b210
zfcf4e57af4f8ebcbae3821772c9677079782c0806e7b84518558713745e6030821490b07ceef5c
zfcbd9e47368ee6c308ea4b2598d885d01b2d5285f0d7ab81a8178596a36a9ff8640da7164fdc8b
za2fb34fc28948f4c0e99fb33e5976c8cf618b37e4c4153a35074f5ccd6c52a20d59e9bbe955699
zd6e757741abef59881f1432239f006d01fbc97c61b57b7825ee372537f0f5c84605d2d40647120
zb6b27b18f33b7528d31d87357378cd9ea4fbb90a97b36217f688b3a357dc37f5d9cccd5edf7a64
z1d097faa3cb7d2d975ea721c53768ac1e16bcd46c633640d04b4b2aecbe78e5246b6a72deaf054
z1f22839a24be8a9f600dbf121bf1989a58575075ca15bec4c54b2a448f4c7446fbd1b44fe52064
zfe4c6ca833c8a59be3a8dca61b8c06194ec771fd79363e8b27223df7413731a88cba14d8da7f48
z3beab42764d89d5dc967d5a1fa272a8b0dd8293ea4bae500f80d8627bf418fe341718474bb1e2e
zf35f2cbac587338d64aff8aaac908a3188e831cf69f84519d63f32b760247bb7132ff69eff6226
z4972fe5ec3f548d9cb4f742f2cdc92475b0ec19ee3259437bb8137eb6c19ff0bb1c19f9d7a2a57
zf52edaa53814c815e02686dd5156244716621889aa4e08329e48e5d1c6fa11a384290c99b070ed
za16d237f0cd28e13a945979fc8d77b63e2292545b5e29ca2e9ed63f3b1e90da61d003cefc11aa7
z327c0da3c152f19d369eb46173b5b9f2e4375b79d890ff8eadfab6e20bade52853a779ea778155
zd694d94940dd86ccea0c667202fb583fb4c49da400dcfd1471223059f0a3506b869e396087919e
z0f1a9fc60fa4598a553614c489cf21152a7d93e65a1ab686794858f7099dafc90227aec4e828f6
z61064cfbb48e3f7be37ffe3d00e333149b49ec5b5f40439db34cbac54fce8893bcfd5eda5d8574
za5dca6cbd182739fa079f73e727a32dc1fffe788da98ed157e34b338845fdf457ae4266350a72b
z624902b9fb8e3f60e58e40ed01b6056cd00056c20b1801ad912a7a1bbfa3cec23b807e7aa2ddb5
z001322a55034ea124d2cdbe55338000b47e2afde07b553b726bc1fb5d4ec12995002bf1805d674
z5326033a54d047db4935cf59f30febdf41818f4e8e6d9a18ccc747c2a6878e289bac6b1b01251c
z268ff9f0f491a7eec8be02ff0c621f9a46c6c00a875229044285da9de51a1d8d47a7d776e03aaa
z5cfbff6ddf5f6a8c838c8e281084704766aeb1d3d351d4cabbe9f41eac0126eba0af9946a62b7b
z3df775150da76625979479e24cd4137779db17bf53bc2536b6f2720f34aef146d478e12c206ed2
zda12e28d3a4dd81445aa9f6b75244db3398fac12dc64554bae9599e2384bee1fa44c0b39ee6bdf
z12411b27604c410280b5591d26152bb30f22b83f893e5a62429be57bf28f05e79bfce1197a7630
zd27b089657023ccf5315da1db3716f1a68e471c4719e664251e48447620c6d6620b7578545e485
z813aebca238c84ba0c40c12621fbc74e6e98a6e5b6819017d82cb1002b8991be687a144f772792
zf422a78b603f217dc8c8a3dd0179674bafe94e7b9332df6e49ccd5267a1851e3902a4d20ac50e9
zb6b75f9b08c0d7dd291e9dc1dba4dff3e6aeda12c0833e2a66244b6d1b434c58b798631d8aba56
z42b6fe847ed5a1e5e0fdcb183120dcd0fcbaa047a5f14f96ec258cbb055281469d91b11576c81d
z72ef29feeb7f0429adc596883920a80eec8b9cfea135c5f20c684ec7b1b4fd67a6e70b1b36b00a
z933448e4c75a61cfd7039f7b8c3f24912bdd0a037e92e4ae90780de91575bc61f0be57d53d8252
zdd3f7a1d2448d2156953ab097ea63ec06c9fb6a2f7bb59c256461dc4d99cdea5227649682fab8d
z0e5a87d7135accceebbdf6a6fc7c99d5c78bd5c9b656568c42f459e8bedada08d525475cffb59e
z9cffdbb5d754150625b0876b89a7590d1f891e5bb96d416f60708949dff3783afeb0f8095bfdc8
zb2812b18c94cab0a2d746311572c2cfacc7ea58d5ae098e99bc82322026fa4ab3889f3445682ac
zff5269566c96601694b0c032e53b71b6e133c9a6258760bfe25ec5904752cca656532e6809563a
z20e60a991785a3e1cac1ff06e2922cc78c17c3b50f05b138ca1c68af7bdc4e062875e3307d4996
za839fefc51aa6283c231c1f652526b9e5b7a1fd7907dfafdb4272450f4ab9919a50c5887e78cd7
zac4e5344c6dedc67c6d47869420ce6027b09f21e6d74821ef8b779f379ccdb11928aefb5edd9b0
z63126f3b9c2685b6999068c12d08c493cfc3b347e1e6417f86d21150e2f48b35c35912139917b1
z384ca57b5d9dc6d2178998d9c9c94c2ae0dfe1a79f76d66cc5a1e6cc4296690a7a1bbdf29dc1fe
zb1a250b55be7086ae04a709f836f11e545821f403a7b4f36ac17828c38dabf62b5aca545ec949d
zd065efc472b1b2f7484494dbb941397e5de4b7621e622dfa58a8615c283d91e9285e8bb4f17e6c
z662bfd8bbe8a5aeeb676ca05df186f49266802ce8f451543bae15b814616ec6661365f08d170a0
z8732cfedff83ec3db6222bb629e5cb563986752a025280fb4c55d8831746e25990efc3a6114dee
z4fe25a0eb75bc4494cb6d1b3eb23aa12c548503e68704c14f49dbc66365022c3551bca1da89bb7
z5d6ab4bda862f6752f4959e9daaf5b2b3f020f960ad4ad9fb5911b2758be62ad17965229bb7212
z3f6f10c05ca8f112456f9c27c0fd94c1aa2856f78341eb9f6df5f01bc3caad178d3c04bef6359f
zc5ac7833c2f09ee48af4a9e421997a8bc255e12f3ac7a7fc299bc2c6d1ac1042b81f5a6ce1126d
zb217463ad96b2de1dc61def914be9dffdab90c7401f3713e7b814c61a5cdd8f708093995f36d76
z4b13bbacc2704f8a03b4212e67df6eafa3fbe8107d53ec74acbd3c7ae3992b7b1ccbcccc80d7c4
z7893f14f9b93c1cc0a7296f4a2dab6f4097b89a51940a6dbd0955f1b5c9e83269dc476435a8d61
z4cf8bc95f9b83c009691d0a92ebee6329fb07e9d41f1be3316bc4ba0b279a3dc992caab32b3be1
z0e93f13c538d396ebd56b3a6aa9c12d610c1ddec0ce1f8819a99ddbdbfd027e77ab3470397ab71
z4bf335568b77311ec6cfe531664e87e1be880b53fa151c914ead0d8f0767f9db754f234f4f31f3
z61373ecdf89af02f85a46d9f6403983505fb7747afbb3a6b882d45a6998cda05585d8eaa631e9f
z8b574e6f9b93f84f9e3fc429ece870b1f50455de8715bb7451d0039b91a4b7a0cf055643a55b2a
za305ea0ca97c70788b554d2e9d2ad526f3fad5ce1dfb518e948177c63c66ccfa84b05903ca46fc
z859576e0a27d3ffca66a0e00d91cada4c266cfe040fe47c9a8325613b62c14a1fa90559d284052
z02b4f1c0a080df6b71e62da60d745069064fcd73651641546e1cf317f87837c6036b7ccf083c2f
z7d50aaabf6415c6b22cd23630481d54378c5ce98d70a347d311249bee386104b5d1d67aa5f6a8e
z65a24ef1e851312e46555756b34698fd3915f96271a1480c1f1fdc66b6d4a54bbdd36ddb1d906a
ze21c1aa75464d9cda7f8000365b42454db95b51c7f346c0581ad7025580624fe9d8953bc830416
zba0d1612bf3731e73f8561b0bf679d6ee046fd858b5f7c7ae653fda15a2ae154f87c9cdb7d1cf1
z10e60fa0b8f3778f7e3d5d14227aa8873cf53bd16dc78e72e1f8d945cf694ac77f99016ed55768
z15d28441badab31b14b6c126271307a2c0a879734f0a94c05708da103cfa5c2687d9b52a31ab5d
zb635e3c7b72d8cf9d1ac1f02234c8349ea91d4b131268fb045aba07177e3997f18b52a42ff56e9
zeaf9cd7feb5cbbed1dff51ce961597de34039e6c3633dfb9925e5e0ad0e3f70b497da9d711303c
zfcbedfb0f950504b30c46d7950c1551eef5a561307281de2592be21d10a66cd195a61ff1c7a336
zf59ea525dcb7370604edb097e832bdcacf01cb9018915bc5aeac025779d3e157f67c3eedc3c6c2
z044d014751bb4265a5b05658dc66f8732014dff1b58d11be576aa0ea0b7a326736410c0138efd1
z55345aa634d3745e0123df31f71d9a0b3980f0a16d1f2d8133c65bf0c99e96469c381244f9d80d
zf8026bb72e80c8d73cf6c6ebc72d60237a72480d7393e16174d9adc31bc422a900c0767eef8c58
zf8793d499c16e378ac74beec4bb599e6d6d3f07257d23d70ecab15d115241ec9c8087f64875e06
z82ca66e1bee2c2123f8925fa7119da416e2876da7e8eefd58a96f546538bf48f2fceeb53c58bd6
z0511f96b7d4d88714118067bf54e9387ec56317116bf7842894dc0192b5697dcd8dcc351c0b6b8
z744ed47d1500f7fb229ad1e4b7f760faa12910715ead46582f34f9a4a116204296b218fbfbeca9
z1c5c3d68d81452764d67c21ddd6675eaec5176c30e3ffecfdcd63d9758894e0d08affacf2409ad
z0aa109219977cfc43fbee8bb4942037de19bf3e5f72741e69bfa27009ee4e91319a2a9367a3a5a
zfb5e008aba2364b8a5376e887feb2b9173d897bebd642e26c45728c65a7d61896e363ca723bef8
z635ce4345671a53de9a7596ab25610db4a74284d23335d42e5f85bac5ba9edc4dbfc51b91bcf3d
zf94a76eab5d3597c2a881c76495c9d1c800e2ab62829959c0b21156c9376207dcd4dcb27047a2c
zc36278344cd197b0a85522d6e4bc79718d2a78ce44e2c878c1615556dcb6b42bb0d1a10cb492ab
z8c0e7a3170e0b8492b8bf100faf2946d8a94cc4c30b4a954d3195c1fffab98920a2af90bc6c820
z1ff7a30b28bab61660f6439e25a303401cecfc12063ef25107d9bd68369b151f88d56268b48f6d
zd7a9729adc8df8db8741b96a7fd61811186c5f3e6591f27741b23597d8f39c4b363d7dddc2d694
za8765f545d3e09be8da59c28d582976c67a5c14567ec61b007854b769cc07f70070c409b545fca
zec7d07df463baf998a90c78a9887763f568b655227dc0f61e3267156e7d0a5997e5c40958060c2
z4bf74e4f90daec4b84497fc1e76ca0f0e5dc9c504ed47d34c1f2d5499b7a3d2bc886b50e85f8f1
za0c8435ca5e9875a57a7075ce87c32bf4b8635bbfc392b9debd90289cb59a94ddf753471a5c949
zff20379416dd54d217483a71e91821191d0eb3c1596957442ccf43c8474a8bca1e245be8e1281d
zd6adedee8b652985d8862d3ca66a0ec6bcfc3441c247133fdb6c05e912c52c778391240c064a14
z5b3dd36dd1f097d705accb377a19b80c6e253ce407fe73f32268392d13dda480ccf6d1f810348a
zc2a9eb05840865eab2f018c334128a1342f66446b8c2a2522abe4a6e23541329555ad76cd36b67
z2f99da1934fd69929d8d546d198bbdf7df9f1207e7841468ad1e2789391ca3fa4a29d2fef5e50e
z202fee7cac6d1a12c0d9ae44b1070a7c63dccc9d15593ad19b201bd108531e494fd40b4b80c146
z9ed1225111b774a70d656f2f8c1e3e35ddd2133af6c38f7e40daadf46efb78708a7ea8ad880855
z778e8012b1ea06c7a1e7c39ebfcd68f2d3056c1c6cb137d6364ac5d19a65a26ea7dd1690a95178
z9f6344d17e6e8f3251b7b9ff030e62d34acceae77bad5e549f8ceddc6c14255a2847516d23228d
z730a7819f0a47e646ce126c8154b69efac63db76224115df7fb8472d764938b4cbd00e2daca464
ze8e8cc4c167bec0f69dd80e0f2da55e0bc2eac9936e200915675a25e447b1b7aef74cff016a999
za0da3273926e3113820a79396cd9125ea04b2ce77da08faca62a41f472c740900e5bf3df2113f5
z3302f7ca59d40060e23f9642dc05d1e40cbb93859859fe24784def02c66bbd013aaf6b00981c5e
zd52c4392c3815b25a4d2ca53ed2c91daa4ce4ae1e5a8cea272f363c013e8bf30448cc153da47b8
zb048b0c9f0709b3ae319bbac13e50c359ca13cec1be0a6be2a304a264b917a3593507e43082749
zdf4679f286ebf937881f09d9ea0ff526d95739439660f84dc1a1fe0a93248de2db475e86773fac
z0b77322932a633f7323b7225d9a394f8b83f803c695a9c0ba11fe91e233a861b924de0264405a0
z600d2f452ec902e84635933abb433565004469a953b7a0206b9159b53faa2849cc396b795b7e5a
z439974c429e7ea03bf806d4a8399394d06fd645d3892ff45f0c54a3eec4c709862e25abe78a464
z5bdb847ce9afde69a3d6ef80c52810212b2195cd696243509146305349d99012a05e6e383d85df
zb695349f8a1237bfc13eb3f1fea3e626f429acfdfd884095a1456bf8f061ae6321f0409f26a32f
ze6220d7025bf38fe3b55cbae48e890f2f5dbf40eeebeeece64f63492f6ba9884b846199cff8e15
z2c49f1128f3ec17029d24f92c3027f2a78ad8d739dbc77c9df63aa38adb2e1c1e65b98af883f48
z71c9203fead37d28406056d87c828ae195d0f3417de0292e7a46f7bf59edbf431ba7490ed1d2b0
zc8b7d5256c96a2968e6ddfb80120f103d0c8bc93ce0c774f4bd965f250b6198baf4a43b8c8572c
zf002fe5c117babff657240d665a59f3be2c2ce1ec1e424781bc28957cbf1ffb21c58dfda0d4f26
z40801586fdce9f0a7089c7e87765d23dae4b5e3e1a4815985341d06e0de41e1dff50c0d4ce5ddd
zd43f458a5eaf26be6d587526971efec28fbd1eecd1e02d86310af170b8281f654c657bbc566ad9
z727336da2ae5ac024b2b49289f75a2d131b776790f9f1d7b8580e8b07271287b732385fec685af
z7f0e227fbec89ae4a05c6de3fe2edf36164477f1fe415d0fa1222057ed85fbb50fce7e69c994a1
z53336747a0c661e38b1909368c0a4a5b400715d8477d3936e98c41b01dc3ed836ac58c01cfdfee
z7a8e0cff4e8f5fe3382e942437f6dd04cf8dfc11032b69fd32ca2731ef7e14d8c8fb420fe87f2f
z55450e0c29ac4569b041ddd7d419b78fd157218c78c50dea67977c08812716c68877c96b72b465
z4a7a3178af371ac3704cb046ddbe49c9958a45c40147f6d4570b2ee396c07c8743a7135db231e8
z548e850b9ec7040c6ecda1bd38b8eba79e4d95ccba92c4df08629da18cf5276477cc934db19324
z6c77e1752645757d2a338e90783fae1d292c3d98c779116cb7f0e9514dd1ce3170042be5c974cd
zd40ef212f8fd09c3b682d3d4c7879ae20e1d20886f4d273238a59b783210599f25c826f5e7b982
z3cfa0dedec2ed9d19df5d78c5d92303f6c498a4c61225369b8108a1ee6abd136541d52a782763b
z0c9c7a36205de830bef38441f46572e462d4b63f281d329e68cdd71d22a7ccb197bad36b7948c5
z71a0ad0c1d67c66071ba30cb94d999b5a39bfbb1bc0d132a38910d65ffc142705cef1ec275bed8
z8ab5ec9d7f09d039890cd8dc1e69b7581bad7c3c88cf6097933c76b15427f1b9b76ab5beda3ed7
z8b79d7fda6b927ba346898c60306bb1e175d269fabdd291b98f8ac5cdd2889fd70b55cbe30c383
z3ca740a745a7508fbea5d4aa0f253a6e17782284662456f10ca8366e88e5c0ba1a41b8b31e3c7b
zcb1090219a1e2b2c7c7485a733e0f2650d44b2ec1cfdb3cef8a34b65517c8a2e3ceff95f915e8a
z37dde00c9e8a15ac97175803bc36e36a06bbbe1ca9c5773dc42a946ab6956e9cdfb20372e77d54
ze8849125711db497143ca2bb605b716b1fb89bc27ce1e8eec1ae90a723fa26244a38f3de33c5c8
z3ec661e0e2f2796e29958f33021b92c8c394b5a16165d3f38b587085356729a03e5bb3d9bb3efc
zfdaed49eda96df46fb4d91376750cf04ff1b45e8e86f8743c68480f9fe0f3619648f138fe38d18
z8acff82fa17ba419eb8b7b1c957c7cf916e93b577060c458415a639150bc4440dd8f5ef99b0fc5
zaf796cb0101f6623de4e865ab4e15d2ee14845d35207b6b1524d7290c5501e404ceaafe1a24255
zd01ee2f7f91fce873b2f784a38429dffe276af348e90acb03a11f42de2cfa9807c59142d0fcafa
zbff77b68125a1fe87123ecce9308ecd7be807ae898835a389d25c67b3570af9a4cb9465def99c9
zdb0672ff833881a6b8bd3d334c317907850a57d065d606290f64adbcd709071f3b373bb7958085
z3fd558a344ce87680d89e2fe49edae8b592818b5980205c50b5a743d1d3e23824cc89001e43cc8
zb095fb84bb0bba015ea41290c92d82a152aaac5ee3226519743f6d5e87694ac659d8ed4023bd4c
z23e28edf9460b3647c615fb95f5b52523a336df9a9de976982fec79ba4978372ff42b4be77c5ac
zaf4ac7087b83849eda53026b4a9e3e72dec59be90c81fcc9ee9d7b07791bb9c81bf6370ee5e500
z6d162a7856b5893bbed1dfd4478317d59620df06efc4792b71950d3e1edf4fc03b2f3734f63968
z198b6058e3b7565de5de6d24fc21244f62daf994b9daa36e593e3b6bce27ae6d58c7d791902c94
zed6d0590e15b7a6898123f1fa68fae9ed91d9c02025eac8a6208b20e6781359d3c62f662f6aaa4
z3b7ab6a1221c8d9f17e88e70f9184321cde509643426443e918fcf13ad50f410d0f5fafba7576f
z921a117714b34aac7b20e659326f64a990d7c5e3e7ed4bc88006a4b90a2effb36667aee85a1195
z8a687762eb2795041f82fd321bb5245951cd91f060c9223373180e38b73bf3ccfe2aed625bce24
z38708c3816ba36215c69c05b9a5c7502aa6807b169760304c348f62644886c295903ee74eea844
zd6a97a56b492d54ee741b9c59f3b31a3e5cc13fca14cd5a4032b7352ae33a00d1a5ee1f9801cd3
z9d7232f46b8fde276980e3d948a65360999e82162f5c1d562f9d20d41a6c08941575b8d1db676b
zf04c38d5628b04489b1b651bc8bb73dbce4748732133faa84f25e74f0de848ebe40f751bad1ba7
zd7303edc4123496172b33f9184e1ea1af6c2ce2ca3e341320af3193b7436c6ad4b68e1c88d5163
z27498f5d7e43dee696741a1dee84f06d38d7eb6c5525a9886e6c54f0db2daabf428b2f9b140cca
z333b1287e890dae4ac5cb30b342dcad4a4dd1b86f5de1bd028d0bc3aea18c8bef109e06c0aad00
za95fdf1ed9690aa2016312c746c6dc546bde1557a5e4dca83aa0df968cb2d7d0fd02c560c2341d
z468be6cf676755640bb0ba1b70d94505b3bf63d791f099af5f21ec369995489c7be795aa62d72e
z3277a94d77c746fdb86b838671b99c9af1ba4eaa1a045b7f8ab526f0a92b0570569ea93d696ae8
z38e1ce653fa07c097b1486dd86974fabb7625039facea6a01815e342bbd6a6426ab13933734414
z0cf784c3352c58b66f7d78da3b30e73249a651a5c9aa156e630e98ce1b96fb7e0c24a0313caa1b
z74bb209a74b4541ed794a716eeaabb2054c1a75e5c311d213326a05a9f005af14abf757ef21fcb
z551c8e381d708f585ba5efd91c59d4d463154520805447079f1de9c24ac229de2c14ccf3fcede6
zf89ed8602b64ccccbd31db126e310b8a0a494ce92fd1282293bb884dd500436e7ba42f246f6f63
ze70cc0d82857749d1b9401c6e5779ce9a0cca7ac618d20dd7abb06ec62d1ec4755348022cf7caf
ze8266e32b6c4ccdc3ae969b46b0d2ed07aac4e653b2e5e08e9196e8eb63b7ef88b9fbbcdb1a9b1
zd45ea827f47b4bcb817e166fe052c2118f11fcc1ef210e02f2980a418b0d511508cd1be6673c7b
zf1a06ae686a6fa813c79c704f953d0d0f74bd29fe925719a48c8b59a3b3b9b8bed77c6aaa263fd
zca5eca7946ae4399a26cc3dc1116e1cf01ffdcb5f3f984f4960b39b60c8d00b18a76a16ca38796
z89e9985efc1e498dd71319d6c9e7a1f58be7da4d77db79a3b3817eb700fdab94fb634fcd9071ac
z06dc6bd36332ce1182b0cbfdde30c51d9adbf560651562f5875ecb6fa5df7629f102af3bcfd751
z1d61f23d7db523a91b949059c6a730bba4d90da83fcef4ffd66249df47e58cf9230d08f2d71e42
z747de68970d6e487e1ae373fd28eab3f2ae7113180e221c70f96c1b45959d155cf092103f97e11
zb7bb0ab8a8fc8799a97d4af03373c9e2ac69d547729063be67ced0b53028664346cacafd447421
z5480ccdedb2af09ec3c65951917c05a74263535f01ba678fdf9fabc78961c6616a0f0426411f21
z378cceb85c759394cb0837ca8f1906254eb9f68260cf5b53e6ed93d8fcbd85dd7755012a668611
z42264e8870ca35075db37795c452fed3ddf582c4f7b00da06e168ab49d82a1264078cf6952683b
ze803cee427fe27f2d97d9f1e36c05a0036b4045a9d5eaebf41560ca60071d9ee33d23690f8d7b8
z7ba1aa24f4e0d82b9110b550258686378dea7311fbc131c8eae97aeda6eaa1419a54437e85a947
z8b08f5a1574d097fa843549d9e61a314e1dc1a45733eb8b5fe2aa5515ded8992ae312ec6ae282b
z0c35cef7af9adfeaa50cbcc1d981893953b47851b5773897b96c1edb5a2db85ab274584b4b32a5
z97e921411511fd0375e1a2a3b138a27c580fe92593d35f00b4cc49180a1ce83516b1c36bbd5a2e
za4decee2d1f4a0083498b3b4ec95a160d832cd332dea25ccb0bf8037d79ad29cfe8e812cd49744
zbbc28625a930a52e5cd99cbaed768ec30f01120f4c60208f24a74fc8fd40d0184953cd419624e5
zcf2691f70e9637f8eff8b305f8fcc444da0d677f5efdc1bc63bb5d3bc8c8d0b54b565a4a156620
zc843cf2f7c8ebb7ec60b7755b2f9c02922d3bb65248201215517bcb587f7c581f8fcf95ecba1c1
zf04ff6b17d9c2d6a04ffac37845fe927e330ef6e2cd16f47ab56c4bd97a01392db488207e644b1
z19d9ef76d8ee2e7071671e63cb67b5addea34724728250f60f85d7a94546377a302769c3d7370c
zd916882bacf17166f618e85a21578602a98a3d8239a54912891088810d8b178a97fc2b12f0a471
z66b3f5b740b8e8179156268688098026866832cf2d6bcad4e2dcb7a70756d666db2eacb3d99331
zef58fa91acacc406135f5d0cb6cef89086d1075f5a396223b20f27db83b8c4536987789505b7a3
z5885bdada58ed689d5ae463bdffedbfb0f021dd7db5f7b5b081a0abd0d82ee3206cb56adb881ea
z1a70ef3d8fa245172bb80536669964691db89e86e7f20fe26ce07adc398bd12648cf7ad7b3fd4b
z441008e35fdd302974f75c73aad5ffb8ead00b778b4252232f2440087ae974485d3fe6340e0d40
z79063caa5e936879b4c81b60510f2c070de5e5c4744d850a41547197b096e463a6889fa3554fc3
zc8571fa3d02d4ef5da73fc65f9dfefad0648eb20f26d24dbfba95f43aadeed86e15b86b106a74a
z12dbed4b5880f47e52a03fd1d9ee3c50daf5658fe44b118a75fa8862fc8b95dd9c17be267e5ad6
zefd85029c83221f0986c40d146145b89cf1f25b4e112f3ae5c3d0c7452e5c22778dba334f2ba3f
zdcdf871e0acbe253f8868836ff9667a364e08127297405aad92440b081d4188e3df8f490ec117c
z1e2409a030853ebfd4398b23e7373688ab29d6a311fc409c8225334855fe2f9481a77e885aa35d
zcaf070b006ca5df83c897e49c5ab46bd99164b63515b865c397363e88bffd0424939a2f0f793a9
z4909b48cc2b9ce5a84078632b42adc97ae7204d3eacb576f4ac22912c70365c13d33c16d486b63
ze46621e4280d37b036a9a075a433645c480149e1129fd786a1ba56eb55ab173b10f603b5976e6f
z954aa01f05f13c962dba422b78bb37d4e9c79f127778e4c4782ef073d705934921aac93f8c87a0
zc70f542b9214d046e9ba8b7a26b89ca7c5fc25259e9a88ed8fbbb25f41c625c1b312e6b035e5f7
z457f1c9c6ed8b7127f5c31d459ceb9bfdd214e75937de3c22dcd1ace5c62dcba9914ba4c52184c
zb7355e7ddf35480be0c13ff771c6cb51b7d9b4fae8b8f395f18355de423e4c7b346cb4a1c3e51c
z92679db4d4b29fc5798649f9d4cf7dd5213ae11f658401c2eb6cc3568b84569ef2f72b33e286d7
z5412704a3879f0904698dfa7e287c7d1cc51d4268cac5cc1a3a949d3a005ac4b4c4811ceeb1b35
zd07e67a7afd5803a238a7822441294c95bb33b08c2090f684d4879e3954e435c2792d98b6665d5
zeec0d2aacf5be5a13706085d3c311b877eb668360544528a15a23fa1ec1d6c740cb3f1b1256602
z5cf7217efe02a133a98fd447ac9a263e53f0a562e917e68e83cbc7145b437ae8d4b4aa5275db94
zb9759465c11a650c3c19bbd17ce88903f1165a79b84ee7a4746b3294b9b9a0d1ae5188a48a8314
z0a45ac9ecb829ad77e8030418d2648ebb48255bd623a13c30bcff3c8532c5440f9d59144705592
z0075c1e9e2087a28d9ac5c51399c7cf3a7666cfa4de9b8625f60431bf8e546d49395d24bb6a9f5
z7df83a069f92bdfcff63675dea41689524fd754c7ff3f2672bcc2e66c1c5ea97520bee4a0b64c9
za52e95c5f23ccf19d01a4122572ee077840ed3692b679fefe25970cfd1f84c2e7c0176f9bef308
zb38efd755ba44fbf844d0cbfcdcdcd40eff49cb917e883478f8ed6c31ecb43f01eaa325434c177
z11bf2b4d4d57b9942c0c09124a89f76c7254bef18d183adc8c788b1fd9392fd427d3c87a2ffc66
zfb5257ef4731929eafe5cf9cb8257f19f2d19c9f73be7722b79a971b07997deb49ff5216320423
z5bec8abbdde4fa40e8757b648fd55789d4eff09b3f4a778c4a648f174676aaf22d019660cb9e11
z29aa590f0e03f4a65bb392a2443441821208338fe1a8f405793b2ea43950e2901793705b6e3b03
z208e7b4fb1d664472f5cffea6a91a30a5f4b8f90f13dd59ddc014c276463c2902d79fbc0914e19
za72815326b9f3998e22b2b6b10ce838477aae00c6c95a6d84e37ec280591e8395d291dbc6663c2
z18fcf306f814b2c8e94bb7db21ea6d027ec8a9b471196e7b0079dd223a4fd1e4d30873530f18e4
zb88bbec824580b8186d7e127c5b72c40ca98cc1730e865a34c6e0043498c76973ab1d0e31ccfa0
z59bcdac0c49f69f56394d49556b817d5d1da16b78a937df6241ea8b0871ace9035fbebcdf1a0b8
ze20f8a595f4ec6d5b00e2eafb4273819c9cfa6feead3be5910b9d679b1c8c412f61a0e8f789576
ze1d383561997bb3a4b7e5e7d791a1a26719a56a876002fc291d0e0d4f6880121401e7dcb0212c8
z5b799379527eef34fe5316f6d44a45ac877c904ef51b6aea5709c995e6324379c8e57c1c13d99d
zf2b610db65b4f3c34579456ebd2b079711d8d9a56a59ce5a3dbd1fc1691c244f9a0ec865393635
zbb1c08e87385f36679fcfc342d6dace59bd2db298f39e4b3edf222f96ecd8e3405c37c088b5ebb
z42103b39eb1c221165bb92b593cdab2932e2836943075c167aeb01fd399a6fab2a896ecd100f94
zcd8a3311d1629a788c8220b0cc1c18d3f75f8a8fe6e18fc7ed2b9566dd7d445a9387897a1a6235
za5c57a51911aab7d88849896d778b96f736e773c83c0efdad7fc63bd21bbb7b8719cf462bd2881
z9491daf45e7fa686d8d9a89ef45d47be2b13d8b85f307e8b64b9b5b940d90f11fa35a5df1d69ee
zf995a04027b54c29c272707be0260ddd445042daca602868575eea58b7b06808ec4bab16867d54
zaeed9c2f73276508d15b2e53d7433f003466c4cfb6bd3e0f14e443f7de484217757675868d98d9
z9f857fca2a9cfe0b2b71ca02ba7e4e54f122664c1fa8114aaf48bc52aaf99d96391ae6f802c0b6
z6866131bd10602720daed16c83917c9e3168eaa9e8b8c7888e490502cef54106714e15d194c8f1
zb00db7d113b20918aa1d9b0a907e68a85ec0ba0aadbe34a86ddad0406455eeee4b63df40fe286a
ze85c1a2a2c4d340cdfe41a7bf6be98911fab2686bfe64f79dccd0c99ac8b1ad10d0c152475f745
z327c700c88bd4c3116881c3568e269e4b9d0857352f6a9b18eb36dbd1e46bcfa08997494886cb7
za7580061b81e3f1631c5aab5e2a1be905739a9df0a3fdbbe05d54bed9b704cbb14e6b364823ced
zc427eccc38f0a959ef14d5e04b5cbb024ba34aec1ee9f282b7fadf8d6fb38441d17e7efb7ee292
zc88717d6f1a8ec24cad9556be70301b1501f202a89f586912152df17a1c70e41fce4b7df0dd318
zf746e960eb7a16cb3ea160ae29672dead4056603a7153836e1840fc6590d06120e4f681edcb92b
z27c8c9da3e54018b062a0cdbab386ee4b343a85b00f07ba34636e292247e78738b15cf1ee6dbfc
z9265638f45db8a33198fad5188947d760ef76f0e9a84386102b7c04315288c29412e84cbb53396
z5b1a48782c2310660d8b7694f02172799d3b8d291c7581f8d8b58c72c2da8952ead1a3aeb74a92
z3012ba4e7910adb868ffdc5ac055b475a5b4a56dfd98151beece83a5be59ea7a72cb2028dd7b29
z016877ac5a6d967425cc94e91ab716a3fdb7840e3694da21a3ff1499a22f941bffdae58f24a3e0
z8dd4d9f9b5bf6225a899f773715ad8629b43983d6ce0264a5a12ed1145c843029e5b5a320fed8e
zd2616c6033326f393a86cb0a3a965efd016981528dec29beeb325df3a21280da33b2c0242ae18c
z20a491cdffd6690bd8c2f42fda6bcd5d62e513b2f0b2a3690a813bd35d4c72315806d4216cd0ed
z521b6e2f03cf0c1a852120bd13dc5d875317cf3f0dcaf76369164c348d857677ac612a99826da5
z4fa01952b89d052f6c78e20ae5f81b1db7c3b41de3923a6590593c7694b9adc396f9d5db5acc5d
z3ac7fe5bcfc6ed54dc597940b1e9e7c84716f4a1f7fdb2db0823d2fd0bd82e56e5790cae49b1f8
z8b6a2b3ad74bd436060c784a7a9bdefd952cfd27f4d5fc59f616409156cd166b644069e740e1f3
z7a3501e8d02e0ba895a8f3af7f08e37f563137b5d87b9085888f846327362961e1aa8fe30dc143
zde7155bf7ebe89459f099687ce4318ecb1633930bf211f165e2e28f25ab4d1c5f5a57c93019898
z8cafc620fce27088a59cce7546015e75271d524f562916edc3ad01826b24b31b7c1f2a610c370c
zcea96d0936f79d6a34ee584bc8e5365f36d9edca7009911ac448b6ea06ec1a89e6d94e0c25ca08
z323dd99a4d6bd8361c680dbeaeeff0a4e8af1f7e5b33cc4a9e56a51d700e8e0ab9ccf2cc9e8f23
z0f485eac7b46a71ea12915f1a5a6caec5a2f2786e49c9a02c2e7c25d4b7a64defaffc28cf8af6a
zbf2de56c787d7c255039509bb3c9b034600e6080d52f658abf0f8104710c08bc2a771f49d642f2
zfde667879a35c40a29459bec2ab5f1f5392d87079a5efb899d5dc9f25883b926ae9a4dc6c3c6f5
z560687c8693c1893a9d6b3e25b8fc0e7f7033bc7d59e7e3774d3e86daaa1e59fd6549a2907b968
z8d454d918bdee1354b1bb697a2a7150d2284a588e99abd92abe5fddc56d27e113c11f352f88215
ze8cd2bc41bc92262ad60af343f6bf96852e18700afbc3bc179cc248490f091aa91840be8fe484f
z23111794031ab9a42f6a91c7b8ddfc8a26a6c33a356a6d9d461df699a48df31d69e438f128f6b4
z832c4668d1381c712b5bb751fed04bd27b355dd4e43de8af62bf1ebfabda14718e390100e2c802
z2a422a3ea6a5a3eec6b0fbfd4edbb7a7060f8400818a387725b13b6f6bcf609545fcea76e52b63
za74e0c4c0975cb21d5bc20b6592e94b5e3c9b1aad8e3e27052713f02deb76186c180e243ac7792
zfa81925a7bfd2449527b1c6946e85f6ce396e8d468e9cd8893fd524ca290d634e48ba4319f8c34
z7e208a7808ade5838944e2291dbbf27e39d00af015a58d554568fa0e2f1689a8febb6d6b4e5b35
zfb5fa2811137feeb4b11b7a7027a2590f0b8faf45d13cdac2c3f18a1deb064e20f999c8375ee19
z60433ddee405003f23bff4dfcff0d47552c29e607dc9cde558c8449018935d30a2d42e5509e5f4
z7d43342c8fd668715a1aa746a63155946edcba05d96e5b134e8bfff19673bfb00cd719ef7b5c9e
z5c2c16a8a9bbc320008e33c8d4da5fc270065ebb99d7fd755ee8d129a09fcb456e9f2baabd4d9a
z56276006cd0ed0df2cad904d81ee46dfb9d17ae75d96afb98c26a91557f4c8d2bd070927a2a8ac
zf63b8808cf050f513674d0871413452a9757792d8dde02a52283bbfc2dd32577569990aaee1762
z777d26e40f1ac09b484f22183ca82ae6c07de98c368158e261feb6729c8ac5f1ec0cc5b72b1b30
za6c72d5bd82dce3702b869a35ccc0fc055e8a0cede184290c7b6dd9cbe9164ac58363b7b97e77d
z1b808b041172296c063ea31377d2f9736c38f0f9b65342374a647f79a3626b31ac633081a72405
zd2dbc2b7487885f5227b49cb0549f076be7cb89b2f088b2de126c9b8092bf5f89f8e8bc83b2e81
z507b595a4f599953c27ca75dc0b38bd26e43cd5cce244743cdbce16a4b0fbced335c49dd1c3f7c
z420b29441ee28406f3460edca2d724bfd039cf64dcc6c1df88ebcdd753fbd3e4ae5c4b9603e4c7
zefbb73a619a295dda23232ede7a28bbfc475c35dd2399fdc73566306f8bfc1666a2be770630e23
z89501f3dd223ee3c6feea1f86d78415be4db0aaf0a41858dbbe2260f46d97f0b6eab67e49d9043
z1a9fc8f5ac177a4c6ec5d90f2d30b96181e8ab0e1374bb16055c575e2e7754dea7fa4722dd8f3a
z333970cb4f2823c0121fd933b97aa728bfb8c308f96ac134b2de451d39154894be96e395633127
z12567f1c16023eba1b42debe03d1988c8d10c0375327aa31479a7e369b281d7ab59578c8226e8e
z89fb44ffd675ce95d89f1b670e7d432258644324a779e59d938d98807a5341849e0a393f1dc50c
z5133234f5c527d56b94c68be67dc98c48362e8b73c51fd7a657704bd94073799dcdd9ab32ac3eb
z1d2fd86fb33aff0073f49500252ecf8fe011f05448084f4dd590fa528a028b1b3a351b80509289
zd3ac333acd7a1e519093a957e3877ad1888f1bd284496088a54969b45fea0e741bc92a174e4d2f
z80d9b8b36e0909abdfc436e4bfedc5b820174dc366c0f8b43cc6e657eba09867d9610ce6bb8859
zacf6271eb348ba365fe4ea898a9c436d563330ce134092928aa175b4f7e2cf6f253f954d65f992
z5360e31f5b50fd360cf733bdcf8081289c9be600ada17baba12001127a2c59225fbef3fb8a2842
z8deb82ec54cd856521663a85914c16f2398fcb835ef9e7b63b9200e183dbd0a7cfce7f436936ca
z3d3d65547885b175dd1ccd0ee99f953f37b2cfa5f38dc5fb60acdd065bf67c1d760d9f7b51fe78
z34b388179bcdf6f3f926e5033e60d460809946bd3d803528a826dfecc0aea5c33d950cf3b1a332
z263a5d9c4ed8eae511620357518d62fb540d7c80caef7432be22bf5442c6e3ecd50dea7c1dfec6
z34b83e76a4398e39a1b0498b3e756f4209b2c86fcddf86efbddb14858847625f7e3dec0b74e7a9
zb18b38f4f09b2e9ef2de937099d042879445abfe8375d2f3d6f46aea721aeff0efaa93c7878089
z77dd3d0f7f1fce1367dcc49c25d72887b03ab235e4a42fded2552b21723b034965b99fc2e96048
zd4b1c52f88f5b16a01b8faab2804ec9fff1530a5b4110695015fae9abba3326920a3aea39bba5d
za6701baf6dbdefa192ae95939885abd635e8ce333ea0ece7b658a78166f7dab6d655cbe7b994aa
zcb93d6d478a1506fa196013ec6a7089426e8ca361ac5ef617e3ac746d23287ff35a229b74f075b
zf924ca07350b4171a7417561e11ab10dce36400c0d32afb49a4bc911c981bfec780523eebd8ea7
zd3ccc73560dbeb2c676cd0fbb5058c977a3e4bf1556cb31247f5d92e9d0ac0827670830ffabf61
zc4cbe36ee4724d554c3dc1cb2fab2484649b76ab95e0bf2b079ffa2173cec59d70896d89fea4da
z9d4c368c6d465740595f3139fe2dc850dc8dd20c9fac74971e025c74eecb987627843fb1eb7d3f
z0a82b5c43a788b5984e58e83c27de46cd591e78269d153cf5764b46b0813bdffa78d454e935efa
zde4f4aed8c5ee476a3d6dcaedf64e20b107ccf9b2630e6edd330ddaf5c04f8a7c07ad7f4cda0df
z973f3399725b576a63d5252b7b893d535e31c2f236352c8d38989e29dd3186f5332aed8dff8cfa
zfff45349c574c5c90e8d73c609ce02bc1c47164f66f8e475aeb10cadede6886db890a7e831468b
zb30e995f78f78c8b6f1adde90a032e064e4154ac03e43e04bede4f514b6faf593acab3e3064d12
za5d2080ffa1b3dfc0940bc311c8dae223d5e9d5614565811bc11b41021e61a0a3f3dbbaa65c58e
zf843bb44d212583ce22df6a6e4bf8fcbfc316054890415e2d5a8e6b6c2aaf394c956a9a6502e5d
zcea28d14249536279b9a75fbfca373371d2c5cd446d79c4a5a13793d8c4f9a8f530169385cd43c
z6279a9c1ea5418db80c68f2e8183998df0f86a7c039364f57aff818cd5a17f24f583962ce9df69
z83d226c2ec53d7c1866d4f4a2dd5f5a291d7e5796fdf53af22786dfde05238ed8cd052093b8ddc
z44d42297f95d63938799bb90fcb60c1add2476a6d2ad0d46381c399a41283fb51e02cb51b41d69
zc5d2438ae395e55dcef2ff73f3d16375ada2bbdb8eaf6bda5e6c095a660298b50b8a6aa68fedff
z598cd00b80a4deb94b27977a270a1f55f00c09018ed10d7ca7659eec89fdfb5fee64a739c140e0
z9253dd4449844d1c0c22f31da9c832237e443a2acd0e6f159aec6dc566aaf5edf5402814c65551
z00ab4fb63f2adee8a4eed18ab59b062c12996d7854b756f16318884dd6e4f19fd87c5bf07eade3
z7340abf1c3ea56a6d012d1ef62151a077e8a3fe4000f3fe466db488538df451272087a3e6e459f
z051aaae8ea63683f5b0402637207011ac3ee0712152ef3484edf3aecb8d980ff016d0ec045298f
zc8a41a70a49c6f2c4eb084d0e9bba71f0a9bea949ad2f6e867e6f5f5a7219844d9f62b1c6a33bd
zc560570b9356951ec5f49ee98c5396b690dbef2405e2007201494e72500a476409f69a655563ab
zee01a4bc4d2e4f671664fd4a21185f841d81ae8294c57d5fb8995ea125043dc215bee26857ffeb
zfe47c421c6808cd6a68de5533229330fc82668e81b0fabbc4ebf916baf00dc6a336d7fda01f584
z4f791392137cf3a25f3a90ed2bfa72069e3ae94f981f192b73608b5a8048b2c15ebafb492cc61d
zb5035f1b814bf20f5630c3e1fa665703c9d01fba5545ff976140e0f597b37ceca784e27291e056
z607ab1201e5e16ec85496a970cb7149301018c288a9164b03dcc167123602225cf1a6a2b5fe4d2
z193f115b576c7a3ef950a8dea352b3adc75a3c9c979971bd41cf442ae7b00fd3bf0cf060e43cf4
zdd372dd7f31066a951e31068fe67cbc77800a8927f4ef3f5c8ce9fb0f515ffda2d846ea630b788
zaf44cb51b955e5b2c6d7dbb6b6664095fb62de3b422af3cd636c872017baadd3107ad9bb761918
z8a242ed2c8c45253a3c5a606175e31bc29bdb7058e882f188d7a0b67a9e71f85dbba5c11042247
zd2da5e51962c48f12621901d095050334fdfe2ab1ef549546f034d4fe8aef368fe9c5bfb8211b8
zc5c9a3b38aa4a6148b06e7574e4077cb759fb2be894f4f343803cd197325be290c31e59cc4c538
z3a133793de70b7bfd37c03d1403047732a9ee0b814c5d2b7d4efe95e1e5231a20d13377f521bcc
zb5c8339f2a22b173930d4c347d0c90d26822b6c899f085ead668961d0ef578b41f33be1d134a33
z536ad48f175e38d3eb1d41c4889c779443b42279c551124ca9eb03d109f6687b932d4736eecbe1
z23a828f785cdd6aac2d017e9f75e2a1cbfbf068f2f34992e8a392f0cd69ea347ec8b07fc49ee8e
zee100f51697b97fa77667f7231eb8262df476cc076b97705813fdd69d39160e5b531d92ce32384
z9f83934fc735c650194550d11feb7ae4edef28178a3a72ea34fa21366b6bf229af9781e94f76a7
z725ce7f8871d0ec6f672f244638b64f13f0874f8215dc2eada8bcbcd0e666a7276e0cf23b73703
z121c135841c03834aad1d32637c0d8c7506f8380b690d8a11d881ac22a8898fe8bff5884bb0fd1
z8e100c4a5dfcc013537d66b39cb39f2136636d412e60d4631038d1f38d0d18e768e887958e6a93
z423b454a7a68c271fba9b0a081f81c2e8365f37216b4097bc23c203f8cce651abd61df7002a095
z2c91f8e2b756bac21f66e9032ab334748f897f96568b84039e1dea6d1b165eaee9d820fade0b36
z1d0f9a89c06f0bee005fa4367b1f4ab6d0549186ed623abe5083aeab9a8d42dbd66f6ba3510b7c
z931ade4d164e3914859e92f640c8a642dad755ecb1d9395a70200eb9cd27bc80b6499ced3e3e22
z1ab1b135e9e866c275b88cebdf45f1e5c87a0c3efddf0abe7e154f2d67d17113dc24365bf665b6
zafea7af25a39d8c1de0cd9da5413978a6e52173671ef5882fe851edc76756b74689ae6208cfdb1
z27d19d01d6193b98f28d75114d221595a07a4bab6ffcaead22e806fe76778d3fd23711dea26e0f
z5b2155b4143b63fd371624e6a8258aab282c974837b6da625857a60654946d2074f3041cf8e7c7
z8391c9bbe8aba95a05033fca10e8159268dbedae66b12ab80235356aa75e6262edeeedf57b4a59
zb5b472d1cf1a46b7db2b66647f729c3e95929e262dda02928665b14c6ac81258e8e119231db5a4
zd0b08a9d2b647255e91b9f80cc4b8439c9efecda60c0523730e6d1dc5d4e53a328fc06340984b5
z76d54ea9e79fc6d4ccae432c36c2259c2e7cd8dc115a5ef66a5d9c2cac0099b3cd0ca0bf6fba77
zdae98ae0e54219ec824903a2b15b105056da3591b48584e91797ee92f7d0dbb1fa3558b8b094db
zc82fd7f187c647a8e899b9fe297ea67bf15a0ada5b88341e74532a4fb3844b3b0728ea0c6a944f
ze78a074dea9b0ffbd574e2cd85d276c369364f820f454f5b7ad00753ccb77daccd80fd3777297d
z8db2e82b529bcec0ef5beb94c96610145b96be64d4057965fcebc351faa944a8eaa6242aa358c3
zc0d87e8f34dafebcc965631d1ec288e2860acf5f517e336853663c4b1d82a045b5417e5329f92f
z6fd46e6030c5007ecd404fe950c49a2928bf22c98fab36b48032a7f7a8631d6b0a7e611ecfe13e
zbcc1a9c51dac3afe889796a2fa0843aeea6bac150349fe8a3b2c8c2ae10f4367073d686be39618
z4e58640db17d207d5716e36629cad88df30bb13d0308493ebccf10d95dc2c63f5458f5046a4e90
zfa636050157aeb86f9bc2d5376963694a0cc2411aec5b8e7b53f8cd38bbbc26a49531ca11f58d8
z2108a67072f32716e09e3acdfa4ccdd100c0b0cdd76652c76fd967d0ad4a32a0583df6968415f5
z37452b00de412c59bab27dde2bd4e86fbd09f0be776a56d7579a0cd3c5d727825e89d6b59bb002
z020828e5b5dc4ea059137741c06e03154cf35009bab9b017c9511f4e03e4010fba3e98e8a317b3
z2a9f045d11bd228c0375319849d046d4635d7df87b8bb06d2ef3ff07d72c1c32a0fff32066dadd
z27649e7c6527d1d4d10eabf385a88ed0a9f9fdef6e5055ad8e58e5fb0a435b66c1f1340f1d7b0d
zf2f4de96478d67a2cbed4237317e19578ef9c4bdf532d69c5be34607bcd9c29c154cec8c0831b5
z3b16088eb38c6f893468242011da4bd542f20bbff74b93624891a7c5ddd908af7a13edd6224016
z826358a3ed88411738d6d5e5e13cf0c58746b91f27f1bc5fc98eed084859f0d59248dc19f3c75f
ze9dea2845ee1a1c77be0a5461272354f012de1554ac32a5b7cf3a42e6208ce4601e10ed8869780
z3a603057cb6e33009cb41d29e5ad9818731d3732a53c61731b799747e033b9f99c24e7ac71b255
z37f6cc1eff2e2d78ca1f4e4823a25e820de99f7604c99053c9210ad00468a492e3fadec9457c48
zdf9c4f2e06a7bf66d642a38c806044e11efb65de7255ee8ffb43a41933d9e5ac984cd36bd84306
z73f68239179ef27568facf9bf1e4c2b9cc8adc4f16a3009879002790d3997150a1c6def721b3b9
z25c15ca5b57721e6d29804a8db6f617a43251636c20a8c76eca769bd7a69ed775e3daac8d86ccc
z9c68e93cc2e79a5ea5f1632cd6832b8f680eeefdd6510692f4e835939938f53f5a1f5a56d7d7d9
z17dda3f018b6cbfcf97d29e960167dd909c7e1fdcc815100a6390ac0eff1b0bbdbd195981a9c8d
zea43e23a6897aa44fb785de9657cd50969b4e87eff306569e50f353d5241b6781d96f66621db37
zbb097d742f0c6c10e8a120708d21086d5d6abdb6b0e9e03a879363076a14a798716da27ce19709
z400dd71124828619cff9e489342099f2bced866d863b0fc05e30110b107c7400d5745d5109efb7
z9569c0051cd4a923e1b002b83eac13c30796d58377e9775b3f5c10639ad67d9ccafe89da70591e
z876f892e7fbc8e731f65658c123572a297ef72d3dc67f0729d56fa5492bb0c9134977dccebf8c2
za1d37c4ea8fa54641fcb5ae2a66770cc998ab9f53d266a64333d081dcb8b9a30b5f049c12fe724
zc0c4d020e76347fb47a12eb784c2c5395454c7d2d183f10f542228917a621def0b94887ab9a0ba
z898473840650661fc5106166207050793f630bfe967e1769c6ce2e75ad830c221c9cc5d90aaa79
z62f13fb64c646b1fd5280a0385520c3d5d3e036b5e7145340842761e18645eadfc4bc08cc2dd37
z45116c03abd462484060c2a34bf2d63adf0a5e6faa4f390cd0f99cc22d2ec855e3ca4de73ac3a5
z0f94b410097e99e16dd2d78011b597ef4ca0939c715a08c12d2a2f48383bdbb2c15adfaf03d28e
z5bab56b0f30fcd3110735cd309c647959e3b614495fd9cfb75257785dbe47c253c1747323bf582
zac0371aac0752e518f0370c8d37c63c22b27201d544ccda04ed2dcc94783517a78a193033144af
zf2ea53f68ee6e8320245e9c35ff8d5652775bff53e24ae198c6c50c6de2326400c2d6224b3de1e
z08b5b2916376f3ca3ba6087aad36554ea05abb08972b344f168116e31b9bf70211000be752f3da
z9f9523db0842980d0475d78b7d056feb549a04f97a268c10f21295effe5d04d6c8483b6089b606
zc5aff15837526d297184555044b57a2f114c3bc2310bd8b4fc580d466dd41fc55d12da6ec1694a
z7450afbc33a2bc6a4fbf99e91672f107a6b8f3afbffd58a8b0077a447bc808e3ade520c6be8fe8
z41c0c7dd73267b3df57b0f3039176c03874283b6caa22fda924eb3adf398765ae0a0c704da72a0
z8bb1bef1d81d1bedf65b124374793cce777274b266f4770a97a7224b29e5978dce37f1dc356ecd
z82f43bb9deba5744e54764536e09139ad1aa5282692fd1b4b8021eb929770d39dc42af73cfe9b6
z17a931088ae3280fd2505e3596291c7de82c590ad447f99f3f0d2943057b6a060460cc13c86b83
z23b1a7321a7e190e4e3e3e130f1aefd307aae70f1b214317de838c8cca22b2386778d69f719b02
z78860002fce62e70b13d4a6b32e7e7e78dd2c469fd0a5659c4d990bb8c3b8a83f618dae8e51120
z55f3a30b95f73e1bbdd3157fb2a37f6a172201de1392bb9dedd080bb0eac137164604864d0f415
z918a05d6fc87a1f888e7090a5230b8797be8088217578db0e265259d9c1729bae408b0f228dca1
zb8ec94c8c8661710972a931e42050d63ae92a64ebcf1a3e89846edddb041ed5b649fe7a32b996b
z737c5cd1bc118a14e735aad3efe81f3c63ccd8d48d2b8a5f55a36dcea29c850721385c6728d1ce
zddbd30b493f82313413fda26f65f6e48977b0da7c0dc72ac7832abb197d83746dcfa2b5c4b95f4
z1c3c7f694f6d783e93dc8e0af4dafa5a2eb5d4b63575a7a1048409d432bb9bf7befa71ef74ec96
z65a2e5e7d6f34f560e72c955f9a69b4dda4faeee196b12f337c6c9b1939d6b18160c1635e81626
z8e5a8db0ddc8110f9fc02d228c89e175ac74b1936e027f0a26cddd91798b3fb3fe65ab441c25da
z9b70ab4c5c732bea414431a79a5f866753d862ef769fd2cc036b4a59022225452d9bbdf54ffe36
z7e7dfb9ec69d855d81e62235cbfb8aac473e6e4276ea922ee2d568c3e25a6cfd03bf6291dc52aa
zef8aae43719d1fe6ff60df4df426eb432fe07f1d8ca4da109512a79a163d3bf94e92f501ce159b
z3d67e6aef2f4113be64239032ec8c043f3530a27c2e2c5e9e53b44096351dac0b56ab563bd9e7d
z818c2f3436bdf413f8191e9a78ceb2fedfa0ecb3bb18eda3fa5be0370d7ff1a3f0dc35ad9ee993
z43564982d9f6077573891ca67775fbf52d536a3faf12938e8dda2d6f58af62145c715e0b4484f7
z3709b58903c107ca8ce07691a41da3793762604c174b86940c42a57c570755b6183b01f81c6600
z8b46924696bc7ee8c6fb58cc8f17df9e3ac8b1df5bfaa44e66460b4782d0147fc6756d82292367
zd3d3f2c4e5e836481794bf16584fb0627702efbb9e208e5bef5c7f38c1919daa9f83588a627dc1
z49c75bfeb9c5c4b3ac98e74cb5c6520b1574cba60244b446f01817ba328ca42211332b5a1bae22
z9b1bb1c34bc234ff8ddf1cdd2e448cfea43311dc0c59a515baba19b009b97581a28b82db31ba81
ze63f508e863d28c000d3b358f665b69815c13212f4c0871a44c10c4e2b8ef8bc8c3a719c1a60d8
z5961b93047c967cdddcdb97c751861da866b7e49340d3d6f83c394574dc0c651162ad88dadd984
z7ff91279c25297f001039eb6c34189b3dbe659275d85f39c78532dc388e7d2bc422d159ed1c396
z2d5f913a9d7119f66285264cf62ee8b17b5d352b37ab632a1fce7199dd8416921e58002c4ee6f0
zc0d98f43c72f78abc9c5310ca9818af1641ae5aebd77b014b260544a81f9063d73eabc4d37299e
z76034066aab835f862a8005e350a34783a7db884306462fd2662482b61835daadbd77d35247b93
z720dde4179bd4743966fadfbe813b1c8ea0a3498f733099418310784c8e93c919a99bc4ea31aae
z03ce85ad16de6e66eec5b7b73c85497af3179e123f69dc4d558bf3f52f4bcd5afeba4ed6ba6f9b
zc38e0b60d0fbda817ee1b1a8334c4833b11f2850b481103900dbe5903eedc25da947dd3b879e40
z918344240705e6c5aa256aface9c935dfb55fe26a2be591ae57f4dea7390e0da83aaa4facaeb2c
ze6ca10922953802afffc662e0c35c6eab3af7c09c58e86180f1f2b64db4045b5e281f47ea299dd
zc7e489803b573d01e02f87c5fcbf106a9ce9f6a5167a5e87ed57e3ef5c644769b4a9ed918224d6
zbdc21566f9f5014d04217a6035e0dad86a1220d95c3c4eb4287fbc94564a35838e65e3cc916385
z9afe021787cff0b497308689e9015ace562fb07f98fc1012917a950effb70259f6f1aa4791d9ae
zd77b3f27c272eaabf5327a4f6001be1ef1efa1c8bd8118355728c425729619d9dd469414c81f7a
zf3cbea9683de926a418a0b7df7b1b422449d7021391245a48bb413b230554a4d5ab754b45fa22b
z173e9478f51e4dba95aa980e35e8394a7c9b75d4b72c81be264d25b3392eb3fb7b942e40074a18
z2b60107d0b9ae969063d3ead52543252adbdc9e85e35254ec1e424122df39f71d3f3fbaf7faaaf
zb02c39b8cb749c9ff7920a414517ca3c3615592364e824f9ecfadd0353c42dc1008f63f2e16b26
z8a65da879f3f845dd45830ae70a4380fd755cf0c6d47bcf50275a8e3b29d67193caf43a90d9c4b
zab0e8250c38a86f7d52c54853b1835d96aa9840ab60f5887d9026ac2a80acce89ef1020be62fc7
zcc98e5572e44dfff83ab7024f6b80b13f9f05a45735707d75f529289c3d924a033c81f4addaabd
ze6877ef34526b04edeff204aed3846ff46741703b0f8ebbef8f55fd537a236ac185b41bc66c1bf
z0b2f05546a842671596013ae971d98db291fb37aba10fb85100d00a38ff42bb384c1071fc10f57
z98aa0989008a8c18a800ce4e09d26624eb1acb8271d3d0644c93c82740ad8787ca9a2d72f2d1ee
z01f8b54ccd35f9cdb950b183eb41970120ec7ab7af04a6539bc7f24f2052f76030036b8542332a
z92acd20a2798d7c58d9d063fec248173795a4cfb2c9938d9a2440be2e5738afd40cd50cbae3f76
z4ef737607c86434c70058b651718378cc96d7fb7aad593145fb00a26bea9909f4a405bf40b3174
z385357f191628732491ff678794bb406f347619f72b89bc0f17eb5c50628b0049bebd0d0753b30
z0092f44c04a0a5acbdf80c48977a9ea21c251750d7c86b4041e07443b754e4cbdc69743957d5cc
z786735f4964dcb4cd6a8fddd9a25a5cdadfdc5ff8ce213fbd1e8ff322307cb6adee98cf0322b12
zaeee2ee19984af684b7688aa75bd9ae39d072638
`end_protected_0in
`else
`ifdef MODEL_TECH
`include "qvl_pci_express_link_training_monitor.mti.svp"
`endif // MODEL_TECH
`endif // encrypted_0in
