`ifdef encrypted_0in
`protected_0in
ze74c34e226135848fe16db9ffd31815111b6d7fb642c521a3f628cf6da949865580b22efd062a7
ze90adae0e65e66a2c36a587d0a790699161455169ed55a01f2084f11770a774ec4c588039b380f
z6de9c5084882a40b79a175f5c2114b2b6d78b070cb806e1c0aa9258297f4687ab308bc470f0040
zb0b1de382961eeeaf2e279e1462520fc31c119af8f2b214846f56c2b3cd2eadbe4099496abff18
z15cec83ec4a77b868344aa20ba7360908f5c0de2a79abf8b3534b883bb12180f68b5d4beb444cf
z3fba8f13afb0abfe8fcc4294810f75afe452434d2d0f1166236c82f76edf1e12979f04bc35693e
z32ae028996dd85737a8f5adc1ebb94f39c940246e887647b64782cd7ab429b0544c173176cede7
z01dfb26b1f73408344a52b7e1f117f12bb9c8077b34876c2e6fdc085981637012dc9754765e1a9
zc512ce062e0b8fb16a214591f5c81e1353b900a611fe1f4886b57940b41b7f2ce99a7b84b04b90
z916f717e73bd10589c81e207ed77ec660a8cbed5b487fa50acde1b055c8870bd8676023f21ddcf
z9c98cc47cfa2d654ff1365d1f45035a045a66c5dfa8279050262ac56ccafe221d4824992a69d8a
z0056c786d54cd57e5ac49b6b8aa4fb7a6065bae21c146cc6f3a280ec9ff5fb2462d875cec3d7cf
za4a6754d947c9e8ceb6b4c9790811631af009d1ba6728b6dabd8dc80bfd8a5f8cd89951b8e4467
zd9d6c892a79c94da04eadfcead6cdddeba689a0850ad6445693322b01dc6d064cde9a4abc9cff2
z1288ab51f7966be250c05a75d1210f9cb74179414b2511b5fc7b23308eed1c73b1aed638a774ef
z3a2f94f142c7a12f62ec09ed92b26b7ecd47ff3ae54934d967a5524ff06f116928de56eb69834f
z4b3cf928d97a885def970124179a048124a7f3edcd21f0a74589369e8e0b1253c995c87638dd89
ze66a29d07ce6047b1dbd08f0d368390cd6f39441c50f191a8d2a5339689ae8ea300d7f1660299e
zce0e190b67691acffe0555efeb52d7f5e2f19a033dbb6127f1a529d770a33987225b4ae3c0bde6
zd4fd73f5b17ab797da2ae9054daaf9a9f1afe5d42ab832111832678b2d09b65efe13b521e5e114
z6e83da86b5b5e4a8b92ab8f4824a62a734e0acc6d51b8f69ab20df0203fc2c98720245ded05381
z8c1fabd10599ac3ee11bf27215b5c6d6155a78cc96c9b58e206d9daacc9fbdf37aa0cba0a90362
z023adef6b0bbe313bd00bed80add3c1b7ef42834743d120ce8a6c07869bac62ca4efa6f946cebd
z9b7aee60235a3ce832da7e1c114f22ed59fe16687c02cf615d89682ec02f592dae32569ac1a6b0
zdc2383d90ebd766d085d4f284cf9779a7b2fd2a168330fa07136c44e148304e7d9a073dab9525f
zdc294432ec769d7960f7ce0e4386f29089ca4a1da02f6085a283eb2b1a6806c7d7e4bab95b186a
z5730e57f7eda41fa72d7b1c630527ae037aa28146fc16484728e11ee79570d6d76022814bf8b3c
zf6173c87051fbeafbd5a4841d0bbe9c7c7d120745e5256d17ef9e6997d690d6d04c5b122d930d1
ze8981f5c16514857512177d32dd2e41f2988d1c900498ec963592958d3392619000031459d20a1
zbde338170d1ae4e597674c82bd772321502702c9284cc0c2cfff1414a829b4b2c4540320d2d728
z8a5d5a8fb817bd943c8a849c933f8e12a15be5a445e54d399d0597591955afe575c40f4f56000e
z380997253644da4559c9c68c5edae68e4cb6febe0e54643ae3e808c0e170bb0f8746c9c16ab829
zaaca623ed50e6d3a526dd5815da902016dc4c55137991e9624ab3ae7ccce535bcbd6aeb2efe041
z885f112a9b0f8a44581c54d9f42d5e440abf73606d4d90811dbc3b6ab5dbe4f50885ccc2ec1213
zd557683cb5e7b95133cddd595b35570902605a139e28f88064bb304a1f28580adfa15549fd140d
z72a046dfa20cbbc3d9f013f7781a546c01ee6791843ecf0a2d41755c3516af3f0cc1043cb9da84
zedb2f925c8eae4d4afc78600a5fc1ee5b49f9e514243b1fd6c3b0812e4eb9176f308ed896642cb
zc7d6d65334757eb51c488407a5af39c59116e77da46fd144101656e902357661ddcb6e908f2879
zb6e6105bb25d746d2bbfb83f4059a6b30ab02d7fdb698ba57c8ed3df9971b72492fb9856c24175
ze19a2d3bd006fc2255e6fdc155229e740efbbe091edb7bbc0596f5308921664135fb070f152c37
z986f396e055078883dcd75d02b328c44a59f527bd636920462a43345c3cb72285e4d1533380cbc
zc4af297c7a963c1dc0f0b4ceb28587913986d8bfa677d8220bf2e55cc88f16d3be3a9a81eaa0a6
zd14bc3742e3461132c79f962e5641b4ccbb246477b6e737a83fcffde1d9f898bde4cbf8c351a09
z3abe56e441cde3ccb75acbc30c83d2e41081fa8c0a7eb4b4d44448eec7947d40d7155b97799a51
z1952e35cb58f71ca3fdaae907938a96391c78974f6c778c55f307ee5b778ffe66f7dae251e3b57
z7743fe1c30591dbdcb8332f9ff0fe11698c177062230c0528e44fcbbc6ec66a41a94d86f6b67aa
z7583a41b7fe93f9a6d6feddb331b414b720d1aa338f1eedce3669e97974ec1f03e3c87f862088f
z778cbb0656fe002562bcf73d0bb1ba32cb4ed2f3f5b927e55e8119c805bc811b52094235fa56ac
z179a38bf50d671abcc5b201e15a1091ea01bd64b832536f21869da1e19cbf4cf3cf6a2197901b4
z9bfaae834461031c7d45b3af6f1a420f0abeb10c9b797573edce46342167a3dcdb244be403c883
z4cd590bf8ec8dba2a4972c3182e2476a8cbc6672395878dc5f659dad6ca65e574181dc515825e6
z0eebf4102e6e9feab7987e166023180d4bbc619fe76ca2115caa67b3b72f9dfd971474f0b5adf0
z56964e11a288afb80727b4d57507af615fd136ffdc970f6fe99e6ae1d6e0941a5636450f2d9671
z2269d5f931746811882293d5b334950eb3df144d7229c2f3376d34d8f5aaa3ca9affc168ba1d1d
z08a57427b706e95c5fa25975138b473142921ff8a3b160a465ebf2ad03f45319cab43833ee823b
ze6fcef739f85a92b4b9f5051717a2f60931ab66bf2c9d811ea225c7e8c05c863148896390523e8
z2bac2cfcb5c3ac7f3b3d73794dc848226cdfd8394b87b056e182ee45d8fdc68623102c57a666d0
z0579d96f1ab0d1b2f75ae40031d52997eba9935081abb533ef98d940564a652b7188d0588d374a
z47c3981dc575b08003cac5dec209ad3518c60aa6f4b85309b1570f4a817c366dd0b940afc7071d
z2e116682f60161e1e8a4366a6d0af033800d5cd931b758359f0607475cdf034c33d78a304ad082
zce7712dc3636faaca7d5ff2ec2beaf1ae734202ef153a3455373a3c25a0071816db20e3fe9460c
z6a8b917ac061537fe31b6ecf19390c3f007bc3bf5f0f898fb34274ca1372a319a1c4d6ab726319
zef8c44c1a148a72387339b5d4fa2997a74306c9341721ae5346711dcd255a8b1022d38017549fe
z6e13112f73cec9817742f4e2c2ed444b23cabd1e7dcebd9b82e1630acd4a0571027de25870c0e1
zb212034cfdbd5f039541b2ac40e10ae4af9af347ca21b5d23c7c7132f6d3f167a438acd7c374eb
z73d8487803792df3ce8a4998c24ef54eeb4e0ef9953b61c062157a96452c29261bda2ea1583d8c
zb73779e16cdc164c84d9762dfd9e0e16b69825a705454817fa977e99444faaa5eb9c3219b5f1d2
z7afcda266874bc306fb3751f03fda5994dfd976626e07b5efb6b8bf0f2087cbefb9691e54443c5
zc5d2ec0dfb5abd4fed4d0a3208e86dd041163e9b88d8a5998e26f02d55a2c56bcc4309c6b3c58d
z9ef9098c7f234a8bac16d7db6f2d82b8d1dbf2264d22e6764599d1fe205d5a3e00c94175b94ff5
zdd2b2b0b3d22bfa8a8583d4de754cb83b8a66749e63f9d2cbadbd3f8d67f041fccdca160659a43
z83f4c8d623e2050e2936bdc80e6a1fa9e0f55ad80a9f36064f4004bb40cabed53e19241a1ab849
z6b2d9c54629e9b3f8f4263dfbf353da4ba8c6107176d9e6d70aca7b740cad3277b8491cde62152
z72f18c3747ba959ce91281462527693f4b7c2ace671894ce809a042daeaa3d7f44e44f1722de7a
z61775868322e6c3a644ceb125f9becb1e38aa3471ebc20d00820577c024e60931a01f16e6cbd5b
z8eaf7de00a83711b4620d4937dec2f5f11f8056714423b6add35e85982a4c892a72d67e6dec626
z0e355702a3e750ee4d8209021a323326236df4deb19bb00cff93ef7dc096aae0ff7282728e5304
zd70183875cc86beb7896a6e41042bae55f709be38f5946bb22b12a5f452c8b3f822669a854b3bb
zcfb36bd4e4fc3bac5de940db34d5648c6558968ccc1faa30f5880638e88d69edd2c5a6b437ae6e
z80dc0398e74dc77cf059a2ec46939f85df45bdbdf9ad20f3d3c6e2649fe346a75a8ae25ba16043
zc4de640645b00a0cd3901b5cba9faea502f7fafe98f4be05156b111e84a621920e032317811076
z1220cfd5f397a5887b383b15b311cf457fa0a5550ac762fc6d167a9e4219f7e413153434fcb1de
z273e69aab2b2388661bfeba1898ab390a10255f485e44db4985af7899bdc42533a004e98e0dee0
z87ab4827044f9b499f45fd791032ebce102e7ac2ddad80064665597c2838c701fe2c2d3a93cb91
zb4e5951507be30285037c4c996af6c2c2249883ca375ed685cfba0110aca8d7daf61c157036df8
ze5685568d84cf8698162b5db948f49d32761b9c47b0c6b7abb2d129a5751f39308cdf857962b82
z9c2b1a7d02bf2c3633d7545b6e56c5093770801c564b231615522b8fc97ae4123ad685db9b9a91
zf5b5b6b14048f292ee5c240b4a032ef2f7a8a3dc637c5d9e578a76c4f7d374e27cb7ad257ad9ad
zd75daa74f00d0f2a4e602214cedf0efb63d32fa992be6187ad04e8c452322e4c3c965c5c00f4c4
z5b56ee3a5c276a7dc7c0a244d1ced163563f23b71ab27d2958623e5bb437654af4c7fe424c44d3
ze336785eb481cdcca140cbde4b23b3abd5be7d7c032eb8766f864c6cd0416202ed19b8f25dbac7
z85e4d0b58646e82fde6cdec30c496a04dccb3f40c2b0b61003707008bd355f2ba4b168fa87e9d2
z779b3a6612535d7c70163c20c8282152abc098f880be62250a7bd1c86efe384c789e27c0212a4e
z70b32bf0833bf0a2367c02e6e3e212bafd3de1fb10dfd61610b06a4dbe63a5740bb356b15de9d3
zcd6a53df468cebe9ef7b2f534356bbc934107ce83ed1ec9410a40dfd38e1317db79a68c56cb33a
z599213086e69eef53e13ca6bf0cec11facae56d45fe9b15b1f51c4e7ba9014bf7e7241cafa4107
z1eaccb1bf7207e44417ac3644d04862695f2ac02a3d9a44e68a06172c97d56be482eb4181a55c0
z66c62c6e87fd8cb7963563690c5ed5872d1ab3c2930713f7c4d3d1218b3d0f30211d26ce362397
z1f969ab1828d8e8587559a65c8185ee0ee6305e8843ac38265df93d46ab647ba001a5d3e59137d
zfe9d75aa7ec6aba49be504226af988a968c5b0c166f3cfe661b590fbf15070268ac2dbde6324d7
z0264a4db74585bfa2a27be2f8a1e20ec50623a893672103901896a216e5f8b1a4f9f396f80b93f
z515959398d1564c9865e922794ddcfeabdef789de79ed621a889a5aa7a553729d1c20c5be9400e
ze190207bae3c6336ec2a4755bce464389fed5ecb3e33248c6ac28d19e2043b2765cd343736701b
zebf25ff8f226d57af55f625c6629b765c73e35f5f31312a3bc9cf8f1e12408284e9dbbb0833871
ze9dce719159c5bb18744d3664610eb56b281ead5158538a2f8b04ff76840e885f2c83ac75c69f1
z1b17136810f0ff968f63b8598b8c5fe4ba16a3efdfbdbb0dd1cb4b37e1a358c6b1e983d9f1f9ef
z380ef4de747502eeb2f0ff7eed64a82f2c6a9ade7854932054553dc6ac574ab685ebe353cf79e8
za7e18ad10ba24fb399090a3fde45a9c3b14239f78b04f53a0164912814c5ab6ce08a9ddd8cced1
z2f114b61be178ad8d0eddae867f3df99229c510bce6725f199a89f62f76aaccfd04945619e6717
z6e533292136e3f359a21d2a98ea46526c49d0ea8fd6bbd7fb099d7e8b125b3b300c76a52d0da46
zc8c497c7a6bef9df7de1dee08903810630a15e8c4a528746f6f484e0603c15b943d7cdf8ae52f4
z2bc6caafe50da73c01bdee221887585401e4ea14f09a3e8e6d1201fc88b58a08b0409716fc0a48
zfc865fa86139adc025f0b1bb1995f4f0b0fc8acac51a20fe2fc177a31ec0b4bf667e3e961d8c86
z1e3139389b2489c4b6acd15e0d6d3f07f7d77189aa7d2bf1e046dae91a0ea2509ce2a7295538a2
ze688458a97aaeb85cfcdac3ae54f8d88c4a39be998a01a48d3ea8676db8bd073bc47fe70538173
z744d8ab52358d3b5ccf2d456ec96caaf664fb03c1c06977a9fc772816865340073bed3b3342cde
zdade2c50ecf068f395016fc99657b913e11aba9627fe82c26943ec98d046a9b1b2fec404f0b380
zb304b7b29313afa05388db5ecb17c2513fb244074c23170748997634ca5ea5532bbc8a3918e8e5
z4c180114b25088edb7460162365736609d3bab429a6420b87d4c3373fb4ff203627893f84f7fc7
zb05c6ae5fa07a47899467a7f72a43b3b3355eb2e24904053cb12627cff5bf63edafb275a2f7134
zde242b591aa60402848fa5f66da9142834c65feebb73462d61930b9f4ff414b1db225326ace19b
z721d71de01667b39573dd5242d6bbd08b66b31addcf6c97406c11c70c2222a71f80fbc2db6ae87
z687ee75a23b67686bec533b37d0fe886de9a5ab7ca47ee2f5c0460f79cb17eae73c99bd8ac7c76
z665396a119bc4d1763a458d72fb5a912d124ef070844e9b39d2be13a288c8a4348aeee02f26eb4
ze3c94d867f3c70946ef36ce6d88d1b2a4e51be22362db89f92412384a14f95c6ee48cadebfc1be
z72c338712568f976a146777acb3917fac25a286517fd8732f9508030f82c1da5cbf8ebb9334fc2
zbf872fcdc5ad4c3034ab4842ec12f4f45e5b5b5b2b7c05f435e8c86197e81b1fbc7f6d41ee9a1e
ze20e367d1f014febbdce68a09ce473d92015df48834918737fe3dff47405bf91eb22ac48861002
zca00d5bed64abb9bde8d35cb20f216a49b6cfe45a30facc232c15bacbcda7d23465d409fedcf04
z5d4429c7326c2ce117b659e94ee0e5afe340e25622b515787bec4a3be6956151114c087a390244
z4b88dde01daef81cfa411daf7d146c32663794c5af88bffcbf1367d76201313395f02a6777800b
ze2a7821b9ced6189a933a3eeee729bf8a274d1e7e6dc45fff6b74efcbe022fe4bfda0d9291f71a
zdfcd8d9d84d44fb4e49a7e6f87357fa494939cc3c3fa3617b0169176eecd91891e3041505a7ad4
z530d751b7bbc02d8b83b2d80d57b7f704aaaf29f217f86826cea4e5824fb54cc1c616a7ef7fa61
z94c7446cbf784e050aded5952a2c4e920fbc1e9ba6eefa327452568c5952a2064b8ae9f6dab7dd
z77bb311887fea55905b5386cf7d69573e7c3b440e7effd4872382b6d9cae8063f61c5612f04eac
zaa5bd56cb85de17e261a96e1b2ad800392d5e212ca548bdaf5b077d56719231d079595d24bc07c
z719f7ea2cebce1ebca33c2799de3e61284e678cf02cdcb0b5e1e1ec6d18754fb1a3cd2a01e541a
z6b95a91dbc9bd468ba83594c9f2022efc316a829bc140832c987bbf6dd3feb61efcfd8370f00da
z88c2b68bc9c05a35e3ad7427685813ebc8fe17f9cf17397513f6e576beb2dea5cd965b2531c931
z91511144e259b7ec4211aad0ea186c6b8e4a98689c777d39739b6dcae3aae39e81e3eb56c0c5d9
z4d408fa46f9044a80dde49888291df49a8fc2476f6bcf03354d2902afa63db888d9d84e7366430
zeb6145dcdb447bdd207e8104d279b543471908bdbff5ae93e5f9bb40b5264b2bc5957a3612a24a
zcb7574731f1620d08683d6cbea1d520211f02ab732b626c1b0b9250c6d13ef79c026ac7b05aaaf
zee65337cd28fefad067620b6eb81f31b44c9c5eb6b1bddaa10f8c25cddfdb87a6ece0c0d6c5c80
zcdfcc8888b3ea0328bdb55384e2d1b3a0aabc9766d3861e696d9bdcd20180907b56c1dff1a1c29
z34433cee057ef2f3db6a922e1ab22e9b05caff7417fff3637b273161397ac83c1a1ba4342358e0
zbb1994b9da9d0bf1829db7b8e0c9619dd6bbb96b4f9f2d7fcad23f3ecfe2f15fb81c16e025790a
zc2124b9f1d9a20371bf8ec814e84e8189a52c1df3a9c86636318c91143af61a90c347c5ce42570
z4d467cd964b91c339c9e193d8b09ee3a4672f5127649758a52cd8efca234c653bf69c76c89d0aa
z9c967882dd936c7b97310ec89c474fb5006e48d538d10c7b29c376966e0fb5afc60a7901b3d53b
z753912e7c248d4994d1b50e66afbc1422662b7acac38a0ff72a2bc7b601590a9efdf71fb7c0925
zb9403ba385eebda6538b3fc03280b9b802a49fb884f8e2c8dee5342b356b704f0a96fbcc79c9e5
z2cabb71678280c459575d02269156a85933f9b7265e3a9e243e2278d98152341c6dcf1715379d0
z5bd79d499905fd4b33101ba8eab529c134d72b2c8a11b389712b91bffab00034bec1cb942867c9
ze36a14429646bbed699a4489de51e5230f7472daed7ffea7d22fbf4fb961c133bebdc90f4d7f84
z752562f1322405e2a2d8d0e35c181600db85a1afc08abccaed62304258ca3357f08b3a3fa2dd88
z1183d1fc6009bbc20decc73d91427b6b2a72f6dbd6e7fc536798d4b22e4b235e2b2782d59b19fd
zaa0c0618da2b924e4362c446c6f7451d14356c7f66cbe126e36e045a62f43ffd3509f730eeba0e
z014d3235500a7bc83eff5623c5883e3a6a8b7dfe3ca280e18cf7af388359b43613b9531d31716b
z64ed1ef7f4d064c0689b4536bf6ef031b01fcfd2a3ad2bccf7c6ae8257cc137accd60311894372
z8657fecf0265f64fa55b62f190a87d4d49df8ca5dab74c77a57f9b6865eceba9e5bff36814fe10
z8edd84c2ac3f47a8cc6e0d10bd872119a27d6003f3162c649c154e75d358711406ee608680af26
zb04f5114fd0a1e74898367fe347a1528e544c811d50f6db82e1579745f62190b3a0071ef6c66af
zf845254c93a0b5b0f154051d446059300b45ccf6368fd9b8483b4ba63745dad32d59017bb118e3
zdd3ee02078104c5c767d52ca3be029fa7ffa1fe4088c7428d843c4d2953faa42b5bf8dd5aacc4d
z0458aa2d675bdc7fe80c34252d387eeb1d717f85fcfdad4c785a251f0ea7f185e8fef3aacb13aa
z9a64bbbd338c44d67c5cd7ed10636593769553355b50fbe0940899a1fa340e7c87c87afbf7a1d6
ze1a1df6101c8125a06ee584dfa4f174c6e3284ae336d8a400a35a93f4fbda63d16cde35704c0dc
z6599a3fb763efe8aa06912a68157426d8992c589a180c1aeb343e222e5f38fa36b06d734884737
z90988c72628df817a45ed5eeac7923fa7788e3c1a191528e92727789234f3bf9caace29f8affc1
z3780d66ba51913773153f6bf207a1c5f8512903b08db84ae047cd0e6d5e1413bcb5475f0259dc9
z752ad98b9fe09328c0b5f15e914b2ba847e1981a16e69529d6a94cb5ecc094351637dc64310f6d
za1602f0aa6f0a40f0509e085cdc9dbb7fb070e6eaa1f3aca1424b983528fcef325b1a489d1aa97
za4a35a604f2782fd7ada8989aa1d4a10d84fb89ec4bb79944118d9d2f7da9cabb9b05840476478
z2c64b62dcdbde2647f141b55c3f6bf456f40d316d958fff354d2f1bc8cb724ad1433c1f7b237cc
z8170beb150b2301f41647071c4978db33e314d48ef6a7ea2e267def73beaf69ef8f9cfeee8b366
z38d8a3bfe91bb0ebcf3aec2a793bf100f094979fce89d95211837c7fc32537805f1eb1d6c85b43
zbbee330751c6d6028967f6a37294397702817c3cc3077cdf9041964bf8cdaabf9ed95ae94d02d0
z7432bd541721a6bef853fd468e09ae9f162433c8c1d2f3a8d445444a177f48ab1e7a6c7f45c940
z5af8c1aef5f6ac2895c9c2eea68b1912836526a0e4b18e17a9ed3f028cfbd750cf1cd57076d7ba
zb2f0dc4fa3c2f67a7e66303c110b508d851737be317853279a3bb7bf8fd99a31cfc03cf8c04746
z3a651222852c14cf59ad383774f40f86990a86089fe53740440dbdf22abe36df162910be12a5f3
zcccc90018e98988a8bb0f1ba64376c10e7010485e254fd93c6a8977a2a41f020e50d00158360c9
zda7c64e7d850c3d1bfdd6c664ff0f4790f5127f931d2e0d478cf6026c0fab43d7a64de942451db
zcbd0f0aca539eccf4ac00f4b3c36de663668519de3d4e22e4d3a14517c5b0ee70ca8a974da03bf
z2066e703d7f492818369e9570aaf4f49d6bb2e8eee0c55a34570f317d4dd28cec1e73edf30db8a
zcccc5257b31d3d72e6dfe5cccd98482710dbd372d54f1f3abdc31e1f5714da4df42a751ebc5f2e
zf4578dd41571b708c7b03526a4d9936a844383bc3b2a7caaa8340b8bf432c9332e9e47d1c87a28
ze89f1941305338d2e1f2aef59e9d315bae0fb9ce528fe8d6b7b8fd48b57ca0eda83020d39a0fe7
z380c4fb6075d6e5d4a963143d75eb8d0838a5460a339c0567cf20a6f2af8e03046ee8f5384eaf7
z0cfce8440762df800748b6efcdd021b6a7192ba2720575b8d4a8bfd611e71f51ee3302515afb13
z722063420c0e73b50fa4b06506db1fd15cb6692fdb9cab395d25baf1fca55c6b40bb98181ad7ae
z2896bd9be286284b284235ef9c01d54ba60325e75e7c5e0855061328229be2b2aa4f5f72c23d64
z06a3b530f118c59efe8c1778966d2bfb339ef324ea74e90d7443578ea5028ca943ae2ea9187c67
z08b981c26b4b822824b9f7dc3fb5f0680e748e72945ffdd0f6daa4c21352e3143d28509b15babf
zc949858920f843d2dbb6783061886a699bc5fdbfb081df7678b73c34b568be4e018d8a6c4a75bd
zb57968505abba8481105b6c1e272e508950aa062d83a8d045186bbdfefe77a00c66cbcc25599aa
z2e1ecf245134e7caf122e1ec447c36b0797e9a2aa4d636dcda863aa034b9abca6b95a800771044
z7d9ab2df08a366de81edc19d4ccf7d939bc1228f6006595fdcf0b66c475313273d0b72831607ca
z024f15432cc7c0d1c4d0b51d16408166ae443607f0d8dfcc480edd24609af09bf8e2ef1d80b331
z801cfeb0cb98a94c50f0f23d6d8ab491a19ce6738125c89e64a1a5fbef29b8079032b3afafe3da
z402ffa43745715132b5259116905c8300a05134d5b7f5de6b1dfecbde10a38ce6860ddf7665c61
z0a3c936b530b7a1a1bda4a1c49635be2fb479ae7597215d7b4de1fd74f5ee1b4c5e8c91d5dc867
z9435d045e038922c06ba900020a6a94ad5134ede4f9cad4ea22f981066ecaf75629a4a51e8803e
ze189a7c18de6adaa179eeae4dd578d977aa8966786b469b5552d6b36d998995760a94be113aa52
zd54c0b9e78c012f58292f60c99d8915320f870ba950a8206b594c5c26cbb788d4c7821976625b3
z496ed9dc9786d3f3578cbe1aa71bb733feb7bef4d3a96ffb369e4e0c80389f16de123f7e518778
z4d4071ae8b6bdde891c2b8561bdb6fdbb40bb2ce94eb0f82
`end_protected_0in
`else
`ifdef MODEL_TECH
`include "qvl_decoder_assertions.mti.svp"
`endif // MODEL_TECH
`endif // encrypted_0in
