`ifdef encrypted_0in
`protected_0in
ze74c34e226135848fe16db9ffd31815111b6d7fb642c521a3f628cf6da949865580b22efd062a7
ze90adae0e65e66a2c36a587d0a790699161455169ed55a01f2084f11770a774ec4c588039b380f
z6de9c5084882a40b79a175f5c2114b2b6d78b070cb806e1c0aa9258297f4687ab308bc470f0040
zb0b1de382961eeeaf2e279e1462520fc31c119af8f2b214846f56c2b3cd2eadbe4099496abff18
z15cec83ec4a77b868344aa20ba7360908f5c0de2a79abf8b3534b883bb12180f68b5d4beb444cf
z3fba8f13afb0abfe8fcc4294810f75afe452434d2d0f1166236c82f76edf1e12979f04bc35693e
z32ae028996dd85737a8f5adc1ebb94f39c940246e887647b64782cd7ab429b0544c173176cede7
z01dfb26b1f73408344a52b7e1f117f12bb9c8077b34876c2e6fdc085981637012dc9754765e1a9
zc512ce062e0b8fb16a214591f5c81e1353b900a611fe1f4886b57940b41b7f2ce99a7b84b04b90
z916f717e73bd10589c81e207ed77ec660a8cbed5b487fa50acde1b055c8870bd8676023f21ddcf
z9c98cc47cfa2d654ff1365d1f45035a045a66c5dfa8279050262529d2cac9e64fd27d9c7de62a7
z731bc808811ded9016570962244887f98fe5440167bd0088f2f049df882af501358497c3b28776
zcdc5426c7f52a851c35106bb93e16fff984784050fc808fad15da330f6f0607eda2d0e0e4b1215
z2ac5b11453f6b6c5c6b428261a64553d70b4ab9f1b396e1048595951af798d8de75c23e123dcba
z74156e068eb331e95842c597f3ccd341bf87af84cccb15a44d811686c10b5caab6338f8bd390f9
z35e3850857fe16a4bd09a1f73b16fb4d985cb91a2a6e022108c6d66aed9c9b28b7bfcecdeb30c4
z21adcfcfd1d3a705ecb82a7cb228b602c508facae7d7277529f388f1ae749d3922daf9cba774a9
z7a2cdbe51bafb7233b5a04f9bb9c3d371ea04be74069b3a4dd10e4f6c35c82f6cbbe0454e3724c
zbf1e895fbe41f8493682f13f8ba66c6752b72d8b80557bcfdc43a34729a2b9dc7b8c72f0159ac8
z0d0ebe827a33d33f251768439aa9bf24495e1bdcb4711553f548d87fe8795529b32395e9d7267f
z12ec53d5137bc2b4477538961388818f47f4719f556358d7ecac8232a83e84ae4caa6f52486cff
z46559e9c94a0dc63e9b6e5123bb709f0a884f9386a9fdc25d7930225d3b0582dbad84e55a3e41f
z60a91f360eda72810b5d65214a328826b6fad412743ba4330adc7cfc90408b61d2db5817a89b56
z303522a61bd236bd56e744cb15e34dddbe1dc92239ba36b643fdc6b24d8eca107e442eeb2918a5
z66f2a3f89416cb1eb2a1d4c07ea7d2bfbf4db240295cf8dceba320b6f12b20d47794ff0dcf06b9
z5c3541707b3688e2f0a13a3ae2e17aae57f0606fc15fba8e5cffd1c61d8b2c5e9da926133c4f49
z122f90e9c6b24b2f099d106e270ee558c085de8e06633a6534997009cc04fd9a09bf7a53d771c8
z063ef5241bf70022af63af82e333f4066fcf0f785704e493e0e7e348f59269175916457995a19c
z801f7423b32b6ee36539bf386ba5ec0eef132ca65b292becae830f8fe20a9719034025198d56fb
z79bf728228952d0df36a3f716e21141c0fded3a218aeb5fc252af538468029dd789279914a959f
z726423f67575e5906de31eb63413a9aef15b6e476cf45ac5468efa82b553239bb7f5be9d77c068
z3d07142ea7ce4a78c837c8919019c343d966d6d1e4b071426620c7d3dfe139dee2a712ec6fb01f
zeb4538ad70efbbeaf1690c4781af517940afaf508ae403fb8d5fb589011b3fab50fe1442a8c851
z12adbc4f9a164d003a4c21f2804b6d3d3575e366b1330931ca934f3525d1a27abf354259dd1508
z2a5edd63b592a778e56b5a53428eff729727a91f8021141919e24f231113ef7a4b4a59941c0c61
zc5775c1d2f04991c2ab4bfb6d6ee98ffacb615d55eb32fd8a82e92d51f6fa695b497285e732712
z73a7e8fc367d72a996bc8838cf89dad6a312a3a7b5a4b5bdc5d68412591451062f8f9a7aa64331
z3f74a51998271a30a2dea582b6032a5307a3663dc54a70c1a7368fea2c7fe36ee5bc4712e2b0b3
zbbaf6018ff593f1cf0584fd132d0515abd487f58218527588642870c243fed3dc9c35f899615b2
z8a9092eba6f9f0848a010c19b4df2461ae2ab77385bc396d36349e57e79881cb0944e49d7d287f
z5af9eb177fd7cee334c826d72523509a26de9d51dea931346b0a9c577eef830a449c2296168f67
z874177cc3853966618fc1a11a939b50634838f393ad846981c18e217305ad4a92d1aaf59cd61ff
z33f513709db9ecda507840e21eb49c9c3a1fca46304c6771ef93625d9775016199ef25dee62058
z3b7127cba257c87bcb56208426ef1e85dd86434761d35059fb121ebd9835f92c4bdec31afe96ce
zfdf6f8ea167505f7e4b0bfd4d52400581905fbbeed130594eebc83a6350f091a1f14f18da0007f
z6bc0187d34cd63c5c9f640530075bc8dbe2e4f7076ff68d584dfffd8507cacc4cf227447667e5a
zc4debeddbbb52fd10380b3da959b3898fd41f59490184511056402d6319f914706f40eda320287
zdb20c68cc3f687a416a581eaee39f7457052d2fe34a3ec25232294183e206b29bdb35f3f46d99d
z47848f0e81ec051cd5b9a3f4d6e212d85a2b2d05978d058b15d23d56b716cdff2a6c7767c59cb6
z1d64681bf8693aac8d6baee7ea722bee3aff36fe353c890475191d8cc9e0f916bf158aec596c80
z0cb431a3969528f6ac296b5bfa690ed5ee8d7fc858ac3fc8fc8330bec2c9d2382a6df2da390b20
z2f5db2e3a0880602de96551ccf5a55c916f8ebe6aa6bda150ab21bc2782d5feaebcf5587c4d10d
zbae04b9143361f06519426b9f222bae12b742def3cf7a14858f0ba473ec8f158b68efc4fea01d6
z9ed092e981c28b8ca7be2f784a16af35d5da1eb525ff817375adc9ff04282760ea2ae6be858c7c
z89ff2279eb86f93893d6b3a0bdd1340dac59e0b86868b98fa01224a4b275c05df9d8e6a7cdf8a2
z804c93e51ee5c89f65ebf8cceba0440656abe37e30c51d57bbbdb381d1d41252b6193d97fbdbbc
zda2b7dcac72a07b1d32e957ff2e514a8efa20d0bb1d3ab44194b1c38e5951e793b10e55259cfa8
z7cf333b642193a969abffa5e5d66e100989a9e6c52425a77090a7a7792a15a7a86b483b353d951
zb98362a8c1ec0fb4955eb0ea9dfddad3607089bee0c5e83454ad9f8904a505c925398430069db5
ze00bae1e855c2dbbb461c955d1b35675982ae9589ec2d15636d4dccd4827e51d13b61e800176fa
zde02a19eac4d1e2f9d2e90ef6c6e5afc7e837ea31b8fe412a081f0b12230346c5000a74720df3f
z7871b4ced55344dbcfc58303df25c542040eb65792aea070028b9c5c7bc9f1522019683a1c9531
z7a2506c45d68d988b35fc0c9db04f6270856b722c3f802189945fe3306de1ef514e3d412c2eef9
zd75007f0450c6431c91874b7b33caf9fd62d76f427db73451990ac469e7516ea4ea226f58573fe
z1534879b5bf659cdde8d2c5f61186f4da949eaf0c53ac30b1121669bcd87be2df307e26d3fd8c9
z7ee793ee274ccca597b68ee7e101919fb14c488cfffbf768af147b3923641a3d4df5340c6f2c78
z0441fe885bb98b40f694cb3bcafd6b984678eaf6253b3596b552387c7da5ed7532bd1c74e9dd96
z88afccc1e716b8fdfdfb84f827fd344d77d9cc3dec6e305b4b7bdb1e9b631df200f7df9ed811c6
z65eea8d01852cf01fa95f766eafbca9fab2816160a9f3561c35de13966375ac3eed714b8c0e8b1
z120b02d5f57d5fba4c4be2f51ce67de57f8148981d130a95b862a43a62229986f636b03516fb32
zcc674cd24e98117c84c97cf7f6646bb900b9b44270ba3f81685ad1b50ebf35c928e0ba4173ee93
z4f06b8acf33061b38baacc8c96cf3abb61eb7484a7015551f2a5c1a932a4fd0aca479dc0b38dc3
z3842c3628f60a804f7a011c766ac07c3142a8c6e1b9f1537ab98053491c1c554fb5b070ca3e6da
z973925659e9f1968ed3d616a4ce57e58eec31611e92cff7f43367d3195935acf198d86b92148d6
z020f529702e95a844d91c35eec8b3d53b9be5df307136bd9a8b2acd7246c3a2f6bba1ccc2cbaa3
z8d0a4cdee43639cc68d0738c819d654a563ab7cdd107c5f21940410b433a6ffc9d162b857e3bd3
z302f80912df071db12ab40047f6b5e1d4561ef53bcc3d01928d98767af04ce9d53902029c1e938
z149c450ccf34c6cafbac7703e02d9e203fafd9eea674666110b70adb9457563238ee93c3225416
z8d42fbdc07f798d05f39ccd0d3820e5e4a8eb5917e8de55e2f90859e66d981c9741b3cd1667352
ze82f52d7acc9e4fa54e6a509aa67ee934e3a66e5f2ced6748af4b626a22c618402efb38c4d357b
z5992edb5e14e00fde220e52d4a916bcaea490b3abc504a039894ed4f4d34a56af42991b415882f
z33a33d5c6cb398cb2445d73b44c026956cf7b6bff581337161a9cdb53f6cfa3da9fb88f7bdf46d
z2d24c2a836b5d3d4646807cd26a617d5eb755c34e5abbc46bb295a69fba964c14dfa8aabecd16e
zeb3fd5e4321195fa9f2b312cf01da4275196af4cf3149564f98f6e37a326a3061145286df82b0e
zda409385b67aa2d76291b9497fc8f79b7815fd7978aa0993a2ea111cdac0d0f03565910977de8d
z465e57a4bba29b51188cb3b25586a9f071b50de0ac5cbc06c2559fdd83045215884de6f770956e
z1a77a5e6f3d4df8060f9eb34bdaab038e3e6bd6c4cca6bfd85833e89e3141fc6e5344289058d6b
z0e3f2c3bcc7c43e4ea4af6caa3f6dbb54322706c019fb1c65ab2d3470fec6aa18b71381793becc
z8be5f55d96f49170b5b330a1aa4a37f2e6e0cfa26455b8bbbf1e9d5fc6f0f914b534cdda30dec4
zbcee16990526ea5b9cfe22e270971561616528f138fc635319e8b85c8097c2496f6d8d85fb9562
z8397a056130b24c3cfb4de47089db17248b641fee3ff190e671b8a1e9b54b3dc92da5df5a9b2e4
zdb3a23f2854a7932000ee1ab5b6fe76eec93123fb22aea550a76b6c7d8a37c62deab3875c9a687
za89a63e4d940645b3e1f4d4ef188b9b7249dc0399cae16d3924c0bca3e765eb9c54a37dc39a121
z763d59d6091c70330c2a3333ae18085dfae2b0e9bfbe07d0709d68b35eee365931d5e9b03a4f46
z84b76e117a72b4a484fd28231f5f74a0365aff892aadc2ac6c130b651ac35533bfa04019fb5313
zd351a071c0245498b8b2b4ff7bddebfb23af1f28d315f24665d103399d91f9a582b319ab52243a
z81186074e6452d3203fe1fd46e071a0aaa67dd95231c7b8d50c17c7bd4feddd814d01155a04a05
z4888269f183a69c5b5009290d15efe4f76968eb5b2b44a02f7b059e4b2da68df3f7f5410d71b38
z8c7ea928b2c02555e7cfe3e1ac1c98d151f076d7c814198e8b4549ab485fcbdf030fea5172c646
zbfec12480e05872a2b4cc34eca482402ac738554aa3b6d21434559d6da43be1d8932f8732040ff
z15add3a15d7bb14e7fbf5c89d4e7f6e81d76a8b681191e4412940219b84daabe3e911a5950565e
z489dc75bbf47384e0bff45f85638ecdc3a1cbdb24f3b0c0c172669a8253c27a51c4ba862d2047a
z77a5c7f875284d9d0f0b01df82f9e3ffa7d479a10005aabd3b5d7a725c9cf6c6069d44f67bf2fe
z6796ae5172693381b1137a830323dceac62c3cc1dc589afb7ef75eb31627eab1d57a93cc1cdc7e
z0101dfc0cc26e31e935dc73305684c31bcd013fa7f21f1a89a22fd54eff7a3dbe55a44cbdca4bc
z508f38a2f4010b8f100a75b7855c0aa9cfda2188c148c55a38fa705c3bb653d08d49b9c941317a
z2ba1a27517b21e78299dcdc29c25d4335953c3e0e46d80049d5853c523c784609f12c567b61bfc
zfe39aab8f83c577b6fc14da83cbe3fffb47ecd0ab2bc3714342dc44e21286ea9e394d7892d20ad
zbe6b711478e38e128b3949228a3c08869bf80dec6c82f4e97c74267920f94212de4ca0c5ba625e
z2e93206cc4a68e2147d7c3863faafa71a8e28305066e034ff9898bda4549cab5dbe09aba765d8b
zf8f31cd7513685edf4dce37396a9a31ee55c5ed287a0b39db7c4ee2c116275a9e76f4124994c1b
z36ca8e3504da5fb48431a366a5786c97a486aafd74a1f4846921aa3eff89014e6dd4da3fbea6d7
z010d500f6e309a57661328cae6e9050b4c1de1c9c846ffd1bf4e07da6cee7d7a30ad3ba32a485f
zdff71bf704421d357f86aca088a43fd041c2fd18e8f853d50c7c67b56af595561a53d1d69698e8
zf1747e932c6ff433f4b1dbc2d1b8f10e286b00fcf7077c15b0ec2b0c896dbdab59654e5d3ae26a
z556562cfdc0ee1b848dd7475825b94763aabdce9673b21eb4bfb494aaadabc9000c1c9356b8219
z95440491446a0f11ef7d820a0d7151594ac25c295cdb454e395f57ed77885b04453712e42e6788
z67ab7e4f2e2cc06cdb381b19a47ffd33a6e6f2418e62cd7a93902fc46f936f149ed78c4becf3e3
zee44bb0900e9af1799c1b9c4d2b87105b42a6b409f49320d7af5569160ac9c77514075d939edf6
z0a6171003ca48ec26513882783677c26c8c874260c2fc6ac5f099bea881079bc1049cfffd427f3
z3b1e910ac3ba7fa817a8bb2b6b24768575202b607a89bfcde69bcbfc3d01c2e6b1117f58a16312
z01f1338e6f70069b34f01a9210e94d9e7e59edcfbc289bf5976881ea00d6c184486ecb9ab1124e
z1e40465465cc86b32805295824e13ac4f710ec5944f6f94934b62fb1840f1dc94349091fb55df8
z572c1cb596cfdf3994fe2bf3ace0605b47f2dc654c10189fb8be5aad7c52cf12a3544deff1960e
za2dd58fe3211a922276e0e9ff08bcc2ca369583c958cf254a24ebf1d68707503bf6406fa640cf2
z1ed06c4156c15ec51d37ce36c86bed5638fbacc62384679e5ecf5aa3ffdda7cff95c0a60299d41
zbbcfcfee02aad025c56fcf39586697c50e84a2d253080725906f30541ef7f43c1bac7f415613c4
zbf8670fa5e146044022a03f46d3c4150bced2fbd7816e8581999f431a80e267d7c2c9257984026
z4c013afe5edac4084cc63a7a5c5fd1b078d06c81e6ac0d3ba76a710c3f9c6dadc683c672b7fd6d
z1191428507febfec0114e48155f047c0df5c4e03b2ab46174d69b14d5171c485bf509d2b59740b
zb1d8b567044e2b54b0f14ec8da910254e2c14dafefea3c694487d4edc77b735907c399232780d5
z073e4c2228c236714f264b3b8a55e6633421b1b38cbeb6ebb2fdc86a8162a34bdd02414ba17b52
z02db24af77819d3f2fdec5fb8c2e6523d4d49eef30ad7f8cdfeff6c442a13ffcf9031cac3c9e3b
z0bdabf60fea5dceafd6a544f9938d815e687553dff54619927b20fcc64843ef55cb40b639cf6e8
z9aab4ee1e72da604a12c0502ba125a8ea5f383d776875e3a6bf2e9f84874b90a9dbadb0421aa47
z4a4ab081724af5e6a1cca846f9cc9225ba6d045e598817a488148ab581b62f3af47ed48aa1f8a7
za2d69dc3dd56e300f2bcd880fdcfbaebbf5402386c84d31aceb16a5dd76d86250b4da596007663
z6d5b02503efbd4ed2b016ba2b4977ac322ffff8e7a83c78eead2c758d7ff5ff652244b6208048b
z8b6ed1887f75ad78d2c49248c2cedadc2f006a23515e968d9a15923c97e59eb204810d5ede91b1
z53c068deef9dbdae20af2fe9bdb73ea81842b5fd4718699499288dd664227346db1b674f2c60b8
z1d296acfdb83d65fa97ad69d736a624e3b938707778944afcfd9c3c25ed8eda1339e232d4898b4
z0ead1a8eaf65eea26ea6f11eb0628da71bf55c107cf1c8188c51928d9bbf0780f708f36a6410ae
z0510cf9589425ab5618e334f3dcc56e8b5e17db91b45fe447f7c94b8610e079fca3bfe06b60e05
zeb731259a589c0b266af70b9169206c5ebda48e327828210f885ef3e791fcd26d2215ea88df58e
zf0cd9d84e0ad74569677d37b676aab07d44e3014f0d08ddd1f06d1a989f0982882cfc2f83d6b4e
z2cb6bb257c49a3e32637729b1cac6c045e98fc3ef7320da30430becb517ab268bfa20538165efc
zbbe2472e84ec44f0467d2a0d8c7d33db60a39fb44019b8ca6474cd8f3f37ef9abf0afc88aefc34
z727f8372637488feb5354257a2be7349a1a247849a9833cd0b78910e2c432ae1c6df1551e6742a
z1c660f5834e3227bf90d0c56bfb75dbb76dbaf1d7d85717d3e88881a4e00c965b8ee06adb913dc
z0873c2bdaa2708a039b58178c344a432b5f9d1363187933bfe5c19ded86db7594edd9c678f621b
zfa2953ff457c08665daf88debc0a52adff8f8961c93e575b00c53d6b8ec942483fb097c495b94a
z34b3a8895e71c101f1dd8be811eb7618a51f807cf716398c9758073a2f4ca878318cd3df0dc1a6
z8bb3b1d93a56fd2a9b5369f60abbad2ed78fbd739b3f1343489cd97fc6bb12d393d585fb205594
z64eb65b4f2e5ba32ce91430adf42e5d8b189c5a62a2ac22e085e103fc88969a845fd319705652e
zc357fad02a683254ea0397a0c0d36d84a1a11a6f72d0ddfeee1b9186a98c772a82154a3ea8db17
z7560b4e938e4dd0ccf1f810ab655f614e573f2860477407263087bbbd6c8ee0afbf8dc21cc8197
za3e576700ebd757f0382313dbd353103ba88d9c278b1d73c8869e369a7f7a04becf1be676a3459
z16a921bed8b27167751015d6ddebf5917773580e40d56c2b22b12840c8c50ced20fec090c4067b
z9419f29ed00054deea673c8dec26e3167790549d4f763c8a9d066e1cc76df396d91297baec3e68
z74864bee78419aea764e62eecffd3028e27de1fdc44ebf19ee0ca5d3eebf1b729f0247fc866393
za1fd58db68ea362cb971a46dfcbd82cdda37e86715e2291e96eb330ccb14905febc250f5e4f901
z0002df40c67f8f2b7ccb3ad79c9edf2dbd855655863e01a40941184820b9674d46264d7a3eaee5
za3857f7f5476ffdc3a4053eee20a5e3159bb5810907002f79b2e15ff02a35cb67d3ef1fb84c70c
z87f982fd55fb7ebd4290b90868fcd5c494f170e06379ce88a3b21a9fb11bf28a5dcde7c6e9bb00
z2750b018289ec555004dc5c8bad7ba4f09e46ece59a289f8a607525afd7d7297ca7225294c44c2
z59191891a0a929fe5280d6a515943b349d9d47484074738030d6326e470d17fa58f799bc4fb476
z736699647ac9a65d966038314ddb51644c50ffde5e40312061f9868cd7eb47778d7bf9109daa68
zf9fe6c956ca8a202485798e2ba6815315b70c52bc25aae7eb22be90b44e1972196f0f76a252164
z1c0b5058e23fa425db9605e37559ae44622501b20690d1c0e22398327fa20276ad9d94962db835
z4b83dbae21ed557a037f8286d9af85577fa6cc20f006951980215ca1dc5b9dac3b78dd8fcf6a3e
zc58bf4715b6e01fb8037932ebc1c0a8a45f18957fd0c1f4996fb18c5da594ddae7a3fc5972cb0c
z614f52819bb4e95ecfc4d5e12228d0edb704875ea09acd36f493ccc6259477715edafff47dba8e
zc71743be353802684c2e54b5010571580a56bb9fc8a5543a7d28f4e3cdae6d13b1a45787c0494e
z8f55168256e024e463f5db36709b194983be7a5f64ee5ac43eff4f71a5e7ecdddfbf666432b9cd
z3edd1df1edf40304d3e5a64608334329b9415a580d3846206aa6f9fe9c86125078e46fa0b8dc64
zcf296cc72e19361c1b95c5d0d4ed7622ea0d72b9182357c63f13023cd9c6b98be966f8a934ad4d
za8202228ec22f3bd28bc7e69b53202e836c7cc3d6c8364c63caf3a458c34143da213a43883343d
za5b082dbdeea1db73f63b1aa066cff06d02770e0d77e7a2b5f6693c7e33f2634ce9f6262570cbc
z118345c0983267a19dcaef4c49b23d301489c4fd47773f774b1bcdbe18be0d4b184016472af876
z54b2426099b4c221711b8f5e3015cfe88782232adc7d109fa5d03d727ebe08ce8b006a75b6176f
zbcebba161df71d3dbfde61a288f8b02ee759eb937d5d404847785ce7ad8c4fa35db90a39ee3956
zca3961f794bff378ca75cdb84f3135c8bd28d74607a8bb6aa37d73064ee1adf259210c5cd7b0d9
z37321b64200dab254e52c34b39b4aa280c2bdd379e6f5a0c81c76b2a031681ba715b3ba37421ea
z6c8a9fcf9e80ade62c6bb41c081a186945c841ca4fa7e2c447bec7c966c881ecdefb4d447b2c3a
z393203eebccf02c30ffc54421c07542b218ca935eebca4c898eaee68cbbf36967170c5c8e945b7
z518b81a2ffc2d37887c796ec4a229c92e6fb21c8286452702dbc3db5ce96f96cf0d3f56fbfc5d8
z7aaa6e8e611b3d558e4d1929ce56f36bb82a6442ffa99ffbb64c85ffae23d1a1c96066caa87bf6
z09b8afccfaff94ae725d289f860cd6cebbdd35ceb3d0a704e044c9da0c7fa4c95b8b2f02a3688d
zc66cb47f1d4fe6eb3cd1a7d60c209bf00b1e0ac141eb389428d11d5188cc83c64abc21a8cf4e57
z5e7a5bf09e5ea0eb202179bdbe724421c55e6fd9220889598e7a90ef49b12173ae93ba631f8cd8
z381f8f98d1ba09a54dcaaf4d09cbde3d54ba636d59d76a6b660509f8d981f67856bf3e3cfa5db8
z8fdd439a8fa2ffbe36499fb3877f03f232103f44e16766ad08007678f06f3d72c4b08dc06f7673
zc58811cab7d21512327a2398b16a1c8c650f040c89e2b14dfa34698826a5845b9e706e19c730b6
z78c5b44f31f3f32ad938456fd0f45207f79932543bbaaf6272b0d67af78bd5bfaee3a97bd93b81
z3bd6cf09351d172a46adf6297d4272208cbb46b115893ab7f3884bc022d7747451b221fe8bba9c
z2d76e23572d7ea412f410c388ef085a11faacffaaf146649934c6a4f52214891a611249ae124e6
zc6ac73d15fb39bf1851d5ca7bbff0c81204e3930c66a089626046eb0f5eb534a5d26e10b495339
zb402b40ba5515fdcded7dd1908b33421b6a301eaaaa80292ab4f0a041e65e728053bdfd86500b2
zb7fe56bbd1e7d77b1eb16453dc3f9548a7a374afb6453cdb599d342669822de768802c5c50db5f
z48902e0bf7f3fc5a269ce32e88847b9e5b626cd149dc3d938392d1bc49cb4aa2f4b56106801cbd
z8fbf5c920f5019c89570006263c3c176723000fc751b7290cb6b316ef150b84402b716bc7af47c
z25bdaa620e6ebf60f0b51ba58c1ec87e49fb284846e809906e7e27131cab42794126c7f8942f9b
z44bd033da7a0806b576f8448487c05e480a6096cfbc076d49d2dad7642382d58d234ad6eabb86d
z0dacd51388c245903691007ed4b3aad87151a61269685f49c788eede78d745e6466d76d04c272a
z7ab2fe6151f6233e6af562012f486afb97b981951b3db3155e49520e4a5dca8306c60b7d73f531
zb4e830269862c3b5f9d9a00e85610f844b9e629f0f912ae35381af2516a501426b1309682a12dc
z2a17d8a2a48f2cff7b0feb27e59dd04673b22fb0fa0b5e2aea66c27ab68057615df2492dba23b3
z41fb93c8faffe6a5fde6412998b61d085fec4ccc8db18e71b4d4f677245ef92362f8e27f4a4e0e
zf4e84bdbc1113b74494d781582199216c2e3a395356d61860defefea43ec454cefe05438f470a1
z37e4d5cfb90381b127e0895c40e04683693eaae44d13b345b70f7e42905b52e5ee41db1b5f9246
z7b46b582979c15ad872fb35b125f2c8903bda5811e06ee788761a41de1031cffc48ba41ce9cacf
z9119d3b2058fc99ea77633321d1ec614118d4ee36b2dbccd09d7cc1c2c109892d06bd5fdb0aee1
zce7bca8ecc82a3bf662872a8fd78db293187b500abbe09187f75ce533943d6227323cb2ee6a8b7
zac91b5ad876af96b389a821e5c5e64d8002eb31c0826630c04e5b2adf13163cf433ee1754b6fe6
zeb42a75c9196d4f199f399915f2762d282e770f997e1e4d658a7e19b99b21488ce92dc21599320
zdbbdf3b35275f7cc23a5961a5ba99127196d6bd17825b54df15db2dc9941df4f4226c3bf7741e6
z2573aad1943ed06543f5d6525366fe56a6e63b01a53f253b5f8ab9075fdbc772546d7302b3fd7b
z96aa78195a91a669b26b651b8b81dc238d02ec7472c5cd46ab297c2ac539f2414a936cb35ade05
z1052fd6daf45f48ff314d263eceae9126ec07e522ff91561c5d612426a1ccfe8dc3d89b8e02ec8
z514c549cc0d590b35bec90ab6c58b6006652631fecf677f2390f01fe4fe17aa58bc8db2334dc7f
za3a5ac6796e74e32c1646b8d0836e88485bd621cbab4d291f228c86832fe99df913fc490e0394c
zff6107b9399a6dc277673e1d01894c9cc3a01d534327ff78f469b4e6781c701ac03e8e73a2384d
z7d671c41b1588afe36c23b5a4c072e3ce30c798fe451fc2af49d64c65d693d66eb82be3f12773e
zba457afe4cee34186907a71c4c45de4255dd9e88eafed5227550a2d93d9b74e3f30abd1712f985
zc5f43a677c90a28b8b3f7c8e7c90d627a01dee7e46746a7fe8ad1040f7e3df8736b147084fb34d
z8ead619010a274cce68e610860bcfbb3a973f7b532d6389f2d21fad29088eef6134b972589152b
zfcbd8b275a1811cb71272088983bc368fa047924fdda6267c3948c59bd9b7825c40361dde3dace
z208b9ba3b8e2bc351937de4f11790dc0b95b35b97ae0b8c52fbffa4ca5071282e5658c38c200be
zfbbed039e67046d04b3f78ef93bfdb0bc5a34356185b3674c41133b8c670e07288276c1215f24e
zbb45b9232e517f7286a185e2bce0c9be0f875964dbc39a5234878d981a175f99a7f0587309c5b8
z1bd1ad5a53231f28ee941ddbec79d68df3ade7e5f75617fbfc451d7dd27175506278079bca78de
zbf64c0f1dc35f5bcc88bdbebb481306d52e0430d7ac325977bfaebf60c96c0cb0146131b377cd6
z0c07dfa05e96276976fe692a43c96310612f76a3dc03e2aa0a77c8c2e81a20b185ce3b4ecc566a
z698412f4b6b1a4e751f60b5cbe2a55b3b38b32eee405ff96c8e782ca96a23ad4f4146e9f5486d9
z7d9337726c3b9c4c8ef8cdb852e06beda1b684b77cf909c53391b78d4f2031cdbed39f356fa6c9
zbf5b0c9727b77cf0e736830e38218c8ddf36c1281b7677778158655e8533ab5f738c998414b2e7
zdb523cf72921b8ea870a98edd740e55056e091769feb3cf2b10b84defbf9d6a4e1ab46b4ab4913
z6bbca34ef9cdc2e457926338a5cb148714c2d465d8a345cd265095f9037bb47ca86af0df1dec60
z0732676f6a853850a5da6463112381efaffe9ec28f80731936139653f0b2beb42fa19656a92b5f
z656dcd166861d94f42708b2e7256eb99331a2988020b62fab90b86ef31c39a124284fc379d31ef
z849d2672f1e11d74b325d78bc74ccdfefc16935f788bec50a52d59eb3380a4a10da06e5f24119f
z21b77bfe6b1be96121fbe1f17e12a4d7cb4bdff505ec1a4ae63c2ab056166e8128b71f0d097bb1
z49389e6f38598407e7bb0e8c1ea1cd8229afb35de9d1f271fd65e2322f8f47a4e24722826669bf
z9292e46ae87e678ea02de6279407ddb30d0bff5ec3dcf4e418eb268db8f7399d1fe474d94168ac
z429819cee05c5328c05d62c70873cdc5f05fd9517262c7315b8c3b11f8dc2976bda9853e05d17d
zce6497b1b37d0c142ab5f5f450861933f879d839428bc26d6f892d31bf3af2a3e60fa26ffa04ce
z506c63a8e11045189195ca3816f72b130a10aa35a229b858f2915d673476cdbad0bd679b262639
z31bfcdaaca93fc154bb62f06eed5787eef26d78b3fbd4978f8aa55f38480e83bd7eac8fdad341e
zf44bef7454d03e9d95bcc6bb55588855f5c197b59254c10e3d7921f2e89885ecd47ee669dc3385
za7d79535a421a8772a56707d616bd2e07eda331af0a5924732ab75d866723e2a5d579180c15328
z43c175ca1e5eb12050ab9362d57693db41b84476071b569d1c1e0767c297dc439fb09c32a20579
zb54f30376732adf24fcb06c1024781ec15315e5bd6e8183780cee7b35785bd0f2e2c141c71fa62
z89d289bc78850c7ed0c686f4f32c3b4f0d2716e16be4f3b25959e987fd5a3416f5a3a0150dc8ad
z4f01e2c79997a8a535eed66c988d52e28b4e448759aa1c08da92ce6b41363f540f30826047cab0
z16732e63116ba9d92e0411734fec9144231d7b101ac65419adb6a87013878026841bc52bf43fb8
z4c7380cd28e2b8050a73d06ff009c25bb41ea954075edfa772379ed96616ed9769567f510a9c45
z0650e9082c2fad1564433e49db7c24e0ef379d7eedaa1f5e2bd671bbb87a42836c3300850bef79
z8e223136604f2711ea5a2f76c62701635d1eb1febbac810b230eba64168db4212cafa7d296116f
z3a097b45ce82fcb2ce595cf3d20bb676af4bc8759d0e4a33e34237df000e57caf762810e6dbd9b
z888b4ebe9397893cdeceffcf5663138028c70a9e6e9ce6b90ac7f784636079db36f2c9844b4a14
zd9257181724b5c56e2404d57522409fe858182530cfa98701e89d34e38f3b3c1dff0840e7c2d7d
z2d521b1bca31e3c27e0e1d540b4739e84d85b9a5d78c905a00a48051b20d742aedfe43f1c2628c
zd87c98fd5692cfe3ca960b362616ab11537a081128e978784a0136462a6272e60729a0e0449e37
z2f83e4d009129fc14a047a56a21d4dca594887709349e53b9604275f36f4b19caf3dde166caf59
z0af413fb6b3f264bfe328c6f2b6b0c694e34d7f3e883c57adea28d6c398c457c626c6b14810903
zca88b8e57711f8551e97e61c32b0145a4865d328066932e03ee0c9dfa2636eea0bc1e09c0976dc
z734a7377b86a075f076b14eefd765b2c437f30a045c16f2b9440a3d9455af254561b15fe1d8178
z04a385c5435f5a9f95fd94c318366802c03ba27123aa380788581a4d12e17ff3b503318600311c
zd79f15da11f0b61fab7025dd6dcce2ecd203eb82266dcc93f0df3c6470854f654d7d6e5a979004
z907ba6276795473e0d2b415c2670b808a322654ac5e21af99961a34cb5242f08030c12912565dc
z7f40a0bdafc9af171772cc298af9da888a0c96a37925fbe88ffe8137ff374d82fd7ded80e025c7
zdf17ec66977b2a212bacaff766ccc214d67863b22095727d1b16c9925bcb03be24140453482360
zc4ec8bcc677a40612890fd4b1eec77319db092cbfdedb8004006884f5f0a5fec8d005b464b2102
z1661a10c83c385df06e0612d67193c87433bce477feeb7a4dcad21fa5bdf8fc6a563d6824f643b
zabe71d259441af18b95f665799ac724c37b0e1012a7864a60c8d3852704b944fd148a4a9249549
zb1d0b484917f2aaea8826b3a9ddbb41505d72076ba5f63f7d9e91c009a71c764b9e6f2c00dca71
z4232b7795b83eff3e2d64b4948e97b6b25241208cafa80cfffd7a19a56e1edf995b2337c602830
zeb77b0ab665c4558961c85339450d1c2649a9d40a7e11ecb96ccacba36b2f7cf8ffb230049b386
z040fb671151a42879970ddb3c75918ad7e3ba5f71f0ca9eb41b37e6e1a131a0559c418ed7a8680
z36264b8ab7929af63355ea6283095d45dfd7d49fdb46273a1aff45059f9632f7f211229fe74744
zb766dacf3dba65651291b351a262ebcef44c1999ca4f6cc2ab1d3998a558d8da0dfacf08380486
z3aa46646018c7cedcffe66bb0b4d8e29fa17844c78986b0cca42ad9178c78998caae244146dd0e
z36f48230b2977dbb67bc034433ca30fef4d64320520fd980ac3cfffe0354d261726a469ec03490
zae752f580609912ac0963ecad05c03d0b72790bf90a4674196095e33a2f26d60e50ec60828c226
z5b59ac4d6f4842629cf1fac32fc3cc6cf9c7327016820a9c5157905489b9ca199f1180484ed19b
z145dbe42d88c77c0ac47c0f5d3861f92470db21f5e33ad5d4756f09ed15341955783b24a1b9a3d
zc738983d57e5352fe6036aea631a66ce0accab9b99cea82b0775c844d512416ae318d2f04e82aa
z63e3304354efd588e9c7ff25f328332bbe82c182fa3f72b2d21b70b9c8f6e79aac1c5de2d0f64d
z2145d67d6b67bea693c87bf4bb32f69da830cdc669bc156d17fcb203b52eea2600076f9b989acd
z2b329a19d516cd86a76051162759b5a12802589694fe7f2ebbb6934f525ca5b17ce66e3b9de65d
z27f41e20b650bcb69ef70daad59bfa372caa5a38c15b6594e0c3446e51110665b0b1aae5c70a95
z128c62218a97ca446e6666e825d213d3b53c25b37241bcf01c82d6939c0f8a6508743aa55be698
z13e6f2eb4db5b78b79fdab3a6e79fc99e36cc2592c4d911ebbe12a3237b00cff0c3ae33d072cec
zda711ad8e8399dae48f4a9bce85b8f6929ea13dc44fa4d196762f75bb49f986d1db3eef64686d8
zc6435378c929eb75b0a849142119a88fb07e0d4633b2f04b02369835b6d5cfc61f781462d8330a
z037bf9b1d89051320ca38232ef978b2b0013a5ffbb02e2272ffac75a27083d1ac72f54e34f9765
zbb116528de7f93e302dcb36bdbb403ba24da53d4b41910d04689a0d66d391ccb3b1f531295c17b
z99442b21a832f50d4ad98499ac170a6b2b0144fc269606464824df6b137ac6644d80237e8b7a94
z577e93ea8b8d5df5a9f0201b5f071a51a6c5d5065f6cc4202e442c400296080afa8a2bdbb2576a
zd0f0b93ab1374ddaa7c11bc64bd5d2ca214f7b888401cb51567c2176b92b4f2a2b4744cbd612c5
z5088f58c4ceda2fc4528e00efab3da9b15d55be6e3d0d4f07a334ec950ef4fd4da82e5d54284ea
z7305efa70a233d540555890131f5ca39ee95846d41585c7b16c573c22d0b41451a5089d6e5be1e
zc2e60e4fc436605185309318a3f0b99123d93f9248651994a6acb12a727372935ec1a4846656cb
ze54343cd72ef0ac8a452006af03f11a3d853868434ee516e582f3b1b9a62962ce70d493a52ae26
z125f7b592123fb6a9ca714e377ba9272acfa1106469dba48263abe06266e737ff075292456a5da
z7a6f4da01d3e0f7dca8db47fdeecf4cacf22e3108d42f3fc57d9908c8832f86036feec3ecb0d8a
za7b63268db64f6e53af566aa4e48bf595a2d3bd0c6af7a846909d6cc35997d9f0837604111812c
z07b648e189dd5343f7ce93e4c4ad625c14fbbe7a755c1aee3b2de340f7a3fd02b0f13cf736ba35
z6a83505231ba8135c760838afacaf7e9a4b0d411557eb19750255ac4c9ccf9acb01a44fc0b0b73
za8c895336906976b73bac22c9c1ea3040c362b589e54b82577c4bfcb0be41794b1ca6e0666f134
z5e138174866f3297a26b596463d51df9ff0e5fc59e91645aec100b804f813b69029f4baa0edc22
z5abbfd87095d84ef6554ebf5c61b7f773d79a756eeb32cd6eeb6d75f8b6747333698ac30c95b8b
zfe6a71a7d2bc163cf8259eb2f8870f9dab5c84c004bdfd06a86015e65147d69499fc5d597a3f60
z127d21f51986921ba2069509281679b5741eb7ff24afd25d9ef8cf741436553a69fd8421818d7e
zca77020c6b7effe8c4a6d6e2b15280b70a3741418da43ff94f47a3631ebf0a34cfcbed147b48a1
zc2b121500c35323a189d78079cd9fd497e9b07e37b870cd8689b57ae007b62a4fe1e40fc7af1cb
ze65d2fbe039c1193294cc37c3e4708827047401a48054a78720d522a63e10826bb6e0e68e70ae1
z4498889f1d3f82f333fd901a4b4c0a6424c7d45a195d72f489004a416a6ef2b801725161a53cd6
z39dcf2929479f5f251bfdb46a2406086258aea3108bf862d5a33224a1fd07e7c7d21287222c8b5
zb866b9b1e14eb70d6c00c7a2c62c1ab8a0bba187de4e2caf2cdbd416a5e89b23b4ed08c9aaa93b
z9cdb5023be2c5a9bfab4ee7d9edae4e84789de16e2fa693563d35e1ca0fef63a9d2cab02ada4c5
z593b4c4c3bd659db37a7a363f1b0d840a35e6892738686e8f3a8fd245c775fdcb88f70fae658e2
z4e2ca6186c468ccebb302df19446f1619e9bb8671865b36b6a6668184fbd67eb99b87bb5fa1570
ze00a26684964bca603eeeff545de3710c6d4f2bb769847597af724a27b7fef890549f894617fca
z1df6f5465084644c7fe2dec58c2a56a88713ec05f30f48a03314a9a8dd8f72e54b025759951518
z904593f6a8aa606e3aeab536b49ed3d5f7f9c74e4aa7a87393325803d51b2abc082a3e8a867eb6
z43b0d448940f3a0c10f1a08e4ad517cfa30c29f1a5199fa10163a36fca593420bfdc91e4c30931
ze63a61466b4c8b3c1676ffb2fba6a5ec1ef271ff4de4ecc63b0eca43bf61a68e8105ac62bc59b6
z06b793259e175c7c9e7857efc4dd37ced929fd852476e7565d27948049c4a667c42841e3c339ed
z4c00271753af6a62e6641199e796a9cde7ac89dbfe356d2439770ca377edd450f871b0793803f2
zf2256a4c92b19440583053436cc51a2a34caac836b1f6dab460de65a1ffbdeda92daef20b3410b
ze077d81b03147a32cfdb678ed5d6d874e01888acaaccc94ea1176327f28c35bf30ca921e4eafb0
zb9d4596c8fec3503395024b455bceb70b0e2c6440614ad4ad9d5c39ba1238b4831f1010777c186
z475a1355e428a14506c8565016b120ca46bcdb5b0e74bd359b85cc7410e5cb4b321b036df66c88
z0bd08b6cdb1827f6a6bf6b83fde74feecabc36ce5484c04b6ac33cb1a474829855a8f87003e09f
zb8108758b61c3ef6dbae4fd023908945ef7312bf376e13c88ff367eafb9971e0e85e93fd194c42
z5a0891a211b0db21c48bf3f9719fc5dbf5f8dde74dd4a1e43eed854e52300f1963e256cf9fcaa3
z23c10c8270bd3a3d68a88a7f0509097f0d08d7919bbed9895e78a7b8a1341abf1351b7c5d1f361
z90798e4c3a04e5114ec8ea74e6951668db3d386c9e9c1da83350b9607b1ddfef0f262c9c5c4b9e
zb546aad9aa285d5067e9f3bbb30f9132b6a1675b0e11347f27c2b0364e23bb013549f52a5fbc9b
z069a775f6139be387cc609b3f86c642a0d7822f0eca38024f45a9ac22f05a0077c43ae6abf9e6e
z5437d295dd7e5c3fcb7ae8d52267f7b7e7194dd66b42cd26603c4b563cfa76d8764a064dad1de6
zce00e33c764f9e8214f1d18b6d488db37514ed399ade1ec27172976b2fb51a76ac1a0053b6772d
z74a02a49c1afc03be8a3b4c690bdedb984891ab9b6da8ae043dbb4e5a697b7b2191ddbcda674a7
z155356ffce5a3bb0537c5d2a48f1dd9b2ef03224c527776bd821da33327cb83a766709cd85b731
z8fe371551308acfeb0d9eac38a64b080edc9558e2d6cff924927e14142edf50f06f5edef6d6cfa
z685342f8ca190e0998276356b97d08489dc4e60540597722ec82e102ce924f4a34fb1e00ed9a80
z8d15b9920c977b101de3bc4a4a349178a0c0fd2ebbfa8dcb99b72b587526c466577727a30b2bdb
zdce9631cadcc2dcb1287108efd36f75f1d9403db4b1c1f1b7ddb0df768a41cdae277597fbd128c
z00b833af07f4de9e1e3f72eeff579f3e65e415128ee954141c32d46fcd6578f2028b9da6bb7042
z9f620a8b80b8e0316d01be9d08d9e670a76082860a692703c29fc35a32969b31c05a6822076edf
z12ec42f3dbdc7a930ce71abeddad1fc46a3c24095c11ad622996519c4d6db5cefe4875ea797383
z03c4702871add4b5c992245204217dea4fec305dcee5aa959bb6a762f494b4994101936781580c
ze4ebcfe959dfb2ff28c305a52a9594e8d36893231c468bb11bcc23bd9c1f35dac86b2a28e9b15e
z574eceb73b7cc4a8a7540c7aaa5068688d152d29f554190067f5f0a3103f26252d7ee82fa1d9cf
z95e3e333935be3a91c2a19185c0a3ff9dd18c692fb8fc58894f0ba883738f45687098a7761204b
z7c5a95eb733263c3a73a021d2706660fa0c940ff2e21d9c7308567454bcd9e1da11b4627017fc2
z40d69aa96db6500f74eddb05c3c239adfa0fd4ffe22917f5ad4c053f3b43f70123cbe044aaf969
z748d8389405a9579ad198ad00d6126c778f4c0f7d6a6d80f8dc4e3fd050d303b0823c6cfa19b39
zdfb25e7b086f9dc7516a829f34e040999c7dc188cef4d13ba4b6fd1eb5c5b23d887a4e199c721d
z9f909fc17bc4e33a980e3c1d41308f52c80615816848aedc34310a7050e3aef573a1727a103e94
zbc8c7d8251eeca2a87781ece096313a5bb44f19319bfe7a5fa8b6f47efc9048ac175238395ba63
zb6d28a4f16d5b4e88f4e8883b30043379b4c8dc6b5b86df759585b21c8122d8692b6b8ea35d3d7
za2befc1b7465b401e2e107d4953581156ffe840576a538013c523be0f0bae98000dd9b85ba57a7
zd99d90dc5f71218dce0993b0a120c51015176634f3ecebef4d24469cbb1daacf1ce42dd000788f
z19c0b409b5d4cc247a0aef7d503d317d5cd2853c1d20c6097de205d5493865f15d3fc3e0463cd0
ze02667e9fce02a3d039f23d16642620799a75f804c26b5d7c9b88e6afd305c4aaf06c291aac75a
z6cfbb0cb068a5e116d709c949242d381363aff9577bd83a6adcd0079123612235f266df6bae768
za843c6b5fe136582dfb4c5a34a543e1300e549af2f52ce2412059565a2cc3ced415d63b8b19f38
ze0b11470e2068c7594db932c958528e703a24fda7e036a97d48270946c9c2508c64d615e70b487
zab38273a5a2506d1d6ad3a20f247323e8cd15ccf78ec39ae0fbe6fd78fa4d16430d85020fdfb74
za333e788dc946e410a4a7e6470705ff800db93b9eafa5f06150716f38571725e0ba09b74d3d19d
zc09d0cbe645446d660a0607bfe08cde6844102c690d26eba6a36b5d22b636b34a4bddce8c65cc5
z112026b4826628913c3fc3f7de7daf61b0791b95f9931cf23f217eed0849370e609407af254c79
z9d90fb1a5271344bf32a85d100215346364f3710c0d45c60ab54cf09d0dd83fb1dfa5390f81986
z21fd6e60c1a702f44cc4aa87860447ef8b5446d29fbd0424be0383434f150cc2c44241bbb77599
z6b3bcb999a2065c0969256db7d45cb011a726a73e3960d6ba15513087f1dcc8596de0d1ebd54b7
z612f6c4e0f1948ab6947f5a4a2dab1ea9cf9c796e2648d26217bdc3fdc65b62dec4a5428f57468
z0ff5d16ac5b3ad9b15883b9f53cf324f25c27a56c7390e6a8edc2ac298dedba96ec95426c3212d
zfded867b86bc8f5aca91fda848d812622d496616dfba543d6ab9b3399a6412f453f037b0c01c7a
zf61d88856c0ffd2c7b958c63ecf47eb95951a7bcebfcaf216e40fb180d1df753df9091becb9ac3
z5b49cfc8ab55888ecca935d52d2e2ed60f4467e3068c3003168e697f93a0ba4766235810d4d543
zb02e036a9f8444d45e85d84061bbebb56eb88bb9251d055bbae9d979d6d1ba75ce3fbad4ba1a8b
z6d22cb18d61cda3588f1c440f68d4dae16d84033a4c55fe3daf14cbee66ac63c41d849cf1236ca
z074270896bb3cefaab6e1f3125a992f1cb1f57035d984f8e086a7990e34d57b47566c814f2a7ae
z5ca1cf6dab84eb9904c1658f152b12b47bd2fbb0bc8b073ed565e90cdd54d5642a5f2fadc20f2e
z30b2ebb7a92a89af563a37bd09bd8cf32963950c67d3efd1d1fb4eef3eae82ff7274bcb80a4792
zc927513e880d06a240092702da1e702344392814bc05bb4c587217b612f6320126a65daec0858f
z3e702b7fef13cf56d679ba5a2a2e228a57d1fb2ef5f2a8438ec30e5e121f58047170e3fcd25b13
zff70bdf4d722e9afb74cd00a33526d514db61e52be82945fb3751277caa1744cd20d3054505743
zaf6501b101f447e9c873228a0c5e7d9bed4d30ab1210283ef5de4330eb913abe3bed5bda4e3c60
z01b51746a08c85ea205d23532aca787544c71d7cd58b24eb3cd5085c88fce6154bddad0ffe881a
z9131daf67cc5b10a1eb6f8cd837a1c12a2a3454227b6d77550ef353888bc28d4560a8dcfc9d212
zed3447c35330b60c55a61f5416a5a31e9df34d32a8f52d9b2c7b2a379d4f758cce1ab3bd09a88e
z7a5dae4145f5b9bcad422e07b9d28f7f47d614877c983826281277c38118c4d8ead92bf3c75f59
z60f354ff576c27893b6fd5fb56b391b7558d46206eb6caf620967becaff97e106e52fe24209882
zb6c2851bf6ebc37d1cc1fd3e09aa3970286f24518f51a6b5a1d987bf16b532b2721f572b7f17f8
z6a4d7cbb15a84d03b9679563d894c48aba723aed18efe6346ea37d02b6861a1455b29de6e1c07f
zdbd4bf8f753c009ef3d0f03374d5e10cbf7a17954b4a1fa0906586450c51683dacacd6a4ab15a3
z3b1cfeed55095cb2833fc5208d80531bd84df2ce71b6375fd3a4dd7e597d55739cc88a6f476d7a
zf9527af421dd8dd6f37db755f847be7d1b4691d00fa9a27bd7cd757f8a3cf64bc3e0acdb543dee
zdc23c900a9873ec22b8f1dea22013bb72ed6ca2e416c44cfd7d0d72028425b80629d34c9736d2f
z5a224a0d1afed5ea948604a53d3ddcb8d777fb6ed0ac7bb309ef63f6080912f5b6f8d0307241d7
z3c63d4d8358948e85f5f367a49e9b97baafa6dc9f3262a13193981fceda496f7dc092ada443203
z5b7be9ce6d9bc09d838c7987cad5a2d9102ece163f36389a89513d9b04a7892a6e96df8c8354fe
zac31a25766809b7d9afac45b6a6ceea38d81681963214638c766ba086194a71381fd573d816359
z507a7820c187f85ca9ad056c85e6fe548e96a02c43c7500df455ddce16b8307762248b5813a080
z1895c8a65553efd6eab36838b4ef8ea667f2e8254f77a9fb4a9143c5c84e3f84d01b69290164c4
zb55a4552cdcc3a5accec4d62dc4edea4efe6e06f92ee6de2bae4a61b33f098ac0a85ee537034bd
z55f9d7d1d6f1fa4fffbbb8db59b44b08c0d6f32adba73d7e2b9d54e78044b7a6198d86079aab99
z72d64cefd8c9d3720f0e72a6e61677e6d174bb3e143ed44144c9ac1ebc289e6ef519a66dab1afe
zbf69cb1d518e30cbed3995196fd09c66f93f6d6954e628355d5228e25a83e77aba3b85af895795
z14898c32f124d43233af262a9a8c3ce1c02db0803c9e735859dc4ea574fe8e86dd65e8ac9909bb
z8b657dda52c6ed1b55e6a4322df8a290f539601a95e14a4d058024a240d5903943e29f2e6da772
z83fee108f6a132815e6a0cce0831b47233da79b11b7887a285bc1eae0fe3b314b4e84b0b5e7bfe
z43cbd9e6cae26183f26e94378f60b8148269a5039a90d5118934357645bcdabc926593e21183ca
z105aea05f4b5ca769be988c1b86c75f0f1c83cfa3f2e94eec88c720d06ef1472f3ae964fb81b4a
z9ef98bcd012622d00a5db8e90404a5949b3630ed8437fd8b55f0203ea1426adb1e7c13e8e377fe
zbb117d00b94973604f9ba96ffebc149643858109192bc7eda911a8225cab433ccd1d5d164a18e4
zc8fb9b2ea0516f6ac62aa5e102301d46fc36306f0324d4e4b97591c3e28d28eac45482c851e953
z635a587ec1516c4cdf4169849bb293881562dae1036ca4a7566949ba74ab9a9b84f2f6f9db0431
za8fdb5c4143ec950d8d4359ec4bb82a4490a10ebbf230e16dc7b888d08ace4062d7f424be10db5
z505196535cf350b0fcfbd3ae3a642b51be29ec08a15522b9584f114fb7b503e7770522e9a55fdf
z3068f7454772c85c45995e0790b9711802362c5bdb11d47e4651fd8b25f3c5ade84ec7eaacc1ba
z14866cf1a9f4089ad2635a37b0e2df24f8594d2b39854e508c90e3fb4eee7e17c299152a3c1076
z1fca6c2c078cceb3cd3b160cd33b4c39f2fef880c28096f8610c79c9e817c106df43546b4e7483
zadab30c4ab1e044f5aadf52416bfb6eaf643dec27e33c15ff666728315e8dccc760bbeb1aa8c50
z8165d37aabcbabaca8f417d396fb306b2c8c8e60544e3b9d6fd32f3b2706954a41557b907c501f
z592896a6c459afeab2675e0306daa048e68523af23e8a02e0b5083783334593991ce98071683ae
z64f15e007314b9a8517ea5d9424eb458d6ccc913dee70a0ef740481f00d597ffa356f1fa7f899b
z2bcfff4a04c6b322a5c2ba8a18a5d77d48a338ca76f70e1ce189752691c5dd380d3e74582af0f5
z44fed56d37bbe5550f461f381f24391063fddda939b83f5e2ed924ddab38fd3b37e7d5f370e687
zc05340df6b7e187e3caee267ae7cecfbc01d4229098de44dce34a8095692e3eb784c0df2995f06
z62c3e72ccdcaba7fd931c1502b9152e6d929d870960782958e58ebab7aa0d3ed799d116c59bdc1
za0c98e5a6032909a3be242687bf6e54d4df19611d7a653fd150f236d27b425d5b84f61ddaaadba
ze99304bc3448bb97f0457dd627801de8a18c64434dab3abe45478fb333beefaa05bf13ef544e3f
z579cda611203b10b8ccaff08f6f342f383ccbd45a03f7a13c10adfaf72767b04674d45807533c7
z1cf45d073ae370aaff35dda189048a0e9634fff0ef42159f3ee18122717c8adac582763887885f
z15ddcf3f74198f2e37e0b092043c695784212fe90d9a15df8f259d02befa70b009044dafc3b2ad
z3de1adcd9e0fe982888b23746376f0315e87860e2ef387b77401458f12a325fcdf55df6a7489f3
zaab558f9e12f4a6588352b9c3adbb4934156b3b719bc0e7afd2676b8086ee2ed6fb314e53e22b4
z834b8a0c8747565b984037af2fbfc4e7e1c261f8ef5d9d731a513a44da2f96cc9d765dc3256484
z201834c5f86d5ddfceb62f8a1818ef78725e2a61f64d866277202ee32ee943fd5c952d8e19f945
zb32db8e06f26411f88a3b56ac5cfca03e99756781258534d60adc9ee8c98a6a39e4245e164a4c3
zaa423a95d9d2ce0cd9e43c9024a6570362158f6aff4251b2f600b12c30eb93a4494f4c9d2e94cd
zccf7278a38785c3c17e00155129876ba889eaefa034c60c3378efc5ff892bd4afbf8921a2cab9a
z362108f288e35df3645498a775994ae057ba512e5530bfc93d46012d337aed3f0cfdeaa815c3a7
zfb8623531b200f1875fc9198502307d7200f86d817db95adc4618e607584beeb01505c459ef03f
zf2a84113b0a208ecaa0c2b08e41719367374c2a085b53e782b01a17b8b91fa6b40298e545c3a97
z8ac478ccf1d01170992acdb62fd63f87c44f6e3977aaacd745b7230a9c1c22a3a481a456020591
zd9d1699dff161bb3948700be2be320cc22db05b70499d5d27e666383937e312b3140f12467b8f6
z37029081b27ed77d341aa05c5dc17f011a43b25f8fb3d6fdb3f4b2f2db70870b5b6fc45fd1448e
zaa7b0b25a03ac63f0a426595691d2f06c54a0906941793fd75148f0aa1f28d6b2c03e45225d32b
z6d5cdcaf495d5e1f387ca4defdee817a61164b84c22748db22c61e9aae5e2e848c5d0943d1395f
z592851b3476f2998cfba64f5523830eac445af9a7ff4cc569e109ffbc53e3274301d9cc6850ed2
z03688acbc37f0238303c3d7f07c92790b948c2f18d75add092444cdc8f75e18db9443b57f6f86f
ze43768bf6f7dfa4fb1f5393994e33af9e5504cc41eada63f16853814ff5317fc525a60a65a716d
z90559db2182dd7c99507935428ec9e60212e62ae06be4aa9b9859cb69eb2ae0edce674bc391f71
zf026f67f34a27c7f62caabb6c4c5bd23d072bd9d9158195da8598debab25e90e140241e3cf59bd
z62dfbfe48273ef05555069546396505c9e305ea20db5d594550f181dbe67f972965f1d18749d59
z069d95cd3879ed69c30a7dde04eb2bfe9f53cddad806f340fdfd21c3ed0ca341a7a86709d11247
ze091bb346baf518d45ea4c5a7889d0cb7505cc392c932f58d1ffad97601757f1b562ce5d933481
z1d7c52e6f590895c809bc7c1e4f2c3273e184dd933ff517f2c932d67eec842e823d06155698c4f
z98de1a0e491b33117ab4696397efc5bb296006499759cc61d2a2426d9a776e284072a73c4b4824
z7e42f275014fb845d87190dff6fbb43cc773df8e66676f125076f4af7679e0733debf493df938d
za80fda9b9ed0e08dcd01869fc910d547278301989adf18c9a4de463a04ad8bfc123d949c1d8587
zcc9f42dd253af8c2702f24336feb8cb7121466debe1bb4f10749ecceda5a0f1533c7d2f9766310
z67df395bc1df05aca85e43c5c33db2a20df3be808b1f7cac0401a12f89dec523d3cfd53a141955
z2f3b3dc87185b6d89adf017fe9b686c1ba7e276bc4a4f808e124ae159dbf55c2c810a0d33128dd
zdc4d94de3c15a21785056bd1b65254f4378930be262cf38c2512f55c0ef3514ee024d995906b07
z31ca2d883157da213342452262a90a5185ebee3a31690d63d7400b2a57c4fd21c356bd8dfb00d9
zb18b336a28d5a2cbc12bf365abd65192ec6433b58ac94128426e815fa086ee363ad903a9a4a976
z480e08e7b5c4b191dcc54767680f370ee61f050ebdc7dcaef08569f99c5ac0beb534a421b30400
zab57a85bff60950cc72cbd4ec691b6e7cf698584a7a3a67390df338a6696cfca310e9262103ce6
z0305f1255e6753f9bf1fd2bed5b30b0f3ceee42c1fff8de84e3de2435cc6542a160b4eda35c4af
z0cf4b9c195f99d12671db1e0d64113757c0970eb6e59bbdd9c4fde493d89a57156bc723bb3e6d7
z7fb624616315a7dfb490ea59df40b6bac84409b3fe1c79a62c4360692a8133934878a165efdb2a
z2c31d54351f310da25975379db874713930f3b20e9779733562bf0d487edd33612e759354aff51
z7c2f9ee5d6ea35899259b9e62b4c7ca752f9614a9cafc477c004bd18c63fbc54089186ab27aaa7
ze2597d886c4204e68386cc3e05961e77d4f079e78afad308a631f19aeb5971c8c7ff4d01b85685
za032973c5ae3668221712c38f47377b059f46ddf91a15aa61e1f82ea5f9cb55796e98c0442813f
z4c5fb874a1477c14948aaa583ab1b743bbef6414a5f44a86091f79b2b2166b9eb3c8a85d90a226
zf8b0bdf147678dfbf1d53a841b5cf68dac426bae9a189496c1326c608cf27a3f58b02a578c83eb
z47eb61e8b7a98dd107bf796fa23fd611be6b150d0cb4687e6d46046c4fbcac6524a453160205b8
z50b65977f7b34248af48cc1c7e97f1bb4ad6eb35e0deb4242d0c2dddc782303305734e105f96c9
za25a40cf195b89e553ed0dc0fb8d79d961291ba172e9c8b21fdd68167960b3dbb369018e4fa720
z740c120114f679b0122105362de7d2c716b9eb0c6627ee0835db848448a084be61bdd859da28d5
z3c6d13309283c14b6ed153680171c7b33400a63e8b85a8180d94a4697cdf5ef2e05e1855610efb
z32b7c791bab5cb05f7259d498359adeeb6a544a3ef7f0a68881bb48b230e664317de8d248d67f4
z68eac7c2758ccc3503a5f5c44ae05072e23626acac88b52449df61cf94c2b5d1f26118757c76ec
zb0cb41870d7c0539c8c010f55f0018aea92286144e541ab4b8c1b7b39ee7ac4810ee09ffefc370
z02a0055c03e99cc890cf325bc29576e02d052c917adb36168a07bd84a9d79e8e94990b30d8dd37
zd7d7c6dde78804c7fb23dee9b7f3746c5054fe71a6db5f15e6b51a8aa8768029048077a9db75af
z3f1dbb037d938a33cfbd92dfb5202b0a0f1092546d9ef60178fb988731811f2c7397de3f86e93a
z2ac3778077ffec073fdc06e18ae452b36fc54a8bd4887d00e71c9f4c2c577438be9f16c5a90ea5
z2ed9bc2f5fa0da01050299f55e0c2af9ff2a43fd0f28959a109315acb39e16b83b29f3187b3e70
zeb4a39aeada8d645490d59876e0dbcb5cc94f5e59ee07e1cd6856036ef11c7dc88104a87bedd3d
zecd155987a18699f92f0e3d830aed79749a32fe738ae33ab6693ce1ceb43321a8f9c4c4b01ef06
z201fb95436f1650daad34f29753352eac0e81a233c436be22d3da8f09b53a26cb2719ae2adfdf0
z980fff6e0e26378dc53f18e82988aabde86d525c6080a99c9be2f4068e266ff6afa0932f55989f
zfc7e07620615dc12d1d02b8800f1cfccd3355501f785aa15242a34375b9ebdfc1947305509967b
z0dfb0edfae33f492c8dcf92bb68f04badfb1a6d7803bf91c5a63f26b61e088260590b1dfc75771
zca5c9c7f181d8ef9a105fde84b60020a393ce7b100233617250a0c731d946d47a167ea5d7992ae
zeedfd73047039b35146f0cd40b25cb8dfd381ec44e6bd3d2bf04b7bba2a395b0d435bce2cc08ca
z258cc3f7f41d342f7fd29ff27bb0cf6953af2f9cca01f3ee5b207ab60dd3dd70b17a57a22146ed
z78eb5a73f7ea388a505d83320b02a25c1f381fa2e0a82989501df4bc7c88ab9cc34c7fd35cbf82
z855fde0e5f8fe20967c38a03b6972582a41d03a85da6dd0a4d58843f3eacbda1a5fdef9c1f985c
ze1241f76bcd7b89b00cff2497ef7b470238018c6f96c3868c73a02dacec4f9062482d40f2cca0d
z4bbf83fac791a0b81b05dacb5d2e90f4a6f52bce39208cb72e4307256b735e92fbbf4fcf8583fa
zcc4c7dd28208e8a99426d396ebd86cb40db29491192aea4264ddc041d0713c4c36b91ce8982474
zc75ea42a2578f719f66194048affd044d79bbd0bbcb2136d96edfae8222a1ec1b890f4ff33cdd1
zaf40cc6fb8c7515b7312997e85c63c44badc4f0ed4a14f137d63ce1cc4d7ddb00a65ec3930099f
zef7d0b9cb5f10bc1074a00ae0e99d445133386000f3f576cc21cf0941f6eb0cf1cc562a507f423
zcb370b82a2aad3f7935f2231497e002480a641848efc5f86022ac9199b157504326df3feea114d
za465b7e6017ecd1d7d8e0c03dc090ba7c40754b4438ab9649b888691fd6dc4f528bf2414f2b25f
zc4015b8cd8d2f4046f55839e7c0c8902d525cb774c1d13ba8e6feee5e95fc275eac481481bf670
z01da07cfb49f5a0b891873e0597c7f75d881b963eb6645d20c90c0419e84fba706ea8d5fb9f452
z8e42f3842d7e1e6e7b5bde48a05f3bcb609d2e5be8ae54dcb823b9505eb762d267eafd0dbf6e32
z0dcdeebdb065055f1c73c9f218f579efb58a8eb0692156aa51bb1e33ccd269fd26fa58dcc8a35c
z4d32bf96c9581d1efea18766687ead30a9765d8f953b4861a3de26e13cdfbc9db17069e0ec5460
zc9d773c692b63bc56f8375bba97a93ef05030041c5bd26b49f36f2d26a5d1da564a202f279fb2e
z2d50acdabae78f4e0820b61952ad9695ed21971c9ca25dfe5cc32c74e3b830d78133bf113eea07
z9d0605b106187f3d8f17f6e6a7d5686bb8def4e622bf2470dfb474837874fe08a67f08c01087de
z1647d87b2ba74e71b9bdb4c2e09cf63835ac93561eb903006afc61c64185a314865eaa6c604b4f
zad44f75708a48b78805170d8bfcd77b9d00cea58b4296c134706fdf3d0b6647b478eb8ad140d7b
z646a497f9e8b1e51069f4171fb4f22ae675413147f29918837fa7d8cbc29ded8329b54cf1e1139
zed0eda98465f88913c8711bbd2b2e11208e315d7eea30445101b9ca14d2ea1b042b361a92a40f5
z258ac7044eb68e80d380cc60f62180195c903659738dd554785f2311227dc4b51a805bfe31d7a8
z5235d5af731f4d27e6243521694a4938b2acded2a21e5718665ca4fe37bac0358e95bcf2f643a3
zc79464007037009f49cc106336c0b905c50d17d3fd42c579dff5e9c1e736cb02b079611fdc2d25
zf46807c74e351b9683b5a3c72adb02cda7807724f755db6fe4f5e3d519d1402717cd38be45f0d3
z741ec8c42fe372fc991424b2f5efcc26ad608643d2fcc7021de56b7288af579dc90406724d86c8
zbf9a79460fe6768552418819aad5fffa41464058c18a40754cddd3fd0cfbb3c56adccbbe756ced
z59c5a85d1438bf1eb734f62b55d9285d8a7ca8651aae162589329c0151beb09b1c43765c57aa25
z5b7daafcd637d062a8c0727a09b1b8a358af11ff5673b1a64db23c857080fd5fe068c838d8033b
z75b6cd7cf09bcefdba3c74b17725bedbc5b063e5a7f5ab4cccb299520d1eef98640e547fa32d08
zd490e2b2d07e13ca3f6c8feaa200035782261087c899acd6715a2be3563df9d6921b4e07b4f56b
zee33629a37a7eff879dfd086d2f145bf50069cad99692d1aa2bb7be264e3ddf6564729296cf39a
zbfa4173f7d9e2fb49ba64712313dfe61fed52ccb52bf445fbfdd48d1b7cf9b659d146212476e8e
zf29339f5f9451a976be2c88b4f05c121081d672f2274e668012d4772bcecec9c0d43971d1dde52
z53f99ec00b04226d31cdda98bed818c27b8ed0a6d759d88d4c78172e63ca5b4bffe536d467da2b
z767681f8c47344b35d6c575f30ebf713edb99db9fd573f8a74bb3d16bb4f0471d0a3aa6cf347fa
ze3d1750426445c10befbb3e2fd81bea58eb1fba64a466d7d84e07fe3cdda514e37432b17a8969e
z870ad6a5f407c2b16d890483567855905468b7d8d856e93e70fb48e638fca015e0c15c2da4f4a3
z3580ab7812e2fbe3e0817849560ed5a48860a5e0a76bef156090e6236172f38186b75eb1dc1e7c
z8bbf4dc5fb3babbdfe4e7c23ed68e6430fc236cace6952724c3d1c5a38e05e716d9e39d3508f85
zb0852ec3e1d443e82737b2211f23bbc43e2987d9f74d799e97654c8bafa9e61e3997d449cb48c2
za87118603c10002a4c151ac6ef720c9d619a807aa0158c6179cf8cb4fb0ade093e0472fd29b906
zb10bc2d6f466055a163d1f546d42f70a928c617f4c21e779339bd9f7264112bfa8d29437f84e23
zb6635d84b98d38d922d2011d4e30421c66b159e1b14255da3832c1fda22823b2eaff506d76208e
zfa8f40f7b8e5c433272165d01f4fb7a7a248d1ece0bb02fd2927b2018c57218b66a65225a1c99b
z37cf048d7ba24e1b5672f73a9f30018192c1a47b5c390b1ba8ef2818dd650b5ab81933d67a72e7
zcd66152f233483e5d40580d560ac912c015b6b15f257dd1235a94bbe50239fccc39100a75c3394
z9496f2e5daea0c00d631eec497f8a70cabf2921b604f82e3d6730e659bfe05e90bdc08820464ba
z5402d19d1f15467ba793abbf7bd424e39c00d62191ae31bb4b5281e114943a172f9a436c676e9e
z460e5f044d110d211f344316dae43358c1da7e4332b10c701c9dabb774aabd05aa82e14978615a
zeeecbe34dbb2890e9a2cfb587bb7394a50d88543ca8757f9ac0a16b8d690d1a0c7c5036d71c2bb
z5137c00bbdfbc71627e33265d25c8d840764ab06ccb380ac82caafb97023f05a7986ba0ee32712
z6455f6b5eb1fd9e342a0978d62b10141e77293ed0c8536a349b7be01e8a9f5a9871d0fd3beb4e5
z4395c4f034e323b671241870ad77479e9350592d7d11bfc9803b101d7d57d1384268135711372c
z4f420773ccb5d0c5417a62a65b2ed3f3f80b797b87b7005003bb86baac68bab549bd3646fe1e60
zb639f4faef83313c4502fde670dca86077326ff0ebff64371e8ed1d4132b0bbb1ebbb182cf57c0
z67072138f2bcdfeb8767e353586214ee7378c7705c8e8e1d220e2cc020345c44af34aa06945b98
zaca033e1f63208257185acef169ac10ca22b5e846bc1163fc4b5c216d22ce67b68483c0086d0bf
ze541a6f03e9535f53f8844c833f89ccc1f2bf1354a22deabefd90ca6953b8791952758bc1d4f84
z194f01715d3e62fbe5e87ca5b5b92a7b7cf2ed770d616570ee68b29c2c55a6d18f168ef7e06773
z70f8aed474c7a41f68bce9eff32bc651b2fd070fba9bd66860b34ef54cb7a5a7bb381d30875a4b
z86431abbc68bfed1f0b09a604e6a9f9b31b893e9b5d8d218fc8174dc817d2bfa0b8ca62c4bca0d
z4c53738c6888561ef8d2447ca08b1b5bfd2360d6b00f846c384f8df425c2aa237add426ac6dd5a
z2f59eaf19d6f26d937546d605321f65a72f023762c6d2af31f939e1cff78456d15b6831a814c9e
z17ee314e9c75262e8520d88c093957d14361aaab6384b4d15fdab664e560ce43407f784760f3e3
z7ddaf79bb4476c8e433c71986380cb257e75db025f423a7131dab2df909a736b2567d36548d06c
z14acf0db8ed0dac50115bba2f3164c51276acee1611c39881bd7c66d61a25990b20745805cc244
z8ed6e26b90b08ccad6dad0fa6415e6fa29f4a23a2a918c26fac058b395ac0257078d9ad33f37d5
zf21f1e6951f9a401c7edda9e3e57b2d356df5c064ea6c150499fa6833236c8aaec08a6d857d64d
z07b969d31a81c7145e8585d589ca779b798d34ceda75e82cbd718bc6037aed7faf731536932dec
zbcbf352fa04b1c87a21694d29436f2da58c948534fc4cdb2f144cb8fb7e3a7c126de45fd41c4ae
z4e00dbefea67b6eae1d3f6d7c689eadabc0de1df8b7cf3b0a436e52851263162ffa34187f713b6
z2b6f1078d3fc4b281302eead0aa1be1a23ec728c95bcec2b6afcd2d0997cfdfe44bed255606780
ze334f90f207f559e1edc4150b571b94a8b85fc8a2e40328cd5cd68f648b1287fd5af5296a32ea8
zeba83793b41994cf0919ccf8d2d5c1de7f5233433f48e49c1a9c0159994e73d8a469f5cf951ba1
z9d4750c47e435d1784a622cb62e043866ecca0e7ca2637ff7c713f18f9162c77f34fc0663bf715
za28afd609c067d87dc24c8040bf6535ffd2313f10b08d3c1800d96e5ee296959c8d6994a3dc462
z877c5d6ccb069475b14717321518d91c2d78dc1e0eac0f56ae53bf31a82f29483cf7c287687ebf
zf9a9035d37a7688b58967a0a9ab465132f25e5f2680190ca126cafe4d25033a26f863b4e8930ff
z0e3765eb2c70dd29cb6655086e961b07affd8b9d639d1bae0159c4013831a6b7bb019fee22c76d
zf7c045b21441e4b52f5e07e60859e65710a09fa745540e2500b16def3be7f6c3786774896f3d61
zee6d906d6f048ebe7a6fd3360a726a7011f1b3750ffcdc6c47f14db914c205d514aaa6b519ce8e
zc3ce2b1869cb40e10f26efae1625c5d211798103f47661b50beec56434be9ea7a3ffd23c2779b7
ze3fea5e7b7dbd7b297b9b258299df29d8815f008bd9266588f5ebd9432f7a136c342769d404c03
zdbf8aab3a78c5a8a8d14f392994e0a2b1f5107b92983468b70546ff9d15d19fd8ed2aff375fbe1
z0bcc4a49a4742d574f61a64e030aa276b941be8518c64e75b8522132ec48a039bc44784336f41d
zda0248618742a46c49499fb7f4e4dd4b8f1f368061a4e60e836b942db6cad2d02629f83aac2341
z6b0cd9d241a8bc5e19218d0f62bf71f878b8a7f27890a91a2785ced5f710ba2e8c50dc6e794e1e
z7ee98fb1de1118a8c4441d7ef67b1865b477d0c9ff5362049e2c2b9f65e05ec46716839f42eebb
z2206bfa49ae7f01251f58c1073d1d99750194e6cabbd70a1612158457a78d1a9acbf51fac217ac
z27d378851732b3cb442df444842a17ec547f6f4bbe26d0950ffb0b283160db3214830e90f7bba4
z14c17ca9f49fa7197b539ea24c64c909c0363e461496e51c258615f7b033b01959110ed04e3816
z74f3cf704274ecaea29649621bb72c42e8fc284d6971b6ccefbcd54416552689b8fd9ffa939fd9
z66e38d44694763529c7e5057c5cc090b33567cbb598886e45f3a94e6632851dd61713970377440
zee56cbae73459ce10b804c0f37391547592d0751687820baac7cc343dadf42525b422784f9fb0e
z4b6e8548b4ae1e4ebdd2b75ed3862b502d1a150588fc138df0fe9c0899d3967152f8b917ca5f3b
z110dc4079f6d87d783a81fd94f14884860d727316a32f78a9abf14cd4f38f6104fd247d0c18929
z3bfa6151707dcc31f1af1b43bbc2401ba69e539c0d7ca8ddeda57a7ba40e1d7a9ccac5310ef919
z6348443c1d109e306cd21a518eeda253220e2dfba2a343a6a6f1c1315faafed96dfa5e7bf007fc
z749cfbd95530ac1d4e3ebb4b719050a2a45b5b6941f7d59c797a8da21102f71c94f1845d06f707
zd0f725819bf8a7348f957ca0082f68f15ed10ef1057cc79cd89cefbd75b12bfb07f6abff5ec473
zbc87cf18a8f06fb79a3756f7a6779464ff09956bfcf6dccb3955cd8607f8312789bd20d5d18a36
z92ce3acb175955173628f847176cdeb21ec3a5c33c963b7532bb7eff03926ca605bb5aa60161b0
z770b637318faec80d7b9deeaa8db7cfc922d97ee80ec49c58d2739d8d55113d30e15b84f1f1709
zae6e03786048d5dfedb2d0137f6509f6c56da309d51836ba049eb8eee3de6c96e2e66e9a38164f
z0e41cfc2b9dd313d6ade8b92b7674cfd959b14b934396e6ed83ce6b3fa20213f42e60a58712f12
z2a1bdab059b67ce860a405240b6f2bd2219dce5ecfc9f6462a1b3103e5ef9b62eb00fdc20385ae
z54eaf76e9b8fce08762738b8048ac2c4fc13ed9580d8a47919f6c185f3a3586b73a1b11c8da7bb
z807fa15526388f452503af261668105e899d728203341ae73318ea0c79f560e9c8965761c47f2b
z0107fc13795d1489587c4511a78a1a2c97984acfb6de1bb2a9dc3a3dd246550912aecd47a2288f
z2eebb9f90e181312d37f777a29e3452bdf96e8f1d7ca53e72c14e2e3fd2844c0e599028883a537
za82beafdbf8d96670074e608aeef3cb69922f88a23904690870dd7c5bafa943897b12bfa9c9430
z33d514817cd4defcca34b7f61e2803fdb62d23fd36d578d46f93a9e1b3daf91cd2903c494b397e
z11ecc51e63ac2d464d9be81dc19de1fb70371dc6bc450e35dc7b36420b4feee6c72d2bc0e5e820
zbb2ddd0e05f572214257257e220f07ffb1e401be17828861860867165f877c3ba4d59f7248c915
z881a60a59413b47ef54e6e064689f381728f3801d6a7839fa331c7e62fa00063eb642407ec54d7
z11e6430628e2793ca1cbf9225677d01baea5900838b2762e6fb85baa4d1c3c2f6abb0dc4f1e032
zba7246421136ab965a16f1c3ef56b22162d54c8660d0cceb137cbe6d844acabca77cd7dd07a87c
z67f8fd06183f44cabe0bd0efdc186566c1869df3f45ccfc0d53273e905bac009ce2b7e85815814
z85a9a981a5b944dec18856aed0977227ac392a5779ffc70bf8d3c2db7f6ce55aa572e4e625e5c9
z237b1c896ed593be7eb02aeb3a8146469d18ec81db1c67e425f04bdb05cb7097eb91ff8984a3ea
z9c614331968df34823870267fac4a4c343a6f6ebb5e0a1355c6a7a62ad6fdfd5d0b3fa72680b4d
z34be4d607c604ed820bd339b39c433afe097f9d1cf10439b589275064b2d6cf3890de2ba724e31
zf0064d1cc3360e5ec7ecb069ab0fdd4d0aa7b7b4f1efa3dd803585de728a2e2c310afc7a96bb1a
z42629cced0c056fd9ae10aca7d01d309f225fb0d65a711597b6e5e0fae0c1a5024f5192d19378a
z25fbc69c3524f314cab488189a40c9c09d7f613c23478b5d00f32446f61012edcd444fbb2b1967
z474bc2d180915b8525ba9c2a0243155bc6642bd03ef52440e5ce56fdcb7d36b750e5dd1b9edc94
ze0975c65cf49873fe644b6c76e002f65289f4d18cb5ae112c3f6ef536551f736444af5f3043e3f
z4c61c282e69c5e1575ba51a2f58e86ebd3af3d6151fb319db80d7188128fcabda7fdf10e3957d0
zeb2b542c60f4fc330f89f7532bf2e0b3e656eeb2965e90b8c51904468d7eec9a2535af6c842a05
z53a0f7b2e5b7ce94beb497c6778aa1993e3eb36754de67a4001570f67bc73552a66f10cee5d486
z39d0f19c035831592a27a701d14a52e54f6c0f095c788a5177606d4424ed2b492c7b62d743d876
ze54d3579c3a89fbb36cc596797f5bba81f574eac8f005e87163137a0771454a8533819219e25e8
z32a0404841a59ee32339a9c99bcd99969de2dc2915ee8325e4483289747c7afee1e1160463a604
zffdb362ee238846a688dadb64e89457ba227a627436e9a68522cd8b25fe74676f8e6e6322f4115
zf2441880ca515060bd64d298b41e9e43d56818787d790233a85221a84d9b131535f488a8421d00
zedbaae8d75b6c125e4b0a58843dc897d73de940a1221f53969d5bd532a16137ce2190816468654
z12b06e2d58c4c37bfab3797a758a86805bd01aaf3a48b25290298fb9482fb6befe79a1248323d7
z96a02cf338151ed93c022a753364b55d270c314c4969f3061a393746d3c35e1b52be67ead5de13
z70170c14be5818cb5b7773390f0503882797f1c1f711c44ecebbdcad423c43383dae23d9dc29f0
z739b65b1ac4351213d9312c8c6c60e02c73fbbbb6e481e5a291ae6852efe1a7e3b117f0c7b59f0
za869bd55252284c3e59845e9fdbb004b3f8d859df5b7fcac6dddcdde038e8ead302d9b14c7becc
z222cb151deb8a4acdaefc7d0b94bcc39e8f5b3d3737b5439b09b5edb61b0534660c0b099138782
z9941eb3f86859034f3c9abc2f51fda1951bdb411facb13343e359b6d66518f276c78cf32c50acc
za44ac7a1c6414fcf57a4e3be57eea43ad88dfea838b732e67e3da71c4f63634f7115b6c9d3afdc
z0dbe698b6c535902f005d560c3863e1c5ca6b6655454c010466c81aa0289233ae571b9ec537fd1
z4fe7947eff5556b6d4b7d9fd949bbaa82dffd78e09e794ded5d6dc50c3d2a2befa6c7734adcf69
zd9543e8226bb6b2e7408c8793e54d14b49086bacd0e64816f23cc5bfe6de2d3fcadb390dd2a3da
zdd8d2dcdf88748882bfef84d52b3acf2bf5882f4a43b8ca66de15eeccf54c8d7cda0bea13cda2d
z677fe554e0a37a9f9b89c98400c97ecc55bb7dde886f3d955f2ce6d6292a397c9338f9cdd00c4d
z55447ecb23d745b2c2d75c378a23bb8bda7cb3b20b5052bcbf8d888397f8745b0a90c23d3d561f
z8c941e69fea94c9b904deb6622ac02c3e21bb4e66a1c0056d7e3da5fc1c7c91130e3aa5e3ba934
z1f76fa81d2a73f488aff7bc8092216cb0066d6d3aefd7677ce04bd286bcff25efc2a3573a0627e
z70457c2e8403cfeccbf210b3e43c1db3fac5424ef241eec2a20e82ae5b38baf1d27aa7f99c46cc
z223027fbcaab0b5d4ee57e406c6660907667ff320a5589c22b8b853b56301249e68b5d0d8f42c3
zddb0b756446b8d2ac489ebcc6b391964a12640eb229cc2fbe32751e16e3387c62872db27782f41
zd2378c6688da79989eb0a88f1126cd80c56174e72c8b3c5b462c6c705b4f3b8e01859d41515b1d
zc3fc029a8c6a29dead0889997f8ba15886ce96004333565c1f24075cc3043a42165a50f08a0311
z5ecaa9ac887fc539e9ebb7437078028b75ffed02087a106d5c1a30293cc3038d463a9692c4225e
zbd2de54def8123670c2e8a8523b5f4c607fa06fd8fb1c16a47c73785076c9e3b169364eaa6d727
z222b1428950130e1499f1a9f7fc3bb9230b6791f63c87216bfef845babf2514a11a19b789db07e
z773b2396759e518a0e8dc25d150ca4378f0a1e2d6c84bdf178a2dd08385ec7a514e87aef72c569
z1ff8668c2720407dc20c1f666b28d0c77c30b821e902edd96b16a5dc16ca8b8d98920a9ab80955
z229692fe4a2a04dc7af0d51273ffd7b28015dc306f74e419802f61c221713ff3190002ae349e32
z7d7cd484ae9ce80a9a736b6c9b9897a8889adc7a5d41d1007796ae08a785f35f7aeeae2a79a4f4
z03938ed9c866e4a862bb313b85d6f1fd1af1b46fb26b8da9fa4302166407e782e4c3c51c13a93c
zd6f2def789a1c8711cf405dcf6e63bf8484a8c3ca31459e07283ed8a1b5dd5ee74dc15f4ccf1f6
z37dbcbf345b529e1fdbc154c88ac02d359a5d285913a9710035f3d405674c23d181678eedd8df6
z505c0db44033d2343de18dca6da665b9e95a9c3cd439355d77a3
`end_protected_0in
`else
`ifdef MODEL_TECH
`include "qvl_pci_express_power_management_monitor.mti.svp"
`endif // MODEL_TECH
`endif // encrypted_0in
