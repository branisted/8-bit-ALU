--
--
--
--
--               IEEE Standard VHDL Mathematical Packages
-- 
-- Because of the restrictive copyright that the IEEE has
-- placed on the IEEE Standard VHDL Mathematical Package, Model
-- Technology cannot redistribute the source code to our customers.  All
-- we are allowed is to compile the source code and distribute the
-- compiled form (i.e. library).  Customers can obtain the original
-- source from the IEEE (for a fee) by contacting them via
-- phone:1.800.678.IEEE (4333) in the US and Canada, or 1.908.981.1393
-- outside of the US and Canada or by fax:1.908.981.9667.  Business
-- hours are 8am to 4:30pm (EST).  For more information on this and other
-- standards, visit their web site at http://stdsbbs.ieee.org
-- 
-- This Standard is identified as IEEE Std 1076.2-1996.  The IEEE product
-- number is SH94499.  The ISBN number is 1-55937-894-8.
--
--
-- The technote ieee_math.note located at 
-- <INSTALL_DIR>/docs/technotes gives a brief description
-- of the package contents.
--
--



 
