`ifdef encrypted_0in
`protected_0in
ze74c34e226135848fe16db9ffd31815111b6d7fb642c521a3f628cf6da949865580b22efd062a7
ze90adae0e65e66a2c36a587d0a790699161455169ed55a01f2084f11770a774ec4c588039b380f
z6de9c5084882a40b79a175f5c2114b2b6d78b070cb806e1c0aa9258297f4687ab308bc470f0040
zb0b1de382961eeeaf2e279e1462520fc31c119af8f2b214846f56c2b3cd2eadbe4099496abff18
z15cec83ec4a77b868344aa20ba7360908f5c0de2a79abf8b3534b883bb12180f68b5d4beb444cf
z3fba8f13afb0abfe8fcc4294810f75afe452434d2d0f1166236c82f76edf1e12979f04bc35693e
z32ae028996dd85737a8f5adc1ebb94f39c940246e887647b64782cd7ab429b0544c173176cede7
z01dfb26b1f73408344a52b7e1f117f12bb9c8077b34876c2e6fdc085981637012dc9754765e1a9
zc512ce062e0b8fb16a214591f5c81e1353b900a611fe1f4886b57940b41b7f2ce99a7b84b04b90
z916f717e73bd10589c81e207ed77ec660a8cbed5b487fa50acde1b055c8870bd8676023f21ddcf
z9c98cc47cfa2d654ff1365d1f45035a045a66c5dfa82790502623b57a3af03bf0f0c0d35b51558
zb8b5f2d29acf03737a9ca2a053b7a8f06800d50b465c41b30eb585f62f3d0c2c5a43bc4376e4c6
z638be7715fb7ac3386a16422aa59b4c0dc305ea4619fa0da6ac0d6418f316c5678252c1d7e2229
z372090a108321271a4e499c12683099bc0d9210fabf8461e6804f99d047b99f98fa4d6614e2376
zdeba3dc8f8aa3ac7d1dcd701694b1a9002d0335a65a877bd739e614074974c3d436279f1516ed0
ze7c2acf8eed1245bca364dd49c6ba66e2561136a76d524c71b149d583d3f79e5c6854b3a03cd60
za99c935c2db6790b7350fd87631b265ba435667b36dd15b037f68b3e4314f9d7ca5f65e3b4e16f
z97ee2dc764097a073aa58c9da06628726f2a18342c939069be2deace1aed9bff856334c18dd23e
z615a8f3d72de0523ebd74ebf32cef0b659034eee95b6eb4ce9b1fc05c31ce3c9c8613176a6e212
z5da3af5fa937cff9c101228bc99c33138f0dc56670f077388e10284be56d87945d5453c632b693
z8d6c16ab605a6998c5b5c67fd6a54e7bb01a0ff0a02918cb0fad9d8c6e2afc458b4f7122cbcac4
zf65d94eb45d4ac3e16b2cb7df1485d4ebd15adcc105e787847c3ffdabdb3187606d1f7aa780716
ze7de5707e7497b4792233bc9bb933a59799528f70705f88213ea61ee26b290a4c430ba1e214f9a
z76d3a559a17c20ac155aae93395d7493930a977be1a050c5d3e1bcbe526dddf612a579df65da0c
z529b62370ece045a3d689ae713356154b274f02f668a22d486d784e24f3f31857ba25867a5b307
z90f26bb29e2b321e30f35da67ad0ad4e46eb4b765a829ce5c0d82f629dd944df828fd1f3efda0f
z65faf6ae85a57afecab03ce9588fb345f610abd741aead9701b1e49df9f30c9a9290d0bb61565a
z0dc8e55882551693e20e5360ec1f2d3cbc9959f5d39a51a64f5138ec5da9e6e3fa01c7dbc150f2
z911965a56f367f0ee90c309e5bb83636e8f5a7df25a232fbc4b6abc1523f47073a50319c67299d
z3ec20cf85bceb08146c2b1031b71714505d7bd2386ccf2c6c2df93d291baf613cd3bbc8b7a4bdc
z396e8d71aabc67a54a0897bab906d6825ec3240424af8660cb64b51eca484b6896eed7f4c69405
z328593c24ee390c04dfd0719a22577c4e84f1513e0a0291a0161712502f45423137effbf46d492
z949b83dc1ca2162e26ca0251b2ab80b431e6546132f1d3397827a4bb541d76b74ed4cc94023c76
z371c609d06f5f9ac73d90714f9590a621b4b30654e6ee28b9fab1ab6b2ce44952369dec928dca6
z43d4c431444eea48201a2629462ac033580e122798c2571e818b098cf1ae2630f6eb2c0ff86a51
z3a94bbb984374ea4c470c7f6e0049c49b3ac9b600cd2c24e213a7e345c1089d988a781057b783c
z737595cdd1719c7556b844ef381eae053062db5ce0f6f74e73e1139260d0cf5fee93ce1af2bd58
zd23160a2b2df8c6c9b2b3c56a84e416827ba447b01c31ec954131679c8d94085c3669a501719cb
zf0048950209fc05028ef7d46f2770c3c0a6cb801cd15d8c15f987e836fb4938adf16120ac10f49
z3d5a8f778340c231b047fc85f4763ad464b4516ac2727ce0f0d51d410f570396f14f25f09afdee
z01c8ed4429697a04c67ce7495a5a876ff4327d76a3291ad3a42c3a9f7bc304d7de317f593a77cd
zc4974e2a013e0548f461096c7cfb4a86dc2ff64bc8d39fdd42ff9eecb9d9b71b4a47aaea0f6f52
zb92b0a60b5c680306b867ad2ab3b5e49ddc14edd8335007900f1835f1809e94d7cff76cc5d470f
z3d618e0a254f748a2ffadd05b3e9d950a3cb9c3ab8abedb111426b464f3a34423a74169ca61033
z846c59a1d4a9bd8125dc662d07151cd54a8c5f9dcf334f9e7cf4afa3e25c640ba3028d705e06b7
za12e6458312fe56dc66387476697ce9879bb8b31a7e0444e94289f4a5138ca2820fc5d8f7acc11
zffc51a886585389531c010a1a4cfb8eebc69087a3788c3b615ae210876f87c316b1093e2a6b61c
za71b0135c1fb3b69e196b8fee4cb590db85d6ae979e1c97522d31f303a4577e7781561cdb71145
zedf46f6ade739a5361d0981d41f163510d270a4f04f3f018d46a6060daf77c3677c626acd3a72c
z468ee409a21598226149097adfa9aa666a80bcf4375832aa8f0cc507b633703e808e9f38c18ba6
z0ee0c0da36e0972a6da34b546b100d4c43c8f98715afd91ffeeabbcff828687202a730b2815f8f
z79e9c3cf37b6b4c11e0ee2835185d9270f4395692b73f36e98c6b99a6097b41bcbab62ff038d4d
zccdefd0abed348f243c47ca220fa7d20d4b3459a6ea221e8d8633b665097994cadef7dc75aee5b
zc7d69c7a857869472c51246d73bde168861148683790a778ca3aa1fffc612e9977bd2cd0611536
z18ec84c993603720dd6ef6f2b0c9d0b43e11e79dc0746ead2855262bdbca5412dacf7e49629459
zb999d2d1863b3195c4b29516cfc51b6abda7aa138169e3c2b34cdd926121b39be8dfcbd9eca4b2
zd04ca2c6a4764682a51807932d4d01e90c5661571b018f95a5c1ada3b375b21946196b2505449d
zf17ee52d83b34accce1be472bf4dc2b857a5d1503829b40d02ac8ab04e606ac70096b1426dad69
zef9437ba60947e3cd1d0bfdf1285443d4c8b2da738ef71af6325dce9ddbf783d2d30659c2a3244
zbe8013d9bf64e78af5876d31e63724dbc214dbdf7949643d5af39c3bdc1e772b4e585252381caa
z5cb2c25cba43919b33c7bbde61dd4a9be2982c13797d5de10fd6a25a58ede72bc3c745fa83af97
ze2fab68ccbccc3bc8edd4db39dec7c0acb576de9ce914ef82332cde5ec271faec2a458ece48d3e
z3a14e1fcdfc0c20072cfc3f975da795d4c84dd8a3035075ed55f2f7d7d36e1655207483b2c9726
za3e0a71a877bd46e6585d406ed81f23ad452d639e41c1a99c7e69435aa2bbd9050ca69f27cbbaa
zd6fd9b1c0297c41e1dab231509dd39cc4a659e6a50a361579519ffd7c95b09588218e164ab7cc2
z426a3e579d8288525c7c0716b272129885aa831e1a70942282641382592cf7d76552f6f05c8b9f
zc09b1c886a60fe60887c6cf8ba98c8e7c679e2aeac8cd1a025a737b1209a930f46580116daec6b
z24ac4cad7805e0988252e79b62a25b19b5f549209a6422c1bc4c04090a6842d38dfadba877e26a
z2ec32cda4789710eee0a47d9d380a0488fb44f8c53a671c4ff63479722b785633cca2bbefc4c5c
z7c2eeb040ce25fb4721c99ae705992aadf7897cbc6d3bc3f7d0e9247cc150cd4e2c73818469f7b
zcb1962134bb3b12fc4e521e01acf11a7a8ed341a601535146d785e8fd135fc016f66dd2c1d2060
z7320d8ac99434ec603f4d0bb5d3c6577039aee1ef67d2bf24ec0c16f8f5e2f1fe8a4482b0eba38
z04e3d3f85ec80e4d4e753b1fae7b75101234e4f0665e76cac7cad63d551692d400904c25b0a5d3
z9fdfc555a742935e8a81c23d8a68a0be495cf20014a1cf0760e3a38b8d7f9868e0a405f648bb75
zdd351585c2e06ec1bee00a343bb137064584a4534e96dc2f3dacb7ca53679f0f7b16d6cada9a4a
z8dfc637032dd43be21f1fc8bb0412e76a91d5d99a985f301162dc459c647133fcdbc0ff1921fa8
zf4e04c1d3fa9179c98e2d48555e25636e0f903711a5aa389c3d2c8963033efd9d13f0eb1a3c2cb
zce0c45ab3b9b91f42969579bab9160f65408ddaab021cfab6b8b3b00f24322d9dec5a38646fb54
z312b7b8676d8fe5a7425353d63c44e75a8bc113f7f5a3f91af3240033a428967a9e067de7e7ee7
z04fb3af540aded31bc1a8743b40791186789c815fc906db489e24fcb39469118e661bc219178ea
za18a1747bdee6e4f0aaf08a763ece24d0bc5367fdb37bec50c920def0b40a26ca57b9b84a9b4aa
zd09458adaa78cb561b0c1ece6915096658e5595fdaf31fc941a856f2760fc0d99d9060b8d0bd2f
zd3e068f2aabba2581e165150b21f7641f89b483260f6f4c9276ff30fc6f6348380a393c7a0f4d1
z337234c7057be0811e48feaed7d5284b175927022d5e88e133821fc37a76eee6b0627e39afbd39
zb9b8fa6aeb3050dceb0fb84166d28f012d5dd99a58fe735e741b5ef22fc5b0cf48f61a64fac46b
z6a592a15cfcfa39043bb82d613ab204f49ee41df55bd2a943124bb0867fbfebb9650908500ccf7
zc4cbb3688adfa819aefa58935c919eb8aae54f0c63a072a87d0737b6d60d639111413cc24bc5e1
z40e8884bfabee380cd3201a27efb2f7d1ab3d1881204562efa3698e91bc4e1390801255f524559
zdb4c2c9c4c9b6b683f201ebef4cf7e723c859eb12eb43cd67bd7f3a6f36a9c429eac32b63289ff
z596e7fd185d8583e5a484aba2136a7d3e019d948d73012bccd9d0c802a8db876c20bb098af04f8
zc587016c0df3d569bd10ff398b7c1003d6c60cd48295613a7c89e83e211aa6dbbc65ae9a8fc0f5
z359f1a08e9ed4db3810a31b52cf6c6ae2c9b03c472075d899c250c6f61b412a8803388717472e8
z54ad41f081785c794e17c090b528183cb3643c116f0c79a0a019948df062098b77b20cb499ccae
z22dd422b83f2c5adaaf72f172de2fbe39eee9d574125b7b85d1b81016d8f2212176750fe8b0f25
z636bacd34faacf6dee51bc2aaf893fd4c51c32912aa5b9b54106ab1a1040c3228ca217d8c2a654
z654a1c3ce3570ae446e9ab0eec73d708b45c13f0585c4f84b8149d9f1d6dade79d5cc7eb1887a1
z59c386c67b91c6cd45c5a0e6505f6cd8b6341842527b3193e4820696e00f2dc98a98a572d937ff
zdb7a106e3155df4925924ea1a5cb893c05d4fc71859c17a2af3540f6b0ddd94aa9be20ae1644a0
z968ff8bf9dd495cd421c78e27cb00ad136abd79d7e9cbdeff413c6c66bd1c3566d9863362345eb
z02e7254c592c02b06e9ae20469c46c9246b5e1e17135a4130f7d6772455cca50141f7cb4d58fa3
z5d62d30cc0026dce306c1cd812df37287a5b85e776add600ae63dc157070e9e96416e79e676850
zf9887e5155b1b780d8a3ee0cf67f5c773157f0c6bc7408549531eb051cf6843fa8fe58bf16bc72
zba2ee42bee5af9aa73c271ef8d3cdfbd8dd65faa03f882eb8cb411969913c67c602d8da4dda2cc
z2a8d39019e977683b3ccab6efaa82f1a5116e54314ff14516305128a6ea04b445bbb01ecb9b1f6
za1cab812dc6044d1a47b4c42721936ed68c3cdbb5ed11bd2bb6487d490dbcc2033a2dc0e20dc5a
z823c75fe516ea217f17989ce3627be061f81cd4754da838d3a94a7a60a22a06ee0e181616074fe
z16a5f27bcea1fc6b26bd1196e75008d28a03f3fa2edc574449e64354dcd7ce3e925093d0ce0f36
z13f0b310d53ff5684d39f9bc1cd282dc27419f7e5c1000ae0e56ac6f64d3f0e7712b9a8e6bcaf8
zf0e447650e49a8d5b98a0e6c28e62870093251617b2031eab91338032dc3199ca065e3a2e04153
z56db107a4d8c8d21765780283f85a4aa1e456ebe6cc72bede82aa26aded9ab35e4288d577be8cf
ze2c2f2f3190495e35283f830730be565c0fbea325618a1ccd6bbe6d8a920875c59bd66bf085f03
zebb2412cf62ade568d5938bca7843a940413f930b6d379aa2975e7d0360d13332f2355dadf717b
zb8a7385f7463316cf86612205a2d1e141f0693e03c13da9a2feba3aa31dc0ffe4c2bfe86bf4157
z16dc5ca8657770647cd98af48dc07882dbec96ed232573844efa55b5822636fa42e414017746e8
zc3a9a70badd8f957b21277038dd7866c6d91e886fb69b6b7438dcb91182b80e8d5533e770709ea
z3f213832457f73a859e3ee916b24129a1a8ed1aa9f84c4c5ba45d6b4f9bcda24849a46618e40be
z48c307859cfa5be6a4b3457a950bffac6f4e85ad2933901c640554fe8bfeec66b952bef71c1576
z11c085750c66d8e1d89adc907cbe2fa71aae62d56abf6754d30c01800eebd94bb8f2fb53a59e34
zb61f9747f91a4c7a1828e34db7c3c8e45ebea89904840f3ffbe00c193aa40700562a1f6610e191
z106a7955fa1f0c72733ac9d7a7006e2776f4a2eb5f01b6c22390dc070acaef4b4d239a60894ed4
zdfe68b2ee2008e192af6e93e3dc364440a593b19c197757a6528a68bad5560b4afd539822cb600
z87bbdf9eaf1d8e59a3a868f6de6b502a7754b3705825077f8d0db935ec1dfb903dd8399a1ce392
z4948dd76872c5fb6d225edbbb9b03624222f82d1cb0de2de46fd1dbec206502baa370607e70769
zf23411850ff4f7ec746c9f2e78338b2e2b38427b8272cbae15571bad909c54aec0ade61c069b9c
z0bc65c45d471ff9c29b5b3288cf0ebfd501a373b42ee52b063bfcc56436022f4d8b746794a8188
z276dddc7091bd9c0daab5e7e9284eb8da5e32c0afcf30ebb99de5029aae368cea78b7d8c749737
z27c9ef412eb47739a29dd9b1ae5c7ebba2218fe233f4b14ef3ca942fc4d66483f200f4a26b7867
z74770eb73ba3f5eeae0445f6a157c9defe073af4c8dd8eee0bcdfad3bed6f5ec0910e36ac4ee51
z936fe6aaa5e6cc78dc5989dfdb80f1130c021df05003ebc5282f12244ad343d416662e4595fd8c
z5771c34f6aa17a8078387bb42f231fc755dcb3245cd004e01f8e9dfa0b23086c70be7cfe84a52b
z8354967a2be8b1705de62489c3d2b7fc8c9105e53f10629d4f6cfdbd44b3331e49ee47da5866ae
z871284188eb209170937fbe4589c80858298d755accb2af1d02f043af0816814b48164a63e19e5
zd89623fa2f489cade65de2ec63fa4df276f99af0581d09c2090aaaee9d5284c71476e7450701e8
z11afecfc6227952fa03576c32a2090a087b47dba79a8eff2e56d617e222222662d49a173ab85cf
z6506d2bbd6d525997250aaa54d4dbe94995809018dd11467279c53f18457cbd9151dd59462eadc
za414112b5727b683cee9bb4a797a0bac7824033d78bd0a9d281f15f56289bbbe64951f3f5c7515
z9d8ff9734abc1d0346804c22681e48e9873f50cd7318d5d35970a10b7c8f7e355a6c7bbad8e8f7
z87af2335c486aea5803b586197619e68a2621a844f9a554d5c69eb63dc4892b8579d1adeaaf7b5
z1096c76365cd015bdfbb329536d4b39d24f328699c4734e036096454d5285d2694d5e8089f2553
ze87ec4ffa0bd0f87fbcc3219b764268c118b22d7bc73e051c03c4f9bbbf5d2b7afe04ac0641b7b
z862932dc6ca8a75c246926fd197437cc1908429c91c4c27c8c0f8141169def8e3000112700619e
zd5f0a5933c9ca308482bc65f8c8e5a5d4c25623162bc8d68286bcb1da6db129a1b9858a3ff4b43
zb4b4404c09e0726b55d6ecc4f53327ee2aa270901313467e60fc9f61bed9ff7f2b4cde3be78a34
z76b7cd601e20af3960a630691b5332b517ae147dc4d3d5fdb19a6f8ccf878422311418e4ece6c4
zfa82dd2a26a3224c6a535f60ed34d1bfa727e7fbb27e707542bc13a1bfc371039a6a6480fcf87e
zef14da208f556fc43ae41b11f2e9b825cd774e407d1dab05479591735c9b96fde9cabc6664a8bf
z4891cc8d93b9b663e61de2cddd3beec0d2081acd4d51598357ec1a08a07d6e2d6aaaf52e7fada5
z190d14324897588b4837b42697efa3f77b61036dae03279f695f8ae351d94fc3cc0fe586b10680
z8f0743f6a705b87fd451ed795b28a6c383e3a5e10b46970a85d6631d4ffed1feeeba2632a10fb3
z8ee90744f35039e7f1e4f722cf7ab038bdb6a045c1e5f20b2152cbf985d2a5f8939bdcf19f22ae
z95924ecba7f5e7305f8cb435b7f36990615189d423470cc2196073f35d5c3e3a853da75936efb7
zc6ee92916a246d233d0c9870c7b0aa524487255d341d75948239854db0047556dda3d6b7647481
zaae65e97e287c52f7d7b014b4d330e73ec62b31fbadc9513274f946966391e51bac02ba2b47637
zffa8a2e61f570ff3cb516740bf363e9f775449f0677787a76b1e9a6b3a9c113637f433e0e7b8ac
zaefcbf7c4269047702f34958a81657ae6ca1b88d7826203f8e25a33f44935120248a894860a6a7
z04d1d085b083d79969a1d32a70ebba67ad23a952fe7bb76f54d60bb1134bc54128acb5e3a86ce2
za9aa17380f9fc45ea63eead65f214876fdb2a6e700b6f85d40e3874f72a230e51f26933e
`end_protected_0in
`else
`ifdef MODEL_TECH
`include "qvl_same_word_assertions.mti.svp"
`endif // MODEL_TECH
`endif // encrypted_0in
