module subtractor_8bit (...);
// TODO: Implement 8-bit subtractor
endmodule