`ifdef encrypted_0in
`protected_0in
ze74c34e226135848fe16db9ffd31815111b6d7fb642c521a3f628cf6da949865580b22efd062a7
ze90adae0e65e66a2c36a587d0a790699161455169ed55a01f2084f11770a774ec4c588039b380f
z6de9c5084882a40b79a175f5c2114b2b6d78b070cb806e1c0aa9258297f4687ab30857016fc53a
za25afc8341302f0c829d94450c399b8ff9b0386c187cb854ee330605b7b59da379b1f26f488e1d
z36e675f0b1336408b3a1ad87d0723054f952fbefc8d5a33eaca6ef5be8f42bc59870a29a5cc9dd
z4fec09ce6e44cac279651402e7e1f590df88ce49ec26ab39f12b4a02855703c6f03b1e85c797d7
za357087d98e5b1f45502e45892e5823d6fa4b762932009620038c05d74efcea7c3fdb38901d620
z36515d0824367e48d1bc182335f158c262d396cada6b0ad58add4f945eee634c2dceadbfb5118e
z14969c29a743830a07124bfa78707f3952b96b0db7af7c9ff36f77137d8c490c4f79328328069e
zd7d5280e4f95742c9841340368b9764f0f80413adb175ecfbdf3c40716abca7b8cef6f7fe92ab9
z6bd2453f1aef7f7899c5365c5c83793cacc7795c269413f6cf0dabad14d40e9285afde8c01a47e
zb61893788ec5060288cabde8fb553f21b02eac61ab0b48ad3d54f4d1d76508b22f0c600861b5ce
zcb30ba708be817b1f50f59c0f6fce449203e7355c1be55b662fef3f92ba58243d81537761af8d6
ze27d7864d2dae99372b2b75bacdc0437a4f7e011d68c3487a89759e3625548fcc920ad06471ee7
z2d701aabf726859343208b0a543c73eeff8406febf277e3babff437ec820fb49d6b78e73bc2353
z884917487d35a6cd06d7d73ccff5f05355122888b886d178a03d8eac5505df521c14d1e332b234
z86bc1de9891c0fe4654d9d65be6ba17e0f35eaa0e5fb8d4ffce747c7530d86192c5a60f63648d8
zec2b11ca4783a37281db3c8b2556885556aafa013f24449e0a06d5242cb51399b3e756b814a7f7
z7d2f3363d024adf895ee1f4c57fb3048cf14f737f4f7878d0d0c6b48a3aeecf0d16f61ec999e70
z8673047544b470019ece6d4e6f8a1469b42dc3022d4e7bf3ec62c2af4cfb08f5a5de608628cf8d
zd4665dcc3f4867d0a07a836531edfba94cdad9d90730ba8b6b2364b0eba1514c0246e78124c617
zf6a26bec02cd6601f40650424a431a340361b2120bfaaaee24cdba68de41a962bafca77ee84e80
za2da1ab25b494bec121443cfa771b7300360491417b42658f3967a20c16d3ac0978600bf5db91e
ze42f8327318524a1e54cc36e7ad8520c8c816f80b84c9f01401149c4b5521b29874dcedcb6a724
z7fd67ae188c4951205e57e15a4bb9686f58a9b570746ebd56d92eeab7dd963999e8dc513e3a4cc
zbe9ed70662685b28ae56c319904211dd9c244d5287bc8c3305cd1a4c2c431d457192b7d7c21d14
z0245708796b21783da99ba1bbe5ec4aed7091a37b97cc101d6723f1ef551bfd041935efed04827
z4274d10879f1a7055719c83d6b8090d744e208e89d679aefef608437d34dd226c1a50945d034ac
zccb76221fddf1fc6ea9de6a99bdd4a14a48506d1af0040a2305db037783d0d8af7fd94ef7e0c5b
zd810d5a686359cbc5a81df8a13a8bc68e95e0006b8a92177843b61dcdfadc53b4aac4005fcdb1e
z5867862308857eec76ba1be7de9ebed0182158fb0fdb5c49f2f87746008edb0ab936d587d3a303
ze07c3d65c1c6601f9c9d6224f36d7e556ead929e45462dc47b08e3cc7dc32fdfbe6f97e0043e08
z3a13cb7a7d843d9a0716f96e44fb89fc4afdebf8f85fba32e31a1623282bebce5770f3291121fd
zfc695d865e90e0f245b92f566498c13f53a270f099b629c3ac709385fb9ff940ce86245794324a
z63eebde0e00f471b533d5f5590889893a26e7cd4bb9093a6e9d93cc141b6e839c9c63c471c58dd
z2ce92c0a29d5df5231f0e77a2d14661623d1180a93346f19ebb273a36638667bbe5d4f3a8fa4d5
z7ea67cc2ca9d8cdc4e3d778c188726b97fbdfcf505378eebbce0fc81da205513daca5c1cd0603c
z1cf67b7fba7eff139c6bbe8ed5435c56ab0466e6d02431eefe0500bb6e2b7e9b1f4cf81fe2fd28
z5cf06bbc02df22e5f7817df7977966fd1631e52687fdb10726aecb458dd81aca4ed71fc2c38074
z93e12058b5f947899300e3f99a057bc37f8ef8ff7d710bd0570818e1fd47e091be7a3aee3b8283
z20d3d0ff2f53f85fd2e6c394d07edc2969dc2df20387cc85b9fdd926938d532a424e90c47e7f4a
za2f508afaef357b334eac7b1a96a71adc41b7b2fd868d61bd2c0c4fe817fac7e49e63c7746a8c4
zb55bf7ea95760171b441914035de0da0bd1535d738d6b035fc29ef390b8890e12d0ea422279df0
zdb1e1c9c83391fd2df385d9797fabe8ad5f9e02b6d9c3710cc41b5a737c69cede823cc7b304f75
zc33d09fc8dced2aa080672bffa7f95f55e4412f34dae1bef8d824b30c7d32a1aeb59c84c369333
z1f7093abf04cef178e51ccfa1c06d6a48dd8277b41cfa77f4133458c77408fd7ca679d409de218
z6b133b407c6d0fdb10849e8c75a1471ac2ff3a8191e61b528cf1ec1b48a3a575565e9c1fce2094
z8d0e90014f2bb7d9574d3c3ceba44876918c746736faeb2d732bf538c010ac6bb0a234d36c4283
zd043f341b26fbe3f32067d2dc037ba9904091c8479b96bbf97f8b971d5c244c34542a44cc7f1c7
zfa26b3c9ad1757c73f726734282873f6e14a73b85217cd9b797229e0d1c9f95359506dfd89574c
z853a92199b3e97f92424aabf222d2ef4b241759cfc12304c8d0e558ceb80b844f4099db0c773c1
z06666e452a40d625812c10caf09940593e31b47ce8631851244b3e9b85d3f76a7228e9f6ae5f4d
zdcd3fea2c49eeed237501ddad5938585adec8b73cf28583ee5b521ced59214f74e47e843a1328a
zb00ce6462739777d8179f36ec66b2ddf6cbf0b8130686a3f318400296279e6baa317968edd6499
z0b350988b6ff5a26394d6dd5acca2edaf453fc2f238dfdbaded4e265280307704b6a9cdd05d365
z040f58e9752312bada6e7e36613ceeb7f747340224e4ea306597f27408f0de3735ad5b079ca740
zcb0b9c026dbca8b1db7951fbc0070918526c17e5377b2cd13d1d696945e25840c296d8b05e4348
z80f465b0897768c94dbfc28c6113a63a6b8fb2b1c2b48275170761874a5f00ce81b720c77fe188
z6ee8fafc20bb3a47791d76f8d7a22f720df1c4a0a13dc8d98e0eef025fb1dd1834cdc923b85421
zd08881cd93fef5084580d422827c3b5888598ba13a8d6fd1b72030e0a07480089fba9ac1dad4f6
z865fc5bfd6fc9e75c92aaac47985deffac790eaf84825f4c026287164d16d925f016c45b6b03dd
z96e33f25fb4b7eacad91f388a81f248f9bf561e280276d3cb55a8f9c8cf128187ad7a5f3de44c4
zbe052baf1df16f845a1f5fb72f2d1068e571dc86e8152939b0c1dabd0cbdc18873e9748fc8998c
z4e96c307e4491337c5d64f9a6bb0a1dd99e577a31f0a3e6e17d5722c65a426a3c5aee367028bca
z0e2d4172ebda4e82eb85cca72f4457d26e80f62f7b1c9483208d3cf340de102ece6bb02780a0a3
z47dfe9c1206c9cb737de57da66456197bbfbcb6983c0db890533c303479ca424533da93b3b3f37
zd318c6e928ed0e0f364b316682ae6b29872569c175721ad25a743d42e41e5c367208d8d078887f
z131207cfe103548f7847762d5f038f7ee3b8a0b7be0419abc7dc93f94c2168659da5d1482b865a
zd63b88d987e120455bb2e7286dd1353488d03a7dccc0454d7977559629839c598e399d02f41b17
z47dc35cf9c94343a8c2fde4d37bdd4dbe13f5c17b9fa746a86d832ed13045a13c76debefa6c69c
z129e90c8434fc1215bbc18b8c465ce709c4a592c8216387a35c341e0f7ae16584a95b314f4b497
z8609b4ded4eab0f36b99919c95e6a8c5048436994381e8637317f0c4adce83a08b52a822f72988
z826f320447e4d110fa5967de14551ec272bf2ff066e69e769f1cf7fd9733767c1eee2f09eef2f9
z9ea652c950d15bc9224c02689355fdb3bdf1d4e60ba64dc74fe1ff59736fd8fc4e772d4bf0bad3
z7c3894f8e1371569f537087fcadd0d43a96a97ec36f31bfb8eaf15d326c3679c3246f6a605ddf7
z20c8507081364decf503c2168455a406271f5533d46c69f6c0200c8df6a81aee0020e015be2114
zf56ca3ed113214a01597ccc7b81a7d07a663ee102ba93f6e0044fd1a4d1805db539d4ff47bb16b
z4094db4a7f088544390623a8ad29f999c515d08b52f8a185ad452ed9318acea5810a7620986689
z6ab59fec013b67078d6b609c6ccb3060b809db40ad3b996953eedeaec19c00a112aac5ffdb89cd
z71df5195f2ca76dbd72ab7d59c07e37354127778a3ecfd8c79b1c43134b677761967594815932f
zaa064adc510005051d440b949a0a317ae9f5ad341c3694144246c58cc1c0f2a120237abe734647
z9be2fd56be3de8e3ba862b35d988e25ed2e6f4317843b67b9e9cc01c618d95e4272e584a15e1c3
z9fd112dd6077dbe01ecb8a0b4fcf2c2cabdff71fe45ef0e205f46e62d35dde716452c2654ce2c9
z05d33d9bf10e94979fbc8c24faff387a9c4c4552f7308d95c69fde0d3fc525230339f70743be8e
z4d4edd5ddd540d51a302b6abbc23a994e08f8f2edc6a1c38f9fea788e14fc54be165989a89126e
zf54ee4e4c5e183a760408804b76ffd8c84ef6feaf7c815ffd619bd4ec91d3024aa93e32569e037
z9dd9ba8c823ff0d16e34ad1cb326cb7170168eedd83ae3d4317f336aa7483ce0750a87ae5cdd33
z91c58382ecb620ffb48c30045e574f9b0617f715aca7bf3d7d95368d511f0af22e8d65ddfcbdeb
z0390b999c3b85e62bfff06a07622d18ef4848a076307eeb9b6c3799de0fb69fd35f63612302e9f
z9ad211947ecef7f17f1e1842e286d46d2b96b39d003cd850ef1857fc06eb901d86bc919afa4615
z7da610345f0e0d5d050bac29539e39f42afb52e6801e9cb240ea6bfc3037fbc439825443027459
z6cd8dc7d24271385b8b5db1971b7d71dec8f823f10ae90d31b9290e9d616947994373f22df1ed5
z3f72cd6f262addc42d1ba52a5454ccc612cc382651e5840d16da5fb4a5859279bd4731214c609a
z56edfb9279df57f06cc2a6f5f14eef3e29f278109164dc96ae2f51edd05d30f20d8513ea4c46c2
z15c8df23c10e7f29d0eb78b3980a621519223e9dcb9f1b561ba5c45f350323a236ae2752e1bc1e
z9264a1819c57e8dd52fcaa51c46b7c622d3b3123ad27444a40e268ea2b808532cafe476b2204ad
ze608908fd6d0a328df67ea2c1a2f942b53fdf34cad81518c65c73e10f29e995d3a83c46e46f807
z103d2b9cdeeaa0e27b97f0d6b7f76624cf5f1683f5932fefddced6b3ff01289df5732ed55d00cb
zc984f9a64a2cb28ff931689882873341293d96cbc02a9a8b69f7fcfd8f97aa5b9bba66970abb3f
z053dd653a6f07fb5b887099acacb8512ff101a733d781d5bf18784204a756f64be3d8f14cec57f
z30e6d4600274f911f7bc0d19c95799ec03fd15883f6e8ac41ae77ba9491c294d09da443a89d1a2
z991b82313478732f873638436f1ce51aa8165a3398af35dd843fc31131b1881edfe92ed764fb8d
z533bb05aa4bc02c1d9007af69ba5ebe1bd9922856e312a2c0d3ff79a56ad047ed4a448003bd433
z355d5ec3ee02d9e9774e422101495ff8ebac4a3e07a25076de00fd5bec98169453ffe1edd2a55e
z4c184b5f4bfcb876488cf02271c908d44ca3ac7c9d61b713303e8c42b387295b0020000147329c
zaa978eb4db82c05b558d38439b0ea2581a2b34c2270f7975eb56c38c60cdbaca423eb76a6428b6
zb9ffe6ce3ac6ac0151da9780f8731915e1cf062bfd4a3adf06bcae0d1ced1e61026dac4babe4d9
z2b042c6148195b048d232e02d75fc38be4ffe62a13314c7cc500877d1056f30eba2d7a06190c8d
z158d41a08dcb22e0086b6c83e375e279b20ae151686f8505a5b369b43a498da4c5547f70ab684f
z9571bfd1a4dc79004c88b18e3635ff014e7a5170b3c6e63c9a62101190f1462ee868e38c9ab22f
zf07909f91cf62988cea7e4b9de06de47cf1205cd68fccf289685e3f15a03b46513264e90a86ec4
za6219024474b05ad504ae78453602ea4f5e9e0cb78b635aacd706a605d67a703ff85de0e3ded8e
z62d9ed70d8e541025632ac0013f261a094af2b28479a09f88a11e67257afc7fe1b55fba47383b9
zd1ebff27b33d9910dfbba821d719f01b5e17685410e86ad2a9ebe49c824a656ac90dbcdc789ec6
zf3f331d2c55e57064b929013b777b0c663d0fcbef99077b699b3fe9cdaad607001b2b785a52c2b
z98e8c27b0724a45e6defdfd5e236068613bab974d680be5c3f5bf42f1f4606a84c20055d5c5060
zaf3d51565141f04b952646a51823ec5365ea34900511e8e80f092c74f856e35c47b5837d0c9d30
z6d7999104c6c28936591d89e8583f7f29a7d156c906995ea704167e15cdfde82cb17359c9dda0e
z5f44c2c049ee4ac875b6ff6ea95aecf5efaa04cecb942ab71498b5f7fac46b7825d2ff8f1b1ec7
z6a291fd756aa18f55a69245845b3320c96fc2579288d61ae79da57fa93a56a805cc48caeb2b366
z7107b256c68fa5df1227599e35d91b73a41e979a25384e74a54a681f7e33b3caef488723df0bf3
z699bb0259ae03bece06c15706b5ee51605e8571ac8e9767aa1780e46742f906069a0edce18e621
z7bf0554fb83b3031f5ca11a1dd1cf9b84ba6350bbcc8936b9a2161e146b82f536acdba32e8f9da
zc75e758f4deb777e5915b5ea7e21a05a7cf0d0786dd25acc0682e59c9e7deb1f20e3815c745856
z3fed503d0ef2f2a09cecefb27568622bd1b0e4ff1ac75f08be09110de7acb44d6ee73cc07fc9e5
z0b8420ddb81b5b77ae531ff489f6917de00ca6933bca21ec9015dcc9d9c53ae995ddbd68ea00c6
z77390ed7cfe8cc2bcddd6fab3446eec96a429024126f07d069809ea29b00ec0403525619b737ad
z62c2a1a785eadc9df4784817fe5a870b83c5bddbe7d38635afe6833f44240eb8e2ecb24aa81326
zb2692debc3495f7053d746f58a27c0f73e17b524530c0545be2dcd18fae3df19207da79b0eb22c
z73a1ab76396018c6c0c8113e6b794ad0921e80523da1b6a77bcda650effa45aedab23936ed28b5
zef7dcad4bd0b2a8d55759483c28668c24ae9487b52cc14221d7d58c97a6129d6aabd0b21704f07
za6d1210a70a64268564157a0644ecae52be7652590475cb4e6a475973a5326b285d328e33ddae7
ze7b90189a60f12f250f329aabd09ca3b5caf4ed7873d2b1a10adc1804fe1f5864caed40697d15f
zbe96ff2d42f183f1e10489a9ae62eda7156b5188895c724c4eab66cf2747cc3d1e12a2a2f3742c
z6090a173a24b8924f15abf197183744fee7b30d2008a2f2730e1efd631056daa818565369d49b6
ze907334b07e32f88350b6498b7cd09ebcbe7832e24af39b8307b68dcadec2dd152e78dac585be2
zb9df8826313ff201de402857b8f3566e89943255a7a87f23e07b74a4b46bf76009d17fa19acb63
z922281356dbf5c5c72ad56a490103b3b87594a8952923011d73e721ad4ce9f8782b8a4f7384409
z0c1e9742e6d45d16a105162422b815321677120f3414395923515ae10076575a49505e70bb3fae
z907cdbf150378aa90c4b61525d8d55f24a6f11c84bd8cc2f1958042e4786ddbc0585c0fdf1f274
z2dc2b2ed4f0fd66d68b6ec5148231f6c202600e943336a61ab64ef2db341051dec6af4a7de6a5e
z1c502713e92959fa10a67da7e1446a298b07f8b195ddce0ddeabdce7482b8c8bb3b15681c69197
z7e7d463eeba6a5236885e9e7ccbdfb5449578f767bd8de35f2d3b2f87bfd1d365f8ea82095ad34
zd17f87ba87b24330b634a86ad6d14d923ea5c3b1fd82e0b11d4a1ee00642b9fc68f66cd3c38b38
za27fa72b7aea7a4f6f1629f8ae1b495c54f5e59da959181060682715bdf0aed47cb498a1c25e10
z7fa0f8188b7511b851c9c1b2a54cbd8c7a39d6711d20f1db271a280255206743f669a8786556e4
zd12241543a6ba75e99d517c7016c5a874b7d5bcb362b0832b975240d23fadb3b6629f17965fa0a
za78982e0d7441e0e31f0969c7ff8933381fb40a334ad108ee8e888d1986bca485eec4ae5e4558f
z7838fa1705519994d6359d42be2ba7ac15edfe4a253986d7f806f1a2e4431d1d339ab8a22db721
zb4a1697b606b3f2b11e70ab6050e9eb12e5f8dde8d154664d6d63f1e891bb9473c3d849c98a084
zd532a570bee89e8abec1e6add916777de9408313b541d62f590606d7029d22b4f9108c0cb8fdb2
z6d8888941dcbeed0ceb096d5dc7f4be18e339ad7db3687d5419d76e7a14be516350872d749deeb
z63fd6b5497eb0193cbbc2dc2941c4ce99bc35bf86c6c2532c3e1abc76b3e8d4df543dbbe730124
z10e4b036e10f3cba092e1ba275a578cb0c4e644bc96a73d5093b97a8095cdaa80b8001e6033574
z2e52ef4911ee272adf276e3155444ac4e30bf029d9518a41118c85c6a00d6bcfda0e283b8fc5c9
z8f2d7224930e33dd9ebf4eed1d613e7df9e54914a5b859887778391954c9bce6f67b273edcd992
z4f16f80d2d03d7a770999f7babe5e68debad3b69ad317925a505ff407e30f860fafb8ea7f02245
zbb4b65da7ae816562cc08123ef543843a2bfa9efb094d0a85e2d12df0eba955f17cea03de6d025
zf177cf04fbc1fcfcd0d31d0e4aaf4833a9c6e7509b37a867fd6dfdf573e781adf4996ec63fb57f
zb811c9aa60cb7acb2a5a55486caca924c4619172eaf16c341b274d519b8328447c2714bf0cd3bb
z10e9745c9d7a90d9af4a3a972160d26621dd4f8f688867cb6e44bde5a919c5d03a5b061a6ad97e
zcd144d4d93c11019c697be967c7bf653f7f06fab60fbfc37040dc23f045a3ad0ff36b81f93f777
z6528f8dc6e21c25e501d2f635b54eecc33eefc5c29503b5d02a2e89bf299f104278a303e8ff33e
zd9bf46e39b361560200fc2cdc2a5f70c2417496140389da3c58990c7c05fbaf91ace35ad1e4c05
z1ad7d34c4cee48e1ec457ddc6bcc3ef47dea8356ffcebf6ac3aa397db5485e9974c77b10df15be
zc3302360086ff797f1010b3bf0b6fbaa7775021338e6c184cf29b629e1afe4973ebef67af119dd
z766b6f43b2780657050da33d56eb34f47e09f1798ba5e55d526c217c041c89e2c5a92c627f7f7a
z5f880e78d0f5aec755cb5c726001b9eb0767bc5ef527ddb764c1f23a68a75109f0fba6c5186056
z3ec7db2bb456dac5ef5fc9a21502126389cd79b3065b6c9eb1a5aab8cd104fa6a4f22b19599240
z8a84d04bf003423dbe7d87460e3ffce60c273d1ab98e0f63026b70ce4695d4829c9c0c24eadf32
zc44b7779ea845a8592e2a439a23335795f827ec4e5ddd6f1dcbdabe1e418d3717318608027dae6
zf11ed0dc88689eea194fbc1a69c5d6fc4ff0d5b79b4d55cf30a232d0bdcaa2e4e329f6b5929ebb
z5d4cacc94b40771a26a1bddc01658ba950c82a8fd0367312247504efd7e623ec3112b50271ab2e
ze79b8b0fc68288dd0f9e2e326c5a25b5178c84fb0e7163242b6df9b6f3e7128d1e69626ad896dc
z64a2151485d208bb03bbdd2893dcb0818cadd801449e1454971f3ded768dfcac3d278a9121feb8
zfb06c7fbda75c7e6d3bb550528aacb54ce6d14130a01034af9937f90676896a379a46959e36a16
z2807df2d6bc5badeadc9846a987fb2e54b2148a7daab471d2d47803bae01d89676a2f430218313
zeb266e43932d3eb149040f64012ea59b848f7b6a0ae7689ce1c7c824f90d371d65fb8671f3bcb7
z233eda163636ab575a6fd1eadb5b39ea57f39d8e5ba77f29a6534f67f4fb1f554b741614dd5040
za7595f99fb08706246a11438a0eeaa460727d347f794c6a898817713cb613c2700dfe6c6d00fcf
ze0e17cdd104125c44d7771be3c0ed1718a0b9f97352f3db0fa1afc58fd89a20e6ff17c63ebe479
z173cf904ec363eaa391dff161a79fb24343b9e3e0de19c7d26f61c3c4b6e7405537a76bf998e16
z2d0988dbcbcd48a4103f80aafb511bd0036cc340e1204d775896ea3751bd759eab9e2522ff4261
z5449079d5ab9dc951452cc571d16b4446d940b58e1fde07db9ba6f124f4ea4e79252f38a4b0561
z51a5add41497205753ca73d293286d5e92ed2d6f583946d60b16fc477c519eebed1b233b049b32
zd7d50d4339672ab8bea77138d06fc9bd9d0eedd2d91a0d32a55bc60aff5ffee7efcfaec4667115
z45f2a1afa95f33234e5aea5ed58e49a44d53ac292a264cbb1249f78c592cb50fb3a9129c215f3a
za0bdc6565cc83a51be8e880433dd86742755fea1820074fa1bcaceb38755231bf32734de346e99
z6020c50a7022b8b054fd10e5a67e201846dfac24f5db7b608c46dba77b2e7063b04bd1d22bc5d2
z7da9aade05cb654e7e61a0599d44ec29cce147024e15e06c4e40ef89ba32f453ba7f55e033588c
ze540e9e1d607bd4e401f16c662c7bf117c8477117901efc95e18b7d757a99df4ba0a200ec4601a
z52ecd1abea97c7ceff8bd10f186c52d6ef7e9d73d59d09b91b0940613b431bdf9324caae512f09
z7bfa10606daa4e3d195c40b6702ed1bbf790ec11a04b2de06f8a55f8b48e99748b634bf2376d07
z8c7ab08a1f18b27d2621ea582b7b8f3e1087d4bdd3dbd91b478ae0ea7180f5b9f559d98c1fcc20
za1bb3300062cd07dd272368cffd9e1dae5f1e46bcc4820b098d2b6e1dcb4c4c2bdcdb5a5449fc1
z12a0918482dba6d4c09bd42e2162c8ac295168c83038c3caea74b245989b7b03ccd022ecf80895
z76e4bbd9bb983f9ba105ddb90cc41b78fa7b372a34592757c3482866e12c0e6854580c97dde68a
z302cf8fa297a988e5ad27fc2f98e9c1d7b587c3a39595e9671ff825b588b3e9624760a35fe519e
z408b4b0651f3fecaaaf1749a3fcf18443a011f9653a8c22c68d34efef19a9ce38b1418d4a27b82
z0aeff5e9156aad560e1ef459c2991081460c10c1b8b2f20f74f778317b805972bb113c8da955f6
z0fa61f5dad06e6c178ed426a85423ca33f9e178855018f071357b02906a99fdeb46e379255aa73
z23b57f72e214d1a1b49f11acb4615fb4c3d09ab09ffd6fcf8cb81bb312ad443cf3658000287886
z74d1f115c925febeddfd31c27f38ab425e850ab7a04892d78dc84b334e650a29bc763a452dcc1e
z13ebb526ce53b7ad23ebc391dd8d088da2ab42f425bf55c0fc4185a489fce5e70d13db285db6b7
ze18d97eca5740dc6224a10bd206bf925224d2961d46167b1dfff64cb97f684e0ee52bacdec1c41
za4412b33e9bdf452bd716366d4d357770e32873121b136b500ac871951b033b3d25647f1921a4c
z3d3ed2f660444a4a6b14b6166e7dc4a6978eff391fd85e9126e2c87dba09507946d9f12f9d1232
zdadd6ef0cb6eeee93c229b957b8b2f0c952414d7332396a455f7a4b75369e92d025bfb92de90fc
zba1cafc6855b7d27a740eaded9c90db8821ec99589249fc614d5bd2013124cf5dc8bffa28c1ccc
zbe25b941ddfc8d734ba7c8a498a01d96d1711624677e0f3792e5a49fa6410c7c3aedb00687572b
z6faa2ca0f04126dbb0e7b364859704e84e07639bc0a6f5b42f2ce36df0648201a3c48557147a7a
zdef3f0cd58a1242a42941420337c990c0533cca65308b57804290d9ad033a47e9ac7126b9f2af3
z57ce91fb598679a7d092adc0f24d522008dc792466b5a2720aed7c00c7bb823d08259942c4f431
z1971de56cd0962b6d13d09135ce8c470c8fe3d7b2e40b80884afff4983fbe753c553f583ac1253
z039c5d483d7e83967cd48999d7152de49735bd0c7ec0d0ca69a763d09d6372116c64554216b58c
z5e1463f01e21d04407122a518103024a043f54fd8262e3f3fa9fb4822ff80d27012e5d8f4f3ab4
z76e942de15b067c8238614681a574dc8dd997ca5dc697a209d157e2c899ac103a8f3aeea0a2f56
zd01a28a36115afd25bff1ceb97339352bbf8b408ba067d92ee7e5446cda9900e52d51249d3831e
z48dd8e48957af67b12dc3d25972e404dd72236d3719e4778acf63ed2eaffb8253a817e8873d396
za27c0bf1fecf00859691fa57c5db1cd23f12e73408e12abae6c89c636e853d7d1353035f9f536b
zce1a37b2b3cb87466152de3db5737f6a0d9cca6f8debed4e13690b4de63e58220271addbc40142
za8a21735b41877c85d7dccf02c2ccee6f826c55dfbb7db944ab29e39852113c5819431a9105cb6
z39261e97c60a1a067d0bffbec1619d4dc3af53c4f90a6bd7e2e83f8d385266b8d198ba87bf04a3
z16579c25b3ab6cda86e331c1e3b1d3f425e8408e2d3d433571add377d89c7f517c8f2a660b5c79
z704990b3c985db68ccd1b8ea5b3c2f6fd685134912a290022463cfd7cb4024b54917b1b990e495
z8912d8d6656d2dfefd2d6625bf926d746487a7455d5f015d3de5262428e6711fbf8c9fb70d20d3
z87fc1a8e1011a1ddd36debb5d0d087c3ad58c3d65503f35ca9d26ee34393a96ece8e73061a23fd
z39538ef65aa4b6a935d9ad7c6c282d3a74a81d92d93e7ea72f60a830d8093154c8e6c68495b4ac
z9beb44b405aaa12414bb9dcff3be4ac3709665661c597f6e54290918a92a1098f68329de57bef9
zffa999f5ad98d57842d01cc8613b90dd7a38012eaeecd2612cc078ccb23c9c2f1f643ed5a79904
zf90550a3923639afd298308974d002747f947771a12262269aea1695006e0836638806b6bc2f11
z45696a0f91e0c6fcd5cf86c03c79dc6676d2d8e8031b763ae1f8102fc13509505bd9c88d2c4a8d
z665cc3f8f504245483b72c18f0f4414c3a754f9dbea5b829f617fa09c3da97fd1c2b5f9069baf6
zcca3a6a9424d13be822f79a43073880947feb236482cfa11d97fea825916107932149ae8abfbd9
zbf3c75e854c2c349ec7f7107d091d33a24658821a598852d4a40e54adba6637e4049fbc77dc7d7
zc8f9481f0731687649a17582aeb3ff59b7732b43997b8cf92734d3200740e01731b247544f422d
z970015588b390baf2b4dff5e529642585e3491ba050b791ab7d7a202f6134f97935ba59ea59670
zf31fd1ce1aaad161384e3e2a99beee6724beba9f7d170dc999d14cf94c00da8eb59e35b980bdeb
z67c3c0968dd628f9e94692b8ac2e0df62f26c102b75b8fc23910ee622af0f564e01dd6ab54b011
zed6692e95cc49fcc3b16818eefacf02ef20989a17f41747618c57ca9cd03df37a02c9a5a19f078
zc5ab3812ce6e4007287563d260e24e130ca7c8545fe212a520c66bce190f17ae18b75c59b7b27d
zffffae20098a58ec2a36bcf8bc84733a69f00a1bc8c1a5a516c0f8e91fc70d9c0210f5ae7c09d3
zc240212e5d049768262c67ba3c212af28d0f8f754b3cc72e7404f7ceedefe1e0a432b8b35b5bf8
z16b6735ff28c02d7d9d08c9788d07c0cfc934e2eaeef78c5aa3bccb3e9370911160e37d5b48fb9
z1d9e61617172893d67a1f04529082800fc881cf1612388ab99245e5964739d4e2c7b0cca5fcbe1
zf0ac8d30ae16fa69f8259dc8836a4dcc4de24d0ff7716f573874d0eac5b4e2f71ddd1550ea318b
zb6c7430792e5e643e8c1799ed9ee6609a6ac3e2ddb0a3bd0f17fab2c1d0cf5d165796eab0aa172
z31e36782857549c64e27e8d522013294f99ac7264bc18d89c9880c9342bb3b023c912cf3caf74f
ze4d5d435b4078900e2ec9775d56865f06764984f849f1100c26c59f04082f4526e109e7ad65660
z32264eb5e838d0a17cf1e3c02059e67467c6864cccd1ab585b8ed9ebb25c1e4dc174d4505cf369
z7cced93a81c0b302a8ba84b7aa711a19783d2b51e0f975a64851234baacc28f732b4bf441bb02d
z69dfdcd0ac2dec117ace48e12e594fdb0f8960a5a8620938a7408b42ffa1101d9d706b640e9ef5
z27d339665559dd5fa1a9d64de029493614b6a92965bb6ce34bfd836902379a2d0bb84d8e93ba15
zd797d07c5d3c3797d40b0b6ff8dbfeaa10dbd9c6b586ee32b014fc2c5c2bb369b9f14059116496
zf32663ef1e1d2093f6e0594ff57cd043e3da011f783e648757f903d114769aefeaf22e64c3a572
z1231a296c5c06ccae86182fec40389dd2478c101e87c8282b06c05b8af0a11b1c23deb82f8cbb6
z066a5e418d7c37eb7f6cbc8ddbbf0bdd40f28173680a96c3339bf3a7bf8ba66d38db768c85c2f2
z236300e5629b862d5cb646fbead98da06b37262a88c403d6c56967cb463d9aad4c125fcee21111
z3b6d454e47020a49380aeb790879b55a9bc06806573e6993e0d19293bbe12312fe2a21436ebca4
z8d5893d97fcb349aa0c9b0b3c18836e79346ca71a447b2463dbebbcf7babd1d27a2ea48f230ee3
z442141ed4f2a6e67f6c7fcfeb6b1d39f6f57dd88415144b6a41a4e07cc48a457b19812d8f25437
zb0eb9bc9a7dd2da7a6110c872bd38256227e262c96e25f72489d64135bef3be8d3034f58694bf3
zba270f27f80c02ca21c6110b369b61e9f271d460fd4fa75af71c3bd9063128ad6549fcba86b768
z433ac90f163e19fe6aa19b859680be2242908980f289207eac0c2e443d4537e8d285e890e3a39d
z74c8de0c5cad1af80d2e700be6524cb7deef2dd37d251d0862685164a5bd2b5629d5d72545824e
zaf3307e52709972ad60d0a3e24c187804a97415f6846ef0c64827f3a286df84509f96bcc8054bd
z2348840cabeb18629632fdf2b61cd7c5e699d6b095f4bfcc942ec77b92ac43d301c02f2760b690
z55d83a499abd231de9958f8d05361d12d9bfa3292545204476a04fd83fd715a76fa6b1de5a0361
z125ae35124753f53feff7e16af967c49256b36ff13a684bc273e2e4c3f6684e43455cf011464dc
z71c9f39052bb4b22690ea61a57ec24c2e32c71fd0922e189b3a5cb4b0a3d7e53caf1e6fd90b8ce
zec9d093e2a41592ef70fe4e2484efcafed2fc5f102a7d37bdb7ca2d6faeaae39af846aeff7ab7c
zcaa34dc59f2ac745820a78842b8d5b09729c8ca75ee34d1b01754dfd36b43902d230982e20ee94
z4512dd512b810871fbbe888b7ec772b61b64b5e26a587b7c9b00e28ecf7b5e67e9fcd43acfac68
z7212dde11aa8c7d571b8d5f7f6cd696f303e1537cf8747484899cf168eca48c2ca7281d8d708b5
zc24f1bf99eafffc26792e744d88f78b4dc9bef7e87e96c1a37aac1a05788d23973b856fea21c18
zaa56330b76c657a81e8dd7159845099da5e984b83ce49ca8a256520301416946f6b0ff8d9cf8d3
zd75dd1992ee143b408a8f43c2626e4e53bc5fb6924a3543250283990203f0e276b47b8fe6d2e0f
z61706b6e4b0df876bbc4a454084930df69809b40e5b3a5c0bccd6b9393c117ba14e1f141c4e8b1
z7e74fb49376c997e73feb7d92dea718501809798bd3c1f6d1252bfcbb1041a3af445e259835138
z2db3d1dfd2f5eb89a1cbcdedc4cc5516a0d0fc4240422f00f478ce07562238d97fc6600d46a3e5
z274a9327f6b376d88d983d6dfa2a5bbc6f617a903f722b8a67c76a0b472fef26d9e3a9e84619c8
z97800dda1bf8872eb5af6ef32770ae8ea4d039f14d5211f432f2830704350228a3d771c8426904
zce9b3ca42786d1186edc23f89c8d2bec1424821f36d6cc18c05ce93cc80458be655ba2d0d19e59
z0ad5d889007dfff9a9647335bf08dcc432e52a627d3d0a65fcc343fa9b129653fddcfe5c38334d
zc3e5fcf1cafb8768bf39bd267c5c39f86208626378b98c88c5bb7a9a86261dc3aaaaca2d3c7544
z18040e1d06900ec35b2800ce4d0bea5fb7ac1f8db12d937b72546c6a1a1348e94ae0289942d670
z35ea916dc65c2b9589768eae889407812d6d05faaa3e80810bda5cbd4fc39903cddedbdc44805e
z7b5b2eec393423dd57772470ccde6dccf070cc830f837b94ac548ecc25b834d57cd36f782499d6
z0c54dd17cfb26c3ee25053f87065c5873b7e6743fd2dc0a2ba64ad503378c0fed0cca75bd1fa68
za1587b365f85e0dbcb6acd77fcdb63663da0959df367a03173412a5ca7a0e758577be8fdddd612
z922887f801831bad15f5fb48f93ff2d3505186e0eeb92e5e6f03ac1dfdbcc9df6ecf8f918f52c6
z057619af92410d4b851acb98182f2d597f2da11dd256c359b0ad90e8fc46b3b427a161d810a557
ze8867992715a8885af49595c3d3b167e74fb69e28e68507ebc8e9b5894b34d0b540bf93c1f0fa1
z5d8c66e308b60e3970c190e9f47625e65b4e84d51ddef5b933798e1e0ac862b7c16815b5692a41
zcbc49c2273820b746a51159e0628e9ca6d7e8cba317b7d50ef93688e771fae8f65efd7c42bc58c
z6c4e2766c6045a5a3d8e470c1eb2ac2ff6d42b616d3f256bccf30981ab5600a61e7b8adf31d46a
za5d130f69ad30959e6674d76faf81a6f26c413a463b4e823c246b94125bf4593e945fa78b0348c
z6b91cfcc1b426572b2c21fbc4a7417d4fbaecddb301e5d548bd8df7a3304342d583b4111be96c1
z1e9fb133d8d838a5422ebf5a403b3abfd4e663a490c717e55376729bcd3d2492706ada9132cb82
z2c321072a8eb6b229d5ee518ea082729499136099e11aaa9a547b038f374e29f9676246e7fdb36
z89bf896d296f5862a46ad2c234ce6e74e876458bc85e130f1dabc7612b788e9e46bfb3bfe008ba
z2f396a3860ed7cf29e81965f1926f1995fa1212a423c1fdab87953605838afb56d1383356ff4a1
ze63b832ad2d15c43fe6aa035858bf85004e1a924bdd4e326c0a9810a1e782117b6abf7cae7c6e2
z96755f05cb80d2fa223589b0f4bddbcada13e5534a63c0ce23ebceb67e485c94ef75676dc6ff04
z22bfe234126892319f60d4552a9944e258a31bb4bc0604ab0b1bdf2cd3bbc8ef7676e40ef7dead
z62120c0e588c54790f8bc4c381bed592de821e3d2adc944435a87add5f6620bcc435f1d3a1086b
zbac90df0fc8abae87084bd7820649d0259ea7b39fb14519a9c5575192c70379c8919db9de865be
z1551b9b27970e340b5847c1887b8413a2128de3b0135fb1784ee7f8a43b935ae4e5277ea83c31b
z1083a1f7f0f5448d7612d18ba490572e7b743fe173ba19ae1ec3ba1f03ff1bfd4a5bbd034f1853
zf951723003e5d8b088a1d77e3bdf5fa015c24d1c60a865b19e89ec9ce1822bbb78da119a10f2f2
z4ea42b448851f11b2843e3807075d76270ff982f735f57d97ca31144c27137c48c61552ccb6eaf
z3067544e0d39855f27afc90eadbca141e5099f2424cfc2d8f41ad0a39be1dcc7f286c130456841
z17a49fbff959a20bb4054149180bd6339c3572c159729c82d7873c99f63869ba48c71c720a079e
z491e96cb21d9f9914485c35a6883fcd55118695ee62bde6f12c1a2e22b7c488a4adfad1e515dd6
z7089122feb7a4f0d22ab731fc5081c4a4f62f8ee6c668c829ea5e4ba41ab4c22d6c01f3d3505fe
zc361580b4335f14e2834d0f321110dba793196e5fa06f3558883c1eda63a6e4a7c682309fb9945
z5f789570e4843d95e0971db8d2ba92ed9ed1a5ab8ad4477d187b6a55bc21720765785d8372d8c9
z5f56a664351a99ba922074b48659a6fa58090017ddd5e0fe126f328ccaab6a112332082e401725
z82aa9f99f2780597d5f4c6cf98eb06ed2711f13745e72bf78e35e30a825fa64383d121f33d6395
z279e4a38c034fa533accc76ced17de4c3c0496615f5f54fd19d949e164ca1ba3e4add33ce0507c
z76fea2d7bec6d67b027d3171146406db7ac60e51211972435fabbe42cb62a881af8846bdd8af2a
z523288a13f8c17738a4bb1bb6a46b81d06968f4af391b6e3407effc3b859005e2c281a339ffffa
z8f2b967ea19dedd6f12e4287b5c25dfaa1f204c8fd170fe3d9a95a72b56d2498dd34d57dfb72d4
za2082a4b656b45a3335055a9a435005dea1a6ec2ff8b648c3a0ff7c6c5b5070fca73e52366e1bd
zbb26c5bbe52a0535d36bbe368a605fe993d8ef8b752f9609b23fd4c99837980f1b3bc83ddeb81e
za22c961ea0ca563a81e30a8c899de232321d96b47e44f414a6c2da84c57dcab3ef29bffb71401e
z8d9838ee24633127d03a731849eb3c33bdf9f9440b388d936826db910f931b76ec53cb2e6d523b
z6c8e0c918b5513fb6c1133046328ba81e70b299de9682b87934b1b9eb248555fb488a61d763fe1
z55092c10bae52ea6faf052f3c4d782dc9846a1281cb55729e30838246ac0fd1097e0122ef58f49
z82ff3c8369211364d4ef42ba526a6b16e425137fdc8eb3acda71fb645ec00a3a2aebcbbe6908fa
za47119e143a0bbd24fac32163d113375c88e58fc5b3552b9e8dc79f013bfa9d0e92761c93f19a6
z1540c96a5c3293823514dbcaba62ea74208b6a9c053ab26bb4ed7e7918ecc0cf149eeeb0862462
z70fa4c5d72580353cf5b223cbd6f82cbbb56753039a77fa97ce1e6c686c295bf0fe1053fcdfb8a
z9092eb618c9e825cfac8c1ef25dac5ec42d14abce37f3a314008dcf770920a1e267d8340bf9e86
z836e9d32fc2fadfb075e1bf016ff682b9771310a473299c11ed1a354a2490f2f2c394da17ca713
z153ce4663b2da07244c4dbee14f6a50de1df1341a7572cf313ce5245acd1b46bae1d8a20c336b0
zecbf74453abc9b65a7629f7076113562f2bcc395541627d3389145d7b2da73b95fbae6f8fb8fc2
ze30598ef1d8d58aac8b46aba0fc195fb5320d057193272bcafd3cbe8e7db4e43e1e18fe9f5a42b
z2560247983ca75c0c85d1643dc8dc6a7d485f738997ab46c9d5df43d5fad10fa969e1c77b627d7
z1046fc6fb79e7f9104c9f8608b6906f5b55b8eb55f95c27acb133332030e5597501f89eb01b06a
z1605b129d39ffdcd720883df9c826018517cf9be531df42e9ae427ea2856b68a08f0fd2ae03c11
z8d82f7b33a8080d844de62ffcee9ff684a97bbd5e5033f062ab5b56fe328593ff1cdba759f2000
z5b503c339c1efe14b8dc7b76dae1ad193b624f07cf0d5f96528847ae5b92d44800313c17f9cc9a
z7d4adb4df2b081de2d63b7086e502a77457d1e6ef43769b71a2650e125e6f9b621eab54da2f793
zd35c2c7c7b1fb6bd2cbbf4b1d06277cd833206bb98eca1496b9dc3f22c17227c4e0672d1cb7d81
z7d4500f58ee92aed5377989594c714de3aade19b6f56b321d8ba8d180199d9fb73d019af259742
z811e3e6c91042b2c350b3b133999b1371838882527c4c1347f36cbc107f5631bced268d29c1f38
z198f84313d3110b2163bb831b938aded475a5718cfb737792f1094e936015485bc1e079e8b6a71
z7a0e8b82c1a0f468e12395fb14764a85e916c7e8ec2edcd7aecc657e5f8991be3ce0edd4ee645e
z1f200e5ea6840378af1c8475bfc36ce6da079742b2d2c88e1406bd7578abc16c73c31789041cc4
z353c69c41d687dbd10455e6cba37094a2645d7074670b198195fe31b8f71a7b3f97a69bbcafcea
z03dc13c901f7df13ea6cc6e9f30472b803cb9201aae8984a505ab8725d96c2eb75c81c1a3734da
zaa07839de9994203204f004eac0d1e5996aad93d719357d7a1abdb05bc75848badcd5d20a09762
zf40f5f62fe640e3e69f719c6ee12cdd4945a8ffb88bd217a23328bd9d0d9642d463dbc75068957
zf2ff1ba03451e588d3efd8244099fe714e9b5255bac2d456b65dda6f5fd7554aa9453f47137559
zb4eed8e29c69edc88c1299378edc7b443b94df61d57ef58f5417e3a8fd755a1b699487a607f654
zec861f5ff855f7148eeeac6d5453d6e112b27df9b8150d59e05e6f8dd558337b6e62c6336a75cd
z2f7001ae507eb1162d31eb693859da671bda7320f91ec0fec729fe1d9a1aa9bd989d0ffb1ded56
ze9584202907c08c695ff5d8bd3dc8baa5192517f86bc8992662b43814314196dea8cdac9741af4
z3f62a31f812db424a878c0a0847521f011db26c72fff25842ed46d226bd00fadd276f92a134b67
zbdcc2bde71db6ac93e580d93d9b9f773d1d04af1062a05d16c944ce031cb71083853e440db4ef7
z79a484b0fff7581d671545ad904364397e7fa70c73781038d7d27e9585ce5cf4e436ec0f4eb3ad
z1e0bfe886c44f857617f9aba0642fb0317c5a88e8874d757014690033502bed1b9031d7d7ec817
z6486f51263f54de1607e2a8d6bcd4f8b3adf101af9186d6a6e04398b85448ef04e0cf863ca7c3b
z9182024cfa7726b525a5c20422430a861b6a526ee29f775583fc1049b9fcaf9ccd0e216ff10999
z2a9c1a62d8fe3f3cba8ed216d303fe509d58df710a6de2976b3311727be7f99d2700086565a198
z8364b26976de4aeede50a986ecc00bcfe22adf0a6a848f9021178d0265b5ced99bc7b757275057
z320d40196d97fa8df155238dab1c8a9d28d866cea08a49b1e3bc54f0f92e7d45c1e0a694d79c21
zf6ba1a3bb4255300fb35527e090b488677993982c24874e050a555018cb0dc39dd05ed8df892bd
zd160c5d77a9aeac186a5d113c84daac4683e909a9d62c2acc93ebdb3eec1e9a7d598ce8fec5698
z0b9b28a0a5540c8145fbe62de248a8ce390130ec6f3659add34f6096dafa1e0b0f890f877fd2b1
z7f2c1577e0bf91e6c769d9d678e10df211d114d54b87af116d5d5f218c2dd9890e86f68d65fd42
z34e5b275375d886ca49b657ff86991fedf363863e79d50df5ee343ac2cb23ad6fe887846a48ec4
z1b1e57a1583e56f25d6a591aa2ae7ac7af0ee21e30478f9301de959cac04341ed4b1476d3f6848
z26e1c2e763f2f84c895013ad507c5a972425b2ac8f91ebe89724cf8a8cd77c6e12d484d9bc6845
zbe3ace383e4977517aa592c09f184c69a176e60b068f85705e7ed2e28b30b3597b559f9623fe71
z73405f452931750228625362f35c6c4c1fab4f063023c60e3a6ecdd36931b6142f3aae7c06e968
z8969aca7e9f34088980fa9b0daf0a4e0fca4e367fa691863853485a0730e901fc428f2c60a5406
z00c65b65816a00f483188bd2df75efde440a33f8cce297923e2f274023635dbc24ef8889d45709
z6b1577f6e6b4e224097602c426fb6c8fdb5f1a256664842ee9f4a432ce0df40260cb9d944b56b8
z103defcc27253b419d5e539ca314e723d1b427db8e97c8f11afcab51610624a9173290bb251e9a
zb356aaa7eb1d5b4fd2bad43bb07caf2889a7ea2e91f79e77a169e9727a2caf4825e79a60023122
zd5c10b69b534e911b0e47c5d0c8b269cce0730456721603e8c2d62acae2619e76264236e0a5860
z1ebb4c770b88eadff3413dab2b8b3de0d75fd9dc902ce9a2817ae300129b9f787a491ee5cdfd53
z134e7a5292c9ff8eb03f02e48855d9290bbe8558d250be1b6524a95e4906cc6c4cfb4125db448c
z24946cd96cb45927be38660b60633e6d77301d2f69669c843e1ce97b66cba97d0a917c7ec852ad
z66f9e96d0ccd6087ff59eaa5f70e9a3238a5c2bba60f4aaf3b7c429f593076c4c2be488aadef65
z901f59d3e3f20f2389aac7915a0635ca21ba0886b251fa4e7f59ef875fe3d7210c5dfa5cfe7d49
zd432bda98cd42679f4033761360d1c94cb5df94c8d56a15b10e1233df4f6a76451e8a55cbd0125
zb113d6edebe597619f0adcf998753b8aa351f1b4f0fe68d9f0800256b659b7b3eda2c11188859d
z06607fe27db43915b799b55b8542db698cf330a246b750c2d99600426051f6b8a9435fda88ddd1
z206b021a1b91b6dc22d34f7bd9796618427c80233bdd2590f95cc2b2e6c84227c494a83b2d5288
z2f67fcea0f710e2459dc2ec3c1a4d367ba06fb10db82e41e201a276d2ed089ba34496d5245daa6
zb3933e36fc2e90e2f770a53f7120db22a9447353e07458eba7449d8d720753b0779438857a0a33
z95424f79ea4bd8cfc6104c89fa8d467d633b28a02719e05095be5b59f40cee75119d58491bf970
zb53d0f734d9ee9c56653a655f3a57bc8f436deda82765d9a2db80a376899af792fc85fe977003c
z3998896c75804474ae94096015f110bbe3fbb284620953db784efc53fa5f071d29266f743779a7
z5222eb24de0f84a1ad1fe85f8c5f59429def6321eb7f5dc3400070da5fab22a721852cc18b9722
z9d0a44acb350f0a8c268df554ca5692142725917459f691797110754b4d928877388de5daa640c
z5245b68cd3baeeb73e93d1f808d772d86a613db0393717685915638a365b0c944bd8463b5d8594
z413e3952b11a013b4a055b8587cb9e90aeccb22197c145c0bddc9beec63a72ae61ea9c3ab4168b
zec864da09ecbdc9cd58b6b4d91ceb92c836bb1d7ef4b03ccce8085fff144ae7e06312f58319aae
z51da1b50e0f907769cbd7a5718dc3aea033396f8da7215cf5a290fc44339b269181a413f38550c
z721baf3260123ebab39208a6b8cc46af83b5d1536f1d8f9a6ec356582260abb3e3c04b4f45260d
zff866b379d53503df3b0dd49453fa8b474e1a9739f2cdd5ee4f3ae098fc6038e49060c4c636821
z9eb5c5e0a5b25e180842bfc4e2e16af16d08bd24defc3870d529f97024fe98c25bc07d09bbfde4
z0aea14dbe825b36fa3513076f55e280cde4481b204e652574152fbd3aeed773b0ddf8080207580
ze8d4a5bb431c40edb3f284633ae332703ca30dba9e5a6aaa951c7a4c8c5c2dd05ed2b5dbc33d61
za75f5e39da7fe15c4d9c4143aa0c74f438cb462486e04c2dc8f243ff09fecdb3606bd399d9a944
z859470773121c3b89a6eafa1872199dd93bdb571de25d777bdeeb2d1c0838b8fda29c949619b00
zbf82e2460dea3fff83ea1d89b7a3a81e454036e8b6bb9ca1bae49d967d618153ad585d05aed1b2
z901094bfa097640f2c10ae0757038494cd54dab767757b3712bb97e75ef0ba8f04ffc29d9303f6
zcecf93d36fe3bcd1eeb66c68525bf8fd80689cbd612625100ccbd93f72eff41f1b42573f0d7285
zd7273004dfd9f0074369ecff194e707581c570b9f69841bd07cfd0f8d6e2702c4b50dbb720f304
z53cef4023ae30129f698f104e0b1277aec232bbb7eb0f6b574ad0eb2dd8712eae6a30ea5ee21ea
ze8ddd15ccc5dd8cf1995ac6d2bcd91919282aa5539b00d5ce66b7aa3010ed65959b7391ace52e0
z3c012eb5fda18124a498c6bfc52f7b3c5289dce704e97055b0121d4692adc89ef168f70f22fcb2
z22b61f9087e6b72bfa2081617ee802fe8864fd4a901a79f967a388132b90592aadaa4408abe4b3
zb07d2a48a2b4ecd8c934e8033198eeeaedd7025a680ea20f8a36f510505ea149d00aa43fbfcb16
z8cbab30d4b7b769e8137df6dc2cb52e2efab41403403788d0eca2832b4f8cf3aa1266618de0251
z7b78c3b417c30a3e5a5e17ded939fe003057b4549b9fd5c1707b202faebf9fbccb31f5d04df1d6
z0808a09ca75bd9aacafd6a3881af78946036c0402fe955f29bedb99ad1d2a752dfa674554edcb1
z983a95d8617e8c21ec2d80a8f1d6f7a1f91da5016b55c4e432d433da84ae32ce4511334e951dd6
z8472d7666b50402f52abe9228867e4a40ef1b5976b8763fa392c40f5a2cfb4ecbfeacf23d6bcce
z08b8329bbbbc20eb3db80ed2015852bce0af0e98b009f3f77b38ac35038814e9950adb6b1b25b8
z564e6b4fcd8c879ebc97344f7a2e3c3986f58bbc4e1ff87e2ae0adfb70c4eb63ce05642c515ea0
z649c0ca16b28f757ef729865428eafefd77d5ddf0e2cfbd99053c793291cb786f655de5f8a6f26
z9ff096acb2f5c2093654369726a26b122574a59c815e5c7f3c94e83b60af3b57c4d1c851594e27
zdd03d9ebaa486879d2c55b322f7efb92eb2112eb43345f0682a478a4fd77e7c9622651b14cb175
z63167d05a56f2b74866bf4088c19655b4c2fae6b9431732c0bac96826288d9ae79750e74aaf237
z0e62f254a124d111b318e816239419e29c8befbff75ebcdd1ca0004506138e9ff625eb01148a45
z2a88562e103e2c6bdd45f8d292d65b7e2a5826804e7938c3a7334f36e18671fc0d8e8addee7f25
z8440f63cff05b99f577c69b40278dbb0957fb7a703c0d312d2d5cdffedbb5c07b545e639d061f3
zc795d017cb0165890579dc82bd2ae12d0be5787b92133dd6410e5365eef475fbbb1849cffb945a
zdffeb1e6d25e35c4bf05b84c6cbebc6e2b39c032ce73c0673f3dae9ffb766912a0e97cef0a8537
ze0e2933c414403accb272ba8bced121320fac3ea573b3349d1fb0003c7de6eb4696f39a5a5c688
z06b3e9b91d9b11b0a9cb7d75cd983359258b2b27d49aa3397b4dd81c6931ceed2d8cde2b1952dc
zeddeb9187aa3a1302d180da5046dc6d0267f47cedad43308825b36a74c3c3b943bfb49a286c593
z4eba6971bd16acc6e6bedac1b6aa4bdf9304c86a651d7d40808caed7bb025777f5069e2865f2ab
zc581da339f51b68c6f066ddd62017c1736914f139871410e2ab3c3e03b4219c260c347b7066736
z0b4927a331225613bcdb70c2e023babe0bb91fea84d48831fb3b7c51b247736e29c236d3fced3e
z02462b088bd6d5025aec9d760db6f0a4bb3b5285894328a59bee9fbf8d1cb8c629706640df2abe
z509330b6b1caf37f05c5857c6a2409c74ac6ce7f4373791e7383856f5e98ad3efcf5854f61da3d
z528c040a187d1e3f7dce3e36c4037b3f50a118628919fbf5c4557154156864f2bfa6f38845ade8
z718ff0a8daa3a81a45f9215d4402c56b965d86ec426a6b1c35f586c12493eb323e8192a57f667f
z2131586228afa59be778f063f03d3f9f081cf57e30252c0b13c5f1d26d5392124c28c19ef2e040
z757a705ca731f0d580cf6f50cc59935b6e95788f84e2453bf8de838ecddf7f54a52ecae1d69793
ze463bfacc649d96cc9cc9ba8d63af06ab71967546f696d2cd5a0b66085188db9aae6cd526cc702
z4390d1ba56bb5b0f170dd680eccd1f8044672d6d5ffa1ffa696ff3f6495d0b3dc0933222a996df
zd79d80bc7d5f80fe4cfab36fecb0c2a67baaf8b0d6125eee7d170e0cc0f674ed4bd7ddf9b2a94c
z31fbb1c6024eb063f1396ec0de53f168821409bc56c7086828aae8f1609e0590c098d435ae33ef
z92ce41e5e21054417f215be47be689d847709a8820288276249056dfb31e46ed7a37ea9d9e43cb
zd3d7f478b280d855181ffc5365633f51277d6f10882e61ad75f6fa421762ed21cca7bf29e2515d
zdf53cbbe4bcc6c36255a8c3b6955d5a6dcfbea526349f185a21fcb6b4d7c0993060b15c8a6b767
z178f97311dbd2c62f7fb00fd5e69929d91c97f56c859dd53361de62b2614e1126d0a78e825f0b7
zc360dbbb0ffea9201c2527a4a95ee2d3f6e06e3b2860e40311142ef3c26bf09a9df06caff8b316
z2708756bfcd804b8b7886ccd20f0c0c7ef2209421d725237beb3a90a5b7f62f68888d59fd5baa4
z8f8c13a61381716f45fe5f5e2610f8f53dc479864a59c6fcb06c4077700b0ce6fb83eaf30d4cb8
z6595e9417a5185c052ca2976b4322776e76acd5d5a0df63627eb105dee6d5e507f5063258c9f6f
z1f27b3a010cc8785a2f4a6bc22e4311f3503e4cac71f60926fc9b29408849ad5e6fc71ce2bf468
za59d611f4ea4535139943669634b909cb3bf7a5b733ebf6314319c6194723ee8892c096201f471
z05e0493ce734badb105e0689af7033c9d5cae2c64a6547f7e7fb340b4ac9040ef4658afaac1bd5
z47dbc732b824deb3ffb389be0c4e182b2f3becd7490fa183ae97c83501ed6b22492f6e74923925
z42a3ee021eaffdc7ff1780278107f7f49cc20b27b10e5cd49140eb96eab824a68b85d6bb99853e
z5183b58813e3f7d520d3a9609e69ce687553534e959ca3b3c9c8f56a7e8742f0fea7c1b264dc78
z63a291e169b6267c465942a68f5ee7cc1c7d2ed21be6338e5f0fb8f12c6af69d4681e43a1f6dab
zdea3d897b234cc098e4027ff58a6fb849d48eb7ccd771df52753ec768724258491257cd7ee52da
z303b11621b9d813464d80e19e6a2f89b33ece3f8d6bae3a9cf9ff33ef666310513f0202f89e181
za6a9e51eaedd890d154e944e685852f5c47035d51d1f096fbef6a523d3833a36041b5f8a852ec6
z398e80e88c87d5bda071f35820795fbf13c1076ab09f7ee3547e6df37f4f124f7139037fe3c387
z6a08dbc424012e6bef177920111e0760f68fd9170f6d1cec2ca4a62822cf8c39afe922f053538f
z15d4d2787bdeaab488413e9de68073820ada27f52aedfbbd03ac83e349bb7c55284ad8a0d90c6b
zca86639620acd78554fd34507cd0bc548a811775bd6521761ebebf544bc61e379458a100a77476
zef413d9e1ce0054d15342f5f0c90e7f7038b6f41b39ac802566932283a870db6276fc8a1dab69e
zcba2912ba55f3898ce69f13dab58d7a7e9bbca9c45c797524efbcd0e62db28960f1c7f8f72e6f4
z50241773bf58a4094ce7ed7d22d5955e3d42e67b9dc844cf683e3f0dea68bb60ab72251a78a63f
zd372d1df8b462e2d30b0529bf8498bdb6419e5c950a8c7246001caf6b3f50d7d492ab807c2991a
z97f397553a590d9f4e84e7a03080c418f2bec98658efbabd0018f3ca4978ac91da6cf129bbc02c
z36254e7eb214553eb783949f71c0c8fdd5d9864fcf73bcf079a7474fba112492c866069033e6c9
zc32973532b13cdec6aa9dc0a670462271b73651b870f40a2e93f806a50466cc46d0ba4fe7de00f
za028782b9e153634ffdd370fc592203fc23609c4d23232760c2382398df2d77a4060d272de0d2d
zb0594b9cc8bffabc98a76f51f508d8c132295819f3cb5dfe3bcba3c69fe04e150d67dbe5269503
z55b442aaccf48753c458e710068d2899ed108c3719d9297ef803d7a4f7a751449eabe70ce32329
z25ae2432928e6eec2ef6844f4b0c39c976d98c57ce1120c94e2f8ffbb47a5c2112ce51ab934edb
ze5420199cf219b1580100d1bb46a4e395002ffd4be9a54285f8a7ef45eba89a1af207b587df841
zd4904fed2c502961774916959b7a1d7b84a301d6e486f91dce139d842f6af18cf35f16cf371fa9
z09b7f8caaff2d0c25e8ed65e53b2f5fc730f8cdadda27b85487d79ab8dddc548c2fb85cce2aaf7
z15bd97b06ebd884f6cdbdec22fdf7cc817de0d75624eb6637f1b5deeb51dfc278a63ac5331b183
z7f061926e70b2ffb121b61a30197ec3467230c3a944684f9d87111c8b695fe3b72c6249cd6f876
z94079555328882ea572792239b1870b68024982ce2e8e6a8bb5d820ace43f2ada334a3aed9eece
z9691901e22d70b6b1f28d82a9e9c7e8f868303f2ee1b240bf347ec941344153aa7fb6a1c925e8e
z7d3e3ad6d50eaae89f02ee323ba8c55b708b72b029e7146320c94ff19a636c24797cb9d35326f5
zebae05d22ca36f2b0024b65f599f77bbd9785d17d24dd8f5ece6076baa55a98dcaf7607d5efb43
z52758441876b18b73a4ac893742711dc3ba6354ecb132a066ed57e689fef084ee9c632290d01eb
zcee40c9d188a03421f2c52979abab5ceb471c239bd3047122667f17183a3ca89c5590f85ab1fb1
zb08edcdfe72a03724b1fb67bc9afd04698d72a198745768b5368fe8cf1edd00aed2636259d985a
za06f3e9c9d1a6df7cc7907e25eec480783cca57eafe976e6b1b81f8225848563eb0ef3bba429bf
z73c5d4ee18901e3470c179c91bc6a9023319e2617f9dc3e460813bd3b230d660b58df6494defd4
zb3125ff4d6653d0ab22326e8834b8d23c167ba8107165445eb5ca8d605f39aca02ae27610a1666
z4af095fe94712d60442faa251b055ca969a0947f81670ba2c7becbbc8ca1714358e26c0e63baeb
z03e1e998d96dd00a3fe3cafc9e66b68289b07acdb9e528c3d6678cb864c438658a267690d22b55
z94141e8f9c54516e779208c53e975fe31dee36de354ece56de13aa38391ca92272b3f3be66a6ac
zfbf77ddc7ee8de867651ef9fb1abd9f40ff5053009afb5402f12a815c9cfacd4d8959a9fdff627
zcf3996cba77c6e19883e3ed4cf1e827e243a6177bc4343cc2da619fab4ef86db1ee38a92cc3d13
z78a1fd0f3b00c4e18a18e7742018b329d41fad50d05956e394cb632be2b279727936d3d3d4064c
zd2f87ef27366170b73ade4d6e6aff6929615128ee648e520bb1b8e03d399192e0a524ab4430aab
z994a2deae25b69169bf0740efd07444c842e890cae5bafcd97b167f109c863597245a343912445
ze5d9ce443968e88fb272e5f7910056be091c8ebbe1e72f254c12aa84b8059b920cf6734415416b
za13d3e873ef1dccf034e0fee1f74a6e733e9da8da82871944338bf055e527af81d7e958ba29bdd
zd7f751ab9c1c4652465d00eace5d71980da441ccb77b209a8e98c932281f4d8c88688f5803e3fe
zbe29aa4c694070b4ab6e9e92168a9335acdd10dfa968aab7dc43240639dc72e4389af1bbcec105
z385fa41fb1d9119a7951a399b0bed6de6a6c6d387d4435b9c60e948e88affa6a2d405857bfab33
z271413613c98cbfe6f290433d3eed9ec2c2f8bad866234142044f8c587ed6d01e28b1a30c7a5ec
z9a56767a80bded63ae25e763424d2854143acedbf76d6e5a5527f7bae031417b9d4b54a348b99f
z28150fe057e159e1afa0d9b411319fa6c659c167cfc4c42464a5e742a2a57877eecf0578513512
z586bd2b6077c0fde6984d4bbd8ebbb4d3104bbb97ab1ab2dfa2788d3da202cb53e779ee236d73b
z9ee0e2c1f43c34761d710c75a8b712ce9235f4a720a337043a4dbba5bc8d4f567272c023b001af
z450d0c232e6224ddba4f57086713925c5081a0e424ff34d9e4a408d25eb3d13eee3caf6df55013
z327ea08b66821fe1216206e0ead327cacf1668f7c90bf60ec6fcda1c931840bd5e9d13856cdc82
z4ac73d4325477bc921a1376cbd3583312513f1521fe6b0bc206c4c45d0bc4f30ac3ce53bb421fb
zd6d51c0f47ce5e41ddc003b6616c776a4b99bf0b694686d1f3dbbcbb3f5be7e6f4b7075d5a188f
z16d621dbbf7401ce3217ad7ba9fb721c1d7386e2afdc7fafd5a1f8031b595b4674147f0d5d0173
z5d01246db12e1bcacedf5509efbb4cc3d0db650f9dd970129d78595b86c05b3509d0e0da5e3d02
z1564100b3c96fd4e0f19addae586aaf89bce416387330cedcdae680308076ab30d794dca0cc958
z44400e75c76293d8b4a35b564c07866363b45e49e59740f77785c97dc111b702b5a0e73d838e53
z33ba1a629e4e75d2ce265537743e0e9cbe8f44ea5a6e1880e6b64a8527647ff41a1e58e1bc0715
z777f817d9aca53fea8b785cd2540e8808175d1b0e620037a87fdddb8f9ebe4cc49e17afb797d0a
z73e5ac92ef1e240966fdbbb0b172e8a2fb5d33a1629bf16f5f9e9cb794a645fae0124bd007ac21
z0fcf8d6c74fedd6927d6877470e6224282b9197758ce20c6d6d0f0da04b8f753339210204ee4d0
z0a2120c174e8180ee2222a97d63b3d5f5d62de463b08c3ef94b17c7093d4daaa601a8fc75e901b
za5a68403d0622b8be83fb863cee2d4d092c0fb83f27d7714e2eb744aae71666b67761173a48213
z99b189a43c4c2981df0de15cc3439ce63fb88f5ee9eb8a541d991113668d1a919770e1cedccf7d
z100660331f96d1ab80284edc59a25937a7d89172eb06916cda42af0881f48af2c990fd18cb39a2
z0faded46573605ef3e971c8664926e067f662234fa8c2829449aa21e4f1aa6b0cad173713f3ccc
zdf3d54dfae7d769689aeefdd86e5c56f2ad19f5b42957ef248a30d0abb4c506669ef84e0feef87
z71437f1125f6d6e3e9119c47de6b52d15d39a4a024dd61142e9627fa118e9d9a0d07b0cd351d3d
z88692fe7f3913bca399e4f667bfef121867906878e871e6a031040a7f24a73e2d05ca1520f0240
z1df7aaf73f681c46e4146552a8b964e19f247767f2815fba43a8fc982c70076df7850818cef973
z8cbbfa9506bf762070cbd13f0f800a8e6d4c84e626476cea19e95bff2893889cd3e449ab9430c4
za50d47774bdaa8c66a667706389ff1a3767eceef6da167524c8a0dab795286696b6af0125f9c2d
zb78bab7d899bd4c14791f4b56888120d19eb7e75e3d20aac5852d1ee573b41cce0dc17dee77227
z49b834da55a6c8094462ecb022fe75ea7f91a11fb25f2fd91f397b045b5395a6a0e10024e1de13
zb886d151cdc974b6bdcadb58806db8fec64acfea804f37d83b0a4921c304de12769ce991921d6d
z1a1a7292fa51d4bc5d9fd2c2f6f932d9b0f7015e585d3932ded57fa21d0a1ac506264564d4995c
zae945b48c8f3ed6988c6cc20ece15652faddd523cbc653543433117b57443412afe6f2ba42015b
zf69e43337e02d04c9091ae4dd591819757839340f0d566317054919f3e69979b1d988d806a479b
ze79cad9f2856e559b888aabef0ace7a2079fe2ec1d2dbf9caa5efc3fdb853acd02bd4062b8b30f
zb20f5c93c5cc0f6e11c5a7e60ee2cbe561728eebd79361bda002692d4362d8fc76cfe852dd87db
zd81c3ba656c061d62d52b643e64dc2444fc6a4649dbe16c1668be8f971f8cd0ded294523972a27
z85ce91d2908e50d7412d9d27fab4f597c202fab5c619fc7becf1f30fbaf6fc1efc5bedf49cf6be
zec70bf0609b0c2981ba77ae68087bede22db9cf389d5ee76cdc0e52974bd82e9823bee4f216058
z6ab090f77a1d5dc69d3a24fa680f0470d81bef581506ff42cfe8389ae427eb427540bc3fc7826c
zcaa86fd5345334d7346777e42b6cbb9160a992fd046f96cbd9fff2db017eb229b8936f396939ac
zb559fea0fd5e79453bc6eecc60e906c02e3e3b939ab6c8b0e5097242af3f15f04df9699b1aae24
za2979234335fcfa8abfe900c6d1c1f4611700c2ac7f43aa48a51cc94fed5c16fb95ef995df17c7
z5ec368fd33d7101d95e79d6f3834c02d88ceeff0268cabaa94c6984a0a6407c79c3f293bda3473
z39cde2f89b25799831a71b2ff5f63919f20114a3857e8b71bc7965ef93f5408f28f2bdf53267f6
zf556df0a148966cebe3507c31452ca9861038da4c04dfaa9c03dd2dc955f52bc0add680f2a8062
z2e78f6734f308c63137099e6428cd1729c793b6ef91cf5c9cda0261b1d22438bebdf72003b7d53
z0f0cce71a1deec6b9cd5cf9fdf8ca8f4bad192bf08f83fa4b12664705fac57085bb01923f48bd2
z9ef7ac6a2f899d2060289182176f5794333594f4e3695cf305c3b040cc64f8e5a21039695a3893
zf58a099784de17d24644b52c098b680ce5bba20cb7b5ea7f84e72a07ff758c03463787ea58d9e1
z0e2c31597eef2852936c8657173caa0cc3552f51d01dc52ddaa7d29c59e80b288cf8c901b37fe8
z5d85acbb7d3966c910e0ff46121834945fa550f1dd7b5c0b4e3c1e1637c0ef0393ea4cce9cf03b
ze9fe66356347982b73735fb15c7f74a36faf0d8a71177c1f43553b38daa8bfdfed7cc35fdfa9d0
zd70c0dfee7b9eeb9c120eec19c96c65db329a5e4b115641dcbbafe51ad7ea618be90cc2f988e1f
z08f7ea396e13fefde4f5a3c5385d1cc158c879f52096c8baa8d3e0d4347b2b269490a7df293e2e
z2b613943f7b440244b4580d1472964e22bc3c00a5f42df98e31172144ba6294ec8881781944f21
z82a81356ae6f41df5b3af9f115263ca975c5a7fcd865a9216fbe92478ec23f371b9023f2517bf4
zaa896b14c491904c68e23576000fc5a2859b74d3ca458abfb3de294ae1f3c09badf1024acc4137
ze8153931070ff36873a694d4034e40c8a4ca18f801420fe5603059d1f9c1aee43dfbda2698a8ae
z86639b0faa06cc1b2a7e57ea6cd81d3bee37f4e7ee012ad2a5984d63d3c5c782edafda73f129ed
ze2fd4cfc4db3cd964673d1d5228fa2d8bede92501d9f91c709c9b3ffac68c47a82c2c8cf04e5c2
z3dcc255c8292d36bd2007f182fa27aa0500e0c675273e1de66d77ae0699b531de291cd00499b3a
z581b6c1660331268de6febf308a3bcffa5eb453238c7639a24a672e5b00d581b587ba7330efab4
za557f5ea58a7d3ac8547aa1b8a6dea2a998446d1ce0bbbe462ddf84eeb6eb8870f1e99c1895426
z5fb18a0703ee1bbdbb220084c3fdf9461d51bb702410c569fbda6131703506878f8deebaf8db8b
z668a990a24b410f96468bae3b05aefd7fe91483e3dfd95dec2c1ebce8966f692788a9f5efeaed1
zd472ee167caedba7b771ca7be017e8ae4367e8abf18a7578b9490c00c4b149d1ceb62c6590d258
z0f73d218447eacb47da51cded2b548c9a191c9e6e140500b6c54c967f0203706aefd2ff12199ee
z93699618f7291345de56233ca8c250bca9816e70e2bc681c5880e6fadf042634eb806feea909f5
z6d4fe14e8913e9dc00a24deacbc3c7bf9c45c4ddede56f85901fdbca039a38209138c665f31086
z3d263a461d1bd84bd818f38acc0c30e24a324bb35ce63024077956ad2199ec0a2ab3fd5eb012fd
zfcfafc51cba3ef22408adbf1c9a2acbf2a1be35f49855568ceb8ddb0c1910c4499f3f26cbaea78
z393fffe6c53aae882de529623335b088cec213fa86d464deb9d8a370e6c7dcefb71bb3f5e26ff6
z3126f6b2d519d07593233a3de7090dfc2303b2833b97156bd39e4dbd107e24381c7a4d9ef4e638
z45ac93c4db354eb29e7be31b719dc28501f79c6565d4b5a84e85ada2fef9889bc2b386c58564e5
z7e805bc1d9ae74480286e9204cde3c99db4d363b54f8bad5f1b213b2cd3f861e634b0d08357b9e
z52698345c8838ab8dbed1aef94433bb0abd84f5b743548c464e35d78efb1c96f88037cb82ceeae
zfdec702b3cf07fd5f79e717092718171879f6bdc7b6aa8c70b76f1b9e019870eb549df7a46d200
zeb23b6973745d274bedd7ac88421e8b187b0ad0364bc54d7d9df61b8eeccd087379812cfd3c136
z2941102b6d86ab9205e8b1fdd67abed83bf7037190edb6dada78f7c33735e930eac90a10b29f58
zf85da64b5eb7b75b2eb8cf8ffd5812405050897f025a08ff264057dab8fbf3d3e65a0901270cf3
z812e13100fab1d27e6d89443197042a5d546d90d72cf985add10f5425c0aeae730dc9f0d9c2478
z5bcff7afdcb1b634330978a8b5755ee18a213723b59f1d3ee7b4995630e45c41d05b6fbb75e71b
zfbd2e3c9c6deb3df65bfd602a5cac2ddc5dd349c9999c792750d64d35da99dd176605d550dc4a1
z87fee617df28ed72d9edb685fd2cd8f1586c2b85a6f9c7f2f4138a64d832b041ca6fda38655b50
zc9cc77abfcb2bb3c9ae164e81fb556d8ed3130e9d3b4d8e6334669641575cea103cc257f2e5619
z79c3eb67fc8e82c04f526172d6b361ced482e576f106343ece214ac00d774e79121d145deebd14
ze85906fa9c9ed270581c47d46bdfc639c1b6f77ff3e377fea0b7208ac104c5c6ed92ec5de08100
zc69509fc665f79926fcceadc4274a0373eeab73acbc713801dc0eaa8cd74cce85e578f3dc94e7f
zfcdaccf4eb9b0cecbaa74d7b9164f99e7d15464a66159529d451982b40658734d1f4079d223891
z81694d89a78c590c7dd7031615813f569c764f7cf8455e5e6d4407e8c4a8c55f06c37263f8f5dd
z83908661285f4ab3c3460f0bd5cf8a2ba2a541d6790d657ed408cebf890106fa3b886d929acde4
z5752f1a3ffd34a6c7dabaa3651d51ca7584611d8e5ad1b5c33d9b22f4730048426ae34a41d6ef6
z8c62793b754343b901c5c14de336ea9a142af3dcafe03a073a5cd620b12cc496164f29e71724c0
z098233b6a8ec134f18fac94cac6228eb8a3e1d7d9821e4f054bc15f8b12705386bbf86bc8735c8
z6f229ac7b43328cfa52c76eb9e6cfe4dad109071ed10cc777fb7e831721da0b973f66ee6cc08a8
z99071f8ddbae5ddd3ad39e04543dd15a5077627d3b4a59a9f97f30eccd8e3f9483e8fb647fd919
z2e0a5d1687eb3cb0447501871dc2c5e754802b3661a6673bd509e958aa6886108683f001bcaf0f
z5b4a49013bddb22a3b5ffe8b5f262e0b84d965c6501322e22b2c4248def785501bdb49a7a09d50
z4f0c759f4ab597c915a737946dcdeb0c969617f095034eb9ea9e2b5d14c0df157ae02cf4f2fcf5
z28e82f6d106a07c9f001a714d2ce847976e1e62c5edb31ec9e1df51c106b20830308ace000c87e
z4749ba820cf732fc3ac1c0fa7d3004feda5ccc8d816ac6a71c2807c86a32344f26b4654e47a492
z078df156063d10d4c0bfeaf0df1d39ef0e1423b027a1ff0d3fe3b9c0541785df6950fa00f03560
z6c9292169ee43718e2434be64a4b6f6b718b4124fa509a1d278f5a448df270559600b68ed5f49d
z8f12386444928602d7ce0181691414edf3a51760339400e3cc3c17c08d91d927c334a88fcfd3e3
z422f9a588bd3d581eee84571c1963c6542099b455f36c8b2b54790ccf82e8a02dfa69a191b1f00
z28a1bbf29afc4b49b85112133816dc31def71e10b51b2cbb77c8103265e25ab06134bb3ba7d009
zee467c927d44e989b8e735ee2f73b01c3927216a2a1fb71a95a8950b899c1884a48b9ffeb48182
z9a9af68f7d04704f4f4889a2a24fe38bb42cf9f5db9b9e8aef0343431a51992711e350d777ada8
z18d997b31e7f964b0cb1f06fc2f1a237f26c3b47744dea388abe7a33cdee9e787191ee4367afe4
za7cb7ac5a89b8dea4e2355b6eff3421907663973f6f14e563f4347f566146fd1d75165e8a25aec
zfc070a9c814411da62c8db53b178c9fda6eefc39ead136dc5e71a8807d69ca4930198ba5dc1c47
z45fe3e57ccfa56b7eba8636ca654c4957e0d4f203c8e233964547330585a3f476aac5859db183d
z68496d2fbdd5d487e90bec9658df8a22b3f4467c34305237112a9623da34b77a3ba133b31b6d40
zf8a57cf1e2f8120ca7957a5fe71455051c5ddd45d5332a4014fb2a7157cb35c982fb2d484d9940
zdf55da2df3b1a557d5db568f11e3b332478638dad73269ae5ce15937f602c0fd1f903c4f2c83c9
zf05ca391c29bd3e22e94a012b2f41655a4e3e7410811a0e7ecc5ce8efd2d90c3c9a4d39f6607fd
zd48344fc0bdb1f39e8ae929fc7bddc3bf069b31d33dda30e5415dfdbecd79d877bd8fef9ef0aa0
zc75197219d85409d99599341871eb6a6af23948c316acd83af436fed66f21afa016a593af6d0b7
zdabf571a5dd088a375f18ffedb68d63eb0cd70a4a72eda51e9aafacd1b33b917802081e3ad75db
zeaf5020081294cbae95cf2c4dd79a168aa7279501c26c00d97cf614ee35016cd706f5a2a7c34cb
z605b4e02c090da001d2dfeeb8db95530ec0209d460fcac091354ab0c08cd5fadc883ce7a721728
z8d9423cd9387ca2a8087753e865d599ea5ca3857cdb7185199dd3afcb3608809b1f9af790a6b86
z3f2972b06a58816edb5c70c63f70dc96925561e1d44a7f7fcd844b359b6346a5b5e4cda4dced2b
z7e242a90ba682892130e98d4cf4f3dfff3852021ebd8ef0ec76b152668cb6e0c92c455d70a3abc
zb71ad191d154b2b2745ccd93c8cfe6dd2626672ef3df26ad8a762ff9ffb8cdfe41b254f382f402
zfc95246045ceab1679e14e8fd75bd14a82701198aedf20a051770e72f14a973e259b91d0a4cffa
z3f186bb62f25dceb0951528a6a2e8ab1d52fbaf517bca7311bfa382150e64e0f15d7c0b25f36f7
zb98d4366567dedbd5e294487db3d467ec8c7b1769178c00a0fda8ceedb2fb5b55c5dd2540ba6b1
z483b9b58d7109e67e3cbaee7aad59c4617d00a9a519cf5cf7dd91de8e150836e852088bce1a2a1
zcb2e0899c7c1d41d209ffee4c33b58ea0fbe1a5c662b632284cad13556a8b5f5e909f86293482f
ze41d65142c9443051d69ebf1c4231826397a8d9ba4aeeb950987e181587ddbea6e346195f86c37
z9294a50f227535fb6cb1650049fd3a76289ede268b13d6b04a490f840292f5da86f62b1e1ffc83
zfa31ce0da4b224a05845edc4f17284498dc7f019ca7d57c5a7371ea8c8072e66a1d109a3e58d00
z6f0144aa7b1bec16cd6e0dc818007db8ad7ffaefa9019ae6e9cca28f556cbe7b60948a764d4cb3
zf2794b710b70fc125839a6137d69bf82602166c0e133338e7f74187c7ad2154ad384605a4062bd
z7e0a5eadd07547371153c4338ff67a6bb8e622e946cec889d0cdc7987fd2e35e186ab8692ea918
zff956743f45f4d2fc2b4fac12470d7e8cbac6661a3df8cf01a56f0c674e9fff244e2b85bb2ba99
zf438df3035193ab1a4cf588e39a15a41bd976adc9aa149803f6399f8f08dd7ce2794f4a99b6c5b
zaae3d5a72ce37b7bf8f936110053fca6b34ec8527e85cc8f82f7d210d1239d73fddadd75cec931
zbafbdde81c47fef70817feb4e772c49a174a41cca8a329252df13488b4eb5c22f0562d0a84727e
zad4cb43954c45b15d958c386501d91535b902e70ea21db519f56350d3c051a3f2968abc47f7630
z60c571fae777d9fb1f2bff18989d2e3e0549a572327058f827d65308574ac4d8d10ff21abc7571
z20b166418aa46a3fe16e8afb774e19113e587beeba47e1f29666d85d9d459f7cd10b3a1e9b09fa
zb1df2ce2782698dee81c16400a57b2313828ee07b66abdb19767c2b31826c402a37e0a9a96c343
zec204465f71cccb73f5da20339aeca32531e97d094a7888436baf3c55a9e4a8a367f3b51f31944
z3298f5d227f541393fb3cd670ae22f5f50a82edc062e7e25479848a560e9c5e808b6e9cb2ec5cc
za76ec76e2010dcd2bcc6d6b438e041afc18d082cb5a2d52cde8a095741c65442a6c67a53ed935c
z96e40628ec1fcbf4f90c6101dc02e038b8201141f515ec1bdb7ae85b7227cf697083f2ed072363
z9e752ba9c281503ea42e402db57506f9f4bf11b9eb358286e75330a8824bb7eb0da46072961bd4
z7f5635d0749809793edade206063a8d60ccaeab075fcd24998c2dd2b6817e0979c6eb755ab80a4
z18c0192e6a1ebb4a510c4444486d8092171312665fd68991be59915e680db56fe45fd2f98bdf87
z8758949b4c364b903e32157141814b88f837d9599e0af17d5b8aac130498c488526858ef65284e
zadf4a4601c3b917f22451095b50e1a8babe4ce8cd846a9991659fabe31b30b08fd528fbeec62a2
z3bb5fff7bdeb904124b48cdd5c60c06b80e14b4277d4a650178a5903987f975480673c794aa0d1
z52480474df600d11699ea21cee815277bbfa45873c526720763d7be2d6d5333d3a59ef157a3c6f
zed209702054213e0fcc5c9067a57fc625cfc29832baf7bb83f6b714775f675db905fb087b83050
z21e28787a963db93363804f681b46ae91d18df249741096816e50b9bb505f6eb97f31b91fc7548
z0dd047c3ce9583dd0ac87a5fe02b207a1f700c6f28ca78efef83b00648f598cfcbad17438ef1d2
z0d9215e16a06504a2f01339f987b4df7b65db46953911ca4945a81055993e5099cf7b5dc57e2e2
zae78333330873f0bd047630774e97d663b83d151f238170d6d035d08e4fc03164f0d02985e1984
z87226bf624f3030be7dc7a3274f71a3355df621eb7d226bd87f74c95f6a81d7389982b92dfcffa
z3424f1d55d68155d34c568cd69e961fe51c50557ce9c2deea8bb4354c3c5a1f0e2ff631090b85b
z75d56568c5fcc1e583cdf07797dec704b5f2a6ee1097c3a1e9123880a433542e61cceac068b326
z7c1e4530244dd9ca140447da043a36c971fd06fca67469ed28dc0f1b7f1d6a92852f79c302f9d4
zadade332d526dc7c5006219ca724e236b35503d227dd00c0affbd2eee47777d9a35f021126ef4f
z35b3ebf4966c9164731a0b9407653a9279779dd5a4d9dff145fb3a660c465638d3a2310390e16b
zd892a7d8c5fe5df3540a8fb7df65586a08f9026eddcb3b008e712d08e52217d8b907ee30cb5316
z38b24bfef1f46ed99a31e601e5cfaa34c36f5da83020bf7492613cb07442a48cdb4c2eeeb1b3db
zffa3728e0b54f527904d417df131b3c584c732d8fa293b4c3625674a92f1b0f0ca977916660d0b
z9b05db48563e17215f4c2feef5988b8d282cc15945f6fd15376e2aab1962b6aeb4bd63bb185373
za0ccb000e0ae404cff6588e09c36f3d39ecab9e7ec1bfe4e595a314c1a891a217280fc15c81cc8
z4b6196b350de7a6e3d55ae14a716172115439dee824c64df7a440f1d22469b6d20bbb44eaf63fe
z474eddbc64a43f4e73498be0eaed2a37acd74d39c63b6017d0944a30d62b8c80414b8aa9b9dd89
z08e284d2108e94f6ba8b08b827ae508240a1a8eca9f4c96a34d4128209e3ca50612e594ad0e007
z8556f24a8a7118422073387fbd8901fd6cf0af5fea3f3a7d5fef7802541f11a69f5fdab7c2c4a2
z420bab103ec80a265334b6166668845ba6d0c04823a4f84c53f9b555598c685521fb7eaaca4baf
z41dfe418e51c7b7506d04a9d1f61b9ffa589652869fcb5e0a250e59d343c0689433f9f599e4a7e
zd30324705ae84777900e95a61487aa8c4d4cfea3c62d9ce6d385aac25ace44a59ab68747e08f80
ze39d62eb89899c37d32384b1a9aa87b55622d3109e6be16e03de241e875162ca4647798e6f2f78
z4ed6693591e4f6401eea9dcb6357aef2438b67b9f7b357ebc6134c4a0f0689025cc0e5c6c59364
z8af2fc50722f50fb7a3defdf7ec0b11f46d4ca5f3ffffeac144795362d72333ad1690ad28c2505
z86fec7cfad8cfcef16470db4237b1318e734102fdf5e7cea2c8ceba74fbdfdac9a6ac1e8d5b13c
z47e77de62b35b9a201f5d5d8377c34fc1d2aafaf8afd051e451bb8112ebe7509967f8c5329457b
zfc4c6f5032181662277aaea249f27bd57809c3ec1ec30ccc5abb2fec99cff1a306e85846fdcf32
ze7c85f7a1bd5a0ee87d21215226fcde871537d9a4633c042d9d6e05c883c8a5680cc53ba7d358e
zfeb0962a6a65085c54a46cdef2ababd3a126e37c5199693ae17cd5223d67e761d6d6cb03272fa5
ze2263b6c83102b06ded5658bb37f3010e41388aa165566181d1c6251975cb1e92818ea9bd918d5
zaf7dc3e0e6c244198500a7b361d040fa4966258d3f7192a19ab31c2393eaf787e7e0c87c65db50
zc2cfc498ca054cae772a22ae5c44c32c319a30e446c1a68f279c9b27ffe85ec796aebf3a62f9af
z019b47e7698e90630451cdefd5dbd0243e073285ef02bdf49f197d2b0771d736af8e14543e926e
z35f16702918d1b3398c73641cdb262ee5bac4f92abecea0691f3f815da401ccdfe5eb2ca3ee29c
zfee6de6f9426b06e377585099e70639f2ffb9d408de7a03ffaafb233c4aa4f1283ddf73a997bde
z616d8bc9b4da6564441790916f93f69dc1505e1fc57749bb2dd8dfb60b78387e562589d036cf3c
z338890bf8aa7f2032e125c0e8c913dc76014de79ad4f22edfc7c76ebbe47612573842abbd81bd5
z1e436e6b332be2088bb1ab87caec3b1ec7c6a1ea351677709f5c90e39dfeede017a31dd6739b1e
zd2700cef4545ca4697a4b1167fb43e6c268e761a97f577862d68abe5250b62f75fbc290efd0120
za6b7f1e543c25bb76a6f1c13de7a1727fcbe80c3971ea4f222036c71362f49220ba08a79a55f25
z88c7b86327c4525a6950c1f6ae985562946e60f5eef739051619e41225e5b847006382f679c4cb
zdb66f1205de49b5ef743166a61dec1d0e3a77a571929cbfa380c16c3f130b9f3e8245feed6e7db
z3b616b1c48c2adf59c2067141ffce13ae050c500f9c3ddfc0678639bf0f02ef973ceb1845205c4
z62026d91548bae96c822aac24e62e712fd18d01f4725b9e0e1264aed43ec664b883a7a4747afa8
z40d611d7c6862ad1e159ef85e474c12ea1a0b67e54534a2c515bd1ced4953a640fa363dce23dc3
z5ef69efdf571b5eb6e1341863e99636b3c3e46e8083d4596f10c5c376354727b46f14982f0aa66
z79c3d41b9a7db485d979b885f4a3dcbbc354c8774f15be92b67f85b266c6fa4c18e0da35abebd7
z2541d8b37c4fa825682fd9b981a9ab0a1b12d06a972866108e46b6e9b3091b7a42181c010e950e
z2b76f726135339a0320871bd887278701df3df585aa14afc84f5c0c733e7284da0171f9c9b6349
z80087cb32aa31e58208221369f25fcd9d394dc274900d7db46fdb16f4f22af858ddf0c6a887ccc
ze3685f87f78bda721feb9cb1782924e1d87c102945157c413a5ff3bf08865bed8612b2c17109b3
z6fe2767d4755016d972ed82c67c5831a9c7dad013fd3a059699ef70f9896e88b36dcf19b80f6dd
zec18c64b80f1040974c0b0ebd301c0f04f2d9a6dd58c3760225a1615d76898a0378651aa36e5df
z618fbff250deeda3a178cc498c2755b7fd873177cbfef0ad6423d2c1209c557dd2e000e446693f
zb3875880a69807fa33a2b3d9be6fbff2b540c72879e1db961ee9b5e2d98dec687bcc06bae23299
z8e2912d04352a29e8a11e7fa22f6bf1265dbf1a596fd19ea449fdf92f1d6de68fa92acd5226371
z9a5d2738565754957cb89985aa2c05d7ef5d3b97c66c5383a42d47ff86e264b20561cbe175e0fb
zd0c5e391582ae6ee07c819db99ec5219b6f65958315ba1c3733b8dfdc4266f351a245845426658
z2c69cafb134167eee0ca1a0aab8edf0cb7edb3640748575d97325224add093c9a1898f34462754
z095d44acef5c0b01b1613a1d17a2ba8b652a12dc7d58ba77628f2d050f1f0da01fef8665d9fe93
z637f426a7638bfb6e427d303376116ee633658058deac4310241a5efc7a47b96544e1ee1ee8ea6
zd707fee7457c66d38b8794c9990a850f2c9ec407085e9460a0c1d0e7f55c216d5ae481dabdaa52
z69b1cbbe3733d0c392e6f6eb5555eac354bf14b0529e18c420dcb19b8d39cb7c000fd195601237
zd56ef7aba4b5b50d24715325743dfad3e4bb9001acb015cecb041e2c64518ed546d0d92d3cbfa4
z6e8e02aebc0a40c3db7be695e1719baa410ab9fe84c3628049c96089e715f88dea2cdfb3dd53c7
z67e014c31117afe3e441aeb58c59460fd1f2b9c0b019db85c6a3093465fca307ee8556ad3a20cb
ze35c7e1ee04dd8c6624b00b333ec3cf93ed319bcde7ee028a02774f1aeb62945c15ad11e4a454b
z258ae8a4e37892ccee48e3a41d0d13da7344b0653bc278c2c53ba24e27bd178e3e7f0cf07bf756
z17c8ada9e204374c76fbd0db0441b763ff230580154f08ed5dd9a707906b29f2ace76fb85af19e
zaf2dd39d5447e5e6d1dc7e5a71c2ba8a4cd8f4f263e855c7dbe24f8e5ff358308faf97a558d2cb
z386cc386ce7c65e37d043af88d4c6b2ff521bc8ac524aac52c6c9fcbc8b3616034221f2cbb7a1f
z9c41c3aee2d1c8021ca1ef7191df0eba32e07b2add1a7fe655ea3b6a2e3c3ec9d537ed1eadeee4
z91ed7b554346cda2b7ef8baa42fc6e0f54fb93d3e11dbefd572a7306a9a9843a79d955874f301e
z5cba5afc12fcae8e09a369e068b436f9322ab937cabac21d09a163ab3361bce70fe023203868b8
z4abc0a4e031383c5872401e2340cd0fd848032eea31d74864e13dd8e52c090a4eb94ac6a954f27
z294d4f036c25fbe8e8915cdf74ff016fce8778faf3bbca3728ed558bd7c0d76a8337addc9661d7
za8973a30622a5de3ed2197f1c2743026d8a3cfbd8b5e58810ba46581ca9530834cb92df7ce9acb
zf2662fbeb9b4b9e58365999afa27ba910e688bab6906eba52a1e36613cfeb091481e51fb97c34c
zb3149414c2b6f6d2d6537d8256cbc1332ced12a787048a7ca6c7be7ad96b5086667d871feb34c2
z5f1e1df37d962624121f43974fa4439ff4447c8dd9fa87b8a975923ca298284f423a853052b437
z26876846aa084bb0ea8455bdbb381a5597c45d59a30c815ebf15eb82af8116b7c8d1f084ed5286
zaba64954b1702a11c7685fb1af42a72155e5a8ef1654ea3133e4bf9a2c56ab044a870e3d8916ec
zf0574280ead04c1c3a9b88e3483c14018b43685580a4dbfcc363942c2013cdaa896500ceb463d5
z0349f4138bcc216647d4a60dfa2f9a2bea2bb4e793c8561abade0304fd76efe21f2c5e32b3f488
z230fb44e1688696b7c554a266821ac0ada6d5886d59769e6a7de1a5b491bd76ea64386b53be42d
zca61a88a62dc0b08f0cd1c348f0b614cb496e4faf98f44ba3028d184705f9089a0cf8a86490d75
z20571599b35af34710c9505f357409bd2465f2aa9fab6d0a2af0b9f03bd93ce2081330d6ae90d5
z39c4d2c24318d6d02c89fe8caa1cf698d446e7e8d34c98f84de3faf18d57fe2d6f967d74b2df50
zcadea86a114ffa57f0bba9fca024cd8b0502ed0860442524406d785bf74844924bf4e43e47e0e0
zba56cf77217e3eddcb5e25df31e93f5a67b7a702b7ac5f0e93df98c81971e98b40b21496296298
z5b98c211b0399275971d05697a47b1c7c20e01b042f40abd7681df4cbc6d6389b26e6f12fde158
z4240117e3667b252c1ff078334547ee9fc77ce87d1f32f003b05adf3d9e13606489930b5d9634d
za2309c2a5fa071866fb64866a9cf4fcd25a5253c716f1ece4c1392c57df133cbe2611a61e0cef1
z9a338e209ded8e13b79409add951fa6d5837cf3fee04e9bc6937a0778b14185cff6ba7b473671c
z9ca52a24db67010b8c4eb2c87990c966fad41bc17aee3c072724043915828f66e0cd53440b54ad
z16da4e755f5c78cf4f38952c142e09083e6355382d926569b8a57a7cf073196652dcdc8dcbe164
z4a5527716dc27f52451b9bc9ddab75cb4984a9504bc8c2ac6ff184573003495c15c70d46d4eec5
zf5f43a6a3a4c7de09b6b41b0bff27b2917668cca6450c966a3e7c9901765f82610721ea215a0e7
zf7beecb8e2caaba44fd5c929efde46741e77c796b380fe5eb06c3d5df135b1356e96cfebd8c73c
z34a2b66fcf4cab698a44acc639a7622b1039b9f606c13a1571ce94ba39786a5295550bd555902e
z282e951c0bcee10e8dda05dd094c8a3be781121df5d21bae8041bb5f1229b45ec46265763c8a21
zfd467c9625535a9c1ced8ffa42cef8ffe1d33022f35bb2650c48b1213545eb79479d5bb9265a9c
zd52ded6a6bc43964f1d94e12dfbd3d67d878317a7ead0f74ea24a9e36f7e5d4ade4fcc7c6d0778
z7580a3adac9b6c9e5af20481889534b01b0f872ed74547ab58e4eb74b4710bb75a5caf3e8b21bf
z392e4e20bbec7cc238e7871f5300adb936b12a712249089fd8410f3929cd8b003673d1e9c9d67e
z0438b4584199a571c760254ab54ad6d0a4a7094a70483306e8cdf735cbf2180ae821ce2ffceeb3
z681c902aa40af4580121fc7808316fbbbe1e6d36157abccf64a0c37e25fbf6dfe888f6cc9a4ed4
zccd64d126aa47017f0a86f07728954ad36fd5ce9fa8757ae09bb12aedad196617e251f39b2c7ed
zfc60b808375debba9081f50c574c80c338a66dfa182017a8de50d7b239b1e836c8fc39dcd7d22e
z9212d294438a9680f43d13b3258f85ff6878736516a96fcc3856b1df2c99b7da9c821939a4ccbe
z158bb0a5f863ff4ce3f7fa242a6d607f1e8a5421009b955b956123c9f3c73e6f8a86ab4e02ca3a
z75e472a44db83bab06438ddf0b0e45871c745c4ff2378fea0a39ff56674ef32da50dc43f0e3fc1
z6faf309e9e057f78b655e285b17274a3c3b33f3bd495599fb06d363ecf435edd3e961d9d6155ee
zcbbdd9dc5c05672034965722c0af727158a1d24dbc1555324c68b8ac8144ec17e752d5191c14c7
zb580694075455da9a2221e17953528c1b4a78449c370f6c224c991364fcea7fa48c1fdefa102a5
zb97d2f8aa82f1d45614e96f1f62a53044872563a98f8620dfd856399db0ec802a2551ae532e46c
zb6f4eadfa8cfbfaf763197e3e25fda3b7ee21204f14a39875d68ebee5546140135eea4a61284c8
zfa5fb8c3bcd9497204eb65b55431101766f620950b57dbb332dd4eb83a9522fc6d1e756df8b721
zbf90c6f144d83476e554254d559fed36e554757066d26894b1d6a346b3bb4431f433a97d3e1534
zc89952a8c247e89117d1155a8685361b91bbf988756e18aa079423edd0565c5fcb59704784f358
z4d0bb8ce97ab322d461cd0332c42a31237f9bca8efe4890656ffef4bae6ffee956907a53d2e17d
z71f563906721d469733ed64c02b65c28dfc98857ef440cbf0d7efa3a0b226e56176e19f02a568f
zfcce8d8510648916a58c4e5ff8818756f3c23edd0d31995952f17ab465191d0ef25f091a7df7ae
za1f579f967331a94300e9978c3c48510064667cb7f28fe884a36194727115d5c86625be19bf8d4
z4d5919f4f2a75e1472c103336fdbc5ef7259632a3bc35274dc7239765f871f876299113de79088
zc53d9b2a3a428051fae9f29b822bd79776d830e4d7c911d3124e1f7705f00de3080929998f60e3
z4222f4136e583868bc69a9819f0018b799caeab753efaf13fc75aa9cf156e0d2f6bd8377a6a4ff
z66eec25bcc0752595bcc1f2fc757faf6058009a7f6ad155ab0404f37c117e3d0a1325979a76225
z52ec4c93f6882ed02c4a1e4acccfc7f73a707ee96a85d7c5f5a4d290017b8757748bacf7e42a5b
z00af7cb391928ccb83e967f917a8fcf470e980f85e056c4461834714fdcef19aa9b71351c3744f
zc87fe1ad0f1b45d6ec1a867f40bec8ccc9723cfd9c528e9bebe6614782c595b5798a64a075199e
z3d4c96756341703febe0f6fb672a680e2616ef200fd64fcb1f0cb5f0fd7d31498323164fe8c936
zd0d5627be31c1325bb9bbd4c96e72acc48f3fd7bdc4fbc78ae57d4ed89f983aba6d218f004f3f6
z4390ff0906344657838789b386374a8c2720d9c16c27c2ea2a8ea68534f5bd1227455e94f4ae5f
z03e2a07ba6e78e399e4b7dbeeff38c78696624e01913117562bf4b1a5fb31dc80b0f4ad7505bf9
z5ed47ea10691c23c9d67c5056215c54cd461624b03bba3c37482b9e6554359609e2f012ab7d3d8
z35ca8f2c91998ed2052bb598a3d28cee045831738da73bb22155ce78c7f842bf170ab2740244a4
zbc7a5b337c18d7f9aa0fa7f760959334de98de7c102872c63dd88c6948e639726904aa23f85c69
zd98f2ce4e1cbe0f298664ec3b313dc61c143622ba2725ed34e1b31a55e69acf7f395c7f42756c6
z96f482f6946def262b2d69a31d94b8e5d165be8611dc60e9f298d330b84549fd142b1fa88ea5b9
z79a39014bfbfb0aca0df822b926e913e4b2b617e7656d0117523f9976e78b9d9738c67552f34bd
z2f2badb55cea7f54a42f22e5d64515ecabf0904948bd3d33d60d48d3d31a24456f900916e43cdc
ze5ce6ff24d49d951e59049bc57444fb7e268f4413a52182162cc771c49c40bf787c24b6ceebd51
zca1fd2cd80c6bb2c4b5c78939bc1379f2f83be6f631b01711677cd1e05e1beb1a5a77b599ec9e0
zf25ac203dd92635fb7ddf452668c767978b68f8a1f5e13a828504f8f32290ce5b4f3086a4f1ce7
z8859fca633ccd1b412f48c42546c84a4b601c6810ea0926936baf03bf88eded5410cceb78d4269
z87e68073b0670ce12326fe855cfa670b0c753eb2ad747027432034d6ec76e2af7e9762d2cd3472
z0e333d7d0e3f87e5805190ef7a406583fc0a3eec6a36e13d59fc915aa53843a6c3cf7eaddde172
zf76f773a1753b85e6730474a57f571f1672e71cb82b9a6ef731e990e2c46a5aab21dd1d0975895
zc4614738490143e038e9a378d4dd00cdf51bcce7db9ca089194f1816b57dafec000580e14059e7
za40acd49a6c16812c99419c4c83e3cb53196da1e722fe71896eec52ac4e6f72d750c2558c361ec
zdd9025771b49981e62459e0041d1911ed0cfde3bed67b2f03992c9cd3b2941c36dee87d0709f71
z6edccebd4f855420ce1d8d5eb3e9b28258847afcb99d2f521021bc7b5649032bd29058da098320
z1c72e466397087ec40d2c90a71e6df65b00f54731ad201786ec72d53da5d5bcbd34238a9ba4cc3
z6ef225dc3656e234d25551916b296b13aefbdaec7246d22a6b16f2466b45a331f6d10f42d68ff5
z63f85aa2482562744a436cfbf7ba06896c2841cf775495d9693ec998b6700d777be7598914f32e
z191f68472d7e03637e3c80151793a21712f3019787de34b1a2ae351942fefbf30d430f8dfb3a32
z3e67f8a1de0e32a8a4c552ea650914902148e376a5c006e5ab3013ba127b8174cc0cdd40139967
zf08decac49d0c4cb414f4a0cf48b1236a02412dbfaf54f9801280a48e8b56cfdc2ccec40c99a22
zafc287541d1dbdddbc15247c2f11af66f928218f262c7d964804c3747d54004fe5a4cd188d0411
zdfeeb0374f9a04c54e369cd932a42ce84782a3d882e9a32773573908bafac0013a61b02c498c80
z7c964df4a4c0f7ba64f1574368dd0f51689d0176b15dc37754cb0046f7fb8a684bc2dd143ce03c
zece492bff7d5ec83d6ae1d69763d97205c0e0d1e5f3f43fbd5630572bf907d7217972cfc5baca6
z16887be6bd6cf332feb995d4ab94b58b94aa857223e39eeb62c2c1d6a62502cf7d5e20f89075ab
z22d92393516212ccb03f0cc3362415d55c13fabf35391f63f8551a231356057913ffdc21c75fd3
z36493ca77848cfddce7873fb8163a7012357d67745c90c8dd9ef523111eb6c8688854ce18431b7
z2528a8bb69a09c1ea14a353b0152143ea41feb9f21db227c45b765ece641813f4e13a3eca9dffc
z5a0cc359937ec9966a82146d9cc01b8adbeddd9cca4cf7863327ed904bdfbb4449d8da1bb65474
zc8c7e3617adda59c39fd339628d1f23158b25381775128681ac0b3e19932b7fa3b12e4221c5d89
zad7429b03e792e66efd71a37b822c3c3a4fda20cf412c945b8b400522440e0f3dfd3b15967004a
z1b03d0ccb585c510873becc78ebeb7178643477f2995e04e8e02a632ba32f62e8ab1d92ac0d13a
zc748b55077e0baa5b8032b08b9d6a246cb79aa4008b264fc4cd6588f5690f1738f753df54e37e5
z22135588a86773b272b5cc67d7164c7e2d4da8358b758f0a38f251570cf1dd160d295f86d1f387
z3845302de738d20281a483316040d08a2ec97e503e55e66eb4d4230f2aa8b0afcb4f0243a7bb97
z21e0b870a07a810ec4b8eb96139660660bbd711fa1a54d9a0e646f66e94524626c8e8a0d45377f
z48806cd2937bea5f2498b5587f5345a7dce5f31b5e124a36dfb770cc069c4f41888f3cfcc83ceb
z54f36bc601e0174503cb60b644a67cc0334386a0439e490c174d8519c345e9595f003169ddace3
z787ffdbd7e75768a187bd4ec2cfd074e9a8824a751c16174e46daa7c044a3fd93adbc21a0c1686
zeb75a798593dec62d4e89231c61af1db0af1a14dde5f9c9f89abade70dad7d5f025922999a2823
z20fed96d7bb6bc8c2e7a6a0ed0ef677c65b954a005433f204c9251c7a7b9783e796f64ceb1dfe8
z78a5a19f9115616e9711463897065ce3d4d19c88447f9ec8b448c4f6a0c9b7896c4fea863bff3e
z4b11eeb4bad3e49b8e16628e24de5f0e33fd9be79c1e790018d9515438812826ee9abc7c850993
z3b2b73f3702ed134fae06b1b7dc32872a67326b6d142f176ff7bac97b07a7fee31e58b5096f7c2
zc75f48988c140f58fa7b9aff65378f73b18207bb492b0603157f7012ab68b82bbf320af1a6e883
zf05c4df63d2de7b7d7fe6236f61abc724aec6603c349dc22df7ac40ae0b39762c888c229ac87c0
zc4c4f90e3108d65273aaab6b1f59b59b4cb95d9fa91cb8f1dd1f18d8ffec0f4ee808aeb5a9d57d
z681f855d093cbbcf1e731925287d9aa9242067a27cca7cf02e0ad95337d93cda5517485bbd25d9
z31ec66a0cfe49647d39e4035dfcad2401e0ca468108e7347dbe3ff007d877a59e848d357e5b00c
z66b33bf61d9e66dcce885dfbd5c86cc69373d6afc683e827ec9cbcbc369c99860eee8006ec1659
z01d31b1bfc74d342259595742028695ad8ff5271020fcae895be75e229820b4957ff96dd933eb8
z6f37e711e3d98df52280ded3dc2f9bc04328fb3f9df97555a8b959b7a52a935f79a3f9000b350a
z9a1e1ba0a6eb250b03641a88e44a9b27cd969259de8a13e195e80c9439ec0dd1330156d74fbeba
zbab0f9621210aec3e4fc2d6b78a0172a16ac7accf9b572832cd491448881fdf71080959aeb7942
zae26759a216cc3a0baf40d42fcd040035a7b0d94b77d173dc970dafa1136d352566582231af2ff
z2d09873b15638b3dd2e44bbf43a822e93e79afd3a32c94101f507b9e8e67001e276407d2b04f17
z7b91181864f7b7cd6147dae69035720e741f26bb9e3b872fc35772fc8c72ffa03d87ea0845e9a7
zba6e400c0558c786256c7656a7a53f5f427ed3e473121f8fabead0f362c041b9b4cda53d9e01a3
zf9f47d66932babf6287a5d0145d7d547e375b306f22fee09b0874b3561ed9875df2a77715db68a
ze3d85099b89f0ae1492f73fe9b5679f2cd9fea5db32501352121c3dd5c6135225f2e2d275512a7
z62e821393d38e76742c3258f261d8974a8db6c45e449664df79a03c8d680ca44039d3cc2cdade8
z1e64e6ef22efeccc32dcdaab80d27eeac3cbd8250a11cd73421f9817c6ac04c7b4a6a0675042d2
zc83a274370e91a2d832ee307244dedf4f89710bb13b96d6313f8c051c4d4cde7cc87f8fe543d44
ze1f26d161b53daddb4c747b6db138a29c7cc4a3d8a5d9751d1a99aa7daa859efad7d96163f7462
z7a18e662e67847b23d79f88faa52995927ac27f495af92bb43ef25d5b699938c0a1a5334c56531
z2828ddffb0676ef14d55e9b58b22e309052e77ae6fb42d377b8966864accb8fd63d2e48024a5a5
z319b460b8c4222993b1191fb2f443e0b887d4f7a67b24b4c80e2a128470cc79353f25214859de8
ze9c0f9b4a0474d2de4ea8a522def69fb18732b9e4590eace30c9aa10f6ca27902a96e7276a4c6c
zcedbd4a7d29a01c0c904f0566a8373884ddad8ebafee6dfa9a348dff949bab4799600649a1e9cb
ze68735a3d9d122ec6dfe6e1e7318f8c3dc9b2ec552089dade401faf1d389910513f89a4ba57872
z0a93d1c55dba49d32b17ed6b77cd6d64fee6b9ed0db293fbb7533e76f492002fb161e0e896c03d
z5a0978d04ea448526373dd2aba16f4543e8481ec831bd93b5a5cf7536f2b65b7fea6c238a23ce6
z6ef0e29100901c4952aff9df8919dfc12a384fc2ff1b7c411d5fe10612eca4a2de48910081982e
za0f36bc8aa47aeffe47f79e5c07ae6fd9438cb18a05826d7d82b02a94c3a023f4477e55819e07d
ze5c8298c9bdda03c826a6483500c4862db48c0d6f4cf4d8abf607d768c07749a8bf082cbab52b1
za3ce1450ccb7d7b29ee6bab4a089e72cec2215efb2fc26af5f15d4c72e4e52bb8c98a9fbd270d4
z3aec32bde329dbddf0b70eb07501ecd560f09994306be82328b53c59faf55c4c69c094b8d26af7
z0cfc31ed7d741b8e32ccafe4018df346e592d3de3ef0835272e992ff40b66e1cb01ec1d8e3fc24
zd52315725dc273d0967ed90135b5d9bac6128068eeaa1ff73adf52bf3c68ad675063c3d97c1461
z27cb026994b1da5bcc83495688fc667c5a13bc1a14dee8a827376787977eba6fc005e960b7aaaf
zf124ada68891f19b46f44c22ce0c6645b5ca6fc4ca6117dd5b0bc82d86eb9fe280ebca571b2884
zd318ee84ea82da9a9ed4b68f8cef606079f066a26296ab6b0b3ddf7c931cefdf21736fe0a49f01
zb65e202c9325bb51350a0554f72959cbb31b93f246b3e44366b804b4ddd281658c638e17a33086
z5ffd3cfcc922bef5ab7c0dbd1010745cc7a6bdee40e51bdb3526deedb77c2fc5af663cfef317a5
z0b4826be6b33ff06629058c1e9d11f62d6ee8f5dcb4f98ecb47f1a2b30c94247ef56ca2a841bf6
z4d9b4c2455b28b5059528f919cbd6003c62b29770bc83455d279ca3d675c4c75f3fe75a28d431b
zdb3770ce9a50e01daa05e022a48646dd307d42550927df93b1aa86d24669a8cab0f1e7bf951612
z30019b1a1dbd5fea8502bbfc3a8ec622b61691bd9ea028f544224dc24200cdeb1d7c65c15c5204
z95e4021883ce16c7d3d66558f4a167c5976eacd352a79d68de48d9a74b85df7423459d26c84e16
zc5443a4daf4a6647e3d825777e7b7a6dd65ea0f4638c3dd0b47bea401ee574d86aefc0d3683345
z7e9414a864b8119ee3dc0e7048abff84e7c0cd3178eea3a46cc958fc06a36033070c823c1c7524
z3dc404c3445e51eed1ed8edd570dbe48fec3021ffd746687d540fed840bcf201793eb33e67b653
z0d3f8ad6f94ea44e83eb08fa2a5e1bab8be3df4f19c0ad8dffdfd6513a3088e444500be02bac9a
zb1bcdbfddc669ff677d4fc5869015198b79936cb7ab01899035b0dd81a83bf07ab2eaf31e8053c
z02aa90ad2d20afc0c975f645f6736d6bac47d49ba077011012ac1321d7c6acc0f6980ced16e04c
z32dca6f46a2689a73cf59d92be97c75138bbf40282e14c40c1140c3899673a2d950b0e00491a8c
za718f6375e67f59e87c328a0ab4bd72385357eae634a5bb539b09232295b147bb415300cb9eac0
z03c1ecfb3f7b9d721413a2d5c148b5d3471f880570bd4b343a6abc789d94f88bbf0aea596c2774
z60b923f36682c8b5f1e8ad08654ff9f5e47726628b8c2e74cbf8468557fad8c8191ee74b76dab6
z2f0a98fb27aa6b699514d7bd2e26118de512f7783b06b2cfd5029252382f14f18f59866c179ec6
z54515dff73cd4ab425abec408052bb7ac79ea495ede56e630d18d3db6528bdb84d94a92a7e8a08
ze16f687a8dbd4ea4d9c6af35e13b562d00bc91e84873184a842c1b029d0bdc1b6cd300d470e44f
zf3b0cb8310a94edf087ede242671ad0f7947e11c645adc73b19e00d7f74c3911ee941249d37eeb
z14a1b327b798aa2b4a466a978518c495864126f77ce8a4e6ccce6f8e30fb026926ee50fdfe9c47
z7e2bb23db17040353f4d3e0c8f53d87090400ef91028d47f78d71a60d7c48191c56623dea771d1
zd916c4d5e1a0fce3b364614599fc85f139e21732e08042cc5c9897aeefc2e0fc41aa54e0cc7d03
zf4de4fea748ad986033dbe28ed27e538f9ade6ead394cb1faf6ef3334ff1ce8ba47bd66fb96834
zbd7031c7913f01ddc53e19f3a23acd44c914f817fe03c58e14df6398ab45618aa565f3b52da97c
zc2682eb50fb02664a6a3cb93dc805a19bd77c350cfc23e8d20738b5f1a0c73f4b0c7661833fd7a
z07e2125e38bfcae73788adc6acfd95658a6bd957b3973926a8b91985ca72204803c472da2cb637
z3f51fbb20e6bd9229330305eeb4b9bc47b0e2be939318f6b137dce7fb57fc6247289d70a9a00be
z651f405a3a6ddfba6da2944d3466cf05607ed3c6c0b629b583727a9e775a710c3835b19e3a72f0
z1db18d5d0b423b9aacb829b3ad7585685d8a5cd128c440dc6b8ec591b2e2fbf9c659cc17558bc9
z4d9de18184585a71b93a718aba0ca257c281e642005e06827cc68b7097951e79d739619a9d45fe
zf11b5477095f4dd6b0071b207e04b73b289693eb820a32ab8b3cdd98f43dc5784dcb00af74e0dc
z9781bcfc8c8658d53bfdfb2a914d603a1845e809b96735b24912ba5a530a88f10f409a439b7495
z32897955c49752b094721f6ec7cbd1262d798aff3e13334cf4077a42dd3c934a0daf24e4be01ea
z0871138ef5fa449b30a0f25c215ce8ca9bc7830bc3c21fc37ede6fb2b07ce06101b58d8179117a
zdeeeeffe5ef8ca56f5d14925606c30eb3df08d8e76c896e8220d36a524cb24a3be878de5069983
zefb4fa4bcdf6f98634d5e9fd2cab06575c4380f69723360611d5e4252720f8949e4a1c0bb71487
zbf43bf2c52f878e14ddd898f5bbc88c637c747c69bfefd8f7026ad983819c67e8a0613fcd90f07
zdbd4213991cb51546f31613ea86d341398d8909fdde7cade2573c7ebc363fe715c040f2256246d
zc7e831b0286ef0b87c153fb95a29d13fbdd4655d61eb0b00dd00c1f8dd0e6115670003adcaa513
zc4faa93ffc899daf5401a470232a2ed3c8b30fcd8143190a75cb67895c21f2600161cb68549fbc
zead58aeaa02d4cc0aaab80cc44cdb519cf2c62773235bb8c2ec4d5d46bcc3e4864f02c9553efed
z3b12ddb877ff9357b956fe2ea48129e9606660566f587c6eab7b7ee48a0a088c098767d54e7412
z700c445a18d4fc813a51a5765c4e6aaa55af5977484dd3f0f575b7738d27bdeb75b737c1768924
zceedb9d6550ffc58badbd4551c94dd29f55d9f9e4d73a37c9e8ca5e29e53f8c14efe165c12af8e
za49b492d8f15997d1b46c248a4c0197b0b2634f51a941a89d590bdd19b8527f430fde410783999
zcc22999a76c650b2d66a1a6230daac671eae5323cdc52919efeb3b2c4cf63dfe32eb9a926c4f28
z67727775238992c17b41cd67d564aafa222a08c902bde1cd489225a013f11f37a46966c6f74532
z325a26c4a1113b507c5ee9d39894c7ae4937af80efc913201c29c1766b7e28037b3334b93d345d
z1990112d77259416ab42147ebe1016c4afea59ac6cfc7e8834c1db07544e04920a7e65fa021cd4
zf5be79b40d286e3ac6d37d7c34f10acb8c52036846bb6aa67f537ab3165e8a2c5d2c8fdeab2962
z57a69cf0360eca233325f2d6535731dd03b0da6234e6d0552c63834528105252d242fd4cbff06f
z1645cba16d84397b499ffeee4dcc2bb1f40c3a620636447adf7b14a35519a8298eb47d03864c53
z6c0ba8ede85e9652ea3252e72a6dc873a6181039130cbd52904fcf1a2cc3a4e31c7b656960efa0
zf0733786a4e740d1e9f4732a8b2f475ca05236be1e9a84c2efd835912bf6b17fec4f761f7e9d0d
z34708c873556bf7e5f82658640ff8440220909a61d6d44f0d022b308f85b660979a08134291a38
z8144342c4039da2b8645626c5f48dc4e559e4cf0902f7d0f98e606f269ecfd1a32f3238f516a34
z98543fa5e8c07e48cb4ddad6ed399307c41d7b5699c3badcdd215b321f25440b5828eac6557df1
z0c6e2b8c78e8bc6078a3d22a51c4431b9877c88131fcf78405c39a9aae0be1eef7c51b8397d420
z861c96667456b56348ab0c7c626f3eee0b470ab97233384848b322e985c551e19eb951013c93c0
z6e30943735d042a17bf9a6c2e61c2f4f41bfa7da920d9a3e2b7828f46f1bad0a90d1a413ddf284
z6d1a2da4aae2436620e0f046129f85e6fc1438f7435a9bcef390821f82acfabca6c6380f1fd3a3
zd7938f9afa013ff8a1bb1b8a37aa8e69b7e4ebe4e2da205e1d9c1e3bb0ab8cc51924c1541f6c2d
za21aeaf3e5ad23cf5c7d62cc3d411bc74eb2139a3d8a21993cdd66ffaef42ced0de8a37b884da5
zb72a1335067ca2df7868cfafe2d3515aa0456c3c010ed6eba3f979928749fffcdcfd5d752b36e5
z23d8ebc24971dcf0ea05a7b83ac98d0b49e55a70731452e05380c75672192566e7af75af7d1e3c
zcba3e9df6d2747f122b96eaf6dad2518a5aad3c9a5287f5236f08ed7297f1cc6f0c21ee292fc0f
zb871ca17b235a4c927624b9585f6f60d0b91c69ae00b98f406163f563eb13a1b5f7873eb516526
za48cac517ebea54ffe3f29979e371e2136c0b2311b9c0ab584e2fad15be2e673ee005ebd24faf8
z80c65ab9696641f3eba3fa96938dbde53b6bb54876c3809324674b519a9599806b0cfdf56b4cdc
zf297d818725ffdd930a8cc1903ee1be2c62624754a198ecdf35aa138ff90e21fac6ef3246c99f9
z97aa77340a58f6eed75677a84bbb2e4a8ba5aeb785466fad3d33e79c37592c5eda424ea5458ea1
zdbcf27a88541dde8c924317a2a1b3b11884e6a8eaf95e93b3b11f042b6919ab7e8d36e14634cca
z76cc6275148232571264ca1f82fc505a0d1f227c6e7ddd1622ca8abbc9cb084732750a34ac3499
zbce7390ffa79983980245b1e2624a9c89f16314c6a2a5ac9415cb80bcff95a812a967bcfd49a15
z52752b8cb544f7347e3047d4d7c5c982ffd520d02b5e37abbc94ad09d7b2c527576b88c9be7a76
zfcc9fb6115fac34ad98751d284490b9594d2321f8c67fb7395c970d0e1cc89dbfc3ffba76ae961
zdba7739865138ee6d953e66d2dac1aeeda19c9772b71d9ab74c9859b7d0b8a64009bb178fde885
zfdb704c128dbac5e4719d7b0e371b5e4199b09300e25e2eb0a442c6be348e71184d92f5b7d4f9a
z501f445a9db2a5ebe84a4b9b8eae0306fca6fee08f91857e87e180653091669d1e085a80140c5e
zbf780ee935c5f6e5e969f8e4019e25a8823a1432f3e81a55874a5c71d2fb0124549e502237df64
zcb01141e73274c8a5b7173c1ebb8b588b98ad14b2e80e830a0853983e79fb7c13ff322271c1790
za84f89ccc0a26ca63bff4884c6e3fe7d0d3ebd9c4538c223d670baadb784eb5693e55f2a731706
z8ca2890c051d76d152b765cc63cd123f856cafe3f24d5c887be9f7b28c629b870258f1bb6c408c
z58d23b3973175674bea334b808d3d370442e846d6851f3575fd526527e10ea76f2f60bf0404ea9
zeb241520ca8137614c4c2c383d7f7746c8b316465e4f631fad2356db65a7817e7801e7b3681ce6
za8a2b82787d3a2fa60feb25cb4a6b3d917385cb48bab3976be786f3607987b4c6f689173faa18f
z00bc2fb87131a7a6625ff1fca3eadb6f36090ec0c315daf1291603490e57d4d371be5b5b806300
z40dedd434d544e456e9d10b1c34628cf452fe32d0787cb1ec100ea4e0e6d1dc63d05f0ed344016
z96cd191d1d8912bce49dcb0fbd16662600135a7c593b061171f819499142ebf23190a526e77500
z22feef346f771c47f2237371895c0ddbc80fda0cd1d0c03726d280d053e39ef32d22fb3ab7e98f
zf7bdf2c6a750269c3bb212b29779bbc3dd82a5e2124c02d67cc8c935c6ffc1529ad6360e9c2484
z0f750d62b6046af18ba94ec90311ca8fdc7aa6bd76c8a275733f018bab04904812ed652930fae2
z4bd7205c0d591eee9ca56a99a3978a1f00019f8cd56e490e4ee2b5987a1c191c42222eaf6074d2
zb5d6d877c7386204f1f52ac8e1436a91c7ed87418c3914b20c88983a5ee2f3d5e8f9bbbb5f1cc4
z9f319177ca6b6ccb0da6d835f695f73cbd4c43a912ec676c703fe813c8e91b394aeadd79d90f6b
zd0baf941b01c3712b59cf2c2ddb668184acdc96784a0b7b3e36a97a0a69abffa755f023983e940
zadd3470d9a79b1a2ea6223e50e5652b1f02462b32e8b6c6c66cf0171dc713f489bf4e0c52470b2
z7c70f5c298f902f7ad246c7fe24e96219eef908c60b508a349fbcfa060a1cea1836b2a8ef4499e
ze4adf7f5248182e06ec9b73ecd60711596df4aaa321a32b2a4152068f0289c0b29b02f67099a93
z53ea3dba1d205d9c0e25bd9cb9c312b54ae2f2209aed46e168b0cd3c25a635647224d80648eeb6
z9490e50d95ebddb9d05b28ac94b2e362e86f35faaa30d4a4f9c1b6b3f747452ce0ef83e0dcad71
z720a11d9844cdfdcb202d215181785a1a9a2b01ab1c2b803b55196142b3fd7602a7f44627f0826
z899430e91e72c2046b37ff9a2f625da2ab0c37a0725a7495ddf35400509d38c85354e1b13376bb
zfacea61b7d67ee353def678f92653051b61fb936e7b29ede29d01fac83ef03284b88db683b3952
z0d9d9c2604b9ef5e218d6eb73ea790406a2d128c689a6538b05aa65595cf69ed8e434b24deff03
z77d4ca13a94f44c0b24b219292fe69c407fb73fa4509a34c66f142e1ec26eaff2000b1df61295f
z686a0c517c209fbd00f20a6cabcef7795d1437212bd822c50879ef698b9f62f484cde3e507ab9c
zcccf07b644e03ac5d62db758ca726b93857ed2d0c1887c2828acc4f9b0e2593be95fd4d11bcaf5
ze5d5d5146e301c043e8aaa7dc883c678e9c4cf4723cd73f3713cf3dba3bfd66cf8b51d130542f3
zcc25c4737df6f76106f71a780117f9599d70e07099ec2316232044bed041e52d0f24afc2859189
zcfdd40c6da68908dde126709a6c6eb3f103ae0f7ff702b11e74c19369049b582dd5ed53aa3f735
ze24c16369685673df399f65d944f5a1b93881b2affcaad2968de194d0c8a1d9491abcc9974817c
za0a91b6739dbc53a2e48da90819d4902fe044b70a824b37dc92d0c66184d2da5f0683d450b82d8
zbe89fa728cac566be1b5b2e8e890c42dd37fa073344b082d1775e8eb9c00b651a0d96c3df02c48
z8cd3ab7548eff251f996e40ead3a2adc7e3cf2e0ee6bf97ba7816e4bb2e88d03de6c7de024d3d6
z63b4ea8593365a689749e0dc2383a96df4b2dcf17733ce7dea5251aebfc68f8e90ff339bef8f14
z7f5ab61720fd1defbb1956a87d82fa0d181415e6beb8dde89e739339d31adce7f7c1a91f6174e7
zb3c3abad1516ba6de6bcad5888b93c6eb73ae8e4c3858a215795ddf5cbb683ecd930f943de8bb7
z84f5423658ba6bbc69598fdb593e1cdb6975cea5b4d0f292994e4cb9da01c70f93449d71005750
za8b9e9c3092c83fefd036fa675c36f40269e167f39ed8301032dbb47441e7efdc7e701526a3d28
zb73ab7092475c29d593b792d546b39ff09c065c2e3f263ba3d73eeeaf416b90f5142867945d126
z0cbe0967c72a1c79e78ff128bf8dd5dade2c9c8abfc3452870d0661e4f3a1c8dd6d38cdf90fa05
z9bb2d916cf00aa6cc429ae1db63bee1cb6194ca75ea3d28eaf5cec80c73f228a6264458b8cdae0
zcfb225c81c191f738d04bfb54564f80f5ead1add35ca92eda3b4d5531e34e613e6f7f51a9aa5ad
z9c556a4672fec839afdc006cb6c1a838417dfc274659e5be708f055aa47f744e32533bc0af9bf8
z7190e97d85d180eac452dfd8cc3a91506b1d79a530ec917bc0182af0314204c62f16444e1f1354
ze1018b64c5075aaf03716571fc0aea7b8ae6864451546c1e305e63d755c9078c587e04566907a6
z43607a3ed176f11bc9eeeb51dfb8ba6996f4b149b46e96bf287b1e59b2e709a94f4b131e89cd39
zb73c28da6ec11a9666af3acc0392752b0d430d5ac0295f97bbea3f5e28ed8c380237d7e5044ffc
z2f06c8dffd821ce678fbedafd6806a8b6e58fc87ed65d35d89ae32179e99ca9acebc7abaf54027
z7602d79aba50752da35eaccdd71abe413b1fa433e387235805620046f08889e7084159e4c40933
z5ff261c3ee0abb29a6991d2554b1eac76a74d2501a4c04dd15bb100ee6886002d9731bd35a05e5
zcbdadee8e2b1d96efd1596f84e2f0a8a11bf5c6962d132ead3dc0992f98e3a8e6366b765a36110
z3c25651013d089f0092599a494dad7c54a4e076070d8327467844095f7b06b6d3e0a67fb4d77b7
z771bd0183e2cfe08f9738a1ff50d72d044b805eb5809fbb36f2cf9409754d946f735d39829ad24
z3c9cfde608b844e2ce33d590f4511bf3ebf953a8cdb8ea0c7811c66c1f569b3fe29bdf465a7045
z1df7e6eca3b19cbd660de2e871b1b59bb6fa9e2f9dcc9b7f18ce21d6de8ad108cb920daed7a56b
ze6ff68ce3b3f729bb4d2e535bad1460895506958ed1560ad525ba9910b5ebdfd46e25ce8c90fe4
z3fd81d4517631d3f7c7fa276c2330847bdecb20851ab24a10ddbe95f225a2bbd73e29fc28230ae
z9bcc80c0f438502916c687c05ed3ec085f027f083febacf5f11543cd2b23ec45d9f61f140bb3c4
zf7cf9cac0a64d6d05fa61a90b6f50a38ed6738684f7262efff28aa3a09f1519d83ecdc798312ce
ze47f9fd52354f587aeed543507b3720f6fd1200b344612c4b447bd1a7f8efb4dab2b805afe6ffd
zf68b61f562922ad9dbd0347f81073737502dcb918cd6e612de2b6502d55270f613481e575485e6
z0fc7f494eeb52cd05deed6b08d5ccdb39c2b57734fbb6d985f6ba69c6b57063a188e719923e3a3
z27b200949ac7c0d41aacfeda8684c058b2b21fdee38b6291fe78bee26b90e237dce0b9b77d9358
z21987a7fba2974176c6b6bbad109ef217fb4928caed511ae3add4ce9909049b9b18f98d39bc563
z65d29624ce110262cc6f9f9ce7104ac53374f6e040ac96f43b340eae4c830d2b6cec29567a6b71
z57ec8351782b08aac4717c967050adfd760cb6663f54d45b62997ad68b036842ff74f39c33aa93
z43a69f9e57731d686a3b1e5a7d131e2bffd262a8e31a5e9324d0592750c723fc9766335ca4be72
z86f91576bbbdc1a1ac09662325343e6c1d432992e6d0332cd0e714ad1e3a52ba4ffd643a48347b
ze7b2d313ff8a085761a067535999894e5d413b673c635a9873f352c3f24240c651c324f31ca99f
zdfeaa3877e19abc391278692efed7b5e1b3fb458f74b510ea88ccaed2d334eab553dac88b71a51
zdfa92fd5b34e988db8f6bf8d7616a2725c333d6910cafbd68950479112b228c7f49029140f0d7a
zd6bff2abf37168f711f1241c9181629d4fbcec584cb45d7fd3c226d3dc1e6af9f8f4d2d145b794
zd2091d891d52452fd79e1080b5e474c91f7d344179f48e3fab139ab070015c0e23a34e71208227
zfa1ed8fafce318a9ae0c5d7e14db38a050e318690be5393c4a3d13983e5a54fedf3b574404a99d
zacc1a9149c6138cf6408c138d9ee63259a6c6e6eb074888f362cfd21dc33f99776ca54d5f3a3c9
zce6459aa7bb0df541de1e6a9bd892b8bb16efb1f60f98eb39c8718cd76e7f8c3e551e190b52661
z6270b2580192e87590ae83d8098f31a427aade2f6431756322fc51e63b59391e65b0e64457c506
z50ea59754ee2d7303008dae856f9e9fe85ddb8f787fc156de405fd2c7a7fad01dcc40b3a9bed31
zb66d4129ac95646aaf74c9c5092ccaf2dfae05d733a1a2102dd1fc589b99716b463505d716f0ed
zef233de54a311300c0a55ac5ba7319fad1b0854b88ce739d9f7e87591c15a7f67d7548dc8543fd
z3efbc0b6d9b649980e6fd361d6ea4fbd740bef0d2d425904c9446e570cff1fe63722d1c8026ebb
z61265d5c21fcdc09e10dd7dff1818d2c7918c95b2b27e110aeeed31be4f86d2a8a281b6c4eeabf
z312ebc186d14962c997c9d32755f60274a48b1a6cef9d612b8fe5ed329486b477bfb392d670490
z8d2806f65f9923459bbed901be45faf85e1d2e0c6985f1a873bae4348481fba912e472ae7a4fc2
z7662c6b995b31f93f5b941aa71fe164cc98ced307493caa407fcc7b97249d1e4ab145c333a4baf
z3325ce186623de981f0bf5617c1bbdebed584bbff5b8cc5c25e647b4674f4755805a546f6faa81
z14f5eac26fd8b3e2743fb13172070f70fe7d6d96e7bfdb0ff5cd5fd7df3f9184b501e7715ee6e2
z40f0399dc55ba7776b1c1b76a63de2621721e154270a5f45679caba14a446092c64b192a620dad
zb8fa7ce43b144681bde829601620cb968b91b091255fc8f0f507c5c7319766c1af235ac57337ea
z324bdf5951d90fd2065512599b3c086e3e7355f05643d456a564051c52f11b3f4b7787f4ae71a3
z9b91caeceb72d58c2f45a451af2c29f9924b311429b1987f154dfb5c3760ea6e94566e84139a65
zcb3200150be4f5a11bf2d12352e06dfe593d779af22a718f51014a6dc2b28c6aaf47a8b3d9b705
zccf30759b62a72830582e497dd14e417c0b131e9209ab70699e0af834cfac52c4fc06bc204395b
z5a0d9e39da649ffc5c80ff673f5bcb4c22290daa0598ea590866f4b198ea241c4db9e62c26979d
z5d934350d416a1dd054bb7996ab5b88bdc8b7a58a67ef0a0229807f0452f39fe46cb5b65998177
z49f0ce51bcad3f9ad6fd77201f2be5568e9bd8526c65b3210951f112aec3a3e57ac675173fb013
ze2f6c51e75b85383391902f19a3821e8c0c1a6824acf21742e7d272bfde9a5e765447ff4617b12
z1add3769990a1e9a6a0a5b4e882142a6f2344b6cd9e1ee776cdd82382ac4359756a239bf15eede
z669728be4c816c91b63fd9b1538b0acb676ddc8abb562be2d2a2f41558d8ba1100ae3bbd150c37
z34986e62815f941ce3f621e49e2b0e38af7fc55315512750c6282d6149aa16c4c9ce0fbdd7070b
z61d43cda70cf888592d2284636bbfbfe4cb3d49ea5bc9a3e2895aabd6fed916f0a5a4cbfe2c44b
z7e89e98764ccea7cdeec04092327666fd9a61e47e32c18bc1698001e3205e3dedcb9692d099eae
zf5e301b07fa89f8167f369eed811483c162534e6c7e118ffabb5e300ad1a1a292ec6d7e819b167
za24d96e434b143f621e76aff979a8ca4a3a4d32dbb82b2eac125c0a1445cef2f132836e02a0a91
z39034ee80d8f54e20c08e682c0bfc420e3c68b39e0fa514b7260e9498f96b112915499f802ed40
z7c3cf2c4bec374d188364df53009637d1c46023b60040f6cafa174fe0c98b5b780d72ddd13e042
zb525bce78e32306832c472218d0338c5845570e9602bdf660cdf9ade83afdfcf1b297ea268d99f
z3c4f3a6f2201444b4547312cb972ee7fda1e27d20237fccc35199c18025e3ff4efd4dd9d0ed704
zbee370fe15d6ca7ce641bd165564c592eb1859300cb4a4f5dcb82389e80988e328297d46e41c4d
z2c3b9b2449284ce883605ee2c774ed14d808406bc18f690159d308d8304d34d7dbe70cec1569d6
z4c72accaa4532d139cfa2fa263dae943921255c0a1448b7137334a80e1214f4c5eeee1a53db2cb
z62660fc46fa3b1397491f902ff992781f4d392ed33fd2b7c9478bec7df5c692d6cdd596a730ded
z7fee1f75245f79a3076e1e2ce82ed14644d00f736d431b2b57bac8231db7e76086f7397e7614c5
zdfbf021076ad160937f565c953dc585e845f97d37ac666bfdef0576d73efca6e8f896b23fa3899
z837441977e84418e096462d15d9a305c462702036d989fadd5b13812f251703a6918cb0d704211
z4cab03ed497d768fb282e01ff946b3b03043f5cb5ac5049a181252e1378d3b533848e0e20ed9fc
z4d9cae9996af78b9a0e7dffe03e4188e830ae843824f2839883430e5a672d41a1a2a4fccc7b7cd
z87b3b1eafc5055539de206c18cc71bb9eedb3bd1748c28e7dbbf7edebccc2fae3ad414746446fb
z08f9d1cfad0e09d5e0159ac8c5590ba540b358283571ce41998412c9bb76df7b696842eed5a9e2
z399b1d3736487b66a0ccc22f411b71e5fbb002812e96b20e383edb22548fc9841ebd0b84e5d1c6
z16a7d0f3c5bbb983eee827e497de8435587b7ee1c9322a9afe2ba10944338d7de7de686eed3c83
z94f5a18d8224f7e91b2f9f0dbb9fd2c8379d57104e4b04d98fea02130cfb023b23756924862b3d
zdc98a0d209be84b6bfa99fdbc74247dac17d7886c00d0687cc73a9ff9455c0618bdf30b43c586e
z17a3bf9788e3c03dd93638d4ed05c7b76c73885d1b2fa1b663a3013c4ea87e2ab601fefa5c6947
z1988c25cd0fede2673fe56cf6362777978689486dc20718a4b1574769ca97a4810b543d5c38800
z9a1b2599d3d4aa5a9445193e1d6e1c1920cfb90a16df0d9b6d190ce35e1355e94034569b349e1f
z981f0d529a5ed629e218c3f328a0bc3bca7c53e8b1a503a7b57762c06aa61f6efd9cf68773e054
z4307ca6f530bec2bf67c85f972ddcf6af34a49d97cbd5dc829653e9536bf7f0073123fc12a0139
z3655020fd19ee0c9722eb14b8123196f7c7a6a430e5cba4c1dbeba306e62fd561e49a7cd4cba96
ze90fab94187c4a3afc4d8088d8991fe4e7af539c4fce9321363ad6525e1470c9982e0ef48b59d8
z7369fe446fccac0176bcadd832d8aacc2df0692f21d455e9e0d79cefb88deca5564adf2c7edc38
z4e94954a84056edcf47baad9d620e1cf758b3c67c63dbb3c196be6a9fedec39dd550594bcedee1
z2f2056bacccb3822ceac30e8053d880ffa49e70e93b7f9593798ceb9bc6c0e4bb5c14251ab2916
z2869c25bdab0bb93a72a2b7df331155acd26a314bc1485fc74152f3b2ca30656c11100033131e0
z38fb093000ea7e51b4b7f0bd73759f9ff1e73a9d58c24096f16431f66ee6cd8ccfc59f6732351a
zb58c9894b3acfa9cd0fac1a171a7323c35b701ee989228694de0eaaf27fdd5adc80c44ff404b1b
z8cc22aa6c6eb91d2b3e45091ded262e4bb4172ce09a399513cc539d61507d64b7ee507dbf490ce
z1f62abd239396a27c02ce3da413e0159f6b7e6e251b2cdcc45add3962f66c886188efc8a3152ad
z6d1a4c54861bd0d8b133153061f8aa97fa47dadc3fc1df4f97d7075ab97b5bf7a902a1c29a9f69
zbaf43493e1df5f153d6547de0b3834ea8bec81c4eeae00f80e9c8ee31463b11dff48e18ae03c48
za0ef6c3142c0ea92b88cd9ffab3f00edb225739cccd9a7a21356fb72ec98ae394e732d93bd3600
z9c483fb292efaee14c6431d0c8887a4fd9d2e213e92e27863b47835dd02f6b73c7e0facf3080c6
zbab001057362a9e91e9486d94cedd88dfac3b324706a4a3b9aa556c4cdde823af2afe5801f198d
z9c1a68e67b9f358a859c13ec22370795b49c128d70107a932bddc2a80d1bacf17cd3809aa7199d
zd5240323977be18d86c5c445ca0ff207ad9a351b6d6ed675fcc99ac275f823d76df2cf9cbe8de6
z582beff17c46e46fdab9615299d55624315f6794eb3e635546995c402a0dc8fc926f16c82d8309
z0e6ee187ac507bbc9871d8acd320f177ca2c88362c5545fc8eeb999cb1dcaaf75a5a97e6724a4c
z965ca882207f77df1d001f97f8222f411ef230964cbd816e38cc7be687480575a979625b4334dc
z97e257d3fbef0ac10a6291d9519f7623f92d967cf2f94fa92d40e91bd67dfc260c11a1ba368b0a
zadeffa39707911bec28f579f864e601d1c886bf8965de0a1078fc276d123cedee28b25e1495613
z7941189eeebb2e6b56c8cccceec656034a23230ee64428cd5f15e883cfdc221972340eaf78ddca
zae43b9fe1158c2e01df2925ae317678f36111d40abd01bdc2afca3011c01f8e175eaae37bab45e
z48359eb618e13557d81ba877d5fa35d2050edf3d88b85665b8b5070553db3b72ddbf6bfbc91722
za95d210a212dd6b89daa17db8429792b03206054f998db28612e0f0439cd8bb55a75c70355b799
ze9772c952132c9fc9c457f3ad552dcf29b99972c9762f9831e14025651a0b75c498c0ed18b7ab4
z9ef56c593c939622c0e2e1bf6cdabdce48676e395a60dcfd4066a6e0df43ab6d25689a8f17294d
z5cd528c8bac5e773aa44de550be748e7825d787fccf71d4bb52145eff3687f3523cba92286a1ae
z972540af3a3866522310b96ea2eddbdeffea610d288e58e5e6fadaab74b3a196b4dea7d76aeb12
zb98cc48623cdbd1184bb4bb2a771f904f775052d0b0fdc3eb13a4c523e7435098bb8bd06fba060
z31a88f74ead69e639501ef237b3c207899b636e89b2b58b67fc61c1d69170338d8526e4d5ee955
z6bb8a0e62e410443483aa8fb30590a4bf115c3e719258cddf2397ec3db33a4c08d2c5e42a293c6
z6a0a3e1f5b8b4a256c7fbdf340412c214b8ea11a54c454a948674d34165bce4d6caaef352bd577
ze23c3deaefb2a1e360d1ccd12f5e287f2badfc08c39af91d0aece1f92086dd79228831f2f44773
z47b2a195a8c41b4366f8d4cced4d7b91b17cb76fbfe789a87f69ecb6ebbaae633a83b3563ec998
z7a93b8018dca97472f66d47b348163b86cfdcdf7d7ec21320812e2b118ccd9672c1e7ba3bb60bb
z24a0df5d093c414f799b25f7c1f4772f141c09aff8470eed364ebead329c1f7f77838623a93e81
zf08e32d78116167f712f0450eb2ae387f3c9dce4650d3e1ed46f0840271fbc05ad0b16923bdd92
za8429ff796f418b6fb4dc198c337454bfd1efe13c5982ac93bc9ec67e1af8cc5b51fdf6efe8ece
zb50b7400923806ac32512856bcec541d48a146857c6b50391761732d8641009f31f6f433ae3f39
z16cf8d3402238f6397d799050591a30c9f8b4383e917427c5dc00478a7fa48d3aaf479add17ca0
z7747bc985b1d731f3f108b00745a351027bba5a5c969af258121999ad667419e7db11f9073fb52
zc4fcbd2b3d9da92e7a1c2adeb8e90e0feb32602bfd999bcf174b922962da6edab75b33f6b1b15e
zcf2e74556ce77997c7618aa9efafa8eaa0a6c65dbe6aeafca5e6630689c582e25cd8710b7974cc
z8e2771bfe7353d09b2f7ccf408ee04ef3cf0cd80e4749082d4b45066c71fe6e147ccdd001c1f75
zfd346ff534419dfe78b783a9351adbec0e257a786512e88e7cc65db966b6e6176e525600a4164e
zc40b7f957fdc8a00295981fcd650026a60007691c1c8f94502cbf7849e8dd4c9ff9302c7a04da0
z894de3a5f204f3a032d440014c29caedefd0660faf5744939c2dc2508c3525b50f0f4111f9dab3
z3ac1e7d921eed6b122f2cbeea528763f3b487f3febb17e229d4268b5e4c518026b6d3afbd12f7b
z1576e53a1df7ebe551d8f9e23f8b5cd05a629cfbeb6352aea448e7ab1541a1839f11330b009f30
zcd6a73ccdb0e8687ec98d77aa21651dd6fd7f9e2315faceacc97fd73400b69457fe0eeae051b93
z6f274f202d0fe3e49df4def8cf2f6e727f8046f418ea5aa3f6446a73f58dfb8deebedb084900ea
zfe92a56b3b0bd1d6e021cb383a6ad636bf7bca3653226be53a191f34c3c55a81540f6d2a26694a
z9613eb2c63c9ba3cce7d91ed033206b3b2c23ae690e2635ffaa63573a3f7833c77dace9508bef1
z0de780b41f8a8a3a0fdfb7ae2f3120863094942da25220b6e6a5dc6257e3bb06a06a62e381a35e
z4386dec85776e008b30f32291e6b2e1beb7fd742b790a8a63c223006bd6e8eec64aae197f2b3e5
zd624de3e7dca622a688cf3266ce975fb2e875d4e14ffc91f6790d7ea8696b4c340148097d1fcd8
z3dd703b9768c1e25a3c1f74fe82231ab59e109a16c3918aeab8278213adb04dc7fcd2cf29c560a
za23b3f79cbcec1e2df14383d3faae8fc03633f65c1b5f203ea29f6e7fdf668e0b0f7fc8864dbc3
zb04ce95e365696e2020e6e4b170bd088af717fca0b9374bfff522409f3687a5c47c3cfdeec8b5d
zebe35ef9fa1d504c97bb96d3c2b0b92c2693aab25db96aa8a5fb35b98eafa7c43b50fb0e7aa746
ze0f1ffca9154d39afd96ed74b3730de1001e31496e1bc6f231e3dcd4282f703c6dde179a892bfc
zd61d03291e329a7d7e1df8192ff0c82b5474f1c78fba6b1f89a4c4f0f68609fcfd296f605f2611
z509eb85195c271108bfacc6f2ffbe3ba551093ae2b56d7d7f078939e0c75df42d3b8aa7d63fe4b
zdc675b0b4baaa21e7b2f5082bb1cd12c23e434c5ce29b14f5f959176376812dbade7f5af673092
z935c625d038a124a70c3496fe0ee963e0428f1a98f5fce7eafa785d95dbe8d910bb7e88b5dc77e
z3adf90689884ba7e6292153e28c47993f9c1557d40defc16076fa73358fb5b2ecbeaf5d5136da9
zfe2384e6a6003840a94c0763f74d05d82494b20f7e7049e6be495adc69a85f561c5141b8a9364d
z23c47fe9d44964698051940d8a7f387b184dbbac7af554d81e3f74f52614955280903a9a7fc453
z72019a9909566000e60bb6913228cc3952485870cf15a3b33ab364156ccef5681276252370799b
z2062ba30ffc58b46a43b0455cffac3e8c1f5783d836374f01114d1d94344a220dc89f3c27c634c
z9269843db3ca390ec41431276b8e407cecdacfba6d99a48fe7cf35adb2f9f2deed2efa3355935b
z74ebd59ff2f2f5c13476eba03d4becd84911d3a84852df0f69383268adc452834a5a3754a307b4
z2a5a433d7df5405f5d80702fd2cd21a8fac2cf027e85b1493f12d437d6627603b20953ab01e7f7
za5733229a8efedadbf15fea55c27006d9514d05f90489e96aa181b464c99d2f8c47025eae1f892
ze92ee5bebf96423b5decd1741d93004ec1e38675be48eafc570e8d692c471729d4fc61604f994b
zf9fe0269e788146d6441277cb312ab7748ef00fcff89d6beee286ae7738b22f5b61a9baedb82a3
z762b2ccce10ed73fe80acbecb9536e8b147ebda5a2831004ad872d314f2a035a14b52fe8d69123
zeef898b3774f8b7af64fec3d06160272f35193fe333c9b5fa3f328fc5d26f24d5bcffd3b7492d7
ze9a2ba227fc2c7cdde86306d1cb4eac1b935a3e712d6e92bcfb5f53d4b4e474d9c9fa8b7f0c5a0
z265ae07e84caef78ba9365a94a1f538c28c60440802aace87b9f8479f1a174c14705d57f615546
zb7a41b3566d58b35bae910256377dd4283e192f26f8734dce274f7fe5932d3375d50e8f82b863c
zf971f1f67c7fabad06e4b4110985ef123124c3f4c735f368ae9df79e8787d403ba04b6f264d5de
z0df106400eca93522fdff67a16600e0dcb5dd25067c1884e2e7752a13a8194f3ebaaaca86d7534
za54c071645b3d7d201c634af0d2cfb7ad8adb099a9dca423abf4e5e357a106fb9502451d22823e
z510774f3bfbfb78aae369eefcc5d2d43d73d0c4830e3efd676831cf277102cfe086a1bc070497a
z24e3b2e650ada1b06ddf7047ca811337253f67e852a17023361f462efa2e74f305dce772fbc0a2
zecd9e14658540d2b646a0b29fdd486146d393b6bcbac48c19bda3c6a829534bbfab2e41ef56060
zf2d4dd7621f64d4953291919ee8572a1aae9760f1844b7e96cfcecf1f9bb58e81613caabb467f8
z64235c12a5da489ee83fc5e4b11656b27b22f936d0b0923646ea4df3af1fe746e474a91867df36
zc47d09d0f4eb1179886ab6d9caf50ee29f8690d67a5997a635fc445539fa562b8c5995b19ba483
z1f91553c36399f791e2886e6f5ec556091c4db75b5cbe45d6517b5f38f99d923f1c498242069a4
zac819d6aaad005342619b66ce9e6480a21f0d86cd10d445c5d07092e4ebaf22c82be0dfa5e4c91
z5c227320dc6f499500897ad9ce475b932e7b054aa685fc48e04ddcf9918a0b2aaff8a79225bcde
z84c5e29858b70c2eb1551316253ce8c9ee51aa7918a82536c9862af7c8d62488f2be95a8f3746f
za0be52c8b964f9bca64518459698935f775816f9d69ddd6a18463caca9b23904fadb1d3296427f
z985e3527b715db7d94ff754fda7a80a857ae67117554d72031c5727637b5d7b9adf506d832db83
zc02378261d243fbae1958ad22d09813658619d51c54f7db347b80919a1c22841a295d02ce19271
z6098b7dab3e22bd4821e988c8975eb0357a6f9d1967c50503b7c280de1a89611d345736e92dd56
zc26ee0aa2110a7be02e108d7d06aa73de89172c26d2421ef50f3ad4e9d3f7c7c92a54643d70f9b
z943e699e5b6b209cce635ad5e251c03385fa92ee4927a1872ee92b1f93ee045d5c905a45058bb5
z2d28c4ed28353a7ccd9df4a50b7df5f66534b471f745149b0f86286273ab93f81a3081335425f0
z04a6a7e41e891bd3b566f4036af350a09957edc2f5ad94c141a0ef84594df30478fe7e452c99c5
z4d2d65f5396bc31181cd70f227187155d65de33f9ac5e0b6f577d87fe8c9a79d28bbdecff48462
z51c4e6be651436f137bcb4a2a00748d11dd30b9976fb169ba8c9b4466f655dd5c98a21eaf5808c
z7ef8e0732f38f291ae96a7f1ad742cb43f110b2e551c7cb0888c6ae7b51576c3e0c1918612fb33
z8cd3350d6dd583f02db4c1ce3aea1e2cd6b0a42aacb5c1c38957f700548f7a6db0f53c9d92ab7e
zd3232434aeee168d3fc2bcb90692cb735ced1d097e4bd65b3cb8d361063eb20f45c923d4d37fa4
z1650771c692d55868780a0dcd62e72ad40b9ac55014870783e50398184eab10a03bec45386cc07
za764e87185cd8d959d1ccfc19960f208f2c2a4501af51b0d4fb2dc315c71ac71bcdbaec214aed6
z520ffdf94bf6751bf9249cb01139250200e2ee0700e466beaa6b2dc3b06a2e3979dba0f3888060
z73de976afd0d7370600c21a4e94897c67790aaac654c1b5f3abf4ac4b4a1fcce195ca84c523e83
z2f6c3d047ee375bfe459ca65ae5b1d6b4872efa4ab15b0a198f424e7570a66cc85c3c528849f3c
z6374c4c13d95b2497361f0bbd4282da2a9addb8779b103679e31222e5acd1088a0c488ea93de82
z95f54b3d167a33fd187163c6f1e37892e57312b3afeb74cfaea423cd7d612a64c291785d85593f
zd77de09e5b4a95140a85747dae99cf98a309739b64ed8e39d20718cf8872fc9e320fa795cb3828
z4256a55a7c9ec7449a9a13a91fedb4d63b375b654281899197287bb1b93d900542020887545675
z6a2f34fecc3c303116fe9f536da3f398b2affe144258f5529fc7039436143068f1c8df45d2d8c5
z9412382e67a59953382ed573596c76fa15689462d0b15f5808c47a8a78518f7e15ab9d4dbb75d2
za4e5e4a3fde3b4eb26ccd2e1ce9990d0e82d02ed5328cee5a56d556aebd933bfc6c8ac77fcbc22
z7d5a892b51fb43dc841296c3719773ec5e58d6bcc81540f5eb0438ec134c14a794ece39c3f2211
za8ab3244a1f6949046769381946236497cdda5727e41f80a8a0d98ea2bacb9fd592e93c3527313
z4fd3c6c90489b2f901a3a43ff2f813a0e34718953291ae6fad60354db8250a34f6b979209e5158
zf78f5d318f224452afe1aac02e658a4862d18b8598e784a0b9ff262d1c05e56a2e79a9907f80a3
z70b5e480190b31d3b433aa7ceb2e09e0a46eb58def08952f10a642caab6cb84afe9c2ca5c6bc64
zfe0e34eb2a637fc0c8542c680e0b945c0c18ccc9b681d09276495aafbe09ed73b70c379c48efc5
z086dc4a3c0c8214a8fd29bb3396f93fc678a97c7097f8a483a85e7137ebb66373e133022b6281f
z8f35ad835f6f2fac0e8407a8bef949c5546dc2b6923ee4ebc5d370460fbe99bff5aba6d6b243e3
z65f75a4c2718c55505e437e2f3fa53a11e69a55ac7854b79b1c84bfc4989eccb8eede935483c1c
z457a9e7430f2abda2b2a8abd4b0fec68120862159c492c8a41d1cdc3930b8ee3e4cda8145bf450
z065c5f8bf7cab74716110cc467202f9b9c12085816ba5597439a1e4ee7bfc4b9886d6a406272aa
z30f1013008c686a3256024ee2f7f1425d2789ece23432f68ee952e9a267e056e76e3012173ec04
zec6445a6048bd5cdb921a2dd512e7013cdf43f4a0d03a760a8b9a4993d2b45b0c37e0f0a53531e
z45883db612a44d1879df8658b21679a398e3f8e18a34276dab27b40de36a936e4b71234c7e9f77
z28954fc646aa9aad4203089fc7f574f390da3c9e8c6fde6838c013e9c30581f51efd4561cdb81f
z30888affab36d745ad57482877a6ef2b91dc302d5f0f4907eae5ef26cbcc69a6e1a3628649914c
zc6fbdd34d54667a934c3dca70b92c02177edbf59d467ab9b095559a98c10debb48887948a863a2
z34c98d95a8f9c8ee893a3c2fe08c3e88d5c7f53652306a4208a3265a32f6f39f86dc590247d132
z040da92d8cf112e17fd860d8e168302de129064522fb50bb59213e90f54f286b69bc1c9409aa5a
z401a3c1a5cb43d832ea840d78a1583598be9832d449c6482ddd1119cb1a094918e985346f4b90a
zb4c48b1ca791b36c2fd20c04b7ac8364ed9971603fed4e31cda0a9f8f6a217699f2e34e12b6935
z9691f8d3c207c250b0052b908fdf3f823582e1d83453da533eb91449d8390a004ab348470a094e
zd0ba52cb0ab598ccef79374196d4ceb22c8363d368d8a04d0f86aef219084f430999c1cff2451d
z685e4fa04a3d43df98f6f55026e18030e3ee766271d87ca0c7c52124496fab71e6ca9880702198
z85eb2dfdeacc015c2d54acee52b913c7ed9153f447c2fe6db4e74b3f8586ae9a51a9ee819857e9
zb043d34def8f09f5643ecaac4277c3f60a745522e7b4ea30c84711a4bc54a1726f8e0e24e419cf
z421d8456a064be2ebb08c589cc9fe4bd9c65132ca4d0f982e86c50a6357eb5ad4e4caa05446547
z0dceaf28621f82d7287286e13a4291ae9e567c714bc1dcd4add9acff6408aef364997173d94104
z6e2c5ab453e748af7db4deaa4498154ee9031bbd5c72638abdb86c2c709c6c2de5114cb999255b
z5e431d104a39bc7182c06d59e43780283e6804b4b9a8530805701a7a594f8c7e841161287568b1
z15075d616aa5ea540f8e2294df0a1e36a54ee126806caccf10334c369b80938b88e140076b8e8e
z426119f1a43e260c86da8d5038d6238185c34ca3406f66be521cdfd638b78e7fa2f69d1e1465e3
zcdd2c3d5e45036076608a005f63ec12ccc1a619aacb07073a20d0fba2429b396b8d9f33691a722
z5a9dfbc3798025e409679022db157b3ddbd578ebcbd4ba8733849dcfa8a94e94eddcd30756402b
z2934d550dd0b85b7e0f385eb3c99c692d1ee037edcad45547b8fe10e3bf0daedeb620f11fabed9
z26e190d24623858bf3e3ebdaec04e216093565b5a25547e0c13df9e1a19631e282a1c7cd799ac9
z33fecc0e7c93b346d383e362ed309496469e0b5e2cef3068f92261a054262efdb3e1177852cbfe
zf4b6abdef5cfeb08873143c409df60e47e9ca5fa3d4ca071347c43b98b5de5a49b61b1903503e1
zc43a8ec8f1a9b961e420ae690c8659cb5638af063a150c55fc28390f7ae29c3e814c079cbb4816
zb9cffc3e7d8467ae6a3ad924789461bc8e4eede24a81fd6cc5d180018f01632ccb6b04e24fc892
ze4bfb1c8246f01859404e3031bfa105ad481e15241bacb3e985876a67edc3409bba2f2938a6291
zfc480582aad66761453badd54a6395b349a848912452cb4f16c7d0e3d6290ff53100fc9a8e04e9
zd252c9437bca7cf4fde5828741f1da0fef4221f4a303aaf2764413d0461096f510b36900d950c5
zbe35ec945776efb08219a171b24d2204b9ae62405c0a93e42b436984ccc83f8e735efa0eecf594
z16d12a0fa08da245da6400c7690b0a0a70e247f9a73cf5d0cd572b32ed46c8adb3fc5192746510
zb49b4b65f0c5ec4867a6fbd863636eed88bfe679fedea918596e1a9f3f6963a333651bee94a7c9
z816a471a36265b4a783f84e49716a5c2ac0d139106ae19d7b983d73f0511d898e3c1bf8d10f07f
z3312ce1fb02ada7fe8edb9136e2621694471d9316db79f78376c8e79c88469b3d5b59cb26b5575
zfaefa3b055c32f40e255193cde6c231410477839dbf36f6cddf8f227dae2275c448ce1bc125e0e
z788e3f14a13a3156eb9d32d9eff8a1e3c89eec5cc61f49aff01ca907e57b5391d14050eed72d0d
z536d3c9425a3f2256e241b05acb88ca1c9ce7ad46a927162fe8a1857b87551d1eb83b0e1a08435
z3858d3a879bfa2b31a2cdf10d0f3b8580b228a3b51b359df3dda919888183ef8c0548f1aa5eec9
z16a68aa4016e3d458ea16298614e74a10f6553cb01edd7b0dbdfca119d08417aabad19af047e19
za5d6e709df3fcc9c4def18ad6dbd725bd50b951d7e10990e9459bf313b6af92c27bf07e41fe990
z1748d053f3b30e41349686d719047badadce9ef07a17d5ffc82f0b0fa109ddf8b0ee0dabf0ab35
za0c16756d878b1ba1c12aa7e72fc3f84d6c9499ed04ea96ee66edb0a73f2412b5679dfb3e5d606
zab5eae2ddc2a4f32ce540c78b05acf5b6176b54927596af1a413faeed21dc11dd62308aa71b76e
z32a3254a5a2e4c73d190952e65e4657b87463ea6f1da00904310953284ba1457133526e9af9aca
z81625975f54fc2f1c4c6c0f89e8f7a86de216bee17fc0607c16066010a86a9f02e79359801a834
z0feabdb92c6ff25c2de1bc2cba636d61a862f167fbbb174c53ce65587b22e7abdbf6444f9dcc9f
z6d4fcb6a1aac0e0b2e01df455611bc2b2e16a73cf6ca29a9fa1ba955ba295f2d020fb19bd983af
z834fffb54e484f58b31464f7b79959f720f8365672c7a7cd037ed81babf9b122d051cf04a54c4a
za0f4667c23cb920f0e35ac2657930fd1994e3649ef1c029b6068e0320a3ffa65693b29692a597c
z4765af3b8935862bc2d958faeaf51b95a2fab92c03a0546fae22c831337512eeabf029ce5262cd
z9c33c057d16b685b1b325ea266a0613189e0d2c0c8441715967df3daf353719a0d17f1da6da442
zc218f334dc3c0357adeb2934c7f8e6290014184e16e63abc1b43892d64ee73bc86d712da4993cb
zd58a5633959d12bece6fa98a1c8c6c4b0b66d4cf5d0beef3674de068f1057468ade2aef660f1df
zdc41a76a1b1632d844850ad73370c44b818604161756864145a3f2d47f254bbf82061c206a4671
z7a7070e2c8d51d7460a28d9bd5077ff94abd6b5844f9653499a975d26096018d85ca9abe55a2dc
zc9522f7de5751f957e188b90a953085b9ab845fbafb66467d82d91dadb19bbfe7828f3f6eec5d5
z3372600fcf51e03e00f89afe3fbe4e825c657c7a793ec6ebee7befb83fec3250f71cfcab158e8b
z4cd28bc959833add0ce0819393ae5fa8568a3f3defa7b30698287d0fcbe160615809e803d201de
zc2a27798e7753b9e753a84090a1d45106b6c6d7b5906cd5ad34e04f42b05877171ea0a49a6274b
zb5e25305c606f51b11ba4e45e26947e001e655ed6c9b2b8624d09c9167fca6a14a1dcdb3ab98b0
zeae8f513cc8c0a131b7d3c25901b0ade3cfadcca2e6f51d0c23438adb9c38cd0ff99d3be4276fa
zdda8576c13e27e83f29ef367c274c014a16151d855fa7b346454e513f783f546f73e9def989080
z6d3449af57dd21134812281899806bae1e5a0daa68d7b281450523465cad3e4765fd95f999c18d
za4bd83e045f86641075ec3c85ef850717161cd78ab4f371dfb1854049e962c9dc9e82f86e82a56
z3186ddfe487245fcf7eeb4ccb74a8aabe82f8585115213dda7b491df69aa2675810de842f04995
z4ef385eb62079456c01038f703175440159f72b02e954b2c547b779d0f6513f864e7e8819f345b
z3e19d37f501dba608e3620fdff76438d2750dc049aa471f1704807e14ae689d1b139984f8eac40
z7e1e2f8f6562f85b0710426364d20d88d34b3e3030de4c9bc54dcf61f21124e108c3a06198ccca
z66a271ae0374412cdc1b64bf806a0bca1c19d5cd68c7bf0f90005050b6209175016a073656f9a8
zf4f6c79122b1338e87fd8895da1ea452cfd642751d80817573ede2081dcd15013b0d15f41abf74
zbe8c07a78f350bc7da87e28efe28e4d3e983bcbe4ad66b4d88a85cabc4153776b63594d52582bb
ze870156a5c8a86d5597f0a79b045d11b3ef8827e9f3b1a2a021bccf65367ff8ed6754fec63b791
z03784478b2b7dae555b3c7f299720b0a734d5d8abf30dd6339d727fc49ed0aae762a48a8547f59
z699bc42148a74e5d23690a4e50419e3f7ce8b429d7739528106d29a993ff6f72f862283845ed6e
z3efe687d8d39bb3fa683c7dabfe31730cc7e1ac45a675ce133613e9411725df042a1710c595084
za56cbee602c9d876d61a08dea898f05123da0d0f366611c5cf7d5c16b85e2bc560e517b3bbf874
z68f46fd39d01ef4fcd1b2403296fee54a72dbc21205a29bfecff2c7ed44971c01e6dedddc4d9f8
z2970b8845017a3fd4d3d114083c4b28278e3fa0476118d44db226c06f5e8781c0fdf8d1ccb5515
z5495f9eddef784d1b1f2ac41a876bb4406108bac4564b8ca50037147a2cf9597a84e38dab14297
zc9149e57e5ebc2508bc2eaf6b5006e1bd8698021ee897758efeb81bd0c3d333511df55da30d18c
z77c1828435902046ca759ab5b7f252df6dc510b9b416743165a615440d1d33a99b96bf8556f67f
zb360cd5230c2b19b082bb1c376356f533ad7554a8010b4e8cd041138bef77a724739f356c5a1c2
z5b0d20be2940e73a5fda7487dcb2bb6577337710c0a93b11d8d5c504f2b8d5b7c21190aea0dee3
z485fc89ba238eca11e991333a2aa243a83094005673fbc5503c57a1b54719c33de5663cfc8a58a
zaaff307ff730d310fde8adca6998aba8f89e317c01d78bebdde19a889035fd003585c983682fa2
z2c979a96ec855e48cb3f11ab42a825bb62d6982171511b1194895fc56ce36b2e44b4de8a7db24f
z0e08f828cb66b386ffa524d215170ce2070881fa3215238f6ac9abfa03e92d1c92522192842332
za4fd8b1a3c0a105d10baf19e04ded9d86ff7f3904f14564be1050862b74d0f39a8504d1e893164
z7026d7243c6276bda3af451aabd80bd8e7e182022b1d9921b9650706f1ebdc0d49d801c722e916
zae353e68fe6150499776b6a94ed0afda1afba782b80320b31b76f5eb5b281a7621198c558417f9
z9722c2c826d3ba5921045f99e5e0af3d71195ddea7ff536bd56db8185642dd99d67a45666d0cae
z744a73b5f6a33e070ce027fa1c61dad0b108c4ad5dfa13964841b9916f0cd3b12997465be3267b
zbf68ad84d76d19b73e9ea834b8d9b86c059b1b914d1bcd2e6efed561c182743c7992f1adb3212d
z3d91e11bafa95bb4a23915eecfc5bae6fd657ac67375249fc0e2701989e8c255dc025068680cba
z9d7d4f9c53615a2b773fb362e9ff7492e619ba5481f2ba0fb23e66555ae1667550e3eca964b0f7
z894a28fa54a9224de6b66ce2c85e92a1f538940f9a205704d0883a661e6e75518b90efcf8ebe65
z70563c7c9c9741739a38aa600407ac2203ad0ac33a89b12feb9b18810317c94778ecfcafa6e731
z76c26408bc7b272964e835dd48f41baa11a6b9ee8b36a18dadcd7305dfbbd7e0df23e3515d2d36
z239596d0765efa68a3285043b981145d06216f1070101e3a74376f6ac202b44df315e1a2831cf2
z9ed4bc740e6902d3a9ccda9525edf052ebf6d1442c09456a1bfc4edacabe9498af3e34e6304205
zb105cf5c102ba4ac5bbcfc03b19fb194c2c4ed322455d29aa7875d605eaa71a708e1d9275e3f3c
zb1e60f0cefb2bd4f4b218453c13e209a49489b58f3453a7997187be149f0327f9cfb02b2646025
z50f6b48fa5881ca2afc3eff44ddbe8e9de012be43273bce0f203d35322029beed4474847b480d8
z0cc9518f9ee9da453bb15e76c85fb85839aa1d1bf7284d828a7fd02fcd81821c9e53c369e09d69
z01be59e972480e326350c7bf10a2f058fbe4e460078d542250e7ce2fd167d545673d6d2326b3de
z5bcf2c34c68f23190d75676487be12152fb4ff4dd0709af76942f4045dd2002d10288e5c78349e
zd8ca8bf653d9e06e59f60cee0c42d6d97976eeefd50d9551ecc3ea8e6cd43814a3453a0ee5a5fb
z2021544cbee82061d926442284a389e9accfaf8be5148030fb9890c0594f839765f0624da32a01
z5d30103d8c4debaf88bd996b045c4cec3c8b331bec3ade863197e795075c5051f18f3ce3f68a1e
za8f40cb954e887b9aefefb0951bf3fe04b932bc1d75ba6125530ba98cffc72fe4152f30be4b804
z341f12aed6c42b80a621fe08632aa4e1a69494f7a0e0ecdec9825d721bd36e2c7e23c13b4300cd
za56ed82146f54d602c835ca35e5a49c778fd2feffd6d5637f4322c412e714345066a7c53ea6e29
z4d08660af057b74f1172d23e628acf0b2c4ae30aff7d37ee029177b0331e86449367d444ed4d8f
zf361d75207bef413011359e444a55465a4fa3546bfe37adc97e06dc97f9ed6aef1cc2cfa3b6243
z1bbab7d2a56c9b75856d834efd85eae0b2fb1e9798bcec0f83edf90f7f5aaa949c47a5c003806c
zee6670227f22f337c6cd8f6136a88cda2dfb881c339f189022050f35f053d3ae198006b3dfb72f
zc110bb93bb264b93d69116dfba5e282ddb13cb21dd8f4fbc73cc189c68a4a7591f2590a62f38a5
z7055885fdc9f6a7d6a4a2940dd85beb63723586352e79dd6c622e771a506b6600176c9b0a20550
zff3752c65bf2311bf8dbf8abab72de6dc4cf015f0eef5aad19f9630ab2635aa8b0cd51db74ca5f
z24922799d3d260f0611a5c23dc4d0ba26265bd64228493c37fa06aac9116a88ddc0d7f76ab2716
z2b2a2119e8ef0b592f2ba5d60bd5345981e43fdb1bdc1cac644694026a857403e7b5239087309f
z9a7550317d955b2b362d7e89b188abc427d618a0cf2b19cff45c4f530a83b28aa3e7303153317c
zf4f26d157f8ee343fc3b96a71d9cceaee0ac4ed25a9bfda6163253d63aacd519969cb187aeed5a
z970c8cb07224a51c2112308eef657ac0a696862aa98c39e33afcc97ca7e0d493bb3a9b31b70805
z05523dac53e62ee5595be21ddb817687566ae5d600cba5157c6df6c1ecb2ff1deb9da9270b0029
z68a51a9703512e3935df87ffb5621b5ffa545bfd99559014c167ccbcb1bafab573bce146447c42
z313ac1e16e26d1fd699d00e44c6a2c16d99b30e33faad15410aba032b6a47ba01d85e2a895552c
z8c1aadc2b3200a5126f1fad66245d5bfdc418791cb7d8061c10230c459c28f6ab34543806615e7
zfba0b7f053c787293fbfb125d7abffb3cca4f2e82f37676f12cae8a3222144da0719eaaa4bae71
zecb0de4bc0a6717f0061550f11f1c706eca786fed8dd760bc98384d6adc9c0b934dec0785f2e83
z70e13e2fdf562240889c4c5243c869623020f2a5b6e21d16208638c23898bdb901b7cea7884b74
zae51264c6eab095989d3a9d3909cb03cbd67b4d0fc245426ddc4521a755f5e0a442e8261e6ee5a
zf2660d683a05733621f0fd430b890e6c23e1bc231a12621e7dcadbebddc06130e1eaff115c8616
z7d7ba6298ba221f689beb13094427824d1e35143e9db9917a4b0bc32322a2ad64759356a2e9293
z539adb8507817d4db4b9db3bd8a69b3863d837f49b3a112ea4c2ffbb05294280016f90e67dc8b1
ze3af0f3db22f7c47e5380b602b727a42c5d0cc350cb070526745352a4bffb3c534c728732d35d2
zc3c16e2aba14577f876d684d5903a33509d114c7f857de0b465755621ac6a10efacf6529ffd916
z5e742d2b3635ffc3ab0ba39aa7cc9b01f2fe26270ab973a2cbe2a41dded667ea9b52991affa98b
z536c80f9b34e9781295cb682f0a54d456e1ca29404dd332e695a9e528a504403a0f3c82ab7929a
z767a8a877121363dd2487d30a78d4e5b3490ecd288aead78b2ee967793ced0271cdae6e91d462b
z804918853ede6ef9b2526c68f906fdd459b0ed5717463371150d047b68970e81f0385eef85141d
z2d3c5149ccf81ba7dfd7c7eda0e350a8b94117ad9431f71f4d2d1b2669323037d44ebe891d9ef6
z0ddfd5b9707cfdac322272d4b0c992456b2344bc8014caf21e2731dc980172c174832c5bb9a2d6
zafd4a3415a527f04ffd52e77c4d87bbca72afab887b6a47f7adb172ac028fc7dda809f62eeee23
zfa2c410bedfcbfb4fe77d065eb25ad00c4d720b607dc844173f768b96bc20b8afef2ab6f97739b
ze9fd93105b232bc1916d84ed9d3c5f2185bfb1367df30af446c69b51609fd2e2bd453870394758
z714d9b18940e66b2470ec5588660039210b9fcead6711e92ad74713db68993706da5b18bc644bb
zf93ed38dc36029757b44e4648f5a939d144b9c4f8932359e0cf05ba335bbd1d27017b01f521fb3
z35919de38debbdfdc37d41d14adce06781e43e03cdac6ce3211befdf56addb9174bb57425b8006
z89fc9b46be4f729c0f300b8880127ee6c38a9874d5554db79c95f6965fda19554c231aa484fd3f
zb82301e609c80596cb9e75d521bcc2119eb9f31355718764dd26588e663b9e9a6511856d6cd551
zea09244d5b4312dd57054e77a72c5209e8a0d6f16c4d48ad751063ca85492e54a570bc9548dd4a
zb40b137091d36585308547c68a49c2754a368f5372bea68357a404cb0e53ce25b2ff2c0ef16023
z677fc9f219e499a36d55a1c211a8408b8eb6f43faa18b6666f21bcf10a86620990e7c3049d6b32
z8c1b4dea31c75fb8bcb0330210023a469d0141b4b17617be73c19c5b48f1d33c65164a9a6972e8
z73ff1ecdceecdc2c8f6b741711280653d3970e485fefe23ad2dcb98c1ba127e6d1b70ac8020fa0
z8021202e467dd903f1f3a4c4dad3e94d9d546f3e622e6759abb6de1afa0975a684dddfc1585f6a
zb9525920ad8ad3655544f91ea4796645dc3ef2b6c7c36892cd94872fbc1696383f24ab2955f2a2
z75c7439a06cd846b6853ad1e3dd2fd70892bd96936b948a13b6914e20e5d3b7df5ef9dc6a0ea2f
z90e5d7a6b24a3039e67634321a7b34314dadafb8755e8c86d293ff1dd465ac5eea9480714ba1b2
z1d1eed8972f808e99af75e18cf887fccbd75c5bcef819a2031fb26c823f48255369e910bbe93ad
z5857e887755e47043db0702161c5f4a17b06729aa68dfcecece6811250ae32e162539402010be3
z3bf2988ad5c64a5582dc5594a7e8a1295a92c2c48275320acc02bbbc8f5337c13dd27adb657bd3
z879792c6c03b5cc83223ef13129a3c6787b7d3d82732eb15030c779d06087e3905a548afa8bf20
z3953e3a9434605a68c916a307627ceede0a90286fedae3aff1badc18265b56c82f49719a080101
z9b1faffa482cb633c8dfcbc1195dd091fededd5738125e44b2e6c53626bac9a4e147d11f6928f0
z3d7ac4aa673f93a93a87c9df811f2bbaa8bda31a05f52190875b6ee2ad36fdb5970571a7e4c05b
z176bfc3d98c4e933f5cbe348cd1a156eb38a9bbbff3c95ea7a541f29332bc736f662264ee6c41f
zc6d1d4752ee9d8080be3b6d16f7d5b2608475f83d9801abe9f6cc27ee9d6cf56792c060607ab28
z865241b31979172e6ed91dd73a3506c80a16b54e24d0d8e1914a744e91a8c616e171d73b5f1f7f
z9928d378c6389e9cacc6565622f26c384d9c2b66bc706cf5f9ad3b55ace6b8d730c53671be661d
zb98743fd840d5234a49d487168cbc7b4d6b359615d960a85e5e189fb47d6f0d16430c12cc9c501
zf06a62de5b6fa9f945c9f1cdb528a904f81506158ac036f7f7cf51cd1c54cf5975191c33d0c683
z96dea30867dd51c05732e72ee205fe04a4230f2b3fe6523e615e066b64b3e35aa78fc30d144f8a
zb62cb7d522b7180a42c9edf146c32bac9d52ab077f552c93a9f1b79b4b306a90c1003047d8b3d4
za2064de8a1fbbbad3fbf7be64437fa9f1552ffde6780f45aaf85ef3bea07faa4a993235ae74519
zdb709983822cba09bd62ff58bef87e29f948c945850b82ce0076387ed5f756c68fe6da0c8c03c7
z20f6f0f2b5851e
`end_protected_0in
`else
`ifdef MODEL_TECH
`include "qvl_gigabit_ethernet_statistics.mti.svp"
`endif // MODEL_TECH
`endif // encrypted_0in
