`ifdef encrypted_0in
`protected_0in
ze74c34e226135848fe16db9ffd31815111b6d7fb642c521a3f628cf6da949865580b22efd062a7
ze90adae0e65e66a2c36a587d0a790699161455169ed55a01f2084f11770a774ec4c588039b380f
z6de9c5084882a40b79a175f5c2114b2b6d78b070cb806e1c0aa9258297f4687ab308bc470f0040
zb0b1de382961eeeaf2e279e1462520fc31c119af8f2b214846f56c2b3cd2eadbe4099496abff18
z15cec83ec4a77b868344aa20ba7360908f5c0de2a79abf8b3534b883bb12180f68b5d4beb444cf
z3fba8f13afb0abfe8fcc4294810f75afe452434d2d0f1166236c82f76edf1e12979f04bc35693e
z32ae028996dd85737a8f5adc1ebb94f39c940246e887647b64782cd7ab429b0544c173176cede7
z01dfb26b1f73408344a52b7e1f117f12bb9c8077b34876c2e6fdc085981637012dc9754765e1a9
zc512ce062e0b8fb16a214591f5c81e1353b900a611fe1f4886b57940b41b7f2ce99a7b84b04b90
z916f717e73bd10589c81e207ed77ec660a8cbed5b487fa50acde1b055c8870bd8676023f21ddcf
z9c98cc47cfa2d654ff1365d1f45035a045a66c5dfa827905026201628cee5aae21fb892db766c4
zb5b1406e11aebfd6dfacc9da5ec03b70c276807a3eb15e28ec7ab1dddec42388b9424ea285623a
z248195c9f894b36317ca6e59c86f11031163f5f52d70922c037057ec3eba50b955600900b32628
zb2250f2b4fb3ed6db7d81b8ca05e994209e236669db511df2c321dadeee74880d12dbd5092819e
z312f2e640fed00f965c7b0e1d2007d987dd08e1042332719768f689f95a8ecae54578598cd4014
zf52c9aa29e5602a0a7c0b59ee67317c72101e7d1c45c07570c0683c158486b6e3157427e0a2514
za97901c629a01f6fd65b5a7f6f7538b7ab683549194b5767ec9f9eb38f388669f93633863ba210
zd15b4f9d05bd96c35341c02c93752c2344db76edf8c697562b3a09dd9e6ea71115a107694a03bd
z48c4beb95a5fdace643d8acd8693678fb3c10dbc716d343185d0f8c8b090128427948cc61f654b
zd79e08af23d1f841dbaa5dc1936e4660e1f04efc36d203629f18a16a4829e3b3126751fa196d42
zfab93a2769d0d4af5366799eff9987e0ad2be0898f05a8a7fe7be72a09e6e962114c35e028f985
zb4f3db4d71c39b999c96003b9bf32fb342a15fac3c4446676fc11b463a9620113254265646ecae
z71d7cf3381b7e84b560f223855b0b20038eec96c1ac4f1af8cb0110cfe327c79fcdd2413920852
z093eec9cf19ae3cd8a67022d07fcd7bc14320c1ce4d9db0e528514c98a62b5d3ec31605cf03599
z4d6eb850c37fec85cf69e6b474e171d53ee2bef5d245d9cea5c101e34ebfcfa73468705933e98b
z1a22aa5b32d9f8d3412392ed7416ae93ef2762a663e61a210309cb52001dcd4a952d8799718756
z65c1db60a4531864be9bdeff4cefb56beffe2bf29fc5f3345b63d7f8ab90e88a20287661fd01eb
z5e716c090119d5d4c08ccdcf8d33e906a8990d677657f34d4716cdbd43f372c20c4a03b754b7fc
zd09a688dec478294aa8052d341050720e84add185bba28dced0c27c13f7c8c7cf2b793b02369da
z080bf6eff0124e7ffd1e395669b8e0fab00d0bfbdb7b4de8907980f17ccc6a990eab828e203546
zc08cabef41d95483de759263a68379bc58694349f4d092ce1c8cbc4d8b1cf9a2a993a7ff3c5dcc
z09f2675b286e7c0bdacfc3510345f25f7fb48b7e6c7f9ce1da3d69c5c34d4db08c56127a25342d
z438ebc9b0fc4b41f387865b25eca0c1c664f5ee46d631b1a7b4d9f584843a2492f0e6a4375f36a
zd408f01e8d60caa0c7ece9914b89550d320296303dddb38ebdcb4c0e7f0efc8acda6e6b587210e
z71b5deece77038173722b7fc945257e2139de2f2dcbf3aadc1d4275bbdb85bcb926eb21d7915d3
zb4505e7608d3cacfd452b687a6788d931c6fee286ac5d74f5c9f498cc7bf8e2d6a6fa197c9f1be
zd7a9bd147265b94b25997659e046511eff70d0206dd77b5e79fb7e3597be5514c639de1d19ad0c
z05f2c3f18ba55f3e7c2c8f092141ffb4ee0f913cca02e0bb1f8f8095244c00ebe259e435dc1712
zdc483bff00a38f281dcf7256310edd6ad95ddbb1c63d82d04456f834dfce146c520a936516a50f
z29a39addeb72adaf9354cedd5aee8b848376fcf1e0930ff8e2955d5b97eac946abef96dfc634c0
z6d65c11e15339bff5a665cced0fff422a2050eb221291d0a204f573861634a82d46ebb13a2e7cd
z54a1d8766affe05b30f533b4430aa6b644138bada310d7e9324ed7ef40e05343d0133ff335b54f
zd0d1c9cf7af527f1fbc9ab345761975776946876b9996acf2b0a5dc1c7ef3a01b979d3c8335fd4
zcf1e2afa4711a10ea38eb5070315628df9f656a8facdea3cc8fd85bf05f0efba585907a683e2fb
z271f5adac55b7d0cbf1f923dc6d77da4ac065b2384eeb11fcbe4e9c4e286b3e0c8397c9338f4f0
zca5cb05d0221de519ac2cdbdf7c08e1a0d16dad14ae8e380d9909c159557fb377b8fce383efad4
z45ffde49c2a441c977ad7fa3d21d5968c4f3a81a3e92e97006f07e017bf15a9ce2ea866c3a1266
z726f8bb7dc1de780ca7405debe14b37ee80aba4e7b76374f984cadaaed3580ce6baa3b3cb72960
zbe04c1b7c04cff28aff46f7e3f9b9bcf091f352d657f97c0a6ebbaa0a3a3001ac19742a265e178
zaceed05f28ee4a98d5b7ca9524c364f47bf2ee066fa1c7b24bd3f92a37fc7bf54d05e1135d49b8
z5ae86802077f20b120dee2b5f8b0ebcfc182c8e312ccfeb7c5565e05e0d92e9b004e270557636c
z0eaa4af7fdf69fdd97f4e917e9286879d6a905abc5d3189863e716f36baee1e21373197d14934f
z200239586e40591852f3643e60624677f80b662e95948a9a41e900d5f6c23f565dfe90df61c04a
z0f7d290023a9543e70690da44322df955e5018cd25caedc3f54092054eeafeec2cc984c8520e86
z6145286c957ce85aa0acd996cf7e5d5af3357059038ffaf73fbca44d913ea5f60761be04bab3c9
z2478e767e0241bda4cee164052e43967c4534469f54063e9bca3b2811d694dc45ca7dbd9937e6a
z773c817a1b807133773e5db0d2f32e689321d06d57ed5a963dc83e3a30211b3cc8f052fc82629f
z119b3a5c9feea68b4363f0f5bfe3725d9c528b2e9ad558a81a9e43ba75ba67931311ed351921ae
z38cb0fda266ca34c98305f40d92421b393f8fe7658cc3684827c0197d88a62e7aea055ecba909d
z93f23d1cd6513ad88c54c83fe93b13bf48352a644055b0115da01c5ba6a14c482bf8d8fcd7b35b
zae4ca8396c69ebe6e229164108d506e0632556aedebc0256e06b028bf00dd9a70dce66c48acf25
zb5451026d6249962f13a15f4a1c215a4f24bd044fc1924dd04f5fc5a7a86b8fc01103fba9e9f17
z5a4b7d916bb85b5bcf91fe3f255906acdac8cb1860eb79ff5032983a578f89a934027ad5e4a03c
za0d64470b622084a0de73abe83adfb0d2e4b41cb5d929de63cf88e7175bc14aaf7bb3abcd35935
z92d1ff6e72e6a77c13b3b2934202d1dc5a371c42c2426645f2c5920af881ff7ca22c0e95d135de
z70c0a78b99b03829ea8edf2e441514347de79056a1b64d02529d6bb1119b515d321b58e739eb1c
z79e74828cf8e2a5379ed097e60e4259b854c2bf84f5af00eb38b920c2623885a57ae81182a602e
z78467b72725a4a106a09a53bd6cf4b69d7b3cea9406d35103b52319b1a26e2cf21b2c2b4321302
zf845a8dd882acc1edc800f7e3e8eb094e9ee738e95fd8fefdf7e58e0509aa6b95c4058c5056748
zc2d1d30f7defff1e4c88aea9dbf058bd92a8d2784050cb4bcb54b881566dfeef527d45154810f0
zcb6498ef5eb60dadd09047339b2bcf92f1b319cb663b708ce0229f187bdcf988c166ec3c72d3e2
ze7eba3d158c68f7fb02ed169d75bd2620e3ccaec149b03f6ed11d192671affcc6b40511bd2ffd3
zf2ee0900091e62d9cf1592b830f40ddbde28a928b1c483f6f9a52b9c3dab361e30aa7311606c36
z808e436d7e7a968e5756ee057eb22c8e2c00c96323a67e8a8e8a2204d5ee369edba6e62286add1
z3f485bfa08d555f9a0f19ae9ed796847f76ac09181af9bdc18835c13c5cad793bda219832ad956
zc64c22d20cf88fd9bb905083011610b8d2b97910ba9eb2c37a73f546e04cd872d3092e4b301bd9
z2b659e124e6144acb1d75c1f8c9a06b5254ecfd9ca898681b502ad6c28c3f39dad1e6afb8afded
z76bf60679879d0519fd3074134254c59eab676eafb0c7fae1713d07996eb58a73058ede0181190
z124b68b7adbaed52348dd24e48e74cf6441ff004f50abcb25b17ca3af2a45d6cf9e84bc3081e0e
za4112a64b02b2fc67026f7843271a401be3663a045f57f151cb528fb20be9986e68c771edf09bf
z1022ed17cef9197b82ec780f87eb2bd677db2efce79a61a6c8515fd25167cea226541494c26567
zad1b87cd50c89fe35f95db2fec6749426580ebc054ca76a8951a8d35339aa4038a1c7c45abe63d
z6dcd95286b0d8b597c2fe08020f10963a518110af9b3c553aed3e16fd6a04b3493ac25b4dc2870
zee37c992953bdc7a72aa3e164622f4f0b4e0398efbb7109010e02330d0b1a60ba5c32e8b6b29ac
zf148bf37d2b7bf29c7ad7a39bb3589f9adcc41b55080ecc05af85172e61abecc619cb7c2b04fba
zc4bbbe5e6eacb2452a3af7c9ac24c1a21b049b9a68cfc54282777f152a15a0b5a5e66a3272ae59
ze5f5af9af996426238d1e07ef601310d1cd94d3baf7985b5f4843ac075234eee28e5da50e880d4
z1110dc18be5e6393d83ea0fe5858db2deb4bb0022ecf4f56aaf0da9bde7a3762c29d27c4d5a78c
z123b51d2ba5ef358fc46c99a28426bd2d31b19ce236c8eb822a4ec0888440a259b70a0fb16213b
z16dafbbdaabdd02aa7aad0b44498772e72562b453dd7656da6a96a9012d4f82739fdca30c68ca6
zd41f02ed0df11ad470316fb34f8b347824293fc3d9c091152cc02d7153b3dc45cd35000917a18c
z2ee48018df46aa59ec64005a343f3c7258f4c22f49b07321dea4d966a6def7147212c2be0f192d
z9cbb75e1392e4ff063adde20aa3f8787b5ef9fa5cffb2b03e55b6929530a37936841ef7a2e2b9f
za9aee566c5eda2b48073d63c3411f0b958b53a8a1f8cecd1bede7c415bfeb4082e2e4464d9c7e9
z71091921b90309d175f21c2a3bbd6dc8b1fee922493ef8f80de2f2888ebc25fdef6deec7b7c349
z210568912611aed3f7aecb456cb0ed5ac4a91e37e5fda1b7dbfed3bc0b40f3d6f06c887a390154
z97eb62f77f6d61b54d7ae41b7778d7f204853fe8e089b83ea420f8d8186f1f5dddb4561b1ec303
zd34f256ac3e67ca9b76bddb7353decd2d13980997a3610e41e2343d52e10ab1866e7243a87057a
z6067dc75f1ce66680f746b930bf448c9b067bf8b915d47f4f9d3915a49b13c42df0fb142eaa64c
zd5eb26f2b05161a938241224413315425a11a1e90000379cefc46eeb83811860e6c26b8e7215bd
zb3c153f9abf9fbbeb7b4e3a64f3238c1e4c480a6b382d8f535190a65db1bb227114f4ec2acc78f
zbbb2f26c63950ff43a491374f1e50aa138c12a5ba0de4e79e8c9cea452e0a6ff8fdac33653b5e0
z9a61890192b0a1d79be66b34eeeed898ecee8ae09c53558c7615814ad05e07ba8cdfbd5f76d09a
z4ae6f9eef26c98e7620f765406fa2b9203ddaa699ff313de31b90ab37690582637ed24edca8892
z75935bfb701a14829943d7c9def07f2027d00504e94dc8e63111f3817570e9d53bf29be385364a
zd25c2d6a3f47f7d4db272c772d9bc4e5b0cef6653591e0bf7ce58e9038368334bbb9fbd1501fda
z29902451166f844e29bb1afd4a874dd24d0403db515092b7aca0cbe7dd4cc0c0b7c2a0e32704d8
z265959e14a780410aa2dfaefb8ecee689603cba3b9e4ac3ebeb367b3cbfdb7129e50f1d1b70ebe
z7c44f25c43541f318402480e85fc0a461b07cb8478d2d58a78e6777f230dd2e1ff9c31281f91dd
zdf33e3273170c55a158bd2b6bae28f967d842c4875f60b55fac99b344ced4d8029cfba8f1f510f
z57a8ae04ddd54a4f21a95625f6dc16ae84ac1ed8835b209248c2fc4f2d641f1fa92b9c76647147
zd0e0c9f50a76e80c69587cef3ac20388ec13c48bd66426c16f51be53dd951026f596e509bcaf81
z45376ab6b57bef4388584d75593f6d7b76765604cd33b84ecc75a6107442105959d26c1d75afd2
z04ee7722e11993477ed32f1adeb4634e71c6a727d8011f0646645ef790b3cc50dff75d2c7b5d9e
z1344eaadcbb6b53cdd909f4582d10c3190fbe896e7f96bacddbe727b843c91da3a2bd8b2b489d4
z085e754bd7ff8adaf468d43a1ffd4e9aebe4e000d27daf159b75d330e3bdb2aa2cf273d804f6a7
z03699704b57cc249afc1e0777f5fb103e86bff3ea3585690f59b567b4da8528a9ed4bce9009296
zd1dd61501352ec0e38cef6e615aeba7a3bf16cee00ccc2c2141b2c427ffe1736c80ba11aaea6d3
zed83bc0d59a175f3a45ea242d3b0ccc1f506082e0e4ea9e4ba9be6195599f99bd75a3e96245996
z2c08b0456805117fceafc0e8447341f538ffcddf5e4c6b733d74264f90cf56008b40b27c422760
z08c0e11fdf40a45a9fa0fae93dc665b1e2bb9bc634e33d33831add7b37bc2893d2b72566b85db1
z24df4192323e01630a2f48342e582ca1393d41f3828f7e8c242af0d4e73e29af11c47120f1e4af
ze33c79638cddc832e3a3396c9b04ed102428a1fac6b251ba0bf9812ccc00173054419f633e17cd
za70630f44df509d0a8abf1fb5d8345b1963a5e3e5ea724b16111385394fd9627431de8f1c7860d
z5c6348befcb92f787e1637cbe05c07aa94cc3b1b64b261f835c79a95320443b7548947a04f2b13
z9fa430cb0d9add36c80e6eb2d42d9329a64a8bddd420e151b0a8dfeeed0da7ff732de01adaca48
ze21dadc54188cecd27b5dd8b0fcf1057a6143bfba5ee161ad5df7190124e5402cc7efd620143ac
z188dca7ed4cde6c7c24d87540367cf0d60f0e6cd71461ed1bcfd6b90fee5c6eff6a86616b26900
z4e3a4c4015a9735cea73163250336b28ba2d9b6617e7e7d21bf17e4fd61468b75009dc58b426de
zc506a7f60d2e96634a42218e47a1ff0e9150506552fdca80d06339f73eaad878880c20a0caee3e
zf3144e8e01d8b3b75587260e212ebd4f6f2268f6bfb1e7992a96ee85f693896192c52e609b402f
z3c35a89a0727e38732b7300239a5cd8f74572d83e55d7d9a3d728f47006ebf2cd536d446a7f1dd
z34dca148622634590cd26ca648752026be81d4e7c64306105bd6d96c701aee661d98b57eebc3dc
z5a7fe4405ef50d9dd16ecd5340e1745a68dbfcdbd7b49bf789e82153cab8cab312a445465ae442
z55e44b3e783f1bbc292299fd4fb5506ad76c3ca91bd8adba034273bb4efd7cb7016da4b4186225
z183ec9f6e7f50d2fb0ab4142af9bbdc10f225b94991871cea3d2c7aaf09f2067441fdbabe5a867
z77fbff46d6d41d039d3253f666fc43b66a617302c50b8d80dc05cf5bd82767d5ca9077eb13e558
z55d55f811a85add921cf3a85c9ed4a417ee53f70338fa5865244c877362207184ccdeb3a38993c
zd50a823420296b3ee92b535ad545ed503aae57daf67393964c5b4800bda4643b6322a2bcb75b0d
z9c29faa6a36d39244c8759711bc77652c554a9de044f9c07b5a9de3f7c2df339b4d6983a8232be
z52970ba8338f6277bd0035fd3b69e11e329d21cc6b2e37c4d760361af76b2cb412b694f9601eea
zf6165193d623eb0de678fb82e4c57ec70f625806cd87d6b0bb2ea1dae5a13d3b256238fb7f9419
z3f4b22f1d86b774dc66284b7444a799ea5f4ce4b00b21de222764da8e3f371b6a1d443e0812416
z26a1a86ad46b422a1f2c8cf84b7be67146b7d5b9243cd8f3e04bcc998c43e9c30c6e98237df5e0
z74f04aede7b20ffa52630624e8810e7cfa969ff41ef162158cf4cf619468190abaa71ba0501e42
z56dfbbeee18227e1aca68bc39c47c6494eb220a02e90f76a6d8ac987ebcdac8fbd761ec89652ff
zcc35ff38e23f34461f1727600e090d6fd77f1211c5c6ab818bd91b02acd01a7d1f525e9fbfc859
z83fd30031f0b5cc79c5b078ea18a574af26e797793ea9990a3344f16f9e88c269ac4bd800ffbb7
z3be552fe07c6c9013178054e076d4e2693365b0bb8f5489f59fa64ac52c3d708feff53f9c4d996
z64248e25d4e32b60886821400f4ee79e6a3d52ba64e8d4f049260964c8c4a498ceb52c33b47cbc
z423bc82e45619fcdd285e582eff098b8b628dac13b7df917d77de73f23c928c15b44891ee18373
z648c87a337c13cca494b8c87d852992877f297802ef9dacb1edb5e03546cceef316b3129720841
z44e952c8dd0a43f81c8bf2ea24d820ce6129adc7902a7a4acdfe04ded5a5eb470f907f54463a69
z3aef401fc53cd85b7c751fa3e89a3e286115b59f5b39aafa6991d7eb0a4d01e31258b6403352d4
z18f9ced8c7e197ecca61afd631e97377b05dcab31a9510bca51e199cc50d3c9fff7a3c855b5a87
zcb9127a5b4a1f9a219ca8d7375fcb4e65ba5d61e4661b91f354df76fdee7b1bf7427bfe065aed2
z51faa8340377a6d7d75d3c5184fc8c832296f3e14824497368b5935fc702bb3655b39c18ad6114
z92101f6b0b3b67aa895abb9dce6224a0949c42b850e95eb9cc8861bee5cf4884a2411377cd2479
z2afb0179567f6f252a8365e75a55e68fa09dea8ccee7302273beabb5708a380e78e75b3f693a25
z9ad7c6173d7235f711b63f3b87d17518bf17b60865916baa168a007e52de485c810cac4b09fe60
zdbc09b63fae112eba6e64b98f00c5c0bf07d142ddff3846bdbe293aeb3d29e02b48b1bbeb94a05
z5cc86474c77499a3fa973a5b110b52af0f1969c5d18cd431527fb258019ff5b87e51bce7d6374d
z6fe0d44bace88b2f969b3da2d016e38fbf5516fe7a823e213c3c46fc41c2556163cc22c31515b4
zd82c7342b3cd694f1c3c099e934599a26c97c9488fdc16d0c53da228224d13da390b0cb8c35471
zfe5048f11b8347d11e4d697a7e4a7af8374f9e5562b33855e22edfda74b124d7bc6ffe71560907
za60cf9993396f8f0d81498259e87fa6e46b994c4a844c35063a19337b78bbdc8665daf58395430
z4e0fab03db965f84b9ccb300793c0f16f9167d8c3bab364ad4c8c1f2a1362e208780e6d8cad8c5
z277a3cc49f8a30da628f618781fd028b1d8f9eef57e7cd3e24a7fed29df41e47f08f2fad6ec8ba
zed70282468d930d3a4ca1b3e2ac01b6a264a2e837d204fd01539c8daa7c115833e84b9c55dd4f1
z965c97f2b7aa0a73e32e8dd2a547f6ad73abb3bc190183dbc250e0a284d2eb681fd94f391edf98
z1e31854fb6130d3a636191417e4075166865721af3e045b6385ab02039ea52d101470700704c4d
zfc6ddc0dfe3cded8f671a77b3342ddff6d850a7b6fb9f02a989fc12a909f5e0435a4d9e4d10160
zbc3feed85a761382409242a51ed0230ef8b12ff6fd31679d5d610c8effbb1a71387ffd8c1b7ecb
z59b11fcb16af49e7b85d991a7d55ac768e54a288639f467c1230a6ce0cd6ea3333bc2dd6305237
za2f18b43e35471d2458f8e4f192fae9a4a57c8327166530cb26e27c384a0955b06c088c7ebe049
zf60731e79008d2613b5c87e3a0891ff5376e7176361e7018c60bd8d380dfb879c054acbbf8fbd7
z85011a070e76b3eaca0f2459f818a1742941901bd8486f92c89cff1fc4432b041800297035e6c3
z104d60f6b8757580fa3ac01308c45124bbab89d1bce12dcf998e1049d86447c204b1d74f6396cb
z4b4c1ec1f45a571721c52dab7d11be96e2737c3109fb05fcca301001e2a4d1ecd391f4a225fde0
zf721cf46b88a9d82821eaccfb349b387b151c5b932f70e732909deb20c18d8b18179c2351cb37e
ze0f46c4969392f4d608cec5ea7b926e801238afb2e81f46d0d9f2a30b15e457f72f03c3041161e
z0d99be29f7b0ed1df01439a07868d345398100906ba77da96f09bff9c40c47fb7a48a5cd023aee
zb16fe0fc7720ebcb1b4e9fc7dd596a27fd47c317f3d2b06ab1153a854a9192b8a196232c84bc8c
zef4c6b56cc9b9b833d0419cda27597ceca403cd7dc555984377faef7c0492bbf55d93fa1ff3dd0
zc615ce907ff43370f9b67d2d34c9eb20424d1ea345ae8d1a12f8187c9af5a26c2ada2cc0418ebc
z587bdfa5915fd45303c1d921b7b6a34e0e974cd04367f48f9a4c3984fd84bdd33e82eceadfb839
zcec3f388c8415430ef5eaa02c49c25f7242b682f2c8f415bf135d01ba5f391dcd94b9df7b4016e
zbafdefd2812789cf60c23893311bf4e0cc90e9a0f9bed5bc1481a9e3e4b2fc4eb96079d37af38b
zb9d6459fbdd25756248519a4b2015e7277951fef5fe1813be86704a9d48fd1060f3e10246761da
z94ef5e3c202f5a25901b861a4de7a8a21de19d623b60bf9481adc9fe5a3637c4c45ee6ab532633
z59a35ef201bbc7edb81618d84792c6c64dd4f02a70832b7549b52888d0ba7cb2adf54f12cb7070
zde9a11941628d2650e95782686c019285af0b1aaad904be151d7bd11ce828bfd64c7aafc465a3e
z78f17224ae4d2f5e844b6deac050c922623f201fb7039a1911694336e5b8b8b540be9a5a96ed63
z3b3491fed45dccc7e18e0cfad6af3cb6e8993f1d3f4c6232e7d25c4edb0667340ace046c3c6bb2
zf541fe611351eba7092bf097079415e5cdf8b71d6db60c2ff10ff049a935055b175ecf6f9b3b5b
zc520bb663702b90bef4b8117cecab8ea9c70229ed9f42cdef34ba596fccbba7614f9edbc2a9f71
zc1d08b9c925c522dd9df89b1446fe0402f727df181d63d07a5c44765bb137618ab88db55947f0f
z304861570194144c57f72e5458410567d3207f2354682a389346a9085e8dff1e312120f7c67bb6
z1662782b7451ca4f8747a9b7e025c89c7df438e27d6df52ec17314c9c82605cfd9acd3aab073f5
z4f2e1d4b1bfac561bfe257fb8b88ef7f52627ffc37956e53305400c2f2088965260f8e52a994ce
z579d14ee53928a6682e490f90bb1ba2c4ac6c752c899142640be047537519132b0957f21dcdc0b
z215b5c29276f620028788c1cf0fe044b23bc06e69e834093f6158f1180f3e1c959419414f50f1d
z489736263c83601d762fb31428ee3ecabd87918d38fd0d9d472d161227c22e2e7eea88da2429da
zedbcb2cfcd4a0f0474962bbc6c4ff6c3dc738449dc532f8b10451faf10023261761bd7b34b9a44
z761c45cea0c0e539d8e514605c254b59fb06a3f8e2a1e324229a77e4f1ea8acbd438d19d383f01
z5b6158268e3bc6a7f259b6fec0fe6293bc3cfeb3ef5fe36e91e0dcb69c11a3836485b3ef082ec8
z942996a462555918a1b908e02c7899406b68de88a71b01c47606a9d2ea77bde5e0d6c4972e546b
z7fd59e31e84ab46a6daca6f8d2d0fe848d59eabe88103b826f78ff28c127d11bdd94b707fbf131
zb9cabac7e5a64152e39484d6fe9f12ce52f2fb1f1fa34d934aab8c38be45f9b6a30e90447708fa
zb020f9492d0ce3c16bc6a3db055bbef91a7cf3b9e10468cd07420a3a0c62d67f0456cf759f626a
z6ca934eb9b27287fbd649371b157f8a9853622ecf01af75dc70b6712160d9a3b38fe94e8262392
z8dec0322d2922d9f543298db4c62f2c76e644f462b5a0f12ab03b744e1c1e7f7c20f7e249ad251
z2d6355d5ab1f51f041415004b5baf77322971c049b8cd3595ab5e38747a4d40abe7428c6c49f51
zc39577bfe732b8791f9f3ab32c8abc6a6fd517248bb62829eea72b3cdd143536c339014a3be938
z060933c87d476c2cc7ff561d8af64dcde70b7f1203feea139960db8f12408947696f8298471474
zaeff49c675c9623cbbd331d8240b50ac398e45f761ebfc17dd2505007be6bc3b8dec51346f69b9
z17b59c11bfa21f146c25bfcf33450352439f819c202e36d4bb437021879389d584b176586f5f5e
za8bfbc1944ebfec769607d4b3cfb6c200cff954287f78fd40e2fb331b3195cdba953e9f156b05a
ze6b45665d6ca19318e0686ab1a506b37ed805cd58e91325d316f670ebb88945e34ccd841789c2d
z2b601ecda721f05fc12d6460ab30099ce8373a2fb48659f4f2e68413656fa438953f59671f04cd
zac47417d1a9b51e3f6becbd35d9b7186f3dd8c75286cf4370147d446e2528b8e45e3ddbd15362b
z5413ba98dde78941943037cc895499b16fe5fde319965b5dba0bc95424cf471fcde8526b7d8fd8
zd8a025518c67bb1cbb385a71b604fa8274d342c25107ad0aab1880d4702570ba0b181766d0c302
za4c365a2d01013a598d65346701982d5751935cdae2352ea9907d7a49a4f4873838d8e38d4be99
z087b621ae2859b24017fd79f26f37c69683de9fa667ad7413d9fe39b0318e5746189b440684be3
ze1506422ce96ba10ced825ed169eea78e3a2c0a0902a169416316b1157fc83b42604271ba97c07
z6c313cffdb3a718c871c4eb7fac9e3368deec6c20bd40edad65c6bc1ff64db6a30df28cc187369
z4732fc4f13ff10deaffd26dca3620a040f26e19d42aefcce75b553f7b35c036a0d6fcef50de7dd
zb741a46f21b5c7cdec96d2b50d4a635ba0b7d917542c0d2d5fa68750a388254933e7fab1f1623c
z540d1538439c3d9aedae1b795325e5bb44ce3d5231579acc2eb7c438ac1efa15127ee36ebccccb
z00dd20bcf8d6165e949c74ef24ad916f7a8577849ec1c490862ea9b12354f0ff690a224c895421
zd8e79b200ee4881266c3e54d25f032ebd0216db96aa341db9126a7cef1aa2fa12d15710ef226bd
z0ea3a4d2643e512f7b86f7d814097b9d80c82bd331e348ce2d10ae2c7e3f3782b8839a58f8f0ff
zf022ab9d5f81623adb19f1fe077755c10c9801f0ce9d14bf7240b27e1905056b72bc80babbeda4
z2b198b5e502718a2ff3b8655a8001b163f55e5479326b0b851cd94e433498152ea234577723f7e
zea6bca1c90f90b9e8b1d51d83be50c79fd62465e19149746bd984e3816bf8a448bba82fa2e8829
z12b760f5c48c72550d0092eaca0923606fc0ca3d533a3d1f65ffb3ad7e5b134b53807375219cca
zfeaa84e967cf15adae2aafd22e0456b72c7795e99f5eac3de95618296401ab6dc77ee56a2443aa
z830a633a10452ef67417175f8a7b8f26430bc3e189457620f9e1606074aa68b2316210846c1362
z0fc38f613c54d048adfc1b1b46ea361a86dfa4874ca76a45b5cd9708397522ec73f8fec994a1dd
z17aa4fd316befa1de5acd0ab0a7cc0ad38f13dc23737dabf1403b91c9d631f955dc9da75925c0e
z13de6097b584b35510efeea6ab4c390828177f128ac5a835a7267b01bc8c5d0a76a715943c6865
zd07d4c4b32598b6b74ee34c0cbc2ebbe8639ccd969016146a881aac82df3446226c8de87519b7c
zcefecca01d10ddf4e24ca4411a4b6a4c901a74f67c369a3bd185ceeb11fdc1097e7e10f909127d
zaf225d75035b4275bb0e063a490a9d689c0d82dc34c783a52c96d058827f8404734097cf05930c
zf611220eb26df524fbbdbee89dbcb50e7c6d0f51ea86b88a7c6fdf7387edfffe40c86568b8c475
z69a2adf866646eafa96ad5e9846366480f99dfa6d74ff28da4dc5f1aae7c54639d93803d6bb226
z669650e1ca6eac2fd3cd4ac526f9df4b236fb11c63a1d5193af023166bf56e85b83b25ece20728
zc5e04d284fb9e1b96004b8efa9bc97ac6e91d2e1d6169d7a91d68ec7b23733a9819203b270cbcc
z23f11211923c38afb3738216eaeef627b984c7e3afc2cece923add8f8dd9ab2b76387e1bf76f15
zb62e10fdd0f20028700eb86f1ce96532b33376f041e9fef9c2e3c9c0613e753de3770d26cde0f5
z07125f6eb19ac77ee3d5f916b5896916b4f10bbd5eb64565bcda1fbce586448f8696f3689d6aa3
z67d9c59478aee328f704a215fc0c347f3fef7465f9a8d64b14312defe2e3240003c8bc25bd4e26
z8f66628b219dd9dba0abfe1f4dee5597f5f49f70ef18eb1ee9dc26e79f9fbc9192dc351d8e017d
zc43664b44f46c3446b3ab47b7524547843ecce26810ffb75f7e7e6b3d6f8cebc477b7c4b960e1a
zf2cef63aec10ba9699be049068df6211e4806cff6521ca9b10540b647a825244bd1dadd95c2180
z307d18985d5d143ae31f5f94ad9e45534de89b0c31a81be79cb77b0d354e2c10d4905117858614
z5961fe3893c86a66b6015a34407aaae9b4cd1695440f6e03ca579f064dc553b3a719808267a2f4
z63f7afeb77a907d5e74d72a8c53e435360ebe9cea06e9c30766ea1df92e128d6d6582f7e3de873
z10941a31bd47d3cba3745f21ad05b0a18f9329effd6b82f620e0b45b38ae9209c01508d9114cdf
z3f16b6bd16c4e5c31db35a4a
`end_protected_0in
`else
`ifdef MODEL_TECH
`include "qvl_i2c_master_slave_monitor.mti.svp"
`endif // MODEL_TECH
`endif // encrypted_0in
