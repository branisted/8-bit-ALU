`ifdef encrypted_0in
`protected_0in
ze74c34e226135848fe16db9ffd31815111b6d7fb642c521a3f628cf6da949865580b22efd062a7
ze90adae0e65e66a2c36a587d0a790699161455169ed55a01f2084f11770a774ec4c588039b380f
z6de9c5084882a40b79a175f5c2114b2b6d78b070cb806e1c0aa9258297f4687ab308bc470f0040
zb0b1de382961eeeaf2e279e1462520fc31c119af8f2b214846f56c2b3cd2eadbe4099496abff18
z15cec83ec4a77b868344aa20ba7360908f5c0de2a79abf8b3534b883bb12180f68b5d4beb444cf
z3fba8f13afb0abfe8fcc4294810f75afe452434d2d0f1166236c82f76edf1e12979f04bc35693e
z32ae028996dd85737a8f5adc1ebb94f39c940246e887647b64782cd7ab429b0544c173176cede7
z01dfb26b1f73408344a52b7e1f117f12bb9c8077b34876c2e6fdc085981637012dc9754765e1a9
zc512ce062e0b8fb16a214591f5c81e1353b900a611fe1f4886b57940b41b7f2ce99a7b84b04b90
z916f717e73bd10589c81e207ed77ec660a8cbed5b487fa50acde1b055c8870bd8676023f21ddcf
z9c98cc47cfa2d654ff1365d1f45035a045a66c5dfa827905026201628cee5aae21fb892db766c4
zb5b1406e11aebfd6dfacc9da5ec03b70c276807a3eb15e28ec7ab1dddec42388b9424ea285623a
z248195c9f894b36317ca6e59c86f11031163f5f52d70922c037057ec3eba50b955600900b32628
zb2250f2b4fb3ed6db7d81b8ca05e994209e236669db511df2c321dadeee74880d12dbd5092819e
z312f2e640fed00f965c7b0e1d2007d987dd08e1042332719768f689f95a8ecae54578598cd4014
zf52c9aa29e5602a0a7c0b59ee67317c72101e7d1c45c07570c0683c158486b6e3157427e0a2514
za97901c629a01f6fd65b5a7f6f7538b7ab683549194b5767ec9f9eb38f388669f93633863ba210
zd15b4f9d05bd96c35341c02c93752c2344db76edf8c697562b3a09dd9e6ea71115a107694a03bd
z48c4beb95a5fdace643d8acd8693678fb3c10dbc716d343185d0f8c8b090128427948cc61f654b
zd79e08af23d1f841dbaa5dc1936e4660e1f04efc36d203629f18a16a4829e3b3126751fa196d42
zfab93a2769d0d4af5366799eff9987e0ad2be0898f05a8a7fe7be72a09e6e962114c35e028f985
zb4f3db4d71c39b999c96003b9bf32fb342a15fac3c4446676fc11b463a9620113254265646ecae
z71d7cf3381b7e84b560f223855b0b20038eec96c1ac4f1af8cb0110cfe327c79fcdd2413920852
z093eec9cf19ae3cd8a67022d07fcd7bc14320c1ce4d9db0e528514c98a62b5d3ec31605cf03599
z4d6eb850c37fec85cf69e6b474e171d53ee2bef5d245d9cea5c101e34ebfcfa73468705933e98b
z1a22aa5b32d9f8d3412392ed7416ae93ef2762a663e61a210309cb52001dcd4a952d8799718756
z65c1db60a4531864be9bdeff4cefb56beffe2bf29fc5f3345b63d7f8ab90e88a20287661fd01eb
z5e716c090119d5d4c08ccdcf8d33e906a8990d677657f34d4716cdbd43f372c20c4a03b754b7fc
zd09a688dec478294aa8052d341050720e84add185bba28dced0c27c13f7c8c7cf2b793b02369da
z080bf6eff0124e7ffd1e395669b8e0fab00d0bfbdb7b4de8907980f17ccc6a990eab828e203546
zc08cabef41d95483de759263a68379bc58694349f4d092ce1c8cbc4d8b1cf9a2a993a7ff3c5dcc
z09f2675b286e7c0bdacfc3510345f25f7fb48b7e6c7f9ce1da3d69c5c34d4db08c56127a25342d
z438ebc9b0fc4b41f387865b25eca0c1c664f5ee46d631b1a7b4d9f584843a2492f0e6a4375f36a
zd408f01e8d60caa0c7ece9914b89550d320296303dddb38ebdcb4c0e7f0efc8acda6e6b587210e
z71b5deece77038173722b7fc945257e2139de2f2dcbf3aadc1d4275bbdb85bcb926eb21d7915d3
zb4505e7608d3cacfd452b687a6788d931c6fee286ac5d74f5c9f498cc7bf8e2d6a6fa197c9f1be
zd7a9bd147265b94b25997659e046511eff70d0206dd77b5e79fb7e3521c625825d366b240ee3cc
z55eb4609f9aaac5b0f544b0400020fa20f60ea949ce57136f63231807fad6b3ec20591df6f53e1
z87419d4876035d5b47351abc12e769ab8c52aadcdaf5fee645d7dbe84fabed8a917c88f52cb6be
z7e32506f4df5d16910c17836c6e7401770a7d1337e9573032aad645596b96cd586552a8f604587
zdb653604c7fb84b5961c903bf5f76522a40967063331973f5017e3820bc9771457ca617c85164d
z263851c212e539ad9ad32cb50cfc9c813a5e4043dd2ce54a6dc0aa362495aa43a33b9173d21858
z9c9eda72c043cb161eef2ebadf1525617f57219e20f032f938952364d0e3e6309e4be068f0b217
z65606a400879f2c8bac7ebe38d49e4b7fcb0a47e9dc4a2f77401d3300e18f4cc5ac579144704a1
z77f50814edb7d5f533fa1d1df4357925054204870c5f9e12ac4cb548552ad08961233a41f4b179
z7cc5d4a1333ef00b15fc630dac72275b01735e165fc6b13822e7dcaa810f5764a42e9e0a8d6e8f
z3ea6c9d90efb6e52081823659f4838b274011a0714b229552e4ad2cbb3d47d19f97ce3248d7fa4
zdf8330e451f9191f2092acce260831970cd7c6a66e6f27be525199aeb69556617199b1d63e63fa
z0c2602f6f1c5532fac31c230c2be0cd3f8e172ec401764777294052e623b3a4c3b3e8d4869e264
z9897f469ade7a97b3782bec2c800a25368d7d56e9236eaa231b128c5f666f649eefd977122c20a
zedc12ac6b7ba80b9b0d060bbcb78198347111222d64449db1a78294280578388ac98d2a76af9c0
z99e1aedfe677133bfaf6ffd0c109187d83907c46aa2ec02ae36dfb6eefbbe3688d3d2b86139290
z6158ce6051a1de2986256eb6844a0b60faf3d5bf2d7db5d16cb9a61ba713a5112f675dafc946e8
z6e2cb0ffc9574220d4dd38d57f23e3fb854c932288f2ed3f584047a1c28fc03e1cf65178aa71bd
z3619afb90be825e617520869b909f38b3210c694c2c60fb5c5ba696bd77421bc1e3a3a13da1654
zcbdd544b3303eca19f5f36da4025c3b0d18d9cedf6c0f8c4db73d650bcc1874a1b9d763fd37e90
z6a8ceefab30f6a9fb35c580c6aa394081d4c0cabb4a8fb37d55c417a1e8924f5e136796f518b23
z2982157662ba441692ac7a9f3a6687b6be863e14cadfc61bb0eea857a98f63973428dccda375b0
zc0773541c01df881bb679aa15d7f0b950e6b46d920c92fbf0eeb72e7090c1a6b69bcb975af2d61
z340ef23214f1f40f32af443481fab69f3ddfacdf4e57a0dd02419c8829d98c267c8090557cca6c
z5adee60b7d6b2a0bcf3154ecba921851ff32f6e6335d3c6ba4aecd8762d52db1b19fe6373e33cc
z991dc17485ea3ebcfab7f03e21d42d3794a725c150022e72f45b460e118f986a0b9572c774f142
z1e6078aacb4748ae4cb865da580f67ed6d1e5e9c69983b14b7542877180e23f50159998250bac3
zddcd6c20d41ccfc8bab3890e6f0328083a1cedc6587dfd6a1b6e40fb4dfd874e4c0986d1be43d1
z9c82bbe386442c05d5f1160e0cdf128928c013232aaedc6c7d86e838dd7df8b563dfa10da32a55
zc5de7467c14baf4a8afe77f3e50af5f978f3f8dea65f4bfc66dbe8f4d924438d3c1e5d3649af71
z52d23f3f911e3818d322faaad1ff4a58e3c6950a13dfd6677561966c8a6bf8f05df302560407cd
zca25b550f8ec905f82119f053b16bc79adbc0f21fe742bca09230e2d11ad62566a73b2521781ff
z8b512ae44def6a019b7979731be529307970a1d3843ea3374c7136264d37852ef88785af9c2899
z48af819069110163f729bca057680ce1dc426bf7ebefb89551a622d6eb274fe77fbf4bfcf6e5ea
z0c0316c32366aacc7407bb413700e59c5497aec8e4d51981eaa4d4c6825af8bf8602999485e474
za5d07fa03ef422cc3ff32add7b753ed0ba8a250e462c0c9e17b6b01aff92238bec5bf342ca1387
z185da7a7dafad9f8b48b6ca37638f646a0a927a514452b441ba3f644896c9409d131b0129efe9e
z4e22a6745df344fa74c179c2b61b247f6b2b06e021f77576608a3c9cfa2a8ba2cd538b5226990d
z294e30e678711ce079679bd14f3b4ba655b806083eb072c41e1ae09f8d8ae17df67ff0572c8dd4
zce2ad646f2664d5db8c667def7d88d52074e830f453950a3b663b3b35cdf6d82f0d4f13e8ee2cd
z437a20bc774d52c01a1a4ad72048648238f510ce55763bcdf51c1c33d846ae285908484db87ea9
z5d3997a5b0d3af4b84434ab3d6238826847b557cf8b065096c42090c01d800bb62ebc919b469b4
za539c604aad7fabb9a6039bccf1901faff9cd755c719403968dfdb982632171923ac5b13902ba8
zc4319abea2c0347f9a4ec5e8c93d4d93efbac6af183c1b1b9e9d64cfc9ae7a0a981a7f4b2e1a9d
z2952fdb7c8e4508bd6a6d5ec983ca786da55bb40aa2e5402ee51f20287ebc00de8732cdc877d92
z5bfc10c1eac3df3eb797de281abd99596151264b9ce8aedf03dae001abf7f38f85513d3ef48a76
z81f9f78883077a2aa3242a58a862ffd5246f2335d9046b11b480563e2333115ce4a9eab629c41b
z24d3964a12680e66bab0d1348e98aeae1ab6fb20754732c3dd3b62683bede3371803df34d3c0e9
z0cf7ab4077670090adabe3bf7d75a4218271aed4c61ea595c9e577279aea9442e81bdb0a0f04a7
zf1b9cd65332b923c073efe36d0f27f98c553194372849f498d792642449a662f37fd68cc42ffab
ze16fbf1b939cf1ad47590406269e5d6397ad07243ab43563f27890d9edf85487e9cf8a95a764cc
z33f917eea1166365ddbb92f329bb2478aa8233fef3b688a29a4b10d84bffda5fc378f61d2e9c37
z62d3037e9ffccbee8ea2c873d40d3d1a0455415b1fd99bced883ba07f1dd8e9e1573e7cdd1482e
z13a2347e5a5cc7a39fe709f3143093a4c80dcb2e6476b67025cb093ae43441851f1c8a43c2c66d
z6b06bcbbd34b95c715d51c73921e25b6ee8599c88d0ef64a6182c11159d1a97bd47069b58595c6
ze9f4751c73c9964457a23ca2c93f3aaab8c108ff8f2306be229cb99f4017068e6d84a981e0989b
z0989a6ed7da49629ed4c9884fa83684fe803bf6bdb92bd9752a3ae900eda200d2fdc8ed181055f
zc9a1712380e67ba05a8f293104eabf96267e13b9fed4ea281fbce5daf533a109aed3bc887bb3a5
z8d9a2d4ff72aae6cfec76efd4b8bce830e747e5c6aea28fcaf91fe4be054f3031b9c617ceda307
z5f06aa7e48a3f4b9dbb5bda8c8a8b116d95311bbb25e6a1d5a936c79cf973433dd3f87b034cacc
z55967dc692c290c1b660a496b7356b65a45eb44b12f4737696133eb862e56594d9ade7ab63b77f
zd3091c691d67a188862147b5383905fbaf71d12b72bb878de46618f9da52c6b743133211d9338f
zf271dd8e940ac2c07e20c8bb0152a14c8657f356474ee5d9e97ec2d13c6414bd1b611f338f200b
z7658787a86e1b754f07d7fe0829beb7beb0be7a5d1554975c8f41fccfe5b969b044d57c51c7d02
z4b0bb14b87a62d031db6b4df75cb180a6c621468f4c11314184ae89fdc4a4cfda466816f9fd514
ze6f092077ad922f558ca61e212bf2c5ffc7769c75953d5c49b391a6eff29567569035366404bf3
z372dc353a441411cc0e724453c898a650a5fb402e2522be4a42eb6eaa15e993c465dd1eb5a2190
zd78e6044eb0b8d6cb351d555836a43de27f790ad6c314b7015602cd1626ddc8cef8b4f1b48131d
zd067a35c74bef6976f21f08d7dfc320303e2f7590a96f2b3a3076c8f621a66572aafca44081bb4
z0928b1817b975c3c6a57f6704984cee3eab720cfe80d808f0c3c93856881c77cf0e7a48519a476
zcd91708e7726402be52bdb7d5e1e1b06dfedb7a65fa4d0daf16db711c722ea34b9fc4a28ecb964
z8ab59290955ea8edab2301a16f8256d47c1efa59d9c4aa17437a2bfc379d043ec105da5c1f4ca5
z805e2cdf3dc58aedc2de2c41986b76e7e1cf123e9b3a89e8308933dc162860cec2350c6a0a4cd9
z09d340323a6e158e3a292719d67f8986a0b6ab7aad015008fa356d1f1e3cd51fafc196b63b9b13
z6f188fb34239a83709fc7a089456ca880916dffc060585c0fb1471be05c6af2e25095546d60a26
z2675d0dcaafba065712e330ffc5c8e3fe861d9699cc3d7a4ac96292507df704d491e4316087c88
z9567c964779aa20e5cd32b1068e73c285fc3e3e220e6b05b50eff88b19f4aebc3a06faf96e3c02
z9c599c6cd0d9b2efd11b829185d54fbf47de59820bf6ddfe4312c6d710032ae67b2e382576c68d
z5d89ff91f7f032f238239325b77adc6473fc96186db4dcb28512a7f8f5c9f5c753f5a2acf23e54
z3746735a0dc06984ce679ad8b020d79b2e3e74d8ed4af2c8997d7f5501a7a9bfb99f99d196b31e
z6f5ae639f8c6577a3b155edd3e89f3387e7ec46125d14b51cdda05a56140e13873f87482e54c00
z0969589e11a0830e32fd5be14b62e1922a600f660502e37d26fde072ec968eae625e94999cc089
z3497edb4f2aff9788107103837a7079084a8392561cf3b5da39d914eeddc614c08ef50b7c9c3d9
z521e1d3886d4a7bcba6519230a7e7a30fb088dca8c0d794c7b5c00ca7791117912ad5069537508
z2107c4f8e92eed5e81aded4943ecf3bca6e5cca18b872004dcc0e3bc3bee007022aa0720c45411
z25dfa1fb79ec4fb96c55a4fb5aa5605a0583acaeab449158db03d38818549c130a400efeea8506
zbd6cb2e88560d5ecbe1f01ad3d1ef36ef60ef695c8f735c1919cfc5e66d2e7a620124bfd43874c
z201fa7d3013a7724720cfc69bc02acd8d8e86cc7ae79f3e835fa2c1cb21ada9a178708ac6a9dd2
zf26d643ee3f5a5183586735d34ae25fc5dfd00ba1f85e78758ed5b8aa24e3c4c684fc0ca7be354
za4267160b4d5664d5188bc0d91a3f3df16bbef0b9f35bf23cbbd599b834712e78ff2ddd4fabe98
zab136f041389f55b01a76a6444004b1131a89d0b70c027327db4b9cf655be33c7f6f326d787139
z0f3bfb43bfa8b2d517513ef6f43fe88075cf4e55e151f2ee6dae636e7d13a9f9318d9b109e815c
z4c7f7e7b9f7a1d8272ac1039b2f0f00a1e0875a8b1cf944ebfcf21d3a558d193c91a8e12d787f9
z4ede103ffc883dab551a3bc210f1127026199886fa176de945d22ca0b1f1809ab2e5654bd6dd17
z911672635dc721eef81a046bdc5a38d7726d17fdfe565245333840d5ea793082b408f120036a87
z12217a8e051222b073fa607c3c7090f112a110ff514fd31175857ad7e8490308463a1c65d45ef0
z5aec974d3433ab5ace77b8df37e89adb2af9158362cc18703c2d1839f6fcd22c55a89430e3ff65
z911906eb0838b43b0ea6de567e5755154da3fc2152565519e48d2f6e34fd311fcf705f5329213c
zddf0ced5ea48b28a669d54317e2467884f83d20dba5a94355fd77be222f0ac1880b2fa0cb0109f
zb615d0e90310a3972ccf2e041d8d37727e9f62c7f8a620ccff39e5df59d30dab7e587cc1453bb4
z4a23d64f87b8d41816d660fca172163ff458f28d333b125de1e608e917eb20e70d00ccda342a85
z8a6616e2947f8bef39da22a36e65d545bd6d95fe61b47539008dcf6737bdf86e5f968e2efcc901
z602947e030f86956344cd9d1e2f0436708cb67b1bd3f7c0a21717399f3bfef2cce31ab8fe770af
z38514e51496aa7de8a6529fab7ea2b27e04d10baade8af97fb84f72f58d8adbf9c1f1a9d057c9f
zb08a671a6284c60454238acbaf729714567c20f034b47516f06e6694c0d12b4252461a394a9354
z870e5075f8ced94da079aa9563b01c2fb9be24b7d2f3fc57d299aebc0aa740bad7c5b77184f750
z3dcce7547c9600c7fe8154783862bb3d9273e2e2fc5c1c6c2e55035926335bbefccbe87af699c2
ze375e35ed49e4e713f7c6c052adf5686249fab836fcfa254bc473dc63c53602f390f324e14d0ed
z3d3b02b905adf2a00a2d4ad95aad9e81d42ace1efe8e2382bbf4fbb067fe5fa4ef878a0c7017f5
zf6f3e50f888ac684477b0cb50fadc7567667b8af36ecbf80c3ab3a0366265a3861b96b6bab9b00
z9e0653cedd7086384e4f9f6a3314a866b4b9772a0334993402a005fdd335a467de6e044026486c
z77573c0a9cc94ef2e9eac75ce590428a918b972e31cf3d7c1c01fb0f7f705e33d59b9aa63b2037
z71d393bf97a6e177755172476d026db457b6e5a2a84f30d4af0e6b5b5954a3c81c5b94a34d263a
z0a7c2007b4a189a2f460176ac92e95e0e852d3096c05df08c048b8c49712e6b8380369b8f4de9f
zb8b5a3c2c4c7c8f2f97692f5a21998bd7b1177e01aeaa48da1194961f8315d843d96b44b625e1a
ze02b87c43e16675a6a7edcd1c883d00349060d9ae7e464e1fcb7a13fe90cef987b43ae281ef5b7
ze22f4b8021ec59bb9a7d227f591bba2ee6863c92b15533bfcdd0e5733de72cf621e715d3246ee1
zd8a61a2f76a0a17d4fe3b0e248a42a954e6503655806d70ffa0b9bc168dcb993e76594e832d6e7
zec9aa7eb6794e1666230e41710a665d980365656259653acc140e24fe339b7fdbbfdb721a08ba7
z68f93cb692af278b31b98ce5592e35b2f3ede50a4243258891ad1e2731d8b6063061e34facae6b
ze56d455be6f234624026b0b3e7249862650b35a36313e85127cbf57e059d1a3c99f367a8863324
z8e6a20d0926d03c53fd17fb578356b97f3f40ce6c05c2b56cfb422e48db76f0692d0b9224d2e38
z7b367536cb37051e55126ff23c7685bb50654ad947dbc83e25f6147496f13e8736174b9c860209
z30d66f3a3a7e55f8301853239774c9eecb547dfd3bb6d023c1978ed2b4bb1cd3f4756e36cc3914
zaa2112051fdf71d032ffb6f7692103565fa62890e08f9a8738a045cb3454a1f6993e2e969d08a4
zc1561ff34efad5fad0bd6c1fdd15d4f5142fe16d78a376fad8b5b5a353f0b7e0210c3064bb9a1b
z1eea1780ffde0361f98103d543004ee5c9d7f00208474b94de22b5723da85d7f68bf2043dbcb2d
z8062afa6dc3536ced6773701a8e0ed8bbfc5f320bea679aa7e7a0b72f14dd663c8bb0c3308915b
z803f0a6b1ac86beafdeb28727b564cc80ce5aa084e448972defd928c90b161a273a80ff1d05694
zc7df253b9f5b69dedc9a95a3f71a121c2a8db73730fe04bb8379bd56a8c1f229cff44a0ab314ab
z562b0d352be87423bb8e0cfe1d955723a68590046e7f7514ccf17bd29a39ee68ddf8f797ea52c7
z22903b3aa8e10b1ff65c9169945a6f8f0a79ee9277f5ea38adea7a6bd4340ec08e690140c0f777
z117e20c508ca07a798b9a7e04f50545c5a0ae2e8a43066ca71e4b2ee8ed845ad3fd27ad95d5f18
zac235e24b2b03584131e9c56514184bbf921f3d3b4dfdbca32533ed2d2bbf40fa620df80b15db5
z2a2c35b625d12f098214f790e74ac58fbfbcc7f84ca3df4714cc50318562a99896d01a701c1851
zeea10891a90ccf708261b6d27220833cbd0972abe4287f3175ac1785ecbd225f443486dd941258
z2634377b46543c3a010961d79facaf7a9eb4f96dc4dff8b42215e7c6450cc3eb203310b5cb09cf
zb614fc384b86f4ff3a71ceda051d7fc34a731da0cc63d996bc1b81d239222200814f193d8aab82
z18664b7258e5e2206c0a6eb89f3c9b001df023fd30c4d8488f8f05e2eddf23837d1584fa607f76
za721003fd9ceb34d818a65b22a23a88ad6db1a1a97c03ef1377057907e8635c7dfb692c40a76b7
z97f8712760b7d9c9d05a253e6634f6c95df4b430c471b8c94f26f08d114bf54d63a0dabb8932a9
zf9a6c7916c262e1afacfd7342de14bddf15ce1bf8e4bfe72e1bd7cfa42cdfd2281bd37c6a7b6fe
z449267af71e2876fa0cfb8a13426beadd03c7fa70391d4413b5923dc0be741677badf935c2553b
z91622d50bd14fdf9c3b47568225a8cc7e13644c9d568a9eb78008d588d5ee40394f0f0cc369ed8
z82e26d9af56af462d99673343250b73c543796cf041b5e0193b795952f49c39867ce4345693002
z5ce6c84a576ebe263719d7f2a1be6735e41ba2041778764ebcf906dbf6bf6634ee52aec3a279f7
z23b22df95d2c5a99aff7cb63c3df0632fdba10ab424121af23a2f9dad9c2d242661d1e34c6e554
z7fa6f6c49b37131e0cf7f6d4c1f60031e6cff528be88a76ac60b0e66f743dec3e4f48ea713c6d6
z683494b8fdd6cc58a0fe8e55ed3babce35bd8387f40d58f8c80b125500378ea2f4a41f9352eb54
z0e9c03ee4727717c1a5421f70c45e334998a6680e03128a1c365d7e466eef2b4e4c17995873f7e
z4738dfab69e3a0954b6e71ca2e528d6d4ac7671306b5f2360ab16528c56905ad2ce8341e5b6b23
z82cb0e45816d1d9670af2fd4a81b5e1d68c3f4740d06621dcd91054c916d9a93fd4016b05711aa
zde17ef5c654646e8aeeb2574154d189d3ec3c668e00086e081b1ff26429fa35eafefe216e57db2
z60ffce3c47db47adca3b0cf70a6e75258c8455ae51e9d30617caace7b422f1216ca2a7cff4ca8b
z0487c02fb0699dcf1bb2adca6e59189a09a1d41ccb7b9149a0ea4b969c552aad61904937fbb23c
z0547c13544d3fd3b02c0218c4617f54e77808d5d6d6decff6a231fabb6779942b41a99e16bc8ae
z96c161a3cd7171214c5caf0b4cc5e0fc955cfa58eed8e196460998779944da3c0cf76dcb0aea99
zabc59198eae48a6c0060a1f2da8f631caea997c0cb7cf06535a4c684f4e2c3f258e50f95a933b7
zea1dc80bbddf7db1180000ecabb0ed589249984ca30203ecf206a0080ea179e52fb0a9033032a7
za2a28c6bbee718f4431db9b8de39a55c4be0eb7a4c691fca66862c561ef99e3fab9c15758f4ae4
zdbec5b6879ca0827358b33c86d55d56f89d23f181e51855d034855423032ec1c90f7233305058c
z6c8e67aefffc4e2b9396d8e02fa7e3577c534c52a750263855401e6c05348a65e33b476edc0add
z538e3fac100d2f659a117a16bc31d1be0f203993c2ff3bf3bef71effb974617e498a889cbf583d
za7248dbc41424df92cd0bb9152923717397491bee43d25c14a150bab80e8c610dc2f98e9ea9a63
zedbb3994fcc1fd1a5850354c326ed018b174cd02c9166d1c1fcba28ced2a815df6c02907754d5e
z57e023d6e6395b3330e69c1a0f4f45cedd559f623b7345f8c59a06850329f8d5fb7ee6dabf3968
z264bac73fb12ffb5fc018f32db6686db116d0ee38feb6a2a845a817e138bcd3ef51bf966f986eb
z6a87383e87920cfb7265fe165ab4fb2d0ec72f85b6386a3c3d211818fa559eda458774d3dc4930
z21369145ae9c89e60ba1abb15aba4492e1cd9e955aacaa830890c9c4a4748f663f454f9d3838fa
z9a43a9d0cf30123018ea188e00e5ea5c2cab37b02a79da5d49604a28228f628687641f9dd6a53f
z54fd685418c97658a4ce013314af56051b0aec63a4cc32084b9fd59790797769421a364404b2e4
z3aa4416991b20f470fcf508daa11caa7b7476952d8d04006a34ca14770edc7c91d1def9c712d9b
z2e2695033a7915e4089cf75b51c4b8e3f8ec643315a02fdc34748b943476eb47d40195143ca220
z8de4042986f0b0000f4afda94cdabcafd91ba1db7c931f53d3a3395d17a2fc9503820853b02419
zbe4c4b89b51ad270917c81249234afe318b13929f8cf1696188139d96fb3c1f92302eaadd9f5fa
zce883e82ce0a160d59fb0c89720c8c9a1bfe3c51771e123ad4155f94c0df45c54054fa780349aa
z842dcb1ff62b6eae664425ea1f236914b0bbfaf527cfaf046692339ed3b65a637187367c2f3382
zb0ee2975aad5d34197ab2d4ad6de25c3e1e0bd1510c7c673e8f484f94edd7a292181b65e742d04
z435cfe29d7e63e960267342a804c8bb6c69dd3b92918259b3aa4233e78fd42b61f68c9661178f9
zc6134ba2c6cce568f90e48333248d76fd18cb8d8abf9275d7bc26b4754bb7237ea7f9edbf8fc89
z33e80ffa5cfa847f10de7f63485a1b6efd72498ef3cb96ef5531c07d61d46622d66cd131bc6196
z0f7eafe97847536c7554325b2e2ee3ed6f5784c7f8de94932492825510b1060b9ba5bccb32da69
zfeaa71dae343ce891f39e90610198d84cb1eccb44272fe0addd443e8aedc8c708913cb60e76ee3
z7e41de8892aa976e5e4d09f74aa6efc976cf40bbc56906204afe03c1a957d12030f8ecc19e277d
zc654b5a5b3d58dad0d696fce7283788a0c1be26f0868e378a9e8638aa982ab0aa152f4713b8f10
zae8cb11a6f683720f298b58583fec3c2116ed793433c14ac5c715855fe402234fe25cf8c84a9fb
z273944db24170dcafdba8c8f43f0db397c459923a58f21d122ba99e7727e9f8bf95d1de3ba7e5c
z9bc896926f93e04233500d8883e2f145940aff042fb2624dc307aaa9114b81868d1df9a2d00404
z1f6ee7fa376d7d2cb406f9cdc72a1ad5fd755c3312ff8156e11f27e39b128f05c593a16a07a45e
zc4f733793f8ea623499eebccf32e2a077d6589fa9b795e2806126ce0997094288e099e402bfd15
z1ad5f7f8e58a98fb71599b33c467456604ef0c6cc70d2f7c1ebca3e4a117e201a077575bd279df
zcb4bb80b3b334c2d838a7e8d8a8b855bded28ebcd8033af90e4747450af0b271202688cc01b867
z6c4e887bcd771e9ed677f1d4b0968859f241572f1ccef59236220e4c47dc03eec55195a7299bec
zeb1ccf7be9d353113b32b9bfd97014f6ec77ce66e6
`end_protected_0in
`else
`ifdef MODEL_TECH
`include "qvl_i2c_master_monitor.mti.svp"
`endif // MODEL_TECH
`endif // encrypted_0in
