`ifdef encrypted_0in
`protected_0in
ze74c34e226135848fe16db9ffd31815111b6d7fb642c521a3f628cf6da949865580b22efd062a7
ze90adae0e65e66a2c36a587d0a790699161455169ed55a01f2084f11770a774ec4c588039b380f
z6de9c5084882a40b79a175f5c2114b2b6d78b070cb806e1c0aa9258297f4687ab308bc470f0040
zb0b1de382961eeeaf2e279e1462520fc31c119af8f2b214846f56c2b3cd2eadbe4099496abff18
z15cec83ec4a77b868344aa20ba7360908f5c0de2a79abf8b3534b883bb12180f68b5d4beb444cf
z3fba8f13afb0abfe8fcc4294810f75afe452434d2d0f1166236c82f76edf1e12979f04bc35693e
z32ae028996dd85737a8f5adc1ebb94f39c940246e887647b64782cd7ab429b0544c173176cede7
z01dfb26b1f73408344a52b7e1f117f12bb9c8077b34876c2e6fdc085981637012dc9754765e1a9
zc512ce062e0b8fb16a214591f5c81e1353b900a611fe1f4886b57940b41b7f2ce99a7b84b04b90
z916f717e73bd10589c81e207ed77ec660a8cbed5b487fa50acde1b055c8870bd8676023f21ddcf
z9c98cc47cfa2d654ff1365d1f45035a045a66c5dfa8279050262529d2cac9e64fd27d9c7de62a7
z731bc808811ded9016570962244887f98fe5440167bd0088f2f049df882af501358497c3b28776
zcdc5426c7f52a851c35106bb93e16fff98478405dea402575c9151230dec03ae58c76f575ef850
z0b8dddbf9156f4e428ff80985e94bed62486b602a882a4a30e461afe18a52334ecc5953e7cf9ce
z5debf2a19a7c03f48f15a486e6e844fcce7a3d9ab1c6099ea29978f629a58619cc91770686f3ca
z58096f06859011a6a44cbde78a371329f69c8cfb385b358ba92bac113f8446aec94ef8bdcdc4a0
zc60d0e70097c1f13d99215d47d7211f9d4d76ae38b5d2c25bbaf798271d0c103ec5c3d44070b05
z9945ed3b33a15f82d46b1473b45f3146eb00f07931d5e099b136a6ea164fa1d91af635b17ee383
zfee5a10dafaf43e0f20ec701e0d6872eaa5d9ecc3990f5b10307528c3dbdbcb37d41bc4f6187ef
z41962bdbbcd223cb28034de8712b33777d5725c9e6a5aafcb85c63c02d937ee5ce3cece713cf64
z1886702da95006b11ff46d3a659a5bcd54b16881c893490e71ca846c2830f3345374aecd3c4fc3
zc35e281bc25c956dcc252ce480d782f514beaf58d9622112452179454360e50159b1493fa85565
ze28248f7b3b5cce993392637beff252575d506823cf066c282959b74c4a5080a4efc5c2643baa0
z2120378712e121eee85a212c36903cac9c4242eea048bdf5a801f52a9b13d1581b77cd50b54be2
z53990671e00a56ced89dac0690323cddbe2fbb1cc077992dc02d5564941cd28765a2b3eaff2fe2
z70161ff01fe234b7c5a63b487940a57174bbb857e865a030f709aaf8f71fcb0a964e4cf6fcd828
z12e3e5b3e22a0751bdc8b98a8c3ea53ec2e8f734bc571a39e58db375eb558e5cbb7748af5c3467
za4317fafbef65912a5f6e797b45e0ed5e1b27321deadb03734f9a1c82b207187d69dd580536217
zf6b8e8d8b4d4f4329047a674c514786d971f4d9e654644a9a9a23eb5616b64030088d565fea8b8
z98eb5f1fd2ce8e5f9058b9483f0a9015ab2c37a98a49fdea88d5af019b621e4f34bf3638a79f0c
z9f7a8723b7ffc357f1170ab883dc0785e260dfcdeade6a6490cf0c3ec7b86b72495a56f0b59f39
z9c6980513fc60cecd68edb36a0a1c5d1b960558aac2f9c8e1186196c3737ee7f630d5082c18574
zd8802772f1c322bca9714c48cead884e43000c618d652caf0756171376fb93d3ee2ebedca68c3a
zf25ce7f21cc21a7ff05e78a34d9e29b75e7826ed627967f35c68a512401d0c69599d00e669d2e7
z7cc3951d52ce2e1cebdc2673944138df2f46141cae27df10efca3cd8fbeb908e5307c25b1b34f2
z7d1eba6777c49b3979eed4b4f62606ea80977e3decbe25dea678b59fe6154f20f8c94d4a46fd7a
z072a39c276b215478681d251020f75a84e5d6f6fa948baf44029129c4b88316a84a3459f581b1a
za93ded7c74eb58cde212c63f5104f2920c918036b2d6048091655ca1c2e27f8ffd633eba76b188
za8f5b8cf2cec170d15967f8c6912042e01fd4461d00640c9c2721a60a3f14b2dd4c04b27bb7775
ze16fb21210598b7a3fd3d7a5cbf7b35504e76d59d9dc87606b44907eda48f7496c9b2728ca1530
z7ebb6d8854bb035f200459907cd57f50e93302e812f19ec8deeb89b9769fdf3b854150916570b1
zd41053aec6311aa0e6954fad57e124804c709856696ec6ddde708d57ce605b0f1be157e76ef0cd
z13e2759bdbaa43c9f3f1a7d7867122b07a957ea37b77edfbfb1c9e0d3e05afe02d16651d17aa5b
z8bf4651bf50ff29f5c34f6b094f44b73064d03c9b4d5cda8f06d9e3f9cda5ce1f51de59f6b63b9
za9fd70e4aa5d9de232e39f1676397f9acd9eb919a8fd91889006ce8143aae776d7e482f1e18305
z02c3ffa6eb4a1bf970a07063b9f801643b14e4d906f0829332f4ee6dafa12648c3fb888d3aa6ae
za53990e1bfbdd470ce08f4dde7069689669a6e11da6626bdce658e007da5839ee5fc8fada97937
z6bebccb5e43c38608b4f54d0b5e1b95a7a2176dce9f0ec88fcfc4d7e18117dc56810d4d4e7b1f8
z565bbfd023aca1a664a802eb8d33b7a838e7b0e3454a7fb8f85f5797db1cbbdd5895fe414c3c06
z63bf1abd5a8949f39b2e126233003808522c6668ca94cfe64a5bec6879d46fae162b147ba92f19
z1e0772b886ef7825b7fc8a9ea9464c8bfd2797a0ebde4e2cbb742bbec73713fd9e0e0f3c5bb5c2
zc03f2af125228a8e28f10fe6c7bef8629d134d46ae8b6811a3973c0b3659fba44af358a82ea577
z86a071fcdf5b58998ed72a5429078cd2da5ab1a375ffdb64bb0be7428434ade8c8f0695703944f
z2d9ba5892c71df90f09f650bc4e89222605509f5f9a63451ca2c333786698a2391dbc76cd9d301
zfc30e4b7cee25c98ab2ba9604da6c92c6fd76a0f1ba6b98e5e15595c6a807803807452672b4a58
z0dcd00a0867a22a39e0a1fe808f2da6bbc7da05eb697ac2addc76506398c8f764cee55a6c53b76
ze2da9ad9c7157da70b1b3e3b2cc63fcec82934fc81aab87b5de16099dd9e13c6530c50ed79bbcf
z357077904656de5bf3382ac34cc5d81a9348dc3a0c03c21d3d0144274face395366c9c161f170d
z901b18d0e35eb98885155042fea15a272797cf1620cbb4d338c17ebeb46698cf38134141d40b8d
zf130367205d343f0f1ba8208f9df79b4e36c358e66bcf6ae9311a2737afd627fc386a848b48f07
z350d3becd650027619f56d2265d8c6918fd8e11afba3ac3949f29f1c873b0ca086234ccc708621
z8459c02ece7c971e10f612103c7ade4ae79ba839e01bcdb8e7fb358521efc4ee6f82f2ad43887a
zfe91230cc490d5d79d7e2cc8d2ffd19578293096e813b141b49d62c78e7a7b0b6c0a6831f5a8b8
zbcdd87da3b8bef5a31d10f16df8b419e125007733ec92f37656cc5ac884682884ac03f0ed9f2a6
zc5ced7278eb06b871e0b87d0d170bc487f8759f32e63b59183b4862163009678854444b4407c15
zb95f603af97f58691a9c51c0b162ed13f00e9a245a25cfa9cbdda4d71f36684523f3c1dd910875
z24f54241e35a3946b8793d44ada1e500419fe6488adc7ad26b7c54f2bd493cf870873db626e258
zacb84dfdd0e0454dd27c496753c241bd2488d1d3a06c22f08de9ca6f5d3643f5783ca5abdb323c
z9020dc5c6febad916fa4f81670b106eb0eeb5a37a5863063e4eb5a5287158184db0059e5344713
z6e3557b25f1d85a710febcaf52cf03b91625056a5805e1204b09d2ac2362bf2e0c4360033a6d87
zcc008efe8dcb15e55b1bd3ece274421d528f7147f239c8520aa9a369af43cb972855a5be502941
z4d83f036239213a8416eb9721bb01b8e80416d0cbcb4a14dc8913d78ed0f6af20294c1129fa5a2
z8edc46c8b0d4fb258855a3e85a9cca9a2241897790ca941436844c62ba34dd2217cdf822a32941
z23f12dba07d4664b701f44508a45e6bbe78c89207968b0e1676726a9d2f9a620e2db2f205f37d7
z1a71575fdb32245df3bec121f7a90bf12afbaffb028486190185eedc08235ffcae4d5b8ba7354f
zcd8936421e9f7b8bbf9bac228c769ce4b7b4980094b8b8cfe87f79a01fdedf59262c1f69e8c390
z529cbcc112a2f1116f0a85505478b06d1bd540bd23513a17b5cb59709864f61df9d91864102398
zd1f8cd58c232500d52f6aa590c453d58afc8529abe1f6f32cb8b15036dcf896bf41f01ae193c50
z5b6d090c9f0824ee2b5697689663a5ff70bec80e6b463acfd120a4d563b966f6d37cfdc27b2dc0
zeff3cfb7d227e3b804ec00245215c79af26047965b38f48c4221d67461fe5aa8c7ab310121cbfb
z4822f19f37f12937497eb601ae397c4e4f7c2fe33f7fe32dac89b1901765afe219dd10d6a79634
z59b2efb5f1c5218c5e74c1ac128e07a5074c7d8e8abb08db34358b0a3b64f4aa14c2af20867f39
z1c635f777079395e518a7f575a557b8314dbf7fe4e3c9ed1b7341c8bcf074d19c40e851ccfe99a
za30532ed51536583ef3e60f0a93e945d0ca53726d4988f9c183610b5a63ecdb658091a90a48ed9
z8baaad847a72f575d2b91127c39c8621287f5a6b22c75ef9b4583afe4156e51377ebf88300e431
z8179d0298ba162dc6a86f7e1a5a3319b845aab1146c467da1a9cbc316698f6eb2bb6cd84750c0f
z4f40ddb06faab5abd9d13d551fa214f463547961f6934066344185fbc480a92ace3965aef171fc
z473df7adf500c53b67cf0c91e32900a8a38a48fa27ecec101a188473759ffabe61b115d36a2956
z1af73cb60143cae1e86464f192aa426f225a629f86df28f6326a1288a052348d2f6d6351042ab3
zb3b7c84e2af2aace96950009f5b986a502aa959e5630dd6ed190757bdcbe16e017acf4bce05ba2
z7d044c9509495e1e06f7883d0b2879aeeffa513d1da094ab52064280e78682a714b0d338a807b3
zdacef2ebfc03cd828508c5c535affbb59caa67c9b4069b0d302a46deb3e1f2613e2e7b55a23fef
z2e594e83152ebb21a44fdb0461855c770317f89912a639dbc5db5bc2ac66f25eb7b480ce06ba11
z3c8e22d2215a3668faa1e5f637efbd58f36bae2e9bd0e30fd05e5337bcf05d06cacd94fc520fa6
za68cc455fbbcf2ab9aa5359a34a8c1ca0b7ee4431f71f381310bd1164c1e656cb02c487d112831
z4fc9248633b1b887f3519828315ac768b38ddd0774b301b9699c45b1c826d8ac6cdbb2b6c8eda6
z8e1842ac2913eddd380411ec8c35bb990be73b9801e6b878305d17518b6196b58dfad91d67f275
zc163006a7218b8b5012742141b775ec03baba82d1f5d67cf49bebe3b7eee802703b4210a8ab2b7
zacfb24a9ca5d792b420259ef9e2ed46901fb99addef009a3f86b45103a30ade3833a3ce93d5497
z955f3fe418820ace9b3ed316c4e658cba4cf5def2755d814fd9410cd04fcb927ccea714837126d
zb35546aeba9bc11639bbdbe92887006e5c868ce5591ddd0a5c6bf6ad1a11f4611a7e3160d9e76c
z50bfc111c3673adf2384d3cf32bc027bc7beda233e3fb2786d2083ed0d606cd37d1f66cf031ba9
z68b5f8f14332090ae575bf2a14b8b011b56a3837f0bcfc53134863ae98bdd754f9203549aea056
zf33a13c51fbf398756d8f1e48cb2c50b218a8face36c2f6697194cf79417ba6f93243ac31ca878
z709ca96fc00fe66d7475251eac855eb6acac73b9b4db47cea38e2db9cdc27b081cb88499791a49
z11626176239a280e9124c5fbe6ea1eeee7c8ac8a70fbaa167b36d12e24a8b44d16a5c3fa7d8e8f
z9fe5b88c584d7dee213a72edeed6b08af08e2e91a98aa20b06cffa5948345416df57c156365618
z49271d818552979144272e3bbc1abded0fb1865113df267a003abceca9d12b5e2b7e4b7975d198
ze3a05c781ef92bb3db6540ec7590a8bda5dc4aa1e0c93842da21c746e2d1b2e49efbbb9aa3d0d7
z3aed2dbf8735bee2ff80d5920837afd5605ed4fb358091c1abaa1ba30a4faad8a2146daee7867f
z3db27f3ccda37c8a3be2fb6fa709737cc7fe63bef2283b72acff91fac22f33ea5c19d2c37842b8
zb253d63802453f191700500afe475f9b1d8f343124d19a14f47ef16c5ceffefe0b990e2662dba4
z51607f8323dce4a76f9e6abb9271f6a283f7a09d30775b4dbf5eb3ed275de35b42866bbe7d2d74
zd65b3c74cee29dff5d5ad7c8b2f55abb0906891059c49f94733073d3301f83c074eefeffcbc548
ze51e5b25c72f06efe98f068b4340cefbf78a5594e24cf5f94e71fef52ac8fb723b96a4f91a4b4f
z25747ea37f8a334c7b5238e4bf40e8737b8cfc3e9d6b60f9fa2f441b4a36c921fa32a4b3240169
z7b00081db743ce95421c280c17720cb674dbcaf5bd1cec0db41d0818f796cda1dc1bcc994748cd
z7beec1f6eee5592b9c9f08d4c5a2e016c0991c7f0d4eebc11c37928968c4d3d2eeed4f5ee6b11d
z8ab9476f2170b31522e0727fb121467b047c124148e540d01a41b6d812222b33d6c4cfc8b6d156
z73862a908e8e2c7e0c745b6c5de4c902b43f03d9eefdda6ca82391be46fd615021767254113d29
z932f73274c47d7191f3428594af14627ed6d35afd247487b8a01332ed629fb71657529a32c9c43
zd4fb703bda135f839cc074c454014be0c5cc1c0854c9388f3a53c741ed0dd24f869c616b467761
z494a2b6ac6336f2209780bd4e5178e1ffdf4f0ae1cca58890480c18d5e4d67aa631c0db9b631c3
z1c8f95c9ffe1b484a1a5d1ee3f2d4775ce82da7b0c6c2caef667c15980de7081f6e4a5d69414ac
z87c30c98247b2fa7bd91bfecac35f7ea06cd6f8dc8eeafa24a516371788b0fd9709e77cb1bf5ea
z0cb893846e12faac0bcf2d041b726300af21be5a0ea034c863d18758035cebfb6a2d2e64462fb0
zc968b8809e02d076e2ad615795b2afb9420a48317568531b7ceeb0c60a871d9b477a691ad32aff
z33acebdc4f42f15917b0b1d911d3c4e216cacc2d458575d63929d82c2511f6ce7cecf5f647b372
z64f82c3f15787d07bd9ec1102943efd3369b8cc161dc3d0b8c83d9269590f4edd50a0a707e90f2
ze579c8d003e6f332fcd71428c3be3a57a16b697558eba115aabbd202db72cb3bbb9f0bfc3f07fd
z9eeefdbffafc7144914b52a327058a15ae5bcdb9145e28c0e820536d670b735cf690a0eac54632
z49a8342b9a2dd070e8590cf928e9598ec3059ed49245e869919523b104c09ce5611f6cf1ca6c57
zaa84b301c246d735db1422a8b5b2694f33d0f5f8a28f5184d7b1dbe64982ec95305b93d5b2f73e
zf2d481d9ae51c8637b6aae532ea9419b01d5a49d44fe45e7dc3061bcf529459c8223c6d300dd56
z1e090fa73200983be4480ff9b42b15eab44906cb5117a05023eca82035813f691caedbdbe4d80f
zf54c193e4558407e7fd5a0f43ce08ab08997d1e2c7005a329855099197dc08a32a8160be963205
zf428192bd41f45b92ecd519010d4f603b8f5b4d0228820c15de3da2c4e9a637e7ad7b4fa0f7748
za8bf4d8d4691f981902affeead4ebde4244dff58adabc9acd5acf98ff27d22ffa42c14eaf14bc9
z6e851fb241af0d5ffe5b2e846848ab58c9b7cf4a3d773fb5cc3cdb4e483f6f60082ba9f4740ec2
z8021e25c296f61b6ad61d4cc362e463a6929ae9d072573ba9aee1620c3088c1045cac372fc3d03
z403970c31d5f1815a9a0f5e3b9ed0ebee0ddfa948e0761edafff388b6f9986d673c3746c59fe07
zb698735da45872253631f089024a4198ffe610905381c6683a52c8ea523e5dd2074bb2f647f135
z87452be9d2454f4fab981c12fdcd66d8089a7125e81663316a83042b18bcbf61141f4329167775
z6c89e33a13ba2360eff2d0e29a8de8e050e81abba3d6cd2b74365651d0336aade3c538e800d82f
ze27fb6d0d6491cc84c1079322ca7c5c9453a96d4cea4f6c84da9627ef75c9c7b57eeebe5f9e2b7
zed2564ca94d888f9e6f9ef8a0c9168a7692455fbe933360d78340c0c856cdb00fb135586aba588
ze2b9ea8a9b99e99227ee8e32444cbb0e01f50aebc760a7d5cd90f08cb5dcd1e305fe45ffa4bcf5
z4c346d708d424c2c6716e12d1d2e515ac7f2bed65fa0eb114235971becba1efc34a4a00a9a6a83
zef9d003dcc4bd425d2c410776b62e9ba3940844f546fb506f9c1ca5db3f2eaf3b46ee58f3a6b53
z4f4abd9cb8a25c05cfd40cfea2f1a2016e4b8f40769cce9eaa9dfd2479594d3d143c4ba89eac6f
z60bb170c17254d8b67e4586d6632d728bf4d66b65a9df639fe315e7f78245da99d56aa2019bd0b
z9ad2721715a54536dc1b13a1ad939fad62516581884a965d59f7cb674c7ce64102c0e96164b8c1
z0251c9e9b4fd6cf888bf2243497a8a6b6b8775ac62db7fa45363b624dacd803706dc685f098cfc
zbb31d1368a5ab70cde14b462e2e28162cb30d0c575a25501bb9121c8a6535fea1bf1b8febb7c08
z1e95bc280b82c45453a41a20976cf6bca68a1f085021a981b837c0a67476606c5024110c6ec235
zff819fa5ea84d453cb5910a31ff8f42fc16b0f103d0aa0c61749c0482d33997524abfb2813b0ef
zaffd71d519d88ab8c00edf44363aff26c25927d10ba29aef7914e3a88836f8a3c2a0972ce9aecd
z3ea2c32a984f9b4214158d7d5cb98ae0f2ca42a170d2bee6b2fbcd3ae964bbf9e4a11483f47042
z50b2461fb3e77712a2c55393a1ab98039b8d0b4e2975168afc3f3068f03117cb27aeeb54920725
z1c55b5ab8d0518bd01b8e771ecfd2ff799a84ca90d0752d59350470d0476a8c37d9aa61e7c6ce7
zba9ffda1480e6fa592b9350ad78be130884b192009ed0196a3823abcc03becb42c8be62bec323e
za917b135d1951f3221cd761e76ecf0c8e0b42e952f4ee8a2b4e96661a0f1c98b96fc4fc49159bb
zae846fd329753345398293fd26b8c98b636d7ec384bf25dd65a81dbd206baa47f8bf2a4eeeae7a
z671d487b673322bf21283c9fbb46dec5a4def487ffc05549b312c12bbfd9229362c2150ae68447
z5793a3f94bc5b9b52b55f3130e78c30718ef07918cfb6d335b626365877bdcdc8f3516d7e9b1c6
za7bfc2078d49b7b89c1329389c6ac8c5e4104b8dc079c8dda01e5a79b1c155155610eec0df58c4
z09eac3d4991b82365962491aff175c20bdc2188fa1f869dc0b7215891f4797533c592189170597
z45939ccde9f944919e3831fb2b3f7482215f5b3f7563589f401718700c8063f0c80f511be0f8ab
z98c73ab4bddc34646868810f26f131f662d20c9abc37f81fa136c1758d64c84e1f0256042bad6b
zcdcc9237fffefcf1e8f1d7807896a87734fd715873f29a78234aeb90143140440a0ca3f3239007
zccd2efacee5789706dca9d3dbc7a25402b9673a1200144cb7f777497046d2f53fb739a39f463ee
z18c94eef55ffba575071b337aa8f3c934fbea1ea30ebf4a59b1264927cc41349675fb677b40efb
za2e6331180303821d1332b6cd07c046fd4189bf57da46bfe70e614b0495bd9a0257177a369553f
zd06475de9e4367e87cad3be7aec65aea72f8bc8fa24c966a967175d6b6d685e1394ac48dd3f380
z7e53551277af64996b9e1ddd50803abe174be7b0480b22aa63cada1ecfc2be0fb62c867166e4bf
z6b6f56c0710a75c9147354992f17b5eca8114b3a1a1b1c84c672bddf9f04b9d09a300e9791aac5
z21ac3047310a8cb501f3cbb624a8fbf48e5b2f30b3659e4ff632b66c73d2b2dfeced233a8f3be0
z43df9ec4f3d38ab75b5af0fc9d218b5a10554900ac6fa8f71ea7eb3fe9384ddc0bc08a825402d2
z112068a77c8dea0b64ee6a52f25eda0be19c5c6c6b665e7094eaa6c82c4179cb6ac64f9da3d58b
zb6ea03dbd7b89f12052a1d2bbe87f7d0d9d6a25be7786a144e980f6594d22b3e6ee79bc2815dc3
z402c6df5b155732352188f5cafa9e0f1113e3fe2e9086b0c38dc6b2d7d1fd6122979960e7cbfd6
zfec7dfb4c3fe20a3483a3c80478852adc66632b3e9124e24cfbbb2115623e9bd75534a5a25221a
za3a5d063f1d27e5251ca7e6fe1c0870f2a51283a1ba2e188d8d6e5dd5374c4affa6a0881b18b8a
z79b2850e73b7c1e702ef2927dddee51e333e1e5dc479dfa949780629b7d5f123beaa8967b52961
z1aa4be09b151bd948caf898c00d1f43c9d93a0f88648867ff5f22471e3d09dd2cbd08efbbd84ba
z35f14c97ded8ef6a21225ec191384c7bf1d8c901dccb85af2d342b674310206cdeaa54bfebf6c2
z2f1d8769b77ad11075048b3c081481d2f07f36ef70abc725ad6cc4e79f6eac08308f708ee5c2d7
zdace2c58ea9f836b6a71e2c23a19280ccd1fef6834a0f89bbcbc0d976b5e25d3582415537e51e9
z2e031b06c0a8d69fa8d87890b237b7e6665833dbb2867847135caec07601b45ab4cd4f3d73ed3c
z9f644f46be4fe01fd42086238887b40f007fed022cd38a5a432d14f81727d91411ab40a795fbd9
z7e3814db9f1ee9803e98d21e1543241e6ac818dee09a7c97ee6ecddd8baccb8ef1029149c31266
za16913a7ce7487b9f097b35ddb6fecc398d16dc0573ced0d80e77e27b7004a04fa2ef4ece1962c
zb719404128e95dd20ce0213ee4b1d0fc6cabbc7a50b19ed1e27706ddcf0b5b7f09a95c2c8a1745
z4773ba3ebc06e2735a5f941a03177fef8eca959d7ceaa47302ca2f4f9de9708e97b2a80d333bef
zc302a348db4830ba4ad058986caadf59a42d4a5c89f898dd8171cb0ca7ae7902f31f66728e6ff2
z2ebed4898a722268795779c8409c17bf25e2f79229a8f7a2b89a2c894de94fc922ab5afd2b1b0f
zead430817883428e1e8c3ed0420e3a06974a3f717726d5b895ea86c8fe0d111ff202b136ae190d
zcace9b70f50d3e716987863dc290f5e9e4287b488d4476c670684ee1d6970a147766d30636609e
z3647f5d3b36b2bb669efb4a1f5fdd2e295bd0bc22278ab78dee1c6c853646e433a0f57461f5add
ze214758112a47b22384580dfa530fe761442b0c88c8ff7df90989cd878ca5e48aa211e73706458
z0fe45b7e769e86c5fd3252d3ade49ad4af426fa71fac881201ed90d11346874a51ccf8d576e3f6
z4bf1b4b59c7667fa16992b0b4c318c2ff5728d61064a7fafe14912f0d71c28cac76831e22581d8
z74e84b84f54b5d729f2abadf83a2430b8d96f53c7ca31b85b31dc2a444e8ff3bcaa276259080cf
z656eb175895b7b30850e8700fc067cd371fb1bd6d1462028b7c5ad3a2eefbc26813321379414df
zdef0212ef281880d0756f6c24e8b7877f1f68a9f0a2a1337351ce221dc106670400f0ece5f07d1
z608876994dc83c6e6af111143c15d57ad33ee301cf5bd5c77986010efb4f78f09890135a15fe1c
z4b21cbaf7e12441ea29be5703f57de6e6cdedc3e2c8d2de8f52d76a12eb77d16504e64c3e540e2
zb2a636f7e1e23f3239c166488df217671304285d74058188abd2bea5cabd684d65f171386522da
z5ada004afca9cdfca91246ad8d68744790b5db68ee2461f864cab6066d6e037b65fb167f4b043a
z502e218b2a038bc41b591af42e31b8602b3488c901d31af9ad0e2c93232408610e8edb10d79629
z9d593187a1a9c213e4cf6ecc933e4fa125083f09fa00b1dbd56fb07b234172e61b2eeff5038a82
zf5e57535b7083da5c41e720eddac46eabbdefc208e0dac9f77d64014e7a965d31f95f0302fecd6
z6606541717298dd883e26d25593f79a694d18f4209d88c89d65d8385f7cb69e6deb4cb57a0d2fb
z49abdbf4577e8a1ec93b274d37fc614fe69ac39b382c2ae2f4543fe150bb3e472f8ab7b7948f54
zc4bf6512ed7eceb9f6d4ceec0fa6300457246ae8db305b50b4264f910a484c33967a1614a951c5
z83e9becf2c7f10788d00a3ed17962571dfcc55107ceca83e93b0ae00cf289b46cd8e7e080f32a3
zc10c6c290ebbb127994a505d6d47cb245a5da1a1643032edd36a3ba47556ee58c889dacbbca187
z6c8b0bef9344f45961f83cbf8682fe0c61c0c01dc8cab4083f06703b9f37e218376a6a28d1bfc9
z0f90efd2fd3b46acba420fe73402607de3057279b8d14a0485fab6834392cff3fa9e464a62fecc
z88ee71e89025bf5c5d4fd8988e2f815eb6230a9d75d59eeac7739e3bdb53c45084a35563f9db75
z2c664afeb47ea9f8a3bcd413a32b260d181ab904e6fff684e4959c716277f0e4415624383a5402
zc2707c1a4791e5cca170c8d94c8f89183de696a611e270fcc29000c73fdccd96eaef1c171611e7
z68f109a08df2a85338b8648bcb93420c0db2dba689b4077ea6489b8217c5f751a186c667bd7211
z04ee512d8385a6c62c9329323250c68ab3bcd8bfd638b527fa9715c11b4836ea34a3ce79383be2
z3835c162b13a0053f4d4d1460a1364cc7964b1b86937892f0f98c4db116eb6222acd39f7a73d6b
z1b2f1e1ff59c104937df8b67407a00ba845231ab32a8a5a601af1e7fb9c5f6eb73e4f14c5d6103
zaa6da539108ae7fceaa3f6bad7132b05e1c77d2ac8b0d66a531e44199ae5983b6c5984922330fe
zd201ff93ebe9a4403c821409fea92ea27fd47494a2e88be284cbcfe8b6f4e18503ac3fdcc84b47
z67473a8c771238ee535d1bcca9f512de99837ec8aa3ed977cafb8e6266ec122b3a49eebc42ba6e
z6410c5cc99b8d3b24e97e6be4990eb24ea7842df229c9a463462606afe07971552c15deea153ce
zc905767246fb0a2b36aafa247062f571086b45eb80d42e1ba86bdf49acbc30539302e870ad7aee
zeedc5cdb3091f65b1def3b13e7650a3cc332cf5f0807b7da1c6df48525148cb019304df2f45bc5
z016dffe679232a6b4a0e484be38f87ea04fae1bb4f8c6f6a0ae56d9f9af62d122877c330e81b8f
z8e24b3664627f0b6c516e9c370b489526fd7579b3d68b5a5417932ae1585fc65bc790ff911754a
ze2e17633b990a845c618693ddae91e1600c04d82ad44f79081839d969bcedeacf52e68bd176020
z700cf58e75616564dcb8ddcd1b038c884a0baabe3d14ed59a1ad369b824553ccebe25d729c4c76
z9858f3aa8962fae19b34ae7578c37ce6bb7f6288eb2b5548a0a5121743edbb209621c4da355665
z4493dfd0869254372aa03a0c6b10e0265c17c77bce25c632eb4ab911c21d18e7957628c1246bb9
zfe871010e96752c318224a3b611673495cb1d9d8134618f0de6a217a89863fed0d5371b683d1bd
zd743a4f15d2cd080d76c327cb0d1a3bc4dbd35d3e3af338d17bc999a3579dd2ce2d18504e42efd
z573c96b71712100c0dfeffb09a6ceedc34b41b8c1bc375612495f346400a900e8cc8e2150b0bf1
zb4fd302aff4f09d68b22870b9741631f2a845834f67cf24c905b811d522cf8cd3144ebc11c699a
z17e5a86119068a7766b919fd22bc554823a7c245497473e7580b7fd2df0dfbc12d76d3e5d9b470
z662f81ab5439f1742b61f45ec71102453bd2fdff3da36b8ada4dcd53b67a84288451d0e021b140
z832b4a7eee90b7ec254cd1b1b86d82b9d1c1fad75087b27c55a7f5adffe24057f4d1c00f20d983
z7843795b52ef86b90d9ceb7e298bb07e57e2f0802a9a730717c5069c5f7e90f56e377e398801b6
z12490951d0b7a237b81ed65bec6b82c7a6934fe2ce54c626d95ff23bf1881233b3090e786a5114
z1e87d81e758eb8a39ddc18ec4544b1ac97300da6b4acabf4dbe884835dcf62d8ed9b36d7dcfa8b
zbf0d7cf90f76e92535640ba010fec907500cc98c588e43629421836734c7e96044def7532c9896
z5d8746b0c83ada5888a0c104d626bd31a659fda49ccb2051e3fcb7e1948e0ee8ac9215ed49a275
z6d33f000a6d2247dbb31d2d880db63ea5fbe115fed9ad610c0419dcb2abf39b1e8a0757e7229d1
zc245efaeaae003156da78582698bd5f523d0555682de08edc217467807eccea997c6f1317ef62b
z5b6be4c1ff0606e7d2959be903522aa883f42a9c42450c76dd6be8d7f6c0a8a71b350279136bf9
z1ff381d3a44694d61934639eaa2415374f899906328261715b58170d95fc05cda0eff1865c7550
zc7dc7147cd26e537ad27139fa20da636410ca160785c59aa72af8c5da0c8c46b094bc77dc7b693
z6e4dfdd900f0f136aadf59be1a577ef3cf3d1bf7ac3a30f7fecae5d11ab98dd73adcbf0a62d1f6
z684f6152b8fb6b66cf42222b382cfe97107b7cc6f49d0f1bd774f230dcc9afaaa16e9a19d74e56
zbdcd854bf4a82d6714ba299c032cade4b9338bb88067195ef3d44b445c27b80f955d4dd1a540e2
z86c3ef5d2cc0f466ffadb086a8f1c2ab6bcfe8903cbcc18eb71e7932ae43ae9f7e2e631a18dddc
zbb926f8ef83fdd135b840cc55f53d49cae59455637d0f6246d1b3f78d38abe6c37a39693b4ef7b
zaee488faed69378a47f17359b10710c45e7c8217749e669d30e7fabf1022cf0282976aecb9c794
z58b6241e363b16185b23e6bf2923416820ebbe04ba89ffeccdcc63230f157cd219578492c1a783
z37b994e3cab6005fcd9d530353d8f7e2dbaba144b9159b664d4601f4470bce702945080603af6f
zc722a405d64b90241f53183f4f11f6fdd655f53002d3531fd8ec5d576ffeb113cd3e9179be04ff
z7a944bf79bbd7abac62981401aacf7a5f9c79f3a3f290c060be5a21d2f0125695b8d5ff5c21d2a
zd08a84732dbbce1b3ed0222dd95c0551e505a6f55f4b15f423622c09495795a2d5abe078222fa5
z0160cee44cb04ea744e823f74b87d478cdd0e945df37e14be6a29a2047ae3b0e73496ee38c1422
za5063734f05ce1a98df56c3c4848e147c84c40e6c908c403cbd50e59545a8f8ee78b67503018ac
z427dcafe2fa57559fda4a64aeb202e9290dd0e054e7e2fa6bd56166cfe79d5287c177eb13859d5
zbe69b5b0cc715c5d3fbb67097dbdc39b3629d80e8096ca09b977f217075d6925130555e1a9fd4f
z89d74b279839dee0ae3b359975a99b0d6fadfb79427ddea9e4a1eafd5df6e7c38d6bf360d8feba
za01ae98126fe0d3f1fff5f347c445c4e7ccf6d92515a1ef204576d29e7c10ca6ff6be855a505d7
z42dcaa33f43cfa858777a826ac8490e00612f8b1a7f9b5c1eb2489cc8a0eac5a4b4a6056f3dcee
z303ad86a48cf5efbedcda5a9c101e48c2e6c6bd0a668ccdc0f2932832d4a3df401363096c9f500
z6cff783a77563519a701ad87f2624fb292e94c332fee7d949bfb0984afb49eb907b0014d4087a8
zb890321d6ccf21e440877c5c730015502bcc37eb49721a65249bba5e62e7e3877330f7cdb1ae20
zde64ec003e3fb7ec44f17f0f3f405cc8a5b7cd27968d10f5536d38936aa58531ca8d039ef1502c
z3ea6c818e3a5b347610e152a46ba48375b362f2adb82f1d6f0c1eb1f5a2c8e836205c418395fc1
z38c21e829ab1a6a44b777a7f554f3f72953d6959232acd1c5821efde0de715cd3f9b1730486712
zec7a8c438146c263a97b4a78d44a0d43ff9302234d47c2b07237872132b1af8bcc28dc72559647
z5ef17dd63b7704781e1406b01bbe81762f9da74676930f7319537a3affe036458ea6bda5b4bcab
z2aeb67f32258ef84f4148717ad4d276125a2c036d6af42cbe94ce42ee98748fc298766d3e3c614
ze6d69cb5acfe098e49c4a9cf7bb1202eb989412317b44d8f7f0ddefdca5f0086ee3a07ad3cc264
z79cf0ff3e54ebf49c4848100e830eb34e8bd66659f71a4c5f812daf393e8621de550620508609b
zea9b88448bd540eb5fa309e96395d7318035e368cf27c64215f35430ffb9e91482ab81e09c5bcb
z5784f3e25cf8adb9f45ef3758637cc54c89ac22839baa7d8c10ecbb450b2ced8a74ba21264a697
z272d3280a2b45299032290487a076edf98027146244faf5bafd70c2db4088f7fd65e67697511ae
z01caa556b6a2f28574d1d509117fda722f43dc7094212edf36796567358e5c566e678ac4860e4d
zfc9d8d53e09dd7543cea1242fee0b313fd809aa73406a5880fc43465fdd811dcc0569eb925792d
z56766bf4d50fa31d7361be4472c77fbfb4f66fb8603b6daaea54d0d3e49d961b742419d2d9cc80
z84618c646fca68364a1be6bc1b2491dddc6ea55e56027f31dc5f4fbe8b4dc52583c4e5937a38cc
z7af1ede59e69a447d425cc269f904c6e93b72d37924578361c55480eb86985ed3ea03d1dbacaf5
z3e19cb580db4499dbc30da77db71cae17c9a43e3cf4cda21f753ec1b0d70cf9edca5907a97658a
zd13f3e8329ea181e0f1c77d03c5a90b8d43aaa2d00915d9a980bed8858afcd19e287ecb03fc6c0
z11b06bfab1e225971e6a5a0992d0a22d327c9b914ffd78bc79fd78bd09ecc14c0b43fc18b4d672
z257797e7e41cba50e93709784629f3c34b22861c08ed4cbbde6bfd11bfd60e5297566d1b82c9c4
z1a13e0776155c32f51a4e2c5ce9509f9f53ac3d44d3b2117049209acc043665e790c4ca3311c7e
zdb66470046bbd7c66e4b892d571959934af20e547408bdcbab925c90f10b221fb96c3d6423a0bb
z2b1937a69085aba7c1fa0ae04910e87c0cea2f37f3b56fce3b9c2dd72cff53aca53defc953e767
zcd799ddfc57a531c7e3efd2c832fc8ec9bd1b9b62944649e546f9337b44ef902bf16c0110232e7
z5fb6cfdaf1bfe35b1a89010865264e83f1ff64209ed0ae9d304b3775a4385cc7386b07c33c5291
z6d2dae023e50e3ea78bef80386187109933442337b96351ecb8eb8d5da87832b70c22ae3370c71
z2357fbfb664737737391e2e1650bede564c1030f9db358e3b52b92534cb6268ddbf075f0b9500a
zb841ab86b00d6fce30753757b88b4c3f434243afeeec332e2e1b9c3bbf604fae94988ebaa1fdfd
z27111af9e47d57509748925a7fd81e58419510cf8211e0feb96803d84518a8194737ca9fd4179d
z1fcec6d0b13ddf490e10e06ea93059385e46ac0a018d4a7fc0377e34a3dca8871a687a132dc577
ze37281382536c2f1c1956b59fbf771b2a534109a01d5e571895dc7fed4fbe6074e6cd39d2486e8
zff397f489516ae8bb1bdf1828714c27be6935be8b77fd9afa4663dea90a7cbd089c25d916b0f6e
z1aa933c947ad0e07fb507e4b0c91297ebc7229646d9d89a7857bc50f9e1226a3e8f9a904a9ec7a
zf719b64e24c3515f03f67b9f9e722f4301c83a94c50eed88edbd8ceffc505be58ce2033e4014f2
z662692b6956408f5b07ca1ccc1e07bcb53d972891f976b69bb4e645ac0132ac1c9fb5726a69e74
ze5a1f67240866b35f669433af7b1efb8ab36f8039f1ee2b03e765f138912678f0dd379175c573e
z79cf08c8d7340d404944479d5098fab89c98271cdadb8be3edd615b064952bad3742566449161b
zbf811109dd69ebf21e4d1fee356a3524e65291d510c0ca5d885e8e3173781552162dd4b0ae84d9
z7edf177aff02f6e7a2b6d6ac863292cfda61a614429b1313a1e3706846705ebf3aba09f1de5614
zd64f7ecaadba13127a914afa139b471a3cb030d220dfbb6e40059807d105d49f1fd7b83a43826b
z49fe28e970d45eaf817ff0b659be8526dba2d0860f77b7dacf50eeb9499983d882414b68437fbe
z9ba02b479eb31a26f1086552699c05164df2eec615eb5b17a8bf0da6aae738c2a3103e0b4d39ae
z89aad5d63b168adcb6adbc291a1c677421655cf478e892faa496985e857d80d34f97eeb7493f5e
zf2f8c93cd69973f0b9733aa7095755189057fb7e5a470a37ebc26d1be9f0df21d183e280a71fe0
zecd03133f507e921ea7c2a8821e291bfe57c545f54c3153b87fd65275acdec434439ffb3921e6e
z710b2e92ed5d99049d297599b447c2103915c7b8eaf2e8b4cb40e39c23e8a65e782676cddfe323
z330d87b85f9cb7bf43a293bf27ce6605ef6946089c168228c47596a714b0e9969bd85a703761ac
z8b16a53fc4b1d633b72b2e1e922277a00903e6fe45cc13bee3b36853a73cf7bb9d2777ed9edc16
z34f1a238585a5ec347168ce72ae1214be7f3e7184c18986d1293b01c32ac853b8df345c99e04a0
zae009d0d809c3503f8f1a29fe2603188ae4dbcf26fc8dcd559f6104c0a02697745934d9f8769ca
z0de0c6836833e02ebba4243dcbf0cf0081eea13abc2a075fca08d5422f62a1730538435c44235c
zf3d50c38e3d7f8c873a3c66e51b77d0d2a97d779a193eb88f3e7ddc6f1929f4cddfad8878eb584
zd86eb743124cc3aa0846c4b59644d935ac4cce8b8be71ea85f0936a7b42e831d65cea97963cd5e
zdbe94add26429df2553cf37a436e6398c3e073a310f53fb4799aab443613f02cc9c185a97cbb7a
z9841a6fc29f391186bda60304519ffe74be84ceb34a042b1194d9df19b99edb32bd2926f293fc6
z316c75955f1aed31347192c83df145460cd506009721e0fade77ea1b208d59d3e3a02f8fe55d58
zf31d026b88eac577ca08db708d3d67e8b13c7c3fca54705b6cfad64116efa8ec3331cf0f5b698d
z33f1bb6d91240e13b965d4b02ce8b344ddfba879ab82bcc7542c7a859d26217f2dfe7a1f5410b1
zad4016607d5752dd3e84fc5a8aada901b743221104ac46dae08906035c054864053a4d910d2c50
z15a1bf9a9fce6a665fbb9015c17b3f60cc56f3ae2bb974bb56e0640f18cc3481cabfd2e2f09c24
zeee071a94d5c695dc9e4b6377b2e4dc01e5cd746583261c9d21a8ed8fd15d8cea7ba6927681f81
z2a728063a34990ccf7e22c3c89758641ba10a556df73189fd60946dabb0e8f3e753744177bed22
z7200b06fe503e0f2e163f39fd0c3e5595ffb65c4494b0c57d54abc707b5b88b337229975f1ca7c
zf13d603850bb77b0efb8a88fe0f54526e49b33adcefe0b3208b53c80bfcdf1453739bad700c2ef
z5e1080a97e44942d91edd0ba4b6ddca1f059c16945f137fe543a89c31a0f057f4842e596434b95
z408e36c43c3be73141a310cc69c3336a611ab28a34f78046bf8a54d36148d174ead6265f7f16c0
zae78e3bebda98b02ba8abf477f0ee8bd38c324924d2bf7eaa1719c933066ed2e5a934b1a932fd6
zcc1e2d38c144f0157f295c1bf153df778410aa1cc5e36560505a9a0171c2c35bcaf66bb013fc3e
z18975aba689dd2e7f62696ea1e78a3de09e926ec43f0c11faf66f2e9319125d34af31fd44533f0
z83d7edfa5dab4e3a26818c8a43818223a989531d149ce7e7317c96497000b87bc9bec25f4ae320
z52deda9dce53530b9cdba9f6ed44d4b56aae9ba655a8ccb656f0c38c24303bf3981c0f7e854726
zc7028b2185d81923a00cfc0ba26582a4e01e750c9e974bcfd8ac12cbc8d0b049b368404487acd1
zcdd1279d04fda86839c5e0118dd682aed5e91a5f38cfa03d4e4a6de78eeb95d9b29e503d8d1e0c
zb3820e036a96d1ed111000f9a25d0b065ae55b8eeb20d46fdf264ca72af9c30bffdae67088428a
zab3ca5bc805c8bcaaf29632fbb6864ce6a2019bc3599674b2fd62aed507b8131bcd173eee60cff
zd7df99e3f355de3918ac02b66d050e94be910f64b8d57a9250eb5a6340b9f7c8dea7b1ae06edd7
z3f7fcd21fffb1ac5456703bc2a4a5c32ed222dda333640bf08917cf3ad808548e38c073c426829
z9f3c4630e3441668e1e0eb1c37fceac31daff2c58b5a07561c32f4789bcd54bdde847211f7a47d
za3ed4fffd3fff32f7012a31ecafbc0d64d8ff32f3779692614f160d1b1d1008186e2563ac6e433
za52db73c9d2f771630bb959de212f9e5bdd9bea19995bf024070efb8abbacfa8962bebf3ac5aa7
z39c130924c787868cd01efe3858796a4f955e12ee3c9286f9cddf72a5e4dc3454f768b1c24f33f
z89f68599069795b9007594eb8df6e63d9b86fac9ab54411cf1e9a28232044456c7bbf94878922d
z72ebb89d202a3ec1f382ddf0a63f6e8d0f06254ad87dd05a6368950dd79d9a09c9a623d1ea754f
zbcb98bf9ccec4afa264e52511f8b5d543c8313169b679d0ccb1dc0a2b5866d35456202822333a4
z9098b6f312b524b53a5dd5f0640a679df800d4166ff6dc502f5b54323ea0ae7b323d0ad483c5a7
zcf5bad7cca4c44c3de5634b5049abae8cb210168916518e55efb6b5dde59d518598c1dcf56d1b0
z160773b0d9b3ff6b1f79845e43690f730ca7a41f478f78c101ca55033ecc434e60fc49d394f94d
za2664fdc50cbe7ed2c6d91bf29b8bf7d97b8a8c926f815e5d4595257585ea68082f5225508b6bf
zb11c63cbdea16e591591a863ea624d20402647b4b653da966bbbfe3a11bbb956859e80edb180bc
z7bf346068d30b85a4b33226db9b570101a6b26c4bc751add36f704ef65b5bc88c62c47eeab4436
z01626bc49c50cd0e6ebbe47dda6258102a0db89c2680beeede35391ef66168b255b154c3191279
z7bc4d2aded47c18db75572ef54533484efbf0c24602243bd20c798106a64884b0d50f30cef73a4
z7aa1bc55a2beaeeb297a0c01b1ed80d86b86e6c713c80de58fbd252a3448751f1489ed37386588
z391d0b041755fda7f725e412dec6442329d1dc2aa7af2cd2b10d41f3897337473900897708d1c0
z9b94459f8fe88e4a035244cff735cfc706fedc83db8ddbd0c51cd7c1c38286403d5eeaeecb669a
z90d2c4013d1bfd18f8caa7b733c2462ac074fbf1e120f8d853ab9c2af16e9409c3fff570e6692e
zf3a509349084f176ff4ccd6540a37a3583252eb5a1f046010b929079d99184a0ab49765b79a131
zb968b35f158279a9aeac4c457160d36cb4334dbbe3b3ad669d85e3512f14be01c33dc98e46a630
z35a215704a835b1ae8adcfe8963586b3c2c69e6f7f194e2c2ee6e2080f114731a46c3da21b1127
z52f6afa904539538f63be5e81448d08413fa758b5ffc48b29deb1934f1b51d1351a24d4085fe2c
z290f60de370c44d28bf64e6f85fb1ed63ea16b88da0089bbd6a3ab82225e1c22e95619c725fc75
ze27c906a533e14fec0f1eaddaeb268d918159cb542573622ab82638c1ac6493a2ee7fa3de4a715
z28adcb9c131428079c63491bd5c5466ae994cd405a1039aae07279351bf443cbfa05adde226923
z340afba3f0daf136d9bf82ad5541302b5813962fbe548adca547c6b58d802c6a38ddb7242bb477
z58722132cdb3512ec1bba28703a1506d66313ac6fe73553791ccfbc8ecb4c59672d6b20f58713d
z4884cc7638586d29b0607933c120d618390a8b824af204c5aa11b966810cf7c789e8128091f922
zd954686699f2df9c9b549fef3c2aa2ac308d471df4336428088b970929ec90c6932136a408d1ef
z924738042e4d3522b54471fa24642c6aff1ec4e54c24cf45dadb47a7afb5ea9263bfcddde78dfd
zebb8cef4b5dff56c01a56861992a0af13072e6225c219daa71a59ea3ec63e7c19c89dbe3a57eca
z30fd3b92e838d016097d555bf877ebb8891d3423ab13c99556e087b4d1560042d74b8e59e4b16d
z83d48a14d3d3c3ff64f1b3eae98617b2604be9440355b46ac0f34c257ca6cfc10a0ca6754d7feb
zd387878febb557bf2f2eb15cc602f210fef71053866fd1b1a340ee976b5998631ff9305a019340
z280341d2c71e304122e18607857d4107249727ebb2261c3560ce746767ba25ef0e27fb470755e7
zfd3ae7b5aeeb6d875f8bca7c88b0d55e8996178991bb42552e458b9f39edf203eeb2e660d3e1a1
zfcd7f4f4e06ebc948f04f27823dfab72c2c653e7fefd4ea829515c40cf17d261481429c5d6ff76
za73fb61d318f6b92c30d50a90937c3b0e260bbaa066cf3ede8f1452744840a3e92a8116bd49d47
z3aee9e939bc532ebc78bcf8feda67aa394d506362dbf0f6c53072a8cc537014f0ae75c04308f5c
z58dd127c0e07aeea01bb7908d8c7057ef4b9c50f5f5c6f20526a588d7bafdcfaf7e0c86d78accc
zb4bdb31f040d52e987d98911f526837fa7e699e3c848c76ed41fb004dc5d931ca6f1fa609321c8
z715d1366c0a9319b50fb29998cd2a27435e01d23486165806eefc6c11be25976d0efbe16dfd8ff
z4c0c3219076330bb55a919c93fff9bbad996e51654075935112796a82e2fb8a9e285bd552420cb
z565992c2f5a9e4c9a2977db8c0e9a7ebc7bf0f98e598afb796c0c6615f70500f13fd7c8b99e324
z20f44d789b6105b61221d432759fb51733c240f798b0fc9a116a2bf726e7b8b778743ecceb6990
za35d8a94947cea68fc1a54f14ac79ec21032cd9a1fb7afd16bfc253758f70d
`end_protected_0in
`else
`ifdef MODEL_TECH
`include "qvl_pci_express_10b_8b_decoder.mti.svp"
`endif // MODEL_TECH
`endif // encrypted_0in
