`ifdef encrypted_0in
`protected_0in
ze74c34e226135848fe16db9ffd31815111b6d7fb642c521a3f628cf6da949865580b22efd062a7
ze90adae0e65e66a2c36a587d0a790699161455169ed55a01f2084f11770a774ec4c588039b380f
z6de9c5084882a40b79a175f5c2114b2b6d78b070cb806e1c0aa9258297f4687ab308bc470f0040
zb0b1de382961eeeaf2e279e1462520fc31c119af8f2b214846f56c2b3cd2eadbe4099496abff18
z15cec83ec4a77b868344aa20ba7360908f5c0de2a79abf8b3534b883bb12180f68b5d4beb444cf
z3fba8f13afb0abfe8fcc4294810f75afe452434d2d0f1166236c82f76edf1e12979f04bc35693e
z32ae028996dd85737a8f5adc1ebb94f39c940246e887647b64782cd7ab429b0544c173176cede7
z01dfb26b1f73408344a52b7e1f117f12bb9c8077b34876c2e6fdc085981637012dc9754765e1a9
zc512ce062e0b8fb16a214591f5c81e1353b900a611fe1f4886b57940b41b7f2ce99a7b84b04b90
z916f717e73bd10589c81e207ed77ec660a8cbed5b487fa50acde1b055c8870bd8676023f21ddcf
z9c98cc47cfa2d654ff1365d1f45035a045a66c5dfa8279050262529d2cac9e64fd27d9c7de62a7
z731bc808811ded9016570962244887f98fe5440167bd0088f2f049df882af501358497c3b28776
zcdc5426c7f52a851c35106bb93e16fff98478405dea402575c9151230dec03ae58c76f575ef850
z0b8dddbf9156f4e428ff80985e94bed62486b602a882a4a30e461afe18a52334ecc5953e7cf9ce
z5debf2a19a7c03f48f15a486e6e85d4e7174c476a99884b05857f3a012b0a263c8826dcccb89f8
z4242e89d1379ecb80b9183d2c39c7912de7a6201464eef5a3163135faa9171f72b68919d60b5ad
z047630d624aaf8c4fc3f355d8d2319eb7297b16614c536a484b38436764df38dd0456c0a0d263b
zef17a97144717e86c83b5d016837f671ce9de93c3d473e095106fdd079972b2902a798dd811002
zfad04c5f5cef1b4badfcc1440dae5f7528b1adaf59c2cd49a56ceb57fa3d15590a334a798d105a
z3960d4ef90bb8062ee8f5f6174fa1f87b389f2d4e69b7ff694d8dde018a7e0ca988412ab1f7107
z756b81cd25f2eae72af484159d3b725b3a92d4b0a9465a6ae33866b7f3a7b8a19bbdc5701976a8
z359cbca50447858523096a893b7a0146ca1baf8626074e711dfb0794284a5a78c0be5af9b30f87
z8124122ed5abcb712d641349b5a837d3ea2b864ba61f710c51ff785fc694ba1ea64af281ff533c
z66b0a2e0f1c5b37660d07dcb96d61ac5cdd581da65ef86155436cfc9e7305eeed13bfe2cf40415
z6cdf0b01fbe2216f02de6ebfe1e5d2749bf07fc764c1e4b2d26a23028dcd2fb2b27d4f3a2c7b5e
zd6e09dfa846777fd7e8ecd78e93eb48909538d6ab4f0a80583a5330ab989b3c177a1d55c3b1ffd
zb34e2b3bf96ac112c257e0d18d08b520d3f03e7b7a743255e8a7a5229f77ef80657c43283168e7
ze8653e77ad9402fef5eb98f2fdc00471e9f7d661b58813167f877a629e1b6b02251a2f597bdb21
z24b1e45feff8d04f9f6392b874e117f6aac39dd707cde7e736cfdd76e6dd26da487693b025c6fb
zd187b498b3062653419025bb897ff85e797ece5477f04a982a03c619501433371f292e4f5a2364
zb3a8b9e5e814a4252a99ce5732cbdc56740fc6cc81e69ca44929d292767d1c555b7069a5de579f
zbb531707817f99e502c3b4474b2697543ea9ce892421a62d14466102c7c2ffa434028465f5f4d3
z5dc00f7ff97d4fd5aa5d70c38ca4c42d3d7b12a9d50a6c9a6bf111b3a77ff97401c16e0bd2e08d
z96242fd716df704a329a558f49e53e676767df383e56f88e8fc1a5dedf730824888542bd457c2f
zf5d8d6ff081afc85792bbef109d9e243b9b9b375a24bb9a361d629e6dba1879ac1a731f292d603
z569328e6c2d9fe3d3f951cb94f8d52206b9623401c1dca50a70e8ad4464d191636b13c3cdaf1d9
z3451b52e872d14285f2464556caebe9e443dd59f387e5770ba66404eabf8b16be618647775ed53
z5b13970fbd31e0714cb9a22d31f7d823f9de6106eaf56e60041c11323173b90fd8e9a5a0fe1371
z075c581a1e7e9b41f75e51b4923d272f2a5ba716e35b020c26aa47673125f901c3f0719065a934
zbdd9b62811cfa8fc6b44da16c3187f33c8a04a19eb438e96b1b1002ff3a947a2c955d8c6c62ea0
z8797917615b463e23876253bbd697f25db7a713823ebc06ff0aa3ba167992973220918e4faa3c9
z635de3427aa6b36d37e200f9205bf02f5b0e74b563a385e885fc6dc0d4687b80cc75b3c67ffd1d
z88a9147e8eb423216fafffe51cb32f1bb8c3f95073bd92f96f4a7eca163cc2e36007865e151ac8
zcc48a1ef39e125adaaf0b09b219d4976909d632b751b4298a9a4a506794bcbe3e93f098ed931ca
z172e30f412438863a204f0e69467144a466c81f11139b27d174113565965603c9299d0b47a2e9a
z144d036cb1fb76cb990855377fa2c59b195272441e546c8801252f5ddce59d43a3c656818602eb
za882a3ea14ccac41342f17d0bea78b1ca5f1dc37106e614460f142699d85eaaaeee323824752d1
z0362c9ce2da2d9a6c57752dd6805eab11e8e62cf9f5985a3c39dc60f2c32f85e9b554535549b1e
zd46ece467675ccf3e9e85b0b1fe4556335067fa5b6eb053fbe07b9f59fbbe19f54133b3fef8f9e
z53599309276022ac9c7a0ece6570e15df1bc04ef1b12d6d1f7b8006728f7e53ede573f94bbd656
z661028e5f21882ce169e5b0f3e0913ac9c93cbfc7a5dc445394de7499b6fe873d1f89c2b837ba6
zfd01a1081b7265d5eaaab0a182a9c7c646d87901fbc9bcf5dae48a86fac2df8e7e0b216557e502
z7a48a10f047da51466ef3bbebc257ec1a00a182611f1a245a183909a1aa1168cdfc8cec1bf105f
z5c65380ed9d2bd05cecf2a3f6247f7210a2a5143ce45e1a497cf6a7ac0edcc5f6f88b398475e12
zba40ad789db816dbad8b499b3a455fe097562055e0f04ff7639af6ae688984f3c8c3d1ca383d59
z744c2c9faa210d7e904a28eb5ba9427236600219e64558341af0c317a54b360d6b144017fd89cf
zdf050850f4416f0ea37b5352abe7c583c7b37b5b7d68ad0452fc383c33d30d3c09ebe6169661b6
z078e1993ea9a0f1af3821cfe282105d74ad015bc1d2e9ec820aed23c977c6f1172095caa2f4196
z7fa5cf9c0bb476afdad816b2e5e045a7c78762316b91fca3c7bd4366fb84d28873ce174eff505a
z8a94a66472cde3185c502e739a3b780407a0d042cde8351d382d0c72cbe3a647f38f8b27d7ed7a
z52579e5dec91695b47ac94a122f3167aeaf498f9a7456f270c26877e244c8f010a49c667a8fdb0
z6bd0273476cd64f80a6ca3c458193e3c9c6aecb555ecaf8591f6db56e98aa4ca468ec66d4aaf94
ze4b3cbbcb3c508ab0450fe2930cd48624a31c65a5a0e73882ba83ec5fc6fb51036ecb718b49d7b
z7e26a312e623fffa16269812893e27476a0fb436abd6ce9bc241cf91278428d87bd19058823887
z051c01c7f8ad0fd9c917e2313790048e20202cdd5f5506b6bfb732f70fa63b76f6ca54d21ef377
z394016199f1e19bd66ec6b92bdeb851332aa9ca92aaab48c65c94b3b239620a9756bdb0e656ad3
z585ce749a971837e2c994608c6d3ed492464ff42b9018b05261d6988e0656d732a746d9fa7ddd0
zb35f692274e5b71a4d7252c16834c8e7ce887ccb743a5baaf871a11165464f07cb24114002ee72
z67bce17d7198041cc308686ec075bbe87db61c5db8bd49d45263b9b14a92662da7f168cf56fa25
z60ddc893ffa86299a371c1233e88006148b31efca522299b783234afc1ea2f7525b1b011e65176
z28fd677fb9ece6cf4fe99a71199e6546d21088a7ab9f81346d1661f03c3407bdea35dc42c21178
z2ac165db3439425be31e4278941f27f02fa5d822ff9e2bb6279562d9d7cafbb1e81d79ac20d1ab
z8afd2f5a84f647706729dd18257e9da6437f7cd45107e3b7b1a172cdd2887a0900927d7a843b97
zada2dd666813c060ea4addf75deeddc3442d1ed8f6c40e2341e7ac70018d25c335992014e7620a
z196632caaae18a9dcc0bbef7fd3a0c5a3c0f67e5d7fbc717701d7bb40a36fc1432306aa68205cc
z1a289416ec50a4cf21a8253c611b7c8d00af4b0ad04da263296961522c2d08aae9e3b384e293b5
zea67656cab7286cdc1b0a0edfdc44a5400b6e10bd1be0b88233d25b612e00f6ad2eb48e16dd906
z70fce9f78c2ac4652b348f7ab80ae0b964f32554eb3558daa554e8ef5f4ac2cad997eee7bda52c
z48fa7b6ff863bcb6ff90f284ca36e366856cc47dee947d08581cae2b617acc0510cca52e84e961
za40b59b7854f9f2c0f9a8aee1420afc7b68c5fffb92a836e80d838df01dabecd1629ef94717ff0
za24532d817a4f641b617da9340ed15bf8fd96ed1f3a9360c80b8ec5284c45362f33e5925b5ba74
zb2376492f2b5072dad48752f7ef385c380605e75902266a68a1d0f20e1192dc8c6b5eca824a314
zd26e66a2917ed37788dc77842c1c717563dbaa55218299e2b7484e357954385d6284cd91dbca1f
z13e214623c5c186b3a095c29893181dafa42c4013e4180064017083a3cc29fd57eb87eccb7da79
zb84843b981ceef7068facd877bf4e00d49dbe9cbe1303a391d13a16984bbc841918e6add0c660c
z2c952eab4d608990813b6edde5d9f26f8fe5e87244b2aab997d66fc0ab76e31740dcc1faeafc1b
zb3eb05c38a8dafda25bda74bee7e075bb08d0ab3de5bddccb459d9f5c5e7a709cfde57d41f0465
z1ef331ede9b00f0e0e68405a9d1cb3c0536a0b94ff19ab8a09bae113377e74260867c484bdc463
z6d1a25547031781f7943bfab8b1354f5394e3411123453036792375c018c4a02fde8bb6921c8ce
zcbcd96b3cb7804cd90ac69d26c0c317c937cf887f21afdb677f85a110e5ebb191396e8c858742f
zf8b709a12dcdf902ed50597dfa8acf8c0816aec07732893bef4324ce775fd5ca34a7242f0860d1
za465e0986d2111ba50a6022fe076e0c40c652512002dd1fc9ab1bd59419609db2cc030447ab2f9
zb35ec946d45afdf94a53d4b912c35f3f7ff9564627a6af604cb047f92d1c73a8714709933389bf
zfe7c6ea14515655000f6690c30097216cb82949d6427192a99165259033b8da3eee6102dd67f6f
z4125bd39bd9ad266d8ae28d3abaff6145ef6a16eba366b846d8060a899968562b0bd4200baf182
za180948ab24fbd58a493931b4395fa75768291dbc2d1275d660f9d5a0872600ea3533e085710ba
z693459e9eb4b38a29dbca0ec6f055bfb58c6908d6fd090f74c9c33ab512d50157e9e49190f67f1
zf6585bc3327568fd48eb8a0508eb72b4064644b4b744e95e5bf6f6b91b945629922c73f914b867
zbe8ff015bd21cf67bf9a255a8a8e74fe72feef8bb2da381549598d961dcee08440bbe493811042
zb1aaa1dc7c447368eba03db4163a06c3a02259123851db0ea94837cd2c5c3f013f63da37cd6009
za4799caceeb89faa2cb42732e1bb54477f37d25dbcd08b56d6465d16bd9077aa92ccb66df0d479
z1e2462e980fb94152e07eae4e8acc50ddc7a48e6d0785bb80f17748c0663dc2466440ae0fd3e9a
z8ad2a8aafda56e014d4ba383cf454c7a0cfdbe990eca3d1de1ccada49ca8c38360857dcd6a9ce8
z9fe77008a72bdd4eac0973fafdec6b64f0ac2366899b93d5973ddde59566bc36bea0899d64ebcd
zf9283cafc5c1b8dc5aba6fc0c4326cfef7fb905584f5950c54537397da2595c7ded6c023a3439b
z56d85d85502c6e4b28dae86d3fc322e9d7ac20f4b6ac7d325f9a1c0017fa66cd820d7cb185f81b
z78a19352cbe4585cb610bc80fefea23bfde88a3e16219784536059621467b497c74d697304b981
ze65256518335f72b3432e33d25d229e75c54fe3632026cb9eeb5a8a2a9b95e2a9d040ffe9718b6
zefe1ea160aa8ece8e85b7fab2532c81dfcbc2906546b5cd862b7f0ec798ed5799e783a9af6e8b5
z4424780ca9119fd0abc0e563963789ee84dd6981d1af634a151a16150d9ab3cc50afb35bd63f06
z1dc90297e17a7446643ea9f1c332e6ea863f835ffb971f3f351a2a0923b0b410fb24cba788b535
z09ec6cb14669549e2a8e8e4965aa2117b4d4d002a78662483df7a7176de6bd2c52e78326f2fc8e
zd11d59c18646ca56f846e95916057821670d7280e78627796bfcb478a7048db2be72110d3971e3
z9672619f7dfa8fe917c005affd3d2f8f262e69023a3715e6edd3ff69691c5a72182c349d2588a2
z03ffb82fb984e95f585d853c5152a0516a8078c33372fe27e38101429259ee3146f70638d05511
z59b1153335fd54a665b407cde700dafae6595482699265a13126c60dcf843a68a6a1262c218d0f
za652a9831689ff7612d9436b06bd67336afb9ef1f64a4fbd3c599b1d7be78099fab89604bcfa05
zc6bce8102c5ba28582c96d26ad4b051a97df30930c4ff7d73d59e9df646dd4ff9e3a1ed8ccebf5
z44b3494a0247762e8ccbf3fda5aa4fc1a62f26b487b17424638d8066768542cf3a07cbfa7d689d
z38e47fdb5410d08ef311d193ffb4ceda0c85d1e4f7f98067d7bd2fb4465b6acef087ab78f7a4f9
z5c1ae5c3e1e44f96213b0fc55198a8dff8acfd1669dd5323b34978136dbd4c81db0e21bd0820e9
zae9260fd18424c1339ee7116d0ce020fc7dd24e655df77607d64366a494f176766e75e662a640c
zf1aa2e62d42dbafbfbf515f61121da3f9e275f8b4880e30d6fc762c70a1c882ab836d5f297d792
z472fb7e416887f5f9de972cf02af10605aae4b62989ef6c97a7bcab42efee71463d2468bcd466a
z071fd3419e31b375d650acab1d98aae63a9f4ab018650cd02a8f68798c05d477cef12d0e757a7f
z5496465a7118653d9f7a1a8759b090b971918e74c880694d41c5ea256df0e6e29252898d69620d
z4162987112a55ee74466b985832599a1827b88e0069342536ffa6a53cb4cedaad655496d6fa607
zfff1dbbc03ab3222dadfdb9f90fa6291e6d3f3900d6dfe7fbcf2eaa96e95cff406c244215f7afb
z7d26746ae7399e64f578ded9fbccc9cc459a1368f87f9f1dd92310b9c7c0a1992d9b817ea24917
z648e0523718065b7674ee58e8fe58cb152c5936dc1878412e8da5291a3a951839b9999f07e3fdd
z1231777c516396f74a2e319b08229118dc510ae9a51c4a2a44749dfb1fb8a7b9477f8bec2b7be4
z381977f2db432441eb815d48485da8f1ffc8892aca3693db863fdfb27dc50df0e975d83ee42bdf
zf0121070e1f4d93cd33bde3115340a743c50fb79743afed648cac0dc1933bfc868ecf1c790b850
zeacf9bc40b3bb267f6f2178df23874fe86e6b24e78dff8f995fc7001407ca1e3ede458c0fe5286
z171c4c5c058f5716aa1ec685a58ac27d47b2d7440faaa7b3377148d9989014f41e951fb4e65ae1
zef07150ac65366607c1bcf0d805c1d225296049e801bbd02b95f50a637b6eb87f4f50963de7448
zd4f8d60d82be2a6fc5cd6743d7740da2e3dd9652669704e345920ab432b9c07ad4020f210d3203
zf216c970f6fcf275ea437b7fba43797437601b49e0759c3bcf9a019553fa5f531b6de615b0b94b
z1cd18c3454817c0370b96c99964a85fc5b17e19c0589292df0b2f641081bebac543d176ba3b488
z25925ee5b9f0dec8d279065d3c2ee1a3afedd47a628e155d8773a90d6441b954c09ac66a963041
ze7f3e390bec2cf2e567788bedc86575be556fd24c1d9b3eccf03073aa24cf63c7f96dec3a351a7
z2bfff769bbcbf94588db23452986cbcdd4dabcfd69ed42d7abdd9936043d1042ba21efd748c9be
zb8cc1990eb7a0712c8b1752683e7b0ef7d7c3a7f726c52741aba9870006270a22ece7ade905516
z2a6d94bd190560215d9b5b246ee1e41ce8fc9963baf97f8353311db7eb7f4f57dd4675891dde99
z2f41a44d6ae4fb35ee5a98ef922ca35f28c5487e9973f574ab0af0362bab83d97570a584137c3b
z71c292c20bfc99f94a181c6525c5989cd361a0a863e9e6ba34477fd3a6823ac4d6446929b857ed
z260e7f0b6c3e0b41170136cae3bdece34915f6e155cbabe9ac3e285061ab4ee900425f6abb0dd1
z5af856e1a7ab9c0597ef4dca8eccda39c21915131807f33927c87eb7e0b4b6c16de599e7e77c78
z38a75554dd8870b9fb1e23e07f9c31fdbb9d7a06f84a3f740bcfdd4315d353ce5853d276922971
z72469e0a17188e98d85e56d6bd77576c970b972fb1e5c470dd414e6c05f8ffdd4758609e583ef5
z5d938e04c7fcd87599bb7fd8eeb632dfa5c1a389b08b3f486491b773c21deaae7e8a9863331a16
zac470ce403cc9710cfad201f1dbda36725d62fb9dff3278e88fd40e61a023295799706e341dfad
zd95c9f9068ad8b9561c5fe343a822495cf7fd21309552432a82e8f612cc06873221b5e5203fb48
zcd77d0cfe1e39ddd617e533f95f671d823451021f33454c38780331664853c119cae332bbad69f
z8e7b2624ee440ffb41ef098d2c0a7058aff557473ee7ec743de08e366457d4bb5e9560b80b8f86
zb5044213836f0603748c60fb800b4bb2f52603ddf788d20c33176ad8e007f8a8b27f4d56f092f6
z06dc3a12a066d76403a67c7da34ab876d5d1cbb4a3e0eeca089a411ad74cdbae8b7a77e4d23470
z63f67d4da5bff1b54e012b097524d13c01ac88f76ed60ab0dee0eb3b1c335b40ae46daf5b13dab
z92549067e2fbc20ad66c0260527773947855cb438c111d5c35ea3cefdc50ee064926e0ae2de675
zfbd6d63c2b905f77d64484a0af334020a815f0b98080d85164f976d07f1fd665064232a5c14610
z422635e483d9167085ef9b962c4cd33379d9bc45c01b3d37ed970fe21dffbdc00d3237ea2ee52c
z1a9a556f76dbce7c43e17426822de933d26834e1a4d99d236c6c0e85adb3bfbe39afb2e001b0bf
z653a448dbc02f6fff34ef8968b06a0ed3e9535dddd09c51c378d22335150dccd9341bf6239c345
z10dcbb8b0c70af73029caa8fe0c7c768e237166198ac4aaf12698255d5987297563853c3be8cda
za33c84bc888b5218cd488f442442a3b6a0574f70fdb040c6208925fb97c6555ff7bdd9e8a1415d
zcd72b17bd24a880a9778e471db532cc5595b60d7f7360d41c988fccf0a107272f292c11b9150ca
zec8f3df1ef73905735f57403e6d9a79b18c4dfc709ce9c01b00767453d0c62fc1651e7588001d9
z1d2cbd6c034840e07a8756243dbaeb29d07652bca4e47ab66df3d5671b17b29e7e2bf4e17980d2
za6b25bd70c1c52451b61dcc9302ba44f5cf427c8099a0460850a0c39e1bb42aab06802c55493f6
z9e10a72fb36708f603633b4290fe078d85e958f367f64c16ff6c9afba5a529f0667f993e204271
z8a61206b6810cd70542a5861a415a6b009a801d4716334fd71865204d0d000b514d994426f34cf
z4b4884b5ac6e7f1b46915e61ad3ca44972dcf47f6d8efc7d221eed004992c966ce311b1fd2ec4b
zd3eee076c717b7f96caf09ff8edbd39947e45d990cd7463f9669bc34e624946a1c6445532a836f
z2f908d5a71968bcb4a10844b51ee03053d6b0c86f7abf1cb1c50bf9bbf196c182126ba869c0d7f
z69a2743929c1bcd3c09c2ec8c3a8a934d50a88d1b665c3dc89cd13085eceab4b4c7b9ecc237ada
zf90201bd6a5d8c4ef747db55a58055629e27aae61a0dd7eb24e15da139acadeb164f4ad792c064
z9a6705815f56f1b5f092f0b0ea72a6548000d8ec126b7eea0c2b4abae1e67d5717bb83a87c9adc
zf8fcfa54e4d35e0d1fe175b470b087020d169e9ae6e274e8e9ae5b5e768726294144cf1b73dcc1
zf0ee9352d2b6d502499595829cb3c2ee3bd233541786778b85c7c880724a88798b804df0b6e77b
zc12a189d0689919eee55b43d4a3c8c6fc6c6c15633a3ddbe19d2d57959d49dda593441d4508ac4
z5532c640a406ec4fffa4432ea2e1e87ec92b2f4f82485d4811a3671b90b5b13005bb8e4e0127a2
z6b3026abc71703421cb16155ce9a2218070c1fbde173340c5d5a6d3a8c7ec4db31243fa29a99e9
z5609885e0483cb15783e1e5f04da607961aa86ba6b2a41f375d7cb5218e3d318e8d608407a965d
z08852d656d152962d036f62f6bb699e3f052c46adc9a08abd9050fa9a6926b3f46271b82b0d011
za70821355a01ba7581e6baa09761ce7571e91f56f1ffa9ad8306449b165be793d6a74b4a9a576f
zaefeb39c8828dd65f827aab94a8a8cde492dd2db217d987ed94c885a679d98363075888eabe8b2
z0663584af4de8a0b3ca3ea58b7ca7716959790c9b27cf8bc9b7410c2fdb78d1698c1dec76d199e
z8fc8a8577bde3349eb3c96406a3ac8455feba6a7033c794ccddf49f56ed3d3c22a35bd4ad9820e
z6993ce51069d9623bbd7a0b129f02889e8b20425add7dcf119c429908fc0cf339f4d9fa907f648
z65e5242b9b0730b65acfd107a18dd870e705b1b815d3a81fb045d3c19a1bb9a9426e164ebf56c7
z8ea6bb0965c73e78fe74168a9ee3402d91ce84238c6a4d37476e3a6fb5e9d924a740417389efdb
z47eefb0edbb4f5485e96e1ce3f3226bbab38a6e6082e7aadba9081a98eec93b114cb7f8e1f2e8b
za8213e52767f01f7dbf8008c5ffef001d8509acb2e3645168c362d95fa64c610344f087bb95fd6
z7ef3475c4edb3bf93bc4ae760a7de6f23cdbc41d399ad92c5a3330de8af98dad93ff6ef5e8ce92
z1b06c32199da9dee03c1c8d2521efd220d33c17c654d72835943ad22ef9c09b66bb9cff6cc8af1
z68de2b5506e088a0d18cb19402b023e243a1201695a6e612038f730f9085848b86f318b48e1b2a
zc1e3bb9606dd0aa0ae170e29a57b0c235cc653ec6681f104ca90b488296926cd6b9c6b6842f060
zf343c4f77c05bab69bb906aa291e624235e25d310fdb0a00e8bfa890cafed75e844bfc5f64fdf2
z6f9848e74f48d4a42bb3a99ddf84ca6abeb0e40cdce2803f60da9c55cfc0d1e802a7736d47fefb
z15be763d8a295b5636341380bfc355196e779f1f39c97e65af27d595c4cfd3c8729ba3a03e6ffd
z7b5fa566d200bbe836c369170f576f1039e44e11482a30d74f308b205261eb5477cead40981cea
za3b83271b38d1ae1887849e4e6f8749e54b7d435ec23e5bf08b09baa97a9d1ee8a89dccd9a966d
zc2ad11aba07c837de09d533a9b8acb7f763c0d291dd1fce14d3178cfacc3b253b9335784769c66
zfdef846161a65bf4758a374b8ddf9b07484441af8c1aed7f8df61ecdc58c52e688e5fa3e3bcf39
z7b4622de5e92bfbc17d58d14632754dfbf1b40c194dd3c7c18aaa46aa7e768582c7fbff22820e8
zecdc5db8da277e140e9d6dcb941a6a88bf5d5304d77ba2b02badef04d83af688d76e36f33f4f12
ze4799380aebdd55f296b94b7b509837391e53fc768284cd62d96b367e857f948263398a0cea463
z797e1322fe22c3a965b47e709bb60009cdb2a4a174174e736ebb5e8a94d12acf527a21ec19dc39
z88379893489740f2bed0660d62b765d76a43466f606bb98b94d9bdf9b30ca414f6bff42413f0af
z81f35c5a32a02965b90a92716562e93b1fbcb00afd3f481a9c0675fa2811c1b8030c8f13e3b630
z218e44db292fe483056adf7133e985fc18a10abf0735561dd3f3bbfa22afced6fa1c95d20f7a06
z72746d0906288efdac9143f71c207e047b6fb36c9cdbf95a246195648822bea247667e7637162f
zdd9ac2610fb593a9f328388f82e2a2ef940c26774f57838f9a1db22e3e56c69b10f0cd18dfd764
z397f7ce2c786b388088a5b4dd850056b2546a93cfd8fcaa0840c4896d0cbf4e4bd883100d0ae24
z065af5e3dbca498447a9f388b7ecc6b3676a05865af9e160639dd69575a06edcb2aabc96b0e69f
ze0288a6b190861ac6edcc95360df4c0749dd463403ecf8c3fc97c15b9602ae70bc935a762a22f1
z0c4927a229a389e31c5c30d4e2fde63d72840971f91bc8a6fb17252b126259316053c330aa3ca5
zaf7a9fdac7f3aed52fe7ea49bdc438b88871ed0036b6899702769ca99355097fec678c14bae5ed
z61225ee3da419de6e479ecfc57ad2fc4fa5a7b1a5a46d172d7eb9441272c6cdf70ea372609d6a4
zff912614f40946d21cf69b5bb38d2e09d9ae73634d743571df881aa0ae0320f36bec9ae75d4f07
z4447670e68d8421f3b3b3f877fbeab76602b880039b0548d9eb1cee1ef8df69a996a940d77bb22
ze339839fb36bbc457baf2ba218f3bff7910c13c5a905d09d4c60d8758d58121da167e0c3490162
zee7ffba2b2fe8cd5814a044c4f431d32d62db51192aa226e3eacefdde8dfc8b07e816f49a94ab9
z7d4140608c4f667e4d688622e788c97e0a71691b07dc1b989d3118c1b019624ddb5064b79c4427
z64b5491a2b5f103bf996dc64a09fecb9760b166eaae9f4908844c42cb7fcac95b6fcdcd1250ec9
zf013d5663bbcb03f56afbd71544133e3473b7826680ccd6cea3cbeb2690114bd1f867c86b58bc5
z3c784964fe371a8604bb81a1de4ecf41310ee1e11160006d8a81d4a0ae4ec3e0e8094dfacb781a
zc8978b97795599752ec883be525fce2c7a02a7f50df20e2798614ee59742af4c295eefbd5ffddf
zf5bb6d1423d4eab975987868f5bd927e1122f7fecb34124d2fca5b412bc7abc5f015dc6b6f6fa6
z3acc1744fd77af5424b51edb0e7867982e0288f27a0c4cd5abcc949804e85fc23cbddb6ac08578
z1ddcc884bed104463d2fbb6a16f2883a7dcd8f1c24c37dbed63cbd7f74a4b00ad1798cde260760
z7c3c420f5e3fb79ebbd6d63d078d21e510812d6dc813d4091f91126c5445566dd3e2cfd1c31441
z545f6701b83b34db2f227bd745cb2866f3264266fa2ef7230adf7e25ce27a09318eeedadf40398
zfa8c6568b04d15c43c6c663963c484023f3068f65e9adf16a151545dfa0a7751b238ff4b6b45ee
z7139ad721f9bf97326e06e36c33acedac89d81a261c4653e5b3bdec58815811ec3eba100967b6c
z8b753f77c3fdfe887858d34527844f13d9ee8807b8ac9a677a63de33d240d33750dacff26af9bc
ze04996e73156b79dab649512ed0f8f527969de944c979deaa10b7f7197a89369f34b60a54fdefe
zeb495b7e74d49a4fa6669201a291304436f0a9d549e34d15c4a391de2ecaf38640960b33160530
z465b7a1a3cac71dfcd6d15ea012302eb5736469da64c8b50dd4e55116a1f3d7b1297b9b0ecc7bc
zde0d2825cb12b4e48507bcfddda2fb2ae0368d30e310fcf3b0c5de5b30b871d9729ac33c2e265a
z05bf0081c09614a2def990115fe54e5b59e302fd56ab784c0e464b4588e1938581f592c163282c
zc81b8916edeade0ff12aebef9707d93a8ce67a1bbbaf67ca53d242bcf81ea720a2b430d780662c
zaee5c8c9e0b7541e177eb8ccfe7a922a8b7d7e17b5d7d66f19b10b307b38afe6faf06a86d41f1c
z28f29e40a01b9617b32e52250f7975de35417c77432ad3350e4437c0e1c4ab2a938690f3931fa2
zf23b39024399fc9670f4367872ac5650978a90a0d49ce1b8efaddb4188be11b7e303e6c1b461a7
z2fa1e904569e9ce89483aa6a74e2fd485213e4c108f602b6d7829a1827931eec240a40395c09c5
z6a1d1e4dadb5965b3c001205ddeb3fd7c0de9cf8569274718e18d21039760724317b728a1f206c
z7e3de52640e5d0dddf9758f1b69e7c6dcf1b31c315a808973cce385d6ecffc5319c3dd14715c55
zf5e3a96b3c6b5a4ef06aafabb06b765b6c01a3caee3fbd2388d89f7e75c4a6146e874e8b00099a
zc989e30ee1450f359567307ae906442a35bc3ffa5d42663f27a234c094e7ced3618e252f7d7608
za1455fa42cc5392cd78022b9bf6ccfd31e9fa9e659d5dbb7c2e64a0e563f85f803adccd744edc1
zf9d74a2cf73dde9b5a38c8ee739a708f590eb4cd68735c4f644ac5453d82831f06c70e579c4afe
z657134d5050423a6236259c66479a7ecfcfd5264cae191d0e31bd3b49fa24d2058d06d7812b863
z46bc1c0bc504cfb02a79ccc027ab2a94e229f22cf64a6465fef2acd9731130421091894c009828
z5ff85f900da4cdfcb4cfcad1bb26d6b43549adbedac2fe528f5a91c996bca86a26509739c54995
z01893b278367a9e704030fcd7b83b562d6cb6f327959ac4b0b583c61c582f7ea1bfad343d71b51
z46a0fc489db8b7120f17ec46b0f5dc3b4b1361a1a8e7bd6a5a6f9481df77b95f05cb3d5ca71fdf
z0de108bc2d5e73dc9c9280b308defa3b1fcbf37e2c22e980424aee19871ff7887b78eec6c307f8
z676b9d883138741b1003021cb0f57c91a80a74ddac2bccefffb28b95ba2d872f063643c20028ea
z19373c114f3f8ef1906ecd6c97b706aafef56f927c1f6ba1b8a5406fd1086cd8e4b532cf011600
zabbb08cd83e58592c86098061769a78103d5c5df1d68b651fba8843b7f15c64d890bbb6f5c8d9f
ze568db3903c8334e49a9f68fb593a4afd3c6cacbb3a1dd632501436341808312d04e2e8cbb6790
zef8db04f2abfcf8fb2f323c43941d82061e2a38e2f0881b12f809cb0ded5559234e2a08c32fee2
z8a106daeabef9b5ff099f6cfc602db5dc02d46bf591a02874e0bd76304b4307c4401eb75fbfbeb
z7cfb99fd0012984f8a0a971a9193dd4ceb2ca5ea79e0507096741ff6f0cd6a252c86a5a81472b2
z069d80246f378711ab9d512d13ee826feb8a073e0280d63f8cddb257334b99df9048c39aac64e9
zc2ba75d2eae9d5c5999381d7b2d00172cbf72d758b66235aaf6febb81b958b8035e3de71239b22
zd2a49c89a9ce0e1810426bd3d4ad85edc12e99e16147466bc5a5b18ee778b05d1be3166bf696dc
z44f27f686d9ffb70258c4afd10ad78ecd61805aec50a4569645ddc844d39e5a96e61938c24ef6c
zeeef21b8add6dc9bad3ba83fddd6b506c3bf6a166d81b54beef6bc40c6dcfc5dca13d6bece5da5
zcab02e79aab4bddb8d120ac593dfd739cb80cfd2e9a55bfe74cd7f2819881c62c3db10dc34206e
z100c7249a278f12a5459215450673095fe6f0c4789f7247df7272f14c5d18bdf9f156135bec554
zf278c90496fe490f05cf12b857ede88303794a8047b81d76b7f89e4579f490dd1d065ba06e9f9d
z2e0beb44302cc13cbe905ebd8d47a0d3b404cc56138c34c73e50f88013ac92f73afbfb1978dcc5
zc722fcbfb6388101b105be62d84652d5ca5c745f4d72e06ea6f3df9066e8a5786f6aae8f7cb370
zda5711dea7b625766ebd27650d81f2cef1eb84b91eb1fbb1bf7a57efaa33c38cf80426947f08fa
ze541cef2b3493f3f3eff430e534c896c8e7b7967422622c94c4c2ac4b6a974b32a57234450a9a1
z2ad919e2a6e2cee2d46e40d71a98757f36f7fa846a3156e57c66ffbafeb0b535d1c0ead517abb5
zc9f3e9d8336e12b9de19d5fdf9aace7c9b1a37b281130fb1fe54a7ace3587457aaec6a88c1341d
zebc63aa7554ce713788b3596a8e66bd8f60904d56d21efca66640325efe0b8bbc65bbefeb34196
z83558b3719094e1ea261068f087f5bf3d25cf6beed1613121472ed3984bc4e01c01a5b5cd4e455
zf56bcd1904b017000719a7ac2c357ce89ac3c25a1e8a5335a753d34172975f2915979ae3eac8c1
z5705d63c4860ccb4bb78480ff13610f2bc053c68210f50ad5c581cda45dceb0e8daa02530b645d
za96716f44f3b14de53d3c7ffc84088cdea2c7310efe07968669affab6fb18a1b5085c884502081
z240646d3319b3ff1439d39b226cb9d660836d43acea2038313554016239f70a608bfa91740510a
z358d7fc57e8ba8af57ceff94c386d3b0db4672c90ca257e3edcf906e3d08c85ec1d1eb6b068502
z8ed05bb0a7c792d09eb91f662999d2714af0f42753d5a317781346f4f49d2e40d0fb256bb554aa
z281396a9830261a358884fdc558fb36056f6045d69ae38aff0c0473eb96b92ed8aeac092de4a01
z67547e819fd056445d661a06c39d7e0a98e04a85b9aacc7e5b9bc7be627b3a364fc6cb8e638245
z2abbedd89fc9a46ff5ea309f240248835cb5aacb412c11543473da4ffad7cb2b7408f971a5af81
z0fcd206ee3ef8bf59bf546063e5cc993f53f4346d95e2702f1a0a4b3f1a03370d266762d2dd0da
z92850b48b1f966131b4d996c7b4bd6aeff8a12b4978602edc51d39cc1e7c400e22cf99a6708aa1
z4ea2ca89d79b5b7cfc40c29875a3b7fbe30db1b5367591724ac233165c8bad0aab05f11cf2cd96
z54a250ed4b0589019de55ffa24977f3a5e7e97264e8a898cd9455074d9618e87086b96409b8692
z9e5b1372689563c66b76a817c70456c369cfae7aac1f583e699f490c3f33e53ea647c86a34e8b9
zbbb192b9ca23a6f25c6303b4f3827a0985d795a2178b418bf87880c4b86f278830206ff4834ba6
z405fbd09355abc40b74a64f3eee09dce38f24183513acd4d05e7e1c3c17aef221abfcd3e916203
z95003fdf4e2aff892a5d124f254f0185b70ed684657a30931bf8b288b924ff1a7292121965366c
ze5fc0d94117bcbd7e68e358563060f8f5e97b519856366e7f0a370e71a5237fab9b5929b977b7b
z79a4db3577fe4cba669230cf2ac8a954170f466392515096f1129ae659b4df18982083722a4ea9
z02e3b63ba342d8a6a0800287df3351d25297911c8e2da8659e1d1d7a076779aa1d33c5bfc76f16
zb6b7df072e83bfaf3358a4accfe90f71a68134ea00469be9aa268282766848fa5f6c8f2e1063cf
zf825e4c74155365a4d9e4131eb13eaa2e036e4182566d788ed851a28fe446335e26589e659fbd8
z0d23e1b6499f598e68fa1493d3f97c4c36807151a32e6d25aff0c62fb2c48bff74c11b023b078a
zbf9a917536e1f05044729e5560bededecf0988841aedf33b7c30479f85ec20b0703575d5e9c9e7
z00
`end_protected_0in
`else
`ifdef MODEL_TECH
`include "qvl_pci_express_deskew_fifo.mti.svp"
`endif // MODEL_TECH
`endif // encrypted_0in
