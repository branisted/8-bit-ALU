`ifdef encrypted_0in
`protected_0in
ze74c34e226135848fe16db9ffd31815111b6d7fb642c521a3f628cf6da949865580b22efd062a7
ze90adae0e65e66a2c36a587d0a790699161455169ed55a01f2084f11770a774ec4c588039b380f
z6de9c5084882a40b79a175f5c2114b2b6d78b070cb806e1c0aa9258297f4687ab308bc470f0040
zb0b1de382961eeeaf2e279e1462520fc31c119af8f2b214846f56c2b3cd2eadbe4099496abff18
z15cec83ec4a77b868344aa20ba7360908f5c0de2a79abf8b3534b883bb12180f68b5d4beb444cf
z3fba8f13afb0abfe8fcc4294810f75afe452434d2d0f1166236c82f76edf1e12979f04bc35693e
z32ae028996dd85737a8f5adc1ebb94f39c940246e887647b64782cd7ab429b0544c173176cede7
z01dfb26b1f73408344a52b7e1f117f12bb9c8077b34876c2e6fdc085981637012dc9754765e1a9
zc512ce062e0b8fb16a214591f5c81e1353b900a611fe1f4886b57940b41b7f2ce99a7b84b04b90
z916f717e73bd10589c81e207ed77ec660a8cbed5b487fa50acde1b055c8870bd8676023f21ddcf
z9c98cc47cfa2d654ff1365d1f45035a045a66c5dfa82790502623b57a3af03bf0f0c0d35b51558
zb8b5f2d29acf03737a9ca2a053b7a8f06800d50b465c41b30eb585f62f3d0c2c5a43bc6b689d29
z6f9564726ab95535ac6754c6d32cf62f73715354535cea443579f83372f451d4891d21f9297de5
zac1a344658e86f3f27ffe9d728c6a706e7710902ed73b2a949361ff13dd2940cf08d3b74372b78
z10e9ffd80ccb06ef3c49fb8765e3dcd1d2aa1d56a0f08be82e23b6ff148dfea990cdd46db0a72c
z6d345f4e4494cbfbb8427d53eed12459334910b5e7b210bfffedbd1cfee8ecc1ba9703e3053a00
z5cc9cda3ec2929308a7d986fb13cbf0041b4334655dd2f82a61519bf5b5978f5745d14f87af2d9
ze3425750db54545996422f144e1f8ae65425e46621c3506eddcd8a6a2ef333b157a8239de3f7c5
zea14ffcd4421d5d707082a5095ee433e16fb3c1d6efcee1c13d3320b54254f59fe6536fddd230a
z332af825d4f83e3e2d16f04d5273af92ff551383e99f26438112487d0228984c6d1b9cf29bfc7c
z880597221594f4b4f83190602e50f26c3e447d91e8acf0cb0d79ff7576dc175346697801ef6a28
zebd576ff08586c0e08ae1dcf2f004362535ebb999f43e57cb90b3354ac950c3236926f45a4ee81
z98523faf87843abcb9ad7660d3f0c7fb3fb8eb67530392fd9393b5b81e47a240dfe09c41f93559
z3bcc5a50d663b2d463180639468664adc3861327fc7d3e20fabdab86680d27f415933d79059055
z9621060005e64b412351f087f69fc085f843538f3fd94ea5b0525bae527507870a7e73f720e3a7
z5afca04917b9f4ad11ddff4baa71041e67b97c3befe69d4cb6d4632c324dfceb831a01489d7705
z8275f55289d601df552b9d6e0545de2b2c35fe19000c9778df0fd32a3ca1b12ccbc392ab47b785
ze670299a43de0158535aebca4b724f362a7bba8e89e299eeac468561a410df4b5f2deda739c595
z2935be88fc6de91d760d583fd1b1ff3dee6ef27358c8d8fa3165b9676b4c72e00be9af82cf3de3
z04a076125d144649567c0b10184c31105a7694408afa7b5df1f0aca54e16c17939504768246f30
z843079935d7d6481e0458f846c22baeaca1b5f4caa17cb71d1c9db32b176b8c2a968f246ec833e
z5739e266d8c3233f15c39d924349630d6623201efc96ce7db68bb1657b926231c19a916a4d2d2a
z68bb6c56fb27211c435fd6b07d9a3dc29444b7111f16c55ffe1d9a084df9e296f70172aca24d8f
zee28dcce2858243d47d30909912c038141c28e1cb00c828168d3a3badac989cc5fde066f485933
z0b9675d007d84bb9a9ba27014d36d57253b360fe6a260f27e3c9f6a7b89196bfddc5986e6d8805
z1e8538606d4df311ea1036b19308ec7e8b7c9deb02704f71a103ce18703a7bbb779f5d1a8f03eb
zfb2fdd4a8cfba079f2fabb4b19a4043d580d8661fb57b0e3d24e563eb0c5de7c32854cf5cfcfb6
z082f7fc464f75762c1c6322daa9b87320aee04847c282044fc543babc3a5d57d47bbeea1fc0606
zbd14c910203b09d750b2a5d287233f71a470fade6f05c465f73ca5d4377fbb509d1eb5115d7bc3
z06544f83c5c9e973bf97ed83c0248d6143e5acea93d36036319dff4accdca34fb75662cb099772
z006bdc2c2966189e1b8d3d45c7e94ccb008ab8a8d5cc285b76a926fca380f617d6958c7a918b56
z2a2739cd0ac8a3106f777605f48c43422fe65e0bda11eb78898325c6a45f7678cafaca937f7d13
z6a8431e6120b01669714be3d62bd98fc7a3f1db3b1d6254abacf51b3cc09a064ff4a0c51a6a261
z710d6bf1fe4fa6942a115737f31cf8d8b1357bdc175242c297eac0833592f753fc776403b48e66
zab2bd7e84ee20d694f11083b87077f09c321f2c5c52d98757e20530ab6ece06c149b5346f06445
zb8026daad08023aabed366337c0f2163750a84344bfccc97dd9f1874376befc51933f369192843
z8c30ae504a12de7aa2e68aaf2da54c165d42e83bee321fd3ca8b333536d63a953efdad2c777960
ze4dd6127945d8aa7db897dbba2e5132a38109313cb26908c0f0dbfb1fa1e45fbf66a6e37056b5d
zbad364b891935d4eff71a721ac059c313a1bf43386ced0b58a6c733d7b7cd581f4d4efc4de3720
z84a132fd4a91535bc974034a6b8a90f5ee11391b1744010ef1b2b3502d290c6b4ecab070a245e4
z4d491a0ae07d338580f1ea9a5116eb4f0732481367f6ecebabe683b8520412c549262b8df24ebb
z70980a7685c1b71e9bb542a89639fe0a74ef9572672850e69403e8df9bf9eb58fcd21ece9380c3
z46ee21a24ada2f9151cb6fc72d6bedc0f642987853705798b8b3fb704b0200afa44e89d2412372
z411b1d7da4092d8faa58a0bf01c106c7fd678e7f8c6d65721f1845b53f4343a05f62a95504e40a
zdf7b658efd1b20442667cd8c138a660a2817dd48c7a70594d23a6e189def95c4cda171b3303798
z562d0e62d3d98fb6dc282f1f1dd11999da416ee578e809756883111dca051e689253881d5004c8
zd2bb9af326adf6cfe5857217a3616edbc48ac62beaa893cf32c42dbb7aefaf5bc5301b7265f949
za72f2dca55542b3149786665b097168a205e9a72ea6d4276de018327100c56ac6e9bd484c07c42
zb9e8ac13050b8de9810746d09da973736982141501db1005c99354a5e84770f12948b974765462
z3b0b678ef26be8023863bc0dd7e96e52d7f11c8b33349d0d237181a96a396bd11294dd59412a0d
z6eb259861464aa11f1f7d3b0c15446ebae1c4fe456e5680ae3f0fdd846269399774f36900e62ae
zced148b84ffc9f8035e60647e1c2b1f96fac298ab41741b0dffa788bcb06d80c2ec51e408c87ac
zcc1fa73057aeda9129cdab725f3e3a8159137a5fa2178745fb1e4247a391296dd2e042c4bb7f9f
z630d3b506fd0613b01d4e68f61ea70322c6ec7ce040491b676058e222cf5a3edf18ff81ad48579
z50a6447923ba0eeb7e7012ec2fbd66bff1decf3449ac899f0c5b59a4ee8c74095bc4176f00b98c
zc3242a3957777c8d670c5c25c19cfbf9f34a4b05459fb43305fd931525689d63e61982e8f87529
z42a194814a50e32de72039361574c012e921f7a8a88500885be0745e0e6f92c8e05373d35f4345
z2c6cf3516bb0d39bbb737fa0bdef61f192522d7f64a3fd5c31976c01320179198d52dbe408edb7
za4726be73fb42c1e3c9b62a6e8916b4bef16e21c65a2dbe331b26ac5a10f61fdff1a63e1671fe6
z91842ceb3a6b8f7261c565ae86e0cfadb5a56f7ede33e99bb6f9d6341ef290478913706de1c50d
z1800c2242721abbd833ceadefc33cb88efd7aba6bca3c9ea817262e49768a5e7f7d52db6c94a4b
zf0f9981f4c9523459d25b23f92589a46f7dd5905779f6e2196f340742b6966b380950813925988
z0ca543d756ba9471fc2222ed1f190b476e284dd8af595e71b264e2a6b07f1b623cb9a746fdde5c
zf861682fafb5173371b619ec3a52dfb9a7c65ec4bd263b2a80b5379f98bc7bbbf17c5da13260dc
z3a22de9a5a343820d2b94296ea40d056066db26fa9bf9d527aa79ef6c216e1ffdcc1d68b278d6d
z2686a73886a2dd572128af355c212da8ed1ccb4dd447fc4201d9ba0d5f27623eafad951993e016
ze674c0ca9c022d0fbe0d4fbf24c6244a549188a57d86192c69391f22933bb4ed9acb13bd9ee642
z53e0023e5b3555fd2a491f077ee833d714d35d33d7e0d35dbe8fcc7e20129c3d5930659f7474d0
zef6b0e01b3008a66606aecfbd483657b2c45aa304fe30f7b53af3e3b4590bc7eb59b797dd7ac12
ze13379b5d8576e5f8cb09ee4dd6ae3e8308272d3b4707d982e78276f983b1964b034b9f6ae2fb3
z508c74d55a05c97571f1e0504843793fd545736fe9a707ed6d4f26c27f4e89366324d35a716314
zc7af3f8412f7819cd96deff1bf01ddea356376059cb0e30c131e5062388465d80e72a19e865c05
z94bf2ccef534e9e9c32d2a47107bb6eec80a45b5572b1e9c9cb89704a6d5d037a3b070737676d9
zbd106bafb9d150e7056d3694c56ce208205a7a2e6e90ee55ff3da97a058d0d26f53f484bff0083
z49faa10168c7bc698280a90a01bbf1c54570bb3e05930a9a821d5917ad268efab1321648cbbeb2
z9bceb61c16650d7fc680ef561526f5e4cfc2616dc959d0923e2d31b8b8c6514463bb7ec76add25
zc77df87dd4ad7ae108986c62a648e7e48839e0fc0f39bf46d84788211de3ba37826bf09a755e35
z22a95ca7878c1ea498a42beac26d354e6f0e4906db9d118eb5a20db6a85d9e01eb2a8db54c4e27
za80a326da5bdac341ced5317050bae8cb41aa88a9063b7f58f49f7488de162afd5760e320d0b85
z2f2477394c8d0fcc3ab00d77ad094578bdac44783ab7cff3b92f6e4168871748c37e91b20f59f5
z855e9368f0ba9efe77a1e792e21ef0edfd6ff690f88dfa6d451b02ee421f1aed942c1d1c1ee5d6
z01d1c7077d1fbf9d2e78fe6be1ed09de682f5e84a4b0b01f49bfce230acdfd9129a137cdb41b3d
z196cc79cae327073cb4572db1563beac768e46e4b569946abf6b33a1d14e3cdded355d67bdbc0d
z5e4c28e5d4a2ee530487536cff6ff41f6039616ca5f4216944eabc3d01a3a88519da4f2ce2d1a6
z3466a50d0a88ea77573edab24c5cb9a80e3ded6ef4421ccc36bf5e4deac53e716ff8c82ea5b661
zf5d818487308917ec14fc4995f7047ae4bb6be821b42349f27c543098d415a83719410baa6c5c9
z82db2039c18bdea3cbee8082a4868c19f2b0906d7819bbca62969d76527591dadb610f611d51a2
z11a10e8a875563bba06790e94967e47adc9f75bf8fccf4dfbab885e4fb609c2324982df4164fc1
z0158140fb45a7fb91e834974d411d4949cefbdf246b1e984fe67c586f1edcd8667982657611f50
zba7df75d5d1e5b8b6544fd2c1af62fb623517ddf188316a44c13672276aba9272ec0c212002e65
zfd336eba0c31c558a7c24fa9b2891dc6e91cf0b15d94ce5414b1e6435a22e06184ab17d9c44cec
ze65c63e6cd660922d5bd3ea5385453cd133dfaadb48b85f768160d92854fa1d31c4c6181ab6e9a
z809fef2adb2e02fe914621695e2274d1ecd616350bdaf369395dd78f917ae057841b0489181045
z62f3f02a43a6497de8ac9409a8d8ee9330423289561772691e68d8b701cf292b3e65aeda90051d
zebd72f9da5bfbec8d317669bbc4271e8fd00966b0f731c78914b66a6d3f0d41600d67be0907f78
z414bb4f68366fd2a4ea53d0625902cdab11ea65c7da74cfb9d36925a20427c55f93497f7fe7c0f
z9eff0ae6ec0a62bfea6f81e12091f8d9f7b2c5e77993f91e44c983bb285e76f31b18ed0ad1aaff
zc63c0acc5d3afd8a2dc54761f728d830640a464d5bde3283834193caaa9baccaeafd7565c40264
z2a47d4d5818c929cb6ae710d89a375df190b0d8fae8f0d1f2c7e1797715cb43a62b3c4599fd8a6
zb9e09fd2a9da1741fbe2b1ded737a1d47680d1ad855e5e057cbc205a74952e6fe5f0f0b75022b3
z99bfc3798f329eb078c51132f88ee38e743dbcc9651b0b7092ebafd1f9e210dfef70ba8ee93fa3
z7733cb8c206d40bcc562bdffd2a8e8d4ec49706f00469692b16341afa6a1d32a3e7ab238b07f2d
z57d1789e0e529fb64140375311099ffc0c0b967180cfd91888de3506cfbddbfb4bc2ebc41c5bdb
zb63f87c84c82bc19c5f56440596df2fe72a0271bc3e79908e3fcfecb2546f7c3a3e073fef5a021
z7dd5aadcbe19b64d29664443d4c149e301d02f7962e3448e6c28f45c7a20ea53cdb6d8e80190c5
zc1f069bbc7ede92805043b544b415cc4ba3736f8193d0acef44682c9cdf97a175209da493b194d
zfeecdd66adead1dfe675d8b45a035808d0720e1cc50584d6b607f7aefccffacc35b41c2ba1c76e
z2acf412b576a5d01abcf245a057fcf4aad346515d979083712d5eb25c3d97aee79b6551aa018cc
z5a7aea0e1a733b21de388cbdabb34709be83f47a1a4fee76c5ba473b66e417ce86d355d9eac10e
z3313f7877e2ceb4650467a589724500fa7f4b01867d77a07a0a693883c1d2e665b7c82678e244b
za4b1b9dbb19cd6917f2361942f32d287030cd9d196704c630fd67eb21a3494ae6a1122a853cd73
z1c1050242132d1edfd789da9181649720c4efa5ba71709ec992cd0abbb9c1f29938e3984427a67
z8f2a5556eb51a8ec3747ab4df0da7d23ec616dafe7df3fa2d84e234bee3ecc7d14d7ca2ea45fc9
z70b3581959f951a0a23a049de49be763ec6ae29868ddb6baa367af13292451c735eaf7895314a6
zbb118d12e017feecf7bc469f9d44b49b7796865d06514f2a2f544f2472847a58e6b326953f7c2c
z906c4b6e6a808876d96b50a755fe5283787556f4b54decfd3324af4042df571d2ab58cc389c31b
zab03b7882e71bb2a96737ea0bd36aa55e2278e4f172ccf28b1fcbf49f244615b386b6ad3c57b7d
z372911edc52c5ace68453594a2c8be3c6bd71a9eee115372a9d0d3e315c913d7f43bcaaf21a46e
z4eb5e7ed5a1c3fb13cc71281b8c87a08d0d56afa1db7f9e36f140fc7a40bfd824d871f8c4c84b2
z0c45860a9d081115ad910450bb6589eaaae20315bfe15f0f01f1d4dcb8ab0b93a3cea3c6a18119
z007dda11ad19130b9661d845982e3a7018ff4995cb1d152b42b508e39b4da64f0adfe5732669ab
zfc20f8ffddc0d1a380445c738b5d7c1ff6cfd610989343ed9e92a346baacab373f79a464e908e3
z52434de4ed548ff6a02b149a89f76c4051aa3cb54f05064a888941f658c2cadcc4843b5c86f231
ze83f5424bb75061d9e874efb4eccc0026de611c57aa9c5a3927ae216b3a10a571826cc72f2520b
z00524fe38eabad52606b3f79410c428c0d6d21e112c4c852fbf799ec978ca6ec38d9fa92128931
zb00c0b5c20c5ccf2cc514685ca7ec3a69ea62cc2e6cff293bcb0c03580e195166a519a6833592c
za032b150e31d41b286826cc1f45a6f27d47c0b92d156b2349b901a12b74d253b4a764c11a05373
z6ecfaa1d1ce9ed7a8ccd2d7debd4798a166479480fdf75237ff8b4320c03035851032f98ac2fbf
zcd348de7317a1279916dc4f5452bb0eb197af816db85363c8009b9759ce464b4daae1aa536da5f
z5cd06f9de89e4bda461d2a7df66f78f3478181d52544d0de7806f272207e2c21b8c9efaa332521
z1acb4adb4955a9bdb4c6232795ab3809ad6d93f94d2dcd22b261dcd1592add076768d83298fee6
zcb0e4bb820d736afa54693cf1e3247df06a945feeed70e6599d67718ab75b18f008a44456ee78b
zacb481c5ba577205d7473606b52dbe46aafed8b89d102b7e2d61fa3819530587bfe466dc9dd9d5
z3f9fd6af02604b715c7bd4c1c56ac4d77b25535a7259f71ef9cbb48b3ed5672296aac5521238bc
z096a73bceaa04606bc627d58fe7b885ed7dc167871c744de92f6f4ce57cf2dbd34e5dab8b812ad
z72f58623b9985816fb587132bc3da50c432f7686aa3480e17198b95157f7f08bc020a5ce3ff25c
zebadd03a3b23eb99b1c08e2573add79eed6677552af22ff278ce4a97fffc45b6409cdb7f7f510a
z3f552e8cb9d4405b6b3036d066ea2b3c6cdbd5775c3ba9e8f0e8877957b4ed84188c5a62e25865
ze1210797917439147fd375f7155bfc8f130d36f4eae150a9886b87bd070642c542f6e9627ccff7
z0cdfcf2b62959fdfca4a395d74f2553fb341ee5f034ad4b9361a284b2a772304736b6c0a468068
zf8a095a2ac47b8cbf4186651706f6d3dc44e6530c29ffa436c0b6a0cb780009b515834a7bc9c37
zc2d9199b38cad84acdb8b31fd31d69ad38a33e7605402c569af480ba775376927c8c87a2b9fef1
z9fb78c82ee6818ed29ea78ec81a42622ebbba545ace2ed3ba1879a28cee38c8e8d10a26dce7622
zfc3ef55d8be8d40d83b8e741133ed7f5038d5102a274e7afbad86a6a7e0e05d213e70c1e0df1d6
z3e6e57bf995c60b6bfaf1f4528e85c274bb848315391a833317fc466cb9a772e14baca4280c06d
zc9262e8d9b89b7ceff9809162d4e9678cd878a4ddfab48a005c20018d9cc0312a630ad178da427
z75e0ff96193b7d3481b8132c19f18a0099bf8810538fc8bdeadc7be757e29cb2dd975a1f538155
z915405ae1e332b83307277b674dbc19b68788ff04b718b7caf7378f043d03daff859887c93ba66
z8ca151305d0e0b18fc1bee0c411a091a7c39f0472127aa3d73e9813ca6ab2a2f43592d9ac23800
z6d5128ef5ccc344aa1d3aaedda757f684e0d9606b8853a4278742469c157c2f92bf1883c352b79
z587ecbe1a36f7bebe2fb8965ab926413292a9edb42b1ecb4f73accb0509260646a5d64f6e96171
z0bc6ed20748bd23048e1b1672e5fe4887aa6be83044bd0dfc87c35ba13aed9b63369fc52ecbb31
z1ab455441dd1dc5ab5f6026978f36ca4ba629bd316e06b88539f16b799f5542714bb8ac4fe4547
z2261b7b951cd6d46e88efb1845fd0c773658e8df96cdcdb104d457932a683935b3f0a3d93faecf
za55b96f02558fd938d4a94ae3002495f8551c87fea537a9a03b7eb2fbd95314a089f068b13ed45
zc3ff91c8bc5f8961a9cf0a0c84571cd5a5b8e5ecc16eef28995b027b7a4007093e3ba5b5e3d884
z1e9b42fd01a22a98c0761cad926fafa1e7e8f2e6e93fcaff57ba12d7fa6b630aff1e9fac474899
ze47de828c14708477d99580927fb32d2c8b654ae0c181a1e69ce3c6ff464eefee354b0274feac8
zd0461d0a67fe29b52fc3b8216a148417d0527a5de1f69c35ef3ebd444792ccf7c89036d9d56f0b
z89800f187f98d9d5658e809ac80f9dec326731802ba28f78a26132ad15082071b7f79003fe446b
zb9e5eab674ca956ea8fe3a2b994d44d05fe25adc981c9b052fa97cf3261c7cd494fed018fbc373
z3f4c1afe719aaed8082ffba144ec7dea0242711db5812be79de5846a00e3f8b7ea6c1b0c703a43
z87900725dc3851af7a0a2b99e9a3df0d264d52b0d982bd4fe48a29ae0b47ad9e893309cd3e6097
z90e8a5398009d2b86d8342a77f828f5e8c3b27d3dbe96452fc0cc624ef31094fbbcfde108d2a54
z26dddf59ebe69b8f183e6de95e7047ab23dd00d4786a83fe272c1d0bfcd62325c380b85eed1f17
zd79caf3696a09d598afe6a0033bb77c988f0350394e6ae45be6c9e93c1b1cbff4da85889c662db
z6c18f30620b3a1272ab0edac5f26bd488da1d80bf0c37d9c626f1e989e026d2b4dad2b7b19ab4e
zda4ba9683685b87018b31ef736d4a7c5a4d6c33f35aaa4602377c21acd249accb428eb218ca051
zcbba75dd965043ede4d4c6a93d242f10e3266777e1e9b55023947f2046d5ee1bc640a8284e2f9a
z078481683bb3cf09f4b8d93cf041e4dcba2090cfd7eb43954193ee15ca3153b88d135d4e9f48fd
zb9561e34ff29c806f4652cfdf97d6a174cc5702f574acbb2dc7ef72a1bbe89de38646b3a28b4c3
z22ab38bcd9942dcc44456eef6c97eeb848e69fc044d028eba6f349b5b0dfc5268f4d79f6ce58e2
za32943fe1dad83043a11405310c5fe125daeff0fb4e085120e1326c4ceeccb8e26b65b650b1323
za2f503500896d4cde92d64e372a8d3d78af2b56a1a144b2b0cd6325907663b40d18e4345922ce6
z5244e2c910942ed54a0e295c6120fdda02f02df8f218f1e24e703b9bbb9fc37b66207b988fbe2c
z6448d4dae6505dd4c25a97d0e354ab7eed7b5187fec62a5b009cd0fb277025880d36b94e10bf81
zf504ffe583494fd28f131208e888a833dac4f43413a22ae86e1611378aaec77ac5c808a06698a9
z75d025c26a8ed2d3c48196c427c8255f8c10de6f147e46ad5b5ffa60c99f30515eb4234b86394e
zb08916f084ebf640168f24a33e2f2fb8bf223710b8940e61ef399e606e506b5a6c747d477762d4
zd5e01fd656e32ed23e7630d32b0801725f87aa6c92ca8868161639251375dfe817be49dd01f108
z1d9697b8a8ce3de440e853f65c3fcc6960eaddd164f1fd5514ca581ca2038db0541b697ec3e765
zf6067bd5c9763d5ca46b3ef9ec47875dc54fa28af50317909566684583a99da19c3095f1f5d0b1
z95e7f90ce2f554c2d2320a50b9e4b58a2236f23c20c1c5837fbd86d4ff86c61840ebf7a245de31
z0d2fd1b79d78ec3ce5130303cc016b7ada7da0133d69a4738946c26074bdeb67774be2a0d6ecc8
z93bc13a9e1e311093416e126eb8b6beaab493e073c25d428a4efb93f01ca29675861faf2d755e3
z15210471d317ebb4173c24e587337bf96b2d16ff7612b5653f58841452747baad46be2570b2552
za7fdcb36ddb09a10cfb3cec2c207aa1e67741763534ab0fb1bfcfac3f65db2b1c45dffb0afafb5
z9d9d45b1101603419b26289a45535f68e43c4f0b455f4c0892f62c80f40262a683fa9277864a9a
z126c34fd06916300cda2429eff263908643b5cf418b230b62ec921c189c96c40c77936b2bf506c
zb3788a975a59c61f15e871d286970ff4ae2284b482cc3743d439b45fb881ca9dc146a368113e54
zbad4d35e0e956113aea4af465817860be88f1295350bb0ebe6b9a5c49d33fd754ad4d452daafad
zc4b15bd9bb9c48e6aa18ec859861adb93f18ad5e5de580e33ba0f73b644962e48ec258ab9680ac
z87b4e1a73bee63cd358e03f9fde7e29530ea3f075b470b8ffdbc03c29d1392fc758e39f37802a3
z483c067cc7b36030af517a9e5994d0e8049d14b0ffb89110342ca5e94d79ae145b01e0434dcde6
ze953f19cf3d5db94f9dac992d725780dd91566cb38bbf20d6703029ff9093b667602bfa2e7f0ca
z2851cc24cf7fbe5b967edfc34571f84bebc56710501e8d7e041f0ba51b24435aa9a62b34030b59
z5a732bedca3fbc8748036efd406587cad07e7081f526d255501730b065d21e4c95f8f2461d434e
z239e89987c5e7184c75fdb4e40bedcc8f5a25fdbddb55752871d8d48b54b6121652b6d9ee56450
zbd27894e0286b711fceb9425c33eac82d1da08978a931770bda9a13b66029933f17876e8099e6f
z1c41ce30e9f63b1d23514576b480df5caa6e7da9fa4b60a85ac553b83ec9a36b22dfa6c9b11758
z80158586162482ef2c684b7926b7f914286e8ca7c20d2d4dee82db7e4ca6c23d6dab765ffd5eed
z4940630bb076279b72b0be5cb884598e639692a7fbd1acbbd2d57adceccedfb188451f00921f8e
z12b28e18e7302bbf523765cda7446940411fef93a1e6408d8c27123aa2c62b56727153e55725ee
zd6e3812042058d8ef3d9cf7abda149a6e936d4303ddff6e57eaf6e63f647bc50cfbc9e651a5a4b
z169a0985a52bd636647891c49e55333ffb4f284c5cab0bf5db1093cc9639b80093bcd335827080
za2dc489bb3dc6c7aad120a198844305932bb21564382689630b4ca4ba08ed72c851d4ad5098e03
z5b3e7636c7d159d253d2f9b39bfc1ee7e492abbde1870a431bcad9ff0bce05860284aa6805ff7b
z6861f10258e422ba08402f1749ebd4c1b016f6a913c07001e1918c583a22fbddcdc42014a96866
zd1ed26acf2e8263012390520754e8ccde4a40d48ac81cd992a43053080033b87ac57382bd2a89d
z16e6fb4628c8d09652011c2d67b071dfc45ec5b1f35578e346a13c5b24253a1927109658b12afa
z0df85ff8be2d9cd69df9ee077b4820528bdf77cb4d79c8cb5d6bcca795d95cb89fd840099f2ea5
z2dcc4de07a0d700b787be387504212cd47d91113ff9121e2a3b562abf5ae8bf0b7d617e4218c32
zf1eedf4f2717e138e5e63c2a2159fb2fdfb7699ae3a5a38730234ba4afabf9c768963d6b43e05a
zdd2aeb66f560d942fb7a0f3e34d9965e8744a2903dbe08bbab1598719ab58fe320d450d6a34ce8
zc037d17414e24eadc4d57656c7e2fba0e7387b3916972571e58e00353be5e9cec70959c20843cb
zb527fed4e2c9fcffbffb0dfb4e2372489819c00db43c15e3bd3e3cc890fff4805e9217cf946115
z45e42abddbfa0d629ff047fcb08c229fc20265394f7ccbef204841641c923d6529bc48f73d87a1
za136a0b0f966206f5e282d51107eb97c9c39914d59a6c9ea61580c130dc7f28abd8e629e10920a
za0243ccb30a3460ea1a81ed076600da1ea14718cf0a8a91d3c77401326cd6e7e7f208dea436500
z162d2436a76fb8516043f4f9baf0d92024ac415939fec269c64ee4054180f2113a77492f424050
zfec6346144ad57ed5fb81f985b61c5564a0ab34f9abb12901523d46b99d065e223efb4e52844f8
z5266e7f9a6b780bf05cae984997c40d23f7d0d33ffa9bf9c0abef7bdbbb57766702873fbfbe4de
z7ce08edacf9adade3f2960dbf5b8ec057660d01832bc07d1e9cc432905e5bce97b4ddcaf56e3a1
z0dcc3fde878f30595e877c6eedcc56b6bb0d47c68c3a7269d6a4c27e1bf4a4a28e16f729b3fe09
z06dc82593eb2b95673f1b69ee6f5071b68e3fe53ca8da7b4391f9388411be71ccde8182b7b95e1
zc366c0c154ca5c35a0427e26ac6e29248c8d2b2be4e2a5cd98d9ba01dd4e650291536f953f4695
z11771c5dbeffb23c1a4bd3b68c854e79bd0f2788c8694d4e7b02825474c87bb95e1c4166b40cd2
z0043c3411266d7eb7e7c9a08eea06f9551c31a36cc1f94fe3930fafd14a57368af8d6410c18f4d
z5948eeec16fe9d6959227dfaa08d025b6b1730c195b306c7afe14e0041648d95d8300dd267fb5d
za515a5991ec0464572f870fd44cc47c2a4b4e01dbe12be934abb4d3b266c2bf5305a549dde683f
z5cf742f7afcaa783d8342b05b1885964fbdb49051a2bca2c7441c82a8e46f25a5c746e4ab85da8
z2ad20f36ae71341d0b1126788bccef568e527bc1743b75939954974cfd0b60cc3b1bd5eb976f58
z0639ef0337a845b39c91681fd25f488ed361fa20c4efffe9c34364fb24a64014bbf7e806b56b35
z6da487cae16c50639b01de24cb1a4a3f501599389c7cdb63de4bf81c6fd755f0cc83e014fe17c7
z7c1c4420d86bf994234d3a457b3fc81be71c1af48143aabfb515c1c444fcccc2a264b59e54f64e
z3aa19f770e21bc2a7b27f557d698d6f0667640cea80230512015c417e53a396d55d554562c529c
z422c8d75b1521ac7dbbd21fd1dc80d1a66fc9022bcfd059134b382188e9e8d0ee8ed1edd4109b4
zb119cd5c51cde75207eefb00850bd20d63e44d8c5875da8249961a067e6c94b87c501df6b7c21d
z2197a401ef224e8848e4bd7ebe587e89fdafc772f03fb806f859a8ad918beb1827e13384c010f8
z73f5cf77c24b150d36b2fdcf531a2f9f5af99a2e9c00cf3509e85ba9c4cace8aa0c3919afb76e5
z4398207aede9a6a1b7a8b62fd09a95c4826025e9c9d5ce132497f5d912c55a487b002a1dc6662f
zae6f53f0130fb679b42eff46f3504a9263f30e1d623048a59e418c51cd0f5e0327579d6a8617ea
zde9147566f4a92ca5fb5a693ed55ae078d989865273122d9ae964dc9fb45ff951e0165b00e2f49
z1f5be331637be0798a360007315bcd6cd6c1c4506f05a83a53a177c22b612b4b54b66e54defccc
zb1685d5b95e2da6af94179b47e7b5febf823b9343529040d9f5f2723dc6b717e8813bbdcdc4b7c
z385196ecf2a3f830d268beaaf49fd8848cc603df88e99e1db6f51e3f8fcce30137653f84e70506
z72889de5168385b37a9ecd4cb70fb19380672c14c9b7f3ce7da0c1efdfcaa18b3e44c7c3a53796
z1444f4a610c8fa13e4a646a630107b80d050360e35e2cdf9f22caec844d472d826e84cb8cab8ce
z562dd18eec0a9c6f315cf750ae7a58302f7dc499d694c90139a7f07b763e741e9396c60e4e8500
zb581cc5bba119e73d4cabde5bd1b2f032430c17985c2d82b174a4372345c64cc727878ac8478cd
zb6b8fa9c442109ac244b4acc939bc0ce5e35c9f3c13da2d2c35f17b5ff4c80ff177d71a4d0bf62
zb067bd5574b0395d4a38ce5871b5f0c88aa740955ca27116adf4b52a4c7695550810a0a5ad2558
zee3cf954ec6b7e7dd6e44cba7f679cd1afed0922746b2d2d3f654165017d09cb40fd392afb4526
z8c0054d85730d67a1ce0253f8b5f281b14a695a833bf5912beaf6b2973bdcc15eb1705debc3b91
z17b10eb6bb5598f626770981fdbbc4ff895c151c49b53b660a34abce06499bc8dfb65fad0403fd
zb2d3aa8c3eb239275992c461a417b61ea90e0a7c7906b8506dc9e1f4782a0366f707685e2cb72e
z49225eaac0fe89ec6eacb8a992409d336e0c55b21ed83bdd2a876cf9ee1009e79e872366806c8b
z2272783fce10cdf8b46e5f083614748b55e29caff6ab10bc4a70cb129999da1e893d4268e53777
z4729c8f76ff07ee74f84bd570e91fd9ad715a4794602b45fcb0f2920008d1dbc5ba9309cdae231
zad79d8d50b4fb93ea08a60f814f21399221376aef7fb510c4855f5b4e1010bb9fadf39f2e4d824
z37f6bc1ff53138682d75f3ab83e3a1eaa2dc253f512d012abecbf7fc509180dd377df36f02b18e
z83d880ccc1f06e23456a258a0ec90b267a86ed92b2eb3ef2036047c017ab375637a4b7192f93c2
z282e5c07a1b3fc52437b452e0cda19c091c18bdced1ecefd79293a9e7976c7d966f80efed0d8e4
z81592b8eb6136bfd60254c77e3525b783b5da6aa15a79946a8bf8c3dc49604b385d77dd9d9852d
z47cfdc286ffd686b7a14946b2c91f70580707727da34e345e023996bb1c5cb239fff3a2152a60b
z8ac320c2ede1af7dabc5dc06b4ecc03e15baa5bcb8b4c89111ded1e9d742399b15a07f205fc734
z9809505a21a6496c17dca7f806c8be34a50bceed141567d51f8d6ee5cde53015bda3066c6058d4
z1ae192e100c313b82edd0a386fffb76dbdd03efe4de607a23b3d072c22843cdef9965a319da4c5
z697aaf4fb0e04ba2c41de5c25f8336bdb61b6b273328740f0ae04f9ed3ed464b36c5f6d1f999a8
z6743e01e3d32d5ce0f0f14398aba0a65301017b04d52d1bea8c6ee96f1c9ae5741d827203258ee
z459dd1e882fd304ace11d1b8fcd85e0af923e4556e7853c23766f9bdc2b87d4ae2f1f1c73d7a6b
z33effd83645f35ac84a5717e1f49b804b197b3150ed0f71b022f320857acd961187b8898a65289
ze5f165568fb7427928ef928ed3f05104380e2b87f7942a56aa82413c902f0c26ca3ceb37a4ea9f
z98ee0975af2da661ffd8fc9e91b3ae6945a127b12b267f15f755adf6e4898a27524cb5dd49da16
z149e712a7e81a9f3414cc65c485ff1f93cfe6133007a479d69e11565113c561c7b047652572a29
z5532f7b4929841dcf9fa660f7c5e98e3e4f308bb52591b80ba304ec0bb449c4ce71423966cbb11
z887c1b24598054c92e37ffb7545ff3140f612ecda4a481f87e0b824b86d6ffe40edfa2aa5ddd86
z04ff7c5ce3e91d1dea4039e2cd1fe882cabf925c84696b933637a869da0b058c17def81ee43a32
zb830d392fc81ccce2e535ca9baf1a05b688e14510a438e2fb5dd23dc3253b0bfff53589f5b1539
z8243b3efca97371b113ffcee353aca53393e899385c409395dab6adebeebeb524b045c384e67ee
z3c2e8410cee9c87a95287594a4e820100d8c8fa1724fe6a69eea1150b46a6c3164a1849c21f9b3
z286b6fa2f40b1350ccc655c0e75dcaf5e33722398aa57e40b7157139fd2e5c0f02e7369114e589
zcc25268c1ef1782df3194555472bd84ea78eff05f0f3eb996a36e0a73290333ae9b81608b72f20
z144806090a1024abb40b762da5fcb402b2baa1ea32816e47f27c8b328040ac92333b085e87a9b3
z69d741bc8ee90425018082f18ddd8332d9e1c65a5f982575a53f3d666b819652ccdd842ebbb58d
z5b93394c4e8831ba6d50846186f3453aa2d568bf9cd54ef7511a588b23d42785d0d2785c8c499d
zc1817b85616453a7cfeaf572d6b59666db1b7ce6cb8b906c448033c0bc96a85d24d5f28cc8b046
z0a10ddf2d16cc2bc146ef6517fdb5d8b349393d2225137e0ec4afcb7af1795838a923a650d8867
z1964d3b6e7fcc42236c7c414fcc775f0cdfd025d2d0585ffc8a6c40a887c0eac3cd9772a005323
zeea32e103cbaae8b2351e4508d8cbd106d4a9bd0718139dc3fc8b1df82885a1d162542d47cd6bf
zf0ec31eb82956e442dbb01b5a8d2c99dcc5c52540945a1806bd637c938684d6a3e72c207c6c65c
zc9bd2e8349965e8ccc7619079f77a061161a20b5e25e8b24fd6815bdc0961c9d897e9a7e39624a
zd156520fa918a1d5f5f6e850886ca5eb6e9c80e8c51602a7dfe9802b1daa78bc298bc3eb97d8e3
z7d33fe2cdcbbda5cf7498f7896873d38b5d43951178161e7d9971134d4842ca760c275643dd52a
z14767fff41254aa8e2d3c85558bb4e3d92737f5c10b2b87cae536ed48dcdb501b54cd40520a8a6
z06c02ed1daf3fdc835987693f5b025540cd97357a219097695675cd617edd11a804b965e9a2661
zefb349048eddd67f7eba24a1b925c8f7c2f2bb67d0f23a696bbfd8088c246b6df3c44147652d39
zfc190898aa9ac31166c60819c4035b3f1f609c80feed3a3bbf78c53f6fa58080cfa6ef9aeb3e43
z06c448cc9c854c4a6f764c3920ef9d7c142234f97298446799345e8b5786a04dcd6183728d3461
zee150b1e00dd16987060dcae7468a74338e1ffd98d9db5786be860286d64bdd7d11f27919844ce
za2eea306389eb9659267c32807a7359784b90bfde186ae37f671b387ed6cc10cc7c2d1ace9c829
z338c5260890f25433b39a044fc471440f77dbb5a1594f7babb959cb3ef06c47c7b025539dc1429
za9e1f5917559e8e29ed0a2093bccc9a166870301f95f7d75fc4154e2e0c8a2558f2156fabf5cf9
zd6ee4b1b84e6736f600087b28f6d779d4079cea48da3c0439c3e5a8092695e3337800fc31bb70f
z6d78542025fd013fdfbd731ac032ce2b98a3d646dd057940253364724bc0033286e39acbaf184e
z9b2296f8b7d154c959f6b4c774fb1d8ae001e27a02490303ff012d751bd60ea83d0c3053d4b070
z908fc4da0dbff140fdbd4617923946ad91a41a963f91fbfd15c0501372ba1537b1fe4a08b5faff
z9f59e276da15b67a763c968dda167abfebfc932a896a357e38be21c32e4bdf840650f49f13133a
zee10a626d03b9f2de75665c13e159effd3dff0d5ba9e19593d3cf10dfcb62ce806e355c985cbf1
za544e517868b55877a71de83c6df2823a053d127fea898bdd9690ddcd5ae5b9624240ddeb59bd4
zc20093a77014978bf8c34686bc85bc2eabb76dba818f2fbfda99962cda09c8d160e0ad8a10ab46
z2fdec4acbfd96345ee7c1b3bc45f8250c24c2af8adf6e0c6fde375961217caf1d1c11c57e6a044
z72ab7d2ca9c38f9ee281bd14e1c3a594a732bc454fcfbfa2928ef6a08b218ae9786eb2cb88ab3c
zadeb38d06d45313396c154f572018f0df89892bc974634246877680b836f7b83c0ebd13c3bb4b7
z5d4b3064db6721748bf9fb6bcce02f2c1b2f219e45a89d37c4c13c1be723742539fa63b115c346
zaa470fd876b6da8880fbc4d74acade5be7a0576eef0c8c96f0de312d0b0a546c3911735781998d
z46207bf61a4256b7ce152be03344650fdfb9523679906eccf2c4e08a63c5391a6d8a6c6c8731b7
z20a13c4dd1fa66c65f9ac66a507e9d4d6043908b931ea234e59a98ce21c357d02ebaca01a4c562
z6dc9b0ba35a0c1cc7a9594ee0855313eeb5c993d9547393e8481a8d29ca8d9a70ba16cf7654dd8
zbee3a773d4fb9889248a06ee4409e1627465fd37929df6f01e62582f15c977146f36751f782acb
z8ca4c15a5fc95e1a54a0cf9a2f22d7cb24482008af24c8ea5b12da6789612e29dc784f8164bcae
zdf2f044a0a38086d0f468b985391407da3fabb88c1e31b8e0dd4ab2e9c5d94c4e4cca0fbb6f97e
zcf8f2f735a007b681069470b40d8ce752a22903ec665cacb8a5097fcbb354415e65c35f0685d97
ze762adff663f34b6c0d39b8f4fde326cc41fa4fbd8cd57dc2666f527189b725c4275dd083520e1
z0b93d63fbe99e92a8b7661ee8d51c5781eafa17b6664c899d2ac0491d0ffdfe027d7a814d60334
z7d3d5185a6fef70261752c50ca6e0f7efa93777263c01873a1209a00d42a0d136745197083f35f
z6b165f123707bbb505d181fb72c32ff0141b1fa0b909a68ed129602cfe060c6c7536776eb5e92d
z43561cc2f7a98910447aba7e7e2be2b517f9165ac49a0c7bfcb60bf5364c4f236c48943c55cf52
zd63adcc767b7ee4299aabe1ad996454632f88023b2c84a27ff37cb1f1cd73a7d1d17815772b04a
z675d1bc58478c441f9e41316b22facaf2f23ac5c510e0c0e4413db61d0553544f19729468a00b7
z8208069f8efb1cb3391fdd809c797ad2458681fab9d450159939ef11cd82ce3a2934515de1cc62
z23e5b3dcd12f2f2a00d66f20758d7cbeaa5c4a2a25153c264d929f6ef08b4d39a1ed26ab627623
z0f0bb701504317709d488de56052070ffe1220efbae20b04cfb14394557656af6816a012f92cf2
z7645d0b21d6980030033a02cfe82389a5b67e52206b04f5f5aa54d632abd04cd9657f26bcbbbe1
z19ffc0444f65e93e3d4502bd28a880cc0d997195b5cca4298c4d0f9fb752fe402c242521aa7178
zf1072f75ba6b9401a4c0a482a3c2ac58d22e7ec74244a087af4144f743435a235a6c8a08e54bc1
z06207c5d20d36a80881df5f9fa3bf504e5ddf2fb4f358c58854503fe8117bc4424ca3f4a3c86a8
z6568403d996d9ccc8ae174d173edc8984f2882f5c23b0b4dcd9f64603b6b6b09b04c744a3bbb27
zf8d19d045528478f9e9743b81225085a67e890dfd1afcae46923b1edf2e6eb73dfb7ec38b50734
zd723ae1d0387fa1be014ba199dc572ddbfa409b2704b1e543398e2ce2138a8a17813ab0ce06c25
z45d53653b8a8e0aec5afe0a993c588b5f1dd12743fe671e8b28157b8c6b06947e3732d1b30ed7d
z447b4f7a2a488b4a28fa46fe268933e35cfcab6e3feaab60fff305ab6db1c73b2c98cf780d22c7
ze9184774f285e8ad065d84a55402f009968887a74195e85cad0da797cc941c917d6a8142034f70
ze76e7114399ce71a83f6c05e03af9abbbb70bda015b23b47eedc58b6b49dacd35cc55416d122b4
zce06db54e67a397f3994ec0fe275a2707f2fcdf68a2a084ff959511940867c05c3b706150c5feb
z1c838d18eff71667d89ec845d3ee5d9813a1b2a12746315f8207ef9b572e254f0c9515cdb9feb0
zeeb5ce350b9db2ba0327562cb1e7ab6a48a02673ffdb7ec2b148b8aaa8bfda16ac2a1bb70ef5a3
z9553812341be76dd00ccd0ab921782da75b0f7d8bfce5884ea26996cb14badd672e0ca17178a13
za947d6e62d1c44f5e3a1476aeadbf4d362f6b9f410fc2b0f65b45d914108ae68e658b343599e3c
zc42a987d94fa44537cbde16dcf0ccd9c72f45d7833915b13ba09f4a976a67adfc19626c304a030
z6b5d6db69ec556445d431dfd128fe3b2ea3f469f84c9a9cd85faaedbc80ebc52e43609beab41a2
zcac49b0cfe355472216cdf07ec6501c11c2ef30c154adba32672c86775db37b43998c30fc9bf87
z059140876ee46e48122f3715363fef46d1c254afdef2c694327f32f36a4acde90ebc527e4142c5
z8683f881da6481945fe6bcbeb90ac446b2654351039bf56ed53b472d684c4cb5b941fbf562bcc4
z47a652618e4cb8622dbd3f4caf8abd1f18839f1bdccec1dab68ce7fa60aa597369612ba79ab3a1
z9ff609c702d6fe57fd19c7efb65fe5d52d4b01c9f27caaa2a51637c2376183f70535a0d25cf7a7
z27d62a8f8b8698dee7f19b5ce364095aeaf0b924f253ff499ef2f0e1dfc52615bcc8df0f265651
zad2f3be4d1630e79eeac23331098ae56bbca801cb5fe6f0d1b518ad57ff80d8b8efbef0c063f1d
z99ec8e3f9a1c50fd8ea26d4c4c43f8c1c776469de5f618dbba077212d412a323483f0b839a130f
zb2bc52871c55427941975a77719d62c18ab7ed7b9ff62d2824616fadfdc13d1b62fa3e559463d6
z821a7ffad402e0e2ea75bd4360175ce004a3c9c7e87d7941861f2b08fe1bdf4d4fd307442dd6fa
z061f27a8e8dafd8a5beeb991ce91f8f6e83718650c99f6d903eabefca79bca80b658f9d4336960
zd2eb7b362c83305bc6bede0a4e5589f13da4e9585b5f228b790fe11149c8698027a7a8734540ee
z006cba701a6c88ad962e8b6c036344ca70103d7db9b4e55e7565a2bbebd4208a2940ac56804711
z2f3f4f99f425900abdbc0c26db97430ecbf958267bf2570cbc0e20be4d8bfbffa1819812951daa
z167d9bab29b97747a7072df82e00c54a58f65246134cc823e98cf25608fdec7d28cfd85bf9a01e
z9ed8cb92683ab9c8778d264e095ffd1ee364bc8ce42bee825e3cafbb1393aaa44d81bbea65e7a3
zf8fc68207bbaa0a970366def7fa0784691ae95c5701a4ea036e2723d95739803bac3ae6f53d0a9
zcf1f15bd0e26ef1853218d1b1f64465832a98c310adf055a4b54b9b536450c7252269e796d8e61
z8d6a3b37710e580e37c18202091fe139acc21faf65edd0ead1577a1c3068a0e44e11f649954378
zcc22efd9f6b2690966fa4f2a65e9a4b5377fa49081b871eab9cb5d54bb6aebd29e4e94ad5e0fcd
z36c53f55d5e225d90ecbb1b55ccb8a049541426774d0fff5da26eb134994bfd4c884c7035b09f7
zada5a5e6f4ea0b74e30847f9920e6d547600dfc5e4fd6f0187365c37ff5c899b3d605358347091
z9bac08822fe1395fcf0a202cabd1393542c4f983890eb1263cc640a458e1a8f965fce1860baa84
z1100c6bbb26cf07f7dd5dae54fd7888409a2c677810590b90c8610ac2cbb9408b21039c9867420
zb46c2aec13566257f15ac39f3519aefd4997bf34d3f630f39e9c7820c3405d140eae491386a32f
z8833ea2db51628e353f1f023d7bcea59857bced045f0acd159faf64c6281b63883e7b875d59ca1
za9212aaac1d4383baaf1b77cc5d425ae8ef8d27ff984e7d9c12b802102c89da5181c822bb4b27d
zd0b2ab868657bd3a1d9cb07b0fc7e6af5ad02b845f1cbc8c179a1dc6e538ea8ef1ea1fab4ab68a
zd93070504276f3ff66b9a21f52a271813c4500eb08b293aae064b3cd782df0dde7d9a98b491e11
zb50042e0d9fb8a27833b8a9df104b1c7987d7fd020e8f2bc44a869fdeb95783e02173845910598
z6f72081904f2971d7a537e48415fb0771a07816e678917a0166fea96ae4dc188e86b2bd645430c
zf13093d1c16688cd4796db00e3cd6795d8ad64bb73c322bc8c9e218debdb4b5cc4c2752e9533b9
z710f457e38b55d3062534b0fc836d341ac09649c08df0edf2ea0e97c8a89f3e72566f74de1bb8a
z899d68d7e98c1116b65ed194521aa430d265cacd59a98d235a9c0a8ccd899ab0bb6c4c20a8f770
zffd57eab7e4d9229d6b495eb6088c80fffb0a2cf184616ea2a4e4e05a002ddaae2a67add48c503
z844e86bf21d72a412eb7deb896ed7e8278e17d3d9b35e66db5068aa1554afa36a958b3626443b2
ze7c1731e0f2da01a9f1ef9c4f0f6c850298911b9e96d7289f16de2d872ae3754be92b5bab0cee2
za355fdf308d87dbf3c80f0d194b0e7f7884a9fd427fd92e0548629667fa03284f69cd88c5db22c
z0771321a0050b3a1a62fbb8bb3f602430e76bad7ff59f1f9dc965d240af7f466a79c29c4c3b5c2
z93ec9dc982c554206a700f8b95f923e9df0d8f137affea58378d79186afb8f9d4e9a00d2f5a326
z9278f48683749cb27f52cf7252d7fcc480f03e3e9711569c3762b02003e15c1a481fe2485c58bb
z5e74ebb84b3cee5bbadbbf0a9a8e6b8733a40767bd1d1d360e5ba8ef53317aa4525cf2cf107d2a
z1eea80e1144087a137fd23ec2400ea45cf93c11117055b98cb80f1a1097b76b4ceffe08d86fd4c
zac6aee609ade269e28f5b5b8a52d1f2d3e6a92a7cbd06949b2d882460f1f796bea0961a2a3cf46
zc33c8c92ffc232cc5131ece2bac8979a6126235ffa811e7fa6354a53a98139fbac47e54e6dfb88
z7de1992607050f672115e90c67e75d1663c6ae5223566c8963516098902fa1d62e765de2bde426
ze7ca016f4eb92140cfe9f1b93cc8887890bebeb12db68ff5aff2a6a22f7961caf2149d6922cac8
zc63d97dda52afb9a7dec785e1bb88fc884eeb542b47a5a9f8a5eb5c749d3a800e7168204ad9e5a
z2de48ac27e8e9ce6f51013e4c63a103346ea4efa3e57c1d3bd32513ae9a0941cfce13fd80a5156
zd901b2159b255eed08585816dca5e2524d84fbbd469c4732ab233e31b9ae1b1077ef87b33cd60c
z205f2283a6394e6cba038985b780829d85e28ad9488c3fa08a3a67298af741a54b1b9648e84e3d
zfa7a92ff2ff79de4e499167447359523b6ec644a95fed3701e2712ece4f9948fa6787f7741c30e
z0418986e94a092b10306e0165ad8eb7e62104cfb3c5c8634e22afddbbe2f41d91b604d9a7eb18b
za8cc1b7c1ad2b8f6d1115ff05e2e0ff57f94c394ca4040dbdac61c5ae26bf0bc2db95e2d686234
z3b75a8207e3c24e8aa7ab621aec8aad52bf6ec27dc5bd82b002d491142629fb82046800a6d6563
z28612bed22ef4991a2ee9f42f17276384a5fa31162619cb23505f2a426140ed31dfca6dc55b26a
zeba22b3db362a21c95c450492497f2b17e6645820583e902cea49aa2dd5628cc3c76cef4293d31
zf0b09b2aa915c6add271d0eb792e1263dbd19743f94941e9171e844754307840ecb0cd94727e4e
z5a7f4ceac241790e8a3b5324622f4c6be82475aebc1f5049026bb20eea77677bb0c710329926ac
z3f9a7c3a2bb7163543000033217c950d73df0b7e98a37e5cc28333805730153f5e4db03f253835
zee31792da3819d0b28ad095762b13aac49484426dd740fe9efddcc239759e3b6893fbde9d54970
zde5a9a9ff01ba610fcfc7c1c96dc3e0877c2ffb401e6e505ebe6b93ffa1b8cd8ddafb3d3b41796
z17232f09f36804235ddb6067baf4707e8257beba5fe418631e5fca1c1553fb51851b27e4002f7d
z386dac435820073a66bfeedf84c47c1eb997e5f9e0b0950af51245fc9f9a0da407e94c9636224b
z4bc11249338a3ae4b7916a8dcfd83c77bb7db9e4fac061fc642d36c17ce0262cf2c92381d91c41
zfd21d049c8525aa37a7cf7ddb1aa4b011a8a4e150f0e793b67001b7704d1e4ea7af0d414c376a6
z8d4b26c2e6cee714ac43dc5288d09830bd8c1c9eaa298f2ba16088b5f0b1906d3b4e0c58d919e8
ze79a9cd1bf17f204c64986ca72a9bb2bb23fd1cb10c22dadd31af2ae72c23816f0e4b2f42e296f
zc14927e869fa44cf5616cdf00942c975aba908da5f3ac1c6cdac090ee1d65cbbd9f3e9b33480b0
zc1e70febeedd01a3519ccb6f650b7301cd504e4f7c423e83c3df676ad95b7f968a67b7204fb66a
z0601312cb5ea130e2ae85bb4b80704ea831db521aee376fb33fbf91e64f851a71cbdb944d8ed98
z17158db023d65ee4241bf48949840ff3eea98ce9ff13951c0b7a158fc64b8805f4e7cbb43ae410
zdd6d6fea65b05f4fe467318b56a5ad97aadac2880d5d43ee9e37a7d9c5bcde634fe65b5571957f
zbc0058f928831e18c36d9c6898656fbe82c95c4417623c88179375312472c69d8dfc02c7449572
z9443fc37c057d6b0394f77001636c37e8489bd25a534a2c443f88c20fa9154fd04263ef78b8063
z9c854351e9d17d5f8e1c0fb16da4ec4ce49e6964c109a698278fa680fd36699fa635599df26684
z73caad69a041599efd56bac4b4fde7d1c9e2af372c9a07a89afd3d84ed592436046c67344c8d7b
z3180812c8ed1444782de262b79c6a50eb434ee9685d671f6df4fe5fed7bf0ea47bbe8fe26985bc
z1264a44424fc78a4b863a981221c921ca07fb6ed4d11d0f2322db3d36a225bb1d3786f92be60ce
ze7a07434ee21ab0c76f5d991122413ccca60ef8054606962963101f81afa77e2dd8ff81b98dcee
z343797808ead027430b9401c83770a1298ede0bb0e452c8fc3019f55c7c018db509819906f9ca1
zb0205875806ba7c632b432420f9d99d78b1549e8136ebb010ab4c86be39604ac33cbe030744fc7
zd1504c9fc6fb8eb34b3766a1fd851f8c2ed8527da085260bfdfb387aea3971800007933feb20fa
zb0949b6746d46cb1c6aef160a4a3dc54f4c1efa6601887ca1c22bf70d473261082f454a51429ec
z867288e9222be79a64466e91981cf47830c2a1500998b4a4f0a3a1869f95baa55c48d2921a8e87
zacdf93fc52716d9169234c3201fb45fffec16a37d958fea46b1fb54c5486258148b714eae06286
z35ed657338d61acf1cc36d3780fd3a6b8d4e9d9e9305107ba1b8638726f37004f8ddc8980cc769
z8b39b85dc38ee9eca570349d9b0d97048b3dba44d308815721e5662e85442abdc604524bd3d146
z5ffaa4dbae5a27e4a5bfdda076b8d803152f02e38ac9bcd8d6d0a31a34e1b96f22dd92426f31e8
z5dcf36dd333ad9b1e60428d14342732c54675b6fa462aa5aadb2e87e02919d08587358b476697a
z40f4d023531bc30b38b42c2d6a6372b91a8b9cf2460050b70dac79ab7f1173b301102ffdc1ae02
z154bc219901e59c5070809fd2d2cef77c354ced6f58396ce43fca16f51174ccc326f40ccbbe517
z3421f4d150459ebb36fa914e310467eb2184d8fc490ce3beee4db6f8b35f39ce6333be9b43e0fd
zcab4c4e803d6e6ab6a4fbaca0bd2a8f1a687e2598b8147d83bcc0ee167db1cca6c3a2c528b380d
z764dd5bb50b0780b22e626507efa94e22509156ca3b8824baf8293b9a0927b227a1424676c463c
zdbf985b1c8fbcdb5d34fa4eb1780279cd02f3997bcfee2050dd99c06ebd2c03600f0d1f1bca080
z04b51a533c8e448890870b64aa51062b516bbb2cbe526849654b01a1cefb4b4858bc4b41e148b7
z7fb7df0ae80b1a98c7117bbac21d5457c16ba197539d26e9cf4eb6e538ab75a3fb685f98eefb8d
z1a2db81f56b1c43688d2d86280898552754732f4747d59697fccda354948f91298d18551123202
z6ce893ce7276db9c2928689f289537905b5fc40442421db3c14416b06d4218f689534e820e5dd3
zf7a51e2691280cae644367f6bc32130d249e9c50d63f79474badbe48e395e211d5664c29c5e7b2
ze8fff17e63cdb9833b3c81fb22c88c66455a91f4426c4e0a1f1b286bc820fab489584afceb4744
zd3d3a6606f037e1f1cc2c93844dd39e12dfe02754265ea0c045ab991657668553b3d4f53891577
z9c5aa872db6387d2863e7910b745b26e905d1021a245051eafb7857aea0d7093feee91e8e07ef1
z672184581eb8b136c5ade2907106d3a63bee39ccbf130e30aa63858e4be354dd4e357cee4e889a
z64a895f6b47db74aa95ead6c506054a46673a2d6fdbafc8cfe768c7c0e8ecf62d56771d7f4a9ba
zf917ed183e0caac338f3bf1d76502fad689f001ca4e35b9d78330fed1941ccbe99ce52ef88fbe9
z6aeb65b6842e4f05a391546229ca0e8b9daf398902b0f0bae28778ceb9193970412c835899c23d
z969fe23d529909fa5b14038e4825193f95480c04110ce16048aa61e51c84f3718393ba2469a534
zd5a7ccfda81ac432a7581534a07dc480ed2eb8e8145f506ffb2ee229eae64e118055c01fb35f49
zdebf647cc5de016b9b4be58d978f3592c7df60ca124b8cd39e67134b04d74c032cf038b0930ba6
z8a03176a9a3c46d14ac7708a4b918bc3443e4531a9f36c0b7dc666805fb12c22ba39e37da520d8
z1f121877486903f507867cc01a9d23e67c1dd76bb1ed305278859d5c5e5d66eee376f123a7c7aa
zb7e0ce53d6f1d39a29b00912cf315b81bd5e82669409ea6d810c3bbec05e2129e6a109273f7a6b
z3cf1e1801a539f67d702594b6d9b4a91d7b47ecc80fe6be53716e31a9cb4bcb7a03a73baa059c4
zcf0038744a632ec56607774848e08f3b979b732cfe56038151aaf8926c2d26b5e7d09672a16734
z35b78be3a27020daf3cbfd0d86542fb33418954e1758fa995e9d10b0d240352455a920fefc276d
zeb2319b19ca3f1cfd2cfa43420743aae99d20de8563e7f89f0c31bad09d943031631e2628167eb
zfb6cbd9e674390fc98b1da0d6bd3ece050c957e7cb7bb5e3197811b5b374c687528ccabdc6379d
z9c9c6b8974f8d3bb47971f2b4ed54b004d18e26a068f755ca32f2d205c201a685680c540895a85
z8711e4d9e27f3a4dd1d8de3032381be7e4802fbe67e9269202a85d9044cfb18bd95fc50e46e097
zb89bc45408426a01663f1b3184e33283ceb71680f2b79c72bba577f9c0531fb8bac6a84a2f1677
zc391ec942457a867c07eacba7c5781d4c1303a83a9c87d749f6af969163fd53d4cf661d10686c9
z3e7377bb9b0a86b69a5ad58812783082f4292c39bdfc0b585204ca9329d0c6dc1a74de9508d449
z2b2b9b39c3df225c4ed78a6d2ef2646fceadb5e0a9945306495487803a64f7213f95a733937cef
z80733281253040745fe46cd7d0a4fd12072bab359be531435a9e64edbe7fd02a921918fe555624
zfd4f861fee2e2d13ae0b4c679705c263d78f9a87094d4e374a4c84eeef05357fabbebc1f881416
z17b1cc39e697eebbd2da8a066b43aae2c4e0440f0d7deb7dcdf8229d01c416419e2f725fa2f4ca
z2cc6ca4eae74a730e10cc6c60715cd9785c6453365d07bab6ff39052b463cc3aabb70edb659913
z8bac80a6e212408cc1643019e0fdf91dedd70069f23b82da4717c4905cc74458cc234635d150c4
za454a38e12c92d5ffee1f6e6c3879fd58efc8bc32bc739738eeb5f295d3e3199582e00db0512f3
zd052449e7e7d0c293430d3a539f0299e8e1204beb154b2f57bb1c59cd7e6ff744b6477f1db0c2f
zebf526627ccedc1b7acc374aadf0bbafebcb8154cf94d3ffe736641efc277f2317953f83ef39fa
zb9edd1f724388eaee10fe313d6a80a476ba24119af293899f9b772d6092ef90f21a00c62c8a155
z0605531f67ab740921bd332901294406066c5df33b36b8cd667edc3dc09c4dfa513b2f4fdfd59d
z2595b6a614127f43e3969f29456e1ecbe66096a3557326d3db8628265f86e1eca36555d8d81a6f
ze39b92e1f88aa1a5362d0c0782098e4e7812cd4f3393ccbcd6fd9f8a0d50d71918043151189f64
zf0caaf4596537915353c74980d5ff0ca2a6ce7ae521eef53c2bf33f7b3323b97072df2c531494b
z97c4c2151e37c1e4a643d2f03cac3e4e3539c0f607c1e72a9e433810d05d2a499084f5928a8b77
z026bf3bbc98f7b18cecb4e5d75f691cb9182524539f7cc6985937594693d6f264cf06e978e78cf
z77c8db27de86011d005cdc0ea028c256cf3b606cac5699899ab5f7434ed852ee212093cb8607d3
z06b7662467a3767e35e25ceef97217533fd105a13a68c27957ddc0369f1908820299041284e363
zcb2cdcd014de5ac66a6c9fd4795c55232366aeeb87ddb9078f07604bfc4fbdfb765603bd1c0c74
z4a7693f4379b41c8173e2c28e46d5cb44ffeafe17fde1fd358a720ed1810a9084c5236f074fd20
z189efe0671d8862f5a0774f04037db72fd92711f8743e576f0d968c58ac657dfd28886240888db
z3d6fe97a168b135609983fb49d93764148ff6f13e6fade2c930e537265f82cedfb6948d3c33311
z9323f21fe5964fa00c510b48a4acb53d7fdfdb793ce70389fb9cb3e32024a4c0df753cf259e68b
z56b3d58cbd77fe6b2a77997626d45b403834ace42a9c11bda241bfb95ba7ada6d2e881fdbe4534
zf05a854b1d7909031f7c560a79922d748c21f14db0d8c268e7d164015ea747b4ece640886c2a75
z1f0613eb6443eb18bf87f77ec6a06da16ec3b0a58b57ca907f7232259793bce64ffba8a9847f80
zc1a6d5d9fac73907365cd845db8ba4c188fa17960868bd8675d666d2b9ed48c4d1ef22c114658f
z50ef43bb223fece3ead45b6debcc2e569396a8b2aa4520a9a6e2b4ea1c035590dc6023cc01d5b8
z622219267c675540934d3ebbada381518e7754df14ce99b4dc9ce10e90db0a4d8784aa73f78bae
z3c8c6e5c061357c22b9afe5409f55228b76a0a8819f8824619b03ba028df4ccfe9fea381ecf7eb
z7d596b7dec4d3b5bfbacb4069c7cc9c126dfe899ebe591ebfda6f4b1ef0919b24d527696ab6e7e
z77d31b730bf4589989448ac5520ab4f6f6fcbaba5032fec5f4bdb04256613a3014e875279a847c
z2f97d5015fa1fad00a87327f33e80ada5213fbd5926fbcdc47a29bb8d7bd8566c1cbcfd2b91380
zfcede2611589cf45706c98df77623bd9ce89f416d123bc7a2077ad65506e61a6e2366a21f59b12
z2f57ea411b62109014af0ea66c9eb147f8f26b6e7b610d962b0284d6fe9450b931cbd2c806f8e5
z00d48f9b79964c35997b5f24ce7364bab474bdae97377700daaa51bb96ab9c7bcbf2ab930b48eb
zb37831d921ddb6a48273fb206a06a076379d39b7eb27430eb249fb2d6b242ae37681d3b4d7260a
z721d1378fee0b24c2428dfba2a9d85fb2f279207d60ec39445d713391557627428a76cf231a455
z111e177095b124f8b52ea3ac42d554ca9b9272fbefe5ffb22d76a421d4741b70ed81bda55ee68e
zf9dc63617ffbc147b2d432de9eb7b5c475fd2348f555f4b0f7e5b10f82c70031b1ccc555d4a38b
ze1fb66b75a7b14dea69cb3b0c5a5c466ef521ec37a304c5e25c0cbd10b51c107ad67dcb5321b58
zf367466f0ffa37a69df73986c977a908ea62a98a39b5d45acc55bdbd7d676d5928a51734abf86c
z6ffae4db34eb026e3da054321ab37d5a63e991af8187a82d11d8e993fa8f069df7e77080bd01d5
z4710f23a053721d12ff36a957689025fef636f2c87bd3b2cba184d831f460bf846ee8654a95572
z1ec39e069b50313fec51a50b7dbb618c5505416c39cff184202dbc4cf29e79a0cb1382cec74230
z9896aceba04fcd52d0d4ce933cc6d40d8981c82ee7193c6b1922b56724b42782df604b6cff794f
z3802eb73560708fb0c32449caf47209fb70fe0db9ec481b1b6db23e63e74b743f52c860a30b1f1
z07d8ad69b8371595bf0050d189fad4f01436f9dd06c92806030894ba46c9b5b97ecd3b74806b68
z1056e808251ad6dc8d7f01e150c747717a653e1b34d0d336fef6112996b0d1ddb0d0ba3133d73c
z13de4d0f99edb8af086cefd3cc12cd6cb9b99c17c6a33ee30e1734c34f76b09cd0b9795b15eed6
z835b670267843704c7b687d2095762d25e678c82bff9733e184d4896805c926d54a560eac7e74b
ze89fc10821cdc351314b6a43a25b71824650ba43e8df1a50efdc7e9fe763b1906e054e4fca0482
zbf5fac2a77485cbd8daa92d8f80a34aef6a79c5814522bdca1f2e1326ba44482dd7ff7b78099d5
z62cb0303f8418e080771fddd1d1963ba23af465373f0a42fea1874116b33f5d77244f30e4e6a80
zfa7bb8bb9a524b9bfdc0487c116baa445afc828e21956f47f2ffe1515f57b7b4007c088ee7b8fd
zecf577d1c6f6f4271429c0a90f5a8be8dc973cd6b0748e84d2dd51c45b625188ab0df1a6937751
zc0d9efd6bb396533bb883a3a25eb491a113bbf91bd1f7c7983bfbebc114aa06bdc2492fd3f3a46
zb93c9fe99ce381da02bd5ee2d3edac69b9a96da657f67ece540504ac9dc20fa959c11d9407810f
z0216fcfc244ad33add943ad8c6a1352bd7fb4b6289d260e1699cd72c2650d331e7f786a941821b
z524dd565fb67a70dc6ac23b85cb516e06654765e3bf279b5f0268f2974171f367607cff96e2a96
zcbd7a1ac17353faa2ef7ba23caab5a39880e05f0303ef741d8dfb5fb183dcaaa7dc8211ba7ada4
z5dd485f738e97704abe9d757c190c29e83bb6ca88d26c90cdc45f7ada2bca8b2896c5a41b73e16
z585a256a3836a694097c16aad8560edac39af923b3fd23b0447c633ce67c98faa4a9ac145a3177
z9a61958d57b37e74e7bef7d2bce5eeb1a8101f8cfad6edb17825c91caad2adf1024cc2e2512ad2
z9166ab4a0ba6f5617874af0faf5afba2a7440025996ac91e6910e816135a47e23813a5e752919d
z2105fedf736df0d23efb0995510a71dffaaaa24c7089b4d85f75d65660bc7b4337793e9960c7ff
z46acb1ad9ed56e880e349e6cfc18a9667341b381b7b4b8cd22987809a3d68362c7b6024297ce36
z466a75fd204427401dc5dc43226fef2068460d67d67b27daa714110a0bf0fb1f08d56a3a8823c3
zb5b183e5ab7e63708eb2e68f3661b55a3fa71c756180c1a310c04b2240c4324c9b730506c0178c
z40c59d2d50f7ece2b0f7f7ba87a6c1ed25f617e0829e0291beccf8f9804a7846c4742cdd21b856
z5d182fbcf47838fb94d29e673627888a6f5b6686f2c21aad9113cf8a1ae271438a899fb117c7ac
z063f2ef511795a3667ff270a8303af978b9f90edb7198ec0466ab6c431bc67bd28b930c9ae5308
za7d6011d2b788fc3c784c8e2d3c754719963d088bc5ce8ce61ea0831b5e4c93b60a9c52732ec2e
z54badfc2ad524c73bb8c29b8b65f681578ef75cac89c1d81c7099661f96cf4a4c883c4576b839a
z06e41b3995b383cfdc9f0457fa0e5e4f44ebe203d98eaf86aecc6cce399e94956976cb10127a09
z58eb5c860a139d0e8ea53596fbe8ac973acb690ea55aec51714a293be88c4c30d200c91e217062
zc16160aba3a4afd137af6c7c2a2cd6d5d890070c3a32e3a5e06d7a7609bc0cce6a5346da62ee6d
z760121c700ab8cf583b3842d9e27014085829d673b31a533a367e131f8547a310d3057791c2a90
zc8030c6b39e8df7de4c78f5b5759a60f6e15aca588630446bb92d0edf58e5cb88c1dc0d41c073e
z218c3b01e1ad23e4e63e8feec628f013bd0de2aba68b67bdc07e4a6b469a6c912a9f96a909f21d
z79e05f4977f3b5e7d15ba7e1805ee516a075250d446721c8369f192cbf1bb9cddf246165b53f23
zd209bfc45bb7a89de91dbfab4bff19f57fe1b4cc71cdc794991bde1e3d26c1e0057f3adaa8deff
zfab2ef622f9e55bb86bd457b45ac2d703367e9fc5689d78f0ba80a87db244386e894f2e9536317
zc38da35ec995e66ecfc6c6a5922e30c46d0c00f836c7d5f8123a8dd732f65cd39116884ca36ec3
z93a3b2f61794be5e87b6cb5a82292f8912619ff1f0b19e73cec87528e69e80f442126f02ac3ffc
zf6e47b6acff7ee5d51729cd11aa70150d940496de6b785987691794012cdd6311b794a2ac712c9
z853700f58f6f5e2f61f0ee618efe3bcee9d3aa9cb66343b6768bd317170bc037b6f4124b2bf5ff
z884c7bda0f493313254afd03555fb180155d71cd4c1e3adcf1e3ae25997e7a7263028cd1f51197
z06a8decac6b81a32d646588cfffe8e274320344e380c3acc7a7a288a3b6d3048d65e471d7879bb
zf9af833e1cdb443f1c20d7e9569de4ba1be44109ee7b04e559180e84b0a7b1e2a761a0b2edb475
z16713dbe3f614a6440434392262b4ab4ea2ccb763f58b9f80f1cc68c5b0e70174bd32db67338fd
zbe585452b1b945f9332cca893e807ae36c7a8ff5650ac3cb5df50f03d1cba7c03c58b5d6f224be
zab53b0b29ad7751e57ba500e313efbb21901f497f204205e3495bd6dfad16d0809669dd2d02174
zf96618122d4d3aaeeae5a61816d4be443298390141b786f3c939640c1b3aa2f7906a99a85eb83a
z9917e3762f856f82e7248e939fdd1912bed7e245019a995c1695ac0b43f60c332b461c1676802d
z0ad4a21d6234d1c2c7d26c9e9b01c152301039c5ada5badf5c0a69e345b13c0931326214f46997
z7b48aa2cd6aa88bd460bc351f42752656c8471ad3dfcd1d8d3c6dfb9cdb9dd9b2a88313592f4eb
zfadec1bc3d588cb20ec284e9d43fe9676018e4723afff59d881639af3fc5c6bc0460c23180969b
zcb23ba1eb0f3b051d30d2322d8078b9cec3e8d9d5e3e7ee0e6a26e72596ee0973a2bc06770058d
z29f51f33817c52d8bac632812358f84481a468eac8bc9cc57af53c0ec7f7ad69327049630442c0
z522ee2054bd5b6844ec69f2ddc2998b01c6145fe9ae533d349299cc21f66551852050f829f2f09
zb41c0be5d0f9743ebdcc8425f1320264b839c440dd6d2c54b85cf6298e5ddaf6152c26df50669e
z482ff6bfcfc598be41f5f6332cfe61f05420ddaff2acf68749802d8261da992e7dc77f3f968cfd
z996b0bfde179c763bfa743b00fe208204420ce23252cb1b892c14534b1cb14b66ecaea488b6036
ze79b261df2efccc123f8f0dfe88a003dee2a917c05b246c35bd2751d8980cf02bb78a9fd6b05bb
zf291b99ffc072bdeabf7221e97c82108271d717c60fdbfa3f6999aaa85a446942f1d944610bfa5
z87d736618e1e8ab688bed35d44332276133c6d6220f0c1013f500f1fb2542f1458713bc5b4d9aa
z07d8323d369d2e7d42f5c94310ea5c7d9ac22b122fa50550e84ed0518d47acc17a7ea990e2c476
zef2ba0c175ffaaba893717e55833038a51af6da7b41fdbdb7ba81ffae3a4687e36f082a48fe5e1
za28cdadd34eaa648239e85e81ac5e434b09330960e736fe8c60e30e8e5ddf81cb0c198f5aae1f4
z36540a6ec1b9a34a7e9487a7eddab9b8b9b3dc4873ac94b7245368996a1d0d3be0cd746f91f813
za2b7b8ff056c059c94301a38832081189db76b7577524c5539769d3a756e2075440398a2a5344b
z7e80b0be46ed4f3552f2b15cc42879fab1713094c81485c69795557d8ce448fed34e7c05b489b2
z403da1504a071b719a874b90974c5767802d9839b9df2c83b2d5bf21042fe4e4294772dd3d97da
ze6ffe19abe0b97683167f07fa4507ba14da629232886eda8b718e8628adabe63b2da1e4edc0665
z5e5462ab5a3cea4dc868acd5a1bc474da65c0395db175e8902a21891f55575c70af121ba6ed6a7
z5c6c22b80607039e912657fbd9ec1d651157466cb4844ed85606be69bde66ba41ed7b9b96aa810
z418acf049653eb577398cd46165532228c4ad834882dbf28a1ef06f6bf1b3f35d1cce4c19947d0
zadcc2f010302e19121b1eed817019cc48aca757eede17297502dce13d37769d98573ebd35c9fa7
z145d7408231fe870dd91d4313d6e949984e0d69ca49568e4ee48151ea89aa5741989545632e861
zb68a32f55fc97afe4e617f27a9918433e1b4a02328eb31eaeac5c3513534179b9ef075a04fcce2
za7bed34331a91c9a8e5b4d55e878c3a0677b77849b931dec416ac3629b64684d53dfd5c2b30040
zc6c65ecb66e330226f5450cd6949040d615ffd655513535be8b1d518e42dce1b0d348f5f4830bf
zfcec8e444c06f49fdd2960d542a3410fae0a9cb713a848156bc5e6bc32552ef24adb0cb8f49093
z4255a3e84480fdb8b82895b00f28ccd18360c0b96792332679d200435dc25f33af6c3ec21bc828
z4435dccb43a69765274c456afbfd11dc50523d37daa4350f3f3b411294b5a4989f9495f9a0f6b2
z33ea7ec8f3e964d71e1fe023ffbc0875fd72fd46011359020a1fb6046a5fb7f4166e7ccf7f5638
z1a1ec388339df8953d2c7bf732d1c81b254616e5cb380c05edd597990f7e25fc9491b134f6f94d
zfae82b2da390d6792c206b3429063a3e48ca7de31fae6dca59074346dd17e27bd42d292a1cda30
z7aa20b2cd1ac2c7187ee2ca6f6b165ddb0a5c72b2e7a5506a105709cc0312b25545ba99de008ec
ze3181145ca25f52b99cb1c988cf08a6e1f5edfc0fe430a9a7d3356317fc1fda88d4323ac33e86f
z5df36f9f6fe54a7c1f73cf3780cf7abb72330a63b5eae050815981ea4126fa7b8aeb654e7a021e
z667f3aee37d80ccb8ccc9cee59ee726955ed50e83b8b8766479441f4700da79fb6497cd1c1d9de
zafefc0370449a59a058d07120bb86ff6fa69a155a6738165f330548e4b4c406b59c6d6f68d3940
z9ce059975dfe46619dc9cd6b6c3683beaec928c5b23a2f33a1fb65bad539e92af2a4b92048e6d2
zfab21ce70c7f09015bc83d6f86c0bd6591e865d187a4e11e23957480dad2ffd7792ecb3028b3c2
z4067b4a122f39d4078ad3ee6d44f8cb8919f9462e4cc5bdbee8446871487fb1a656a6ebc27502d
z3c9dd92b7975458f3ca1823eb0d96122ac0e364111e2fd733f5f76050e5aee055f36d09724fbaa
z9080ec1a0e7929e240c0f4e1c3c0bab077c81f6ac78b7c0511fa48fc49fd3f61e9b442f22d816a
zc58bd6355dda97dfeeca45a95c14d3cd5f6407e5baaa59c37a38805efbfa50ca2f6245a34c7292
z78cb1c1590ee2a28c25f754c36940ddc6f7eb0efe899e13d48ce077682c0c25f63ee6ad75e9771
z37de6210b036132229e35216192256e26e473713ade1d1281174ca239c057cb753e99bd1bf61ec
z663a0ff80916b63f101371eaf0c6c2b3e353ace7961989400e818cd99e5a6a3a2af8ea1ec103ac
za6e07c2498d45c163ff511819f50e918d4eb7af1b902104de522c4e916a8d37fe918e50ea7be0f
ze16d0e2b3badd442da2a15fac1d9bcc964611ee7c3207acd2fe52627ccb3dcc9ff685be9cdaa58
z6b763750b22562f0f688891ccade41aa20e83ff995cb58488da79a8a30546f24e926b8188455d2
zb77ae49f2103707e6156230f460315baf74ef524006e5068b1c962aa6a521fa868b60bbb4d14fe
z78ec7b23724eaf224c5fd084c7a532eef84fddee3ce2ca6ac0c77ad02b02069ec2fa1b3468b957
z5495fe99ffca550491ed05f2aa948088cc2f54bc13719b05d5656d185ad079afe55c6c0c53761f
zeda3e1dd94e51441857e87864d4cc87121d0668fc627be0d8cfe49c80f50b405634f1a89de848c
zd8eedf6d7344b85deee310a97532e3d788c5a265d60496a27e285df5bdb3b7bab1c55c36fff1cb
z428b50f6c2b3a665eb43b2f2c38cbbed24033dbc93cc4766a574785fd21b177cc115beafdd2a46
z8b289628efd9cfc2d27c4561bfd1b754a52cc18cc7d7a45f0db330ceb03221c8d3438a4c6ebe1e
z6a7c631c4fac4a0beb82c9f01d226f39238faefe0c863a123fc5274ea8ba7647d63713a35e4819
z08dfa400c6ab9db67517bea10ceb18fc8d13d9ff8c6ad2ef7192e313cade87b14cada36aaaba98
zd9c68359f733824d9752ce8812ba7d9ad68aaaa9dab4ddd15a1820cb297dce152c6af37a86b9cc
z64cf980ed8a931b66da139ca26581118e7328fff390cd91fa2dfe184ec494d01e4c23db7cdf391
z863587321c3eb4246a712e20b0d423e5e2b3cc35fd7a66d9ebbe184cba75841679cff0c4efdb41
z58c46afa364e5763b88d57865af7a53ec6d69321bf417e7d3e503f9c6c8cf0b498ba5da389edbf
z5b173f80c5d1ad7065bd8b4026f14a711910122c63b67e0d43e8a478f7f1211cb7c39534b57935
z4fd6f5432f676bc83874a01c0cab48c298a8e5e35f168353ddda824dbce63352ae448b151fd88f
z102c58f429f82ab82ddf4df67f8d37e3cb222db77d6370f3aef12ef059bc162f68ad0c479ed8f1
z715ac0f40756de8088cb059c9a26f057802c4c0844e1a472aee6a22dd236804e1e1e36ce148bfb
z651e6cbb01dd6b40e54a015f7d6f28424199f555c6797d2298ea7ea9b1d611e8e7a4bbaba09e44
z9bb8e74b11bc86ca0dd5eb44dc3a541d21115ee9f12c2ead7029c0cfca20cecee768a95fbed63c
zb644da4202675ae48dd21893aa7299bf335c3d88f4cb16abb8ce2067649d6a0a62f00077b847c9
z17314f25ab562dc1c4a237e38dcf384d78344335c6a220a2135c06eeccc041a08b9a554b770c6f
z6df9d693ecdfbecd48cde29cce4000b25362da9155346817105c6225f8ded77860e966d98c5d6b
za79650fd658788ed6e1e182a66c315a28acae148c86541ab67c1c80b65db852bc5505a8325516e
zbaa654d8ad65d074af08e36fd8151e90ddd33e181c67213614097bef680137b2da827c89a74eee
z821afe8ae388d7a0fc090e8af960d106d06156049c1913d4e7867d654b00ee51e7772e4d2265d2
z85a9688ab1045863d573d040361d5301f403400ae40fca426f29ffc1b0cc44f7403b9098f575ab
z3c155b466d167b7e461e9c1845d6c1533cefab75b29e65babfa117b323c8398b0ffc234c7a49e8
z073199fdc82b5fc264a5f7382ce285511fd244263e8dbfc66db1f358f0d83e360d98459f1bf872
zb3343d9cd6c0c0e9d39b0210d65ed1590615c69694f8c59f2683f7b3051cf44ae68127a8592d95
z59d9a44e963b5c112b3e9f14f066255c7401205a1e719ca12c71b00a4614312666d29489ee3cd6
z6cb1c509d33fd092a61004f629a6d4f8b13ba48daae0ce4086f88365cdf33ce31028189aaea014
z62c8cd09e78e6c42915e34b54e85fdde7ce42e7acff0df7cae15a1f87e47f92203e601b5b90dac
z7afe802df90a15c17eb65f9afcabfe4d95f7eb667c023cef5513c24509867fa74af1a8e6cf8fb2
z1bd1adb1e994731616c12613d2b80f478e592aa574a097312765af24f7865f96ae8a3cdc0a692b
ze3d0984c5d47d689a886c00770664856058375dc7968c23fbbfb54c7953e015ea5a1c5a8c53dcf
zb677a7dbc4df46a49202592058c148ef7fb3da2f3b71b961ad9bd1edb0b3283e9a7f246e2af78b
zf3f138fe6bd4c5709bffd0faf2b62f51f4cde9526f2becdaef90fe499232244a8716bf16daaf5a
z63e156256aabc343d9bb3d34e3cd87808928b804aa455b93833f946eab22ab9bbd98146060e921
z4f3d1a84e03b0aac578f37564184ab41442de9907c1a1dad2487583b3b5fd980af892a6f6e449a
zf75ea4e3f79d3bdc0230ee33df249ded5fb642181711d723626582842c24a67ceb5fbb89c83e67
z1ce11b1804ced9c43611233323f4af4249ac44ad716fe8f0bf1c71fa3a30b95a742c4cfd2be183
z6bba476c0b03f7e98950a8a00bdbb27b27c6654e3ea71e09c265efced863e49cf8cd4a29ca404d
z8618b2c639dd177803f38c77823e1c46b3a292cbbb2894c31039fa2648d2799739ae98716a7348
zba57f84cceea6e56b7f0a3cb0ad726d94296f507743346c99463c4fffb6bae3a5cb9067725e070
z301b72c09feb2cb341e39b4e6ce814366b3c30fb2d5dd1b39909b7153119fd93966b032d02c480
z938e7e394e2eb2c13bd2725bef48deacf1c24cb610f606e54586a896fa77d56e232b68af39ba36
zb3ea83244c77588b04365eac360a1d637995f15fb8104226730925fc8048a38ccf16b2b3dd6efd
ze3b88f6e70e3019cdbe7eee7ad1a865d5b3c1cf08d9db1f4749ca3262939001a5eca02a579decc
z079c905417a41bdc5d2f0e028164d53474f4f6999812bd7619597d8cd6d2bdc8a9a7b4fec9078a
zb666cbbfd67efcaaa118c33268135c151936e984300ee26440a7a7af180b17f0a10eed62344d01
z11a1fbfae803735392280255298fe6f03b8ebe2a98fd4069ee7c1289c7321f066993493b5d8407
zebb1435d813d5a8a93782ae40267010accc5773e60a68e1779f8ca84c73abab825a028b0af9307
zd6693984e8cdd8e557303b155da4b575509893922c42368225a1f7585e8f28306aaea3055b9771
z4d3a7bf7b9789f4e17316865c296c1ccbe0b09687a9fb9ce1ae814a2e8f91cc35017133ca8e058
z4b306220b5610935f43b1841f45dfcf04a923d7fa47e5ec079728222d744b31fee26553b4228d7
z1777e9be911baecb4d8631aeaa12de4878fc5a0a74c4743743f801d5218776bdeab86934fdb78e
z8a9f458a6302ea4a8bb607b47b480e9e438c43b04d6a62ad1b54df72ca8dfda6ba6c96aaea40c3
z5d2e188a8eda4842d9b8ca703b4a7a76c78b361f93b10a90028b1b91f998f923744166bdcc5d81
z3fbbeb58354e0d1cf6f34892de490e95ea693bb0dc999af29d83974c4ef255d936f0b1d382c759
z877839532fd9c12a95a069e35d8dadec7a387747b295836bfcf8f791e59996bfa713c16d30ef56
ze8ce6b71848dc3cc13c11291f42073c734be35d9dcd690c4cf2868773b2138c292ab8d2e274f2c
z36c34a925f2cb83e52659d1a4bddd3469e1f490717ab5fdd0b60f3e9c95468320db4a70ca25f9b
zb9d7ccdc9ed9d1c6f7cc8e0fa4
`end_protected_0in
`else
`ifdef MODEL_TECH
`include "qvl_channel_data_integrity_assertions.mti.svp"
`endif // MODEL_TECH
`endif // encrypted_0in
