`ifdef encrypted_0in
`protected_0in
ze74c34e226135848fe16db9ffd31815111b6d7fb642c521a3f628cf6da949865580b22efd062a7
ze90adae0e65e66a2c36a587d0a790699161455169ed55a01f2084f11770a774ec4c588039b380f
z6de9c5084882a40b79a175f5c2114b2b6d78b070cb806e1c0aa9258297f4687ab308bc470f0040
zb0b1de382961eeeaf2e279e1462520fc31c119af8f2b214846f56c2b3cd2eadbe4099496abff18
z15cec83ec4a77b868344aa20ba7360908f5c0de2a79abf8b3534b883bb12180f68b5d4beb444cf
z3fba8f13afb0abfe8fcc4294810f75afe452434d2d0f1166236c82f76edf1e12979f04bc35693e
z32ae028996dd85737a8f5adc1ebb94f39c940246e887647b64782cd7ab429b0544c173176cede7
z01dfb26b1f73408344a52b7e1f117f12bb9c8077b34876c2e6fdc085981637012dc9754765e1a9
zc512ce062e0b8fb16a214591f5c81e1353b900a611fe1f4886b57940b41b7f2ce99a7b84b04b90
z916f717e73bd10589c81e207ed77ec660a8cbed5b487fa50acde1b055c8870bd8676023f21ddcf
z9c98cc47cfa2d654ff1365d1f45035a045a66c5dfa8279050262529d2cac9e64fd27d9c7de62a7
z731bc808811ded9016570962244887f98fe5440167bd0088f2f049df882af501358497c3b28776
zcdc5426c7f52a851c35106bb93e16fff984784050fc808fad15da330f6f0607eda2d0e0e4b1215
z2ac5b11453f6b6c5c6b428261a64553d70b4ab9f1bf3f153bd631387c118a296ca10cbf0349426
zcf2ea5eb241fa84c8ecbbf7180f10eb9ddd4966d421e6ca571b198ed195474578ea51160ffbd6b
z0f73216703aef2bba31d04f6d0877540c760cd2535de4136d5bd4771107747c34c07fab3aaf6bd
z67c5eab3938266c996e67839bfd448cabe88dac2c17438997a3ee0a0543dc656070eb3dfe7c0a1
z57e24e01799b1ae1652a0133882b63649084f8bfaa3118d244afc7add4754b673391576b226b50
z3f1183996cb6c7aa50dcae3ab472cf58578ab5f1cfe4908256c378b43534b06ce7c49d652fe037
z4b9dcb973e82556d0e8e17a3d827e91bdf67c5a3474825f153107407c6eff8009f2a7a43fabfbb
z9aaa142e720d087cab66d83008cc56f7491e9a22479095587dcbb5f35a41a9091c9e504aebaf0e
zfc91f5fa18bb5392a828fc464263edce631f47a1220e1d3f7d4f53df54a96d88ab7c4410d4d1ae
zbec8f8ed8705cda750c8df48029be54f05a4cae60cf5494c5d92dbcf73961f4c0dd65d062cd4ad
zda89ffd02c8af7f34ee909e4721a1973eb623509212c549ecbe2ccc2952602ac3dee6784e63fb2
z533eda1e6ba2a4b8d70a0cae128737ab2c7171ce5211683003e91b9b395d7a9d9e9f098f6d88dc
z49110d66ef5c63f57a60b437654ca0938ec3e1fada5ea48c3684f1c137903046a4990ffb9af4fa
z446bb644cc2efdce2bede3891dcc34dcb5b72c753100b4686c6e680a7a8f191fb6a82719fb60db
zd49bb1cf9ee5353aa125c778aab5fc573fcfd8d0c9cfb63ea136af23c6487f318e208e4f818dc1
za57fcf68713c6a169e7346d64a865157dd68c2bcd94b58c55130d4d1ecdce187b18db1dfc8b96b
z784e3f05f3a341dab3bc17fdb0bcf85013d23c1beef3bc345e2d440d0050d35ddac2ed9c3b8c4b
zc0d9f70d1a26d2e1e9e1d1b7bee17c8146314e69b623a8e74e637ea9b411bf51bfb1bfe36ff56d
z5e37d717b40ab290c0681e3fd8feb846d3606e9f1e98c64f5336ddbaa0a2dd3a6a148a6cf39704
zcbcf9491a7ecb5890a72ca3bcb8a89d3d8896e3ecdefb47427c2b249b2e12504cb4af8bca4d451
z7b4e77f9ee5f115da9fad24cd22bf44e2df618c0444d3233723736a3d5814c2e3370a8f94a75c8
z686b8aa5d3dd58f44107d1f2d6842cb49b7d43fb2e7c46f110d017c4044b2fe634ca92dd50f0e9
z71c9582c60fe085bbb0f61a6770314b47c8bfa0002a24b46c2bc0a3a4c4661344eb93bdf363547
z9e7f307daabe3196ba931344d3880309a02048f6f83329c3b6427142201eb49476abca348e44b9
z68591de0a3f91eeaed99c28ed6a2bac1e989a159207db57a60c063b8771f182cc05fdd3f1fbb1b
zcdb662d647c1334c2cc954028eaec1494779b9a9dcb02f2f2d6aa3bdcf16f3c968bb741a745f0e
z69c96389a9a7f868fb5521b2dc9898142295fc4eeca271d66e41dc27f38273cf31265ed5778263
zf690ae07ce6010a28f8fe1c6c14d580faad1d0b6f758a63cd6240fd4ce3e02b705143a53d5272e
z4f3adb35164b12dadbbcec7986a3007825abb4c3a3469b0b9f7b0f89c1d9307e443d5c1963a6c7
z9f3318825c20ec3170ff8359e2e50b0c38b8d6e4ffc8b19240e82f9786f8c5954f4c727bc952e8
z548e78ded095bcfc7e479c24106a6f37c91e37ca8975b603472d4bd54a506d6a570547326959d8
za1f94d362983170593f1f69bee5dba30f3663332d8b4fbb20a14c9059fca2a6da0df46980ba9b9
zaa53b7f3337d58fbcc3a568525ecb14d7a2fe89e25e7dd893fdad1b2667dc1f0109fc092038aa8
z141ef33f0482d9b1885ca60f60b389abae25bf265877a22a3a48e598d4b8a46fd3111e22f87549
ze21499e48a55856193b6c41c5dee8bc6cc20c6781b120060f6b8abe267f53ec226d2ee9ffeae7d
z3aa6a3a6e8d059806efa33eb3339367becf473000320ad8b56c9f81aa94d4e5c05ac39da54739a
z00e74bb98a3a89575417b170fa441d2e2faa6546f30c573a8fea16c3bf6fda675396c5db7c115b
za3f4d583424910ae7962045799a050461c306367d3e081c84fe781200d92566f58f54b4c058a7d
z3cdbbae9739ffb0a3e86646f0fb6689669ce2004a1ad838ec66200492a1ba2e1696fce00a123e3
z8b50e65c690ef194d7aebe8e70cc2cdfb22c167f5ed659d681bdd3d1a156e37a9942414ba19d7f
zd70284e73d50d841d58b050702421da36f11ceda16e24c67c7f76df4e01b73b0c6cbf522abe88d
z0ea74247ad253f7884c59b9f84d88ecdefe1b2573d071c051db85a4d487903b3726bd4eaa97e5b
z1612513642acb5a778b47c9f304c2b31c5ec8479ba1f35c07088b9080d4f50e67940b4c329190b
z4e10e529008544419507d9a2c98df7b0aab97ca1e77dc7da4d1feb617ab4872fc97750e116b701
zfe7cec487134a3c4cd1be4ace6a113c28eeed34d639acf9c6922bc79b98b4b22353eaa17ae96c3
z207e09044d91dee6de0ce1f96c8bae0f02881d68c2090b2ecf22d923a64fd7453c6664b8ca77cd
z5fbf41179852483fff4d961247d09c3c568a8a66242737aec3b94f5d714f004d058b5a432fee7b
z2e68f15939225aa68c2a8b77011074d3585cc76f343deeef2bbf79cb2f658ac4414d0c40a39c28
z5af0d1fe67b21a8ed88923e767e5d5422948fd1f6aee9e47bdc535b1872deb7f3c613a2682957b
za170ad7ee412b32764bf7ca44c7b624e63db2279419416e511983fa20034d1e5bf79979a5a81bb
z6a40213777fc96f2cb61e9acab132182678f208e2c96f8fb5a25ae592f28c08400ec64e43b6001
z1f0b5e7e5294ea04b42b63e4ceec020d73fb49858584819270baf0fb8db11ca4d873cf628a5137
z75f2e840cf30afe535fed95488f15cf67f93c271b1bc4343fe20f152bef318845fb490d5246311
zc578c4f21993fd5c189c691dfc4b10bac12c85d1d6da13b93402af1dacd16c317b3251205c56c3
z0c0b651566677f379fe67873d7dd9f074650ef128b2e763ea75ee9d5ca6cf8bb345cee7bfe956b
zf0d318315f0787f9a7dad89dcaccec3e2d33eaf30560d8ae08c6db2a31265bb277da0aa71b9297
zb9fde97f88123ecb4b47070a7841088c2ce3fb88f48c807fe5667a50e13207a0c43fbd6b031807
z00b6c16261e70873d2b3fb38931a76bd9f81a2a73ec0c57fb8a65efa02a599cde724bfad9aa664
z03cfd35ed5ac00c6b1f406521900b9b041c3e54b38c422ed53e439458d9c29dbeb2a3cffebc66c
z3a6d505e18d0b6e69f3417f52abe46c655264aa1fadab66e67f1a87d676da91b44acbd73995f5e
zfc0095468f0648dc8689c6f6cf227da1d9aefe654aae8d02eb4d7fc2e94c0c694b0d90801db26d
z5a480038f6831ad8ccff779b31e19d9fdf56ec0bde0f3525ef2bb166b604edc8a7e80c9c1cf744
zf026e85f75551360f04c152b012f87ab557b68bb9eb70afde0aed3b97ce27e395d4378e4d0d215
z7079296e28f7ae1e0a8222deb9caf9fe4cc32db8da99ff693ed7b3ee488f58ef69d6a9ef8f34a2
zf2ef6b0e3d8ff3b54118c622f8b4c34c53705da030e35b34e48d132fe6b93ee20fc68828408893
z69d117a2fe2d348db34cd0344eee95981e74f4629fa150bf42c6286662b0dbcf4f5ec0b09aa5d4
z4dc29c7820e325e754e5cd6b41b61c75ac4da69b82aa15a301a7262ff85f892fb77a8ee6398c10
zc15111defdadc9e84c43497b87408814d3cdae1300873680c42c9c15dcae3a4e2d748cddb7ded6
z35af72199b4847c2a2d27cded8b06d6c26631fd6e5971ce4a84f40cfa6ef0b44210612677d1420
zaaa3b60787d4e8d84edb736f473d95f03473f50083340f1fe85262945b29cc090692d76145c73b
zd8767fb36ab51a46187ee97ea9ad4c6921ad1f7f1ebbc2638d48254663066be678aa0f390e59fb
z80f44d22cc95c417f23dc7029bac2ffbd621fd7616109aa47f9aa5ade3106ecc4a420daa259bbe
ze8018b6c4f00021d312fc814c87693339d26418ad49bf6cd485a82eeec8ab1d17d98ee9a70f67d
za55ce4a7b2803781bf3460536ba77ea87f75f3322d9004a0b1d581f12b47dad0e1d57d93232414
z38b78c5da109dd8240890e5f955683a977cfc79f826fd5ff3a210fb89e7756fe43960b67c14871
za4c7ac9d7e4e30cc2b792e17fdebb5a05f6da3113321fc5a223d9f489f971a3fe2e9fcb468ef10
z9cc5e4104e2e1f1717dde03c29ba4f8b96707b59ce77d45306ed4aa47bc4cff7931151c5947122
z4589caa52a48df6c18dfc97fc0eb5a8c101f0fdb176a9c9abca3da65de424d62351909fa780e4f
zde7c18d270724fbf24620b307d4797e59140380e9fb6885afd7de35355dba41efeb6dc0e99cf00
zc16f6d6951e98113de82d8f93a759946ae10748f3ce569505d0a2ca0ceda3f9139149e56a3799a
z73883185aaaaeb23eb761d4938c08e4c97896f689b390358bbbbdfbc349975fc884b954e74ebe6
zd0982d94a92c9e83690ce81eba12e2a9d3c77545ee835365293236fd2949f3cf975f132c97904b
z1197e312e6331ab709c28baa7bb2b9a8ba637513e66e5431212fa23a64615e20519b4a466be435
z3c95647ae07151079424dc0910e4284b8a2313302fb0f000bf24cccdc7ffda7ade54313a1f7242
zc986aa0aa3db3995b5e096b4bf0bc2e53d6d21a94a76b9c7b38459423cd91ae2279b8518c34e60
zce9467649ca3cf652a2ceef9f2bae24549f14e58594cac9b5f6483e63b4f384a116158e65e0be2
zb3329af7a04c9143c6c89cf88dcf71fd5edabfa612304304cc13de7a250470557b0fa1c7e016a0
z920b2c3acbd75e466d6360db73979d704b48e9a2ba1fcd2b721982abe767990dea0a5c55009932
z2884af288dd6539e57e5b7af0e1085de571e4987bdb864312a96b5335a04d4af357c08288b80a0
zcef1b73d6ba3f61cd6060b9a9670b6972db9978e4123dbfcd97853def8196d89f588e0c1a365d8
z0491cc3b3540576ccfe85eab07db09075f7fd2ed1f43db0a718a8b2e54363b402ef0ae8cc2b71c
z1d10116ca338bd5576a2c25c2f21f3561e7d926e9d1d8f9642dc7bedaf04cdfde88d7e0b54c125
za1f13340ab6a3ef7e593cf580218437a1792def2f1abfa8f440eab11268c51337260149918887b
z91d55da3c89e70067e30c2a88979e641c3c45bc21685692fe6413b7b7b8512fa607d069707023c
za0c42ec4b3410d62173fa140580019a67f058a201d03e021e7d7e74c169ebdaed2e44642954d9a
z432e228796914bfac1d1479094495f5a615f6a3f3dffeddeec3fb9d3146567045b7e68fbf00a99
z47b39c09aca8b65c4fb3f8f54e65d2e2c832e4cb12ffeb7700165c856641608935fe28bec7b5d2
z43b114c7d2c5b87647f2adf6172a73243eb5d9167e82373ce221933e21c8711644189026b44e2c
z82f5bc79c8cbe4d66ec746f55ed727090d37b21b93f619b6bc0babdb550267d33375ed45a0d155
z31f825f59f8355e5c6af1f47b9815e0462bf996aeeffcd813b7656949605e01e4692be1a296609
z8df80265e846427550c5ed0a4791b152eb8c1e0175f311a545d2b80feed17cfab0f61fe5991b5c
z7d1a2528d020744418f70a541f0c2c918e97a411a44083db6983682ce7374db66771d8a1689c55
z96dac730c639f39bc51b9d964c30284669a01b835b7390789c593305f4209c28185ff8c57f9dd2
z656660f957627bdec3a7761a1a8b7ca9e4b926d6a004ac687de0640527d3686e869c5deeabfb83
z0c7bdb854ead75d0ba86820c89bbb93251d70c73959d446a810356b0061a16c1a5baa3de16d8a0
zdd22360adf1bac2a84a73603af99c4894e0482c3402cc1d96583dc6f4e09c188c6b2b8e3592212
za2dfa4580882b938c3945c9db3057e8f83b657fbfa3359bb88e4bada299d4a4ec78a6f0b11eb1b
zb5cec3f5a9dbce36b4597879216bc80d80e2589e933921cfe1db1a90736a747cd8c706983b2ec8
zd8fe2ac2ad8f1abf7db3987e05f6668f95d0172d62c01fab255e8bf410df4191fa97d9f0e316e2
z858f1ff3a988d40d7c55d8a0cb12cfb4c85135f6ad40b170c8c307849d9bd171b3ecf861ca0a3c
z1baf3fa90fedff8446ee02e3a09c662d8700272a0e0db50bcdaba84ede665f068a3d19a0b599b0
z0c425adf2a4c93b3d688a3b41af4fafebdc01b1bd7c9cbabda2dda001d372911160bf477a20f96
za02c5a2e9e2584a98710e39bd8632396e953a35095637cf7b0f0faccdb6544dac1b551b3e758e4
z8f1bd826ac35952cdfce675715a5f0596f9e2e646ffd7c9fa363ff52fb800b389d2bcd98487cf8
za72e58850ad1ec45f272697159c6e958243cec685ffef7ffef54ae1b7bfe11b364411eb8efcb9f
zf37661b317941c165f4d24c2342b1df6c68c59c12addab66145112d98c20c4d9979a22cfc50af9
zfbea3c0529d1d54b336ddb656b40f97a9ec0225742c65caceea00daabb838186047fa53f54e55f
z6abc33d7bc4e48ac4efc9d977e9259557a260dd52db5ed252bc74a97b4d30a6b51db50206b6a7b
z59c6341c43cfd1e85f04c0647542819abc55b9bdd899b6b65ce85d6c5637fc888d8fdc1e3e53b6
ze6de11495195b457766a4a92f2b0d0e1fafd863a097b4bd5ef1aa82eeaa5ddb463dbff086ceb7e
z608937188f4dcce647ac68c3e35329893ff56f2bf5bda0b1be860cb15b822ce1d619138a0c7729
zf75e5b15240af6f7997e8db9d60d72941b1c89c6e2e3c337e2cefb5a6ca0ff9a3fdb9e447d4d6f
zab13808e8165dda8d6f0624d9c59cb85fb42f5cb16ad2626f5f341a9d737fe0751a6b6c2a7b4dd
zffa8aa0a70d4a97d324780e51f7b0e9edf04487c3ebb460c7eeaa453362ef2b5034b809706d06c
z0cf3c3a98b77b96d054255d40af1a4000f8316712a5804705dd67a8b3f3352085d0abac1f5ce39
z7b2aafa90b4db1a9bdd65bb012c8eea08bfbebcec9665e185b082d644cce8ed400992410ffcfa6
z8598b51f0140b7a87b9a281dfd41fdb0d7945abb6d9e87dfc23065d3e6bb51e4eb1bdad443b6f7
z94abd69a9ce92b49f7ea7140e651fde24f586db2a4e69f112b853e5aa7ed6cc40d1cde41100f2f
zef427b7646fbbd69e2ce9a02d2fcfe23ddb622a91428f222451f18506d52b78524f1479758b006
z16da26c246ecb099a6c0baacfad175c4ce3aa7beb484abc6f0c394c95246f0300ab9f9ed27fbf1
z259fc4f778080bb2486d9e61074fe64d348e7435ba7a1249904f7d6b2b98bc52e1a06ac2e98a4e
zbfe664ff618074d22ac3e158e8da46c843548a8780ec693180f6c351c6c2bebe2abe4279ff7739
ze48ddb09b6b5eea29c18150379d2d59d6d253434361624b273c0c98be6f5d6659d73d36796c06a
z7004c39179bb9c1659cc0d12536da4b7f37b230b04a03501b02639857b4afa5726924dd97c6599
z25c1c73fd836ba86e06a6ec5c92c9c543ffa4c0005993f9d97621fdec18b04697c3bf787cc4437
zea5a7c7f008e25402bea9ca580fda70683cb20891039bc8a6a96cf40117d113d924c292112f915
ze1719e366178bb63d747b862379af9a052aa51f9e0e9028cdab49b9897218ad602b901f020a3a6
z2ad631921b635e6e5bb963a71325d425dafcb7d45fda69e23a06959e7a318ecf967f59fe078292
zb6a7235422895840045ecaad41ff4021c8982fd9ec8f5ecfa9d05848b7409938257b1fc28e8c09
z82850742d232e6f5c577d8a6c5a25341eb46c271ff98b1db1b972c7988432eaeebd34f2430505c
z20bf51866e22bca91b8130c1603f4903b86d8b82d810a9c7b9d4fe7b5e5eba221e250851a3d9d1
z16f755f40ada3fd5b90fd5c88363737912c996a02ec2b17e50462aec3d2894e0290dfc69aaceb5
z843a6b0e1f89da57f59a5a555066088672e891e169af66ad51138c3823fd6fdadb9d5deea07302
z33af26136a74fb718b40a280b81eb5d0aa82781d72b0c4e474e1cee4ade6539bb7f28c0c1d8b2d
zc721f3ec2200e80a1f4655fe0613f76f9c36d840fb650ad8193a01665bbf0f011caff3187e61ee
z8c4f720fe136c7d9c9e36fa1ae26ff1ac263754175e5e12f7e584adeaa4b786884593623677749
z61c9981a264f1c9113d0379b3da3e51301ed1fff5104f99ebe907fe19f0c35ea385a0a4484c895
z8427b1debc6994f25f02f6e014d1fb3e88b31fec028d576410168032cadbd0b57590284e969db6
z5752a2adc55a69b926690e4e66bc24bb9bb1c6af5e79d5e1f19aa4b942cc11098ec127f332972d
zf23dd699cc7dec7be7e3437fd660861b37717a377adeb48dbf94e53e25862e41438664eeefab1c
z511e05e5582a9aa5e9efcd3025d7b1cc5c3f671b9254d0bd0bd3a8320c97cbd3dab6ca0512a4e3
zb059743d984ef9da59fb007f4b239118eafa65ff32a2a5f8bdab1dd877ec95a6581ac2272f9373
zf0634384fb01ef3e7f7b1edcebd2046d80c35441b350494b8696a200a04150281222f155c9f557
zed322890d497286df85b690b98dd58e449119a4d06627cd074a99bcc51eebbc2c71eaf33c29435
z07fb799f8116277db4b6db7b8163251d1fe5d616adc57db21e0952cfe304f699cd848f631653c9
z244d0349fbf483160f764da249714229d5b9ecdb84bafa433da451eb7dc8484af95ce8e3cdda6d
zf89768de1af46f8aa4c2d3f3cf6f99965efa233e8b8de0a85bc47e8e477579763a97aa9981fe9f
zb4ae1dcb51487dcfe2ff862b007cfed291e4f339e965d221f8ef3e8cff033e2d002e105541e49b
zae06811a963aec929d17f8e5413123ad03089fb91dfebe86bff236fef9272f5a7f89bbd79381f9
z055c112c1037b50072f05b513f9dafaa45e3b8de2347030112271f7a64daab80e0dfff6b3dda6d
zc8e99245a4efd74d3ba5351d6c125e5f5e292c05a49ffa3b8f681e98749918cecc97b442dca1b5
zecef521ffd62f2713e1da869d403d3a34f5c8b3c8073e8a459f72a970729c2997785a0ed332fcb
z6faf8eb0a5b591e81e186a962299bba3890d22cb773d4a1918eef23a9d5842b4ccdf2ed96846b9
z07b17011a807bbc65015b358079d3fee2f95547d5785cee1ce33c8ab5633ee2d71612769713048
z32ae62e9052c3eca410293f2ea73081072d318fd5281dceb02cdda8d34616d6f9a2084f28e03b1
z70e988fc6a1d95b931cdde4116ab64c2ebce36e6873323301b89b757b6a8b038474452ffe354ae
zc8a225d91a7f6127a33118219150348e432343314162d7550ceb113886d4bdac769f097a7d3c95
z7d9ac8f784a65537d453ab85b86988b0b2f6715814f3071a92b1b937233a21a0129ec2bb48d70a
zfc8ad0e5a4722b0dcc6870b314442304b290cbfc6f5166cd4e1e4d464b0ac7892a6a551184c498
z1a0f5e80ded367b326f57639e3b699c8138fa8cc16b427ffd331635c81e9a121dd3775a2a66859
z518e40c26d7cb4a7060ae56671c6cd780f94eef3bad059a11da8c70acf7a138f7af61352a179c3
zfefe29cd3febbc24defb71a78bfee054b673d0e80e4660b57867e01e4960111c0bb0f16a0b340a
zcfa101f54e9a3e310cd28df30390bcfe051c42f9ee450fce2689373e38ff0afcff83153b0b84eb
z8a8e5a4ab0c5a436eb66896907e1b65928fa08f708fffacd6bd8af7de1a748a307ccbaa3d8667f
ze929e95631ea3d9b2f872a0f517b2887dc330211c6de5edff2bdf45ab63c096ab9761bc53784aa
ze55a355313858182eae176324b2f974833dd1ee431c64d1e4d670eed1ad780b30d409858599f89
z67ec9cf14762263c64c47d56b570b1ad2a42f85cf001a2ea4afa0e433d69de070dca85df6d64ac
z559ee21c5a412186fc9b093e33f202d63e1d395c258eddc0eb8fc38b432d4e41472c516166a3dd
z0e33c0f174db01dbd8af4e14a0f16036947a7897e7ea2d975ef0d64a91cf457892836fda593717
zf453fda0257e2f3d60852243ab24469a75f1ada362c089335b33eaeff2953e2959de19b118e176
z25cc0f0f0770549d88f25e657eac75596fcb2f01eb721d4bbd6e3e3ddbaa0814a3367d00f51d89
z89c6509303fbca0f2bfce70e6aa73368e9b47e8de6cde1788274da70e635be303c6fed0092c614
z906c13a06a5298a82c2417734e3731347459aa5b15fafca8fde16966df634b9bff6343045ac32e
za127dbdf19f2e9583c15e7566f41a63d3cecb83f801bc084340fe49ac96675e0ccf4b49c9c1b10
zf78af2529410c3649e512c377fc6596b2c42fe5cb265863421b73af14e92556f02c2621a42ee10
z98bd57e77b2bd601a670f8b39f49587c7da5b95347ad27920be4588a967861cfe527c43547c645
z194f797fb2f84068a3517afa6e1a88d8e2d00babc5594a249a09f765384fa8be751dbd240c9449
zf6b76cc23506dc4e9dedfea7c7cb05658e30b59fe59b41c7673c4959d6d8931a06273dfebc69b0
zbd0e66f8a9300cd46ae877e3918237036fecf97a1f2f78f484632872da54c39005763123abc52b
z3eeeb2b4537b15c92731a21204a81b15791601de650670585f1bc069b0014bf9ef06831b749d19
z1bd24e5ae497e4ff3edb6af32f27920072b93927ac6f823defe7e2ad884f0fdd81beaaddd0afae
zba974c69dacc0eb81944005c90190403ba0f456b9737d3bfbdc49a02fdd5c60e658cae730d9d5b
zc3b8ece03870a60d3116097b36911cec54b9173a332fc0d039ac4b70519097ef44b7d2f0d7fcf4
z39311f73ec69ba229e438d8506a7642423e4c2ee803414138074a4c0b8649cd3c80cbf2b818271
z1e0c2d5026dc9b9887031d2c4fa60ba4bc5c839101b9fa67cadfecd14864fc1f3b84d23789aa6e
z00abcd5a719ba5276902952c5dd578254f495bfcc2faae05c7073cd89e48b46504ddf5ab794d4d
z6018226f8c1b7d12fc5fcbb21125bd037cb04051aace931bf666b03a2e1f431f3b4d843c353934
zade6fc48f34edbc552776a5ce10f028c3415e36851f084c325fe631b32ad90e43a7f3fa14aeb19
zd29d88bb547272b8fa70a6ffe684dd7d9dbf6589179c6de1c07f64298e6c6dcf01e5fede782eb3
z01e2f1cb8800457ac3a386f73ca3422c17f9da99c0fd46a3c1ee8f83cc374c1cccf07c0b2ef2d4
zc472509b40ebef4b544c3228bfbb9aea1629a1e64c8f4b122a4dd3a9bb4524bd955722dcaa6243
zdfdb9a75f18c20bf81b4733d687002ceac164d5290a28f99c56eaaa53192bc3eb2e8e02ff8083b
z14c77284a6b155ae41dbe3605780632898b008365ad152354c3ed3a15001f2a9e4507fd299fd2d
z81c34dbf82a55a4b24bdb6a58465b3842d0499fbb7f0af8ade100220996b7762bc7bafce9a42cb
zeb515f009bf4828ae3581383618b0e0e3709eff0869903388ce8ccba0f9325cf6c932a2ac24ab7
z30d43f9a35ef64ac5b5c79285dd2855e05e7b8207b789f47bdcf29f982674d2e2de998fb08e177
z3caf7bdfbe84bb763da7c2b0325aa047b8c8256d37c558d33b2effb494964aadc57b61e126bd3e
z430e88f3ae2e991655d07f7ec00c9f89b706eaa57bc90326255e7bc6d3b9bb202cd6a5f86fab91
z50dcd32549ca44bb553033c0965942aa2eb1c151de6564ef878d3a9e870b7bec28476f4c518c30
zede58161d49b99691201baea2a59e4339fe12bc0400090e567372e2263e06904464be207807ea9
z2b1438d814057258e2e0c0ccad9c9d08e4d936f9fb505ff61c9b2875ad357b4315fc38df5c0bc1
z0e136c9d5a302bed6765304505ce2eaa20f4d31e17b873e42dbca13baee763a2a8b68a6f520c2d
zc1a7a11f7bc60828e06576f5505488283a4590955ea0b47b34280c4e45753d32e239f6b71e0835
z82143cc5272c1866f970ca39b8267f0ed6fc7d419972cd1fe9569d1bf193dc3f8d420d25a5fc73
zb28b993e4d2f590a9fd36ce5f6ba84decbb7c90bf313f1b1a51c472babea4610461e2fb1d91a3d
z96909fc4d64d2042b82f418d2cb823826b86aec6e9805dd3633587cb75507f2c334ecc15473c1d
zf9ee7a331f0422099b1f96858de7c0816429695b97039f8adf6d6c685a4b9c3e596b43a9dfe77e
z26c89949d070ca6177862c8901e8af9113009ab703b6e1944a7c9d70d701c56035aac4b130032b
zbf41946427f5c7baa5444117e8cc5291ac18b0dbeae2b04bc970a2961ffc2992a40842ec904990
zba7495af413691e1e9f4efe4a0424b8923eec846555aa56372f294c07f147585afd2b378b01656
z4d6fd89369d8f1eddf1ca592d6771232d0bf72d4fbe3973b0496424a43dadd2abef98df5027359
z4a61e4503f53219866340a784256896eab9bd9b67950f1b31101947b2d04a9f4accfb774210fb9
zcb30fd6a454a20e813d77ef29345d16845363a02ccc7b17d31f46f13e2ba94e6c6352c27dd191a
z40bab4f2667adb4bfe8443706b90c3945fabfeb0d8dc750c9eaf76a4771a6cc6a595f0f1d84ce2
z97a3709ac37f247caaa4ebb0bf3cb314a01aeecedd3acfab785d7558eaed8ca961d6340470a918
zdf4fcaa531da6ac7bd0c6e19d3549e1edddeec644f9cbae1fad80939cefb2dc7ac9a3e9a95a62e
z14e8ad7aa7d1b911586cf297d077c6e4289d83a572b04dd78940b086ac982657beac2126842c57
zc59e5c79e568c044c1e7b9ba51676d646c62e802ea36a589c14c14d739e83890a829ff8069e012
z50143c0f335cb55686a34ede7ad0d59409b608ed2ef96ce83547b01a0293992fbcd50594c385d3
z1e3b579d2012d3c2f54613152ee088963c7938c562b0682004f1d5db6f6f799529f766ffe1f919
za6603ebbdd0f5517badef39e5d3e0591fad68f15a2421f89db6c4b05aed955e2165978d04323fa
zbf4213a545d156524346493c9637bc65c2017da882b43d5d13719655bf0bd5e8ef415f8f16fde3
z18666f5deab9011d284905d6a2fcbc6d5a135ec5fe732bf5d47b55405b6756c3fcedc2a6192e50
z1ec6efa807eec7cfd7f797bea53f6f46e7664970aa166e829cbc124612731016a4f653263a7fe0
z6500ecfdbb8155918b7c67ec02bb8af36d574ef0e851ad7cd19f83d88e541fac63e6679adddee4
z358c117e5c974476de99b8b94f71448e449d538576682c57a45dd7598df17b961154513e1a730a
z418c28d2195530b76ab9b552459da7598572c3915e71f682ac0959c23cda8935836316ac23affe
z10bdf44390d0569bcb5b8b565e9b5a8c1302fb44624b6a50a685e0fda4e062c3727442268d8299
zfc82c5613810ee8def3c83495abae64fe060fc727922d0963405b24ce85d14a45c8d882b6437b8
ze39980a28fe11035a08587b8a2d545abdd266c29333f3be1b173955a00903eb308896252173d02
z7245e6410583039deeb8a7ddf81c7bfce9db17bec5383853e4aa330ddc390f3540b98ceb839faa
z65e0e66540b66618e766ab1fb32e570898d2e8d3565d02167deb89f7c3a61caaa168ae44648e66
zf015356b4933b57a240c2f4d10df92ac0b9aa0fb6847a9cd872bef516624bf11db0fa0c178678a
z416305692c72fafc108cc9c3d9cbd49ece5515a6875141673407a16cdfe238a27470988de76509
z9c7b0656055e68c8dedb87b5eb05577e341e082401894e1286014779e8535e8babce6abbbf59b3
z4f7e7d72ad64e139cceba40841eebefa93836939525e0be383ae7018b9baca7f8437bfb6b2bed4
z81fd28a7b45dfd2b59aa93764e47636f04d813146041124fcf2bb0bcadba7a212f466e0a917c00
z8528f8a36d18686c9445fd421e69cfcba90b7b77b84dd8957b78bee84ad072a32feda744b366ab
zdce0085bdd1798a489dbcda0d99ddedaf197785cd0f93a02ed611c0efbab747c6d977e5642511f
za15ed55311dbdf247529fba3c8b115232b0f37a6f2f3cb85e19a43d03de4a627c1ce139565542e
z85a1a8687e574d242bd7d1f1275503ef19f8b96f6bf51b48616b6d5b8dccb33a5468fa5a60d7fe
z0d6331c55ddbe68b043c88da1310b5aa23a18f578e055985d6f46066a2b9b9ebd638a394182756
z96bf0c83cd5df626b64e164ba0ff708e011c0203cb7af5b4b796b87b33b41f1917c48bf25247f8
z8a3992138b9483d59a632013cbcb6e178c558723f567753c46002023631cde6abde4deac9072aa
z5ad313e52d10dfa2d4697f7c48d6a7e8e20ec6ef3f6dd52d623a15802d8cb47b844bf3bb70647f
zc011abf9df0d247d0bf7739f3b25d121176b8031a306e6f31f1c2aeef4f883c380551a78319615
zed3c3838cc716110e21115cbec788d524be54e03dfaa4ca38a2306976b1cfeb97bed7dfd42a483
z7bb533ef85b2e4dc32828c97caf245977e720ccbf7b8473bcf53dc70f6e250386fa2e3db7f7dba
zcd5532194a9a9c4c8205b41ac7b134dbf16ee7a0414e4ddfa815bdb73c5703830508509c6e8edd
z31c4a10366cd061077975a97e8e717bcead5413a80b67ed7ff617423d1e5fb7520b1ebb6ad5d57
zfa7bb76badd8c7103e7f7c265a855cd80b19730751cceaec8ff1397422ea289b45ccfd5b96c094
zbfad7893126bccdad203ba196f802c726ea3fe05ca2ca33b33980dfea74f172a244678474e1003
zc7801a87a26464f42c5966a5c5b169b219f3bf7e6ccf34a1199994ee2d4a43ee30f7ea0b3ed137
z6a77a43234cfb4817bfcc68d5e5e66577d5598427dd5a00b2084ac53f299fc564c0a8ad59e58da
zb86c7a13d21d2d21eadbb65eb66479bbbb0801dcd94e47a95069f077fe2f64b0aea431e740405c
z0744c3f2b78fdaec8599f9bddde321269810e4294691da3cf250f84b7cddd208d27d5a7f97dbf5
z4181264efde4ea52e5bee37517f0f053bb09906f96e41d505bd04a085be587a05e22a38c156490
zc39198f2fef827ebd1306d2ac462fb6311b4e06c1b0b4048dd92d5cebfcf808478d9c8d23f4e35
z79d283a354b4a11646fd37e91239fbdbd831de28e7cbe1e20a0996f52c01cd5a3c79775fa63a16
z8e3574be588fbfa90be5a9db9263474588e84920abfdefc7242f5aa0c0fb5c7d01e7564ef041d9
z052ed629fa984655718051bb53a280271d2654e48eebefbc3ecbf3b2575dfc194ab21083022719
z73152a0088f364cb40269829f840d00797fa6b6ac70d9aef44521f9bed0467406ece749a1f147a
z23915157bdf19d0baf1bfc3ab7db71d0bfb2b5e44dc3ea559582fb04ddbf863fff052993d4ca7e
ze7c2fd82ec9d2b679beca2dcc90a4f69d06e599ac2d0a0b21e4edc546e6eeb20d67c09a7f265fd
zc54e02bf959d6c53dcd5093980a46f264338f2c459adc5def6704d5eabfef4912102c8c6f032e6
z2bd75e2bbb2cdffb22983e7865ef33a667769c9d0d587f8b00e280b23829d0febf045874b24547
zf5f41d253c1876cea997647e57d5ecde490f845a3704911925a15c42691b1a41a8337470b3f619
z86ecf579cc80bb5d23aac7484414bf4a420ae245b59593c42ce8f89fb4e007fc70f6e119015a58
z43cc46fd571780473e527b7a18b267893a031a9ba009a771e9e7a1717b2be67e23dd352a31ae50
zddfab9e2a710ae0412275a44ed2a0efc4a3e91e2df9aca385a4df9298a24cc0b67da6a4d7ce0df
z27ec351b0d07995c60d10c4dbfde6715395d77450fedd16962f3a2b48db7680791ba5a84f1f325
z4c13df9ad4faaba5819c9fb149f4eebac35ecb6be6ad052e683bf644df84620bc2b7ded3b65f89
z91bec0227d28b455440d0090aa069e7e9b92622c6dbe355a47077bfb949b1aa5ae5523810d6050
z142ee5913624fc06bba0f849841064e86983de17220f025c4f214c79b6db519b3f3d033af8c3af
z65e8dfabb4634fccdae2b94fc1a6c591536caeda7a358b2b2e79c99c31e79578b472ac3233447d
z8fbf839408f0f202968a6eabea74547f918fad507b614f41059e4a4e3130eac9476cd1f2317851
z273d5e159bd234c4bc29a2df6119fc03a9859c775d6a02b8e817614b7ad1913ce2b5c7215dacc3
z9c03693d9666ed51d0a6d672b437cfd5d9f5456185a0024dcaf7c928d82f20ee16962c7bc21a54
z7bea003f73e4f1bfff158c55d44890173a9773971e65aa273e5772b01a1a7ed68b21cb9df83eff
zc001d7253744df9e1c2f7f3a01d151a05cb2b7f8d9ff52186bb3c88449dce645be67b0dfc210d5
z0a1f9cf04b31a1789f7eb7374584f7f3313f7116e612f7f85b799f8837af5039fdaa6cb6a7a7d3
z137e56221cea200b5f2ce8aeb715240e03bff8ee46851e48e3d746cf212a574135e1fefd931af4
z8164e73e744836695efe94b58de6b195f3134d32e0879ec9b48a2013c655e3496fdd0e21b6b54b
z58539bae773afdc02cdc97695f944f71ef5197d7fc89b02579ce381bee5d3f5005c5fbfe416f25
z245fbe4d858c3b4e876fd70fe30e3d6220bcaae57716657778b92b80ec6193dfc30abc5d439688
zb34d6e7e23f411d511cea99d0f44bdf86f83b0286d078b4d331d8121fb4b0038613c6eee722f53
zeb513b1f254b3d170d3467971a6edb67c7b7a10466e3bcdcc173d97d261120385b68406fc3a6fa
z48c5b82054b81e963799f81b8f2a51d67df858031c228a6413b818f9c38a5bc967b41898483acc
z62b00a4b40fab7b097a099ee1b0669487635cfe583d3f16a349d0a79dc1f90a44e6b142e1780ce
za23ecdc2195f1b7ff7f194c3a963403f50c0dd16fda889177f3348bd08ff4498f8308f9e3f44f7
z47cdd9d5af256d7381a304d41123bb14a264cd097701cb6e76e8c21e5259b30c5d21a24b8e9010
zf1e105001ca109e63f9654c21926fb346ed5220d1f276da6cb78037caeead604003780a02811ed
z3dcf49d864ecd493240323b14a1de519f6b65b2eb77a2168304980fa920f6c3622ac68aca0c2f1
z0694aa93fd252e6562361cabdc11b9efe49492f6d9c8014972e55cbcd2d9a70d94f7f302f898e8
zc82b71ebead2fd192fe01e931cf9a5ee1435eb3208d753c06886750fb2d288c236fd0c7f9069ba
z0d086568a34aeffb5f38d10e3cedbe9fe7fe9f87c5977c38951b1dadad5f0f1cd9112baa550687
zc83642167ccddcf53768f400f607d0185adf89dceb7eddfe060610084160e1f18409877b265f5e
zfc0848694e348ea2b553cdda61f888497b16cb26fff0035f3044c0fd38c6eb45042283e49d9f22
z0515351462b73200d37bb1b74a67318dafc089634c66d7dad325390cc6c160148bbe25cb244974
zb1444b800adc9696e7e090a5c63aee40b75977ee15c5113dc3a0a59e8749752c2fff31f61e3a10
zf65dd15d7a9844426abcd99b2b9a4f5134a40759098b2e229fc630595ebafd947ce52017a3c46a
zb18603ea8ace09949c4bf0d43c99dce23674a03463bf63c32384bacb2741ff2ad559204514abd5
ze72b50ebb37ffd465643dce38fd087d72c7f4a1e7f4e04d3358903b6c8185439d0d56ea7c6d6be
z9d36a7dd3dcf6c06199bb3db03a4bcb385ab72575ef7ffd048c0c2c7ab57dbeb8d74352eb096c6
ze450da640049a03e7457e5f065783512b3ce4bcc6e83623f17af6b4d5096eec01edf292a1dbe86
z58c7a226b37dd7861062790c04856e05d13fc46feb70467cd024bee404d752ba5ace1c5a92e340
z60c58cf6099b1c5e6d222a18ebc39979f107baa655ec21be527772485172e1a860b03588b9289a
z6c45941a93259bb4a0d13ef6d54db27e885b1022f15ec24ef25ae37261e3b9f77d6958b8cd6303
za96b452645991fbc20e381692287b520d704a741b48c9df65ed0cb1cb2f91871c94ea695acb406
zef1a19243f258071cdee83d9c3da18cfdaf25b77907089a96c76d7882cfb12d48f8851e6d12213
z9ff26faffd5e28403de095d22bf1a3069205df9a117db9371ccde35411889bdaa768f5758a4611
z0ab52e54a5229f5a15a2037e98d12453a703dae0704e27aa1d5f5d3b2caacd2e5bca4e43cd8fd0
z9e9a309d80677306ecbec0adc11ea52298b88096994d41eed9a092961c77b25c44bd573ea3b948
z2cc4526dd3560ef8e1084e210a3650248d7195ce63b55121d9c3d7c0740313fd9ecb93ffe6cafb
z75de39d2eedfe88f35090618ff8b9813f7eda56daf96d566ec991a1b9fd48e3cc9aa20cb18fb67
z72a0bcea626e5728b96fb723463f0c8eaec111ca5ed1edabda8bda9c32372615fddee781470345
z44707103f1fbc4216a3f24aa32c448c421f3c620e1c3dae641f73fb93ee3f0833e9a41b0b2da40
z09942525b1c69d8aa50cd02158c6454a19528ae71fdd187b7c17eafec532f7954156e033b61edf
zeaba1f95d9c55c1695161d2e5d65c9e0ba65ed7fabf06bdb9e66f744ad9874d67d46d878588dfa
z93717e0b5a063fc08181760dec361942d59c2aa62d1105c5d185c55924198b7d50e147c8b5c12f
zc5ba1f827fcbc759f8ca4fd2e9a7cddcd5b733cf4d924a1345bf8efd941db46d79376907c9dbcd
zd2b32f4ab814e076cdff43876e8122b0d272094ee034bd4b5e8de3bac7fe7ca039454dd8fd3fd9
z3bed2363d6e382cf2b635bdeb7a648394181b6234df9977ff0890af2c0c088f45247343aa8ac21
z85ce648b9bab53b82e4abfb937f5756f6daec9ff3ede5ee069a4b228c812e485c053827acbed87
zdaf295d5b7c1453255e8d08fb0d34195a928fe935ef23bac81fab2854e0d92f5e8ca762c069896
zd3276688bb749310a8eb3cd11f91f510cf04637c8853a53f9f0f0af9fe01d109aac21a6e39f4e9
z92b5eb0e3e41061217ee948613646809baa90e8cabcb181f28585f6e66b08e12706759a842abeb
zd3a19f6d23bfca10e67360869224db5a72ecff1aeb5ee53f3fa1bb71a2fca69987b4b22dfa730d
z7c703f0860fc40c5f24496adfc14cd6a0bb0ea323535ef8e49d58c83ecd5dfbcc9d2321ded3661
z01736ced0d73b4f17aeee9029f30a7f7840f01ff4c8f3bcccb781f3b932baeb3d8e92e3a7bfaa2
zfa8a5d9db37a2b6f296866524fee6823f7d94151fbbc616ee275c132cd3594fa9a1fa2160f5a11
z989f2ea39ace7ef6cef0a785b5f44b748a500688b0caf8432a10adaaca75e5e64fb1506b016e92
z9c348021982301e913abd480dae9bcca894e00ef32b053a99cf2ab9d6e3d1e4809435c70dac7bd
zeb437e89c31c65fe64e0a996d30de09cc26c1030cc5bc79f441e0af7ff369426be40e1e75231ad
z098860086e3d9c24dcb9f9ec690a313c252bb5f504ccbac644c4dbe0cd6878b9b9fbb1be311266
z06df7f0ed1413b36e51d55d99375087053f0c3c685fc3db7500101b3deb48c2fc8507271c7b7d3
ze3e9d052bbc4c025da99db0d443f6d957765aa6e720739acf85d0048cef69509e7197dac436b17
z0789aabea02ebb1db6d9d95793a2711330bade51d4cc2658b968b11f594b2680da1c13cb8b7dc5
zfc2c109ba3845d5b65873cf5784b68d0798fbe0a78e4afcaf9067f67a72aa9d9f12e07e2d3ed63
z7a6cafa928f50bc969d3d3272472faa6238ce8f4e0c1b864a09baf1d9a9aaf6cd944ae4eb70f62
zc67e8f903c817123ff8fed0d31ff744b89b0a3fc131d840b8e9dd1e20f47cdafe3cfaf7e9b4382
z5ac0bf42874c1fd7db620e1313efef1d8ac731619e3255ca5611e2ce4660eb13af0a8fa18290d3
z2823aa9d5ebc52628206562fcd4f3bfb25c7db98c2b4b1cb972620e745e86c9f414b4310106926
z844d162b5eb061d55d0f5d2b324922fe4110f31a17b9dad1ce834302ba88ddba033deb0be16f57
z02c151cc817704b856d709debc14f76f25e02125a1d68288be9a177426433c1438f39ec9aa8d84
z80064faef4ecaa1d16dfb91706dbe9298d90a732d56c4d2dd183df00d0beef2094492625f19f4f
z8decb7322bbc00ec0dfdb93310e70b8f4cd73bfd2bd879780cc3be8c6029eadd5dceb0360ec48d
zd4934a85919100a1d49bce49b138b2a80af870720323593626c96d291bf93fd32420686e53158d
z0fc6b03bf2aa0f04059402754f3c763ff80b64cc8e0055d21bde711baec75d73cd8d3a7ce44e69
z84c2c06af7dda61b7b5b73302a4a733e125b64d365a21c310e35dad74bb0740e2b292cc4dab598
z54b5e3968339dcf13d256fca1bbf40a54d5fae5effdb211ead1d2f34ca3e764d27a6fc56fc7fc7
z8cad3c97497cf5b3694b77b10dd57a1d2b0a41bb4d66e30f0e3bf2c9981ece8cb8ceb597065403
z4e0d5ae9c6dd988cd721f9542bf38dc97c079a8249f2a27d6e1b5cb8c7b78f3be582d8bed00bae
z6f6f829da8da343db5199bd4e53748b96fc02327339109d335613e817be14ef83b3bc77a65dadd
zebeb95dc4d11929f77cc42f2f7b3700b7467bbd6d89e3300148326a926c609b22a7d508154e376
ze2edcdadfec775ffe32240158da9b8a1ec6294dd6136a701b9690f77b2acfa04b1a37dbfdeaaae
z89e0111b67d1191e0e5bc86a282bff3eb8fa4b76c679bcc90c18ddb0f13a8c862900dd254dad5e
z269ea67aa3a47fbb22e87befb70440de95c623fbedf66b7f8db81374e1f7f6a436a0b10a131b71
z8450a3edca5a5171a26ec2b78e4af0a89a60af0c8496b11bf67e5764cbe578fd1ae46a5d4d5059
z8d033da0129802dc5bb85401116c536cb4c24a45459ab7ccf07d8f0ce219ab7600d5aa8b06b1ce
zb76d7660e5baf1dddd8be458bc218c85a398564dca3494b4d5aed59a0fa83c803f8e1dfafcd91b
zeeabed16e79c8e1fa980e1913a6297f74672aa2d022cfb8f5c9ed2e248a8b6760a0320829e81cd
z4c28d7fbfcc1e112c8ca7081f02bd8ef023da92cc45925bbaba449d4be7e9e0474fd5f447ecd4e
z82f429a70292bf317c9339576b3abead8431a38b6a229e470a33b7a4eb49b0104f897ac447cc4a
z1490540c31cd3d9f3007ad4e396c51ea74c31e8b72080b69668c800e72bb6327dbf169bb80113e
zd5f4a547fde3c553c641c2256ef5e0f662ac69d0474802781205ec37b3aebea80de2514cd81edb
zcf2adb48670e97ed87a86ce35e9f6b5087b7ccdb0c3d16f8f2964bace617b7210a8dcf27f97704
zc08f9be04e1f717a9b10cc81a6899194cdc9fb650b7b42ac749de4be8c638bd63e2200914090c4
z7cbc6a36ee499456fa111638dcd7116a310bc55e442dc280dd77f488174a2d6aaa7da5c14d31d5
zb8bebecaf0eae3c401b4eed8ff4ef9123aff052b44786e9119ef979a45f5780332403a5d83dbc7
zcd3cc2fc197f2b0abd6c1b75e3fde803f7328af5b6f12809ce848df604814a653617b02095331e
z3d7a1f4b93d95c49db96341cd13f7ec384bd347752d1e467ee9d7d9a683b2d15fe4ca6c890ba60
z998d7e51fb10b33a4fc20fd63533968f668a1020f4f84f25c9265330beedc5573f2fe6c830759b
z82dc4c55d2ff7793dff4f10fee32265682b2dea72f088fcfdc59af6a430a8787bae8b9c7b65905
zde38d8b9ee86efc8bb67f9c3ba6b9b6761d004c2ddbac030ad9ed6fd0b924247fcf62cba1b747c
zc3c0d16abaec0e445eb2e7e173e95f93283922632bc6341bf28d143ad6d611ad68df1038b74f66
z2ec4a31c12ae8a1d4ef58ce4d96143efad61958dd9e2ab07efa405049e0eeec86639ab518182fc
za25de7785fc29b1e3489355db3801cdc17beb5c15aae46a3e6cebf1e77e5683ed2113bdef07cb5
z0f373d75b4eb568712c084185ff01dee6ee4e1fd160b16533eb49dcd6aa9992680a5c786ea86ad
ze8a9bd2c0a890b3ff326ed162651cee0f7a7123c57ce01d676c4703b4b78698a747f8ad7d9fcec
zc568389a0bd7543e0b63c50f084556259f74aa7062da6cccd8f4256a59ed1bde94b9de545e0346
za4006cbeda2bacc1b4b2aa75390a409a6016f9e1d4a7e76c7b3542a627a669defd9215bcdd6d37
z0512f399bad487e0e6cb72d9bbdb69a612c5e6da49349a8e3f626feaa397ac49ca74cfd53fb330
z7f0c0557db43c31a51d901b2c52d7d1caeb2f3607e3163482a7056d68a3609f85360e4b790ebb8
z41aa1962f61dd9b7b047d60b010f30954c795bd4ea85c797300e888780ff5480aafea4b680c4d5
zd6ba1f4d6b2c3d3fb0c456680c52a6904249e8a4b8306c09f78f518e0cde4623485ed81ea71922
z7955e16f05c173fe363824fbec1db1065d46d9968d293a5d12d52bbfad08064a6ec95c5be18d06
zb1cf5c9daae059b5f0e8b104928186d4d2bb27ec128980d1bcc67eaff08e981e9b932c4d93dfc9
z3ed24804a68e77e2b4cc1b1b28571acd57b7a67b577eeef699706d31dae19c417104b764f3d2fb
z2261aa5dd4f25ca3ae6b8bf1e41f4a92fae2942f3b185e26b317df23762759c781cef3ad26bce8
z06313ae4ef2d052c3da1efc6179384ea64796d73cb46f5d63b2ebffac7eb1ba2edd0ecdb87fc02
zc63ad97f32dfbeafb4c0b0be95eb1a5ca86211cf7b669e43c6432d79e4766b36aeb0c7b0222c62
z086809d6caa7f6b454842153d52e8f6cee5f6a4d44b91ac223834db8cf76390e1a262a87ca44dd
zdb3494145167bb39f299bbc85850eea8d41235e6c0bdf07f38ea75400ea5e2e7ec99bf7d84344d
z9a7ae3df75ca8317e8905a20d2791f9489972252199a12c93ad95cd87320b124f028dc85eb92d9
z04c6c0d2d92d420b21959e24061b1360f2480ae86501e0bbdea9158f6933f0f15b212c8936ceeb
zc35abe383c0e7921e4d681913618d56f963f6d025fb8bf422da7195111c059be3206412fb0d809
z1f887bee09c088a62f439157328e037ebd9e02e1ddb0d5f2f8a0e4178c0d9ccc28564b1164e107
za3b4f86704348ce6bc8bea9873e530f3b3fd91d7adc0bc9f91856101a79ef7b9ee237948987dc3
z3c111b4f47dada2b42593169e65c3a63a127237542ea0bda57a64bc40d4abd1677e4b02d473a53
z9fb7fc969bf9fec96f07dece669c0a0672282d76443a9ea0a4dcde9b3ae9c8cffc9d4c726f3372
z592509aaf23ded8d6f51010427ccc7c8c08f86b2644bc1f9ff983b3aab8e329a406a060cc6e3b1
z3f78406643799fee6a193e3f46b709d34009822a9915d6b812a41b5e604f592b879c573048e7ec
za6ce28e6ddb2f9f254a74ea46e2807411fcf69dacc171907b9ac9ef34f99ce7a3d3d0a27c31ca7
z57586711d888a8f00e426f101d77c339b0311bbfaa1b570d5cd2735c9c4ff16a6ff5ff9fd41ddc
z8c7949793310215fbd676116f111afe52f2fc2ca630f45e51624d677bfe4af136be4af5c75a71c
z315be6cc4995fd39bceed00376cc68f9d9dd9d39812347573163f7c03b9b4eb2fc99f3760d32c1
z441ac69a5c858bff582c0cebd50d0b50a8689e2b8f36ab0d9ea3f6814f369727b132bf9e9f3744
z938d849ba59a74e8ba8d0a244c49e4eb1f83ba77d36a40652478c955fff0749adf85b8f7f1fed5
zc4d17b8152491c3ff7914b7944c68b2731e8fa1e81c8a13dee67e8e25b7af9186d1ade0dd97a87
zdda263db03161cd13e126ce8bab6acd43c472e78d03b894f1e287c01fb3a216029c3a7ad5ba9ce
z0fc0c20c671f89092c33098833043543910f16b8102bca968c9ab41156cbe33e0c9f8c5965ac27
z6b3e54c9195197ec9fc9975209173173e4dbfd151e72e45404d6ad03436bfbd303458fa839561e
z670e538a7b90ecf85f135c1b3738c788b805db7df03be63deaeb1460389504d2c6256cd28d2757
z4548f0a4bdb2c247a2f8f89585417a36166e7e18be4bbcecedf4dbc977d956a7edc55a4abc6b24
z0e534ddcf96276fef953363774980e63087448b310142c62708956a80be43e2bba3d480f94dd43
zc1eae9c8f7947c2748e1f0c45b14d0670c30b21536e1e083957ac4ba874506840dbe80abfb70fe
zdea24003146342cad50726409930884e2a1ae25cb6f07a57a740843ff385eed27f544be2094dae
zd3e0e36ce51ad25e55b31800de450aff12462f870fff2ede9175139fc522abb0d0c0c37e0684c6
z3932ba2489f655d9a9294db54fa03a4aadfc5999b54cf75cda9401807eab0bb1a20fa4f0e5e805
z5e067e6ad6b5195a0cb24236312601d0788ddde63a89bca3c7e3e0cd2e60398148f999e8c19ad7
z6b904a2cfa8d91fbcb407ae54f465f4ebc39e9809c1f06ae3656f4abb80fb1e68280c32cabb47f
z42f06396d02e78adcd22aac6d95edae00938ac8a11ecf6c1a4a0f02a6efb5a4048dcce97bf4d16
z543d8f4e43a3007ca2f6a36202daa4966af0b0d678d6454af6cab7a4a0888b8abb39dd2ab9d046
z44330e60ef881aa958bbd5bde2d1006ce95f528fb04effdfae2a67e130f9fe6507780f33ec41eb
zb8bc58f2da1256df8b16c66390dfe29c342a0c377f1a8d88af73a8f1e0f9550359ca2c9610cb05
zd240ded5b1418aa192123f7fcff7c3ba375b1c6dcc50f16cf7a42a22e8f6ac159874c95ce8ca3d
z4f6b2567e9586a81e56e15f5b25a01233dab9acf73e76ec19b1b08efbceda823b79ffbb9ab0317
zb323e49bfd2ac15fc1a77a4dcdcf75188cda6460b442871e3af156bde16d7cd5dd526c59e08037
zbade18766a592f081b9ddc11d150e26b862afdbe365520184a371569a6f42cfbf19ef4e5f1e128
ze8bab29ab35839f03154c865f4170bf87b53770e58d3f8f16d07d15eb54010752c88ee89385597
zff06afe2278591f917b6b9991718f0d433fb2bbdb78984390d6e513eae0b26829d11359dd2d77c
z577f48f6684dff83269ebeb763a8c58fb6e813796e6616ffc4af4a20c0b7edc5574495dd68b525
z285db618213ca136bc264ad8e4f57deada99cc880de500b5845f008e36d7364566188def586fbc
zcb1b53cc9c8e73199429b021a6dd660e34ccc28b29915a9b4335c33576b1ca235725196f0f339e
z8cd08ab27d15bce70fd41e4c9bd8d7a96f18d31a81774d930d51967e8e937eb383208ee4223e99
z34dd05163487f617718f59344a9dd67f4a8f2e65681b33c94c28167b69f916c1a81176da8e6756
z142826c1941864724d547d94bbce81dff8d97d33bff79ca73c145eb3e50506bf23e6d469b49d11
zf3a61ede68a2d9d96aeca7655f55be5f2d4e46afd069386d65b8694ced191586b14e592103f7e9
z0084aa417ddfca5e889920b46cbb6437806a4ce39712a35592daefb4ff2413d6edb3e8a76a46fa
za724ad3466cdfdb7e06499c9c858522e18ab6170c01cbd3bea22fbd55fa4f5029b17492a501051
z44face1fd67af20bda6db647ed9c1c16ae1610d5fc3010c1c67d0db624c26d73a70b87c1f893e9
z6f50c1a9e64b4102f86620d3639dca590554d52a377531f111e730a5deabf4fedf422e787c55f7
z7e9509e40d9e442a60c441b22d2cf5049360888a9631fc1463167b7313f789d090e5478ec0dc5b
za49b03a9cd07059cc0663695b9fbb7d6ef33b7e9b8b39be717efe19f9a5e519fdaa1d8bf11ac5b
z071ccf9d8db313783aa4855d48fb8a09c8a43895608d857afe9cd62b7fc112c36be4c98f8d0381
z76b3181b49d8629f6a0eacd20a094058c2c187c505b73e6e863eb9fcdf9b6a9e1da3caa5664098
zb5c2b2a1d9e37c3e27cb188257ab537a260eb4283a050d483e55885b619c07c5084e0e1556e7e1
z70927992ef319a4f75f552b18593ddc3f13b21586fada87fb3bdbc64c87e1995cc9159713d7299
z91a80fa67c2e9d33c0a03987e5263fa6cb919e4f88ce826ff264fdaf9cf776aa6b9dfacf5002c3
zce8ed3d6a98385d39e9b2f70baf0c6e3266937d48141ee7941393a1e1e917c0da2b83e6c2b6186
zc853f989d0d559a9b467e4b508087c630659b8ed77e111810bc1c7625dc05808b8fe040e625efa
zc9ea572b6c29062e03ce1ce19dab3ce3b62f41db0cf74fcf24e18556820fd5be90431af2e00876
z7cbda70eea1c46c4c8faf17398295ee5c89f1c5582b4b052141b39908203002172d7e4ddaffaef
z2268cecd48ede98eaaf6bc923ea880ca48956fb4e288bbfb94142f20a96915f974b730d699f1ff
za4dfa1fcd70f7389c2f7aea72c5d93d5125cc644fa567db721b5d605db9f04382e33a3e3e8723b
z6c4105eac78d15c175c7d8008679b6d7d1b91671aaa7953af6426deb0d4d5e441627836419c1bd
z701a472efcff34d045a5777b7eba166ca7c51470becb89af02bc90f4688678778545d60b01ff41
zabc8a347edc8220cab67c1493a0f4327c1a193c93ec7a6da3ecc2e09bd5add9ffc3cdcb17d2ad2
z27a415f9176c709b1790f7d72d2326b6ac093d090d1964da5c7a98d7e51d1722bf164cbabda157
zabe1dbf398b14ec7a004a73a79ee60813ad96b3a380654c3f23c9fc5d49911d81ae1c8fef387f3
zfa7a9a34779bb0fb900c2de5bafce6801eb230ace434387c8f5f00c6117ba8b96feb1c23716875
z1dbcf6102dd30628713eebfdd5ffe584832c63dbba8fcee7218936635eec862caa12b171d5fd68
za97847b844354bd2cc119e89b0a685dabbec902b11db0f9f38de736a7f7f8ba3a08be972446c59
z4bd9ebdd3a7a5612342c36f02d75a738f5c20fcf26bc0959864fd616e9336b3a8efe5e053ab5f9
z7b2ad3a0987bf8611e1dbcc1a654362e0e62dc7d25cc174f9451ab85a7874ddd58298087d94565
z71be3b582ddfa2eb8d7e204292b0da17c0697d487461c6036aedf8d73be37ab3f77d07f6ceb8dd
zd4f367327e95470daf0558b3b8b2794a7908c2a0abb5526f7d11111ea19fba22179d9db76187ca
za352797885f54576b83e8457625f76ff6740c8d823bb3b765a9a966a29c0b32b0f8ea392af4a51
z5ad558770edefeb1a867a8fc4ed36c610e2bf283d2caa33992199efd6e189549b24b2828d17102
z94cabd4ea63a60cfcf0c0d0984ae861f806353aa0a660ede1f84171898f6308119dd15535bd488
zb46205d598db5599d174cb72bf3fa2cb36a4f6406ce2097b8b781a3daf583093fc562c1bc4efc2
ze9e65660586ac77bb40da5026e669b6fee5aedf5f289d568f8a426efbf89761a9d9eabfe3377ba
zf5654e753652d19c5b0a2bef13d478e55e3018233885a8342a5e0af5241b8c0bb1c61782727692
zdd0a1b546d8c8594e6a782b0b946190d45535e04d8327a0aac7425f9119e437a5b4ed171d4975d
z8b7ba7567d4e2aa137f645baa077753b9c40ed3a3aac0279cd6c29797731c179ceea2bbf2dc626
z78e2257d5edbff467f3194580ed981ef357de6a64175698d9c8bd34a5e44317684c4ddcb6445b6
z460ad593b57641c39088fd5a6ddd1e9bdc9f0fce59932db5c183e530c0a2c5f1e4206f5f2bbbef
z3659c5b97a0d4a95d5e9c6ccb95dd168255f405b271ea0358a6b5464087b6e60d6799ea184da19
za1a6a8d41e99846cfa401100057c0843b4c7570b483faff61c55e6e03513cf05d78630603c7a70
z68f28c33d1b0d08aa820ffe699bb1979fd6fa996f86ad839001488422d8c7c977cbff922c0e444
z93dbd27a5f1410679217d20e8710303640420c30b4c86b0625308732d6405e0d7c31c7fa46df21
za8453d47b8590f3fe30f8263f33b4f77311e5c41f8e7915b4e637ee78d4a390edcceb33ba82b10
ze782795b1d2f68e93f8ccd9770c0375f861ef7b73d8b147c8855703c192151c29141f075bb7ea1
z3de951ea92301347203375a2087ffe51a52eee1106f43f89452794c544a0b38415c905c630e465
z93711f76e7457a4529c5e3bdd1d19e5c18fef104fe089cfac7cfbd49cb4c98198eb0257515165c
zc158ff3687ae674616839b9e5f2cc6f59cc177fec7a1c2e8ba89d30268dc7178d5cfd45b12548a
zac4dc243942ea34d6eb71d1140c9fffbda9d0ee1f07fc6018585d144d4743379f9bf564b6d07f3
z64b45279f5792ac2b3a1539c15403677987572198a5ec1b0a89748c4e0958fa02205e408799c19
z166a90f9045d0a98f26cabee3e2ea7cc4b78c5c880fbe98662ee611c599c2886bc540a8faaa630
z410a2b27df42b429c7baae5fedbb2b113219ff42fbde14f592d5193135344775b2d8d759802751
z949c7bc2ffe4481c84783d31e18022d177e6a5beb3239952705fa04ea418a2c3053e8f7cce4146
zd9ee525d00836c282c21afeb9248480e7b12fae6ac7ed875e2d4957608082e1df56210d750f40d
z36f556b13305892c7432fdc869a6d7c96573369e11300ccb0ab8dc3c4ea8bb73bc21059a062f95
z22faf80ae382e6d11dfdeff0fe8e5a8f057c9dd87930c1281f7989966deb816ec787639f390c26
z475a9abd0aa7f290447481bc6fe28ad2d616b79522fdff972383f30e112a93e728747e6c188825
zdef47bd5c39ef1cf07a61748dd29758d6021a3c79a02a6a6a5996674686cb19839414b1643b2cb
zc5b21bd1e266f7ba46b3077f6d13a2ee7c6e9079cfa7403dd050c26df706d8a6ac41d960bec5e9
zb5b75b411aa3464bfa3fc8c6101f1dc77ef20a102ce1d6873c9d3564451ce36dee15173debbe5b
z7fc215b24f41639a7f05d135ba925ef5460243d37c100999f74f3b59c78ce9b3a7d855aa810721
z9f9f5622f9aa0edfe1ffeda06daea3848eea219a41d98c8f2970a946119bd1a92ac5284db4348d
z9027d16aa698504e67a6d1888cc037d92cb1d0c2266cd523bd1c64372aa17bc6b0800471b2f494
zd885058e15631ad0585d38abeb5ac6a271f778fd24ae07be2755ce42629c27469f25aa0ae38fff
zbe5f2a6c62fb74e14e9db9c55ea2539697a05a94eb6abbbbb47fa3a1c870be7e2ab5e2c9657e48
z37c0fd016f88aab79cff0293253bf3faf760142d6389b617e9c476d3d3b2243e69f6f2f636b370
z96342187899338a45ce7adcaa2347e6307ec90a89eefbf248e1428a430009fc192e09cb330c50f
zba63ff1337791a8582c33ca5e2ad330de5b67437f1b20c11f8bbd78439973926357e239e158e84
z2887dc89ca6de090beb59f6de80a27e65a107ae1636bf08fb9b0eebd041a9fd5ab742228508e1a
z4baaf7f4ced9f116244d85b27e60486a12aebfc3c2fe5e4003da700ea6aeeaec82c9c12ca910e0
z021b517181b4489f11a98db2faf92cecad2c5bf7efb03137c472b2d7e969e2f6409434bb10e594
z4e78758f5a94401feeb724428c37b99d5c6f1ede318a82a5165a05247bd3924fc1104a2668126d
z680aa65e9b97b2c8080118e2c9029d74c71d36df3fc6fc5b5689d0fb60774445ff6e224259a797
zf76a74347ae2b9bc8d79fae808fb6c429195bc5eb45052e4b0e0dbcbd8922a09247a56c4419eb0
z80dee30d13ed332fb0ed1a1156936d3360fdb903320d90699a7fdd125f40e01ed6030f5aa746b8
z6beddd4d4bf44746a8cb17bbe90adda6bfe05e619f8e9b635fe6feaa47e181374da1f3c7db8516
z278e2842c465c0c272413ee3924608d157035e03c3328d8d9320bb04fe8b8edd86a8a175f5a18d
z3cfcf01d75cca9ad0066b0707d2874179d87a3ba2bb8e539f3981a211cde6885de77d8c9642ce2
zcaa48074cae6c873e13a3776e992c7b5d9cf0408937734a4b813d6fb4a36e2ac9f7b9894bfb03b
zdba0c634161d939ccecf615fb7336c0ec39e3cb993affe0a395756332dc605e1fe80701bb02638
z70f15b0a5bf2c355c69af3de0c45145bc1e52cc4181586bb9a942b592ba798c720691254d60093
z2a1afdb83bb4fa9a5a4f4b851472ad819e64ae46b6b4bce619574e302233dd0d3d8864f35f8168
z9352726037b7b608865dd497cdc81e91b6f25d44b877f96673abd880fa16d60b51339328e83770
zadca34de74f40c6db623fa8a0d964ad4189e12b2173656c1a7698546bbbdcfe67b33b089c54776
z834db1d5007b8266ffbf74f6580c48650867a6c7e25da46be3eba071d315fab94ffdb88a856aaf
z40111e33359870da319dd946a1b543a1336775b32ba6b7aee8ac70227ab8155a6fcc93accf9c3d
zb09a4d9103c7317d79f2bf6f742d051c0406c5240326237aaa918b3b07d06d610c796a6f2498f1
zf4c3392d01707cf365ba6bdeb9f75a036d880a5a463f9220e38b9ddb1e03ef2e82a2c979049d67
zd21edac900eb9ff3ae9eab98c3c4f3c1dbb794e8c70dd6f4bc7ba4d1dd806cf8e2798f9037ca1c
z9e5b44df73a057f1636bc6686147a5d914ab3754edd200b4208d7945d3b10760fb7b44a7fd4037
z39dce75973ed46b1c277508649528fef9c258d6c6e97891987b7593b141185c1e7c27ea7254c5c
z403a203de9bd25dcd1e55e06193009e84bc386e3a0ce27ea51da777a8134101ae034237451b796
z123b22f4af2ea4601a0343811ab0a594a84a44b9d7f66dc1ee89e4bca15d6e7beccecfcc6753aa
zc5640d97e098b9d02fddeb5a6d5d0ccc0da28ef5e466f675f1c601c4e42ee59821d6313cdee14f
zbe3b3d07245718cf1f27f5f4f99f75eafca7dc6d7ead6d916fad09d2115da27f1ae08d6bbe4494
z87aaa490948a8008b8141508f0147107a70a9a6138c37aa5027aa11ffcb0cf2235d64d1f101859
z61e509dbd131e74598ccf911690ea8934cf4ca4244812ffc2fd182ac27e12af6ee48575d5bab2b
z9ab366d08c2186554e147b9d1a8eeda806ba5f595b4107b77fda5c7e5eb5ec1d5fb8e87a23c549
za2c89fd3a5e9546f82fb4811e376b8b364c783a3380731ffe31162055f65b311f8988ce97ca2bf
z005fd554a0153b1b8526a52fdf9a61b59560d1a1685237e338e992669494a7daa2d5932866e08a
z2cedddfaeea76bcf7036b987681396725aabedf7403ad08d8de55b955b142ed73b5f5362e20b23
z2c11387a8e27eb940bbb144b612f75fffa066f3b0892502c9e0967c8e09de11480f9fdd4fd342d
z960785ae053aaeaf60c92a2d58bd02636ce277e53172156f51dd8349ee6983f612552358227149
z651d5bc5ec98cf95c7a8675f7d6ff4a2b1e0f033e35e654ab82dd257b7d1d0201209eb16cce16a
zd9cead4bb5cfba1938df20d6d2ff2633e81eb00c4213d37f9e766b2c8c441d33c650942bfa3aa1
ze365672d73c8d0cd66a0e322cd5f0363765494a77169b0777527fea2a2dd1dd1251b873f139364
zc58c02ee7c713df525f720fac51a1b87af4582aab7c3082ae9a71aad0255c2076860a356c560fd
z6c50b3bd730ca8bda4298a6ed957ba4349abd2986cd6e6014cef0fe736fa803bf069f557fa5792
z754afa923ccecb06b4eec87505d82df0468c60eaba8a7b156f0752b072b8592f430e6f660a6d70
zb8ec95206df9aab20b7e06d27837cf530fcc89bfd794178fb6f6dad6ef3c1803abd7076e7edc40
z2da6ce43d2ba5ddbd0cac95c6a48128d303bc6ea15ebe8106eb5d0aba05c7cb0193c9daace4041
z18ceb6097f1561365ad0be6314208377043844fc318aa5efb83d593c1215d7cbced8397e254641
z014339c5c1d04b3df586797beb44ee55d8c882e7237c664992ff6d0742d70c186723215822a145
z95b947f2327acaf439558c4e8afe01fbca361298565320ce51bb8b9475d008f414a62143204d24
z70bcc17adc7211d4f42d591015c2e51263bfd8a278aaadb683b1e466678c502a4a0d141e2e6324
z8e0ce1244403be2fb5e4a3d55c109ea4526dde1e7f7d927cabc3b3a60df6b4a75fea7fb0866d75
za2964758ac5ee047041c66cad7d23519377709f3d8e9bd5f2d79b947548f0960add8062bcbe4cb
z4238e816183c56bdc6011e7b4292b1da0be24c98f1c2f508f339e056cc21d7c6076d56b934b824
zdd5b088a3c7405aba7e6ab2189f6ec9c56e7fb06d5bedbf8bd3407e083823e2c91f4eae53bafc9
zec7f7320b9960e80451514afda9fc5d0bd8fc293df8723b3202d7d675034608bc99967e9a16d31
zfbb867dcc8f1a43c0bcaacafcc82cc8850232cc2a553dc52867b402f4587561a2dda596afd9b47
zb3c2da06433a252e166a84dd5852e8f6ccd5901278063bc7a2d1f1fd42cced114dd2fa54e6ca36
zea4954cd98e3114d6e00253d1805ad9bba6595a14e3bb6bf044e871af89cbc9b08b56284db4d13
z980228993ed6550273f59bb3316d06630be0faf197f3e031ec2b58bd1607d9629c237e5daab547
z9fca1e27272197c0b46dfddf49b4c4a9cdc646731086dc67e9125b300d8641dafa47bbb0971be0
zfb11e3599af4b8f789c8d577444f7ebeb452b2b12a32422f9c20a7568332f90ae994a45ec63f80
zc9739c87523a991243db589869662fdc0c935dd9d5439e08b754cf7ba41a521a2baa4c1962b604
z12608e77f26cb00d1199eabf56ad3c060decbef96546212b14266eca0a5f9339b9cf268c7e50c3
z1088a27a9c1e531d71bbdfd00c6b9a63e0d81311bb84779930e705c05294aa4e36a9be15fa6b48
z6bd588a16a2ac5a20d3e66d6b3f9fd41c48789fb92872430abad567c2b545bf44d4248cbbe2976
z7dff5855f3e077b1c7d152248f99f8a01ab626740d2788827b65ae319fee9cc764f587bf70b61d
ze4f1cbfdb4f480b1d78e071a6beb7def13a14c0add00326ad26a42b7ae7132170e02b2181b8dc2
z0dbebec984b7de97f857d5902df86acdac3e0a5b47fb7a0b35e9bac15b33c58e36777aba6bc8ca
zb8f938c276a8339c6fe9e544db563b02aadd2ee8bb3ce3a722c15e33bfbd09964351410600a6e0
zc29b12b6aeca81b7b7996126a379d4dc5389c64ce653fb6a809cd4def093678e0988f7f2224fd9
z9a31c10e74c5609f7ced24a74b1b97e5592c8bf95d23661e710eee8ddf7a92a879aed5a98754b8
z4358a84ecd5e524d97351e954cdf73e83501b641e642730fafddda56a683e6721063d1e2a56212
zd48d024179c296e13ceb2c85b7775b72f8512f879e06fb63acf8908db3b79423114b8075b1589e
z58f578d3dca7564f5b11cb9f96e9366bfec9d645293af8a9c173f4148ee75d851cf237df69daa1
ze453b7c0ea94049062a100b0d9a4688e8889f62cd4851c205c297d58663837d2ad224badc049b4
z0a2b74e1d96ee46be577796bf5de217a432338aa76bf3c337b5d079da70e561cc06b9ae49b16c2
z2a096d87026be08467d4c5c362defd78bf93438c3483b027308c8b69244ea0fdcc6801da052e29
z56f84a490d3ba80130c7c192caebf3e4019a8f1d27edeac2c294d6a178b18d62195d2d78339ff4
z7ace11f85387074021da9a9609011f1f3fff0171678bf3f749d4763bda34955cdc9cbab7f4bd84
zd059684dc846aa6aefbaa0b975a67ca85a71a65bf9141fa430e2cd68f294758dbd1062cdac2271
z23070afd6bc63e321445abcc8ce008730cc6187d1b799d65c6fd8ad226f8e4467c07c0568a2ed7
z5951d293e5e509dc1e47ba59ce775ed3a38674e82209225b772158d6813b1d156ef72309b05e04
z00a6b9c0dc8eb80ff9b201cf24e53eab6f3aef01faa8a013e2fbbdf6c2ef07789de86af5806763
z27f6d27e9deb0527add90ab8781c6f97f3b10e0e196e1a9b972194d1ebeb274b1b3308a3d49050
z97b5cd327ba96de47bd705f94807b5e006fcd1fd95c89100cd2a18e88e600247ae7b447445fc11
zd0abe1c7d9f0541a7bb40a5c5c4f79ae0b702dd1383d27f2dc404574dc4a2c526abc96e2a18884
zcf01278cb93ef12dbe770a7d74397fd649e4254e62ff1700be4362f66fa8ac8358d2b5787b1a11
ze9550377769c6c8a196cfa930effc5e6ebd72183a45c807957eb8b64183923ad865095dfa9978f
z20af18ca25d5c11ec489c580722d13318394a5ab3e7f2c3a6030fcd9a84245f743558a83c94fc5
zc84f8abb1a6ca4db655a4bbeb477bdad8f846ffc97f9a26a08e8e7e45d5ce64740dae9ecc3d078
zcfe0eb2944b5fb16bb7367ee2d45fe22fb739a5b20b5c3c6f1c46d80af71e67c3915a8dd985e39
z5567df8e6cb3037bca2d32ef1298f0eb147eaa7085df3aa8e44120d41aed9ac0369b1294377552
zcd466f7487fa2c0c115605331181ed6830facc1b4e2eec4d8be309cee21a236bff9165d9a234f6
z98d135a5cc93a1be1ab6a21b8f662c01befb373d28658d837a150c09d64d2b8d590fb09d90175f
z59021ad2e54799e59115f6a8a22f46401a1e09b27262e5a7b01edf5f748b77a63d36e9108e1eb9
z339338da9306742d05ee6d4dfab28a92ac86165e57631899afd9f5738314246f32366a381690f7
zbffcf7c32e2d5d4897c0d7f7ca430a262e38efca683cc909148ca10ac711e93a64dd8a2b87a182
zc30f1946828424a2da2acbb4dc1a712a43824967134f6e01d5f8a5f1a1312aaeaa53d9f2147dc8
z66b04d7c30ae01ef50209c4ab431fac3181c80080435e3d384b54c9b756cb19583401314fc01e7
zb09cbca38a61c15b1e7522923cdb6a7e5136d59f0b0d83c40ed22f482ab362716aee7ddd15ab9e
zf3511a47605d9d37e267f125c9fdc6153197a4dff9c98b47592d68a28fcf1c27e98b1dbde3badd
z28214c729f4a9cf8f3153e31e30bc7bb03ff05f883127ba1c2b38713ef749a41e31df9fea0ac5f
z459e6a9d279e2084f1925f1676f756d5dd6356f32a4b5fb1563fcf85d35457a3dd3d79d94bde38
z7891daaff4f141d9af4f0d4e7859ea0f90d77851f2868049b6658298e55e96e18ddfc80da60022
z18404f8817cd2c129f33d9839df5ac117abac9ceb485464adde3f0f2fb1ed53fb4d3cef82f3526
z35ebe0802b1ca19c7f97cbbca22cd1b70a2931659a1d9e0fbe057a8f91fa32c46ac3569c6f06b5
za2c29dcda91ec7ee568b0ee510ed8bc2bd1138d2c3929db2fd7c8ffaa6f1bc57af2f27deaf37d2
zd6e6cd6424b6531d2896effda1da36544a3f65e07c379f49a55c0b3da0e6db976862f8d81e8c2f
z31718119d5ed5137716fddaade2252659f65c7c55f05a9250d67facc584509e491f245e99e8411
zc82ce66d7c2120839324e10d3184ee46e7b87669eb5684dc3517f4056e6372c03be1720ca5fc86
z7d0a9f4df463065ac416141aa2764d9e2423ad4ae436758e986035133e5c98c825dd86df6c22b0
z5dbfe3326514db3d64203cb6af585542df00e560b4b524b29aca4a47b8656402a9d993db3f39c8
z4b3c2a215b6489f300a3100947c9566266619e53f5d0e3b10a19a34432c8af59b5eb44fc60bf40
z25560b140c9777d16af83d0ca24a4480d884bf782a9f1e92be3efcf2ee4137be9b4a4b92d7df28
z7908a86b99b2966766975a21d7cca1ccb188b2ab716438bcc8aa9264e07a2fdad8ff963014df8b
z54b9558dcf0c49feede0329e4cd32c245ad01cc53050606248996fb8f89ffb6619afddc2b2bd48
zac8625a21acc462b461c7b71a20e8a2c8cdd42cb7b2e5ac9e28d09a7a3d77d11e1622fa813002f
z511cd63ea3a41eaa3e2752f707e2f19d022962d5f17dba0afe369b9fa551c1399849aa116980f3
z9c6f0681c262480e5d46b582f808bfc897ac535aa9388750c8a94140ddd22a805f4b6220f8fd3d
zf1ad4e949d69a73b94930d8c84ca38fc67b153bb41e0fd247e1a0f5147825863cd3272eb16699e
z7f897a0593733f4312a1899243d1ccbeed2c8c39f51a9dced5c53d1aeff5256a75e4b0c1094a75
z8a0cbff052fac093954e195fd056199bde7cdd6fb90ed52408b3090f92f5ff688fed492b0dbb44
z3f2c8e7d35f596bde0f28c88c9dbf1c201b085c31099c953675dd13bed0c030ac98d62edfa3b50
z59b1f63e98732e9d7d3a77298d0b0300b0291a1a73d2f9a0aaa3888ae2b7f97627f61d1dfbcf0e
z04609a276108d8e2c484ad2a5d8b2b58febfc3f959f4650d9e515b6a006720b0839c37a991fd8b
z1494eee987a878d737da7e8c41f4f04586469b7a3e89b440e9e286d367552754cd6dcaa3c4423f
z5e240f39c0053fd51c01a0e38f08f7c58974e47bc63ab51653b03c94d3c6f4f7f0bb2b86482ed3
z6de0e8712717342b951b162edd2185e598329a79ad1c2ffd488494ecaf64a81fcd8f969d960780
z383842c47f5ed09a39f342f8883cafc7b41891e5ca674150a48ee76712213ac2bfd82373fd9ff5
z3633a7cd4ad2c8f5d7f6d06973896893631480dd1bf4228890575b266939bfabd7e51a1f7c0246
z7183925029d2d85e06d66f1c4cb9d7cfc0e59915a57849f8a78283d1249520c82836fe7c629708
zd19a9a8f186211b74040c58172189133ffe3b790c9cc581d38f7561451ed7f53cd4c56f4a916b1
z89ac2d73de40fb88b5afec5f3c2d848a041bae0a1be8d4cd040d0c5ef91c0d3d48b24bcebff7fc
z80c17244abd568d86bd53d7b453420f8c3d58c1f62f3591159321be79f933bed8ff49ded5c6e87
z0543773c91db9d2db4c68adab378766d45419cbdeccb1a269218babf95d33c133b5452c9a43891
z93752311e4d13a0768d7124c3ab86234b2574e089000ec3b3fa6ed4dd2bc645d2ece75d2dc597e
zbd7693ea8f4c74132aa5cfa7df27138f65a116eb0541187b003eaed4da2e4320b6a8e7645cab3a
z379c5fadd9b57d5b62ff507b6fd619b39a7df132d8917969bb24be791e4e874502f661ba22f54d
zeec1afd33a64065fb4d8c9bf2002188d8fa91e10a9d8f5c4d471bad984d4cfbff37ae3119d3caf
z3e52a18e27d30c91c42fd7668db1b5f12ca35975260f1cf6685d6a5270ec3d9022d01fc949efe1
ze3ed002a6abb8aef3f367ee33067c2b0efd981e7bb4ca0ec41393f1d18583ba51fe2bb49bcd08f
zbc7faa4e95793218556f1b4803f48118376eeedd06d09b3198a87813a86290681d629899dc524f
za179e74b380c7a95e7340b06aa7e6510a26a3393f2f443304f718dfa16c492a6281e998372abab
z4ad313b63e9cf73c3fac56a4f24a0867e49c196e0b91918cc895abe2feda3ef54d18eb7042d2dc
z465ca6075ddbce3373e2d5d0852d5953f80a87e89aa2ab3c2548dc974d30573c991b18c248ee50
z57a3d92a1fd524622124ffa6ed6d13434f718ad6b9eba45130adbb804001ef0817681b3d63b05d
z267a05d3cdd4f4a944816b0ba1b88c0a98487d7ff8ec695dd692eae7a840c6f1270693b3100863
zc6dffc714f1be72ee20cd5d027c5bb89c9307944f2f901e585b55ba11d769cb8578d4b4ecf196e
zcc83222c3b883c77df3175d990c4074c646dfcfb942f58330bed155826001cf1fdbc18821aecd7
zf745037c8b819fc547b75802957bf2487f4777ca4db8c73731e7c4419d51a40f7b7f18d7cfa5a5
z28f20a6034c5c1556694340a7569c36cf7ab470f9e82d56b1f8e66f7decea22f09545d2880f261
zd925a127da0c0293d7edfd95495f619e01564f04d6a31cc06bd5a7990ea067b5ce40586157fa89
z89618d26685c2137affcc9a4bfe911f328fa463c72f2c417c6b80383d8b4896d99bae1d2170116
zd88ff5b95cbf40d748ec3abbaeca6e3e5f8472640bf949f2fa5c302d4b2d69f146f67c10e45b8a
z57e314f954a892c30300ede7a75665d17d296a9c01d1a78420bbd63bdb1b486da87f4b77219eeb
z72132416db405ad33667f3b6a83ba23b6728e4de448de95bc7228b932d0bafa61aecd73d526860
zf3f0f2e9cca986d95b28bc3b52b3636dbfb7e767fe25eab13fd44cd2c4f7bf94e1ae7ee55478c5
z8ff74d1d3b4929589e51c3693cc05b51563b21d467b452d686c3b3c535ed499ae500feddabf799
zb8ace4f9970216ff7af4f1e95924a1d0a23616df05c114727ca14c650df9e24d4beef5b04eba0c
z42c98c585c579af562c22e57e55057909597493238eb0dcc9dab274ce7a922dba6237431016bef
z3138a724d81a1247acf7f87700c762b64286482e38616e46a8c2dab7e96294efacd9855da78e0b
zc10c064e6909d5fe0c29c63d2312d61df96b2ae915a5d857b315bfe7bc705c9cdf6a30e3726fc0
z0a66b58546b71db87e0645259ef683c6b444a4e23f86edf791459830ecf88c832d9f35c12e3a2a
z26f97369848104c2e6530a595d12ace9e7def262bf6843b14b8b183629aeae233c94d90d176168
z6bcbc80a4e38c9fc338f8544cbebb5975a40322b282323d36f0405bd6c3fc1914957bfef32c916
zc31a8c7ab384ab545d774ce49e7be9e20d33eb3a08ef4a87426d32d3e698a9c666d55aac58a337
ze1828203c260b6195b92c6b574d7a7405f5a946a9c56a74479919fdf74a9d93f871e8ca52fbffb
z39e4a1499c3fbef03550c1bb23c7c1776376e9a62d56f37db46693ac5e27c26af065647cb262a2
z29c4873d8290db13c3c2420c773baf879cacb18ad87fa6ba116b3280086b11ba632ce2a222fb41
zd71afc3e8ba2933c7693a9997b4e4cfb64f0d76a7844d49e961c334b1eadf340059bca0bd59394
z30929b618c634b2110f256bde3df0395d9fe021a566b50a2d8cc9d3c1c16b96d93d5bfc1e83935
z21b553b9e82bfa9c9c3044cd52c96e67dc79f1b2e4cf20c0cf3d067f91661d1e7cda1ef786b5f9
z61225a2303daff8bf2c4020a20956c5c2073d099f04e12c80e01bce4733079d8bdb9d3e1cdfa8b
z622f07febf539c5bbadcd3339fdb255b51337fcf1512473e96c840669b37cfa88e432bad4c551a
z439aad3778a8fdb5e12b86a8b10a2e01c029bf0d6bb4b83ee6c00c4797f212c99f985b0c62d908
z8b2d95d1504fa68f4d0d88026a1da580048f80127871d1a6bf456552cdd64f23eba565ea0d3619
zdfa7bc6da62f31ed8c6484cf39a79f0a395f7b9136c8ba2b56af6d640e078b7c8dc8617d652abf
zfdf23501ebb394977b639ff7c92ecab3fffb1128c83248787e50ef6b63263ad5fc9dd5a607278b
z853394cbaab907ffdf94b3b0ecddfd2f62117216b35d3ab6106cfa0f11fd0e261ca87c6fac640e
ze7e467d940fe5bf22b3a98159ed3679c7cfbe3288e1a73f95a6a193f9204a9cbf60d59d0e3b712
zfc175ac5f4a19244a97df02f4047865b066ee3544793357008fa4290bd28437ae9d9f7738485b1
zf4092732b4af1ed1a1e1e5bc53b0048aaaa63dbba3fe599e706791e847b0fa418ae62277a95aab
z350ca6e2640040528a2a61ca55e90a0f5568a5078bdabef313ef3081daa424572c04422098ca4d
z8d5dfd1b64e17e5cee12b1b7a682a0db94d6c58b9bfba9be27d796208c7357b6c6ab558055e8f8
z2349ff5dfe131187a4b169e8f4ccda4c4d0bacfe5f0a12f5965f9351580e4578939a71b0479437
z34650817d0274adbfdc0bbf94866c4306a9c2eff05216e81897c26adbaeba2b4f5d9c7cb671a81
z283f45d8fbff90035628805c547694c6712b3bbd077b4eb30549d9532719cc213f612caa875d16
z0eba728f440f9b82470b01920a5486db3f2adf47895fc36ac4148fe0473dc815176da4e3d4cc76
zf6096ed2f7b44a62647012809f0a751f94879e03b0a0ae34a5310bb4bf33681ffb03246e1cf6d5
z39ce3d292b067b197705dfcdb8fa8190c19bdf1d346f9562b2250daa8d3c11a709e7ff9202142b
z89b74656e7ca490ff850bb5fc5c1af6c731e2e27c4699926bbaa14f5f8a86980e703b9e0179d0b
z2a4a9fc4870c07119a0e538c53525b5e81ab7a4dae82db3ea05d29435595e036c49461340d876d
z06d7352d0e5f1177c27a4b9a8f9855817f2ab3122c5df1e14a8084990e678fd044b19c15c0451d
zdbbee33e3b95ffd3dbc705d0428aeab158feb0215017a26a9521de0652ce55de4c202a79897d8b
z369fd58e6174aa53bbf6f2ff804ca14e3edea28c0922bdf2e83ebcb0f20b4745d59b87c58fa9f0
z26c171d9d1601cce52ce675fc289ee5e62c402a40584133e62896ab1275e11334a8b3e91f95fef
z0cfe857ab2fb845b277c39332aab1b8070d870bbd26adfe400a9d91ce2aa2507a2094834cbb5e6
z0520d13f4c566cc5cbb29ac399b762ebf2e6dbece6a80b6dc56232b7e176c234ca86c76b074108
z0a6561dbed8aeb96f6cf8fca2f32be8ae42c92f6a239334b087537ee87bbae2893efdc9a3bbe6e
z78ac78a2f63255ed1fed61083bb957dd4e28d1cf512b4b4daf15d0c1aac70842552c320f9b17de
z759bee64daf20b3674f9752871043c3daa784825bd2c56a546b431736794dba2dd280ffec303a8
z4fb18c3ee1c6f34eafddd2621df60005885d30458cac5e940bfadc5810e69259b5aa9fdbdd206c
z8f3d42b0ab5cbcd55cc7388627c449f63fda165c097c42395c189d1fb77d06dda38205cd9968fe
z323a2cdd40619bd1ce5c73f325e22d32b58189cd1e8fc54e42944db7e689c52bae907cbccf5b68
z6b317c357c162eebb039aefdbb06f5685cfb4f16038b1fb4149a6052536b17f530044f7b67dfda
z40f528ea2695a4c9be3c7f3a30d6c3d47097e2e89993f5e748faeb8e26ac4f9a13bb44a4347952
zf4a715ca9fc5be65acb1ee2aa7d850d3be69ecf335a23b7f69e7d668b7254ef5a29495f8f908ff
zbe29f914cca35ba0d868fa02ac3323c6db47a2d495891ec03defdfd0c090dbea3f8ba667931a97
zd1a34ab3d7947533e9c390149c89575f7f6ff588708c01fb7db133e7f905e74e7ac7409503ca2e
z080c75e03e10e97ff81f1973234cf42e4f1137df88a0745421c0449ef6c666b7d316c587ff6f34
ze0f6e2cc8d16ee8b474c995ab53ea95b90c680571f8f7cc12745cba5ef2806247d0f1328c0a39b
zd45537492d7a9e1e9bf5a91a2956802ec1abb11e0badd52645a8a8b582e518f0bea90761a5f644
z1171c4740d73b444fdf8ab5fa921733f44386355d315f5c7b519e0fa64242960be9c40e9444014
z784c9f54ecd91e2f05e87b9b9a44c938e9a997e4e28468766b9b966c5b20cf310976ed2ac21e23
z0b86023d7f2a25245cd6ad4d5ea9ea7b267a4493581373ae380f3997b6c11838bcaeef2da49f2d
z771489ec32e5ea7cbfa67ed11326653847cf5f8b12e0961b29b2be65b3dda841d44eaec3453bf6
z180b27551eebec3e1e87565063299f72e2671a45ab01201d509d60bdbcaa6bd39163ad77b7746b
z855895d7066d9d37113a3ddb335d7043389898be63868cf7a963f06f9c6e53fc12337b38cb8d9c
z31b99f9fcab0fdb7b9fd91e139c7887df7764d1a3dde78e11cd4e4ab49d468792a3aef9550ebce
z2e2299d23c91dd4d346342c5657dd88579730fcfc466c89e1ec04721d411096b3023fd5315d9d7
zff6f29ee19424883d5503cb32c36b0804bc8e6da7ffa594938ec468d0dd3e4f14e3c959a6005a2
z95760136a240265040635f2cd64ddcf7cb075288f42bb806c19c1cccc6ed5935f0bdb38e7f9d53
zb1a4a8a9ee3ae87a1da8ab82901ac2ed9773c76cb47d7cb2d17ae981bcf6cb4ce5d561a6eb3a4e
z02c2b6b7c7f0fba0be9c49b2f9b31183d44fcb580a746e8cdaefaa29021f6d1ef13cf9ca9844ae
z96577d9bac447b774dfd0c5f0a3cd561ddaa840543583ebf9780c2c259ea36b20b290b9e0ad518
z5a4b6af8eaf4fb3a472d005d73d379f44ce12032e92411f91280a3123ef02a088dee20b6189530
z8dc534e4b3bdce918877133ea90f65693744f3b68a18aa67d9859898781b1898d88b9126d23be4
zb8dcc8f233a0e2d7e661c6ecf4c1e7e445a1abbe96affff16c047d59e2b98da38ae283a71e95f9
z165d28ce4a6ce36d0ee08c6245a3712181d536286e795c497456d7a15b78d1be7c8d3455c2a603
z3a95079565e02d2504701b9f06f6a94e9b666c169839fdc6cc07b99ea23eee84f7721b75c6a20b
z6152ab2c611bea2b5d32a17ddf6b886baac9e43b9f8b45640874ef6ba14b74b2e58c0cf7470624
zc1058f2fb4c3a6c2930f4cfc0158397bf693304e9b93eb9d1ff6cc08403421f039c2e431b080fd
z761474dece3154c0c1a8372639ebe867c6d081f0fae001c735a57ffec9c7101959fd6768c122f5
z7eb67359583e086c7bb93f706b72777de822c92e68cebd94d09e051d68dfe8b9dd8e495b6499b6
z609664e0b72a80755b2f834df3156a37b6ce74e0cf5fb6730bd40d1fab30dacf6dd6f14a939b44
z4df9a1dc7785fdda920a6720ac8ab42af40b32a4b1cacb0e4e8752b449bf6f7776458bdb3fcc70
z0bcb9dd774813052fb06f25392224ee2bec00b512d493060e3227e790156e68ed20397ce43464d
z629d8a4ac0fb37e10e5589668a7e13c749b5a4bcf02aaed723bb9f93538bf49ffa80519a937121
z13d5d709151127bc617be2ff10a5526f2aff52efd14c13cfdc9f98d3cf5f57b6f79a93659fbbcc
z57b54787a96a491b2593536533ca0396b963f80e20d5b8acd59b8e6620d18bf8713f0ccdd9e799
z6c8d1ce4b567283c61f57df184536769a5e47f19d129a3c793561a296f23c6cc7f4f54f59b101d
zc1731b79ec4ae506ca54f905f18db35349db376af7494edf018768f806d9101826e8520f5fceed
z13eb299dc97961f32747c410b210db359322e74c4068d79f5557714482e440b556f014ff040ad3
zd30c50a9373526b4ce617d7be7db0baa6029871858d662d4b2b204883c618d2447531ffe465bbd
z57ceafa2834768be05de03450f86474b2b84df82c97efb3aed5fb56cf0267a9d6ec1da1bcaf702
z17b40935ed186c8d4845631975fcdaad9a90a8538d4a4600d6bd17ffbecf27241303b29c51dc83
z930d44aa47b4fc56057ecf13af2dde3cd68f248588b042276e26fc69d6039d154d4b1a937a1657
za77dc006b32c785e1a0a519a0aa14c7ae215c51d61cbd795f1b13038e3f1eb9a1c06b1d9eba925
ze2da01c8ed93ea3dce981bee5a9866136c0839e07cfa786af9dcc8feadeeeee2bd831c94c59eda
zf9723821d804559e2e5729a9904b3288c02c3164b34209b46dbcf19507e62a5fc1d96901ce8a62
z2fe1496aad2be59be8375858a7b26027352af0ce160d6ea741cc6b6219f2ea11f6bcde4ba9f436
z830d2da17898be3f1e183bd099c57adf88998d91208a4c43f1a976ef3bf2370cff849afba85943
za550cb77315c79027ab592bafa879f3aebeb475431a895e726d44764782352eccdf05b6e6a2606
zd7f0e269846e22e66ddf8b94da5a7f03fd1d9b7e596329097b194b9b8d080e0a352bbd0408eefc
zc7eb44cc7164a2656c540fb0154c3a14fe7042bfb7dbc023c99bb486a2861d86264a0c7fa0e18b
z6860f0727384fd2f7472ca011ea8561759a8a6f6e9adf3da9a683d1cfd1d81412d99d1c162a221
z7f9f97ec7f05ca741b9252748b672abae9a43b73ee2df3cbf0f02a7784005e8e3dcd35a19d406f
z336e227c3795253c19ff89a031225c13cbecdadde6d699cecd8630122aa75dc29017a85c77fc26
za2ea7bc3a9ce93357a61a02165e6d77f3e5ce0632772e16d5806154cc683f053b79106803017c8
z41c452513847cf512098db24427acc46099b96da63247931b53cb99aae80264935e75e58642e7a
z97e019642a181777ad417924c525faba085db625c081ecb9554ec248810b7303ae4385ba7efefa
z226a083f56f379b181662646fc4fa2dd43b8080832e46f0c5c5bcdbdd8aa3616ddbe25611f6018
z13c9d4d224caa0832c8a4a4266d0e5e21f0ab3deed589d726dc8fb245ebb6ac4b388eaa925d942
z7956cc0e99bd75825c36f0e8cca22901c00d11b0f24d0d79db1c464ebb7f8977f0e341becc9060
zf259ceddb627c226dca80fdf436b6033f9a9a662c5301ecb3908c1d07ed285272ea5883e698d00
z0ba296066773322199d0698b4ca4de1007377a5f24dde158adfd22dd77239e02bf23fc73cc8ef8
zdb1ccf17f10fc68647c9e8893b12fddd8a39f14af6fd7c46e68e7bb2bbe436ec438b7da8257023
zd18aba16e256b77234911d2748acaf6658e85c0ee3502501b98c747b3e100c651f44fb4f3108b7
z204922ba46d40561709d70b84e3afd24e2c0b9e95342265db29e8fada141cf393529abc06e325c
z542fa324f5007d712f9221a97a1a41a128451d49b30a6adb18aa14bfe4028686da552de941e0f2
zcdc61ef73a7f9fc86987f0d3591df89af3957073c503aae033e4769ddffead48d5198290680254
zffe4c9511524ef6e1fb8d72249566e65a92e340c3a9338bd1e6509b72fd32095db265e06239e27
z752fdf0277f20a59ae04d397ac8e4745c275ff0dede3ffbb7c5cd0a53a028d9020d24382ef47fb
zf6fa2b36094a5d09ff9d424b91448e1058a93682b62a178e82d0e171df57511328e044ff86a19b
zd57e0426ad796a0c967f3b9c2370cef4ecb121cd763d5ea16bb65a0d7f1598c9a2346b05677124
z9871bfbd966ffc88259877e5b21b5adc23d0f460563b849b027ae43c0b5f267b427f48fab25d3c
zda561cfab0d9224f2d6539960751f3d72efeed03b8ee95174d9162c4e9be094de37de8908d515f
z6312f8d1147984cb74604a53ea9106322da22ce47be24864277b888662a6f1028c6eecdaaa6cbf
z2e5f9e7d76aa5c93acf5a5ac41f7c40fc854d7e4101379a638e3cfe56b414d41ae57d5070d8810
zafed744497b21e49df15db6342e35e298935a695babc492e547ef27acc3c4847701af174a85a37
z6e7bc3cc9f77c3dd619a7cd825afd946ecc18d07cb2bb48f047477dccf9ff0e00fb2654c883463
zb8a776eeef29d30a021ea58981bc83d9b89888223fc4cd494bccbfa02760869aef0a1bd96d02bb
z3250cafe61050c0940a5abfe1531c2af284ed61c36fae4372224e2faa6c6a646ac1eb06d6cc66e
zb6c3525f65be9d038eab10beb8a36b18f19ede92a9be0f510759cb79572896eda2126b5d46c212
zf2175472d86910151f7b633ad63dbbd101276fe33815a0e624ca4277595ba044aff18ed6177b4b
z08ab2be687f43ab1a301cc64be5ef64480cd961c7f17c697cf83c060641bbff44e6b0cca6e997c
za288df0db44d7e430d0383c86b939bb61bf99f7d0e1b25ec16deab6a37d0067c884783121d4dd0
z0b7932f38db252c24fc5ec60be19d2a6cbe8292034d69faf5ebc8a1cb1b6d59e16222e0396ccea
z77f07f61ee1c16b3a80d4e7125d35e8ea2c3db19293b34389eda8d9a17a869c142865a4377c344
z01e55e799168a3e43db3e8e1933e7d39ec0a743b6ca223295dfd5665ea1ca8f07c1e371e0a6fac
z1a58f880711be39cba7d8f55259eeba942f362357cc6dcb8d0eea3e6ecadb25a766f67c87b9d9f
z48526b07eea285ae6811574523173ab0a56d7cdcc546c73a6a64bd6eb6fa7ccfffb8035934af7b
z75da4f0ffd0879fddeda911fda130e9f77bb26b2ee09105fcae1492ffb42bf26373eaea8ac5dce
z62cfce8e85c5acfde1a748d4380e73604f82d6f73f5ae9bea19e59507bb3303e0fe05e23893b64
z803294610c88b9228aabd584619675b58deaac9a61cdd037975ab6c824982cecbb2efa15acebb6
ze8b424713228ebeb5248afb63c86e92868d27b3e905ea43c433dc3420a12aae93efa1d58e46992
z1208cf9ad8ed7bc0a76b3808909d4dbc49e7242e24037ab312cfe704b7bd6cfe81e548ba856e1d
z3d711ecf56ee2fcc0b91b61e12d5961f2aa3ce7aaf52f47111fced92a6b30294cb5825129f9e13
z6a6b4ebb1616e7ef87b4fc5b74b444dcedc11793123e65b9712aef01bc3d8eec45fc778dfa752a
zce9a55d46a6059c7e106d16cb6a85c00a51b0e4c8efd000b8d6758b696c41e3996f034854c84f0
z45920930ba2b368609325b70545f9d66b6f7b6ca37e9a1c69b87d23a94b16bca4b09ac00ab9c61
z0e4f85632e1afd4cd734914325491e083353d9bfece3ee90ff60e49d199a246db7bbb234385952
z57430b629e591f6a9d7bd1d6cdef4e6f96ac29a1ff7b9ae7761bc171482b019b7877574634a7b4
z7ffe8af1cad3be5c81a1a2a8a4bc8b8cc4c1496201fd7732f7833d2c2795b53490937a1d61b645
z6c5585410e4761d64be988b2ecba5488d2c499033d7d71c18fcb38daeca10b8c6eb6189f07011c
zec4d1a280d208eb4864bf4af461ceb2f5e3b28d264c86d898b552d1df6c38dbb5cbb572078055d
z1b023d2bdf4b559706b7ebef6a14c16e0b621b901c47a32bd0058be94493278edc4ee6c9313b06
zef77d989520e65c589ec44e4258ac4b2934898636b47850196bf87a19fd5cf8325ac3d97755ce2
z917978a29e8e7167b22ad8a1500af3f85b691cc3b2a9ba1459f099a95ff792eeae5954b8dfff96
zc08d1769d4c40024700f23f67655523a32c42dd88818d250ab561cc936ae7704730c3351eb4790
z689c866dbc7ff29ac0e00ed71a9c17b327d1f5d0ff52c311b5c7d81e7adaf0c891dfaac26c4c93
z6a1960e79db6aceede2801961cc2b2c6aa6f269c409420ce5680a2e5fa5a9e3f889dc62e5dd02f
z4d7432c468291222261b3ad171f510f9d96cdfdfb2ded13f0f328b1e64afc5b0ea7a974c12010f
zd393495a02ad1e1c7cc0084e5a39dbb7dc388f6aef5bcbb3ee90684ab9fb3089bc1d2badf18dd1
zb3cf2f149f722ccab1e805178c504ce112e3225b58425039e9f72333d998a8ae4c5f70b2e871de
z9d9af2536fea8f2ba0e4e89f098b689a80cc846e43f7f5020c9a00a89dcea9873d4c3ffe5bb337
z227e31779a94509eb7c73eb246a4280c40b77eab59330c5f1518ca48f0c2ad2f4c329b2f1d4cb1
zbef95f381cf3b6818d03bcfae00b4d7fe950a9bd2faba58d4bbe7bbf6518b8cdc85614972c0ccc
z6f16ae2a055ced3b584f58d116b28fe12397e343f91bdb00e0290f3dba6ac07ce472fbcfc2124f
z9aec1307f5fe9b6bf70d2f126a30f3d53ad12e9ed4268299a0fd25d450b8161ba3ef221c2f207b
zde67f6457e5f63120b862345166356e0f04a4d25369a760c1185273978c430901341a272febc6b
z63f13e3bc96f8cb4269f38a4a1a58e9235943503369e7bb4bb8030776a92ca8c84e9a04569091e
z33c4e9b06845df18b917f2559bf27bcb412b18a2bdaaaa7de425160ebb3b4f8909c418709e7106
z56fb90561316315d9106641766f3d237cfba00e38bec952306901607882302af4235a01a3b33a2
z3331d0557d21175895bac278ef2458898ef6c44301c5d843e97d14acfb134dc7f266fe2f68e852
z8db7e21129dcd9c14442753baaf4e96f590fe0cf64467cef828988bd2ca6896761fb51b7673fc1
ze74821cf24a1a24fb2794b51d50e0263cb2d2b2cab03529cd8f9cd1c3668a25ce96510dd933a4f
zc6ebace9ca03502185f79cad67f296bc3687d59f7657be943e6ffa60462dd06e3dda7debef7119
z1224d84a47439ac05b3f46540d8178ff0f78b3e05e28e741d6f7699b7d3051dbe3969f6c0c3353
z450c2c35a2e4beb9c4e619d5962a8f424da15d7bc524cb65d1ffb8b1d64e0f95a85e5440c045fb
z66868367dc7452f92b87c391dd857431bf5ce95342b4f1fcdf5042c1d0b1369248899c3b3cff5e
z8c111d43a2f1f27b3b9999727fe04252a5dbfdf6efcc98b45d2ce74101948410a5a9bca114454e
za63e5190ce027db97fa0281bca5785bcfdf0acfd108afe0e5428a5c99c13aff875943a12e89b0b
za41426544a9e3c38b901f09ca884b8923b4fb6f1bf32b22d85678251ba6644fc114476cde0e4d8
z940e6abfdceb3cf131aa7600bfb177c8cd4dece8ac7b5bcdeae756b0525e9e29b0eea073270f0d
z1d0e97701cb1630e1d3f7a2fdff39cd25afe0fe9d8cfbf6c06b7b77d2759350bee7d5a33f440bd
zbea1ac2545eb27c5e3a9bab41ec263efca1d1d864ad85aebb73117085e6cf0cd4775d7d5f636f9
z08981769059a3339a8a316947292f5e34d2280e3d3c0fe2ed7ede8dfda795424c447b73d4dcd7c
z8a7323b455b6dfee70de6c0207f56c331f1b0d046e9a457f12e05509c8868dd815d9253d3dfb14
zabc13fc32d1e1d25d02b0a426e567753fc199fdae87438ec7b7277ec922f29b0ea7bcf91d4eda7
zf87fc125fed913e58ae32563619457aefcbfdf398babdcb8070b480e33980e754f9832a377bc79
zefdc5c9c510c87fc9a3a4e07ffc4b53633c97c8d601fa79cb9971ee56f498ce1df89e71ca206e4
za1cab9aa47af2dc1568ab75252bdb915ec082de89c6622002edd2f101c9cb274c6095b69dd8f54
z494bad9e774bff72a7491619627eadb9284b820c2a43f135a496ec03d7ea0659a25bb89c8a0822
zb5a13858b70c3a50ea0f52571481a98fcc41713dffb8f61fa614a0887c98b4c730d807471a7b65
z456b40a09552f3b5d4d2998610556028e3ec1afd99ca189c58429f9702d95e8ad4adbe56b86249
z2279d4f89dc23b22f24ad28246651ba961b9e040d90b5b832dca81d08f07fa568aa97beda40a86
zd7417e6c76ea8a55786eaa53e1ddf96f596a1dda79d5712e70575bcb67187cfafb98d3a3bd7a8e
z45c92fa3f49e9847ef5cda69a425b7545504e5504f79659aa9dc074ab8023746bc416381c93a15
zf14cbd2d9663d254c69c889ea41120e85afb0f0f6046210501b5fb3d82812dc4889e37416b6b08
za0db4c0f1aa76d16fc1cf900de1e7170a589fb51013de43f75a542249d6988a8b7a9f872ed47db
zcaff3335f18fd63a8221adead98144d7a6ac6aafad286c230063bf964b89e309f415b0ccf16363
z82ed46d29ea2903160f1fc112fb7be07db62b22fc10a7472d9b8b5ed5edd506b07625f7e9b654a
z4708f0419bc0d40c24081a730a8ea9e200662b086b9135a6ed28942825e65e678fcfca036e0e15
z8a9b74e9806ba1ef274a37b582c4da73c03de6051c872f7d5afd970774b3e993977299259dfadf
z3dbe36c8cec63d6cc6972508d5c3ba4ea661086604b121b4cd8c102929817f17e15beb6147bf20
zb78818c1cd02ad778395595acfd41a454aaadb536176d5453ba853f8997f3bcf83b75bd38074ad
z111a09dac6dfe7e7eed8556b15c61bcd6fb02cf3f014d0a9f4ca063ef63ab02003ce960df67006
z7950a5d28ffaea03f561e07999a8010e301b9df97c1be414455079b68f4887c8dc3bec82d229ae
z94af4b1021c693003a01ba6b8098327d4b0bab81aa2eecdf06298748fd225d20be3ba92c850afa
zbb7693f036fd89f37bf94f4842bd8ff959fb173fcdfe605b70ff98980e4ac74185d4ba86ee4b8f
zf97ceee3f3e7e409e43cbbeeae33aeb7e320c426884e1b58445042763e2f3f8af83a136016859a
z27d1521853926534c380dadba9db30fee43e1b9344425615e6aa7c2d86db9591e6a6083c2eb599
z3743936e22533a3bd7f9e00e7aa15151a7db7268f8367794494779501368fb47aab75e536386db
zf2eb946315b54637f14f61f2fa1ce9bb65396efbd33b884b232d1d56b2e2536bdec35a47b6465d
z0bc932c73aabc2cfc5ce84ae98dd9e22dda81afb0a368003b02d0c5a25987bcc43071660939c25
z1bd8f2ab1344c2d91e18a0d1e23378cc0357353cffcebb773eafb8510498c70f3a04f0f7fd01f4
z9d79f88bfab450e4c9241f0865b785c7d34cb057018243259fdda333eef2cc2efab6baf46325d6
zadba85a6e475f05aea89fa642a7a8876eb1c5ad586c94cf6fea0efb10cef9ea99c096f785b2958
z9000db6dc5a269c1766a1657fba476c126a6ffda26089a9562ea54af16424b26df32cb08ea183d
z192e44282356ec73c2a280a1b245264548bbc35fd70460f2665e92c45d462307a489ebaf212d54
zd149ab5e7faf66ccf1144f8336b35f214ce8711b8f4b852e739cb44f7182399685bb8a908282bf
z4817c921920cb6132ea0ca958a86e1e6adbeb928dcd3a96c581f11d9148b4e05797eb1c057b1da
z6a63807de320610177d2c3a64774a6e50caaec381c538a5f48ff2571198af0c24a4eabff06cf32
z3b87d550a3a4c58a6cec6aa98c12be0fcad0e36fdb6938eb90a8b20e4277650e5b9199dba15b42
z07e011d60db25106599c62fdb4a5b040ffa3b0fc0754e5e6e5570eff918cdfc75b2e2ca549892b
zc977a205d5f040fa421077189e98309207b175682773659b6320630f773ae98c4d1e4b1a95b803
z8e723512065fa32ec2c77bc1b0d400a426250324c4e6ac089784c9f7c7a7ace615c395435557ce
zc8e50568d5aac2a16d9fa5007c6ab2f45e4905f66d6e2412249c55219d5913bb852500dc309488
z79b89acbc43a5cf25b109b55b5a5b68f49809829150ce8e05f752ac2277666ed95e92b7f6093c7
z059fb9dcdfdc223a84bfe6a4ac25cffc7145f4aea7def5db892d304c559deb3632297676a6a1f6
z68bee3bae2a23d32e379b75ecd6bcff08b8dd479e226589a56577cb9030233d8e7d9046d96c7d7
zf904c329cfff1ade859f3d4cdfcd281e66dde24be31ae6cf782a7e689d25237a5094d1aed50f3e
z88bd11bc3ed940c457f4738d93ab687ff8214c1133ff8be99ba7f314cae521c20a9b343f4e5ac1
z180d445b28da80164d27e4451a0f8546cf4ef7c4a4a31ed5138912d407b5c3a6c833b3a27c3be2
zc72936735dcd01a7ab772a114f43f5b67ee300c6691136ed213c7e49275316385f6695d796efea
za2de7a3425dc5c244c47b3ea0ac2356f7f9b5c769928a112c2e263e140809899ef0ebbd52fabf0
z8dab22d9e9250507f68882cc38015c300c8581b6649b89bfe2e85946b79f814dd498eb2db8e187
zaa3cfbf4ab1d33ef52d018088f16269dade72dd404471156657443a6076262d9a0d00b904d1455
zceea5402f98d4d3ddfc8a896edd70e64fe0c3ff356d0f8c73e20a7062090a1575cdd73de412a66
z546108095f3a21dcdce1c80d2539bf3a7b375ebe02a207b095c73831c4218c786f473674ffb52d
z880c3b57f68d6117c69a58bc489c3117184e22904ce6990b4d3408e33ee2610a7c956bf728ef34
z79909b845e4b04cd901ff5a6136b3b22c8c086847279147cf4204538c0d4bd0c0e054832d3b2e0
zb154c4e9de008d52ef6eb2ea2b0a280c11898f40f0bbbed6216ad285d0076cc940cd36c0c33fc6
z537f62177d738347a6b78582af7f45e3a86d837d790f38ac0754354bd7224612c1c1979b15a773
z899389d990091e222293d933f04f6acccfbe40af387f9072e40a0c99ed968822978f78c4e0f202
z05c6fab6d59554d9f4e66e9d3b46724ea80f523054c19c2b4d362a9625d27d73ad5eb12f293596
zd09d719510d9858b42064b3a852cd63bd84c7c4efcb703e7007cfe867c55cb8a39ddc689c77b8b
z4ca1afe659188dd171d35b456b8a07141f59a55b66cee76f196f4a663a0b005ec6e3cffef5735c
z2a1b4a5785bbe6555cb5a1bb69d89fec21d5b287b2262eca314f52487f0325a859764501cb76bd
z67fc6784991c82ea61290c00a340978854e54a11a0db53c8e2dbf0307dcb56d17becb091560702
zd17341b15b34e88b90d28f559262f6b2a9b0eda16caa55b50eef8de213d8aebfa3b22e765d9ac1
zc99e8b56406ec37da80864bc9667530ece58dad37c89e63341fc63465a3ad01e5dcf9cb120e57e
zd2e93094749b7c79bbf839d5852454630ec38c1265fbb405ba4ba4ad51768d586b8175057f5598
z7fa64fc9d1f44b04a3f01c6e0d0cbfc2e1299f6d3259c844b138682f59d72412d417b98289a261
za4def951ea439bae0e0721924ad5587d11c95291c3856a19405bfe6bf8991239c449f7aeea4019
z4aadb02e61282ead454db46e75cb5b1a74d76c65a24fd0b4d1035d0abdf5f5f2cc2736908a384e
z7ea73135c867edebd86a4c8c24fdbc25e560beb3fa49dd688bca2a583c2d84a7ac60278f9f7fde
z362be7f7198e9e12de5fe0c63820061f228b6461f16f6c6ed770bf3794076da70eaa2f0b5295cd
zabc3e0bb87b654c722fe66bafffaae7a3c722dce8e09fb9f32d142c171560728716374db70a9dd
z76bae8a2e0c55fa542f6a65517a2178eb78896359dee5bc774c923221044c1b036c1592d289523
z997952c5c85013630893c18388243cdba25319cf74bb97fadfa0c20b81ca685ea6ac6d9d709110
zfb530271487c215d882963f7b821e6455d6ef7a7d13d3d97cf6353a176c000d7af4a68f4456315
zf05f1e908bcb77703bc88100635dea5e2f196e3c8151e9df8996bf54384a9b11995f65f0868fb9
z307ed10ef024a623395cc9b413829082d6c1232ec5d5c9a436aa56706d9348117c2a679764e39b
zd9726239bfa9d3f9669b150edd9abab38943b7d58cf7229bb9f38311cad52530b26d71732b5f65
zb0b816b3342fbea079324bf4e9e0bd616671ced279571e6663e04cb9272c5319c8ca5fb54d0266
z5b5079d83d66c74ebe2d9673bfeb42eec6f32ac7538e5062b16aa642dcb0ff015a0fcf4bd3537a
z62484981ee74c62d8482399d45e2814704d0a85d7b5f0e52a63f5cf3073b3ca2d875a97c019d90
z9b02c638345579075e87021da7072c700b700eed2d94b2d05ce8f5cce6cce66c9521286bb1e0e9
zed238229ea925f70071f6a6718e06bdd56dcaa9c0949ab2bc94d8318ef4b3e8425c1aea8ba09ee
za92513d73bc64c23aadfbc2febfb43f4cd7a28947cf841e83572b1972373ef1e493f8434e4f9cc
z622a7a000a331a6e6bcfd08e1f4bbca6b81f41466502ad10ddbbf3ffdd6fdeedd2d0f93c8a8152
z2797d7e7f05de718fd1a4bf46f812e463ece03528a727302ef5c8d7ecf95126db03c178679a401
zcd3558a6c889f35d25abc681855c842a8bec641ddc96d86025a4d9cabb752d409be862c100d260
zb397f4d2eadf39da30763d7a1da3cd4a9feef0a697912ce116f8454c524ad7de9669aed3ea85ce
z7c93ab931fd823a656a1d4fdfc515f30ca098aeec3be58fcdc2b5b09ab3d31e0e49b6f29a54bb6
zd6b2b95e0b9d339214ebb85dc23be3ad1a2c16bbe136eea97462fe107d14519fd2e7b4708f2365
za4fe64d844371cca6bd1cdb30132690c903ac18d8529ad06102a02e5ad697cdc22f7a66355328d
zefa093226f7b3ea53dd4f08f137ea3c5d753e9deab351a96a06e3648d675b825ec3fa10f3a5e79
z25e48e3896565ef61522e701742b7885dc1397acb6d473d16f3c65625ef4e2e39cfbb1cdefd4e5
zcee126d09b5d5aae755580dfe055eab200b01a2312a11c2601fd55dba95153f0b2080dbad08d28
z7c31e3ae5b600c41739d8b2516f06c81b09b3391adbb9294903675543f18b8a0450bfe5e2be2a6
z71839ba1048e4cd38ba49ddeae47d79357ae7af6238e1bc89c36f1263b54898b183a594aa04c5b
za6d2cd1f96631dd0c13e5b668e1ec725a1fca0f188f54e9d9b591be888069e3302127755c662b4
zb4828ac0a0c80b50e19aab8ff1df6b30b62d6c323d9b3641da78e3c7653d8f0b8d3ff2c3e927f6
z1f11e32298de7df3a7716a02b65c8cfba47ea975b9f43f5d900f854130c363121e0a7d246464a7
zdc42c3d33286f21ac05bc776761245cf0d895f565b9d484f7831422812340b07f476e811f89c1b
zaa677574dd9ec3c536c72485e0f16ab655b3bedbc5c48be335f1affc9bf389c5bf5112e81b4c0a
z5ee0a987e18d17bf2c89989c4cc9f0e4684dbc7dfa5fafdf9cc50001ac919425e0baa3fbd90780
zf3fe59596bd6d41f31e87e0283434e8684cec890b63f5595462c1eb443c2411f00530e1c66cef1
ze665f1662edfe80ad79a5bfb1425bfe39c4e208a987d68380c33248fd5558f52151e997353cbeb
z1d4817eeb427731d8f67a886732a0f641a063006f012a23b181c7ce77af9a17d3cc64668002d5d
z39784d1263702e80f0cdfe8f6a48762b13cae113412c47f3d7f2952009d8f798aeb5375a940477
zae42c64e726f4a025bb27c885fb3c452673da8f636104ce38c720df9f9b27faf80889177ac6e73
zf22475851d2f8660a1e2b68d8a488c05a2ee325781989c5d1d06833bba0de091f94a895a927d43
z9d9f9c9c3dd921508df1508ba4af8fb217ba737bee40ab49cf6da27d680faf9c5c89d90cf3def3
z05e47a01a3eacd5b9c08b632c1022d151c24e732b537c88b99b2680fe640c154f319be9345a56c
z06df3831e38887612c09c6a1b49d88cac4bc617d227f728ef014c04dd8f7a03bfd2facbc28717c
z048128caf59d6a96b21f394d5f2d108a36135ebdeeb79092dba75aee229a282f6d36246e9c26b4
z782b675aacaf2cb7bc0a9681ebf3f2e4d0644151dcb4d08225a721d1027884baa6797a9d072442
zed60715b9207a26429405066e158d652da00cd3a5e0458bf2378211945f4e55b669f0021bd2d56
zcde0e67803c3100db6dc702afd8b0e883eb6eacb046c7560b120f7c82ae6cab510957dfadcdad3
z5cea3d06e1db0664017407abb9b62e5d6d52bf1103873d3f3a3f053b58df6a5c864ba3cb63db0e
zf8a65c5910b3f4fb797cd43e8962ad9733cd9c19ebcc5c906c987056cd999929785c0346c9fdff
z6eeba23951eae2b0fd64a6fe089d1335c482ba3b8cf77ee06d3b874c490405978f9a58cfca70fe
z6d72b2c16bcbba3cf296645d7dbd44f7ca346dfc13ee41ab500b007b388acf7271fe64dd8eff59
z5c149354d7c4d796a4a7997c85a66b18bd8fd9aefbd753fb12e29350c9b6e07eed92a3d4c36fbd
z06d67c1308f84fa70812839d2d728949c912fbc4e6a2d6017315300e9a642ea2b306e961d034c7
za95d3d68207ab654d87fbb70fb90418fd73b0b68a0e9b2c31f412e6c8e5156a383619e3f2af8f7
zf67428a6e2046a1624580e822d5befffb3b6b7c6c20af35337565ec1370dc794f9c737b2a9f2e5
z5d045e379b9e121ef1ae33e35b520f4800e2506bfaec3475a0528e4385ffe16df622c8b5f31045
z119fd5170bf84cb30fed219635662f24092618fe71e0cce2897aea40aace10e029fa32e45f7f6f
z266115e2744fff78fdfaff0b5ebc3f8aedbc00a904ef9fa8911ae11b22fffda9a69183d5efd352
zec46ac3cbb21b27df635267e573ce1fc677445bb4c7f221e90b4321c9b75e1ef85b2af27999261
z6b23bae8a97360e632d3f22649c8963a98a86614377137c89c36c43bf499bf0a430cb4d0abba02
z34d6cdcd7566f095946ed1c81b1187117fd5cb6e11df6de4e531128485a89e78790e14b4c2cf87
z942bb9f436e70c18f0871cdb1b669a1b5677931574044ba81257dd488e10e4348567aa4825e841
z18557017f48d2c62c26cd54087fd492c374daecfcac1c5023d31f26ea96702a700659f8016daed
z6912db3a2383b3958f0d1de164071d4ec2e4eff47a830a3b22c472879236b5698316df14a4ade0
z9362c5fcee26158eba792c3c641a2f0ace4af1ae4fd7186f9747d54ed6b8db0e0672db4e3759b2
z8b4abd7a3f2910ae9f320328f0c9a93c1f01070472161be8ad7737184f7917145e287498090a0e
zdb898573e068e59c5b6007148a84a1cb35b1a97ec5c3725e97d4f1e63a2358862082e8cba76c90
zf61719eed952c310b2fcc5c7f56afedea801a803ae5a4758cc92a08333faccf2de46b84b451d9f
zfd3cc785f994a7d4320a22ce2b581578d590ed0dbc4fb72caee34a1189f7d6b452b6639eb5f511
z412f41db38a921baca29954103a429cdb8c13ccdef92048cae848118351bfd584b4c18bff7d711
z3d94c068e27a0f74c42d7821e74b56c008934bd7a7f66f262d2d1189a4293750090956d0fdc69f
z82eb18c6d6cafd428db65a5fff6718ab75b9ade9b864bc9c277f37be26c7fb9937a4e326f16568
z0aa851adac643ce70c57dfd70206a5102e79e43d0370ba90c7e34d4cbd501d6cf2488426f8520a
z63a7c74389b416d5d82a0c59cf95680e8cf3a047681d573a778ed8a57f80dfc29a2bc9b83e8ec8
zee8ff5881895584936414d2d2c05822c597601a43802729097334d3ba58a6e8c35c938122170eb
zb61b4a10d4ee1d79e32c8050605585c40c0fefbfab298c99eaa147d28aa9bba3f31b1467f8ce5e
z43041590747060bb3375b98b62ba03c6cedc68fb5310b2379f624d14287aedf62ea81f64fc8ca5
z6427c4c0b329d9e1def4b1e5bcf7aff9aca4edd3f58bde2e7d1e733bb636c4b6d8f90ec9246aec
z83c503df0d82dc70dedd83de8e27e7824d842269fefc00484a20d72d9a25ffc12a9987323d0d78
z1d869b04ad071729c2ef276f9abad92ea135beaa53f801edec8d5997cb3670d109496ee9dfed1f
z9e8e38d7a65bfd8227041c31c1b2d207fcc19a62a9f71df60c9df32f79c831683ea67eab48476d
z2d2e4d5f67ac828fcbca9f4df49a45974c53681e04e610b0b6c36ad5f03ce3366f98d5b856f887
z3a8a91a4546d94f1b4650b3a86955d7ed29000056a0fed62d04d2896d7478598e61e0367a603ef
z737b6ae4730e3ee8534b53202814a121417ee2ca7b4002ba95c9ac256ebc21e3686c5c26513b1c
z82bc5a59270acb22ce57654112aafa081b8902af1839afb8b6aae651f287a16f7a1a38db052a30
z3412982fffda67027893445e474dace943920194b7b40dfae4c0f294f0f4b0049f010082b8bdfb
z7415595c02c813a5ee68d2b827629dcf909ab4a300cf0928a94afb6a912e513b923ca180dcd17c
ze7f5dad325865d690a34938be69f5460a91169d9a3c53b811352f7c31b6034ae339c0e0259e066
z268906140f1281baeb471fbea84ca42557c4c3884bcc13e7da6864f12246f40979f7a8e6c49a48
zd0138b4e92cbe2b09152aadd433383b9fd02f8caa0195f7df6ac81629b34e7dea53c30261a8bb2
z98987132940e5eac1520625dc6831ad58262730fd462eeaddac7d89ec1735222d276e9c9312f11
zb73ce7fd076deffd50fdc61d7d0582904ee44ea0b2e3d36616c6378212f34c935516f6f95f24e2
z96977816acb130249c802f54b353cc60db7a3181b89ef5b66ecb1a9c77e04a478c139f4108b974
zc86fc64511d1b1f77ceb6db4eca43386f256c8c8cf033eb4408ea64f5af352bb596e421c880ad8
z2c404faa8411224f8ff35715b29b1c79284a2e8f92c1f5ded9c32216dcf399284c1a6aa087c10e
z19c6770e467ff1c3cd5079f32b63d7d4f86443bedaceb0f4ae009fca230c7a8f07073598069a34
z306d24d0143e3ee5fee9b9ee5739263c40f4d2814ed6c2bd29a8bb65100ae819e49a958af0b98c
z51bb0ffca5cf2906db2bf530a12531edeb8a717982270583c320827646df51050c9948abdbad48
zdaedd6171d684afe398def87630d2d199edb996f6eb496a175a578fdc79dad0b3b581252259e7e
zb5303558a0ff7c5686ba38bb0eb5948e350a3c75d8a0d622c661be0684008072df38a0381a092f
z2bf8fed04d680b2065f5fcc03c9f2963a462bd072625ac0102adadfe78c06dfc2a1302ff6546b8
zf7d3f068f751d61eed3c1129a177102f4bcb49067ad8d5441082a29441e68f2067acac0890b839
zedc0de69a7f06ea3722220ab87de42f5e428de19756aa14ec6e96af9ea6c38285ff7e2672d9984
za47429db14da1cc2560b7c17062d7a9c176ac1da7fd6cad77221dc92f0796facb3234a683cfee4
z761dc37d3e0c2e4fb1e2d75b6ea01be22c85c3cd83feb0f2f7319a65fc795a1a3241aa4031ccdc
z2be305b153e735d904faae4ec442689cd6f37ccda417d1995db7c5715a316f22d512aea8da01aa
z01a5e9712ccefd84fb258ba15ae3d83d351d74c4b5dc9e8c195a3d5bfb2cc96a1a740c32ef158b
z283a6800c26d5afc9573837e15d846d3fa1f537a51f92320f9cae1a0a233d5d3d3cf8303f1af0f
z767101c955b9451a2053c5049d38d08a28915c953be5f17462bf8776c22b1b0037115cf9d12105
z148ab8088786770c0bfa26f4fa06294c22c7df721ea7742724465e29884cd96930b26a88da034a
z88cab41f8abc943d8e53b19c4f0c22b6ef3a0c4a132fc95a42ec4d22dc9e1499e60eb61a2d972b
z2a52238069e76db2001a8df8ef04a95c6d6bfcf05bfb53665a9d16f1f12e72533281f545bad323
z639ddb34408298b66478004c3e258c35c47e0477add189fb2faacd4fafd208a65adb49e8355086
z60bc20e67afc7f90ec1abb4f1e2780dc8fa74a438f9195cfc5d0041c1ee26ee62b225cfafe01cb
z6e82dc725b8f0022abff25e23889631f816fcc73180396b40095b13ef9a6d05028e2a93792f8b1
ze26001ef7036462d8b2bfe490ba4205fc1a3743125ecb284b8d465d6f6e96955298b9ce6cdf70d
z91b228fbb82e97b76285a549c2041c04abd8aa0b9f2fe3b86c77c0fb11aed597c2cc15a3c8bd9c
za0fea989b136b147b60f441275597490f22c5149a47d77693e972c1cf364cd767dbb83dc25e50f
zeebc9d9b53401868dc21aeb91c0f42b0bde3abb29ae41143476d325a52ada404e4301a063c2c9f
z20bde3f62a4548edc13c4c5f1bd4e00c09cfb26160dd9227e272b427921a80fd962b54a44cc3ca
z3546bd1b98949bf3dd6a9b08fcbe63773fbf05290c5686155ab8e5ad372243bb1ed059e576c7fa
zfedf1149d19ac014bc9f34dbae75e1f12e82cfb400297684494c4373cdd531cd86b0b44ce7d3fe
z374bd57eeccbc7986a025643aba5e11ce649363b3302c95fb89a9820497d36cd7a2a33a9d856ce
zfe9b277d3f41a5bd8ad246f72bd91f96ddf1af173a8f576969ff1ca66110dfe0535b7221b288c1
z8881210c584f46c741246da67a82f3706906d9b6733f56ae4cfe7e3740c339e6c18eaff66d3547
z6e1c7d0463c24e430a5c08db86ffe5beacbd73d93e852b7cc801efd1cd6d157cac94ddb47b481b
zc0e4c71c11104f94415f73be77e71b0c9d8f8ea4410f5863ecb541496a11d79ea6fd7a01a0e472
z70c3eee34181caf362761e57d0c8b619f0bfa1054bc3d49e5b9efdeb8b177cf7acd8c04ab1ba6c
z727a3e52be2a9b6bb3a685a3c0e5380512a0777b3e1336de2e6d947a6412a04d5665bc2f2958a3
zaadfdd26fb165f4b98113bec6949a987bd41b23c40519f8913e0f2020ee15e4fc2b669d3a3b491
zdecdc7e3c81897b38910c0ad90fcccb0a9d88fbad145b72f0944441a2fc782a24cacfe289ec82d
zb75d1d4a5fa4bad7bd55a1b2feda48b260e631f1422af93c900aa0400ee0734c2672f1bb9ff573
z1b52ee3d367c4c6bf15e46f8511a275afacbaa5487bb66625b5bcbac538ea70ce7c74f9b4b5ead
z52b8ef4a752d75de8eccaab73736c5f7c0a000f752ad73d7329d7c38816db77384525e3fc97e2c
z36f37d52bbd434a88393c06592241aaa8d44d6f4a9cb4c9078ec00bbb01d5fd3bd593ea8be5925
zaa1e8b33dfae7f087be37084209c48f4f282661acad99f1067be28c158744bc27dc9e8911652cb
zbb68e7ae775dfaf8c18f141512d2f22835ad1bbb505698d3b6669f549341d3647bf1e0190f3bb7
z7733c592320d9ee9a5361de11469d309da32991e00e12c1b4986b3d3b3c2008ce0fbca1bfadad4
z8b0cd87b8e89537dc2630d4a4c1a09cb73506d945c243463cb598b6e9ed7f39d70fe06043d2a39
z34f70b94d927c1e9626bf046e367f20d502106992eb2c20767967b8ec9309b17648e5038121bad
z6a8433e6ae03f586e5caf4b2488073cfcb3b95877b4840ef130b3efc1cd2a597ffee4d6b8e1971
z5257182f73ddd6635ce3cf3cf1e73a59dde8f1395363209e77a13a34d2e3f1e9e38764bd4d857c
zb2835b6b79b2184c4be5b3dcc04f739d9a91303291b72805a9a8a7c620cfc0bc9f403aadb58618
z73407b9250690aa0c9c42c68e4dd2b3ac6e7e867a6de2256b08062fe6d9d1fa67e4ec004d65d86
z62392c8468b84761d8c56b33e8f45b4b738221e613aee5eddfde27371a270a26f4de22d485be82
za19a0b8f4b999a36c61546ccc2799d4115629029c6c849e063ac70dcb1ec34074a38510c0b3f2e
zde94e10854797d611be37366076b9ff9ac634376e1eeba0e1085c353d3da5d957eb671d85fbedd
z21d3350e050a9b6f69b29e1df215a10f181c81b5d80bebf4ac9b7b57e8909974a349f8eeaccb21
z9ced94e1ff35346b9153742237a45c7dc277ab8fec21c4a698bd0f84660e99d27962f920029540
z0ef00849f8aa335b703bac4f51a0b94513186a255969a830a30679526d7cfcd1181886d59e918e
zd17322ed6dea576373e85a87c495964e711feb0e67e8b1cc369cb9e1e1e07be12a15a3e8e627be
ze269d94ec5ba52cfa51ce5f99d6664af8b168d5df5e8ccabc91e4587010842526dea332c5adcc9
z144d7dd51022bbd1ec07dd6abc5a38ecf0a8510f70b78e1e5c896651e0a38f2a2a928bc31db57e
z612b32d4782b5c19a632e5afc830df3de24425b6da41ad76ba0275c7de1ce0fac4a127c0cc5b57
z10d39744f4256e934644297b031f37c3dc8e97ac1f871d49884d6b97a7043561999c9a7129c9df
z52d39150ea945cc6c4bacceb891465aabb81072a490af4d84d29e4020107ba334a96331c183915
z403e8355a12c3997200ebcb1394897383adc72c6966859a657837eaa10f87fe5578e38c4f749e5
zf94944807e248c59787d4971e2a5978a0d945f0f80c707f0862177cd73008d3cd047ed564430e0
zc643c6328e10a61949d8f90b68094b3b364ca548517bc67eba92909c22f1b568c600e7f9e8653a
z6a46517bb6edaeeae9d01a0b4cd2187aecce885277d8bf9f6e28fd744972a6e6195bc96256d6af
z50e55ed0589fffdb3e72301126162c980c822bd544fc4bc538b9fb2ecdce35f0760a818ea5c106
z6aee9aa41a1c137b4ba4969a811932990af1a977a075557cf63131c2d3fcb468a177e44f3f98bf
zb56fa1fb056582f9e81e7133217fc0d58934bc05c0fbffeceeae1806ffc27c854e0f1a32bf306a
z8044cd15136a952218f5ed80401b3b91f193eb1835b71d16a129dd668b4c322d232dd8297d5873
z1246d95e45390dbc7ca69c5f9ea61b702626325b0afef64c43f121743f912c7622484e18895437
z2e4cb4ba8501b0fee9ae3c7b9873c6732b1db9cb58f994bd22687c13c24354a7abb2f156e36688
z0a280b10e5fa6b74d0a328ccda4772dcb921d1fc1dbe99507d39eb58fc0ecc9740ac043acb19f1
z76bf7942878f5e50762745c2cb10b15a856523ca38c14200cbc5a4607012cd7e73f6e42bf12a8c
zb8e1f062ee099844dfeebc86173be904020a092bb0c4532c0d0bdd2d089f0d2224eed3bf28a426
z7d01161df67c3e0912e2478b26906501913c0e9ba1f4f57b7625b5f62fbd06fce0a13b83b920db
z0475613997fbc206ee52ac352929ad00a5fdc8c4d6102b0cf588ded0aab102ed8edb5f0f310d2c
z5c860eb40775671e2f1a8ecc2601eacb272815f1e0cfce4f5c69a77a9240373c3ce4867b486998
z019b3d812a8162247736546c9aa51a169a6b4006c3de3ff548445d296653e91a8fb2737e16311d
z8a11aac39023085a5c3b5c161e8bb34379d2055a9e0053c684865fc7c2cc13ea7a80a953ec03b1
z8f0d1fbc9770b5254bab4eacf4301fd6b8e3662fb15055c5bdfe1e5c99c5b38a8e678db48b7383
z838c0ca892b4f5d4753aca1e8d57b5567e081e291750170ca725450a64f29c927251943be29b2b
z245dae77e4bdc178c9eb9d8dc8891884ec8c86c41b895a5af18fd303b352c616994bbf346f27de
zc7ffda8e6e84e959968ef5182caedf78ffb297c465b081a79366457e2f62507d181df4a9e0b14d
zf4b0288e88e2f95547436050821aeb6a9f66e650aad3f771f5c8005a32dab5fc7653e5c6656ae4
z297e31cedbf2d9cde5a60b16f79bc8ffbe01e8784e38387e187e62a5cc542331c53375c16b2b6a
z49a6b51ca98192e4cce87f82556ca497c050a784b5042ef0f50462fa2fa61978cb5b33ae90efa0
z71cd919fd8211cc3532a034997edec13c0877461ad047161f07f2956508eb5d3f78d1eb04c9f35
z39db3eeeb1e834a79d39677c66dd642ef5cf7f3bb1f6976500bcfe1a3b46cc614d7c816d894426
zc38c2aa0e615856ce726325f9d399330f64be397c6dc95aea3e5bace611ca218d9f9e84c594ffd
z0341e59593914bf98bd06fab9f1b0d4af99d5e4f852079cc485962542010655c44221429ab77c0
z19976135525d81469b28b2f43e32e5bea2c0c8f9540bab5b81bd9462ab6bffe1e6aafd144d9403
z06c15f015b96bff004d1e8faf4b38c8ff57aad58cad3a75615981d345fd7aa0686b9cc1cbd963b
z3d521d598ae3ec0c84abbe5ed8ff8dbd48bd1ce2a2aeaaf62e40bde8df996fb993818c04956ecc
zc10dad5ecf09d3ea63cd641be14c2ac1bd3165304e8beebb1e07b536a2659a9215166da394774a
zbb3e5f08ae56dfc36072d206b8deea81a22b5f9279f1aca6f2903386997af33726bc9f7df1ae31
z1a3c81734428a4f6ba8e517e480f834d88753910a6a99d3f5e0bc4eecc786926888dd27f5da300
zf8ff5e52ba53100634ea01fd41395bbba15678a044e483daaa1134806f97c5d0e5268b5eb9d6fe
z088dbbfe025432e07ec058594be7ea265c4b91420591475bb4e1bc647e96200c2ba7b16b5bf018
zf0792fdb034d09f80764cff8d29299e99a4a2825205da2caeaf6aef0a5c9b3fb00e36b8999c7d9
z8721b77c0fd67dca90b51433b1880cf3c748ac22ace8cab21f5d2e05c88d8fca8b55b09c0cfd2c
zb4d4d2f699c062cd1b063887cb3a4fa44a3d18694344484c22e48640ebabfffb96b9e5365e2dfa
z88bde922afe94d001fc7a8527af6fc07f3bc8554108760836c61eba5d3b730f9cab28833c96846
z9f06839ffdf9d6b4961654c0b63d4ca304557b1f9115244dee3b73793bd300ac4defb8d2d6830b
zabf08c30b879a0d2059dd4fa8f86207628bdc3e810e720790c07fbc7d27c50846edd4137e73662
z63fa082183a70660b3f21d19504f4056887179e9e86644ce543f708a05a7a515102cc5d8c3c492
z0e8d11683aab844893b4e5f2e9760d212865df992b6f82216e16d03f26445634b462214053f369
z80ed8f4e905067f48f77565f38450278c4902da27650628c27494fd4e704e4d2ebb3d796ff9b85
z9c7f87ac88f4e1f46634bb90c8c93b95d436b0f55d938750279d6b97aa146b259c5be00b9103ce
z4a3464722e724caab0b2c94f080249d06edca165fbd2c4d716672fffcec9c54601b224a42e28c6
z67fc3d8fdfe964874cc5ff3346cdfac8dab7d65fb3a05aea5822bc4f518eb26d52759a632f1026
za3bdc693b32db8182ff56a34486f8aa92af28e44ffacdd0b50951b6887552cab68d7b36d415e0a
z103f0a391a8058889ae06b4073dd58b570b0ef12d790705e973977bac6598c71351143173e1033
z891e7ad15e8a9618fed96f420096cc1efff3c9f0cf9c922e3e91f9c6ab2110d5554215f0922ebe
za1fa45ba296122b876e038102952adfe91ff1d5147938262bc699047340c5078339edd12f3224e
zc19c934344cb52da09334c7d0c3908ab9dc4e04a6fcfc8335725240c8167e51431966131defbfd
z6b5f9bda79eb31e61bd3012ea6cf2ae8ba5a287f2b29b1843a9a20aed6a0334a7ddee1847e7396
zb07b10d3d358ddb07a79484c03529b4a368e397497903b419faced95ca6eea0d0aea8fc70835a5
z7f0c05d7076e8dbc79d5a2b9c4b63905360616d112e62cd3968490aefca19c746ef3048ab70de1
z7c0f44ab98fa3d6121aadf314b62af0c34e173698306c2a821cb5782f4ce6e329d4ed7271ce534
zd1e51350124ea475af99416eca0488c0b114acef152de02e64291213615be790a57bb7c8e65f40
z00f4d04f5f62b2c6c3464033087273cd4cf80d34d65f16bf48d08a8049a7a02f2f3a14b3b2c49f
z2ec2c9906105ba3f89f6221349bbd03833dbd29f3448a974444eb9a47db053ac31086f60bcecbe
zf60ec194fbdf8b0a53882f918c0b8be15f1820c40344c2e0c66fe9f75c99168cc056803ef7c151
z31c470285eab34ce193782ddced163fd00897292ad0f6e845bbec4f27a5ef5cae4806803c98d4e
z6626fc8b6a67a517a32f96b674dced44b3e9ac1631182643a0d45d63c641bc3d1ac5bb63a1780d
zf54565a1d2be323f3038ed5669031a98386d0b13a0556355c6dcdb5ac783efb716a95ecfe38b32
zd6efcea1f67dfff99180d91a0dcfcc295a5386af878938bf1fa542ab34a7cd29ad66fa3806f2d0
zed56a3ee90d04dbc57eee039657c5ae4a1cd61987db7fd1e6ba4ea053d46908e41711f9d235fb4
z51d2fcfecb80585d4ccdae22e9bbc66dbab4ba818a7097c9b4b8f4809afe94ca5631c3e6b7a0aa
zf3d23e705bba8bcf74709b3ddff6b804449424d63310c9713ccbc7c0816327e8a99c166d31a289
ze3a41532f17508bd78342da2545db558e5a1ba155e8129b7a2c2cd20cf7f3d53a84cf3d0e17121
z607f84d6b65c1460b2ee2e1354ab29c8ec3848d1f67120d3e7e69f12524ef5e17505bc79c56fb7
z3885152a58c908b24b2dd5ac2b8662013234442310f33bf4520d2fcea87039af66b4e24f7c0cdd
z5e121fdaa81e4f52afa3ba85bf70a2a7a2d4a4872c2ccaced8be1211f1a2ed99c15d762635c864
z68a4b17f25739d3f841fe9168421886e2e8221cb591063c144b2c2c2d755265f6d5b9939fed713
z0bc0deb848db7d18c2b52422482f1c3a0ad241bcbaa4c5ff561c0b4b4b9c134398b095efd32f1d
zb765658313cf7c01df2a45e70973f55b20d7ac25e999e4231bb6dfdc1caba1755fbbbde4bfca2d
z2955647e41c15c2a55ac9c56e9c396ccf14b246474656a81a6b9689149bfd8166e7a627eeefaa6
z3e28bf214ac3d255c1f3d3d52a10d91cd9d5a8e13d087aec0ad5076636951a82b1166acaad8a4f
z81af5f3a9ca470e01bb6a2de5c3d15fc53ed0e1985327c0551e5e3b9b8fe5c84a70a27a92a4dfe
z2e02a332d0c59c30fc9beab754230d22edbcefc1fa35721c61e65858840fde9328e8d31ab0218d
z38e8db5110b6b054d39d1fc9091fc00a0d8a80f722d8432c4afe237ea7fdedc3b80377fd95e234
zdcb5551c08dba101885262843e8e2e7560f553d934b3da45226335d6d89e91bf8903d23cf7bb1b
z21c40a55e62c5c57b95bf185b51a2d488da6af29563326295af5aada64e733355c0f832e990132
z60cbe070273510cf5c31b6092b87d620a690452e5c8cb14fdb6e25ae5dd52d5283b39e01f5c2dd
z9f87ad802108515d8407318464f229d36b92d9526b6ad98f32ba6c5c6939144f61ac9f337ed197
zde7a10ecb6409703dd682dcb5ebc46f50923697a102cf797ebc28685e129df253f5acccf946b22
z1393af90ce9236f97442714fc98e3aee996ef503743bec7921267a85cc4411fc9655b90bd67a80
z6a9cd623c8035bc095aa2b921799695ea69db93351637b12a7c3c4dd699f7c032a4b78d09e6b75
zfe80c20c434b3935c8fceb5449f83b39222d55a534206b36b2acf8610e6313e40bc364fc58eb1c
zd88d50f8d4f0bf807838a77d9fcb0ddc80ed341b09649bfd4821bc384c2105b84d735bfc099a5f
z2534128d2113cc6f298a917f6a83f1ca05ab3e5931d8bd4de2fde34c38a5f1c99759a6af9a47a8
z770db0d206dd42382eb836997518b703e27fe85bf1eaad1c028bfee99cd2893cf3e6c94f7c59b1
z5ad8cb47bdbbb9f4946982e7e2250cbe69822f3ce76fbfa3ac29bb5ca798bd95ee871909ac60d3
ze3ac89ec3653dc1815c7aa4da41f0397de0856af545fa9131ac247ceee14e2a7729e3bd460928f
zbffefb507e13b1b6f5675d84de86f824f31772c0552d7a45d3702f5ff02c9d536e2a185ad38912
zb04d09c899fef88a4be75f0bfe157cf8bea653b9b741de65fc8d711552bbff8966996ab14cdb9b
z8477377d832493fcbf5b2de110bdb90da00f31f4c42711a0089a504c531ebd8fa22421a9852439
zb58c64ca113a34104390d5939c0ee9b95d4efb25e2e539c77a4c23d672e8633f00e4c1b1fba363
z3caeff746975e5b085a8500e8841b4fd61b42df3eb824dc1a3dcb06af183f3284a3303aa8ae945
z95b119ae756c313b9a004f4c2d88dbb518610fb868d0170f9b1159401aef7d2bea4184220734af
zdde8a58f2a03bcb5ad91ad5b4ebbafe5135954d8a5fd3beabeaedcbeccaf7822ba56eb8ce3a106
zbe9f1a4358e662978947b19a24f16f4695c07606e7c2e0aec89406f9e815d16af602a3ffcce384
zf37ef8c7a315f96e8f51dd11a800e65ca7b3bc02f29f3e1cefe08e27dfc24b7b10651509f136ba
zde9cc660d35c8d456bf6c1103012aac49f9172ce4c21dd9da75778b1e0e0c17c5cfca13d1b8369
ze4d7defd40ea81e992e8323aa5dac54f16e173db8bf31d10f4fe2611973db81d8cdddea667f864
z7bacc8297c09be6c5398301f06dc42dc5ab2ddaa42d30fa68e0a94e795d487aa1b338814203e70
zc337608440bfbed320f53ba2c91cc8b2059b6b4036195859ec21abd9955c789558e2289d91c882
z36bc56c7f85dab4d4f921e73a829dc1d0e3dc207aa91e4d1c485f8a1274fe1f7e88c530807326f
z21cb0ca89eef590ba4ac929d29cab38a49fa7a2ba6decc898e28c5a1c935c15d4e890775230e2e
zfc6f887182e098e4a6c1f6565daa0b437e356d2391285cf174693d0c86b4137525fa8409989c5c
z55538f895596ab86845a2c8a05081a1afa0b9da72118575cfb7f65f7f47ade5bd40c9746fa7bf5
z6b03a97f4eabab4499852e4d71514455a3bd4cf31b589d9c7145583bfd95314c014bf9a08c1c83
z62e049b425efb3ccaea436f9dc08e8bd64070563e2cae185558ba9ecf561897ac6784134cefa8c
z99f6bbf1c129fc3164789d5aaba4506fcf5b9ce542884b1c279a495de666b5fd01d79394acce3d
zc8ecef79933bad9bfc5539161cdc8f85b27f911cb82de647b01ba925752588668344666d7d84ad
z71d6ac6f7fe608faea9c9bc5a4809374220389d097343c164c538589d72161682baca9fb002fef
z24458534adf2178288394f3e2d58cc6572939aecb0fe7b95bf02995b6d0575e8e1fe21ff595eba
zc2c2567d4e2ea1237bda4c5d2b615281f0d7ffab26921473bde7ebefa6cb9d6362c426c69750ec
ze8b93bf246a933aed71fb2238b1c459b1c901e524c5a95b970429331225ea6c653833cf15b4567
z046272289587da2e160e272e0d6444be7134d0db630828f6f5611877c575cf02dc237fbed9ebe9
z89819e35e16a3b67c7efe93a0115164283388d4df07402acdd9bbce40ec738e70185a1301785aa
zd522d01dc5e6d7f7d333abfc2f18a315a0a0ccc8b4d17fea464ba51979a765f59d24e3aab017de
z86f9d2eb9d083aef6d230acc22e9f9ad6ccadfa808395e6adc5dbedf2e6c994f87bb0a5df4b086
z09f146a5ccc20539a8f9c0416d1a28f7b7134c4c84db0d023ffa1f187914849ef301bb78abd866
z5c7a6c849ab17d47283b098f0e5ee55a7823daae9112954b9be1530226627d87d29cc59d4b4885
z89ff1c47c4c4344f54fcd45e6a5ce1e17664b48d130d6e5cc61b609ad088fe2c3b44fee69ef065
z0f670e866cff038a962b3fb433f7ad9eeda868a56db034c23d06492bde358298b50d6ee239a865
zc6d5fa5f1a5fd19cdea12a1b504bf8ea5b568ee5e740d665ac2076e3b14256753e3c7a9de9e3c2
zfc4061f057f5498bfecc7ba195ac6d78d47045efcc7e52814242dc6601af1d6a6b8b0d4b229286
z7416304b58202e25adc2b931352e2eecec6c4343785fd3d746342cf29451bca6ad89755a7d83de
z6abd619caf98e84e958b376a3d21862c92ee82e6d7fa72808e46a0911c7e49f7cb0663d0fafb89
z654ebfd4542da73d5d0ccc9901bd8507440561c813e31670ffcb88f24f7577fe61b2ea5268af54
ze6b1a2bf7377d1734c3ebb9583d2e0bf8e3f4588c752bdced59b995294c3ad7abe0292915093ba
z50202023dd7557b9a368c958eac8371388df2b4a4d46b2b6c2041f77ed9c6e16674e23a185fdbf
z5365b308120060a93ed708a04b0668f905dc6d3069511c6c4a0eff6841654bf5e9b6e955def0c7
z99a8f1b77df052c911528d5a7ca0fa6775237cf30f793b1383ae66407180340e4960edc3bce6a4
z38ec028a7ab9a4281d687bbb40f6c5e4510e142127fb81178e6aa61b90e3ad5c2aad25936d8ab2
zb698f25acbd8f5b8a8e55e093f9c16584676d88842e612aeeba9345cf4a4ab590538cf6437d6fa
z2ef0650c39cd06e9c25d0622bef480e0cb47473cc2fed22b5fdb9f5e2f1e57f5f94b4a00778aa8
zc4c02cf19811a8101fd76d55c2abd3e6fb677bdf23d35541273df321e0e88ec7ef84ae511e1c1a
z2618f474d795b537f14c81ebdee999e85bdca86bb74d2a2c9c476f75b545bd43bf3f7d83e04871
z6b62b55928e083e4d7470bcb0edfabe567c69b518b39fd0732b6f9197d7433e8edc60ffc9069bb
zd3b780525723cbb05548ec35dc08677923ca8906376851f89e2cb09c63fe530a0532d63428d169
z91e228a3f9def2471ca9e187ce59e723288570a922e166c14c4aa3959406bbc6ce63fff05a976c
z36fd3677c267c8edf800a6ce1bb20896cf3f5ebf7e648dda0d266a22c930806891420298740780
z4a16b3e63ff8bee103328ec3664f8f6dcbbe0ef4a7f1efccc15178f812e9a1ea99fbd8a7b11f47
zbd5adffebcd2880c3a0309fc9f01bcf35776005697c06d6098c8ea9d68f8d3f65c36d9a2c60356
za39d73280260f8146f361668e984716bda9aab5332b1792836561d52413fa01d229bbafe96ca2f
zee2c1521c9c6ad26eedf9c4883790c16300ad409adac4d524d0df8cadf1d0dcb44be3d4cdc442f
ze438a1b7b9fe36252758a167fa0efd11ee1f45e889d48a4749b65965796811cd832453bae8e6cb
z9b9d5a018ac7a0fe65b9faf6cc30c8e37ef9523e283aef7154d5baa8fbb5aaf2becb9be3c1e8e6
z7143b1eda40ebfe7996b127ba737c26698e799c33a814f77a8a51d5f051c708062fb556b016a3d
zc1b74b9de9d75a7fc07c4fb6154b29755a6da93f1a9085361f5010d0a3e79f376513cd9d048aa0
z816180b0b5c5f0127f44949b34a2800bd272e7718c155453ed2dbdedee808d1f452c4402bf1c3c
zabbdfaae7bd736fb62fbd04dc9365dd965d0458f55e25aff3dfcaaa1c659da98c14edbf273f8ef
z8c549675f665350c828e09b6cca9c396ff313ebd37d9c8e00a15d87413a6fb1ba9cc56d51616dc
z94967a7ceb0532a55dc5858402bde686c30e27e76dacb7e13abad1d8ea4ab62aaad6c1a7d18ce3
zaf963a0641c1bd0b278330196ac8cf1f162ccc521a65626e0ffbb25d505831bef2f3e0eb7dfc94
z6854690fdc271a7519ee326b7a3bd75f2ef7e10e7f83adc5082de6252850ecf67c7e8c2bb11d4c
z6d02ea164e704035207f6f1b5d0275254bc6de36bed7a059b1d3c719842d0dcab9a232ffacae37
zc0c80cdba420380c267d7852ec870bb6faf01ddcebebc4af9637e7e8ce6983baeb4b870a6732f9
z959e98315b24339387e1f2be09b52bebd81247b1b9b651461c6d260266b972a3256d10234e6a41
z4306363b46a66ca646d893cfa1315dfe1667790fc295a1d8073fade605b3da7676588042917e48
zcce5765c2f322f566bff77d99821128e065a3e956d8f5b3ce7b9267c34db1755ad3f359bf8bb54
z7171e86feac2e0625af6e6efa2ec8d8c264cdc5b2b6147a2a3e8ed2159cad25828cee2f705c02f
zba6d13fbcc65ee1e40499a97d1b92a668c1c632091fde03a25044fb0d257d548c4df1812f10a6b
zff42def4dfde32be9eac4e13009912b67d541d5d83635ffe8a74d632dbd75918f1de759ef415be
za6d1406092ed3a85e3324d5359da8c733868c5375182459f4d07fa229e9fdde69bd3b11d02ec11
z493041154954ffdbe7b55144b271e2b6240363b8c3e4e2911bd7d92ce8c58fa70f89e0f1a356bb
z2e6136247195f00816a30883e634b905ff69b94a182e38b16aaad3f4855cfa2d54d94da71bc26b
z9217bee161094d7756475d07ec39a8b9973b369df66562ab530f401d116dc217305d6c974342dd
zb932315a824a30020754c1c9d2d5954b659aac5537f245765d0e94b246342c8d2608d4f86a2fd1
zf9a71949bb45f2b671dac488ad70c56b0da7a08ce14af4665eef81ab92c708f789e700c72c3e58
z6bc9a7c25e5ff30480058ac128cdc4033f6c719ac6e3b6742e4d3ea63ed8fc97f6723237506c1d
z2760dda820176815798098bb1bd66d6029d2835a4e100134b4858d5729011d57448e8696af5146
zee77660a0870ec7f228f20bf705692d676f8d78e307cb98d3ef3f4b34f2b627fa48d95e2366204
z209943eb9fe56ceee113ca5e3a1429816e7ce9f764f98c320067d75142d7aff02862c42211da81
z3a58b85e689aa2cb7d16cf1bbf73838fd57d21acbae43224053940c6f0214338fe74a6c052fc3e
z4bd104b8bbfdcbd979c1cf82c320b6d8196c9d9ae143d46f80af909ab23a6abbb743848b854180
z8d0c40b0a34983c70ab3ed8880ed2be0c43b1b924fc0cace04e990cb4b632d85fb2678f98ba384
zf201c80690315c643929e5b4c6807571219df078107aa161db1aa8207683d025cadd275ab3df85
z69f41b85543064474da6410f7df881f2e7402128010d6d5dfb78bfefef6670b7a036218941fc38
z7893cf2bdda78017c354f92b01fdfa16063b8780d99f198613512c4a8567a8c46be4540f1c9cf9
zb5535f1b0182a2f85cfcf3416229854d485eca85519c2712f495f828f4f6c5c763e932579be495
zad8d42cb2693ff18b08ceb3b414693bf8e4ddac96d26f0367290c53d667880dbf2d027c91897fd
z69725f52feac5de99574ca88ff374764665b862fdca68b2a09f5b59002c003d58948ae3acbc1ac
zb5e2029278d6b7ff92e91bd59d32c788b626dfcbfe1e92f93f468cdde21b2d53add82885272ed8
z877fd70961f69ff936b26fcaf13750778c1640de07f24ede0066ee9dc01ea7f56e9c1f25bd966a
zdcc50e0266517359110646b02992c71f14cbc3b1c9127424863e8c08d5a1df12cb617288637cde
z2ac3dd924870fb0de29501e50854e248c494cc3e8c77775b5113f23d73c6211577cc07119edfd3
zee7c88574622e77081669e97bc704e8b5ef03379e75f2413facdc095a110c87c8d959e78d7570b
z28226fd88e040187f402974d03f7ff3532faa17e7b8677121f24849209a428a922fd096223bfaf
zc269ffaa7e1839e1c0025d4dd402e7da6f32bf0ebb53e2ffcfc840f601d0bab25773206acfbbe9
z91c307e06b73a6a880f20103fb8fe1a781e54f68ac151387052253d0f86ccb2885029bef5cbe45
z4fce717005e93c2b19f5bf65dac8635f04d364637ef0afcde8981704cfc690a4161b621e0ceb03
z2d92728117f86ff28fd329124daf5c3364f55269b6ad1a1e503de812da2635616a3cc5e237e046
za2a66f94577106552a861cb01f9f5bce23c50b3844400b029410ec84a0a5ad46b5b082baf87c2e
z8b0f81b2a9078b42a18ab0d310936142cec54b67054b3e99f042ce2f72efab41cc9ae75672e043
z30a7dc5292935ba4b7c196139ba4c3e569a49b6f5f0835896f0ba524f538ec049e0fabf268a54b
z8be7caa906458b1c7af145689554191f318c72a213bf5788ba029a595273bd0f81a8021c7a7930
z4baf1e633cd4c086d31dda2c1900ebf4b0a0624cc87a5ff53d5704575aa95ffb94d7391fb5d5c3
zc0c0f51b5846caa746c93ded4ec2e29a6e5c8d6fade3e7a857437d81dbd41715063bcfa2b1bb72
z03ef75edb847bab6986db6e0ac519b946f9356a346eed18856390d84b7d0da2cc48b59cef8d126
z05f9db3ab5d602f44d0918048457b663504d7205052fe2f20e1f5cf6ab7d67b41aaf2395420083
z903dd3431db26a1ac032044551a946bb6974ec78d6e8ceecff79aa10c4ec6254a50503e59f0286
z5c9597785a2b63e2c56b10cc7884ff4cc71465a7a8e5380c2c7b62ae75752086237f06af1b91f0
z3a68b16d6ce0345579dd00568c8624b84f1df9ff7a75824db50abb4612b6128adf16624a0f0124
z4d588c90570315287aed7ea6524b2326745dda436e0588ed33b7c2b322af9c74694b5a30505269
z27985f2f35193b61465b8a8610be4461fd77e96b81384242286e500eb1963e82924666e9a4596f
z4ae0f3e9571159cc7cd2f18a8114593573f0bf0f231690dd722966200446e57139167dcf667774
z253735552f8934966bec0069741002d5dc206e84175fa50461fa3fb2bfca3756179b30161f7ec2
zb236b0e746945b1c4238988ebe9719c9e3ca6a6b38c29d4157acd72aac83c1c286e8ace4f50b41
z935def56ca3a566492baf6beee8691eabba934025bd75ee90b150c60aa3876c48931c98037d56c
z983b7e1aecc3bdc91209657c28d6e0945f355c7a3284655b86f5219bff9d694a7697d4e21ea139
z1aefe876cfe739e2523c3301e573a59c9ba911eb10baac3157b367973b95403b7ae94cbf1d9df3
z381b1afd6d0290f4a4b4d35e2cf6e23327d5f29bb1d0fdeb0a4f5ce05132371d8eebaff002c33c
z17426db25d056af960b05339bfd261cfa4ce8d041180d27a120bf0ca3c6bf06e02f00cb3e891a6
z965f3d7e32269b55dd254d818041056edd77fcb447f6f5254e96a5c652a25b84db0259659276f5
z781d1ccce257a2068fdb53b5e740dfc5414939bb77c04f350fa70aa9aebafb800d822d0f440548
zcea99413bdac4f88716fc26d2eef3808d9284be63666a14b27817ffecaf8420cf664f4e31043a5
zd9bd58698ac8284b7a10c0a8511d4888894ddf20ee1c6f076a0216c8bee9e42469e10565960c51
zf062d2920aa1fa811c5a7f882fe2ca8aa6fcad8d6a8ee52c9b56cddab77e7404ed3d232fe8dfd1
z4f98616f6747517bfbaa83c781ee332bfc9614ff75070a48e5c5da56ff6f75e259d7f35fde41fe
z713392a9cb672203f575b20978968639f240d494c00456a2abd59083e29e971f2709f83f6fdcfb
z5158a2b73106568c787cf39bf116704d6611b6abc8066e1be39d6f753ac7e0c3534e1a0beb522d
z5ebec7129f4ea88f3f2a2c0c98deadfa41676449b5663d07de8e0eb30bea92fa399fa7bf3cc607
z25f4ee09d5037f09a62eaf3ad39788fe9003d26d38faa7a97c378fcad64da83bb62a79d6d35cb3
zed50d87b45463003f66a250d3dd7c07755c0da56f44cea9edde98819481bf223a2c14731efb2f0
z1007c99edad9f69dd5865a1a788ba2b4473e77db2a23eff580d2c56c9ac026646441a79d897152
zefd6617eb618061e08ca98f16216e45fc6d2068e1e7634e96c4e17b6867af6523f598f805e7812
z7e635657e9df85d29f2848e359fe0a446494aa429331358520852343fa828e758390c12795f752
z85d7780467ad9a3caa9e61b263f1390002b95314dd2e91e227acd402b73f50b2b71a66c9dc3952
zb95a24ad9e13a79b6b888b30e1870a027abc72a42638761e1edc73833962cf206eaa821c0c0afb
zb51119ffde01bb4462e53de2cbdd4367533fec1540c76bb6e31d3773b5943fc998a75414304152
z40d3797ab4b2a336cb35adaca0d3d60a04a0a7c2721d83b849aac4e73bac464c0741b3aff99d47
zc9d8155c2b488f975efdbfd274efd6095c9655ab7d2f8b552c68c125ef030f8beaae050f6a5a89
zb4582d29e4ea5b4ac26a5ea8f340693835bb12411b4d8f3d02388f47b2219cc728423cfb5348b9
zfa2288607d4669e1b43206a9418a67f9618f66168e987d67d7be0e94ed92e7ed5a9465eae811aa
zcdfb5e4c6d1968f07979f592d8087dc82e9a6467146c71406cf815372ffa713049e09cf724284c
zfe5d067989c06ad1572845594cd1b4e953abdda424306f30f3e93c89495ee1c8a4e6c36db33016
z18b9b4630dde308d1c1848a73158ce5e66fd60fc538f0239d0901834ce79123f7aa80da161c580
z99895a4294ff69ae0630c3f0ac89d77bbb09e49f5f31fae06687706023a996ae03f4abd04b04a9
z6e9ad904e1796383af8d25fb1385540e210a9caa646044c25365698bb2f685376b7323031ec62f
z8730ca5f638ed046f1b5d5499fdf9802445d2afef31154c22f9e447135a5dd7ed9a0cf4eea9619
z433888f0134e5cfb55b2c5c4fa3372fd671f70c8b460a2edb1ac57bfe6d41ef6ad41a7c3bc3ee1
z5082f71c9972a664443d37bcca43ea693e38f0414c8d761a183630e99f4d347d13a723a3210c32
zdc82c0d97cacc30bf1842640f25e3703c24e365be2b08519c3eb295d8be029268052f72e17d249
z8af91d8e1a87166c75d2138bf4d79e10ecc6d8c6cd1a77f280b0ea3306f911d33918598cad1db0
z30c840bd261d8fd1f4983daad330dbcc4c598b7a34788e1956b8c620d7785e0d2746913878de67
z06b762f33d7d055fb1a78405573a76dd7a4a3ba6add007734fd4303eb4506081ee3b339d2fb9d4
zda1ff7e3639456f5c724f6ddb81c58237c8e41284c1e7cae9a14d3064e5d1857ac9b53fcfe57ff
ze15cfedaa39d6148214729aafe17c8e318aba9061b5c02e878172cdbfbc89785bbdb815febbbea
z3ed9f01ec7064e43b26a2cc1a19f6b773fc419f1ba8708cfea6b7e868e8a8af6f72dc3bc24f7fc
za57a75a4a7124df3b4c887316a6dd158f91c125e94cdc6840267575bdd9e0f290a1bef0a984586
z985944c6ef715fcedea1672a1a878e846870eb2945dc49954344398206a440d0939c68d80a9b00
zf3b844bfbfa20e6a9eb9d2277c6047bada036ce6988d48fb570341e8638729ca71da94a5e30a8a
z3e9f99204028eaaeac605625faf7b831a63edc0ec1f58fbaecf60a0da93df1d2abb8971ba9b78e
z53ab30cb228e16c8e40c3f0241efaeaf146bb37c90a5773c698808d9167c4d8241d36ee793c1fa
z2235ac11658638c36a69a66751ce2e09a31d2d5471b68763513ef9f6fa9b4696facb17146b6e82
z5fa9cae9b1706212058c6c703af586f7ebba329729a71856b6b0adf0dc700117cf28c71f08bdc9
z191620d11f2c1676a8ae66f8511347086460f1f2117754051460e40fd8924f201b0c6636023033
zf08eb7e5f6cad7aad8ac89e6e383d06644a16a0dfdd82f832f717ea741aedf38bc7b6fa0bdbe35
z6aad39fbee86e637f5d103248dba101d8b05314f811159ec32db5c1b7b7f40e47006768a5b43e0
zb895a74f7b0fc958fbe61dcc4bb2d28a48e468ed6eee7c9839108153921cf90497a17a5c55c0b9
zda1c9326460d5031ef9fad6938b7f3c6839e134632ec0e93733da594cec57147d164563748efc3
z9015ca2546568d891d12d56af3dce4cb8a7819dc21a10a08b4b63a609f096c63b86ea30c764d0a
z5893f4f0f580108888c5e5348982418b9b71826823ce8c649cc0cf080b46333538b76362c6c96f
z1691d9c1f5e8550133a4f91faf47f7ae27bd8000ef1e95b56ab7ba09cbb6faa3dfe6a2b21b49a8
z05fd4f953955c6af47cc1b336e6552bff50b23ec2ea030537822c7901c2bde245e001efe9d7d5f
z480de4e873e9f782390c4b5f73e5e0e53fc6adac0d068e39e541ed7ba04f1bd618ed5c93d1528f
zc77d9af20a733277439d138fb4cfe022409f365f30905871dfd5fa8832fac7d2fa799173040dc7
ze2a1f0b387ca69a11bb85fa6d6bdb5c98b84735038db14619402a7e54c3e9d9f54c5e10e736dea
z1fa706db37841fb31811ccf395e00f3345707dc944d0a8a59f60b0159a831dfd74d614f0ab3f02
zc3955d7a98da6562277664aaaebc672c14bd014ac0a3980aad8aa7ab1298dc9aa790c33da4cf4d
zddf1d0e2e84f7c9803290cd399ff8b18e2b203092985413ccd86cf4fabe8b24e3332280f2dbfd0
zde64cdb1a3821bf9dcebcf39ee94003456788597855e4d5396572134d450b6561bbcaa0b2a9707
z4854b7e61a6a71fa40220da6d264bc48915980547d3020231952ce906e7c6fe974a2b0502a1674
zcb8c8f6b5b1f67b4adc79e51b5c774595f3fa66801e653db734a63b0742ce589296a9ab92aa466
za6042c37635466e415e48c884c217f0b073fa78d1a49ea0b5738da48baa2f1a0c4f4f9cf857105
z246b61ded6db32abf63fe23c2e4b4bda62a1371bd43edab33a2ef7ddc343009aaf2b199a636303
z6ceef9ed65c1c3c9b91243c9a3139f954d046b1d2dab1039f9367f5acf1feae272f91b1ba602dd
z0195370de6080ac7916deaae2ebc25080fb38b6743d0c90386ddfa1e839ea6f9cb0da87bf7794a
z93c2d17a0f21d615ed7417fb9a1918e427ce4339916b95fd136529c4202e68bafb82406b93bb12
z647c808246086517e30075918dc05b3244c722120cc0486949c88f940a08a2143dd7f4f9c666e4
z3457dc375f2257c6ef3a24e88814a17535207146d615858dc8a78fc90dc6e3dfad71ee418b4583
zc09817fe022f2bc7e7d4431d48f18405b84ca50e3edb535b64434ee5ac0adab30a0eb8ae6742f1
zbc946312dee0a8854c7167c0bd237467695507fff2647a54239c2b304c59c72356e447baa75f74
zac8de681212508f52ac39db790f4313f0fc1ab37a17c217b811f9a477d3dfecac312a89e0f0e5f
z344b37a04120b8fc7076f3a703adfdf45c09824f109653b6e4d1babc5964f7889bf9ad8aeb28bc
ze7a6d43ca14c393271f064792c23a7090df1921a68d5296e07bfcab9f304631ff8eafea726ea94
zeab316f8dc6243fc6ac95b20c73ee23834612de8fa574a5de7c7b07f7f11e2e70d39ecd4d17778
z948d0e9e8ac639a4c624da85b9e7d355089dd03c6559255ada7805b9cc2840b41aa762d35021c6
z6623fb7d5f0f70b1c2c15c83da90d172338e860050700073a90d397bcb0e89eccf1d579cd4b34a
z8837dec707c568175bfd3cb05b13e684fc9d164e5812d5abbcd48504defe9439e43f8d66bbb13f
z087c719bc56bd6dad8dae534a7e432937a29d0e51d5125a8b86de3cf4a6dae1d3e5f2aad80da82
z89ee2c4b90bada9e489d72b0da0bb4cd21090f3bb4e69e9a2502522501809c9015f21fa09b70dd
z90fe6f2e588e8b83f4050328ce466363903af2f07fba3e6c14f94c51b5c275e0216a2fb2e816e4
z99e23d1b4634fd127c4d90cfc01454f8efa5e512a7feac7afd5a70ef5eeb4fbf242d5e8f066681
z4ee285bc254c642d4d24f64588c2d31ad5bcc0ce2fbf1308ca67777a9adfcc3be3e3eaba32406a
z621930399e5debc6ecdf85fe85726596c5b06f0fc2a632368a3e4e36aa2dfa5be8c7f0697d252e
z4f9d3ce800581380a16ee73488127ed3e120f685d215bd1fac554eaa5ec458547820681cbb1fa1
z0d0982bba6d156e8b7095bbe0281bb26b81112d718c943813a722d6053801dedfe8898304641bf
z9d274690c4ff69ed13918415a98de99d87758248c00ac5f5d23f6504555cfa5d5d420810c4362b
z972a8f1bb00d1acc9a271c51cc21a1d809f3d2da319db42334843f1c66e38f9b6721af55d24824
z85d313ac0f93fd5b664fbed0d5bc9cf356ef42fe4120217c58267dcb5dc9f943392ea0dd0b04c6
zae4ebf609b6d51f401f79337f1f9a2fc58b550c6e158b41c3a6e7597bd7023d7abde87dd294150
ze193ed4de4d46156aee709b6b4548150e6934b84dcb6297ef55d6fef67588d1f023b55da0bbea3
zf22ccc0d0880f9d3ffdf40c0d53ea67a8c44ac7c8adf5a13f464dbc9320f76d8c53c212565fe04
zc9552f68c062317d5bb443b33688bfe8a44eb4e9b16d7ed1c1647a344631eaa9787c1025275775
z237a1f03611981f3458ac7088e7e7d684f902133cb190e71fac8da12e73836f93869395de68de9
z607c76aa2226555b48788b95cb55270533801d6228abc662ffd1f66f5549b0aaf85b6f9f6f2964
z2c861a3ffadb8bc6b9a52ec2f0a235246c1658236147ea89cca11b9739b146b2b1fcd1d3a031b7
z15783ef63b8e9f98ea7d61c006b3f475e8b6faa99b6da6878526fefe2b56087a18c23cdadea621
zcddaa6571439646b6f3bcbe7f5f16fb768b1bf20737f9e7bf2f88b7b9b348eb97539125ffca031
z823c8564d7897748360fecf472a9188e8c62a59978a6c4b01657b2d75d8226f54d2381f7413e4c
z62e506aafbf158e52717b873ab8173d8b6d4542679da71a164e2aa2ac0afdb0a8c812809392750
z7d6e365dc928459db17ef9e2ebd5cf5d36f7750dd23614f7c2d1805b8d6ab4a6373b26027fda05
zeba7bb67ec1c78291b9860726814adb3d640b57abb8d6851b9e530e76c244535780d7fa5956027
zf952779ddcc1e40cee2367840ebc9d6d5bcf22dd56fdf04291fdd042cbe1b35c604196dc9a696f
ze1a6bb03f12740b05b02a96e0b64bcac39f1f69e28f2133d00b2624bd447db77cf52a295c4ebd7
ze2ac5d81b899345cb4a928ab6ae70ee9bad000460012ad9e37ced7cc081de3f25d682a808cdb29
zeac1bd3dd00db098bc54ab6c9c2216156237668017c1601b39b971d47b02b9a77de5fabed510f8
z52ab4ab3b1d247234cfc19d04bbb35ff16369ba902c6680e9a3adb27a8a8afb381b4ffa68d2060
z491a63d4d6cf938e6dea85236db9b94f36ea3dcd4163450dc4aa9220aa52d7b228bda25d303612
z68d011a19414d0080fd0346998e735b15d482a93ed22c5644b4091611536047588fc6df2a0e62a
ze9fb2152b98d60fe27cab87d1ff8524da59c3dda540fdf8249c5c5098c59c03dcdb10d27ca907b
z7ae2a7658e880355aa06dc9b5f9a3fdeb28e1194d157fc748e2889abb772e72580000f14ccde81
ze99d93f258c874af6c66fa9c4140d08f2fa1a3d24f62dd86bdceb8ccc2b8c78375d9d0a7fba542
zb244aa8e373f206469f6c62d7878b3f353ab54233623dced7e653a564f8a708277ded464f5c2ba
z23fcc8fe87175ab7a352105dd764f7f7a8f52f25e1c38f6995fdd660786704306cdb845dbc0e19
z06421121c8e33d47d321cfe5cb91991c3f502d411094bc26672020fd2bb31d4da73f7def48f36b
zf89f799e1b5eb9e161e7a8c4a51a4d54621d7ca9dc65747f2b97aa175cb7abc599779124bc8384
zd60eeb7f8f3466b4f8e211a8d761efffc970f5348bc7359756ee7dd742780651307ac48dedf177
zd9b02643f13be17ca90b1daf902dae0b07f04f95efdc28515506c90e67faee58eef7a40680031e
zb6b810c21f6586cbf3c0d23ed609be1c02112558f98bd19cd5dcc0bb27d51b6704b51fe111554d
z8523ed5f81c039eabb29d8bfc58e73a2a9c246138afdea7ad2fdb262d1f5a0fa831d5809e26307
zaa18cbd72e3637ba7a9c6e2a3fc4fde18d22f2bdc54c18b7fdb238e9b67ac3b43f32e629506462
z10770f5cbb12de82c411b958178a6c14c538c9ab3ca1ad4cbbad4e5320c35766fa713c75e06b54
ze6323d1773b59f4bc76d988da555e8ca0676acdd7499640dc19a030ca58b8f847b7bec3cf3cc5f
z8d9d8947771f859ba4af0e7935f82a12cc29b0cf560996d91ee3a070e22f930840734889be9282
z12adbed16bdbe433f067617cadbf571dc5adc0f92e2dfabde016eafd56461cfc436589f608d4f1
zd14ba31f0fd65a48a5ebd658975742453c117049905a324b5ab68755b2be8f50e030254c7670f0
z7356f203c7393ae09f4d1c36c43895b3e7be86659ce446247f3e569f5ee6f32f8e0295b93a40b7
zbfd3cb0a5c070d52aeaead00179fb54687044dc677efb95dc906da8a7c6a3421a63adbe6215cef
z245430cb92f87d3bce02644bee6fd14da3f146c3cfebb91ea087dd2a926707d3b033e30372b674
z7865b1206d213b0e2bcd0fc24d1c0f7273a16d490ac21d23b9b81dfcd8ab07771d92246b5756fd
z11de35cc63c745193b97dd19e27309cc323dabb8b7a2557f8c3e9027712bed51c4c29ab62ee33b
zd4d3e7c2779ff586e7b5e036291420308754eb44eadfcd87a48b52e7c462477d15b695c858721e
ze344b28fcf897340d9f1b6c10eb94dd741e4b7892eb065c5149d16c69c7ab35d6a295f4e1cbbd3
z81543384acf7f6633f3504b14184517910a094afb0d09f210d424a7823eb5e6beb6bdae07720e4
z55389ac9e212c0fded769b8d5244af58579677fab132ca79007ba62adce16af44b30243f96f52e
z4d68680e9022eb453d68b7219f04bc3de661f539b00b6bbf64c719fd0b0c84d060f04cbda0d80f
zb13500d4e9a7fee43446436cf8fba89d593cf839401483b5c48062be993a3af866c1fb13fec37e
zf0e2cb98aa02ff67c75b425911ca7eb514b2cdcb04c3036d0d6c95601d44a006d2e0e02848607e
z8d4d10b157c5a721ae4668b767579a0a9cc6aeadc4a00cb6369cb6a2d9e23e1062291594f5e3e1
z7f54736851383b2cdf03a369a5e069de3ff1502a4fc8ada38b89196becaac0f506dbf81ec70b24
z2533a485455b45140118254b4373adf4d3b5f24afc9cb08d239ac56731f759d06983c28867d1bf
zac6befdd3e55bb64e3fc155a98413702558983accbae52dfd275d742242f82475df5a53dcea9cd
zbd21ec2ba7fc9fc79408ed6744266a40417dd98e25bfedc6ab1c49fe7dcf4e45ca0280030b44c3
zc045056cf469a4f31f76bbb50cb8cc0d902cd07ad8f2dfc70b17438886b046490d4b36fb8b5670
za1dfb5f793c4388bf9bad90a6404c8b1c034b8dbc12b93a592b2d23d5c47507571525e2387bef1
z2899ec32511c7566f6fd353ed4db5e3e75c73a3cc99fd6570401683676d54c1fb714d40a71ff5b
z39cb23373359da1dc46411d2ef2d460163f92449c706d654c3ceb18cb460a43062932edb786cd1
zaca1c308f57442ae08d415ec2c022039bd7a5c301e879cd7636dfd4d8a1dca06b5686fa9ad3e7d
z031995a308454cf79647d840038904f67d72865115c7ef25aa65e34c0ac85cbcc10398e47cca90
z87b83ab817f88fe8b1acf348f39c23c06e3acdc1ffa29e3e9aa1d5b365bbaa082803818955e779
z4da27e38a8aacb9cba5aa1506590f6cffc54ae5dc45c172814b7f6ecc9ca0e28d32291d6e86609
za93ec685170bdacbafe73fa2e703ab9afe97457c0044234509d3a2495b17e875b0e4b9ce8e7768
zc90d0abf5ccfb636f71125a4ea9798c04dbe444ba29394e99c99b29237245374e06653275aeeef
z2876c9e8042e0319daf08d1990e3b97bd77e0f07df8f51b170e56d9b13c097197b2bd157c092bd
z77a6b40edb745d98e3e42282e6d257cb3cd20add7782a9010fe324d78467af9df4ab04f753f274
z6ff2af4f1771694caff290b54caa467cf84c81a76d07cc4dde7c2d757c10fcf16c2baf9cab3a67
z2a38ed38b2c86c2c47119caa5f371858bb6352b5d3d54bd16d5dbb5fb7ed32f3440043a3cbb3f6
z10d338000009266af8479c54af813431058032b8f35ce44fb40526997cabe7a1ae7e806455d73b
zc38aa51c293d442e93e029f0e689230e6cc1eca4320a3897ff71e92c3525b5369e8a651073aa57
z8bc19d5228f88d7e4b0006b3d38f43af57bff70fe9bf35e5c77c5cdc607314063737da6e835251
z087bfe4db6992aa3c1080c1af63ab4ce228e8b68c6198986c1e9bb0d522cacb9d7cce693e4c8b7
ze533d162aefd3a203da663f4b07ac2b1554da67267756b6de40162c50ceea4a7e53f0e970a1f63
z17d9462e3096b972698f8b8a1842bc6dff15b3bd5be46607fc52a7a9bf19d8c57f24f0659257cf
z655d25adbefd31b68e1a27c3b96db1b6af7c40c9f8bed0271de732031cedba6b19592462a77fda
z99d3e8d8653ccde80ba4d7c8c2ba34b41c27f0a656507b1a2307822b06fccf277da1b73ce9d2e6
z245b0d4a30da0910903611a5b4e014847e4dbc0f9c7f5f382ef4fb15957c79dfc809355c8a5a71
zcdb870fedfd00887cb6d8db55c76e8235b63341569ef5372226165f0b109c65c2e4adb33a6d16d
zea8b8436887b3d7a0e930a6c127371c4ff99c1122c55a3633e5992492a14e837e104bd859cfc50
z46d25280965f758adddbc23ff70160aeab478e910803ff12d2780ee76a33b3497685b12aa0ffc6
z1a19dde4bc130219da6be631514e56c3529b50c43670b6f60b88df4c96cde77b1cf187f363701c
z34b667178e088126aa71b42c1cf7d5d77a10927de32c3021395866821fca8a93a8433f547bbd49
zd06b0397d9d082aa8a8ad861a2564e814272f78ad461aa10d8f61b29e3223a6e068152d0c8ade7
zb9e805b331183a11581ddb19ce9d7bc3a67604806bc4b6249d59b77a40cdf308b813ba1f390efb
z18fd44ba16ff6ae4c27da2bfe9c447b1043815de247a84def4f2cb3f6ea36a4d3361297687f52c
ze0b3c9e0cc45aec40652c62941d17d4462151fabb9f82a1d101af8599cdbc08052cc73ea35c7e0
zc1e58025f331c4cffb3601edbe788a7b610bbb05b5799002640c30b040c4dd1117f8251383f50f
zacdfde19c9a2c46391b5231efe1a798e706a12591ff39fae27a1fe0efbe6999c2f85aa6f8fb03e
z184044294e05c2b9f2b1a5437a2255fc0685d8750f9def197c55be5c891bb2446f13dfc2a34d80
z57d399334de63404c2c8d42ad6cd837c6e13f91829d40a94e5677e5da01f4c886841e910c12271
z23cb16e49a5022db96dec0f7097f57d00033b9eeda579456773097ed741b54cf516b5a7a6e77d0
z718196eebcc5978073b3b188c142cc1b25d6ba2e7f3e5607aaecd5ccbc824d86941c0718548ba4
zc6b73b9126819e82551ed772a2d28013b68e9d6f6452c90b09322e4740aa68747f4af0e75d0c75
zaf8e43a5745b23d07933fec04d157b63e9fe96d93dd78ccc6bfd0bcc584b1b478526e84a004451
z2db4e9f21795a7fb32546cb82b187b9bacaa2b0bd574058d6176cf667fa516801280222ece87b1
z7fe55114b19032ead3cc75cdf5e87dcc05e16bc3796e510fba3221ee4949800e14caa1b7003778
z12cd4a9699c22d376ca2ba023302754ce6008d09c7b2e3b5f58de3698a4c92a7b265c290b65f0c
zc0264fc1aed3810655720cdc6950d77d60c96d3b0fb49e01d04d9971b3152b152466f7fe63a70d
z650dee57d7973582719d42d1067d0bd145e45d69352a117f4a0d24781f5fc98e0f57da89c0dc48
z182b041f34ed5dae200780ee1701d26aa65fadc7ed2168b4f3613ae970056919d9ed576eccdb48
za80f9546f69c8a3d3ff0578348ead5e0721cc555a51ae59a6708e1d57551b22f5ab36fc4cddfe9
z06d6d67ae1e5049a46cf688bc8b65b96f6f0b9dc5800d5adf79279fdcbdb15ef14c491847db98f
ze36558f67917079d853d0b6acdc954800dd719ce45bb0a82dc5e9f0d44b730f69013705c16fb07
zdde8dddf94dc20a828941b91d488e579256a00e6a525b0185b6fe159fd9ab10a775ae22db657ea
z216de7e3e2c8ea6b4b27f869ec2891c8b5fcb512a76f6bd8746d2c65f39d588ea15731e7c43cb7
zb52f5e5d4f2fc0abadf2ed0a9759d07c923cf2df764ec984edf14b27e4c3a272503782220c8ebd
z37da14cf3435e6d91afdebd89ca15386ec52bddbbd693e8f979d72089b26c647e9669a546de959
zf751c8abbde5fd34e6a08ffa2846caa1d2859c126ab851e358cafcf047716a5bfaf4dbf267a5bd
z4b0ee4e6ab873c8511dae12af04b34ca3f3894c1343b701768a826d9cade771e2dc894802aa984
z686857baa0f4a5eb9810e44a356f880642e9ded8efb9c7475b84b4f925bcf3ac8eb8bf499335ea
zbe985dc5ec6b5d599dd693c677b2f223585544b215d6d46e46e6aa14f4a44b3537714ee45c5b80
ze2a8b284b4ecbcdf20d88fd64f8cf7aefc3901cda9c25ce1e32aff2249e2b17283e5f61e63cdc5
z6884e6b6eae387039b1a073c146d18f423dffd8b053deff25d195c7cc543bef6ac9a1da02b52b0
z0543a6e518524e44bc93c631ea758b45679644cd27936e60785aa1443c6994362e84a3957bfa8e
z8282c02cf4cb537403bfaa46c88fd3ea798c67d8d25bc8415aec418b7467ec629a44f1ff76bdaf
zfaf35453ee4a0942ba436bf377ae454eaccef4e9173b8da991d966c1fdd495e63f0aa4e034eea1
z4637db2899122bb4388ec149eaf87b0ea24d348b7c77b5a0a84db3642264d87ecdab476d43b2a1
z7fba1e50a06c2d299e1ceea96c7609a885ad30361ad1c39b4cdcd4983aa18995cbd65d99b918e5
z5f835bd8cdeeba799d8c2755b9a1c6607fcee676af5240927b5ab2d55acf3c9d4c0b03ea2f416c
z88664a1ffc0aeb979f8a7e71066fb205521a6ea4082d7ec674fd802e5bfc9fa8230cc4962f6d2b
z50859874a8d90f525dc556df40f6c3d26946d3396c074068212e97bc8021cd1b3b6f69428851dc
z99a7faffcafdf8f8c2d5fe08daacc8bb6c2f9eb6eddf3851ac4985675bded530d0d107e0ff8376
z66ffb727cb3c9357aac979d0ac6ce3fe445547b5653a3cf8cf282bcaff4a52284f2f585c9d11be
z671172e61d1d508eb3471d9753f67f6f9bf1030896ba3e7f30b660521816eea2b03a4b3b2d4885
z43c1c76e461f0ffa9dcbad60d7c03b5846040b2a31034a27fb29c06d9e145440643d29141d6b52
z6e5c7439a1b93fb44f2c5fb91541d9c9fd2f83822c38942b1e25571ad83e97247b0a70ccb44f84
z73ce09000b57ee0d7196acab9c7a4d160bf33a73f29ede11473526921c3380d5ef4423efc2c6d0
zdbadb0c7d046d4b13a2f17bac8e039e743e05dcc245d40170df5383befa42b04ddf2adfe77217a
z82709aa9697da51fc1a24f3dc02fe945fb3dd1615558ab1c91942a923849d8f4e1613079aa5922
z2c6a6def657d1e174fc226fb3864d5e994b6139094270a9fb0ce3527399756f3c525747f610853
z71fa2eca217cf5126851b21c6bd9f6ad03ebbfbce6f6a94a0257c90d704f9b7f0b7fef026f288d
zdb3ba96a0a563ac7b415c8e8fe7153fa1a82896ecdc9c10321347dfbb4bc5dbbc33638db760dcc
z319701696041a5d50b29869eb8ab30991b25010aaed1d40528516178c56b494a2a757fa8f8ec7c
zc452a61e354f552a4e34fd8f7efcd589bbab77127090d63d49abcafa5bb0aa4800c2cfe29e8e50
z1ed767ecf0484e83a444685ed9b0cddd98292758206252e281517961aec324aa3a19de525f11e8
z716f0106233477e4efabe6b2e02740379088e729dd6e74f019c6c63e81cc8403306c692b42e617
z367dd4afa86e281af285a81649ca620d9bc6eb73d150e9f72549ebb6bd3f443cdf89dcf147edf5
z2eaf10642f03ff89a0f0d5918c954fc1ed43cf6e2129f0e091c98e6067c79a83fc1224c60677fd
z8ac0b4983cf1cba0315bd94a8bbf566b687d92f56f54914a500ab18d22c39a940e5109159df9e3
zc1f07213f7f3b7c0de4442c5580601fca6527b281ab66cd7fc2dfdf9bbaf9b7334317faad4d0f2
z87c6b8f643eb475a1af4f19a686ea2fac4f2d62a2c96a049fd2fcb6951f39249c6e9678326c28a
z6042a53360c19b34ad3cdc27b0ec5bc0914eb1e550b9c056a5748633975af92af3dc71ef2b4d7d
z6c2aa886cf4fe1ac343d8f8be8847ae932dad1d59335cbc9b06192b8211aa5247a59cbd60b43d5
zf2560ec2b8ed3efe84c30d488d55c451cf47dd2e96913a2952dbd50e942f3e39007fe2cdc6d430
za0c56e65ea287f4cd41ad9e223177475fcc110f87c84eecf22961adb9356af4292bd14d25cda1b
zfe8cd1f1807f427739ed5c8e5e902c7353f057604793df493a517e707ff712508e8d797ce10fe6
z2d894f9e81150fcb25b51b88ebb12e4eee6694f6137cc85687b8f978ff7167a91560b8aca54ac6
z4bc63d671eee8f5841a99faacc44a59a25859728bf4e45a46d7b9f1306d1532cc19bb476e31962
zcde3cd1223a2ce572bac1e2959076272c9e46ded7ca778557224ccfd1a9273a879f91ea5041870
z85b996f373e2602828c9ac3ec43d85a66ebc1cc095d7ca5ac28efb59b7db203d6cc8deade8df98
z370dc263c67b40702edf07d1716c0b2e5f7ec806372d3c3411f67e84da48a9986e0743774200c2
z6cc2b87fe09c0952a1e5838670fba0ad80d2eb64b83614dda7bb9d9a06d56f982a6c21a8524edf
z4ace40593ef770ec4a22a162bbf6c7b49f69915202561d393679c7885ba6cc14b122fd192edfe3
z32c3601e902a806442973cd166382e10211bc46c053ed72f25686118821f9c9aef38b42a0b8fdf
zec1ac84e8ed965e496d855830ee5e2fa4d2f0bc362e6c166592f385192f13ba8bd72e70704c636
z25cf209ddd826c3e859329546035deb09c5e59c33a675d3d4be875d013248872e8e9f68029cffa
zeca9045d1b89923e031a7a5d30ecca4f94a9483b43bc02d8605a3011cc8d35871743d71fe166f0
zcce5ba73efbe163a1f78b284c735094ad400698fdd36c8e195bd0ebd0c482de9dd4be69c129009
zba6e32474fcc3555c14ba51d2b9ac684875094e755d314923309ee7560231d657f817bb9f70142
z3aabfa483ed06a4da3782d441098dd06f416d2057fa0c25cd2d6f9d586cd0f86a89d5ec4b84c32
za00c788c425a03732437ef8834caa03d8605eb68ab777853f597d5b19ae776beda66b37c048ba2
z8dcf9dc6f0075146955bc464146588e067fce68e4ce85df71f61d959e546e4c37f8faba7ca9c55
zf1405fbef6bea6b2f4792cb73e22aae8b0147f976bbea92137df3a6a3c918b147aa672436098c6
za511f246bb9fc73bf085eb2987a9c42f9569a180de1a220c3a4579f51d66aded18eb5040e22d35
z11261c2b675710b0633b06d5a702e056fcc6bd965993863b9c982a09c74bd47b9e6991d830390a
z6e56054ea8a12740019cfe20d131da99e893e389b7031566faa9f7de7d9a1561e46715b647f0a0
z5171be93cafe4e485f1bfc8189a8a0267ccc55b315cc6e945a051e54c18cd6723353d187072e02
z13df3952e19a59df8ddc39f2b92024d18e3ef77db2b4a78fb33bdb06b0baa0a5b1f39535d707cc
z4ad78f74e7a1afe0dca076496a1c079c53e0e02ddea8fe7b3f29d56782afdc487d92b807eb688a
z2314667940bcbb1b1b55136cbdac1ee9b8f7bb7fb39cb92a2229f92c748218462797e1bf27edf7
z5870f08d51c16050e59f414af0d0c98244cc2b82342f92b8ab18e91736ac03246f2e3fe60ca5d3
z819a39c9b13902243790f412ff466bab3923e32900bc6a03fe20965629754641ab21d19fb48fe8
z5c207d663f20b7812dd9c9172680b9252f71fb4c125465a6e4e13e3bd8950f2b45699eae0d2251
zf82b021db899c8053e38e62777b6d77951876cdc843fce4fc79eb6afa480e90857a4a93f1e59bb
zcedee0093515311f65e58a3f571a469f0bdafbe15b25b0eb1bc055e74ce458ad77505953fadf66
za40b6cc0079d78faf057fcdf5fef37d6be587741b44ba6cb16a283e138de27d36e92bfadc74fca
z244c38f90c802508ce6eb65b68217761e34ec8211af498da732ccd840ac26c4247bf19eae30cf0
z2aecbdbfec5992e840f8c83cf857c230addab137d9b2912ee82d384252592619964e266cf8dbca
z90f4aac81b6b6b81607483b8c91cf4896596bcc2a6aa983277b5c646a3734d4e003190f4a7966b
z5028dcf7b2f6535e7d39ad5ceb923c5a1935eb414e66ec7a62b195bab6a64ed2aca25adc85b569
z443ad7a0708f9795ae66346f53cc63e1c7fffd3c9b85190896c6d53341b785cb65473aa5d30eb1
z4aa8d8263e382993aef2c63a15cb97f8b0e5db59443106502cadebe35132e995457c0065143c54
zddad5a5b93fc3b41586a24aca9a0787d0f966d148fc05c4fd5917e700e137e2d95c741c3051550
za0eb5815e7c4915551308173c1250cfe1c9c6934c3a874864c82a8e26c8604b06c29f6fc01af00
z351c1d674c092698194850b0411b6c45af3b75f2cabec788cd0528a25bf6f825b9e1a6311ab864
z73b7339e14bc74e819fc6a913d89100c3007440c6f2aa7af5e4d286e670cb7e964708e3b44b2e7
zbe85aa68cda57a328a493783b912cbe4644d204ba1cca5e7ba13d7a2205392e9388ea4911218b3
zf2cf3944a4db6210157689469dad102bc6928e42f47cf5d4633cc34546a5a6fb84540c32c6a76b
z092883aca5300c4406653c6667fe9b95aa65db4502f81c4dcbee81da1efc4521e88c34ac159f7b
z745a135669c7e52cab192a403e1b783c0d58ba2851be3d370ed5f9da1593c99649f11c19d6c22d
zddfcfcca3c10865da967b39dc123c5212ffc482673b79efd7951286102a2fd9a6ede7423829f10
ze88c8fad07a82b4fa97e07fea6f27e45121a3f41bb1529576e400fbd8e3e7f54ab85909250b842
zcf2dc50233ebcbafd44064aa2fd34c7e0a055120beade7f201d2c758d8fa0e471cbef41afcebd1
z1d1ccf11c1dd29b3bb54ef9b37730129634018cfd77245e5053656da7d80f2c98f4577b04bdc8e
z6f3a988870ba566011c8d29561bbb807337ebea542fa1e4f60cd78f88b5f57d086aabc44ec099d
zb88b723ca6fc84b2b28fc04ca0ccd06e7d88df4cf3e3c69ebf135aaa849ab3a83254cf44a58fa8
z202ec60dfa95125124dbb0ce5f01fde4289714b8a07ef6b7424252702232d3b15af1abdff15b3d
zbd6b9b332b4c41e3d3f2269b06a3961df2cc9dc5825dc62179b9f0a740471db6cd19020b65bf43
zef49412c16eefb277683642bc73f2b89ba1f20bcac840abe5372ab06c8cdf8df698c1bc1067ac7
z3567416c9870546abbdb9d1e4f43c36105b06404535a13aba08596516c8fe9dc71317db483dff1
z2c1dfefcf3da23efcbac9056019076aedaf51705edd30b226b9a08bbb2f454774f47bbcd9a95eb
z26a0b9c56bee82163cc8425e23e06df1959bd81089497b196638698bbb5aafd103d2ea75752d44
zec6096425881b67ebd4ec46b2be2d9c7185d81f22057fc079472109d1b077c57bcb365182727d0
z87d1881133d26b5fd1d945ef5337891672e1a1d94019d8e0c85b34d6521937b199709d312b15c6
z171d9671b7d31854573f62e5f7b25ca446c4c560f782cb9c8d3cae5432dab5c30ee8d05a128262
zd6996e8bbd9c24d182444484dbe33c120fbdf01b5c3cd1c9e331555f4cf79c6aaa5ac3b42d3eba
zdbeeddd2f7961d6431d5fba8a45d51ffbfd16b515e911875c0b67ae94a65bea0f57e48262fad4a
zb96b5311126ff7d4aa65366dbc31549328d2098ec1aa08eefb5020b3599ae402b9fa1d8a86bfdc
z2cc158bfe2e530575e4c0e2070ce0f9a7134b77906cea5e9f79fbc7055e14eda17e554d2d46a96
z0c9e0e3ae0e0ff42db3c3d28f6a5b237b2bdb452c522be52d698c7b46fce1b6b58d5adeb2da184
z6deb23b954df3b9fa53e0d0f57179b2247953e2a4eade2afd387a347dd0021bccb46c6c9ec0e8d
zc43d66fce21c5a99b5fc9a674be4645a2b7c5831d7fa63a84bfedadea5aaf62cd802e1ef2ad5c0
z7e8643ce062fae5757a12361b63c1aa5dc58c84be8d9f8becf4ce2b9859134ffa3bcdee1d3827c
z2aec93aec9a73eaaab87f8513d03c2ed70be6d8cc0bc255a6a8165bcd3d8080dff226df8a6dcbb
zfdd867a29e803ac0e82e513a9dc859db31417f4ef89717b8aa08e4c0fc58c7d75b15404e5709ad
z55a40b84406fae0ddd6218ec65dc8f9d0210d229ef8ca55ac84c5a510d35e11d004abfc5cc26d9
z8ab1cb2415c71c201d847a29d193fd1a91a8cf8af3af0d123fa8fce61166f70073ce4ac8449d07
zb29b9c17a635c01985660b03883e9f205b2eab9734bea8f96ed912574139e63608c26f2930a128
z47707637c2ab0adbe115c9a59d6c49c3b13315e8b6ec5a77cf909297123133db19264373f7ba2d
z82bfdb879ac03e21405fff2603cc7409c6d2678f0ca80c119e47673df6ea70921ed7df1ee2d924
z60d9c43722103f59575d7f3fe0d2eff6e846f1cb3c341d01247405c9b475924a91447301a0b5a9
z21193806cd82204e8e034b05869772fc15b222a2c63263a0cee0d50cebf3db001cfbbfe6f6633e
z4cf745faa6d235a2dd8e092890fe00f82846fcb83a37472e029dd8c8f37ba9dee1f00b48a5670d
z06a74131c0a1a314ccfb86527e5bd48741792148f2455de91d7552f8570e61b76c01d68bc5b5f9
z7acfbccad81aed562d649b2466135d2c8255d8c2a3dc93abee9165f9e994a41921c5d108de5461
z93554132c26a1a9d5796e61f762ec49a38649854b67e77003dceeb03abc2974d67d6b5deeca886
zd0a3f0da75cb4805d72e6c20d92560d40642a369422b9451d4c4022445138c80e8560452d49c64
z2c094d406183531a959949a8052e46d6ce7cb1368e8bed3b80431223e8a18e2d62cd260ff571bd
ze3b4ede27b060fc25995eec801bac5ccf486bfa7c7529e32585fbafe4a8cbed79e70c94a6b1f4e
z8c2cfe8d7cf06a37fa3369c061d8cb35139bd58d74a1e0c3841dd7eddc9d0bf8bbd20638aa517e
zba51a27cbd4cd689e1b62654d8a664f749438cf78a9e6b56a838399bd36c05a4c69176e99e1a8a
zd69ae27891f3a0124ce850e07acc01a9b695cc4ee658f6943710d4b7e47f2df560a1c1664764c6
z6ab45bf02361604dfc5c24ec1f00a5fdd4a478fda52d413a101697dbdb61f8013d1e7fd28a1232
z9123b3564cd927198eb61f3d97b3514e1d9e99779f01f7452ab3e29886e8b5d482ca551a735fbe
zbea1499949f56a64008476a3b73a20f0b07bc27f9d09e9eda6b49e5b7f83d3d399567864460bfe
z8daf0337e31a951eab94746af5c2273334da50dc60ec79b8d684bb03b912f82df17db7e08587ee
z59e8753b249bdfa03d78a72c26dc548ceaa21b06296d13856185728003ba2e77ae825d526e760d
z9e37bb163dcf92eadb60b5a84ccdc6ec1ff8604d88c3bedf7fe5c68b99c94f059757fa1d04e73f
z157d24e65bb3fa419deb65791510f4b74ce309bf8d96e1a3168c3698ddf98c161d01a2bf2984a6
z85cf4beb2e69c787eac51b2468fe672ba236af9fb7e57b0273a46c4ceef4b0ee6e8b1529a91935
za88e2a3b9b1e709734e67d2b50131415b781e4b3c17f761f3f544cf3e3a771ff0c25665dc947b7
z058bd8c46b1df188bb8acb547e66a6e4614b66d146a195084befac5eb330ecf56d5eac9de1accf
zca8b1e0a299ab010c8aae037b6af2fc0846629db4583e58c9bb2df75a6f8b4587566662081ab84
z186e0068c720076d01d611f76e2f37bfed4b7c9a843c56a51fbd4ec83c15f02c960e62df6f67b7
zaa48a8b8a1875a96ba06ee997620118572ce63a3eb341bb70c3a7bfe4006da01fbc2a383640992
zaec5da3f55260ac14e66de0cb57b56ef5a153b0f4c00bfa06a29ddbe264bce47fb9d61e3fa08e9
z2b5c8884d5fbb8d09d2b0d812be756413a7a11e28a1720a7225d8ec0fb7218053bbba1b12523ca
z32f165c5ce6939511eacf8b1b9bda2140e0eb8e8aa05e2d509a666d72d4244ba3cfca06a6a1b23
zd2d3682fe55fdc13d2523cb3493c5456300a403f02958657faf8f6a002e930e2da11a51bcd3812
zf2fc5c128707b17b94fb5d70f933048de47adad64b2720caacb28ac5de5ff98c9ecc79aa1a7afd
z6ece013449611fb90cbf77ec74788459d8b94ee358d0c80d08e387da4be2e925992ea526adb700
zffc66f07fdbfea97afe3276b32e34f293a86b5fcf4e88e47d866d7372d3a7e7967990c7edbe16e
zdeb521b9a611292b867717beecb968bc6b2ac858273cc26acbb4b789726dc690b1579ce8a6f19e
z1b3e9db345f78a197e2de59e96d01f9665b8abfdef297420267a4b0ffaa09442d4d272dfc870ef
z3b6be2159756b482a17565695277a9731b4bccc922eec639bcbbab9f58c64b49eeae64531608a9
z400db8ba7d11e47e02e3e98b33347aeed15671709384b9566be4c2a2132632ad15a5d6e5aacf8a
z0651695918ee06d33870988f073ae5ad2e8c6ee5d856876637f2b3369177ff78f6c9b36d507e51
z59f7fd245750855ccee3dc01f25229635f5e9390bf2841b34d39408922121c6b837bf4272492d4
zcc008b43ae1c7870f431bc28655e572c0b07a47fb513e6845ca9cdc772cb442a1585ccc8d6ea1f
z22898bb736ae54123d45d388263ceb7d6742e40c8a487927cbe76d35187267df3cc78aeb308f54
z3c4ba33fa795282cc9562bcf669a4870bb06740183b77fb8db44e9e717c99b93702205d5b341d9
z30989bb9d7244e72a2889c14094816a6b5334ae971173d945d24a93139591dc30f2cf649196b05
z815450aff25d40ab37e3b8905d7b6f7762d62892a6c18568ee25d54ac880ca3ca1659e7fe8060f
zea041181c702d78690bc03d0621445595ff488cd123fa797cdd792d8de45f5814d48e3504148b0
zfdef24b3387c2350b90f4389f32aec23be0741b06a5fcf880297aa255e260377c550ce577af08c
zcb8c705575cc9956531b708c6889eed6f02173e68207639e79dcbeecbffe856847912dca99d984
z61963ba0aa734b9dc173a8bd71b563f521c6cb8e0c9473b22bb2393c7c46be04e25e11cd20a8a7
zd000033f625e7ce97b9cceafb02eeaaea418f517e5345de2541c02461e66a17482d1ad6651c61b
z89374942827346890d98936e5fd06c65ed7c5088861d01b82a4d00f0b37966c1bc9a9c8435a4e1
z58a4ebbd52a2975c7769c650b67c21cab9dffc60bb00a8c721df5365d60ef2e5611900cc08cb86
z45f1d2f7dab550d5eba7c8d2121ddb041f2165da4f999d77f7344ab38b566f19ed2c3f244fc908
zfd1fd7056ea6e8ad51088b66090efc744dd8a9084809ffca9f550589cf0bab78a0d3d5ff4082ad
za286e7e4c503cc17fa296e1774f744611fcc0d3eb6735993853afe6a1232e9dcf36284b9a9add5
z0977a0b44a977a705a4c0adf59cbf5b28d225a28bc2b604a3ad043a0bd6e14be5e187abbb1cdbb
z0290f55d9d6853529b4639a0c48d7a1dd786eb995aeb08ac42ad18f7b451b8f164f398ae5f5c0b
z747a4c1dd690d1dafba16c65a7ec7f9ced2053f030c6bc749472d757a8669cffce68406137c39c
zc6e424d9452048148be8bf9c3e399ef40f45745ed05af50bc0b192b7864178226b4a01ab4ef5d7
zc7974a966ef44daf5d41024cee7dc3067911392a32ef6c8a62442c420a1d08cef5f15d525cfdac
z231022da126e8b92f13b6dbfb9c973b8205c86154f59c9e90642b76452e4dfef3e07c0f63592b5
z87145711a5445978037bd09bde59337af4de1762284fae278126c25c4af9d6a2a385634fe964a1
zd5407694b2c5e11443eb5795117f34619895fc81c009b481a0014f421029d51b24ffe5dc308994
z6e56d35144cfff4ab55a002f5513bbc8d05a345a9b76bfdec901f0fa8e9c7faa6d901da97c3e11
ze27f8a206f73ae3bd95266b77205518d59d724f6da0fa3869af16fbd8d4af9512eccbc00500961
zb866a08b584c3f0ba22c6923f4b092c8bc3ca2d0aee5fa2666f86cef6b9c177c2bc45d39d489a1
z1d34e92c475d37e623ebaf22a6332aecf4f2324e539852ca9114fb628e236842e131ee3b46d7f0
zd11ef8e7508921ecb90c892e9503ff67db9888d46c006a8cb8c3fd8a9a761ad0b4e2efb70785da
z8a3659209d8d05f40836f8ec6039c57db9ca57f7220bb32deb8338e859f3bdf9c23876e0d7d81e
z273b819da5c2cb852daf5895c0c2a4a5e7dd92a5f9e7920d646b9d1a50f37b32c5ae4b7eabcc17
z7a733bee2f7de056f0da639a1b5983da10df744ac4521896083ee1a58507288716e884a0e37dd8
z5bdc044439acaedddca359f9a9bc093841b5e9d7bd516c714e750310e9a22d18641d9fd3c9b49b
z66e48b25b78258703ea932cca85f6f6e479334416f05a582053027be7c44ab32b53578b34453c9
z3444cbcec8d3f49c653e24774cf5dd7a9f3888e8241cf06b722f2a467d74728cf2d7ec6d8315bd
zf6df7c0bfd9bc9afa1a8a9d6681b96c9d3215ec5edce515eebf4c503d2ae53eb7e6ea831a47e71
z064fc7978a772953bd0fe6a199dcb7df39bf3b2a8ab9708f3d51b03e9bc2ab232859add94f4bc4
ze22a49bcf4abfb00354012aa6bffd4f5bccee947a28933e963b3a67257843316f3c4de6c14908f
z4e8943a11ba8d05389e890f84cae5fab7f094b5bbd335f8eed61130500e78e8d9aaac936299c92
ze4b30fa588634297c08cb8be663f652fdfde07fc4f95448346e83e5e61b822f0491953f27df9cc
z9ab4a6ed64ef78fb4f9b51ac6d84a1d0d4ae24218d89a2c406c52d70f84d8c900e722cc4f7cb15
zeebe90b5f941a5e92c4d10b967bca68839a4d21a7742140d5b743fd322ea4bdaf3d521057afcd1
z841e36870201eca9ff6d3830296154ae5a21f19d3a4c6091ae28df901f88afd4c86b1b617d2ffb
z8daedfadbb891c209fc1f15bffadd4f6bb9338854a65f7c3504258b556a0252e56c078e58c5a15
z41c2d306e9cabcd4a894d83e3dccfac1a2e03da36135440a5026ffbe21a4872410aa9be3187968
z5dfbfb491d1f4f088866901da6a11bbeac614165f5cbe65c6b9eb8521166e3ce3af3c46f3fbe24
z21bb45e3ef1e3611b5d9091e2b515cbc060aebc609df61217d99db009f88496a8fdddff2eec101
z8c6b9921cd9d4b7ece38da3f9f8f9fb89abb662cc64f5e5d56d25ba4ecf0d48993d2583a8c50d9
z2a17ff8d4269797561feefe6cf9ee6a685a46776000916a7e046507041d22df8d2a99e65ff7fd2
z9b0f7f18ea7692ba2ab5706d2fa028014a131d41d20be0b349748408d0d8675773fd31b45e6b3b
z867b4c0e9642b0600a16dacaba26ab488027663393123f75aeb730ad89bd2dd2c5fa65af24e55c
z250c3ad15b00830cdf3af80e0a6485ef19c398bdddd29d9c8a718df752daa066f5c505ad20169e
zce1bf8ea8492318106473d7b942e48752737981d5ce40314719a51ece5e170316e79a414ac2a1c
z4811fbfaeaa40fac97b05dac19500725296be4f3836313de53e68095f48ee4253ba4c5f33e9d16
zf430c804d7096b9811f4ec4a21e2515c175037cc1750287e30e4cd4f74103d0c7600cd5903304b
z9f57d059b45b657f9392c6f1382ef592665fdba6dbcb1b1b8a73e73a87f2c5f6eb89782a64ffd3
zfc5548dd0201139584bacd86060bddfc2d8d68f6d40084cc9bb227d9f10be8ddd3884ceb642077
z1a8f9e61a0a4c65ee3fef98c3655c0c5461a5cbc4cd5f2cd7b1e218d4a71e961505172b8f2b931
zaa8952ad376de681b76913b5f4d9d3ff41bcacec2ffb80213e22cb82cc482d2d076b01abb34cb6
zca943ee78e54f8147b293a3c0bee5d8f23cdc1a06d4c49d95ec815ea8e673a32a3f1e68a0ae515
z7ce16bf3fd51f5705833c7a0f39752d2f052bd44139ff6a2f558372fe6ae653f08a1c786a02987
z83ad0320ea59e66e83f3ec6bde1c2d692e27214566e98c3af3a3bdcfb51d83bdf2d41c6d9f90c8
z9fe21891ce35acb51678c04c4f775703972ddd2ca7049ffa3daf17e69eaa4cac7bc5b05c7135a5
zdcd816eeb24416a51618c8492840793b6e8bb1ce5d672c6d05879f593dcd53e74f32941c787944
z9e829c39ef29d457c44c6fec78dbbed545cd1b5ff886ee50a591b8694c7b353836fecb23cd6903
z508e301054dff08a758b54bafc55a34b177cb3714abc86c7d1eb4553a47798bf91b1b00274bb6b
za79a09cb3b82919e268e631296296b0d2afdd2124320c4b26cdc7f653565b2308166ba1f5216f0
z31f059cddcfcbbb718b5aaf3a6c301aad82e740c53a727ab20abcd69a8544f3db8d973d561e1d8
z5586ab3735bab73b19f0d7ebb3fe0946e4766bdaca1dd50ea5381139df97ecd21b7ff8c2a30ded
z98466b6c62212ca09dadd1e960498e3b67209c1c25bb9a6cb561908e09e23f3925aac244394c6a
z60f5597bc307ef5423c9393ada37d6f19cb278e57cb41fd3db0f9f430322ccd34ff444e4b7a35b
zad7312d37c3d7faf054f457169e39959d0c582b0aa84353220cec977bc1218b961e0256a94c9fb
ze2a1025854b8ad76d19f38675c8688e0329850e107784ff0fe6b41d1d475ea4cff6412a7d72cb1
z59c0f60dfe2d7bb2e7154532561919445f280a8c4a276f24ae066556230082f87c0ee9a8c66cf1
zf4098504aaca73b8a2b9326a6e7809e0a954250e024ce5ddc62ee6ddadc5c26c14f223b29fbf1e
z1f017203c66daf89e0e50fd66615b29bcbacdc8b3c10b456f8ecfa91be3a2e4bcd3839d5061047
zab0717c8db5c576666cc2a73d972563b5b80a08499743580ffd95e23b00a54e8aa7ee2c6489966
z77c94592cf72aa1e1d35dc7afbf21b1e253e0cb15cfd91d31da726c1960ce567aca43d6b87856a
z2f9a4d6d01d18dde4d0e1e61f56fe8063ccb298d1d52f91df040d53f5639c0c065b644d6dd639c
z06b65300411cc3ff8b0a399455e2237569b68ed8355e994c646ee9c4d242f63d01f58433e7cec5
zc9a4334ffa08b9ecd741bdea31cf910c08ecd8f4ef791dbbc935df745947fdad22143ec1e465ea
zff4772604b75d5906673a0d176720bdf2face604820ac0b95e2ac1522de7a5fbd9a272159c436b
zaf981a49f2c991c0ce70838f82d77a5eb2ea13b899d6e38b60b45bf99615ff2e0e897cef0269b6
z9ed3d193ba3c1b40b5db8807436b64c32c809582114297b6967bb01a9aac2a8fec00faedbbc9a0
zeb50607bfea6de3fca4a1acde1e2615a1837c7117e1176fe0555e3c22fccecb8ca62923dc1dfc4
z08f4e0318a021f2a07705c971127d1ba2e4dd756581e8a8c9aad1d6d12eaf1570e1f477a0fa5c3
z48ac285b8bc78e7afa715cc3a13a78b609290354e909ce78a20c2a54c3985dd7865324735d7685
zd8670d594d0108363f215d9f03d7ee55591a8f6512de99c8e3457bc977fd1d6c33b62a39557ca0
zeb7c272479da0f1444be284f0a26b1daa6719b344a836bf34ba445dff09a6975d7993918ab2731
z05da5f305d38a28c3a76f3da913aa907a093f411c390b3a4a07ae57ae91e2d3e79304bd067383d
z93c7e0f77f931dd0c0124022d7b0cb6d42a47f74b0f367d9e64322f20cdba0079f455393ab0122
zda47b7a4beb54b120fd520e9b605c03c7ca4c2571647ab53bd90c32b3a6e2f2a61677b89877689
z062605b2098b066c94854e2da2a3e843d5c976acf87aeef9285b345be773e116669194b696d7ce
z7c255f8c72844f7b52562aeec67164e9db770fa63c61a253a61bb410005fdcafa63b04f7f84157
z082697bae4a7d470099640139a2c2f9f7db105c080ea2ed55576d9ab31ca731e878e8ef48b2ee9
z9f4c5445385b757229d09c79f1e621ff28e5d3e1f778fc7f0e93c2ff724d7e3a86acbe9bff2e50
z6380150bbdc298c183e91f35cc5078ec8d4c96e416e943d9a1921e91a9336aa6f3e5a61922ad8e
z74b21f6b9c37b50f20d32a6e57581172027e0c3f1ba88f2088e1c9c6c56f1c56867a0a855d8058
z24d8da653e6f9597b9f566febde65dec0cac7ffecbfc83615d7713d4644661f815865145da3262
zf9273bf1fe8f7dc3d90141a192dc8798a94a797749bd3d9680d3293a80c9fd1544aeceb6d71b93
z00c6290a1b3e5a65b4ddaa43ae7ad4097a93479f3b1fd40dc50275ce56198642bea3940ff0c386
z21c13711d36570b10eaaa19c9f096433bc5a66c63e40d03dcd89784b97998457d01ef3f882cf4a
z27e433fc72e672dcabe04f8872b02b546a6ccb7e95ac1cfc518c4ddb41b2e496c0c38cf9846dc6
zfe4368c4c299a309e1dd4962d7516639866c87a72a13bf63f9f9ed67dab65c44b738fe596d34f8
z6b1702dc24922e87eacec2b8c2d7f5bd03d63550b4ac3012907223cd6e3d489c703554fc0e68c7
zad50da9e875ac2ed79aebf45d74a3847287f530a9b0b3f89290fab3150d6bb968e221af23ae750
z3ded96ccfe8184e3abcd438d05f7d085b8c6371965ce485b42cf5a35ebd05ac9a94f9a33222d89
z98ca5f885caf665e1d6ca6206e70113e4e2a28f88147c1ab20335abefbb867d2d049a9f258508f
za530336711974702172083911ffb3aae954bf58f34250c77d89067f83fb291a608336c37ec5267
z73116b518555a1a736d5fb420c99bf26cd05cb4b9dbce62e87946dffaebbcbc99b08ca0c8dcf4d
z8f2ac92e5205f75028277c788883efe4a41c9361d37648a224cf5f5e231456b86b519b3d633ae6
z8a83e8963a5874c492f88bc9429228c2f974bbf27986a2b68b4fb68a7c8e54766eb543f76fce66
za8d45620ea5562584196690e2c97a89dd957673847fc9ba58e57da4acff7e81a12540d9d6e1b40
z36551d5a9eb694dc09d97981d938e92c0d867537305e4125cee34eab8a2de9b526a1678dcfd842
z303580835eceb5a5344a882ba8d28080ebb945ba1d4678d6b741efb6181ea796686c1c94a1f474
z1f07ce674f64e49c2f7bf3754219ce0bd8a2bcda94692282317ece1d189054ce3cf6b91b285e0c
z2c0bc01b72f597ea45d25c508111666bb952003cfc0ec51d0afcdb704c0cab0d113c9e52cfb0d3
z7f4a992e916e187a3821d3a6b4b6457051415034937a0531ae53fec191b19e45cec9a2c2d16bd9
ze64ca45ab519723239b45df6c328d0f51479d433f6a8905f65133fa2abaa23c03b3432e26ce3a6
z05f8c068202db0978b9036d16397f0dac55fa53030cdfec29f36cf4dd90a96ea09a1f9fb803f8f
z337c97ae99b09f0f839e01c753c27a176a4702b8b95ad34cb3b31d02150101747cc0335ad03031
z1929981186e846ffccda5551118c4c5e2dbd853afb669179fa4d8123afe85e6404386f17ddc4b4
z12ccfe6a8e38bc2639dd3b90aef36fb0b4602120957182672991873fb2fc6c40798659b2f84f20
z01a129a830cb6836795ac439f4446251447ca64783c649ef8aa3a5c3a8a32eca9a0dd37e0a26d0
zb4b78e15050ff94ff169b68ad9b7ed3066c7ccbb69eef1a796f3540577385331e55b7335812e9f
z9934796049e976e111e97f710281a00083dfa23b2a1827d95b89170cb07b61f68c5828216dfbbb
z097f4047771b3872caf3a5f3053bc85b685319e358b43605b6bad060f5d782f68161f6f3e8abe8
zf31cf62c0aafd5fa76e0f99311d93b1061970c58e65bfe1c96007d282db2b3777dfb8e7fc3c5b3
z5e5028fc41044b98a35d1d9382c6fde8501693f374d7e80726a6edfc8369f2fd5d57161b9cfa93
z3fd16fe32130116fbae6acd0cb0e36a092d858203b3a54982bc034301097c6d6ba511a2db9669f
z11e67e018b7f82e206f57f0fecccae8cf8291233406355979456c07ec332655f5e92a3c70d3450
zf5736a22965c553b1e8864c1cbbcfc9386946c3454324d6a37ce501401dc5407c531d177099ad4
z5a60c86024a8873d01a389083a2cee59d84a6d72ef1c324165306d7b2b97981c5f9e2177f19017
zfbfcd977f5007eda9c1973cff9c0f2aee919d7939c8c27d46316af440a3c538d88f9f7febba72e
z73fb95a36dfb2c2c1a65aed0eeb891a94b40683564e746ade5419b24883e89113d667d5f282468
z7dcea6d99eb4eac29301252ddbcbf09a825f15171cd1417958a752db611dcec8870f604ff164cf
z7e795c1a184a376685858eeb59c740bc25fb8d13a3eb353ba305d29ee1ec8188c4d6cd31e01133
z17f6f63a2c7c4d7348daa6f12e7a6dfed91ff7b6ead1f237007202eca5015968941fdf872a0339
ze8aa60c0c2e5f84c8ee4f1475c1ef03942f7473d7d9b395b7193b74beecda6442856774382ed6f
z28bfbf8397efcfa2ccfed370a88ef23129c86e846a302a741aba5f04193364d34c876492dc6201
zccb9b7c75c7b4b339c05be6d0b7453f54f6404f20638a4109bd95c4e975b34199d521fc3d099c4
z0a0852d74979796230ef0cc73ea018a9069b7fe99adc20495c527a6b3d8ef540298ddf9dbe6b2f
z51298adb47beae27e0cb45b59bb2054620a8f010c5d28fb488a8145b57748ff816a8a4330b0015
z30a68d7e40e44977418cb6ab480dee1814e0634a8d1917d16799cb069a837e6301b71ae00dd68a
z454c6718367741bd162f0dd5084d81b3e6ca964fc0770cb314bb76a923d14ab2deeb09b0b8b0b2
zdef97f4e618fe89bb587fb2643da1ed53685c5c3ee4fd745954332e3668f5ff573202299f882e2
z1c4152a7e129133d961709a1e6fce7694a559f8a53605dc6c890e06d7c27753c666cca689af096
zc932e45f184b1581fe40f43e617c0ec3a87dfb3dc7544c046726f0885336bc20ae79476cbdfc4a
z9f12073fe041373a5e45bedd067ecf9fa5ce5f2527da79922d38eeba5b89f8e2b95b21c440cee7
z67a2b24e925808a8075caaf1404948d165801a117249661b51d1951dc4a2d3163bd26151189a15
z4c1ea8220c18d97352925acdf517da760e821ebed41072ea03768962fdc1b5c8a30d6f18ccfeff
z0b0f2374213d4b570653f8ed973f0af76295cfd9f198adf4682c5c87fa69f9d19ded9025598eab
zde086f7722913237227ea73b0ab7a455ee130a8487251e46fbe2c0548ee31d4127ad5ee0e0d503
zf3c6308242fe32741f57cedede8b17d012ea2daf0e8e39848a11a78dbcaaf7597a1d37d43e7778
za137b4ee261b3af74223bb13c7cc3192206bd6e219f306043bdb0e2aeba7e6af186b9c1c49f737
z44b2933e1c907ea3036608b5a6f025265fccb640654410bd1068d0eca0697af4104289b7ece2c9
z17a28bba836051be1e18a1ecb9d14399e0f7fea3314d5e9ccc1eb0a71e9e8c8b013b0ec74bedee
zbb1ae7bd56644aa9018a29de5bedca854a7590856c6fa576d9603e3e905e9e9b27fa38ded375b0
zff0dd05eb2edee77339dfcb94c3ac4d34f2f9c664cfe33b985736078fb59b7a809205272a2ecd4
z0500737aba510cd1a5a898fe52dfc7d30f243d6e6af1a3bf29c213667c3872372a5adfb071db58
z673c30ea934672add3b7964b10388ed9f0528ba202b71f016018976535aec004b25340d7d6c7a6
z527e16b6a1dc2c5ac8e46c368304a0e1301105db74060f0936c5da7b45e4b57efd123648db44c3
zf19acab0aca9609b19d48c20a194a58bc7ef4da079e06c8c607d2f7de4098f34b7ac84cfb98991
z8a37075833775355be510d24d312bda29d3c7f5e25ae7abe105cab6201a83fe049abccb004cbd4
z4ed830c7b293abc8a5d19c815968c131478af92961e7e10117e5a5d5ceff4aebea691c7da49a54
z1e4c3e561e245073fdce05970c6c2b12cd50bc8f8e15c8df2e6ee8cd7e25c3f690789b31e1fd45
z53fb17dd70fc475afcf8b5d93ead8bc20cbb152ce961df1302b8698fb7b98e0e1fad10c53309e0
zcd0b56b988f16c2aaa4f306d751a1d79b24d2a78598e48294d8c5189e5f3350c9fe3aa76ded0e9
z528992663584daf13bd342307cbe69afbbf6a057f94e2d96c8c9ac74541e9d854ee3d4bcf24cec
z162b235c101032d6195713cca037fcafba6827b5ff14798ec75980d51f7a64019495dcca387f07
za8e8b384787962e788ebd3846ccfecbe40a2801a0498d980f354e67abd409c7822eaadecce2612
za49cca8e8097d66c3a91ec964d5fdb9d81fa48efd64e6a7aa5e28024e779f5fe92ba9117e48d04
z1cde876d3d612bb5e0cc37478132d04e80ee63d60adf83a16c7a983b704e6ebdb1a226198e41c6
z1514c3632ef48a2602204a0627925870db548d9b47a3996535e3b11bc717337f601e6f44d7656a
zf7118907e19a37976808f51f6436ce1022bc563d8405b49e476a7240187b73fe1798fe75c3d192
zd18ce1930d9c3c0d7d4df9150a91c05f80308e67082c8cd93dba20c0ed32c1d9964db0a6d019b0
z3898149b37864d70c2a56e5ee8392cda2bb79349f80225e8b8b9ebd1173ea30a95399038b8963c
z602ca5804d43e5f1ac96364b5a18f584b8da14d88cc2b72a2d6324e22f60a5fb38d3f809e86ede
z4533162dbb69334fdeb32f8ea579c18067bdfdea654a696844792268c1c7ee981e85e7ffde29b8
ze5d97ea1b5039188408605ce1e8c782cde1ebea18385e3a40f36c28d75e0aac1ba817e5ef88763
z04b6f6c2a3a37d370cd7cf85dcc53142393dd620e7059de70c5440224cbb64f7b18e827ff1be17
za4a8516d780b2bc2eafb87b7205b01769d3bd892aefa6f43227a31ab46b83efa6044bd6a650fc8
z882061e1123fdb579bdb88fb56b7498aa2748c2dbd5da7e43f8b44b1cc8bf15d48c7936c56e2a8
z743c1c976eee414c63efb9261e94bdd15c9508af9e246547db69d17ef1c9e60b9a125696e30a11
zf19e2a72401c96756ba411ab632e8049ecfc87318f14d2d13ebb32ab8367729be4eeacc4072f5f
z6a9719656598180acf6efc9ed4572d0c782bcaac70228af4b494c5c087207f9fb449642d5b34a2
z32c7bec44dd8a625f6d74f914e885950d748584eb5a9eab1f101179f8416be3893ba0ea81dd03d
z6890a932ea95fb4a2efb30bbf5144c8c2c9fd8bc253487ea3f2d24dfa431c7512e7e12de3b6c1c
zb83fb43e5350bb9a5366a76e83d971d3413c797eed798a93da8b4912c5e6196b392939739e908d
z79fefe6effa5b0ea7ff90e7131d04c3a4b3de497f0bdfcd8894a562852ae4f238c0c03327818b4
zf2150106af88673a9d7b2f30f4e92718ef02b830e82753b97412b8ec840480f701a70d8bb710e2
z6337e0d4b59329ee5f079130b0e41632299b7b2adf43fd72eedbe5f4d2307ddb8a762f549b6c06
z41b08e0c74d72454d217a8e8a68db39659c3c1106a6b20b2e2dbb3169981da90fed86494e95eeb
z9c780583f2bfb7372db86041fc38c7d8c40d53ce808d9dbe1ae5ee7424a7dcdf147af8fd7be1e8
z377abb551c22e1074f659d907546ff9795fcc30d2d352fa3363148a7f0389d8bda2d2406c42b20
z24f11720591a163ca033d54458348b44b71add77f66c7fd9439b50d9c1d358fb7fe7a68461f53d
z62a87dc316fa659861d5bc4048c7c83484b5b51741067a9eb601127bcb3c1507ad8c7eef4340fe
ze4423a9f3f3a7b02c5fa97029286e0c7a97b99e35df1e3257146151348d5fde6785dae840ac32e
z05ab45849ce7c34478af3c4ee2998cb21642123029db35484ce45c524848f67b14c28ff7756bd7
zb42fafadc297832142057e535f8d0ad5641236aef52ecfeae398e27e7685ee62e3bcfea659173b
z11763806bdc8a8dd87e27485dd38de40075cbf6e4055e8a4de9951374d9348c0e60e2e618e44d3
z22195155c583975d152b2cce6a1182ef557286c974bc67cd746226b183c571fa26d79c587f3193
za8515b21f279352125e4e45ed20f786ce6e70cd859b567e043d115597164254c24b15d4d57c834
z3b2a45651848d3ef6cecb78189ae9f651a93b9cdf8402167bd8bf161019097aa037beeb2710836
za8fee2695a1d68708a96eec2025fe039d5c1920fb513272730cd5c5363e594657501132f088503
z54937a35b3ebade7721978734a1ade4ef7c291f62dc2842038dce1620048859e6514cba321e8fd
zcbe53d858f532128a704f72cc484741201b67ae644cde1f7e443bcefd94d3b702685060da96787
z3039437a51d4940eff3c29028adbf15e75a2ca1dafadcb24dcc13eef9e650ba2dccb21e5e0b3a0
z0ed869dcf77ec1779d234b7c789849a3428cd5384a49766c64d37775a5829f375364523d046df3
zfdec696056e37f7286d1e2440710afea9c51af2aac9cd6904e5b860eb6e4ba47187558608e6088
z6541246d42d6657abc3255732fd7cb4b4e75f93ffa5a465173ca8d1a4172200b520cc0100f9e5c
z6d5a6e7ff82e778c0485b9794b530cd79b2113aa6f567b5bc3ce4a977463b6aef4b73c0b48ae34
z6c175c95090fa3da7cd2acb0d922e9b366c59e26bc14bf521ff8186fb339cf8457c658f26e10d4
z72a9aac25c3c7a4490dab82bab02080e60b2f0f97d33f08b71106aa7553b34c3ef23c97f92b144
z48b0ef35aacc0824a4cc4bccca806a48206efd19d182b4d6be3f5494a7e7d8f723c0a0e8edeeea
z00ed231e982d1f201bbcd44a26f8adbb6071f3d86a27bd3d7f89cdd53d46430074b72981e7c628
zac3fc392360ae9d58b6e677bf6ffa9fcfdecfa563c5aed4584a314df572e37a5c7b9bbf0c56dc2
z796a5613b1e0215d3f92a7f607252892aec100d48433f82580bef249b1ee4d9a67302929437409
z849f9a34b63ba2f0404788e109e04efa1a9022d5cd2da4aeda2592965e5f2ae8fa1706fb769e43
z14bb1b34d18ad1ad98ccef371201e7acc96ee24230c863aab4979583d9a9624c896222adeb09e2
z3f696420277fb5553db425bb4343ed6f08737171e9f81b9ef6e8fa7cd470ce8e61c7dc31b92633
z49c72e602c3feabffda3f864026fb669f68493b30e7c877ad1cd0ce45b3768c083deb5f5c8627c
zbf7086c0f9c400370b0bca0bb88eb1e2387ba4782bacb300699634733dd5ed94740464f1c8c712
zccb938994bc935d5d829020b4189de4bc2a4cadff2a23505765622f89fbecf4f5fe4aae1b66625
ze9b7cd83bf71f8be473f5573b1b8966c99d579f0df9214db9dbb1a0229b816ccd3e4150f569814
z1c854442e4b4b37ae414a7407e7862890388678251863d4a6a1026ea15e10fa843f862b73ce0dd
zbecba7b27f64c8095fd22201648570c2f1141dfde8eee5bd909353c272462bdb80ad838366c00c
zc31e32683b6dc7960ffbca93a4d5d7bd98e56d9d589fda4984b3b174b414a23b4cdaf2b593bf82
zd00e77eff6d93788d890613cb73fc8f96bc83c244acba2f8a5dca7e74b3c8651484c0b2e3b339e
zff0b20c46d7ca05602d1b5e2c7e0e12a40394829a8b991eddd3d2d119b7d1fdf7989e802e23966
z51b518f88694b654b242ad5c01b580945a6b84e17c8391072bf910ae59b442e3ee654a7541c7dc
z92fcf9c739a2012f7a7c2064e0d817f5cd267738538d56a5dcc3c13c05d5deafeb1b477e9c5190
z2b7488a5411d87598259a215f76d150ae0c3d0bd677ea8a3922a3b36f065e53cacccb7085b6ceb
z8c3951ff13964322e646d431e020203700173363a70f152149bb31e14643e145e9e970fae575e6
z2b12da8caef2b28fe059d43be15d4d58d6c4af2ea2fe046d8b6756495ab635685aa46d497449d6
z75516a061ba6da8fc436888a863e6a05fdea4d40f9134fe9c046ad39e1d1ecac405afec5e39896
zde84f932aac4a989b477b7ddb8a17325920618608905044be0edccd2c48ac5f5a20accff8227f4
z54c5b8ff4f30b8a2905fd7455af0af08368f61e5e98774e2b4925b035e335d284c6753b9a06d84
z4eeed4184be726f223ec50897bf0c04bb476eb4474b7f991bc97f4546491007cf96efebce4a1c2
z7ca5af7ed8d1b0ee2d6479471604398ad5a63cb3dd515d858da362151b1f5cf5fa3f3db78ef3b6
z8cb45ebfd9eb805288e34b8f5f60469edb49278c803999572c320beb027060843b5b320842f7ea
z0357fe877878258ecf30b013616dfdf52b336912968f1a0735234e4a7466deba346196aa150936
z2686c8c25db99b01ec89384b1d9a2fa3c70a412e3af189499441bad4d363d47eeb9ee75f185421
z5f28f37cfb2d65a6cab331716e5ed9d4491dbfdf1264e7f695abc072513717590421b88fe608a7
zf5f72f81edb8d05b8844ce09b7c5b42765a759a49d876107e84ba1a819ddfd26f300b4d8bf1e08
z66283d67bf3cd196ffb754f3d649e3ac03abca39ec4f0f6c1d005ea9cf5cdb8f0e32e6698875bc
z10e4a8da25a28b23842291c0f2aac1318d61e82c602dec8527ced33708ffce20055c03a185dd69
zdf0212d375cc752d65910e65770b7b9fcc1b5765326bc944a19736215854ed00ca79591bf0e08e
z7749f72217f00f50f15894b15b68fdbc56958dd597ae540c625020b1d29101c4463cbdacc29452
zbc2bfbd69453634c5176329ffedf6858c676683bb7ad4bea7bde4e219c7b16992c33cd0ef04942
zd188a609e1811411402bf694f413f24f324ef1df400985bbed0a933c3af69729c6f731a6e21bec
zf734b21bf917093378d6095576195936a0e7d591cf19e62cfff01ca8fe653c1128c150f6835ad7
z4aae72a91243bda7b75925101065f41a4ab262110d54063ff264d359208f0991f1cc81e85c0467
z343c8541aa38ca06317ac56dcf54af6715226f00331cfc4c7d647ac03f382fe57b3952461a14f6
zf24d0c620da6b007aa684aeca347891e5a9da34828c5074a35d86e66135d0c64ff61dc0ec488ff
z96d4bf11cc173b5668f3181c230cecc900e021f84e0cb21a26ae76b2941fc40eca9a87ad90742e
z6ac63eb74fef7fd1abb2578ab4e1a406881cb53529dfdce1a37c3a5ced7f2790478d02ccd5a648
z549f98347f4ae057635349ae15049a6a629a51b646ae511cad0671bb480a90bcfd3e79d7516b57
z125399d9b2883d9702c669ee4f0264b4e7e21edc5d9e54dcc66ac393aed1003e43cd7b8c4776be
zb4a8b57185b1ed5e2277ab29a160bad72374de79efbc8349ffe7ebfd3c0707c3968249ab620e22
z89168bb48f4e77a86c94d96bd96115f8f6ab6c33dea9c442ce27200d842cac7ae94090ef34cd31
z96694405de7b40685a80042058f40bdc29d7e871a580ca9daebcc4ddab1c5e5f7589e1fd1bc66e
z18e20e61ae7c7ccf297174b8d96ae1d50b9c3f5d30d7b8e9f8797e9c5a3cd7013d2ffffd788f8b
zf310b9f373aaf7d81bed12ba1eb4b5a242cf2f4aea58c529085835ce25eadb07fe52f9bafda4d0
zfebc8472331677de20351e5b62e55c9406c83eefe636804ec8e6d7fee2f0b1e9447ef104c533e7
z5e9314165fe8627b7823b5b0ac368b543fffe64984958636b6ef61fc2a1c3ed08652e2bb964eac
zd4987be1e40dbcaa8299d3068db2ec1c0216ef2379be4e86ef066261e89d36778f572b2a74c3f9
z8caf06fe547247193b3956dd1bbcdd7ec901f97f54a703f5345317c1678bf57883d1d47be4e745
z161b20f8066d9b493f3fc3bed59f127a94ef02fcaa1d4642530ecbcb05b1028ff47cf48a440593
zd6b63af117fee2aa19644e1e8baddc6e936140e2236e24b5ce0fa71e551064ab5130d6ecacb763
z8ccc780b2e38dfdbd940337733cadc6978eb4db3537e798ab499d937e914cf11764f10d9cd395b
zef4f740302eec4f806d1f6553780654594c6edbc46c06483802e390679ff04e8e8927687640f32
zc66391037431f31e981690372287c3ebba50ab753f7702ee8c66ef7b2e803efd9e2c9ba64a294f
ze2c323fea6950dbebc795d7e38dc1c0c10aed0db6e4312c1748a44aa45a517d820770a7eca1ffd
z360ceb2db97730ca3ccb8e7508223b83dd5eec602140f71422f12ed57ecd38e8f6e97e7d793f42
z2b5b85de6ff7c32f11908e83b7665e20b8b5e1758cddbcb2b3f7c7ce0fdf9a8e35d0c574b7121d
zf41ec07a9f9ea522ab58115554dc064d12118606c4642052284e71b9e9b42165b8cf0791417267
z94427fcc1f5fd09546deb28ca538bdce985e3ca8063cd145212d6f50862e133fd7c9eca2458567
zfb61d8e712c252286915b97515bc21c7f19bbd208f2031a6290f323ef036b00d269ea4c400fe94
zef6906c5164abbb3aeeba07a90e856b3cb197a694c1c754e7ae07305d36d5e3dde09d7a80bf8f6
z5db96ff62b823b25a478d6141f50651ff3abfb6ccdf23a185dd027fa2821156c74667e5919323c
zc8e2a4a31f6ffc559177f9f3c639480ab874475eb57023c3cfc783c17050c991b0ff9507dac017
z893cf9a6a8dfa9f1d0215570a2de21089bc5575cb79ca9359cc63c03b546fcee592a0f35dc9235
zc24e7c689b8d6cdb54f098944e60aa3423621557f809e44546182dc8c21d94bc4af0611dcb4cee
ze72ba84ade6522af996fe55ba85ef70f39f456f0dc1a10aacfed46b27a03664a672f561b5a62cd
z32017a88b8901cffd115cf7ad19fe321af4df7feabd8d84e1b5492e6810ffaf576770107e055e9
zea7002f9ce7888e2382eee05b0c14cedbdb75618cf63fde7f5ff246adf013fb5c1d1ce207ebb71
zf1f7cfea7e4d7ada80c112ac9e38f727193fdf32863388b81afcf47d6be24cb0576363cd782b38
z56be0191f21348782ebf86cf68a1855f8f056d27ede458ae4392d03f33e00aa1a888ea7d80903a
z02cb0993a6886184eb5c34e2f74acd6c5858a3e092b4a4c1948c0f9faf8e2f7a72d1770d1a0acb
zf57bc10b6bc5e3f3c8199b876e78c599532d5cac59866cd37d08d49a191115dcce92345aed63c7
z00e3d6d7c8ba8997face3e1c0ca193899fe09b481a33b5e18343b5b064fe542f79c47a4aa116a0
zbf6d85b8cc64bafca8419944e0d8462903399358ce0114d119ce3bb4dce6d41a885fe76f63b38a
z8990487c40dd0ca6ba7781278535994b8f51df33f8f9b1f27512e3f4590f55b4816ebda1ab597f
z61984803d32aa9ea9c03789b1dfee3f0e92482bf1cb2b0f579838a19b67dc6dacaa41c7f7f9868
zdf6ce28155c85a6649e3155b785819cbb51ec871f56e73f780a81d7f26161ed49f315fc8ee90a3
z15fc154ca645314658f3870710c3f48217232090e1b9f0f276c1417f94942cde8a164c6bce580a
z81c662842105285cc5227be600042a28ebe76f867cbba5cb9b4af7a6c37b88632620540769e7ea
zc3fba738bc6d19cbf38f333292b4bdfbc15f2f5aa6e9b1039d2f22139a07570a06a04fc14add37
z4ec72b13ba56fdbc340872f7ffd4c89dcc9835fa095380226939ed4d7c7864c7b30a4f6051e328
z344ad9d6e3a59fccb434b6a3a8229c815bce4602fae2348949466b3f32eee356881c25e7ba9e63
zd0f568ec172e4918776fa14c9ce2721dafd7da24a8f51aa6cd13ee452a816c2d61015087ab9605
z8d2f2964b0682a121990f0d1a9e5194bed25a351e3b979717994a5fd36dab3a1a044daa610df3a
z96390a6a2f393d365776cd97262a977efde69ddb29781fb106fe632d5b0d666e123c16e3612332
z0665f44259b92c14c027356db56c2d62e81767bac837e9e27b28fff4396a2cbaade657b5e6946e
zeb7adcbf8b859b8ca5d500ab33406c0d333623e5c2e33003137172e5d8db32a12dc608bec9af7b
z3281447e2459be167251982883d94b99ffd035b131fb89caae1c6db277d4b2ff34e466f09bf622
za0c2bb312bfdfb332004e1bcadc202e1bfa93a77aac8d6385d300c59bf2594bb91b286d190a144
za76da453103ae733c3aca933c0af217352207cda511d62d00598f9247e5dbbac98c467270887ce
z4b426845cba6a52f19630538a22c7860e7e4e9dd8b268410cd5c5c17276654ec28b1a464720484
zc0a41c3757d8ddad8a25407608418adfd9faa7182fc636545911a053af8fb6c7997d35e27b35fd
z82aed4c473c7f2d9022981dc9f9899266f151321aa379f5104fa9316b1f8f179adc3b360bc1349
za4b06bf026f4ea3e6e24b6a9e9521f217484baf56558778713b5a63d8e709c675d35523b351a3a
z68c5948ed7e5f2a95027942902e4f6cd5291ffe1fb4a2c2b8f1bf847cf5ef59f2ffb2c2149e3aa
zb0c98a8045b410f569b3f0bff6f3556e29cd882ab5f66410c93b800fbcd5fb81f417dad1cd2080
zb9e0051ec7a7f0197699cb6a9913b3c867c1c535d322858e7ef90ea552f886ccfb1c15cba396cb
z058ac5b320a79fe18e30ba35d78871f43fdc858243bd39bb21a5eaa46d57728f1203fe4f162bfc
zfa057a1936a11266074eb76db4bc0ab277cbb78605a0e47d4e1f955b0be6cd780e9d2710586520
z56fe33480ba416469956f51f337b6e7dd9c1d306f37d36f4394b11f09bce2ea4878d80b4db5db3
zebf8f4d4c99d5be71ce38946662a3ed29b2977d084d0e54968ec0761b460a7805bd622f5de4aa8
z43f4e29bd8ab63e35c3297a14fa6f8de9ffd2e24e5dfabdf818f7396f0b7777128df42ee008baa
zb6fb8cff781699d33725d2025a454540891a4d03c725084b0e8d6eee1c73527905a00f65c28dab
z1feb224ecb7253c247ade09d4136f5322f7179c57862ff1c196da13228d9de2261b535136e57e2
z9e7f795dc0ff0989250ac788156d0bae983813876f9c47f6b9d6cb8ed0442d8e0268724d2d964a
zd4421a49802f1e029f6f4253b82537c930e93b8a4fe7b1ae2183b76849fa45be2312a28b5dfb67
zfb46496e96960ca5157435f3db045eefbd5db8441c15aef2e1d84ad88ed8975abafab1d1b08e20
z1167cb98fcaba5057ca676bfacd6fb392431367642b775ad467e10ac7777270940e2f131665755
z6f16535e40986ed6a21e4b99122f97b995f2717535547bb2f6f5ad88b1656ae7e49213d40d818a
zd57c3cb10efbf5f2a5c90669deabb4bdb0e05856065b1c87504237d8a1d27b1bdd1bb4e980e5b7
z46c24001f19beca2d018e4d894bad1b1be5e674427d9d4710a0d028e3a2b679bb022a8f2f05148
z9d6f68765f87fc66e81b2b60de2f2baa4f008e57650be642a07cad293194dceb7df2798b016883
zd1fa6537cd133b39c662536a78912a3ee04e6a5663ee31aaba785c4fab8ef14412084c55a3c4be
z239f0f98b169fd2b70fa9847b246ab12a054262f425cd76955f12e37ef96d295a3870c48e09cfb
z6fce4f43e4b8a57013b416c083676df5a8be23a10997d5389bba83f95b73afc7c999c2f23da62b
za1a405b59c9b43b2222d4d28da713e413ab9ce2cdb3d75686f790f54931af38545a24e3f9befcc
z5dec64f4884fd9402199ee19460c33c13e60887d3e1a8aea1c167010f80f91a5937abe61a86cf2
zc5d0309053183add56688b41e5736edb73aedb9ef6cf6842248e37bb19a397a93dcf8617aaa338
z07a7274ad34826a4977dadac76cbdb225b6a99d3d6371437d7bbc27645f2a2bf687dee589df96f
z8694571ab2bf4aba981a9d4855650bfd4c16ab11354011800f4aa348c956d17249599ccbb615be
zbdcc5917958547caf1b7ea6d8620a1f62b9551859ec2f5c04a6dd36e90e18a6d7211f93cc0845b
z89bdf3e41d2bc8cb14524d25c2c13e6b4967b22c2a13db27bd16c81ae6a270cc1bf0624981fc1d
z12b3022da361cd1a592fb25d89dae315d9cbf4f4774a75c9c0e1ea726c8a0b5130cb50c05878d0
zecd92756f01fdcfa77aac526b774331d3f00bad8e3e62e83c4fefff8e3827dfdb3975531d280c8
z0377fa19a0888e5f475cd92a690f466bed344dca6a037b4878101b6f282b79d3eaf66a6bc076e7
zb6db3cc8f639f6f2d5bc3e4bcc6d6ab000325668197450f0d3c7bd8c73818a3db49cbe4568aa8d
z35b93e70e3da40edec9f064d2cd920f02d843eee8a90387dca8c14650d2ceb662d10f11c34b5a7
z155c0fd6366070daaa2cdc64e4ec9e3d723d4aa744b88edd4fd2d9f9171d514d2323a8ff665284
z4347f72e1d16c814bcfe89e4b51719ebacbcbd1396f7c1915a2c68cffe1166dd29dc11ceefaa01
z41da86e54e02ec7e44effbedda7317ea3276f5c72031dedbe54f9c42eb557b3e77cfce2c02fbde
z20935eaba5c3ef96cf0bd27f136409e607332bc49537369bd95f5874c93b66e463f786fbb3eb7d
z5cc4ebb2a25e19c72b87cfa3012f582f1f2cf9065b318c44b0ffee9f7908735da971e22dbdf042
z5138f47d63514fac9aa1ea36a05779e960c3a44b2df039d6f0f21539ea2d72e095d2eaf2fe9c37
zde1616815da8dc281d79fce106f0fc5ed731d1ea8dadc8bff6c4f02709a632d6b19c2daeaeee49
z314ac051be109b58535fe9af14ee392c7b91a329949a07fd21edcb28a8413bf164e1c09da49f77
z4c700bbe1fbe06d94a22119a90691226982358e55e2b820b2ff792f4a37fde005b350ed41e7d2b
z469c5b4ef10bb02e09cf155932ef5e7db4eb8d4ec1a9679ada2513efb6831465c3b2ffce450823
z807cbc807999ec271b1af7fc3b38b7096bfc80d7d0dcb49bb5cf17852bae6479eba1ba77f8c509
zf56363c04054f7f756fdcfa413412345897b715119b78a6e35a00af3b1aae72c12ab6710c47d0c
zbd5239f24050b22618ffa6a45d849be1ef2ea798000696785dbdc739bf5342aaad0af82fb03c11
z3a206225a45457aa0f4eadd0a990d247ee79bea6b509588d8ab6a94adf7a6a4f5ffac88982c919
zdba9f5f89eb94ed6a8c36bd7814823672a4905e1152fe473c422d6389b0ca9eb846f82fa23383d
zc707fa855138c4533c631c66546049841e949dbed50fd720e5e70185168e3109f70a2e7882b81f
z26a422f2a9fd4e18aa694ed17b311278d765d199ecc5c2edb6013995e0f823d08fac718bee421f
zece3d5513347889a851765d00d2fe61a29b2633627ef6db1fbc66e2ed1591627521604d3b5b6a7
z37dea78e3c98ee9169b6404badb7c449f3e67bec5522c96b9768d5a574897a48101b0e91f76e3d
z9ba8eed0e5f2969e3291ac2954210050917e8072e18cf365a6f65fb233e675d5e7b6668d417122
zeb3c02b2d25db0e0a05050c1c0179afcb8aa914eb2c286d30e6f6ed1ee8c1903c01493b10c323d
z559e928577d923cf3f123c56280724bec9733dfb5a4385d94ac86b2fceeb528865ceb4e1260bab
z2e194f44f1e162c151376faf44efd387bd87fdebad573c8a1e61fa31f43f6092391dc8ccf7db0f
zebf37e95763859b4d1e24e676732ebc1984ba69ff3d975575d3696926f9bc5dff09664a6e4620f
z208aa5bc2a5d0a4effc526d3c7d9c033a03bae4427d86f1a06e13715888f4501c57dbaf979f8bf
zb6edb628984f59f6f38d1e6fdc5aa38bea4ad9826b1fb0d3b972715b88224a1b075f785d1a4d7d
zadd85f035aa0c2fb1d9529ad0924f62f28a6ef2829216798a9f2f346e49af0f815e673418c04f3
z1ba957df4b3732627613c61531c13613769ecb57480e34a9435d70d110bb46830abc90bf9a5f94
z441c1e5429d29d88975189f3797d553f6fd7c5a16b20d02dbd67458b02176c0435d25b6cc259ed
z5f3fcf2d1a32bfb632a946cd2e71d923fd073467db8d135c9309a2bcbad49586343ab91087d5c1
zb2f4a970c68feab499cdecf034e45869ae84b39f160930814be39d66ed7e12dd75b84999612399
z63c3e10d3a5fabc78bf08ce5a000ad1b8b8576dea243057ac25df1b7c8b7cc36bb4ba1c3e38b19
z45d7ac674e9c7ca29e0638ad3fee46b981d7f60b9a70726829cfe1fdb60dd5fa65ad92b9394e8a
zeac1d3d6cfd67e5452f14d8ee2933e1833d4f221bdf624d5d62347779f789a0ee178e2c326dc21
zb6ca7e947c1b403e3b5bb3a2b084719dd809a7b7d79d325c4a81a9c720c0afebc7b59beeeb56af
za1454fff64b9397923a95a66dbbdcf525aae87d425b0188b33af48186fabb1596cab1fe9b562db
za914654e6f30882c7245140ace608b216ce405477d196d439613d2bc423ba4370a85bda0a42594
z4df0d71830e2b0682d182eb1b5ede12df1d25b94862b6100e2f26431406ad3e4cdb9b5e7e2eb24
zbbbae1d33d7b102a8a17aa67c7252c8c6ecd96052265592409e6ea7b47b74309746217333709a6
z607b012a8fdb36d1d0b4e9cb7524fe7f3f25e02a1f8b086bee092d28cdb483935c2d9b6abcdb35
z38e84f165c1bbd2519313930ffee03590431d7ebf3a8702a9f73263ff202a5eb6edccf86dd32d2
z3507296a18b513b4dcf844ae0a927ae7e85c9ee06b9a78a280d2131e8458afec5b443781af33ae
z8a22211c7df8a1e541a1dede74f91884bc5136f29246db69ca3e5a8ac32c6082f20fe80dda13c9
zc4a6a1452f33f2c63bab89f50986f87db73f7414d869c03a6be522a87b1d10f93c81b046345827
zadb4c90bc7e0fb2f081127fe9012d2eeaaba1aa9f808a0c39feb562f984a822237f40159224c43
z54ade8876e18ce62a61a8f35781fd3e579c29d3c676f4971a624b0517189df8f08236183202365
za89d0d124e5b63ed00610ce72224c767dc4c1484b6c239340027cb3f24a3e2f87c48c48509c27d
za21bcacce293e513b5223b68bc5446c9ce3dd92e1839f3f38dc52d8a335390403a6b4fbf618d7e
z4907945c9ad9ee08195d6249492e98ca673b50a5fea7b8847dbfc5ceea88ef3e2f89d6d335ed9a
zadf6d98e43804092c8ae12ef0032cf97ed0ecf49a8cf9c54d60a2ec2a42365b27ffdb81ea30b58
ze1ed2c3499edce3fdcf99915d05676b8ee9104446425809ee3f0342bffb3c10911f6a4e3d984a7
ze9f86dd55c94d8d84fd6be3b5db847ee03ec8c8ed12ca3a43b0370b7ec8a1d464a36b6d3fea04d
z3bfb083a60916d5a8168ac346e67c87843d9dc0932743984489241cd45778fc38a94a27865f659
z4ce12f9ada1cad35010292d2fb35b6064a787ff4f1ebe8e448c2b740fde1e1e0007cf883696bd6
z175fd355d7d38d344be7072187e7e6800de0183e039e5339ffab550672b99e6e15ed2a7609a9f1
z868eab3799d1d4a6172b0cadb9c3c0c63e1b7b81c07d195be88e09efb9eb30d36a2eaa7bde6f0f
zd2f83e5c4732fddbcda17cd3d5b945784aaa96f3992025b0d10e954e1aa56a6a39d3355a2223ff
z49d27340041ea2cc97dd51093bd4abcf3d8381b0b7a947632b0d98fb96a5f4b54009c6479326b7
z944d58b2a09aeea583fa06767a7bfdfc1d8dbc11892d50d7fb6a1cdfe1a21a2b404e35cbb7824d
zfeb04cc10262f1eb09357446d6cad73e70eb6587c6137d8e9635691d9ee7882871a7181c06d083
zde9e9947c5e4d4f6d40d7e6dd09498739242ec54cac6c1bcf3e5794fe2e9f466daa26a978be210
z04a1dc0faaa98413b78107372c800d6c9221b9406f6abb39aebc254c7017db9e827f5005697fbd
z4409f3d3a43bdf1679f9de82d9e0e88977baea6d49d3d529682baa5dfe85bd5a85b79c265301ce
z74750269e5a61d64bdde7e16d9bcad506cb7bb4c6328bf7090bd888b1d00139e01d28c7e8321bc
z7e2881003495e38faf93f600eaa664d20adb6e57f387f8d6fd7a3c01c0f02fa9c20b899a830079
z60c9d7bd95011c96606892b74b02dbd9038e95480a90b66a5501ddcea5f24467b71487dcf2cc06
zfac81b7ae2005a6716afbdba45a2538c7b1b5faf15db11f48a2be8ba0efe52b6ed1b957130cdce
z039dd292cc2d411358e6d8f7992c1fe68e98db27e68a8c89d2691886b4e6e25790ed106ed05338
z0fe7c170cb06afa12fe2b09435385bcbfb248c8dab54f4ca431eeeb4bbe3104c27b3c8f7ba662f
z230bc448a33629841c0b4d01f6c4d63d551cc030fdd8af60a31561d3cccc77dc84b6acd57cd7a0
ze0413ea431c73a8546e36a39397336e5b730d3b550dce748fa30d1e06de289f3d3f80c3ec93836
zf1ff9069a4e2ff32a51dd1a59912f6c0309609bd33aa18ef075b9f722d1b1aca9ab774c39d28b6
z026b779a7a227cb1e786f102fa6922102c530b93f9463fddfc36fcb51e8a35b0886cc3daf510a8
zb29fbeff9d59ad2b760d1af5b047a201e170be98564756906f75080cf7e3dcb04dfea6c2d0bb52
z8f44b54db74a4ef0b04e00bbcebc7eec00fdf5755fe99423345fc47d791f936abaf593dc378ba4
ze301ecf1535994ca73a248e64e9cc384f8925dd33a1fcb356fc5c13e465cc320707587bfa70323
z73d11ea5b0413a533fdffed4eb1a1ba551da931a6316dfce632f82add0723145602afef528f483
za4d30709c7d7ec270385fe9354ec33231c47d166feef77131e99e09b9d25371cd6164473cae908
zc0b6903809dacb7e7bb102e7ea5f240b8135c4b0f55e47e964fa1ced983be7d31d6258d20a703c
z72b7520a87cf14ba4dad6513dca247147d5a1fba3e0dcb9fc9ac8ace794df1952c9f6f42ab1bc1
zfbf0828789037d115845cea08312654bdce53db564e47239efc30c9ba33193af6b15ce4ffb48b7
z257333956570828cf9527bfb6ab4900b18355607f035cd5225a7a86e93671adf9b4d74b1ac7d87
z933cc44e9cc89e79ddc8bb2b82d1a0bb2b69d5acb8cf8b2929875b56645d32078524b9ecd360a4
z0a3b786a741acfa988f7506c75735b3eb52643114039c78383887d4a0dd9d1be4548e2e25748a8
z9fb0c0a81fba364ea2985d7091cf4e6e56eb1f18035e90fe3b7176c0f67d57189603a9df02ff5f
z362338e2b966233bb6f8e0c27c3836a236ffc079515e8ee81bfd88f7a4e626a2418347d3f44036
za0261e19fa542c87e509724a01bc97a8ad1e00bfa246acc37c0588c7f74d7b65977a397aab7081
z374e901316031c7d320d3de89aad4a4b0c3a5b20a3c79ad9eacb84b2f7760ba86a285423526e40
z08acf9dd8d1e545b17daf33be27984296fa79bd4d3d6482a1783206efb5b6fffcff7dce31d8c26
z62f331440e9025e8ff95cef00d565656f35adcc2b88f85c287bd1d89612f81612c967def6cf055
z623fa5ab190002c16098bf9bf44acc4cb2c5e1c4cc794007340339e600f45491c0b2576c30fdb1
zd5f0ddca642309111487546af85551e817822f03bd5c0d11b1f557d77ed3be2602c2f66cf16316
z2bf3b77c06c07d767a739633bb2c217583099412623a5fbd9dd575313af43cbdb3ae62a53a9e94
z1ebd01f1eaecaf7278d8f3b9327095895a5157e275f0b113d026867940a25d0de755644dc4e4c8
z5ea1f01b0bcab2e5757864b3058fdc1141c2e1b3abceebdc29255d9a304660163ecfa8e72be9ee
z444bedb9cbddb96248fc16bf7a70cea83ac08ec65e779b015a1e308c9ff0ed2fb84557af8459d6
zb1372c55fe45d5d0fc22528b0572fc7ff400c58dbace1bfbf66659a9f4eced1c71f46ad987373c
zb11036437230d0990740732270084d227dc7a2a5de454bc4d6b2a0e6448d1e0c05208b6573966b
z7742b59c1bc54239c18cd58fa64bbd6ca1656374e6d018349837f7753f2ff9557758473b227221
z2858084a00f5d7e0ff821b6d8bed67feeb46576b4ff774a70dfb358e204bf091d8d68cc1f9060f
z6cbcbfdea0bb9a53103884d9fa8416181374c86394cbfd107d4ee0d68257045269f581fb52b7d8
zadb2b5a0a2630bc78c8abf6d05a87ea10179ac516263f458a98189fd298986efcc4f6d521c2298
z257fc8508eafe7e7b5b95d847b19061bff191d0a865a7212e01fe713e82fd5b6491a7164696a53
z67c9295349d370186c4321ed59a73bc35df26de687a0549a6c2d7b1f904a5cc1c74135793caaca
z7bac4d6c19389a798018d8cb046ce9a28b3ad2167ac41bafa28612f0b97fbdd7f06245dbab2ad2
z8b34d1abb87ff7f269cf75a1793c05f4eec84ecae6cd542923ed5dd1a15ff640b7a3e25d50bed2
z2775825d2b8ade9757ef4ac4dfc324ff9385c31a92b92f3cf8a139302812d294b735f22e5e27ee
z7caf2e1a5f5460d087d3954224b3ee369bade4ad10a2a363b92dda065a197b7a6cf2ce6c569709
zcc089e0b405c4b12aed8fabaa216881e474aead94a17ebede27b21ef367eb13b49cc499efd8aad
za3fdd54e409f21b5ad8a5170bc730093d4cb9bfb55430cd0396a5d9c76e66818ca795771063b6b
z13e2514f21a0277007748ebfb91236d2d4b8eb973fa20196df1db6d97a5f8e7cd29dc0ed81a7e2
ze6f3816bdc7796d0eeff23bf2da3baa14f4e9219139cb834ebef1b353f85d32af1178c002cc703
zdc07ed86dd6847969372ecac60c1ce974f27ec72d0286dfd75662dfb632b3b89f16f0d8a13b356
zc259c21231dc25e540e0b8bb3cf3e5d33db6ef30834c92cfb25dc7baa9f4fc803311cf7b0cfa27
z8b603508e5a0de319b69d8f69ea5e1dd210edf0af9bf3eacbeb3a8748719fea2a11e606daf3640
zc401db88a0a3060bfefbed55fed8ec2be1a167707de709130ed0811d2e2381b01fbb9f908de682
zefd3e03b94d5c6cf4633f29a336e144bc1e7ee70289aa95eb80f55f8742ceae4c460172bb7f653
z40407f85d9f03b2d93eab8275353b422c72f213a78f678b5c68113495b58ecf316e44cec1f6579
z1b59b27f2cc6b71f7ae1b1f13a9b242197f5ba23958ec170fd78416dcface313098292431e6330
z7018e14a85c6ea1e1a84c784b72532a00db6786a663f4e8b64c36c1e77c7a1dd4ced6b75e8692a
z1256dd295fac05731c6f513a8724277d4baba5e9f4b7394b01d5b06260ffd803982bc240317e3f
z5db24962cd8fbef252c79213d1e568c2f89f80102cb92f35907bf41b5194f36a72f201e6f1e54b
z04b8d08394a811ae3334f168cc4af13df9fd613b0a27c31b11c531c90398485aac6c1be7e079ab
z37ad4169e099f91556096c49a7b2623ed12082bd96d3bc35363c79b243bc418f473629f9e46737
z7b4d2d729be1543d9fc778006afb4e406e00714b12dbed6d42167af83bb5acf9c4778ab9254ce8
z584298e2578fcc3f6eba8c497d9df906590f6ff5debd995823292debd761eb635f8b60c26a975d
z12cedc57815ef7fb79001d1046c53d1c58e4abb163a858bf4c900ddccc2875384943746fe2369c
z20a804166f10384fa040519eacaa537bc5b9b358da5fe10742e71d36804d05405d08caf13fb7cc
zb4677f3d4e272c761e3e93d52414a582749e9493e16c6d67c1cbd5bfe20caf8dc30a79484690a3
z6e9532ee887553cf6846ba0db7eda7abcd7fcddf5dafb9614a1d34e236fc5c34099ae58cca18ce
z73f2f2b649638d3204cfa00958818ee65e9f782c1ae966471793a6a8a6638252e6436f3db0174a
z4ee51421399922d4aac805e81f93d089dc99446699411ae6ddcb7f28a60940d0e257c9e4bdf49b
z72fddc4a0fe9d518889d70e22299e98814339456412fbe7d1c21b3a98ae2bc0fe5d8d6c71718e4
zd2320b2f7437037e6f8e8caf96626a0c25ef9d3844038eaca39006493e818df5fe0104b91e8491
z9f1bfceaa8be91867de56806b24736da227bdd3437b18b1f5fde9a7941e61f887aed226176b044
z118e46fc8c315a50e381543888da8de0b9c3893f375e10aeecef389a879bdc5348e904dea2ae92
z18c8e75fb2de1b2f30be125b144b713b721b709ae2bd05007d610965b84e271b9ae48e2fc273cc
z14844d527628b0f20af6209ae52bee2db670286f7d66615fbca6e0aff0ebaceeaee557ca6d730d
z4257dc7c3b7b0fbdae10515343a131d7cb811374a208db66baed938a8877f4d495c00a02daf7ae
z34a82d901ad9a9c98e0c0534c69adcf5d5f46e2647841ffcee0193d9ad2d2550701622442c4ee6
z21eb3b13255c808a1bf98c29a19691fd1392f86c874fc4750c2d2aa5e896a781bc44f06799082e
z26d9be36dba41f6ecd9e53dfedfbc1ee637e4066ee1455ff391002f48951cdf3e4f46083685705
zac4203e94ef5c6e1c8e94426a896abafd3846fa33827c1af970db3a7a630237a078a4cf0aee5b4
zd28fbfef9dcad423fd0ebb8aada624a9e5d5475ac668261c671d61fc569509631c815d16adae94
za210d2e369da387198a03f7af5b5dcd1576fb5a96f615c2ef3af3e4c11e16c733595867823617e
z745c01c353fcdc7a148aff820720f5ffadd364efff13c14f08ccf7d0802ad62f209f1624321d9e
zc486dcf7139ff46aeae7196d3e2423fce14428231ddf733c04a8bde38375df4c047c3d607ffc5d
z539dc3fd32818c2a3b4f9d6c5d4593fee7d3afdf848a9a3082d0ba9f9302f00f2120831e7d92e5
za06f0bddf8692b6ff32fa468c6236eaed3b17387a718199d917bab5190495c3762e2b0a53dc57b
z973cb5825733361519ba202d45a9d2dc092a954a328873f4f7eda7386ce6ea87dadf81a19b1014
z38c69fd39f3452a1c7fedea297e7416f701334cf786dbb06f604eb425aab8cc2ed70f66276466d
z174e7bdf91ead652e934673e81f0984b6aebc834f89e53d51b87ae93399f03427637dab945547c
z620a622ce69eb91ec6788f124a3353bead3d348304e0dd07b1792a0b39a4dd91497c0345d8601a
z39e1fb7cb9641edadacb55bcb23199047da23c8306e02d299c0e5ba6c7813d31f88fbfa6d926ee
z986f93b15a0ae41a6d5ccc0f6ee93af07f0ad48a31c404d706357d3734e2dac22a560bcfd20253
za7f5b410241d5d8df7be61153962692f6f4023281af8251951443b9434a7f2617e3795a52073ed
zc51f9dd328e83cd847328544e34ab9652e6db451906f905ad4276f3fc8b9890f02831b79ead33d
zda7d81adcd74b4f7e2bcc4bf9345d5aad40ddd7943190485ec3c48523c410c4dc0ff2e6e15cc00
zc28ad22862915921505c6acd18a5f71c98ad0a1250ac8f419ef91d190735f7aa965ec0579a43c9
z83dc15cd377b711e38cb654857c676673054eb6dc6e391a887bb7890878861d30a16940eb4aebf
za0b914bcfd608f010db3aa8f04dd4e25623676ac24810343220b8ab7248cfb1aa5cabe11d31c43
za2cd7783af8e4c804ac0e2933bfcbc002567bcbccce261eb9b35dd5aa9b143a9bf98664ba7a549
zd9d0f5b1eaf617ede03d643f3c05c589174b6fe228ba8aab87c799ed73a00f9378146958cb8ac5
z5ffef0e513914611f3fa190373443b09deac5d2dc6222fea82c459e16bb1ac94b61b885f57693d
zc44d92577480cc33e0458e8164ff8d3051205bf591fe75437cfc1e54a311392c35ae33e6a11bac
zb0302bc28bd5096d9aff651cfd41d66eb647e89935c0105f70dd48efb2543d9b463121484d0251
z9e9cfe485ba961da9b9dad451dc1ed0ac131ac545d2152402f66e2327e44ff93d9b44e30d6de3b
z40e64c3e29f3a745cd477d89ba59d04da335a7b229f40e00e474c19dfb1c0e444612679881f80a
z9d9baf83a012442c9c4a0cbf5af37fedca1a5b5fe05d3724390ecda22daebc25ce934edc9858d8
z5dafa8727aa4587979c661b848b08d1337c65a15eac5a96c1abeb539648d4ab749f791e5d72fee
z89b7465b4547cad5cc25e07af08773439357536ab45866c23506eba5f9568fb92774014a792d27
zac8b18d30439298805133e25a04d0a74392b277a9e4d2be5c4ac3363bc7eecdc550f5a541fb44b
z10709fa151bdfd76adce271e2ea467d9deea5d9fa1e85c76ab031045a4003babfcff5a15edfc13
z462c8a7ab0782a2040da667a14e74c576977a8bd618bedd6594ca6c32dfa0e554f550f8a062658
z73eaa63f505de08f6fb69693214c972862f0d1d02f5ab0cdfa9c38b2f95524421015248f9b9efd
zb2831863e35b5ea8f9e5ee4b78a8861321d2faf8c82d09ab4fc7d06e065552bd3eca18adc5421c
z1b77041565dafce21677a82772f2db44c4355f71e2387ab59201c602aedeea2f931f7d378c30d9
z15d7affb573549dd033668a4c0906aaf074e98fddce78865ff0591c425792f87dafc76730fc8ca
z244d6a592647e699cb0c4b8f0dc0318f4bb9f47002e40cd261580cadc1656af63dc2118ff4c791
zf19e96c50810c01c93f73584213c85a447ef8ad6ac904cee52bb1e95bc934c03a148962d71c531
zdc15ec7750b14fbe438ad861e6b78518bb3c4345b5e8976a2d09f958ce8de870e11af413119715
zabe6c63f6fe4e1f0f4637ec74e5e1f5962a62494393ed4985d521448fb5d729b5df8cad9c1ec96
z07dca73f079eafe21c0548f10cf51c47a5527fa468c1af541b5bdc0f2669c46f0c38bf9bdeab72
z84e71730d26def63b0c77b25928e55ecbfc180e8693d44b6163fea375fbdbac9b09d8e3c58b7b2
z917b6fff1efb1f07d867e33be6f661e97a430459d97450076cd40bd120b277bf0f4f76c57c79c2
z71a7d0f74209b30cf954e1304b2fb9894fbd693ba31b3a4c156d8c22ff9ec9ba32c1a3d5110c0b
zb858d7e781ebe9ed52687f85a897505c99b6e92fcf029a022c3e2c22a5b1c5fc5747d7ff9f1621
z8e63a6c72078ccd0f3b5c6f9278947989077e3dedf4bbbe0fce88bb3b0998588389de15110ccae
z61d71552c556efaaa37a5bf75eb55deb66248cae43dc15a88a9b2191deb315680e67c01521e424
z9bc6e084b301b00c222672c2830e56c6eb0838da0055a62a5bd138d62c56f2e7db4d9b29f45029
zf43526e49f0c52a47cd0554411f976cabbf7417a2149d1c857618145850666fd0444745619fb75
z0a52057e49706875f42b608c1425c5d77f387572130b177e8a83dc764085cc2431a4d94cbadad0
z8b3a06a618f92e42fda949972c270e296f6ee4d41b68ecaeab295db3796879621b7d33f46c9102
za43578947e6c9c472620025b6922c7d7296ed1dfc94544f9d37341a2d953c88e89e44bd4ef1878
zc083b6837d46327fae6e7767383d5d223f153c1c36b0c2feda998952eb308ad79afb3fe4f03974
z51e8906cad9d382b879f7a68daa659c4131a394b883feb0fdb6f6090ce268a137f428137f9d944
z918d7f0365ed1cc2ca0348dc0e3abb0ffe2b2336970986a9be6d90e7b6af564861c69187b208d5
z708763f42686ae72789d0c6e79624cc5a30c83e9562be2804bdda0fa394e989db767d2ae3e5ff5
z6eccc18c65baf07f85c1d4e4c3997bb54b739b0c10674d473d57a827c8e52b06faa8e6cd6dfcc2
zf3f1d7b8119d1369be14a3cf980ad17bed77d1139e1368a7b69947f72bb5d8f828da5fb8e31e8b
zcd4edac2cd068af24f126dcb3ee00d12b4b4f59b5488dad1358da205fd1201819c71cebc33110d
z36075bc4ab3a2bda58ea580d3965ec7ef84b787af7f0f7b6ed093cce5e6807978dd2fa25d3bd4d
z64ee9098803c089861692d7010a6e1d07c554938349cb560ff315828463eb9a412c35885da7403
za50974ac1c9ecae500b74c97b3de248052ccb2166099524ba5550febaf8d9db6513871e496ef70
z24a13d3cf8a38f1601c67458cc55f5bc7e7531b916c4e6840b4836e91b2ba6781f207b1e45f139
z82d72d1121c210d81c4aae837139e07253eee7e2839b49e5211f2f867afa64dafd06c3d632d7d6
z8976dac16976e198044c2412b39846c8f7d76386d8556189e17da26eaf4777fc86678b758fa2de
z1dd17e82dc2f40df2906b03249977ab93db560d88aae91d8e45b9735ccc84635e91fb5a3866e5e
z94c827aded5e87963a90494c169ca9d6d7e3638e7c08d48c6ab54fd9467a9ff9e0fa5ace4108f3
z9cf29419505f319e93351024812cb373aab2520f4e899d488db199764be186fcd59074ea21f157
zcd00c2db0e6364fbde33269f93fe37c5e2c62ff3df25304db67e8bb3cd6ecd9594ad17ea454d71
zd9a3ad7ba9d4cec0a70423ec39672509390ac552a51397b7ae874db31b0c0f3ed2cc2194e6225e
zf129f9561de57f1445836ce56dbecab8869d21e9c3b5091b999638fb4ff546a8002bce5114afed
zf50411f98cbdfae4e215877c40c3a8b0c288b66a94d9a1046f163d15c98d3276e309e2828b8269
zb192250049850fbe94210f7173097c1d699b06caa1a34f6190967b5728c3133ce792056f6690d6
zb16fc1cf1ac7994783a2e16aaffceabc593c0190dba9a4404d3ce864c73140f247ef1145adaaf6
z2a1737bc84b4436b5568ac937adc14ea8a2b55b1edec03becd295a78d42c2c53967fd533c9919a
zdb77494a5d7a54d3045187b766cfbb6a9bd1363be589713cda9915a617358880f049a12ccf4958
z2749aefc5051c3b0cf8ee3329a66b3b32f9919a18d7bc2fe50c47bfbcb74b2869fb7eeaf80b1ad
ze3cd5c81328d1762564f4a9e71a8d6665d2657785d0559e2e614f0885a1a016819a21df5797413
z5fe45d821350adfbe734d34ee428fa2b25cc087d30ddf5ef8bd6a0d27b34118d0ec3755c88c35b
z8988861a094198d402d9c8d81fd8c06a57500ecaabf95410ffa58c1c8c8c9964638560194ed974
z677c348b80b95dd80fd1167709c792623da6d897d9cfdcc84493e757b5daa40c49082fe070004c
za96f670a573b9b28e925c4cd7314df697eb52cdfb472d3ff4c4c9be35144871dcbeea24b5d9520
zd6e5e2882b690971831677f88d0d9ca10def6bc52dbfd71c96fce75f7cedaa688c1181adf56d04
z459c3f2b8d11728bed674b57adac6697ae4c3c9fd767d7a960fc82de38f311e42acbb07bde53f8
zd8f8a1eee5b1ada8c146bdae35085918cbef237d3fb9638310b41003064e71ed402ddcd028aed5
z09af84e7be0429cf86345ea609957af713dec3b00a07eb625de41bf472dc9a6508ca21eaec6fae
zd0d9eb9c6157eefffde6d77e454b6f17c238f946f7ee7a8ff81df74dfe82694b8fd0570f33f4fd
z27bf0c7008535eda63786824e7ee16160d323763e2137fe5bffdb7855f4b064729ee96bbc1d7af
z407cb39925332dcf787d37a6d132a4972828a484749ab04e9a5e424315cd1a48aa6deb8fa1b2c9
ze771437e97da3025c8067108bf6f9650780a1f62dc4109c23726386a0890e1f9557cf4b3e873b0
z719410b67fa10a561277c259623275dfba56a76973a47adb2fedae70691dcc9c448d37ecd048ba
z854017b80bb4869c78255d693d8235cb584bf77884792c9e99f9f76f8340de1840d1540bdcc8be
z70c6e440e71c348254831603d51ba8bedcea8f217a133c76fdb447bc990175b1106008574bb1cf
z5e2a982d753b8544f78fb0f6be8023d169740af68bdf74580f72916de82a5c428750423f1c668b
z79e28cc4e00be7ff83c8992fef6b4fa65913f53f591151fadc6e83941d3bab224720f8d3125b6d
z587ae03c481ce57e2b6646cd4a29c0a91c8cb768149eb92a7fc32c95875643a79c13297ad62e32
z3eb240d53cfba19b528cffb6eba994051946a626ad03c999e7b82de8b09d76405a5ed76cd48391
z2435624834f62dedc24b4a6f9a48861ce50731c187fda3ffe72679aa084a9e70dd9d4c09c25dd2
z658d3f3415afc08996fd2d571b2d2ab8ba3009ac7f67e178e1a1edbcd65720781a4b5fa740abbb
z461ff2323201626796f52a634b5f475d4dadbcabaeb14153e7c4ae2c15375db2e2ef2a17ba1f34
zefe0081a7b924a91f37393bdfbbf3edd3d7188acc206f47a755f1c265af68912909a7a75ebb350
zbb4a4bc27c89f144617eed8da4416d7556d7f45a6ef067036803bb56bc771ef0f9c5c121572477
z3a002629bd4d4cdca427ad2ef83c39fc9dd787d8dfc94a8ac74577f8bb4dd2d61ad5e274eb0ff9
z87fa2aee433b21b0fbc06341eecf7b7243bdc4709cfc7ab82909e965ffd3417e091b35b00c78c8
z6618bc3747c4b44728c1bb88e1254cdf05658af6dcc323f72b9cc3df33559f4b46197785ac057e
zc28458828495c5b9547f35f679112d125ca6f676b1917cb3d3002fbcc9639e355ff7e8bce0a50a
zc7fe957bbbcddeb07cd8cc6731dc86c8b64cc8813b2103c385a001d2c4134d597644f9cbf2f9df
z7865671ea7ae7735c8341abd7037ac8d0f8fab1dc0ec8ce6df4311d95cbd49867705781b29a22b
zfea129255ae2b9dc89d58c7495c6fc205b5c33e6c8cf6585909e0bc0eab6993d9a648205a6f67b
z29de70d775700d082df6372a94144b7a087200a7d7cd57e518acabfe3858f34f1adcba7666dd0a
z5a4b1d2375b147a973a7f2f710ef58a5a6427ba48e7062d50ba17fe44a6ff116a8475b616de440
z1e86f092c28be13297c3ccc07370db60db10538997c2ae1e89dac84fa2e7bcf8d60cbf8a41b6a1
z00b288723f18fd524d2900c6c2c48712867252144878fa4e55ea70d571c06180c6e5ee3a74483e
zc3c3844615acf64a2b7a8cb8db65b9ef82ed03a2d638dbb7de11e098f564eefadc9af8043ba527
z33e19b9b9021da11310371711d05a7479b66aa5180fd32b06a0278bd64e0f65cc1586dff075d36
z7062e223c8a342261c96d3b7259f9691c92ece25369efbb92415e4e58a953c70aab74c84582028
z9a6dd2ff9207fbab8d57f16c48a6086b6bb720486fd743d90b297cab7589b54a3a29bbbdaf236c
z209b6639be6a15794ef1b556282231e07fa1caaed78a3c32b419e076ea7040030ab415251ab278
z42aceac62c627a8c5211949740480d154ebcb537b892e4969e842eb62f3b2b918e0c953aa1df80
z2fbc7a4ee84000d9c5ef576647705fd82c015b57bcfa62336a8136b7069663f26d628eba6dca58
zcfd97a943ba56208832527346e10fcb59090993919db64848ab1e83a3f8ba7c4a6321fc3e758a2
z146b6f5f46e5387cb14876a5511cba3fc3454dd145ceef331ced942efdedc9b521fc9a9ec92d60
z656de2bee746dc3f50ffdcb067da04b40d78f1cf69db202ccedfdd9f438b84b66aa41df2bd147c
zdf14d60401b981c887819fb166f87e5032f5360d7270bcc698214fb8b388c781a51119d58cd6b1
z81504e38bccff508737517e02c4637c08f449b57d0f853d543c5f799a6f5e868e5cecce391bbd4
ze51e237e01cdea7380e7cff5644cddfa66c2e358855f035f9fc6ef795f8a1301a42822814e7912
z635ae969d2e8811a247efb3b94f9955a7d5e9d0a0a0cfaacb1dbfe87340db3c4cecbd9e704594c
z4ab905358d5b86a9fbece444208826fd5a4f9bd5e866e14213e5d0dc54d08ac98ed9c659dc681e
zf0ed542fc5de0100ffee80d49702263355b96a3f3cc35d7a8d290b47534f8a7de699a6c5b0399c
zdc1b8cfb9b433af4260cb747bded0625ecebc020b3aab11deb5f23b07fad4e0d9b2d95fb5e0d99
z2f061982283d05280f736e5d0a64dd32b2f719bfce4ab73cb3eea74730a43a415d0c15ff786f7c
zec63de7d4033edc2589809b5aa77a0835ff61c8f6d72bf969e1d407d8bd5269ae605ddad36bfeb
z4247acda4bb39fd5c144575e462ad016afd5d812cb63a3899e2a6898b1b09e945d011c1365d30c
zf246945464b1a25259badb8d1974ff68ded8558d72c67a6252f998a6ee5743fe1b2256f6fc6580
zc15c2e13815097191059776287e4ce300096424fced1b2debb1a6a836b9d8095758d945cd16996
zf170c1825bfd076471dd8dd708f3489885014bb8b4c65fea2584ecd0673845345d051763ccc2bd
zc22b4c2c9d2a7e8320a910b12c79611f6d4c748704b4a6e8f78571568369264f33824bcae238e5
zb468e9f462a66a8216655f423d74796d21d2b7fa000ac7bfe65d3ee440674498f23a5e51a62fed
z7866fd66cec861bffb06497f59f3599df97555eca759aa02fb4e1dfa45e81e5806ecc7ea7377c1
z7ac5685b4b9a1c5ef7cb48c96e0f6fbdf4eb29887898ef3272b52c30b42ae36bd3329c21bc9109
z7f4521b9dcc16a881f94d68a8ebf8a1bb3efb96e07c7472930f14b8f4b63aa816cb1bbf6d09042
z243d812a9437666ce0d89737b010ea96e85a13f75d91a40c1b815ae0ee9ac4f116f2bf7e31046d
z3275eb77c26bdbe89adcec2d7d46d4095f54241730e521cf1575bc29f04c67a9bcc3ca052547be
z980198787e9c1e7d0730b1b1f8a48558d79661415f3bbc640a382cb09a0526b60c6398507309a4
zad367d8b9580a69910da9a106ea27b3551d910b34eb74cd07a3ae3de047a3f5d5cca196e7ab97e
z0cffa947ae25e88ba4df104a21614e676c14e1447f636ec1506b4af96b26ca840aa4a6df6d1c54
z607be06ad3f07e04ed15ccb8fa48232d8aa2ba72bc44299db14188e825753c7b62ba41e8d90a67
ze03a290927363ef34f64b9f8f294ddef2a08bb1fc33822ae7f9400186a13615fa7906813846efc
z946d1b2c09b5def7cb2f43bc50ca47b256b3a3e1a0d74d2d86b1178cb1180250b9adf51b13bb69
zd38363e2154ccb3fbf9db8ea6d8729073b193533ed7556de200fc7cb5aa243032728763c6f42e8
z95235942bf63c265f02a5a114e8bd7f95b5fdb44dacaa7190a4e65a3b180b56909334ec363064b
z2ee8b589a9f822170652d09b3447f1f027a4bd64939cf640259aa9e5bc6ff7b67fa4e6481db9e9
zd2ec8eb7ccbfadf82bc27db327fcd30d3fb63c9eb2c3b352155bc7cb3f1bd92f47cb85ebf36128
ze1a6136c0d60bda31c129b5b53c99d072a5e4af0fcea3fa4185414c2010e6a4e740ef5cdbd4d30
zfb789056635e7f7dc9b2ab885a51d9b50f1137443e1e93d6cb9ef54478d72c79edeb0d564967c7
zc7a9f7c01750b556c29a7d35e07484ceebc0e995ee6350aef04bf609c6df47926572fdcb2e5543
z03663c8915dc4235bc0abc9423cf2391cf968e3d4fe5470776d3d93d34cc5c71f4f028f4cba0ff
za5a99139dcfc6a055f10eb3c44b1a08e50320ee9b285ee1c6ba999651083e5624e009ceebb50f1
z774e8cc1a866646b8e1155c26e2c2f2d33793512b79e0f1fcd13d1507e70e794550ae70d37d753
z7b3704ea59ac856a70d44d56709a3d68f9cfd390201bf4e921a104e87aa76b94d873534e84a5e8
zd57583cb598e96a329af03a83aea651fc0c29cb1eda059b76db5d7835cbc470b1ee9293bbaa871
z88c2f13ce94658d8d2993c1201c037da4f32757270b7ba027f551add0377995429625db04d0448
z73e74b189c0929618d5a0393c5e66149118b5891e74318c78ee82e1f5bf0992e158383901244ae
z3096c85a4c81626aa4802856a6a6121d9ab0f18ac65fab3d376c74cb0597672acddf24bb3fa514
z63e1a35b13c2836ccbaec676da0f96bcbdeb2b7154cdde3c0714c6cac2b157b7d4593e66c986e9
za8f63efc45270e32016764e40dded39cebca909cbdf8b7cee953931b9aba143e46f86617fa1d48
ze5d398397ee3e98d5b443d38725401cea678f570dc997e0fb37b022f4858799af10f823549e946
z05c1fde011f26fc4d8ef054aeff0a5771ab000fb5fc2570ab90e0afe7be677f338ab9d8c313b50
zef4e811b53be47b6c98af3d7ecbb85fcb9a389a76b7bf2a8e1554cc593f5d4734d74a13208c539
z8e34695091a82bda0f7293fd4d1d548187c644133a3e50b2466a45c583232a1b0b15736401e9af
z8fc94ef843a2b515c28f6a3300510d9cfed468110b046ed4bd47d837e4e4a841874b500addb496
z99edb5a192f0dbdb3f0197b67172d261b96614e1dcbefbe083e4a9748ac32fedeeca223865f92f
zc8410744cc5b83bb52727403aa281a5f5a25b7290790e7b30a127606f55bfa0066b15b503b5693
z79bb5fbb4dcad2a5a26c0af7e759faaec58208611a525b0d28ba87b455b35116c5817e8531f16a
z50293212c58b85e0310fd2fcc3f2056fcfaeea229b6643039fddab821db35fdeb3a1fb757eebd1
zd470920c4cf6676221eac26c18a5925a9778e7b61c7aae43d02f39522216c649e7f626529b37f7
z31fa1a1493bdccb72d1d61cffd7467dd983a9b43ef97ee4733ba403cb6cb9d1c5b0a0877972557
zeeea2fc3228c1317db43816556d96630045b78e26730f59f47b8fe9030e2301043756e13427ab8
z9d4a8970e25abf852d67a600a3baed801e2aac728dc4a31cbe8683c703cc6fc99443daff8676a9
zed0adff6c7f2e317e42b819e5025857f6edfc64bf9779c0eeae45aca5b638231969219c3236a44
z6d17a1b3315cac8474244b7301b7c1677abdf0e87072796533b7b52cda5e94c78d551dd1b3cd78
za86acc4c4574add3652976f79cc38773d9fc26675009b785f5f229cee062eff746d02172675549
z453ad2e5d287c3e8dda47e4fe58985d5600521eae25c8266199ed49134c3e05780bb4d8083e842
za01ff285cfa6e54e8599a52c2a47dc122de5d3d415b51d37bfd45f56ec140f7dc9ea7437a196fe
z71df9e4bda691da002a9ca3de239707426e13000d22ddb7f536d5f6d56f391756b1a3fef004174
z9689dd1fd3d16588ffad0e077f1d8462e425a02d39fad1443ac0b577154c8d22c91bff46e4d798
z02be05fd1cfb5bab93f919e210ed9464c2c2e70bc0421fa98eedebebc9767e1599a8ca144ae691
zbc0f88648366b34fc29e26ea5ec9f352a7649c989cbe8de9e209049aea1772be0f9bbf3dc2bf99
z8fefe5928deabe59f483164a731bff8f8ef127bac75ef33b1e8b9b883066b736e8a18f06f7b837
z5a97c8216c1e05a93beebc0c1ba6135572eca7503d6fd6917ac5bc2c566577ea62c019cc47d10f
zc3612b4ca43a657d9095e1dc4cb16aff5f4585fb9b32ca668bf202b6c3583a7a2a6e25bc0b1f11
z7705d30a1898fb4fda33e800c9bc48a13b70c25016a95eae629c6100aa16506c29b79292bd3d9d
z279bc00f2d648bf76c813e90393423c332d8e5400c3d565206616ae98f28d80897beb5566149f1
zfbd5b7b09573c589dff891dae0f151c3e74af93a7904ca2c58e485208b32a032b7146d1438cb2d
zaf541058900772c3b4cd306a128283bda2e04eb80c9e0aba5579763af13274798b51c33e649114
zfc005483cbb86a7cc70a207c0109266aa90e5819e5029752468101052f018320f051723672ce5e
z3f37b06f62bc342f64ec1942d9cf4d129c87a8cdbc7925475f7cc036fd0567a4351b400a94625e
z0ae656f62174f668ce94e6e47c78e9272b51546df052e21e75bf24d7e86d0d83cbd8295cecabf4
ze05d79730bf3301ea33ece8bfdbc26cc2c8aa352c12203a88265b090662861fb84801588f8c331
z40448f7b6f8b468df1dee0e75f39189695175479fdf8530cfc784493ff0267d98bbbdcb366ca33
zaf8e05788af98434e002ee2b387ff05fd9b2629d07579e120746daa31660eeb72dd06a9d31b2b6
z5253d550f65bdd936ff80f3f60ce2417ac44ff98aa144f526a3439e37481c39846e433bdb146a4
z24f25b49265d2250ce138c5c139a43a0170a8feaf04cfe58182660054106655b0d76b503f976b3
zb3e537c1877daa1ad2a6bb1f8859abbb6ab785509b31831fa05983ac657a64b73e124939016c94
zf2068e6b84e1a2e5fad0fa9f5f07e3807ec8f6b358f1660cc6730fbce1a89565a073f425afc3bb
z1f798d24d2a0d776184f6e1097221aa9fbb614f246b366ce07e544b7e68b90d768827221973f5e
z407c2899db5145f5bfdfa2556edd3fd83a9cecdba3a46a3c2c15d3c97cc8deb09d9f112e6a0870
zf241450574ab5d9a096bf21ac5d7706b951dd3d4f5a8942f0a20d143169cd8fdbf721c7cd66c25
z776a064584b88ff535eacbcce9de48793793a1b5ac59730201a25bfe25b1522e6a2e3140a33322
z0a72cf225eefc9c86d2335c40b294e78ab3aa26cd59cffa51bbd485f749446a75bb78641fc9de4
ze3f99e70feead6c61afb8301b1cd5e11a607e74b956659d791b36dcb55691530449d252d014abb
z0f5e3e013246c8855994545448b8aacec760eddd9927d3ad039c8624288e842c6fe22ea95a6e8c
zbb51511486f8625ac10229300926098fadabe1ebdf4299883b89341fe7ed88daa82efb265e3f5a
z9d79f70005a468a4ed1cc8bda667d9008f835808bb0e9ad8c6fdd57e5c65973ed6644c9951d7d1
z212113dce683c1e3bc9e99a540bb4b1ce575de7df1c891d91d34581da26450f85fdfba826530d2
z345bdbbde39afac34cbd66866aaad8fb9eda02bad99477f1f6aab7ccc59879fa7124af383858c7
zcb1588070267e3fbf9152445a7644b0eaf88d456d136052c0673ff79d0d8cc6dcff6e1968d0551
zbda5314ca69eae36d9dd3d92aa76dd56a74a420836d5d190cc72cd098369ea1ba474f2389bacd3
z6d58f946e81121015fbbf5bfa1f92ec58eda6e9cc4a018578a829b54a75887ff79092642f490d4
z4609ee5877a9291df21dcc7ce372c430d0c86de17108c4d3dbb487e471f981eadeefbe7e7dad7c
zcb41b833b46b86d430562a8e36bd3b5c56f1cff8c93e88d2982cf5503088dce1b9bdc3004a548a
zc55154cbfbdabed9f5932f9452e227951ab5468319bf49bfe1bdfc39cf6510232e8553c8bdf6f5
z7b1663093185dd5d048288127da12b678377099f5003cf7e18c0def731b82a25ed9339d8d782a7
zf288bb6ced52f2aff544ee98e4bb138fea8653c6d03c0be44ea8e38db23ce7baad0ea3fec4b2e5
z8bc0f11cb62c431bee02b1e1de2c217c580e981f429dadd1d5fe31f562150c53d16f48e21f4315
z392994f2c884f2542730b3aba332a48fd97b8540f2261be5cfabbdcf18bab7e1a0d80f346b8eaa
z7551d7a5fbdc9d45fdb8528c05788ba1a7214b19f80f974126be390763789b5a90520a7dab5c38
zbcdab89fa9f951c04c5541fb453fbda694a1d952b0c5361796a408cb1d8cd155363364ec191237
z406b458d8326d29404a9d6056dbe314a5c9567c915ee9ebf3961943ae4b8a090c5be41bbc94b2b
z9c29058ade646e173286281b6f382bdd0f2a2051d45080d94340bd0c2da977c4bd7ab8b93efb24
ze12c7b5728e1da4b4243d834da674d86972f3421ea817e9ca72fc67c6eaa5b22e9cdd0cf22fc0a
ze64648cbf847dd3afcfb1ad0d3a70dcad5c6e4ffbadc053fdd367b69287042a8ca091abaf522eb
za1fc6adfa8902ec878994bf70df6c80bff1b48d85b764c4222553415e17d7274c8432e8500a0d4
z4131b4bef20be0ab6682d4bdc80ff45a66197617949366df32a80e56d938903bffbca5bb35db02
zc23f268cc6705c1de40631871443eb985ea54704a6ac05293429319e76ff01d93adb0f73c2092b
z5af3374fa63dca2e9047494d0ceccbeb739c23f35f039a30614321e8262046483bd2ebcaaaf76f
z2c6ba0d69cc56a9dfb7bfcf890521c24c99e1b3da7468abbd270efcc91ac60e1395ea18c1eda6f
z3d87ab1e96bc96e03bb2c3e10725665abed36244f53ec65097af83f543c7b42b22f21338d24d83
z5efa7902f13f35e472cc518673f4a8a034c4127984fe22723eeeffcc1f3c33e8da2a85f7f9d090
z125d4dc30ed828b220a6c55c67471309be609cec27cd1888ed0356f365c6b871760e1298da4a0c
z495971552f992a0b4c0807b31c86c7e06e96328ca662ff984eecab8f1b476ea69e8be915de9711
zfe6b71fc0250203398c4493e0a4232f96ae2dbb42b46c2842dd376759a2d1e58c522fa04cd8497
zc1ed916a097c4631acbf7f4a655be71618241c5311c25494b5aa88f1ed3541856aedf7ba1c0b5e
zd55c9bf05ece1dc3a6c514443fdebdf9acf42e92c9e4a7db80790bea3363a3b733532aad2dc3fa
z0d8b1ee795abdb18ecb2d65ba83ff75b0d4d0724ea8ec45d1a12a47b8735f773e0835ea89636b8
zf51f6da540fd5233b4ce9dd98c85df8118cd21120acb93eb64b5610bec4c17b42cef952fcf2f18
z0c293facee2bc63ad2a3bd74414cba6c0b4e1b5b8fea0e26738eb74d84de228df7f17ff49d9491
zf6e55e0d3024d9d496520b75fd00f8711908df40a53a55bf5f0ab9c09ed1c6657ea10e7c43a617
z615669ed589c4686cbde8d9aad208571c402a24b5fedf29b64a07c0174b1e4381a775735481088
z446beab8772b348cccc976cff22fc6cc5e34c7adb4cb6b9ffde2ecb303ef4f3806c512c21b3f8c
z98497bf68a82e10fd04ce9ad7a8d2461a09d8cb02e24cf3d270731a89feb5f9edccedb0df20a2d
zeea4fd7a1e0231d43c2b9ab2ed90726b496f1b7dd3910658bad86589466d560791fa75017a4b20
zb019ee3b7da43ac6a9c69f8a539f44a68778291176a4fcdf93f5b00f97e4497367ab81e4531174
z7f129a7f8097e6af49d672c943b7b554fa4c7847a522a2e0004bde0dbb5b402e71b42ee80d955a
z4d06f6924c8abf4c77b0a142c57265425d51a27ad164e53be98de1338d59387ae638754a1acf8a
zadceb93a28242bbccec8589758651beeb18943799d3de1bef569b626a3efa48769730a3cb45559
z0cd42a4b6176d453b7a252f064799632a86b66923e9ebf6d04af275051428ef2243e74c9311d7b
z13e5ebf5a54c0c456af484adaa0f252bed74bbcab213bbb15d7b185d722cde8a33b16413c9dbbb
z9825838b46fe000d27c976460afce9e222db5d0ce483fc8b6be02419fa09daa214be891b51a486
zc9f61f0d3e235a85f6f0523d8ad2ee823573d6bda44f4a1324c9f1108f360841799432976dbc20
z27b20e819b3d3ea1c54d057fd86da0c152b7e1bdd2a1a4ba231637550768810cd94d3d639c7239
z6648f25d843a891c76475de47b4a70b09f7ca43937c9d37eaa25206d10d4bdda08c7c828ad23fa
z7ebbf517d757d3842b015736ceccadfd8eace7ca3330f9a9d135dd170a9695d2ab6fa69c0d53e4
za4211899c2e3406affdb82fd45f5c4a05f7988777f9746bf7aa1e8378675816a3483a4ac1877c1
z6ed17ea9a70fe980b92717d271ec0fbff2d1d9b0999f54f959b6e1cba42fe0b49aa467741ace9e
zb1ce0d2d8bb4740e04a952fbdd48227a728c5b6394da9da5e48f1f06f6ee8a35d01932b0234efa
z630618f4fabc7757ef98ffb9f373ae0998fc82e00ff4d78b979885a0a01791807edeedacf594c1
z49696e43704a0dd89e94db2c5f8a70cc56dfea6c63456fc0ea866b6a6145e7d1fe11864d62ba43
zaf5de1d288eb65aedfbeda14c2f2614f5866c73deb174528c5df497bfd925d8a1fe458233553c6
z84c519b9f52361cee68e3fcc97ccd350955e1e276fc8cd8b074360e89246f3790e5cb215de6caf
zbbebddb7f3e173e8e2ae98d5ce769881ee02685545616695fce2240c0b451ecf4c4d5ab4418094
z28c7a7ecfeda27d1a55cf88e4e0f72f6c43c54aeccf7fd3092847d1db4907c2186b35d4f0db509
z0b47cbc898e13e49e6820ad90ea16e7f8d672ae9b8220d5d2a7e2dea8a956e187e798d821e80ad
z0d0e9e4205c8fee2a26cdce411dc64828bd1083b2c6e4d99a6db953c14259a0b6fc9f1d4331e74
z238a257766477bbf0b24da366b91f148d2f8c164d76ba146927434a1b7faf984b9f484ce8b3123
z8f9daba70d4be2c5ad63fac8ffed431e4923858c475ab5dee59013f1d440987e920436861678bb
z8929e99f30452cf4f1f1b7477576708f6645d3117a3d5f6bbab3f55493c82311be61729a20b797
zac3bd7a66c0a3c315d20760a99da6d1da3444d8c957a8337531f2a3eaec992d8c735c9be44c2a3
zd993b8c09f206c1a14160fb7eef14b2200f6ef7dca0662e58096d6f1ad0966c5dfb52a080b026c
z2d4da389bbae88c426c2c75c3a86149955a009423c1f321d85c815b8de98f7a5adca203bc7b669
zd0407c8d66400a2322b1a892d499ef63a76ec3b6a30efa5b64bb606b1a111cd5d67a277777f146
z77a2c008f70acff773f717255cbc0ca66e751e6b8dca864244c07606501109ba04e7e4a712cd3d
z37a019cfa6f4d1347423cb23c08e7232399b88eea6745c39a260a18dd45bd4cdbdb38cb4e6eecb
zc1e3d1918e90e5bdccf287ef2db1c772f31f407a4da5d5f120fde3e69fcaa939b126572982e26f
za4f2b4b11b186fdf91a9807a211d4db21e399c85445c23714c94c69641433aefc681a9cb041f42
z953f8793a15fe334d340e688cc18e95a342418fa22d0c9cd2f3eda8b803961fac8f8fb8fff88da
z2124b15b1746308dab334f90a69cd72c25260f4e0a01f99bf706b9a0ad059c8ea0d5c22e34c068
z0486b3069d8b56c3a1b76bd7b0058e818bf57b00006cc83b579fd47dac7e3937aabfe4de464ca9
z00941b38f66a4479f0b45cc5595c6d242f226808a8067645f9ad2f8305e3e666abccb9a040f7fc
z972714ebd51870f4128249e74304787518e3bd1e28866d3e4f587eaac1ed9161f26c8ed95aa602
zc081dde2319608a1d5a94f2c437a961a7e231b59b9e35233ad862024c652bcc9e31ec11ceecf6e
zc17af1924562263db6add458b4485bb3904779b9e358b18d38282c3928bebce3bcd161c1284fd9
z1c8916e60d7234adc57e1d17a61de972136bd4f614e48e9a49c54cf7a773f04b53f0d43b6c93b3
z8532a5bf7b871de7ef4d53439d80c99b2b3c4db3e06a6201fa69a1e60811b6b9bb9d0232bba6d1
z723de620ef705318a8d9e2e7bef14302031360ca187e7aedd654720bbe998ab9a6562681afb1b6
z4dc78fd3c5bbf7d8d4b3a1791b7b51129cd02fd6631775834aa24948e748a243f514f2f8564c63
z1fbe3b353ebbf83d0c17971cef586a577b0cc80539d803760ddfc95639121752bcfa1098155ec5
ze7090556fecb0f4df188a4bb112c7fe1575a58ac5a41b6877f792bd703ace9ac7e046c8064e3df
za41448c7d7a2cc7a3b2e440f2a438628d8c6010e0da342ab029e8561fea807d7bff64aaa63a272
z5461c74f3129e40521147f21818ba6c5f3949eeb991dc06407428572d4bc014076aac51021b3c5
zf14247480cd21f6b07794621c2902d7ff7d60fcf49a1750e15528bc8c187ad774a02b3738ec15c
z9ad4f075c829982d690dc59f85ee50c1a0ef1cb9c15841997f171520bd520e546fc0697cc3b381
zf593610d930bb839bf0cfce735e1bb2f07c50b5756c8ffb7b13801780a3c8bebbd34d824bd5545
z077b9247668f06119551365f53fe8f7af92b61966cf59aadc10e209d4b72d88da9b57be5aec679
z5d4e424dce2624280d6a37312429c80e8b806bb88f97aac4b3b92f4bcfb9eb785ad54bccfd24f8
zbd625b0406678d9eee04b5f2a42657722c1e1ef091b71e4c83ab2b5a2f276e3e1871b86abcbe6d
z1df53a876b327395bde6886d2f094fff47ac82edcdd5b5df629e90972cd08cfa0787d24da1230e
z49e4f010f708f055fa2ecdf2c122324d25d3d5d857497d26382a0ff22defbfd2633980f4c59c01
z2966ddc78b21fd0e551162fa8ecc7c076c890526994fbd40b65847e48f69c2f41bb0123ea5b4c5
zce9decd3b7ab3179ec6cc93955a99ce8db4e62c24bad0a2927236098cac944982be8301e5d113b
z07d1c56ef17f302cf032cdff0f9e3bb4219a519372b8edc9ad10adb1cf727951e62102475ae2f0
z67afda49b436846c3fde0e70604ca574bf7e7171df09367dc7a416dd7800d85c47ea38ec3ed237
zea87fcec842a3ea64d62825c07da5b4c3e53a0cea75c3c310ad1a9f5b844c58b365f8287729bde
zab5d72d63fd582bdd4d2d9f4cf0dc19493a9c91b2a7e3c43432b9fcbd91492ad17db30e5f5ef40
zb0089147f649732e969b5aaf17490afa8e935775948edf390df8348821554c1af279e0e4a678a3
zfb959e69895ad687eef461137f1babb8535cf76deaa398d65f4bd3cb41515c4954da8c5ee6232d
zb4925af017196c9b4942507007a9872658ab2cb4006be3119caa0377d54e565948d91902dc385c
z6d614b3e8be680fdcc0858dd4321bb67dedc9ae54daa057e80ac0a906f7b567d5ef2c604b40ffb
z9f54aefadf603110eca00096dff57501c2c1cfa194d846755906d7f2d4fe791a49603df7a78af1
zcee1ff7e66a9ac66bffc7c659249cdc6d41fee15e37fd0e42c06e426709dcc6d2265e829ea0211
ze01183a78c0d92e554a09720ccea3435cd459df8b7d2f3807837506c95482b9f12ef2bf73783a8
z6acb9e6874d9a22b700c386bb11e5d75467ec0490b639a9a5ea4ce6c46df76426dcea1d5d71c1b
z4d54db8e8fa6effcc32ce5f7bf65a2ee9eb29b3f22d650795db32a3160cc11808335ba76e6e798
z1d11d3412cd6a37c40974bab99c9befa7859fd5b62dbfd6efacd00d52ad1f3268c88d26fbfc5aa
zb46bc264734df98c3e13b4269db14f6af101b44496d293b31325b61c091c9037bc5c5b21b861d9
z4101daa639447ea6f8008dbbf15e48c8e8aab0f289d3729ea84c05bdae9c8e9921230206decf60
z542853aa660827c4e6bb531cfbd9ef5a49e7593cef7eca379c9bf059accb78c571308d9ecb82a2
z331aaef416082c8e246967245d31d917c2f57be9eba30a57e7a034d39a35fe0e61f8686a509b24
z351e76f8f634eb93a211f8e044f02911be1f56bd4a69e5cc96a70a96a994ae30795c73a60ec264
zdffebbd42a493bd47e9851a80b44203c61e53c909e3482608273d3cb4f00ebdf7a33562ccc6a78
z8c2a985eb9200e3e667baee7282d2a96a026ed287974d1a12e7b6373e2478895e058a141ff2314
z7590a8d2bb46429c8703ace6ffd5a89de8f8627c92f56ca9d0fcf6bbb57660c3c767b8b6f1d8bc
zaeb1a6d32c9bff8dce3087f7c35b7a70cb30b96e5acfb7ea2a8e2a2710174fb429964a7ac4306c
z7f1a0bdc1f8107d439faca9e02cd2b4234f0a114a10458b6141d169cc23ab17f20f5d237ba3e79
zf7ea9c5c7d1e29ce7b5516de61584d81187ffddb47260401f286b7c181adc40a86b2dd92f74908
z22638a18e83986399f9ca2826b82ff7106ff1870e6da1a52b869cffaa84d27b6b46b1c4e1f2002
zcd55d6e0099b1ed3cc0078f2fa48633440e6bda4036d84859189924c5b408b57afc0b448dfafe4
z23893a6efa998222fa943eb7c9144479b4a8bbc9042630038348bf9d36ff927344e3f8b0db9dcb
zcd1d01d65b36660df6a9e2778341e224ba7610c61cbc790e63e7a8ec39c6289465344f4b10b2d6
z31bc4adeb7265dba5d246c79875ff530686533342a064ac01ec9c7c0e89a7512891be8333283ec
zd54bcd5ee27355046be9d9fbce312377fc4a00ca5017988044ba911397f0eab7a3aa4c4ccbc7da
z4de5219305830e292bd036fd581cc97fae79cb26c67a36f24b4472db780c182b2504170a2543f4
z73434fd786ca65b992b7e784d5e0c76dd100ff55dbd06cb036d582f1dbf06d6c898f1981b23020
z6f65f7c18ccbce5b69e6fa0aeec43a450dfc50b9d9876dcfce250b7fcf9a9dd1e9cabd269a1e9d
z3de09d86decb8968f1288c9b40c18847fa716dd6338f42ccf835002f11e6e500bf52389c8ad8b1
z13f78448c7d3bc7a0f3eef66cf39bd5d375e5f9d67ba5637a01275fc5f42e9b0af671c358a6453
z21756a1497cc86e17c0cd1fcbcd0bb7bb6591b652a4302d6e3cecc23898a60ae0ad133c63ac43e
z8600f46d59a1f08231ba512a98f92751122695b88a8615decb045bedbdfc1261b9c8e7c0253df0
z45ef233780323c843ea653c85663b8af4fe9e068e24e7d0e51009daccbfc7dbb68b7a1d453a1f6
z928d7913320498a2cfaa6a038c23663274d8f791f087f3b5db2a8a5eff3a815851e3393067f6e2
z92793b7b31fe95d1264240efb98a3b8280737b608fc077a3b31fb08a2e089071775f17ca632e26
zda4872d3ae912a59c8136d4ab1d21755223aa209ff429a598dce77093c17ffd304e7774cfcb248
z3cf8012427408fdb752beeaeac772081c3e01fde10cd547cf42cc5ce83c18be7a61a2b59f451b3
zfbc4a916f06ff3ad3e15be417ad65440041bdbcb603d991393214403eb708ccdcda5c16adbabea
z76aa53c5972a0c2166623d4ba2946956afc5e0ae6738f94376b97fc8c848d2bc654278e7a99df0
zb412652a944120bfb40a93a4bb237a2a94e81755a9d8d2129e90d422a96a0df78c9c52719467a2
za614b4071d50fae07a54ec62d1a6039a0733afdbd5fea9aa66bdbda1e6204bdb6747c7870aa0e9
z98eb7ef067262292f21e993a53fa7e0bba2ffd4fb368958f6548fb0147009b7d352f50c9a399a6
ze43960ec6227b5757088979c0ab19fe83d39e4b7c34a8c60adc9d8835d7c3ba5f86f0e1d7f1cac
zb5eff296bb5d34c85c5c225590e5f19d7b870089620b7939c98b15bfc39ead28d3c176b1efdf52
z2ee9ce363b87b05aa84aa86ef57dde89ceda5fc4d45ca2b05ebfc399e27c963688350d4d1492db
za53d353e030d029b0242f15515a7ec7eb7e208a51964f570529d2efd3bbdc094c025e15bd0f56c
zc68b24ce18bbc82a9e620cb6be710278c2da726c3b1fa119885c8967b548bd78f25a02876d1612
z2fde1bfaa820331d665f62e1579ab928609e14f332e388418da582bfa60bc3edf4a983d602f4e4
zcd39efdf2ebdf9e6cfaf0fca958af7c3eb07774c6ee5fadbecf99fdc33ab1c974c84459d66be6d
zc13253ed3183e0a599594cd58c5063e49b6ed474dc2b09826d0b19da639451f41a8a4e8de3411d
za1c9a32fee02eab9f6e479bc17c9db0232ac21e547acb914549c7e65b863db80b03d63d2cb7a08
z311d49f28727fbea48cf2c27820b9a6145602b6c400d26870f28b2bee44c8c7fb7a14b48ef1edf
z263b52d8a9ce169ea6eaf70936397d48fff230bdf059f5efa2fbcc95add269870f0c17b475d5cc
z82819ea7d7b8cc8422354f919954105aaef159955d8c7a229f7423d29d544af49e8acc9e3769db
z3117ec3f98410f4c510439c4dfc7618cdcde6634af6d04f88c10a351df27ef84c7279e0c6ff8db
zac97b37ca71d26c2205b168e9813baee9e3bb1916102eebae35a4a872d2ddb26d514bd41172d21
z0d96f99b7fe43dfc4dad0313b16bc048c65b0cc95e2921f1a1d498a4c726d02813407f63694dbd
z17ad25109047b0a2585a712e66a12a861abc581d6f984a68ead7d9f73087a7c27a6c4ed3c5617d
z75a13b3449d5a728cf5d9a305e64b38f2934d5fc80c797a214f51d908c4321a596e47f5d3401c7
zfcb39718301d075bc5898150c1d94210618b11e3b996b9d7718fc34bde41fd425e8af37a53af65
z66fa545bdc4897e6e538275516bccaeddc1b00711e7b140a30c4725ddd62711d7be06f9dc6495e
z8ff0664207fe20eb552ad89722acfdf571747be48ffd20cb0abecc33ec89d8ae775154ae3680e5
z340bc4c0072ebf0252421881ee3d993a21add99fb618bfc561250f95cd8d6ac841744246a78dcf
zf3c89cd089dfee89e5bdc02fe33c5474591218abca27666ffbe83503241236652e97e8c074ded5
z513c9246d001b36a4ce6c3800d9711fcb954ede9f2c5a02bd37aa1352d8740bb138f2344c0b54f
z40bb6e362cd5dbeba4a24254aad0c1eee09f0e1d2c67666baa971bf6abf7d7b344a6f660bb872f
zb97211f6644b9236efe56015f0846a618b5662d2013c8040ecb49b17e5129fea3a3e270f1aa38f
zcec0c7e12a81c1248c04791ea6bf4851544ff2ab63abf6b4052a61afcd929da05934a57dc69c12
z59b2024ea5bc0b01c35a39b8458310342d1932978836fa06d62e6f158d842f169172366f07eecd
z1cd3c87c5ea4aca62c1eb85f44c8c9ec47040cf5620d8b2f589f6483bf68b718b2516d8127ce3e
zc5f6705cbfa6143d1f734c3060ca4087492434c95a9dbf50184ec7aac7f18c3f31e6a468b0cf1d
zda110fc172c7361b774ada8127cfe7c01bfb9d962ff335ab343134cef94989c14c24dc00b4d5ef
zf193411a5a9e99af243cfb7b98305fc95fa3b182557f677e46807f7f8c6a78fc96c314c20d0364
za6db9d114cd82dd812a654cdea2cacdf3234b6476f67db799c59b21c4d7410a9f0413ccf111c77
zb0a95b03096a4e5871eb3860910ab295c62f499dc25c09e7bdaee9206cd89e8716e35a73eb5239
z333f06a671258ef4833e3667bfec774303b7aebe0e311f6e221e7e85d1d7111f626a40cb79f94b
z69be25c08b45fb752f82f4b0f8a0c6fe820b22912c52387b13243598729ce5a02cf8a2bb39bc40
z210de1729a4fe0bf225634940e3fb82167af2d02a14a92d042c42466e5e3deab6efac65493fdfd
z20a0f5b7ec9b2c2270969d8034e8d4b5302de507438341b98f10ca1b9b92c61447bf378e85cbb9
z3992d231266d096e37dee76cdf31fca992416f7907c53a877ef5edac011a76ab800067fe80f078
z10a23e276705e1a672ebe6c083890a9194a808bff2e928acdf9485ede7bb10104f24480c602b99
z96d4fbc8f4c74dde25ce3a63383ce6cf1fc0da192a2483d79b796356016f2edc9fdf413f247e18
z6d8e4b7d0258377c0ac636c24490809fcf00619f3f1d410f531335a054b3f2de4b68efad87a02b
zcf028120d25e25c8047b357f0356d423772069b8c2ebf5de10b8983290949f578299eb74dfae50
z1a814c281503fc480d924b02e6959db590fdd47d4eb04930faa4d982d12b0ead61e2bc288780b7
z513d6e298503a792ce08aba8cf245f526aa536c6a5ab12ea9b22a76ba054557738936247766b15
ze08f659229d0a19c9e576cdf8a71172669131acec9d56d7d7b1122956453cbbcccb75ba3712dfa
ze48e3e9d131fc5fc176cd944364e0119998639fa674115c1fbd3287f75d0c9e84b947d777ad419
z417e63092219cde142dd11f64a723b0699feaa125d8d3414e14f5ab372b4f6d02c2757e35530ec
zb0e8d4d62df3503afbffac850fe94edf5a8d74d175938cdadc4473732ab3ef91997683a5e828f6
zf8dc9febe2137832c4794d11abf65821a2794672ca3581dea85521d7c577a2a01306df308fd83b
z9459f50a47162327f3f68603dbe7461da90c5934ce11a9c3299f4fd05fc1ba90ae0e5188306a37
z6bff5e9b970d4a878bdb3e4fd5fe1f6fe58fb75f8d41111dfafd45aba4e2cf60448c6510298313
zdcdbe49efef76d495c110e7962f9a9f1b07bbc3f44cd324e457063e943405e21233870de42d965
z10bd834fba716ce10ca56130f91fe2aad9729f41ee34d8a65d82b91116d011ca7b35eca5abdcf0
z2931b4da3b7f68bf7051c2a5aceaa78b36cb7e33f42a3e9fe7a0a3b93213ecddedde26e9ce05bb
z097f482cdf7fe7050310c2447b75e5eba8e627c90e930178ca008a4a1b5fe2bab20f08db44bf7f
zb6bf38ef9db48515ffe74f6d1ad3818a29dfd623cc23ad3cbc7a775b67d5e4cc03d109925cd5a0
z9ba3481a288f8a43ceea5f50ccb0fa525a2fa7a1d037430fb8a6b2f43c7d2ccf534e319e451daa
z4e1449e72068ce6e810b6b378dae7662b8f6cc9d44fe4d3d9d2268cf98e788eeac9377ef3372b1
zfcb6ee706a0388f0d6d707ed618eccb7ef08743f68a97de96418a4b5d7d01773dde972dde13413
zf9ded9a1caf99417ba29f2796db871c8916c45179aa7d353598d7914dfe030896086572f46cfdc
z8c3b5c481761f4850285558aa29feb9613deda5e366e85b102798e57b610c963c0d2d86e6e8074
z30973d808856aabc1fe0b634164ce462595f896930f555cfae2ebc2e4b3cb4431a79551965f48a
z470e45659ca1180137d785c0eb1d70ae062f1732e48f27a6c8f3ac12459ba167b38c27dd27f973
z827105609b454b823ed9dadc28e04b1eca5be2646608f8552226ceed9b50e2e374ef9c5d4da12a
z693c11bd5d8d7c6f851e1b9128d52a86c3f648620c9fcd45ce3a3950d9c1fe61d89b08e28b4f39
z5a5e5ecfc97c604df04f8caa549ea24339f612b8a929a6acef3739cde5e33266d83ae03789e1ce
za8c2af72042ea92a2d9cf99855164240776c0f7e8e06a696341917ba1e9779dfe634eaa2b6cc91
z0b6f12b8816e38340fb6ed566176ae6465e55007dcb483430b0aa84d15e9921eeb6af76eced303
z56ff8983c4b1615039506329fe84f447984b7d39d668628e1df573b53eed440775bdda534e4f91
z7a61abf1ea417349a0a6ee5290059ebe3e6f63e7a5f9a08cb2a8f4781e94059ee13566bedfda66
z5bfa86c6c13a90cbb9c0b97aff64992b7ac9075d046f1e55792c1286a05483c6e3dafdd9db26ff
z20bd46631cb5dbcc1b25c1d215c21aa9b27ffc62aec5607e6ae8cef2640ef77d5766bdef47318c
z2ce856bb5bea11a31cd18f0e791c833a33cc4a7b9a0afede943c7acadfcdda7ea3dac8e810b096
z6162327e050503ef654b486c5a4b7e4e4c707d0f0aad38ae26b6874bf829492e9507b1201240ad
z109f03d2d92bc76bb466886a867324fff7cecfc93d77ea5c4f561ad2cfe35e4195d2f145a91606
zd023842393275ec8284986df60dfaf2bf96176f91f14acc9ccafea4df89f742445fff31a15bcd0
z9ff121e513a46593f9d6e725becd1305dd08cdfbefc252ac01660b1c0f4d5dca00148ffdc0efb3
zac2785fd9de6d9693d20ee0558d09eafb3b550563864d8e1bd5335db2d0962758e688d28f692ca
z70c8a8b46a240c4ef5b101c9739fcb3614b48707dcebff881ba71a51493ca164c0aaf0c8bd840a
ze3a2de3246d39c4ea0efef06a2bc64e5f2086b148dc208589a41425a667bd57821db01139d4344
z3a33113487570db81fd8592cd065893e10bfd3ac8410ce30df209f416cb240ff689f48bff7fc43
z1ed8e83b4db361f8a8c480454a8cbe3033626a00684a2dcf5b8c6c6d0ecfa721c15be81bffc288
z03e8bdd86a39cf9f4b0e18813352b909462d91752e1c349438fe6e515fd3cb3d0713cfb0f57534
z1c30e36e0d33ff99c1842613e9bc8b676df446bec07b5d463d3c27514e7e1556b9705905aa7306
z1680bd2fb4288de43c358641d7f927965cedd229512b4a28d9af72140bb450e4c13100d30c0d7b
z66e69ec0f215907716ad73275ae096e005b04fd071bbc34b9bca2f06b70ab1d93345eb4145ae0e
zbc7158e9f055a3b9c64f2547a98afad679673f016a4b0b313cfb71638f0409db88c95b8b750d5d
zddde6aff9b9cd1c6590c4ea71bd3c05b698800e44aa75e4cf0de50d58e6427f39f6dbd980e17d1
za1324dce8ec9e0e9953793976a46ae08d0a756287e8d0accf68fa021598d600f5d2ee9b3f98787
z80baa6c5fdf67378d25454612302a29493541589ab87c82e0d933bdd12ac36a199793a08d11fc6
ze415565b820fba44172210bbd1a31520c41f62233718e126db39c7b47fcc391ac14d439fb398e8
zb5ed63ecf2777160dfa3f40866493a1b1f5767cf7560883f8844b9dd4a68b3c3566c4ceef7d642
ze431fbf9ffb09b2a26c6363dd003254f522820f13a8905ef37a613b3fb6043e070d9f526f01876
z1082cd805cb4a98a50928a39d9bd6fbe7b42ea78150486dca246d9728c03f12210cf1d86beed5a
z3691169212170d302ee4195b35c702beeb6ff8c3f36fbb76a109b3914c5e633e953adc20133016
z9817a80fa8046bd081d5a5ae378f77a37a82ebe38cf359ef641c2efb3fdaf4b0ac44935637efbe
z63595ea96dce0463e2294463ad605ad260de3afbcdcbeeb9f4985ef5329823bd7cec613f651ed7
zc927dc60a34b58fe91cc23ce4843c49ca3724eb850a70af6f1b0d1095c3200fe8581b87d4f122c
z9d06f88a6a84886a142ba51d01fd61b45241a0fd98a248b3b4612989a93b90f8106cbe07944cd6
z2b7c4ec31d2ffdb39116ec3ea7795cf9bd1457d4e4ddfb81be53c49152e95251a1ef60d7201d0f
z8ae062a2fee52efdd3dacedc0d2668383d6e81552e4afcf424ad595bfb5bf0d08002fb9582fcb3
z6bd076251004aad04fad6a1f52dc83cb67b004421bae40602c10fa87955f06d24eb509db48090e
z2badbdd1e41d13f046a43357452ea3e87b1d2a630d8e81091ab6c1926e479d86077d4bfa5b314c
z3a4919c0be39ef110a9d33944aa62a56b5fa843504f4a7a35944a4789cee6462eb096447b82b08
z5998d3e7be7aa0e6f6aecb483973f25bddcbb08c7f6b7ddd06db58fbf3c674329e782b199ee246
z0525467bc8618480464dc8cf75d4f5fd426adff7b102048c69bfa37558f8d8bd1e71558eb42926
z8a76e6d4b5ce5574c66f72fc602aca39e2a7b1a5590c3ec145e337f1e96893ed3ecc0df5ac23b8
zb5d19a33282e4f026f7c688b4d66097a4d57d7177bc71622e78638ec96336c80c404bde475f5d1
zc5f513aaee67d263aa76cc7954e33049f3f81cccdfa2a5fc52eda919c4467f36a6eea08d81d2f4
zfc005ee2804a0d1b2a12d05248b1d7c68d6566d767ff7042a7327bb0dfce83570f206a23269cef
z3a2667e73ce9aa069a0afbab065f4febb0fe841e3277c5007071eb7352b20db4a0377bbe6311dc
z2d9f12c4a6820cfa6e7f62ea96ed38fed8e21dc3fe976840ae28cbd406c8f14483d68ddcacff4d
z389e713944e387bc06090ffa2826910795968ae3458f7d45dbf40e441afbd921e1e71d7e687a7f
z36a5353af0a2a2557a7a5f059d37bc21433d9638a11a68e508591f33352b70fb132a751b55d0c9
z22e0cdab9fc7e7ac9bfb2f288d3490c8763c8eee12b68899e7b4c1a219860d3efcfc97e7d24cc8
z41aae6cd58849058e12238051e8cf8ac6ae489730add67986ec6fcea2bc805a1b18408d91a7100
zc81a136fd9174deafdb6cde803752b7b9cf5993b104d29765d0d83138d80a75dca2cc308d10601
zd052db646a8dc63a550b1f92862f6731cac9445bec54cc790e85baba0b52aabdd66118b4dcf7f5
z61a8235fbb89373e2717854d8fcf26fb7bf3328b818f422659f8b29ea34a91a00de59f1c66c9c8
z67e4711ca4c80b129092fb6226668d4023d5c70a0bfec28a0ca497215dbc02de82949d6acba35d
z193189734030511305a05c5b4616ada665eea859578c19fa2b95651c7005c9d14b9116491394dd
z1e4af7d4f772f9687c8b82f096c106f9599ae2e4a9850c1bc0cede63ba306707c84f73851af8a9
z4d241a9e0b21f55a1137795d5dc3f8feb8230c032fbd2e842f8842b419a2859574c84074b9577b
zc5a5386b5f226b6738cc6eb62a7ea08f80a9fb32d3dceded60f5dc1fd11a9cc2599e778f052369
z1ec909cb0275eb47ae0e9cd06f072af2bb6b89581c0ccc7e17e5fed09d3298612afad1caec4042
z95744f81adecce183b330f578a7d20ac4c2fee39d9b3e0eee88ec9537e4c58b7bf34fa1e904059
z9be26394f0c55e308c64c675404b88dea34067e377a5fa6224e55fc2cc5b65471ba7332a587822
z26f2197bd09b8efd352d96c96074445b74acace092e606839c12ac8889330227c0d2395963d4e9
ze6065f27ddeb5b3fc9ec9a0c6de9b0ad2dc9fe6da1bc3bd902e781f97ae11303a08cf418130d26
z87d5404d82ea77499f463a927a3ed2d34320dab944ac17b0e490bc3841dd7a1619923f06ca4223
z9bbbed03371de65b28d98ca08b008ae32cacacce5c67cf60e7899ed3ada457d38faa2bc653dcd8
z7fb66ca79784850dff06f87adf416b8657544660bafdcb21b4dcdf40f795a1eac161db286a0940
z7f1838d7ed0d00d48ba0c53dbb82ad561488b7068a6262b19804d2850584577d7f1a5ce87fa117
z69df27c94bec8a4a4d38f313780928e8fb0991e93a381912124894df7f4126666e6885d01cb30c
z3ae502ac6c8a7ba6e7c1d6be1ad9f0210f78ccc872d7f64c64569daa6061376b81d2f4286a7900
z72fd33fda89f7c28c7cac582f80053706776c6afe8f79545807c1797ade3d71312bceddd823cea
zb05624382cca836349a026c99a7ab4ed0e81aae11befe99a900b44bbfb5259699992bd132183c9
za16eb8b1500028d3a9aa46ce8bcb5ab562d573f1532aa3aa3f345ee30e2751f23d33d6a930a839
ze3a5e1e84a5e2a07a49071a9c6cdf68b5a7a077c0e49235f28142d7d099f84511f1c191943428f
z835eb70ad396b08040560b895304118c51fefff580a8aa7609c74ed2ba91ce9e314b29bf813f30
zd1b3c36b40b59b6bcc74eee72ce3592b327604538e87a68f79002387c19ca250948fe200f6f35a
zd82c6504b86746dd71f1cd13d1509d2fbbeb88835618d436576becac749bf26d86e358b4b56e63
zedd47e4ec1298aadf70c0fa0dcb2c717d00888b6ed04d6bc4bd321b12058e0f64760f822ab74e9
zdd2ba933c81153806a91e776ca4742c5ee0b85c01ba9236e17c70e5c36dd0018496f9af3d1b233
z86c93041a3a8e5d68b08d2cb26206fe0fc131b18b65a54865c0ae3c722bec70c95a6989c346fec
zc09826648d227585c67f5058584185caa3c7040ba76e8b46ca0b0177b0251c6c1d9ae94e029243
z3c7096e86e8ee2a99e301eef50a926a20dbc5c695bceb14a61453875dd0390cb19abeadcb178b3
zf544d6d81b076557b8fc3e797b5de727681b9595b04d8780c49f011ed62ffa4d9e1ade704c06f6
zeb55eb85c25cb1c2fdac5347fd0a9505ddfc664a32bd76d87bacf195c15d9f4ee1309f87f39086
zc30ebd3208359ec833a32fb9bedb3a6fd7e3d92b2b209e5cdb0e927f33ccf3aa1e07ef3d15d6a7
z88e0f9a5d65742060208cf512ea6bc1c06caa6909d0ef51ffb68de7923b8bc7008bda708c5da88
z3958aba816b74503026f184f7e862441aa1040cf340660efd16ee0002ef02ba85062b2cb24ca9c
z735f26c9baa4a7a70d02b045b5bcf45e99e512821daf824814ef4375b27271224b19337a411e4e
z8f15cd1cc79cf979cf079cd454620fa245dfadb8536939b1e41dd0013cd126972566badd54e9a0
z80fe632098a6db92c406a072600a6c8a3a52ccdbdc7eefd119759d52875899bdfa5c93c6568cea
z263c2cc5ab0b2fa21c5586f7dc1c1b06372a15ca5370a2f99ce316e09ef04d8510026b4a410d24
zba9041d84dd03826886afff800779cd57b33941bf35c0f2a4aa34fa5d9adec3c48e9d68d5d87de
ze8ff0071384607cf0c38be5dadb5bc6a43d13034264d4de66664dbb948b8ee234632aad8bc2e6f
z0aa363f9691231d6e24b2b938756c923fd498b250f30f0ea41518149d7ab50316f2d71235f9442
z8e8f760b73d1983c1ce8ca56b9acf32393bf92f99f8338bc0a24e7acf0a1798c6228a20ce92cd9
z759fff494c93d29f72c671d2d0ddd602c359ec4241543ac4d70cadb6e37f959f9cb1f550853d92
zecbf57d5c11d23a0ab7c242ef95db4505b13fb7dd657a0b98477903d6c6d2cdfdce86edd0ac57f
z645ce21d5f39c48e948158a58b067304c79412aa49da355a1a9d776dbbeba2678f885958947f0d
z8a435923b3c29ba2e0a38ac0938dcb7cd5d0539b428f2a45b48a20e2abfea7fca51e7296da60f4
z5da3772d9d899b3e47afecbf5aa2e60302f6f39630794fdeb2d3471159e25ecc839f0fe29c2206
za0c70e5e264496c3684c6af784dc9ffdc1951462f0e70b8ddbd3c27bc848cf9092aa53cfcc49fa
z7e255722f4efa764c33b8070856d3c126b961851d89c32c7e7c5dbad4a38661f7f94b3db23a4ef
z1da0c3428e181e03fe0ca54897bf4a005f20f7dbb5f14a1fd0b1293e3b6692320f68c6f75c2a27
z659604e20c50b30e10aa99871f5ec261652563951c18b10e182d67bd692ac6586e3d6668f56d1e
z53c96a371e2ab744c7f1bb5d5b96c78d73c1f5b18e856e10637ffebc1b00827cdfaaaa4089c9aa
ze081a3f09e2bcfd858da70d973d7e50fad1e705b61715bceb5d0971874badad08af8212104abb6
zd789586839b7b85ac79b29791d00b69821e9530dba89474f689410f44b9ec3eee90f4798b84556
z6efc7e36e44dffefe71bdb19da40b2102c3d7c70d8b510b01e3b69081a69b7887a5cbcb680a8b5
zb3e8c60fe7a3771c360b44dea8b91a5992c5bb7605056ddabb9eafa0e07f091c02c15d3a145d94
z297975e33a89efd74de7eeba5e2d151dc97da0a5da36a8a0cc1e0046b11aceb7ff6b31fbf95c4d
zbcc6e2d7cf4c8300a942d7f8a531e8e4dfc6a88f03d5b298ff1681316474dc8ed8797977470570
z9a8906d63b8bfb3cfaa5b0ba5a35845cbc8229a4ac16a422ec57551ebb237600541eea67d3f61a
ze872a0ac0bec075f3ce18b981a7ab33924bcbf32addc732e71a7ba35f9adb4ce112e74245b1003
zadf5e644b52de64c0afdc811323eb81882f28945fac3d3510b665781867070e8a890c576f626d7
z68fda2082b9b587fced7cce5dcbf88fec60b92db59664f603759c10bb3226a606cadee19f597ef
z1c03f2d82396111eb1a4e6b29d222ec365c03645c1dd7db561503ce5fb738f9f8a9a0442d77f8c
z3f901a3d043f9fadbbb3b173975c491c940ba9505a7dad71908e427b5eb6ce5a001a23c79c1dcd
z0b4683ef35ebe2ae4ec4ba1664fab548194f476a817f068eed97a203b087694e90f3a5d140f5e0
zb36bdb7ad978f39c1f7db461a6262fe9996c01ef2950353e5f587369400cc79dbb3a68516ba1bb
zee8406f873574b589abbd39be9e7118be11ce7347900f681111d4b53228e5487b30531dbc0e51e
z7b62856302c4b6ce347f2b169a5b452f4212343693e38c1ba635af765a14402759169062c81a57
z1b9b222eef96dfac9d636b6a8909ba1e1cc50f3b91908cd1b8ef6b2470a2369ec4e07e88cc8f96
z263445d565450a2cf4dc71f147aabec784122a218ea6418b8b6158c6fe0fb7df0db32c49f7da56
zb1cdd1cf75f1efb5cd0a907884c76bf80f225e83fab79ef4476b7963063dce69173f42eb8b2fc7
ze80ea68e076aee1a76f1a3d141e5a7636d72211cd918a40aa586823d46d957e08b54db4e436c6a
za6c93ca3cba929e8d0ff68b32b125c4f96a60fc98d22a62cafba29439e87877e9e04c931f0fffe
z97f30c0cbf8c5e344c6e6c6a4115e807b884d355bd9054793dc8912690bf32e4627a9b7a194f43
z2d0c1ad6c809f4f46fe267481e44139697c81f762272b0e08e8b41b42373352d774e9f59dd1d34
z60d99583cf0e413390759970b99c2afbd8b9aed008e06d681dc16c6c701af95c5c682c49d7f071
zfdec3c1737447903e20ba1926d1710929c304dc4b815f7a9080c2a4fe2cb85c631ac5f6ef1eeb5
z84704ceec7cf1dcf1ac3b3ed4852d82bef936f1084dbef2f51d6fcec8efc43a4520a2a0e876641
z81d4c09429527f8b54bd010d0d889ffa9354d45e2ee1a1dbdcb48511a642c1eedb34794f551313
zea4b7b91f70120a3f83be535dd4b5c8c334595b31a2ff9bea3a4f1f2557210591f1da6df59692e
z5ea7db522c258a79b49a1687239b41cb28c3279b48c844375ec633b7bfcaa9712dc27cb12c26b0
z274f898144dc687d1c46524ce96b3b600c5460c6f4bb182bd4ab6711952741d01ac612b8f5e16d
zd9cece7fc99e8a304817961a83709e03b9c4ce5a82129afdacf5bcd6139c4da31b5ccd9c803a2a
z9428cb2ec4d3191d619da53814fd4fac973dd2719634c304d8e18fc949fe30de94b8978c7f7caf
z27dd42eb1b61ff1d7fadfdda3afd2d418209bb2e2a816c127def54c345f8dfc4540ef0342888e0
ze42975bc0fa1cc728bf245bb3f4d311306aa97d21b2831d89178725f9abf32754abb3755c6b362
zbc6dee6d04242bc354cd4cbaf63e17a39daecee548bfa11fe58cc3666c4546b103be4f114429b3
zddb54eebf1263be5206eff081f14b0bf22f678ea8f9ec553a90cc4f5076ec969b1d8d70226b470
zf98dc692eb663ae3f6c62133e581370455a4d420522040c79412b1afefd383616980ac62f9bad8
zd5496e9961b03c6c9074416ffdb4013a648f7bf367ceafea82c16001d5f88083f4e91f3f5b917b
zd5f3c29d374a2cd22f9eb48ceeaa91d03d4a9c826cf7b376e2e92bbb7f3cfe9c59001de4a7eeb6
z1f3a24c15bd2cb7933c00ce970e8e50d981d56c95315e3c57c35a45ee8261183b66ec2e3236518
z4b60857e8d945aba9db23283e678a7f28be3b91820e4d19e2c043e2aede96987ea8f188b6906f1
z6cec2baee28c392f1abca85ee2b3a54067b946e3254cc6e6b315d0ac97641ef5522ae27b81a0a5
zdb5102ae6459992b3eea6f72dfac890b63a8eb90c42b8739fb8dee7a8d7e1e175f84eefb33a301
z8b70c28ff31bc6d25366a28f0b75666a3db9899e3afdd0b580f75da183538d3c6b27bb54dc58c2
z7e75d570484146e01b88080a9feaa150aa6e2e72b0830d101d555a776164fab5df31e289d51b24
z2d52f7d36c128345d8ca6b3a8864b14a3ab07fd6a001cfd14cffa957a7c28a279be208fa506d61
za0c2a2d376717197e568891212765bd41670a572d5685d823df09e08a6ec7c3d428e492c0a24aa
z0a6ecfe452c509c5c76e19f5500c230d42a10e10d32473f958700f2c4d5c05422033560a1f7edc
z4220f718a044657e9337adf014a2ea397ab2735d73cb9a5f9f2de024b24966003a555b9d895432
z95866dd199a70f5d674a2afd5c4479e69c5d2ae59a3d84268de5630f1238a17e9115bfddd53bbf
z91ff17a2ea21da15b6514457fc9adcedf496faae6b32d22ab34ab6570704c84e3cdf0d3da9134a
z569d791e9df2b1ae695a42b5fcf5fc95bca6c5483c7983aa7e5a7ad1073dbaf1cc83798c056224
z7701218c844f62e5a349d1bf9f077521da956d623584b75d01897890d61a9edc179d57b01a8fc6
z21fda781d5401025de2e963fda53a296825a18d9a119fdba6767bbe9e90a74e139f929e0f55bcd
z4ba3f50335418b6ab6758ee9d1680bd36ff6293777a163697825b4c3dd53202971f9b2590bcfe4
zd09e034208c91855f2fefe5502a4e4a64572d3ed67ad933a4ae14794b656e18bb82f9c99526308
zd369ae6869e5929df970fa40e16839c65df2555f68908c87ffa3817af832f7f44101878cbc51fe
z377fdc0dccb8c0ffddcdcb2de4318c7582cd73e1f0f377ced5b97b3b341ac15db69e0c826b8665
z081965ca3c4105d0ab6b62790529f9ce6b173ea1b016eb4727d2db7a5a4dc07b888155070bd67f
z46a309a684c232b520788683e8666fb09f9567440a104037cdfabf296eacaf745a7af2c1aa6fe6
z5592239e4b923d0d7f72ecae75fb5f936c869c99df92e5646699fb86bc242e69adc4c6d7c881f1
z872da7ae450776f1bb1bc90fe97944d325518743eef40fc7a9c42612785308e5c7dbbcb6e3c775
z338d6755f4041c5fb2c3920b69e0d36e84509afb15b3df38502263464ba1d717663e4cb8f91786
z4adfd1edc6f6a91a9dd9a5800a9f680e194d3159e69fc3ce39e047e9943536e09846da6fd9cf70
z9b0805fa28590530cf6c2d13add9d9a144d2c66807e9918b3f555d884e2ffdbd2d7d20bf22692a
zee5c9e9dc5ab6b76a864aab78d90c95e7b2e227d5b8bb64fe3a3dad118ed9a26ddd74d0d488de3
z5a5c4509d7ea0a9d5e2fd8221e55a730a583f907dc1ec208dfba6c12c956cd7cf5f5ddc144c42f
z2978934993e8e22cd2a0cb95de6dfb83866830d95ba0bce2c1349bb4f772e36fa84b02c142970d
z6cd649f4e443f2d0056fb25beccc302dffc0b83fd57e39a8ef87c04548e34f253c368dc2c9cb24
z067541829c3b5d92a86e88ccf51925bf20be95c35cc495741ac1727a673180a70f47e0611c531c
zf393447371639391febf717c7cead992a0f61e254658e23d741b046d58b34bdba30e48e9916a85
z1a24e83c4a7a24ce4238f237d619df3f9f51ad3ccff4769b142c9a7d9808c8e9392c3f69234126
z0b13ac2d5464464e89e1d8ce128f97df8d42de3a7ccac65414455a864c0fbbed5b5b9a7d7a9264
z5573aa73a9bd264c627b2a6f030139488e03e6eddf3f9ea5f2c3bc59b1fa31eb0b751224e6c649
zd2a656b6fcb8f987dbdd2cc1c357ed396070baea9bf4be350304e66ca4d0aae000506a7ddf2630
z3229f62083fb4f0e45789a40ef036a321bfcbd1ea4a76a4cba48c9117dc4d7241cbd9259f745de
zc97d4aa099e446ba09c68f01ef2763e6d86aeb33aa602739b408880a4b582d48d47866c937a0dd
z7729c7c3e788700e4f949602d42c6fd2d769811f209eeb9f4d9b5c961573b4cf94411ce60c3f54
z2f7999253190bbc5619a920cb8a35f0e3977f1075ccd5443c2ff8589202e3f9ce394a5285184c2
zba275c4fc3dc07352dc6a4918bf74cc1a474ea257f20bdc6f689cd524a1290a6bd0ed0aec2b175
z0efd354f8f4d26a93abdad0ff27a7b8d13e2a825f136a7e2f5eea8aadf33b27dc9df25a86e4731
za678a2b7dcef8ce2be296b70a6b0e153ecdf13e2e0ef06e552d7484adf2f9b74567e43ca874d73
ze0a60b98c4787f721610142285d350de94ede271d1d187199771d3be80467be5cba6c1f20687d8
z3ec49ae4973f4c71f1b6fa59b06fcae32f6dd5eecf7fbe840526c4cbc329247bfa160db4f9c96b
zd9e68820b855a39899701ab232b7ebaf76d09cf3850d9b1e3177ba9abced19e010186c3b66f573
z14202c699e9cc5d1b916184d0e23d27287406dacde8684834ab8732199c10f1d7cf3038cadce18
z7bf7e0782c1a99f3cf2d28ecbf735f1b435ae015119dde721266bd6cb05835d8648a9b91625949
z3eeb1642d018e920b2a1847987230aa2c73c797686ad2059d7d66e2c6127ff98affd1fbe71dcd4
zb6b3185e2c308bc85b6020f6ff7296ece5caa9150d9f1656d885c866e176ea028adb971ff2fc2d
z1d3992fe206a384e6ebc0df4197e0c502d4f9712979cba0261e33a3766c7351eef9311e86b5b26
zce464b083db4e47c9b902994d55982dd265e9eed199c09710817cb544c80e9c0249d341402ef0d
zd4e30d7a11d3a781d47ef627caa553833969de2b1ec30eb5ae42852760f768a83e0461de471acb
za5ee66634b1bf0d7ca05bfea3423bf709712797794557ccd6fd8dfd145a2e13573030d8d5f1557
zd0ec0a78740e21b6e2f4d29d810d5056539ebb0ed43e0b74c4e7a4c12a6ddf9e8c402edcfbc759
z708e2219cd38d2fc358bb4adb0b5e9cb071e5f33780024cf0e96a87518dafbb9d0f5912c71b2a0
z252800cd0f17f8ca82ff978c76d61349786827a52b3f3e98b45c645afe8d7faf2c4f9a97603dd7
zb62a98ff31825fe6ce027b3cbde200838924a155b97ec9931e4ce9e1ebe7fb3598ff6deaa36d0d
z5b435741d90af6e6f2a04ecbf6889a4c58bdc01417e24b21e456cbd9d1fa1f8b043e8f2d018c78
z9f1306e405ebc23b6610c5565dda94dc2b3b4bd10378cca8d02acf30575ff6d0a92e2d07bf34dc
z8f158ae2bbf8a2dee97f49a4377bb8e2cced413168c59c2dbf657fdcb2629bd2909b744790fb15
zd37572175a88a8360fefddaf62f668232b053a2a82ea4f45a897904d938e4fe2ae33dcdeed876a
zcd6296e90c380939bd9f931b26b843bd292176a1d0d26386bf1cc09a1f1475777ad26c26f10bca
zee12d8fbb8e3a9aed0b8d9d81a378cdcef2e6bc8dc9a2685714dc55e07c697d89c4ebab28adb38
z02149f650586b6cc65196f9f65ee929df50a6fc3fe3220fcc78d8e7f51c507ee3e2687021b0e15
zee95786853ae8de776b8f7ea65d9adaa5d800226a943e2ae8deeab89709d971db09ec289cd8a24
ze4c1d8feee4321b747032f7df5ce0338381c72bc41c055d4000f3ada1eca6e70d600b46d45253b
z8e2ee2029e8bd7d1e9890fb7ef2c475e19dddac1a3837404378d48edc1f9c2bb1e0a10e8257482
zcf8f15b85ec2fb22a86e873e6fa549359ab33194d17f0dca5779a08440687660c6d545cde2f58b
z5c3f7844cd1fd679a20823370dfb8dcc00e5ad5a081dcca8003cf7da01a30ba00088d7aac06b65
z7424f57d204f6d4b0b074763e9fe257ef956d7af6e70086054d49e07ae7f7bc1849ecdc2f1b319
z22b511a3aae238f03d9e6f586017b9dfefd98b7bd7a1404ffa551b89622fd707e5e74474bd2a0f
zdf048a5dd96fc72ebe05a1629c0c8e9199d9c0904d2410f3fb71d4ef75080f9e3bdae469786463
z567bfddfdf82199722ddaf079294935f5ae65033b4100eb0f26c5f8e32b762784a1d387937c404
zcd968aea34e682f6a74040a62c9a206cafe63bb6af46b39fe488940b52bcbed78dba5d17572a53
zf1369085e7059bddc7deed095991b3afb1b1ffd70305e5d450c63411e73b6ab9478796936c9467
z4f488f9b66aa82c26027dd8fcf0bacafd6c4cb222c1a4c14f1b17ccb320cf455dc27fe7f8678fc
ze0c21e6b7b9ad2907e66784f50c9a8912dfffd8f4e44a5131698daa879807e844173bd665c591f
zce90d57cb81d32640295271adfa48fab8df4b1a94b8acdaa95910d570a5e2336de513c5b911410
zb7b688ef3afcd913f36e60563365a40cbc9bd96b7dadebad4feff135e9cc22dfe5089110d1db7a
z3baf0fce921ff5097f18c061aafca31fd256f345698043406f49eda1c6d7fc17219b7c693c9d8b
z183d5d73845e6ca8e3be2eae38a6f192eda88093c1675855f2c6d1cc88439da1ad07f3784d6e5d
z40497f7d6e008b8986007d441defcc996a1e6ae857b99e08cd4568fda5d691358bc9d6ac923b1e
z9ef3c59708ab9d90410cd225552112937f0d383cbf12e0326e48abbd4a4263295a96f087a0bafd
zefb6e46f5989694d1df3bd05440423eb3286847757479bb4177b3cdfffde85bf70be5d2dfd63d1
z33df209f27ba40b4c53787c290b374bde62eac1842f44654b91f45a79d56484f67bf1e508b656d
z916777148a7cb5eca44198e5db9b89a7ee7776c93e4a952c0d08b2a7cd095c10382ef399e4c305
za1629b30e7b8fe730a3a54f0376025e5a54821d2e18d3d5727827da0f5c714464a0b264c16b672
ze58e7df3f604ef8212fd7caf0782407e079577c9d6f3f462ce7f9985008e16ec0e9972cfc037c7
z4b45c3951ced8af03aca4cd1139770c70b742fc22736b2d53c714421528c9e163dc5bfc3c6d37e
zb7be1567eafa0d113f3e0d2c4e1b7002c4f281f8c5a6207e008455d67fc593ec226c2f5e9f1739
z29e350a183a20e5468795049538fb693c36019857b34a0a1484b9f183507a85700224617b7734b
z9f7465a4eef5983298984036c7e3ee2bf806241fe18ba15f0b2ea1ea6ee16ea81d0ef3360157c0
z0749aa8deccb1e3613d7848ef425569c06fd637b54d74a03e34ca034ea21d0d531b030fac6af6f
z78b08f7395a6b661414e6bd4c025e27f2ad279f34db026ac9f3d3057f4ed2b34c168a76e636989
z823baa7551d1183662a5c2fe215852f488486b0c054350366b7357f83dbb266da6ea437397546f
za074d23a371217d9e8110b7055fc6e1bff12bd7ad384a9dbb4584cf8cbb330a2f6444f9196bed0
z2fee41e48bdcc405ad837b892d5c30dd8062ed55bff5858324ee8770545505dc64874933231392
zc6a63fc708854928949bdd478edd3bdf60cc304fee184095aa70d27955393f84ad73fad0c1d747
z9a7830e7e6f93cde421176361ac4efa0ece5db39ad141c41e9b69312b566144fa68f008c84e940
z29c50d426d7d3ea0dc988af5d0510bd44a562f35775ed948d6ad911683ded15dc86977fa559898
z492865ec8d6f19c284140ceb0d7e4158f756a76cb6f5fceb35498e9029c753b62e815d7423cc54
z5e2ff6c1f99885cde0bc25c13eadeabd59738987020420bfe5e390fdb98dd1f6fca026b0f81720
zb5dd89e867279b8c47329f2b5a0aa72e9300eb3aaa0b47443c5f69f62eb45f84a7253463404f8d
ze45f5c14b24e8567ad9b34e1b5016f2370ed4b327157483ab3d383b810675571467dc13200ebca
z8e3b573e5303abe801bf5ded5ebc71d2427591b584724ba8f94b1b504418244a83798d167ca6ab
zea80c5f7a504d792748446de2320bdf097d61d81fc2216370021d239fdaf2cb1f5df02cedd5372
z28561716717408bd570dbc90ee5526498a08eb626bbf2c41ffabcb5db85e21dc4f50abdad4262c
zcd40a0bc2ce0c99f3b9581484e03bd361308564c04d19dcfd8c5a4c96d614caf5ac8acd6c12d11
z6a3b04dfa1a1ae9e0a3858a6d110bbb9411fccedc99d3c812305eb3abcc513802ee2e4f9a51a5a
zfdabf0ee4ad8387a76e18af941161c0d931f25f489f62ead42a64b7fccaaf530f6d77d42977c81
z6841e17cef5a9a158a568d68e2e870c22c79becbebb12a667ad8be283e7d947bb47c92d6b1a6ee
z3bc4ba40a98531f65a7d1348f31347bc0557b730f6009e26d7c511142c3f0f0fbf5a0eebb0f749
z267259d088db33a3de605ccd9c482b947ef7e9647890831fc4aefa2e92a94ce291e54be0d2abba
zd33e866db1cecc397281fdcca4b22597f960f5b490982d954b99d84cea5ad7a3abd1ff0f7228dc
zca50607110cdf3176dadbeed009c6947885e48a10824701e724b3093be724afd00cacc7b747343
zd594eaa3587f1bf6ad49e05c709727c4f136c8d07cd7e003a09f91da18d2687d1f78143ec5db20
z96c62d8b62142738ccb4568ffa9e251d29d24dadf7567286f13361a6c6d386041495dadfcb2f3b
za1d654327aa96f413cf524941154ce0d22203cf1ec043348a08c30c24a718ee2e5628ad1f45398
z8eeb04cf13441634cce6c76eceb34e9ad971abdf7bc96f539d7b5c7d317f6dd878da3b7c1107ac
z1b84a45544557db5048db4ebcca38068de48193ee46788430af12e4957526d77bcc1f5d1a3033f
zbbedf10f67f259b197c96cbf304e75fc7f7302c1e4184f2e613e720e21d095f11c3841de28a4db
z79f6e18b1a5801ef2c71f4305e5d488e2464ba9117dc54db8cc95fd07818a4d193fd9a70eefd10
zb846eb015b7a745a654d1b75ec530f60ff029f773e7244328c6edcfc99257138bd2474fe88a7be
z8c5ced1b64b18b10a08c1c821512adf8c3eb9546416fa4f73cea93b862e5de46a271aa4ecf6e1e
za117e087e3bcb0ad0990c763785e4f763e0ebf9dcb710f3cfdce9c0f0327820fa9596872662cad
z34acc5803ba2c9842012bc639500f1e514d3256c1b31fcfe3d3326a194f4c599b40a098eb6e482
z8719fc2d7ffce358a9fc3f0bd9f13e9b2bc78bdbc63bc921a8e1b1b9055da823856ba1e3c9532c
z422454b63e7ba6107cbd14a3e23f52e814e2c65d05e8807a7f407a36716506110945aa84c6bf9e
z0e572825d659ff61b373d46850e1df5c0a04e985f312b249c83b406aacb64724f07cc43cccd0b9
zc3690d4ee616910d4c7b504182f5aacc700de580065004f887e011392708124968397e8f6c78dd
z0dd29fe319c1de46424781072d9dbee446168e5768cf49974a2d718927b6902aadf040c2ccd78b
z3f29bf36245989f220ebd9c3c3073d4d89068f2a951dd0932fb90126d7bafa63c4f122c27a11ba
zdcec6cf1b14e77e82c39018ba99cab4673d4aa351925beb286143ff2f0548d4146d44654368ec3
z9a3aaddfb5c09807de92e25417d86079ff7d78f8db39e6cc5073cabbd3fd6fbdd469762bea34da
zb41e496c30d62f1c72f02ca0db39e2ddfd1bff4701bd1ed9a154485087167ed42175f4f47b0b76
z2475d9b3317711d673194829e06b48653a6f43b84fbd88a221e91dffbbbff456b8b690a811b5cb
zb024423376a1e828ef693c16dd534623f9547aa071780c7b691af5bb63134589399bc903d358e0
zf472070efebd91b935f1965a4fb5e636bbaa50db7af43c570e8dd0564a7391e238ab55676b83e2
z5367fc4fb5e694cd7ee26c1df6677c113ec61382493fa2b83a3a76fa0dc56c2011a3883220b19a
z03969fdfdaefffb26a5a9c8733e91658fed56b54bf672ebf0977910acdd9d3a9651c41650e3f69
z01c455941325d212f66d78e3480de467bddc0762a1424af62a04bf2ae3e70717907bb94190cc5e
zd457bd161612f1ec329e6722f55a7d4a2e007062c31421f13648bbbef950d96aab924b5b74a790
za20cc7595034cbf35df22527ce0bfa314418907f8fcb1a7abadf7a26ab7e3c76405d1d861156ac
z4aefb1d819435af6f400e8e458e0ffa5fb44cd57bb4bb98fb75e625efc58457a7796b1278251f1
zc441b078e77db890b65424ace534c7b3e0cddf5b7f9207f07a61f94ef82039f6760cb8de2d7891
z1d034f27bcb31a8b4257b6f134f5eb9d621f513167ae558dac961dead325f295db44a4792d3f4a
zb425b77412e8334657707fd8816bf7d82724fa1b5f2c275bf5e5622e84bff1ad90154af20edf06
z5416c101502d767f2f54bd20d281452a3ea837c02de1ac1b9f57bff3fcb71672a982a9fcc1c8e6
z8cb14bf553304ea31b86392692e8c4bdd5c015abeb136559f4804bcfcaed94e7bf7563daebd3eb
zbb686e1e95c28a0e3b5dd76490efd451172cacd5bee33e8f29f269237861e43723fc59b9c62325
za9a52cabeea7ca068286697400d8790904b45988c11bc4c0149ef954faf50b64b846cf10902ae9
z8334864788ed03b7e9435a40164c179e05057d0333adcbe4cd1be2d8c9ca896c157c6c83c1b03c
z1a50e4c619a3fc705c4696e2195b34518816b5df84c5414e34872a9f0873144983cbc2275e8884
zb88be7181146fda87ba060514b730374345884fefd5a9a57fc58c87bae8447cc4d2cc0b245013b
z88c131f7f5133700b8949c971b0cd72f4654f38481f34f6ababd107ab97f0708b546c5a566211b
z562c0bc962b8527053107d0903af884463788df79100601defbf1b4b5d5ac4e51b30eb6dafde49
z6d1dcc3eadeb11cf3e1181a1dd6f32ebcdc539b85e80cb34628e749005671db7db90080c6171da
zd88031bcdd61d6ed23d6a45f0f93cc2057ed58dc821c79551604bd6b59aea82057bea6b7f43322
ze014ce3583352ab41940a1a56f99f962af388dada44e2d7fe172c6ca1255e1dbda3b0de197a0f8
za45ae7a9c8f01a082d9e94e9b1cbc0fcf7c11fe605193cc8265d549f8de4d18949e003e2278aff
ze387b2bae7628fa9875633f84c09902c890851d99829f8ba9505305939fb9f764e7cff9d77c8ed
z288f1c684501e35c7aecd0522a7133671054e9e2d973d515c4d61b30e60925d7d2e208093917b0
z63decef7a184396bbffe63e1a50dd67671c3e1e6e04099b1b3dc78563a3babf956e2c323bc707b
z6e7eac93b971af609304554b0acd8073eb41795e04f397b30c65df2aa9d4d3a08615bc5ed6aae8
z6ce3c9775f25e6a99968da3e0c2f02a69d4378577c42b4bee466410a5ff91f44d817d1b25b9638
zbdeb6ab1c2777c904d46e0c435f7f587fc5275b5428c277653c205dc3624d974e85681bd96edb6
zde6e002500cfbcda42be3fe1021a225a6375ae28d3a2636c60d22bb25bf15a493e66e8ae12ddcf
zf6ddd65180427a59bc1ded18490195aeba216b7821f5efddc9039ff62673cc2b5689ac6015b75c
zcecc2742d3d0efb004577a9116556742253d62cf0eb1e03aead1974c3046ccb4bfbce5c8118f2d
z9111403d0211b7c7e566beabdff634f05b4edddf0f7de9ae687bf96c2ad72cb6f0763cf83e2aa7
zd6f85a6b40606822539e84a8e16e2728cf9997a33132154f1344dbaeeb30ac83718b8ed54598aa
z88cdb3582d28020eed1288b95fe16d0f9e585b14b1a76e979e42e5f013aa8a4f8d4766eb2853cc
z7d71d2336ffcf42d0f567c7a1c19ba6719659f6f27a583dc0eea36bc7fc6fd2cf5fac7cfd4aefe
z491ec496d8e1af841fb3c43ef93fac403bf5e607b489327e8e86104e308e33ec3672f5fc345aab
z2c6eb5dc0afe2b370124a8f767399761bcb8318854b970608146c5929d6b3f9ff793a386bc7a61
z05d58428d9df0eaece6afca7f693356a64fd24c9f77a5d54d08b117a6a95f46923e3291a64c212
z8e4dbdc49adeed39491a29afb2c64d12165c501f04eaf9816296d4312484994de1be5a3859ba95
zb19c9aa43d9527054efc789e4f2c7a45b12b4a518aeaee7cd6053c75adf99d27a2f0602ce36e94
z3da5694438905e0f716f8abc1311887ed3fb7d55908ec5fc636924a1cd9601db9d40cdaf0696d2
zc15e94400cc4aed6af1259efc4393182781e64fc235c327aca4d8e9499dd9105f38b53d1617678
zd60324e260988517d66443e63c0be152c97db48f376fe9a6eb6752494d93fb4d53ba85e1ff9dec
z68865fb1b99d1620868ca3d89004f7f23e5beb796ff9bdab7c53e34809fd479702dcaff13e0819
ze711d657927cc05bee887cc05e28ba9ecd1769d5c2165a56635a8fd84e4e235b7ecf7a2c679d2f
z09aec17373f779262deb909ddc6162fcb78a097e22814741aa2768045270dd5e8ffa591393f34e
z32eeffd8e5422c8e044a539bc73561b9b1cb6ecb20ec5b06553882a548d6d2ed87cbf9c7755b56
z15b40478d825496086cb7d4f02d45ff80bcbf6a250b202c7a1b29e10d9c5b6a31fcd90da17f9f7
zcbf6963ca35db203b22e1e0be2c20c738558a6a696caecd70c03052abe8f4ebd749337d8bccdce
z26140cfd8854fd5a1bdba68ee5787be3658753c13564227f56491c03274fb8e51d5ca8018d37c4
z8d3bce483addf671257a823ccd0097eeba2fcf5a96fdd14267fa64fb68d13efcd8541e964362cd
zef3beb1b528c0e1bb47a96a61beea48cfc980876def941a29968438e5d4175d7a32762a402cced
z42693318e215ed27faa1da65c4fde7299d5ddfda6236edf2e11aad87658ebb1d6d20e1e9371b6d
z837fd84b24f70f6a797fdc718065a04c8188f1e4fd48f0c304ded56ee275443c43158fc87cd5d2
z52c752d269ffe159b546f87be0a08c918c721655ce48453837478996f84377f707ace7717edae7
z3dfd8412cc05305dba3a4d2efbe78c90acd6f5468a36fd1ec510f3f894dbde2e7ec92f5709e4de
z275652e453eac7b8a675e7f6e4979b77a9e3e88a207831bfbcf93e9654308520ceb000a180d4aa
zf5055721a9b9e6ad203774e424924348ad84418f7abd3fa6d42d51e8f727f76fbbeda071284e92
zc9101ced1c67f3db8da1d35357571a6ee3d603f8d8db3dbaaef4dfae877e4ea712567162e13cc6
z853ddfc66037d539d581c0aeca45d25e808e1e1835719a79d3c68584be97b4c2a27b8b283397de
z0c3c543a9b5f810add8e9680710a31ac58ed957e987c47b37bcc8097ffdbb91a3f3514b7c29789
z260532e17066a979c3ac8812b144e96c45856b05c673eb418de7a57ca99b6c218849790925d3df
z03cace3617451eb5e19e2dbc23e3b3f63f061787063894a8b7834201bb52c0e2949abe66004974
z14b4c29aac8a76f70e67e263a31a6ea5f268d891af2a84e6ef63f03b1a564558c6c39410a5ebdf
z2978b9a00e657a90487fe7726dff03eb89a99c45663ba2b47f14003d7a541cdf225012dc171a34
zc33ba0abeeb57dd8d77cd3b1dcb1ef1ba600d7227c09095fe84729d633ea567c0adf71fa8589f1
zfbb17040e1feb20f50a3139a75ac5f04f9d5e91d8513e2fac3f0e2eb9719a46605934184056cf0
zcb3e8595d15d99bf9b6908d77d490736bda4a6af13be217abb4c2d16e7d7c22cc01413b97996cd
zb1d723041d8accafe467341c9e98b21d35ae6921265c444fd6aa08608c472c3318bc9c688f1bb3
z6c3c3c6e97f898767e967de004002eb4ed384fed8eea8224598650250f35e46eb85cea0a66d0b0
z59b5ac447f23ea95a780f659e1a7fdd7181d08b1600c5e79a4b330f3f828f8936988d14f2fdf66
z3968f7d109095765a531e8c92abcce0f1ee8cf0571d88f9be006a6b74101177e0a4367d99378ac
zf1f5f7d6750b9fd5e9dfe196f3e46f222ff8919b62323c3331ce52ed6c668e7c8eb845c417e56d
z16f0d1e67b93f8b9fe7c60a48f9db1ebb0f99115d7fcb2bc5ea3880338659bb6714281375e9480
z47e1b70c5a69b798d4fd079bee1e7554e74771cf8a8032a19a816faba8a00a73e5644b1aaa6cbe
z026f10834e90646a67dbe6971d3e9c70b917a31c11720a1177c839877533a298da29c1c908b439
z6236ac163d55135c9912ab284fbc733b8cbd5bdb780057c46b233248ad7081b4f82be692f2dad9
z38b5689e2b828fc13af7645a11f6f0c84b975bf32549ed1e7d0abfd59e49ba855e41f955a300aa
z0cca3c32a612872a4f2d63c1bc42a76021cc5a536b6e34172786097d280e73ce7c7b59f58fd890
z364c18758fb0ffc061daae2b66a15113fb53fc5168bfe7263a27aacbb05cbafe9dc783a9b7d0bb
z4b8ef4945f3c5eefb49c267e518fdd1e0bebb1226d6991ae15d1a0f4e0937d6de518a4ee220b6e
z38f4e44a722834b97bfe62f819328bee44722d47d7c9defdc2d42de43ad87fc12b6cfeea8d0ca9
z58a9a7c4776adaa01f28fc806d3651304a649ff0d53591fc885f0691950fe701fe8e5978a41e51
z4669929e279c6e3cf852918facf951314148e6cd76bdbdbb6d1d80ecbea5d0d50edb6aefd720e7
z9b66901285021687e5dfc4ea288af1d5b102af9388b3e56f8643edcfae69ab419b75c3926a52de
z2676b912e3e40ce6eeedf437ea4d22f6596f9fbea038f0e4e0212ee2e5a6b0aeb83f11ff3fa8ea
z6f57e5de65752440d7ed0afa0e259ade6d3e06326a4fce9f528730a35479340b4aad62fd7dbeec
zdeaa7ce87f08ef9aeb5403021b64c6a861d79f9a0b62d34ee5bd70986c96f72d89c6083d4bf2d8
zca867c96982850be03862bec8bb0f900eddef8ff7335129bd77c88033f9749fc4efca83e85283c
za9d70a4c71b08a43ca302f517ca8a8e9f82d8b37749914fbbaa8beb0c80248ad7c69ba9927950e
za05b5a2df33ec7520063872248dfaf06d658710ffc9a7059862d417c29c1a01eac7a8f18bf0589
zc131847c84f5d0467fbe4b80af4915ab4aa8ebacde1cba0a946642930d7ad28acc3b0be2c267ea
z769f504d58b42b51ed464dc19e903c67ee52e2a5d659825a48ce30d45029b968af707bddd48e62
z4e5bf2157776fe69c5a7458e44056bebfbd4797193cdd68e1604b0b87add0682dc1d24f08a7a34
za99cc7acbea53ed278f6216c99e072543efd43d134555e06941b77d5df68ed55d7a705ff69c3de
z6648b2f725d2daf2c24f9e8171de9b1a5b01a96e4e140839abc43e919856d1b98c4c5b60d4a4eb
ze4735670915845ee0df069eaae374cbbe625da24fd027dafcf356cc52979012a9a75ef33c1b12b
ze2c86d4b8c163e043804ec4c8608977ae3d4db7ddbb2fb5a4e312a927646718cbd8ab8697e3ad0
z529e6b0657541c8e23233fdde2a489d60300298fbe4d0cdbd53caeb3b2502e15b9f15834b1920f
z72be85b495d3b6dfd004118a977e5e3df5171b3047eaa9a751151bd5eba5991448a8ff27b2e240
ze64f11c67f32781bbc15d9685ee6674ba038944b8670c9d353459a46405a15a2b35d220c476f2d
z55918d9a3f650c63e1b77d4e4f073dd201dc497d02fc7e808180a464e0fe84259820fdd73d7f49
zc0709bbaaf61f8d3b20f719b028711405179f7039517b8f3df3297f690a8a9ce151bc231d6272a
zed164c0f4a7f62dfded38edbefa1d7d2210f94c76beefd1a9abe470af2b8a7eb0870ab9ac5d14f
zb38a81b41222eae3e3ee296a75139a9d806facebf0d9965ab2dfc3504cc20de7e349bf58eecfef
z2ab72028d746dcb639cab52513fc37aba3a54cef1e62d467dfcc1e761115d207928eb3b7d7642f
zd152bb69efa023bc8afb11a9ffcaf8c06ca558668e71b199936d77b90de13d8307baeb1cb84ffa
zdd42787f4f53431ca3ef4bf1df26032c532eda5e44ad786c9e828c0f31b93bfcdb83ca3de8ac8f
z132d2cbb00eda805baa04049eda35bb7c155da4da92c4ffd1b83b75ef2b60ca80f55936ba45797
zf5273a841ee8a09991e89fd736911209dc54d8179d966a17cb11efb937b60407522a37871967df
z48952717f3cde2d215e1c5cc4dc71160ba12168e0c87d04f4fb328b849aa83107e96892b9938c2
ze83163c91e062afe2cf8f8dd6e6615aaa8afbed2d17b31e7c6b979d1fec25e6533141c674b548a
z551c331caf991b088340729c853dd00396aeed1b07d817d0e040dee8f9b3345f9a005fab6bd85a
ze9e728bda564d6094d972e20db22708b89e41c979ff1b6d5a864541d05acd1722257a1c2a8a2d4
z09f36fafea1a70c91297e280def24820346c228f85be3da985bb61d0a08ab5cec9cbd5fb4084dc
z303e9a74e9dae58ffbc90b6f36dd806b21761a06a535ecafc5eac0888a785be69763cceed11068
z20415a64be09455b2211a1dc920733c6805bb4f05208a82cb044a9a11c0f2e6bb57830a667cfeb
z1fe20dc329db3247d30d29d7e1cdd115daa25c3fef4b962108b755bc189afe92468cddce1fdd3d
z205188e12567aa7d3c7fee9043db025b1bfea4aab137486205128b80850e7f3fd46ebb0a9c70df
zf96b57ce7c9fb90cf606e4bd57f854e96f01c02979f13c6374b6288b84f161cdecf587b2e92238
z0ec33f272b1fc3d3ac2c6676a49c703020767f811f15851dff55810bb668a57e545b0d6d5de1d7
ze7404dc8e1af6e77b42d6a9593bd7ced61ff15ab79ee8aa2099841a3b290ff69cac92d534d9df5
za1ac47015337faaf34c775380bbc838c8c4d919666574fa1ee190d4a5973d2047f1160356099e5
zf7b25f6eafb3ba59e76c74d470aa3376c22bfc0baa57e9ce1d5eeacd2504bd9f7cd30faf36f14b
z3ade8425fec7566c22d19e941718b6bbe88ed68de45c05d3795d8f9ca0d7241f3568fd89ec1d5c
z0e0b39dedd26c2d833c9a79ba3b8ab29a2ec023f974a3e6d32f654fef77328243a9b7c4d6a4605
zc47bac02c463824b0c075fd57ca42c02e077f71a1ca542e6f1819e8115264790b8805f0ee1231c
zbf95faa1d06df632be148a6512b9b8d69b1bd2854dd942429481821ca733ee65dc024861e75c6b
za281e5d2ab1f43b6d43e5e62422517cc0e24c9ea4f576b49cbb969622d7072d95039891e16e22f
zc0732c57dc71571586b9b34255c6101d8e2daaeea5b44bc1028e8dcba82145442c5071e8c4ec6e
z159d8e1b37daa1f4c9a4b9548401f3548b5b02890f6836c28dbd25b4b2965f5ec773add3768bab
z21d5bb8d40773ba54e15889cb1f1845245c05fedfd70ff2a531fc605e6c4b67e94e7701da1f8b4
zee748617bc3f1522e2993abba156eb3dea4cad5e7cf6d704e5dd1d18dc50e8cbe2161d8633b813
zfa2328fce0d998050d1aed11343ac26e3a790c28179d5ab9e70da1ad97eb55dcb835b8ad48d04e
zbdd7e15ce9de2ee08e90086fe45d201388c544adda3b2c442e56aa5005f3475a758bc7fa130f02
z73b233b58d3d218b95317a84b0022a1ab394b9a82df4884fd9087ad4ed6ccec4c5b1d502fe7c87
z1371119b19845cf83fcf1c6a5611d6b3dd645a160fa849680f1bd5f3391bf6afe96f8006a34a7a
z18409f38bec597e52e7352b303bb4ef37c5a62bb41f95925dc1f6999362d097d7db871a947f45a
ze059e40844931d12eea8c554e92d554674ae5ca80bcdf5ee1e2169855271a38504d889cc8bba49
z0d8eb3087b3ea8970ea2b02106a08ce23e275976ae3329147de28ef667b6f1f7f70ffcb56750bd
zc2c1aa80fed47afd6d86d148541c7384b70e0eb57003ea980df1db47c636a4c1d9b280524492d9
z49f94d54bc20fec616e62e84ba4a44295ce5cee983d26182d69ecd0c95fc80d92572fcddcdc457
z2ce0fbdf38571223a92c4d877b90ad2a578f13f1730796403e813e8d30deab64cf1db6549fd2fb
zc6cdca66cd73befbb411f2fe476e3c38e414639a3e004a7a2f0960d7303b49cd1ac3f3e9fa8f46
z3e1f2c94177e3063ad0b992e47821b6eac34837603e0aa9e4f447365d7bcf8dc50c46c75da6ebe
zc06daa4d8c1c38ffa8087ac72e126c25c6bce70d86ada582dfde945c199d5d58c1a2dd1622c23f
ze25056c3badaece982cfd87dad0989f5b5861fa53701709827542e17c0623b234d1aaa46924816
zff0065af644ca4c398bc23b04ea3209d07591613747af5c081bd100fd9b703feb723abb7cef1bb
za1b7eff0eabc37cf9636b09edfaa207bfe37f0df22b438cceaeeff5975035ad16a066ebb9e0b4b
z69fb94119aa980e16406082b133a6bc35da7eedf4877ee8f72941335e4f9b0be4a272553599f69
z93bcb43b126d7fb4fabb5997cb3495f633751df9721113f856bcf7c65e49febcfc1d78063cd28b
z9feb3a77a37213f8a5cc7fc3cdeb1f5e17e456b5151acc94c71521e56fb463f7a6c41ca6090ee7
z5bdcc7745ba8787c1f7fe901d0270d7547e9187e1c2932c855b66e7a8d0f9e0109274b6b714d10
zefd2e0e1c69aef8d7c5da995d80a7a2e63a166e474ac7d8e1e56a599803e43a9f7cb7e327a0161
zf644dec737fc8e2a8038b3632fe1f63b43a5bdd98d74de059680184ff2effba1517c1f3df1c3d9
z66fcfa762acaa162b6610b4e26206da4836f664f17b2494cbf91c1bb70f52066e0a9b851ef6d50
zff91c43bd17d4a906ab39498cb028663cc7b87dcc51ba15ff236c5efd5abffb54244635f43ad40
z8e5b4d442e710c935950d5a7767229c5927c022fa6ed0773f851ca95c83376c5d8c065a573cb4d
z6385d324e09a4ba41df22a7db9ffbd3eddac9fa1a9f97f975deecfaac11ec44b52b75e6fd1ffb7
z4c9ef95140ead681bd77ef7f6eff7230ef548d337d4a50ef5838ee500ad83a25c9bb428b44d904
zc3186b787f93b1010cbab334f132c34ac21379ec2ce56dce63c4172616ffcac6c3d202ecd9d578
zaad34c7b45103934373dcb6e5c0c9c4edc9ce524db2f4baa635f93284bb75d37180599adb17bfa
z997f5a21448a977dde0a169030950ebc4b958295d5a77d0cf4bf2f2eccefb4f1d2675280ae523f
z31bdebff67e6bd6204949b2d8f5e5ede3fe6141e1c62133b740c409f59736397d588a179fd27bd
zd00a929daca0005d726e442dd1ec39f5cba7bee6046d76ca488c3ee7f07166ab5a8e8fb0815b1c
z238ac098956f348c8504b7e409606ce540376bb77eb259d434c07e59a6778e371517719a80e707
zd904c9fd6cd9517d6983e39fed8484730a7cb23fe0c76c2a7edc8d900f76f442578c234dfbd9d0
zfe2393c5178225ed01d8d4635f6b727b07fe5f37366f0c77d894bde56a3f3a159e852a9519d601
z5548303ed74ef1dc0d9a97f23c7ad27ec2fbc3015e02e619c94feec7848ab9b9cd85b117d0a865
z0bbaa423c1134e44e67ad4b85ade0f71871b526972329da832732eaee30e42726eb4c57d28ec5c
zd7688a61a8a49785775116c5420ac2857c208ba87e681469e22541744eaa6fef6d26a785ddc215
z27a03de471b0d4cf05f0dee2ad650b11a2271a64078c8acf2cd2629f382cfd9f91955aa7ae6d7a
z18be1a06527825095308c818a0c7260270b7908b04a97edd2a175b4f2dfb420ed903672c9b1548
z1856f87a2d1483fcf9bfb8f86be456353fbd5c1863ef1b5fc72beb84465ff4d38c903f991af3d9
z00852e448377aafaa6f3e2db06454bd05158b90a3c6a9e3a5bb8eb75d3a9f4481fb5ebb15c2c14
z76ee732c96c5b3b42d61e9ad9f40ca7d7d59120000b97597162a8daa6a30b1028442de2fd9a5bb
z8ef2469ef39c4b2b7b6c2621de0ae36e4871ab508329e7bdacf8cdaaac2b7a86c5b6ffe2fc24d2
zdfbe8583d66667dcab51d868324429e127d6bd8f59ef8675b3d1b543b23fb08b3f6973f57559ce
zc07a4f824a957133fb5d3266e7647e2fdf5791c1cc2edf908e3f64ede32a858955186d57326345
z8b58ebbdb6e059e95e192f33379f12c1d5237844fb0aa5fbac1e25e44f5d170e88ba34ee223701
z0b2a747a2840079ebcad65d5d972d5feeb578260d087546c61cbad332a2841059a98619257d1d3
zc941dd1787b3cbab41a41cd4505bbe21410e7235a24532e0c9d8648a00d387b073e5b6ba6806f1
zceccb34b1d9d5feb0a77c5b5837552b1277051fbec4538ff0e9156a52c9dbe48f713f546fb41e7
zb9ed0de4c2b8f50ac1ebd47d39200c749f8f618daf333c3431090d84603761ba80290cc644fa9e
z4e4e53151ca395b2844fd7ab6ac591a15f70aeeaf3ef621339e74aa1dcd590891ca25d144a4ec7
z295710842e6e946d9cffaa139faa0b7689b00f1332d9273193d7973f6694e6748d19957988b21c
z313007bd1b8163fd8e78fa092eb7a893ea9103f4e7f6404906e90b9ac1d08933242fd0ac58d3c0
zb49b255f6fcddd6ea8c67b8c84528280289de08fc5d6a08ecb691d37f40d6ef1521fcfcd78c07a
z80b5d3a3fca64b925b3c35af4d3bfe300dd6bc3643b74a2af523f6b29f6c971476b9a7458309c8
z9675e26bb807d0acd432f7c71137ffcff890e3975dea7cae51ecad278d1a892eca488202c5c245
z6c9c338c0c2f74f2b6d5ade239c69c2ccff78fe7053bbc2731e975cfa5f073e08bc22e282600e8
z18e2af65b84253819287333c5c9d9052d84245408feb3d235d70eee279776dda322c3a96457ac8
z9b76d6a2ffd30ef0f9ce31792a0c3436d500c3cccec7b4d572b96b743a29125d82895e32f05257
zbd89d95ee4bc7d245e325267c157417e8043ef6d4eba89f95d2e5d9fdc83e4d6d193528964ecac
ze6069133de73df20c047d1baf14141de279f7f5ee7968c4629779d0f2958395d584a8cda49dfc5
za8228fc3c9df6382414ad8fc426a562af17bb45b447ff04a12393c2d3650daf81883b29bf9f7c0
zaec88f5fa751835f482eddecae8d6efe84dc0b92f4e189ccf3cd44353fe245d87c06c626bb870f
zd9311030d337acdcf6f3d34c070ebc87f4e16a748eb03e6922c40ca118ed35c9cdfcdcd4d7b8e1
zfdac6f0047141a68afa5c7e67ae85d3472bff5ae7055b2dd60402e6c4e5e8262c5b5f371469df6
z9266c4e1d6956938d774e66506b022b69568c4c9c2b92ab96b4cd43f561f9c84387c2468eaf0c1
zfdd9c86f1324a50a369f418c971f928b8e4a627a83d6d4cb9585a607aa0eda16c519a631395ef7
z9349f79ce9fae3414e2244a87bc86d70d0f0796c7b46becb5a901710ee6de9fff9fcdf963f0ef7
z3e787f30e3fab3701ab44cea12aec1c087086bb9fb866bae9a17e1d0b4e228a6594b50e64a523c
z9f9433a58cedc389918346d19b03ec85b6172a948366a77b3a289e90f5d03b68384b5de78aa918
z478e19c610c2cbc28e8509c7ab4bdd8b82865e89cefcb8ab64a6d8e894e349fd8a25eeb8c91df8
zf9bd12d5af2fbfe35b742f6f6be9d79172a9463a3f2c119f970484a650271a8f07d8b1e8d109c4
zf13f0e42c56b5449ad58035ee3352e6c0080ff238e21dd2ade98722ccf9d19f37f4d0cc1e62d89
z9c04f93aeb842d364ade13890d95a79e85f9ed5d1a48858fd70aeaae42672dccdd4588e8e28c4d
z9fe55e3c01f0d899504deeb01f7533e17a7f58313d1097c3d422874d421f70d9c88f0bcbc3303d
zc208aa3eab384d251056caf887ae979b820c20b3326cf0c5806b79a9527855a9e76acdd5373913
z15b6d762da48e710dcb27c960136f377b72761c55bcaa3d71c867089336ced43071b24d2b70364
z247b17591b02bc50d2d24bad49e22400f4024759a660b242dd27bc9985e6b5ffabac09a669cd14
z4fe50e96d286575aa3cc076d25ee7639dd23259437af3a745e301584d4c6ebbdf3adf7f8c57df9
z0e9b206be07be8373224f648aabdffc15d115ec66431a33a753f4708f3faba1b22b75ba1c047c9
z8fd982c2a2b0addb0be5248a767cfd73d4d2b743689d6324b63c29820c23cee4d637cf30b641f9
z59d31dae063c17dbd263ab0c6f19007e5591a3aa7c66abd649067543af50fd368e37cd1a697f72
z7d550454560aaf6296e404d3c91120e70592460ba35e531237dd58f979216530f29902e1db6ea2
zcb32d27ce93c0b463ce2418a32e723f529748d7c8cd8768c4d1bd1e2cf9ca18ce53b6b4919f709
z81725fc8e7264eff8f3b8c7d8a1371d7600d84d5a9df78243a24e8f4413f9aebaad62e5af2612b
z9610e6b986ec8bae7b83ba8ce55e2bc28c6b2c56c863675bfc63866dee8446284e84924b11e8da
z7c6fafd74f0e038c4fae62030baf686f8931ebfd641e247980eee4f7f8469de4b101478acbe8c4
zad9a1b8ef2672a8d128ef1c599585051835802211cf05ce9eb2baba4766105b329eedcf4c479fe
zdc28e2c1acfdfc44f734cf97adcc42a858cc5fd0fbf768f20016dbc8bf0e45f1cf34fd2e8994d8
zb397ca488e665b3808671bbfe66f1f653ccd3e9b5b6a25756f61535ac85834991ea42c85855fcd
z81aa34024f36bafaf37cb8a03d88164ccf9f11bd309d9a1c07edf9e8b3de3b6980da72b010ae71
z20001a8fa098244c8aa6eddfba83aca322c57f37e0c360b0792efea921b6704d126a6ddc554bc0
z21846b5cc69f14e4a8342a7405d782bd1601773e7eb01ed8fb737f3df29f5b91f158d498b8fdcc
z853d360b96def9acdf9e096ce82b0423c3d8ed85ce8272fa9e617c65fdc50675f6e7732324b698
z23c3d32d5b2e31e605b9fa8df7b7ae13cf79dd4de8ec0dbcfbc8903042b899481b1c4623807449
z4154c0fd7980e37d2e04afe1d2d36f12986a213bac8e48f74d8dd2ef3f34b50a7bd7746ebf2f90
za90c0d4288524758d762ab3c347784a8e9a9c065b3a9a21e666c4e6c4ebc88182549ca30feab3e
zb7b90905d307096802b4d60df54adda35582be3a0a367da58b8a484d78c74ed57222420eeebc7c
zf32230f101069a51be53e26e7f059f3c448b6f79eabbc1e977c12f261baabaf307c00b89c17802
z74124fc8ec6e295fff6ba27ebb3e3f1bd823f2d711275c2a548bcd90937952409f25e6d75d9276
ze67bd100bf06685f8d35a338fe366c443fc1d2221f1b8a7769ce25429c189c6fb178f1ca9a6b93
z50ff31cd9668e2f266905dc43433093eeed859c18656922e9ed698e926291315c7ce4cf41e196c
z6314c800461e3ab9c4abfdefdc5322f3fc5002a55c20934082bf2f643824228d41beb8fc855ccd
zaddd89ad6e3e795ab6b2c4f94e7b90987f0b5d48a2f2ed62525887a7108bf25e2c40c4695466ab
z2c949c425a08340f414e9b3f8b87c28e13f7d9917038fdafef5b6769e001bb2522c7c35d7aa7cc
zc6c1b1573501990f20921d330b90a1aa959ab00f73f24e92f1aaeb0aef8a4acafd0974eee619c2
z599792791f97ac4278c439aa8afe5a480e6e63d70067bcc93fc03dd2c0366b69403bf4455ccc8c
ze8e7783bba4ea2c7f8481318f52e3ca1207d4e1c6fa1c21e67e49a3d715d38cf5a4573200ea0d6
z5b0c335a05a0b92bf3decc770890a43ca32e5d071eed233ca593be20c7a9706180788b23b80bdc
z8e5ea8327617af5319aa1235bef9370a9be04607d46a618401e8adb1f7fe8c04aa7524425bd22b
zfe2437db5bf3d973749e6412763777383e7aa4293377e1f2363617b62f25f106b748dbee2f83de
z347b496aef3996aa06ed570a457d167c854754107083d4d79c6e3bc728ff6ad631c96fdf32340c
z0030af9fb6a213dbd2fbeaf4615dcea181e767accd02abf9f145e50b2c39d471fcecdda63533b4
z3840d7a176e8c263c55c6cd071f55ef3e5f0b76518aee53e4e3781c769a384cece58e63b4ca9cd
z46c1331c957d02701bf7065ff4010bdb2157a05a0cadc57374227a29257b972f384bfda391be8b
zb54974b9a9995a1a826c6e96b8e8a442b761a193ece13e47ddb2f08d1fa072d8e22b0c499ad548
zb49ef3b2c36bab52d587ac917ead13193b0c91fd8ae909536df0918216c134806c151c810e02ef
zd61b1247cef8905282b4404787dd311f5a426099cea140b41ed5d1e5599344e2ec55dda7f37ed6
z4a83c6f8763d4a8c099bca50232c58ac16855bb7e936986311b7ed062e825382bb8b039afd3322
zb9d14b8e9d7f867ca614304f2c342945ce3f80423860fa898bfa0e249564d8eb0af457e2d8f2df
zab1239ebfd203ea86ed2697cd7de0ea01eddb55ff469b517acca8dba6f828c3e845c2a45d68822
ze6a4543d8204e71dd345f108d8bf3c79b28b2c940f68039ccaed7a3419c9c62f6eda86439b6028
z8fd9ebbee34795d64157be80f199f6ec43a023d073b4a12d9a67e63eb518fb257c595b7c21f2ed
za9caa3e5236726f7aadaedc30e229a0a66e948b8caaf41b421357367df6fdbfb3c1edddc127b1e
z29c3482e80b9fae641fd249eef89a8c4d5ca4c4db2dd41130ecd1e56dbb2d08d54d620d84b2e27
z45ba1fb66ed5bd0172b22d1552d4e23bc960a0abbbfb25fb27b80030fb7866a4c46357fa178356
z2d85e4eaeb76d5e68b459a4113ea14ee6801dd09425824fb5a09e6acdd3b933dc8eed1ed8fe007
z9ccf3578185ed55fc910237e2b5e2db8a8d0b8d8558e49019c2fede4518440a340f7a28f0de0f1
z5015b64c499a188c738640d32cf930e9daeffd5acd83c92183534219337923995310ee9f0114ad
z166ab0f00cd8f835c3210591bf53264277a1c3964ef7be13725637b55547eb5ad1a37be2f3bcda
zdd57fa171f4a4c56c110f403651bc43bec61a9949947b1b65fd6a4c1d5b55979647856d05f1d82
za46b47a5a3ba3bbf921a5e2fa394ff3bb3679b51d6a852547d510eb5a7d6a8d7aedf3a79c42a1d
z7dbacfec92044541e3ab1ef08463a8eb82d38af238b215e38d2d95bc74abdb3e7e1d3df3d48d50
z6fd067a6c4e8c62097829391b81236cce296866c56522f9ba87dab52818769d7ef482af6d0613a
z82561f76ab1b1c44f66f7af8abd66c56b52722813616f78b5582206a5262e308b66a34ac5c08a0
z17a884b857759ce2bbf19529090c7f7f0cd41c472431a17704c47923c8c7b54d7dce119d1be9e4
z9184a8368b76824cd505b771969f87934817b04845b0e692cbbfe507455a6141b397c0473d38f0
z6c771907f7991e84894d5a16ec4fede66c934a66084fd87e4aec340ea118bcfd8482a651996d3d
z61828d1568f4f5a06641514f260de9086171490bf10cef4a6c3ba1bc3b44e0cca1ccce8c4a9901
za3dadb6dfd0c7e86848ba90b1a1faa1a3665ecbcec4f303ccf54c8b80e90fcec8ec5bec7e42578
z574e441ae50c50cd14fd50a5706f534fb3c2c8dd345bb9dd4378521121326390b33147dde99ff0
zd7193c00420246086281eac629b1661f1fd80324b8abdb652466f0543c3577614e095547c5ca62
z0bd5874b35679b715337de8179806ac2b7cf88ea3c247081c0e33e4b29d305f93827cb0e280c31
z9aa551c3df139e54934171496ff27d51a8366538aec6147181623e77a35dd2a054f48eb216c94c
z7bd60dc29c92eb879e515b6b2cad8e357017700a866d7c809134be95b59d271fc1eea01a9d54fb
z3879f8bce1428604a4084e4cb22d40ff66e730e6f2ea60a131afa15d3a74a8960c5385e66fa83c
z4df4935e182717292e1e4b42c09c104bf1b707d6dba2305f00825add01b29b87ff2b5391399c46
z1c83d7bbfc37522b758d34f79f0aa7215d1da12b618e361fe2314cdd50948d358a97fe18802a0e
z9a65bfb419a2d089213af326f27b9aa75e70eb1489209dc14410b82796a3a4ee4355945997facc
zf2358bf5e77ee29b793be5d55a7eda0cfdf512459d27dae9c3b69e3b7238923d0e18ebee5ddaaf
z0a0924fa30c1cea1c70b1452b9ae1c219c48eb86a1d1c5974c28d6b2f9f98b5838580d17867441
z91f76db4a280257b8da10c5e48681702542e0b6518fd2f8f2f725d96c52dd12b95864a37a11b10
z07e1dd4190457ed29d3fb8c06ce90ec26e5bfca8f9c2a067322f40faa33ca8a3dc5d28753f64da
z957f0635454dc24cb2e182264689499dd1a907e4eccbca89ed874da46e387f1943ede1c9fc7c2e
zf098ceab3eb34dc5f6467924411ed57439414c7ba11cc89b805587f4e1fd52827688f80df83b69
z5604deae03a9db0fd32553385b7d5eb725079d346b6834bb82a9f8db8cc9ca93ea87dd66add853
zdc87ee6eed31853e38ebf9c3cd58cb5f769f9a71b166372800a67b073b68b2f6f81f8825c5a9fb
z6c1de3b98690480b54cfb0c6d1865fc4167212e415a9272c12c07b978eeeb5c810742476ddc7c2
zd83f7ba04193481b4a9a299dfa07d5a1672e82ac49aeb7d58cbf9834ec97fb239166d8e29a07b5
zd54ba08a7b0c290a17a4afe713fccd45850405380d6936c6090cddc6fd474f151725266e558936
zf0c64c6aa7dbccbc7bca41decf599c7cc989126051dfc327fa9ce7109954d343eaa4464a290036
z3d4a86f29a7848bab06884a95b384a943bfec5521f85deac3afd411edb3105b06a9784caf93783
z41d0a805cae349aa17c746c2a7e3f1fa5730bddbeee2ebb5e3642a5162223c70bd78e4c7abccda
z00b892355f2195304593e9f6236c20f1f01a7e4c2b6dd10d77097d341f6909085e946882d25531
za7d7e9e71bcefa867ba547c5d6ecb0063e5385304e85db5f17cd5c032723682920f9d90c9d0fae
z2805368f928ba855ca544c984c7311809c07b91e5a2b10f0ad469f0ce23d756f02af7278d4eb2d
z19903c7cd695d8acee2a2a7ab10d544450a89fb9aeb433dbef6426c5819b26cbc20739442ef935
zd27615484ed1462c13078c5c889f50669aab601dff3992ddcf8fd2c85b339d7dcb157d843f013a
ze942af0236255564951bc61c75d438453ce7251e4cd72f6601be8236e24056cbbd5538723325a2
z8b247f8a99a973eee388fd20119bb9e69139c20cfc2ab988d8c77d046e45615fd1065765974a24
z1724235ea168ab76338a26e29ba7de2f258ddeea30aa4498eef305b5ccb71b930f681c067c3e2b
z32af48d7da4db0e622071b9ecffc58050d33e6e3a39788a1b532a3d247d9afd487102a0a5d6400
z42b5395bf63d67264470b9cc2123912b4e5b0c166f3d28422bee66c794e1ac99ed8be9544c633e
z5cc01aca1ecf3acc43e4616676d81a6a6a047af3674e2119b73d5d76875e3031e6851fe842e963
z1509cb270001cf9efd1574027299e7bf963016e8728faf6e67096a1d6c6952154e2a1a1d50db84
z2dd924418a56225f0de3a2d5605a8f5afbd799db88e76338eef62ee0fdd55e89f28d5fe16ddd37
z058f0b959d7187e019727d4b5596aeb399133d365339f0869b96e01b9b88892ac533dffa544899
z96ed65e678ff214be9e27f17ac91f391278a5a16af3cccae998d3f27a64815f2841c34e11d5b0e
zfeb79be082bb5c0f4eff72678a224edba5c9c8ee698859f9649f34b007d9e571936f36bd106aa0
zb1920c34c2777f1ad01e648d4566e616d736095728bf0f48b2e8a05afa2859807e488e80ba90a5
z964af8d67c78b41b7eebea5f534e614a2e8cb0fea044c1adce0161863417e30e29484b406fa00c
z69aeca6645f2c56029b7ac1efb6829783e4a95f24431d9f0bf2b93bc1dac6b1f7fc57dc8bd42fd
z85ae6fa90b6b3d0400897069d4f17a61c21e194ae1b60feeb8e8108b593dcf69907e86588a3c25
z5c42b4003dbbb8d151e7b39fa73201b9aac6ed2eaa055c57ac5fa1ebf826ac002fc94a53f217b6
z3d86b3d43dee213bc46f04b752d64f7767b53145278cefa6011c874ed5ca467ef766d8632009d9
zd07e5f38c54f3920d12e652fd53ae9fd25a8784361108a02f215bd24b5ba40c36f525d1f46521e
z4ae46ca0585085eafd8113bac1c2a285b0f6aa91df0cbfc55e331e780a9e47ef9cce3c9e5166c6
z2944b1242049d69bbc3c3cb079a35cc3636bfd7cea2d81a05c7aa5f9e3a25454abbcd2a7d0c0da
z4526ff43c52556a0d941635a88e8c9aa7816a3853c1ee2559d44e42a0f51f0690d04282e9cdb4d
zba7acb12c6b47990ebfe89f1fa1d349839ccc6e53591c814429c3e4e168ec3892d7a805ef98afe
zade3c404950c6aa7c2a6ecd88c413a757059f261097bf7e78432ba24308194e92c0e01447a476a
z2c88c255c916a81433bfa738d986831343cc73cce4b6753d4fe0c465fee634ab313fef34c8bf5f
z62ede72a9e1109e97b871268658ce6d4f63a48d89abad86a077ef6ce8b499c200e64d300743e1f
z51db092238c3878044151b572bd3e60f8d88ef38d952a87c7baeb6886767620be1e3598310fb35
zf5f52e1a84fcf1793e95015f30c289c28fdff20339e5dda16c703c20ac2e0c7dec473a19fc62d2
z9c6d212b2a31f591bca97b321b91e17f645a34c568f80a14d26335b6d42aa360059c451b52028b
z0a92fda662e9259d30bb352dc9a24d053536f503281cbd973f46fd13b0db41a9d21cfae583399b
z6768900040a6d5012fa921283b6a7776f4a808137ddb2b257b1647a5b1eb44e00c383352d28215
zb0d96f0015e505262261de82b5438752acbd46f25452dcce9a25e50aa5ebdc8826ae27eeb67d89
z317deb5de84cd43c9f78d7f954830afa62d769e07564adae5b1a70daa6c1f31cf2cb74c5473a5e
z234810f3943e1b485056c6f44967ff77ceddcb43f6c3437f483f88235ba5d39d005580ddbdb382
z62450aff0b636c394cb132c07ff0e624134d012579e4a8a9ab72e89edb74d0655864777ca1add8
z7a43f0129eab5a85f79dfec749a211896f9265ab3a64e6877b45ad65345eeabdef47103c328f88
z7f6aaf2c0eb585ee4d052796a697b21aca70b592166cf42771f9c71410e91b5c1e9cd744616378
ze8164c948d03b64f2d028f9b97f4c5cf1b3070e459746ccbbba95ba7a5e7b6228f6317319c998f
z27ed89406c106dfbae7e70e5b6689d8c6e49ff2023ed463bce1b8016fda5c00958f3696de42d71
z0c8f0b952250dc8b39157eb31d09a9e00c3c4f9554b5ec18b2408a9e6ab042d344b791ec2def04
zf9f7c9b1fa3122a47251870e5cd7dcba1456a27fac706d4ae20b27ad61dee2c1ff481c8a6cd843
z000aa2429bb590cbac92d64d343014001cd8446e6220f76fc0d1ca8e141427bc0856e8e45a4e2e
z5e2c3eb4e8e801165a3a3877564e476efeb2e723d5aaff62d825375eb8e5f7db00195adef7e659
z67e74c124cfabd9015bd780d2fc8b71f046582f9c84c182f5e7731fc33190b283a5df498e5a1a2
za3e50e4c8e0cc3709672f082c401dfe982ef7003fbeb521e1666549452dcfc1d9d574556fc6aad
za237d467d8b83445db9c48e253346ba29293eb64e3cd4eddf2103f4de0ffa125c4bd1da8ca054e
z28f0c01f53ae271643a26650cfbf3468c828daa351f565d8fb69805ab08ea82173417edaa43160
z62a5e22515acaad199159b7f12d0abdc5e08832aac66c65be214905f9b022b315f636425370020
z7d84845f8c2682b32414159a62ccab9dff9044fe9eef1c5a2dd5dcd6463a24780569b6b1eb784a
z1c489410555629ce4a989f923374f2e3a871f1ab13fa9ab0f92501e0af4a59990d6cb63179462d
z62d61d5e087364837302ff4e968737c7e3fe7e5972e51a651bd9542b7cf5045f66c1e1b64c16fe
z784c78cee9adf110e22a88816ee8d64d57ad30551c4e1ec9752cfb512aa0dcd82f6896b3079902
z8313ff5115ddf88c8b2aac2c6fb93b5136b4d0c13d9d41e687e4bad5c97f1701cce22cb2152005
z14cf18243d939ab261befca09d0ed94657db43dddf187942b68a3bb2d6f18634915eefeab7b84d
z93bbaff688083b7c3011c6214e33bb401d9a413191bacdf47c28f768b640de744cdc4875697a56
z23d7cfd1cd156939a469f80038d90b53c07ab3a6d8ff8006855e828d057a227c8a923876e7eb20
z9d87adfc163587c158fe0435ce09dda441a185eaf4142c26200dc435281603386df644fafce04f
z161147f15e8774efd7182498e93325cfec9b89eb2d3664ecdc5312070961d78dbe52b9e76d8def
z9997d630c75b66573631f99ea1819b01d6af1be20c563b95e0b8d73f8203135df4d169887bcdec
zc76df6a385107ef27257fa44ffd84e31506824728536bae90e780ac97ec90b249bff01a7e13568
zc9a8e1473014ce337730e2c80f150d4bbdda4482863863197edc2da197ff666559561eb0ea31a5
z540e73c8407e4684d91c35ba4d8c3293b5b67c2956208d9b3ad982179af2c7d949918345d478dc
za7763373ea7deaaf2922b64860cec822446e6eaa60ee9ac3ce5699e8de0405720a003027b3d2b9
z1c381530557844f8f8e149d788b4c760b06b204bf6b64d5745f209f45a998cdf2860e413682cbc
zd7561fe23e9491685525d2b0b0e5440b6264f0938a201132b2d033fb04625c38f18a89701492d4
z266e16273ee3f62fbc49602657c08d868d9d2cff3e6a3590787c626324a36331425fe1cf07dc65
z14978eae7634c1b5fd992cd55a5a5d4a74f28db34d53af40202fb1d2bff7140c73d315aaa1964d
z5e4f307ff1c8a9bf8cc26623b44d625efd65418bd9f015f3cdd123a299a402922796c96cfc17b5
z11b12640381118df09b7a232c95677f94c059694dd58ca042c2995aea2c75c0b309049dec53e0d
zd02874a5120f50ab72c668d024b83a36e70ff113a4467564f9b0388f223ca191b3a50999c45a3c
z5f2a719f0448efd8ed40ace872b7219dfa21ef6bf674ffb1bc8ab0a1eb37d1e866f2dacd88484a
z818b809bbba64e531d277afa80111972241c5c4978b0e535b5b406e8349457e9257424a85a3904
z7bd078a42f2da4f69f399caf5ee33cf4fab4e2ed710fcb4522fa28efac118452e2bd6b1f50bbe6
z091375d9cf76f9201e10a77cab8ffc26ac69894432a3573c00474fa23f3dc7dec373505615f5af
z4ca4a24662ba47e119cd42fe1cd2b8e2d3f76b5253e7bb51b26ae65c0838873a052187fa06630b
z2d4528cc60b9446fe612c6ca6697ecfc2a9bc230ab03a458ac52d793efba02fe5cd81886dead13
zc9a6205be2fad94c0b4fb047d4325c501cf879cfeba0db9f10d0ca715c93aae358656feba0a026
zdde65a0be7970cd1b6e93527cbdf921db9a76b97f5112cc20ae15f0221a7821d60ce9eafc1f04a
zba4850ffb898ee794fa8509d96f3086e84494f10de0407210b57e09705b122442451eb83b7eee9
zbaa3d93aa16fd1e84203ff46e6bea290b549f7ff326ec9e08a1ed906062b552cee9f1d0d14191e
z57d53b97f17d598f6ba13838788bd20e577202e2ee2f36cb10cc01ab6f38d0607fbb2522f66b38
zd30aa69c2ff013f7182620067f844bde5cd2508173ef255f77eec86b0a16d735dbca8da8c9ee17
z471d0a9308bd59036ee5b73a4d134843fe5bf9a5d6caf47a333bf42d59c9b7253dd85426e12b57
z9dd1447e12c82220be4c5f9ac7bcbfb5cce25c2125c5dec85998a8a03019a79f69b9c568821ec2
z2204297f3dc8acd90470a3d7e38023e81f926c34d635cb6371eb231ffcb16ab37ac7c52750b1c2
zbd60d42b74f1706e0d9d7ecb3233b36d9990f676c4d81ca1ce6dceafc3e192cfe7a7c85d580661
zd8a9420c9316a870acc6536fbadbdf173a29afaa89df1fe177b01e3644b5a2c78555621c6aae94
z4e8aaad1f821c9d5fd16d5bf51abb564284d5245620aba57cbd9923be4c36201213eee1b0fa204
zca686d3f04a4be4082a9d952b457f94592ff1baadc671b09b739c0a0257488d746680ded8807ca
z0274179d250ccc0fa7185b46a69b07ac88ddc028b6ffb1519ffdd556fa45fa4c9a5d790df009df
z7418bd020a1e7ff05e6e6e13dc19e5b57c834e36888b6e532f655beacd5c30c5eeaea1f05903b9
z36d798b72bb6cebae97d1a215e999472630f8891c7bbdb8ffdf99ca238ca36c9080145bd17c034
ze12de27a99185e6835acb1a6a18b516c83f7b3e89d4b893baeb1583c92977da48b64e8fddbe72d
z59d399a070ef9dfccf7a8cb697e96258f24b9a56c7e02ae9985abc2ecd4301ee11d4e7cf09cb8d
zc5c7a8fc92909200185d9da0fa63c7224b772a949a1bbd1bb57bb34b2f9ac754db4dc151ea61bc
z5418b52de4a90d0f61b006dc2f9f2a55b9167270813892a8f686e2e6b0842271932cf940fed754
z578a4b35b70f1bc1b932ee7ba2e9744609a80c74dbccd760b43e92a698b98f72534b9e0d51c29a
z4226195065737a3f38316940ad3faba8021efb35a50f3defcf1cdc681a15d2d2863ae97a31b2a1
z80bf64602e210c9199575237a53032a2cad7e2c19048eb502250f686a8c8d1a8982e68320d78bd
z744fe13183cfd07cdb2318abf77e2b26cce68f4f7b1b50e2f0ebdaa705b883d67824ef6d87b167
zd894651e91bdced846117165ab952355445c331d47a92d928540416d101aca94544405911926e6
ze865f383796e04b516de31bd3003e150a6b533476fe8de4ebbc1320b0190ec2f6190d8b5454c75
zaedd67ac300030c7f3b8afbb1fe96e0dc28bce980e0b4f52e5fdedb96350f0b2343ca5023489d1
zb1d67abcb2ffe53799badb1667147fc149ffc4157bbce7e3dc2b3bd2ea8d2aeaec656d45b53931
z2f7bf1b48f3bfc534a01c845fe106fdeaf95a95ae26b907fb636bd16afa3300e0498b03df6e65c
zdd5e4e418222df7f4a103187edee1c6cb271ee9fb8e3823f23a7537cc4cba9d87a6dcfb283d2e2
z709e2faf6a51d485fa0111e822facf6cf1ee08225257e1123493b629c5197fe81d1851b5b3ee77
z727cc349c5d84fdf72fe100a4f374da3c24b755ea6af5112056593daf5e4d86445812c4a495cdf
z6d47bb9d84b19cbe7a2231a3a58b5dd5b9849e1d4b1bd63e32ab871322fad3da78839d9e6960ca
zd6b03f1f61265b7ce757a218691025bd6da0cc8e2fb912a4aeceeff7345da5c4adc2dd959db690
z588ce60ba79fff1a97093f8f21200ea1e0bb3663599e922346eb81a0b4c916ca6fd8b1a6fa84d2
zb188ddb917808ff00716b0a88d5c5eee3e9da2ab156aadd85cfa72f9ae4ac8752a71cd96660463
z7a7c1f123dbf9e3145eb42dae90943126bf8e4d7ff8a6dba952e150c6d8f2dfba769aeb737c24f
z4e72064319c2d6a64ec566e859fdc2b220242cbd630304391a99e9c811a97bdfcfb364442512cf
z84c6b82126248861cb5f12daf09a976bc475970cc7fdf39fd823b06306efc09c43dcf7054ea6e3
z326f10b60bcbae998325c1671856ef53a7c2d32f11da08e3cb0e4417272fb9b428b179c38e2432
z733ffaa9ec2642152c7159f1d9a2f0251343b5ff46f2f778a8b969ec02bb3897444dd87a95abe2
ze6f900f218dfba08d1a14bb4508c60e673a2130bbf5123a8acefe6506bf4bc536330894ced0aaa
za2d42706a1361aa327f68ba3f81aafe22003d62fddfc462cf4908c231aa461dfcb52f72e416ed7
z5b6f018aea8ebe5d885e63cc6d8526289676b03010b3a828502a868d4ea7c3354e5dfa81938f6e
zdff2d5da7db8e7b1173bdef72d0417d48e93aeab6362a755412ebfadf3b8e7b7aae2e8f3af1607
z2edbd83db9420117989b19ed7afb74c62f50803ef692de1569a6b0612659cacc53ab2c68674e03
zd97a4c64c7b670600e209c85ff85417db7a828ea117c565b23daece1061f334169d35515fb369c
z2467d35e0a1bee8a1e099ba571e4f2a81519944ea603276df5b047157f8c8ea835a7a8cb05ee6a
z91dc159dd474a952706d0455674822c2b91385e57284874b74ea148da94f254b4f9143a7cca671
z728c6dde60b88063cd997f9e35047ece9475a32cd8f2743acd165d8961fbdcea8de1e0879f273e
z581379fbcab32f772eee6be18428430d97fe20c2cd341a7d6a2b02c277fbe536867bad3f76b7d0
z62bb64f674a7433389ba84d7f9458eda592999c1e1e44302185cfd2a0a0471298cee2857a03306
z7039dff37af6f622c8215a536101f40b227794d80d5245ab6365e65a058fc0ba5f35dda49a15b3
z96a19206d142dafae0628e1f2d7878e02c353e709dc0dd077cbf3008025ae287890a7d5632fac8
zb139ddda06f1ee4a1d66c4609ee87bc1f0d585f644c3e4a095486f5ee8428db89dff49136672c2
zac659951ef9ac61fa57045194c78d0b54457a28e1be457440ece1e025c4f0f5cc4f4102f1f3961
z48e608ead9df427d28b78a7b44978b563b5183f0a3b16bb9a3060d73ce3c29a13b960d7f1e66a9
z3eac672bbc1649ab25ec56d0788eabe23cbbeff4b69c79dcde2d81a0b947802ec1a2ea8fead1e0
zc3e48d6999bb37f22daeefa0c25e9daa0703151be1e5952d53ed3e28f346449a41b2f077399ca1
z1b8f7a21dc8ee4a30f266e38e04f248f9905d0f4f2877e9b1c250782ff5f384281e365ba340f94
z1d10f16dbfb33946d53577c7e1d5f39df6e21d642ef91bb37ddb4c135086dc62b012b3e1c9a22a
za12fa5cf19c05ca1a6e221e3634d1471182a3e2c8615cd1f7edf4b9b3cc814cd955e8b74a3b4e2
zca54ee183a8ab20b5f4b3c41803d92e7be33d3206ca845eb606f958189a725a1bce640b82d678a
z08ddfca5176cb12c7239a97996e7e5614c51bd0e3f93f33f8d22c573b3ffd9724b9e821f789be2
z12b073ac0194a75ad880c4d49ea653e5ecf8855ab3dece1d38acbcd7bd0c922b5d48951a8487ac
z3bcbf31c030c9c75688c4dc564f810433ae250ffb9fdaa10955da179af6a8f7755c3ecd987b9ab
zebf4593b4071e2caf243f31b899a1ee82b76b2470cd7e76be46afbbb61c4ac15a649beaa16a7e9
z98b4a6d4a393f88bc00119cd2f047ab266b8b072b507a4046cf87d4df8c6cc94efab53ababe260
z59089dca3fd464722e151482297f55c283b8c54228f613405476ed354ebb49305b62e1e12ed970
z16508fc6d072fa400faa015b76fbdbea008323786dfc25779ff4c766ffa030b01636f950313eae
z33caf2a4b8f5255d936d3dbf7f991a688224b5d6b7f5eea6e350d3a6487fc7acb9d850d166d911
z70673594b493e446c2635a7307822824257b0cecde436423abdc6dd7c7d02abd3b11a690c5916d
ze512d7e9053883550d29bc3823a14e13761c72e348b7545a5273be963043e921419549fecc1107
z52a176112013d6ec4d617aec65666a0ad431ba0d306c4627866f4f4c6fa06daa0454a765dcb300
zd2390c0c53e65269fd7efb0902963d8acf5a48855511268d135c74aa19b14d2f07a3f1e6dbc7f9
z37f964c574ff6d37ff196486389be94b171253e8e1c71c0f791d74e70bc5c24baaf1f375b7b1d0
z04e424ce90793821bf093f45ff054590efd0966b1ca10c6522adbbf24f4470d9ee4a7a749db2a3
z7dfd5f559cd1ec13af039884aabdd1fa0a5d604496302bd51e9599f6b5309f4450976283c0dd2c
z19e72a8234259f5c7b6fdb2a6fb92b302508a8159f183eb2b464daf98a899f3fa44819b7c77ed1
z392344d68c0b7af8f3843dac4c8fb8198a72c1ac0cf8823a1f0dd87776cabda7c7199fe3feb083
ze19229bc46e5a7d8a37629cd53b3b9e8f824d364089f35f5a3a6755fb05a70781515fe418c5ec8
zcd353f86824c23e3b21aa1aed185cbbd04d6e74f7875a9b92317a21b44e27988d3d5433ae3ea2f
z749d44323ea5281607ba8bb2865d9d9819d54a8b6df4b02a17d61c92d339ee79aef9990a3c79a5
z4f51ddb2c2bd1fc8f1ea905921891b0f32c917b2e16ed3a3d02e65efabc0fe7357d7530d1a1a6a
zeeda286275b15ec9300b3a823f0b5fa3abbff3ee413db2455ccd7617b6587e506f373d96ee12b9
z64d1c2250760390bf455c9a5b2d7d90fd61e2a5682d59be0e89acae9a77183f4f0eaf22cabbf70
zf398b443d03b12c6866d4f97ea1ce84955ca62030e6896a2576ee69203d2fd7947bb39fab40897
zb0522405b46c0ccd94fbf77f8aec01ef5e27523d38ee74e31a632bb9242e5b283adf156b29750d
z855a97cbbc675350a814a5c8f186b6695f759c643651b8c3796bb5bd12fd6e6e2c3e4b88df07fc
zf16dd566fb552c86292cd5a1b8a3e375eb6508fef2f00b74b1eb59ee0f310d926391b4337a87b7
zb39770a8159541402c5fefa3425b04ce0cc9f7babe232e8fbf8ccfff2dadd4551dc84ef7a8d86b
z85c9180e46258bc8f53d8aa6e9a1d39768b1e936776376577ee925710a24719418243988deb9d5
z97ab8d7ca36280b35e9cd14c00a11bd3be3531700b3db479bc1d0e6ccda1c802c82915676bcb9f
z505d7c06a9500cafbd6c72a4d7acf6ac50ec968cbaf01b4dee6976fa750d1dda77406e68c0b1d9
z60c2783006ccfa54b83a370cbeb34a9eb85be53f8faf54326b22d9066f8da274f25f9b46acbf29
zb7b4ddcc96643f50f6567ac63416aac24a6b7cbf66b5e84756f2312da16c62b0b4a0c0db6c7297
zb9fca15e138b5aeca7f9611ef4d29c74673fe23665786a6e1a8741ec04dc733b4252eb52fa2fed
z4a89522db1b8f288b1c02f8815d25a8e4296406665765903210a344fba25cf05d7bc579282c745
z1f077bab455794733e1bc207e49cfa6a2ff63d8e5646c197c278a3ae31bf5a2e22fe773c6a0a9c
ze09c265bc1c36b3365efcea190b5f7a2371573b6a8ecc5a57edf8d83d6c34c431e7c5235a5a5ba
z201c128e9726671d63142c2d4aec98577f80059554dd070f4602c7cb0fbfe29bdcd152cd947be4
zfcf3ccd002b1e0b4efc39526fbd8ae6003fbb2561a01a6e343ef2a85bab8ca3463b7ae3c3a08b9
z072a5012d725b568ba4723c15cd01a22a7133e7b5598ef412765c6c6169144a827f682b0d85dfe
z6b4974c81343c7c1132cc40b026e412e34252aeb1f0825ca9970655c1d210f7e332dfaa74f566f
zddb2842e47733732b5f5eb3079fa3a6d3435f6f4d76a6d4ef1a2e7694ea55f6bfaf358fe1b607c
z920e2ebfe66020834fe14cf283e9de9ab9fc49c5dc52ba3f708f2af8bf8aebb64819576ed78dbe
zddd46574c24d4709ad38013000fffc27f480284949bea44479fc0dbacb94e922dc8040b3f81188
z5ec6059dcb770f145f77614c4825597f72e9a8d0b3bae257119a4ce3d7ebe8c180ef32151c2c3f
z9d70381b48b2e3d2f6d10f749a5045e23df5c87ad8563e6b86b8b6a78320ee1c985efbe196dad3
z83ac21265d67dc198fd712fd33830a765e791012653e6d7c41cbc721f07eeff7faf38fe55baa1a
z4e0ae20b95f1d0cdbd1dd1f44e9000bda08dfd7f8c1ec3acd6687332cf6f3bceaeba5e7ad20e26
z8b3d422e44a1baeb1ecaeb0ed0e2a5d18c64ba3bd31c719f718c20dc1c0cd7ed022a085d5fbff4
z948e359b8ed3c50fad5ec8fdefed8d07bfad6af49ecb33cd28f5239c3920d4060e1e236d5101da
z587067467de2e6cb9924559b26788b6b16a544b4ef9fe5db6b36a125b46a66c91d23b606fc1595
z49eb5f8df7e3c1d0526cd501d5787e68c3a0680190b248a81a04496a4234bda84f773ee72f4468
z09420f68ffc8331762aa8cbb341af1303c1b3eda38e2185ba028438e67222ba1c9a485c9867aff
z9829aa904641f44000c6b1dffc8f366f5b94618506f8df3ead7b0a20ae32fd3b37666b6e5a1f99
z80aec52b5c52346e908066be08952d4fc6c52d11a52a3d1c783204394e26f4eb044c06ae60ffd0
zc1c7cd8a1d97306d5f9d2f08f589207e46f7d8c7b4a9c7bcfa7227c6387d135e25dba53a19c15e
zf19d354cca6b6f6ce30019cb246c115a0161cc67e5dcac8d587c43269251e706e6fda8f9ae997f
z10e10e7a0bcaa009ad937afbb0332d922b339e0a7e197d653f67b31893ca86cc4c7d5041dd7531
zebe157bf37464fb21184af2eb1ab9b02ef3c636e19e65fe383361059728a5b9ffb7b2028c76751
z1ce099419fa52ee40c6cefe3f492893d37c7276de5b3e877d14a407d98997333958d3cdee7cc6b
z79c42daece21da3120ee23d2fe3c7c09be4fe46646da48c6daa7eef69139ad05552557d2c18792
z6476aae69f0e0e56aa2f5b3d3bbf47b3dc6f4dcd5fd311b2af159c753b7729fe44814e8065b517
z5a7dfceb14c2005f43293c64b235c05dc2bfed3f90917d783d40fbe5bcc549fdf35cb99abfa743
z473c5f0e700cb45c9a2f65675b7662cab4fd5a3d94f594b6c457f34384360bf7cce62a72bd5bed
zc1f6be2e13fabf6e1caf9cf8d78b5f13a940f8acac78659e3cc0d851ee13b68282da34e6f2dba2
zc3b9423f007d0609074f0347af27dd32c7b5ee25bbc1eac0873a15258e2d869d1c7d387e0f2ac0
zd79d9873d7b1c20ed7d5e838590f3135374d316237ae18175bfde4617a71c9074500ac3cf7bdb3
zdefafc35759672a281a8aa794e4907846f509c0ba78feec95e49d413c33656beda5a6b4966ea16
z29fde1eb5a015b8bbb4701a8b6204f3e5cdbfbd7d03afb6a23ac785d2bce2e934a0163d503bb6c
z3cf0fb031535cefd5e0f0723fed5ab0fef490895d09271eba553449c38ec54af52f50fc165be0a
ze307a1f78d109811c430491dab5b8d0cc31f38134a2e590290c2620c769d525c2175bcd21889f2
zd242c30402247dddcf33f243ce961084a35f3d89d09ddb415a4c9b152aee32d646c42b9e5c5ddd
z4ec7de0a8f506fc42a05870ff5f67046a93043ddc61e1c3563483c9e91bfaef2d0139b1f8321ce
ze4313fadbbfab5b3c9908d645c287f6068464597a8e05c4be1da3cfa7a27f5c6916e5da25da7eb
z070d33947ba14bd47c2e90bb6fa2215052741d41c9b6bd981eccd5034e97cab6ef042dd8d708d3
ze151c1525d9b4c4810a07301f3948114e83dd6d93146a6e3da5ed92483b8e3cbac6464d7157def
z6829122e3598cfe5af38cdc806311221ff0b95197acbccd93553a754be9de0e6efea75ccf89d10
z84479508c1dd7c068ab5c3263f1bb9c8b52b927d4ed0afe8c7c8d61ee4addc50846bf3be83c4b8
z4afb6ecb6521e748e45f09c48cd2604404f442ce765b69dfe2a1cd73259cff63c70db864c23e0a
zb4bda85c1de944b2349bc37ab2e7decf519301d2801af1474397b92619140a64928f2a27be8d31
z89970c00eaf7b3e2fb1286bd8d40577c8252d4d47010a4bc1dcf6d7fed6aedfdace87a95c09f89
z06f117f99dbbdc6e2cddd5d5a6a5aa4c47a67232a44397ae4a8eddab66ef1abc47eb9a1245c61c
zb3ac2f79bae5d56029bc22ab1988f8ba00575d6d63fde7468fdd544a2d4ba22dff2ebfffddaf6c
z952782ec3c1d2690c930ca375b015f055750138e5a9ea3a0098bcceabef525f55aa7a6a29014dd
z2879af39e5e073b390dcbb8cc275d7ce92dd3392daf0b9606830c1f28720080be0737b0e893d22
z378ade50600e0c907caf7cf8b9a47cdd51ab7681f08d53c255b4e526aee4e4b8da215545143f94
z65008a83f09a2b9ab698cc2202a71e4e2a7dbd65529139a4b4660f22cc503c403160d30c3f6c11
zf31258ac20f0ddca97c6bf4bf4749180a99b039c92502232351877059c67426a5b7b736a9dcc5c
z3416de486241c443ad5b4e66d6c075e52ad113cd0dee9b8a01f75cfbb9675c3c0b80f695928e51
ze3e51c2af9786add1219352e12276e3c55bc0b6a046d559cc53f7b355decb5f5fb35c85838a331
zf644a56db648d0e74e06b25f04f3477d4529c83b4b3a1b0a5eebc46ac4095c26e6e7889898b5a0
z7f5285352c332a9d79ed7e0eb4fbda7b3e8e99dfc6c54d37026a307ef896366fe483284f5326d3
z00d9d150a22c6340b2cb9269ab8f42609146b5bd362f67f8998a0a2b2c76cd159e7f9d92cdbe8a
z0a369914b2db61d3a6ae89570d3f89247bebf6893a70b8d9dbc27802fd18a5afca8d2c4645bb8f
zb2224bfa98c4cc44e680a3219e5dfe92d9ac626a9f71fa7802e17de1b6d0a091b8d401663cfe53
z3fa1105b8e7d033020d5d287c6ea5124107db5a162e2b1d1c66cd28c4f36459cbcf9db36c97aa4
z5fce468cde79e46cfba74a1c210eeae5ac079cfc15ac4a4948bec2ea8e4a881a212e1d50af50c8
z78acfa6ccc07bf03a41acdb7bdf33a74fce3e022602778ca28fecf3775fc2d00f9beb828f2bb20
zb70d3b404b4f718037aae6a2f4ad8c54e1061631128ce63892bb97e4432bbe5441c152245f5d0a
z7617904f1bbf72f43ee7965cb4dfa58036e1c46ea1da6c0dd5ae6e4226608c017257ad69f5a41f
z1f4ae710d46041daffe6ebd7058d940648175c89462cfa3012fa0d14897f554018a3d7b12b8c1e
z7a72bacfcdcdaee1e02cc4c28f29ce78b14d0b6361b6a7d84e2f96b144a2407c6393db323d3431
z06123720387a3ce4ec250568020e5653eab514b4356db8e7f93431b9d3c2569c8e9bf8983269c1
zbedf73925f7a79f49f5c5787df922a224a86e0a54e9ffac936468e2eaa74a08a8f1323f2cb8453
zcc59126a3ffdea5eb2d6e1b71a9c7651c3b95258aab8e42d720571532df53998596845f90bfb03
z809ba704d8d2d790596359f2c9b88c8fdb430955e0b1f360dec209380e0b48b53735c413b1992d
zcbf34d05288129a33e095939680b39eec456d58dbe8588f89ece2c73314e404426584fe1381fb4
z3951f1970ae6f11c7b112f961348e23b85f6f641ad13e2c3c48c18ad7eeae7e552f867e974334d
z09fcb9dab559daecd0202dd1748fe3c2b56df7b0de841a866e6bca58d4c3fe61ab75ddb89a1e32
zac13ae139b1412fc3d5c3fefb39c2918b5e333ea503a7f0bd1d07d243316131508e975ea6a1a45
z439101d0fbaa5c5f9291acc8a9104a892f7155dd4d495e3272e0500f8035a27d3cf66f0a7d7d60
zb15798e86c9f5439057cd00f372bbbeae5fee336a2be96ab0fa7bfac55855271d43b642825c10d
z66e15d31245a38f66357adecaf6eb29a7bc1264455e669d16be18b62b5e14673a148f3b0fc0441
z9985a7b2901bcf176fd7fa2d826f5613e569bd6f5deff3063af6c39cc1e5c029647e5ac5ff7860
z1c77f46931c76f5b7a4ea1791a8e01ed8588d5e06aafa355ae231e5a392f7e122ef9fb59a9ca39
zd6a12c0245080c20d77bd23fa31241f282bf26324f7b08c3eb519a7b327a7aa7fbb518e4b69d56
zccd2f0841992f76e763ca7be7ad066cd0fbb44a6b2d896686e4c624d0980e5b756a0031a9e2154
z2b848538f9c42fc7e2edf60f7f2d36eaae73826efa4bddd84bb517541414afb0ae0e98d4ccdd0a
ze80fcda64cb65c5b20e6665234a45e47f7ec6a05406b9dadc734910b71c220e301a3a1fefed1e9
z20cc0f733e1d6d4e8a66cd07b6c23de009da0f74ef52f0c80ee477dfe476565e2d841aec8ec60c
zec4d2dad2ee0ed91fb8b676866c79104787a7236303327e5a5efafed1cc6bf10c0fb06242d1407
zf118fa04548eabcc55903227b0d4afc6c838c3449eb788c23e4bfa48987e3650c337d6a27df7a8
z09ab418873654e792264da3fcdd7f6927e18f575c1a1839254145f31d7d6e7f23657a91a3ac8ae
z6b98d63f670d47d1bf3b228ac4dc15f4bd98292bb1385a9e460ed0a0e6171cf192aa57547eaf1a
z53fe8a87b9d81fa7c38a41c5df28c2f8b33933cefbb5fe5ada681757c4d802ec94394e226b0e50
z94edd3af438351f7bfd32a5f61518426213c37a66a3ed15f8cd04f90201515f7a43080edbdb238
zb691e28377a28f850b7b40a95884d6fd3dbe956245b38f25ea80a6cf8a4415b1699e0a8dd22b8d
z9f7ee0417ae17246e19484bfb464ab11364fa57ab78ec525da2433a9598dd60bb3608263f68bab
z5b7dbcfc8a854ea81bf4e4a85c7864a349a8a8a3db436e39f2ad60287f8f1a268ce2dd3c85f295
z2e7342f3c64394d2bc419a6e3beca886f6463238384c653a9738826954b6d577fc08c05040506c
z99b4503165af64f0ae1302e449a2d1fdcf787e0a3913231f244cee64b131c908808783313e274e
zfaa799032a92fc5d4f169877d840db9c9233428f51325f2ef625830b064aa842b118ac0934eebe
z380d756e09a6580f0399ca4cbdc615bc68783f4444548baf7b82132d2b8895ec160e7a15b12019
z8ac66ec8409f288c8d14961751e714b2e8f65e126df6ef85b7556415b38b435d8437aa0b506a41
za3ce37133c0a5dd634f00d3b61f67f013ff7b76fa2ee4c3d61c87c5f5b85ec6d43ad32624652f4
zad76047c6c6f766b066301d2b5afcbf1c966153f6e310e219a95ea3722217e84891fb0b9dd604b
z00f40391c1ea97a5f5156962b02adf4eb09ddfddf5a7ab519531d9e993b3209816f0039524c7b2
z258a180642510ff8ffce0b18db46c87ca84c27db6ce6df084ebb449ff5902ce935acad36334d6a
z933175d85781f05588fa6695f4c23d11255053725d267c2cf3984110e53bf3233dcf2ddd59ce7f
zf70eefcacf89fa158d2135b4179d890b1b0fa0b3aab290e582a6eef2c52188dca49001f0117b8d
z011c21f2a75b4578398c0ee19ba0d1b655be89fc090ab9bdacb2ab425b821d488c8d83cf91339d
z05884714a69f87cc270c17c3dda5d4becfa8bbac87fce800de4b99230e30a89c839f7215222c47
z732a054f66df8e8efb73e64779285569c001f448188d9827beeea5119ebbdb88c126d549e41fb3
z1c77febde79184bdb410d22643a24e56a92b804fcd1ebb63213d4ecf5ac553473fb6ba14b2eaf6
z88fb57e0ce04abe0cbb0e6f7d1cb80c6d01a69fab46f0ce2042db61bba143955b8480159f101cf
zcf360b55607587da1fc28499cd18b0d8c23c6fde83ac8fba2e1970dca105ebfb637d09df21f9d7
z8659db821aeee19bce89cdcf859a60f07dc42a731a3d8f65f03d8dcfb68f6bdff71936cdeefd68
z6c6219b28c8659c45c6d5c8ba5927e976f33fb2053f448becb7eeb216990b06cacbb2950ac05e4
z08c1662b132811f6dfa7031f91ff114af5eb4ca33de4b6c669d66fc8714cf30954d30a75f8529c
za000768276fa807884e165e52afe2eb12871769fed96e01b457070a8db9686d9ac1e7d93ce2646
z30a220cd493b728093729edd07a0ab0f59ab89e188891cbc740f989d35f5d10e41129d8782908c
zd7f8e85c4f6d55369eb3e913243adce688fa8d0d66c1d4dc06545e90ea5106958bf5e0099c18c7
z130d7b5eea83b07e61b32b5ed0d3d1525fc85f0b499dff02df4f2b67f2779a5cdbf57dabeff29d
z9b41228c35f51075b5831afb8818876c7d818b98248d7242e72db402c852f0940b099915143fcc
z9cd5f91887aecbbe43bb50303a0d35f3f2cbf28045801d7bf84054adfac74b8539ad79ea23db4a
z5c29ad962d4659d4dd6871ddab1e1f7d0f1bcfe054159c5e210bddad32ef2519bfd517482b2a31
z2cc8d76e4dfd26b639277fe494892e1a9177deb58e0a6401d15d39781d8ed93e9ddebdfd14e4a0
zc38ecf30dbc0627de7a04e3856627a1ee90f85e3421081758782efaa366de15dd547df5aa2a339
z6c023265bd807f7cb0700b70153b6e1f7bba7d0c0417eef2aa29320d2d00c4224ed53d61874c18
z2206c51d3d296f13e6d61b33e95d04975478a636f611ab65e885a281af055a478f850879864206
ze0f03dcd7caaeee07497da9447f250d3b2774253c1f794bbd73ca2d43fa65d36f4fcbe2203bfae
zea42d4f5c05ed18dbcc605e7992aae5c2133c523bf739c235a904af1a3bd9f3e6063319d54814a
za119804e1dbd0d6e06df9aa3e6ca8f4563f042357acc674f8742e3147db18cab33828c139777e6
z842f5d484b32b6b0f1aebe08d63f6e9e0c6cd1a98016e337cb4bba1d133e65b67c74c42a2f5fd6
zeb05599d9629008ef2ceb16ea90f97cb86d7856ddbb5aae6e10db8ae516b6026da50efb96a1f0b
zf471a6ef587c166520b784d410f985829ddad4e3d11e6fa59606a64532b0c39036590f2fddcb04
ze96f107b160bf1ca570d1a3cd270634192563f779e0b3abe19794614b3cb1c687c84a54cf4afe0
zabf4494b0fd1f321a0daf229fd3ac56da23fc8f4e89f2c79ad9f5535b5c2b38b28596737fef7aa
z131089c6592293e93835bc473b922e11e3b9c832fd423bdc6e62036931ad752082bad50b6db2c4
zaecfaf82717149ea71fd6890eac5abdbd77bd10c60b0b2d1a5690a9586f073e33044983961a338
z2ef9897b8bc1fd4384b709a0a1181e3291957cd52b7dd2a096252fffe832c5bd279728b5c9c696
ze1975977adc916d6090bb632b1803118dbcc505548a4d1ab8552a150874a133c002cb794dca57c
zd9817088d605199523d97b1cff473d29f8408137e7c95f26331cb463be714bd8c2a9eb7937b2b2
zb163ddc74e874920a172f429f6db8a73054fdaeb2d0aaed34f84be977f5aaec255f2d532aded9d
z0751de041127814c73063565939bb5d2b1060f3b980394597f86c9e2cb2cc73fd8f1defac49ff7
z0444c7540722ef32b482b5399a012bc49c6464acd5780d03d2a1514f73d724d1c022b920a31c11
z4c8be10b7f02327e7f700b5318673aa2da2e42a1ef1cd791d76d29a9a5838479b4350ea650f1b5
z048974ab785ec3b9700e0dc417b0aacb8fee737d7df033c91e04e93f1820b68daaa86a9341ff9b
z9b657c03f2a699baa09fa35a39fd624f5446b85c0696b8c9c98a989b30aea81cdc3fd948fbf4a0
z6aec675d7d3e63cf7803e05a2fcef10de9e6a044344e3515610a1e3b36373d2489b2812045caab
ze23f8d37e6f2066f01fb5b40bea7f728dcce9a5cf5de0ec0cf03ffe446bb48ef38dcf142bf0a78
z916032e6e69260477c797ae065afec695b96c5834e8946a2429d32934624d0d307ac9ccaac0588
z61244fa365408c56905a07ffa3af15ab0b44d4011df59eaa162efbc25f6b8a4fa03d0eafd28df5
z9c7b2f5281323354c6ffe45733f302465075e3f004fbb7b88862ae83ef918e6302c89c85c787b5
zccae1df983989a7aa042a72c7de62377c5c70fca43c3012e8b712bd78a8cd108b3ae4dcf46931a
zcf14bcf0f5c47b7d1f2b6dadedf8f44318fe72c6f207dd8c791f6e2811869e42d2cd572857151b
z7783868814f627883eaa3bb64fa2bfc43551101eb666f968664619c6b6f9dee791debe57e8a518
zc53ac77fc85687610a50d137d2f281c51f84663c7f90f384bf655939cb168c5655e562df53f835
ze7f177d78b87866a8c0710e52d0daf712756e5fe314b3f00fe4515f48290a025b874d216895e77
zca5d1f6aa0a6bc84c74817788e7aa3e14744af7e929abf7ac7f8d83befd75111e3d8fe58b17934
z8458d0900d3db94d3fa4886fc4022b8056343059a83039fdde3f2aba3722bf752fd62103eac981
z0468d0901b2dd23c5ad5497aa021697788416a354e9b10290b0f1190b28f628e23dcb45fef8e35
z332f7a8c1138483a8311f694785b447519a166efacac242593f27d78c5cd22311c16a45ee71588
zcc062f751e1e880edbc11d51decb92f24d55e43c6123340a5233e25b32573fcaeb2db7810c0374
zedf5fc3e5f43cd8213d34430736deb3bf3fcd54dd4c06a5281c9def616492e0655c4ec2cd966b8
zbd9692b834aa9effb16e52ef44bba6d017b8c63487159d88b2ae9d6a4990b987d37f22052c888b
z3ac5437dec727ecfcd40cea5abf9ca05cbf4ae4640cbcc69356ad61114f45600cba5fc2f405ea3
z8838e64bd85b23a79f2a925a5de6f03ae3cbe23909961413a60025d0e7d312206a585a6b5e87ad
z81cd468932aea6e3325b6fe1299c9f84a2bebb5a321a6291c015d6bad3b8685db15d2cee3a2ac8
z523f93ccf6b3cfa0725cbd608bc4e8ab6fa5e2f7e2919d73cb71eab5d97625354639c0926c23c0
z6686d2c1fec3b380c035a54d557b271cd8b45412048357bda97849572f9f15593a087ed0fe86b1
z9dde2ed78894ebdc668017dc845ac1f9e478cf6ba695a9683b5eb925b18478da76ce70ba1969f5
za205739ee164a862fcdf0b37b6e0edb9f32d55b0a02bc38ad4bde80b013268d8dead155ef73c83
z35567fc4a34816ffa4c702eb46e68bab2f1709f217d61536fba6956f22a86de2a1e03159b94801
z30fa54cb6f3ed8be6790915e4011bf72bb4aee82704be5cf1e7a42f01554ea3fc858868dcdeccb
z2412840a674726e8add97c42a3186dc9fceb42b780887f4d070d81f782378b84942498729581f1
z04b3919eed515490df7a205c80e791c79ca5e1f74d6fd340535128bc27b8ae54a98d11f94fc952
z4cc69da5c7133ac3a90cc7a22d0fb70a1e66815ad19b40f18be9520d81d7a71a27f7b3d0411426
z3617786a8d50b5b2f3b811e553ae9b19a9ddb90133bce41c84e8b8bd411486e46e9b9521091ef4
zd76f1c4e11d6425a6d499151bc0e931abd0fdcc88f3ec2c77148c2cadab7d596d9cc1e01770a79
zbbcb44aee8b07c152e8c871dced32cf6fa54b88d2135c93bad1b20ff54e27ff5b218e1549568df
z775f0532fbc80c35c9d071ff9fbfa8b096aee48d73d932e619f6f824f77cd57e2e9ffff5785eb6
z4bfa0b254970ab08e509fbad0d018b59b1a16bb5d8d28f54a6983d4710f66967909a1a608425f3
za4f066a1a43e673fd84851a29e8e122fb45dfcbacaedff63c821478af1d660e3d5b1010cde2268
zfb403bf5a730524f02b2499bb8c89acb6031b3036ef2e40b4be1775bee792dfd8ca59d56449137
z8b518d19ee4b47d23cbbf637efc085394223639006bf18665c799ae4db1c830dbfbea98259530e
zca366efd4f8c5d12f38d1d2422ccafebb7ab4893840938415ebc647004ceb09c375b7e3e096db0
z16681ffc017b376ac4afa2741e20e974b5f079fb1ebab323db01de874bca4c082a6bc299226fc2
z599fc3b32b4c94895db23732acc10eaec9e524db4c21b2392d40b725cf878fb18eb4d296624484
zfe6014bdda1af0ab174ece66300c9c7132e9a00849d6bfaed8cb38a7b3d7326aa112d7c3624836
z48b1ba7684a2c0e88ca77b99c5af2e169bb359c553a14491385607b7f12dd661f19ca60c721353
z4c3aa998fbcc2866eb596b5173eb2701f1b161d2084eba564384cf1a1051f48c2f5882c1ec44a5
z81b49336d4fc9bcf9d4037563b3299efc1a3e8aa27e337f5c4e09528f1e0202b549bb30c56956b
zd2a796889c63b6f414463cd4a896f71e9ff30ada88cdaff8ce6c7fb7a4b9ef31532a453876cae1
z8209bee17b59235b7fab96b9732e21c49f223a1c1ec777c5a1fa687eff9dd0933876469fdbd8b1
z09a800c999d145f3ebe61b1a243b396f6a3854d1f3eddfaf91d8e9487239b9203fae8fbcf36a22
zfd05e7f32b7a5ce6c7a6647cd88a89dbef069fa3c5a519f8a67834aa263dfadfab2f1dd8af2f2e
z56d03f87701f7a03c7f36ae0403eef95668f942de4fc10aa2debbe0af333edd3b9027c4b962cf5
z36599a990b7d6122d44f5470d0f3e8eee79c3da68c85dde2805e052904b4cf0c3edfa350725110
za285c812df4a9f0baf32d52999b177e33468abaf17fe0572cc148e43a1456edf9f16fe9ef70b2e
z592c37df755ae740b2b1e3ee70449ab33b6673fd506c31e8866d3eac247bdba095cbee842bf82e
z6575f49dd95f0c0c24b9bc4d26afae3d901523567cf5c6f113365f1ed18120ab929cf90cac14e4
zff61827791d3aba7ab459ce486ed1787ab8e117d21338a232b77bc5ef5d125f9388187a514a7c4
zbc847c3a9f1b0c8666d8eb65d324dfe5f0376688d26b682c50cfaa7d0371a857e8e6ab2b52fa6e
z697006b47a4dd5586606b6a9ace803504d092185c71c316015bc184152ad562b3f694481e0aa91
z5f38eef2687d8ebdd9939db0b808bb31f7587b4586d4a34a8b2a0009d40ead12b76c8cd903b2cb
z753c0d808e5a6ae2cee63a7e449cc51dbc320a2f1a9c925c49e4a8624ee4f7000adc1f88cba4b0
z6a786084257ccdb2d76e1c5d3b1b2e7a51759af7229713bbe99229bc56d69a1be0d09008070740
zd1cbe24bbc3bfb25ec561b9c48e0a9f872eaaad77237e727680e115ec21c181699f6ed40b43194
ze2c529754b0e98fa87f5d7f6a7e342476a23a1a2c75923ba5a707d57de8cfafabd9f41010dbb11
z72e2d2e1d516e94b3a93427402df2ced2405e91778a59c65f8c047bcaa589c7de438e48518650c
zc82be310092fd29650b02f250370b7013ba9089aa8de5d8fcc137afd1c90e05967da8051635fc5
z16dcfa9001e422507e5e5f0f5046d8af4a7f42bbe34f65b5b6cb12dacedb9d9aaa3eec572a0c0b
zad3f3d0ab2b29264d54ce7ff3975157259f183de76789fdbd86ae6b9a70f78ab35d4b3bfa238f3
zb2183f42faefad6afd6af21f921efe2ac93bf9fdfa225553f181b6feeb84fd8fe58aa1eed92b49
z830451d4ffc13b58f30c23c3ff609dbf7718dc7796dd73676786d9051957fa360f71862504ab07
zc07944229b6ddcc7bfb6f09f8e800802291218f2ab68df18522e000e0b307053e4c7b8f9a365a2
z7c222233f440cd9d434a69b6199c0496499769a5b037c3372a44e34c9848c4e45af869ca646f4f
z51146a0c32e2cdf1ff9e4842daae8e6490828a732eb3aead0d2515162a62f008db4fc98ddd4b66
z7bff7a80cdffadbbfe31e84f413a42fcfdb9f90cdf9f90b49e08523ac3d45c70e9791a761b2f79
za83956e1acb581ea54fdbd2069867f2e741f7a039d4ecf03943d39b2fc14e3c122ddfd0f67d9b7
za42a6fc0ae5b35389ba78f798f8400e5716b68d62e68400b4a07c973940f43ee26f5329c72ab63
z907d3e520c344c42046ae80a7417005374a90b6aab0695edcd9b40c9525264ae229b2a4f97c153
z88b7acccc34add57f47dddbec162d9a79c67098ffb747ed01a052095a4f2569a32e75d2aade5b8
z5c588b61a6cbc8f32e552e75d9dcf87bedbf97df05b355a41512392cd928880fbcdc3c7b27dc19
z4b8000a5b833db311795331f874f55e13f8912e5ddb021934bfc70f1718c0b0b2f735636fec909
z5862b86bb3f63434a301b33bde5978dc7188ba91c5a0e89e477f7c975c8d4c46a33c614bec6538
z406cee7c42be051e69be8cb0a055a924f4e17c90a99b427fe282d5c4fd92d02838ff254836667c
zd2e0ef97375a4130588737078580be1e6623c52169dcd86957f3c05e8b5c02dba37e2562423591
zc0c66e21c2f0c8c2a33419e8cd96ac7a364eaea5a91070b500a391ea0313a989026f55145071cf
z175bc967ee41ba7f9e6ca762086e9d2cabd2d28fe9fa118ca80dbe2adaea19f9f7650a22e16d9d
z105fae9022b2b45d71986d1ebf0b21bbeadb019b215e09192f85e3c34d5936c8c5b5df3d8bece7
z543875b914a12de7010602b328caf088ad8f46adb2d4d30a618a8cd78ec120b8f700d9a41190ab
z14de33de73137a649229808fcb11199bcddfb44b154129a6149d0b2160fe013e1b033f9a7271e9
zb1fb3d8bc36e3b7d70919fab6d2a488e96fa14caed03f3151d1f9d36fc13ce6209585685d67349
z5f38301d966446d0275cef094af76fd0be1e7ae3c493798d0a118e32e47e759bf4e8f082dc5566
z25ff2a9a55ddcbfa8d756f832d69d8442ca3f1bad13a5fa55e1191020537f043fc383f96e6edfe
z02472ac291bb5a0797721f867b5837ee9a59e30b675cc967cdce5f1e3e23e49dfc74cc2647ef7a
z3dde1fe2d2b3dc38675b79abbf87518307977738953b7e51508ce5be0ccaa0794f28b224e21ae8
z74949dcb9a7e0a48089c6fdb9aabb1bdefcdb772ceaa07c9aab309c173cc811324422d7c65612b
zb7a61c45b5348a94e13648bb467860b3c994b0da6c50a5475d1bd8d43fffb8e6548840da4861e4
ze081e4c7ad30907530a04cc99a21ddbca6d0452c8f83275f4b425dc483dfc18518a6cc13b2854d
z7f732b99a0ae0ebbbc9147be584953984fcae40937a55d4fe5cdde06d831285820eba5600819bf
z8132322c06dcaf870affc225579c4eff129fa813988327489ee4bf59cc42be5cc19ceed84a5456
zd06dd4f3ccb76db28a0e6d1f2b31f44fd340c138aa973ef45aad1ebc867ef711669f372ec833cf
z6606e61dbb853b0955b0a7b4091238e0604de7edb9a83ce4d33c1a9b6dbe2be3dd35fc3fa5ad05
zfb32eaadc8fa6e2f5563d889042b46ac6281abb368dae0084874b27ed67a05e4ffde090b1f39d3
z0a84d59275bdf65247aec7b3b9d013cf9f03069b87d623bd0580a1343ba799ce59165c4e9b5b84
zb31b501c12d826ce269dae60490fda9cf8ed0f7c72e861c2b159c4b98ca2659c43a66c5249baf0
z736bea1996245ece0ebbd2d9923e7e4c1d4822efa27fa06e8514199d11b5c83cbc14d30c470233
zfcf22faaa99378132b5f36757b91b45ecd37f2d5ddd889e9382dcca3bfb858a85abad1c904be12
z8793562dfdd669fb4d29bf78d174833a39313b43bfaeac4e054430ba220135b39c595c9d394f54
zd1885ce8f3cbe19ec4f4c1730e6995b6e5817df436c62274fa3c1f8dbcdb186205d324452ab58f
z99454cdb32cd6edb3f80d4c53024c2e126627a07ee9247ed10d89bb626cb1983a84d0456b4f426
z331e76dfc6a5b91a18f85293b3e62435848b0c808313e1c736223bb027e5940f19a2940a19d5f0
z13c3c606427a0fc09b2aa18317799f9360883fdbf9156657e2dfe4f5b131766f1b5991aa6403a9
z0ba958c9637764460797cd5f9b4010125e362bb63d202a2e8fb1e31505088598c6b86d728f13ae
z299ba05f01b3c2c287af4663b6ca5fa79e6c641241f4472a06503f47c8d4fe74ed4f1b04d01032
z2e000a395e8e1aa9c03ab9f7c95ed8b93ebcc88eea43c8b98120c6045b52328c6deda5d6a677ec
z057e373802bb5cf4dab4f812911d74c9ccbf7242f519498ef58405fcf1b81b108e2f0b23392adf
z2159a52278630a3f8d2c01adc9413b83f0408e6eb7cede072ef776ce73cd5f9556d109ee0e4996
z215c861f1719c85573631b5df3fbf1ff924dc884e40a9cf58768f4e5847306ee967d874b32b1fb
z2b4731da89f30cacd17b3fcd06b4cd43bf10e8ba8ff624896838a813c9748bd41eda38c4127cbf
z0c4faa93c1d9294367a97a052a28e8d7aab10e6f7ad47dfb801dc402853cedc540de45aeeec7cb
zfaf7e75ac2ac0846cddd13ce7cd214c6a35b148e0bc0fa2db55ac483c4d2db472d178ac327fd35
z755224cf1742f0daa812926d64dad4790b73059fb085ea954cc3c31a8bf5dc37f6bc8a5b4c8d31
z5b8c289623016b02765a53aad5778884552682aa7ad20dedbe30c78c5c81784931b27fbe4aa8af
z4f3fbb624e311158a848351c75dacc0134ef2f28a36fdb1a184f99a716d4cb2c96b2e00dda5a72
za8816db7952403474c87bc43b98359b65e290745e7f240ef1ce15c3dc6fae5fd3b9d249a09af3c
zae6c53677d51b9e72a4ab98ce68b8bdbd04a43e8c8413bbd363522aabfdfb9e1dba762b5a44f38
z7bfdc4567eecd5ac1dc5ffad75ce5e1403c1481f64905f1fb0d6eabe99635b3cd4600b2452ffeb
z53f4db793727bd56d7a4e21c9eea0a27c6236099c6b13e93538f751a669b76c61ee540ddf23497
z441792b84ea4bdcd48d3d70884193f5e4b0993f643536e85e24479be8a389a920d90c45e96da42
z94f1b9f1d7cfdaa4597ae89503b71d9758f783072f62cfa04ed3cceecd1b789a5132bac6c62006
z7cebe572c773f8f7e9afd75100dcd596428d0ab98dff7cd279a25acfe268213b9e1ed16517f8f6
zec5acb52505c4bb88d9b8c7202b8b2b8a1bc7d9f7dd1586eed8cb15ad7e66c87b7c2dd1c6d4130
z18fbc44d83bc16b497238adb3c7f779a8e676fd873ab2c78b344bb8847ea76444850f32d6bd052
za070496ec082d9ece19aedbac1fc2b1f473a9d3f7c6acb0d7ca9dbdc611758f540d37745329f33
z87f1704a2547b525b1ea009bd0d10cd740f513a2351a9ccf82efb43ee49e9232de497fc6c62005
z899e096a160f00c654d820cd0396b113146f830eb01993f936ed1f28522f2cc3d690c731f7aaf0
z31e15f266d26c084950ff49766031d05a8eece31feaf8fbfafc1b4796c6f6665021c136a4dbbe1
z8956f78a32749b7a7f50356626183d9b21c4e7a5f6be1381a51b3a01ec5659b78c427d44ebc621
z90b2d3dba818e5215afb0c89303a8fa33556dfc4d7f580fe52692197d4b08745b094db1687b28a
z195af7a14a90fa7ae2ae33946ad2ba26a12a4895c7896594d5e30ceef77571bef3466c669da056
z164fd2c363db71cf91d1c8a756cd23ab82ab020e100b748ab6c8c6f3764d228168eb761bae5710
z558f763c643c6368d99a7f5b5782b52fd1ecbf42dd2e98b66fb4f023e466b7ee7d6ecdcd0a9ee6
z5941a5b996fe44c9eaaccc1d858a39b916fa070a64a182caca214cf88edda87dac06cdabf21c79
z7e44155ae5e478550b9a99bdc18fce8cff9198f46fcb33f9853ad6082b9cce90c7830907764a2b
z0f3c6a1ba9bc268ae93b694358d3ee46ea79b4fe2b7162c8ad64d69d3e860d2bd8ce24c3043fce
zcb06aaee747ec38ca3ca8a9cbaa3cea6a292d1407a9b90ad1e109844738c987ec51e62056f1d23
z5434d0f3846bbcc742958849c8521aba9127c8cef2831e4539a2fc1df6a4389413130acfaa66ef
z48c547bb0e29fbe77e720b08fcf3d68b4808d90aa1d4b37212e47f4c68f56a472aeec170e46245
z3438cbf9335638704db05f6d85d4189dbc0f6ae3e4604031c2a6f8cd71ddd30614412c6d22ce62
z02eb47cf62c855a48648ed0b98e8ddbdc9817f2a1503f49d084aadc4673ed5d36c305eb535e8e3
za721c0cd512aadb78a40ad1bb9fd5330cf8fbd0304bfa87fa73db3fea9546059c571890f785fb2
za5c16c827abf071fe42dd8a92982c045a66c282e9cf1c609d06bef9f6dfd4c913d6f902df7cfb6
z5808c70c2005e3879d2445a71a48085f731d8a80b9489bbe164f21fa4298437033bd84667bb392
z3ffcb8f4cfd8621181671b7cab51a179ec85f3ec7effd05bef007b5f4c807d8b530375e25b1362
zb1bba372081b423f0054cb1e44fcab622bc6985f6a1918f4c3eeaa17db9d71b4b4a0a68295fb98
z2088f34f3c93089c94b5c1a0bc0db7868e64bf94c18fefcd0ce1c1d50d3e3a296d65c438081949
z6a9858e2d3065e60adcdd5392ab916c14e9ea0a9066661f48d0d813c45b5e11932a9669824c324
zef94385a0030ed56f058bbc8991c8d75dbb643c3e8f054413f4579fc849873d5a779fa93cd7016
z3f24960bf61f517a5b9ec37f96d65d24ccd34b22b7b3afb665e6d64918eff82bd01b5bc709f742
z8c26e59036cc545687106d152c4f5e94a9c2a1702e830495952b37658fff4243a4a724aa338226
z8119234c79b1726c5d67bbd452b3e269e47512367f2df28d500e95129f132c94446eee4aec3394
z5f84a2aad961c8161a01e9d2ae3d601c14696aecb06242da933f2152290469786e70e48dad4e77
z35173c8f33eb30236ab10af860c4d2ab9cced0b5943625a754da0d3e99f3da72e0bb9910ed9723
z2c54c23c8a914e9ec6e6bd3e47d1aceac247c8ee72e433b5708a03edc8d4ae39087238537ec9b5
z78e53ed51d7747e407c3c4cf46cba64cab1d142ba7d08cfdeb10389113a95de19843f3e2407786
zcd4126bc7e76bdd28ec5cec413af288919bfa57e8a862fbd9af47fa55ba3610717b26bc12b1aed
zc68289d6f0aedaa60b61a4f012cdef01d231e9f804ff30740a03b2032e47a2334bc4fa759616f8
z6258cced05a57812b41fe9997773c2fbc0c50952933d0f292d2a303e7d84b7f51faf70043e06c3
z87592d7f85697bee9cf50a9548f710221bfba340003140e92be80f69b14370ac47ac24488f9683
z6b9b1beb3f920a4ed9e35ef92ed8937101d8562860138e91fd1fa4bea80877a392ad1b83b13dad
z7c9e0c3931de6634dd76d7967bc1b8b3620a52c06a9f558fbf1b0322d6aa121319686f6b3313f6
z20ecb5b45c22ce07d6af4fed91314850fa4d16bb4123c459763c28255d8d911ded575d9eba98a2
z476f10a53fff2548083b55502a205e41d4fc37124440985904fe7e1c6dd4fbed9dcf8dfdd8fc6d
zd2b1b98830e4089f467e1b952f6813544f218581c976364cf1334b13d385b47ec9a82932ebbebb
z270de22a7e0ed1af81a6bb3913059edc97863e6e8b1420cd8d70297c55b64a3547f38307cd014d
zc5f385ad546e30055e049e109b4d7c7bc35653dc70ade36e4fd2a760929ad74253acc78c57c584
zc8fce7560101f0aa2bb289622f534c972ca35d27299deed23d80c37252f5c699f158353c248173
z165f2bdb7444b6fdb024150f82c4489df6a5dd74322d218e936c77247a305ed7f98353e49ba083
z5b0ec4889eb99574623ce74d81dcffc86eaeef69c795e274c662fbe66cc9dca05a0e0f9f398826
zd207c461ef056f3f86dfb890d13b522e6a2b43a2c1109c2cc4e4d1fc4ad49410a94d632a99dcb5
z7d351e23c3ccde4076121b25374b4cb5ab1c5a9bc768a3a1c640b6bb6660ebba80e2751f9441b2
z637494b65aa81148fa646fde06720fb51d69ba24d72ff3f9fa21ffbfc9dadd404dbe2c15283105
z1d8291df436dabaa8b9ee47f8bcc5f3b314180541b3c366f7b1f5a13d7f351524958c9f69be810
z62166d6b4fefeb5f4f54dff78b155ad871212d44de35384ade35b7da85e442cb64993cd6a4673b
z0e54a7e044e17e287591c42ca7229b10bc9612a5af6c0f99ca2c9ea956a25acdf77eea929b46e7
z8abd3582e30eb3abf4b4555c66c4a844a022d0f0b4060e7f9e0134ee26b9979d7606fd18dd9995
ze879160a6b752b42f73e4e8ce1b8378241a30f5de84efdf0a2ef3df8891736d157277d5a200f26
za52c8a7dfc57a98efaa3a159471818fe7e4dc8813b976c61fddcd0676a79113a5cd5274a88bbd5
z9db2e1bf8d33be71832d915f7d5970f7d574e5fb4ef15a32f8da01c6aeb88e68080808dc6f2caa
z87c219be1bae724eb6e3f876292cfb752d041589a6cc29cffd07d9f6444100c23785fee312cdd9
z66c5b7b6523c3ae119d06327bc73abeb02b36a26a30e71568b795f51dde91f4f61bfbee3bf00ff
z9b6d8540245d1b627d7bc1b183a2d0f3a6964c1a2cbb7d5d40002528a6325df3b7750fd0fb8d75
z3640c72eb800c2bfb2f860fcaaf1ce8684338d9463a8ec2a6426f536403cb9f42c4fafa684d743
z1c189ccef7fc4c74945272b92749aa99d0134335d64a10532cbf1cf26c64c413a69312afcb296c
zed841931c4d48d0bb7c3ace20395d46e08b902ae547b8654c53fccef9146d7205cbb1d52fb2dd8
zc05f94d0f52e6bc97c2cb35b49b23ec77eb8aa2481b72445bbf704c037ff76f620589d9c9d63dc
z53b8f2149cc51610367e78353489607c3e4a6790709539ddea62409a9df517f1d51640b805911d
z603215d00b82ed2dcb83b65a408a1d2c1ec947763ee614d587ef4293f9e49f10128783fce4b59a
z8f588efee1d3f234ecceef5194f3fda47be3c8b56a5103a7b83c47605c7f0d4cdc317dd909e64a
ze8eedcb39d2a32964e140ed57c13193e760e6e72c1d08b208f90fd74a7473f611bd11be8dda170
zdc216f8be9aff7628615d752687557c870b02d4bf91daa12167e5066127b51fc3b275ca8834869
ze41e95f6d2d652a571cfc153898b7546c87b6e2a91bbadf0bea17c0491cc6119d12fd38da3b47f
z0461b78a230c196a035a213e2b249667ca13cf1f9984acc37bfb39ab1b01300d2252b2ab1db88a
z0aebace35a2c4a30a158e5e8a68dc52053787d04c0e17019c61c2fa0a100c786e96b918d701685
ze16020b4d72288c3dfa368891a9df7b3508227c5b09c066fb3219968d022ce1ab21996858bc7c7
ze54baf8874adc35ee2504fcefd1bdcd0475d5c1a77a05a2bd4ef4eecd4ad1cfa3951f3ad7e5a7e
z31c91cf04f77bace4897d1b850ccd98805fd86a7ec32dab57e06d27ba7fef692ab060ce2e477c9
zf19da87ca115205e90aae86fc7348e482f5952d14439a9ce8c892bb68ffb3759001063536be6c9
za290358548ca7a6337a0f56bc6caadc2b8b8507ec85cb81fa852707f5a942371669960422e12f8
z9ebd4c7413600a349e79f4444fbc6628277fd1795222f9f697bb5c7fae0e20a777276cede746f8
z1db14eb27f7c28a9247d0f228b30586669bf7d103bd83faaf033d923b2ede11c9461f6bf68a015
z1a90ce9384d7404d7074e2e2d9a40abc97b15e1d6b2003c8f24078a8f97900024266d6ac688da2
zc845321cc20eb16020fae58d3fd1ff770d19e21bf2de7716b97606c925cd4ed8b1c3cc1748d955
z553839572d53ebc9da837db7d8443719f461da2e0593ad9ec9360236a736a93d806cbbf9c42901
z7fbe2d266d4c9df6ce16ea83d9cc81ff8eaa77d3cfcc0628a51ab36fed26b00903422bbc0dfccc
zf5de9658c4b4002e9e9dfc15c94ee836d12c3d402257aa71f9d400d0c135072f83fb8317c6dab6
z0074f8822986ac0c4c021147bfbb151c1c5fe8aa92fb30f19a0c4f819b276d06f0a4ef0cdb9a17
z04798a0a37b7b4ad7349f52de252e8d5d79691397887beb5549539936861c137e51ca8b9d3b4cd
zf637240b49cfa357e62422d4dc86903c06d8210a91ddeb801d7cf765161198043ee698b1544133
z55cbc9b87f5cc174876c728598eb13feda92707113741ebe274bdbd5b4ea97b025cedf8864ebde
z77943ffd8efd8a68440f8f63896a176428d7c66312e960029bd3f01d1406a030068cbb8b30d79a
z650195f7a629eadfb8dc51efe7d5cabe6b9a0867beb92b06aab0c8c4b3340ee3fa8978102eb881
zcb56c990a52a33ac71c7a0471e3d9618dd20a1f69109b8fd51d2599b837ef42d53931b05f0ab7b
ze08d60676a8be8a5e2e2a9bf2b0f432f5d8edc6abc04eab85a7962fb19f866821aa3ed4dd5495b
z9440e870af5fd2b7889a49aeb88276f4ab8335bd2a161365dbd863841df4b0063fff91f30a4a4b
z8121f982b520a2df33bad66073d0b1f571a98a05fcbf0023335ce553fe8b9d34d8dc05860e67a5
zed5a162a48b28b6efa11d4b594736e6567f3355b186eac96f5728342a9d3d419275c928b75100f
z21124a1991f174ecac234347898ffbe55ef3c79c7fb3dd60985754ff40d87f325dc4753768064b
zf0a790eb7195f38408cf603b76b12e045b235821b06079438f48b634889b6926de25a354e3a8d6
zcaff91450973f94a374f256fc19cb6cbc260e20727da628b88257e71861a9c3d1e2680fbe9970c
z1434a35e76debd9a871b532fcec3a00d3c7b6674b8b21034f6dc2e7ca2dd383296e1db1104fe52
zf0248868304f8d8d09fd0ff9dbd7213138a7ad19e6e4e1e327978076ea1cffc68853e2cda4969b
z36b545f1df35db9cf5549e9194bec2ac526981c2502104768dc4400502c42caed26a005763dc2e
z2c1d3b6e265e92a900782509bfeee5ff23281de85f686ce4a353406d08eac43dd9f1c953543634
zb2ab20369ca12e46a860fa50ee49c52f10ab12ecf35154af825b66db342c3d2fd55afc91384482
zd34b4a696e8196ab703c9c89554911d813589bd67e90b41dbbd2250c5a2ece24e1a57321150640
z0bf07a5de3b05d50c8c8eae7bf4d45b226705e0c6216f3bab244f30668a0bd6559b073358d1957
z619940ec9086baa6c9e6b7f2985d40a6d0f93fa312c5129ff9921fdf1235e49e507f4ce3d28594
z0478b23e0cbb6ebfb62c2fbe882358e872de7d87b290d8a3d41fc01f94fac6adcfdc592cea9953
z61b467a9ce576f8753256e7b64f8a0594edb64ffa2c53d42147f7ff837673d5cb88c54ac1c6aae
z08dd1e849d79664fb964ed1868fa54b8a692ff6bc630110671f11e34b03e892a6158c19c619ba0
z6b9bb2710e01835e4ccb43667b31f3f81c653206f5923a22a4b84791bef43c6e8400693412940a
za739256943b7f05d74530b6ac727214d4611ef17eaea66aedc3b8e6d95fcc0942e87228cb40be8
zdeec27968363a6079ef360ed321ca197dcec0c201b9544df512b41899423dbeb45fe9f5d921f8c
z192a06af1a199d495b190e20e377295919d65af5b7cffb6237580f70315d246fc84fa2b68390d1
z66e53fd4ee35863b5e2451a64db9feb0dce08cd2902c54886c45830f2b1cf29b2dffb7b3da9d3a
z5df7cddc69b28737f1e0058439a4b61c332cbd632140b4b31df2a1e34fbcd04696eb867e13aa53
z1ea258d6c4c09746c81923bc6304cb0568b86f74b0a04d58f787616e48687b467b15b4f4c903a1
za4b4240f2048a30b7186b81b6a3d92a2b168d64ed8dcecde9ba2f0e24f43099dcc0085d7e7263c
zcbc7022e81615d4e3eae1c223d5fe923e276b56384bb83cb725bce06f147f7f96c35c38157c464
z954f850dbf25d60c3437f0ccaf16b0b61965d0968da9c6970b036afa04d3451a609bf5efa279bf
zaf68b6863fa67d3182531cc32ffbbbfe72697d03a5cd8d965ac1f21ec417e0ca55d84dec12aea7
z4160e3c4a195d2b364c7a8015cf8ecd2204f9cbe97338338f051cb5fa2a5f05d944e8ea853367a
z3ebca236f3f917feccda22cf7dcdc567c2b1e10cc224eaa0e7daeff440d01c547404118e61f587
z6c0b05f06cd04d149156e322e9be5b0a161e6eaa3923c9645be7eb08784c212e62426e362aa5c7
zeef63beebffe6691af91fb28ebd1c00745ae117e3f6771421d3212fee620f3ee792d5a385864c0
z330246576c0ee502e21127feb12111459b5e69cc231cef7eb4dff85b9848540ea04036e5a91b82
zb8d9935713f7e0844668c2f33564e58cae420e1e6fd9bed0210f7b55b9e4cabfe8cbf6e63d6e06
zd4fb2c10fe0552338d051dcd0022511adad94ec8727008465c7dbe473f4fcc6398e1243b80741b
zd76b4e90a3cdd0f2db8a559fc80a191e12b5154be85d7fb975a79dededcf22c249226b94febfd1
z9093b32dee0916088c7d4835830d405e377ac1d2260d9bc108a9f62b73fb9d5a376c7e3a83b501
z58c8c58f9293f68c75ec0e10da61a64914132bcc10e2c726199c7630bd8ffa9c4350d7448bde4c
z9e4447f554e89e6afd32a9d08d38e5d1d353792ff7c92aa79847c85c264ff7593ba8b5d9a24b3e
z38f00f7390f4439bdc20e986491bf036e3a27e836dc10855561cb1ce9e7d3606d2f998d6b81464
z7d274882afd8850b54270e5ee03cf30b578f169af06025a1f5806c174ef74a9bd4955b99eecc73
z4ec1f12d5ebba401a3d6fb30d49c6c4c07f42088dcc0932561f8fbc516b2949c6668b09865a90d
z980f3fb9bf263101f76886c659dbf095a788d7d2155f8ffb119efcf3e45c789074c36a5b36d324
z1bd9280d1e27359813c77ddec4821cf6bec5c7a17966d5a89d87f29b1a468d80278451e51cafcb
zf13cb464ea0b4d6227a5aa68c7a887668f16180c0def85af27f133c60810c08bcbabec19e8b039
z1e847635be1a8f8ffee0da6ea9e125396035e34dee346982d4208243b87267a264e0d78be49480
z8fdcaf8f6f478d224b53de95202c4b4e5824dc6c7aece6b31df577e7b0c11eb44929e67d47ecf9
zc88d22cb47f5582783120417cb22c0a64f870ee53fda05ff885d2d2dd927d9338367d05264f3f2
z63d0cea8d030c2ed61dee823f8b9aa577711654f2aefec8200541e258cfe9560dc02148536294e
z6369406c78618cbb01a0a7305a5ef1f8770373728865c387e16766789090557d0c569947b43353
zd1d9734cfb67cc62d1a36af3aa2d5f3b45b1fbf3746ee6f928ab4ae6621a93b117cbe1ef2e2ec1
zf37e0467ccd814a4ee48d5a19056cc58f1346ab1cb906095661fe4b2e36ef699045725586f15ad
z7735f695ef480f33d51e3e6e6a1c5970cb0f3f7dd84aba18d1ff738638528dd5a1582fb7a5794c
z8aab731fca7e9b4309da85a6d858f4c3ce54e721d530c7880d04f3dd0adcb4597fa8b6b8b0cae5
zd92fe07ece48857c3c1066506dd779600f388a258cf81645753956356b719423cfbb6ab919944e
z19fafc732866dba14ebff52fad52cf0e734483c6fb911da4ae2d29982f1c8e26deb98b0dfed54c
zbc098ef286646270c2777f7081cb734742e50eb158b978d97b6a13e51274d776f3a154f5571730
zbe9d64f6afefa7cd26aa742e649e8ed742dbb52090d4d155d00086d40bc86f996fc38e97eac516
zac1c07efd59d2766baa87570956248cdee0ed9d480e311915983d78b84091cc160dbbc60fe51a7
z241f5a1084959981df7864b62f7264af70d923fd7eda18351db27cd7ecc410f59c5d2fef11509e
ze622fb13baa704f9d01ed693a0895e215678c746aa1ae7209b8d425ad92a69b92380ef934adb02
z18827634b3c020c34b278ee96287ee63d81fa31953bf9592afc1d003d275636c63a66a8ff4f5ff
z5d6f7df57694e1827cb1608722d1f1b245bb79070c2df83ce8327afe8150c41091a120b2ce77b0
z25b4bf76e6a2c0e66bbf8628bf9e7583a5177d7c3f6f2a6ce857020f91ead54d15466350543ce3
zbd38ba8ff2b9dbd0f837daa20de5f1137ba12f7e8b9a0bdf91789a324aee65254cd13ea28091ff
z889944ea62bd83afe18940599d0c9ebf4109d3eaab3c7a54ab0a212d5db1f6e70a316b40baff8e
z2cd1555b187f5385c33986820a160cdfe41d0fbaba2096b0ac7b21e60718fb92f339b9f5ad42be
z53763668e6edb45d5f93d3255c1ad343c48f87ddd314b067518ff9b02ee5ac0d14d9ea633803a0
z36a81a9c527597ccaebfd2e81540142bd1eae22981db420cbc28e9ea91a2889d30e895ee83b1c0
z47844c08b9ac248e17428cc5e8aa4dbbeb62f657db3e505a0649fd51f9563715b69e15de036241
z81e91f427c49c30763e6f3ec529ed02594227423165ea3f32bd639bf3d1a4909e35c1e5f1a349b
zb1a329afdc7d72da35eb284f6acee180dd6d6615f98b0ad490061b959ca22024915587fe865a28
z6379b7a154ba9ca619b9ae4a257bf24587e998f4eb634b67b96b34d1de24799b92e11748f82609
z52443965d529d687ea652d816080cd742461d11aad73da9a376d2baa4287a3ccb4d273e30db734
z6581a43bf7cbc801560a44ed17b3f07d23806967aa6ffe3ca3f1fb0ac8bbd9227381bc773b4c67
z622fdf83da599c86a5c91625b12e04c35822faf56ff466fcbc440151c007dcb27dac6aab45d86a
zc5222fdf42de25007584e028f591f076159dfba5e034a2b23dd03d3baee04439cfb4c19f118bdd
z845a048a94a59fe277c926d51d56c93bdb8c384102b871a0d5c243a54eb9aed5896aa5c87f2238
z4f2f450aa23371dc995e60d80e57840fb8964087c1422a2684735abdc2e04629720d0c05f0b9a0
z191b81babf19776f9d86cafdffad07213d94886c957644aded2651dd17fb6f6024703dd2e60ac7
z988f2e5105742a28028a8bbd9bfa6cd30bc6dd13792ae6db1e68f1d07a768e754899ae3c43e03e
z1ddb507206ade7c4e6302d12d65ea28bad285e793c014ba632728e3e45a82bdacf20ef0daa459d
zbb0fee2c91899fa474812e186ca8eb43316124beee0077fd075ce05d2b86eee727ee56325ca0e2
z36519e954a1f2912a8912e10144280c2d1f8747d30e5a9fcae631db48f4b80352d23277894ac3a
ze03594c8379ee229f4865fb82bef13de36b6269c821e6893654423382cd3065887a0cf5456b39a
ze2ae6552c14bf2934b644ac9b8dcb846934c22da6d6804221c8db48f6589ca15d42722a6a50295
ze6283d45f09be6505638240402015998f7daeee3565f02b2088d3056862384ffca5c555a2d6833
z43f60810c866a1a605bc5d7217bea01c0960ecd3182fa39ee3e53c87fbd7c41986d3405f09ed80
z6c3cee4591d3e0b3bff503ec5ff1068109ca602d096a77c21e661f0952d42c377dd24e2d4231c7
zf54b58e37483984ef6f5518a2fdf5a2accdb3416c1022021e6de4da5046721c214d145c291015d
z033b67063c89b22f9b286134e55e57749f95af31892db90d971811dcfcd5c3c419eca15c8e4730
z22bbc6e5e739de50f9d70d550643e117dc5ac9190d52064249a08f5c4912d80c4a3cca6970431c
z850be9adc090fba6e56ea9bd3dd9389baf81a42dfac8d0ce93f379a35c2c72e21a5f2128b3626d
zb005e948475eea35bd13a67245c46e0a57f83aebcdfe1d77631e701c94ebb95267d0db4065607a
z61ea0904c9ba270062ee7b5dce6b1804d66a2015dbd05aa4fd785b86401e93545c214f6c788ed5
z2732240ab106a9c02910b08bad4a666902ef0b0a79fa9c6afe435170ba2917368c0340fc339258
z32c8b58b0b94a67931c4351b838a2e57761d8475f42b0edcf5c844dba6da95803c6155286535c3
zcbef9051cfe8e87c30ab1216a23e171d19e3116c8f755b96901a775b7cda270f53458b657a7b6c
zf2e2bba1b59c1b73b9f0658434fe8d24fb9b8b3dd74526205683b487b615b38940c059a6ac45dc
za14a31ffb0a1cf13312602eff5dbbfe6f6541d203274ca49b88ddd3adb9a7452e13c119cf7029a
z89ef757b1f19e7d01695fcb26b0d7975fa66665a8f973cdd9d2d4566963204336389dcc3d66dc8
z6a976a96000b28e619af87d35ecde0b441b424dda7189d8b50036487372edeab6d242246e5e8f5
zaa38c5c75c6ab346f3e28bcd53145b83fae5f178d2224b31bbd83abad106d2aa572de80ff53ae9
zaedbe7dbea10e7fa6c29be360efcdfa5ea190c765677c4752c59a19182253696e050b01903e08d
za096498aeb39f47944ab109c1b0ee6dfbdcb703d794b6e55eda4eeca0ddfe23302d3685fe0dc61
zfd2ed5a341a445cf772118b4c83b3acc4d92703f739c791e66f2e877a6a83d1c0f732b6b7ee930
zf029ba06507b2edfe8419d1324edc1a3e6794ec94734341a091100c470c866385cc21b2293db78
zc2c477a7073b61084e7c28b1e109d48d3aa9cf2aef46d791f718856c8172e565d9fa1e26c8f7c2
zd4691bf38761c643244103d9048cd6f2391723cdec8f91c4ad47d683fddc37795c728713bae722
zcd434ec722488019fd946219664afa745b2d6c94f51c45d43c2c62de2072cace1d1d52bc466c93
z18a38b362e47e70f075cd42d12a9751523086a3bab1ccb3b58381afa6d2ad0d3671a71aa3daa66
z4dbea5593082d9f4ccb87f2615fe30f98e9b18a9a2d593ad1f1a566f69925a19103c2bf04d9491
zeb394fa074551464a3ec2cc759f3505b6a352218f235bf420dc2c736d8083668a68ad337c33c51
z2f86abb72bae5e28a94c076523ed62a342bd910e42100a6249460004f778c9e61506d4f76612d1
z8498364ec76f65d8e0f517245e326f887934ee53a25736debc61bdf8a54739500a14eb54e52674
ze56ac95dc225d61945cf79e8dee1f4b192d2614244c0f34bf2bf832c4cee1391cd7b4a5895086c
ze2c3a5daf843c5af77d827eb1326c480beb7e619798147012a32f3f9c667c202d5880b8b3a0753
z448a1b09acdac46dde6559945b187b7e32b97010a262aae8b3b4dacd162ae9ac491735bbf7352b
z75e40f40baa98b3108805a40cd926024babbfca4deac0732da980a05c540d85aa2a88c3d56d98b
z4c651ceb02a14489d840868bb0de6c1621ccff8a14a8f87c3703d5344eac566061cb98593b3d14
zc9e89ccf46a6e4923b2b408b7d8e3652e60d7f78d4aa82a85e3c8847a1f2a0dfad1ddb7b8dc34e
zb7dc5b9ab31542fdc02bc097d545f3eda557301a944f0500eec404111b5a351187a92d5679e852
zf481935e9c489a4a5fd1315d3be57054f7a5ed6c592ab12ec116f62a0100ed45d407468036c1d3
z575343801137655418c54bd2d88986ad0ce4a23ebbb473b49348998f53c19bfacb3eb82c243b54
z529bcb652ad01ee6634abe581a93a0ef22406bfda05abc4d42f8959ec7756bda8b74678e82fa39
za86828102e68a0ed1f2f3fec92b65e92d11ede60b656e5e8c2b34990cabd27a041e90950fd3707
z58c75748519997c0c45f19d4911c3ac47294bbf2c33ffaef26e0935458613886417fb124a657c7
z924d7dadcc1890f6b2112752f4033ea967e5b3b26a44bc5d1e6dc5f3cddbfd79ec0a35975d561f
z0f394683299052c231f427b7ce9de93e7b6e9c5f3c7aee9e41a16d14b5279bfe23cbdd81ccdac5
zee07c600ec9f3f7c4eb3a4dc285817c0c5c5a6b7b8d1bd729b5e874291ffb002a82c0553dcd927
z27b6e50a631518773a4183a5598876d175794bcdaccb6d6972ee94b7acae5fc96236873e549a56
zd6043444f55644bd11034c0b22902bf520bf1269b435636a202cc94aec7479300e748616b9627a
z8e97cc079d84525b531c61fa11271ffc66ceb26b0aedfdcc541f9ddd5769a8856b52535ede7689
z81ed534fd9767b47510772da9d0141abcfc437c9c3ca396756c3c731631ec4cdbc91a8daceeb4f
z2e87fb2b73e4021477b8415371b5dd609e205fe54b2c31e243794314d48964dfd60b45b8194665
z33378a2deb8b34659df6e1481ef60495dbf53fa25402bc428e03f3d30642645736c3a6e56bbc19
z49902c7c0eac5f5fdf62cab69ed787406a125c4b967a5947a7dbfff6fe9b3f4e7d2ffea9e27503
zadbffda4ab1b953d89d674a9a21b046d8897fa1c820d549fc063d2c49bba4893d96891e590047e
zac7c7f1d05801ffe5cbc74f83336fd2362467d198b7cbf2d44ee0f9427a4de918ecb18bc3a247e
z98b1bd967baf5337bcb50b031e43fabd7acb6faa7b2ac0fbff184e47183907a721f59e46671c3b
zd383b98d6fba71a45508d30f2ca8634d8e60aa5a3677881b926bc1fbdf84f1a987e88f05b61f3e
z6315a63231622e1618760538685584738bd9001c14d1a313bffc31f6dd6a3ce00bd692d042c193
za7385b2aef3595556ecd1831f284593782cab15d2acdc185d592c030f8e1beaf6aca96158a8fc2
z727fd5b553185773a6967d20b0771126dff05212ecb526e7073f7a5ad9a140a26ba4c259d3ede2
zd5751a75d847888e67a8724afc2a66db33ebcd5f343b6e8b6e6019afd21bbb066b931af902086e
z4d85eec0980b93b05b9822df36bed30721ed21ac9e8281613ee2ec045455dbf0aff87b6c00d03b
z9e0a95dad1b837e410756ab43cacd0e8c2f56fc6e3199d360670961260a44ad65cac6385990374
zcac1978f57450c9acec0f46fa61f971d16cab9d8d79e003b9f1e9cf821c0f7f69d896078a0e00b
z773167276e556ded3b0feb09af6e22f5df13882404e2cd76642b55dd2087a11c86253b78cdb9d6
zdadb2c06cbf9b3dce6d1222ca0f3fb04b1e37a263d6e8f50c2779329cb7373ac3bbc6c0732a7b8
zeb8db8639dbabb09b90865aeb0adc98de91c72a4e5b6ce673d4adb57618d0557f1fddc2d4c0207
ze0fcee783761c97655e21aae320e0eb1b2f50e33559f34641829629aa5cc0488521ae2168f165c
ze7968d66b51ec20ae5dade206f8302a0887981cb1ebdc74d0325e847d99f405b5df0f6b5e0677b
z163cff8690c05a2dcbdf4f94118011a02f6c2ee60988da39b5a31ec52b6e272cbfa89dd5f4a0b8
za042570828b3cd52a420e243af4ca3624ccc79a26cebd9cc7f1c26ef8121087eb766e479dc24ff
zdeabd40ec06513ff15fbec94c6175541b7320573cb0507e7a1ad81b12db122a91b8cd24d88a510
zb4e86154911f95ca0a221cbe332324fe2b036e623b5b608776f24fa62f1dd0756f2b7a952e7461
z66d6b25b627654f857c137705de88250fa605e2b23f3b67ef48eb7a51047a4a933c9ba8785d13f
zb07ace54bdf990e42b608408e79f067a52ab62ee0fdc642c7cdcd6db47e0d79c18d3c7a4b49a96
z44e30aef431fd7b08492fbe9f1f931662c8d25594f69773c795354d5dc57394ee0090c539b7c1c
za841bb39f41ef44dcba2f342dfc91c641e2bda5a72bd431c1e532e77d938cd960b1442562eb74c
z96a0507c7995bdc2db53a588399bbeb1d3da2b989745ccbc4a4b686c41e9e73159b3d9b8c7fb95
z960ca5fae6dd2074821327bad4eceff093b862ad412d620a83786d7307966953c6c1cb109816af
z4eef67e92e8aa962bc9fdd98c76a038ccc537db660d3499a03d7e2ec10425d8cc9dcbf1c44f4d2
z1b2bac2c3238c24e4b7450241d23ddab7974d8bebf8b4ed93b27eb26c4f1f95fa151ab618b81e8
zc5b03b25608cbe929374bd302534dfc197892d05beb9c8937376fa7830b6fce8a939e6264d57ed
z5bbf0f4141bdc55b4450b55a3386dca49840b932245929949907c4912d38a7627d28a2d38d5e02
zd8b2e66adbb93d9dbda080c295a930e50f50c78ecb754709608b7c7cbabbbcf7c6079e8afaa6ad
zf563a519704873e04af488d4a03b731930ef0d46182274533e5ee73f72ea09f43812f03f5cae38
ze51a43415377ff65acbfa9d81356cb39f3a3c3e2c060b3f11cedcfb3b1dbf3ea9baaa8ff44c573
z47271ccaeae193b034ea6c49c07788316c2b6f1e67f237245d524187b75e0b8f26094502b9b309
zaa7d67931c73cbcacc5a4934e6ad33e75992b8f5d94940b8fc3c5b75511b10c59863e43470f514
z594e2dab0376f822e0f2367506176096640c5ddef42f94c44ac914e9826647bf1a75a792503042
za4b289c0830bfc995b3763859370e1399dca886025022d81a323d174e2dc1ee0df41ce85e8208b
z44879f9db8443554800dc3d36f33e874fef02e81a82e34af294199ba4defa726c2114982dbca53
zeb0165dcac1fc972ea9f9c444e7f2d0c8ae3f6fd5f235d6873a2fa690fa9df2a78019bf396fa84
z5b9cbb19286796f00246151fb71520ea38f59f56e1c0d28616229e216e734d20ee119cf936a4a3
z8f876379a1a0a5728476f1db84710a1ffc8ac8f1747245fb0346d7b136a367d2c4d39f1e692824
z88e332360a3e3d95361f961e8b880921549d5e3dbfb6485fe7e80832d83b8e27d396f9c340a2a6
z7423804c1aaec3b181277b0d93e58d7e0710d54b395868ea9f9b9b1a3eb68d32983ef6b058c6a4
z90d639a9b2b7ef980b5bdb1fa427ebb6246a9e3348eeea1b36be06535e97ea3ae9801ede69978a
z42bec32a514d12a2708c140f834e1880c47517771ce7d26da5a98b2a66b08e3cc5607d3e643c2a
z1c4373b3fb93b56dae94eeb3e7a6238f7c188d2cc4aef06da082bca4affe5146d6d72539c99a0a
zf8733a42ee3b43d1318aa25c7816a0777a217018e1000c3a242f331b1bc157ec7de14c60ef74df
ze2d29207f1a0c452fc9dc33cad55e2f25be4c3f8865333b26095b2477edeb43aed1044b7090f40
zaf4d02e00c7f4cf1cc6214f183b2fc0987d9639fa649813a2b030ce1d0d5bffcadc8cae5c17257
ze61b6bcc34aa8bfc03212ee0ec101a77594ebd416769a536f797b3fe1a3b42b8c09c5f071ee100
z227ceed96489eaabf2b6c317dda5e041035cb3cc5f4e3c5d83169867f4d93200bb002dc756f6fd
zc1d510bf16f59b8b94c6f2b36048e4725494e00d51f2eec247d32757c0da2475bb924000edde3e
z5a82dfaa9aff6f53ef7cef0a7d73c66ba2046936514c76050ffc18be9e5909c863eb2f69904418
z93ef9ce054baf602074484fae26db5a9999247ae75f502805310926768ec6eae03a001b5a6d8d7
z42dbddc1c124abcbccdb86b2757b82c7341e6068241489450b7bd1aab630bf55e9f24d589c29eb
ze72954b5fa103e801bbb5a08a4359f17747c5ad05aa08c43dea467cc9b635fdf06d67941e365e2
z1a7896a498ee12e1086f3563a662b87104f209bdcd6d448e92da55ac95786dba044204f5caa130
z5f61c86411975347bded3d7626b29fd88b97ab41468ae39687ec89721ac56170a001408c15aa5c
za985c80f669f6260a8ec678623a188245ccd6a48628805ffe40fe242192eb6365c76f5e9e31689
za6c3b999ca275acc3bad9f9c86e78113108fc75d157d913caedb6285b70b928ff7f9079f8ad402
z8cc64d42bbcb13c7cc8ea96bb409f2ee34ef595f77b55e219a89ae7775101aa475291339290c88
zefe8c6b8f7b1bacddcb3415dad685ea296884891c6a7cc354d67f58b32c480a916bfd766316b31
ze1477210e3be3270c8c4a49828290080e0a26dec6a2da81262cf5f6b99ab643e266b54b0fb2879
zcb817b0795d32c887da4e2a9bf855b836166ccf70094df4f867ab2796b3e8f2d468db35f5a2d3e
zf27e53144439dd3520942fda68c6e358b8c1c7dcae1af38e38fd0f7ad35daf585ca01b011e60da
z06b62b4b242c72dddef8bb3dbc5f257f06072313836d70b36f66f97a1741eae0b5329b2db3ba42
z9aa2450bb411b0cbfc7faae12fcc6f5ecb7ec9635af2415fa29997452c2a838f5f7901ac84f1d9
zba9a9c833be8a4bee227baaceeb99c7f34c7f073ffe82bf0d29e5e2c4fa1cffb8a451e177f083f
zf1d70f84f574d22be16eb703204ab8357aadc65eb243bab8878494857b86a32043b3e3a73cb13e
zcaffe97e8984a92601e6615fb74a494b83046516a3cc99c69417f93d9a41c5aca12f0af83cfc52
z1d1af0596b948afaafd225eb656489a095b7744d58e86254204b89ab25b7a6488df92f55c3d64b
ze0d92e95b4d7bb0d3bcce589b16969af23d7a0ac5184cc93077f82a0abbf5083cc5e81ee31c765
z223aded853808128774aa6d278a634f4ec78912fa62e3daf079e5931e360d28d31ba68fc268d81
z4626f25e158c11381f43efde7e50a867c4712e39733d09fbca410a1d18c26e84043623a72023cd
z5ddf3638fb6e9fc11e6fb383115fd6f3cdb5eabe166346c0cb8d354fae00c9a3f1ebe3231074ba
z40fbdf0279751a44b0cd4864e1367140e47ce7f93b7f3aceee7b1bec370dd7d8719b74d175a126
z650dd08767a725fd2b80c74ca84fc457ee811afbbda489a1d3a0cede60a9f29e363ee602cffa95
za19e3ff9a6b44c732c4c0791a83679939d9abb323d2eec9a0677310f3f333003b15b66c29dc3fc
z72233ec24338272339e59c96c0fd8ed9f6cfd671a1cd2001c8ac80955670432dfe5120a9e7ac50
zcbc823d29d8616b5e6aab7080a033bd17487686d3777c395bacfc34ffdbbf9335d1c6cfd363eb6
zacb0d9a7842a91bdc6ef42ccc1cf8dc7966f51d44686a4aff20a0b7a7e5e8782e9b7099241de7f
zc1c24c64d99c376b985fab8a446823c81664b05d4c52336243752c9577d0cac6e19c5488da5d49
z813d5cf1aa51e5c105e5aded255847ea5a3ba4b7497c355bec36fffb487caab3d9f3cd6af4778b
z77107b49d25b4414f181de3a24d5e6b31d15ce9e4dbdced834e9a3d4436527a4c3ceb95a6f50c3
z92e375e57cb4fef156e6a39b76ce1e6686edf82a43a2d5316cd769df3658733ba81aa8e942f2c1
z9707652f2f9414d97997df338736bb969c26d7d314fda2ddbc9fb1aa7f2dc56744f64412941566
z6612e46b59f5ea328a2422fc9fb858f425da217d069e1a11686366c7981ccf57a02cc47eac8805
zfc53dc357a224022cfdb0ca4ad5a9774bdbc5d99da10ebd4a94ce6822d9219d1d35841ce9ddc38
zc239cdb4fb67c20eb377fb0e65041ea764869449e984df8458877b55e6ca56dfdd7aaeefc07f12
ze403b5f7e29bcb040e507cdb86bd15076f9074edbb5ad1cba14ffe16ffd204a040317c58086eab
z3c44029b28b92275902b0841fd66514b50bb1ee2396d9ff13b9b29196d55b7fb65502cd744ec4f
zbc8d41a613aba60cdb431d00663e9e4d5484ca32d17cb2228346b9285b7952d861b1a15029d3af
za16d3036e2d9d53c55b9ccff09096bee07ebf55e74ff87937b608f9c5d02a315f18e87808e85ce
z6e3829baa9843af392c1937354a02824e26e3627aa9c9105a365f249ef85a1ebb7813e690cfb8e
ze3d07ab31bdae115f27e8a2d5f72325cd44b40301ec46f7bed1bf41f9d01f8d62d739275229ee1
z159f13ad41c1bdceef508d4a6948865263a51c0b9fe59a9c1be5adba03c4ecb9b0b514012cd424
z7d6da6374cc019e811206ccef3264d2f551fc9dfd763551657f7385029f1a0a288f93f4bb49858
z1685c398505f5c986d71fd38ccc274f713c269da9adeec7b86378ef7e069d23b226ded84f4225a
z358c617a9c8a60649c0e0ce517595a14a73fdba99d3799f4d9561c815f2bf03485478628f5405f
z6e7b2836cf58372e0f493d46cf70934ccbd64e90903b2f391b9d34cf7cc85b2d0e95f7d73fd63e
z5fc005e3021bbf61ac323af4858f8db222d67b8d506888359fd92bf9586eb51e601a760a9f3fd7
z760ce0a1325d47f120065bf8a9dd8ca5f7f7e68209fe522a32342bb4c1e128394576d36a7ae6d7
z6d57ba00d99e1e8d4f8daaeeb29b54e88761ab4511fb2fdee2b3dfd09b25be84ba5f3deac4f6ed
za33d9b6be6b3d41b530c07d6ae25251a32ca284aab871547290634099a3ccfaf402763cca736db
za78cc4064438cae19dafbbef2f54c10b3ca2238cdb97096f5a44a4107994d7f4f7eafc4bf38386
z592e50cdf9e6f75b181878ab66f23662c808e6422cb6e1dc612e159169aea8989adee7a5548da1
z0ef7440d0e44afaee45fa703a713f8d8a06ed5f7cd24570210aa2b58e8cccd73ae539398d6322e
ze8a6ca48a41b6c7c8c3464a3c7fb7d543b6043b1322a37564be395b9c0aa4eec73cefce2bd67b2
z9460f76e77e82f18f1d8086ee3bceb959e43a4ae401d1df26b0258d12922d0a98d6c679ac7bcfa
za2126fec4aec992a3dfb16c44982b284b9b943ac6df0be4145337bd6ead64ba1c981decb2621ec
z0cb6d7f13f41bb45add0f9b47e292edc1c4d6b975eadc966507649fc93a1c1ea04795685f518d8
z6b7b40a48f2166822563398cd5de8060082a1c4e8b70063a3b69f804cf1ef587d4bbab069464ed
z0c4d1ea7008d84efcdd57f8920dd8c995d397622907a277e8ac8ce08b85dcd057ec171fbb94096
zde3e4f511fa25bba45d4daea7955b0bb741ec70fb37f9839ea1cc267cb9b4d606c5896b62cf67e
z456a47ef0ef30c6c27a5434fb26b85b531223c6bc775c1457ec475721bbbeae294b1cafc921995
zdd298d2315f5afce07ba2b85f616a96273f86055d8c56f12876eadfd22b9d754084ff8019389d8
z827d30df03bc01fd2eba0a0421c3e7c4f7132d5e9cebdbb8d6b4b22688aed40dadd36d762aa318
z6ed74cbd6f2691f813e74687accb7fff5f73dc90a1bc23aa6c5db63fd4495922d90c530ae6f283
zb290741c680327d0ab1bc8c703c389dce232923d839ab93e41df4d390d60ecd9c67acfdf39d3c2
z1319c0f423dfbcb309e79ab5166338a67b4c76f6a529b3d1461d83c85a3361a5eaa093f2ef09bb
z807171898892322f7477cdf3cc51ba0f5899ce35f48014aaf17255a18ee2964a7e59468f216968
zc393f327089552e03701975dd3da5d63ead8e0f304747f80e0e23f374085b7dca5468f1281fd82
z1ba11fa14f8bf55d77fff59d80e55c0b8944b452f57eaf0801685058b5fe2f3d6a76fce7c8f537
z1936332ed4c3d2d55ea563b32878c2f866ee6d03f0c593948c68541013d0d6eb3791460e7dfa52
z2800ab53895f31b6217c0499c384262ced6e1c1f4f16e7f42728eb7a3f076a8b9695bb093f32de
z2669e658220b8f1f51662fcd9c0793d51cd678511d8a243c2cfafa113e32440d77d8211a514d7a
z041df448ab6ad504c93b5029414bbe9b58faf4608a978bc5c79e88fdfdb52f02724312e13a3f50
zb3bb6ed3a7f9cf3c6ca72553d9a0335281f47dad9f29fcc46fce14f006663a2d0a029013fa4bdd
zfea14d2dc295412eea648d09a18128afec4dc2898c79a02cc5ff38cb61779f2f55c4b1539fe50d
z1735094f7ce6f68d035de51351f0eabcbeb04687fe39ecf7a89d80ba9ac6293de115c7737ac4a9
z93302da8a8df43e78e2f2c04ed567c3c582a69545c3d819d1ce74787a48e51ce83bd7579aeae30
ze3ecf406ed3351c9415cef777b2586184425c5609d24cf8dd02845e08b12c69a7803881c9d23f8
za7f6c51739a00dce01833ba0a79617147dcd17577fe706339a8752e6f7a0e66419cf719d6594ab
z15b895958e142ba726d8f098882d21e0bce55fcd1da24610d3e93faf15a3c04f33a6949652782a
z11dbe6c1931e3e5c8336f65a4061cda87dd9fe6544b00845a7fd72ef52309c6a184c5638b75dce
z6d681154f1527a30725fbf94a638bd11cf56e75ca5b530f4aa34a435247b3db550a1e043d180e1
z2b7f58e0f348b5c5cbe86a88dad1e2a7ff7ebba80fa5a4b7527bccc64d3e60668287b0fe922fde
zebe85f2c36cedd67d0d8b861c71c711e8152b348f30bf36cc52e6729d90dcdb7103f99cfbf4672
z09f7147838202e56ac41760cf514dbeabf7dd9438ce0760dc7c7436d92a659c522978d02959500
z87a0d830715cbf9cdd9e255b04ff694ab3cfb62cf4fd49aecdf55ee7e31af9e0b9a7e9fdde6c32
zf9d4bf31e9aaee069609cac9566948fde4ef4305540504b7ebbf17e0e9384de0ea4dfbd1060ef8
zb29224747d7349f3a2c51691fb27a9c943af4c62e2ea305e7f6a3788518c138323902f0083aee7
zce1ea95109391b6534fc328f1d69a3bd32f679acdb187c6b20f917f4e7221d24eb0eed23f2e012
z01a8fed9d5391f7c34127942eb135a7bba0521b414416300e7636f33a8796618264234437a8003
z167c1fc0fdc72905cc06be5a59fae0ac1924ff321337a7ad8d5c74b0f600715d41813241acb51f
za4ba07962277a5695abf5edbc35329dde75bfd3ccdc195e99201ecccb4c724fa6d7df06cd8a971
zd712fc47cd99fb3513edeb3745a0a5254e7da664010ad161be15eae9c2077ad3724de0e931eb25
z1118a5fb74c05dfbd9f412942af92d350ab3cbc78a3cd41a8ada8c767b93bfedb5a05e97b4c362
z2a0c53b1f1ebfbb8888f65c590f841d40178c5334fd06cee59308caa512373c1ed2bffa45218a7
zd010a7beda1c1854f6f4c8f5a958197289982d2858f8828f990664972ff11a3a51587abc33f751
z5fa1bbd16543f8cbd4cd5fafb9d90d69b90feadb33d5b69126bced8aa41ddf5809e498852e21bc
zd263226be601f984e71a9559cdcb51d959c74eb8a1a812fed6798ce11f77ced40920ae15577092
z07868dac9749e3528b710e044391e77453c768c9f7cbfb87db3187219b3d893aa8d9aab825aa5b
zaa3e27ef7bf177b824e7abbaad8e96a4e38c91997e07b20e9d61a2f8bed2103b9a4796286058a5
za221a0fc809a88c021ac6a23dae5a6752b526e530787241eef42089a9f6c1ab09804dc7875939f
zb2a05ada72f08100906ab1d49b8ef8efd8028362a25e00325f4aa7fd4c7a19047d62125a873e02
z6ecaec3e1a51bed3f050e193614f9031e9b54a320852510c167a5b834c149054d9a15bd546479b
z27c2139b14045a6d2605173d654e00c2436b5d9ffcd8e2f1874048e29b442fa9051b97b992f41e
z26fb310242d9c59ce57dee0483f778a7780d970cf6a2b82e020ad5956b66804c69b4adc02aa716
z33dde127bf94094c311331535df578cc15fd5cd48b44e1afe7b88e0bdeb9ae20f4490b7d58c617
zf2d606b07d27d16112b481f35773613896ce24cd22e819cea61c2b80f46050f6c0b81ca6c0285b
z1b5303e9f332cad6621be4adfb991596372954bdc336149b69c2c73df89c9503ce7d1e0aa905b4
zf89db35d20f10ee178991d7219cfeb99c45ecf93d523b269289bfed697dcd24c743423e9a0de87
zc41509b04feb4da0596930956a7b7e70700bc5481984c64885fa7803be09083a892342d2cf5bfc
zb375628de31fe938ae6aac37b17aec612c8b8d9e5c2cc52cd2f734557ce84dc3ebe15fa8ede975
z0a33e3e2e417700d44f9023542428e88f7a7b55725f7cba0bba7c4c83a953c147fa40bf1ef5177
z353ccb7ccd53901ea7ccebba987e2b3f6902f8779d7c40c731233cb82e6402ae3049b2e1044923
z12b9ada02a310767c11f5a02c75dc4da916c131fc8f02638749fe309d552bf095973d5dfd0958f
zfaa448bad5f330d8ebc69eada25757a00da3dfa886b527057d0335eca172d5e44c18fb45b31c22
z44a17523bde60edc93ca59b5cc08ec607a99da753c67ed5c7255dd8f92cfa4bf9a12e2583fe9fd
z60e015e1702e3ce7f5b226bd427ccb0c10ad7541d4c0ef3a5c9c28621ddb50172393bbed3e37d5
z71e03d5396193f795cd217c0c51f934d1f35621ef4b2ec545b92795efd3d668ed1c7784b0f79d9
z05eeeec4e0b42a1cf654603802d28e4ab619f3a736bd5b0063208bdcd953713ffc109f27f1c090
z78046c186ac9e4fa8f39d3d06656715e0a8c0ab2f26342beb488fed83ee0676e05db30c4f11a51
z51fdae89688c9d6855307ec45b14d5f8572e959104ceecb2879ba753e38855e90f0d5b2df3566e
z0bb6f9a1c55c9221f15bab0e3876a6f05e88d045f199527cfd871191b826539f932abcfe849c3b
zb90f92bfcf07ff4fd7e0388fbaeac9c7b27bbd3d8d5200e29699caaee349a928a0aea97e9e4733
za2e20346372e07e753f27723d7909165d1fe10e9b5cddef257f83956ac51a8ba8b4dea07b15c27
z3107a43fd73150ea5f67fdea7c7868f81892de43f15370d4436123c3df9d9c67aa2c1a1f4cd6d8
z352a7a9848e70b9979c2751f85374bcd3b04041b5487a9b03d6ce18d0510e0a4a583a6b9bcd6e1
z5d1fa5f80fb21772aa0f0b1fb19f0504c4ff65c816394b81f669b1c9242daeefe85db0e1b1190a
zcb5da4777ff2e977a64bc589b7b5ccc26c4c0c3dbba092ee41a1c8c3f43a6b13a51709b1a34fdd
z9e3a1cfb6edb11efa338f2cf1af3e077cc80dfb8aff6b4ecc68a0297fa3597f005f615771720a5
z03825aea87d4a38a6fa06de5033bfa30db4b81593257ad4fb9eb041be2183ddc903a0ded788f7f
zd6a5ca342d0ebabd1cec0a7f2c3dc2bd938ad3088b8bc8989a48f0bc2805a3882768983e88a341
zc71f15976589161f6ded932f3731e492371dc9d5cbe3332b5a878c4ac6ea19fd9a60d3497e4836
zbf410d4985c5699bfe02cde409800e1e588f4a100372236469e12521fc5f0cb68ae31fb8ac824b
ze29c5768aaa5d903685cb0bdae6560929b745b6407c385b7bac05f568146b94135add1a5836361
z7a8c8e40d83dfe25a59fe3bcec9ddcd59cbb4f47b4f2f2e34c016072e3f5a6e40877ab7ec42498
z8df544af3aa803e8e0c41354e90e3a3761aeda8c7b0d4ded2e2868ef8bd1ae6724c9173b6429bf
z36ea5d9a5d9c1bea6073e08ec6bf032c03bbeec31f7e6453f783d35223a367db21225a05b4ba9f
zb2b163a699f2f73e4350a5893b560f67b98cbddad4d8fa19fd583b5bea3ee55cd74decf7d1085e
z173a22b726a22a492af0a23c35ca90b33f034cc23add9e63b1f6bc2b9efa6b323b792062c66458
zae8259d0f66b9bd1b9afb3feb49544eb0d59a0524b4a9928da69f16fba6154153d8d01520b32b1
zed27112783ff6a74dde39c8136d006e4040a59e57adfe1b4ba10b825105ceb55024246989522fb
z7ad6916bbea6d8edf5b030d59e77aa9c6d9ae37cc2ce0643b0e5ab9c5e3bba156a44003f4b4524
z48260a059a7aa5f0a34470e868fada5f91d431319f6dada623c8542dd253434fbf6a15a6cdaf28
z4e312d80f600d441b2afcaf2ecc2c73954058f2b9125a9bc110a06c8620b0b825009ca17ccaca4
zc227bb41dfdae6f98b004c6b9ffa45f68fedbde07557043c36cb14409d2e68aae8af42e8f3a6a8
z38795717259f208b6f846a399b86180ee97a056840b72b96b53b6c73cf965ed33a6d628df2e488
zcb2c21648d1c6daa6acdc791a53b6caadefac634d1aa773d46a6fd9f0ecdea5222925d30cb28f5
z176cff387fd0a23a3496dd02b0d2411ff6327cff0a5e70020d78bb39953dda5e194a82e4532562
ze22420df76def824431dc23c5c28ac1797044f97841d4c186ab2b55b552175b11eba19901d6735
z8a85c6b4215f5d4c755abfb9a11fafe6bdf3dda06b465d09d529f205708024b1ca11e7ffe6a466
zf3f32a891b768c0494f04bfdf9a12522e1f0acd8d2cebed5e62417fa2895fd67f711a804adcdab
zd81c7899478a85eea0f9bb6ca741ace213d17ff635d026b04ede4a35b1dd1fcad988a6ad22ef61
z9052d9f6fc38f219fcb31fa0de7dc54b7765f11044a70ac1a56cf992fcb7179d593654db195d35
zc0350c71898b2c962cf0738ec0de301f590d151e39c7303afc01a319eca9945cacbd7a1ab13501
za06d248b95460430100383d1d6061aff7ce3def6c7ea8b806c979da177439b5da6a100fd585c84
z363df60abde61e5023253b75568ebe1ea3ad3327bbb720b2b019873744acf65c5d2638395d4b33
z35a96ad83abe5dd324a417a36f07361929bab8c719bdbd40ea1333a7723b0c37265677d2c586cf
z240504060f5e2a6a88a3d3e4b302c953fc69f9b2d4f21d610acdfda322404c7e3d656997a9de42
z16ecda4d9f6d4756e7812edbb97e7bdc86a5c7ea3de05dfa3538d1d0fd4655e8579b79fa2cc88e
z3001814421daabdc89a2f03dbbcae412f99ea19bc7e79e09bed450187ad93685f4382989562c7f
z4f90401d5d1862018d8c174891429c8b039a0d14b4f77d5ede553c035360d075bc2eec3d6dd507
za221dda0b13eee4139825ad442db810044a4750d6bfc8e1021dac78c8a54f9d95e3c510dafdf3c
z949c806ab76f46a833ed8c54562d70d539d28dddae3201c7486143da88efe337bd4c17a4b3b15d
zc83a2822409db89ead09914dc0434c2cc8334a324d096786d3dd96cd3105bd0635bcab36e69930
ze5e51ec3cda6165d31c5cfedb46007f7241cccf0d5aa86864911e6b77e352ec607514493f3d70c
zf04e39e21aa26108c3eaef991eebc904f17b44a06c11df6bec1b68c10f01221d030aa80eb6c599
ze497994b8cb5e7672f3cb0372efa9382cabe3c60250d24bbef03e15ca2030b711933000ee18f6a
z89b60ad4555ef644105dae96ddb862993ac28062c4e1e0883f7d7823628277667ac73a3c553541
ze799ee64820dfbb47f8848d528568172ed3807727f0d4519333aa81329808edd301e02e4f753a8
zc6e429e055e8531649b3654094995ed91bcb26ee9b43c10aaa7bbf43db378cff086423e7ed5c86
z8e81458774ea5783ca828cd7d7b7a92a13311b114f33063ddc3add0e4396ba11995e19f088197b
z1ab51d02663ec7f2765bbb09b71927f32f729850c7a2919afa7071c345937578784a88a87d857c
z005c96b0491b0ef8726a10fe538b6357f966e9c6f4d9fb94b44728bc3b0836a6d7d8b705dce9b9
zd31f48f5f649a99ae9a8000d4d4f8c342906d38fc201b57f44ce95a5d95ace57306e96d8773753
z7bf929751e73930d1dfdbf5fbb490a967571d5683caa2479684ff859480dfefe840218a878919e
zf443bc9a3c41dcc0e7bf1fc83747681eb7add2d784c10acbbc9d211f7f89c4449904f68e4fb890
z28b22b7484dbd04a7dc662ba1902ddd5fbca05216f8eda70eb818f2d6de99013041f1bd0b324dc
ze0f4a7a919eb8a6fac104aec3c61606883ebdb424dddec6ba36a363525315ca2b8236deb831e2d
z27d8bc7df7a981d233b5855ff01f348f00c854a6e68b46dc5cf825cfec4606fa0acebc30c0bf26
z17e6aff516996f17f0bcc1264906b0cb0848dcbc90170e170a44c861030fac3549702e1b1a620c
zd6d028bab5bd596a10990ceb0f1fdcdfbe40cd2a808ca74aced50d916e2d8e2db58916afec934f
z1636af3844c7ab605754064c298275bfad71084c6375832573429320bc146914437fdf816c47f6
z5bfa895c7ffb1bcbe97a84dd0ccd340c35b858d7b3f494b7e197a94aa95c95ae064542deae46af
z7d2dec40cdfa0784ea7a758605b04e73068ed07c221ed520d0b633c6f3b51f446effbb40a89c3a
z3f80465f11d858fa5b7acbfcf036ab533e83d540cb2392fc9949469bb461d5de88b80c3303d29c
zece027a53d15fc55c5a1e650b42846ddf96222b18a7a739979c3242588239b044ee34d275fc0ba
za1dfc011fc774ae3c980de09569c42fc87074e56513884c975a6f659c705dd9508c1fab2f8bab6
z34952254411f4c3df793a68eb43e052c074655c61437c20543ed5afb4f2779dac312e4ca509bfe
zc93e929584b79206f1c7bf4b4320713a2c5c7876daf175ac0380259ca850ec9f46acaa342995ed
zc91199bdee8b3445b3dae1e3f1227689470e2074d9bd6837afafe48644641133faa89b2b6c02a1
z7dcbcc6757595cac88a0a8dc81710fa0c04c24db59e3d4f28043e7308eebb95cc0704d31805bb7
zb49f140d7c672494b8e6ad1938ae125070f212c3c129c8a3b91ea580d552d3caad91f6a984521c
z07c8cbc06d8790cf0ddaddbaa018cc100007dfd70056091ea8f25e92ea48ff8c3e3f24c120c0b9
z3cfc6b11a26da8889b24808b50675d6ef4a5965c7fd08208544d3d1c5d8cf5b3a0301473436fe3
zf9837103b23d68b959c5bab42f58e7260b323d09ac7dfba161ffb681a90b928d8427840a28f59d
z7bbd56ab5f369c9f32e4f87e8891cfed04a65791fa7bbf1ae91b4f5dd146107b46dcb39c2d4798
zf563aaf0aff1f9cff7e55209f2a07d672d8522624bd30c77e5217df9153f7ef885892796ddc3a2
z0e70962939f3d9d65607f08197c297d5f03b224a2d69659076ee506a39c529eb792e4bf8df80b2
z4481cd87880d166aa79d9f85a27a2cb7ad9d2f4fa98d07400b1f033d65c6573f4e9219fc6bb3c9
zf92f8ee698f20811f6e0ca0e2ad9d126705f85b420c012559309f13fb1ca911dfb44f47caaa52c
z968b7118d8ad9b2497f041606cf1e8e11ec3f57060f869ba219a921d996f1165862cf536187288
z20f51192f595e3285de5f96a549d2c5c344a6e7226360d9395289299fe87580c641cc8ebd47575
z03f9c70e2a450970d693720e5fd82917b767c567ac30277c8d8d74af245295cd0d18b33b4908c4
zd1a0d7fa4b47de529844c801063ec7da36f0cb4bad6237d366d61ca398f3d44c4e7a014e3318c3
z6fc201de16e24ecadbb60d75e35d9073c192480e9bd4eac8439ac3fe668c560bc0879f373588e7
z03faf3847d4a93a32fb5c1b588f57b3d50c5bbf5315697922af7e1cf312de95022828f67cc71b8
zc9d81461bd0f799e03fe4e2e8b538489e2b66c0f299d414c3ad88f0fb58dbc30f7957beb41c44a
z3afbb952607966f24c18f65bdb8303dd7a3d7994ceeb71b77774d432f27955e7137a6642884ee0
z95ecbda9e1ea6fdc1e22fbf26a26135aea00930452921a1a9166891605e7520492f4457aa3b481
z90104ed21af6b9177b7871b9024ac863c0b598338207e7fb48dad7abff339e1d6fe321b1f72601
zf48bb4f00fb877ca171a3c4eccf0d05f2bb4f8808d50b4be1e18eca07719fc8fffdf778bc18f89
z5e9a7618efdb5008652a3d680226a013154997cb5f29046d523fb9f61119069df98c9c98079ee5
z42f40ef88a77455d05e6607d2c463cd3ddbd2837ed1a9f59d72d06b5295d6597a7c4d75ccb9845
zb51794ae7012a3e51dbe12a9b63971c137f722f314ebc84102e00b1e35936615c2dc81952ee69f
zb1456f8dbde2da7f5842a02bfde06bae056d2fcc213d941f5055c0b516d396ab5e287e0cf9c2f7
z5c2fa2be32362b284bd66cae8f5a9b4fea637a5840e2b48f69cd6bf61f839ca6dc63483d5b6f72
z4f4c5b5ee01d6d95c7f4f2d81ecf3d82854d5f41cc68620d608cdd5155a37734e92b802a7c9666
z8b6f6b50b514221f2018b94d5a7f7d0ad4254934d3adb57acc386128ca2ae19fcb03d9390ad0af
z760d5d883ca9863a38dc2fd612d9d115784e4658b0ef28c9c01652fd44aa81b1839e009c0feaf7
z72ee84046fa1d15417aa923912f75f21ebe0601d5af0bf2839d71099a805cb728d0a8a93cd804c
zac62cef7095f5f08a7d8e27412ebf3f05aaedc791d130c150bfc938a068457d68afac4f2790525
za9ba9e81684213f88af1d1a44598115dcf687812ed01a3d52fd7837b32c8bd4a523106ab66cacf
z7b02ebee51c1f827dcf9217bc48c5c41cc1c1975dd5c97aea16ab14034ed13582364c3fabe3dbc
z2fd83f0ef4fae36aca18e540bf11e363b643b262527b69b3198a4da532922ae46ea7df82c661cd
z21d9c7f0e2a489c24cc8bd4172a7a12f60decd5204a2764032d40709de5a2b1779d0ea4933a785
z54316dc8ee692dfca20fafc921de1e801443c64b72dc388c0a344fa5132c365f5042ff912440ab
zb49cb9d8591182ca5ae113618b48436b04509cc8abf4511aa526a2e5216c085fc586fb75dd51a8
z19095207f17a2f0c381fba2c186bd7d5cc1a4ce6df528c4223b72cda3f04f55abfc79504bce9be
zb6828f7ab75b080dbfa44a0cdf7a06cfbd9a2af013550808e868e49dedd989a4734ece1dbafea8
z8d78d6776bd5f59f344238fe956dda214fc8c3b866126ce3fa7f9fa334f163ed5b78bbf59d428d
zf63ac345072801fa092d44f039fe54dad89082367867c7a4cff0c1f4de02660691579f000fb88c
z24891d38e58272716735ceb068a8376d7bfdb766e1a846cfe2709e950ad5f0889111a617b75a8c
zb9ec1a3c72d507942d42aaa1e4f6ff13cb5633ac9474e804ec9249d514168b090906508c391b4b
zcecb1c25c8099c58d45444587f3cabd2a182c9015cca511a535ba6c92142033af02c72a452fbed
zccde248184e2fab3b42ed687f249c1eae2efbaf56be55f74613fd41681821b31e38d02df0249c6
z18b4d9fcfad7e54322dbc035a797146cd3dc60e0a2ad14e88be4a26f8b6bfd66c549eeb9c4c78e
za3d142a9fcb98cf7eb0ee253edf0f46873ea33f570ea18eb67208054f7e230d68fde1ad1bca1ca
z3bbd164201f92f70ecc1a3b5332091ad7400e0d08b7d6d1248748b97df7febb186e48768e4d5a3
z35cfea3f02ccc62e84f938bae164b6ee2db0079d1a224e7243c1c2561174aef24ee373301d9e50
zfc48ffd97f36322f979b8c044503d044257153707394a826032574177f8dd56f9ac06b3e1567fd
zde1453d850324aeaefd40c3dd900b848c87e3f00af58b5f9b99369ae3d3fbaa62a31e631b4fa69
z5e738171b35962c49c06393f27bbac4d21cb2e9e967bcc0c796b122691a915acf5e9934c8e6a4c
za0f55608775c3b2a4bfcb1a24b3621f8c4f9465945e345ee3ded8c2b7b48f56dce1499dc44dc94
za1dad4d0888c74237be0e8b969473c61cfb43fb465ab26e4357099670b4bad2654a86aedc47722
z7e209ed958dda6d39b5f89ffecda991dc429066c197744aac25bd473a5645c13daa8726b8424ca
zab10d1f7bed1b5ada17b483b0243c1e5e5b21b112b10d78cf84aa28c265d426f4f6ebac32d913c
z33668579db03e16832dd80e7d2ded1d58f98cbe5a807743bd900889f8959640513447ff9588b4d
zab4cddb9ae67577b96e992d1a62241e6d3466021c3ac0fd8d9089a91309dd5713edd0822c8c029
z7103d587a9b3716d62252ce1e4051fe5217d4d6da9ade0cbb32941aab7332a33fd90819a7120e3
z20651e68d6fa3f54dfccd3c2be23aa8a8afacb53aab71e82a907301a203c523b06d27a9cbf1d01
z0a393b43963b11d4ebdc5e97a4abcdb33c975d5c87b4c5741646367944515c0f1b215068bedd2e
z8d489cbbfa0b864e1709d5b47a0abf4f52e23c88e7dd2cedec82d8ebfafb1e30752a43bd9beda7
zb0c236c80e2b4b8e1678c3874af799457a776c91458e8925591c85fb6785e4efa74f5412856531
z39082a7bb89d8ee1dfb3c5d4053d36729986b42d30e27b6369145f8c8e19bc8be2febe2df5cb57
z7f9cd46e161574c6564f82ac79ae3caab26343d39630a047bff4b69225b33ab80b0cf3013a7ac7
z68168ede03b7116297567a3e97a84a84dbd9b7b30e69d34e7d3b185a62a20060be6d233b44d676
zf2e32266622ad486ffcdfb169b11a2f54757e5990c4b11703675f44f7de495294a3b76b615705d
z4b1287e555764376c718ed24bbede07a84875cd9443dc7db4a14df5d8cba799cbd16db056a2d86
z9ffd376c178163e72138c0fe71a25bf13dd1bbe87b438d259413cfd1e08c501f6ec3533ca79ca8
z8ca68084d99ac28f321f0f43cc2f1ea8dc146fc11f9a50455c197d5ac5a8780299e9ff85cef7ef
z7eb2521d1a40cfc937319f353240267471ac03e6d6ae3409abba9162f1597a6c806062d85ef12d
z60a4768be3399198cef44d05c3096d3bd79031a686c592214c9bbd52645ed58fa020f227bb63c3
z9dde8d5d5bf5637de7afbd093f5d979aa02985a18e4e8b77612872b18f060d468f524c970150bb
z8bbb32a851a102b2cbfb9e7ffbadc7d240536e6e7d755ec6cd6c16db7c6fa1469e0c38a8381cf5
zb3b502b20edc789341a3c514d326d87c216d91f5dab76159a1f321b611ebec3cf3b2be8301df1a
z321f71209bf8c32c272ac09e2fb400768e9591afaff62197e8fc2ea41bceb7742a13d2d45ca4a4
z8b75a849ecda1cf9d3cce1ed96f16ed078c03e3b20195bac1b280aaa68678465633a32b86767db
z3d6ccc1599e5b44954a418d370073b3bc1a8c657ac1c1fe71eea77eeae5ffca3a06749eaec1e98
z88e9174d283af807abcb3c695066d9ac4a3289891575d6d15ebd1fe2e2e0e1b7e4fb258cb7f1d4
z4cda72612c413b0909870a989098df78226942257f632eb78d1ca7aac5f53f7f73225952103d9b
z1e1a4c295e71d3c43fb3b9ffffe217814554d853b1915e3c1977b2f2417299adcbdea838bccfcb
z203e0f4b816811832cc6b1e1818f98881d6c603762b173bf20ce688b80b4ebabc8015a4e1a52df
z6d3952052845dc1dd7ef1c9d6016ac9a7663a18ce6dde7bee37e8cbc979aadf5b612c4de5fcb6f
z2bcfa973986e1a510326b2e5d5888e7a3695af3289fe58356bfec6884c38a85f27086a6d9591b0
z3dcf349c62ea9959a4837f50d8f392e7afe598098aab3adf1e53f001b7da50de2b76f4553a7f99
ze5532dd708a536758da1182888ca2d1dce2a982906444b062f6f2677aab2dec1cbb48a38f189da
z85a1da94f545cd7936bb21604e048f075186b1cdb4f26fc4ef457d1f0ab488e168dcc5f7913852
ze486ff9234ed0b8413b5ea10fbc199553ca754bb1ece075decc4eb881387bc70d0887dd690c640
zb7d3a533a473bdfd8cebf9ffc43c418a49e3e40dee0fbe5b09708f12f62ba63482564dc20c5de2
zb4516693e54db3bc603bf561442de834567952431f40801c28ea72e1a2944f14c96d0ee15bfa19
zdd70961ee9a7a600f9c9ca2fe4c0c567c38a222204774e5bef1f838bbe73cb5cd1c87acf200b09
zbcb9029902814ff1a14856ee8254edb3f8738bbd66f2faf2f27e984106428cafb53d6496d7d246
z285a241553ea2e64d4726ae6992e57cc9f39fc5e0fe6859bf814525247dea8eed1070b18c6c29d
zc2d79c263be2c7a481dba94e5370a46c5fdb1de540b35c4e6a8a693efd7c79fb83f00a6fdc398b
zbd3ba0996ffbed4ad647dacb32e3277584704c29d141a66e79aa22bd8fd2cb0e0386283e709dd4
ze817e9d7dde1811176380be89c69445d5305a880ccd1a85660f8bebf095d9ad0daaae59511e79b
z67b74a75be9b4a001237211e348915e7c9d0a759bdafefab59f3a4a80ad7d9f675c47298864c85
zd26f64a28f16473b2a7709bbe5b25923ca68d6b93a7416924550475d5258f6ee2a639269fb48c4
z963a6c1d33cd01c181e433ed60404c7bcfc2ea85954dd1abeb01473aed5cb8f152e255decbca37
z9cbb8d117b56eb8b3e9f5a3ff383522a96e9d68400c106388c2803fd7d12ec1b9ae62d6cc1b993
z660d1a13bce9dd2afde38fcad3a07675a22eb1122aa1e6441a20a37a49d1dd6a051d823c22b6d7
z4aedd09aff3e7e6f664d351379f04a241b8797a32d61f562de4c8f85324c58d1e0d17506bf474d
z909955a2932b8d402b6cf0d926e3e1c3e5c8743109d5b9c9c5150f6cc634529bf42db0ae80d6d2
zad40487d4474a9dd0af01136843ed81d06e37b11282d4ca9132ddb970f3b3385d7a472317b17b9
zbf3096492e84b13f0ae3391b7f84d4a2840245f0bc5c29a1551412d51800b934a9a1ada0e7c559
z8110920ba783969ba8c465ef1249cefabd0abd8f6f4bbe7a5a02b4ed7d16db87ce65ffe603d078
z42ef9727fe7e0e1ee3cff90f42b3031c8c5472fb0235db06b2fb107cb93d252e342768866cacc9
zf71038bfd99280d907da108c49e9da74c37132776185df484777efa5313340dedfd708e3a92022
zd1abf69619f7873620753d8f06718d6ae218bf533f8acfb2910d4f7de2c47591d2dc9248f73d6f
z2a65fb8c43ae74c405787e1855597c844b987baf09482ef7a2ea1a0b35c36287dab3f5ab4158b5
z7cbf5d5dce4c7065fa5383701f732a7e5d683f68e86a595795bd7cd4e0caaf8cefd40782281121
z9a8128b15eed312b1d56016ad85cd25c1b22a1488898d503280d073d79b63e22b892b1e585c9e8
z0064b6f03400526d0fdb348f1d65615ef35565d51010b4011fe650a0745e3d288aba3216c7212f
z070b500eb4df9eb91c563acc55a16b8bec0267caa082dd9cf34f7e09b2dde8fe9d1f6c900145bd
zf843ee3e5e80ba39a195ba86e821a736808b9392d8505699d684fba0da01e5a9bcd2461b64a20c
zcc08c8935e951a0204928cd7af7b8029b917671d6e88163da9d86be8af699bcc7ffd98d7633959
z02877182b466a55de23a47eb80abbd8d9b6e43f81949aefc6c4b575e55f27ce9975d1febdf91f4
z939345858bece3b34cb25bb0e2a3ea6b112f436db18a9a176eb9103ef8fe3482e4d79926fb7a63
z6e4aa2c86ec728bab31382450f2a78f849a3540c7455093103901e87dffb79a74badbcbb35b7fa
z223a637bfb35a73a1dd5bff84f5c4ad05c25e2e0b2d888d53c7e48d372afcaa8fe2130238f0ea7
z0358c09079238c4650d7d77bb465999d5707924557d427c9fa80106748494f40d5b387327bf545
zfca31d63018a0bf6fb85d8b0b95bb64f10c0b38617d6b9cd8c035e3fa1fcdabab7f12281fecc6e
z404d1a3414815baf6ae77688c64c77c72d0ce3746bb6565ae2ecb506efdee0fd60fdd90282002f
z2c750f93331c12e0b6eb48281a94749996769d008045335dacd0cfdae71880ce4ac6f0d260d05b
zfe6a13e445a71591b8f0b212bff1d86750cb8eb94d121e670d3b5245e2c8883ab9c6a20ab18df6
z1d1915f445a037acce4ee3b7c5febfb048bc5fe5a55b7fbc8a4cad5d2caff5003c7c934c8fc158
z6c9049aa80a00e11a9fbb48cd518b33ca31092dbc0f46f21e7a0a318fafc7ef1891d205ea9bd27
zca5f85e1dd93cc97fa9c3a16f2f7e0deb9d13a63003e647cf83e33d74e88ea3b2f3c6b0d1b067b
za78127b9aca3b42acae70bad08d8c63d2401c67b2e35b18a453c3881f3baef81757c1798a0ce1b
zfb754790b8c18a9fa5dad94c4e5afabad08edb5043bdc4afa8e98b7c46d05d539b27182c266ba8
z83eeef68e2013936eb8b71af2fcc167464aacb51b7095f3dd402edfcc2f98cc2f3680c4a78a056
z1890a065ba9ddb4fa0f8c6aae7b4c42795aa1c084de173b5770d9e43e49cb78b51e10bf3c37fa1
z9b67e790dcceaf1141d9be488fd8c217dddf774e806c232507b99a907a54a1f7d2775e3977a3a2
z03ef24388b249b287bec3ae24418d5dc67e327efccd0b619bad75dd0f948b5c56140e65b8644d0
zde0b05e44420a29fb5e71ba450610f106197e21eee461f0511a54e0f990763113017e6f4c9847a
za6746d4a8ec9f7144add573ce2c10b94c3334c62e89a9cb7eac638ad659d333016ef05e217cc11
z953a57d24a5bf901bd9a4ebbd764a1e08d0ac8d6d86161ef9aecf7e0d267771aa8b4f5d24152b5
zaddcda40f4899db89e8ad1336f81304ce56841ffe0ba5347c7187c2f0e7cefd5fe1e51daa35025
zc4652ae6e3ecc08a2ab5601bff25f87d98f9dcaf86294cf4413ed99eab734df373694d9cff31f7
z838f495dd78871f28749e8e3b3a68fb559f1e57c010d40ba0634258b544702c9f0678e4690097b
z085be42f288c0883e9557809aaf5f4ae363e8cc6c19081a2af05eb85d6873ccbe2dda45155fef3
z641fd631cbe1f92b274e7e8da75c463d443dc9a30ec6e0ba84fbd6a49b4122ef110ac5435fd336
z10c5d8ac7a18351456f4d0f14ac9d3a0ba615526909cce286b5e0e4302cfc5fe991b191b8e8fb1
z097ab687c2fc4d9a758c9c0569c4d975d0c968a7bf3669a79fc02936d2462675f99294c67d95dc
z22b5ab3dc7eb061aa98aa26923b7cfcfcf9b031fdd3f68dd6bb08a0fe580266a5f6f9b147d4112
z99e484584c66f2b5e70007cc320b950957b7f3aa50fea4c1b4cefaaa730c7174b13c08ec36f7d9
zb700470fba31aab4907657cb296fec44a5e7330643c4a9272f6790e3f7427901ec94b2af6e1918
ze549180c126e38b3e832fa1a24047b518dcd4e725baf245c956fe2fe902d944395941f82a5fd92
zf0e00931e7ea2055ef85db410b77576748c277650c3cc91ce6dffd3ce6fa753d87130c00df13bd
z4759a25cd7bba98ba15a0a385498fd89dd77538ccae658069ff1186b4848e74b750c4cd7da4dec
z3caf82e0fc70afcdd5ee397a4e4f47ae8259b2da38570426b54d0ea70bfa9e2825add45175da58
z8b222a0f0a64ccf30eb6f90197c27d99be8d3988a9b8025c998e619d6b17f71a4f72e5733eb218
z9ade1ec301efe48cc05bd99a98c992dcad80836135dbb6b9c17bf552f32b703df6ae5dd2f4895a
zd012ea0f9a132b214cc0961fe458e0c5ac87d92f7f07c7c42190953888c2bdd5bb13461e450851
z8fb74aae0bf5495ae703f9bcd73dad8d3813054f4044d39b5dd11b0e89a58b35f116ef238482d8
ze07dc1bf70999476603afd3173426f6d87ef9c3949e3e641b27c9724e4f71cea73dec5cd77f85f
ze89b0bb405a1ec5204374d3247c10cf6676104f30abbe48df6768fd853f02efd965b8b055c2908
zed77cb6e6b9f69faac0d71e9f0e730a4a4feb76b17e506951cf845bec002c19015b499a135522b
z1c81dcd7fb60d0de8480e9a913f2b3a6fda331a6b7da2dec0561b2e71be0c71a44f59188939334
z2781cb931fa167629def7a3f8f44de99b9dfd153bcb670a412a2273e3e62fb17345aa687398c18
z12203cef9b58bb5b1c2c00e5a1985a1be9102ecf045382edee4a7dbf5ad88f5512b185ac835f46
z39b0f0f6cb999d1ad42f56fb1cc599c0f31e7f570d4d355447a25adf847e169c3cec83d2fff795
z00c707247e812464fd1bbcde965ee86ca18ad6d37b4abd63cc2dc3bb5167f8e80bfbbf1cc93efc
zf54adb4fd2c10a2f28cf7bace88c77db1a48a562e7d3f6c309caf38cd2d3d0a4f0536bdeaaa871
z5805324996f25b72f471099163a327f171313bf731e2dc121d32417f90d0e54e5472dca64eccee
z31bb54e66e40eaf64fe1f382abcf71ffc9dfd4791a898a46ba9c113f22158779c237e361ec2e29
zc0e97fce8c6fec309716f5dd14cb8f3e57e52a2645824697c41b5c6f3d76b71ce2ce8ff0c7e2bd
z95063d3ca965da317f365761ecece11a62c78a3d12f1eeeb8172a799cec9948cafa71265f9eb12
zf05dc5bfd26e4b2cf816417c6b8b974d0087760344ce6775a46ede63c4c2aeee71a9f364d214a5
z750fbf327b4e21b4cb5f1247cbac50eb64e13c66fdc10394b38c9f12b9262a365455589e56312d
zc3e8b31637a3f2bd215ffaf6adf09f2a1e84f09445ddf154bfa4a6809f62cf1f4e19d924af2912
z120471038592e97489b6553391cce1201c4d008f716e7cd4e66fc86adf4d07c8c131a75d9a0a90
z3aba9d5cdaa51f78ac78ce0d89a70fba421259e0551b6abbd247d0b05329991a23d567fc68d5a9
zef557223ace9b8ee8a6a4cb0f7efc49e2a5c967b81acf712bde93c23769640e53d6bf4421418ce
z22e8a0c57e4d08a3ceff87ed06a0915e4d2cea623a03486b6799463595069d39cf00b9f6736f25
z86cf2f5ae459f76084fd73ae99e0950b1ae13274098cc54756b44d0d7cbe7b55d00550fbb6bc12
z40550bf78f501543ce11fce78f8ce60023a7967f51481f15d618bb7cb861eb05a718d8a6d1c786
z941cb41370081f75d7ddeeff7756fcfff4b2fbd7a708942c5f530458308a6356fb472654285b4a
z34c4243e331c8cda922ba91e6904867b31947c7c03cf4e1071fe4163da07795a7d4a2ab27152e0
zf633cf710aa2f39ac51e836f3d8791e26ac4503114178ab2cdf71e9c66022cee80c27b713116e5
za3a6b0ae5b1be8384f16f8e1d9c3fa836c1729af1769b6352dc1de3981285d3f7be6383225f8b8
z1f9ad075c287d9f5b6d54eaa11856339f80470c6eb5917e4682f5cfcdc3c1880dda2b710febde0
z1a419addecee148a993096deab4f2124acd722ecc3904f51bfc86e8614277417b46020fb357b92
z384cf4909a6e7fa9c0163e250079e4ef24116ffff8234863231be16f6c705c370e9456c90df7d9
z3692710f1202f75e5ca0e3df53139e5d159d0a3eadc014727eef36daadb4a02314a802f8dcb8fc
zd5c645fcf4fd3dc66b588c26a08a262a5cd3fdac4c5a3fa115d777a1103ec948a24eb4f8d1fb99
z09aff67be44b92686721d53622209bde0d16759c742825cf1369f79c39f3c00477bc8f21840b32
z46f61ba38f60ccd9de6fc9a19d2b74fdf593cdc49cb203e5d60e62596a51b22a01df91e6de1759
z19cc29370629c5502a09fc3ebae569860ad1a04a8ed126c8ae72d14a6063de8a2497efdb3d5373
z234152e66da4c2ec9ad1c81bacef198928d369bc2ea5469054fc0c8348374b93654c14e66c4b81
z9c950c2b1188159a5d9be27fccf43026b774e16fa1b124796ec4ba797e8affa2d805428702cb29
z6af8b9d0f80411501f4ca67ad9833acba6e9e37b3d65ba836e94f89ee20dce32adc9837bdd6250
zbb0a3ec48442cd3d37fff3b1fc942b6ad5bc97cacc309a9dd8089020f1ee80bcc24a1bdc1a54d9
z9ff91026d5335776ec255bb3e01fc85487fa508c4f98e784ebc3ef8b228a59fd6ebb2408382bae
zd3b008437b847abc498acbaeff538d93ee15fbb3a1555205858df47e094a043827a43f90ce570c
zd546e9804ccb903fe10792ead7772000ad209f716efddc61c43665d2b0c62f1004d5ceb33e3924
zbbda8a8649e94447d335a8c9abbbe168e98e63baf48b692c4f0f88615e5ff735678052bbd11784
z835d6ea8f121d3d495e49136a33f93014a86236d0d45a3e069a087f200ef202b103a11a416adcc
zaf79b2945c610ee4bcf28b0712c0bd769a6ea971ce7d0138c6d2eef183ad95551855e7032fd3ab
zc5a9faa9128bf5de4f262b0edde9f692ef5dade1f9af04aab39e4b843119aaace945a74de3cbd3
zb17cc6cc4a75ef75458c12e975a885cced1450c770bba6ef399176c21f98773c11f4609ab34ac2
z140be5e57b6553b7a2e7d5bdf07cd1da0ef9ead6a2255cb5faa49b6518b7ee55b8970774896932
z0baeb3d88f0313ed5d0ac8346d41514a3e1d27a4f44ead4b48f8b8b8bae956017f0e2cb25c822a
z6abe3f446a1055b710e2e8524b422ce994ed213e783f523bcd1597239586830508e0c104e8404a
z80bf29cacc1c0c8ea624b42066b453eeb61f747ee7fff93139bb566d27e858578842dbd988ef62
ze77273540dcfa9b66c10fa8670ebfd1241d64973cbb273f5244d8c7e37cb71705af94713b69ae1
zc6989d700931e4cb83e790a55a3be1c590f65869a2d70b7ea749faa3d9ad3feadf01a385bfcb86
z1aae083d5502c45dcf56828c4f46842d0c57335025631ee6c731a46fdbd8fd5722d07ce89a509d
z29ea2ad7e03fd221dd7738423764ed719ab64456ec969807de33b9b781502ed28c58f4516877f2
z5e1464e7f61d836a371bc7df0addc21e80e87dcfab0e9a8b6638a146dee0d0029f12cc983c27cc
z3adc238550fbff7a2618e0c20357de790c4eadc134d61808637531c473e63e28bad6cfd2b637fd
zc25644dfab0218fa9b3a8783088444e87153d272d2bed1b9eb0531b22a2ceae16fef1d86246199
za21f80e0ba0798459f0739cb751da7dd49fc74951d64c6c94fe2ad279d30558da7fa900ae11cdb
zb3eced700f2bf790f8da2fc8e6d9d81ed69efaf6a8a76d934214a7f65f161930e0496de021c9de
z916f12e5668d23668a4749914bc5dd233435cf19ba965b9a4e8cc994531ae431426a717f7d7e75
z523619b07c3bff7be20639e6db518da609c9b4bc85904276b57b62acbbf8e9b62f108f22a9d465
z75633c4327094a50f7d8942c12c3dfca9625e672af0dbc5b87eb7fa575c40c8725eba5cdd71ec7
zd6dc82df5284df5a7a20faa9493321c6a9dcbde50dca5ab1ea472a918a8c4909670b0bdb5a02a2
ze3b1e0d12d4eb3e9aa58d36ab5eecc6a923fbc9c91761aa49b985c80b3683d2bf834c610d89403
zbf05350d2eebdddce14827289d49cf4b918162dc8cc7e31afdb746b2cacb86b5de1597adb1404e
z6467bf092b0f2c3013dea6cdda49a2cd3c11a51983837f450100962f769d1c193c612a418abc12
z05e22a3b4e2ca79000669bd179a5ce3528fed2c2a58610bfe71d4a0af331a310ad3b57f1636c6b
z61bf4fd7a609fd10c1b6401b043ac624c5b87850f1050624fb879fc2a33a7fa743143958e3d7c6
z8843e4e3ac6a2a1331340bf255f97a3e564bd57613674272b17e8c70263c223a3f25e306aa054c
zdd33db180cd5c8acc7e7702bc21ac7d93059eabd240cf6bead245d186caa2a705c6d01aea05c29
z2fd96c02d89962f1a48e85dcc806891952c400984fd765359fd1fe2b41e3160b4ac4ada8d9e0e0
z7f9c1134fbaca285d33adbd261677e385b6f3be349d3b1ad320b2299faf1a5c5cefd903bccd6c7
za8db173cd9f439340f140548b379fdaae0fb294fb9cdcc10ae407ab4ee11f5cf798f61ab48851e
z1ea576a18f9ce95c4fb7b2d31aefa8c51a8b05f11f02382911b14c10f2df2a07121e78683bcadf
z007e7faabd832a8dd37c6504a2d88971ec3128146be1ba921af5b378d39042a29398abcf8e5153
z750f9990b1e021adfb807c2d833c7adf6054bac7643338bb30a7c6b71618b03bef33c6affe1759
zd7a3c770fa899968258696e61a59b0589e9751e452935c06ade5827627850c2aeb92a93a7d0b48
z0e2e60481bc3958cfbfe1e123e5c8b44583ee695c2d7aaba1d8736afaf7b8688bd1cd4d8e8d5e7
z60a4a321d32a6ef3a7fc938b2b07b370faa4d7d211a871d7e8ff684af8e87ca69c7dfcfa3a263b
z5ffa4de51f5bd5d6e631ed1320da15306a90864086fa25284465b4b8c0ba8e758c0549a26b0668
za0896d6acc40033d93ae894b3afc42883d57cc7b01c8e63b9a2609fe3785f5e8e8e0debcfa2330
z2210f22326ca4e5bf7f269828531d92f61ed513bb5c10e4310d51785f141047ebfb8f82ed15a69
z160995ca7c35b2e06ded183a6411f767cc80a862ab08c7b652b709b5c411278f1604951a9831b2
z969e1e9b3736f098845d4e20cd2ad02e18fd2331bec47cd8eaa4cfcf959137456048c93bcf5b6e
zb2108e03b5ad660487c18202b2d3e34fae8908c48323cf06e3f324e47ccb0df7e2d5862b0dd55e
zba5279dadbea4cc8f5048eaa8108f176990d0d39b3b309ac19abcfd5e77a1302e1d01f13301b1b
zf55e78cad65ac8abe66aeae502ccf014567c7f75f800949117d46733dce2e457dbeff109e81122
z93059273b2511050e9133b93fc0c90535598fd81d00eb4218e601220369030ba200027f164d9b4
z0d126b7b0aceb290210025a89de60c4a66a91ed25650671502e46379140dce7591048b6c40bd20
zf52c6d274af8ada330bc57fabae936e52d8020546123e204d807331ec574f889e2f902ea749ec2
z828017a9dfd2ab9979db35fe970eb32fb7132bf0c69900358cb109db627a4d19278de175d73760
z9b731db58a5b4be253656468b99f26cf441546a2a5bffff3b5626783ab2f582cfeb66add73a9d4
ze3fa11f39f7b2ffb77d007cf28f378120436be8a2e39af7c9787452b2599a80ea23bb2e0f24a75
z2512737aa178257fdefcbb483cc332c204216b0fdebf47d0c8ca9118d7a106254287751728e919
z2ac5fff333848183e013fd8da50af2ca595a22b5e3025f46c10bc42ab569cfea763e9a7ccf6bd0
zc83a4dc6bcaa477a55f4d5ff37e6d86149042822e2ad421c5e142d6f04e39e979cfb9466bfd5d5
z40abf787e16ac028eb0216484f2526c72ef4716fe2a9a3e73f836a9ed82a747f429c371e293aae
z978323a9796a86a13e5b69541bf5971ab80d97479877b39ad5d138d06b1eed6fe99875aff78eca
z9fe8e893a3b8362d6f30461658bdc8f98b8a4f86da08fc040e573c326ab4adb54f537e0964350d
z31e2e35847ede289f4584d9106d04221e0d1a3c190f1e15306741cd97bdef209bed37f7bdcc575
z03f5480859f632c07d5edf6429340bc761466d613f9daaff548e2fbf11b6dd4e0fae4b24ebef00
zb02778a3a039d011eb5f86228e6a29904317caecf5e09e53ee6ad4dd0514fb9e8a96292334570c
ze6127f9d7f65212199bedf97c230f3ed4cca88d83fc04e4ef29675384a161b58139bc490c0e9c9
z7790c5c9467598498d2fec35030d3cd0df265be6f0587f08e97145adef0fab4a563a3e314174ad
zbe7e712382abbb79a40d2a38b65971dc6379dfbbddf31a11c01d7a05fb9f9ac65d69fc9e6d8903
z0318122fde5cf12e94697a29cc610465da1e62b99358ea6bd5faad52a40ea58a81008eb5a9cc2f
z4850e5a2255aea1036bb085e1be72baeddc45e7b5a57e6693521a3f20597219addcc1fe6d8c985
z0441df1cf0e4213444f7f60d17bb85168a05982b0b81b0bcc1b49a55bd6923b32fa5dc154ff342
zaf2f7c947cd391fa137589c9cb89f247ecfab5b9a0071a663ee11f6a412a5854eeb450e563dac3
z7a9302dad3bdb87dbefa642d1aa93e37181fccab2c0b76470b8558898bd17cea4be8901089817d
z49baa510f8da0e6ec095591158936b027da4d2a302e8fc9a657f822704c46cd5b4c90529421bf2
zf65d04ecab6c281f32168540f914872fe3f1eef326aa39b45aeafcf52541a38130ba45e7510960
z5d758521588a7cfdc24ffec2660491a3f447b95b0dafbbb527f355b83f9eaac9f3866ba60f675f
zeffb409ed406b877d5df3a50e27bd576052f6be3d3dba97a3579cd92bfbe59aa078c66578dc0a2
z51b892002bf4fa589046c59f6d9973cc43336b26d3eb5a2a947f34c07bc669bd08d54965786ef6
zb21fb9f4a9b9c00905ea3e54bf188f6ec4ce7630d08e5f9ec3b13b4419d2b8c68a10dd8c15df14
z2736d9588b32a36e30bc68b632e920e7ce124e7dd1b507f60a8b2231b46a4097a491facaac5621
z2114a45d9816598d59e7719f2d8fc55453ca0a5f60c81b5f50cdede68a34b6e3834ca253e7e57d
ze69da6a7697801bfc3a513157f8698f9c8acba7b0181b9b60c0dcf90e1e4bebedc57c2e62befdc
z88f6272772fd93a5fb8472f725406a60b5d7f5db0ce1d8595e90f8e7a17d8696f738d432c5cdf0
z0d31574bc383c7c279ed99da9b43fcff0ee56ecf8d5cd67d60bfcecbb5d0548bea5bf72f6047b0
zd17899d02c1dc5470d8268f64f5095ca91e72c9764c9688bb3d532c88b7205f509d9ec27985c05
za8f3de5bc83d0bf4d8a35bab5a586874258b305e9df9dd7f8ce5f9ef9229ae9b7292adc31d416d
z3c675bbd8c0597184eb776c296aa905481dd8455ddd8ae17501990ccf69fc0396a4d832319a1d2
ze632a03f145082fe2a9b7adf31f79cc633b1c46758d7575e8a904ee953002fe9a1b86a7a8269e1
zb9dc56769db207fba29f631bd00ded4a776664b68a2cc2836b75e190064f28ca4a147164411a4f
z9e10fac5adcd05c19188988298b25025c7e1eb2b030aa4171ecb84d63a902bb4ead23cf894b8fb
za6f053aabed92445f58fe9c8f7bf8fd9edcc5cb568fb68270fb258ad3a3d10d77d220dff91053b
zfaf8c9cdfc9e9dd4d547047ad4b1f9b1480b17ee7eebc848230d4d6ba1322b51ec1902ce7b280c
z514ca991edfeb02bcb148c54e4f0d3562ffc4bc1822c33af08020f16ae9db28e3774a2229b3bce
z151705f088a8a6c40725a88ba408b87925044183530a2edef19b53e0c5a0a6dd0c0959dfdc3d58
z7c785e6da3e0b7270f40c61d00f88e5f9823707a749f522ae258623027b2d1132356b0bad8c6b2
z4db4fdbb87e5285e2406e72506a398ddd54b7feab1b77a5814d0ff217555e7e4f1166160a52400
zdf2f9b6c659ba115d53d4f6a7027bfb6d1faebac4e3a74011fa3c48c6103aa8a6a3a77f614c596
zf7a1ca76992cc951c6a932aa6f0379b73eb70e588472a3b892b54a416bf2b578e6bde9929ee824
z64030564020a991fa8671338fbdb251dcb96a8981d2c6f2ee78b6bb93519a4d6207c49798b9c84
z25e338a663c6480566773e5accb2d61418494179a5360249628f6f362b2660593994bfc367669b
z10a72c5acd7772ea7aedc6f22ff1ce8d1a87b80a3b27fc3097821ab2325fdba2344dd21c0432de
z3168f0c2b26a2e3600ebced57d2a59fc00ef8dcacfe33194fa85907e5f648154da45051e5a3af9
zda0bc2df3ec8a74f2dee50bdf33b84306a1a5230ef3c6d52370eb0be9af6cd6930e6629f713068
zbc931fe8a1959e6db81397125931bcc20846b60994c73773172ffcc2aba7c1394718ce346a1065
zc0dacc7e0f832927c1a6bba2b93a7595645fdd5b1ff2f480284ef4acb0e4a581c23e9c81c8cfe2
ze5b5a0b3dcaffb25f9bd61cd27f7d0ecdfc16665f5bac582c63e2a3e124c3598eeae6a5a28d676
zcaa69d59bf4419b5685ee668c6d5eca4c8dfd16a29d5bb1c669e4c2bad14d16d045ce1f592255a
zdc51eaf8e9d26f3726a46e2849819f94489d9b6554f305d05145894da1d31176a063001d5b2961
z44881718bc6abe41e551f77e710af6b2800b6e7f6d97aef604f6d541f1cf70d50a5b4431027dda
z5bd593d34467c0b96e0b3d499711003248e8fe9331a8fc09f2680ea08b39a58c5db05a232378f4
zbe623125e0534b87b02e624c8f44cc0ebf9bfc517e30cb4814229f926be6ef4c70aa006960f0c4
z28ef3aa599faba1e0933c8319814e66701b06339709cd7eee427c834f30934c928f10083771ecb
z18d4524d4d7739d6acf767d1eadba7ec7539c0665e34f1900af872121e6f147503f3b5874f784b
zd315943e2b7d2ee2e3f217fffdb157b7da9aac075a569246f133c8fba759217c144db3d6a17171
z481889b51e813d527c017e3ec408e5ead379ea39b5a19c156965ffb1bb42dbd39b701737047668
z4c6a29debbc01dbbf61f04e418efa97e35349f77580a7434ce0641b05b87855b33e1120339effe
z9205ad340cc92f220fb7d856ea02c2ddf96b1b9104114d993f9cd48f6f46450226d062fcda9617
ze7560cbbf42d797fce98b5fc43df18c39399d12b3300207e53deb2f655d82ffe13635b2a46afa4
z1d89b0e3d0fcaa34040cb3f3bf1bd26b7ed6086a3d975f97f7958d2651d69299885634f9ac6283
z6c8693d2194c736a6f741608d9903baa2af0694c985430a460fcf030fd13a0ccb5d4d583fc9920
z8dee87552a7a2ce70eaf2431af69730cf246630f0307cb1f3eacec9e065826c808e3d06a47c396
z6ae3893a7ccd4011e0f4489f35ad6b12ca7b50ae687c72b2f612653321229ac76ade1fa66217e0
z4a78c07998437b84049912b16b2460ffae3472463a9ea33690771937eb18df2613b5d868378572
z254cb7e0f0e4cf2119e71228476321cd6274443833a00058646a39050d5f4922fc9b3d9c827cf2
z97b6b4594a888466625cfb14ded6da2c3994218dc393e914e9321acb5d87812bc6e9d4bdd3a0dc
z9e46c06252771efab53012423163fabd75ddf04f73e7e9f2cec6335bf1cacc6855ac9b9ad384f8
zde8cefdfb6e8fff97424891b9687a473e3e8a7103bef4b3500e7230519e9781c69ef366b1906ff
zc1833b38e104f1341ca6874c0842e2ef2322bade7197505496d25a452c34fb9f7d269a86fd5f32
zd3aa431e55c9fc40c6a2bcec1bb99a9d0badb0f50598df19c9643d571412cb9e222be1af758910
z440a4ac9c952a5bca71db05122b2b904101c83eda53dbd5d328f03258d840cc815daa295bbb61b
za345b0b0d71b6426f9002063e50dae6f68f0481eae0ff768b86141f4bf2e09cb4e7b4424b31dae
zb0d390e2dffe172b067960ea0765af9ba2545bb70ec06b27a70158fdbac69009e81909271d9343
z447464a0bfa993bc68bee58e53114b1776128fde618c128007d47ba2037a7fb5d728279c48a009
zd3f104a9871be00aa159c56fd5ad83b256401ec315246969b20cd9acc8dc174d2d2b0e4c67caf7
z7a4a8881528121d08ccda559ea595762707821c94ece4b955d32001c737905a65f84bd3f962836
zb46c61ac6cea48fcc2e01f69b25475bca1b35243495eb76169d13c2bce838a3287c69f5b9ef7cd
z7523c352d371d64ea9ecb52d34c952fb7c06b98661729ef788c2bda6fb4fa949313e45c3b4f79a
z528ef0628fdac65fb19b27c5ce93324df72582dad6c939349ac970e5d1c717f5c1ef4664cbac0a
z3944fb00d73e7fb25b8f59581fe2a0008bd8a6769f669ed5eb0edfeb4b62f528adb1e3c75381bf
z8cc8e692f06fa9f35248229d004a65667486927d761ee31a158cb748efb834e1ad20509faea6ea
ze56c8ba5d43220844d8b6cf67128904d1d590d512c7231700320ec630c2e7bff710af6eec57a32
zdd42fe26ffbb66ba3590b87e3fb42d27901cb8eaf45ff534ff73f6af5442a2ad83691ae304440b
z48bde122d41d95c120891f7e44f2d38e173a12291c5ecd25adbb36b6c70750a71a654116831570
zb56949aa76c97c4934ff945bbb2840457426a052060d49c8326a97085168227b25a1a484db0ccf
z6c02c87f55e4d1c2da2105b2ad69f21171fb6db78a1c4ea27a0c80b13e975d2ced433ef4fdd69e
ze63f7d1ac70b9e0f077aa13758351d36f1643f0cba9fa007b1901c957affff4739ef1d76d5b289
zf74c6e56e40e5a735e558fa4de3141c1c826e8896bd7d4d9ee4eadc4563305fc93e069e46ba1ca
zdd1852f938b0bc760edf320fc4a157a9fa6bf2339b312f79676fd2fd317318f47b20f465f6feb2
z28e2094b3fbb12c1e113117b2f504070831b71fdf82d30276b5528eecc5ea121801fed443d5078
zb5bb588b68cf69dd3a28d9df84ab4c163f4ef4189233cea51caa6d4faeef8feb07803946ab0966
z496533acc2e8950b577932bb505b5365b9e7becf21054e238fd5ab7f037d25ad4e8b01aa33b97d
z7fecd9205a40d0b4553711128e145e6e227e36d725f0ab7d2f805cac267756e425f7e3874eda25
z660b4cd97be513148281a2a8a90f7c2b17c212dbcec832cd85bf642ffff92f544f26019384ecf8
zad2cec0e8114e64a829b2f050a5b4161f46a4e21c72ea33ea94adf51d8120344999dc6ab439356
z30b3282b88a4af44f5dea88f4c2f8e6b8433fdb33d6fd4843129878d1b2484edac807de4f86ce2
z2e91efe32d7b6dd5dfbd4d1ce57e9524d8e52a44bc21f1a28d32e44254b8f94b193709c9e20433
zdbb0f904051af031fcc3ba00af501c8f41bd4d30ff273866a3801f56abfa99b3dc6a38af7d4951
z6bf2a17e9c12177ec270afba671620b867bdbbd77cdc3c14720cc6d615cb2ab3b71cadda2fc98c
z00c605a6f30a10cbda77a89ff1b7f3cbc29dcf0af06aaefd1676541c218b719fbfb54829542907
z228c3181b104dcc98079babb76b746629f9bd18e643173a1716bd4a706ffa46be8b70db9320ed3
ze23b5fe7f35f4164a6367e0fe8ba056e1661a906c1ee72b49a162f11d795a55ff413260ac8747a
zfcb22fc94b4498f89cf11ebabf0903946799a6abde645bbdd6c34c9bb8b3fee05f1e017ec812bb
z8657ac624032c75871864941b017a5e5f7c4fb70bbee3e62cc36ac1b0ffef57c586f0afe4e664e
zba7c2379483742404f0662c0f960e88bdcff77aa2d4822e9095e9aaf004212892f93ac81a1bd75
z4f7be4e64cb0a9cb77ad223f8bdb416a0349c9fab2b1b920fa599ed9f07548c21f9e06934bc7a3
z5ad0924557776222ed16756cc85f6c7699ebc268e232eefb9a19676d7f5ef58f07c5704576eaac
zad759325e0e0068a180a4e768aebc9571ba8ee21e852db533ec2e2d24caa00e02dd8fb4ad9e64f
z277cf94b8ca0b3020b8b64d3565fc7c24ce137a092be4415e2cd88e4616d11837efe6e5e4839ad
za44cfd6dcc35fc7c9bbe04205ed58f270ee506cf53bc5dacc627a3393cdc4129e36227f6938618
z77a474f500702b8288e0220a4ef05d814362460161bd3bd1e67eb313f21fd8098e9e112a8650f2
z98822c09c7b456568e716e747efb9594a0404fb3c8df02006f0f5f978176385df8fdf1e23a1305
z776feae31f7b72ef4cd2bfce16292d173cb5b80d9434acab096caeea90ddc875cdf435a9a19b2e
z31055284e09be0fab4c1177157a2595bd92197e47c935b42bd1f9e75c139e534b972bc0bb1a8a1
z34fc0697aca7bac7b519f34321ab3889763f693a7204d48f66726383879eab1094dc7d1e92c07b
za4d9e218c816ca8dff64fe50005ddfc1ad86c270850b1d990d41fed3c0858ddd77eaa5b96055c8
z451ff38c8920446a91d80ac28d2b9c440a5f3156f30fa0366afd711437ddcf8a7ef8b985f99cd8
z2bc7fcc660651bf4bcdb34270a1b3d734e5b237f32de4fd61daac2483a52efe6adb1e5d0bb3e38
z87907e714adf3d739f8a8beb46d7e3be2070a8503b073820b8b7bf1f97958e62efa5824c3577cc
z5b2dff0d464d8ce338b13076b3d13d33e09cc2ad6bc104f6508271db00d14fda02cb339766a2b8
z0468abf9ece6d6b811681a5c74b6bd79aa2e172e0f0eff9e86e4599e498235866f953e2aecb2c3
z364de6226720d0a45f33e577fa570bbc788987e8aca446a70959c46b72358b61f861d9022ad06e
z637ed18ead1799b2a3b7ce79f4dd2a6ffbc74a5edb0219aaead5e831150e6447a10fc0628b6fac
z0f156d15d67fb4acce92633eab5bec2a385845dbdb18650a5406fb4bc7a4b4804afbdf21b3d55c
z6975e0dfc594f17c1cd462987c6c590d12ff629fbd99298556c13e7c46c10d02097b479d005b48
zba9e9942fe9afeab8e5b38aba9f83969abf53b355d5786643deb501b2eed5e5d0f65b182c2eeb8
ze3a900a9456e251c5716c37d2e01990e9e0c20bd8cedfe01716ecce46ad981af58759091f445d9
z6c8282ffb130e1e22ca78d838fe32f5773d9651c8421cd6c81df7096c904144d8f82f857886c61
zf8f168ca87c7a39a3cb05abb7f6c12879932f2a05c5131d712951277632ccf471e941beae8b28f
z6496e29d199d86c22a7cbdb09105283ad825104f27fbb98e4d207685470d5af2012e49fd7cdc99
z1f2fee6f564bef1ce3ac3d9218590d6c8b52eba5fe56e92db1219523997761632b1b2cb4015b54
zb0fb8652f9f9877b0d40e8be8e4508151714dcf82de6ea033b9c19b7a60a70252191002d49ba13
z552dd0c08ea9083ab2d02ab4a3e59ee2ec4a16018175e1fd1636f8b93c30975bd7502b523f9292
zcc99c2e19fcbf588014d2a5c267de169a7815c6078b1b7aaa81873e6523289c7d6fab2f0666185
z64bd4ffea78bf1d488ff6ae67e9f0b8e782d6629883e23401a664b5f2ccb556fe9c88149d01622
z3c0850bf347fe22c88163f07fe0af8a43c5f68bc6d608ad31c1ec90de3bdd781ef8dcfe7593c68
zd5ba9f2a3b88198a23a7054234b8522a68116fc8ca56d29c735424f4cfb89fb683132e0582f243
z88b36b80c995aae4457c886e88b9cd41ed809f30ef52a185ea57474f48783d1a01c8c8d80bbbde
z2d6b93e96ebacf1892f80348a66b2333fba952ff3e55002773778250df0690656d8c695d5fd7a2
zf2643eca7003e777cec1dbcac1ffd7c7714bec73369bfb1c5e57c23e255633df055ec77bec34ec
z06b80af459a40f7ddd1701b450f906a2a90258dcc411fbcb92eced6342d9bf129139d1108d0bf2
zc50f4ff50871698d6d6b5a9fd5a8aaa9d7c47606ad3e00fc8559b99b3247129564da71564256b5
z5b81f6a6d9255cf82ba824c3c898446f7c6fa8b56521c640c54afce4c05fe9fa14e9075fd1e87f
ze6b0512497f32413350925311f6f582d246647046d216e3c8daff5a0ce0e8b2f284209c2211c3b
z6a37bf627c15de0d4fd38a6466b20e3f42240310a2c2c7138cd59814a424bdc8ab34409fc6f1f5
z135fde1fc749587fc18169798d6f36c75cec3bbc49190e9f1e11c6ab69de9ff256a9df6485b248
zb03259e4273744b30e074cb844968aab742b6828348bc255978a778b5df1e5fc4da35d15b5d3d1
z19cec2cae18f4afc5b871cfbbb75caa213aee49f38527b947550b9e30eed34b744d7f5783cd8d3
zf2a916ca303142b1aaa2b0acd9e488a62c5264b3d54218f4fd8fd2ab1a04b5b14c44bb5612a3ad
z281ff6dad36ca3227253d163e520cf9925634f8654c74a630edef151a0a39df33ce2e657e22498
z15ef1f3074a03fd0ba10936d2cea2cd8698c6b34f5483e9e5237407303ec98a940d69bdcd27531
z23a625d76cbc4cda0b04729286617c0813e50a2545acb79e6e2c230979a992856dad51176060a9
z3332746203844eef73a18dca0944c1662837ae21a9c32393c7d3b09549e8e878615dec56c51ce8
z1f0dd424c8a93c9b339e22916fe6f0749f2c9c450006a9270b99599ded5f248d45f2525c233d12
z6937e185bc2c797d27273e0282df12f6a6ad22bbcceeb05620bf78f05a816448086fd7d276a2c5
z88facc0eb9634c7f9bdccf6a42aa875074645a520c8ee17439e0b06afc7f4324ed903376957244
z45aa7d13b4905c063bf4c7a47dea2763ef73706f3db781964938a3707fb5b04d7daeb325ee2bb3
zce99dc45f276ddb4aae6ad574875f372e38d87d4885b635199f57f06633a310c260fb415a0e0aa
z3f302717815c6fc050489e3d1e7ec09637feb5a2a5f3e2fa896f4c0399c05987cfece0eb6fc4f1
z4e18db5c85cee1d810dcbc5d71c89637cb2ae022f33099e40b61eb499e9f2ff2a601614121cc89
z593d401505fda7547f5a19f79dccb538150081a793d67806369bed9548384d267baafc6e8baa9d
z9ce03156439fc85d4b3f7466d240ca74c092e3802d49835f62579b8612a29fa3f1f31971f9fd08
z37ac4340a72dea00deffaacf4672b79f3be97ae20f42bd0ada63b73b11d388ec1d3f9f8ae75307
z29538bd84e0fdfdd1eea4fc97b0edfe5883081a57753173ab2db4278022235215b835c2e1b8ea5
z51a45523a55c986a2f28a4ec38d2ccc967a5a0c89b70da7fcbd9dccb6d9f30e4548395c5f0728a
z2d46b32d0c898f4a34c495bb13668f77895c0ab4647d1292e0d327ad69f135237be54d26d60971
z6aaeec4144918548ed7c9ba1e9018f2851d33da608e6d54eac1e296c34db9366183ceeac23c690
z7682a0fc4c852d726c384666a48aeb75a7900eaa40082a23248ae7893138c7594ccf3e4f207ce5
z819c2aec44302ef3da01db7849267575a2bed30bcd88c6f9d4dc121fee286ed425d8b262b9f8b2
zbcfd343393a8ccf5b88bc9adbeaa785d83271bcaa4f49390c25c0bbce6671fb1f167601d0b4931
z9dc33f4bbfc3b8120dbc188aea9c33b58fb3fc70cae769f757b1672e81460213ab158198c76778
z3695710c220cb3a11e02a7c65a00e00a9701e08ff09297d2e4b6cfe9713b09ec01c936ac90644b
za0bc485937857597e6444c1ee71b1a1d99058601fa524cd149cc7198a9bee849051348ab840eec
zf938781287acbbffda4f809530fc1c1dbc941376f55671b19c1cc9d8a771b744bdf23aaeedd683
z5d299f743c0e1c8f999e1e7af6001487c608f018f23efbc6a3d4750e56e32a75a1d5034708d530
z478e988036f9fce1519a018bcb67105b80746f7adbd72051b8c37d143b3636ba5f19c16f6bf486
z3304a71efb86ef4689a3c01f8d71d029343f330527d0e05889828690e18ab99fa7821a31879906
za7baae02684c5a287c0ac30079d21e016a252202f0c355f8751020389460ee4ad0e37594bd1ee7
z3e3f998f9f3ea99a0249459261fe26458c3e2cf241fc873057c7405a482a1c352c4b6772dd4835
z06d7261bb093d4b402a11b78ce18f6e9e94767dde6f6f39189db4270f8660bf1aa48e1432810c0
z62f14e80c9cdb380994ab732147e16602b7bed3c7e90d0d888371408ca27b264d308b4200b5b37
z1093ff0f792aa8c857d16a529753fade0ba2fbcde73da4c87a5be6a5c4adfaa71d864e8c913c26
ze7b4a5af6c287d51338ef9391902000343ce7e588cdb464a8925554771e6965abb2e2946bef041
zf08d7aabab0433ca63967499c35062611593bb08e298877465f003916581e8c65ccab681ccb2e8
z9154b3049dbdd3419e868c0682fb712b5d3abb64f1f2c9577c1b7b9167a49fff04965c492ef2f9
z16304c8ad4a0ca816470ba60afc10141e9cf0deee209d64963b0d10bd0b52da6ec7941a8cc7f96
z88da6a24abf9751e7b618ed2c9143d84c22318410a60fbc57fda6758ebec200ec4f030e02dc890
zb560630389854b9b64c7be4ff236c81dc272064e5bf197691808d6f536e92703a3a203e7a8a5d2
ze3cfd33fed7bfa75b9f7eb82901d643f71f30217a2af98917c055a3c49829262bd9cd524ec96f5
zac1a66fb65676d5ec428d627f1f8aa1bf8d03060a3c65bbd29d5d045647605cdd47a68b0d7a10e
zde10d9635582b364ba527d78034abbc9779b929f7531456d6f749fe8054a02b40690ac7e6566c4
z4bd4a9b27430e65d7ad31c1335962fb3bab2036fbc4b434f14fcf448df40db0a84168b898c11a7
z1f5a1adebe7e23bbbe58e0492443f0cb1259aff2b5fa83aa5ed8df3f182c4ba3f0e4830804cb16
z7246f723d576265168fc0bc52180cbf0388467b5e1040a817b22473cf6c630c5a28b456d589c51
zcf1244b3b933b4ec09339312c80a5ec17c724ad738582b6426fc46daf6cf6fd0393ed278099d02
z88588407555d434adcc33670d48c3b77a363319823aad848360e8b333376c1dc6e20508c295670
z4ea00af157d9480866f048a4fa1795cdd9abf0e1def797ca9aaee55bc100d1b7920f2d450b4d7a
z4c541152fa64e8541eec825f0756ac015ca36d27f01b72ee23881ccbbea47d3a5ee8dd3984cd9c
z7db230c3655d8b00b3606cad8dbc10c403c0a42ddae76dcd10704707d10721f80bf6f3742f469b
zdc496b55b24571e821cdf3202f3f9f05a5b5a4439a0489ed8a8cf2b01f8ff28d57f8b054842a47
z0d3482b1a0589a6aa6e2057008baa4cc07017d25248b1a0b72b04ec09cbfbf8d45a0e4ecb9f1fd
z4746c418bebe69d0abeb6ad81db056be0804adab5372b56fd42fc26b4982a274c02e11d9187e18
z95c1e436892247d61db8ee966c48ce828e48391505b8eb90d72cfd59fc56c5d524d86c876e8269
z5380fecb754a010cbc84369035d761341529942b7096f3ba1f7d8288b326ea73a1efeb5cdba217
z402180c61dc8df9e9f3ef65dd2b06363e489081d2499af79e5dd4c108bc1a9a3393fe647a2cc03
zf50460fc181fbe0bd49c53eb027ec2fa406220ce21e89489cceb4c5e71a9791b69bb0822e06af3
z6439ab0adb5560a75b1b0a3b18053b72954c6edd130d033556e9eb477d41d34463a294d1603256
zb5f3664d1869bd6ae0eda09bf8aa95948e65ea247c39bde0058d75e7888cd85e9fbbe6e4f010b2
ze26835a67c72dbf9389672568ed161f530b933dae9a3626bdae7e7b0af7d5823836a8bc394475e
z5e1b7b95f8efbf42d8ad18840bf1b05014cbeb59207d328eb7f4633ccb6eb8538bd6b50355261b
z792bafb8a05c6cb1e8e94d960c00ac239941e4cf24bf1e3d34675963daca27a5fcf0f50e4fc949
ze022b24fa224f11054c8f9bd21467a9ec17def5717b042908febc44ab70a379fadb4b01b48e23e
z9809e7ee50d7bcffbcbf3d820e6f9f9116faca5cb9fa6029a24559fd3441301180635927d68814
z792cc37ba090fab9771915bb4a91ade4b1be748432cd75554936207c369134cdeab8f40ffe41f1
z937aab56bd8bddc4842b3601ef6371092fe383e7ff62256cce2d64935e00d7a6c74ad53695d169
z793e07253342296a8315f23acd562d29643b0f74ecd4022cfdad2d6d8332f0c00649a9ed6fa219
zb774ab5823abcea5ed5e8260e8981cfee12800b8d45f75a3c26eb997c4deb1460cec92d5db6457
z5fa829309d58716566579d2d0a5cb6cff7f97c59b0c20e2ba37b939195042cef0b3b5520f95f5a
z4b308e2a2ed41e9a2fa50ed5ce1e3c25fed3ad8d5db97ea59249ccf4a386cee325a3588f56e416
zca793ba59256035fe6d736e0a47a5c216766b7eb21edc401a48ed395e438cf8b6b86ccb37cb21c
z5ec8643b6f90cf0d74817c01afebf266af86c668d79b3d02c7075d5dbf20bd9f6809e6cd48884b
z3ba3b836d3bebb8e19209e2023550c7e957ad3b156c700c549c4b112810f9f85ab46f880565349
z552f411c7e56ee874c08317c95a2a27eb041def6e46f13c723e0c8d47167d06b1427beb4e275cf
z0befefa136aa5728b5b9892b0839a17091294c719b2337a7990517502ee940782477ecdb6d5bc4
zbbf5ba1f254aafb4c0afdb5939a4877637f256403176e4ad8e7a00f37624085df4a24a73f8e809
z1fa6d9de7c26e06b182032ed5d90f7c559e7da082704e2e447386c689fd7f1c10ef3824f6240ec
zeb4782e4e7ebf24047ef01e8c30f31131065cea70bebeb9041cc06a8230446579ff777efeeae5d
zc2c4356e4093e9fcbdc1d47490c1a6f2d6e2367d4df3ea6c9558dff8cdb16e3c6737a940a93dca
zff38771e655c1b96c5936a330ea2936de41d3b518435f2cbea3e95141de91ec365fa4cb3ed6590
z11e80e5c56b9234392f1b0b670e8ebaf5189785e6166670964b3194e387cea793cedd76f1a7a94
z8af4c82a687299c944cbf93564de8086402f1965864b389f2235aaea1bf00c23d736a2f7c25ee5
z1b5f896b02d95e1dead14e2af16c8c8319bb5b1349fde5bdc330130df333c996a8c34748516d1d
z00ee204af49eea35398c44b4f0863357e7fad1b64de8dad30d773eae2b8725203eb2fb086b6347
z24d3b90af959bfab7762e9adce3efa93372aacc4b2bc3a2692bf555f308792d671bbd607a0e146
zaaab9d554ac9fc332b2954992b1b666f979e7cc4029c2805058e4fda7cdca12bb01a47926cf668
z3c4e01db47c55e9c8beefa0b3612f8ed3aeee8be473bd40c5910124ae98bd21f4b1da2d6504d30
zcebee5b442bc3ba8d64dadefd9330d785b96b0eb8ce2745757c3a8e28381b6462335b8801d7b05
zc91ab56d209b31b5f40b00100efeb531660e243c8afe2de323c5e0e4dc5e40c1a2aec788bae7be
zad6df54bf15741ea61c20c00046ab77a09df036b6ebd77b43f242ac4ca7c6c3ea4fe39cfd53a3d
zfe7af0a42c3cc7f31ce79af6352d9e5a514ff89e994124b35474c1b982e6d6f7286f81bcb16875
zbe2e723b54e4c1fbd1f871646197484b8458cf6429a4b8c5a9736019d42f9133908ee0627e8b0e
z3bcf082978e121ca69c112d5f1c320f32820c1fea4f8079cd4062fa02ac0432cf6500aa17f4523
zb647cbe6e131edf28df7e8dc953c1d820582ce11046c8be7198497eac6b4551f58c67ab22ea1e0
za6640c47318f304dbd8f89aec559b6716580dcb13654e332ea3f62a2114793ae0b9e453321ed5c
z133a802feeb5dca9abd4fbf175ab853c4ca43ff302193cadf36d3c82198b1ada3fd2d105c5b394
z80eb8d91afea0635fd59d92acd0b08d6656546746a79e5e8944a34ca1d08e5ce391a76d2553e32
z9328feb8d99086e96425831de2370b722fee03d76f01ddd3e15fd4e780e2ac27c590e7ea0ff94e
z52c8c6293db3893d29ca957d93a24e5db7b30b3fd75ee6193d953d20cb3f542e36e4e73a2af2cf
z7a6ee93de1806974e0e843650df4bec20939804d5ea4050f0e296927f3c2e9c6671b8bad742e74
z984fb6c088c8e469c7780ea829b1b6a5a907d2aeb2c745f301dd29387ab5808a490d2e6eed8082
z9cceff20735ab9e5fe30330984f547b6ce071bbdc38d0c18acda422f2ab957efb292556939e1c4
ze3e0b7ad9471610f87e9ba7c0f33bebc787a619d69e42c655410da53d280bfde3b100deadecebb
ze2c1bfba7e8a354dc30b07ad26864e07d09ac6ddb664ca7dfa737e92d0c6a013e1ef91eb37209c
ze303919bdf009931588ec31750acdc98cf4f938e1a9d2d8cecae3369531c67666c8a4a52c7510f
z334ead18cba8c040c2e499f9133aa59b16231ab35c628187903a657c83f05f255830a74e55cde7
zd195936cd2f009e3699c905573b8e0c395cb509fbdac91754af3248fb63cfe0fb0180833fee711
z7821452713f5f62d7611012298a9dbb869eb1b281baf89039456e2727d9980d98ab88bde30f649
z5c55c828439c14df048fd46fbda8f7cea9f8e8d62795788f8bbd091b98666ac99e5dfb52bdeedc
z09b28ddc3fca6385c3aa794cd9023596ec9d47c52d09257df52e5e4cddba58218923ec2d01bde9
zae89492917b3ed611a0b8842dd9c6c18d8d61b503cd499e0c2fd1b5d99737f276efbd8b211bc6d
z12e0abc7f7897c58a416f7a7496e6b09d6f988415b5b4d71e2a19d2c6eb3146854994417f56f1c
z8845df5d48b0e9e4f39f32263fe0788b48197df2ea6908d870ce9030f04a04a223527e7f9d8772
z569f4e6c3c0fecf8f69d57e16818f1f02eac924b9a5f5e8ea7c95b506dcb8a637127c0ff895662
z7143dd6c1b7398b9a5ca21fe6b1207f8613acc8a9c2e2ff77586df8b9eb5bd7a9872a7656bdadb
z5ddec2ba0d712c0479eb4fd3314ed90276a7b8b48058ee5b9fbec2ec1c2added119d0a3263ebfc
zf21be2772663e38d52ff511c88ca47b1649049feb90c3f69ff78adfd4a6fc9e94ad6eb32ec6251
z40f9af7a55a423b154ab112bce1b9a3bf43f1934728d7848d5cb4366ba42bffa5a702c92c3374a
z6dd237ee841034e4c76aa728c23ef4324b36337bd87654d042e77bac9728c67af534a7cd18caab
z9dc2cf32ae007d3b97836c6e5531d08ed1bd65321df98844655dc3e5546fc2504785c4b09e211d
z0ced8bdb12648908f41e67ae19c4eab2614127fcaa262fb76252ca33978681b9660c2f85aa74c9
zb020e5e2001911e73ce0ff9ba426109c3bf75f571ce0dc3db6d4f62d4382c15639c7b3c665537e
z4303009c64410d4219c46f8e55224d4984d7ae3c4fde2f4172bb58c6eb4550059c6957773f2c88
zec53fc4f2f7efe0696345fb15691f1fe59e2678ecc3f26ac16885ba5cc4724546d41be56753a47
za488eef36287c75fa022427a9e7ae1402f27185863bb53ae51bb03646c966ede7503d3990c8e2c
z85fe235e5752ee068c2ee0e9a7cc8a665276da5a8b78ed25645e34a1006d51149c44b930e8682e
z8456ef3bb4493f53e9090d438dc17239a6cdf5ce7b76420ef685b407b8b21237c2fdb4702ff4e2
zef2d1ee68c777c2ac8f3f7b472c3968d1f53c7620102bb8fd245ce44163e5ca4e48a984e4ba814
z1251174ff7529e21fd8b644d742c8567f12128a67377861ee573bdfc1be3626de3b0fafdcf18c0
zdfaff90a3499f0995f9faa3829aaebc63d8ebf233b0fb23f18f2681b4294206192f84fd9f14c9c
z2bfb588e9c4f5190a16d8ff191dd9f45d4bd32132ca286074ef0889624bd4dc1931464f2b6b88c
z918fc1ef0ee9e5a8f5fef1962662ad0fcadbd86769d18719914a6f5f5c8e3459453f34a9e30e9c
zd9889d776c553f57cca22688ba78bf49fbe3ed77250edccab14e31642ac5325b8f232fa6d5b431
zd22a8aa5e596604c69418aa1c1d33f5562a857ef7bb760afa5022ce837b848a0b6b9603fe9f7c9
z320aaab9b770be593e2004110311e347bdc1ddd7c828ebd939db528ccb88fe9bca743f345ab206
zbcbcd2e57ddfaf135fb3583996376bac2f8ff7e63630cb34744df9ff0dd1b0a65a0e5d27752674
z4a84213044ae7942b0943f095f8ff81345ce63416f33f792e5b8ddfc1ea279f39a0d3907ffafd1
z53d91ea72da311b11a251288eb14efa2c22d0b42edebb93a7296f66b754319e32448ffeebf35f4
zace297c9c2df9213a343f69e395f74fd2997ef78006485779625cac40a682c2e66415a0592a6c2
z4dc8c79919d1bb107b9bc2ac944ccb0bc2c81e5ff03c9f1c615e2e55b1e62df9fca084df58a460
z630d0ae202592ab7f2a538df83f7b13996dbb422722483280658bd146cd67ba475b7e6bb138ec4
za3e35f55d8bd135fb890750183fe74e74b93c2e23bf7d6453376d6de96a62a8461393523715057
z5107eca6954e62188648172bef21276083eddb1cf89ba0defdcbe7fc249c7422c4ce818872de69
z9a50c27aa7b6af210539256b8852d97af3c7e3f15d020da13021c02b4d82fe60236ff77df306e2
zaa78ea45b934e26edaebc8b31c224404571ec0a9ef35416e5c53154ea85cc10ea9f37cfd5c9367
zd238b81a791d2706e4e7a5293376450157d88ee8dbc05a2112eb4c9e0aed86891733f7688f70fd
zbe9a3e26159d892501c28782bd0c432a898b5362f25797469617cda14e29874b621082ba3602a9
z16650b6ced4a8427450fdd3f8df29a874bed351bb0db2aea070bc4c1ea6be644f9038368d902b3
z6dc70d1732525e181ddc9cf7483b45905133bde931d3a6a2f8e878d246ee7175064a0d8c4fb4be
z50be9b9f9a2a10bb07b6af855a68551a479095717a284a051707e417e335665ff3e36a053ad0af
z6e626e383c593fa30a4434161f9e30a995f805a664022e6eb8bd4ba85ae58c83005ad0d2f65d6e
za0104cca5b7a4b2f6a00ab07ab30ee374770c799ae53634ac81f9bc47c31bc5ca4ad472a0e8ed2
z0636f68985947808b7dd24331647ee50fb3cd3ce23d9dd0b15927a563122872c056976e1d418b1
z2a579337596062f70d96a4b83e6f25752eb6a622d7e594c824e368a70e953547d7df10d0f958a4
z39cd4408ffbab0992b307a2679ade81ce9721224a5013b76c8b09eea1efcba47d9e780aaa6d4f5
z541da71b9a4ffd253d92800e9801fd9e4ed5b03240ade0a3478d450f51cb9bc48bdb74973b5cb6
z4eb164b90b480125fb0d477ddf8f453b3ff20bb944e6b7406793e05582d81a28aee26e40503fff
z471573bdaa386910054c07742e7673603579953b864d676cce722af0785450957192153a7b3f7d
zbcae199a9f178086f99b79b2799140f38e22639741d07f05aba2ccaee3b662db4a36e3c3f8ec52
z40e8e1d01efcb6390f9871f29aca336e81b82ce1502253a90e9143e3b1f8eb9933fa9630d9edb9
zd6724c22ae728b2de80f581050dee9f1044b6865b48c90232adaca83262a83f15f4ba886f001a1
z49c15f9a480d7306ce3ca805af5230d9eeaab6a10a5681038a391010640b7d54b9c39099e68cc7
z57ab44ed14fbc285f8265a0b6946388a88446b15d1e6543c2c628724e3c2460c23b4674def4aaf
z0e9d4c25fc60102ada64cc0eb69f6b03bf750f2b56419a58e26fdda97b9cd636dc09606e24f90e
zd805368a7146e9431b7c0f803703cd7ead01d67530aad27cd5d86c953870b3434d839061c44c2a
z4fb6c4dd9d0348b99593e8c73e557d678caf8a87ebf932657184c207b6ac8ba5f32a5f1fd0534b
z3e0f32c9fdf4d2fa5de7ecaaa50b3f6757d969b0e8045656486a550292a65736a8af6ae67ab62b
z582644d4f5c49acd373cd2bf1610281137ddeac41be33f54fb75e8eb31c8bdd89ebd6f73e171f2
z233849a7ee956881b8862393708ce0baf3cab59adc45564e333955a5581f32c42d3705144afce7
z55db8fd78a3459f97ac3630253ff754789c32032b045dfb35946a408f1be69d9c07adb5e959dff
z977bc8d4b94529851a91aab24467895164216d22b5ce7094f3aa96a9cd12806216b4417c303c20
ze22bd171d2e0a1963403bfa978c96e032b429c0b87b51e03b09d522cdab180fb6c15d9aa31f1d8
zdc38d204a73254a1548c535f818e8ace09ce05613a429d08aa0919515123f6b8dee5d4ba25e582
z9e588eee3129b2296a8c3415a9de2b78e4edbc89580a80b35dcb77dfbb54fcbbe4c2e973f54f1c
ze05c7d7c1eb8dc7ba1c67d4ea6a5342f11d69cece1f64e25c2fe76faf19bba7e0697708de2f7c9
ze3c9fb7a3741592f39e54832219deb691414740ee65fd2fb6fff199e8ddcaa0576b84746c7a649
z91ccc3bbe1f8c849401f71a583929151df87019bda2c9814412031583b87a75d47e5d67939a88e
z0d6ae62ee8cc1d273d6771392bdc54f1e6e24ce9e863b9e1379431d68941990c266021e65d6dde
z6a15408c43c69e0c6b6efab8afc57fa4c21b2f436643b0becb83b1d3d2936330df082ae16e999b
z75b44b5aea5d678fca775d2ca7468783d2a18c3c4985b8158a394be95dfc039f4e57b3b74535f0
z670316e4dd5020bac604a1777bddfb182ae3da09994de6821ad7441dabddedaab109c87037ced2
z6e0025bf78e34578093ff943e6831f14b6408bda1e436e8807dea91e2d097ab7204e76ec9a501d
z45fecf270d5d24b8a1d9abe9725ed2cc6468c2c1f76a408db4d029afb15ab80f567e294640a260
z78fa5818ed86afddc41c4f737883aa31e09ad6bb1b791c29aee0ee47282ae8ed8be81f870c0b58
zbd7b4db0158af0e04b79d7eaaa1b87c88b0d0c25bb3ee038efde152566b06c96cac4dcf7ab5f52
z4f22106a8f545b4d7b45cec59f8a6e13a8a1de4ebfb2c5626768170b226dd8e5686faf6ad8fd7e
z020d2d3424a8f1343f9581541f5d27fe5249d3e61d6d0870b170b59a9d0275b481d660b5ba0729
z020157e27708882a9819f420170f305970b018bade92f9bd0720bf07be7728c12a71c047195697
z0285da329d37297776e8bf1c10c8db69ddb50f4ffcdc76a46204793a2ce48c836788aa4aa79c66
zd4300cca2bc8fe6d3eb59c71d64d16e0cfcc4f38cfdb62d171ab2998c621113f4be800604c118e
zc5247c3eb18a3d01a75d859c4949865b7f0758ce853108d1d801336bc84c1df37270c4250dc961
zca3dd7e6cc58cc07622dc9391de2729a5abd8d018904c762c983ab678c212cf9297e8f005dbf1a
z894e480b4e11f0c256f40d7e4b2c7d483f0a4c44aff5cc2c631908c01c59289f74d904822b2b92
zca630a2051ee642f6d7d2a78305abd711ac247c74503e57616fb7da24d3ac3924d1a8c523e419a
z0c660fc1293de4fc92b48c5559423f0e749321f54e9f5638b649a544b0914e518d3e1ca02fbd01
z34008f9655e4ce3254145e89ef0cff28e4537046a30b443b157efe5ef0c98c22b61a24c505f9e5
zf24a3cac28ad3a77ec5ae0de28f95a18ef17f77ed732b06385f136c924a9675674e21c1eba3e77
z864b482c610eec05cdfb9f7bc6478489a2fdc4f5a4d64748092ff5c3e7d7f504423868f526f5e9
z0b7d69c1a5ec73097249f801534e660329bfdabd39f3337d6f2f7edf8988570afda7efe9aafabb
z24ef1249d7b7238a3fbf4f6e7e35d3bb885da0ce15ee5a7aa43754d8fee1479341f1be3fc2ac87
zd43123b74cecca52600f03dbb3cbf74403e1302c97840a0227ac79ea3bbde2849246c1ba5864a2
z5ab19d247077ce3e7f0fcb9e1d5ebb815bbbdb01820daf6246bb54f16cd080a0d09daebca2a92c
z726992b8b486f75c0fc34e182109a2b2a44829c6d9b320f7e81f2088aa96b542e8469ab9397b39
z2f797828e696a01d1f2a7089819038b8b450d99dfc5eb88788deb44e46db982341b4146675e052
z7e0e0b587907064bf9c1bbcc73f93db633c271eb79a72c00c26fb73bbf60801317d19af939c8ac
zda5f22e70eda8a887f6bf6f92557b5bf832f9cac9a298f6483c65ccbe74ebac6b370aed3a8bf9f
z5794e55dc23ec72302c932c8468ac20e92c580424372a1c117a5838f65de4fe57858869be3512e
za9d9a31bf1396f2c26c748e02aba710467f57bb56faead31d6fa9c58e00447e07ce435fbcdfb19
z2b0ebfa8ad39d33e5e352e998d60a1e204a602adb9d550af31cf5af5252542c76c3cff306224c4
zfa98a8109b5787419975fa856eedb96906353ff3fc6d067f302792a9aa18eb47c9b6ce010d3b8e
z4e66507e9c7f62b2520d7b0971095e12fa0901bdaaa6d807f695a3e571af59b6760e89e061be8d
z9d3438394b55835dc9c4fc72bac8978a9f00df6cb11645bdb9f411578d621e9064cf06f8266003
zece6f9c88c6d31006448b90b3fd8dc3b971156b37c40e4dc3e09ada45222197f97a343de09be23
z60ea5b0f55db65a5060733f52b4ba4e64f2b65f25772e188bbe3a937d23d006a9cb4437d50a665
z0609e7f5bc26320c13d90ce61176528baa5fc1d1748021335302adfef0a5ddc8b3909104609e76
z138db16e607b0af21e5065f87daab25b429bfd7df5ea2e22a3e7f23326fa9ccfc701e86664a795
z1ec9a9e9f99e016f191b76a70f2849fea673b2697d4188d4d7d9a4790e9a70299a911fe5ba364c
z925e16ef644be073479b3f729642e8ad5c44acb62bb4ea29c512b8a17773bf63ad921c8d47b0c7
zbad839e53ff89eacc4555181442f4e0b96f9ee115d2edb53eb2857fd99354123cadf6c338d04ce
z3059866dc4462ffbe7f98fc77f7d27bd4f32e881adbe82110ff798d9f9740a7741d3593e9b5311
ze0035c120a4a013686feca3e6d428f89edce65ed8072c8fd1912e9837f55bbfb4d61bdedfc9d0b
z37aadd56952de07ce954f6aad8408719ac9ef56523e9b8e97f52852cf8cdb82d8df4dc4eb796a5
z8409c52a6fc6a6254c30e340c44c224ad16de4e1539e915056e2aeac8eb4276be5d497343f39a5
z94b989775615383d657b40c27c97b792c323c090c682e58ffdf5bc90a6d8e0d8fcedb22fca5c36
z8585a44ab804812eaf0d887c10ad96398448566d7c54e78d90fb282b8f85eee09fd8964ce14fa0
z0fb4cb4bfed60ddc17a7b721a904e1d9f0957e092d15d1ee5b421b244ecae3f63efce8bc4a1a77
zc9fe2903d02ca22539da2f9e382cba42f52e61cf841ef83931746b1a348922d2cc767a6624a4e0
z21860fe00df87ff1897e894fb2cd6bff16e90cb7412eacf7fe4d34fe05322638e9f658476cc5d6
zdab07a32ab3eb93484f45f0110af63b7cb996346d37d3e55ae516d060cd5a8f80b783b4d20fa6d
zf8dd3ac308631dcab53c545be2e2598d77d3e5eb243cc69f2b651f937b0e680e0596a67fa2f532
zdbb94fabedfc02d660200b5707fd3dc8e230a8b75973acfbb2216259e7c0fe6a25ec50a9ce30dd
z99bbfe46acc74f93585aa9a73b693e9a4add85daff98c93b0517db6062251db9d46deda5563e29
z73fc643d4ec280de4b2698e65fcd9117711ada929791d7aa0254f0acfd588d9c71d4f61bfab03d
zb1020e6c6ffac119b6f0f987177c9ee9654fbd2db7390c08fa24672026e96534956da70fc2b16e
z58f72efe5bac8cf2fe94c07941bcbe69235f7c8e24e74e3f774e7fd9d0221cebb92cfc80602149
z1a3822ce4fa77f63ed53be04c54bad277181b25f09894bae458ca6802599262bb902f08f2e9f14
z26daa168fb6f3e527ab98d78713d29d948ec8868c7a67ebc29576c1780fd3e104a2411f80bb41c
z0df9e5ac5f6aec312c925f89c3de654e2510fb68a4c7993bf92edd0f42b42bbbc122a2568b2225
z512eeda22a4088325efbc69bedca0a241f0560f6ad92acbcab89add54406b8c2607464bb867179
z218d14911fb21d2a13f977f1d9740f47cda5769c0e9c83fd04721f39885e9fa47df1cbc411da62
zf50f546b03d9e9437bae28c7fd86f40399f5f60d58dddeb171cc770136b459d5e3fbf8c6a5cc01
z84daa97bd0d4eaa1a87fa6282575a849130933fa1ed3884291839ab521943f7568d041746c3e72
z931c7871961936a3a3fffed3aee25ea0b5952370cb72f54f62d70ae0c842ea7113eb644dcc0d32
zdfa7f207af466368375f4fc82204d6102f209948e956d07b5ab7f9af0fb18a5d46b652dcae5ccf
za7bde84a2987b713a24aff729889d8adb36d49499f61c0d3eb865ff4f85373442d64b5b261c443
z0d4aacfa0f8632a9f11501587d0a4eafa63a511e1595c6a8ee997a49cc58a65df5867f10452d4a
zc56397a3b2ac291fbb4e370b05798b1c15dbfd4ef1e74c4a4904bcb7b90791dfbcd92d789f4b2d
z073f0f3391c417511eaffd4db35941e74b884572f51727b2f15d80ef46fae82cfec1d9ec6aae60
z111c6f7363b628c64c56ba13aec23a82ac08fea4b45317d9bd55957c07ca615478cef062271438
z770b4a44dcb77eb9a653cc10eada1ee6200c1ab09da02efce54d554c5d824d114221e32e90646c
z5172f68249b2c900f8e6a8f913c4846953d46745c11db984bc993bdd4e55fe977fcfba9c1c5dee
ze241c89d0ed110aa3063e579f4dcd01e0c761a9fde65c4c20f594bc554465f675bbbfd82f5d16a
z9e767307181fc56b43e48e9d3d899e6b11a6a2a49e649a5c0d1062281daed40f46322e9e091c39
z9775f7a69c0be10f546e62e1ff62cf660c6cf5de5b4e7613ea65131dc04530cf2180846b2a0701
z7d9556317952ff26836490463f2a4d0325d3ce01246263e2fbde025f583e222e4eb0d19da7dc5d
z868fc7474298322225e92531413d9c5ad80abf853c71a1be44eba3bab132834d64f4638bddf3a8
z6df9874db890327a88c24a53b8c58f9ec9a9dfb8ce346841e7d9f928961534bfe368578cc3a138
z1c3a9285d7a4f732ce4e391689ab367e9d5a85263c95193c8691935476a0fc341fb26c3a36170f
z3b8859983601a5a1170da01da2a9b53e6c12e480b065f121ff1f125cc152c3d959494fa499bbb1
z917e215620c80024b2fbe0bbaa64c75c07167171b047f2fb3ed85bd42bcd83658347289dba7350
z2a2f800421827bff6afc6b95ca5aa166fe6e789b984209299fc62215cb2fc4ef4e7b6d1504da5a
z2b59c4cb9c9e318579c418d3915cdbf033e7a705e30269a047dfccbd74d64bdb68e06dbfb48a42
zafc465305cff9dfc57e61de1f0a0c16e04520d229a3165d1aa1a46563e7d68d11b9674552955b1
z19706730648c22087f5d8957fbf51bb981bdf58b5bf89af1acb51e0fae57c001d8026bcb9aa375
z412f1573319e85ffc2f6754eec235efb530549aa9329b06e70e1e6b45034f6283e36807f8cea97
z7d65215b34b68bc82946a8d6092d689f42506a0008b53d09af86958985e9941537bd053677747b
zdc6227021ee0847cb80484eb7c589aa5b55b04df443a3d7336a4aa95020aaf4183a8f32542c86a
z062b3a83f0152f227b8b5f6d46d53951954d81c24e57faff474b8a4c4e9df0c668fb21aa169bcf
za4d1d751f4f2c3eab1d230d5a03962dc50301b087bc195528a63fe7243b5dbb9623b3523f3f2cd
zd597f59319d2dfef68663979685d2d0354dfd0ddaf3d09a0b214a3c2389c7ffee72780aae35f98
z560b15f49def00a746a014ba64160f0ea82287acbd1fc7eb8e2488854737849a0c2fa28a9216f2
zcd1ec901a29b9f492da73a60a07c2e5f2ae2f64091fa67d8168a4b434d4b2b916036496a21796a
z68b6c2597791bcb3e0bacc0e4f4b840043469646116be1bb69296358eae371a200998cb3c68b81
z432005c78e76a9ff6b890e265924f007ba27900331db71f943635cf0da8474d28be16844cb015c
zeb94182e54d24c6be8fc502b62518640eb1c27051493ad452ef245a7db5dcc93a56e7d28ee1d5c
z6d13d8b632c55032e45c406aa237ca301b3db39d6f1cfc3c50cd8fb306d4f6103c5e60046315ab
zf49b2dd323194840865003be44f56572be97e283384d816a672bcac2caecf2d02a21107858c845
z544c37ab91002782e03f6f8ce5b4412bcc4b9b1d9e667d7a03a6f853ca099d3d2a0914da6e165b
z95e07aa65556c2b89b82ac8f0a21fc180783dc42687ec106dd69f0b33848125324230923f96de9
z460ba0129128fd26d85edd3c86a334bd54068a60bf5b6364b210ce9ee72f99c90ec7a80d974f64
zd3ae227f86f476fdebace1af0a5bf2003e9870c210db8198a642311b005ab681459a40a5621bda
z50b9d0988306c952574aae1bf3387bd42535e0d42a9284bf702b594dce7bedd5c6751d72738b27
za57904481fce9f8eb93053824516a284f34dbddad65123b0a515476ef334edda09ff5d2616191a
z4bb50a50d2882b1ab021aef5eaa1ebda9b6c478c9358551101cf3ba908657f13bc5cb917dbdf2d
z1112f15f0d6363cd193bf50ee626699f6f64bd54fbf7b47381e766f2d100c99623fbee5e5db30c
ze6704d48ffe8b8863c16d8de666b4b60ef98ff63f42b8b690144edb37bf33e57e07e5a608142f2
ze902432ec16dcead396a1846e39cf58365c7168131b4c3483082035839c3788cac09977dacd02a
z3f84cbcc47ce7f6ceb836c3ad374a6ececc7d4b65f5a502c80263f00ce2551ee546803f97e7c38
zf4eeddf9e076f3f9fbc68c9789499958e8ef9040b78223330f7cce6fe06c3e01e4499b6d8447f6
zf616b59cbf4aade9396df3802241ae066ededc7c99c7ebcf0e2853889e707f4d83d1f7c0407cb9
z7803973974fe5b046982d4ad2727e192f3d528a4a80bd3e033f458d33b33302d0b185d468dbf1a
z2202a01f49808885d554aaac5c2f8f5a3f091b3e7b3ec66939dcc2332fed986a34230bbe10d547
z8b37d4c9969dc4006e4d03a82bdb5bcba2fa8e8b54036e5795e6d1492b0c7df00497b202395a70
z2f4ae12b0ad8920aad4ca28535d655c00b60860a27718e79e3f4d748f117ee05c403b805a4e02b
z86834c7d1553a784bf08393b5641d115fa99e91fdda19d2f1ddf2d203e68a723769609139443a5
zd8fb48f48e175bfd9e69194eb0bb8ec07ca4c0289c75a56f257cb3ef722abb31e4598641e0a232
z26c910670bd9cb050266106cfb94e5c37227cf1e49e569245eacb8d5dbee59ad23374a42a18f7f
z5b24d108ebccf4ed90786922dce0058afecf3edc0e40731c5ced10890a114a9fb4797e91b9ffa5
zc3562f8c0719dcbb97bc6fdbae25edb379a5f6fd6a6e0fc517fff7d22f26072fab456209fc93cd
z3d112d2f7617128825d459e1a40e9c5a7719d926bb39f3acecb960849c61788d687a27b0d2a051
z00d404f055512a5611c7036e2a9160d5d82deb50ff86f803dd247235476ac22128c13266a5f8c5
z11bb61024d598a622453292c22a741f82d5cb45db187f4280ae68f84267977af302f164713dcab
zfb5057f4101e80645dfda728f333d2b0beabb8ffdfa65597beee6b83165265bdb81b6054ff899b
z4d8f693a2f9212aa42d958c8c524901c0f9c64c8fbf9324e3eb01e9a3462b2e92f7cd5416d72e8
zf9709d062c773108e4ca1a529d59b4f0ae90c4f5db002c62fde0597c50d5b6b38242a8caec6ced
z4d00bdb44f68baa22a9b32faec01b7aff22e992d6f7a82537b14f44fa1173de0b72d8f680b589c
zc429d1b84c03f1bbb3b7bf8249b1db54878c3f51b0e795c7da36661fbd45dab0feb31b760d4c6a
z2d84faa5fe972a7bc8964c83ac9574e53851188332d4327501d77b3d3a3774aeb55f0327370145
z3a24933f5472921c93d79b32279ed09332b5e279d5f1f0909964a34ed6fcf932c167b554c53f91
z555bc7b52c4c3f9d5b1c17e958f4fa12844daafa9ef4bab3c148a80e7b3d6f2a53e7f35f4e8aa3
z8662382129fe958bf4e26928811c8b389c0791c55b218326f6fcd1979150d1409768831643cf94
zc9b66596cf7be04fe6211a7db1f9160a9ccad4f7ddfd7ef48cf8a9b1d49dfa0e4458e05506f72b
za2b2ac56066cc13bc8a45c188dc7ac0f7b749fb6b83bec0b3e47833f1cce5b60ed522de3eae475
z097d75e117fcce2579f261eb468d5fd5809a2c059aebdf3f175bb7e1d4b053be8466ad85729e96
zf2b1f624dc5fbb05771ec3911940cb2ba9b2052ef4fb572f736f5e9e8a0028cfc52a3afd1d68d2
z5a7ee524ab501799a25719f0909f452ffe68e5638f97dc750790047fd210024c21d0b762971605
z0cc87f5ceaa7818518e72f47ae19bace40e16ebd4c80e5c7f6a475e83d33eaae5514991a53bed1
zc5502d60d15564ef96c21fa517227a2d1c15f7d691e8ccc4d89b3f8d02aa9a07b9147df68fa48b
z1bc0f9c12cdd75741f85ad981910d012c511bc9247b775b0dacee02302a108ae5ba703b160f4ec
z1149e4ea47a4ca3514a24562ce995655cff75ba32965fd3cd83b0508e65b3b8807567364acb55a
zda588c1f0749170f67702b6fc6628ef10e302447754448685a96c4e8b8650e9f4ff481b33e6099
z64c210d9c05b51797e9cb75e9e8f06df79828d31283b9f68eb7a80acf67261bf9d67892fc3e6ce
zd1c10c25009d42bd909c58f19ad5092dfcd0b5f2debc08b796ff3157c90dc512d02f480591544c
z9cfb6a4f0675a81f513986fd4de0141c2caab1946e0206766ad2b07757882a12753bc7253c42b8
zba4c878671c35d58111064cf97fb2275aba7f2785ea84029f3d09314e5c625f7f896602035b155
zfe3defe6de29bb0e1c52a505f489789edfaff4856c56b112b46fbb8c48b056951a8e37a39990e3
z177b16b99b9e9dcebbed5100ac67b7c8ffe7f729f86c37413df1917d3ed22f8cba474dc189b88b
z564b44ea3944a8b7c064af324d84caf686da7e3a8288eb142bd259263c191e3e428445be93551b
z7df6506b2890f75c58923d307ff13c1e2e2fb13eff6a101c525b9e1efb454148c3a6a075b9e933
zefd29356cf1fadc63a5f45da1909da1cbb8d587ae8fb1e9a2fb52143205d619f62839589be3061
z0fa862808abccc2df96a0f74e74e7154d8b1afc4c7dced994ae49fa23414e7f3f8da5d94114bdb
ze953184473abe41804048e6c595c45fc72a5eead71b52aec6d48d720f8bbdb0cca7cdfa3560160
zeb88d442258b012c549da189cd74080d8df462a2a0fc0bbc7bd6cc2764349f452d747972881c26
z4d0aeb5dc0d0d4c52607966dc34d219ddea40a3177d077a53c2d1b65fa3e5c2a1572a702338d26
z992d69bde5b002f79ad56a3cb986fd748be0374041e108c3f378be933f69df4991badd31918e67
z9394bf843abf5e4b6020378532135c00a6b928d81f0eef0f76df610834046a0b9936a0e8af3088
z9b38c1f6a77decdd671ee1e3daba65147882fbd0545aa3cd869e103af9a4f13c61e947d48672a5
z89ff348e3e4576dff7b11b970f12730ffa4d15bccdafa63a68bb830fe585bc848e3483bba073bd
z58f2d0cee8c20ed4786c21bc9bba56b0b918c747be6f5bf4d59021c6ec96d03aab5aecac490c69
z8be3f0c428bfad75cd21b27be4fc506bcba55205e867b8009cab73d035e03df58d46dfdf26227b
z5f39cbdb14de18fa238bb126ee48e2e36e45b302eda16ae4ae61d048f6015333390121177984ce
z5f8494847698b0f4bbfeab7a982852eb094d533ff6b19a60a1b81935b6bcfddc0730c941a50a47
z985120618795eb1bfaff4445309579afa46293286b4e7dd84a05d104ae1bb453abb06e100a8f36
z6f4749b760a025742f8f6db8b68fd9a284b1ffe919122e809490270ee395238fe2671c9db1a8d0
z55933ffc0ac00f25788e85b8ebabaaa1fbb6a6b57080b0aa4fbb0865f6fc6bad4804fdd8ca0501
z79949667a773604018c033a0480c4035bb7a60fc6ca3b6037c60aa24996b4abd9ac283a18dc26e
zd4ad97cb103df3ba1cd262f673bfe30e4a2e34df326b9da6c48bf248a5084acd41e630f68493fa
z0290ca3eedc1a8efef1eaa25e28bcc2075b77fa90adb01175cea8d69a414242c576fce30526da3
z54b6c86018fdc80dfa21a2c236ae4f6161bc8ab326f1a42ffe68750bf3dc088c0ec0fcc684018d
z5781dc960ac8b18a1caa756f114f6705449913479a6266eb16d046ec32365da61ae9b46d38ebe5
z448e658695b7b4f470a80e9d1f696968bd377292dc2668da36382e998bad2d750af4f305ec53a1
z108d26cddb2316506e206ccb1b364cc15ea19bced5b282ae8b21f36640fb547fb46b72e47dfed9
z88ff4432896d7187ea86942f5feb804a0fd2e776e9c31a6307d51d6dfa27a1f40f7fa432558b40
zfb9f490471a12d6184d6db683a8b36177dc6629e62e475097ab8f27d18b65b363e9d8d5caf2e75
zc56e3c1b4440a22792bd9b6afe424c91592ddaba19995227e92b3d937d294a211c97aba6f33482
z399bdf312198761ab643a4532d560bf49621833d3d57ad26d28a233d76c34acda84f052fc5c353
z970d8e967a0bc6098e50567c8c7402c1af4fa23c43848501d699148b44730f5efcc4d2e22ec743
za31d8c5177618fc8423c2c0d9de7598bad652a784a740a88a117db493779640be5013a88da4fa5
z058638301edeb69710fe69cc5eda4394f76db61b9901316bd2ed16ed181d6bc1d491e75ba23d1d
z40bf9338ce6618215f1782df54c61b5b448eb72dfc60e376a9a006e9576ab37f0beaa554cb2c3c
z4db028abc4bf182097bc6f585cd22ad2d5d3545d8544f9dafcb73e1ee36329b3d5a0d121578c80
z0349d799f85138c1d9d6f655370ea5f048ff17ccca3e79dd02d021c79a08709fc85f6496f8789a
z298e63888e792920a120314b37beeaaa1aea9880034cd19ef4d67d760607a48db426b1675ff401
z060b9c36bceaa4d6d831cb181776f51cadc696512619dc153d60ea5138c6c761ff111f632c903f
zf5c2187435537fb8efc479a2fb901f618c9cead35fa5fb35a51fd14e3e3c993e378cdc0a7998a3
z70cd8346a20e360519c4a6621d8bdcbe4a7c3bbc909dbe01c18d0410d77dfc2a38560669a16483
z97d3864b37de695eed1ae350f79b87195be263d08d94bdef9e4f4ec72a6f183e93b02cad7e8511
za924683f1929d848abff5ee1207178c357bb216d485b07a8b351f8716a79c7280f33752f0e7f5d
z005832753170704f0314cad66e5e8d4729f057e43753c8f04d5facf7036a8f5830e75296b23a15
z7fb4ac8131102373b48b95456ee853eb312b2a683b7d9c653f80fb47d601d0d89b935f57a15412
z592a274ed0a9c49cd665b8538cd53af1294348c8d9f07d3b6fe39b033a4d16a9876690818ec0c2
z343f79d8cdf68216e2c2a5902c4a49a39b1d2c21ffff17ba8052ee5e3fdd96115f37916b8443c2
zed122b42457e802b092fc7f7384839a1784cbebf56d357e4c335f915fffa344f93c1457e4a31e0
z5f7bf6176d49ec515686a028f7c76766c598b9f059eef5383e0be7bba30b8fd8e3b38a48c83e4e
z9f1fdac855d81438b02d8e3e3cf56523382d6f6f796d790efa20ccb2dfa399b60990ebe8942d51
z8f353ca3498f38ca8b905dced5d750ba5b229ebe2830148dee9c97e87c0b9cdcc665841c0b6a42
z1ade7a1e9325cfd69711f258612cf2fb580b8085769e4e933b3956e8b3828fda36680b48a6319d
z1a9afb7455fe0c640459ad1606e283d9ff3731892a9d329598bd1b2ba535c6664af7c832027c92
z521064a35b0aef31d9a581e94e18448d9333f136ce5679e5d2514a6b567b892e54104c8eeed785
z001207adc0f445bbb8b2ef0a4a0e89194a37d4149959e18754b8351ebcf651b84e8b30937f03c6
z88f555d218707b22aae4fd50ae9183f1d6f2f90156a09298b179cfd55645485d70e885b3098bfa
z6b06816b77463c98e4be3765c5b5f7db3ba4702a527d97d15b0f78a37706b7d8b7ad55aeb97beb
z0d390cb71e5b389d2166e769dbc742539bccbc517f6682560deee1d3c883d14641352f429201ae
z334c1d4b3bf7c984effc1d5fa076c4226172732a4eb5a6911e50426b23eae74b22a1fe3e362150
z9ffdd47cada63e65fb2028462a5403f1ae1ab6a365ed2a9f5dc3c61291b1195a3166a4749fe902
z999cb88787057b69e1b88db4fc0172b1e23a69f85f891dc316626d1c34659b23b8a4dff0d8df26
z464fe1af5d29f33177e5b23a4df783e5d16a115be600ffcae27d59bfd39dc610e5c02cc0d158e2
zacf6b1889969a1ee1a8c341ec684db6e9aeb1af9d43f31579f681cb4a6ec81e906f9092712e4ca
z3ea9bf489f3c6e92d79bfd5bdf32f1bbe15e3895a95f2a53f7740acb208922c4991ca9c71e409b
z3ab870f026c6b5043dcbcae84c35f9e5ba38aa6c2794e29598e8e80435f17d9a5e2ae72b0113db
zbcd345d86290148f4448a18f7b03a512fa2ddefd7cc6727a22b6500b768dbec7986eb12ae128a9
zf546d8a9c24d035a0740eaae5559e96d0e8a1cff110b8742ded36a32db2438e0ce6b4f2f36296e
z2e888e918b51dac9636b97be7b8520aff32863ea46cbc92f277387b7782075264ce581fe6cf9ca
z8ff17e1a6d710aacca82ec2637db69d8ca884ba35c8506f22aa4594254b57f8ac10b80eb7a2534
z5dc2cf2719da9ae1d4d928d4892e8dae8f20cd4abee8232e07820a71ed59f8ea252c3cccf0c736
zc4ebc29c3180abd50a62ced933a9b15073fac053910f6a9421fb2a486fb54726828dbc86de2e7c
z03f3e2cf2dd4846dd33b1bc1187fa2d619287292e3acacae7e1a707f4ea2cdcbf881fc6a7f9a50
zc9eeece8d974b174926c7fb78b85a3db683aaa80ab0498836a71ff2664896367d2c9d0ac0eb0cc
zd0c25be10657a5b2851303d70ba0ffc45bb8c4f75f2848f229cd3f2fe056e3df0bc548f0913ed5
zd8a5ed179a12fb9cb9361f2546c25482c5535ea9fb90a68bcec24a28679db940a3adfc53300ae6
z72b68ab7037c210cc72a445f59be41ead9a05c330c463376149cfa15e518e7c66794f10bb18682
z41291e1139a920e9eeb4bf88c477d8f170a4ee63e8d772469cee1028a0f0c3d0a58f078ceb4401
z91a5f4981c5bca4e2aa6bc27b537d7bfd1b2fa5bee12b5928e334c9b090fc7acfc6d2167caea7a
z9a9db856499bb0bbe051be8b998a6c73f06b9e0b62d6add8be5ce7c5b653b1028d3abfb712da8f
z2f75fd82acf15e5d41861c075d205dc351428a0edf4e6421a5cd5f5a287f30c3edd2774cac406c
ze71aae34f22ba7c4d975800b5d74368793cb6a8990688c9e592b955b05846a0b5ef3c9bf4467a6
z92df4489dbf4056039fc6e2ce051595248976e3fa78d5a680771da6d56240d772bd4c9ed8850a0
z24a889db335f7b05045df52ee69fda95e63afe365a20f7a55c6736daa5a3e23c1a3ebfb4c2f8dd
z557e2316b17acc0ba089ac393fc676331da356b44f0546ad00b1e81599f238cfd977c2153f930c
z12a9f09360d74665da22fb01ecc3fd910a8f10bd7aece84348e87836612d4f5a1192be5480289f
z5b54acf94c3e0009c2679d23e4a21c2a6869df85bec501faed2e3b75a791fd73de1fbe94980855
z3996377b5f563c04134864da47077a3d170df7910f0f9c3bb2f77036c7c416f884fe602fcba280
z7addc54319840620778388a5dc44daf76ed1923668d9be66e41f2e58b8481bb4f3eb2895986de3
za5ab02c0460d904cfcdc25e8623430635d8ec9f64d95560642f430b08810d551ec929928f2a3a6
za08d47055239fff72e729dd8d3e918c3eb6b4c31756324428158b98189ba3f059eded2f25a464c
za8c3e72d6702228ba96f0e3f16913a928125c9e5b3d63b7cd6a50ae6300210d422de9c0ec75458
z9ccd0512f29e54031faf0968e758bb138518417135f0c94cb363d777b42625dc25672d5304103e
z85bcbd4ac96c9e40564f55ea040162e7f7b615b38511ac15ff945d5ed972e0e00748b398687142
z4e0087e29e1a6fd870b88cc0674f72ba762b15473cf468c86b9d043e4630e958a0dd3032fc33f4
z7f6bb029985b4816d498ed350d5411961df58645bdd46e031acbfa3edc55853c153e29fb365c3e
z2ddaef9d3b27ba9dc26c79e3418505afd06fef69d7ed5edecf525de293f743dece3bbb7de8f0e2
z21d35547482ce430931ccc9327b5ad7b7bdf4df9d48a0e6cc3a72458be44ed2a2d060e4a3f53cf
z3eb775760373e37cae3d6b1b843606369649dace798e2c865bc832b00481671407791841348398
z3e7071aa25b24a5cc712251759b59d6e804bf3f9936c0423d9938c7f560737e02af39f06378255
z657e56ceb73468828ad04685b0635b1d10c3885470db23242a4257d192c67dc102de4ace78ff73
z0df22c6923540faa389fbcaae8940cf61e468ee508f4bd13b086318c90e94a676a60807104a005
ze62a0fa91ffe31a41f85cecb3f1eecebaa6ea5b05f96346765a985cb205cf469105ccd1b1224c2
z8214294d093a2f2796b8d19f08543b562bda3b8de8de4b019d98e7810599e26a16623284dd13a0
z9844462936de7c80c0f069c23f42b45cfcdb2ec5b7888d9f5437ee29ef742fd5628cdec8c92041
zca49ee5ff2fc1f91eee5d4ee94691e1c60aa75e566378b0144512b0cf5337e1b5935b8e3e7fc5e
z5625a9bfd97329cac453bc2a7cabe7e73e90d8a368588ea2713eef07b9aa5e9021222c5b6ff2ea
z978c0bbfcdadbb27818e1c7346506061cc3acdc3a3ca08189c6682ee0d4a12cab6e6c3b0abf08d
zd2bece67cf6c3257c958e0278ca9949c60e7abecdb4bcd5bd16ddca8307347bda49a683954d256
z1d26b3b7cc9674993be5ba60c79e47fbf0fe41489bf6e697ea6e117867a1d621bcf4f8e0c3ab1d
zd4f0e6328a149437cc318a3c95316dcd5364685f9113982648d6f69080d71329186d0031a9ae94
zd0abc1d972d181a44e888bc307c1f07936f6774eaa4ad4f2b46e158f5f5a305e87231cef934720
z74473d5c8394e72d6322d5e571953b2ff70dc435bc9c3703b8560246baf08acec9738be858d1da
z616039b41b91e02115ac481ace9d6791c960ca7b97c806a5530ac75780493e5a0c94dbcb5bf531
z1d625433a48795881dcfe89cf96a9ea68e3aacd3f9b4b397f776d4c68def6661569dd90cc2b0e2
z50175177e88ad507e4afac96c76edd5b8cdb0bffd5cf7237ef78c8930a7caec4c63572ba6f84fb
z97ebd9d703a63b6f10612754ab61159fede66308f7e6d977690f6073351b74cc2416756e640304
z16918f682ba18573745e451ef29f668a7355bd5c3072cb401bab37520db3a4e5a6165e95d87772
z06562cb032b23e13413802801c66fbe99c34bb95eb2c34e4fdc64c93da8a8fab1e1b939460b36a
z936e51e7137da3e9cfb4c989df2fda76f53c633e116c42173a00ec8b7357ca2767857054909c09
z36a553dffa487ecdede468de0b35d6551b5abe9cd37460ce4ce3554fd6ee34699b600224e30765
zc3a0c7e619f3211b6bcfd13a4b28771bc22025f230076fec7a8733a13fb40ca2c080e678d71b1a
z3f2099283369201236e93439701506d18c7d6494e430e55dab5379112f8a8918ad0c774d50be0a
zab2093a05d03b4c05aff283e5fba7aa0e3d599f9fb810d4c530d60519a98118736e0cd3d811cbb
z4bf3baff7e29a52e3caeb041b344f4198ec6272a71af43db505ffc4a083ec25fb2f0589740c92b
z3c109ef56c5abb72e9c3761b62c62a1330a01e496991827764c755cdf2453302ef8f12da730586
z90dab587bb0a739104275b99b6b49446eee4d4f4376f8f51348911bdef93c89f5d2729b3e9e0a2
z3f633c6a8c90eac59a2bdb4e77370b9e65feae8fdc9fb188a364140fce42c0e154fe9253658d01
za5655b3d52f2064a3177f02d339ffcc4b26e12e2e8bdac2957aca6ec8e8eab4517484024350ca8
zf30680d0fd615db4788536d97f4c2700fa519d1f6f657c8fe90bac46f775fd38ff191bad849de1
z536df455823bd127a32c9a77ec90b5862ccd6540c9a019033bfa0269f0756893fc536d8077d9ac
z90e5c1699d5a0efffea7392d1b48bce6f75e733c702123b158628d068cba6d135d1b2a787d98c9
z7d63a223fc87f1009100ce1f97a5c639daef8142cb772d8dbb43c1be28ce5e2ab01903a0dc75b8
zc1ee5a516bb07e1e2b70c2c504be8826a1527f940408e0a72b355273adf30b79d449d5fbbd56aa
z47125525252e5bd660db9573b4e1216575ffb5eb3017cdb690f54d80f51655467afe7964a23fe2
z39b1daafea3412ea53bbaeddcc950d926b143240bd9a89d164a01154daf4e4ed141e0eda9d55e5
z44b07ec95b157e676ea3d5033dcb1dc341d7fe345ce48f0f810cf535397ee8133688579f74a984
z7cc7c499ddf204843f41e44d6a5e8dd5f0c41501aad78b413aa73bb1fdb36bc4c4fd6a7ae21e35
zbe9bfd9eaf98c2d7d3bef411c05089224d646c7d12d8cd997171752e0ff384d4b4ea9b56fdda9f
z06171b02d1235a2f789ee83e0575cfb1f31eacc6e4ba1a0d52c2cfccb4a04f4629eb32ee914562
zbeaba0b053195c3f6026a91af128840b5c2ef0a19f38a36640ca1f2889b57dfdc05ea8b3fcca3e
z6caf277f0debe8e04387db8d435ddfb276b8a998a70d0f50a09a0606f905f0f3e0634ca5e91e70
z82aad375b0b22f5eb800609d5d5d573c01e8fb372d111c35b58ee412f614edd3fb9f2ed99fc790
zac2a0ec5681b8a61e1c6a81bb3928a32bdb1f33ea87b47ab9295b072a12248aa1431f1b66080c2
z5d5863ef4972d0ed56e44b11a1cc014689327e0ec851469df27eb53a9f638f949626307034f1bd
zb6a00b2ead4dcb305a0d3921c78739e2beea3cf3acd3e235e5b1716497d7bd2b2e42d96e288336
z55de5602b3ccf885c9b87364e6f605c898d85251e472ce8c4fd20cb0b44347a3fb324577e4ee91
zca727631c88391701552aebcf129808b369c037f46ddce3edb7ffe1a1078a18bd78a8e6bf9f812
zce4ea6fbb992cfc97b224a9ad48439fa76c6f3023ccb3a990a5de7b7f0d06981012d1b49c42bcd
z9d2028f8200209e69b8390e7c00d425e52ec108cf22276b5685d5d11131ca935e451984ed56682
zc5f00447631878a64d4787eabca7e6ca86433a4f6dea937e7fecb6580f9e86ab050a053677c4b3
zde90356e2ec0af85b3151fd4ed57d532757094b7c3889356fa7c96810135ec6f3e5ec6ace64bab
z40234ba85c000ffcca15dc7945f9f51e23b9c6342069d457bfef6539ab9ed080ea60703e4a824e
z2844241112a187c2a22b16c7d234f7c4eb0a5e2fe7668699dcc403198dd4fd48ee67a296ee4e2b
z50b126c51a1c66af2535da62920c926d9ac23a895cfa97625f1e9eee86aaa5f7e531cf5c227318
zefa6854ff0dd22c937d5c227560fd468388dfb1d9e9f8040f459f5f3bf6f6aff2fc5edf3cbdc51
zf49b228f5aefe39a328e1b500f35528c638eb47784f4e99944e2984c73fd489ad181eebd626427
z64888a2204b6aeac2c445c8ba7b0cd22745b3a8699f4049d36a77d35480f529d7aee484b4b79e3
zd483b905dbb2447f852976748d33e625573bc78672fdcfdfc9f93c88b6bec8c951d4e68dc76727
za08126f8f5ef53700afd024ed1a4b6086473acf4e12269b3707513218bec780468c97b6b314583
z05f81d7fd9aac353ba693a3cd598b3c63b80c5e690203ea7ac93acee268eb22f60a760ed39ace6
z27848089f1ff0bd3a19347c77d0bedd26614f6f9af2305a04850dfb8827d678cbb32467680df23
zc3a1cdacc25abb13b27207cbe2d0bd5c1db7a0a7f314076690093c890191cfdd85d1d5b7285588
zd7aa5ccd6e9a3368f526bad7ca7b033961d25177b2555648041e475e9b8a2c670d37899fe5508c
zb567c4c7aa9fc89321198e8f03f3c35a8f24b234ac0aa1673e12ec88bfb9eb9056685ba3d61f80
z95a0c5c60fe16de03f63f4fa41b8dfdd52db900f55a7fffcd0ab569838c16e82d080cb7295c3f5
z553bc9133fe8173758fdb946d9dc8ea52ca8d0f53002e016d33a7905399af538743607194662c0
z29afab91bd97ad7e365900d7d6390ce5fc481a05bf07e69b45472de1d4a1438098444613f55e62
zb978d6a8075cf521dd983befb0650e21b4b5f42d36080c98c3a833238f3dd454a98385419ce068
zca45f0b59bcaa10f0cd5c0f943ad0634bc8ac8cc2f460e981620e7b5feed237db59d898294db99
z228db1875060eb4841a4bbde91b584cb8577f9a65558d25149e5b3781ee1fb4da882e90607db71
z35f1817a9a069a1e629f8a5639e2699656f36b890a548336f808289c1f9a78f8fc464f610b028c
z35cb49e07902ab1a62c20cfee64af7f59a28ab798140a73a36f92f4f3321b28089aa0217a31fd1
zfef3b98e814e6f4cfd1c383129a7610ccd50c3ca3b18a7b0ea48fe815fcda6f204cf37b4f38415
z6f1fbc5afd3c170ed81611d145dd317c8877b6514665a7b77ac5d336b56001913af2dc1c5e641b
zf6020a820e647c77c435ac5a62fbb01ead80b53166d66de6d685346b59faee7b5b96bb56d62630
z1a1d33ace3c335fa955cc791358c40821ab49d433a6eb789d64c742282717769b2837c74cb8d0b
zb888448e5f5860c627d90cb465509884a67e13b8e57ac41c2354c698876ba6f932fff51787b5e7
z339e164f63f4cec479c455289f4b348d6ffddc491cfc0e72cde29ae67956856969b48c5c60fbe6
z5d7629e70f7d9538676b76dc990163f9d415e155d63fa6522a1afc1c842b99d1d15a82ac245942
z6d6f392506eb98dc9da19a3ee595e53dd18cb6a875ab9ef03f2b338bffad6cdbbd3c0fc01a26fe
z288428812a6a838890d817467f1f0109dd2f0de485907f71c7403b03da0f11627e3cdde42d2548
zbb865e59f22fa6d1ee2b1750e4f069c3c08eef61020767f4836e41d572d84f8a7729a14a414881
zb58459656741621f765291e35452d7eb7c3659fdd2bd0145c2ab899f963b159b53c7d4d99cb1ae
z30330f5a5afc2858d7a529fd98b53bad66ab95c83791938a2afc34c72a6da11117e319348ea9e2
z59366c3538394622f8a0858e893f5da58d51af91aadbd432b9d94e13cd02b01f1b3035ea04beec
z22b344884b56e54be5bd959cd2ffb934139085ab5d21e97cad9ce7d637ef34071279ac9080abe7
zd438723e8bef4f3b67305100b50a9315c01a671281486dd441946bc94eee2648ed145c5a6fa60e
zd6602cbb56680aa6500152be525f94976450764a122bb9241a6d96a8c1e13dd14c6d6ea0b07d6d
za4fca941866e0d4b1b23b39a903bba47d942cb938dcc2fdeb4d43d8ec894de2aade8321ecfcd11
z5ad61c30fa9d0c5cc8d8e11264cc91f97e8586c6de1c6b8973149440c9a1ec3e6f5121ebfdb12b
z67cc0aab154ad87ca91a62845c90a3dccb36875768351711fafb7c15c2a4c5d96df4c89acca71a
zcc2aae83276c19f0b21732e6c66f815b886d8dd90f6c5b4a225b7b8b1a6cd25ea81928dae9d43e
z9483807ce138fe61ae07539b6e9ba11eef4fa937ee155f797ecf30f3437f7c21eeebfcee69c533
z5ed14553a3f8ae5129f2d3b7255eadec11d38aa225d79fff55a3a259d16f3f67f61800e06bb66f
zdc1f2a9ad22543652696bb5fd306d4f29194570b5c641ae53727d0c6bf2519a175aca12453d4af
zb7494d6b83cd811b9bb1734c0e73c1b8d38105427a57e1dbc48c6e86350bd4974e5fc50e89efdd
ze513545fcdf9061bdf49b7f81a7f5d086a201d7d86b9400387df36346112d47e69edb48c10f796
z5e043deb01dc4b1faeac5d918b7aa6ad13de9fd2142a66cb2e87c28164a74202dd7a4a0e1eda0b
z1ff43241dad4cd98928fd10206d1c62794b8d47a8540651965e72c31db381205d9053afaf3f13f
z4256ec64432bfc73f7b0db7d57971c77a6c05d5d41bd2a4aea536470e2f9c6de5d39e76bd3b0d9
z60556fc79152fa16121839b2af747634d8a5c25d5553eef26f29915ade8cd8f95cf4999a7bc1fd
ze2b001ffdf558c86aa4e6741ba51dd0843fd90397d2a6774e79455a33e4340ac33129c8b422282
ze804c13600410a8b3c8b47fbfa1009a5046b2e61eaa5c649b7b53fd56441c9c0fecd155cf51b8c
za02b5010d81db247f8d9d5bfb3267ffd4e2fdabc07ca0e018f094bc5f31f477234d43a7ecc2a43
z9e249ae4cd0cd9cecb70dfc492900a7fe14d04132028e867d8ec6c4fe957e08e9c63fdd0c27373
zab5feeff94ad77bdc61569d79795190c4ae323f710d17873a3fec7fce00a27cb184ceb61a2a007
zd9ec82ae97da017335a7f09eb170fbde72b56dff43693b195f138014647ea5eb537de8aa2e30ed
zfb8a12fcd80ed36bd7d42656fded391a027f078667ad3c1d612030446cc969e5bb53f1b122a5a7
z927d6e90af82c551aba32a31a95a4d32be3315713cbddb9f35e1281b685e8d632ed5d2f922cb11
zfd17a7f60295b40b31f94656add2a4b281774df77001b382b1126f87d6df68a79b984f679725ab
zae71cefe5600578cb3620e61e9dc34a9358945d12fe4549542b84c6afd06716d048990de231e5c
z14bec55a624e57e628a90b06dbe853626f52da539bba0998446993569c339cc12fb704480d3c68
za3bb4e694e986c6f615ae1227723ab4782b4e7b506fbf5c8b9d552169b2640f7802543370eea3d
zd3cc1139e07822041507572431b3673c2b4ab8fc4fb9194c44a1121d42e46e68c2973b3742397c
zaee5e37675b18ae0f2bc06b0e5f922472a24898975a8cd5d880119a3c6b441db6dfb49a15c39bd
z8d3e4c1ca82c89bc813fa2f26b46360afddcf3335721363c6a57cc50db206d4f178e231f5ddca6
z6f9ee4be18faa0d7200cacb95aaac6814a40607ff074739be7babb8c1632b48f74ddb9ebf74569
ze075a0bc1ee431ef8c8880e01cd4ec55e533844e8a6c26271c39a65a2d61d7318fb68c97d98562
ze566810eb06867ffa2e71986d090693f7df18c523964c9cc3170783e1e3bd839d45e9960ed22ad
zec74edb7835a7e293625f2ed00821f016624de9f128aac7dc8cef6c2b65027afd396049ad45a09
z5439e67bc785e3f753bce1c0024d7328e7d85594ca7ed14b780fe7c081396754364a8f2d59eba6
zcbb23e24b9e8a01a3505efb9ee7afc9fc50436bfa4d7713a1b173ba5227a4bb852fc52425fa7cc
zffda8341c0a6c3843c7c078b6db1cef58fe70876b29b973871edecb5543a2c898485a7c384a8a2
zdbc74243f387d843ae75e18db968416130d56f44b37964834635b6df59c9d45e83c736d11330ce
z94584ece8e0e25ae4ffc9fac19c87bd90f3d08322adadd64396d78708dfc19bb792a6037e6912c
z65f8117fafbabd2c7d9cc09ff33cadf93352c2b9bfe0b0fc1c705cf182c4f3dd584454d35ac2f6
z278fa6b76df85699a4cb16a7073bab5996ebb79d6e865f1097465e83d33f158c237cf5398b4142
zabef759f985707cb2c0cac8fbd6451abfec9789feeef7e4e4d2063c23fdc3437e1f5b97b58d6a7
z78dd9e81fc4f233eea56ed4d7ce890d39e0f7ef0adc3bce31980cff2e2cd3eb2ba4b9c57f519d6
z2b17a61b5c8cfdf6eccfbf20a3d37991231108462ebf07ee389621cec6fc9521ff528a34cc7dc8
z3fda976bbb0e6d6ecda5f7bc5473c9f5581880b0aa1337e6e26d54b94e2347ed070162e589697b
z1feb856150c4cf6227e2efdc321fdc411ff6a3c0ed1dde761bf6516d2d4afb298ac2ed8cee4aee
zbbfb47cf9474b1ea78a62c98d23eaaf3d8ba62772348ec5e10fb8488c5e1562e6528e59b5b4d6a
zf08a3ce360cc78f20734b4bbbb2d83cf9949d54412251c53ef048bcfc723d3cd75c279d67a0a74
z28771e6060fb13a9cfa48969152bd39dff94eaf028d7f0c284b49d31d19d77ee4210ef1a546cee
z8b09621b2ab9ab93c6ce30c02e8f2b6323db4c552175ce833edb7b4d577c50a22d899afd09ad98
z3d63e853906da5b7fce833f75bdec496708b690eee44fe1a34580edf2b45fefc9a4333b69d5f1f
ze93afc028ba42d53749315998d4d32d9d63bea4fb9d6beeb17ebfb044b47a895d6da6fe2e4172a
zf23689292bf272f30c01b8520fda6f77f58f8e8423807c9392f4e222e94fa4ea589fc4041bc7ea
z5042f154ab22b2bf8679ff9497edbe40a36a358a4950fd059644b2dab74364a97f56fa292c2d34
z8177a80553db3a428797e2dc525b3dd66050207f8584333977fcb7c9c6962154e2710727d1753a
z80b4eb85ce472ef90f2143ad7c5badb7bb2c3016d6b541244c4af00b5ec3bb3bdc64b72d0763bb
z18cc04494feda02725d5165248fed47b0d9ccdbc9019b3dd664f84040fa0bb6b26dee51936e577
z89c96522b06f8e866b050ba5889d14cbb5cdd73b7300fcf0e2d08d57903f6ffd28265527e392fa
z626dae59adad00a7025c24d211e988b58b04c670cb8643e2986f755950b2f3984d226318a40359
z53a41a69f8bd66691a9da07d92d52f4401791cc03f4578fa9331d73eec27e229eb85e80200291b
z94c98078b240605571d208a1a1ee1036f7d05644087bc09cadd306cb945bde3aa07eb9ae85333b
z5ca06df70e6a56a196bd5e2201d346c7b0f83d0ad5897ae9e6b983df337d2319ff93197b6161f1
z08187d94132c7510fa649511d6ba968821e3fadada17e590cc58c44236b6edb48c12b9c4495eff
zfdd773807dc7ac6c5265a75a179a7dbd1758831eadff1158520c5797fecfaf065d1a7ad6b5e2a2
z38c3ca7870f47be3cd2e49616552719a6475717e7e079d122585e9132f504dd92752b390c1a733
zfebcd92977ec018e00c92a7602f0c1a7ac158aa27deea3e1c1dc64ab291afbc0a54dc32424bd2e
z473c6e5d8581463e6e20dde858a410d3ceccee73968989e74ba7173e708a5e33dd9fa58214dd55
zfd50f14b533e71de026852b42b8303dbafc11c5f0bc9d8e3e01e643d333dd4154ba4837740269b
z2e1f8758fe68a1de353bfe3975ab1f692c9b04ba9cfe158c11ffc3ef5e5ddaddb34b7e6a607583
z74a989e930f60d46055c55724b52e1ce32822ba31af04836f17345d5613846ef02d1c0c891a1c1
z76d6d0f7c2d7eb78018ae417247c52fd403c8022541ed06262789a4ddcaf82555c33ff53e2fb04
zad0ad2f9578d368eb0dfa67ee68dcdf757497a485053859f683d64972ce945c0fb6aea7745cbbd
z7d94b9c2fba0739f5a794654f6b0ec1a707764e06ca09e4ce5c414b4d39e36ef6fa67be89c2614
za98d84d8840c15c61cdb2f988da160fdfad863b1f9811ff2bb85213e0e7c23fd56eec35cb94351
z6413150985c31393317bba039fa7aee1cc3ce8d56926f3b87faed181c1a782be1064ef913f2276
ze9e18fdbf12cdeae98486fdd660fd0c30a2bbcbe327e736481afc04730f7ef75a21590c0af3686
z2dcefaa57b560cc941cbf99d798b77a972bec1823a3987ed4d4852507c563d6b208b19d87f15ec
z59323e9cc31638419fe837e15c6d79640ebab2d552b0b509235b6f2ca06ad0b7de7f2c703d5e9b
z68f649d62ad8e44f4d4350b298c9254b7f23a0fb394de20d9ec033cd78692df366c5386ef8158e
z6e3c6dd4384cf92258b8c98002ea46dd29189d22bd00519333752ecfcfa4101b5bc6c13eca6956
z1f0057ddccb584259b14e503ab8b38d8cedb637b205633079009f61dd2c4ab4a602352f38f3083
zf2030a2f775cc3f29c4ae28ef7b8a40625437b93bce8ed27bc8193518ba512ec75d1076c19bd34
za2805283780a730efe61dc550993a6326606dd843e65193c18b7ea4d21a002debfa84b9364a257
z1d5165daa96fbe005cee9a1eccd092064f59ef0d91754ab0689137d7841b53c0beb676e2a5b26b
ze40b40e4cd3b44b995c036e9d8630f7ed414fa3b8ed25221e5c0e05e13a76ebcddee418e79ae45
zc3b165777726a7f344d15047e0c31c8bd2774c72118de36960bb4edca665fcd8a6bc26858fcd19
z7d530e6a3b72f0569167ec038a99a6520f1d93263da0b3a3f94802deca21345749a34e968db001
zacf1b11e6fc933e6576d90bc58baf0bfbd5aed067e156f74718c611cb109b22a2fd4d232ecc334
z52d4e55a1d1cff598ec26364f1853fd6fc622bc9b903b02490ff370deb80f0862464a0cfc1b1e7
z059a888b4150a0b779acb0c5e5240447f75b0247118b7ccc4eecebb3d952eddd74bd8538884d48
z1c54166939aa70a175100d6391bfe56ec05365c2b7a5e02731618042aa52a144d0fbf454c8db79
z62451054b8e485de1087b1c5dbc13622c27a5f7b7b07aff397a47cb10f96ed479efc96a93c56ab
z1c8207630da2d3abe40ac5639bf9d59f250a91f3f413c754d6d1a429f6a2dd6089f6e85a31abec
z3c654ba0c43e0f4e5794970012019f04b0f72bf87a03066c9b2f78f38611c831e45c2d78dbc9f7
z6f971c1c953da2509c707413730c63b56997b90dbc99d8f4f76d9ce366cb8667ee61f0f7559913
zb2e669eec8a803d78d27397d356df50a8a0592cae260e8647ccfc8252c74d59e933ab9f7e6d4e2
z169c159afdc702604e54f0d639c7644fe14b38452478091edf40a4f31d6666350cb0db85040540
zcbde7dcb5e14b9e4d65d306bb0e2b3b9729d09bcc36a764a84d26067313f2bb1a980748f2c9bcb
zb5a08565367afa1959aa9d0b7bda03f0979c7f6e7075f55bffbd06736eeb6244d1583e677ef737
z097f9ecc51fb90a351b91a4df87499d7a58ff3d6c0a710889d0a94888c4b590465dc337c8a87a0
z18108763c277dbbe9f42759762bd6b5d9e90f646e8a89750b5c76d80b8f66d5e20419b8b4353db
zfde5fcd1d6185e661f0102cd57af1ba1bb96fe20603c30f64dfe42585eb71480789a2ffc738f8f
z43124d62d7562a1cec83a03ad105c8ba153f0a0b99e70d7a1047da4e0e0f8b9376f1ac8e5e69a0
z5e85f00e76f7e1463f232f2c504b6c50433a5d518e1ccde68458476b285a6e4a839034d6a9af55
z7f2cf0e77eb5899cdacebc1dbb370c0288cc6f0c28eaabbfc3e37e155e0ba6f862b6e64bf6f838
z85a3370060d508d661d6dc7ae40e90aeb5c7793717d524d1952b1ecb84a09e1b7045e2c97daad1
z1d68ece2d8f4f3fc86f6b6543eb64458f9c2d9d5fd17feac9e9b632aa21e85c15efe5ba0759c47
zfb960e5f023ec77f78e03dc379d9e62b89c2efb64ddaedce6b89acb2419c929105e8e7232be1c4
z5c6c46be0e7119504906610eaff8e7947729cbdf1c7c3ddbe4d09317c99493b943fa449fed44cc
z5731cac2f58c0c932631fd325a81faa7c5cf55e2beecb77fa80a1c0face808a784da55e5a0dae6
zde88f385e851f037829bc90ef36ecd7de7e5d6e8022f7a2b6b1860599907a3e1c39cf31be511b4
zcf0168105623dc752cb3a3c464850171ad0f8fa5eb467fd3c561aa7a74f927eda27095a29fa2df
z0e7fd5ec9cbec7297899904097911bd9826fd53f9c2fa163d233064d05e7fc530345170ce2a7fa
z40649fd41d7f06a991ee9ee2c4dceffda05d6c41541f098e300bf03d63d97a622532d5b6e005a6
zee3b1126514c248c25150e078591ba16fc32453fb2bd4e1e04b89f9961a7647c0a34d08058ace5
zd3509b387196ba519932dc4cf30006f1f80dd6d03f7afd8015e773839199dc6cc1e0e5041dfd80
z85e8acb5539f98caa1734deb2a5ca161ad6cf4d2601e6b7955538b19314f9472ba95d9b3da1df1
z97581b8083471d3af50f077394527e733488ed89c37f0b3d6cb03f6d2dc7dcb9db62c911214851
z05dc84bc2882958f9a900944bfced088e05c5dcd5e6cc3dc0dc9094f8cbc2647f1f5b533177f63
z2d8d2187f9036e20b8aae9ad935d60d217139b0b0a1e375d5d3af24f5eee9520a70fad111f0606
zd05c6e653738993ae4a2c9fa6d0d63027a6af0128fb23102dea3d20deb12a5f50d8b46aaff7b41
z7a9ac6e36ec397c44ed4f320f6bc2616373d7e9ed2d49325f0ee34f2a388fd30ae8cfd24a5dee3
zf08555870ec959fb2c841db2e7eb009f70b43def6b33cdbe03bf5f30048ec057ae70517609f0a2
z20814eb3e8e59a0e0bceddde39ac1956a871b9acdfeb2d421a074293cbbfd555195e47163a0d42
z4bc718a2a5938baffe1dfaee37ec38d03ded7bc2a2ea2f7a1ffd6f9e080b58eb8e31a9ef52e6ca
z79c1f885089b530cad170e8d207b7e33897477678489726ba45b9625d88fa72df3c9ee36c63b77
z625ea8d32d1d096798ade82b368abee2765f5435582ab8f0fdf0d767d218e02c5e1de9f8a9701d
z97002d81b37e9e9ce4604a6ce13cad5515f06f74da75128d4fc66afb1547f83187829f3c513d45
z147f87c1095e4567a67f26b696961c779a4dcf6129c1d9bfd3355942e7f7464bd0c7915fabc727
zb00ab9044330f906c25c4f27f6e5a1f6dfcf8dcb29b5543004673403678585fad9d899f1a6727a
z1ebd4bcb7c6145408945bdd760dfcca6be84e70798492ea4b22bea1ce03eff62e55d164259285e
z014f41d9b59232ec06cabf1983a10300aec1fa3152c07cb36f5bf96abc2ec3fcf861867836ecb2
z5ce48b370240a98b7ad1bf74fbbb6f40d194410ad07f1d188a558e0f21367d6a56a03eac7674c4
z420ff2a7f5d2d0ae1ee75841edcf8237f7d30d7a237f8a0ff5fe519855a7fdb85e0f7c6f514b4d
ze61e9be8075cfec6571ce8fc9a5d6cf79096cb4fdc43e5bdab9d922e6dbe0dbba7d108533c07fe
zdb2475d46822c5284e01c314ff88c3517915aa8987ac85fe2ae79584e4f66e27603e08f76f499d
z5761d4d6ea76b7e882a640051ace66491e742b38def85e985c0b48bc3d59e67accae59cf3de42a
zd9f40d629f7671608a40633dbcf7eb0beb97f1ee55998fd07b0fd95d3c2232bab47692ba536bd1
za5c6528e0a6e5b5be5543a666abe5c01629e3c089b54497605c8e43a9a7f60e1635d199cc9b587
z662d0ce094cda870a280f18816e2cef9bd9780a8265e8979ba7017110d5de390dbddf0e41612c8
zdcdaf1e80087da68e8f5c95bdcb3a38e04e970042ee6262d7c5e3e3eff7c03bd35aac91dbb32aa
z64b9c66adf79cbbfc1eb25d4042d5ed2fef879b3aadc617016111c6a150acb02bc982e22a6f017
z95dfc2101ab462afccbccf5eee7cd2382b8f15398cd2ac854f9cba315cd42b496b8f876f7f01ef
z7d42e70fce79287a43134468c4358a3f5feee724954de0168152153a4626d88e549977e70c879c
z7d91fdd3e677f1cb52f1f829c01ac0a6758ce51cd5c6de4017827c0e8a06a788f4f8855a6d1811
zdf11e71daa9f2c97dc42bd1734c86535e58c2bd3a16e37fcfa76c78e5d91c6fc48951ed17fd374
z6905f52558b7f23bcdc9ec26195b5c8b8d6f254d2317e8ea627033b429456382d025278830a7e6
zad18b84f60413debe763d3daa57b5bbe125321b06e44da7346fa9b0706ffc19859772e1a14ba50
z8cc7f0e5d38f70a28d33d731d8210e08e2928d757a1bce8d3ea4266f127399938338f675cc79f4
zc02070cf0dfc4f4a1d144f96105087c536e2fe1269bb6188d551756d14abb275d6b30aadc98273
z2ba25fedad3ae282e877ab66966d9531895374e74a29e714264ef58da0ac131c2c02e086081012
z6b614d6e6bcc4512fdd8333e63ce31ae82ee0252b0e2e08409e0806cce4e57384cdebaa0f7e093
z51cf69f9420d1b83965dbd1f7559c1aef716c294cb5721bef5a367fbd2ed2c4c44fffa8f9ec6c2
z4868062ceea68c17bdb731fa1ffe03e5c6c0a5772424f8d18868780ec29771e73e934aacd52b0a
z5e7823937dbd78a40531b7d697b2e365e5bec75ab004428ac6b1d77cdb1de0cb1f6b83fc789146
ze340bb92c43c26ce9475e3ea0c631cb471eed515a6c7b8fa77216a75250887b8b5dcf23131002f
z6c65b5af714b62d15dd138679ba2862e70e695cc1265eacda27978d4a19a062717128f2c47fd17
z308523e9d435954f24e66f46dffab4a9ce7ed1d287237c1b7486e3263c21ff28290d2a5d5e53ad
zdaa4f0e1822138c7c13ad294b8bc0db10adf2b114ee2fad77c19d2d1b294dbd1aa3cbd648ed7e4
z7630cf38eb8e4af0a0dd14c052de8c2d9e2fa0968d6ece48e7a906429c487b744c7dee4d20620a
z08b95e3dedfac47d66e6865f75ffd1228c858adca12807e51761c94ec766a8e16293f02374b492
z4eaf828c1a720d62659c180354970716aa5008e2917ec193ff81cc56cbec2e4cd401f43d15e58f
z7bcb26eb7a24018c6820b7814adffeb2e573e4ef626c473f32573b0c8671449ed6b7c3b90e4879
z6f476d121fe2a38d0080f5211d9b4797a8b39dd191b46c367bdb1ecb57ad64c79a0946e4d86aeb
z07f977edc57baec36b007cebfb3767fe90e437177dcfd13c232ba1212b4a571ff89293b0e7776a
z85a34f230d65059c053656e8beb9aef168534533b59325899c79f46c8ed343b1fcd9cc77d0c668
zcdc900e9e1ea22f2176ab5f31eb6c37a72245c26900263e2e0f797796f8cadde788fc8aa538501
zdb3295cc3908bdbce60b1b73922acc06551e21eca39da6028649acfd3f5f3f532bd374e6f5da87
z10a789c2ccfbcdd79567d011494b2c91be5d8f6ee7817d05e58ee3be13a364269bbe8c46a0b0ad
zbd2f8990e0ead8cc658f1a053436ab67924f6f9545d0872494be87fbc27bca30053292e5720ca1
zb8ac77c051506cee4a20519502cbccebd390080cc70fc1f03034ec4e0a32579a61f327aacfdf97
zd539757b1d4a542ac2cf194dff7612dacf8db8a3d86fd98f08347d1a6877ca55019ab6ae031a1e
ze4c14b4434b12f68c0f0832106acd5193eadf3485271eaa936afd4043713a0cd1da1ac53755f52
z75b0ccec1416848db639b45bb3f60d96add5c37eea3c53d57c2843571378b8bbb840aad4ecfc9c
z73c0936be0423afd814ac3b7cf23f4576764d5cfe475d5d80d67f382395cfcbe1459c2a920955c
z03d09d7aea062ff9d060c98715783391bfce20b35d6298f319dd4ef8f9e4f5bc9feb123d0a42cf
z82fe870429719fa18b215cbed1f772ed2462180291b270a30dae3ee0370ef5a899f569e9d9f858
z430d7d5823a3a7cd28a78c9ca536b2e1caeab0b1f2b3407d2c6dd239e5bf25acfa68f7f3e090df
z01c947ad28604174553665a7b183f98fedce23b1a1a7de75cf961750de4f152453067c23244795
z7600b46afaf321af3ac55a047d6e091b4935a427cc5d73113c62871fe26ae39e0002599a1dcba2
z4c8b5599e5afacb3f036f183cdf85a43e508a6b906da138c0ed8c108bcd4e92b436f184577dfa5
z6087e5659d5f1734c2ac6edbb381f9c584d4a398920968b0e37cc31f0174d5ff6faa6035e18b43
z84e4de0007ea643a16cd36d86238bca852467ba99025704dd7144b2cc51a1053a96199f848b76d
z783c1ba28f9f2edf40590e601abcf7bed72f156fc5ff4a864b9d768c8daf6eeabddd8d8db729f2
z9f84eb1d734d64cbefb4049c645567182d3519a0f489c2a5b79d6818dd67ffb6eaaac2a6fe09ae
z4b6f076c57014bdca2370faed3df28409efd3a5f0e21a8a9a3ce5845965bb97c4ca883c548f40d
z9c9dc270ccd93501855b0b7bd1452d4870877c98f1d88a6894eb95c8cfb7e80ae44792649a01e2
z87c8377b3c9ce8451c57e0eb33ac96d3b39a1c5a1af86533aadc3743d5dd5ccd13e640371c8867
z754bd4d16d5eefe00fee66c530a61468ca60b38ede6738ed8446575570d054dff152607f1ca9e6
z5410ce588906ad4b62ccc959a26872616a0b9b302243185b8af67cc4e18f0591058050980c64f3
z55ea2850b6283107f09da164884388d4d930f24626b0dc9426b2b8173a86e186fbd9ff1e4f3f3f
zdd6d30b4a1ff31b7e9b02215884bb7dd894a88a6823ce79a9927c826a16a05e38484d00a1b669b
zb58381caf62030f4fbcb23eb6e4756d9bf9e8f453231f3b3f6dc8b3e6dea1f8b34cc533d7c54d5
z1d8ba2412761c4f6bd747f875c8576f6343993f77c6f1bb8d7b23cb700da6e575d2024674be4bb
z2b4a3e18abbe6dce609a4811e6969663007e2ab672f3da89ad0b824a17c9a92bd687576227189c
z53805baa15a558666f1831bb34d044635bdbf34db04bbe04c3686fe17a6fe51324a4102b8b51d0
z258fd464029ed4fce995796b2488fa7e9d08b0116c1a91c91a91e22040c3da4f38ea69b5f0814f
z657f46af000c325e4cb960509e2d585209f3e174ad69d97f994cf3b2ec9a3e533ec89e836e0238
z14990ad69fb56518d2ce4e0ff14e9179f6d7647dea15fe0c0d1c28006512ddd867fb313d61fd2a
z2e53e6dfd00fd21db231d94a6800ba30bd70e7d10bdb8a071b1d0d9d08a40d36bc86c9611d67e0
z53e8a2783c125411e2f62f2e8679d9631f922d361c2930529a23111534b1bf493ed2ac043aa507
z5c23719f422307bb6a508655cb15772ffffed6c703a37304a858ff2161ce479c485df61b7b8fec
zfd6c806876ee88ba40d4ac56acc36dbaf3edd80d4f3156a59d8b204be6d2846d0a78ecdf692c72
z48f616048363987c923c8d86452074ae1e44c2d15ed0ada7fe2678bdb6f950f27b9f18db73e445
z0743b6167a4c34cc9a77b1ce1036e52d71bc3b7ea77ea60802770874b37f0ee74cff2712dec282
z1f16c846b46869b771265764c468eb32c60f7cd3afdb5788129c50fafd592d0d92348f60a8c201
zdbd109c3d39b539ba49eda59d0778f341a94353981af8ed671027e10b22c8b30568e817b8aba85
z0f8a59a89e7e7608feedb920cf18e5e66b824f8b65ba58ed467fa9570443e3f59daa5a217d6dfa
ze55d8d437e07ffd9b572f3c8ae90724fa5a2301f54b3842dfa13f87ed67d143dbeb5d6801e6282
zf8e79f3393cca29d039a8515d472efece3a06bbb61e364de0f1dd2d5262925c8df8c9e13da3526
z48579acbcc5a0673ae04490cbd8c413d5cc98a338c2325f2521806a99f379c18d9d38d22d8d736
zfade079861b47d67b7324ed931e1f644c7ddbd651087b0ec6921c41eec006357af27837886fb50
z0955dafed51bc39c0237bf3ad9e54f79ed76b52c2600e8f3b6d53046cb5c0df96de682536754c8
z64c24ca9b86cf5e7b9db804e222b1b040536d4349eff89e903841e172cd6c58aa38d844da791e8
z73dfe45acab95a57d3ab75c1ccdbc356fb4f5256f0952cfa51323645f33c81f9aaaaae2c9ca5c5
zac6b76b55f153d9eadcf1d290368c4f9114d0117df81d82f91ae23d56f341e9ec9c2d53770296d
z329f4dcdee1056a51e1cc65687f0d10b0a5dbee9b020133c34d95f5a119472d7377aabbdc60a1b
ze5b07535b6f679b84cfca48dc00f6bdaa4cf496e9ed470317d885b8e3e05003d51f78d2397d5e0
z3ca1da220c719aa6b0d981aa3731bda481a7a2e43cb6d0d6a0e27576a600ab6fe41cf69b58e55a
z76139a24c654ac4995ae93a859bbc75b24cda20b597bcc53220944ba2dd2b8aa4be0ad221b04bd
z29a316076110a52eb8ff0e2a9b8298eba142809f718156d665eb4e635ba0e999f6ff94aa552bc2
ze0425e046d6b244281966a105f9d5998f1a8a43da51a627343d3a5cd18b889370975bfa2c6362e
zcf0651b0453f9a362ca56179fd7c42e01b1686eb0bdb8e57bbdc6ae5445e401495408156498fda
z63872a03c7fc56a4692d4cda2c22aa6d27e41b40f45fb18a0adbf77ec635eb735cef58ed043886
zcc59aaa30bdcc5473be81aa97b0badbf27229aa9b1d62d095b1462497ab455eb4484c72c72093c
z4837b8e1190ebe091267370699819c74ab47cc4616319305232eea0248cefcc3e5a0afcf540144
z688d02987b96d686e9c24ff7ed4e42ebb7f37184c7e1483351d196f56a1323b2c40fc3ac27a100
z0fe94dd9d961bf1cc52a2f4c2848c6f4582db5a98f0ce098b92d826a02b8147038fb5ad62d1676
z49ead32c9ec80a11fb494190ade20c4d43e39477a6aee8942890a06add5f652a2d90ef135215b2
z405c79f9f94ff01afadde71b6c0e3dd6d3667f714869efd5301530001d9a35384f4aabb2ad9803
zeab5841d0a654ceb75d7f94eaf3cc8f4f1785df685a908856ad44ddfe52c9d1c4c012b10e84ab5
za941c9f4de608276bbeb9c17bc017951a3842ba2bf7311ba98fe56154b01d8e3db8c6c979550e4
ze47d240b84c66bd8a99dd07501cf47afbd087f11384eb21813733069326fce78e9b2b4cab1453f
zedb878464e96527f7bb9e1eb6589366cbe49679068b34223b5df0617a870ebfd355118be261ff2
z74e1c3ba9695244cb6a77ec930435ac362d22020df385a63f795d427a35b5d7aa3c49d4edc7400
z51bdd90861186b5349b0e754f80b13de682b3b0f45b2c849355fc8916b6801bcb966815d2b1e13
zb0c79b73df280e703013feb6d5d79de51cb0558aa441db4b260e3a3c9085a41044f98a08694f9f
zb8ccbd341eb0977c973b224b583237474fcb91704c3599db3edf5a685361196557824046b83a8b
z71fb2192838d795b5b8833e9b8b40d1a68933bb28d41c44943b62f37be3bd1e072f46c8ba04745
z93bde6e528a4e6590b9f0b1e9147138bd1a3edd05e5a13d468deff424d4f928ca385f367f83b50
zf0f40e1a65af2ed808a7cae9b2312ccbba5bf2a8c1af716bc6aa184f9064f058fe8317dd1fd1b4
z193f39c260d685b5396551ed27e34cf300b0a9ef04ca53500d127a72662f53e1082b710d004b1a
z1306fc381c6116551fb8220d67ed063642d0226cda5f07004f2a800859c3dfb9e54e51e9f21117
z994314b5e579459de80a89ecb2754d3ad084fddae8da0931675417403ab01d65df9d307a865921
z4afce4040fc6dcf9d75cf7b0ed8208ed1e2ed33cd92b8059e83dbfb13dadca4cfee1558bdc70da
zf90f0239157423cb55f74b896f688b80543eb7ca771aa2119040d8c6fb4bdb80d2d06c66eb6310
z44d39b82ab4058faa0f87eca8e882f4272c40b6941ebe4f995d9ff092f15ed87aa60ed414a6571
zc5f35ff6d6fafee9f631af2c4679fd5dcc8e97b9617a9c97d7c391d61cb17c43623e58c1fff92f
zde44b967c87154e8a786f5842981a9b69ee43b0fe2d048a035d25267e967586ddfeb29204c13bc
zebae45c90f269af83d08344b1ffbf2cfecd3711c89cf4ba417397d41c37579625e927ca90c447b
z2972917229f4099773bc0c91203b515091146a6f31525229ee79145c0f664e3f2460f9b443388c
zd7cc1c5f50e2d48562799ef77d0cfee530262c269213fb5be7a525a284da9ef81bd0e891c99a67
z8b774742c05d6657af7f764bd61a653efbefba7a475cb453b2ec9fc0740d09972e1c7a15de05c8
z074ee87923b2491c25c2802d0055bb9d1d2de5660cfbb4f8c75841ff0bf09edc7e2cfbf9a222ab
z9da6e9ae0d6c40ed8faf80435b4a5067246ea1bb3975ea1e3d240be6a84f2d491bf99e4bc399f4
z58bad80aebe5a500dd6762770b49ad2627f7957a764d2ea53b8d025259962c7a2e12b22e7eb2d0
z64f97597dbdaf086a9dc83ad6290dbcc843ef6bffea8b72dcfb0eba85d19beeef7b4770a65676e
za4eb29c093a1113f05b3096090341b704bcd0a6c210c301538eb318aa0c9c1ad65596da017a07b
z1d0fd5b69c4e4ce55b4653e920d22957def2b6218e4bd6126a66b915687f1bcdf5ea567d4485b5
z41c4f3b8038852e1ee0b84e727569b24ca16a93948a47394cf736fb0e8011bac8cdb54e9077bd9
z04c372f145a938c5ced1335a84040557fc309193bacc17467e5fce931598e75974a33235ca950d
zb8ecec1f136c5febe4451c2252b1611589ba9bca59b03b0c9b83e7f1357d9d1d93cf581cbd6b15
zb727e982fcf7eb885a8aae3e521111d17ac8e3d3ccb02cce4a2edb6f6d310f773d830ec69e292c
z3ee74d5a5933d67db2e324d627eda7f0894623bdab79c8fc3159145aa4390fef0dedad3c9fba2c
zeb5ec2798f0bba2fac4c68cb8e41f661c1bb9ae3c7a9ab2bce7c6b3a3c4ff286ac7e643684b434
z57d8c1cc5670c218ed1064dfd7ec134ffbfb44377babe779fda4870fdd265148b6a2fcf9e0ca85
z6ad7b13f699540b5c80c892706dfbf7d5997ac1da95a6e51c7f59733992e6f8352ffbc362a7534
zc2187b866c3c1dd55951ee8c0d5d04896ec8c5c7b25ebd7d6da71665e9d0209a4241b2568d13c9
zac4b5043e3dc172149b952b382f01d497ea0ca66172ffb22b3da0522f559b9c36f92c13cda3946
z11a27c2eba0ce7ec55ad3d718f76ef11d91ca64f7f4ce736f780f0cc4a47498e5552113231794d
z7d792e341019ac9f83f0ddf9df524f0932f698616579fbc7f48263d1b9d685d6457c15be4da447
ze35a7403287830bdec5a26918be1830a249255e9cf40c230cf33e6889a04593da3027603a99a7a
zd34eda70945fe84e72536506a1578f60c713f274482b092af2a107aca99db1cbc239f3a6b5e539
ze9767799b90c4edc2d3e911eedcc1b559c29156fd7b516f5a75cf225bb7d4485e60dac780cb49c
zc17d593a2afb502d7066ce96971abed3d7378db3630713e0a21a427363fa12a0a4e202a9a77852
zd248c278531733528b74a63a2d0fd8e269895b16c02067150c98bcc80979fdbfd799f492c07f1c
za23c42b90cbb961119dc6e7af66b5ceb46e4903945795e31cfb3a383be70a13437c2578eaf23d7
z9852bf8db26a616fe1a11061a1381ce63fb41ba632cede186bdfc66a2b041e089436869d30abf7
zdf71ba015f3c1a9c57ba68a2048e1f52b9c023eb0f721ea3b16b42c99aec4793304d38489f1d03
zb453d56f0f91bc1b6c8d99894cefd4a88bf81825280e3842f4d850f1bb3def0573d98d5dc9d0f7
za11d24c5bc0985017f8ba250d834b14aa4ec1915488146dbc55775dc1fb4c1b1eabdc021797099
zbd82562cb686e206fc5bd6baab3f14add1e68539db5453ec4bf73914ae7ff950f917553029a6fc
z32ed347be57e1ecf1e374692634033c280412342fd453b1f2feb71e337d341b59ec2ad15da619f
z9a7e0f657426f560ea23e4d034feecd371b4b95aa43e1a4f14c9ec44d6e1b8f2d51ac5cc668320
z7ee72552fec4d7046c79d92055bf9d3f65b72a72ed19fad1c52dee0b031cdce627c8194fbf5bc7
z660abd00d10640dfb60d08dc2d54a7627f5cdff65e61a01b04bd415e0cf3a8cee0cf187f4bfefc
z59d48d039cee73cb70a3aec9b902f50f98c5943f3a4fbc8ee3554f06047b4441b1a356ef9da8d1
zda3a48cb94cc6c602f84f4b78a6ed768f026cefd3654975c44b52e3832419fdd7585d835602ba4
z718b085b92c8861fd654ef2674a90b0fc8e2c98bc01fe048d0eccd87a67f9339f406f125d2c968
zf6f9d97002447c7e0071686d3ed2ff29bae208ec30abdd4b16f3b6fd16e6e11a5187485d7e1c4e
zceb277c663ac4d943d2668b99278236f579f36f53b34be8dd044e8640c982d92e869349157bfed
z4533a1c3414728bacb9fc7a113cc3a206f10bfc64cc9f0fbca47628fcf0efb09aae3fc0aa8198e
zae2cd16c17aa9ff5f5ac9c8b8da628643100dbb08a7660c2306e463fa2d54e4ee4d4286a2739ca
z5227cf152b33a65a358bc5a7b0ab924e3c6553ed4a5d0eb3b4868941999bfe57585e079f117ecf
z014c60f6f41f9648e9cd12c8916042d4a0a3b68f42f0daa8d20d05fe003f86239fe429ff405b3c
z212a2c653d5dfbe66a7052ce120e0591c417069668256f3d98dbb7e9b3572fa3c08fe4da7c5615
z645ffdf8f2f37e836837980799953abca4cd6c781d46f001d800f9a169636fa4591e55fa6fdc59
zc4c53bad5fe6fb3d4c3b33f2feda0389dc419f0ad7f98e24e4fa1b983418736037ae32f76251c7
zeaeb8a5d88ccbee872f7dbbbc26af07306ddaf8b7872ea624a34d991ec292a78ec7adff2d6613e
z2ab8c14c795b801150f982dc73ff16c5e19f127ebe7148f6c3406a89ce4a19afb344e620daa8e4
z112134e4877359bf121a619b680cc05f51164e5bad5a9681cc349b92f5cf2139708869b3c3b878
zeb91acf3f7c3ceeae7404516a0071aa44ed3622735b57fa36cb3a610c4d6734f0170b774277bc7
z9cbb564717e5df68ae9dbcca788340923a2560e3d7a3ab65c275cb67571fb769c67ffb1b2d8f89
z775b9d7903e76f6d6e879e0fd67a0f6fc4ab33bce44f8d5bc6ee4272f14be5d177e782fc8c1700
zca270260e877b16c83590b2332a89c47cbd0b4219bd4dc956b2cf6ef423a0ab80ac32b0ba681c1
zdfc8d822cee6b628b0b108428eb25b0ce3fd21f37281bf5ad6bd419794351d7ab7357c3510ce11
zc0c0e376306061d54f00df66165c0d8fdfc8f9652c2c19683c9725aa9642931ef035fefabe8c17
z47f1585a8fb2a1e13fbe07b953f0187ffa04f6acbdbb001cc5c1df10c3675b39048c6ee9f52aea
z4b9f3b9455774c9b7ec1bb5414f64590df4bb3707d5f004844e8dedcfc15adaca5c7359c718abb
z738b5137fbc1043c0037b03ae0c6190bfea514edca58c0c8c94e60eb7c7215fda15d1231fff5bc
z61d92fd82c0ec8b04311c2fd974b270597ed4224fd5160c289ba97c8bf833ef332e33a63d9ec76
zddf71766dc6c08a3082600e68a736320a21a0dc096b33200a9b4bd3c01881526151663b56342c1
zc51333c4f41dc2c908ea95a1569977290af9478996918326b191e80979fbe28c0c8350fdd3eb8c
z2c7115ce7ac1220629cb8a6fa6f7eab70c36951d71b7d1666e321cbb11adb20c1579c6f6425e11
z3184bbbf147ebcd6dce7d887929bf02492149df1403ca3edf1e1f457a7efa1db27818878b518a7
z34ad925616ff1e0b039a0361c7fb3a16dadad300c96007eaea9ec22a1749d252ae0f50cb27ac33
z60fd02f72c3219a93abb8ed74cb58d6d4169e591aa9939c54e320117ab7e2fc5809eee234a8c47
z83fad0af91df2dd27aaba8c79d5616fe31083322e764d0aaa9a4afab4ce5d7c9c8b72352182b68
z827f773a6e234cd311abecc52118da6b7f30fa00f15c3f2ed85896cfa83d504649e6ccc1a6a2f9
z05e487f538ed76b97cb7bdcc6d7671a6f88fe4a93cb83a74305c2b88a52f53a5f365c3e76e98e9
zef47f24faba2f71f13d4b21fc29c5e687c97a09d6e52869f339f4d31aa8b371dc9a1cd24f2135b
z3dd2c7dfb65c4eb113f098d46c04594e93034798e0398539eff0efb7f970b4ee01c24443eb59b1
z990b3ede0392b44d891713f580bdd2b142f8916a22af0b705145e78fcc996f789e8a36d6d809b7
zc9ee0e58fa4cc7ac4e859c90ed0923c7736896520f13ca02f7589e918cce8a59f7262f38023347
z7e6d2625fae384271fe072a0fbcf99ddfbd4635fc81a9bda05fec514258e3fa74a691f7cb3c834
z1e30b910495030d215fb879f54de0c59de2330c09646b41c2e868a7708c26b15eb52ea5ef038d6
z05d5decb3e09a40beca1b7c601971bba4004ee52ecb5823f91371dfad6b822132b65222e03712b
z5053a6c24209cce3e3afd04dde8ce4738315a8e1f555798f67cd413e5d93a79cda55c4cfadc5ce
z79e5a1d53c5bd7a90bc2c8510e817e41c8d38cc40c75e53835655cddb84c6c8a6ce83b1084e46d
za4270e4599d67c774f027644cf8fe919a41b1555d6873956e98707f261787bffae85b3e9d7c64e
zb74e3becb0153fef15c0fb25efa1a1a683c8bee5859f2235af2ed4d8ec3ad0c8c3c6c4437bd4ae
zf82ef23b275525a5bf3589a7f7240ff5c8e705674252ab57416a5656fba4443b7b04e726541324
z8e13b45ed4db34e44e20807b521627c0f02febd2a0e6a0f47efe0e63cfb412c3249925c1b6a880
zd165d94e6e2d1a826bd9bfe85882f315fcd9cae5ac5248cd0d07434c0f0f6193cab62b2bd544b6
zb32e3018f22b8c504056fd06ecfc119a00e9210069c67c30cc2dfb47c081784aa622804d226f84
z2f1d100fc5349424315aefbd0c923c2b93c2955571710d37de0a8afa2f0089638d81ad34eaf84b
zb5e5308e8f3c173e9851c189fbf085ab516b11511011e41aad35b67df41ffa456ba601f593e410
z97350bfd4658ed0dc9e0bf7c1249bd3469758a6ed01585d48ce352adf14760c78199dd471eb20f
z26ddfad52f9f2f56b6b488409f5703408df49cc9fdfa87a9a3126a3c8460628aadbcf02c3d4b8e
zbe7da7aba9b6804866ac21abe10094e8c31327d4adb62b3987c815300ce8af8f65d15a73a82eb3
z5fade19f05a47687701e519a5494b1d9f0aa9109561fd045f2e2191941c5b9023b7353e2c787a2
z6aba8367fa158f5717af17d3f96ebb0843b8e882d5f7f23aa93e207f28fedcc937ac1c8336dec6
z7bf091fa6386097f44ef63e533ade9ccb649d9c3546bc313707a649467907e1f52f283aa16ced7
zc55b0b111d426eff23d097bf7073666c10381de81c436234cbb62f356f51ed1f181c7dd8678824
zd0538bdf9211d75986cb53dd888fa7c1fa3b9291bab5cb26c26968c9ec6a156763138cf8174b37
zb4ed3f63270d093758fbccada7c18e7bc550c2a89464d9a88d51f795e84186ab553651aa57d4af
z7d4a19a3ef26e37425d74fa61a18b260f2317ef517842d956a0d4304cf04bc4790d52731b09801
zfd9fbb5cb30a57695af6497d5350393eaa4ea77161da42e839923e1bf7c086d8fd47fb76a7e254
zdb16d404edb8ec8bf7ef7f6f2e5eac512deed0ec4ea3f9b5cc3c3e1a98b2e21c638edf09fb8242
z0f47f42582a00d2f7234a9bfdc1b84b6f832fd25374764ff45f6bc5e9d065804692c1bd52be569
zfc897219922daf620bf060d7ef198e6677b1acbb77de8891f473e04cca61cc7ebcd0dec352e8fa
z39f915b5eda5a610d2617f1eedccdac909c68745e88e4a7044d24ac90d9601f92a51690469af57
zfb9f6f7d6f83c57d258e158b7b2441868f86152d294b1a88c5a04730ae6faa5b9cae46a3f021ba
zf88d2e38e68ddf9f3250fed32f2b0cd9685169bb376c0eb9d38ebd2f259af499f9dab4047fb181
zebaf7a805128b44ac4cee12912fea359c40886b4e601535fc55f9ac87b6ec720cee0de49c9f5fc
z835ff70992810b4bed262e9eaa07ebbf12023ed118c2a12e7a3a37172ecbfa2aaab9d03d57aba6
z2bf93da1ee8adca265892fff722197e55d0212cb1b2cb7f0f66bacd4ff3a47758982ee60ebe37d
z57117c2ac75633a1cebc9d5ba4d6a8489ba4a1c9120239f271c220a157a772b757fe434d5118a7
zc9d863233bf1a59c46de955761da19c8934287207d8b9da4b56e12efd62dd62a6e783f403b10f5
zb66da0880b08947a1c91b528a53efcfd32620b2df82c8115ca26ee13a49d4d3094a23fce6c98c5
z9d30bdd8d055e8fa6ce106dc08f0b72777fb98ed3d8f805c05d7acea9269024ada6590374241d9
z795b4b8d0e63984c122db8af1f8eb06a35889dd45e5f24e52cbb4e905229b2aba91c5b52c23039
z5570dd5ce2dfd74bfad022c2bfdd68fa7087d655079330c23dd3e650d1215af252a21b3e3fd913
zd9b6c0e21e1b3b48271c3374bd9735136d5685081f182d04df72867ecc96dc1ddab1e8ff606535
zb70544d5b6be5d2c5f2d81fd7088a1198118fd0e29ccce171bb6b8361d51428f5246542c6894b6
zb690b9004ec6b96945478808a0b3e4ca65fc6454c77ee17186f95c6607d3babdccb227c621bb7f
z7f95feed64f9d7513a354c4ec784ec66da400f41d69f0bbc02cfceb5aa8cb169339524f88a3125
z1af16c02dadac072452286c8e811299629018db2ee0a720b5ec6542183e48978e364b2be5ebd35
z656ed48f6d00e6078926b9b705b248b226c73976644939892e52aecd761a951637ec8bac0d831c
zd78b5bbe11b713d3e4b5212b8dff344101432c61d442a780af70b1d1fa60c81c18471bab9e460a
zaaa00a80555d62c040fa82e2f6c30b829e0337288d464d0406b43cef4b9902edc9d9d7c2bc102d
z730fc6e9e1a2d14d2445618794038f46d8bfaddeae0331ebde43e6d7cd9b82afc4da9c164983e0
z06d41d458181b34881630ea6e784c3a78858ba6d3d0df1e2ef863005fcc7f6e1401dc43adbece4
z4671a955f1bca54734782a130060b44e17814188e4d6c2b1c656bc0cef00533b6fb04d2cbaf332
z9d33ee209f88ac7a9b96bac7358cd4bdc700c6af7d30c615bcc90e2488cd09dfc397ca045223a1
z9e85c80ba28a4df632f78fbcc4ca197a78d6728ce0990d0c4defb5d5657edfeb81fed5fc6c8924
zc1d247a81dbcb9998dff0c89e62acb0ae8c866860d4fb87561fa3caf814d642d624cb3833f94e0
z1192fe4ac1085542abe061c62e2f0681a0f5ada8f145521a26eee3ee98bf631f1c8df6887f85d0
z23853843246efce34d862f63bceb23a245b51dc1a51fa85578710b8b528af952f7e494e2bf57d6
zce3beb0e652944b7db249ddfef3952fe01a2692d85e60d4ead6c39a6eebf19b09e552acaa3037d
z25baa930cf87d8a4d741ca7a12b82e6dee3af6683d32789ddf35f6d6f0e64646f44714f2c03bf0
z6aa08f8217639339c7fc01812c51d119aaad46acba416fb0f892b0344836f8b2495b0e78261247
z17eabe381485da7b6bc445d322aa72b05ca047d41483bcceeb0ec96e08dddb59660315f35f63bc
zec6b8b190053fa7e52b70b599cb749bc98523f8f83047140df477ecb0788d3d771862869fc71b8
z028085cada1c30c2c23a137824fbbf69567f0f1ee0d2e61114c3348002396f8c3ef9aa5c33ea40
z75d209e58b4c74fc0f76e1181e16986ac77a7947807d4f4de22c083ad12ba8ff79d413e27d8131
zbd8d894679b4972f8f2ce37a0ae78cd0f8585629cf76e594a340ae6ec9d0e7caeabbee3e18089d
z3c09e4e16fcaf7d7be7dbd167883bd5d3fc89b96c60fa2b9a17d8f9ce3ac1ac30abf80df1034c7
zed2be2bc9c58fc46b24d4afe7701a543d3942b786e828af26ad985bf3c899c78870a6485feaa14
z840b4cbb93946d14c6d5fd488a7ac10006fb4f9e0fdcb22c0196ff48b44d51164e70d2930ea12c
z57690d918bb7983a9b0f9be2dd1dc29f54ab6bd3183554eecd43ef00957560d0a7854cc0655569
z6f2382fbd5a8f33d04644dc69b03e79495bf96f934a32a16fb8c61acabcbb8eec6831286c0c07c
za1c7722e3a09f62c952892e44a69521bb53e5742f984b0d688bc098c4bb3a25a1a199a960cc449
zec6e526b3f2eeef23eab202093e51729b78ad7c52d0c043488acc9cd512ad3854615c815ed9347
zba94adc4dbcac49ee6863f2c3b79f19f9c3e2927171e0241c61d1f2e2d7f9ba31c5f0d460e6147
z771a556169360360dbb47b4320284cb1d510ccabac7691402d366dd0ebe5c90a2050b2a84af6e9
zad0cbaf0b4258edfd17d48f8f2f3102d93f964eb566e2cb2666e9566a97c9b3ef94e686a9443a2
z046dce12eb586b05b0921c8b0ab491fcf7b5d59e40ae50a487dcd247d0c0f7b005167a047df401
z87b2b547c08da8c331077c1ff8fe1b86e08a6b72df36c0ebab5828a8448615735ff7bc7c65044c
z8a08c5d9d027a7d4f61b9654ee255d00f52ec54de527fdbe81ed16824b806aff4bc48ee82bf004
z4e32a7aeacd9529249e4fa01efb0bd9ceacef90dcc8b503d238e868bd9c29d46a429bc675fa529
z3eb2c980c17bfc9c2af45160f94ac74a08f729caaa5259086c75e6f2d34432bd442a82b628ceae
z1e2534a08d946479d8c0647fe7b006c5a26efb9c8b3948c8f517eebcc4bac35ffe98d5f1b95b9e
zf61b3c4bf8a787afdacfab138cf105618d4e78b987ccfd1a17396d9ec02f2857b6f9cdf5a90a8b
z7c849750b04fe7a464ae27a82a60aa41af6eac6c70c7146f9ff40bf65a02af8bc441dc35f0e64f
zf063ecb1681ddf72511b2e1250768568ff8c90247eddbc778834318b0ea5513d6863cb8523550a
zabd38132da1f20ccc849fd2238c99c3e13fdd4b1b2dd4b21a8b157386ab60d2c501bec92f36a3e
zb76916806957fdc54bb5d9de8cc4eff5428cded851d46272b9507f80a7261f1ee523f860050406
z31d3e040d692b370c5f5bd076450b599d56e37886ca32134cce591625cfd14b9289664828da9cc
z311a87ef147a91cb4310a81301d1b601093f58a8b92578525f18ee332120e4de3a250c33543367
zbe97471e6d9eb7b796018c409011f27ea6ccc1ea09e109511b8cb7ff965400c8f93a70f6c57093
z08d9eca0fb938577a7c698b18482e3620d7bc34ec5272e917ee04df3ba1d3ce37f40b602eb52b8
z88854f277d6f0934c7626660790f9e838d33d1bd3802e6da183578a389ea9fc790a63a3f68a6e0
z9bd14f64f3bfae77fee02f9328bf12d86d9bbeb227648251bdd22138a7e55a85979b8a14b00fa7
z4af49197299a62a16f9e7f3ff1c2d6e8a6171c002d5c35ec4f3126a67b5bc5ff0c50d069059da5
z3fe8847803448007e3663911b4f5f3a0b59bbcbb084dd7b88e93346cf2743851f399c21460cc01
z9c08ec32baa78b309bfe1c4e5643a15128443d808a42dc19c486bf839721b300453afa90412532
z73bd61fea0e88de57321bc48e9df0bce57271d971a48fa21c2ece9702faf26032fb99e0eeeb405
z10c87d3d3b47931fdd4487fe22d4eb1d9fedb97415fe2a92d4f473d2d1f9b2053e7dfe29203ced
zd94befe70c6d01e9830fdd9a2d637d2e10028bcb487f42288a17895ac0bc24d349b3e6ee0f063a
z4e6a86e17fc45f6807b087f3149697e1c94b7136f03830e63f796f5463360477147e240de6c9d2
ze3bda0619bc2fc0b7aacc8904761538621e7c0c37d44fa2d1e10e3b541dac4743b48fa065c1249
z06eab75dff0ed8f1fecc163b8ca7cd7bae2ab6a2ed87b7710e3e4eea7523f73ec4c6e7cbc48dab
zf1a023f19a0698f0d837068413f7bf9c71774393adbfbcdc30be7427699c0180ad0d2e044834e6
zc1892fbaaf123d0befb1e1fc79e3acfbb452335a97aefa284a26715fd4ceae7041ddf7dbd390ef
zbd6fca666b9dad1ac6a5b491d5b225da94e5dba9760c773853947c1f3b6a9f370e77dec46e8709
zbcadf1f576d2081a5f987127e28c80cec5152092c1a8d66c291433f5ffc6f01bed9a5f76bc259a
ze6dee17e9460ed33808e246ab041b0cffffb29de1878ef1c5d7d27bd2944c0625f727df64bba9c
z9cb5b6e93267f29f2957a1cc92a7a7684a96429a03899d4f03a8a3af5bf86f9c8264eab88f485c
z84630b6e9b5dc3cae451e7ac964e8a88ac108058e01c75372d84ed3ffa3e741789e0bca5dae335
z59e146fb39dc3abf3117b2453845a66a51c0f09a9cd419c2cc4f2e17271fb39e7cb576b54376b1
zd5fc5fbb78bb45bc1ef88e7b14d01daf3048658729bfb2fb336c946a7b588722205b6aa272afa3
z690fb87b00f6ea215adf807e21b1def893b87a3bd7c5521a248a05e0a1eb9459390ce82b7daf18
zb84b26ea766c4eed6896f54fb287e9b440eb2086d531f399d8f26e04a4b609af47ec28a1fc1030
z98490a9710f9516c9467930e7a1d4640f38b4c891b6e93dc0e520e94cfa70975beda93f13eba89
z4470adf9a53840d18b9ec61c56d91e7fcd1e880165effa30dbd73bb90f340ee22ae281e216bb81
zb330e0286d60e66e7ef0703ae8af065c78853054ebf8d9c52184264b5ba58e15ce71e66ccf8a19
zc9678102b518cc9c23e6cd545274bb9fc0a3fca414b0c2b105075102080bf24ef7ea9082bddb96
z22fab09f1a37e3f9d99e6506490e06e8cd04ee4065532f912a29a916172035ef02fde1dafe9fca
z9db157f7c7ea1931903574982c9a0ec04c2d10d8091c29660c4786414dada6e08c0b693d7f17bf
z32185ba3ee9f7a3f921aec2a28bdb4d85e29e2053c5b03a8c2bcc6bcbc03785b2d081f7838464a
z106986b5116ef67963d1bc993ff8e8c3311a16dae1118557a155be0ee1ef215ef5e34ead6e1a21
z7a51c3c342d23ec00a9e7c34f117aefa010f2a45a4870c855745f823ef5d1b4b7d71de8cb887fb
z00c82ee5756e13b359e59768c501d1bd4b4315e9e91e804081d2a273d7e5dd726b1be4c8b38b54
za0b8a644ed2e89e552f76e0d0c74e032a1f6c97568ab0f96849dccd61d0f4ca75ce08b55193943
zdff636516e288c682e1adf1b7810af9165766135ca22f9d82f241a86a24a35d7d60fda95e223d4
za04e56e01bb700f6f0366f6ae4e61ba58daaa714007b8dd8eff1f1eea59311e09269dbb6c9d8c4
zbcf1d62e777c6d7d58e002cb84aae988b01be44a81077570be225336239b02737cab8122c7ecb9
z6aea75a5b2fe00fb7cbd8c47671cf5797d9c26d94e7f8dc5e45cf692e2a08ed784b815255034ab
zd059be74a1c7362f6062aabb92e4dbd9ddbfa65bfae0bb6252f7b060361a0bb36249da6d441131
z8723b613bfed71e31836aebcba3da2b17a3786ba9b1f50647ef56eff045d4ad5bc7fc3e4f6e356
z82aeb42be6c34dbba3f7d52208d5f9cb33763d617924b4abcfdccb776a07a669221463b12bdccb
z90943666e5f841772e671c31301a4fbeff0fa990ebd8dd3ae1f950e11174fb374f2fcc8a098ba5
z0476a369a5382d12ac7130f475a645e252064cee7e46e9f3898f557f9a7b05048561f68f0c1ef8
z6b26f7c3c62c15b15776b1d84787347f3739d4d5bfea779aed816f2a372b794da3e7e1d39a4bdf
zc618d2c108e769e942e13912bc93b656b3a2d89f832e0eeadd2bfcda09a6804bd52fe495a792ff
zf5f4f2bbb0dbf5af89fd1d55f9cadd063adbe2038dd532eb08199e9e5478d6f22da5e5a0136323
zc4506e0f8b8b773232969b0024eafcf5c09f7eca7ccb3668a9039ef10cbf8b0d04ee7b689e5baf
z840a79c7316548f229f36f71ce65b593d41c5f9454fa751a4837288aaf8b18408c12944cd5fe16
z06f6a6e0e6d2a3bd38ec73442859c052f492ce8f9f328c3df0bcbe1c91b86c2e6c62176d5cef93
zeb8a0a180e3ff8a557178c6ff18596dcfc0e4bce68666005ed6fc5ac633f5c7ce734bf87620b5f
z8c34ce211482a2eb478ceba3df4862b1e91d8bfdd1f4fdc02230ab1200b644e0a36986608466bf
ze72f24daa25d8164e7d6cf4334c0442a55d242c8c5fce628c6786c9c13cca96ac05d962561a669
zd176e723e0b77724c33cc602a6bbef218ce2051d70a9bda768cc58750eb152dd1f53b2cfded0ff
zb524d6e41ecae097cf434df7ede05b0c3a136a658c01b539a4deafe3708558332a4a6de7a44604
z56b8449cab3fca0841c2f88f3557f0889403ce85a466a52bf6bacaedb30063e944b9a60dc5c27e
z686899ef369f4fdaa2e5b5fb79ea35dba059886f8e07f7d535f9de84210fd37910d7a35b6de970
ze9de03cb56e4fd963c96f90b8fb46241911b2d67bb4e39b9fe666ced6c9049bc6b12d8e5c8affe
zdfcaefdd1f81a77666a80d28b93647fe6c66bc0c2fa7e1768e7c4441ebce75657b23171e0550e6
z53a1de6f0e7180807b7732442ae7a15446b6e048f2b6bf50ccb6b941a33f3dcf4819aff719399a
za6f4da9741458d0e1caf13096cf298f7a5e3f0d238d4c1593980f08932508bb94c329ba23cc012
z84eed2a7e1fbb36382ac3381ac04bb81991957803d00da3800c301dd9631e1804a9b7577439f9e
z9a272365500259d8035dd1c1c808bbad29920e6773c94c398e3d66c55f08aafd47fcc302d3c728
zac75d3c8c143f39f58a5674fc5417a373fcfa4e119e33a41dffe669a239bbfa5428cd6f89a365c
z32e8f54c887c0e9f66d1f89adaae7979aad2a6a3b95149cd1a9ccc2c46826e962516728701e3cd
z973b8aa1fb405965c9de6ce9d1bae5d1716b94114c82d5032ea55509f7f77e1b8ebc3033dc394b
z821e11630f8d596cc71bcc75ea3856844f057e6e760d1a3ea398c1a0ced4dfda38943864087f87
z55a2dabfe5dd11ebdf7f7b13667beb6de5500de3f1737e77a18e33098dc3d5ba1e2641df4e6ac1
z5d0839f3d645952a9c4ea8758043ea9030e1e69d057f755ecdadabfbc811777e70e6c310341cd7
z521779447099397bb37018d4cab02b83117ab0af02d760be2db011f7425d109a40c23c4e50a395
z97ba103f8822c3e29db549b38e50d5cbc38378bf0edc29ebe68ddf85f0fb711cd5ea87855792e6
z776ac8363a697d7aa06ac1530fb25448be8bc197b55b2822b998318b444ce60870973dd6b302fd
z681e3c5a3e8951422f651680ad93d0b926b4e21dec1dd8a2f293d81cef24762a4459f9c1bc76e1
zb5892e29652cffd0910ae1e9ace48439c565be95c675d5df3ca5e05a1b26bf00933eecba3e3452
zc64605f5835644cdb3627a3279c1873de890398a442fa567df1fe23e8249af69bcaf2182ca6141
z13f8d1eff5d3d7562a004f10165152ecd8b2f3d15fc53d8b641315e895970de0a510838950e3ca
za8cbdc5f0829e0f34106e08aad22a121eac69639dea46b92df26d405f9f4c36a243b800f0bbb08
z8abd4f0ecfb6557a3b3de56e1eb35ac6100aef7069cdd0759205d527871b3fc40c0b43a941dc1d
z87159988d277e6d430c8a5df0a2acbd26d33a49e169464f4556444c6993a8b035d212a9f93919f
z269f795affa50a9378c95865e112d1edf75c561459bb39b53154334c9504b75ecbebfe4146bf8c
zc6765685ce08de73afe80cd71ad421d9110713bc0c0aa82e23a76b7d468f0da80689443bb59b73
z0abeec1edbc2240ba09c4603815c820fd2ecb6db70dcce393a2b43a78e71a78f0dc22308680ddc
z001cfac2de9981cc0659977a11f000a518a22a274f8ed0b4209cf54ba6a9faf42457c118b7a13c
ze9097a6df98083e3ff48ddb5bd0a8a7511e88f6e26e7c550cf3ee34a64a1575845916ee41411a8
ze6b76c3e51e013a6a781cc21547bdc46223444900fcc55dd0748bbee0299cce65337396f8bb482
z6e882028ecb5559ad9bef46ad7caaa058333645f0ae293cf8960943589d0c54725195919fbfb05
z693aefad74aef389085830be1d7c1ee10abb5d21ca20b160fd2fd41fda4448a7fc98f2a762ff4d
z87f1d423542e45517a1b5828a9c54423cb39565cbf505c86f276f63aa6a96f166340fd71cfbf3e
z43ce49dc7462572f835697367af97df045692ad924248e41c0ab744501d808f59742dce7ad98d6
z0545aade7e939f01d127e73a14cee0628ff354b79de7690ae4fe218becf9a5963c78ff3e536be8
z722a5dc6f3fc8ac1c967553e2bd3dfc81a2984bda650d0068954c3473b512c7e5a133af5acda18
zc71ad0f5fa29d6e18850c30bfaf6cfeffa4702afb121b6571da0045d7f642f4283720d283d70f0
z29913b6a8ec62af887102e8dc1893e8327c714d78f6aa0a56dc13e53d8aa0c1eb7fe7eabfee236
zea6c24a4c3e731739d86517abe47254df21759da5147861d9013c42af0c432ec5c89898b199445
zbafe281ed4efd770490e1d425b0dfcde5457946d26a9a8e04d304a3bb2edb8f0d215a32c465ac4
z3ba0263b865bcc20c0990746c367d1a45b669da93bc6c216a23afd7b699edc5714243df433cbac
z773a387309464f3dd5e0ad612ceafac6246b06a8c55764843b1ccbf03b659377d9698d609189b5
zeaa55e1c56395571d6bbe7dbb3f9cfad5e4424b0232e929ac5c49bfdd619a52b7b14142ed41283
z22b2622cc1ed2dd628aa05381c1f2a9960a51b96d2aebae9bd8e8f86643c8da69ffb09c3235c66
z74d46ea34cbe3721782d6a5911b3d4cfe7258882ab02191402f52a0462f47ccee21b9307d985ff
z65684c7924432b73f98ace11814653831f68c5adf995928e97fd050ae1dae537b85199d76e1785
z09769238ce807449184cdc8243817809ad046ac3462ba1eee386ff5e5c2968a13b18b64f4d0462
zd7779524d9d72502d95a7619df7eba256816d5edc069ef40b2d600dd2dca2a77c1fa6655cb803c
z16146f69381b2e81e492d25dcfdececaf64006cf59ad609dfd717da17cf90d801aa4cd2f2b9e0a
z1a03556a7d035ba9815a8b79194232d95d76d5d51872827aea96e39cc2d52d4f171bd6a7f1ffec
z8024e936bc114fb93adb3a04cd8d957518545501a667672139ee313c6836d1949c2ec4370e35eb
z1e05aaa73b8d66a338fb07478c9b6e9ec67336637840427eb0ea042cf2d1b34cb36d2d4c218ecb
zd20b39f8efb29e7831e22c75e2a1e7bf17194a541d1bc11b4ab7e497396a02524a4937b41087d8
zc88c6269ae417adbaf192cb44b5cc9759a4f2d238950970d75b7d48a023ce8ede23e083195f99f
z70e4fad0aac9ef753b6dc3e87c943ceaaffc243ca7787c69b7ef4780cac375a049086613087bd7
zdf1d47aaa6fcedb40c129abd5607ea76ef5d7ec95d9198043ede84bdb50e1077ba819fb80653b0
z8426327f108a3b713d1319ee6a77195e2314ba934b94eb3d9e306423f3c96d850e98d84ec7018f
z90da1ae40a0b106feb8e7e20e25ecc708babdde85cfed316227c539a68dfbc91222502d0313bf2
z340789b233d234d558d03a5c0deb12adb949dccbbf79f9455474ab2626ac85d9aec29d5294c7dd
zf2d972933b8868a117f5c5c169cbf2bd4ac0d70f11f01f05ff35979ade7d6a86ffc3a05df6a68d
zacdbf5989979beef5137c5954a7b28c55f64375f92d16ff78088923ba6c6e36cf49ab21b6c4723
zd72a222ceee04f0cfe9b6f842270487bfbff127f4da7daca5045d9cd2093c551066563ac514b8f
zc24e643337e29dea00924a3ccf90d9297f6363471510f9ccead1eb2f5997ecbded301b7b836236
z7d9fa90b412898b225ce7bcd6b81db2c4d757ae95c5b62883954406381501d69f1a3f286a00e40
z6d57aa81c60fcd73c1b657988b482e7334d31227c863a9b2c1b41fc0b1722e6cc798966a96682a
zf0893432f5a656a445069a1b90e2caa69b2c5b03a050d32e264773c3405fd8f48b8d4835d3ae95
zd4b27ae5e5dac4e3d5db9b069b999a83e81bbf9bd7adc8386dc0c337a540f05c71ed4ed5d2109d
zb263dea7ee57164c7a9197ef7f796f2becf9b2987a10da462af2139c8188ce9c3ac83ebbbe80b8
z62c48ba1f572b90e1e9ad2e1c1cff32c9ebd9d7799a96413bffd7a5d97951d4f8d3d8c68ac49b9
z256c481b1e8cffb5b98ed1144a42a49a7412f28c3e8978ff7b21c98d042a999b4f14626017796f
zdba87378b077737b89d1fc94ce007a0ca984165b4c483f97c9d6272ead21b639a5f67552846ad8
z605e4d79da5f7303e10b75ab9aa074896427fb159f560531615e81b2a48c6d32695132a64d7b66
z70084ecf53a7b43ba8bbe280cb189a6df798b342aa88ad90d3cbdba09276f5cd8f7f4b57a7459a
z503b465bf398a21dd546acfd94c7a9798f744540f6aef90810ad5483b6a5d1f5bfbcfc5bb72e8f
ze61af7d603790234f55f08bf35bdaa63d4428f6ee5a07138c64230f517376fef6968aa04a7b896
zd7c08dee442f50bcab2abedcfa022271241844ae201d958a04b7091bf8769598e131fc12487df1
z4030625979a90ed6b32874c883dc61eb9462d7e8eea7375a53eedc865aec1ebb4237f655423425
z8fa43f38572fa4f68af103ab556b36c015601539adeab29b73a8d83ceb2fea6f847866ebdc8a9e
z8fc58364fd8b958d75e50738c7591e1ccfa3d6897f129e944e0cc03c4b8a7defde2ac9c710e709
zbc9446ed7530afb960d95114d7d8fb6529f53659afe5b8f50dbd03a9cebf085e62d7c710ed4643
z365971b913d900ed008914690974e85c1f1a09a30bdbdf906232e2613d5ad017bb4728b6d9164e
z53813961c6e674cd1acb8feaca33e2964cdb6028a09e4592ba69dab300e0b8df4728105c5befd9
zed17538c88103139d7451b46a3aaff8952191e93e12d81524ff94a2651510bd150f4d55bcf4d14
z5fdf55ff9d259485e6c371f4e7fce4c1728813ee80e86dade180d09f13b7bd1e4c64ce081c665c
z51bbf2f5db1727526debc471a3d13bc5019afb3a72e696f6d723cc8bcbeefe09a31feb41400c70
z479e5a4a019c1c1fea9d495371b298299e66d6cd923bb38df0af4cb78560b69143515fa9dd33f9
zc2fcf4066c598bfb7f5bae6a6d9b015eaebab0bf9fa4cf629518f96117f8275ac36db975aa0f67
z92f7e287113114c1d6983625f0e4b4cfdf41039ec4b86f0b4d2c48a62351d966d90cf868a66640
z474a67565f8b37cefcc2bcc19744939a269bbe8e05e45c140f09c4eb029ff0eee42584c046bb0f
z370dd6503b232faf9ee952db07f16dd430ad19ea06c989a2289c37762aff0cde92505cf57606fc
zcb24a8b36230386e31136bcee1a9604e00ad43a26c3aeabe425e4c5ed54f1bd7d8c4b304bc31c1
z9ae5bdc64bffc405f5584054233a0efc13e9717f265e114a90373e0a09fd39d1ae84f623dce6d8
zacdc5edf617c7c54075e824b6a7675aebddb2055940523f31b20687fdba5b26f2a86bcba98f962
z4ff49a798020911858b6197610d751f9e75e4af998ff72dee7f4cdeba634abd0feb7a9fd0342e7
z45320576e7f824c3449b11f66278ceaa49c86f4963924fc68a249e0e3fb84f5e66530756b259cf
z5ec67dd43cb0c3744be51412132b876880bdcf27f58969f07e0c9ec2abfa0ab031ba644093ccad
z59057051edb2e14dc74884068b194b78e44bb008c6e15aa6e9bc3c35bcebe9b2c548836acafbd0
z7457a30267c5f15a07ecaf9768da3d68e8f3c7b17fb455f08d08aa939f5c8d8fe8bba77499a39b
zef924dac5874a6cd5d824da1f38346bda9a5753b4762c8a9cc4a2c1e18692afc2e06c3ae64e29b
zc6318cbe7dc2fffddaae2750b809127dbfac6d27d8db1afbef8940c074be2544bc7e69969d3be3
ze9e09c724263fcecc25ae5349bbd78d3d56cf2bc9dab8e34847f8c264407613aefc6397f62f26f
ze166601e3fcdac1555d54492582579e94c30e13c6ed7aeab27b7c0664318db8cfc0ad4dce742e4
zd44a2de5d355d9236ffc0b70369ff279bcffa7dfc41183865a8c396661164d09b96c3bc9e54f01
z2c24b6e7c227fd85cdd99c2a0d4bbd39953898c82a45ff0fc17f023bb03cd899678b3cf503de4a
z8fc6c3adb7f35c929c71c95ab3aa8da4cd8ec276143baa2ee65cd13d92f89a208d854f28a0482a
z9efba363698a727f67cb795d4433184fec76fc519e6aeacb33d2c10568b7bda06ab30ec2d06ebd
z6cdf5510c8b83830d387cd2eb902e8186a4494be0050917dd88112c974631dfb576f6c3158ccc8
za445508cd8f967bae165e56cd6e2d8740324c6aa18cfc8f4eb06cec13bbb54f458023df515e247
z88d39d1655ef7ee8e8a7257ff452131040b4e201eb13efdc4286e2c8689da1cfb744b3d66adc3a
z61b3e923b552c0998abd24475a1deb73638f2970e10c1219cbd3e9e627e466d5dd0703d354e44a
z16e5b6333b22246d090b243413b4cda7077c47e446914148e2ee55b263b946dd61bb511caff7f7
z033a8b9f01ca1cdea4ff34b8bcb88de597597985d1d00ce02878f2f5c5730345f7f89dec964a37
z4bf0045c4cab50471b0bc91b6e3cea59787476e8b2e068d0b3bb915af1a47756e82f3c96d1ce1c
z98e656582a707b4972adb27cf576392513c5dd0b8e1507244439e2a6bbb90d8d8c2dd378feee75
z18ec4bd9bdbbc8074ed06af8173786c90c88d3b6f114fad121a41a26c9107a7319b23f53d16df0
zd90253294bfe709814eddeefcf4b8b380fd1ea865fd33f1df746a838842ecae826c4751c5295b2
z341b746a158c99445f160186c31ba98f70aed6ab0535f732bee1562d88199ca15550a209559476
z1d350348ea6a3cc89a4e600c48816bf62f54f60fad762f01a5f973127013cd1811e9ccaa8c585b
za6b5be9216b5c8ef44bd686939854866d17553cfb4814273095dbb7e27a39bbd401074468ca817
z870ab2d1d9ee3d09f2e2d65decf21727cb5040cf02f807dae90ea8f9080652be93deab43d5dd64
z33066bcc4e0bd03e6a083668ae65028347f5e8a06c06e48b699fd087a2ed340425847dedd945ac
zff4dcedbbe986c20a43d6b34727cac4921c10f8519e6e98b68710c07ded529ea09606eabb3b286
zc108f697d82adc9f22221a0d2ad9e097f5cb733e64dffe3fd32f40d214c7b0f092992aefe4015c
zdcc9a3c6a7277dcb490433b2dc0324edd96aad8a1a7baff74844d18fa406121e026b196dfcd04a
ze1f9e26c6cacecbb2290dba92eaf113c6cd4ab3a2c041c5be850875d16cc66f1e81b996efe9320
z17cdea5751846d080fae7a42b9d3337e8aa4a899b5a4b97e68870caef09a208148b9deea94b03b
z9d40aa94fb938a424d48a2f7a73b72c79018a8d9c1e731f49f5f07069f726e50c0bb4aaacaa2b4
z043fba5b07b7c1b511efa0b534804f23ce6e3e73b45f212a9acd199a08173bc2039bc4e2b2e256
z796a3ece0032901bbbcdf05f62504f2c03c73adc35c11f0bfec0a8fc14a60b776f7055f17224f1
z5d10a4033b35c46f0a0f10949a964fc0ed86130386f1ae2c3a96894d60c8b4aee0ec9d8038862c
za4089ba62d94f1e11e28fce7715cdaf796ed7e2c277e6f6cd063dc03eaf101d8d1e1f845e6d8ca
zd3a0ea35116a4c965a5f08bce7391c31325a388628dd01f74a346e3032a1c0b10a4115d39b93ad
z6756b9ac61c96711ccfc86dcd796d49992b09ae34086f106c1ec26a76555698d1b60a412ba2825
z59ef2d213b936e76d65f3b2bd9bbfe5d82284dd5b639101b26ddc255b8ccc9155511d34de5b59b
ze32bc336fe1c8bee1c4e63cee5fa8bc9c26299277d6417610b05552cfc000862fb419c76a7af76
zacec78edc8626f6278e4af596e3ce87f5d8d23b4917e7248649907ec0b2c0b1b335397dbb9f1fe
zea293a7fb22fcc64909ba5793ecdf6425bea1cd4de720bc221f4075051a368ca764d2a13083a64
za96b081ef8e19631fb6598527dc2b2fd74799817a0ee77f4fe44e8d3c175272c43086e4f10ed88
z7802dcdf2c45e63a08fab5a9e61c0f841be4826bfad5ccec81c89838235d82e827071a4e98e94d
zff6f23020eac7a1fb8feeb45c4fdfb11aeb21968a5a1ba4d6229e39f3325221cec7d544e14d221
ze66569bfb267132f7750689eb15502161fa32112482ecc0d9c85218d75b0b9ac6b047404be6302
z02787810b435ecd0a0e194c3d2082f1c8c185a5b89789cd62efa5594dde0b24eab8735b18ff607
z6ee6ac6128b63a596495ba9f4eeba8136465d33c920fc136a3d2adc9a9c6270ec2757f3424b48c
za863531a5596a00a77456731fc7d52c70788ddc9df1855f13dfe4582b4756c7c4fb740d532c2c1
zaba366a400e8e47a0d83b6d7b33732c1387145aa2f4094bb8d9743e34528315d70e6f75f7e4a23
z03c344f519581513900a5ef832e0e469b337fb0097e088b9ded80f4443de7a9d8eaf06d54992d7
zc9027b24b40b6953d51353a552eb3b111fcdfbb40ba267787bb797a7309e0239c75913c335f1b7
z3d8a5aeecbced350eeeffb7cccb572748887cd8f64f496e71f809a175e4ea06174031363c0ab02
z8808c5d2bf14e933ee5db503e794911315afcf0120191505908e19cd8dec70f6294ca14f41c035
z4e1c04e4217a9ad3ad934aec65f76f7c061cd4667310db03334751e3479e096952b746cfef3a0c
zc17e95642cec4355ff15f584ba762b8a624324a5ad131f5c29a99fb67d542fcdda316e99ca3817
zb3a8ab4af1048c42304d6805ad56180480dbfb93033b3fda8cb2344f88b25babe8865ec7b362ec
zb6db2d69569410a5e2291d4a3da64ec891a521853d7ab1650d8874bec4d399f40bfc00fa6b7dc4
z49f828a070971407648b3c7731cbaa67a8cfe2667d07c796581e4cb6e86bf35928e9958dfe3f8b
za2a724f573fa3d7928783ce6542a1fb5b09a6d308e1478da435d66dd88316c92f0b57aabe51b1a
z4c686da1b81fd73d73daf46a98397f3feaee2ea33f04ac10c781a92b9f0fa7891ba60d04e1ca46
zaebde0c3537711e73dbef8aa687a6d457c743440c22cba205ee3e1338679c462f24e2654073d69
zedbafdb537f3b6c70210f3ae53875a1686ddb1a4ed1f098f8f68d8d102cb217564eb196e186521
zde5e8b8a61ec02b93bbde6f278520fa806d86b9fb60da6d30c7d8f34577a8dff005381bbf3af5b
z49b474aa489d6d90d27a55621e1fdf604a9c0e89d6f9294fc4e94f14f141b55ac27824cb03e501
z17fd1c679bc1b22b43057697cde378e811240f3c91d450e85d244ed0a73d53b6453eb41108c1f1
z9777f82c12be312717b86d8a7de7273dc2bdc116c0b0c235324a06e3abdcfc132d856f53fb5772
z72c5ba5e3db476bbf44528d9e31623bdb47b594ba98f8115ce2e6a0f25cc0a987185822a79093a
z1868732c0dbd5cf77b05bdbc9003d7821dca209aee71ed20630ebb883ea6f258f6a7ffb46da3da
za7eab65f57bfb079f8e314546805c03047d331879d9a209a1798394bbf914154842732e1048bc7
z1ffbd0918cde448eadba0a114bca77497c3f848503ab23f1f908a987d99bebe0ff0e52b92414e1
z8d65a1ff5b4ab1988e7c0c2ec8a701d7707e22a7c9558036680d102e6ca7bc28a498f0db15c238
z76bbfe9ce565fa177e6313347dc48efd30808b4297c1e23e9081f349a2877a0cdf300493dddef4
z942ae97ee44b04e51fefb7f4a009dca510076d89797d03f6173a27cbcf603c2c80e2dc5928ded7
z82eed93117eba26996f3730792f9e818d65ee1d29a4cb73b0462a13dee529d7ff83ea7287623f4
zd0e17c0e2bdb10b5104401501e1f599cce4c91f9a4716e083b3bccb80ba4e8044663e800a17475
z65eab443772a1ef7e6c01bafeaf2f92714302283cae052bef506302893a508df161c87854c7eaf
z4b35c4488857d93869fb932152a834b353f15d7d29f4dce92577c9187c9890cd601aab866bc0ab
z6242842338f1daab602edb5af8524015ee7a370ce1cda257479d0c7f813639864eabca6822572d
zf50f70e1e4e03358c962606f00cd6c6a22bd2f172c2962275fd201aebc2e54c3d5d6287651a854
z6b18cc0b8cfc552f2047920d7898955f546107fb2dd291fd3aa48ff348a6b6491d15d0d608ba6b
zf47baf96a98ca2f968b1c20936ef7cd380a73745981c36c0f3a31cede90893b97b2ff9e05fc3e9
zb6ac6953ff3c18ec07be3db9727a66363d872e8c8ec38b2715756c4e216877abd1aa5316078350
zfcb42add9bb08ddef9e9c13e3a8f66673ad14b91456f83c025a4a2b5f26c51690da49cf4fa0106
z1a8bcdb16a7ffd738881327163ed5b87d72618346dc97f6cbde1216cc1630ededf22037d1111bb
z297e10d286fe396899d79c7fb1ae9ea3fc4904884edfe18552c08e673608a25f8d2660fa06bf88
z658e5ba8daad88af7ecddebe94d8f5e16860f948a5d5ee7b2898c5165300b933a2fe606278379a
ze774226780d178e448e6b75efbef21a6ed5be8da3d57d762b44a65e92bcad1b265cb8b51e519e0
z18159fdfd595f8a8b1c0ff13d0e484113c6cd87f2e58c0273618caca5da77e8e65948cbb21e216
z73b65f4b3a313e6d8ca9fbe4b1d3126bf8069f83e81538432918c9b4ac6e9ca98bbf29a046c84f
ze7bbafe9d37c6a793245229a2233dc33688ddf9d35470753fdb1aa90c4235b74ecad734b763f54
z60710a3977537d029d10f98832c5765576149d3115614f9ad3ee5cb79ac458b45363cf1f00e4f2
z8b7c8c1be2c6d2f9569b36d186da34ea444186791ae4463ce0cb8dfb5dc29400b88aae6f91f2ff
z4f8e89a05438d5b0da192bdeddf9c1fb5333c7ffdf562fcbe88e00e3ce38336255c660b66ad4ef
zeb72ab80f9b2b80abee20ee4339d564d47e3e11a33e954aed5e92796b6b7b115874e5809277480
z19341898f60f67aedfbce1d5ad87b1fc669874bd994dbfac6fd13ddf249b2f6703c0e2b86c3d6c
z896046ef31f9fd0f9dfaac4b57dc744368050e905b0b7f4febfe741ed1afdc323e3b3d64cdef06
z6ac17e6f6c9a702df2079ec58728eb6350adbf6e1f8bc12c180a9b9b46f7bdfa051a4d6ae0ce5f
z4529f4cd7fa65d8c647bdca0d81fe7400ced14341250dbd459c37f1ed83ffcc875e1475cbbe459
z3f547df2a3c0a5cc1df7d2d1a7e4a407ddd0f9b6a661f542799736cd458efcf3b6972707e97d25
z0b57be110347aaf62bf8b77ec8d6987732fcf63357a87fbeabccb30c4831e99bbbb6c031573332
zce25675ed62d04633055a5d7d6fa9f32a47731f4281548850891f3c35989a859052faff985af69
z2862fc4a0c23e3be69529c6634f8642361a90611a6f5a90391ce8ab5dc9fb85084615c8cadd30d
za931e9e0e16f81c00c3ec819bf3fd2f2a2da01b152f230a11fca787c1e81f7a210f6b8aff08889
ze980bc2d67f90e6f75e3728486dba8ed3027f0b566ab7445c7a37ca97a11116bac00355b104fd7
z18df3d725e6fc6b49500727e2ad92d1f3554befb85f2d33eeba0d8cf27569dd2db68f6debd0ccd
z83e48dcc2e52d4eb17a81dfeda4a94a75496f8c40369af4eca0ce820345f3517b8f9a3a2c15f03
zd05f9d165333ca8711e24ecfda17700f631e17d2e36129b501c7aeb986bebed653eea0d0a839fe
z4e9e37434cd32a6452f5e2c84ebd330d5219afbfbf60d4feabda063c64ae5e925b36e6a2eb7667
z9bd2bb9acdc73e65878b924983f2fd6301d4da36ed58280e052c23b608fcbb9345f40ad75b5718
zfc65fe29666e95a9d31a9f8a2a1b4f92e851a01a4cf27bb9cb120b16792adcd70ffb7549ce691b
z817805d6205d37c95406d66ee71671240954f931cef55a0edf5bf60be603e275bf35c8237b1838
zf9a6814c20c02f8be11ce7f89ac040e475fe324dd3cb9f7239b4d9276dd60c9e83d9c68334d8ae
zd0b1773b745fc196f1c03a8408e4f6700c207f9db373e6e8c751609662565765a98dfd2321bebf
ze735eaf8823b71c45dac42df1d8a045741ce26d1a7256951a200908dbe93812bbee62d35199047
z57f70ec2645042874f53b2b6cda84b29bc0ee94de31ef0bf07e35466ef9f480df7d571962c3de4
zcf53b86f0cbf6d31aaf37f0d274aa645e838861f1a5e31a31a8ffea45de18d81e594be53287d2c
zb671c06bc8df69ca61b59a491478088608e9e87c8cb1cef2afea302a7c645e1b857cbd7c217260
zfc325ebd9fd0bf6517f7afc7c56ef6b82962d9f0f14d39a57de6aef8f9bd589f167c16ec42ddd0
z23081362eb096e2ce62ef5890cf54b32ed51cd1d0a9547fbfa1fe0db61599647d9f4c73defcd50
ze0145f9c5ede8e1f565f18817c829545a32c0927b5b5d7e61d0e18591e397a43d919068e1e39bc
ze97b7aa8bd0631ccde17b9f1f2099faf226d36cc4dd3c02df7e5f83756a84459b394b77b669a32
z6585aac6544f9f59597da6688cdc54cdacaac4aa47bc4b401690319ef88f3b76c399fc4e45b6ee
zcbce19a23400020ea8c25308347a1d4b1a7c8592ac391244a065867dce5a03a323c18451ba6144
zf09a8e48ddf9ff222426b60d17536b4e2b58153cee70ff53f00ba989c72de7ef5d065258ab8c8b
z08604a9236f40834ff7d322b11e88b76a729c8072f81af1df7a77170921a1aa3f99808ecf9adb1
zd37f0a2a025d4ac6dd31ff135f190037c2e43d706bc9f647e0181cc65c81e9f97e4d53545d6b42
z6c73fc6439d1ec5119c0db1e34840e7eff5c14fe91e8276e5b176b663bbb79c03aeea9779ae29e
zd6af0148d2da3eadb7a31ecb48b3e3f6e08f6b270c8c963489d4b4297fbc989b8bab1f9408b50f
z5de95f8d3246048ea36d89a2abcf580f14635569c2d4e7fa451e82c3da9e1ce6b0ee909ce1cbbe
zc24f046aa7f3b1090fb62387b60f5846ec2a2bc0f844332978d1ade4090ec836ccbba549b91371
z1f96c57eb149cd3ea10d26f948bfb9f18d95f62bc80429efd1facd726f8728c1fea64d2a502e0c
z1896577963dcbf52c87585ae5fcbfec2bc476064f3e33f9aa33eb9cbe8dac1e01f71eeb1d782f1
z842ee79dd1bdfa8ad9f0309cf3b2629a8497645a2400396bfdf43c359413278a4ac5e3a540aeb1
za3b127d723e0e936fc2d3233af003ea68babb1fa48226fae9dd9b5b4698dd7fb7baafb36acced6
ze62ac4159c8ca66180ea5bb67c5090b34d32a0befa527b7daa175c7d29206b9906a77447a80f96
z527ccfabd2963cb9a0d5322e7c0f23476b65329f64e7d87b932168ff71ad81d4c79e195025a3f9
zebc6094071465516499ed12a61efa1268bd3221fb9efc790c1dc8c3880d08aab3174bd1cf2ec05
ze8a1f6f78ec4fb09b5feca14849e2fb010605bcafd753827fa9dd1e790a96b5410d0d25967057d
ze46462e2381a04c001bdd2b3b521e468fa80cecb0c9a65df42c560dbad0f058ec44db6f7e4a744
z5ff908daa8dfb8dca0398024e7f953f52182a87c2e5eb86676f1d93886fe7de4f41045e6994b2a
z8516dab7d2037f636ca3e79263d1d6d05a914a699efbc4e0fb158b9e25b1e954e115e4ddcd661d
z710972b64655b0f24d05b4f7d1f00489ffccde0b298af3d63c714f52b088fbf0c6e1183d48debb
za6479659409b2eabf4ef0ea4053189eff848422c1c44099ef8cd920ddbfa65cc6cf862c822e8e6
zcd34b4295a9438cb309809a03dbc0a06d6f5f1b13ff52ec7db7f8e9b6da734fc3c0fdfadac98d4
z73325444303d75c8d738aef7223086e064c5204dfd72ee42fd9993521374fa155a978954a072c4
zccd8dfb215d1d9b046513f2af5b54a0f25e33b9a60f237a8ab969db1ba775f7e2fed26c1900cd0
z8192121c043aaff8f6d0e30900faca433f5c9cf434be1540ee261d087e52012bcbe569d2c027f2
z863369cea80aa43405a39373e8923e7b09caa8b721856b56741c7f4499dd27cbccb9ab11d38ef2
z818af1857d9203d615687fabc6dfab9a20495b484d0bbcd38af07245a6248d179794bf0a953fa6
z1379762938f4103e6d8cbfff7b861474037935416e61c9d51c62fdea58026ce6b83a9523a844a5
z55eeaa09e2bb9b6c0b55c0e724dad0742c4e3276709617040f3a3fd52ef8a7d46dc4e6b7888c88
ze5c7a3bd7a7afbccaaf0b1ba0574431a0ce5e9dffe43bfa08a0976c964cc2d71f12373c28e120a
z0f470b007650e6b18fde2d2dc7512ba9876f06df718541cf80e1c4b84e40770bd4924ffc504738
z767d6cc3ed00e60fcf356de5e6ddf2a005787decc241c5dcf5ec4358e70effe4825504c10a3347
za206560a3564d32986fbc54b1e3bc2adac417b40834854e199142d0b7224f5ad231ab6937284b8
z1bfc53bf44ce274625aa7e441691a83a60accb10f2459004bf5f87eee1d183f17c9841935cc451
z42ad81029f5e8387cc9b1496c319ff4befae66d23732d9c4f56add08b26c1ac6de7e56036928d5
z6e01ef5ce822da39a8b117a547da30fa8b15a68d90ee6beb9d7360a0884a300bbc37efa910e06d
zf8e2a3798705b425080a9a9cbd1ca06f5b41dea7026ec7bf0229cab459716f444967d6f5a3db76
ze9da87abb3caf1f61c6999dd8e6b6db3d23e5f20e0e6afead9a6d38d3d069969273b4f6c8245db
z10ee0eecc2fccca3fd7f31d4ada78e569f1a190662f08b4ec9763918c7a3894698bdfafe095a3f
z77216627048bbbbe386e9bef9ac4d6e796fa0bbdff6042651103e4452c0d710c95fe9977a92021
z43605d33cb0904e59365f1bc3be334db9487a34d92cd96cf1fddaf0dd017f9cd4fee6397ae79f1
z906932dcf5f1c54822319a8ffc02425b91eeea2615a096939c56e4965d8c61f56b038a0265fa64
z86eef966874732e49efe700c18cd97c4b8e688ec8e3227a42cb8ebb54c1958d76498ce798eca9f
z217007164d89928356eaf6feecf1a512634f014ef8c40aa8c43ccef2dde47c7ac1004198c6cb1f
z2914d704424e0c1ca708af4fd0a158084be7eb5184eb62a4acd6a017da6cd66fb0a51a0196d570
z1bc10ee2c88c58a508c6e98212ac459cd91fe4832004e671ddb4b829edf36c10b7bc4924494fff
z9264869cd54df77ce565045071ae38d7f36b90b84fe7611c11f891e36b67377df513e549440a68
zbd4ac6209892e15a8b9f8e8eb44d0ad29f90b8182a9bb1e455e50514018bfca070e4f2e953c8ee
z1d12357dc3b264da1e127c673a1e2e948558c811d28f41b9753e6dd1044208983bd982cb0efd96
z208048acc0892ca49c0acf7e7ccee538fc55e67f53349b0d929c0c7e4d90068bb6ea4635c2f226
z72b418ff6429c98b3ccf109c1b4919b7f268e0d5eac324cabb8a8e78f312ab8c7a7f9673e11704
z23c3bdd53e11dc4b6f50513917843d4cfc540e2035c82f7161b62f013027a2c1f7abc56760a13e
z78d253ebfc3397d705b9a264195f68b93b001496f60e8ce325f767aad0aae49956e77b16c67225
z0dd2f275ad4632005aaf6c4a1dc381d8ee339848c73307303c451af9391b1b763374ea65cdcfa4
z82c1b4b027f1f21034317194a7694ea4e0ef92369f2a2cfd80245987bd5bbd8e7459722631d0f3
zc3c542ebc6984ac72d28c57f4e7b66f73eb8946b7b492d21d0dc91bd69a2f569f604f95991da5e
z42485f352213be78184de368a2eb5905494613ca76d2705015fd8c75fbba99fa9d1283681ba222
z36fa32bb56305bd32c994f981fa8ae5e788e183eda9fad7b5f863f2b401077f66b39e3a6b0e21b
z48bbdf2fc9c1cdb4edacf1bf52fdfa3d40c1fb967a53337f567691ba48fa2fece131f265f01772
z111e0688136d585e4cca55a6a482a0cf9a8984b243a548437f2e0c3f6cc6620533528efb6ea49c
z179ec1bae283e59ec0a12558d1e069150d81e906e557da45c8c0827466fe2abd93bddf39912b64
z1d79a7ccfef012af3426648c376fa9da2a5b68b558a4df0809296cf3f44eb91050752d9419ba9d
z7fee8ec7cbb399ed7807ef2170ac5c01262535cc074474907081ef608d8ab7884078c7973f32b1
z947ac5acb86c85636ccb3209fde1d6ea514ed3c1ee6911e37f656ac731293dbe569910ba66cd50
z313defb8e483a2bd45415c1b3c575d4b8f33d8e10da89f9b6cf480cbde7f10e88dac0a5d093ad9
z9ce2fc7ba59dc5305870380b873a33f8bfcc977677934347ac374a40f3e62e60e9fcfbd1d54166
z7a9913829f3d928faa108d641afaf445b5eae6530e5f77679bcd91b5b41fdc93f2be79b503ac67
z1a3a8ee1b119480786bf69263a72318fe4cceaff7240d11245f59653fc18b601833ccf18d59b23
z4ac15dded97347c8962213e7f67b97185ecde6ae4dda76f996a570ba49616fe90d5c5f2c2da665
zf80dd3e89d88c8834e911ca03dc312bbc1b0df2d2014e31264a7dec6688aa69057ee745f83ea24
zf48d9347fbe5c2ca1e3e7bb8796e36cc77c898dbb4a4fd759396ac649bdbfe49bee406b23f172d
z2faa1a860e19faf66fb2813bdede9495d31d35a2da0c02737d6e5cc0c163bcbb026ca7fbbde25d
z696480fe66d1c0ea0203c513b09580dbdee7048baec9441b3b63e79da9ba6fafdebe4f6684bfef
z22da108c18c2d3b6a0f0febe47a17cdb07fb428aa80b2e083b02b8aab42808a17eb0a225087289
z2b04843783931b0c3ee5abd975e468b55beb81fdc14e7ea4d3735b5dbd9e721745c88dbecefe81
zfc1befced01a55216f24ce6dc3ae483662a6eb5477d7ce5bab00972f8100ea57bcc74606d9fd90
zcd5cf50b1264158b3c398911b547bfb0036a57ae7c6abdda41de43e0e28e552b1f14a1e2c575ea
ze31e7c1f34535f3d9287c4094ca5a0fbd06e6061ebb7484b3e49a9c47c87d6210f45982f6be48f
z7a80248956f77c54838627c6d288ba49d637a427dbc0bebb82ba47fc1bddb3a26bc27f86db713c
z5d182687e0183439721834bad7b9cba4806aeab444a1116ebca12402dcfd895db33d39c35cb286
zf9c96c6b4361cfbfa61a6878a4ee360e57a35765eb35a9e11badd0a5fe2df45b9b436cef1c7d7e
z7ea934e1221c4a509f58d489064f2a646ab9fca084c7269b4b9e98c7bc2924881fe3ab0320ea92
z4c65f188d6424f16e8047316eea9205e682f467bc6d5b0a68c9bf309df2edbfc3de2d578596072
zfedd451ef0702d799569ce883e07ee3399939c1f00a6d9d006e95ab061c0bafecf7d9c3092a737
zef5c183654f5f8489699ed0fe08fd6711286e89c192c00304c8a22ca9f03011b1f2697c4f278c0
z38b507da00ae2199f9d5549ce5d0e050a81acd63b555564f3fdbed823bb1324b83cd378bb2627e
zde59234a668383f3fd7cca4387eb800cd1036e8566e0aa6d4416d284596b23f2ca26ae2d28428d
z940b5a66f63f8083eb70251aa1a72c0259658e4fe4ecdd590db3a3a6efd3ec7182476cbd0de3ca
ze46a86b690ddd8c581ab96b38c436e15278e1eff6828ee06e1cfbd9a3a86566cd55f4d5952da64
z450ebfe3d24fdebcc01cb68893eef64d0340422f3c7c18ecb29bccbdc867ff9aa42e5300be637a
z96ba6faa6694fb312212f19c43a50fdf11bb969032bcf4f803f8e0ed7cf0ea7eb8653f4e03b0a3
z23a7d18f199dfe8fab7e1bb83e7bdf551dbf46d65e7e9b9e2d615a91f4c4ba58a53418c2e8388c
ze6b3f1b0e2c427cfea0bcd3ba7630671ebd0947e8af331ca9c64cb53223540810853ec970cf72b
z12286098cb5f12d6f24a7c933843f2c3c3b46c726cc2da9fe3749043b283a0b9ace9fba61ed720
z863752486cf3f6402a239aa416aca488a32364ff9bc1741a53746d001cc9b2a12a795e5bb3c3f6
z80cc687902f094c65396936ba87d0e405f764621a94fb2a107f8707bb77f09240007c2e0b47cce
z89714f831d6a1dd3f82e853562c7cff35d1d0483fb2a471f3ca07e2e1d913daafa63615f07e0c1
zdd82f89bfc3795c053be89c912563bbd317ea9064e3e1094d84746194a862a5a9da3ff8a1c8c37
z25b724023d8a70a997274052616093b7d779c5a5cef07d5c35126b718d8686c483ea6a49c27ac0
z958edcc2a72ab148f1b0bb68dc6a115afd348ddea0498c874f257b32bb74ebf26f5bd76ac32ea9
z6123604f36a7272fa791df36adce4a40b66e1746849a7e3b5ea15e171a02f227f6f6d1d546f5a4
z53a608fb2b37955a77e033ecb1299b2d241e3fbbaaec41d0a8c7587be45ddd18f74826f77d2d26
z60c24d9c1dc1a4ae6de3c7f0079c010140be2646c4c71dbf2a6637f84a738c5b6e31f1875627bb
z78545e8ccc19d407e2bb52cd5c58c12d490d33c83503bfb5a0b9584b3983f907b75c345c3b2998
z52312afb54ac8d4c5d2f072aa9e6eef012b86de56743dac6e30fc130274124a9545b86061c02f7
zb0a3488577992d7797795984ee6c03557ab145017baa34a35a765712c01653cae59590b61c3c46
zdde92acace00d5821c1ed402b5bb48d57bd0f06cb6200c1bb1e5a2143ef891300a6c8bd555b4d7
zd71d60d778edcdbd0eebf1c88c5c6212021639951b9443b7e5bc0ed7bf60a79001f46fc2d7cf38
z9817ff568ff4b77c267bc91461556c4cb9d135fa8745aa49b00d6760c5dfa0f6aee9e854f20280
zaa74132bc70769c8c09985efe8ab4c1338b5e34417272fa182ca83ad0b57d677554890af07d9c8
za3311ca56b8200b8e9cd4509e2a87ea8d378f2c477afe8c8a5c0275e34bd8460748bedf13e606c
zeaa288015c17073861acb22aadfc0a95581c8aa6fe024020fc9eb935ed38ff4b6f8557c0f33d45
z36157d38eae95c8a5e33ddb269c33b352c95772f49199ac763b41b566135285464a600e8f12a5c
z420b583383bbcc1d5337d60c16b34e1d3445d99712de8aea7d34f8c33ecdabacb82249ab88b715
z190d9b18146a399cbf77737a54b2a522c615ba35cfcec7c0283c51b16f91563ac1d967aa3877d3
z10397891d46dfa2c2e62e4f5223347d05c90f9be88b11382e463fa0cd5df20dd35f6324dbe2f8e
z6919e57615d12d5f7121ddc7a2f87112b9aa516714ff45f227f5666146f379015618157080d0ba
z848e37e23dcd1d33845d5640e4eafee844f85440af3ed1b0ff20c5a3adf545e95f76076975c166
z022c921bb3271b215eb7305b0bc828efcba291556dff1e973deab3eabb5cca231e8ca3d683ee3d
za9e16f5c55f3e59ee86e76031b4cf8a5cdea2dd24250f48ce8957635bc9ff381a5c39a4e7ef256
z5a54be5021fc378c5a9dcb4b57ed4dd1e6df94af7813823bffc467adbb6190b8bfe5f8caefb8f5
z4476650a13df955c5cdd5423e061444ae43cb16f7795cb8fcdb18f6151be18e444f0c15fe9e504
z22bf7fe85faeaeaaeb675c5b33b485733255a7a33f8c35e73374aad68e4c2dae1819ddcba46e69
za3c495f71bcfd8a6d83f75b6b1ac7c0aad4155f228e8828d8267b2cc2b5a3fe87623609287aed9
z110e40cc13c8a644fe8a2520f88445145bab0cfb1fde349d07af4cfe4ecbb2068b209a6048fa68
zc72e5cbafee79ed70f68da2d01c79259305e9c99f9f59ac61b31c0bc1c001abdd8265c04a867b0
za9a450060d246dd65127ee492a8d36f3cb5bf1f620c678e1f9319c336ee4170ae8f6974c9174bf
zb9fa79bdcef46b25dd86d3aa3520a46a40eac903e6591b3739b4c89db4debb1d7888ea4c0235fb
ze3069d1aff496e7b248a130ee5b58053e4d192d78ef585fac811e6b4aff627ee57a1365e57ed09
za82253ae0b0db24b83581ca4be4b58a9ecf13d1faf66bcd3b7de3b9bacd0ef62ab04745d6fafc7
z541adb8afe99157a144c273b0075dbb65ef7d0877f2ee8b88dee29d792dc28af6a8f9061edd58d
zb4d1f1c71cf44527dceb1ac6805c201633a67edf47066ea878bc6a5add0d56b3adcfd9a6113b3f
z80aa6a8147c818949ff58076263c17a4dddc52b66bfef471ec3568c57f961fbc43e3d56a6f46db
z8ce210a03c6a6ddd14b3f4fabbb54de6c9577740a50948efbfdbc5543c102518a0f95fb27b3a16
zba014807e65f58924d80d17fa7ccd46b9ef40f554ab49bf264db3b1655797bd2468d23560ee6ab
z0e1a49e6437c0e948dad5f2bbf1d405bcec19fbe50c44beca1b0a7f82c2e2ea1babd97034fcf9f
z9541e419314a390f361f0c2401c40787a450428e60fb99739fc5fbe779f7b4d8776882db73b255
ze65ca9a6880b3e5128f113e2bc961c034b41b0aa01d6fe205490e5ccf3b0704c6a58b1eb72cae8
z263135b47b9bb6189a0dbc8657c97e6745dc056e144397a7a09ae540b2a45351f464d8c1a82a63
z9bb207a5ec4eecc5fa749f4cdfb28ff38790df132fbe50c552358058230c8fae07067928887fbe
za30180017c084f130f8a8b01f2ce05052bdd44b6ff805b8b48080e41347679cd40daeb0da01a77
z78bd7d3428cf1d186d2982bc05ed76a202c8e24ccac6a7e6d2c47b26a1119b539e8962492dd2c1
z2827e1ece58eb2470c5593b89ce042afe04ab6bc550bc4126b604b4fa0a14cc680c742e4fa9118
z05a66edfb2776260e66f05e39cdbb0cbe4d5470046e0aef3b7dfae1bfe7cf1b8875be577ca0987
zdff054b8ff037d9d73f58fe341a99b9c81818f1d883b0bcbb7f944ca04da994671271be6a4928b
zac8dd81dc1b8c57753ee32d4d5e3462a1502760352f8551f3e01e5c5f31170f3b409e578106cbc
ze4e2e007581501c441bd2691b08c596f9f8b88d6f55ab7d895b53bda2e0738892bae2cdb6ed4b4
z1ba7b444b7489044c1ab4d7dc5965bb0fa821a599dfae5d420d7d2a0e3f9b8e171e7563df50d87
z5bd8491940e9e19e1ad06b1d48de852d1572a0555d11f837f5745a3d3a2d9ed54210fdbb3174fe
z7cd8c74fe401d3d075c372671f39664c9b6a1b1923f0bc69e60c287d69dcf4429ba7207a1f3e93
z4a45d5086509f7b7e3dda512678b8efb8b402a559507ade58fdc7dae9bbbc80cb03508284edd4d
z87bc7d24a334f829d5ec5efc9cef8a87adbe452237d5c776f989bb4370da1f7f51ab0e64346d37
z34e17991028669c7d2347c0ffca80bd60913f4435938db1dac72dbbda7f9209f6eff7dc6f5bf7b
z65cd2d8df08ca3808dcb202298b1c0ddb4bc06905793cf2af88a51f8812f0f69524d03335fb4fd
z2d7b2e2ff581481304ed7c2c1fd4be4589612d3b79ddc07c81d2a00a8007a9b63c44f584d4bdcb
z3b2f0352ade0b08cbd1f3ca675d0df2b66f03be12b0d27b3fe567c79fc2696113f5f5353190191
z68a7f508f46d9e6856d5bb763bc12b62f2d569c21efb0611d82b513cdb49b4dd920c20b2d23481
zd552b1a9b261c0975d246b1fcd4b0e50c540ce8950e115269326524f35f6eae38df8e920d0ba53
za52f2f20e37ed748a30eaf5bb9db20bee7ee86d5d80f7a3169507646f08756432d9ee73223dbc1
z681a36169f27850bb838067b39bd345f991a78addc36813cac2f4db77ac6d9a73cf019f17ac435
z5778fd8d82acd2be8f47defa94544a5ce709cf25660afbb8b802c9964b6f4f143bc0b43f34ce32
z975cc9cca3e6fd03f90cfa1d6f3e5de47797a5ffcd0fedb46c1988bdf43d1dc3e21e479f82e99b
zd653581c9eabbbfbc5c0fbf4071bcff73ac90bc7ea69415b7803477c7d8023a16f556c98b4f13c
zbfd4054aa73c6abcc0edb59bb7662c6634aec7d05850ff66392adb072328dda360c33784fe71e0
zf60d980b45880c534b955d442b5d8ed2030c92a05c87c4140d21e5f44997417e18f0d1d641793e
z007bdcacb83e8ad67d9cb49c2a6b78d93466d0fab03b83c68e5d49f548e0269c4ac1ed02e83845
z8feeda4d399f1377ba87663fa911f728a9943871a9a2a3cd1839f906a981e8ef3592ab5545a16f
zb7bb3fcff053ed88a3055d826c6bafea24e72fb23259f576128617b1e2ab535b6761c63f1b0664
z17be45370b510de6b1c99802ca9684e2211ea4525e5c7486687cbd1665e77121c1024c94865ba2
z88be999731ff1b91dbe314b1d0fa3c6c1e0c9e94843cdef852b8ab29532feab1ddddb8e61903b2
z3464ea0b905e4e44531a337ecfb08ee815dc36ae4c3e8e95b941fb1e543815768c68172061f5e2
z8532d620a96614cf2410889fea6dfcc4e86d22448a1a9118e4e754b579cc907a0bfb04af502a4e
z258f8f89d9c49e07fcfdbdd1680ccc2c4f2ab5cc84638208e93f33888cd66d23aeb17fbb6a9aff
zeb4562d7fd30f1aff598f30bb744c7e5f674562cec6c8dd173a44107276cf242e0790771135c32
z2a4e1becbec7257361e4728f2113b9be0deab85263a04ccf076d69f7d0f09ca21a555d7ca634ae
zca534df999c26afa2ee8b04089b7c86b2b93fcadb10c879d16c8cac9a86fa45fdf3acdf07b8ef7
z917df36352908b9173ece583578ab0f2906691a0e5a68938cd82f9dd966b33b87c7deb045b8e98
z3e71f7e386102011e5c462240512d6a41369ecebef9d00066c82007348dceb3a5fb0b7afab7407
z302798b8ca5b275ae18baec7795bd3a4dab2d347c2b211d635d81ae4e9438e248430bda8bfa576
zb181f9b314aef2eac26515ee335c19ff2fdaae8449c25f4a21296607a10599a3a3ec7bff8db0ea
z9872885acf8cd7036f3c95b42d6b23429e3606e9d25d5c6cfdcdcf6f7b5b3cf479e585a92f0df7
z03ef48deb256807b7615e5fb0155a35b5bddda876c64466464196da53b423295f690daf516e2b4
zead17ea1b2ff5395d9e9eda170a2092e9ccddde1469dbe6b40a259bda3ffb38fca4f8366880655
z7dceabccdcdd134ad483606b5e6c2fb51ac096ad7d1fe2d418838ced1554a34353747578ef8eba
z5c094dcdc0a00563d1bd9c2e46ea4af37a753c7d2def5d56ea4d23c119a4fe35a2ad2d50ca6d3d
z6b2c802855a001d9ddd354dd5d234f92468df512f08004bcf041f7490797c7c6d8cb10c51ffe17
z1a74ac84f95b4b9df1c889247f3e6924a814e5612c13b9901260d8d0b7051fa8e3bc21f78bb7e5
z691942076bd7363d7c1619cf6724bbbfd69fbbaf88f5ca5328b13ef1460e16a7be86f844e36188
z0392323af17e68aa5bff406216cd9576c1d1e46d2ea2901f37ea2d487d7b7b2e668605b05dc6f2
zed2c7d5270af3099b9e9afc3aad5a7baaaa7e20eb1bfcc0a56ca7ab8e0655296df2a5164893b24
z04a43b3926037dc6e2675d41732e8c3f95b6bee4dfc8916200e5e3ad4d9f4d84bfb0e2beff3f36
ze3534f1d1ba5cbb60af94455f24d4cd462381fa5af34ccba8efe9185ece653adcf7a70147f42f5
zea57c7b3956250c281cc2fc0a309dd71843b5c0abeb00cd9aded9436a54838ec31eab3e1bad5ab
zc753a9c52e41d1b48073cb9ec070b8fb534d3c4ccfc6cf359ba5f1f9b63011ea213ea6f8a2dbec
z1c1b35e4485ea303267d8917d4b7fe114253c337d7f8910e9172f367aa6db9ccd485d4e38a92d3
zbdd9666cf3192a28d77ba8317402f4bc67d99adadee160e7f0f66563c829f50f64f27e77003bca
zc60a49d59c9647aa9864195db65cc8a630f90300aeb8216c156f19351cddce6aff3108906be765
z26199d9524924662db9b54a2912d3f63fe93a13c4e7c54f12f2c91e60ea925b54344eeec240e48
z9576325aec3f2612e7c2121bba43eeb5466df578585c460cd5423ee2e36134fbb28916c73bdd67
zac479b48dca17e21b27dd551fbf4577731323bf7eb7e304db7b4d3025e2c389a13ae124163e563
zdfda16bf0c6efa5288c58fe0bd83098f924d1c886718fcb9b6c594235c29f4d006f084e0731212
z1fc3682eb6f5980680e4d4cb747c5025d124cc455d142a029355f155c556887e243535d8c44457
z48fe23ba3d1cbda0f364268d0c83d1f316fd2c85eb7368530bfc78c98dd2c5ae558ac27d2d5f4c
zd92f26f5aa66afb972666ab0d9ab9e5476d1cd6c62688818d7c70d5668d2db96e6c70c02c78a76
zde82e3808e218dcb9be81b74223c454da8949bfd41b74969078ae363a4002c19290c251ca02e8a
z8da43db6332c65bfbd69ac8347c4cc09f5d1f4096be48cae6235269925620a38aa27d982930b65
z9414266544d25e724aadb8146262039ba9f2ac0914cddf6f4c08837ff1531c8229ac8bb07b0dac
zc97dae7e8cf135e369bbc507503e3999b42f11146590347bb40513d22adb412c4bc976fc0bfbce
z333aab68969101ec3a40b1242dbc4a8cb440c600acb3965c8b4879e866ae51035f90c80517450f
zeca8738351edf585485462b151957e6e81706706aea0fe7f831c5a31334dc624a54bfd44220657
z3346b7a84190b973d5da7788b5771bceae1d85f550fb1d60d22876ba43083cf9a3e4b6306e914f
z0d908940d8811305db281684b16c50a855fd0b1d868b349ee28de9ad991178142bc56e247b7f93
za89e50a654795795eb10ce6fbbfe0037576afe5f9df7122e53cf51da7a1fb4a414e11bb80306d3
zd74bc1f3ac8a1926205e6a7c7a9b88bccd7aef942e3f162691ffac10fe1330e26a54e0c9f94b92
z84218ced748005cdb58a8058ec81d3fb0f6889db90f9d0f3f574d2e23684518e40122d89d41f97
z089f6f478d3eb49a4d94677c891034fc09dd30ae0453ad9422bef4f17d0624f718d98044957a7c
z62f55dffed9858123ac872306f2d8e740a706f1570a5faa452b91e49d24e17d426305b160de783
zbed0ba4c3401a11ca0a55d990178731970d8522db0d39bb173a0f97d24cb0565eeb865cdb36000
zb4326e08e5bdd9f724dfb5c80bda2ce4ea81e5bbf55afd9f2950911afc031c6049e844b9ee2e85
z8da635e86d953cfa9ba6aaa4551689759170f912f4e2a90633f977ccfd3e95761f883c2980ed28
zc39eceee01016f12bdb2ae31337c47c63a5da892a8ed52a4ea1eba1fb464c32855688b8a66ac35
z9fc6c848e39c22da59220e17830239ed9a8961248489e5698eb3433aeaa23d17719b2c6ee51ede
zb990af60b8e4e6de00fa9049bba1ce7040d1201326e8e4c365b47b8d5044190f29c696ed783750
zb1a98cc5f2780273b5ca6e723cf820d0723d1ce53e7aba4250a2e8083ee3bf46cf80e8d0abe6f9
za06c755bb40bab58e6384436652949b1a3bcdee12d3337ef386b76bd6a0164ad3c4ea4618644de
z176b546f518fd03e695069fc61824938bc85d49c35829ef37f08ed3818cc56be36d34e4b6f31d5
z3733cd5ae6499ab1d5fc4fc3a077fe62e14400a09e7801d7ecc89d3cf88506a7e8d97b3d637f6d
zd4c393ef07723bf60482dd7e1d8e4b62cda011d800397124011b1dbc771b8c5ee6be11536c8145
z17ff797c998c89fff5e32ed333da8fe2f48293abf7702c15ec8586aed5b63d606d48adb78b81ce
zd3899d483a556980c62087f9424820f9b35e5b5e14a2b7f1853a9e4b6665e7609bab2aa33e7ccd
z71645b27abdd7cdd630122a8beb5376cc884a56f3da4be48191ed898531eddfe6d322cc906b229
z588276613acfb37ee71f2a5d76513502ebfa1b84ffc13f437c3ec81741ea4e8830f648f254f4f5
z03a77916b05d2d7d4e66fede818bc01f322d4e3336f75744d80161c2a280032e3a05829cea415a
z27c5a283dc7f93bc07d9aafa1613b40da60568e909eeadfb20cec10f1c96333359f282d422311c
z0fca94c5b5b9456d23068339a35b651782daa8cb33157123b58e38dd2fc18099e4605870da540b
z757ab27b97bce8e2ace800b64c49c35773af795197740c279ad6ddbcb73b3034782cdfafcb35b1
z7c559b4f612a0568faeff73fb3044baa4ad06a16be29bb55bd869a808efc9a9168a193130812b9
zfe25ef8119e670052c4f04c8d8515e02b14b27745fdb63385776723737e9d3aced85394a134801
ze534e79fdb61a5deb7630e18753232e1f16f67b48f5bffd3f85ac6a4d1d02aefffee75c3240922
z39a19896dbcd9f969c89e9b7799e90202bb4047cce31220ccb18a41cd1f5cfb8735495a38fe8ec
z56c75ffb9e0b5b0e021609d4dbfdd2476ec2c7153f70a16d0abde351690c07b6aaa357dd6aac48
zffeeb301fd6589d23d4f529810f16e02643d5e328bc7cdc3da7d40496eab0ef7504bd9bae0f187
z17d4d6eaf80a9f25956ec37f4da8ccff86f5033b4735d63ef8a6b92b8bee8ff918963a87b74755
z818dfdcf163f9afaf9984d7ed3ee1e1545db2fc54010dba438481b957ca43885caa1cf0f0b681b
zeaad29d7bf76987aa8299293498bf76c8a4d03556be59b16d0b569bb1509365039b9c6281442fe
z706dc49cfad09cdcf8905502a7ca46f6f38fb2debb48c48a9d4f45ed371c50d1b69e14b4463275
z785e748c2b6b49b2ba6a49fa9212d694ddc447eae8d63e3db385f4664e7cb00c555b20d6d13d96
z24c5617ef8439f3c520eaf43a0c957d67a8a6ae0c958076d6f6fb80f6e137c00ac11a3c0c95a46
zc03405b03bfed172f0957794943286304e5ab4315a3530cc419e6ffaa654ea71c517473c100d4a
zd205d306b127a05b994bdc09b7dd64f8c3d074ec6c8335c2622fdb91b0b72103ebc41282824fc7
z7e0b0520a3e70f59e78181be5639d0c63344e8798a21792df55e744f6c1cf435496bf90d30b87c
zd9e1c33286116e72c7dbd20ad1dceaf05f034ae59193260f3deec7e79a27dbb750d34b167ab013
zc792929355eefd8910d5959053a041e79e938c66c960bbd6ad5c980b083dc8dd21505ce450f8c9
z021892756cfb3c79c616796768fa6463336c3198d90f4ee0fab7a0b037fbeed1d55e6a1c71d46d
zcf4f575eec3d73afbec1a0643b3784e83bdd106fbdbfd5a8cb20e083be19a38eceeb758dc594c0
z2ffee0ca8190f2c3a022ee090c84c99aacfbcb3107fb637072b350e04d91e74de6b26c0397433a
zc3762fe06ee25001abff7a6296ca528622ee41916e6b7e88833c2de636952ab1796957ee6e5920
z85f336fa320258c502c3cd5a6d8de01c001db2d1d67a3012b76a58d67b941cff949f93645dcd83
z40e226424654b5456a3e4585265320d90bab98eddd6e8d4217439ef7db0995f41a680262039541
ze3f07f4d97e7dd30d0fa1703bdd88395259bc65afbe28105e393cb89da7cf43594f38d26437a1c
z002e7d3acfa0df4f77b7f194e1e0c3dcf8cdf47594a0fd3e3b667ac5865b583643b37c42e48655
z04d73e51f2cb8c7e4829e71485f4950e4fe3101ef1992da251016d374f0726e3efd1852b3614a1
z8b2ebff0360531cbdfdb9d5309719797ebab5a093c72430bbd1bb9a0ea7a2e93bb0e37de7d92d2
zecc966c68b09974dbd5a67986534fe88ffa2083bd99e078caa71f1e8fa29b9cf4d1ea4e0526a04
z0ed344146845f256520e116bb7e83bf8da31f06584c5cc9eec115b86f473dedf8699b225084b44
z0fae72386c9f7f8dc787171071cefa5813a35a45627ab4d70e6f8afa4571d2a194462f73b150a3
z7b5d3c3e0c116b8cdc6e0f0d7748ecc80f19638738420450f4a08f629f742aac73c8dfa8b465e6
zc2ee6474a89b552ccd2215c3fe20acc46af7a3fa798e8b0f078e78753d8aebb172aea866e61901
z19128b79a3d14eb5b2e4385a4019b167f87d04c9358bd2ffb9b869a657e736d355ff4ca0cefc1e
z963bc26585d633914d8c3ac589cef8eb45662ac37ed27e5ca5ddd96dddcad191923bcd3aae7e9f
ze7ed3ae1c88c5a6752886b088c9b21a538c2451853857963162b0d51a6e84afd4ff6e97ec52045
z4d52359c3145b6a5b601f57c4aee734b8079f8cfbae619c0a27420473dd4258b6e12b673d6b489
zef49c5593902cdb7e8d3c3eaa5a9648fd13fd0398cb0cdb7fe8ccf2b1ed38c32402c47bb7f4abe
z878013180803a5175d4252ace15aa8f462ec0336de488f861483802598a283b6e2b9834729d1d5
zd609fb408cf6a68bc7b1f0533a8f95d8f0b13924fb5b231a98892ef2a5a7e85679c4f47b7eda5a
z2bd75ca725d2c61e9503aa5be3d94a8b70f7d84c5179337b8811e9d4c917dd5e68e25df39875a3
z1ce2028c5e65d02796c86700f2afc70fb8c8ddbedeb8e451be20be4e6b9e1b00452506cad3d877
z32e51d9b43844e17c1054385769529fe26486daf9229288ca1b14c4ff4db4b22d6cb8f27b33a54
ze881ca64de6cdfc206b4246b1a3e6fbc2804f215bc5eb3020901aac6a45c50431a9b78ef3fc55e
z4e92d43f98890285a8c0b79cbeac90885d1463c2068e726998ca0717ad1e083b03833c218474af
z33ac13452d190ad09309c5121998dd1b0ab19cc44a22f211ded19ddfa56b99f97a825a16c6d34e
z9b2672e4de7f8dfdfa12dc691f3a28fb91503b60eeef690fcf1b7ae3c5dded745b5580729261c6
z84bc6a16ae9a1518de3f3966d564c209307fef0025e1141456d03d97a941090e2d85c66e6df56d
z63d810491dd768f0123988aaa7233df5b256f2e94c711fadae8794b951da963d7500041b6e1773
z925d005615b6b25ab7dfb37ec3825a27e4f449df371d575b688849f7ed7bdb7f41842acecf5e97
z10684f2c8e484713e33122c238209eab7fbbb5324e7e7642faed8cf898f6d6296c483c2eb99350
z705a73157d3cb21fc0b84bac1e84bfaf109db53b0dfbbd92e90660af30db2b70c937ec3bf62ffa
z95d16299e3344fcd7a58008cfab374e7848c7d15047fe3ca4d4d999b2eacbc33af50649d505072
z7b4130dce9b969d152d8e07df47c4951365d0fe022d1397ed17a5efb913b1fd2887e0bf960e2e7
z0a42419523035fea5b60453444c0f88a731c529b6fc8f670b0748fabf883e3f7b5f114002e5f25
z9382598033d7685cce2b7e1b8e4a3cee57fa9346a04d84a157d7c507047ff351caa26126afacf6
ze85b3f795f355edaddc31718e8b477465d87b3b7cf62c87a54c6719f7a542ca688e5a03987187b
z397869d9ef685eff9c08482403ec86a46e2a4f38311cbd2a9359c9b5a3772bb841aac63b9b2c81
z0acbe0da717e6c87e3c240c853b2e152dbbe8e02e05d61f919ecf1c11299f55f98d507232dca38
z773a617c4123f589ba322408f8c9f8255969a1c081e5607db0e0eeca1d3c9b5170a8be87f18e0d
z254b9e9dcf6662e8a870e29e8062a0968967329dd7990e426b82ef1e3500bc56517e7fe33af2fb
z414336a702adf1514b7bdfb1bd7986b15c99cdd42ea57e5e9700c62eb23c4bd16eaf9d9e254a0f
z2f1e00acd5a8c2f44c8c6cd7db5924f6c38c48220619f4093d2a68b400f3fdbe053ab8b236c24b
zc35a905debeba8e399306f0dee912db17e4b1dfa3397d2b916c4b788c081d3ccbb994f6b2968de
zff206612ef14ff89f4284e434c2add0bbb562fe73e3233f46141137cd5d37e9cc55519fc9d7297
z28ff05566c1b19a53040ae38ad36d71724059f9a346932d21f055954b7faff9467f4cc0a9c4809
z0ed3d2a956235d5a7f4f125695065e392969c9cf4dc663e2dc2fb8fb105d86babf7affe783d45f
z7d6129ed1cf21c1c1c9a7f42039030013e4d2e3fce25552f4a12e4e46b427ebcc32ee1f33cd0e4
z8b85d010a9bfc71f1c83ca951d62a0db68475882ccde415dc5df40d7f77fd2f8d789954445f2e7
z5e68d676bf38ef42a3de4c1098ca27715cd18c0bc88b26ac5c7c1b74eb8a0d70d98ae8538ad79f
zf99a2c878313d71ad1b755ba61c18ef2bc53eabbcd503d7ad85df562136d21631183abf6e7fc4d
z37fff4999d78c2107a06d5e7c4346e44b3a55aab1c9a0fb3e38f11fa365464dc38b8fe3b615005
z9be75c5fdb6c3ba8b422373611ad6349ceb819ba1d6b5138f93e279ae41ec0e5038abd2e10420f
z4760d1b71d53bb10e795e31f45cce770c980e082fc6592ef6d61e83b875eedc2e33c71fe44a172
ze0885441744166115b1a954ac89a44fb39e17b4c9f4efb2b521bf14001e024c8d6dc55e02b02fe
z7fe2cb04799c21172cfd0b2643dc1c6d325befddc333015d5473c0ff81fcfe430b84e04eff8811
zf5a21ecb81bf395522d7a63fff65e34e513f2cd1153f5df912ed0924f02fc634c3060efd60fc14
z3467870d41733d4da1db9831c248888d25e9dce56e51aba6dfc32347dbfedf55e983b58bedb7da
zb567d217ecd3aea2e87977ed2e61a6299063d914e5106854d96f433f6a5df61cf6cf72e5d7b7ed
zb38483fbc5cdcfed9f18c1727315e27cf0e7830a09d3058fb3fb36378f812cd7a8a5ac52b1444a
zccf149396bbfd5ba3eeabc594f479377aeda9805789213dc6f74d88a267888e675bc7e2276f1e6
ze19ef7acab0c5c8d7332bb5111bb94c993b97922c20bc6c2307e898e3c9695c5e56e155065774a
z4ba0ef22105f527fa6a70b7e2e2773dd786505179b97a538476aea13796889fb49f7396d3c5fe2
za6234af2d4e41da143558b3adc61510dcebadee220e8aec740d893c7888811eeae5f791a1dcbdc
z320229ed0edc299e699f7689493ab566ff6e52c9eacd3d1fe1c758d9a03d66fd335722bb63ddde
za72e5a45b422ed6541dab6e2bf7c84158e9a312dc3ad84a494c512f9852f52ec480d0c203354ad
z14babd480af4df552e47b1b0de5ebc4b88e0873fae805461f119017f51ee4ce4049473c81e22d5
zdebb672ab020e66785d25c9bbaeed0704bdb733a35fb94d4350fcd83cf96dff866725007e4e7ea
z841b3128821e445f6ad2016b012c73dd8106bf114eea987ee5ce2c38c69a05f369b0ddb7e958e6
zb35ff31bd05acaf4544693ce6ba50784abb9e16d1bd33b0ac1ca04c99a7a79a6ac26ef85bd8df8
z00c0fe8ad5b13f90580ee6b0231c7121ad413b91facdfe280fa620b6dba8dc75e4ba99bd9123f7
z75a5b3d4bb3727a0f60e4023e3ac1e3cd8bf5985f9551b4ea57f532ac0f6068aa6b3e4cc43d4d1
z78a0ee10fb02b59f640cdb8f550199bc5a194f844a96065e0589f9eb6ae90ced2596796e5107ac
z0f448dce92473e3c62fb231a60359a7f18c17f469d22e5310ef28a78898b2e97afc7f7e9d4b4b3
z7846c2e94199e95b541296ea8d45784badc7bab9d0c09b4d76a533c686964817c52b2e9f0cad30
z28a851b20c25607ba269442b50145876087e8aa7fcd51e1f174b17f35770ea8b79fefb6cf79885
z5dd2d859fba8ea5fa9bd4ecd19f38296c5fcd7ad8d4851ff0914e14893d88f5db6aa20a08d7060
z6c95c2245a124462083a00457e482ddb5e88bcc582b9e28e794f7000d7bbd7483204aa0c7d1043
z3995a8245b3950306cb8d6e23866e07335ed777fb78b8e73f1c1815b3a9de7970c362a1d5aeab5
zbae4cf8eb36de77eb41549f3db2dd970d3aafb55b503dda6e739fd21dc3ded817d69a179b557c3
zfee2fd769076063e47d4a79a03c08b09d0e76bb299c08c326943ebc6e21d283581fd055f0bacac
z19241bdf5fa8189a6443dc70796df28f52d58509872cf092a9284ac2a93679907b05603fa7a82a
z78ae88a61274a0a12a3309d308009978640b567c83557e5d231027d8e11ea9bf012e50a2bb8819
z6bf34592596e06019daaf47d92a3dfd91bf0439c07a3d2858d9b280cc0b5b622f791b228112a31
z63c66fcbefa884d3415e91300f38cca8afb9114ca6ba39be0c5cf081b9b4255abc6b63b1d5b540
zdefd668033fc64131670dbccfaf8a2c1890427a0c08b916ea640cdc37c4b1c0cee0412072af4e4
za337067bf1762ec69f72a4b15f15c63fa56d1c8bb5ddac04cda9560ccbfcd22c4a9ff6e81ceb41
z3030c39506545d543589f40e30e507357496ba12f65809e301968bfd56142f94255b9a27b57352
z74eafdda0e410a9136614ae846c36f023961fe1a6e1ba841878d66865e47bbc02bfea56b179a6c
z68e463795fbbba7b60c5101afc9c66a92252b7905c59492e08168c5d095e3cadfa6808d1f3c2b4
z298a9fafc1fb306af9b20bdd67e331e49e1ad9b5bc5faef478a49ae1c2631ce2a3d7aec100ac59
z060eeea2c55cba7738d17cd67732b465b59307d9f84ed05b5c638c9ff28ff5e5d71f083e85ec99
z7fc009240143ca0cad2a216fbdf076fde7cf306b9832f3ccc7d9515a5890e745d3268fe0869b94
z79087f9207eb3ad74a554fc49e7f300538a7cf4a772d82b462d682c3e7f404e5002ef15836e880
z62461670c5efbcaadfbe5f2e7cf8c357ffe1e552ca62691c10d367eb64089b3cc8d4842e85241f
zecbda0ac9bdbd4cf864f3f01bf113c817ebd06f14f1c69c161718d7558279140e5a811a22437ae
zee51649712de71316e81a2561c38af1cea6e2d84ddcd0f6c72287b89ac026d0b713038614c4f17
z43752ba1e0ac79d2d750b6e9f0139d31304d3f8e993e5a5bbcd3be55d35a6fc9ad86313097b809
z278fcc183298c0fd388b02c5b1b56eca8ee3aa2363dd33ff1be7cf70044081fa03f678e1d17b7f
zc9da2f7d034aa3b6d7da7597f8dc60057faee9ea7c50f65063189b0f609e6b3ef343e278cce14b
zb6cf2651447bd3f30a01a98a1f500bd617d7e9e3474d2b412329b5b556e2965bf4eb24aa84ae3d
za7c91005f8803f9146cb60e03421e3de3a0d2b6f6b2040288de63914f03513df64be6a7926216b
zf71a6388b27479487c53550db4cee1bb644a6fbff326b08a5bb9f2101de1f7e91e70a25e8eb741
z09e53ceff570ae5d403e12c8c90a4b9b437490adc319a1b6f383e730bfd02fe2dbb107347ca400
z203490130404957692aeda328308ff8aadc603c93651d9e55614cf67b38486e3e71f5002ba1f3e
z70d5277b8b73b0abe2ebaaac2b7831341a4b78b4c9ccd5c9c06b71faac286095e56155450dd147
z984e7c1ca48d8e43bad87997b7a38d2ffcf7291b1651c75a29895c478af1e01217564e25fb38c2
z35cb87cc0108c859bd0f785ffa940d1325fafe43acc1feae3cc49b29b9bc0d81edbb45c31e4f45
zb433bc28d416f7b2c94a01ba3fdd61868de479fbf2be6f0bf647fec5196f9ab20592c89e7e7272
z55f9f652bd3a31ff51f95b233b1c317a7ea80430b9ba5682f6e62f518767ebadd4777743ae8a39
z36ead5a0453c8786a3e231a8bc68957ea73d92e670c6defba80f24fa49a9a5bde989c4aea6e4d7
z7f77f3347c1942749473d45cbff5012e78926d701748e6e9d23eb6034a8d4c7c7263bbb7b10c10
z92babbeaa022d0d8e2e48333207e9e27d38a699f8655745ba1e41d6ecfbcd9379aad976eebe8df
z9d1b7d06c426c69c4e950da96f62936f5780480bdcab9b44a0d12c7cd07ccb388c308213554b56
zf9c8c3fb46d811f38d406ebbdc95a0cc544bc54ff1dbc658a83bd934b52e7c3e12eead0e9ca025
z565bfbf90b81a555177a282aac41a259e0c7a02c85135a436e01d4e663f45938bcbb6b00c0bb2d
za5540eafd9743b2ee4dfafded27cba684f09e1a809482b051ea809a5875ed234e83dae5c54fc1b
ze771ed69de0580ebc9ec76850d340ba54acd8345c7bb61bb80523ec0d00fc64eb24246b1974389
zbec9d4230bcd20a977bed7ea3ccccd520f0adab8616998824e71df8b669d71f9dc75c0b3d5e238
za9525b42296c916ba708ce595e6e8799d8fd50b621f5296740afe2fc81f57794739f2de3217445
z806e3d6ffb9caa011175e890acba231ba1d95026d207ee3de74b3a95048f8390156ccec32f85e8
zc04130899d280db3ba4040fd309306edf21c3d3dda1cab650793905748ced20bd2e9c6b4256e30
za3a8e49beadf58eef233a85530ae76d187496686fc546e10d155124aa867011d1a4e66f3fba698
zb53757760153be70da537638159fd22bf15e8c67490b93f2ad9d7b292d4fe31616f99999db7202
zddc7c448c21646dcc99fa07dbc466faeec3906723ec7b6efb0cdf1aaf0b6184fdc3671fb798e86
zb1801f46553e3ab187fefe2641f2aebfd6cbc064143e8600effffd885a46e7621b758447357c9b
z655d55dfdd3b749c7e784898e5ab15613107433c837d95e454f7682b7625ea579567978c66ec62
zdab380160a87add41226ed3592e2214d4634b446bffb78048e78eff1192ce2af33c3edabf74002
z195c5db9c1e51f5dd93838eb648444f2bfd235b609496e80689bb19d67aa4d589404b1388b793f
z6a570c8cee00fb77669d09d4a1c533628235df4d1b75f9a56854d7b1755f1197ba363a6bc94f86
z1598f2cd60f5f04140322be1cd74928bd18d3ff90f31c59ce891119bbd0d54ce69617bb30690ce
z9cf11d3e88297772a4dd925dada540fc73ec010dd9e6a0b5fdb037221db035e4e56d6b784de8ca
z533966c287e95b38b1e1f87176f5ec036a25efd2de36152193b7765f6d9224fda1177106331a3b
z77fafd3beb6d2c0d86691438f62e9288179b73c2b6c6d3e69b444ae2d171c97960ab0fd060ad21
ze0d688ba1593199a6f9b2aba09811723eaf75ad55d6062a62aa427af1c8a03a30f04ecf9464124
z7cb94e1c3c788e384904c2236d93aa4d4e6f0f3c9a9f47f6ba7fa5c1a98ef1a19730f08b1d3ce2
z313cbdb077c705a703a783bfb72b407b93681141872eb8ae11047ffa8ffa6976baf4c11c24d61c
z57b7fec18600f2681eea3a97052aef56bbbb000d2b113834bcfaa1c7a4cdcfba21e527f1126058
za369ca48938b960db399faae7334e197d3563a93650bc19061cc35bd570831d9d6d3a494152f99
ze8fd4d58434c25f55315be6d711c06ffebe0596806cf7f0a9e59288a9ac512baad7ab4db0551b1
z478810be47e24cfa600e02756a5cbd05ca9d2020728e12a7285d2d60a3aec5cca706c392dda17b
zf7176920fdab6bcabcd227c8a9f580373c91acd7bde8666e7b8506c352cebd2318c7dbdef5274e
z6a9edb56f4a2ed929972146d1c40a5b81bdd9728657c39cf7be76677793453723609d1a421e943
zcc37cd6ba794f087cfa0f4a982d1194e6a78ef9f5be4f8f082051396c9ae67df6a0b886fe107f2
z70f0c6e408b90101e456ff8fe3386bc57d4877417da4ab6752f01806d065391bd048c2a01fddd9
zb28624e676929e67ffc2d8d6e4c9508faa74c77da9c93945ff4e50586b4c4eab55f5d26635c45b
z89ddb5d59b77972d1a4466f3ff440ee2d56aa58390ceaeb4d6cc41d7436f38de481dada8c91e64
z9dec8181c963d271dc7b2b222d6c51d91bde0f4ff9b63eced4ff32b732c7f1e5e6c907d426c4a4
z58ff5f8f5334c16679c2a990e72e784e7eb8924f8dc7f35cb7133f540b484ee07a3f322a48b0ec
z1291ab5ed3c967ea49b990d8f2db75d52492742f13d1b59d10d8b04d696e2f55fa5a32b1383b3a
za9021a6f510536799ff9cd0309905ba13cd055ba22e032d9a2d3d768ba46e9c185ad5ee60fc37b
z8dc10b66a60468f9e132fbf8cc30f7c5bafab371ef0f1d69d9c8e9c32036f874ff1e797568c9cc
z67e09d272d4ed03288d449e725d65dccbda1fa97e7ad8105d31d77e2fb55982d3cb58b0447caa6
z1b8b96a1d71c9218dfd26720670357dba9d5a305b21b7ac47169679ef637ad17fd8302f981c63a
z4b811e1a98ef9c54791eb2299ccc97580d0c48a143dc2c8d3f334503ae67d6882dde50a1acb7b5
z280287c5d69d8d3a78f618f0caf7c01c544a0e60abece7bb90868007ef2b7d6510a78717ac12ec
z811db890d9c8c566d8bb6d2813f75c24cacc79f9b24ec397b18cd57fd41f820aa475d2b3e4607f
z258de4753fc4922489da6a55a0014faeac6ba71d5357de35025f5fdc152fd8d50f548e8239f36d
z85b9d47b3ee7ae88442aff3f7f4c09b8de17140b1c004759106fb5df85dc43486cbfd19f1b2877
za5791fd94223ca2d0424e4c0c9590d4993d08cbed48ac5106b75dc0f4455fcd9718f62637aa287
za44eaa10044d9a1b4188bb773f2f35de962349be2c9ce9a49f4005519a1f1e1c01e4f575bdb9e8
z56096131319881e10d95166a508fa4f13badd654303e4c8d6f3c69906632803da450b16b16cd95
z2262b6dfc8cee4b61450edc46480a8ce9d36316ed268dee069e6894a0d8f811f957672437a11da
z37709984cfe801c159bd983a5b318fa0242b1862c48ce9f48093082d99db0177e325503b3fc423
zc8b93b6b772ae797482366da71fcc4c3b413d03781b3d1950ff3a95d3c4529e8b73cc5a18fad48
z5d1dbca5d1dcc343b734b085e99d01af2dfc659c5fc232f194c58e3501529e9dcece7c89e1deba
zdeff8bf0ceb95fed6314903ded8d36d39b1019245e88528b4595a16dd5ba3648e8949e6b22d91f
zeb54ae8b36e4cd14d16d8acd56aeb90a5f421f47e2d29e088c12394aa11e954c8875df1b0025a1
zdf8614173c69d247ab396c9ab205ec623492bc1dec5b7ec541d21208d42d132a05094acbb32042
z649fd3e54200e4a4545729feac647213ce16c5fa1704bb9280a99a54dd120f500fdd35588ba0e7
z80328a5e35474a8a6ecf763c7bdf8e46f6dcb5105d5e234655596bd184fe15dc2d37c807159d85
z06951e0b1d49fe21224a10e9fbc0db7c86b77720c98913278a9ec70d990078cd779ed7596b196e
ze0c791c9db8117b11e2fe4090d48ae41cd714fa5bb1a7fc73a4470d5a2cc1fca0494e4e4c83965
z298ffc2cd29744fc6f99e5a7477c9469e90b9e3fd4d9bc62c341e64105565b00e7d3145d10665a
zb2dd95175ad220ed605f68b1f1d52969fa3dc575b711e5498c31ead6e5b730285b4dd5a51e14c0
z710f985b423e4496877e17462a21c40587c2be631a262c38f8f1b9d0a9c90f472005655e566196
z73c8937e0fdb4a423f7fae863d4775d9aa9a6c6f70c0aab6a84974cb0aa039f635f0d4abeb06b2
z3c757051be83bc57be73a61865b71b0cc6b1144bc165d4232eb211072618997058ceb5d128b9d6
z46bd71ee05ea92b7bc567274a730087cf89450d6faeedf36ac08ca13a10b1016bd284dc745e207
zbf53e8d2f3edf7ddeffb885a31d18619790473a0ffacd187a67b887f2ec8c88a19eb5ac6673840
z508b4929c473781415110081a9f65a64ba5b707a17f0a444351dc9403e4d54ae860d1657a71bbe
z2c2f1b2a733a9c95d759fbcf97308173a6e62c8daaae14868c28ba3373856798931535ecb8739e
z69daa78bfc38e97a09fba9411bc21ddcce949f46c5bf63c205964fa89d5b97fea8cd61c2ff3656
zcd8a4eae6736a901493321d43e2dd741f33e2ad0a814108749978f675761b569bca3a63a882413
z01c5de7c627c412e623ec51c03014c7477c45e2262d2772a4e3582f407e9a8bb045fcf2379ecff
zc8abf38e956693dd1e55cb04abf5b94ab0386aca44259d8a5b5da3ee7718b0b6cb5f7c77f7d7b2
z78738b59ccfe05a3ff4319a810c1db68a9c25965b30e41bb461700dd17f2a52fb2b1e70c092675
z4920a1f2c1f565bc300b9760d5e3a12c1a0edd6b2ab4cce6d2ec838082b3122d3a0f08e1247518
ze257c7e15a518555a62df3e441c968fc3e0182cc0ca9b1b475e390e1ced9779bf630fa227ca86e
zcefa4f5c9e6efe22783387580a7fb2180020142a5141f3ec9b7256ef8f11bfe5b2b24b7278fc4a
z319a6383117b39db5c01f205d4ae32b94bff83fd530410f8f606878d94611613274d393624e5ae
z31d65de5503004ca71dddd7903fc120037f7a8fc8bfc93191550312979ec8dbbdd757007d16394
z62ecb320e378134e74d1cc6e53351c7ccb34422e7816fa5d8c31858e387e206b4ae05676f25094
zf8872b39f5769b352f2594cd534da7b1a9059c20679517e6b293c7024fb1b5c5baff252e58d0d3
z949a6e0f247fd4b422431481e0a8b8dee2328188360aaa3b9f9d5301356d72a6f8e985498d969b
z89f4b5ef1f4eda6402710431c611ab8d0035a518ecba1e5167b1fad6a2e85113ba85d677218607
z7167a494481ca641ef6f9dc15bbf21af8a9471b33c0095b882a3b69fdc1a8a4a837d2bb15cc2c6
ze88c19ce873a6a1827e524759fe219e2e148ed63a5add5662aaaba71fe63c454242b2c9152dd14
zf4af88742d6aeae2ea354ad698b67d390f6ce56b39ddf8c47e10f4087387b37394fdb27c732f17
z8ad165d761db7d55df19d3ca1bc8faa57f2a4674e715eb259d600f39ded0b1f98d80343b782c23
z02f6d5f1f207fa40b4c6d21907de5dc1cdcaa373d008bc941ddfa7af506bead44c3d4fdeb489af
zafd34eba856947de033ab341b9079231de05c980857d46ddfd504fb46d6f4cacbd147e007489ba
z0c57af12c6ddf1b0d44f7fa6eac1bae8521d012c1f8e6faf0768f92b5fc6317ba6708fba04807c
zc3ed5ae988575a483a26fac3dc2c8d63babb02ec8e050950b3c3bdca8f7463183a823650c0862b
z1f34a655b11842b7b83952ad4940483d1ace1741ca3e12bb97ddbe3e7262b672454e2673957c5c
z706673e1bd352cc1aada15de9db402d9987749d66223a0bdbaae72438b48544fdb7094130b2730
z61ab39d4b387b7ad8520a1560eeb2faafb4498b969f5ddfab6a462db1946453560e409db4761ba
z55a203599af37b9c01fe0c7dad19b6424a9242aece6e6966eb7a26c1500116bb703edc535fa98e
z55bff11b31bf48baac67dd92f13a0f60df3b12a67259e6ed7edbc23c3a181b35e5052da28ee68c
z127fcc147013499b868d809ef097422be8cde8808563684a3c8aa4fc2bb8dd80e65a5eaccea966
zb7897744fee32dbfe2a487ab954ec7801802b5ad4c0f708571c848ef6715ccaeb9e41f0e4745ff
zca3522aef862164573e8cb19a8cb42dbf4aa756a773561c6eaaa67c6ca228e6466cea8963d6f93
zfd14707ed387924b96f280f1ef1d6dab09ba6d8172c68cb27f5bae483fbf523533f4b7ec450396
z614ddc3b292aab352dd1ac19c20d139391230b4d9b8b80e07612daf5511f8755c108e31a8b74be
z69260576be46903745577c0d8aeea224fb88ccbbd9073352493e5900c6fcef2345bad80ed55716
za88c35f46907547e52c8ed62479796f4146189e0a1797f5d092b451bb99b87318f4442ae2ad9be
z4b7f21c5750c1e3200e4828665ea3b6f104707272f21a2477ce36513efb6eec77cc75d18c4816f
zf4c608f55deaae145959833d9cf34c054c96ab8ef3c9ea64a52ec07b50b1c7366d7bef6d02b456
z27e6cc7e8cc6d372e66343abe31a92742f38e038ecd81316a084fd96975868ce7ca4372949fd7e
z9842433dc2e1f95c2b09ad4904c857e89cd9c7d611887d8e88c21516bc9d417c520da347227b70
za294aba7fea3ec3e860b925dcb398310f4ca3c32c8d7716632d99da9ef817e9576fcd62fad2c2d
zc80009759414987ce947c00e39fd8bb77e8ee1dba152987fa67bc9e56e0d250ef3e0533fa9b910
z14f5ad52f06f7ffaee3f777f50d8b7f317363b4ae04c0beb7a4d4692bcb694b9d25adcbe947147
z9f597f83fb1a81a811418a42176b47a04a021735aab45f23837a3b9d4317c73d45b0303d20eedf
z287da2e9407f2777e52f8e435558f63ad2a08c986ec4bdfc758e969f6c5f57aefe91ad96573fa7
z2d16d49f3f2dc0c0edb5ac36905f11923ae48406aad3acb184c9cdde29b04e2aa6a588f78d71c2
z44cbf246df4f9dbb2be15743ae47c3fb4c461b001f7d18bc8b789b589cda20ceaa6ef708fbaec3
ze7e6ceb09ea49b427340f490d776afd9abbb8dd7ce5bb1ef262e37b83f285cf9f3f8710a1d4f00
z830bc03466331d247a4ea9edde2f5276de042751284fa249b97409e7d19dc3b729bfe4b70608bb
z70a8ed775c4405a3bcc31ed1505c62155d1d1fea1eded6e90435159062a337e95fe4a2613ac702
zed2e3e4d77f293d8cad11a022550ff0e40bbba3c7bff6d5b0e21dc84b410adf0258e02bc51fe14
z3dbc7f345729b77d61017b794d1bbea6b5e61ba03e66a8f467bd88ec49ecb82e32a2da4d9f56f1
zd0ece66cfc9638145d958f76be496eadb3f1c74e5b1d9350c40cf18262b613e9a5a04e6054f9be
z889db825bc77fd89afc9d34b5537cdbcc3450db25d8798950e6aa5525150faf8648177568029d5
za02fdee5c7823585995900a1eb26d3a61d4ab4178ac875ef7d8ab2e3c58df8d8fedff45693bdfd
zc5ea3447de61817a7897f9b9d603ec0df54223c2c4db56d581941b86fe50fdd074a044cf9fc3ea
z03f489092ac5d18bb421a8139f6b55f627c71f5d7929dce5873a1b1d8473fd0a1047ab9be6ca11
z642cbfef9949ccb333dade87ba2013036b1842f6a92c0eb5132ed15b15b58e50c0a3eacd56bf29
z88ee901540a2b73f043b74f51aa641d9716cd72341bdda09f710781976178afb406c765099d398
z05e3955a3cf84abc03b5c9076bed7ec261ea3b934c82e7aaf78a4bf4ec3354c41ebcfd0fb4a62c
z8f7e589803cc1bf1575f8b87510290403d2b579fd0487d842421273277d070062108ed827be45a
zcc9517a39f3388e67d060b2f4d56567862a5a170dd6ba4febf8496932150eb765e0f9c8d252226
z1103b02fee30abe84e658574d83d86c6603fd6c7938591c91f88abc80c2002a617fd2f59dd9bac
z2f558df0c2adb09477afb4067cdb77174921d320d605daba538ae8acb34f42d8dcf35db6fe2d1b
za5cba454a0eded9bf1709ee8afc7f967da6ca60ed93b34c336ff7f895f606aea159ee032aab9c2
z2f55f21998ca5f9312360fb17ecac8b58651bf7d0be8495f23407b85fa1c2d998ede12b473fbcd
z8bf05e3aab98c2efac0022f31a33c6293840a2d125509b381d26214a16027073786c11cf55228a
zdbd76052a0a08f9aa3f7f7aa156c64b1279b8b2f4852b3f364083230bdafebcd55b85405665424
zb84e20573e925d77ab7bfad165c7ad013240ddc57411dfc33e318fbfb140a56c183fc8946faf7a
z1c20fb15e42169c8e2b7509176e05715dc60bb2bd5089ca727768552b2ac8c879a8f8c75243218
zbbd99d4fe7b1e897ac67287f6c644e8cbc7faf769f846a2ce1d974ea047bedf5a7898d33b005b0
zfe02391f8d7152d487044b4ec06ac8fe5a14e7ea0fffe9c90e580e4391b08bf3abc0fe4287fe89
z6487c1804158feffe89a9e26c96b91e4c48ba379783e23b7c0963733e82463296bac8fc1cddff5
z3867002a954daa648be5d27a7b43aac3ff6661fa5d3f9cc2c35094cd6d2e36c0a36d5799dc7959
z1da9d0d94a152949553a3f8ad8a8947dcdcf0fb37bab368f0d1271f10fa361ffd9b501b50329ae
z38dd7ee9bacca12aea3fbe238189f7274cd7a321a329c21d64e1800b281b898548600a8943eb45
z6c5006e66273d9666aff80b57bb3e822c70aa87d23859728e2d89327c8555e51a33266dcf574a5
zbc9dd31f8a4f8b73a18138c9887c090b99f765aa359c34fd6737dcc4808c5afa9c29df8eae9796
za4f0523aae94459cf506369a49827437f574925b06150301fb3eb57f603d2074693a8c0cb7c35c
z1adefbabeaf4ee2522afd8d48e82cb1029ee1ba8a88ceaf47e905f657d6bb41f1f33e0f5b95150
zd82c635bff0aa6ee68b2a7f109b46bcc3c5560d3656774244aab0a4d1e31b84083ab1bab2f561c
z7113e74aaa8b1375297aa50c03f0ea85cf04105b3358b3404f6d035db79a5d8e312570cbc41565
za32b43c640c8234c4890df6bf03c70f69c3256ae02bcbfaa681304a956f7a972082e7f8826bbaa
z32741964431a891bacb854ddbea78d630bf13cfcead29b7452db2a7bff46fdd87099e3269ffbfd
zf96e5a6d8c84a423802e0725df472ea52dda14af5f199838e219b5a2a900efa11579ac6b39465b
z300d1779e2b7c8e551e4fc0577fbfd8d46e1db3d718ff9ee97aafb302267985072b12eb71f951c
z14ca78bb5090021a8223219c42720094eaf8c7c3345723748bc3e70a719d4e0c39fcec94311c60
z761f4f82dda766d4831167e3478ddfc8f8a49f428d68d05adcb7fb642e61f947257326a34a7ae8
z52d53d9200b3a10de905c8b829c1cad4634ba24a067e65dbe868bac746b87c44dc71d0fc7d9306
z4d8fbf6533b496bde88937e5b6f80695e935bd99e744464ae2285b226d7b4434803f8edb2d250c
zc7e60565e1cf0fab2aa4acb71e2a01c1903099093160635ab4200cd2d8a66b853e0f6bb6204483
zfea60151819ae28957fa64524251bfb30755751198c47a2587bbc005cd0fdac00bed89c3827a9c
z77542b4b518275dadd0c8744d9f902671feed7ca205cd366ec6237b792e2e95c38a44cb01ca541
zf2792f01a43f57173233558b26de5dcbe3588fd823681ba6284fdcf37f4f6ac6e313f8ccaae3f4
z48b781d6f49294c12e62b74495ef900f5285a9b3f03b85210a81ba64d24c9311bba20e13b8b4c1
z4084e66f6405c1918e65bd116bd4fcd8fc3588b6891434255490a2aa629620762c5fcb0add81a3
z2e43098a899457671a133d04e434868827e16f74a2381e04007a58170d9d323b4f844ac285b6d7
z82644e72fb50064d38667f92a95a1703c9699b4d10eb09d8274eee785dae1a8356b04526d5b1c8
z6554e1b4febc4b97619aba9110e3d2d2ad6a311adc75d43bd9f71b2468ae7aa641a3db3465a675
z6f44f510ed2fbb4ace47034ebb445bce9a1c8a88633da0f7fbd09bdc8de1bdcc425e0c58a19807
zf5bf876ef1739ee89a05cda124afca12642f239a95c76459b6a1d0541061a67fcfacd686437920
zf7f726a2b92178ee30ccff12c9202f9c4e066f404aec33a2c618c24fa87857d6573ce6e9cffd7c
z1bc432e43900d2fcc74ec1e5ae29d34c4fc6d9afbc3e6fa87ba2b298bd838f461bc8b86962c297
zb68ef0c9aacaf172f4f301ed9dd22380834b4500571b204ba39818e1b40cd33d618c79e3e500c2
z97af7248f1095b48256c309fb5e77c7e05ecf87ffdc3943411b13ff16f9c443765e6e3d56338ce
z520bfa69f40267852549807261e7b9a242a53a2e4b95902926940eb02526dd764bcff34e2907ed
zd627d9b50b70bbbb31fea9e2b0fcc562069f2af860b2e61ea9888504d1c675f1fb0994dabbb698
zcab6712a82df2293db3cf4a6d5c78a272c1cb01cc3446bb42f2cd2633e8339dec97d021520d0d0
z2957dd90173d3c5c6191ea045a230bf90a3beb9be38bab319dd3557ff431057bbf2da7fe62882d
z564fee706f6bbdf7aa6e2b70b809b22f0be99942adb1c1f687207613319ab2b4f3ecec272033aa
z9807431bb5ef226b67294a63d72c074962a6df0e710e8bd168d7a99182a4e0da93587d4bf0a4b4
z873c8b4ccee74ae5ba8e721e02da19b578e1838d95b260e7d28fe3b74c707d0bbf6307c69fdb98
z535ae4d608bab7841e84885abe8a9f1eb9a229b508230748442f2c9ca6cad92610c81827768462
z7f498e8bb83ecafcdd1cb5db1077074c43bb82b07344991d377c70b171b0dd40a4cc2e1ded925f
z2bee4e13bdc6f94f6f9238d55b368444a63e05427ee1b61ae46dba984b437bf7f1347f159c2b5f
z705967b5b3be88af2ae4a8f378541f26fccffeaf8fd5d7931e492c58260c56ebbb4cd0838cc4c0
z62546026b9085c6a1e52b4cc76549ce80192e8a1897eac822e96f86668070fbe63b43b7ce2917d
z17201749f1f5b51d7c97f731c7c4ff4c77c5afa2ad2f60549acdfb5d324811a01073c9ddfabc6d
z9384ca0b2cdf2b442dc4ce4b1ea1492e7c13bb7a60b55b77227fb25c488de4e121c780c1820225
zeedcf3ba86ddfb6b8d83781ca5d16d279c974f448c0dd2486258c3637c51a265b9915d15cbb64f
z2e0e9f5f8f6b1994af8d4a934341c94cc3e6564de6347ce6720a06336665a1de38953caa47706d
z0ec745ce8d62c84e9622060458bad1569e1c15d4906c2779db9ca80486a734a0dc488db667719d
za441ea428ea8b538a8ef11ae2a448958b5b2794fe76aed8e86af6a5f157236ac28e222923dabd5
z06619befbec5355965d274d1b15e25e3f01dca73d3ec66ae0c14ffdfd3cc4eaafbe8bffacabee4
z43dcb67b67f70dc491bfba6100bf23edd511dcd75e07f895cdcd8429ab5eaa2b0ee33fc60815ad
zc3436c67759c60003879b7c27f68b573f8317050cedcea42b50f46a9fba2766c4ab128cfdc3c62
z218335a5e05dbcb4e34deab9587b0e66855ea4faf74ee6dfae224c5993809ce9bbf26f97216026
z6e081ddaf99798b2707fb88cf07a6368bc172ab47bf9bd367948b1a70d5510c6bd807f86adba7c
zd9c8e2bfa930de6705bce05cc85343b62df7e2ab3813a25c8f3b748fe10645e9c1830cbe5a30b9
zd5cca156e50badcad3e7630e3b4d4580aa660d0308d0e4f1b3ed7312c64cd64a4ffb6adc263f97
zb91c2f49cdde3977da7d22641c658cae37a136fbf9adb8c7ef7b5bd77827011452b703c97462ed
zea94ea1ffeebec58cac2957f69bde6d22864f1f61495800f49a4e5b836d355e86cd296a742818b
z63d709bdab16d9b618796ef37c4120caf0281e7a6bd00070b3950004638750fc34a1bab8994fb0
z261892c69bb0e9cd38ebbea88c9229782b90a35ebb6523cb614d8722019d7af9e5c83447ad2359
z4ec5478b10e79af7978f87bfc8d20d819833c0e374d08e576efaa5d84944344d4a367a6028e427
z869eded1b34442b683f91507d2490428aedf10f3ce9d449d7807ce6ebc5f9c1c24fd878d6a53dc
z9b28fe871d199ec9aaf64ba47a73414da6a52bfada7a816950d3a48b6838502dbf320d042fb15d
z96d29ff32c52743ca305344278ac1f2986cfc662b1418b1ae91eb3166161cf140e5c174499a12d
z27f6d2226ca3043551d6fdd4189af3bad6c274a5f8bb3f9432da97900d5ea4d2aaf205275491fa
z48713aa349a60ed6a9637684610faa5396cd565dd46dc916371312d4aa37e8975bb956d0231fa5
z26a0866884a7aa4777159674be7e48ad8e039301e5f3a4b2b714fdcfb3b5503dc25d9f0b8a6c96
zd4ad816ecf8cff7d56d16ba7a4e13053160e3730b065bc9c089a7927d2e5d3e5d543b5f7e54c74
z4e99886f9f06ff2f756f3f1f2694da02b7509a4e6116d3d47eda3d0fdf7bf55bcd871513a92409
z401f3f135258a470a39fd829c6af8ecb9ef5a3ff9f19c6727e4c1fd4958604c68fb9bd7b7d0cc0
zc4e4bfda479a25abae0b8613eb66f1fc59667fe32536b5c46f8f7179c85b9d8902e637ee2a16d2
z0cd54af3815ed37fb491c227f793d868ac07ba288cf4d95a73fd6ace79e018f8531a4122f11ed7
za618eb0addc2ec50da4ae42c43b34f68295d584e49eb7eccc2fc965cec19b71274f655886c77a8
za63a88470076a2fe005300f80abf0980f11f662505efb95856e9b02778febfdc62bdfbbec347dc
z16d39dc024c3ce90ed2dd0bce5fad638c29a2ce18b52d940e8968d2f94a7b3bf59da57eb44a0c9
z895bce8f135266e1f79fdac22277e043ec6eb78946bcb1045699de0640a1815fdfe387f6ac85dd
zd5b00b94594e55b063becddd3580d7ad08402ab40014ad39731632c384d000808c7bfc6fdb436c
z59487d58c14d2ee58a29a848d96891a877b993f11b8e6edbc1210cbe126a061b5ebfb03e1bf0ce
z9a163729ded60def98eca33ac27f28c8eeff5d0e668e879081fa8262471d32209800e7f04755de
zb1fecd5916bc29bf4dfbbb3799f6c288e865586ae38501798cd37be4757cef2b1d6170609f3b70
zd18d930ace70ac8910171e23688fe0f4d5d803143b1b8d8390e57b40ceb7024dae36f07b9f03b5
z2908d0afcc56016562c60e820aa43afec205b13247025211e034028608b3685d77b0bb4ac69a69
z9fb61b0f49330f881d8581b64e8676485ef98a766cbc75cd1bb818088abdd0934ceb2ed77b3fb6
zc48e8365edcbb71787e76a2ef870d6a419cd840fbb36a7c337ad5772bd960c7cc2e14c3b30d44b
z13119340f0d86993503ecbe3d841b8be109d6b65b303561a5886874a2f5e5575e41b56fa5261f4
z669818f59d51ac1157f2dbbbbb05c5dbbce2fe0839ebc76af17d5e44342b0682d639e6c50f8efa
z4b18af3f803d4fa3fc184491ebbeb2afe6a9dfe1974c063f957ed4c1f2e3ed535c657eb0814b69
z7289283abf1211f06c824eb39545696f7cba4684cf0a34eb0e7896978143b13194c8255b9b63da
zb4c32abc88b486a277f2bf29a3c0198ac9d7dd142a1e7293dfbcb739aba30988b5b7a80e8adbff
zf77030689c6a25337c186a4956c530799f0df46902bb161e8de8fd1fdb06dd6ccde4f51cef318f
za2cbd966e386fb7cddea65aae486e71ed63b66b0cf04c44ef9fc4e5a4771be9d964c96f1409428
z0f5c8b5280bc4f6f4602d19a438d9d08df94e0706c5fc2cc373520938421f46f1bca71fabae00a
z8c871ac030f571656f483750bbb7cfda5efb67768067fca654e373ac695e632b7b0de4a0e6685d
zc3865a6e3e2efa67af5014f74de3406b4508686a5741a33a28557ae9df021ab6b313fd42c1338a
zdda2ecb794c904912637c8eaab658593d187ed44e4aa5daa6b7c05d527eaa750e7b7476d94a909
z772bf78d3103046dab2125b4685119c6283b1daf499865172e0ce8648c15c4bc843376f37bae6b
zb6237861730f4379db03987e83d60b179eaf362bc029afb5bb80f4c93604e6eaf33b28bdb8f9ab
z71615bd15233ff00438da4db57a5621debd2bb376afe42f020b00197c51c79ac3f451b8406edcb
z5b7b83f20d2f5a0257cef373b7f51914a1451dc46d635d8e236d3f213c6f72ac65bfa9ea61448d
z03da97f828d566e34d484177b72a62ff237f69b2c317f9f12e5c513bfc7497f84b3766c3c28ebe
ze988732d6a826ca60f91ef05036846bb577eefbe84086e679247ca8ae291518e9b3f0902b2a7e1
z6eda35eeb589a54d623517dcf38e79a8ecf2b1da3c27c253afb9b77134380ef6263031b356e601
zff1dd9439e0c2a2e537ead654461035aa5094c50133fbdfd75e2d9963b9242702ea3160e23c15b
z711e39a799e0d24b9e9f8eef7c5138dac29de701e39a207682a7b54f27e9e99b55d8f122a90b38
z80d5036cc450fe05eda2c52095e2e2fffcc17e28184bcb0e173a6fe72116b1ff0e620afedeb6a0
z7a69e909deba67b51e96bf1d48a4ea6ba7844f4558b7c72e23539e234cca4e37e78e574534e0ff
z10375ac471d652f53754cfe8d8154b2b5c3b866ae7135496083c91c0386e353b73afe6e9d7be38
z827570084ba0f8585ec2b922c417a43c7203d8378cdd031c9f4a6866ef963fc7687a7dd0e87664
z190b56c0fe158d23caa1428b0a4f39b2aa613f69150377feeef94de438342190109432092eb1b5
z5ff960d5a9172f77d55046156aa6d072583b8db18c8da9c049abb3503c1fd21e07fd038860c97c
zcfcc87d2bc517f4420879d853d4c23f8c39b81bd44d616bbb557601d8a8c47abba364ebb1edc7b
z26a6c8760838affad06aff7224ce72747c78eb5f32b692d8a9c91887fe8c4a970f89b85cc9c7c2
z6fc8bd681f35b7c4339b1082582e11215ce83c4ba842a8cabf30c4ce0299449bb3efbb03bc4538
z24aa19e7e9c64ed87f6a7764c330e765efe24b2565f3c0e41a9d52691109319e0b35ffb50c927d
z335ff9b5c66c40ea4a6a7275cef94a27fa6a222efe501ba5b95b670dc574be052dc81b4a933804
z266951d5359de335cb1fe7d09588deead05bfdd88af91035285a2c235b87105ba16c7de1d82393
z7c16fb32313848650c6043b2cfb2d8774b5cd686520024e96309095464b3962d277cfbc612b3c6
z1de910c97ebc719788909a634b479bdd2f877e99bf9eafb2a240155b8765be3bd08f4f0a158dcc
z977c259656e0cecb558010735302893fbdfb766c9c54a28d4a9928ef5c6fc65f9ab813395391cc
z308cdf8513c4e301c23d021736d0febaeac3bb5ff3fec080a9c62705a57b007ca017ec76e561c0
ze21a0fc34e8303e9f397b6f98e539c965800a26891b898a934f1d01e5f1cc7f854c802cecfd790
z5283be8677c5162386af2a172541c5dbf3255f972bb40272c35b55772d9fb37db0ba502243116e
za8a1c715e8ba7b3eaab3052406cdf92936a8e0d98011adcdfef8ce88aa625fffe452b4cd692946
z8a3fda88754e10f48cf603b00adbee4652501fd4693199c30777d391c745e22ba3d9ac9b00716c
zad1817656bae40e99e438fbfd907b36883966c22f21f98ab7d06b702e9a875ee43dbd0c2657b50
z3ec51edb542770f9e4efa39284c235c322ab769247ccdd33fb7c5674dd277630fa2c36d307d068
zf72cfed441c4946f354935cd5497cd314b0c890c063c214332f122e4b45e5b170281fe9ff9a25e
z63c3925c14df24380a5cba31f353e7081c601fd66dc401aa07ec60ec4f0653fa2ef1c0eea78b6b
z4315e02fabd4eaf85030bc44dba008a8cf104299399e4fbf3cbcf6facdc6ec6995f1ac2e1a8ba1
z0559ddea3bdc26edb6ce6a818d5cfccd7f71ff657b1c669ba106e0bf6ae6a6f1fa4d8cec5b39f7
z28b9a0c0c0007dffd2fe493a6c28c4e4a5e1d89481839dbab0d0fac81ab0266b16b1ed256051a3
zf283795f490fb1d2ee35cf16a985a85c108d75de9f6ca82b742e965ea15f832ec541276027f6f3
zc138fe5a9ecd8f236758445c9a21824329d1e86c66cc0d2bc82525808db8b2b9c6d046d940e905
z2fd9b0d288c7166bb8efccb83517c22829ff80c3c73a9dc7d636178c6af7a687bd1ba45fe6b031
z141d84c2c62bb2693e404243d12d848f217f88168b3dcfde4ce8b9c2b70d578c439d34fab7c7e7
z6987ccaf63cc4610207f522d3a3178d1653371fbdc84e9e9b9d546bd11dde18641ec2704f0f7b2
zf973d987b7606cbb695f2bb430e5c4090371149e572393c377b8296fbbb91f023cc799600768bf
zde99d7113167dd93f11daa519f0fca6ad4b5a27f5c1ad813e5564872c97ef7d11ed591354d2d93
z84e43f4da19b7e8acf41bf1d4e03f9464c5a7e929b5dd94f1148c94ba4771fe4d81819e919faec
ze28d773828a3b2f49d714a5894a745d041433f439324645bb7b4d3e4777448a9ef914142391eb1
ze3ccd391e248a061d90b35ec9c6e96161ca393adecbe3e30019c462ad683ffdf6b2836649fd4e7
z0bd8f3d247570b138d3dcf47bc7553e1737267f6861442707d9fb6457a30717a59d2ff3024508d
z94d3ee55330fa24858b659e9f372634b0a53353ece8ccfbdf5a791bfe80c835938039cdf49e2ad
zb79279bfa4fe373d475b5516c155eda6df39a976920c5be1858bb15e082b9349c3066affa78d09
z30518ce5277a5b20a1e2adaa4719ef382356dac69c0a701f86f9c47d32297ef42ef1d91bda2d70
z16d22e8b591fb00e234290c45f1edfd6bbfb11badfcef06cd511611b9c107fb1b2af896abbbd8e
z35110d5c18ddd44ba1f0ede85f8cccbe25fd1e07e4d4c25b83e5b9c1d46c488333bf551d218fa8
z1308225573a98a5493f795a49454bbcf9c7181bd35569a77bb51bc9f2f1c7766396734e07cec17
zf26f2326369901f9e9fe99637fec0cd7651521b54e1b5c2fc797959527f06794cc8936d345fc1b
z16f6d7ab7469ec600bc5587694a02739bc24c13c208f7b2cb131a9859613c2c0b658332e430831
z2cfbf4e3d8892e6aaa302573cd846615556887c4bcbb79e78f342629e78880d65bb70268bdfa62
z8f2b8b90a597c191128de230258749babb27abbf269b62801acefb59fce7fc44a08b0cf096be28
z06d483fe6e0f7ee703de88b4d107584e6ba85e14f5c8701e1b1d436ef25f96c1b1c0ced144ab8c
zbf43eb8d84019f485414649afb7e51329853f98834fc8d839aabb99f3129fa4104bb9c5f9b695a
zb0eebae30d957e21d9d517c5a30d6495c71b0561d21949e68ad5dcaab4fca661ac963bd5185e6e
za1d021bddb346960097a1ff3a138dc67ad855aa47b365ed287f6cf9cb3fe99e603fc4bc648d1c0
zcf4f93eb7729a924351639ee8b2087c18143021a2ed06ea55737ac3572104bb27ed89e2322028b
z56a6cee41c0261e87bf54fbcb50cdbeafc186b797b25b99c181a01891e6506f7774626370f6ee8
z8dfc5faf659c6819f599b3fdc2cea8b73fc545c513c86367b14bb0f98b983aa8d546063d999e45
z8f6b7a231afc9f5affb3777d7a457ccfeb89c37365c131a27f8e58f4cd9633b970d7b6600e91af
z072bd8138b35ba46faf5780840f17ea0d6fc9694a10eca32e7494ccee0f8b589540b7d43ffeb2d
z34de5886f524218b9c22e7c3231c1968e3b10e2e8d575c1f8709846b7644a4754256296b97b321
zd6a2345762778244b666b97b286d6373fc219c943c14f293c6404c433f29c3da19e2378b3b27ef
z1bb7b709f4d7f3bc0953e64bf8c47dcb420f32188fa9d09fdbfd6e81b73d331bf7a0f7809d6bc3
ze8974299e8fdd87131194afba6d9f7578a6610f8b5df6ca5ec3c5eb693f313453c9c23fba90da8
z924c42e935d9b226bf789d3e617755b24ac3f1f0fabb737bdf3f45d64887aa786ffe55e61814ba
zd1a9ff2c01ac0acf95fbd1bdf8bcd34a9ac9f5330eb4c75b46fa84807c9bc20d8fa40a509fae88
z3dfcbfb77559de99dd54e543e4d82feaa4e671b223343fa065dad7654816454c720c4d4a679caa
z6e179c9be8f3f1a7b65dada43da2cd2ac66f6f3ba51f24dee43f3be52125f3f20043fc470305da
z830ef265d7c66951694e35a5d240dd38d57228e187eceed63a84e690a053062452f72c5d5dfb39
z99a72bd441d0e32b317117297b2adb1a291a10736d6aba4977e8942458d82d288035c8b4ae4248
zdd7ae1c827d6e0da3f1b874c5a73ff1201e54544e3015e0211713423b2b0894701791fdf52d76c
za0359cafc6faacea987793f30be5dc0715479b416ad25923294700d70a99fb6068e693959b5c3c
z627e5c14259e89a24e34410511db737e1f8e4c9d7bb7addf315f0bc84f2d633c2113a7c45162cb
z61a98031a4dbf72f45442dfc8ce39c6260ca4faeca65fd4fee4dc54d25e3ff4b5c6ae14ddbbecd
zdaacfc735b70fccd81386f02e98fbde007a0347643e16900b8f37dd43e2b8b312f204262963cc1
z5fa57da05c325833e37d23b77f57fc35cc3df9e0b1cda075b1092955d942d0ccf2c7b7c3ca0c96
z127473bbfb0354af55a1396bd47d6dde62c0b263ac47f934953a8f93d78966eebc0e33e6146666
z63af4cb9da951b655fa9483d91109e7b509dbdd587869a5c1f069dae8a834cd6f48a1e6024102b
zdd9f5e1e4ac58884e0d2c5356c21a96eeeca659ecee1010d53ceb4fdde008ac57e97a1b83249da
z712538015282297040af020e2cafa904d5606ccac14fe558ecd436643224e9bff919a4c72f7f6f
zee71182edd70dfe07459012bd23a988934617a8cbcdb227e3cd0f43fbe394b92b8281b97f1ae84
z44e93087dfce0303ef79b2888959e4b0e43b08c10fd8d33f7bd78b1e48c883491e652bb4b9307a
z4f49c2e0b14f0a90bc5b51d1dad65fdaf62409433df9cc0a6fc326a37c43e0df5551ea49552f3a
z044a3ffd30c5a032302462facf4651704bc875b50e0e3119855c97ad9264538bdafdaa8770b6a6
z2842a2adbdfc83138851c77501231a7b1f82e091de21ff73d54f76d1700620f36640cc4aaf370e
z93e755f349713e97a925262caff6f642848c1e7fa36ee1bffa9cc75f3a8cc4750f3adf9dcdda0b
z89ee0d466c7d94e72e5a23ff12ec5bf92200e284e899c734cf13814d7888e03d940dc49be44221
zd0f10fe684c15ce9d19001974bd83fca25128203ab18d7ca097a45b217c1d879e06fbdfb84eec0
z983715518cc7ce4729d876d4101206dd12e72978ad6ab17383e88d7f08f5076288de9ddb81f564
z2f18c2e960ea33f398c7290ab11e20717232968d78baf4db2566041cb1947915e395e1eb92b9c2
z3710c7b5728e204329642b28d77dcde6f65c6de51b8994d38b6e5446ef777e909d2ffe1fd5033c
z0aee7b4cc05ffa1ed0fea5d014a46e7cec5a88e6e8a16ef95e17e98cde47f1872a654e102be4d0
z33cacc8edf4197b067eab13f56c57304beb463c46bf4d21a55e748f6c988b7f343f5b5da0b24c0
zc36bdde7dcd34c102b39792db6a7f4fe729508053984afa68a594337e734edf24bb8a5b4794095
z1c3138083bf850539a9b274efed0096bfa8767097271c62fab40db7c3f2e7a5d545901aa067cb5
z45ccf705bc3418eefbb5bf014d3cfe80a40e5060177fea998541afcea68d7334457e2d6e9fb1f1
za9f06ee36a6dc48ca926ce5baf65008f0ae92b8cb56b222e69ce6a8b0fc11f14e6c2169c34f168
z6159eecaaf4a7d50b0a686b9d70d08764215b5ffcccd299ce67fcac9e4392ccfc19aba5c537ea4
z21f72d78733d0e4bf53ba094282e7d8e615480acc1527b4bc70d87f208f237abd4a6cb6b313855
zf85e86dacc4ab026afa3479b98f2fb6201f462068e89b23777234f0a1343125e7969d68fb24118
zd91c5798729edf0d120c201026f3522c415abd2f4edbe4c491f14270aa67bd64660566e82de8d8
z228efebfd2274480169e90a30d4e07ba995c289b6b157ff95df869f608d20523c0f508cdbf3430
z749acc39c84c4b2c172479012c68a4acf157810acf25029d6c57661f559d5c6de0b875618e03fe
zc66fc878905c808a5da89907d72c757fa5747033c4b9dcdb7ec39c52e60fef752f6b21e23c304e
z5509fb888cb1a2be28a2a1e6174c7c63cd23ac7b8b11566c665287db8d63913e14d740f8296cb9
ze427fe556746667a52c5f7d215e8175daaf69b23719e14a5f04da888bfc54d451bfa4f90eef12f
zc951ecce96a64011de56a480bf2bd8c7e7e37d2c44c09689e9135f7866a2ceed12eda01d6e1b32
z1f6971391c3b1b0e8beed8c1ec84e6657beb433ac308a8c8fdda91f771aec7b4adee16e2a07134
z9b1c51ed4e1a3e90cc118683ed52ab8d73486a25c3d146cadaa0985a6c4eb5ee0d91db750cd22b
za2209bbd018db908e5ae509297f37e3c359b65ab2dceadb3179c5d196c8a57683a2a1c937b12a3
z8f49b958b2f38f5c11f7fb0915107f2eb3a37240243b9a444a5b599832c0df9081be94771477ce
zaf29659397e1dfe10fd5c9ec8723cc635c67f316036c51a1797d1ddcb36dc665057e7fef9f663c
zfd00b5428913225f873e8e0557472e2cecea3402db6d20ebf3f855c7f15c6ab9e3a75feb8a5cb5
z9c1f444030be58e0acc20d8d31470a17888f81634a7c1e27be671771105daee3647d6dc9b60758
z0401a76f3ec0021b042cb1fcb594417fee00439dae93a603b72378e67675041ef59009ba53a813
zb9ed8f2524512e9040cf4e880c2ab7f3576e9104a581c5e7283c54ed0e5fd58c31035b0f570018
zf5c41ab5f601248c9e9ca7f836ea5d01d92395bdb5197426c26f1fa52d1f386ce62b56d27a64b9
z4c92c5dfbab0615c43d115f7ae6efa7bcff425875d1c3df1db00b2e69a89497bcbf3bd7c1a1619
ze19e8e91b6edfe41cff02927940c1d3ee2b93d93530bd1755bfbfc4feb33f05c1bcd2f1ce082ed
zf2be11b9856d865ed7c00719d3053ff269486596257b3086937deb78c982a9a170c922a16ceaee
z804ded890ef6c051a864ac4d3851a6e30f55867bb968839ce0bf205ca51ea30bc52ebb9071a5e7
zdfe1d5d54f7569d6e2d9978ae134b054c0371a4e29f07c7ddb9e0c7df723299124f7358a8ac3bf
z444a7e7770a12e97d11c0fbcf5fc677b2868797634a7b5b17db664d3ca397f77275a373305b909
zf7276828adbf9bbffa4679c276aaaeb6ea85e2cab0a64f98735c963100ad11e87bc5b790f66ac9
z11b32d8c219661839b622a2baa45c818b04a2c7e5da630de1dce0d05800cafc2a29643ce02e8e7
ze91bb854e528472d5f8a2819f7a0b64fe2af1d443e586a9177f98ed3bab2202204850388dedd3d
z15ac0340049d4bb8da0a8dba17bb677426fd0d33d690b5aabe9c5995a5c54f782c80877b49549f
z585177161bbe250c04ecb10f566b711b5d7a7ad3c57295a649bc857d8d7a48884c2deecba4ac33
zbc7b21c2641af46c0b31c34e1995d8dd3505be36d0486cec4f2f57b16a44340fcac5548be78f75
z33211b266ba88c86b1e05a45819d833793c07014becd751d15ffa399217ad642eca098824f0013
zf64745957be98ed3c7aa9bceeb4b0af78d3b686169242e504cf719727c195f5cd3c256f63d2e7c
za30391f3bdd8da90f777f236f454cb4ad755a1ea0de0528c1f7968f15be9191125c6429dd8448f
zbfcc33adaed097fd69788e2938fb055f8853ba10bf8a8f19d13913354e80c1ea67694a2f324705
z59f8fa683a5edfd149dc813f8c64f4681867834b198be9a3f0174700943ef690d88681c2109caa
z348060c34911fbba3cae2e1477b960fbc6ccf855c4e3b269d75c82e7ab12131fd3a4b5aab4ca39
z82dd4bd25c4cc762120a6bc7420d4777eb74d13aa0d13bf490dff6b87255a22da094fe06e6ac04
z5b57f221a91f6697cab1863bdafb43f94fa5dc2d1cb53ea2e37f2582a62e7cc351bf3357086ba0
z3ab14e28cf9d42c482658bf7b36115e26831d88a653b5133fb4774f44785cc2343e369557647aa
zdf63377c516376c091537ac98ac1ccd2e075f91c084a7530f637a39aba901846aee6fac3e74441
zc3790e4bb9f4b314ab796dd58fe39abd855b2039fc91563c246a127afda058cd49169213b13011
z454d9617d3c17b7e5cd2118e862029ddf728ba9788ca02df1ae5741ed169383684769468b6fb83
z56cc6c22f96bbb5da32137098bf9a1a5eac5004d365c144cc4aa2b0381fb9bf080e152a988c5fe
z50b44797463701ab182e93ec928ec3c09a7b96831bc33bd4e9dcc51365cbbd060431324d2d2415
z1dfa247e30770036167dbced202c8159fd1fffa8a78af2f60b9e08359ab95a0c3845d80dd2a5d0
ze3afacb45e97fcc96574968294ad9f6841972650191487d396ac3baa27868623e4edcf2d81de5b
z2072e4454080ab8298267917983c00690cd6f954c436d41c95a31eacf329193d761391aec2852f
z02d84312453f28519eda8330acd7deeb6160af2922dcbe7d15ea8d92ca642f426979b1d5410b33
zc8deb378c389ae4585454c6514b371946861012155ec0b9670f7329668734a7d6e634d0a7f3b53
z232318163b9b73f3e368db71907150a8f1e4a37d3e415f2ae84856bf6ef84b08b553b81e71782a
za446c3e846d911ab8cc05461773ae4bdab156b2a9cb0829c977696dd532199b66410d4b6f89d43
z29ed93aa5327402a0c2e47a0a6d8c1ee1622e491bf05839895f6396ca4be8027e1ae13e47bf7a2
z050dadef61c39b67f2070ea64bc9928ca6b8e85edcf40de696702cb8b05929f75360d42697a835
z56774757e815a8a26638182b38ccaa4a902f465f0394f75ebaca19c5d08404036a0d3c30b134ec
z67e5fb7f2d8f9f1f2a9dcd994acfa16ade63b6ab5b440256d97a5521eb9334f022e2a6d7c04a8c
z8a3bc15560033f0068c947b217098d8f40572deeaaf3ec74a4ffd814d589bf564c0ba36adbca6f
z9a8a519c858b5e2688b5ea5365320d87a768a7a1dd4ba5b8491386c206a7872c86085017fd2570
za4dec5402cb7597f66492c0b9b4942955769ec36c800c034a2710cc38ec757dce704c123534ec5
z72323b7f2a58ca2de149b64cc8d9d2c1d79c479d9431a638ebcccbf3d1bac9cd398effb27c182e
zc240b330fb0e175595c5bb796c7c771abc99b4ca4a55154c780fa2ec0d995f1436809feab63efb
zb7d0882295874711c01a04063e25b233820ed33b8f9bce1147f87e20b41c34dbfeb498e2734fb0
z3106075edf99af20256445b255ecf4ed4f6d51ff2db89eb64767795c82e2520a429ae12ecd01a1
zc63a3b330e39fa54d0fec7e18b51afddb08cd1684d50b39fa447a40ac7628be27550f12a599fa7
zd3cf871987ef627e18e452874b901eb6541d733ad11d7ef428010af98e24e7b11ab5ca5a4184c1
z51f5f1e362a447dd5303ba9ee954a6b26a827edca3041d7fb50e558e9759d4a7bb2f4a62f6c913
z4cc1c9a1fbd32b96b22439110f57155da266aad78b89881317e2a053b9377304dbcb6fe392e08b
z7e1ba153ad6d1d129c1754b155160b2cf9ab7560026c791b26ab56eb865c8c9dfdbf11d6d36e3b
z96a3cb4711989784b28b27ad55518a94ed04cebd30e631125f4e4fa96e75fac603402b6bdc9eee
z2798ad3e4193ef808aed664d3ef25b3bed753b1dcd83f19a8c4a1e8c1372ca6d7745aa92df0bd2
zf9e4f330bcfd57839f7285ab820bad648bf6e556bbfaaa84848b605eac693846a8c406b2f813af
z2de68b6d50b783143ab7e9fa0640510866850b4545cce2feb217042873e3605eb4943d35c479ff
zbf95645e5c17a20b6af14e4eaea38131a274395d9b5e2838335665a65b09054a4d3ad01154494c
z336cc277f0cb8f6a198a130655b54b14b3f997e4fa5f4754b5d23237e3dbb124fddfea323fa38e
zf1d54a80bfd914d3db44bae525130369c652c88ae937fc44d56ab925b0957c3f3f869273342b2a
zf0f8d9c703a422025b9c8fb2da1e2cd765344dfc1595ff4e1fdf0c3c8c8012f70c45b15c4fc558
z2ca9106cd5b9159cca49fc056a55e49985d9ad4546b240acc9aeb1949828fc6ed3785b457f770c
zd064a2a448b436db1ad87568336b0fd0f3fe185cf2812f0a292ff6169b290e02ff86410f990ee0
z3241810b15795c14b1c8ea4474de5c833f2aa99c5f8db382bb9a4a3e23e0b91901dabf3125c217
z07756365899084dc4c0664c1fa86dfe524eb8433cd623d9137455ad1edc9158ce249c7b2955b88
z50eb546bdf9df5c81d7e978ac066d4a41b6081913320f772c94dc7e0bdf25031cab5177b7b6aaf
z2a4f83b4c005696da64b0f0ce2a424b4cb8f7add0d72631abd1bfa572aa485725dd26d09ba3b91
zb840a3f568714c2a27718788484ecb4f6b342c4c9ed860dfbbfc4a1e1aa720cb2a69bba14a74cf
z55b471fabed39461dee697332d260654bff877ca6bf7774a3e92cba856a758efbeb808af92c75e
z1f33fa9743f0b1fc66ca82339f538f00094474e257e3948b8d4f31c600d791f2459b7e06050569
z7f9273c6602d0d17c14d5ffbcb8985fc45afb0dba7a86e157e65af5ca50dcd45128cda6b2211f8
z1a2857659d13ad85cf81bfb9a848405de59ce829517c42ba435bdc2d809bc8f108fd5304327b59
z4d71b71d92473125b1d1c3ef1bac5e6b6527bad01643666b8de5ea4c417c35f035e05ce70b5a3c
zd4384d051a3af221375a36bf21c1a5bf4ecd86e6354c8eab20beac83c4a9f1529c5d064d47f8c7
ze6026a13544dfc055c7e052e631596241078264b25f9e15d271321fa9ea6a4ff5b7fcd13d20927
z711f9a41e6f6692837d3ad7aebbbbcb683add3ea6053771cb54d4d0f9de4944d29a7e8c482f298
z2863023450b2f8a444c82cb39e0516e2063171c892080830a284a6917b815455caef91f37107ff
zc59aaeebd8d260e6498d9b342ca39b52affc24ec100d14d9b90342b31838e761466d0473fb2fbe
z8c69df732413852d87fb3fde27378f9b38c0a26e914cd066094fea6d718943161139f43287a97a
zb4430b8bce319958852c13288d28eb72c2183569fcfafbc229ec71c7b6b43d930a74e1a2ab1ef9
zc0545ef8eb9c633d1047665f52b6d53daf2aa6bf665fff473ace4227bd4f37ed938c2513febc15
ze3920d4358f31a5828f44dd96e89f0bf87768417860d5f171d3b8ba5c43b20fc2c3dc84ea3c68d
z1bd028c1b244e7281d66a8a5544b18371a3d09e9eab34455e9e60cc9c0281e5eabb1d9bdb2d2b0
zef30736a9a5689c6e04045e04d3411419198c4794649679b20a3015fdbab5875fa9ad50c0fcced
zf404486c347c87bf0b381cd5add472a8c0c7357857c593780eb89f6644eacd9ef36cd3af3d17f5
z953052639e978d7d7e56070089b085169b1f8f8d236de78d6be56a2a051795d8f50a9a0f053906
zca164c8b863e3f166c79ca344adb154340f365599ddb25a39243d3808c0f4f9b7546a526a40fcc
z58b9cae393fe0fe258d4bd17b2e0892b7ac1768c5bbf2eaab9d8a9015b39f853add2f54d0edff9
zccd0ffd167b15c0701474ff197246f51edce2c6d86965bcd9a268698cdc8f8c4dd4c4783fe309b
z82bf6bb5931d77544ee9f3a3cf73b274be7f3150aab84d0c47219cb0f8b3590b43afb7e95dec57
z2de3ccf49fed94231df7768198b5ba6d4ccd02bd1c6c0e70c32213baf96af468049320fc686024
zd6dd0b6859354b4dc5161b2d9edef2a2925d38997dd5fc453335394f4aa695a9ddfc5826fedfc0
z5a0c9eb4da524d2de7dbaff284c31457fd38e3d147d2dfef760eda726fdc063c34aac6fb928612
z857d5a7a49a7161896e12737fa9cd18f919115238d50c7171cd9eca0721e9ae269a05823e1ef1b
z638370af0ad9b450a26975a33f48aec9c543bfe8c75d10a0335222f8b76151ac27071d5c1b45e5
zcded796b257065f56c59b0ee2907962be4710ac1a1c29ddfa79f1f1ecf0d7be15123190c0945b5
za354a8098f8beb012ea9fd0d9c7a8d6f59ea9f30183b1e6cfe952f896ebddf366b5ff2859e2cab
zb8e41d458574f90210650f879302b16c2b4512b2adff2f2c521a40bf487c2248f56cc189e47f3c
z0c2bbe7ac21c7442cb467435a81b1e99ce006c0881330712e53c52e4351243da230fba4f3aadc4
z9d89566c82c2c8b2053200f3774042adf9db35a05ba1a05dd6fb61dc35212b0aea1d42c5ffac79
za166bb70498999bb6b9a3f628d0b2eb460fac04f66304a20bcbd2d834479e1d313744338f39e0f
z2415644705e4264aebab39872c958f73bf25ec9aec68fa8f2bd970d146602707618c33874214c5
zddf2dfa4d2aefdc98b57aec9a8f3185f33a870a4e8ce8034acc63275e2a3c8db9ac0f4b59b7546
z5e1041fbc64e259e55acbbf4d62678c86449437c26a51085f62923bbba31019782f766bccef6ce
za1c7592ea24d84faf39bfd469a72386a144cc90048e9de120832892feb71a469645558e65c5b2e
z2c32db6642dc0679cf9c3da1fa5db1d397bc65384d02ad5f53150126ac0e6f15b684da2cd45001
z9d10952c258a0ef548f692cc4aeb993d85043e189e8524478cac5d326e1ae711970a58234c71f9
z162828dde9055ead4bd2c82405a676a11190278e5dc2dc4c3867f8cea12a1099a2badd358d157c
z56324f7ca9b0bd9902217954e81e7728d9dc4282c1ccf0b09aa1df93c2dbb22734c3fee120ea14
za030cbaca6e0429ce440caee2d0b786abed9e13f6e5bbf6a3c1f614cc2a69d21f052a0516b39c5
zb364ad551a4876187b1fa0b31dc25056aa54bcb651d0d0e763a797a45c198883f08f76f0b8ae9e
z10af36678b99de790630ce6bce9637f28e851ba7f9f3051c3584b0e2e9aa73169eb7848f02d67d
z3a5356d3d27f38384125ddbb3f82441d8f359ec9aa973b75ee7677e6b9c613b10862522a5a24fa
zeca3a886bc01ffdf93923eb5d0121725ef8becf24332004768c94635e0cd32ebb7b4dc6c0a6d76
z801687fb885f7f8defe5379f3f4238eec42a7c4dae4255e0c7cdb3f4359121376948ac9ad404b4
z39d72e9c57865bddc255d1256f2ad0ae5f6dcf30ebab17f970adb0b07bf248592b1250457f50a1
z87c04b2f75d188c01b63667bf3022e6fa1b15c53eb5bd3d13182636729d2e82d1a990a28115291
z247fd4bc36cba2d4607c65a2ff2e4379476b8c3ee7998e3e256fe6ddbace86934341784663afe1
z75b3bdd81103b3165da6260229239d8c41945281efea53b4748a6dfc9e28c3cd608894b6bd2d0f
z2bec02afb76daa418fdabe6d380ab6ceb1e4e4647238d67eecc8db30661a9257836ba80f491a0c
z9851284ff1fda2e9a48080c58069fe6f5ec43ce8298a9e9c54fca3c61b0ab7e29f70f202fa4621
z31d37a68a837333a25e3c1315f43f48c380d6c8cdc95acc51155a8a3923f579b1c60dc1faa44dd
z1f0c51e33b7450e76da7666e628b76cc51d57723288b510b4cc02a3a6f6bbf2aafc0ad05289b80
zc6b76cda44645816ead978fb757bbc5cea9e9919999abd550ee18c569ba08920b2eb26867114cd
z12a48d96f4fb4800ec6d1835de4a83953de2b65ac1bc8a05cafca9f5770362eac67071ca21740b
z10a49647f1544dc8fbd69f0a476cd53e5df366f9c59c8b0223d63bbb294af6607f1ae2dd5297a2
zc118c2fe1323b9be081c07bcc460921b2e4c3087021e5ff9cc07530abda75ab389080b3438e079
z1c6806abdc9388fc5045aba55554151a5a2500882181c65293e7504ef562439af995c2607b364f
z9c0aab2c3a9ee7f87556593b9b42b16dad16a8f0f2e1b4214c05413ba692156d99160d7b60485d
z20f23516551f3170b22f3333ba3548d1bca7e0f0b1e2149024de9bce4b746225cc1d5c633f0564
za76735d1a0256b5c4dab79ce3e62e515e9e589ae194f2f7ffc07839a64a0195c54bfdefa764f81
z9bfb925ae887ae2f9007106862e49d8429ae82237f1429c672aa361121db170d31071286fa9b89
zf0bdda34b5efc11c82dd7f268fb2cc34644f50258b0c8b11eeebd9ae5e5fdd55ce3de29ff5fba4
zf574adf9181330b5169ede3d44a6d2df27a472e85d33e7efc832987c8ca72bb49d61d1fe5d16e5
z565d7e62375375151a74ebd932ac504e9f5afbf64c200b88e47ccb352148be7e59f71484caccf7
zb764005d3467e8d12f0afe0b5e362c07265a049df3b375d0a2f53e98632f3fd13877bb752255f0
ze608c3dee493b471201d10698ead814f0635f68459c277001992694ba0035cbc815324425e9a39
z553675339edcc8d304bd31236c4dc01afcd8c2141cc87c79b20b6d799cd9d145a3a235faea05a7
z4898fa2c9ab8c4e795eebf3665e788281ee215366439c7ca731e84af365eff73b4f86692ddad8d
z37926761b21db34950aac01910a99d0ff3937059515de3c0a9128b9c0dbf31f998bbdd0f279713
z81bbcf2fcdbe40ee28195257295e0c8a91da32e5da9b3fa220470ffaf6ab909ff824b2f42ed0f7
zb1a138737cf058144cd0155ca0a35a942b2a21b8c1eb9b89ad0d757c29f523b6bac8d67430f451
z7410e75e93f73ccb54d44365494366042976047281c64e3cc80edccf0daa5897ccf1321a5732b5
z98ff2734b35f360f9ebf9b4bc86bc138ac46b9392a7a59d9a8cf3461dfc3bb326095be17cbc98e
z6cef18766b41f47e1b9514bee6b4ab82810035dd1bc398a9a20cadf4633d0f21890cc1e7985be9
z83cdf9b4e799dd9cfde7554a91396d4063ddb00b2ac549fc6c7dd74edba40d91aac7a39a764910
z95c93dc4411673e46d82d7b307fd9c92fa3f0ddbabff0c49e98314d3deb0a2ee23e23effc47f2c
z16ea6163720cd9f0dddee7efba9a7e9e642b952a4bc628441ce41a4c71ec4782165292ee0168ac
zdebb5028e286cb1658200b8e0cdb2f8db60f7317ab08c25a49478674a303b28b7860c8d1733d1f
z9be09dd7019b90541c656858de5ff780ee31f4b7e0c5182ced9529ad82e4e6827f129550f8bdee
zc397a4ccfa14fae6ce38f4d6fd1f5ce44a128f31a53de1803011ba179a1a0beb7d81a457f0544b
z64f2ca1f55be2806de0899c4a6e8356fe9b7fabb2789c4e4fcda9c4968a0d989e8f5fc71d6de3e
z3f29bd40369622ef6e7ee8d3d91dbcdcfb03b7dd05a329f17dc9fe1198a49c5d2e3e1523bd8df7
z76ed8af7a63a0036247ce7d9fec9537c39259337ef5b34826746405b95a8bafa80d3505b577ab3
z4dd7b3e064196b95bf451beb0aa85972679d19f7cf9295e9faebc39d613e5bfd850888d7918919
z1813085323d91855451b5abfd82f743dd53f59f73c4255e0bdbe1de906f392d0c5cd1a52a65a95
zf975cd4370b9bcbbc9306720e854ad0537a7d5b176f14576c81cf5bd514d7060a4edabbd18d9d2
z2f2f443b0184a5c0b5ca860db01f460fbf66c62dcdb9ad7d45d8c961a1b69c5bce8aa793bf8b2e
z6f8cbb6de2e75edae11bfbe984b0af0e2fa20ab75d9a7651d33ed61b9ea983b7c766f3a5cd6dad
z0650fda4b28cb1ec1ccc723ffe6fec12d40a5162277f25e754a354fe98f4136640550903c3dd6f
za4d9f98eac01d69f859414c1e514cf6bfc15fcbeac101701afcc0629e47d1a39e74873083a1953
z0d8141a4569e5c61067fd3b125456576779a048e93a2ccb0f14aaee6776d068d1949505112ac17
z315863a75deafa05d1eb1fd04624944adb6254523d757a07a8e217e655b8f3cc8b6cc3cfd531f4
z140e1cbf20649bc955445db0b3705a5c764af42e7fe73016852f97d1760674a20bfacf6bfe8d5a
zb7dcd3156bc38b90e5ae43f000e1720ead2e8a6914c64a9047b2d82f75fdf1293d95b0765c082f
zf0a71be87dedf977b1819927f189112a580cfc2022c6723b3a583d72310c7c1d881c040c796afe
z73f383cb799f457def1c73edfc019bb7384484f334a787fc73170f104c3c16dc4b1c80a219f795
z4cca0f8936cf3d9ec9188d1fb73f013171c0ff58766df249f1bfc600866cc46b7831f74746f38a
z7b7cca289af4ac4f2f64b2bbc92652c7035b2746d5d218415d9f03ad35a81d015c8605954d01e0
z78f2ad3e93d0c2ae77fa5562a1e41afb726baf45075fb73a104f4a4357b0ac722b29db103bf9a6
z098daa5221fc21d76806d2f8f17b6e9d312b260209898f27a0bf56c6c4f2cdb6724718bba56890
zdabb18d0f41e92a793ee40cf872aebf26f73124e47aa255393d27f3ff2d5546108f116c6d1a574
zfc8b120f971285891be57574e47fb79ea91e64779c24b2293af8e6558f9973945db20f40719994
z0dae3aded8a043ebe206aed337da1329ddbbb807dcfa63c55ec65284c0408fb1ebf34088d92959
za058b831ca5ba4a33d06bca08c9de6d055d31ebf3fb673d7d64e329c7e8f38bdf2a10284a1fc97
zbf5c1c39ccd2f588d00ed89491bb76613bcd759b9e026a4d4e4c8029127033dbc9da5037c649c1
ze9cf8df4ecaeef53cbe55961a19f8c52169ccb6eae802a4717ebe6919646c8ae76071d77477ae6
zd209c730342f2158a75863bdec940749dfa97d8fbbf9df2ecc869fd15da6cdd47d47daa244981a
zcb301dc49bcd396ff2c1a67d7edeb8a86ebc440bbd56ccc8ff278dcaa5774552a2d1bfbf905f78
zddd01b82993ff79b21b94a74df10b3c85c9dbdc5a62b6ff52bf13e191396310543ad460db64f98
zf2516a405f06213ffa270e7efafec9e2a2261270e2586b3d0e3c46ac03b8bf230fbc6bfb5c457a
zac79dd7de4781c5759b824cf2032324dcae93ecdc56ae6257b4522ea9d87919f1b2def53d876b0
zf171f1774c7d770ab83bce87abb0878f2855cf39deec8f0687d9f755db904d7b0418be384409ec
zf686668752966dcd49fc0325c3fda4470210c7cfc7baf0f1d9bbf788df0ce74b6cc4aa459e9f10
z22ce58c1caff1861d408f62ccbb5f4a750f31b67fd5f2e8f02842b18dd95d534b0783350c2adb7
z2acb778ced793968f99114bd49a67eea5b6d98489555dcb6e43a466c55f432296180ee7e782c7b
z628d7a4ca5c9cd8fd1179905235b8e7374f24db01ff0879608649cfef00ec740993e9bb63aa505
z0ef50d601156f53d4acc6b3a79d935e3b9472480795954ea67dfe0520355d88610da110d61a2ce
z9a72c992b22986b688c8d2f335a49cff1bdf03f15420e36ee2609a918bd98594090e6fc650a903
zcfd6b60db47fa14255176db36be42c7882771220ce562771df54dd6a36bd0f2b9db436b4992e41
z99acae10d11d7317fcdc04e30479f3b3d77ac721ffb24a9f03a7da6ea790837993889d0bbbb661
z29e77023b3bc17d766188332622a94c6f577114fc40b278435e40c9612a9f861cfafc12f27e02b
ze2b8dfe77b171c50c5fe441895e7687ee1dcf364f32ae7190346cf33b6f5e0a02bbb7f4a1b1b27
zdb3729b90999843627f22226f202e1e2e79f13a3eded0a90a46fcba308d4fc6123490cfb130b13
z1b0aa6ed9e6e3508d7538d85bb0af3adb3f1bc05f86ba5d143c11e32595b4c97ff7cb07ae5156c
zb5d7217481d59d156c3bb0155294eebadcd1da2e6694524aca3aec59d7142ace2853cd7197a093
ze73fed6ec7bac5ab504eec9ef23f46d28ac04bb67c5eeec1884f50be8426f53053cf3379ddc2e8
z2d219576907e8f674ae5ff86b654f02653c0587b7a2fee4c8e10512fb9b16fec9da00f86d30ffe
zc7cca65a0caef6dc056e7595c86bf9cd56737d332960f07a2c8e59566d0c39b09f756bae98463f
z09dff606f4716dfa125064ce248020ce7c1076f9fcd11ec5c349bbefd210dd4db329508af3f596
z5f0f8386eea636ad44d53047299c0d594210a2fbbb5c55a9e11bbd13aa02bf227aafc5d5b77b14
z261eef980376f732d4c500300bd4841e359f2a8ef01787f3e606fe06b00d94b723d86bfbdad088
zdf6c37807cf728d2e5c46094ae572ed0fb674b12b21058cd7f2a51e78ca9e22ddd41f3fc6effcf
zc1ec0590345aabd6cf054cfe99c0ef72d74bd49570a02421dc36e7e56328b3d8f37b23b5cd21ff
z74465de61d71e746cb630645e9063487a9e21cf679dcedbe885a445b513648575b43d5cdc645cc
z63752febb50edd1e046dfc71ef27270d01affb6c2f3765691df1a634033e206044863596f8da00
z8752bdf9a3d48b57e2b1691726edd87c6725569835539dac6fd5c9f68c4e8f49984a30858113bb
zad5cff7b8ee5ad730261ab9371ab6b65c8b09fa08e70462228d2d43ce4dc459dae017737dd2822
z0135d46df01026d56820681d4d43514ffa5f032a4003516534f753d8d98db08362747c0ebed211
zc0466768c63092234162867a09ca310656ca4ad87f3267b4f55952ad8d0c7feb343e5a39aeed56
z295138a892304226f09c7f2a9cbafe053f9930c2db8e59dd604e893190bcfdff19a76f6f2698b6
ze3dd611c9855f126113ffdd58d0ac91be76c43944b771766fcf8b06765c9106d85ad67ee96e610
zfd420b271dc3e26986c3efabfe4fa6deb1f6415df63b78c28ae3d3bd08147d009dabccdad5ae73
zcb5016f412df8eacba65a324620abe78021066363b927b78dbc81636cddf3d617fcf18a8c0b3ea
z2d0ec02a130e1899b9beacd45f57f808bd6a6e8e48876f5e43f1c22512884f4da36b72372a718b
z7a425b0346fec000ee2111267217a6d9f2fdbf2b071f84c0cff966a879f6beba50fd4d8581fb72
z64eca81ab1a42d85603aa1090b84153395aa5fdb443a48e4d941fab142b1aac9dc85714bc6a86c
zb9fe88de3ce733045e60e81d8d91d16faea6b50dc3fc6b7c14b4b5f4b81963a4254bc9663fc0ba
z743f0d637db0d8f19392738d9233dd33c7b2c632a26d33894779a6bf466ff4fdeda1df0b9a454e
z610a2ab0e9fe55c92371017292261ec1b1bd095913ae122b4bc87d229b8ad8ca265395fb9a777e
z937cca95b9e0b70f62732e0d2641812384658bc93b7cda425322756196709f3f3b653d4ec5943f
zf874a61263a5a99295a0419f7ded84b9faf7e84778a018d3922bfee82a5fa6fc962c22cf20eee3
za0f9649d16b1b29f9ff8373b19fc9268ed32fd082989fff32c380fa68580016a858332eed88c0a
z051c1931afcc5619da0697eff9d9c21a1918a1adea832512736d4cbb82d1e047c31481be468eb9
z9908e70b251d4dcf963f0ce9df826ef6948a8f76c098d59e90fa5e6eefd3b0565384631c2ff603
za89add74d839a9e4be85683bf84aba45146dc9664ae63ece091c07fbc09c251f1f4691919be7a2
za3759b1b0fa3bfe8d9f0f5396f734e8c96a42afa676514090b5b0d79cbb4defdef6d358962a3fc
z047d727fbe5a47bd5187cd026c6bfd62b130e6dc2e07dd5a54a26d38b8ee1c9cb0a6be448a690e
z526c6ee4e786bc38f87947504c5fcfe60289ede5cd0112266a35524cf86a5b3c88fd522e302a79
z5c3fdd627eac244425bee8eed0ef816389738fef169f885cd36313f34655a9c994b4d559801cc1
z0af436da16818f87c9e8a7c6c4fe3adf18dacd256123c992e1f06cada4c71383f8d5fc7a426b36
zef0790c9e8244362e353b1553212920a83f25c481d0264340be28c6b3d5e5a3b7f38f980e7ddd2
z84aca9b75c4e248a812162d63dacabe8a45575b4af1ffc119b2b69bb31f516e6a3eb900d16a175
z93bf59595b8448a9286dde9080070dcb1af4e937a88d84bd9e4bc7bd2dffb7bf0de036efed80b1
z2365c8e972d32a32e28949b14c6dae078df3694785fe2f7cc45f500ab93ea6d2621d310ba9bfe2
zcb284cbcfe0cb536458c39f2217129edc4a8c90be2294121c81863740e1cb8ecea2e8fd4a026dd
zf9b0234806a0be9a203cd635eb2d89b02cae00d4ffdbfd0b12fd98246c0867520c44398f13d0b2
zb32930f6dfc5948b245cf42531e0df669697f368373e73afb6100f331f5e19fb63c6eacc101662
z72a85b5691aa4bf3255b7d630046ed1a03c01a095d726091868ba8fc31cf0bc8cc2dcde767c6e6
z3308274fe5a35f49a1dc3a3ee54b6f80e53de806f2052d757c81d5f8011cf2ad285795376081ae
z812395511b8c8400b772848850de81f5282a1a1d2b4000bac39a11619d95fe3b21dcb899ead219
ze13c3b6fd8f84acc0e18b3700e68159647344bb77cb9891b373b1acdabd5bb3f164dc2ceeae5df
z9dfb42b97ae9a81457c67d430de7b50ca1829477202f07432f2ee8f0f6a4fdbc44784d0440e59f
z2d15c927cee81bf049ce6b90bb88fb4e000e32bd37dfe9d42a267b4fb38a6e2751ee5493d3ebd9
z6c5e41eeab4341036effd1ea5c81e22076787ae11878456e64ab7a5b2151594abe9c3e02ab20a9
zbc5e3e459c098c9f97790d6b78b6cd6866bc81a47b645da228a7b00ddf64e1164b0b1a361f6ddd
ze6a51838ef92beb9909937a6e26a89f70ae7dc82f762d0938e4f71610d6ce8639d386545b28fa6
z8fe93b1a70325a6ccf135dee2b5f5ace89bd98915e7738bda1809231ea2b3057b37252a07ced3d
z2655624ca18ff45d38a814655c3ff7fb78e33daf203755b8b3521548f1d8d317605d5c48dceb4e
z0de6c999ecf2d30d2146808d5e7c40302b8a6fe034f221037301907ca7dbb956cd8e9900be75b2
z2be47c53f0a947f4c73ab2a7867b2d88a4d63f3749eb61bacc88747b891578800853c26f799ad2
z398549a56d1dfbcf975a9c5fcdb2d4b7242a6f8b699c976730bc6d98f82bdc05410c9f44973948
z6da8acf4dc847150d3523dba9864658e55fa4bbcbb800eaa929574dfb30c77dfaeb7d51b2e0b2b
z846511c3fd871295011e21a81d1eb92fdf9456101d6bbe27c4d8b3ef336a72fd15e3394a4da393
z11e9e7a5fb84f2c540b91aa5df00d830f37afd7822af6bb333c674e93df1635dfce1403db759bf
zded87fc299f3621d9b579475349a5e7758300b28399bc2214127193b30c107d4677943eb176693
ze002fb365a527f3b0c3a5a857a7197c0740a31712084657ba9d31f847d6ffe9475cf3ab301fa3e
z77a5c7311a6e6b1a1cbea9fb9795ba40dc65bc88debc482f664385451cb512a7bd416c03e2f04b
zfb4fcd3c7230921449099838f6d2ebff09a9831799c04d167ce83340649216bf81469a0d158641
zc6327156c2b781cc644ceec4b99d3154159c76156d6fd044d2fdbc7c71622dd13a44c5632af224
z509cfabd1a64a3a6c7f6c53ac71e5c3ffaaac4243a92e7fc5c1af03e6656889f1bc71d90674ce3
z8909701dcebadedc7527d9630fc03e81b6c599851a601841f8ad93ebc2aa03587da07692cb61a7
ze942f147680a0b3094f89177b176431f8492dfd7b464b03a93cbe626b057599b73853c54b7a774
zf63b0ea32daefaf0ec39b6fb0d8f1fd9089510a2f8eaa529ab876512e8122e3cd96a5b1a9a9fbc
z84417cc9f932494162cf51a148d35000afbf684d6d5035891a7165d656a86d12472ec043bb2fd5
z8b963dc85d80ae5de4345652a6ad0c9d3752044f465a62ebb420ee97e54aaf72e483cbabca4eff
z11a470f4981c6e89e096b3622e64a6efe4b6a57b6e813fc1927e698d88ddbd9a3e72813fa87cdd
zbb21aef57eb188e4bd7100189186ef8e7dcc73de65069dbcd34820294639532d687cc85f219c9e
za22a50c6091b9c51424264cde0dcc2076dd6637a4b715563124ec6dbb26bac9e8069a754492210
z3679367d4b8df2b871db618b419f0e2e248172c28f92b74c05d6ff14832c4da4f6c780a695c29c
zbb8e68b39dbd2cf050084137a182642513fc316ff23214e198a931f74f19cf81818db6d75f449c
ze80c01a464094707c1df2651bc2692a9313d2b5b02d0428cae9b724773aac5301699300e83748c
z3b5961f71a9e05ab22c140736d2f425ee7ef53750166b5e5ebb1f6e32f28675acaf40960fd66a5
zdc15e394a36f73782b0d61798a384602b93389dac91d246640569911500f3dc5009fbca7073ea8
z56bbf56b79c88748269f088b4e39ec3fa175d964c9ef6205e70ff760ce0184b280de9c6646a62e
za72e65a9ac737df509b7d2cdc556e6f1a88244eb57ee6ef1c4d4bb8dfb0f08051064498c66268d
zcc67629cbbd934551b0c9169cef46fb75d93e94a3767f3e018226d42921fe1f473c7fda738476b
zb6350ff173a656d62d0a03b0deebc72942aac9dbad9df7f5af0f22c920063f86336daca120253b
z0f6ec0cf3d5fbb4261fe907847ce979dde231e1a4c9461888e9a0237f6c4258a0cdae451a8947a
z98b3a2e203495f19975175e11ebdce07f495f4e0dfb9236230c8c3a2ab286171026ab44b23fcb9
ze88637f30c7045753f05d91692e6ea643d71a64e3029796b2fbf863d53ae70821107c6562b7fa2
z8cb25d54b39410965af39143d3c563d94d5fd80391fbe878b3c3fa5e64790ebaff2524a0eee0f9
z09fa2b14c7182a5ef6737795267f411e617bcaea8e24dbf41c0ff8f4e74241bd830b01629b4c7e
zabac4e5375eff529d8ca57791795b0679615646b5050d619cd52a2f020342a529fcf030141568c
z298ff8bb9f0a0d2381f024233def7bcff8aa99cbe11ce9549d02fb4c4385274722e7bcfaa7fda6
z681f0bfd8b17ca33498379fbaa6f963b2ec8ec56fb5f9c73356e209165d069262a257badc66186
z2d467f5c381c1a700ef4074be12e6717ab103b14c7e7cd3c53a8662dd19b3586f8d62ad2770cff
zbb122db4609600d613a43403f81ef2939bf9550ef8da0e6c3f66a8df0c1393e5386349342cebff
zdfe9474c61140f7db1e2e65036d5b8d24d329e5295e39dcda571fa8423a6e2f9634f21dd99ae71
z747c9da221d801f6be0af8256042c45cfb33633f53f7dbef84999f4afff921aaa565eb106a885a
z490c669af6ab2c8f0b5d5ec182882289628921f5066d373707f1a2abf511c523776df8a68eeede
zc861054f09a909363ce2b7d06e51c51ffefb3e0bbe934ce60a83960373407e3c4c1fb8a8696740
ze1e5e9584d9c9ab621cecfe17f1fb4959c43026d5d6ceb4fb927bd3b2d8429632de329d35d19bf
z404e1830387a8aa81655c7d8bfe40b1a44e8f7281be04255c158aa06396a7a5d628e573cef7d51
z842af8377a6bc40f9eaedeead12458399a624589466f03a17bd2f35bd37c948a52ad64c22843c8
z45eab3f843340e06ab54884946b5c30f3c87bc4f16556fe0acd52ae98cea4644072441dabc1812
ze5dc028ac50f5c5e7683517b7676ab5615bb68b64847a81e282fafda45a2d53600b13d0094b1b4
zb0f6e8c486c97db7a0733f1222389ca7d6963659a488b8eea66eaa4facf1f8cb60f89376edad91
z0dab4a8096c362280bf4da32c50704380f5523fe8309c484073c92cc02bb1ed44f6a1cb02f6335
zd0b0220e7a66ee864e44a3229f47dfc91bca95575fa4916c0007cd02fcbc6b29c25cf2b446bc1c
z3004b8727719592efcff67f512d925ce4f90a14968e45a7604f5a16912b71ccccff041a1994160
z33e3e120afde57d7aef9f07ed7440af59ea4f5742d5b1abe4cd1a32a91bac3ba1983f934ad2a98
z21663742ce8215ee7320bdf5f572150deff69452ff49e41c2f796d2e64e8dab7e0590b4f873465
z5ce8b7c2db0de110b55ae1266e698edfbc893f61f29c04c4cd4d78d00d6cd591ccf9248ca99299
z1cd1c34e1441645af899854a4058bc3058aa3ed047b51628c2703c44003a633b5181eb37b008f7
za8de519dbf7e2ad1c8bd29e971fd7f904c693b7f1bd253abc519cdc9cbc116d9df47d03ba981e1
z194623ee30fbd73f8dceb31a655f208df4811a350e9f4977aeb3b3eb26edad7b73f0421f8268ec
za67047903d4ed5794b33cd8d2fa98012fb92723a4b1e81f1c4a37e7c2063b38475de24943e96b2
z11b962ab5322d6598df7a6948afbcfbeda8662511292cc5465813b2e28e20a4343571738ad2ed3
z0ba882d05b218bc9ab6c135efa96a9cac602c6fc779290ae5da088457ea1c5c4169e33300872dd
z3f42f29125fb85f4247cde53cfca8deddce34f24bb3bf3bd338496e10761c7f2305d8c1dc27370
z0b5fb2b1aff3833c59286a4e27200847967f23dea7cab089969fa92166cc2bef552226de94c594
zb6e5e9ebd979b8771f3680600f15fde859f60901f29270903ab70abf1d5cfff66373a800207702
z63c6476a48d3f0f55b1bf3d90bc1e479bbdae6e1b4930a412573fe714a0f3d93f923a178899d68
zad221aa3ca34902a43bceb705a5ab7756f0a42b2ef7e13a408abe03f2d9a5fb6869ccb170b8434
z2b8fa6e7507b8e473fbe88737f3c21c6728dfce9cc512e7ebda78a8df20a8d21c8a11123827b47
zd93ce938cf6af5bdadd4cdf9ff4e3b645cc77390b8584d8804685c9b1cbe504b1f3ec42b60c56d
zb245bd3bf9bd332b0572ff6b49c9bc608b5b371315409636b273ebc6fa2245bdc9870b58f27a76
z3b901fa9c3a3f840366151a7f33efcea97f6a636f4dadc7f24caf688fcdd2a355ff6ca465cfba0
zf61a720b5d5cf443f31032c96999d51fe28cebca1b579a60d8cf9446ad426fb100e433baccf707
zbd0c70dec38169bf1459d80c7bcd74481adf327c9da0f7f6b5058984cdca2368adc9f431aa8e4d
ze77f8e4f9ae8f8f2ee43115879a677a045b630e6c3e62ad9aa0649c7f5df396711428b7cceee88
z42aac2e0d6dc4897720f67164d5467dca1b70ae24e8d04b6a0e0d396e63c14f3cb75a9c9bb2446
z585576d39f1189256756a0c59fa3a37adce2696a5e44e6a6974ec5a3b1a5e03fa4a700ebf0ee69
z7013799563f19e8ae3b0640ea575770e6686ae44ea8838e6e2011c092d6105d83d9f456da5b607
z9ab50d937cb0738c0f26991e20375d3e0c2555359b5747b81ab42c01954b653535642e3c3b213c
zb6332fbea73dd6a235c256061a3ab901124e3ad13530d3036a3623a40bef986febc58e3de80fdb
zd394b00c019165f38330e572fcd55cf9f5a98744f2b5e3121281e80d0a462ff81a2010c8635c00
z2ed5024ca6e13673937b422ad6be8a3ab1e043c6ed2cb41b4939e53dfa6836e26b19e57ea01d19
z3bb21eb32456c88892cfea9aa051dcd17af12eaa02d7439f29cc1d394575d0188d79891fa7b207
zd031d557a5503016a4e783371b42b2a041ea26cac0634d2976ef11d9330f604e03671ec8d0770f
z25d0b311124e0082fea3c9ebf4a95abac8931653a6e611f40518b6b2f291338a5b2023cd4a9beb
z3b10e7e8f057b0a09879f276938ccba11bba918edf4d2d14ddc88677c7f20f99897641a2711cd9
z48cb65d8ec827e2225326c68f77d4b274383e5600aa60f1c1195ffc2d05f7ed1152c504c5822e9
zcf75d1c2f472e01ab91f8cdc01d9b2dcefc09fa8d958c01e59504e2d2e72725a17c7a4ef2e94d4
z4f3d9e3586892a140513c7411b623a9a25c60ee513b7da8070c55ffdd8538ffc1f9062aa730985
z09064e915c34347f60c37bfb9691ac96e7cda21beb9d00071f4e40a626f459ebe49ac4ceaaef36
z0e1f9fffe3e9e555c9f990faa4e73e754ec9df4272e4b27f3f410d3494f0e4486a8acb320552ab
zad14f7ee944d9cd5a76dee0e29e229c19d3513a9e9778836c947a95f01a53e8b9d5c8bc72dcc73
zb5e460150dadf48bc3550979c57cbdc52b5f600cd4c49d158ca9792c93ee4e6097e829fa427d38
z0e9461047fce5e200f1d74819c3899003eb1ea213a92aa47438742fccff6ddd7e42609831cabba
z53e069016aeea41ccbf87ea98b72ac5ccf858f53a66f235cc9d7d4744190110804608e2bbceaed
zba9e6c0dc13f33be1fa476306aee405f25c104c3806dca87133e1ab18fe78f807492cd83b36a9b
z08f360e58570331334feab2a34cef80cfa9466904903de9ca6a58c3c4e8e26e18f1dde746c0756
z4edeba68fde3b2a9d2fbfe2dd936edbff1ef0eb37f8726eca5e1fb05cc20e2d3f023231c35ae18
zd5804fc6e6f20a3453394543c83630ec8af5bad6dc74d59348a65ad06506ec5f7ea843ce3dcf12
zfca4ef98df24f6e3a9ee1d374902805c750f7d1bc61649b6e889886e6167084b0db7927797b719
zdff6336fb5680e2ec70e1a526551c87a1cef77fddee92503090c8ef821290cb733a737f6a49405
z9e67e1ef72f2f5963dc252d3d8216ed12bcc7da167c6ddc348fc026bf043c3de328908bfcac318
z11014644643fb5f8f6c7a724dde77808a4bd5f80dad33a0b9898bfca117f09c3e100bc3cdc8f0c
zcc0a88ffba4b5c2e3d1e11831c08e737147b18bcef199bf5a2bce1b2b0442821f5e210d3594959
zeb01ba291fc7ada11cf4ca44ae9e707e1a09517e6e43ecec5c1872b81551c4bc96c22530d0a8bb
z04e9bc821b762a7aa0ebc26ef406a65d2a006efc2f7b09bbc7b012d2ece565f7e981d31169cc0b
z4095b3fff3bf983fd393313e202309ce8893722c0c450aebbb55ccfeee127dd5436729b9063456
z311a9e2b89980bee01ae7d7ad52cca912824f36c703e7f644fc518a817125bb510ce4a519413b1
zeccb04102c359b59f68653c290da7e60cdfb04dfeaeeb1588802b3eb41a172ce6c3e201c7f38f6
z394ad22b19b6008fe6d5a1d934ffc5ca9797852af63912515d817f89a01b2a25596b82785298f2
zad370eaf9e52ae42a49e42db920a3e8152acc963ff76c891dfaedc2dd135c3acf6496bf560f35b
z03dfb036708829bd1f7735118728df4f926c16364ec2033ee0ff050844bf22f0912499924b21d2
z0a5f52d0a1f558c60d3fee32374007be336a8a46167f408f2521d34bb0e5c7024829c5590417eb
z48226e1d0784d919c9d3cc07379750ce8bd189a09e0b6542a7c0bcf72ea7372bc8b205d83e4117
z2c5a265c0606fbc64d9c9d8557b1ae6f0989248dacf67d1273c182439386578f6e7b783e669512
z76c7e6fb7c95135e76066d4e4a99432e3377b6eacf100f2d8884bf16e03be0d034e0c3eaafeba8
za1dbe32be99a597ea778c3a14b2b2e0a2a49dc9c2ca8df4fc5b2b8e3e90f2a4a3be9276bbcf7f4
z48b28264c03fefcd592ee0654b1bec73278dbd5fa373314330f38a79a019d23963cbe6b1e4ce80
z6bd5f59d834f1219611d075c012d529b145fb09b3eef054aa4fac079afb22fb7d928deb7811dc3
z2bdb507364a241513c08653f22a4b002ecb16fb30aa179caf1eaeddf15d39808fd1c0213ba187b
z9031ca22f0d890881ba6c2de1c0f3f3fb588d41ec061322b9a2d6a5ae5eaf1caf36745c2df0f7b
zd2d95d0262a1e922247811730dc5ac94e3d09643a98ab2937f8babdda25d640303ad7fc1d6e61a
zb01fe0bbbb2e8fb4852a7b41465ca577603837e42b231a3802d5930631c3668a4c45e3cc78bc7e
zf360f7572b5efcaac8957c71f242a2efe1b86216ce502069b9a34245003bc82c896bbc9c870638
z7f0261dd7873a4ea27c0cba7dcab72805ac83632c4cc056aec2166e9ddb587df942e89abaf69cf
z99d3096bb2a298ae954b2ff80acf5b150d0ac397f26e38d921cd4d99dd2a9ee88942c5feebc653
zde56db832d86b1f678379dbc9f49bf81c6562b219a23868815dd03898cd0fdda9dc2e3dbc623e2
z57707ea257faa6cbda8af6c5b182fd049864f2869d83f4b5839f8246cc5dfedd2b7ece96c27eea
z5d82034fc8a4c774b4ab3a3fc1ae8fa2e1aea741d7a58d1e7815cdd520b9c23e9ed98c188fb7fb
z3a6922e92f248f554474c4b8a43c0f2b79ba465b2aefe30b21da270ddaab544e7d41d1f7b6cbde
z8e2abb9dfd58d195a1d2c3711be1b9707e1835c93325aaebed0fa96d7b4306b92834b5e4f497b3
z9b2ae608d81802750b18ff7bbd953cadaecb845678e0e6781efa8e93fa7824cc0a87680d5ec03d
z37f996a6d0c621d3d10586174c74fa93443522dc15122ca1263567e64966a2ef72b78f0ec29be5
zdec8391ad1e5482b5f104df7d53d14431aece448fe256cadf61be2ac2e82af9fdef35e400c1588
zbc2c94c8fdf00d63b4b9777f6faec328abfaf6a085a896160f3491eaf3d6ddaa79e3ed16f448b6
z55be39946fa520c94df27280ac0ac4a0549e233af23793ac78b5fbd515a771076fb210819e84d9
z76cf9ba2edf1a14ec05ce5daa81eac0d368236fb9273fd7a0c72d3ec69a564dfcef45bcb560a6c
zf6ce093a57fa4658ee05e22bc4be2328d5bbf21013c4c52fba727c9a6979f448e19416f42a882a
z19e7161b061c0b5212da33d7e81fa2d8816017f44dc38f107d69d66d9817ccd89f2436878fdb6c
zaef71ae64d5d6dbcc90261ebca11c6d9e24b6a0568a1d05fa07bc8dea3fd30468b8107c5abd959
ze53733f3eb260fa961ceae24203441adb5268092234798a9e18306cb17544939a1321650490b7f
z4b38323e120529d671cb98e1ff8473d5d3c4481afcc02be1a5f9b52f6aeec2000f408dc2d3dc03
z82e5c89dee91a590bd7bb423d07c5819e6e82817ac0e9e3b112b0a97617be7b91d41892831f9f8
z159c638878e4c1610d0e1446a13f96498a28e54dfb5916bc7032dbfffc516a0690537e4a0da4bd
zfa411b39708f534b89600ea6a160c341514369f4b547c577d06f59e9fcc858827e1c3404ddc27e
zd79444233d1426a1c17ee4a14cd2ecc530428cb389d1eef5780ba7176bc7e4ced34e085d3e3103
zbde1b3837b4edf94ab51092e087e5d4afb157ccbc8839c7f28e5ae09553fe2860d068d793dbecc
zf3bca32bf88e06378b4fc274fbfb82faf50d6be6206e008b27312c66abce92a0bbf7254c239404
z6f9af5fdafbdf110dfdbf187267fe2203ec90f7aa995a43cd875547337794cd4d326bb581ec60c
z7f0d59b072c6db81dcf37e4ac634d7c5c289443297bec5a4622df7b8da58e8f81528e4d266d5c4
z683ca712db06c2209b1e015d2b6585465c7db19efd0b3d1a90832c528158fdb5cab9d70dd65e29
z411a0bfc30169c20a38bcd1073123b969ebf44e3a34aee120cc400e6d40391020ff9118311ef94
z66cac633bd0a5dbb86f8287cb1d41913bd07691784c44b32ec9b6cedf43a38ebbfb4f07413b518
z6dd27065dd6849a77033c231c1f6e2bdccb0fe24569c96159718f3feff01dc900b8659b744a10b
z7c837d106185a06c0bbb703fbe5077b7c45009339dfe984e9e3d6ff44fe74967172eb81c4c962e
z529067b65425596d3f9f612108a6cc45441c422599d0f29966e97922d0774c1e10947f6030b14b
z4b9a96d404402a217ec37b9f46b1f44253258dacd9f7527e0cf2f06216f556654f46eee1445747
z6bea30e5b60bac6e7cf2b39331ed0b5e52304d65cb322c63ba7ac2cde2dab8b8d6c5c4b67e9bd1
z1224bd888da51f3d98bc0ae23705d54ba8dea00d06ec5f6912c48cc5cc470a4e42d345b63f09d5
za8525b0337a72a662fe0f16eb8f2aefebb9b4ee7e7e7d59621f6b2f4cf4403562a00048a7e0545
z62e630a84812a61a264b0ad345fee3945cd79955769cee46ce43c649fb26f8c652a23ae924cfec
zc38d33464457f10c36ba1a126dcec6089d19b8ab84eb2ff395060a18571c5bcf8cac4ed899af88
zf6a43ea4c44668bcb6a179244eceec55996f3c147091cc780f1468f353c6cab4dd8838fb35f40a
z05ccb6cbd0948b7d544cae4def59d333c3129cfdcdef0d532251fc144fed0428a91cfdb5d33ad0
zaccd49b53c74e1af92ac8df1aaeb459d602ef1b85452b6d613b1487a8e6fc7587e77ead012df10
ze8ec311c51b94813455002ea5d60d786a4c3c012803a87fdac4215ef5cb6b86e2ed48ec89ddd43
z085c95ec699312a600bd2a40d8539322ae777dfb30379a60e9263c504f64b2bc4398a4e6dd90f5
z47efc4e99c71ead64c7ab96e1b4a4ce13b4132c0471b6d26ac93eb6e5b5ecaa623a27cd51f7431
z39a9143c7afe14d3fdbe1d566e3551760fe7ef71d82be586d6aae61c9f0e86dda40be58873bb19
z7a36517d9509e03e65ce3555fe1e3cc2827e635ce0115ec9af19ee10d0396993126c5ef356c724
z69f8dc981102c3cd646d6681ea772ead3e42603e8b64b9056b65f0f80982e2964d4f6848c97588
z90b6b533a4852bd78d3efd0ccfb7a37460ef322e3f225b40bcb24a6568acd7ea3592651fafda5e
zd1e3dc7fa9e8a0cab765dbb86d46751957a9699afc750525c53e8cfa6e04400bf44aad2695a7af
z27706358ce1bbdfc0a97315f932f93de5d678e7f326d092ce660001e33ca8d7243be675b451063
z74621e8a54810546923177b885e60d49805b812b2422eeefa0c948dba3984d7df7a837f55f3fe0
z9a0d50eec48cd0178c8041d2304993e0036c18ae5a8d1b48cad34162dd8af446ed8a22ecab38b1
z51ce209dc9fed793b6dc7a5769314ed2241211b6e32c27108590cf44116fef0bc7dd55b01a92f4
z7c66adfe490b7c54b05718de58278f598794f5fa3260df8bd10669bb00bbbde4869173bac61d1a
zb0ca8719c3f946676d628ac3acacbb4867060472844a95f0b9b68923e43b8cf881361aa72db792
z10e3aa62294e348b0e077bf2d2f2185804779837f82cf3e99c1eb2c7c22b802bcfa3efcf4ce2df
z9ffc9ca694b3a0a9ee510c2c99d2eeea7cd93d606e35a6903d5925dc3ad8d8d574ac99d0d1e5c3
zfa44c480eb3c9932e4133769b9c5029c9f07cf3e62a15bcc1b99bc1f3b28a5b62f5bc15a088cae
z47ff277c9cab4a3e2f0fdcb923042473c26d4cf86dea8237475b2b1304ed86cf543aceeee94e5a
zd0d7a525f70e375726e66d30d9a9a105a9180cffdfad7aa2d4f6ca53056051b740c53db0aafc23
z3d4de9db0f24ed3dc6f038c7fb6fb3417855ee960dddcd4aff6a922f0364d11a07a004016144bb
z136c32bb188ef4ce85f7df824897fe21af07061e7adb0fe34cf411fdd754b6f814c64a573eef1c
z28d1779f2d5c8d6a1ba39fd3d7eb7783516721934171bc26720a023ddf9c28623b4ec17ddeb264
z9f92f5654d58d49382c4bb7ee95f7aedc63ba17ff597f554379591f18945740afdfd67ba27a742
z636119a8b3a2177a9bbba68148ef877e96e00c89fc224377b8f20ef840bc8809d7e81fb9d74ec7
z9df4dd0d96ff9c25e1d2c7fdf5be489fff0b6ec888228c65314b9e92c52c5a143cc97c1d994f9b
z4928cb0d4855faec310e8cce608bf3c939d0ed73fab41fe6f80a02957f15015c23f43ffccc9c22
z1c39dcb4f233f398e548d7a2e8da5b91e066d25833f2d80d3bf793095670e3dfe26b94c1c83188
zc7990c39568f89a621fbee76ab20623945f51abfdb8d8b6a960861f2d4c9aeb4a1ea965e953702
z30d9003c156192781d4d669d959cba064371a60b233ea71f6be0d6c1b620ec30d548bdae726237
zbf64ad52ad50ff10ede408c99a66277c1284fc0e932c9e6a46100c4560e943a8523eadf5e804f2
zdf95476a42c1c0aa7840c42714d1d390b224055335d53154e999184b2080085d9dca84bbf16b15
z449b1b4c9ac7ea2b6b2214f646bb02643cf12bb72450a8e28ac0cd26fe8b9c98096d13ce21d63a
zc3f864ba4aff82009360b6fb5941e01b1f7540a0fed6b61ee5244ed08b2ef3c7a875ebd6c7d967
zbcf5ddda30fe2c52d597ec998222e93251b9ac932e8066aff7b953bbef5da473a2ff14e073395c
za4a149f1eccc347e7e23dabb603a7d8bf4dfe8db82ec9f8ab77e11824dc96019c58b653470448d
zd290beacd71719ecced8f68634f21afccdec6784ad50e8da85ff717b02a4851bccd54d188fd889
z6b02c711b974b8e59576695e4b7720e2bd4bbc372e884868c71307cd63c5d1d5e40558884e66a5
zcc38bb08830f58bd34a564948947fa9700dc56222819b22b42eec85ad72d2ae298bc55031453f1
zf69624f6ea2c9cea511dc8179826dd7df1547296a56e5381c45974855293020b3b02513a6b4cc0
zd6230c5eb6f00afb00bfcc7481937f5283f684d496845e72a672c2bf9abd3911d97a1bb5b9a125
zcecb1e19e1cd6e8415642e8d5cf684df4b8fb387b71dd5dfb376631102795862f22f7d0fe73dcf
z47bb340d5f198d173b1d0e3adb43200ad57d0d0b56847956c2cad5800b08a0c9c40a74965a75c9
z77791987ab2bf7833cc69cd4d2ffd458f172105dfff1b64c440a90569a6d58134475fc9e52850a
z81fb2ee17d500b9b1f25ffa024e7b0f0723b6e2bfedf648aaba467c21dd850824830676209c8d0
ze9daa790a45183a0c98e6826a8cf25d627bfac3636ad08f6ec33ecbd4949db9a1282f036bc5f82
z8896409f47b5ae8fd55f11ba1133b94a96130817d1adf8ca44371962f1d8b0d981ba57bc18c0d7
z98971865ffc1c039eaeb3fedd301d755e9c2cdd499fdbbbd3cba014df1188e6491bdf51a37f036
zaa9735a165abd0b552339c2c0e03ebe8d64540082b53f17ff40e7a855130f4234d7505fa52c14d
z31e36faa02e13a713fc95399b421b412f4ba620afbb7f8ba8907bc61dffb18c93f790688c55a95
z7a697debc1eedd7c102abbb3620ba6407592d699cf3deaa5747bc5f03ca98c258806de734d99d0
z6e4b9b06ee71c2f037ede097805c5ee42928a903f278b2eaabcb5d006f1627db44a1491bf395a1
z84725ea9a8dfbd16e1c0cb7ae77b668e21cb240627b657f1b80a21ffe46ec1f2dd6bcbd4cabd5c
z9580c928ac12327e850652adb7e48c33ba2b022de30be984807a05e403c543dd72ebb9360d2d1a
z56fb52a10f495f87ad5210ccff5bd7e2a4e354dd340278d364e5e9cb7108a5f1b4e05af7a83493
z468e74f1f41502e9888fb1371394a2cb5469aa9a6851d6eb48d4a8d435502e0e66ce9f72946ae1
zfca26d5d14b92bc64672d9aee32e4af5f2d25a51af0beda887cceb901651d06c9f8dcd5911588b
za3610d0e9b5e8d0cb22b7cd148c8ea716d59aa1452befa075e9146b4f5fd1dcd1addad14783a72
zb8c9cdf79bb41a956a794cabdd578061550cb899ad1774ea41c2ccdfd296fb5478b29addf90ba6
z96db72e661f9fd2e496a24d29cbddaaa15840da376f3c48173b236b148c418d01a1daca4568634
zc4ebff7037b276356839ab0ee0acdfc3e8be10761fbb33d8f261bf8af83e4c1411a1433c562431
zaf1383ee6ebc9df58005d3b37bfe08f7a7434a4a86706d3290081a67a56815c45a600fa5cb9f29
zbd764eaea130441d679f150c5b7156be05f9b7b4b89df8c4cea3d6298c6b80c0b21cc38f296b36
z05d520a027027f4503a97492d72e420e69e746b0cc0342a03ddf640b72e2fe538533375cf24597
z90b8f54414fff2914c785803e7730939c6b800cfc78a334ba5456902441632801ebd611a956dd8
z986756a734a5e04f8f56535e68e787570d739959200eed30fc7fcf41a54cb64281a41943da6993
zb1b125839054fdd3153ccf38515e2a49a0758f3ecf4353888a2192435bb4b7426f951d6cd1abb0
z85a78d021d10cf8463cb9ad9bcc99d8d938e79e9689cfb2543ad8ea5a78335cf90516465428228
za8b5790f586859696b9b37ad8141873b373fae0b4d54c05dd1116bf44d1aa98cb2e458522bc358
z4117ebd7a69bb42895895b3d57d0ed42f5af4ed2bc5a2309037f233b8fd12987febc449757d501
z1a8c7e49186b662ea4a650073067349f18274522fea891ba4d3b79b48f547e5041f6724bcdf4f3
z4363d26b804fbfca43222d4c405d71a4c4fe0cc90967fc7b559ca51862a704b086ed38595e171a
zab66d025363331e82bdf1f357c0963ea1dafb6852771356aa449962914980adf9a1b316d7ff268
z5f36baaff5d6f1030ecdfec1df14241443cb928f394323ca55ca4eff6da635ae69ae93951e7c21
ze588f7a22d96eae23a610571d8cabe3eee9b191cca29fda45dc0661873623912171022425c2d5b
zd3f6d8272b2bd4d3b88d6ea0f97fb5027a7bafcb469dbcb4fcd8d371d14e99af466f7488db1e71
z92211af95480f76561f4ca39463873d5bf6b7586d5f18a2104cb274f02314582e72660d339b434
zf0f9e5046cc3d434033f65a9e5bce5ed498ea32c98cf85e02a10c153a9ffaa6bf2109a6b5035b2
zdbe4146b71f674edb759f8e9258cccb62a7f92707693f835ed3712e387ace9c400931f14ed2300
z6b26f263dbd46ab2443729100828ac0e4356eccb5013ce90bdc982fc35024fdd9619f7594b221e
z28fb1247ce96dd7fffea53b5b0d24b729865208aa90e6dc7a1641d1c5830af52f6ac0306f706fc
z2b29a62ae6b43a48f38d550970bb55a70ba2b5a639747850495171a0a095e8c2146184ded47a1c
zbc23bb4d36f810899b4c238e91e548377d235f93c76d23e0f9a49bb2754d0911f0d46b97aaa4d6
z96feee30359c67507976669c68da6a2950ea00a592cff8527bd11546ab3e37776c349d111a5c93
za95c147c162bd4912cde593b7936c9b075f11c6cd11518b8bb294879eb73411e107523ef957d02
z7db8fc4b2e1003f728070306e6e4dfda086613b442f2380eb265bafae16a4648c94798a41da82f
z2c89b9677324e90cc7f3e1235a1bff185d6ab7b6603f38e7b2ac18120f5567641f4a82930222a1
z1e1e4f5ccedc9704d068f8fc43e0f9944d5bb9b95c3cf03a618f5dabcead71069a89468239ec96
za18267945fa719724195341b0e1a451dfef5e971ffddcc59acd95ad1a66179c6236587813d1611
zbd72c48af91f8e00a7b95ab96b1359fccb1b65d6277b45d7a5d4399d891fba0fdb28d96b327c17
z57bb36c222bf003b8c11700d02ae0a98049e990fe82cf65057a385d970292869e6e8d4a8b8a906
z778ee4cd745ec5ba3ca1c8b2b34e6ce404b48fb9de965c456a48ed540b6ff4c34ee303633e9b55
z76b4beb39caae0e3f90e8c3c5f8fa09d83c116b482e7282acccea26d341bcbc2e69cff96803051
z1712caee391a7f1f9953f6a7355317b711652360742c841dbddcaa09daa7dee7da47d8dabf3e7d
z32ac5762f17939f328bf3e6a8d2da23e1b535700b517fd0f3f3dbffec752f7a9738417ccdc51b8
z70ad4ad82232f8ef01ab14b7d57626fdcffa906776b35c464acdd5861eaed37b5b4c903989771b
z2667655e0c40b1a523653d01ee8e6a43d84dc8f063ad1da7cc974e955f5655f36692618be0fb7e
zb0b9f9776a45fa7ab497e00bf0c2f57acff5ca68f8415a5e9054470be2b6ff1b64427b55aafc43
z819f6ecd22f49c9e436ecfee6911d7c3ce9d81ff6ad3fc035cb244bb4dfbbf34033229f904d582
z9fd05a742a92bde1af04790171d7c9a475c84d5a01cfdf8f8c9dc1f029a8888fef76aa9bc89a49
zce4cd1ffb346d5f4992f8153f84bda0176fc29b88b3b058b2787aa2da63e4bb54c9c8c0d7bcac5
z715c67c2ec8e18061a9933f756357a93b1e9c7f1b7237473c2f5ebc1512cefd465ad6ba3a7a153
zd78f1ab24b565292330c81212b041ef1c2cb14de34c017d27741504507e4a063e0abeb8af09599
zcde3ed361fbc10a73d6baaa0e23b6dab494da646ee6b332b226e110c68c23095e05f2c6e5b6efa
z8610a3405756a00593818cb7dbeb056796217b2594920d2841978354f9739bcc9efe28b267bd43
zeca357677b422954eabded27af880adfdcb84c496e9cc61bdf4b152cde108536681010f3934efe
za521d2f34f38734ff14e0404b313c7a0262df1e47a7369e85ca9d240af886061e5859adf51923d
z516a94cfeb27316eb26fc2bd57bc04092ba5297091715aca2521de26c146337a85e116e1fcd2eb
z0b154f46789d01bc10f65a9b9ffdb7cd6f5bb2dd0cd26f771c39cd5dfbef9e8ef3b0dfe7afe1ec
z2dabe6c35e44207fa0210e705222fac45d405ea3e49f869d37e4ecfdec58944b86da12e9a20e41
z0f3c067a72843c4c80086726e778ce92ade4016fee634f6872f0b33510d0ed3e4c1fcf6ba22e3c
z84b944ff4ce98d1e9c600e2a3f0d2943c77d99396e7279dbd93b2c5ff3a0eb933f678d956f6380
zd6b3e5a54dce90d3a504352b3d27fbc2ee1294b3bc4ee1365bd849bcbdc0c2963f7e349c90977f
z04bc42605f36a6bad300e270734fa16e2f5d69eb21917e21bbf6fddc2dfddc5ceaa7802ebc95c5
z206fdd87d1438070217b8d58de675aa65b641d69c48e514acb65839de9314622589b857f794938
zd79dce0383be38c8afe451cd1e49281843317d025d1a28386028eb80ddc492945c2089825b29de
zd071d0132613f5bcd76db83997c0abf7d75cd00636028347e9a2c89138acf3766df65ef7e74d5f
z32b96e8f0fe04e8b56b558da6a386e06e6eed89e51678db3dba0cd9dc26859055bc97347c56494
z472c34d7a6284db2e18fe91c7de47d605d9b08206167cfba53050cdc2b67d1a175d90910445cb2
z54c35c9d939a6a30b19a32c1ef9d8253f3d047f6abd0a629cc03bc9870dc8631e35bf306efc04f
z8a82c7d58df97e7d166e58bc45db97c1ba3e5cb0362e95f13d3205cc79a7e871ae6b938b314e48
z9ad2c1e980249b7ddf0a8de649fcd989cb16cc3c83f774f983d2dfae42b921bdb838d7e943d88c
z7d1be0db45cc26ee22d5e06c0bef3650afae6d42efba122a9f9801b27bbdff3baa020d13d9a51e
z791aa8bfc2693d1bf1fa2610ce05e2954850be214d82554e68d08d2147e3352b75ae8a7ec92518
z5039817b8fbb8d3c310a7a16dffe8ec3a1c46d20f22127e7d6318f3f593d396d0e6c4f48a7382a
z76a98842e7c31f720b0d462eba8f6e5184133eb4f45d86ed16a68225a11a50adf9c5821baae15f
zed1bd5d86061db22222d9d305250ff171cb7ee50d4a157faaab9710b8ce81fee9c683bc17538c1
z8d12b2ce4fabca2b3f26fa690dcb8e1b5426a58aa6a0f3076bc42e480d67ed4a0b907818b628d5
z421530fd49a53cf03935aa06ebf5392511c0ca132a101539961a4534f2e077f27a8d3e3ce66f84
zb4a4a96c7cde2ae81d64e286a08f80b710094b427a604a8dacb2d8855ef64c4c8e5d16f3b183cd
z1585483f3c48a2d17f46401a62002fd0411a9e6427eacd6b91f95beffd93ef971e5b0d4e705ad5
z272b2cbbc07d417f7f6b85889201a05a7a1d3733427fef052a4a7b9b064f5e9a2b5ce3ca1ead19
z8108f8064deb25d7262dc979de93929804a24278e803deb3d6e9e9e2ba9164011d65e46847f0c3
z4a5589f74f1702bc298be74477ac99815a1ca67f4a8202ee89dc433e22b3c8580cceeec8fc312f
z4b2deabaf2afe2593c8f0b1d895173ad0e6085a3d85ff93ffeecdc9ee4fd2be48f702d4450147c
zf4254377a510fbd75a9e8fb25206a068321a367a5689af98255a96f8fb36d1040ff46fa370d440
z887e8f9312246399db3690eb32e701f35b3aefb9dbfacf711a2ec5af760ea9916312bc12ef7325
zfcbe7532e61df65659d3077e131c863f676c93d9eb06deb0e1ad59c2f434e22ddaab4c3fa21e25
zd280c78c8d3f4df32328499998fc60dd7f1afbc9020415d83903fedce315d8f4f33adf7b7176f6
z941566cf2fbc323207cc37771ef4e3d5b94df31b291a990998d468f75e0ab338a7d06697efb6e4
zf5c9bf634c5350030c2292c7f4dfce4364db14f66411451ad6596b2ed323c35b65b48781d59ef7
z44a1e010b3245ac5e0721aa8828d3bca5450f296214b9051c62e86a6cf1d19bc90d135c0ff3549
z9eac9c91ed2108a8468cba421423e877648fa17ddd0525108d42f0cbc6be3fdc5adc878107828b
z4bb493d1a7a25f6b75b8f01ebfd4849eb6ff00e10a9ad707accd1ca046893b636187e4da8caf80
z674032093b6212baa170d5bf43fd8c0ba0418fdf246b015947cd189f75cd2225d76e90b49a03b9
z4aaee374d03884c7aeaba058354f747a07e80fb1485f615eb062dd9c801e05ab2fff9bd70774f9
zba21fa06d4b630fccb65a1d95361f29e6e6d71712921bd08bfe4eacd35820e10d36ef774dc1283
ze47b258a8003692eefb0b70f24ad6f18be28f2b28ef6b7a3a3e65372106e1a673a63b68b70ea66
zdd7a7f7f01960e5d7d9a7e18e079f190bab8f30cf75d00f349e8b515b02310c348cb418b7ecfff
zaeaee896657956420a64c192d5372ab4b05f0bbd945ff5d38274f0b36e9ff3d8cfec94c52d053c
z47241377b6e89b547de198ada715f352378bf1bd13954c52dfc9dce20961963083782b7bc8de33
z4249fa417c1e9a7ae1813f7957398a604bdac50eb96c1afca5ad847c2b0a8bc8d9ac4222421c10
z89d12972ff195bbbaebd5ece21e1095022bad9de340d8abe18fb0864476335a81fbcfe42107c02
zb48e4a4b619019794d404c531616af211f751fe0b58ff0c376f5676e11982211603d28e8e3d13c
z7cd02524b476ac7ba78bf7899530cc9235daef3b545a587153fa167c28f6da0c4c3f6feeaf58bc
zbc0d945a753f88e184ca74fa9786de8c4d595d53f3d9b09e5736fa209c9596152555d19eb68166
z7a355bce5b48f37251346e633c09e97f7ba21316e884d350640d683b1da900e087eb5ddd075d3e
zd64a5fa9be93258c611a2f313615d73e5a13f49aa0b7fda3d6bf4d3b8b1c70f849157d0951656f
z387f37a69c17c3600d89bb53b0b34888c5fcd868a6533f2221677642e8a3b2e9bf9c31237ecc16
z12ee58e5c1911d94a3daa027f68fa830e842c6382f40092bd1511fc1d1cba4bef4d0dfea7f97e0
z85b068574a21932220d69ab943590d61be23d039bd186aef41264f837a66ae3ddd7980f314922f
z6d75b6d5d60cabd5790c5e11060ac0bbcc0ce8d213cd307445a1693c21cefc26c4e6892f3c72c9
z5d1d985eac8263c7aa84788e242a300abc9ef72f988f734a40e45ee36312d89a113ed2029427e1
zd4a5dd317720b0ec4d60d252c2193ac72f92fc63875ee6b0b5c0370d6b35dd90e0a9a07a704459
z78de1be36a8e7553aafea49da303e85cda6c2fc5638afdfa293b06c551b5db872cdaa93b080eac
zece8253929919c2937cebdb806d07b60b0db3776ce82e9cc58f477938512c0cf45afd5adb189b5
zc14abbccfdddd85417cdd2279b149320b2708a44d9aabb7e47656e4f941f6b79eac268e954763f
z8610b505a2a32e521b0e1481214b194c08ff49eabc4629f6f3dc739d9c6540f537879fe841ee7b
z5da53518ea8e8e7e21bc5f8519742c02d014cf17e724921386e41cb08fd85534752802f6337a8c
z24eec95151abab61606c4e73883879cbdd9d74a2836659301dfc8900fa86caaa8d80eaa1f23f89
z41cf3ef3e9df7eb503a1facf59b0be7268e84a2a37a5b2878d7f006c130e1f4269ee2d5085e3c4
zf6e629d3b5dff95232aad4cec206a7719675aaa2739735ad65d6f3917cbfa8ab774f71f909db24
z3271a9b688d0cc181b65d70d9cb268e7384ca9da966b8808c4d8a87b6a7ad2eaef1f9d5ac1efe8
z2b4d909d11a7d12edf152d4ca7bd440190696170d6f923fe796db64ab3b3883fef9edd33f05a4f
zb8d9cdfe096fdd02d33895c925715ab73b834adbee6968166da69c9fee2746c7511faf7e09f010
z8d984e45be53e67da5d9eee1cb31e963173c28fa6c9e3a8f1c8273c4972d926c7025baa1c97e35
zbd18c09af6e083285a3736078fc23b29b19e983040fc9046310994b4423674e6393d7f8d0ebd56
z8a34f3cfc351b2e1e9bd486eef8f569616d560b3d2be34a2681c0969cc79d5fe2640318d80ea68
zbe51dc4d508d3c6e0c8cb2f7947b6e830b8aa51efa6a09296392889cda22066782267a9813dcfc
zfea836a6c5ff837bdb570c2971a02dd1af756124dedc223ed8c9093aec2b27b2087e5bc07dfcfc
z52e5b0a95b5e6454a191afe5258b0507ca6fe53d931942e27d20266414bcb4fed63c1bfbcbc9a1
zb76f58fad57284e11bdd931a24f19cf8519da750f25c7441846a6cdf06742233ddf2fb01123c5f
zac2d841b970fdc5d29f951958a5c2451ceeaa0ebc69132ba6132cb62be1ec6c052d9474046a76f
z96ad14af2958d8e86d200a9384b3c176a8b494ea37499d2017a589344f6a449472c246b3355a0b
z21c8a3a639b6eaff0d23af20af4e55d7b50303dcec7b69e11fac150976e17b8ccc5b41a5b7be43
z3ec6c26fdf68ae4b8553f323bc60add79a896842315181099ebbb2e8948ae0a35667e39e06dd44
z3628cf972290b620e0f694eee9ee5e0b8734e7c363c7eca2a1d2c720bb40e180ca89ecff40a599
z6607cda81ac6dd7599c5082f8f836c30075492321e3fb5f14e385e68a085ec5b22c9263cf54d20
zcf89d2fed5bc506d9b8310294b23708fd0902e9b5c4f5765ed2c641bed83219baaee2b21eb5890
ze7424662f53347abc6b6eb7e93fc00d18ff2253edb070c48f13ccbdb41ed5e38320b3b724a6418
ze71ed6c33ebec54df43c8c9c990f2c8fada5660db21dd6bf6a30b439b39e1bfbae9fdf4ff16670
zf8f73dca78d6584e1c68fdbda7fa19e62278ed5e878a66041fc11b1f23a18206f9464db7b4591d
zfc8efadd5fa85a9f48d28a4ac6ca4e369fc66f68dd1021dd9ed6413e189a21f5ba2bee9c74db1b
zaad14d83a6ef85b77d3ea6517e2ed9fb710bf2b1c25da4cd5d75d3df35f3687b04a429e158de44
z0c76361fd320b6a5d261c349dd07c780ae5d783595c074f8243a1d9e9e596f4dcd05e4eaf7886d
z7cb6ebbd1b174532e19805a5a186fd7bdb269c2aa2e800654fbb4689e672ce24a12d4335111236
z11fc066143528d3db00948ecb93b72e730e4e886c087e13204344558bcd3f0667c42f72d15b2a0
zb31edb25b8870cef603480f0f080b298557dbeb6eff4f51077efe0a37a202fa181c40971139497
z65eb96df0f1aa60e1c97c6da94b3a2ef88f06c835c7820fd9399c614ca9c2d6ab512d46f7eeffd
z2cf933a8ca42dac6ddbb5fb5d32c91ffe96cbe31bdfbc0af4dc31a482770355e52c4b6207c52e3
z4ca7d603b3beba074d9f774abfa32780c0161bb9f65275c775fcd3b95e6b258c10364e6d2c00a5
z5d9cb150696e25cd01ce0c299ee62cbab38f6f7f5d75c19d37dbada883cebe5f01de8725746985
zdf7ded3c64dc8304199b2f0efb17113e8b1e38962c32339f844e64bd9db82b44afceb72872bff2
z950a7a910eec6b975af0466bddbfe133a27643ff8ccdb1b58b7ff8d91864f7e9be30a42ead0482
z80d34af5d1095a4e73e248044bb7435f20513c068033ba7e9eed20ead9eb0d215f34319ce905bf
zac01cd38b945eee31b50d6a2b1ba769eb2e1980ea5ecc0f9f7661b1189681dac29583ed77bef85
zdb69646480da0d8413fb7d7bd675a81e3b7b9a06faed5e3c97a2409addc5a5974453cc15d83319
z3c4689e23f34f9dca4a3a16d259a0c5cca57e3dccc407d86fd6ccd2c2af3fb751cdc1c0d2027da
zb7bf7830130c98dd8d7a0f5a7aa2c0cc49aaa24cf8e494de87b2fdb6a52924545026861789fb9d
z86b051b240239136d897707389c35a2bae322c1ee33588beee4ef9312b2d18480092e073cbc642
z5af8d5a969e1c967e47df647932eaa66b1a52c7ee7496f7396a1788980564ae2ab75a56239ff9d
z43a6a17a299bbf1b7eaf5d742287c11bbcadb59558feae9e481cd036fe28e40ae31df18ef7a477
z09b1fd41ae6dbaec220f4962407b25744b0a1c196299b3595b75c56bf5e7fcb2971192041630df
za2e97494d6a84e4e95fa426250ed34504daa648c2b904a46035d50292fea06ae33738063e34ab2
zf90f48c262fa7aa3b770ca3b00eef6b42c61d0caf4d0f546e671c0d638f2934b42690a29d7f330
z894d8b2ca04deb996de390834ca88e69f715d9c9fdbbb9674bf0940d1a0fde89f066ddf0a14e46
zdca7e6c37320cea7d05071d64e4f727b0b6675fdcb7abe0c9d53bd0e9652b921be84e0decb0acf
zbed7d5ed3a0977c4f0783edd0d6c97e9437b3e2328871f3d65409883ec7931419c1746356178cf
z9707a2be5eeaa855580397fafad3a434d127f3115a63bec9480be47f92a837473b0d8013b49977
z4c78ad9af49806c4169563cefca2f2532a6eef81fcb457f1e5ed3244430d451a6064b2a2ede76f
z7fd2846c90c9351a0eeea0f8c70884f12e21a91f70f63420adffe4059512cce8f73039481205e9
z68d8c671c29c4a20f43f08fb4a5dc27367dd37e2e8eada5c48a65f40dc9ce7f7094ff9f4f83073
z66a0f6f0d8c42e2007ddd63511c1e256b78ebd8e88f084a9a6e86e2b8b1a11bbe5cf7b4dd72a0b
zebd4780fc1c8e73060dad06ed10fa393a94a29cdb86edfe1c0b4716ad44cb4acdae6e99ea19ad0
z5ca7272c685787cbd62f69da8c9bc3ee55103ce04b861df061e0685ddcd7a3c5fe95608544f74e
zaac519363bdcb436cee6406516ea46da6d77550041133ef58142919309d8481d808d8acd9c3a99
zb80c93f1056abfd8e07a45dfa915e4b413bfddc0965759cecdc67f7a362211bceac861c3574f92
z3dcf14b026afb5f862c15126bdec9fb3a30e0a1b999eab70e2222c4ca558ce9255520af77b9100
z3cd698ac79f9b4365be9def28f55cb60e1a82da07c3edd6504c4f4b3359575a89407284c26158d
zf7f822c635e019b14d809e35b05458f0bba16c70d617987fb9184e8bcd6d55d33215525b56fad2
z7b67b7d1252e985ff5e8a1419dd39568f5f78a378e7042388c798cbba0e042e2145397bebb231d
zf37a68f4891b707111c0b49c1fdcec782c92972682afc915ce4c4cc5bd986256b68b69a3b7e099
zf235622c66e92f0abebc24214351144130314487a3bfea08259467031697ea88bc6d38ac98b239
zc233c37cd26d8e82609ae74339d590d123ca55ab24f386ef5c86d34efb6ffb8cfe97c5c9b630a9
z84a21a396a4b3ce8b2fa32d59e5c1027d5e431f0511f7771e968af37520a8523eb4e1d45166a2d
zd2da8bd5f92b7692419f7c0b8e595b5829935c10e69e8425a4bb42fbc0e3ec354e5077b3d60d51
zd76c25ea3d8174aa987efa273dd1e5eef8541b863d8ebd1fff426bc4db504794f4f0cf5446c41a
zbd3ed6cb49c858e4271b9673d131f64f57ca57d3036144124bd4eeb43fd9ebf46cf0b361994193
z4d9771dcaab459137993890d5cf9bb5e0a365dddb3ccd04e630e8790f39650001685fac513ade7
z92dbc4ae7b127fa3e5197945128c9101473a7cd10f2d5af072751b7380dcfe5a872e07f589a131
zfae1849d0fbc15a180a673b669d40ff1fe6ded24a7055f1f4632d13061e4e58ca99a1afefb2e29
z8f92bfe6e2518cae7b77e537cb1e20f908bac9c74f3d5b85e2e8e7ed34191c16eb45e1bbe7fb98
za0ee50052b77c884662353b245390b015fa7de432c5c528966127330e741382d2f10dad76a5665
za20e18f110632f2b22881c903c671a26a422f27e890e646a308a063da66ea434f62147b2795a96
z662f10becb26646768c96e05beaf2e12b0383aa74434d6b8ef33aa14ce82752abb8211d0b9fd54
z7b75ce4591784ac65a779443f05f04a0b21b80fd85d7b08fbd649bcf3c4c5048f3c414b2005d79
zcd112f1e081a9089dbcede44f5ec3f1863d8a89b3718eaea672e903a5445979d684f2ffa165b14
z9fca0f94e4cb774d3cc660529f0b280af2269f168588fb6ae50b3176fbe015760eeabbed461ec7
zca0c3b13ba03abd5661ade5f79b5c425febf8c1662cc5a8e2bbf289776efece23822cb40a78165
z3acba7f2dcb849d7b600cae6b1b412cfef915b196a672c694cf528d0e8234a7a984236eb04d314
zac8efb7ab2c9f354a0b2f752c6035c02e4c93f73fdb6d374397c50070a6a596f7306fdb7cbd5e4
zc28f32a2ae85f5f923f260ded24aba0858a016294252d665394f5c17712b4ca5a4c3486ac9cb5f
z26dfbbd1c0f191dffc9e2dc89c7d2691b28f8ea169277275b0f3e8efa1703291c496b878d5412d
z7277bf2aaa343d1b781020904897c754f8601e14c29258d4ea0ff34b7c4fa9795fdb1872fd03d1
z1e6ab5cf7cbb1cfc5b67c559d17f0dcb4c6113b4f243948ec9f9cb7ebdbc5535ab48bb4df84ee0
z27248e308b92f9607f550f10d59fad2cd0c5b3413a99019d04755bda9dc11137b7a6fa8c335510
z0f3dfc41d13e66c5b93d2490ba0bb337c3b72624a517022777e1f3273941b074fbb92b93276187
z1404445baa4bd9ff1bc9b19c55e85028f6ea49725c1950d6fce993c1e458d2131b050adfa16421
z7648af8b29387c6481f1078dc779d0d7f1cb65b0605e14e9bcfef9cf4575d7eadc73cc12058000
zdaa9153c5751025fad3fcff654af7dd1d11c30930e4c3789a4104f3144fdc66802d8617d5b1a03
z4659dcca60e79d97b3a87c53df8a6268c1231aa3f47f31b904ffa7f7552351b0901eaa0d651cce
z4c6625859aa3d4d2405bc33086df2b96b49271e18e7be380c818bc5319ab4e44bc257b1cb8b398
z5234d32b5aa48c40aabb6bc7a5c174d8ea0d5206fd58064e9bc7eb0d9cc3796c85afa2c3e08eed
z319a10068a60c584042988973c38d54d646a82e8e6dd4fd6d818816c867474f0d5bf26522cc37f
zddaea23cba65e7a19ce8afc228410d2f0a16420f0a91aa14267fb44c2d7a4cdc07bebd831cea2a
z4bdf5a394c78ae2250f7c186e1b2a8b6a669c9de8a3cab8d5646e793c4a28ac55592e7efcce214
z1d709ceecd80252e42ab940b77ebe002bb0b8c4ae471657e6da34b05de5237e0d01931283ed073
ze0581ec03a0c73cc7e29b91fcbf8fb9ac1720b66b99b799458d55a93a61af8bbdb59db75722ec5
z0e4f4fe4da9ef067b51d6ecbe36cce5bdcb0375ba2ec774f9a45806923056b1f6d70f5551129ae
za570f9db35363264a93d70e9a6f17fab5e0e7a1fd3362d3a8577ed699046702efb343122c8faaf
zf7874b4b75780113a16f6aa13096b5d55fcccafd4f2cfb887369ce0ad97e859bd1ceab5b4e38cd
zc0c09f7786abd21f5272cfbbcb1c832836526ed546ec0a31ef41516f4df62780fff3556bdcf1cc
z57616fe1e00014936ced2ac2a9e90964946819c0a4c2e93f05787ba802ef76595271916c840719
z04e9233095a8ef5fb5c59a7febb2c453bdbe12e4da2e7f16e369c3b5ddf4bdb8ef0951cda1ea19
za8954f2ad855b3ed771f4b9eb8d48f450c086a6c44b0dedd87acf01879ba95c1bbcb5c8c12f3b5
z89478a27367dfd448893452bcb69aa9606599518321b68f81ecf3946c6b18f08d5d10b9e6a6a07
zeae3294a86db1d845c1f6e31b366886d35afa655c81c63172d30f0ddaf762d6472e69348a21e3e
zdbd0c32f4bdcd2de468574c7dd335a89df7e9727e20b1cecc9eff309f65459eea566da12582219
zc45a175427f56a23ad347282b499672404bb52d7755722241763ebf9bbdb1e9c8b84687121b559
z3857953c09b27f7f4a53c5627e868800cebb9007e5f37aaa233eb8026cf0c41105dd7c952587bc
zf655ffd1cdc2921af7661a9556c4e74ed1f6306d6c971ff8db319a63ec18a3cb032802df00f005
zca2b2c571333877f267df8590bdc533fca6b6d16ce0d8b8453034a887947b3e6eeefe870936bf8
z1c0583d3e2e7c8122d3c6c860a2c3c38f24b43991c8951ebf933b800b6fab9a270d48abafe98da
z65c3f25c2be3741ab5ba7bf1285ff20f3e5b06698fda821a60da9fe40e43146492bf0e7de1c51c
zf27fba4894066ad5ae7c30f5c2c5fb947705609c2a8ea2ca8662f4c5484263ef7cda7ccc6ee8f2
z9fac872291f784c70595165c6378458a94ad47b9cace0070bd99287ebc149f0cc303d4529eda55
za58a8ddb389b20399a64cade97b552c8a791081683b2be7fdb81ef7d5b09a0d21603dcb1051e07
zd2bf53ac36acba0864dbaddd358c76309e9323c83c525836777cd1b638f874107c33add4781eca
zf220314a06410b6794caf08006485e3c718c227da8799957aaaa658e936c9d35431f831eac3d7f
z1b701ec7121954395d7c98ab2428f5342287dc57a2426019ce52645d098c92ac05805a3ffe0384
zb9c577f76c68ae34d8af66480317eb33d4660aec9738b3e03df1202356a3562157ce70a8c595df
z896e27643276e46c2d37f0b6141010f80e8559ba0d82b4dce3977dbd6e62db13e8b28913335c2f
zc84c0acb2b3b1acfa43c29da1d6b766c952bae4a66268eb5e5c3867a745a56acda933ac963bd2e
z4e99fd72630e647159d731ee819f5937ef5ed08b40cd0e35b839fc8b1bd7e71f4ed77470c1c6a9
z7a7051d128e0595ad51caa285b0d9ec9b0b2eda6a8fdaed6756ca6d53b124d90f9ef27e8c226cd
z412ba5c9240757eec0a5e94aad1c6061b3ca1eebee8b948c7d3ccea3256c5c86badad31a5a36dc
zd047965236ae3095e4916624ce381fd26e501562c79867dc25ed773e8c5f6eb73bb6a8ffdfad6d
zb559b63764504524b2f3c5d0a9265201dd74c316b18bea54e59a5fd8e9c30f3f043a9fcc245e64
z5b5d3262a490f17f5d252308696083143c7d7b0cb182bfcac7709230525c02875ca9fcbf7d5ce1
z8b7b41cb466fe52f0047dc601bb4479c9ff707198c9ee8a5942b7041ef1e8cc6a8ffe542532425
z6b27c7d0a8fcca0d00aea367460681751d9bc56fc8c3b98070f07cc646c2699033598664e35718
z79c023231ec21f775280bda2092645a7d6e616103347c677d7d99693dae61f61a6ebcfdd7be435
z8e847c82afe859f3edd6e7370d25190e4def2f61ab28c8713c858929974578d8bd38788600c190
z7a58aee7dd2eda6b9921f35a45fede27b7452c8b0d1c823c3d553ef7889a85f0c19f79a335cc0c
z9434139fb6c1586f3979dc80b329fecc873b50661eed7d238f1b3cfd32f71a6c6ae11dfdfbe992
z3579e06ee9fa983f90c09f349bf74351c88db169e9adbe467743673feb9039ed91e1a044d9c706
z60ff1b5f6005ff1f47abcf24eebea3ddd3a597868aa2dd9b77f5a819edb6c12854117581f2fc5c
zd79e949100c3f244b89a18692083640231effd1dfcd559800756b71e5d2b3999ac81ef620d7cce
z74bafc1a302de25779fb871785d62e7f45fd4c4ce82c72b19e0e6627d5070b37a93c0c01333d47
zd71dd39a3214736975fb8596287d3eb700bd1923059cd9b18d2e008a1eb36bea4a42fc2df32191
zc1cabe593b7d9bebe44006399ea55d1ead841ddd626895f7786d75a8c0183a53849e73f9b3c927
z3adc7024e8fb43923cf2cb5e4ee6cf56bb3ca4e3ebeb4469be917b9dd918b4ef2018f7dbdb8dcc
z68370ce7b0df1bac8fdbb145e47161dbd76961fb25c5de9773470f74fb4f3c89272991d2fcbec6
z829f10e2d66474da2d056ccc52f5b0fc54dfe876d68c27e3252e40ce6169d586e6ae730421827b
z2881a88b0ecf3219f1e990289131e2f6a89e492623d4dbd801627c68ac4745caa4e326c0093585
zca155357658c2854622f22e2266aeee10d5ec53f066154c1aa1fb24869495219c852409d69cf0a
z16874e2683adc1925aee10fbcd5b1aa96d3c43e1afe0f47afd96ba1ef246ac324b6d39c6b94324
ze05bf2eb87a567448aa861c522434c5f959ea6dce7b60b6e05ea9ade425ae1418eb8eeaff4b3a6
zaa3d352305dae86b02dd17628b888705951c931e2ac0ee6705ad571682a05ac217dbaed5e080fd
zc82a4a5c4fc451a4f3a7b201c0ce68e38633a9b678e35975c7cbd82c15d1faceca1c3ecd816363
z96739a4708ec5cade61de7d28202cf5c14a56c9615b035a5bbffb028ee9330ff2537d91ca2d315
z1c48a0a56c8e39101ce440364c8d5e12f9715bc3cfa9673fbacd54f3fb031983a49b1f107035c0
zad3fa2d3aead1fd85086d34bee95531c44d468eac296ce386221343dd516c5f58674598fc8164a
zd7ddc7a8e6aaccf91eeaf1cfab3c8cc46a43a03cd1e37efe6b3e42c1919c7d2126e00191cf34c7
z8b661388f5425f573612f8ee50d0b3a253fe14bd5d1dcff42af8858d4d661acdcbd7c4e46da3ca
zdc5f50921c19aefc67cd6d2c5a1d40107cd62cb34985f4b58df2f03ba85b491623b399f97c82ae
z9f6bfdde6b7a8bc8a3b821e7e8a2cf3cbc8caf6138882f3fe8db400522c14d72956ac81faa8b56
z71d79ccc34014c109b839a4579a7bb12ebfdd4e5b956492529b2a38bfdffc01de8c94424adc31d
z85a537cd881fc25e5a25ed40a3413d24b52592c9cc5d62960ba3d2b0f5a66e5aff03ec58c30ea1
zbe1074df36838f63e53ee641f8e2bc1031992dab3e1665bf1e8ba8aa66394a5c463bdeb8ff6549
z28b1ec7587446285bc42df51273f87dd4361779437b8b7d4d813f4e3abfe71bdbfebc9d430763e
zdef334106f6e7549f8f27c208516502c19dae45d63e72425ea15210584759e7c694152a5275caa
ze2f464f913582a8f43827bb77cbdc22bde938c45d037d06ff18b980134f4878690cd41d3227cf1
za78942ab08c700085afb0b020f49ca7c388e3bdf46301e998463fd6979bddf0f2d262f29179989
z1e0ddf64b00b70f57596909a617239185373cb1530be597bd7ea41c622658e0c3952baa248b7bc
zfb92e1a0ba51b4e3de29596c204a26f5f6aa5089606be706c9e664f247e05afb26fa4138589dc6
z0b15e8cf4bb375e27d56cc7be5b2e9cd7ebf3f5394218d3b58cefc9cbfc469b6e58fae68862ecb
z9041e19d70894a36b0604ba00ab33ac0d50385104ddbcefd083707f62ca4bfdbc3559d5096724d
z49dd539ba45fbcdf978df946b31bf19b652fb3e71109b0c42b0b2b0c6df56c5c3133f7729f55e7
z660b9f3f25d5becdfe91cf85304d96fd3d41387f9ce1deefd09632d379f8c58f2913fc432985c9
z360d8ffd8a357a45505da01ab146b6e0d5937cfcb658915ab6b0878dda22dcd050bf1ab7b994ba
z077235c329b9c12162b5c4fdd6e3046884daf9a95d43e7148db62db20cc237d38239ad704b8de8
zdd323e27093a8d744e3b1acaa59e62354117f8d0c1b3178ed162a059c94a5aaf1e38d300305db1
zf6b6940fc03006363edeec07b2610412b602016ab8eaa3a14ee7e758b798496cd114635b857c93
z2e6c0d3e59840ced7ca545fd90ad392c8e0506fb22a9fce599def92bc954e3ee1a81865bcc7afd
z82754ddaf2b279a85183bb2af33364fccefd9e0f7d6f789f136559995f83090acbe504b8e02875
z49eef3478d2d932694de366f0ad2f8961e48796ac31a40b68ab494735d75106054b1b24bbc7b0a
z12265c9702f22c9bb8e1ecdc62ea4c592e9967470489500b9649ba1a38964838beb1a6b89ef723
zba6b34b7ebc795c852f70b5317319725bc2c9dfc20797faa944a20bd5e9ccae344ee2fe772d474
z0e5aeb9c5cc5792ac4c748e446f6fc42e722863433ba71110fb51ed59a5095278da1f1a8f60454
zc550a4e9753dc10542adedd7090d26f73abb706e1bcd97b64c62c39a9c966b06d75de50c29f903
za1ae74087f57ba4fa836e02cca19737a070bae74e485a782d6056909150e55394e24cb786a734f
z39c7fff2339020d27ddfd2b996b040ecceb6180d6e39902964be50fa82bca1f4369f334a3ec9e9
z13e73a5458598a3ee7c111bb3fc15224900c8fd932fc8aa9a373f12cab6345a90521a363aa32cd
z55ff6bea5f1c8906c921abec91e04bea74b64fd5b499cdb517125d38be9d3d14af59923d1b559a
z35e3e6be3220f47dd7a2d76ad63b8aa697f58866734279f098113f2370b11eff8cbe5710b0a003
z5602991d04dd757fbb0887fa3e53c763f1c69ee156c6af14cf5120201018d30791a034015edac5
z7dfc3d9d0ec92b7d9b381829e5cee5df20169c00ee1f27ba263b1d2ce251dd052eb7ba9ba30f23
z98dfb32d91d8031793b1f4cb3792c17f7a363b2303e443850ff1333f9a92a7c55f31055083cc3c
z233a4a5382df84b07c0c2a9bbf2ae148b86ffd461633817df69f1888ce968f922600bec12bc050
z3b52e6530531e76b73c28cf1c1218cc681d6bc182c166b06a01d7fd69859ee5b91f4973814e2d6
z7d0d2067b408f9b991d41a99217dce5d825817b7fe17f48f1e719c4dd35759fc03e5ab07413af4
z0f88aedf742583d144f1b2fb32ea76ec9c33a308094cf8b5ebbfd1a5debb7a63d6e3f89beb2e94
z12f85f5e2c9c0d93a92d889d88f4d15d542cad83f66f606d834f5584270f01144591058e43b440
z4f87e9addcd7df692bd7f923dfbbc706627dd7c918e9c677116ea1322ba255175c6c2680d4d540
zf85eb819fcc2539459c36b68877d4e8edf64c886a7817129c3826414da97eb22f8ef8273f569d6
z406becdc5aceb434200897fe3016b91726e310ce739ca802eadd1603c89c029e1e1358459e2071
z08d9bfd0f86ace4e81237f6d3f64050bdff7af4b09c4940f94cae1c16a5c6f07115e95d482fb00
z367fe5a099e6473df476d9bda07e96189b8d60e6876018e2828e09fc7350547abb845b62a14844
zec82948794061e45528343fabbbfe38113d12123fac970a347a2fa397e62d034a5aea1f2d1270b
z16fa71a7529be2d068ec636f0553f23bdbb6dd9a15ff2f0bcfc7e22b6b753b0989c78038532907
z49bbbaaf3613c7af2e57dda6cb53a681b6eba610d9dc849da4b2bf25dfb50e7e13cb9e92c67bbf
zab7271f7482c4cbc513d39fe739fabdf82f9a86b367ea6cc99d7b54ed1d7fad158d68ddf04a23c
zaf7bac4ce03e723d5ddab11cf513eab0aae2e979f587252a89c3402238514869ae052ef0692ef9
z04fda6ae603c129b8447fb5f20558909c4ba90d97d179ebfdfff8fe7aa5ac3bb159c6735725f46
za094fd97b0beb6ec246028554cc1668cec6459cd57a0372a276d505d11b9b1f67bdc2eb1bf0062
z668a02bcd1ac6eeb103356c9abd48a8998fa4d48dd48a0d3009c15fb9599d13a0d78db8a75600e
z2c8d009ce9ebffebd7f83ec63bf83b9b652a4be44496418aeebcfecb8e88e61c81dcb9cc1dbfea
zea020cad18268e6850f17567db6ccf7deac9b3ad8eda9dc7fd74f9ee35667107f9015ae5043c93
z32d7ee8e58d408bbb8696ee75d4ff022c0109f8c3af45f77cd159cf3d3cb3955cf41d6cae7253f
z5e4d635ff04bb5752799fcc5a72cf9eaef9b61ade40ff7dc05ef5f3f2ad3f025281a2607eb418b
zb0069867c6585c434c77ec69e9d07e9fc57565702d6261b5501425db8cf06ddc37ffbcad643336
z8a22267d8abf94306c4ab96f1a1aa77ec8b1f48a993652221b365c87fb72e862ba86804ad9cf25
z097b32045bf83a956c257eb3fc30c4c67c48d9e7ab5b6d1a7ff3eced3a5bc0efc5356006c804ab
zb98f7531abe1700a873a7deee7c70d6bb43904ed8615bdd9c599a86afe36a9c7a2a0a3ace4a1eb
ze7e65b79f16273fdf55eb05841086b31da2c6e37ab4f6ce537771e6daf3d0a2fafabd914a5259a
z76d6410d81c786a427561cfbcdca513e513d89d890053da551ba296309197f573ddb9ffb78c26d
z901a736840ae057fd52cf52fc4eed9329e7d0110f536689f725a0b25546a079ce60c5ebd554841
ze3ae6ef68769c5dbac201a7d0767f6e374dc2e5e139890648f1a47f8920c5b1250fd9f5ae2d24e
zbef1e0f9dc30ccd371a40c4619f735ae0ac9603320a12a511ffbe14404ef9b00bd6ac877850fe5
za2c60c93c40f49e8a50bbeb25c44c27d68cbbed1ea2faedc7f038659d5d5ca71d2d15bb4b10497
z496770a8e5ffc9c45f6f8c794cbe3421e96253c2936ef84e73c31b90c381e8d4cdf1acb07960c8
z1a34a0f196f505e937226eebb3fbf287a0155ddee7f5e2a5b5a07d9a41d51dfbfd32f362a5784d
zbbafc5690667bb66ca9f56c6536078906cf351d0891c8d4b39afc2d0e01dca790599550dab0050
zab188c08eebcd06923f33d39db6f02b7372b78fa4d2f2a495cdc1321ac6239504d8f2aac417462
z7b3521befd6111c18f905c6d1d0bfb8ceaf4a872b5e82a01d0b345b5cd01d008d191e509befe73
zd425854aa30c63a5a691d61e4388ab1db6ac970f46d51358f84476c9a173e3c852115ff1a26340
z68d643b389bc995e05d8eed4abc15e6b66b86c25d11620ef503f350dd37da1e287a5047fcc7331
z9165360da756d2fc6eadd2111f20a9dabb967b143e65aed262db8d4db83fbe57afa2f5ac302fee
zc3be6a08bd8042e2a83d786d5e7a24f67f4a30ed26b78aeab6ed161cc570652707b8f3213b16ba
z9957e8e936c016adff6f04b0e667e940f95db6199204749bc742d0bc12f2a25f95119a74236ffe
z270d84f4ff559d6b0140939de8327b016c79483774c4aa410973a9366f735133cf4eea25407c8e
z4835d7d7b9f2b33eda9bbc54d947b8d5415d38605792354fd91ee1e7094a0390cf3d680579f41c
z6e05da547a4ef1e03136e1dc3f5dd037a0883888089b436e95b031795aadc50382b1f2ade92191
zef762dd247a41eb46b2f48ddee8c8f8f49ba0950df50165415566981b1b59d9269aa49a5a7ef57
z9829f97fe0f608b8ec4cce39b91649783faecd068e94694e3e57d9dbf418f638b74975d8ee4672
z8ab38cbb412f680b1956854db4371f9754c38d6ddc50570088f0d9ea95c515886fe65e01a4e12d
zdaca88992059f8d498d6dc26d9cd0a0cb8137206b3bd472870fa5c485305a2a01f3078bec5771d
z8dd14d9b1dfdcb11ec491b40ea169909ca8d340013421fcc7f2856d04e8969810b4a46426fa912
za0de751784e41fe6d66c3e001048ef8b018e9c5b2d92abf6db025908e23126dd4bcee01b7bc3d1
z4feddf3d3b8b8cb71ee09c8aec00488b39697f85ddeb5190cea9233f5fc6507497a2ab2db559ea
z6422dcdc4576dfd5d4b5519589afdc7aef1c5e265541c66d775c3be72221f67a7d8b16daf891cf
z32eb893c68b34b3d1640119ad701ef1049776fc887aa29b20bb4f25ba2f79c931bd290b2158153
zf933b67318b7296bb7fa7d02aa2581c1b54a102a9d352723b1a9dab20e339111da5d24aabf7fec
z34faa10a3e00efd98dca3f787badd331635289c1105bce17cc0b9e968abc8ede108044c168295a
z48108841a6fc2a817174f996b90d763fa24ae13fc7f8c3dcf59b0b0734622d1d96a2c5e5e7c82e
zacd86772c9bb6260a29c9428ce0453a57778d1fe427ccf6ee5af3dc59ae9d7a287d296f4160c8a
z728a8ba8e71b4df8a3138985455b654e337a2345f5bfe9bfa55a40279ebcadf362744dc65cfa62
zf74fbf96bf3595394316cd78c2e3610a3e90f899352135382d6f652799db5a2290ecdc7490c466
zdea2057225c2c023c044f8bd5f7b971028a48548c08dcc6ab726524e2321c58d7f725a2c711162
zcb5e9c2e911dc4d0ac5a2b19a28bf3319fc8a02505eb4e007323c8c7f88d4ee82b8c3a77b42ab9
zf4643d83efc6a97f84aa4430deb20ceef2c128a0a7246bcf373f9fba76113e1703efca7e2b08a2
z4bd8d80cfd106514cbdbce00d406feaa6bee4be44addbd6b03c9f9baa6d8257ce3b72e1662cddf
z19b650efae7268bc9b4392a2a1b321fa7dd88d2303e2aa27f314b09e3ad5fdbe3da735a3128dc0
z61c810f3897d2ccb34db6c87cd117003c84a50b1c1fe37ae29f4cf0f101def43a3d2bf8e3e9ead
z088c5d7124a8194dcc535199eb29f186cf7761689b75f23e00dae93f6f3d89132ae4af60fdad1c
ze41bbd08c0c852a927b63244b1d8c92757a55c0c3f07a1be3068d4c9e8245b52c52952db608855
z38a4824bf783a8277d278e212e1de44a248bc719818a05549c7d3467fa5c84c09b279fc63a548e
z1d4e085710557aa74e495e45b288e6f3a2b31afd233ce44a71c23982763a5a74fd23f8284ac4f4
zd0ebd4aa4836e2d85bd245901c057dc040a2653a406729ae0578387480ea060c220813951bf14a
z56326d6cb2f82e27d46b21474d64011e89a755813c93cc293de54b0a0b9aea06642f15796cad73
zdf727c875e4c8f06c45023dba7a7df7aa3b652a6b8654998f4744ab8586799c5dfc23f8851288e
z0e18bfc0df020b5bbb10b4f7e6bed3535a1738c72f1c4e60a246a643fa0140a928e930a88fdd67
z308c000ddab04b4caea8c4f69039b772a77522b1754a7d8dd2f85f6ef0188adb5463cab02a62a7
z0f494c0c9883412ff569412d4550f0ce7d90994094ad47925e2ba4aef8fb115992a783d086daec
z7b088c55d14ef49c65a77f2d0e677d2e159c1869037ec82c51ebc1a3a52cc2ad9320c1a865d7f8
zc2b1db59de66e62ce19c91f98d580fdd93ba19840d775ee5894be9cc7c754da199c076964c409c
zeebf4ca6b19e2ca5e21ea5b524847215410ed0106f59e9a87dbc3ab925a2236c3b6b563e5c58d4
z41a6dfad91d11fa1d0ce4851ac47627a8a8bee2510e072a83e54d3cf6f9f25b9dc31e812b5912a
zb13f76f1e76586ff22770487d8a4bf109c739a99b655eadce2461abd5b319f6a9abd2a2c6775e8
z7cc786629fe024b464f98a6f8860ceca6e7d16593515f295b9c03e615102a14a71e65e88ec8907
z853966f1ed744beab521121caabc0c7918f29f8c5fc7cd9c6492eb0404a8808ceccac55e50cbe1
z89debd1007837e39a7ab85771b2ffdbafad135776a166e762f73092f80e5fc0b1b1ccc46499723
z84f6b3d920e4c81da0a60969f6cd2e909865ae7d9e53a8f53544bda605d37730d8ed11a98a4ff9
z792949e93e36797f2ce0726e6ba1b445b1f689a5294c7603f1a891614b405155403a61316cce82
z641428d9a593313f1f83d7a2f27abc9a7c0b53305fa302a732d48956d60feb7ced2f19acd8084c
z4b10c76148d290c6fd57babff01eb964376d8196af81032652089d0f4f8e7b110e0f0b5c849ba6
z2311dd9358d07833f274c11d1b1aa5b9a98a2bf1484108bd7b43758e41a63ff592bf503a818b40
z5b824cef603724aec284f4ce3ad19af5b7c4da58fac005bbf8a4ac93a98406eed2255f5045bc91
ze0eec2a9dfeb05ada36a74db3987ba8eb509e30ecb039ae8dd6e8c05c8207693ac818f24ed1f6d
z8c4ec1cf9efa1281734f6cab5c9e1ebf1edf3b5d9686e43adce99aeb7d845ea526dd4fd85118ae
z1f9b460d5b4afa2f6bfab9bd9bee269a8d1cbced9c257f0a7d04fa7cc730b17962f29e59f61125
zd0b0b536957dbad4cacb08cb5826ed79ff1b5f7d75f4313b8f1bd96adabccca29da34bc726b300
za9fc8bc11e29d8187d1ca5c5fd5e207cae1da6377d173d074ae88645d977c4528f624b1fd3d5c4
z8227146f0dfa53217689b759205c3d81aa537873fd75f41cd53acd3f1d1f09d9657f4cbdd35140
z73ba757db3dfd5673272490e5c999bccbe3705781ba5a397ac7714409e91b35c91ed6f72a70f03
z95157e70e15f7c93b867c772ebd625ff6ca0cea86d7cbd12759ca9ffbed1e2284ac9137dbaea49
z5dec62c221f3220ee4d77f0dee97d869b2991ed4e7319cf71184fedde018bec16b1b25067fabd9
z6f2ac15be02be89cc366fe97455ac159d1f2834c092d8ef93073e0632a42e13971699493b97b39
z0be4faa04a3c0f5c03c8be45de6b3bce0aa0d0ac06d327ffa34bea6b91331b55c09ce01a7a7644
zbec333f041025802ea0fc087e8e120a8c3769b49bb7ee784372737018fdeec6436fb9379d6f7bf
z0b4b7a91af0b05cd24f3f23999388247b86a3d91908399ea0b88b0876b0a16e36da5543d6dde57
z94c4c7a033265ea761c8bac498171d5a7fcf7c72deaa9719a937e93d561c31d4a5b4e0cbe492f7
z8ca84e028d66554be6d613f037b82e40cae60f632c3b7b8c630f7b9f9bbcb91ae41c80bc767b9d
zaaa45b8af7bbab71b79e8c87aebdd9811887c69eccf5fe07a9a205e7d7bfd250f5c059c2dad0d0
zfdf9f21f8de9e0482448e27b6d9f649aee91a6c28ef7079df2f23b88361bdcb370e43cfebd8766
zcebdda61aa20cfc9682bfd21c0d8bacb6c69fd3b79c7fc6201cbc797515d9c1afeee88e5a592c1
z5e5c9024bb3764e8435e2ec6e608aed7aa14bdd832e5931e129e25d0f85a802825256ebd3badd4
z0f5d5fa2a79b4e29145767385d93120ad674c43c7455a93d8426ab0ce2bdf29380c2c3ca7fe1f0
z47492033c83b1fa0fc86cfb1e38dfd4b762afdd9079c2061cea33a0adf492cdfd1e67c04acca21
z7eb79941220c63d742bca28d3a3b3e99d659275389b530b7b8e413372521ca64daa595fb9494a3
z2f86afa1bd86810d5a7f89b2977b5c49eede91c9fab6587f48c88804a395e4cb5a0336938899f9
zde012b0a7f74b31c5396662c2e420afba3b33ea125235573a7c4616a5a137115f111327bca31ee
z4163bdd66be3f9b5c95f9be8fe1c03ea2bdee0e41e8985ab6eb02996c40e92444de9e34593607c
z877af01edc14ca39b51564fdbe5e00669a40c60158814b504b1a030bdee9ac43f5179f090ec641
zb09869115910dfe5169198b075487fa0920605e17f7bd0c7e7e8b90feac53a98f0fd05c376d897
zdd3146b99c1fab982f28d5a5678860a98a4ee89231b73c51cf6befa160e4656944142ff62dadcd
zd6075d321538cca53f7463fe42d6a139bfa412c2157c7ee19ae60b90c272d1f5e6dbc143d120f3
z9ca8a26fb99b6e3d5eca01842f2e8c61ee8ccdc9ee2900291520d22074c546cadb1b991527bb3f
z3f0f4182b87bb2d341d7d42fdb4adaed88b51be834a4159bf22d3fab58e55af106f4d23d4567ca
zdfceef2f4c733901c9d380075a0b5aefee7ec5bd109d39998c213678e85282da8cd5bdcf304601
z80e1a473e81dc96014fc0a6510c9e325b7f56b869e1a0fc01a9150d553ec0158b1055304fdae00
z15c814bb74a492d036d2bf9606a4901d5c8514d407011be041957f81b31d3b73e030e2c401f6c8
z727f3b2aa71cbeb1fea55e3e2a71c1fc615d0a83b76cc6845bb3e453ce948af41db8b93e7f45df
z047115274d44921033666c3e0d24be9979044eaa0bd401f863456603ab49c2b1ec5ef37211a65f
zfc2c1f5b26c62b794bd8e601f224982171efcbac05c59c3dff28b7317028f64d6a4e1c00686e15
z9e9389dc5e3c2d13b6e4d82915fd2096a46101d9ddfa0d24640947ca7e9df00d142846895cf159
z5bf53ea72aa1e1a1a8e8940ef7a9f1b509be5f34aeba9ffd25a6ea13390e0c4a709b4317476022
z83f6943165db9a034a5149214d6d13321a568f6253879955e54d029980c690dad68b1021050ed8
z0c7cb7d9d8dbcd27545abd8d4cb4c98de52ead6192bce079c003db6e2f664aaf7f5862e28d18ae
z0f63af0e6dc656e75d98b5cff323ca3ad7e98ae18590e261edcb44c3a4c2f816b06dae9562bba5
z712244626ceaf6acaed6fa94d230075c38e04dc6caa98558de7c97ec443f08fbf74aa02fc4aab3
zd6320f4cec4492d4e46d87691f80653bc0f1e2a993fc060cb9811e37a78ed50fbd2eb988fd7fe3
zf1efc0184e7309a2375e7a06e38a52a4aaa75a5a8db81be933082a00d0ef3081d513732e2e7691
z19d059042195bd38a24d08aa6cd2c3afbf6481b989cd8f9a57161c04be85346291dd13b3b2c9b8
z5eb08c2b0e7d22b90ed2246c7c928b3c20004b8eeabbe21c325436ff4ed6f88a886f6e2b4b6eca
zea7cba26ebff652f9df770f01bae925730791c23995e5503fc830ae813f66a5e768e7973ef0d13
z909de8f6508b20d92656dcf775b4179063d4cbcedf17d1f11fc2e840c62d8d9471d94604abe36b
zbb43191530168555b1968cc4010f46b67ee37e5e3254fc3e61f8965046caf45f4d996c0d556fcc
z83a24d6839a8262f4ec8f0e38ba250b09565b28c1a4e2ec25cf21043d3fa0b998669fe8d19333a
z4ef1f515eb59925cd858a5f9630f1d3d1fe822b07e04177c328c86a9dd4de54298a4028701cd4d
z9098d4abeac1fe4e53db8e4df1f4cd03ce17ce09be7c8139b451fc1e813fd56c5d27237cdc21b5
z2bf323b2590223ceea4243ab4f9c7357456578c1e20de64d78c84fcc279c26ef7a38824a1f82dc
z1a30e9ed7616195ccb9eed8ee1ad3098275d7b0bc2e7a2b50c67d97d6eab400084543f6b4df2d6
z94f2ce9f5e5642cb6a3093a4c2d21fb2f1c34f0ff6eeeb2f74f7e1d5cd42b9a7b248a826c2eaea
zacf8fecffe878b56936ef03980b57f2186a59fc893998f9fe1e3a05831159f60bcd50568cbb346
zd6692bbf5322e28007b773bb071c4df47556cd0412b9d85b62c7dea726967a1b86f583784be1fa
z8256e6b73bce691cbf112f2e3777c38a98ad74ba723f478ca56c6b3f1fb004ebd71fb02e8d23d3
zb842fcfed2845abac8c5c6c881a276b59aacea421648921b64a6cb680ee91e2230bff69f2530a0
ze81d92cc81bc2131a8abe22583b18d24fe268aa6b3ce510ba86de71c51012c0aea0ded5e819675
z2b14cfec8d7eee08a94beda94a3d88109bea954a52e7bf19722ed2d80c246cdffdc8c084451202
z36190dab1243cb3ce06a393e8685cb6479c1d0ab9a8388edb4a2257b8765d7ba32572447f42ef8
zd956ef80b60db4dc03aee607afc7b587a533dfad69a02c845e777ce678f34783a7877fc1c06cfd
z8391185e1afa26ac499dd1803a90919a05a429372c99ad54d87cfa5c373adb3dfc5afc0701cdca
z54a93b133442022028c12ef0cd11104bcae39539c6bb23c5cbac1888157055c7cb88aa855ce713
z4029b9eeeeba0fb9314792488d1a7e298521c3e235216ad3a7c96fea276becf1109463ea82c353
z0708c893f8958f31e92cdbeb738a43f6b17a6c46b9a8446bf92afb86a26c9f3ee78fa10b0d329d
z57804999c035b2289e76c31d7c7b9e489ff0c87aafd8e79ea6fc7e3628bc60a4fde79f5ccc4353
z962284464ec5f084443d8f67d9e673c5598e6f222e9c0113016cfdf9fceaa988dd576e4a3d479c
z6e53b5d7505e9a2b4614dca4f0a13603c991b0c2c745d5d35ff20cf3b9ba868eb3622195e3c2b8
z8097616ec5deda9b235a2b632b6a2c5ada75113b9a15fd07557269b1679aee31c9ce1ddedbbe80
zea779c62f0b7fd28f073bb8b1a3bd7b1323be2b9b5c7d1d16b85a49d99b62e1e6648045e0193e5
zbe88c5152bb99eae4721a9a5a1858db914d26addbaab57455f9e62c04312b9db50c551a23ab9da
z177cfb6ee8694203d4d82be98139bb49722296c65f9d1dc529809a6b15b740dffa7d0ea8512303
zd059be1e870bb8cf7ef89d728133215fd180ce1ec173077594e203a79dbf5cb809abca1efe07d4
zb502c7ec7c0a0203c237cc0a5bea0dac6e624fc4c68730b6142f71e327c2b4edde9ee08c25d51a
zf189db44b03fb0dde0d052c9525a66e18315e12747c0557f90bc61f0338cfeb0dca052cdd52eac
z1a31e6ce46d3b805d08318d46ed8834dc68508def71c264e71f61e41c459ad56e14b075272809f
z36821c6dc4b8f984ab69e76b90c1e79758c8b7220cf7242204db5ef27e2d8919a7e60abaaf4b87
z88cc5bdb66b2b7829d8a8421ee58a67be044fabcc6c66c44a31f7430bd39dbd29e42ff7effe0f4
z383bd9659fe1fc3be6a7fea9572f052c67392c9260074db293ad07a44f32d0dacbc85b263dfcc0
ze454addfcbab48d044f851bbfcf15c606df06989e73b3169304b1431767b3ba30a0a032bf00644
z5bf6276e6f004e222277eb7d7d069493f6494978aa5383b9e3bd3d1f9ef4a43226ba4857f1975c
zebcc91b9a0c33ea7c02c03d90c5ee5f1d1d2156f5f5991903a83f653092557bb6fad17bef960eb
zf099f30cf3e65549b1ee0c9f1ac09b2c1fbe38a577501e5b37bec8672ae8f5d4306ace610893ba
z45ab3f790990765ef5ca9d0cb29a562240cb862cbd3cb6fa287ddf1bb3db20e8d8a262aba22bbf
z91dd58f9e2176f0f66101bc2eeb68361939ece3dd578707d315d277d94b4970147fe6c2a7b733d
z9e66436459cd2a3f29cbdfc366b52470432e6867d64836c1865979d0f54cbf186860bd02dd21d5
z32d9b0e851bdfeeb844774a26df757d4846d0c05a45c55b10536596c630ddba0817af31ed9ca6b
z7eb1beecbe15a25898f1b2af857c6dae8a4fe4e029d2dde5ede895c707686c7b14946ddf0454bd
z06bde760aa0714b3480066431c97642a2bafe662c5f20254622310a7acd413b8119a72eb8a6d60
zf627cc15560436068466c4958544167c56b6ad498da3b87d3beba920b087abbf3b08f6c8e92e6e
z6c5aa39ee14c5550572c5f8f7f4088c1a629ac75710f9041d41f6d2452cbeba4a2f5b130a0b139
zbb8583c9f3a713dd78baea673d280fa34dcc2b56f68d46a073d8c0033743ee2c2079d413c5a746
z719005922815f3752997f0cb243517aa142b210042abf6d321e7c3795b2da7cb1037be502bcba9
z85da5d5551cb3fa3d06ca2ceffd4c23ac4426cab9f28e71e4ce8e4d53331ac167d9934560cee25
zc2b55e5d19cf1a3882a4b5ae75be8af472c27c642ffa33bbb076e50ba66212a29fcd3899ebe945
zfdb3dbf5afcd438b09bd5c6a9b07d7a82999553df7074e0fad00eebdcd03a469b28871300bc3ac
ze5cf14fde26ae5d7cea94d0d6ab3ac905bebc2a53d8d952446cf73463a46ad2e4e6c5d0a72b97f
z8d52cdaa00aa30c1988483b3a9c8c33464fbeb82b0569c146f7a5e619214e90ff775a490e8a329
zde9880dc07dbff3d1890f1b983cd7f7de37630740278891fb367c1965b4575524283059f999620
z2dad3c5c32da8df10c48b19c5f9ce1cedddec8775e2b4b3a51a97da008bb043182891da968b47c
zc079a7f871b226f5d0abbd9d727cfb309741648a5494e86702986861b4a8c69a93904b3d1d71ea
z845d8f890fcf088e4bc9686f97b33b0f77082ae2d0d40726feccb9de20ab046b627f9589d3522e
z0e8382524a132f35943b5f778dc203550f151a3d3eedaf27a8cef39458af32d06d3e3f50e80d39
zcce29f5d6e480a3b9a88d7e355ddb13b7e91d481b7e5382b50907b02b8b02be7f2e0acb3e2e987
z3daece3f4d0f3beef62fa8e4322a386d89ba637ffe31b5aae9e62087cdf6c06743ae679216cb34
z9fbf13e3e9ddf15f184e509548bd19da5df9a137b672fe389d4e57a1a8f32f934d63b67d0f61f3
zcaf0483d9b19105315c671c29cc1b1617df132fbf7847f85a45843a1ac2ccb127b62eb333cb65e
z6dd705a97d1124c2fb9c1e160f95911a3d39a7af88f0335e17d432000da27304471940d180845e
z00faa6105a8b6a4143d82bff7f593a752465cfcdc8be7a092c8d07d3d2472f1a8e390d0ac12b99
z6292f55435fe39472f05b835017c7ecc554cbd1732a48f732e3a023277a8562f4869e9216a9f8e
z09e8bdd6030a0449104437ea7cc81b27d020b3c5365aaf80d7ce54ac308697ad28f22cf30cb63f
zee8a294537dd31e796ba8dae9ccec31c961ed3610cf1505f1d231b2d92c625a830e45a4cc08ae7
zb3198073ecf4e5c9977dae85fdd2761e38075c267e652ab45f0db4ca9da664cb057bfd28c28040
z3aa6a8a679180e45f89b6892cfac855794da2b9b83f0a1fbc8973da27c090d7ab5771538f3947f
z16a1542cab722d1669a139665ce4bdf5cbe1521e9f0b34e160b8e2dbd8632f1d15076270034cee
z9e89601609fb7b7216f69184bea7d12b30ec493ea41934b7636a84fa8985de1791532e7bac17f6
z92fd881e03a729a2332716aa4ce80cd7719df20e7b79b763f8428e0d168e6a28b68de6243c76f4
zc459df38e4c05ddbb7b22e21741131ef9978adf7dca2681aba442de2c9e5e2087a192dca7b916b
za48d26fee8a2cedb4bf66061603f97c33525762997b23cd560a62b270b8142f220d28a342749e4
z37c5198552dd3150afff69827bf21fd4f3f8bcf89d5714aebd850f6e32d092651f7c19709036f6
ze2a8b3a7c7fd7724c2f07bc57be61d78e09b72bfd0571955c1756b0556642ec99d391f6435080f
z0167ba40871873f5a3f476688358dacc5d150d160ddbc95dc219cbd2e5fbb3a01491461ee768ae
z09335f5ba8861f34e4dc41f7cec259b170b2fbb36edfe838e2cc6d8442123d302853d1c1799dfe
zcd086dc23d33b03cfe2eac77a0c3f46ba2c70d8e2905f831736180aa6bef6addd78cde1834666d
zc6ed46b2fbbe0d43cc2e01caff71cfdd97855752f48558655a59af60adf01df1ccdcf88196c04e
zd5fecfd6e72e507059ebc4d9f65367426c31662d9b64d00b685f85f4f56682f5476cb49e42b417
zf7f294c76c170972fa0c65ffb19764b293352b9121a47380495c599813a81acadbdd05766c704b
z8ca889c89510e68e60a2a02da464a7ec659b7d27b44f8abc46d92428866b38b7e29df3f4338252
z2f51e4ae0ddb4645808d3c00aded8cd2b9c03b2cefb53417c6c4aa9b78034b431962a247b943ae
z102ca5083e249d8dafc336b7fd6bb50fba457ce3999bca761684115ccb3928d6c12c6b355293f2
z28801f3956b8de2a5ef5d28a34675f92921c3dc8472c67b19a611a281ec2c76cf595f58884535b
z515978ffa78f21ac071bb84d25611a51e5e7085a3617ff750d330bc5ee23019d6a499738919e8e
zdc9e7f774916bdc60788abc0eac9c32b67976255a78d06832b13f8a708577e7e3591a523a6a131
zb83daccfdd996ef534e4fc3fe7d9f4a106c0511eb56bb23752439c2d24442bc9407a0d8ac5ff4f
z214bad907f43a0a382522737a8fe5b8c64fbedf642348f1483b90005bba9d06a8daa381fd7f6e7
z861513f08c98834e8bef52edb4b57bb3bd6bee55ae6d971cd68223acbacca1f26f6107c767e82d
z110fc67229fb520fb9f0faa6407e26f1b41d5d580da647cc3bd0e9cb3fe3a54eb273bbfa17768f
z4f4904d7cfaffee72ef15130575e416fc2aa3d9680fa00879901680a5b7081905997cda6a15c72
z108527eec8f8c68e4e751e706b55341e4f23396aab67c650a5721798d1fb1366e7bda445d0ac13
zd805ed713092629c1f241619022bfb925379b61d29472dd665e5c108b6591748d43f3bb2eba307
z5b72d84cd68b1ff3ecf77e3367eb5e4af9adfabf5f32d96370f621cc20568b84105e85d13b96e2
z02e798b8d64c43d27defed3cc48cd0b92f6ba0085bc5bc0369ebcdfaaa52fa5afa6e62cd4e0edd
z89018fb94185fe6a5ac52931a36df9d0d8276c399f381d984742c2fe4e1c72f1fabe9d0dfd93e7
z123d0d32bcbbe516b5acc70c48511d5ecb9cfb93b7b8f513ce6dc47931d809d8ea977a74e6154f
z8be00af7e692b3e979de7ff29d40c9996a4b12b4e84c77ae45a21151b031e65f57cff046c12c25
z8c72f957be207f28febbecbd2304917e91ee327570ced5cd8e26b058acb626f582a47837adfebd
z750ba431fba65d9f68978c606bdbd32325acac6e24d4f72d1fe4957edcb16d350bef66f7ade8ac
z7bc97e3760bc9cd3bc1d4897f803ab148dcb70433c0e67c24d023662a296692804ae5435c91cda
z2d3b4124e2fcd4ba409a61ed4c096da5a21f45571f1a88e0c00f08877d5974144df6944dcd57ff
zdbd47f771423ca4c06547c3aa5bf2dce08b27fa1efd6da2f965ef08c589e8448b7cc40fc867fbb
z455ee2d2ffd6be8d5f6ae3bed35d52644c950778384b8a8f837c9ffa9f40efa282bd996631cf30
z90a48b60ed2a455e8df8f1afe92cac9d3f2449d58bb1ab16718ef3bf2cd346f04daae94a09c80c
zde2c46a4de7f5bb1c841bb0265c7c34e1fc9b737cfa793ac03919911f1f062dbccef35ab674cfe
z338af533ab819f05d24d3229f1d7a2f099f4b3dc7af1f15b939731841852f8e61c660e809d1f06
zd8000ba05b578e5556ad419764b20de9703db9c4437b43e4d50bce10713ed4cb3216034ab3f255
z4f600df2b145895e55c01cf320df42099e624f9c85c7c8b5be691a40686205bd64ac21541091bd
z3ae3ae39f6f22032239146e8c0925ac96a470810f9473ee29a287c0aedea9cc5c0c8636942b466
z2e0a6c69327ec024830ec8c5e0ac1d6ec2b3953794e09bcb6b7ba31a59afbf5d5861a373275b66
z4d2ed935b0e5ae24a425fc13c95d8561a3c89bddb0ef1da134e33153f8c2e38e8d08360b6d454d
zbdda561f9da2980f636e3d340cf532b4312cd5837b68571ba597440e5f198b64b4a3a8d561741f
z9788da58fba1bbc9a91afa5614beb24602a033364036f1cc2c41178711f3d179f5ffcfe42ccaee
z8045185691627792043747acb820ff3c75d6e969428c643fead2adda25edf40794217c6b823969
ze5d5a4a25a6635dc44357ae6ead2eb3c2b9f1b9466ee5268597666f875c206746a8df4dd3ebcdf
z9062a0a8ea1bf2ce76d714a3081fc44b2e1ef2e6f651ef57eb8dde5b915fefd539e8f989a9b0cf
z3a8d8225e3093f744fd9808a33ee6b6e1d92a60a06e61223708c384cbcc00f8ec30fd73add2653
zbd2be6e049cc33ac5079e51932757085804db6b8576dceabf47f1ed99fcf55bf248d4782e7d059
zab7a9a0c2b5cb2d8e4ebcadec86effc354f87e43920c707125c5773e4b106570e826e36e1ef678
zdd3d7932bb33d6b54a0318d4f78aa8c901b7b608432a87ffc09c3e76eed881beba35ea066ef64d
zd7c1808f87649ea4eb9e53bd174ffb5c5d190087c088b1aa81e72a4e0d1472a36db5851749a683
z20ffac1c2cddc604b8d374f12617282de56bab6a4d31acf6c30a0048f9c25e739510ddb74525bc
zc29bf24d6dbdd84dba2f96d0b4cce96b407961e94af9bc1fdb109e5e834efb8d0830e51363bde3
z75b3999188fc680a8ed59d41a9c8e585407b8a4fc0e3f5e73a8b8d242fc39f4df909ca7f96a647
z4941880d137daea825ba66f21cbeec3682c98ef8f4f107c5d6323c3a722cb6ce680f9e89615e32
ze653fe77809a6062c6fa8a09f66d31bab8ecd23bf66cda81deb0a5bcbc404a7f1375da166e2cce
ze561584d68c39414bb7303f68f70790c02164bcd86220174140a0ea7e3c5646a3bbd69f595a26d
z15d461688e4b5da9c732690ff5de5fc1157fd1e3beb4797c4fafe3562308c1e2982c155c9bd247
z3a3a7f946879d4b8bdeaddeea0f37f4aaa88c1e9f6b4cc183191616ac85dd6769a58992f5c5dc2
zf895435aec17af5c5d4393ab851959fa7f59b18cc15c422a13c70a3eaab88887720ed855a189e9
za0d3e359db41950b712f6b23b0d1b9ec687a4d32863f4b7d39effc4ec2cc306d835af824ef0ba8
z126401287bf5cd3e6641a75a59e9ea0cc5d36c3ed41cad3a5567ecf7e6ace725db991a3ee99e7d
z46cd18c64ec10624057cb9d9d7933f2434ed29393489720e74e942825d6c9cfd98a2481ece5bce
z694bf65281e328a6844eac68fb816993229988f9bdd2877a2a913999857b929175f322faae5f3a
zb0733c44d08012391f56de9c95dde7284c29d203c2229cea4b11e2d91f5ed9d94239fff7d22142
zc4eb1971ba8f55fbf28cbfdcda61ae0edce1c55c744070f6bb052b77fe57a3ac86a449d75461e5
zfcb579017ecf5f2e74f20e8c2becc581680b1864b90bb94c7dec17d89768dcac2524420cf03fa6
z90134a6f7f85ef3c17eff8f5e3b09276d942b89bbf240f55e1a68a9acfe7d1cb0c24a009889d4b
z012195833bcee2b5c9ef5d55c374b7be2b99effa89735da88267004722d003573344433091bb8e
z6b1d911d19fbdd67f846f14eefc3768bc35f4aa5fe2a5cdcc6794e00d428f649f7237eac67d34c
z1bf043c8b20574dbfc15972eab752cbabdd3551c16c3e5a58ae779cbeabd2406341f434cf27fe7
zb7eaccd53cc7040cf40302efbe1111e54c73b0046ec83fd3f52467f7f99f01c71aec5c191d0ca9
zda75fab8deccefdb08d4ede84343ba402ede6ef34aba1cf1665c2caf205572ff37ca881dd97976
z6a12b4cea33ceaac7d4d891499783c9fc8a3b00216a6fc293e766b498a6256c5637363164c0dd9
z95e11ed2e3acf5b1587dbe7015e6f014f687349906b3d73a7612647d6fe9855c007571770e9ac5
z92857994d728270f0cbae1ff148a4c69489d4541fc5d6842523224f1a86b4136aadce862d9e001
z1875d0b4b95aca170a698ded4ea1f9b069e3aa1e10e76fe898dbdc194eef87eca68faadac8c189
z11cf1de5ba09a7b841b24bd5128b966258f64ea9c641de77e90bf01b6db2c81bc4b7bde7037f7b
z35a111d50e5882b44d99409e919d6eeb6b4d724ad75f42e4067fc0143e06ec947cd4648fa79bf9
z5313d661c6f7135c3be32d6fdb3191b3bb40c54ca2c2a9a97eb9b900edbebcdc6ee8e03a066f92
za391cd9266c8e931ff0b6a39f7c46005ab86c18bce860cf8f7d019596941cf299e94b10f2164fd
za272c1731a5f88da524cae93223357b28b8156806810f0ad14cf73642d1313a0393a8b56891159
zc3880d7edeb9b757666c4881445757c6747bece8c90f975c0c2e31ceab37b6f7ca2431800c2a56
z4bd2a756e5f6679e50e0458bbdebd8e702fde67d0209fb8965a3b3c55ae4bb66a4475a3030ff94
z9a8ac68cbf8471c215e8788adca31dde4a633f0d3d98d742fcb43a68ec43a7542fb4da94de18c0
z76b8ab38fdd0d0051e455ad0cc74da7a404f203751381a6164630a95775dcf69820acd0eaa8f2e
z86620617e8b3f8130823a515b3b26037aab28a159705b799cd0496777f11e1498dbe81b72ee0f1
za83ca8d29b3f5e8f10a04e0eb6e1f8c5d0ba192b4584dc4407d959097fa9a9f552a735b0500ac9
z2eab0a8576b5ec80ec7bfcd5acab30429dc01056a1edda2b3a1e5ca562ad58b3898e6c6d433e97
z0ad6d9daa945fab20e5eed6e5ad606c397f9a467d983422a0efdb81b54c874ddb8a8aad7e374bd
z6609d963d41d9e0fa5bc66cf031a32a5d1601105e446fe829b16099b8804ff4027cff71ac27088
z253883038cc06df08764363e9b0377a44bb56cc2ffca6e6a8c12755fe0c4c541dcaeae06b2562a
z81e36ab434001cd907358bb089d16f314b847f4f4c595dbe2abcf0f4789bc4c0e312de084f313a
zb52b543f3787d9c4bb943562f0ec91f87ec6333b874f55a541e95fb555d9e9e4210441a3befe9d
zd1a6f2ba19619d39bcad0e3c0b620b28215f672297c129f2b42a975d1b3d7186fe0a958e75b351
zee64b77b544aba684d473c3d631e869eeea69b1f1d7bc647a46848475f49bb40b0c128b0929ea1
z81262463e3467e77959c5efef65419a8996bcdd68efcc614ad383b56b8e7823a3fabca540f5e55
z06bd5344d0e5abf73d3f1c30e8208e9c26587f8bf7c9d2efdbabfbd96182bff4f56df171c21364
z1cdf6605645e4beaabe27f5a8c677149fb8ff7f6425b6f93a503cac28f1c8472f8c05ea580b3aa
z7bd279c210ca63f4b3f7bd623e2a400d112e6cd598d9e602e99bee1fddaa70392e41f4f272caec
z511a0ab5de09e1470bfbf3aedd33df4e2df183d77b24e577ce238b2a1bc79de950a4d88f5c6e24
zf6d5a3f46915c03c4b8b85d64a8ecebb13a0a4a9f101dfe827d7dd0e7d6e82b421f7267af8f44c
z3d9e8891be1432de1b24696f94260debb3a0d42cb5c207a0133e16024da113c752ef3cd2245d0d
z25066b8b70cd237c80810fe19c0ee6477bd032d5a5a20be11fa7daafc8a74ff9b00c0bc6cca6c5
zf2a16d22976aae0f7d1140c73c31944cc5b5ace634df77e3fa62380e70badc4ab1f37bc3321111
z94b4bf548c83c36e00b15d1aadb00059f3727cb1354da0c101be94e86a45307052e31177febecd
z43e1e7aebc7efb922dc199087d2b2423423b85cd38ededaf71514ba91f172c85cc63d2a85a9b81
z077e9cff8bebdb5c76cbe839d08aab6e8d9cef01b9c263de31c998fd8652edfae3f94a741776eb
z3b228e920578fd134ed9be9cec26e6f0860a609de24ab9b94d14be9dd05ee2df6d373e2ee3d9f0
z259471174c8ea157d7666b8660e5ef5e11458c0cee6c28d36eaf6e112e2d47d1e47410591e02a7
zfabe57a93c82210d4c508e41f116a259631475df32468ec68a9132417bc048162f812cf7edcef5
z6ba7e83a140e02175284e0f2f3689e8c0e4d5fb616539dd31ee0cff675a90ed67972886a080cad
zf7f033cc3b9c46cbdc46ff038fc6d4d73c1d0960b135bc1095bd9ba841ea2af2b0093fb60495c3
z1eb9a74eb7254cbdeda47b7a67bf8a504c2da08510cb42d3cf30b4eda6dc915619c3057a7de4df
zd9a5b6d8d8912b74d81fc55abcb5745981274e66dc6d74029c5355ae8f10ae63023638fad2c489
ze2861e0f614e9e5c69c82d69b35dd19d89b406d53f9cefc9af8665f2cf49f31e2993fec2832e4f
ze3511f759b00924d7b75bc4c8014cc64a582165f56c8e2cf70c739d4a8e05f11f28874aaec9b28
z7065fc7806972d883d2d20a1b4d5c37be7fe46166093c2c1419abb1ca2ee4d27f1eca3a170b960
zb57a72eef5f42204dd9f448323c186673a2800663721e11050f0901515e310d44737722212722e
zdbdf26281e994ef8c27a6154eebfd2a461ffacc8930e29eac52192d5212958aa8ce6c0706f85c0
z9ca9271d37d78cbc8a81c03070ae22636048fac4cfeec6995333b869c2322e78872cc75d04d337
z3b0de1e15bfbe12ee0678b0d92901c07b5b9739870fc7ff95e659d72cc8129875085e69f32cfb0
zdd2c85bcea8a124bf2fc88219155d1aa817d974c5bbe84a2616db55b5faffccd23e77831858a51
zc7a9f69cd1968cded6fc535d13c9309c4633a39f484cf83b63a76e5577289fa8515b6c8d0c39bd
zacfc3e30d217c7b1cef97241ad60501dfe66a5a133cc15bbe6f8882e1b6b10ea4911101c6f4d60
z02d1f423d4eaf819e75bc6e458befce3238c5b5c5aa02a39d3066cb6611995f81522e7265d7de0
zbf7edaa2ae9fc1b61053eca17120ad68fac883a7671c0033bc45c15383a8b05b27e1882037aa93
z9e702722af538b47cbdb1d60622684747d94365636fec5a8d12480df021773765f8d09fe7692d0
zaca4ad51adb4c995e4707ce323a1c3e29c272decc8e7cde12131e8d4e2869cb4f570a03b30925d
z0c0673a152732312f9cfcde1ba21ab7fadf493fd3bc30350dcb706c653b78f6d53a07bae7c15c8
zafc2404ec03dd1685d2ca98d838f8c9d97fc67497a6d3e52338fa9b47c28165578b01560737d31
z3293a07776e89fa57c5eb10e8d751d1c432b9933e819b0a4ca431136bdc02bc8900c8e71023e72
z9b22c4bc5f5e249b31d5a81cf1bd15ab477725182b3cc28046f038f285ffd81f7decf326a74880
z55b3a84b091df8a64e506b74eef14e85c5afc674d63f3dfe60b1afadc4877c9b53a808e4f33d24
z4b58d3227e42756ebe96f7dd614744c759aae6dad3979c9a2a24b9e6db3c702c23e7f6c28cfdb7
z7d10c61f6c1c8a665f6a137edd828c0ac4175b0f26ecca4295ee9a7540fb89f3114d349fbbfb0f
zc9cfe01ff37d4c3b3ede184c11a06be7e0a604e4e2b5e9ed4fa6dec71e626fe031b59a2393d7e8
z5cfdd7213dcce3c04daba00cfffa78ddd7fb0ecc1f2bc466c178a1fa6ba5473bd4f6f287b47e40
z1179c3161bc43836ba84a66a855009cd278b3767840f01ec6ae3d0addcd81d23ec271bdfb49e77
z5ef64bdac999c22d28ae19d98c18878ad4aacad2057e4dd9fd64032a135fda2ab2c21e09a2e1c3
z71aa94e19fd472c252770a0ac781cbafa7287721cd84d78dd7f84190261110f3db8dab4c632d22
z7d3db5974bdb1654805fed14d71e8e96489d556cc49fe8853d8166b2597b3e2d343706eb830a93
z699b5ec95bc51b83df6aa07ab415a20d028c8f66f2d6dc245447df71813c287e470dcf46e0c195
z18f8b92c59ffc24a127a3bc32b6674beb86350f6af967bb8935cc704e845b0c04d84852fa676e6
za0a330acd1deb52ed05913e4d26a9ae38ed2661403ab7941bb88c601e20e124d3176290d957d6e
z478bb956e15324deade85dd88d58555c8c6ca793413d077c4f60be9c141ee79ab4ae374ca8d0bb
za7ae3297bd63db05c8ecdea3fa1cc66981a0be06e31a8436da215f3225714f90a4aecc305ff69b
z8043269baf08064d07a93a0b268bb135a971f7bcd1025ccb6b140a5cdb965c1192e28061a55bdc
zd4407d98e7edfae76f87534f1ebdb5c02c8964b08a720c11582f0d70b984a65b87ff1e6480f738
z151260887a452242d3a4404b5f916627354c81162349de31613e647a4d715bb2f54a3814b0cfec
z89393579de569f38993f46f9ecbee2c39dcf89dbdd01b9d425f9cd53c52a2a75afb20a647b1779
z81ef9fa0d2cdd37c941342ef735f420a6f1a29b854304af2953fe63a54b6c9b440e03319d40b80
z5d7295eca4a62df3aa27a55d1781b49f0d0ee55b99f2eb164759bfb664587e1835f3f18cff3f45
zedcf3a1c130aec32761a121d3fbb868250eaf5b2da15ca295abab7b21d3ce2e46e265521e92f5e
zc93cf6c4a32778e24b29b936189bd728ca638fff6f6a3bc8d4de524ec1247a6a07877efa3004e4
zf9e5b12408b3f61716eaae92dabadd8166b9bf1773191d3a6663c106df9f274db21e0c0e34617a
z5cef91e247e0985efec76d701dda51206bca21b9d9dcbd8cc239a7c4dce287878b74f8cdfa211e
z5be71456ace703ca312e3059e101385e5c53b90764f10283f0022dff5f914940538f9f50fa2d01
z25c16859769363fc923459defdf88dcb91f2fabbf26cda69e31d027c2d06096f8be5abf320e189
zc26eed97bf5e867ee67ed57b973962181aae94f4271e1ac9556b8fab8c8cc71b1c114a7bd8e609
zcb085251242c366c8c0d4ce1b9a519027326247b05d456f772bc835277a887a54de6537e6e1324
z2ef23aebc2cb9f98384300b0a1b21076a129eb83401ea8e4815e25a48f8dca396e60e90885cf75
z296695b938115e76aa42ee6dcb5648ee2b3b5caec35e731ebe2fb60627db538c3e56fe8694f665
z0cca883240945cf70390ffcd9dfea946cdabbcebb1bfd0de77dbe723fca2ebae6fa00498bd4287
z2b1ac95e52c8db45913c981d27930b66ce6f62324da48b173becea931c71409daad1d19bd66735
z1303cf8f4086a7abd355bae6a37b5307c26fd38075a5ea7e5f9807cc3a04e44f07f0f3d1540d6b
z8995418cf64fe1e6165911c780cac44bcd8147e56e7c6aeda69440075ff76a0c8f2873751bf3f2
z8c7e3c11957482f83752c9e1374c0597d3f2ff5229f52cc25c3059b5abf6b613b4b58ce32455e9
z422fb5804d89f3dd34bea90a1ba4dad38897536cdc42d3aa45a82c2b9c47d21bf5c58756d3f52a
zef7e83ac9c8d86bde744010359fbd0862e56c9efb3d7b8c737d1e95b8170b4c12865bd16ce0b15
z1aa23109a15f6dfe076dd3091276982862bc42fc28f855c542b336a6f167c8eabe888f28aab745
zdc0de8279bd24a2aa0cd99f715495a930379c8f8f4d9fb3ef5f4cd5b5b9ffa05cd0b62b885c22e
z93c84767ecf6abc586b345a5be57e6eda6b98a1a0dcd13237ed4c81e789dbb78c1e213931dfc9b
z13e4a3ee94a0f41f0f5d7c6ac73f623a058ff71584b1d8baec6237c100038931f14166355a03ac
z25a040c08ef13114c555a0413016fb994fbfe47716fa31aee713404abd011d8913de9d662338ff
z4399d9935b446418452d75d17578339f24a9130eb4115ebdf953892854d4c1725ad862d4d2a019
z93bfd6dcd7b2a370a6ab09da6afee91689863bd69ffa6f778ef84df0f98cb25e3c07ec8fd69beb
zf60291d99b831d143aef80d428d510f62a81767dba9e07d9a9e9a6d2373ab201fba0df80d50d4a
z6224ba3d47c7e9dc3dfd27dd033a9945c0c21c0d750941cf24cecaf742fb4cf4ab46c8db297d37
z40e690e9f5d7c36717fa578e486135a002a9f3c5a780d4dc240e825d995b73382946be73bf40ed
ze604668e231764745c2c651ca83558679c445a7c4a171f4080af0c706ad9b9e7d2a01d473a2c0f
zb7a9b7e8c963b456a2c7d2acd51069fb4763072337eef2506dc8bf4b20cf1269c3ee4feb87b014
z4e09c1dfb390de05247642169510ae092d4e58ca8805eac722ea1c74a72700da7ca8ef3f6edb3e
z33ef746151027ddea1782ede6abed6bdb1306790bf1f44db1678566e33ba4c1af8db7b87b445f4
z7c1177002476445f11c2d0b740d374e9ef6e21b63cd5801be0f8b255ca408348656028d9c72ef2
zd6ae81d0049001752e4a1602272d21f265b76b0df5be27fadfff5d0f71a14aa1ba0af0e74e7c78
z025e56d5d174a84e5ef22610eedd1b552c44651eb4f02cd0b008cc3f5b1714c6593441a0e19c57
zac0147f0790a8077075bfd3046215d0be3dc70dd2a656331448e8842029a4ff6db763ec3c50c5e
ze42264c21e0cc0d9eda8d03b0e4fcbbd4fb66541628180b0aecacd9aed91ddcb6a33de92065807
z416f78f7dc2e678cc97310a5f6d3cae29fa2ae8fa3d57c6ae0409b86e73a9d125bcb6f5b3da1fc
zd948bc81e039466978285bd2b462e3ad4135cda37d8eae19651e3fb8171e0dd7d08359e16eb3ab
zd1e8a0698d326c84b1fc3188fe02b62a816ca1ed297749f767ec87923f7c30520db5401528f14c
z4e2bdefc710c293fcf46e456b04ee93d6514d8e506e5f645c773bf6a80b73a13e9feb6af539161
zde5f71fa769ba4138b13b2aa5f0331762ae7b70b5819e30c2763fbe8ccd07f3167e198edce93fb
z3fba93d369f11dc87faff779de1b172fe1aa3d7493afd1069208530ec340cdb813f013930d7bbd
z6fb44579c17d5f1dc1a223ce4a519a56d7f4a6e298ae3efe0cb617f0057701ed1cd2f5a32759d6
z071a90c7002cbacc7f41d089630c6b654d29de9466dd6b535ef95b645d39f53dfa594cfb39fa63
zdb04173456f87ae56850998cbc901b284b677ab9c8cb3ae0fdf9ef28a02e127e3b643eb83bc490
zef11bf2a323be4fa25954f90fddef04edf022bcb53740e629391a8bdd7f282239f830a648d777f
z41fb1a701f803b4ddf9f69b73f19c56f5a4b0a48859f1b5a71d220545581e15e454775aa4c8f58
za1e84567aa14c66f90d0e5223f3f8ee66ac960293aca56df7d2f290025dde9531f0fb5c9b0d949
z9c0c32add9e541ec99fb773af3bf7795d3e75aaffdcbc2875de01480d28ca3fbd95ebb91482921
z5f6b0c2c216b9bcc993e88bc2c05ae75b0053e8966601bed132fab9aa956094731488fc8aaa875
z5ea0a1f2b68011654511369411d8686660c4dbfa13beb9f99add62a276662f16c7c68f33b33ef4
z6be3c2913d2b2ca2248815406f990c72e06476c4c2391a2a810113f81f879976a4348251346597
z7c1e610af7f8c8d77099a26dcaef94874722bfab41a1f7ed5aaae788d9e851e8ef138064ecc099
z972ddc5984f3bdab51d4e25d49feaa32eedf125c2fe05c81dedc2b5ddc443f211f19c298b669ad
zebe4b07466e8383fc792fefb9159e4803cfaa374fdf7e7b48361b51e0a2688706e01cf65c9e869
z22370d960aaa701270e6eb1072c450ee51aa84c30f50b99210cec71de7a98e33d820639de170e9
z3bc962a618adcbe65c0c2bec4aa8f27a6801faba4c3777e851315c5b1cfb5e1342104ff6b8b6f2
zeeb763147fcdde9f2b6ed287d15eb26c9524c8c30a8a950894a90a76fc580a7b7bcbbf0e7a1a8b
zf8caba5e0bab537d62c47ed64ec1be733c04cbfe4a1e288577aeb58de4656e61e2285ff18fabb4
z276d83a3ee0ec3cd6b51a2e68c711192bdfb9e2113405a1696c413e41d7074432d88625016aca5
zf5712185d9cfc6b45f00df7bc9419f5e1b7493161ff84540fa362913baf809092a9a5919437c96
z65f1913b77abb06e8e388481c0860f20733150ef621dad4bf51080fca3ed69f295a21db077f0d2
z4e9806946de6e21e8cfb83302f80f0c559e8a4b17ed1a17259c16d5be01bf2f0d3dc1b82456cd6
z6935f449e4c6da383eebf3d65cf1eb6aa05e07e212f264a19e20dd164ece81fba154a57a385afb
z030d21d45e708782185ceca51a853ace6802c2f760d1a9f76a9d20912f3e4964d11479ae90a40d
z852319ac931a883931b4f437fd98dc569033097bb5efb34a9f2ce671ca48a3676888710eef1734
zbed9b54b6c3f9f1cb5d054fd3f645457aca18fb84fa604ac6a5a2b7a2c1c012ea54da0be901968
z43068748dfe4f74e4e07bc867824e8d79b3c5f450244b0ee2bb94e6d529645455039bbac0fc519
ze0ed102385d0c3e7a39292db6a57c8e5bf000ba18878734fb64f89d82655facbf223492bcab279
z7a0631bff106280e60556920f03644b7a1c8e3907885fbb8aad7d7a3dedc696f0406330b963c97
zb19fbe539913a4b1cf419678838dd2892d28060d747955e009e018fe8cc44b6c2db8600dbda60c
zc81135f4f3b42ca06b68f5b3d4bb8908bc72be6100223ee7c98227782db0239f96043185b3d2cd
z3921d0ac94ae656a61509ced5640145dc9f05d8e44716ad66525c490b57d3fce4163c90a1ce5f8
z23ab6d665d1b0bb1a7942d8f9ff0637d8e40a7289e784e9e623bfd8610ece3bd76680b940df18b
ze3c408706b6c827320d738aad7ba93a4a4f911f3cb209c17cc43c203dbde17b2fd29e605cea0fe
z2675e69d1982d4ff8ccf6ed984679d777fbffe30892f1d141b9ea69c6e98b061bd45bb4f0c2d99
z4c33081012e0ea4765036a4ab9e69702d59536715214bc3e5a3df2b84349bf1aa2c676044381eb
zc53cc39d40ba6431fb435fdbee7d215a67e0780e2fbd07b6fe7ae0c0ea373e0703e2406493542e
z8ba62b152f6f16063732a33de1f20944eee49325021078b0aed1fc72c598b58837a0d6e182a887
z83e4dab292ac872963428650b5d1b9e0c9f8b7741459c546fa05cb77fd05c62dcd255148586450
za8825855dfeca9d0c485e9acc5bb465a306f1de3563a2fd651e32f1c279cb2ec9971354a414547
za37cbd2fe683057fa9f3f6ac63d70b50bc3504775c99fc778be5444009cdd117a2c0933aaf89ec
zbe5264970d4a4445ade31e4c692a28f68cb543736ccc1a4a3cfecd212abac256da600043da9310
z3b3b5aa632f60c91d3eeba6ced40f546848b1d0568ac14e6aef517b0852119cd18ddf0393cbbdc
z5306491356750e3b6cc53731a55598091cf3a4c7142f725a72174a6ffe53d0bca1f162b7b6e2c8
zdc2a1fe81788cea2cd21a3e5c0865f8e7e6dd423f67162bcd18e621b82e19f994c185693789c1d
zf8fb5eb47b9d66c65a74aebdef48e56f7e34476ae42f4033e42d0587b69fe5234a10f84c59f548
z4fc6e4bce24c8d306634b00fd9646cbd32a2ff992dd89561a4efeee61e01fb4460513e2f1193ea
zc407731159633171eb7f99a7215697a1e70894f382abb824085b3b73ef7469a710a6026fc4cf23
z98979f177115ec3ca2e9681ced66af018b021782de815a4bbb7054c5b4fa0ff0aaf92e7369acf7
zff3e8656500c02d67a5fb3211ec8fbb77575935ab873cad8426b2ea8cce56c0e3dfb94af0e57e8
z7b0838686bafc38ee7a728894ea7d83fe486b2859c47b9e059ffb1b833c8fa0f22a4df9ca52714
z0f1da992bbf0a439f1a281deacde27e884c14cb64398bf2c4d21c7cbd99f72ead962cfb3f0a5d1
z162e2ca84de10434ff8d57886fbd4da82713d8ad728f9aa058240ba1729c8a9d034143dab783b1
z188e755f2e45715e7bc50be4effe44439e14662e9f1d38bb43676869b323b14d01313b21cf4e5d
z82d5b91f7c5bf1c734081ebd88795c701d43303c2f11cddac94f11ec8db22f72e608e4c0f65e66
zd4d7d97dd7474ec86596dd38d89834bccce0516d87c959e04bfc58dda91a81ced30795c1f95fa7
z179089a534bca205c0632ebbc6dc058c670a843cffdc99b2a412469c44315870b775454b66cfa0
zcaa33469cb045c898ef5238260171c0bb0d68b5603a5bfe02518a65e79638061c3af5b0faebdf0
z857d657daba1e63e8c8b106a4d2469ace75a9835ec026c3a457d71dcc50f6800ccb7e42a2db39a
z66bf3a96afe24db75143bc68dbc885aeea67565f6b25fbb03c090948f708369df005a5b1e12366
z61ae29c81acecab627e602ff0d0bc5f607d1e7c5123df45e43f30325bf62d66a88e6f7d8c0a3c4
zaa71ad4287621dce4471d28cdebe54bec0c288268b1fc237f58c22d74860f09051e10e97ecd3dd
z170cc33e4fe72d024ec6396e4b172255ad2ff484615349053335dea531c279387edea769037221
zaeabd2bb061cc667268e22f651b290a06415956e8c19e1b141dd2c2a8c3a40f1288f514a19fe31
zac4cadf26590f3a960ab264b045d8fe57544fec51156b4f2a730ebc7517a65f0b48f426ff1407b
ze25c3b8190f33c3ad291cb559a6d6d8db2b1382e49f930c570029b286d9aaaf7c84590d5720bee
zbc0cb64209f9e21a8d624af74bfcd0e64590ea634eb2271c4181aef9802479a9f7703d8f9bc962
zcd07b6806fd6b59472d963d16bf5730a80658ebcd39d78c9717d32d17ee0232921f971fb2d249e
zd8c80c6855f1768c7741ec5c5b8dc992eafe4ad13052b4b3c36061741d38ea6a129df7a2923782
z9515d1c56adec85c5b67821e3ff606409ef1b2ca6d795a265a016c2156ea680872bf7915a1dd7e
z874ab91600326b091b4fdf7a8084cff808cf2064c71e85facd15fd0b5830bc9e61cb5bb6b3e1db
z4ad178f8c9c119afbd48393e3dc2382062ac547f15c8340325cc9bd97b5885618eb3adb2b520f5
za854bc784f30171cca80cd666c34e19f2eb9a7827816d6b4da9a7f2e51bff46d3351b32a947790
z6af26540d80ea35a7c161f3f4fba9a71cc2368ad20e27f566db8ca191583bf8316fa7ca0a24c11
z862e19aedca0fd75f730165e683276d91294e272ab3cd7d1fc6083e8069df6d6461f1a4460e4b6
zd51f7c67e4bd4b25f91653916c84772badc76bbde4fa4fc6585dc36d0e9002cb9060ee99563e2b
z46dcc44bc0fe65d12afaf6bfd3b53b7e8a717cf4aa7f789ca6a81c0dc7b66d02f72bba96743893
zfb58fc9c13fe38b4be213a83c52f26b5550730b9b750998b9df21783c8438cd91fb349a531f49e
zbe784f83bef12fa05214873582b47deefb2c65258d05824a77fd484337f0fbf83eecbc4ac0afe3
zd223ae3c6fd0b242fb37c94bfaff6b52cad6604774f5e3f056b35d34cd410e0d6eb4f76809c967
z4ff016e88d7fdfe23c220590cf4475b8914abfb71d945b23fb6c5d33348dc63fdfbf3beda12f67
z5fe6bafb8fea2a7212bd310778135dd21bee08294f51cd78ce5e1028b2babb45c6b3ab6788ff6a
zf2bf50044480324769a23fbd14d66f3e2bb455215b517268aa58ffcbb634481dd3abe989fbe47b
z4d8cca94d073fae1f2d300e5b3d0e9d744740ba8e19aff622b711077af95f5f226afc998068699
z6c5108f75a366622a0d3420eb1c4c05535d6ce086d682f65a42765011b8ab24900667cf2b8853a
z394296ac5a5f5d4de125fa22010b3a701c34caa08a3ab157c4e3cd17791c098e4e131d4d9c376c
z6b0f146631a3f2b14182b54e20b368643e7f8615b569d8d610dbe52289301dff7bc0219a7ad611
zdb0bba79489db11830c1cab87d0d2e7340dbcf2625ae5be6745668f0a4f1c11dd64fe8f952bf02
z35a536fb3c89fba9a257d7325640859ef470da447024d539235612ad7a34286bcbb7b01d94151a
z4de78e04f5409657217e7473f9cad544ad1e7a545ee2962febeefff9e74fa266aac87aa66600e5
z9c4c74688e4f712565144abfcd7275e2da77847eb3d8b63c6438a2c03da9ede2129d9d02729f83
z575d812870d8ff788e1422877b0034c0c6809395f775314043986fb5e3f91431ccd7a8b31266fd
zd4b7fc690062115a2269cab928ed1ef3dfe1e15bb7fbd016c7fdab948a63ac307c9940f11f43c1
zcb90bb7f78d3cfcdd82a0f635a4eb8eedd112237e6c2a6f8fabd6c88e471f9a0ff687a4ff38467
zb1917c764c482ec14da18221c528864e6f0752e43f909b9aec033b6feb92cccd5455e7242c3dce
z706cecad700c305451dd7ee6c0d1c02b7e2b96646d65a44264d344653b337acdad487cb920730a
z5fdb94764a197de17f68128b62385b611283c0860e9e5f8aac6f9ac02b34cce6fff6b571113230
z3b17cb188e26fc4fede38d80439334a1e2414c6e612e0c680defbfcaa9bddbdcd2572173f527cc
z2c254f5afba02e5cc84dc9de272165146de02d310ce69c964999195d63da22caae5a5ccac6a477
zaf7ea3031ea0ad5069d27721ecf82a07aa15ed7b01a76afb300deefad5d273d1225b780cbbefa7
z0014804e557abf3d3df0ae273d3d06ba9b0f6360e66d2363947f548427c9eefac90cec956bfe1f
z406e2671409f4fa1ae74131d83b5d7ee7e2f58b6f4e4bf396cad59ef716f0d428704fcba97daf2
z7573e3f2720b2a15cee9f768c1b75b2677e61094ee0dcaff2844505d99571b9689310e3af2056b
z0c9b62c157a762e599ec71d402d1a4a8deaf23770cc47b5c0cb4ee5ae27dd405186a5248fb2579
zf151bb0a66747f4d9d4af648a2ab9ae6a49fcee5ce5db6ca89e38169a649169c93ab7c2ba4806e
zd9e04dcfcde653f66dc3100f74b2f9840c36ac02f1fc39fe3c232776d3fc1a7f5e25a03967cbf4
zf44eb9cfe9da72a9286a58c4030d9e143d379ce75f7ec1bc04d4d4211da9e15e6b120232335c01
zdf42eef510ef3376a45b3c3356e246580e6bf2b96e8a27452bf27eb2d69e803b5623cbfe330e59
z157accc4de96352acd0d6b0109aa8de44fb74f71b6b8b0fc130762c4480156c2944878c80d5e0a
zd183add05567da0d04f6b88817e7e5d7de1c97f7c3fd539a191d86e3cc9f8ac739a86b18eb70f9
z5a6f80710f28f4e663fae06aee72683cf26404466cea56172a21a8c5a0fa1e483eaabfc98f061b
z675b255366a2f078c24d2958d37c6835268e65174975ba8b22a1781845ad9a1ba191284853a4f1
za35529723b642371ffa1bcdf901a6f3a85b4a07c65330524ee45c5f10640a0ae7af789ba65b4a0
z1016cd0af1acee4f9b70ed5b298789413421b63cc6b54b40f6fe1f7fff49a7defff514afdc0652
z60089f23fb4863a491356485fd6c1fe91731bab04ab72a9b50726563b0cc70d2eef7463319ab40
z5c76de12b07ec8c4acf00030e7d303fd34e940ba60fbf7c5f232c8bbda7ecc4b0c4157a0e83b4f
z18dd754b7df26f3e5a71b16e3a24f7ed009fb3876c500d90cab9ed86b7dba96e732d421688f395
zf86a53e60b8509137beaa3409352b33ab88186ba70a76876c799f617e89914111d0cfb327c6c61
zab531add25348344e71b808c8482f3be4a602c259dea6f5b48f419ceec4023ad618d86989ec9d7
ze408b4e859575d1fb7de537cdaf0fa75f20d9f9bca8119e67313483ea549ee71171fc7edae088b
zce91a1b747a5e2fd72a094376657cc156e4bcf2771eaea000ff0ff0c76e055a9f39cb50596bf63
z886e0db07ef569a01888e8af6f1dca48caf55f21d31bde32fbe2ab27997c771e266219cd226d29
zd9b1bfb392b8d4fe9f5903372df5f4acfd11cf3f1d6aa5aaa0df0850f7977b7c51fe8c52e97a12
z7cade35f389b27eb3059f274d8e9cede8301567b4050e66294fe7b96adb08a218963a4f691b198
z5603c41b0e7fd678bff418e07009b00512e584fdaa6245e5703f1e0d8dbb2ab53c0611a58e2188
z56e9ca17d189505446ae90860c5d87e3406da21fa650cdb77d1d09c42d5d28b57ab14c9b6b739a
z940bb14320a7e6d4c3a82ad6e2c74da95159f95326ce473698ce2b0ea5902880e7ec8dc6f86cb6
zb62b576faa780130d6620ab5f37392c3c3db2e596a40d376de6506be9d759d2e3353df15d66fff
zbf0802babd0c5fee08fdc64bacd6e04092e3537a756f12aa987dcefa7d250270c86a6397757127
zead2833c15b4a74b9b68a646ce63474755455a9a077c4074893cc1c2173d99b5524968b3e15aec
z88cc0afffc48d8afa5ea09d7bccf234175e6625ff0e7535d5713bff440349aa78bd27dcf0e1d8e
z76a908277c5763a691ee96e094cdfbbd54787a4d17e7cb65f72989fe3e6f91440f7fe940451bca
z002becd37c2f3ccc8c389de032b476ceb294006ab7480ab7bfd728a2a0f493fe42555e7d058c9d
z9406d8122e405d2690b6764494fa5e43b111a0589a7cc80a963b93ec13a016c2cdd5edafd9aef3
zb0ab6ad0054c28edb6b2e51642734e1644f962ea6d7995c251c5998af94c1c06ba4fa1bede5568
z187174de6ebff37cbd68220d88912589919a1e5ee335c6d58684fbdfe336f0c6a08eee5b927051
z95c1434ee53988f797b33d6e2814237b3e03aa9ac96431806e96d44b8fba68d8d3f07bdedb1612
ze0923d6c945c1aa9b4484dca8badaca8006ff1fd236abcd6a143abb145a6eba27ce6d1c0fc8add
z5191c3186611bfe089a6361b83717eedc620a604550b9809aaf358aa6f8c2342aaf6e31873e0b8
z9702d1d026862d8634154cffb01c3ad28db22f09b5d7b891bbab58975d41a62e6ab62a8aaeca65
zcc80f5e686d8e12e85353556d0811c48688f99a9c12377465d3739e38a73676ba0528c4d9ae2bb
z2587356a51125a9e0c0c6c5775d06dedb0c4e7b47272d16236d7138a8635d2076d0b3760811a9d
z1a675b71c713560697a96ee9db675dac48c2edb89df6f662183b881039b1d1ff198fb4e4e778ae
z6f998064b2c159ae410193630bc4a9d4f714b34bae9156bee5c0ee1fce22370367a26da3910724
z5a0e5fce146def801c20a3faf004d47645d655c3b72a08ff71af7097e68f6759f1baa8b34b759b
z219c470f29038bf4abf58dc939ce9afebdb46cc5531fb36dad87d04e4a2e84e78a4fba0def40fa
z440b333752d147069e42c7aa32e0d212a4b9edeefc88e78934535456ceb0d1b9d083ceb96fc935
z94053751c779109c23e2ed9b3f8d115ea54bcac0dc996598697e56d0d74a73fb122be15a17dbdf
z9a5c1f1d1d049e60667759380f03adcdb04e942860d27998fc9d2d630457731082cf840935db3f
z176094adabbb8548e453881b2b72fcd69cd7b05e65bac11e64ef4375b045a581fb04623d5793f0
z49e8a17281ebc103eed1f70c15148295a5e8bfd2b7395f8882c8b070ca3f870de1a8dcf171bc69
zf5786881f864b5ff714d8ce881450d141676a7ed1dd4a5c8ddc9ba01ae7a4b7e181f733bf80820
zb3d69370f8847e783b655f7412475fd50c460cde18ed6340b882191e2f46d1b4343c600ce5a6fe
z6c8ecc597b58cedc64560a5c9554b69a52844f2dd6c00f599ab5635928f330141c7a80e820f61b
z3b0d1678a9e658f0bde313ed2163698561756c90541b0a9e2701dc68029e7eab8b76791b3e9409
z13b18ca8d31ef3036abf2170bd138714c7d98f7ff59820b07b49cd40ee0310ca0a7a156c0a8b8c
z7fb326339de066315a9b101efe97a3d00ac23130c3275acdd2239152d39a42229c02e299742c94
zf8a1b232cec772ccbe9aacd9f1d55ab1c0da1560de6714f893b7aadbdc3cbdac465358a7273a20
zcbb5c51b94bd09517747975e152fb7f220bdcb0447abb05a68163b063e22ae0e7151b7cdca4c1c
z8a57bdbca53fee8bc54776b8f3ef0a50c726b83f81dafa96f99eeff364c9f956dc4e224dd216a0
z278efc786da90ffea48d2258d6a6e63ebd90ae8fea5749416a6619ebf2cd9cfdec47c8c955ebd0
z8067734d8d8e90ffcc515e2366bfc02786b7a195f61efe5b81f1d68e27e188d829f8060fce7546
z1990af96897cd545fb0ccd3e03226abd30fa9d8754480fc33d978d8699ec4fec101f56eb1f8d8f
z8a436c3d06da113b9daf59f4227aa5a35ae4468bcc0004e7f6e42115a61c53f53dad4eedd57493
zba634e396fdc10cb8e6d792129443a2128439fb33f68017f398d521599b3cb2d9f6bb39125960f
zf98848836ddde92a5b3725dfa98eac9f564703f11a4f0459ce7fd5f3f2476d620522b6c39b3a49
z3cb29a07144a720c9508f5778c0b03a385f18cacc58ec6a4834c4152bd404f247b2b18a2136dcd
z7516467abc29a005f08c24c83201716c9dbb0c3f100cb52449b9663c8863c2567a9f139345c835
z266f8f6ab2cdeea4cbc9a5f8827ddfd0fea0e59683d835b09c794e48add869bbe6d6730133cf17
z1ea1f887d77559e39222f5892657013aae807201bfd7ec01ef270721201374797ec760e842d080
z37f69dc70343a02da61b5556e772fab2b5f91582549388e288acd1b64f7cbec082d3c136ca5262
z671ddf217d4f08f522990940e44a751690f1fd516e3e6cd829097afe29b10c4870689ca6909bc6
z09b214a595fbe8ffeaac52b840972d210403689daf128eadc39f99bb0b91d22b16ed139ea441b6
zc7a422c3d9d8e5e1e9a9413bd76f19e2406f9ca97ce5055a1b8ef56477f25c4fcd8adba44f6281
zd93738aa6c95b0b8b3aab87520c7f8452739ac432beed1aa47d7c402082a045d18e7edb996319f
zc24e89a4f8267f66c4d30c9c49235fda9e5c696d38f34f1307263e6f7e3621cb73bce5e7f0280e
zad55436060b77af367b718c4bd6388628bd4f54b07b4da7ce4b1e878020997dace43a84996b9be
z8708ae199b41770d9f81de9cab8eb34087597c4409c89e442bbea0b94f20ae63137e38c611da95
z5ad2af3cc9f8223cc9aad239feb2aaf042e84cb4f0a7ce70b107eb771c59d83431f39e5d1eca24
z81347eb786e8429b1c8364e430f1ce798a10dad5c0fc33750299773d7b19ff51bd7242709a8a60
zbaacaf03a0ceee45b2f5560914882a48ae0a3278412231a67bedce8c266bb55973fe18dd081f1d
z217d77d046f221c628ab8be2470e772622b715a635e8b67d12bc332a0a56703342a207e16cd96c
z3c3f8ef849e0590384f17a0bdc4b0cfca67ca394461d75c30f0048cc06a7d8a74025ae69062f6b
zcd091316d77f84359a59121f6f01532354fabde3bf0161b1db2484e10ad93d092d5b4376e6a1ff
zbd9563f1f41851d0dc032127d406ed0474aadc95969c8cea2e13f685da565fe9b30e272361ed10
zffe132b1bc22f4919c62b38ea2c0ec4253a5c9d034c18c8371acc9658a6cc1b59917f9867d289a
z01ee90c210ae11acb406097ed7ec5084fb0afc70b585bbda7e0f7ab525ad86828e5ca52aa84efa
zf9536bf686331e080547420bf50fb0576c839bc6254b2628875096a0333d0b2cd5f3d28cf2f942
z020cc3721189cf337407f605d004999061e26a9ff337b59d34359641ad261c0d91a26179a10e8e
zd269684a103ce408972dc53eb0a637f9b27f5cb058587d01c145d61cc75b6d6f8483366b5c47b0
z7d71604d7b06023f525c95deb279551ab116b51259e0e43cfc24d39415577dbdafc10ea68f43b4
z027ee19578215ec41bd63e7fe4b629e2292fa91083191839cf000db1adaccc00fc412db883796a
z8c48cc511e24aa0de96d000f2cb22da8986b8d179e487de6334aeaea77896437ccdecccacb5639
zbc6ddbcf5a2796fd05dde1ae04a3a7cdb2c157bb15e493b7bc8fc81e2d6d7fa25039ae6efd4b6f
z11e8890610f457ffb67a622ca4f6f471b5520f6f5a3525006f1552c034edaadb677cc5e2fa0648
z40f7f2127916687c682f0bb11791f5ced9fc79ae083b59c52063e1362a0d0709ab15db73723341
z4337994bfa5f16698a3c987da51e626012b420aae81373bba5e393c839f0e9fb8efe226e36dda0
zf5b4420986c4c88a74d2d7a4c1a3c76595f47900be29e6a73ca2cf51cf26196523f805619f2876
z40e3f7cdab546a242a82898fd527f748c2e85999eacbef8609ad4143715c17a1adb603e3e19b4f
z8062d9db88361ba28db8b2ebee4362fe1f495c6decf4d8287830c370f8c859408dd0e54141051c
z6858577c3b11f714f41a5a0a508d1ba532719c5638735dc1561676f843d6bd4237b7886eb29d2e
zd17dfba0e63235df30fd329eb1b2ebd5a0286d79a1021e0075e41a68e399ed7d59dc2f3bc73957
zd00cc5a34efe94be10701c12f329832bcc761f1560e47b3178341879801f2fec46e20145efb54d
z0a179851e46f71ae8598cf2912650481109c2a37f61c5c7e8a7694c6289c71ac727287e4028e37
z600394d6fb95bd1c012c8450b32082301274e2ae78563edd76c7877997e1e97df755cd718d322b
z53e83b114c2f97e12e9eb74f130a41ff195717adc0ca7ef9072e5c4750f84589103633b556a255
zef698935e690ba8f56d9b223bd71c57010b9b9bfbb564806419de28acd7c13010123597676bb48
z4e9f4492412b3b073a317a94b76596e096e7ef6c1100b37a319da4a8952148edd319bc386cebf2
z6305190720554bab3b230391479e98a274462db314adf3431b8a1a78bd65302d89e11f747a3758
zb4a19952c6ec2cfee29a875402a4af310ae3928acc38312e5af7a7d41f373c8287b6ff56b55a13
z10d0b2d38cfac4d23e2db340a1efe2348cc696457452c496321746a0a57347054d95017f1cbb1d
zc45b8d84f1554cbd26fc629c8014789d0f28ec6c4afaf763d92335eb1096969bfbff48f1eb6291
zb9f85dd55d0b9b48aadd8022191942bbcba9132e384637eae6a4bc32de89c0069b92d3f22e6131
za447f79c9dfd56865661baf5678f9fa5a817b3b3b61272ab600457565c059aeebe761757f9ee01
z7f9438a40dfe44bb0d7cd3a24b0d17bb1020cb6c2fd31b58f3951d63fcaeba837a193e9a2a6e02
z678d624de61daf961b1f7bf6570889c59d9b6799e0a2f80b1b898af72bfbf6efa422dee3e1564d
z6b5591696ee5328439cde8d01d3d8f454a963fd955101c79da34a4bea714ce6d244bf52f469aa2
z98c213ebb10373f465c9d460ecc19307a3ded9dd16a5e35333310b0d188dbb27533e06e0177f90
z2d267468da022b34f59ed146b9ecb58ad3126bef06c94de72f13d70d59493323723e88c2376dfc
zce75260c289206a3796e48f4b47efda9a7fe6149b063c9c07c718362d1272d5b30b1564580fdcc
z7c2f172adafd41a3ff1431d1893056c306b6506d8f862dfd9dcb3a69d2c7582c432eb0bc98f597
zaae306cd00d6e9b7b1c6207454e11378f4f17f350fa6a3fbc71a73c56339399b276405fa717f85
z24f3d5c6f998b6f372b94b48024a2fc1d41bba62452ac1819e71afd8d9d802e0c90601e74bb9c3
z1f9bd8bdfc710179a1cb07659cb02fc2583a4fc966ac42b719d3ee5d848b4a576f9bf1a5646981
z6ae56b00e2c4d5666d9e21d9f6e24cd155c09d8008e542099a74f1e234f935aa1fcf5ab6c2efc5
z2dba43c05e9efdd12e15a9459652dcb721808ded90051c5402a0f004ea574f56c704e71c92668d
zac62c71154073fac1594303dd8ac6f3e9ff95703060e7a317c43b501baf2e9dc31de7f26ec742f
z080c9dd223d5392a6fc7161beeaed33710d65a061c4746e64c603972609d4563ce34314df45b79
z2f58f18d93bdc6f4cc0c84afb0764c366fe75be05a339a4247afc1be4f46888e0544b001d66c4e
z680c15829106c8a6171318c96f442a399731a19978ff5dc5e56f37a8805a060b6191c4d522c863
z34e7a3b01d60f94c927a440e9d0e1109fec8184628581eee2aead3494f8977f5a2987118614bd6
zfa31c8bdbfc965258b3446019ddfd4dcd8be68da839dfd2af37f9ddce2b058b9057e9b7e803183
z330497cbf596d924d560e10973c8797127e66958bf9537a37fedb0432409bb61c7bbda1a68d368
z52e4fd9f5b00e28c065c2584dc3b0522bcc46e5f70a639cd50dc4bc20bb0b342ea81093ed488db
z8043e56dd23b4dd8dbfc2a81393c8acd80893837d2bb1bff5e9f6a7eba44860a775dfb5317ed99
zfdd1c12cdcb7634bee56c32201dfb59466d7ccf629cc0c050737ff29c41927a76c9c5fd998f6bb
z0c39fbf7b4190929f1271721f26661401e9dfbfe57fc1accb2266a199bfed46f3236963674dc74
z091733a747c781eed02423978089622ccd76251472970f6db06c08ae25955f59f3a09175858311
zbc016728ed6c5b6c12cf1a0cfb984367c1d30f356f233ceb3484685f864f91616a8be1c8585b95
z0ae612b822d8f68b6ee547126032c3c8b86176d76792a5a08f712ef4e9120cff3f82b445b43a9e
zc129819cbb20b979754b30d55665a8cd28933d1f31f507667ccc14c60b4dc5b5523af4f1ac43b4
z274934758630e52af283230aaa09b148fe1236501ccf7414a07ecc1c8a2826ba9e9785fe66f4c9
z399bb01c26eddae2d7148206f38da0a84db7ee671291ea33e23e883d568161f93d4597bb1bff49
z5e81236967b521683e997ed0641d8b444a0ce23ad496fa3f5e11c7af74ef696ab810aa1e63b065
zad1ad60a14da7f9aff7d898cc58d57b5f19c160d72d89bac6bd71d0077c1f38449e5c2af60d40b
zee92d5ddced48437782e8d203241a8e8697e87b131240ff52414e4928caa5eccc7bca240bea0cb
z21651ba5ef09211515c5affc88243016b03ece4b5e22a764533ebaa2dc7a773058d0d1695ecc69
z46391c2f93a585eb731e5ff8cc39f5f4977733d390e73a5c1c1b3da6ed5d0f01397416bd4d82e6
z3e68fe02a52ba2d8808417fd5080c91613fad310a51cc547cf9a5f1b94c59d7d882c95fe3de18f
z7d86070415a6203a23e687010d007897d74a69dae51b792406a043cf1e8f9fecab3886050969ba
zc681b7d2eb8778173ce261f0936f23d3a6f074de5902f02b66b66ea8e4690d9258d7d3abe58500
zeea0b3fd25ed5b5aa61299c86e925ae8545e46bd23afe1ddf174780edb6eb1c4c04f42dc2854fe
zcb65d275f193fcf6f3df6e5baa7a2d4e7572a74f4ac5673a0351d474732721d707ff3553a32ea5
z039095576e49bb5dbca889992e259cf233f9a33e88caa4db0cc9c6e0baa57bbb41755c6c6d0764
zafbb9773b1cde37b4d009d1e0d58d0c1d86e09ffee313eab2935336fca4dae43fc839c9e60a722
za92bd0f5baa24003cd3293ab73a9df1e6852a94f8e096fea3b5895387f3b1f7def61d5f08bbe24
zf61d4b52196eb37dc9e4dc447f3137b308a873260922ee6e915e8a19644c23cf992f1e431400df
z82d909526b535fb5bbeda5b5b0611d0708a65444b54196e6c3bcf6c4931544308a58610f877f16
zd4f0baae2da4c6a2fcb34927f7e522f609f03c01a4d47aa1f1bd7c979c7ed037aca52913d7cf70
z752420aeacb2fdc0144515ee5b2598d48fce242f40a57d8c927815304ad2893c632f96ac366269
zf7ae948481b29eda444da8004eecebf15dc19a424629d874f0d56e51a831082221163ecb807213
z2c85ee314a251e4382fc4b1eb72e947f68b0fc4c1c1dcd28bafdd4ff3e2c308b0d9bf475c54b1c
zb655345247f22e239429374d66ba480111122c8e8f3b84e90660d8cec65ef7d6dc3fd018e18045
z6b3fcb7550ff83e90ad6970975c69d4589fce3bc258020090609b32d328a788740c6f6df88f638
za7e8ef66e42d027369423bfe4577c4160a9ac7074fc771aac85e08d1caa3e8ca77cbe143a4a737
ze5aaa93d36fd3ca47829f1bd9c1f4d8ff924aa06df5fbecd93145bf1f772ee57692b610186267f
z0f179180fbd03bc09e61b54108d0d63ea266c672fbf0693ee73f349a751c9232034299cf8ca3bd
zb8e7ab0ae53d5ebc02ee89a2ddcff4de27d5a8fbbfb6444edc01700babedbd5a505caf3ffde612
z497d0513804da02e6eb527ac2de84252163826fc5531e645002b6e3b0f7f527cffb9d16aa72607
zaf600c8cc542c75f1ee45692da4cabd54b3a951d7e17214fafeceb708d867fb3ed30ce8a437d1c
z68771e30f365ff9096128f5830c7f679ca5b69923caea3fb030b4db71829286b03f5c6600cb0f9
zc5dc3472bd3ee958bcceccbfc6375a13bd0bd3513ccfb1399fe7c2cb4c98cd8cef81cc3796f45c
zb600e3f1dfa5aa92804c71dafec2a35ae86a811aea0038fd868819209d923dca16a8200dc6f74f
z5bfad97f891058527db48f652bf2616d8ff92d9a59e3cd48126fbd906ec66c77ed7d2bf8267fdd
zdfa208d4ccdf188e8b0649307fc6f7cff0783b55c9129037f19a10ed26f946fd187431af83226d
zc2d15346bfc4451e406376c8be152195616c422a3f1d0b78daab00762637a3bad1342817173502
ze4b9c37ef4a0de624da155ab98693821cc179d34322595ee95ff9d134dc4dfd39309c9b45fdd0a
z2299ab676bb1ab5fd5bd9cdc24774636632d30cab986c8cd0dedc911a4feb4e46a1e1c6082207b
zeede2c80686de05c459e31fa535c59d3c654ef705d5c94d415e6c6f5cdb050a5e54e1e1ea5aee2
zd46528937bb9f8af06e1a42512407c758367942c3b57d9a8ab5277c1ad74674e14bb2e6a539fcc
z56532c10461e67a7c4f20b290af2a58a2db9155915320a8208df34f72af8af7c75db83f6eb4fc6
z8e94873c87a7462c034a8403dad250ef0c25179cd1639bb521e24c95220d80573b38e4b570bd29
zd67cd712f052ea9660cc621e957c1b1022b9a4b9a324718575b429be6af90419c402a186f1b0ea
z5be1d6e694fee6d0e731fb7b07dee163629d1f2ca44d61cc63956fbab875c3e5d4fa77deda9b55
z90d05f53b2d533c63f1c36a6455aac3222faf44ddf993c3e16856f8f231da2631d7fb842396107
z48c91675444e999bfc0b950542c603cfaf6a939ef7050a0b0a97388212643270b5a74412a1f9d9
zaada4657cd85022715fd67ea5dcc393d2d42c22fded04a8ba3920c5de29766efa5212ca52878b4
z0c5b7a37548d204abfe4ed685dedce5f097dbc10c64d9e71c215766ab1647166dfaa6df2cde2ac
z8558d2054445782585f4d29651de95573619fcb4ff9e0b0bf2690662dc430c8edd961fc13e1acf
zfa493cb34a9a28b09ecbf27e27cf4dedb868b805add83943b0be541511a00a4c8d509a11c732a1
z6eea2face4cceb3550638d58bf463d5126d545596e2e06c52430a01ecd50b45e3bbe4b4d3e86cf
zb977d69270c004ca54cc282f374a0ebe829d10f324208057c620f41af6aa5a8a0fe515994d0165
ze153b6778c47ad369105fd77e9cacc3480bd703a19cbcb5087e2ac4f6f0b8008cf0b3e95a132da
zebdadad4a9a4ba50ca9775451814305a41a9757a0a7a069f52eec3263c199075a22879eb80f459
z74f4588c5fd96506d384b5fcc66c9d0d49960cd2acaa7330deeb42b2a4b0d9cfbe822018bc93fd
z3f6d9d6ca75a9630abee14d543e08dc2bcc2f0f4fddd9328d0bbc9fab06e9ba361a4c673a321ed
zd1377a434463eee68d38560f2097ef4e0e9628c007c400aa2445f91dbb203d5687df0389ebc661
zdc056464b5d3a26f8b2dd39aef9450c0787c7bff643d7fb1496d95bb5ee5de446c3f9fa4f1d8ed
z18dd0b28f1c1dd4c4d35593d7f0da6d505072c706de9a497480c0aa28e3a05b1cb78abadf8cdcd
z23f5e5cf00edfb394533437e04cf8a0440e4fd8654c2b316b670449f49b7cc5e7ba1172ee0873d
z526e485e3c465c77b83c2fb09e8fe12ba693404d299dc4c5f5b4ba665b6e806e9c2d0b909a82ab
z9518796a2b4a86f9ca8b0b72f19d89c2d90d13f3400074cf42525b199020e95165869c93362d69
z0948566e002ec0f195e26e2f2aa78c378f75b10ebb5b7419a1efd9abdd8d851e09134a10415369
z70de608ce26d14f0726e5067c904a5186242c8152be660afa40a002272d8b3d483cb87e8fe8d4e
z1eaae25f893d9cbef63fe1bd7441cc4d90df4b52bde6ece40c15f0bb6659d7afc2e8d78868ab98
z2ee177ae7253af4e6c6bc9bcb86671504caedaa66a67ee16eca7565519223fc13f1ede83257acb
zaf6ff96093a360ebb2e17ead2d6b8a207ebddc09e083f93e0ba0e48b9cd8c4760db5a125f59a91
z52ef106ff1e674556cf3dcf0350291d832d32f01733bacbfa314649dd3c36e2a1d617698c42165
z579dba04ba2dbe8d1e2e95304ceece34acff0112912fa2cf39d30dee61fbba3d96860fa1b3a791
zac21b7340a9460cb506449cbc5d99bf681d9e2a4310a171ac4e0bea1a2d79955698ad761c03e68
ze192402e633ebc585a492a07e7edcc21d4fccb2a070b5378af0cc3a67913380aafbde852c3b927
zb4e159934c21112521f96ecf5625cb707b2135a5a643e12f97e3eeaba0db56e27d851c4c3adc90
z12e045f7b0a9ac1ec8aded407fa090eebb513748a7a311e915a41b77e90d9e63bad78f6f34c120
z88fa07b3ba27fe2c9c4a9eedbae7ea25c4fa0333f344a75a142d7717346f2293e34c09ff5134ea
z57b118cf999d13996a4eb28e00f3c40d9595abb309edcddaae2d46b73fdc3850588a7838494322
z2b72b6a0d9d427d8e7251de63a58e748e5ad4f4d9055b804c99352ef1bd96b504049d07b45dfc9
z91229a236e900f507946955879ebf7dc00252a0aa7ce9e3b7bb4d34cbb0ad3539b224f4a7528ec
ze93369ab7766420b92cd84bbca1fb318c98bbba62f06480453d55b68fb021847509aeb56b407c4
z789d36cc2980aa8f0fdb03c4547e3cf2f5f3477c78959a7829c1efcb0f1b38091533933d7ef03d
z13ae59eeafbf604fbc2dee423c0292f3e1a8bde3a354ae9985e0563db1b1e171352efe208d4cef
z31214bb934734e894acf90e0754ce1f65b86f55218f0985b3b283bd7c3909d35d234bb41c4eaa3
zb5bfa1671d36a6515bcc4abd9c0a1f1a5cce9d93d993269bf4019391feb812fd9a215c18c44884
z5ebfa67fe0b5a36bebe5094a2ccec83393460d2a43b2da1007c4e335aa4a5dea2f825d63812f51
zf3cb0476d8ab576b40f78371c4eb65b0acf894330c5f71bfed47d23737b180dd617649c686e076
z4bc2ab0287ecf96e429bf73143a8df5bd61e4c3dfb7c2b5d6db52150ed68a2bc5536b34fd27066
z7ac468ebe62bd598ddc81c8c5485ce7f4757421ec7eec481e45826c3d5afecdcf73f0d909418d6
z056d9a788a4be7c285dd258bb40ddc3e7c6352047bb653dbf1bf9c4d2d8c2ae09b6282a874d5dc
z462960284a7708fd05d0c7deb4fa7e9ba026eeb138960c8bc79dc883fadc4db8012cdb19af5e6c
z0e0d67f2e4f2d94d50acdf023e9313dbbf97e6ac5047230a4f93a36572bfeaa5ed368398bc2bf4
z804e1ca312b12f21b29c86f0e9ab26829f41cad0619ec7c7d5162d2f0828906c021f1aa1d16909
z97b839c93c26276925729cf9a743eea730da8109dc9ef1716ca42278f4dbe6ce10045eacf1227e
z1dcbe0e04e08755f9d3964e1573f203fd94eda7e6c25fbc252a06feab1adf359bd2ea41e67e3c6
z4fcf2734894e4c5df7f379cb6c991f5276abcbbd1a2a9f3d71a8c6b0cf3ad6238da529a08874a9
z604cf6dfd03845f29a61519655457d1658f4555af4c98e6718b8688681526babc8871c3df02c83
z56a1d4baa0c54662e3c2cb2d753d390f78095e080cb2b8cd64287a0a60918f54cb4587a3c9bb0e
zc91ae424fa037076ded81e66c681d57975b3f7be0c931fba0ff2c90860f9820e4e363ec11873e7
z1b469f8e2af18af5e66e46f15fa6a86d20ee60f16769195334a1c9d5928df4ef34fe6324e7a2ee
zd6045fb405400c82f2755d17b17b2bca2bb6806e67bf0db17f5ceade01f1659fa259261bf6c601
z067b3430e45acc8502b9edc4a47e25104b03f8a6bdca0ddfe3d140d147a612f35140e2c8ae8890
z651e14717da368a1034dfcfa33633be24e60bfdff3b5f4a24042e70ef70369138236a6c4c2312e
z61c7c38b30dfafc3febc7c0f2b8e0bb3a7e93c99c42a23e6a410d50b5a7793a08f71e47576fec1
z38b7b2d5013fe233c217d2e462f6603fe16cad8571c56bd3451791b1d32aa7fbba395695ebc039
z8f59fc5bde2222017bdf26541522d05f272ab9b3900dc866b84f832acc9ba5cde758a50e6091ee
zbb19fa14ab2bdba1a45f5d12d925f904de669d876bca0f2f255fa5db31c5d09a2a4f0832a8eba1
z0a851a75bc1b66aed173732d9fbe6ff262ad2b768fa89c547144bf6c6454f16d2bf8042122b5af
z965dd82eb3b144993f520f3ddcba46d24502aa3abcdd666363b1cca4456ca009655e9d9dea9bdb
z50da19979d0f358c5b63a9b641016f3f13a527126240806b708bc10dfcae420f7d2d6dc1e7b7d7
zfe44f72a333cd7fe5dd909fefb4b035d74098664dc9be6afa7e822491f78eacdf3a470026cd86d
zece48b97bdcd7964a531ff71eb1e6f3ee772fe15eff130781ab7386610a3aaf90a76d967b96faf
zd051b153cac155edd9d0ec355fdc0d826cab244c08a61d5b7fca82426a0329768a85e15afcc785
z301ed9b459b0550295977183a51a6ae197f32bb257ddf62b7c79643d92f24b1feadf5e637a834a
za4425c8d1b2bb96aed64a5361370e39f90824cb16b4a28957fb2403ed8f4ebdf37278924e26f14
z02a7b1052f72af61af7e4804ddbc90bedf41d91064c8ef17d186f53355242c4f89aa5374cb1fcf
z8ff914db91983f3c607ba8fa466dc22c7c9ae399c217480916fa87eae2534ca266ca4e74657e40
z93cf2cd30ea4f683174205e85a2d3003a875127da911507b683d82134777dc4e9d9c197f2c3236
z5b80acf7061e2557169b622293f4bd2aaada185dbdb445645e97703afd70731f3f4337796f555d
z72bc6423c59e39dec2b66a62bb5df76a9b70c5854fa1661cae37b854847160643cdf6e144a6665
zf93ffd596813cd65dfd2a60d6f8832397873e084239e3d6018a7e73bd08d655c058e5bf3e39fba
z801fc6ad1a79abaffe58d2dc13affc9cd2b49d34e15507603281c673b4704cc46d7752e58ffff8
z8034390cea05e9ce34190fa233b8872dd4125c1cc8c8603b1c0a189464586448597533a3205caf
z1d7310cf0e1feaa7574ab33f695b52c3b3b7a0f215710477098cef27f5ae47ed77039bd3b5081e
z49bdd2b5110b0e484e44a3ffeb15dfd1bde5e31cce60e8f148f99c7aeb7c0a43aadb1c79fc1705
z045323c178441c2063347e4a75afb6dc9e7812e28a437cb8ae7e11a15fa15a6c0f9a2b7ebc1315
z2e80012cb647a86b3cc65e4aeab7df2be74d334f1a0db9c17ff7c466b0e11b20f155f687b14340
z255ff2cdd42ab26ddddb23880817ef8feffed2a8fe164858b0f520617939217a252bc12fcc1e42
z30abd65becf4b0421f86e9d8a5404a0af8feecec053e1e84137ef158a55304d86d0f71c55130ab
za3985ec7dc04075ce49eb77c64ec89fbfca1132c732c35f8abd5328dae55c26d6c2d0453974bac
z42fbafd4abdc3ccebf1c71512c22fde69bdf351e442a51a538617b400f532f41a424356b28e8fc
za5379caf4aaf897aac9ad7cfdf72883285a846b940fface05c0d402da3c81bee71daca284b0218
zc7471587b4aa6412245c441a839887c0c10d5f55bec8c16b40267c4653e3995ee7847b4d5b04ef
z8c31c1b8b5604a26225822eb099f1786d0ed2fdb8f56b07d92430e1f8f724a6a8117ebce4b8145
zb15cc2699b53dcf4d9f264927ec79bb77dba012c72cfe7214fcd61c46be86566d0ebb789e37247
zfe09cee966edd030540f0ce002b3d33653dbeeb0ac457ffcb3bcf6cc86105b65b1261235ff1403
z52de250bc490f46d05f66b92c8c021b32126e640f2a0771b65c54441d52e45594414319ae3b563
zf015b83c508c6aa95507a1c6148890d94f0d3e27f5519e07551d8595de09edb21f9493f75bc238
z26652cae52b5b4dc3dbb6a59c3c251c736412e18ae2f8a3df5f1ae205f7eba0945515438c6ff6f
z6b4daa90b0a2eb4307529e8c4a033ab0a6cc76eeffb9f6d03a777a4dd63bb69e99ddba76cfde8e
z841b271484724c5a11ae8b7b51bd1967a8291bbda1edcf8c6f2631fafe634022fbad49b1dbeabe
z2fe70634a7a41c4fed92e6b4543c8170df50be4fbfbb8bcca767e212b4fba9c8a6accd60cd0608
z5611104de9a205353e603bafb5f974a3b834c65210b10760be3b8fe2530ceaff437cd3645ad6c3
z18e4abea69514ff72f263b40e81440546b778c96cb91b7010d09721fd1e11a92607b039230ca84
z0da7c6406c718fdcfad5d28e4d831d4d5d4503d10168d3da39e0bb1a9cbf85ff5c4fcfd9ad9303
z7f522126587d8b008e4252a4f7e662d175d7358dd460803e5bd099677e6605be62f8beb626685c
z44956522670e3fb0919cd95f12f9c653c5f78766a5c362a4016ebbbd13f889c6f77aad80006c4c
z8eeb435f76b4eba246ad040d64c4ca18e1316182327eef89d535006cef88cb96ab57b389db3401
z959b90cd0494693721485b22b8230aab90e8578a728e8c16814774ee077c99dddb4e266205032b
z5f0c75d701e9efff1e3e83ea104858b386770e4a29a841c34bf5c54150584221b0e051b82f331f
z77c38371ffd637f616be41b440d849810822c6fe3f34873526243e79fc496661c1834efd8205e7
z57aa70746030dcb4cf3f1895160ac53e547153f7c489471b4ed372b618a757c221ffaabbe61318
z7e942a112364addeb705f5e234c7527ce71e0efadd09698b0bd416b263ebd507a1d94c1745e034
zefa2739dddbe424408f9ecb631f3934af1c0a933d62b9914bc7a0eea662aeeee693d24e043b8a7
z387ffe87f21599908f6d12b159a6bb6860964eac92626b1bda5e5d729f2869337527e58e80c8cf
z6742f47fac3992cbbb9a56ed79214ad0cbad300fbf9a8e491806f3996d7f9d0bb5c84e87c265eb
z182192981b649346662a2da16a141919615407ffeda9b3a6cc17e7c73a10480df0c8789e92ec11
zc791c0a267a947c03067903804c79cced303c4c2535b74b84f42237c228f4b8edfe6b621297c44
z59acfb38247787868dd4742933872be9afcbfab6dbea4ea203cc94b50ad2b634e27c385461e7a5
ze8f8e6287942801939502bc19ae59e71418fa1c0cbddba6f427267ac800e842b15f4db3bd29319
z65c83f6039626b18d903dd843202f31f8c36b95fd41c600c2784a2275f1388a74997737a828d49
z3b4644e778b4fd33e0dbfeb53bd0aeda1f1ef9c19fea0fd2ef9c1dedfd8711c404801fdaa077b6
z0378989534de04f50de40ac9d298bc14d0e5b1fb33fca0dfcea995a8339450929f727fcca1e733
z911571ea573f7418688495b850131dd6b07e339245fa230bb168ab55c10e1336a089c37a067be7
zd50fbed267e4982bd508f6fb3a16529f2b04d47b02810fed35982628d10ae686f016798eee2f1c
z94d38b7a3e0624ff4074db43a4b6cc7a76f8e6930fda3d70834009188e3a9c0b0dad03afa14cbe
zda3c0cc3be4ae5f3c127aa4c45737bf55d38708d11ec374a4819822c29e878343e891e51045ce8
z5d826cfc80b76ddb4916b109cb90b3a7a8129183e18a42709f8dae54535d81e2d95527cbd3e733
z06d80bb977e3bead608461d4950805d21b5b63f693ff0c467f87a813a4f4e5c8aa771cea3420ff
zcbe8403ecefaf2d48ca61e597c71d2dd77dd517e611cfd979455cec474d7d1256249b2c54506c7
z8fe0c16de7fbb5a29c50cccfe7b282554f24c3848981a81ce39a9104a965494d2f3ad615b2df3e
zca4dbd73cf6a2d86845fd8d071ab96d161c73fe3212a787ffa3e0351f3a7ecf066879b738b960f
zd59b8370ae1a8e969a83d8674e518a2f8d9b2ddd4213ce51de3646685684d0be167a0fb207e868
ze713c1c580808959501e5d50eadb0dd5a07f6c17ea5865cf42fae9e5551b329ba58e4cc439b609
zeef9eed6399aea1f27bf806ecd3859f972c4f4b9c0da54247dc8689aee62dea1cf265c25d9b116
z9d2eb97308a1331fb2ff447c45ea4688a233bd149eccae59d7fbe1cb1407d4127167e2c157efe8
zf8bd3620d31cf08183ae72544071b3a55a8300204644d94731c53a5e274b5becc053fd7ebea9e0
za0e55bba7cb971a9c1eca1241adc7760a1d77f0733d2bc9f84463f7d3347ed40899b8181aca0eb
z4d401637c32243e1bb70497203f3f95755c9ad2a8852a194a0e765791787131a94cd25e21e00c9
zf7ed9701c5f0c6108331696ca63806daf3deccce30ae67af7937ea7b3d5593b1cfc974e0dc852d
z33800c47594e5bfbcc68aeb5ec1064ee402e1d7a64cb64df9766c2bcdd72bbf5f99b03a9bfa1dd
z0740e9dd300e8cf64c2f7325621fdfd589b3d87f3ccfecc6ff6bd6ca60a1595576510bacd3fb61
z8b075e400872bd7df61602d2223febb525b9ddd636a2532129f4ec58882f9bd7afe10661ac1efe
z5ddf8c25f2b4f0f8a18f7aaf26537c087238161bfd7fdbe118869bd2e1e853d1e83c845dafdbd2
z55f74485af0d589db142ab7154bc42cfaf0cbbbb9be76710ce8de9980899ec901cf4a8fe693bde
zc8e1e6193520c7bf3ae40cd676c5a8850d261d3dde5c5288bdc3c661c52139b18972eee58fc979
z7d57276bde0c38d791d90eedb2e470d79f546c220786fa1b1baec634578262b38a1622d3d027da
z2f7e4968cfc5fc083cc3a93716acfcbba4206b3bd78389d41d48eb5332294baac7b35f7387a676
z20eedee5db69bcb46717443499a13f3796ef9378e8afcbda57dd603f0b55f217e9a7b8eee0e27b
z9bd724339144ce061471b13dcc343893cf5c30fd8a54003c3c08899aff63e3599b547b8b3f0c74
z798ff07a8daa2687fa5f3c1aafbe274e425712d3e99a89fcdcc17b81701bd3672fb02b52add333
z37eaf78b3782f5840218bcb23333febc381a96318cf37263425b9e15624c917b2280bc4e82ef8a
z39b31276523fd17f239222a07d6fa665be847e42d6407dda62a3dbd3de4432d57b7e67b5a12038
zc3cb29c0c82b7bd8d4a2eb09ed9bc56596c222679365102824e0db5e3be90b104314bcc4e79107
z66bf6dd240b3321a0ac244a131e63a2f3b70bb25ec244c04d2ab09478df63e55b8539894ad15e4
ze7eb833ccfd42225015672349cf8d921c0ad22290a40b466b2fec624830d1da3e08eb4bb570202
z2f495bb1cdce5b73b74446f41b5945cf95d2eb1786e4c41d1706e729627f891a3bd7c5a3acb763
z5c4fb01cf71b21b48dd151af2d70661f4e9e7bf1a1cf440b190428defb616f03cdaae9c9f388b9
z6f6e9f3ceac2c2a3118b12087a0f88163d419e37697da037c5bf7e796e19c1056a97c40aceed12
zdde4a928ff5e36e026c192de73a9afcfdc0dfadcfc3dddc3c055b441b819ebe3fbc54f0c51ca93
zfcf6a1b78ae6ae388f62cca430b576ae9d2b66ae766feee3f93657cd4fdf28989e9c7b273d248a
z32ee7ca57198ef981c105fd528b0b0d30ab8dd2932033cd5b5bd5fb92b03e5a0bf68301e4754ab
zc1022e7f5aea28b09e2d309b2da491451c1429192bc66a7a71641b167de8a1db54c85dadfc90cf
zb3b781553e48fceda1c5ac0768deec972a30af638b97ce691bb1d95dde5fe1d6f659c6f58162dd
z30e7cc7050ecce53a1792fdd80b613928b4aa44c89e2ce7abba8f7831d6667052c9d3dc60978a1
z96ead25da8c7653c9c3321a10daccbc3a65dc626356564c0c0ab0903a80c5c2c817f3a4abb5fdf
z380eacc81954a440e649ff12fa8791b9a20fc0e38d5c62f04675ea90c972a18cafa20bb1746d80
z4a11e850d61620282d39226054e88ccf7436c878b9bb9a103998f0ef6095448c484a7a7b07a90e
ze6a8fa0f7b3695a61a230e95b2870cdbe4318b1be2e42c5303eaf0e00e8d3811708965abc0ff34
zbe14d55bfa5a00da654cbfdf51de421368cc1a0ea7762b76184786d0c76315168e14cd8676b7a1
z83de9e894da48368a669780c7b371d013ca6120c263a1ce68c5f997fd72496146b4c9837415013
z53aa060e59c1b7843ff95a84b98ac86da49257068350d0fcb8107e45c4d2d7903c109ee28ba7ec
za07deb69aede9b16812581e538fbb8234d01e9b372ef72d0a712168e4733e0b9d7ed226be5ebe8
zb4235e82e05cbf4d86bb0a3b8c86449680f0d2807f5eb422baa8a2415297274afa353aa4684f05
z4fa5efbc7390dd673ff914bd3dec4ae62ebc0277de90166885f2e07cf807c6f3cddd714418bd58
z8f4caca8a4669df472e86e5428ea158e02d7281220199b99fcf1217d1c58eb5f369dc8dbba5362
z75685060e1b48037f378d35f000a11dbc857e4f5d685b5d2a5a01765a08195fcc46116700d1680
z9b7b26f70b3541ba6fc96b497e7f1674c13450501d10585e749bd743440091be4d2a503cdfd2ea
z2bb898e6b92a400891603b026da5b28036cdfed87ca1832c462267927538df32e6e4a427f07f6c
z21aae7c2657039c1254eeab9a6156bb41948c19ea0bc062ca9c6dae418629978335c32cd2c2499
z462a45ad2f5f52b41d6abe402ed17ce9284252ee6f97072915fa33dd00523abe7b3307b0cb0510
z4f376a40b49c497ff7c024316116d2713a83065557e06bd1d23ba2c02d37f4ae184dacf634eb46
z0801e5ab449e7440cc830d71096f730874e013864a9bd62e43c066ea864c00679bc9e2bfda7b54
z7c4ca22ef7e14fcd4e915bbe7ac23e5c7228f75cc0bb0a5103d054295522479c029e224a191d82
zfbaf5599eb146990f938948d86ab09da45b25fbd8bb03d53cbce32c17bc2962548392e8d27bb73
z1620ff591f61a3cf73ff2bc6380fa89ca612d0cb68ce9b8ec37ee5bced067b0d51dc88daeb5cef
z78eba8e7a708ae2cb6be8a13643f257581aadbcdc7e97291e26de87bc5811ad286567df1c4af52
ze9df8f08339341e1392c52a3bf5501348a50c922eb1274a547afc0177062e6da258ed0ecb0a4e0
z50cff4f08ec283e95179775b327ecca2e6e9b47b2a168c887fe7e2b5a6f14897af490d79d49d8d
zdae48250cad928545ccda06ab9a638efa5f64aa16ef6708842b812a66379c945ece01db2b18898
zc369fb482a51d8f3f216cbb817efe8d221bcdcf2a3e9e728039c6bea008f958213ff5259b5909e
z9dcf0a527fddcbe91a08fa75cefcf808cc68de9d70f1c1525368e4347b9d140816c2880f09dea0
z0173a849b91ae2f35703cf3ccb2c5e35541f79cefd3ee256525cea17cf212b4ee9cb2f3ef8b13f
z33a7b5f1d6741f673f6c6aff883b60bb7c419a18ba4af37659193e6d14555e7fa522ee463aa342
z607280458ae543f40d10093f13803e2ab321088a78adab1ad9af290ecea4588fa87994e77d2c0f
z9e9a219d3a212578ce5f896eb3d11681caf4db4baca70f5f02a96bce195aec86689a16902cbd6b
zafafd4671d089939b01c79214fe38c2d9cb845bcaff10084b99b2112a46cde844546ae6facc522
z201bd3bfac9da1556150421e7c078ab7e118bc1e35925fb29d7b97e8df90c317adfdb8cd6f45ae
z2b87bf9b78fc2af4d04d8efcaf46aa4cf002281e15c1d09e97bf0d977717a18e6a83f38757537e
zd292bdca19aeb27f7eb73c8238845c8f842b34598d004a40deb530825c2a0104640c703c9cbe14
z89160fbfe5d49b29a7146aa67b13d7773c49d56b4310893959207d2ed57116f8f6ad279fe1bee1
z1340617205ac432f7a8c2b4927cb33ab0cceccc17bd23de7a1ae4be922cfc0fd74ee270956fb8b
z3d04d4db624e212a24fe94925f49ac064ceffbc07148db5dd1013743a12511cb4606e99df39fdc
z860bdb47c31a131dff0edbfb4e54ca4a5e3166160f3dba1c5a3036de6127d3274c395ac232cd42
z52b148d61c95604599e627052ba5983fabf49728170f207bdcbc5692214844e6dc59e17ce51f51
z76039e5c28e4f6fc24ad7e95626ad3c72f41c1f90828ec5174b89583fc0e4d90bf6196ef151cf7
z7affaac511f08e2175c6ad1df701fda929549df16175002ee62acef3303a9490a762360c0580e9
zc9361b55fa56719ec8637a87654c017b304e61178b36b73adda8a9ef48fda915d973b308d7c832
zc7cc49b144485c353ebcdddca5f7fc5829c72dc316468511a7b83675cbcd448b51bb42c85bea42
z46bb7ff61d1e1832c0bc1514049194ec056df7be4221fbe26753346099c0927f4c847d0e2d4dca
zefbfc9d56abf24fe1ed785625538e1bc0e5fa5d5b58ffe26a1e4c6f034c02dae6b6f8f56aea9ce
z7d94a0c00a930fc447b1da38f9d85fdc75ff04859d3728ae04793f73f46afc5e47705661a1591a
z7f44f35d7606a741822176e2da4d96d66678eeae6a1fa9f9dc39f8b4818f081ffca7548da588e9
z6845812ea08a8a1eed93aaa23b5abf43b22b3fb81cd821fcedfcbe14f2c5400f14655b2b0dc949
z756855706d4827d77732254d24710cd04fad244f4bd7907b644ed4f88c99dc675399246038311d
z0837dff0cd097e087f1c7d6ca00a9e75cff21697fcf615f760116931c478d8e24444a06cc283b3
z378db0f8b79a63f7f48351c19842404de1f4cdfb59e25d23097917acb31b60f82cbf2f5ff92f38
zd10f5509e151ee735cdd4b9434cb568a3a9fe2d533ea596ca03c0cd0ed791e172e4c1c08e35078
zefa7f2c227145ba27eb2c34467f38828bfc5a2ca791693341f90a2680447752a2e989500f72d04
z3b3383a5baab523b4a7c7cb4357b729cc9135cde67c0bd7a1bbc5f26097025d989c8f718db117d
z3fc7758592d4c57d9c50067ec62c3a8a4f6f3424b85a6addbcca1a762a7685ea004ff9b947d06c
zfbbbba63104d186b9b7751735a6ecc0ccec9c7d15b06e5a1a3d3cdb69bcfe0da388a93c4dd764c
zb035f4467fc4b2bf9d879c4497a8d1158e62b235f419cfaeac712328a3e34bd1bf682337a6b38b
z264121a6454c639df41bf22bbd0bc358a3990f5b11abfe97040ec23cc7b4116d66d8dcdeb19c4c
z3e7fe0a7c5b2e006d5aaa4e0f6947a6842e08dbe96a5dd57c1c337ef1a32eaef5b04bd0f167f40
zb0fa372e2914d7a395ccddaaa9a849d5a395ad8ed660f015807c6084f25b3493502bfccce2c61f
z0fb7571cc962ca93cf119b7896fd2c589d712adebad4eaf86f525c1051f98da7241d72b17038eb
z91e7eb8d00b77ad4001a2a077b98f302b8eb1b1783ed2874924d6a43f812560b8d844aea481040
z98f56f602dec0cf06cd2ce8edfdc66f72ea276b2d01f9f29a25c9e43534d8dd072d397e8e11048
z957ffc397b20ddc744ef110638e0832cda3ddae2510ed6c324a921acf27a925e4df4ff6c967a21
z2f92bba9293981ffc73bc4805d0932023925d39c93682c45be9b2a34ab10b3ab7a0ee7330e4f58
z36fa339dc01041c7b2f9724c97050c312bdc66dafe02fb86a11d811a99ebaf4a556a98d79d3882
zafa39ea814c92419498aadb75a2ee5dd404e86ecd6520fb42ad2e1248cc2c9ec44d377fa2ce3ef
z5d02e3b2076fcff18e17fac67cb77dfcc6f5fbe97203015499672078787d5d7ca6a689ccd5224e
zcc3114fb2a6b20f62926fceb2f4fd1eb474bb8be08577933130a15a83949ad80e35cc997adb373
z73bb39bb3daca8db42294b8e371a75837cf8c2e0fbe65e2962f3fa73bc309a662bde47ba13ffca
z0eec4086f84bf46d0427aaa8a429a67bf71e21530efeeba18948cc2fa382e6e11f7bd3caf8b11f
zad19787bad96b611ad5d845e57c2a7bb5640d25cc2b80dce512dfb1128625a2c8840c5fef9b34e
z546f78454e137d8a69a5e2cc5f08ef10ddd77010cf528253a59ac8f2a849377375b07ceb1d93ba
zbad7f9c047b8acdd507ffc05bdd8eb44f54123b153f867712ac935005cd5b98787bc44ef8e439f
z0a607787130c0331f9c601878009ea886ffcee278d02bf2fef49bd69d25281f5ba25f130026aff
z646a3f4f481223e945fb0868d53d4285d59e3b091691f056ebd80cba18f366149cc6cfa1f2c507
z3834633513db9c2f7af884ee94e6c8001951fe30ff595f7777717f9b0a7cc56e037711d1733d8d
z541b2f90cd6b628733c5d4b24bb0b427e588de150a85f11e81e47e36faae5f193987e5b8455b40
z9a901ad0cded5a386cd2c88223e4135135173298496bec5fc41f03bbaa08fd7d6e976512e57e27
z9b4eba17f819998ccac360334b39f0f7b239fc3e0e2950707475ab9c1772029fc32366514b88cd
z2987d6f0f4f7cf00cd9419a3c95fbf15a37265517d281822e3e59cef24813c1855f81190482a13
z45de31ee49e02520253027b6eb1eb468fd5da31a1a37904f4fffbc61e118d628c4510d3aaf00df
z1eedc67d4c8e822f3e622e22c9bfc089225b168539e462a96bbcbbfbcf0e1515f551798d758536
z59d66adf34b645e81e61a9bc45b04119f4571d0d0b44170f6a837b254cd76e5a24f1563916cea7
z8989e14d42bc784de1b082e911c7605368fed0a772fdbdb734ccb67b11b7f936e0c2bb8f27d042
z95b57d11ffbaba58533cf8a66eb3e77ac301bdf75bb75a4c0c92780101a300584f4bb1106bd283
z32c7699807002d18798817a2f050c941a663ce0698fb73a30a2ce7050c545979f5ab52909c3c43
zfef9062fcd000ad5c66b39b877a9311e3d0382b328d0d9b7963e03276738dfcda91b0bfb22f515
z3d973aabdeb45108ec2d70742c7dc1fdf7924fb4462761a2800d0f2e9d4de0de6ff2fbb1b043ed
zbb502a7d45a0cd6f67bef83aeac27f4c2def14a7aec838b0970ccb8ae1275120c4b7c3aec27952
z591165e63435499752397c29eaa718c054084cc3cb48e1a7be492f523b61f8ddb52bfeff92eef0
z652dd21954db61356c4df2516f68067ec4ed1475492663a0a647dd8e6bff6f13ab52587b69b9ab
zdf9cc3360cb38ae21478f6a01b4c830507dd1898ed889417b78874c06fb0d7b17051f0c277bf72
z7056106c8137518a0a4b6b8187771395c5d44f115699f3034bda2b941ea7c067524ba01afb05a7
z78915b3c70c5b7d9a9c713f235b4ff5f82825fb22b64ca32337ef47f9f4fd2865fa12ac4c79326
z0e08c3933f575acaa3225166685249adacd053b075e3fede2cf3a39a3059ad36b429e82895eaa0
z6e67b36100e6ee859faa78057c1c593c46a1b77f0d0e462829a251717561272a925bc0a7d6653a
z97af410bf8b0db1d5bfc6a233781d32b3a2a3464e1d2a056e6c6362258b9250f1a74dceb1e6759
z9387f655a23cb22a038bc7c79b3e276870e26b17b36b8d7a6a2645d6bcb2557556098e2038675f
z62e42198f8fac1ae7ab5ef9619e8145f1e562d71eb43d7a410d895156b138ebe4c22f889789f59
z024576ed05193b642a3fcaacb6a3e70e7910d3a8ca187d573f65042994317eb27070e1c78faf54
zf13e8437f7f5026b7af9a743524d53e2aa033d0f7be932c500006b66b26e57a30c48baccc7cfe6
z1d1c0cab71a364af0a23b392e74be8993e85afe703068d420bef0fa24ecc5e67894490871817e6
z769845ed1ec1189517e0dbd3787bdcfb39e02ab6d882192fabdb08afa92c354bd3765ba99d2ca6
z3183372803f14555dfdfd1d53f456524953a14a8b5a94064421565b9c9d80e1b79ca6c3b30f14d
z9d879b3b7d6b582e659998bee3965c12d0b6dbc537cf4fd938588e318f366ff603f70f23a33841
z35ce571cdcd8584f28cc9b998c753befe5b2002d91501d801bac19e2df7d93fc2a526809c84bdf
z3722f50a49793e1ad3c52ef8fc7689452c20db6db7706829f57f44427552691d71695770adbf49
zd65010a11ac8a930d5e7751e97891a7223064720a2f46266ec4ec3a9f4d0319ac0eb4baeab82e1
z38ae70fdc563c9866704dc972d991c84d077eff2115210fde94e0c34bfcc6dd7b0d4652c7d649d
z24f3e238097e0b69566c8afccb771eb1d177033663a1adfa71d5d8cbdc768027bb604642162dc6
z8e7b0717940f4d74b49053bfe0b17ffe26a7e34cf7277b3db04904f46d516d55c132f07ce4b44e
z7b4e0045a737b1572df7bb2367fc583422df9da5b7472de35abeab84e41b91c6f7a6c598556331
z1d2f6d0afeaa919fa01c011a2c88ad00a6b1eb2046bfd8a44c2b1324a8f3fd00680957365cc6b0
z461ea943786840e85392eb0c677b209b40cc0e0d0b033ea9b8454b552a4f151f241d1692b49fca
z6975ac9aa8d0e894c925b5d9f687ca125e4382f4459aaa2d7de42193a8cfb25b941b5cab2351de
z498d3664e6c0391244dbe7fab4d1d64cbbfcfce95797772bd753fa78f6f693c8c17be091936e3e
z19504d9fa8bc8330789e296f6ec1bd6f1f36c69d4a5904c3c5632f9de4e8bf66c117f46362eb85
z6d0cff5f59538fd72904259c65538fc135e3854d083a4cf50958dfbd5dadb071cfe585f6c245b8
z896f4c876a1354898815791b3d2d41c77903d57a1d2a1d0a6cdd326e2e57aa36a62bbe3b1f18fb
z8de1bccda54f5b29bc6d073ec671f7a182435c70b8945679a7941dd7d6f8cf9432a6469223e7e0
z400258c8e6ce3db574ffe3a334f57592c3cfe54f46cefd9179da2a5bdbd4b8b9a791d53a4f5e4d
zd8ef45ea1c0159054aa34f6755946c9671b52998a671ffa923384462bfdc8eb549b005f901cedf
zba26d977806bc5a032793ab44f3743537908a6eec96b7591ba496e7427f154855604d5eb4e8e8b
ze8e1462ea4748d7150a38841695f7b688b221f75a1f48a8793d8ab3761587eae768205dd9f8fbc
z5c69b6367930a071644354d0b3d3eed8ac75c57aa3bb108c210cd8d4435223899d5cf962dd514a
z29e9dd3817baaa00a20a3eb7d494502960d5a6fa1a603ebe1a978fc93eac82a155c2ae98797c29
z2fc91689d2a35f47a04323cdd8823c8e1c4b8011f1c08236ed631e43cfcae3e4558b423832b56c
zb079584304df21b45cafab672ad368c6f69547970bdb4d69efa2f8cfe7f7eacbf8017cde24ddd5
z14095e18e2e2f71402192e549e10cc9587b02a81604a6bce0ac5134cb40719a9f5a47806078e17
z4e2075b2c9860ea24047bb1c6e53bf027b7e94724584155faa7063a1840029826a02cbd3900669
z07a2e6b6087e6fab4d5d211b971df7af87f05b9033b97f5821f7e9e278a8daae82b56bb399299d
zd832e8d2afaceb51fdb1174bc16d464ce2e1d99dab9feb27175591dc5e4aa29f41f43ec7df9402
z0cda4d4dcd05650d7935e9f14ac94c4ae1105e2cb64969c1e8301f0d16ce003064dbd70339df7e
z24445641bf66312880e9005c702a3df95706c515e75a22c08e1103104b43dc8c729e82d346376e
z0004b4dc4e3c5ca68ff63e3a7c8de20832928b94269a3862353f87f900cf71225b8ce52d78be4d
z7a4ceaf0c1eab0e536e515ecf75cdc8a8aeaafff59292a10183a3e8346b1e7f7844dc6c5db6f39
z18239cb201ddc5a1e57cbe1d7f5ddd9949c9cf3d6f2532b8078794f37bd5e53ad1a81797df8313
z799c5ea13a89008417acd62b6a8e9ccf84b29b1e0e056a4fcce1871c6ac9d2414e380c3e7b30bd
z77a0d03a446dc0577b384b9c8dd486755943c7ebcb0bc14f40b17b4d1f9de884680a465f486b6c
z70f7e93be12db4f1049ed73f105831b2f89708b9fd35c7b75545c8535046c9cb67b9d317850824
z27218c5e741d01ccd9b586bdeefa293cffdd3a2c315c25e6b3b8c96cbf6f09ee63425c0ebf293c
zf4eb2e13d657bc8a4bb44c696b95f940bcd1a608a1c6583e7542b2531726b4e75edcc87c700ffb
z6408907e25d74226f963be72ac5047e5ee315677b65d478e0457139e7b5ed4fcd53fdf4d214f55
z9580ea549f772c5c06b9be9d596c3ade5ef72051a4142ef2c02afaa48eba1c86e677fefa56f61f
z6a5f8fa2cf861f1d3f6045a4b324e88ba0ccba07bba676a0fb0bbe94f3c38782b96670e13bf7ad
z52410dfa87f93d3d01dc249139bc17570b7c6c2221a26f5638c05499375fac94f6c46b0436447f
zd585847b3dafac299a42aaf1cc0596e7fcf1314d5c74240a8f5ebb918a1d263d3cc8d0502568b8
za29be858606fdee51b5198117d1ff5926719cf8854063c6f32db50ad0e957ca7bf5f9db97bd835
z77ebb841cd2b7188e6b66ee046d8616f93cca90a922404b245a5e5770b406242080734f1d2a898
z4999891e9718030d0297e7824e17c0510a8c250afe4d1f3fb3f8ee5edac1cab027e83a7ece3094
zc521373612c13a17ad13aa6aec65c7dbd3e21005fc5e9483a57ca2f460208f0b6a6330552a7196
z22112792b5e83a3eca75d34fcfe5d764c81016d97fe50afe39b928d8e0d8f0a2121574d121ea85
z86a1c33b18d96b4e037e6cf966adc022bc053b8a9ce3628bb49833449e80c018c5f73ddb291fc6
zc7655c36679fc106ad80a7d411b8276f07753a0eee89d02417e49718cce43d28c86660dd322030
z34010c7983d9c73894dd087452ed8d2774d4e4b553c2c683073516ee05426a531d4749710de816
z81a3ac25c86f02922799a5db2743556eb723cadc2dcdfcd70fb212d75d3c8916bf688c7370fd13
zcc1859d0d732aed5d404d05576c66018a872aa3a1f35571df327d62f474d3cba878339d1e6aef6
z81701a3ff0fb692714b01b2654591974a03bf74977d10353b3eb268f05495f97227727a2ab686a
zbea3eec0ea177ba74e4fb1f8cba06025b6af2499584355ce08311021f4d203156f34a05ace84c4
zccb48ea7e5e391f49ca469d7e9595ac401fb56f9f8d44f59fbd58def46301584eee97997360558
zaa2e860b5e13976ca5fc9dea973abf930ebdc5ebf3e3b95da5898f4cf86f1516cccacb53c8a110
z77aec8d7a4db86fcd0b2e9a2a9a087d44c1d8c95b21fdb9b7cf47d0b709d8e1678feded4bd0376
z131e3b07c64a77e510b18f2322468ede136669e47a4e19ad3a53181158bf0ac696bf92653a50bf
z0bf763596f28661056e3e8fa74010628d8c91c183f80fcf5e73d89e8389cb7a0dcfa6a01b40539
z21d7c931de7625e4381b3f60d2893a043ecc61cbcb222b6e7de26ab668858d0537850d14741af3
z9a25f3ebf38ba09c2d75eb2deb993080f0c5dff01b80e26ab397fa12d012aeeb5f152dbc626b34
z16eaa2fe2200d554c1300edeec9737f6dd8d0926fc11be770cf797f0e8f1a60455c6b8bc721dc9
z4dd716004a417a879962b5fc936bc76646a61d38f507fbfbdae06ccff3b56b8c41127e8fc7941c
za95ca77a7803b6481fdcbd76786421d54b9456525d429d130123bdcc7b7f78426a02783c7284ef
z4bd0dd8c42cc79149c255412fd8d679314586a786328e05042e810d4c484b67039ab4c437c22df
zb217710541045120253e3193693caf962c33fa92da6fc1ba7a853dbf272483ee83b50f7afa9ee8
ze39d4924735ba943a4103c6c27221a517d55d6b7bceca0770a11b6db4da6403b3fc4ca3f2cc467
z40cb470588e3cd9752f02d99e35fa9bdd6afba34163b0514723e63d8f0ee995e0d77ce2ae86813
z68bab2706f7dbf70f1f69f9d713644356eaae1dbf6fed23ce3569f713e06a3660d13a7e1e1c747
zc5143215d67bdf437734f13b87588d1565dbc8118d6b49ef61d25c5356a91cec563e0da50c6f6e
z73fc378e71081c697bc05c927bddf91c4442ad5c993f2bba07c689a7d978b9a5aef428838b12cf
z551f1fe66c8fb68b689913a8038bde8a82db43925b008a2d7a808ad8ec0f6cb526e0e6219b5a0f
ze51ebf49e99492610b1d92fa1e7c8f2bd9b1fe48f218a975c91be71818df8ae4de48cea49e4e44
z6e870018888e6487e7cd7e95cc6feadb492f16e443f4e417dcd96398c3569757fa7b773ea8c4b8
z062b405780209880aec3febe2e636c49eafaaac954bc1b52482e1b71bb3f91e757d44dc81e6c9c
z20c8bdf4f21bb1bc5c2c56595151d2320ac69531a9ee3379d42c07b0b5c231ab9b78854addf45c
z5a3fe226beba877fbeb771d91993b76538c452fc780f4c637a0c462e5132a4b94180413fa4a2d8
z7802f2523225f5758099c8b7082435303358e74d21305a7370498318baa089e17efa2a3d759cc2
z141eacedb119b934f070d58c6946c6529ceebfc5854a8d0c03467012bd7068cf1b7c976934b0ae
zb8a55ab34faf9693e3daa9e17a2472cf17fe903f63a9a5ea181dad7f67bd0697361f6948b4ab87
z30a0ddc43873aaeda2d9da208da44c3934a6bc10f4e0b728971b287b03ed559a110279de0988d3
ze29d8bd6ef8acff8a8d6c0ebc760458154984d69e8bf525c0b7e1b863113132155edcef1f7fe9d
z55423328d5c751e11b48519754e5f6c9e3927f1574c537414b7338f0de36f6c717b949f3c20741
z33c8c9076fa608accf69050da8ca682a838e367177cc5baa4cd174df8ac9ad77dc22f0cf27af1a
zeebb50203d2d1174bf47552b8cf63ba93855bf275758281a517adb76f511dfe12913daf032cc37
z5fba3dc91315f60891613e2bb98d3c8ea9dcd35ba5f7746e4635fc5e2fb787424443a4f8b13cfa
z0699e21905f1a07c96ee2da2b4975b782f4601eb34727ea5fb4c21bd49ccf4021ce12e40f0bbf9
z7f2435471f41f0a34f1bf26ba4c489e568c526194102f43c08cd79f434b88e7ac894cd1ab8bf35
z41531299ebf8f93eaf640d1767b6e70206d32435107155da9dab66ee88be51624289064479814a
z589018b913f60f042205c6f0e4fb0e180b67c664abea7d3f658d4dbc6faf63c8bd2b8d4f701e18
z11dfa6f7dbce6cda13fc2c606737e4f4b2395ca7395c5b94c57dedac44661c2d3d59ed337a93a8
z1cdf52c2d12a0a16b13ff8e9cfb52bcdcaa6f4d448681480583cd0e1b48f22bac51a4c6e63c20e
ze393e53b8b1a80613b36610d9a7ccd7d361c44c30f240e0224f832628c803408e2f85a25f25f03
zd4b66e4ba1f0c570280f0735ef4417f0c62acd98820647b35b2ebc96fc3cb5bfc2e46b818f7c64
z1523d4c57567a807744b785a23f83ed362f205d39a686fda88b4e95d3d48b00a2ac393459388de
z9f6eb4a42062ee7238da86fa4ba615edadc5761606c41b1ec3d12ddf66e75cc3f2df98c0429c52
z48027e3331d7b58308fe000d17f881543cebfcd4becc7adabb368408bf326c3c3867a65304dc8d
zc8574e766541cd80cc82be52c3ce7f71cb15b844d779038d59edbace27d97c006e7cadbd2fb7d6
z7de9367b933b552b74b9d32f37b1a854e3906a04a5d98b4ccac4bdb10630dd51627d18360b8bda
zeb60600e742fc4aaa3a819a8db9e1280098b50714274a55216419b2c67777fbc934c0df583b6cf
z6a83cce6c94ba8cd379e13e78730887d8fa745c2847d987a185e74e47d012ac5a2997da970473d
z53909c8292be7f14256365258157ad1a7d10e6193fb8e209e25507487e894ed5530b11179c51df
z12cec8214f7bccd956bbca07f172e7ea44be2148bb0ce7c4bad27867484c3373097ee2ec5f2200
z8304c10e965202070c9618de3fbe7bed281bb41f3d6c2c75fefa85d2b4b437edf1655c1d0f5a70
z1ef0899a6f9196f66ab075149679ef88a750191bad506f83730f4e95218f62d84b7efcf9570b9e
z52c8578225608541f4b1a4481c2bd6c827853a1179523b4e46bf85d345a7939368cad98bfcefa0
ze3171e4a83d8c7fdc5a0c2f1c8d126895ca3c7820f6bd2d71ef6b55b1471882fe8f5046d7e1921
z6dc4cbf8153737635ea802c493b07ee8a417a26bf59658197f1d742253c476ff054729d9fd6939
z2dd2f16601f5ecc745e139c62795017ea8aa3ebea3ce3a858f5ae82625e5942e78c2e773c83e46
zcd345cdd9efe249dbde18206091deb2aaed3a8e20b4dc41b61a05358a56f5889868295ad1a32fb
z335b7381f1d04d84eb38881429f7d584021bf0c1de0224d4df87f271eb9f2c8f02a17d5d87c564
zca7fe536425b8063e8b780de927a74a6d68e55b476944b01e8c864662655a8a52b2599922eb524
z97caf2d367239dca41be27236e603bfc820d19b1a157e568b8a7b256d2d21ef292152c3892966e
z0ff04c44755f859bc5386bd4ff059061802b3136430fdcb6e357cc0de6b3da8664e3b1d065713d
z000734a06d4efedc0c71fd01a9c57aec39d13c24ac192f020de2f2d1c1f38fc7e24a462303accd
z77a6540753fe177863c828ad04668c6284be59defd01435d7fed345dc1b54bb5edd92e87985090
zd88aa072c8364c5a211b23d44752dbe85cce282a3a6375a18d4b2f572a603c7f5255e38e2ea981
zd6f468fbfc9f7f6c906a11e4cd3d9b748268842c2b3dcf00d0b639598f0afdc37990d95325d236
ze69df2d8b133c17a7057f8157217a71a28f0e97fd3c640d104bba5c9bf89e127005cb5b016f76d
z991e453397df29d572e28c7d66f5ec353c7f1c5c2b2f124898232305e53865323950396de47269
z5dc463f327a3b79e3f0638ad8a812cc46fb151eee510e0c96034b011c702de4dc3b33fd29bfc3e
z08bbfc75ab2ba6096c245605be42df9da0db0cc46c9203c999c497997fdd4b63ba043bdca16e5e
z18c3b12ddca4354b58809c0c31d97e35c402acc09db6c08265bbccbf99672ecc1551aa35d67a59
z0b98ec0eadeb130c6ba725b136114fa602f00bc3c1b3cc2485bfc0b0b0283ebd6c255095ab875b
z12289fd768d55eda922c52310eb9498fcb36391bae772d789fca6757dd06f116c8d8d54ec71648
z3f489e4178eccf887f1ed263fd0e6bae00d887c415009a1c6ebb0b93136d7673ac1dee86f5e756
z4314f3d8c32880d954d57f91645c2667b909179877e5abb46ff340c76aa0e3623c54fc2cf2a447
zbc758eb529aecaa1bea168803acc654784eb5ab55f36483a24ac5d2ba823fdbdd4ba747a78e64e
zc09222dfab32f0fa571c17dde7876cc600afd7f80644b8ae33a7a041fef3e75d6413029006d355
zba9780f6e4a0e633fd9f7e77227df1c0f71331986d7eab4526f9ee53c8c80a4143ff1c1c68c885
z9b592678f43bf89e988700ff8b4532fcf15930649732feb9eeb462e822f0b8d98bec441e5aefd9
z203499ff158a765ce0a2495605cdc07f0c7bb0aadc017b14e318f499d4026f12eb1dc4646cccae
z49f9be4f362a3254f7794014f17ac1538138dcb182484f240e78be1ae2d5491be87484fec216b8
z968429502e20ee84cc7af24acb441c0c4f07283aa818c490586d5ce0a3be937b10e5983d0504a1
ze4a786a9b79872522f0016d911b1ffd2c4cd9e8408bfbff9003aca8e509a1dc3e4d5fcb34cef9e
z4907d239f43744c6fed4c9743e3ae1c56c2092ac645f47ff9a54c2f1a228957a2253f66170b068
z430131d5e50b69e336fae5e43988785697932179c4211d03a47a1e64551aa1441ae5cd6c531958
z135e0480402083c6cbba3db594eafe876313523dae4f1d0a15681758a49cd09e562cff5faad4aa
z5e9db37b961ef8d414b372637b2ccc8c673d238ec92a1d36ccd9acef5adaf4a5906b7be22209f6
zc848c1550778c3d597410145f05826c2874851777561745b2aebba6b5b110393896e5f5356b290
zde0ba06c9e538d80dab1fdefda2b63ad86740f7e7e93deaea8699299400554b6a2dc249bf33a17
zb7a3cbc499f5f1033fdcc45d0b1c9c3a69e81baa7f4db578f4233f747417a25661958df9a3ac76
zc67ca146599b6f6a1105ec91447185d70343c8f8176c8c97ce95b4bbf351e5553bb8aa28a77c10
z6625e6dca19ebd62c5ec9692bec030364211c91703a3f97fc7babeebd746eeef557e6befe41942
zb7bbd4c31f2bb12a70a8be80d86f3cdc2debeeb3bf8b753c7febc1242499ae422e2759b5d0695f
zc7eef382f5650536e8065c3918a4697df06bb5dd96c3d142e1813975700f399cf347b0961de47e
z76a1c63de25932aff25bd6e57be2f9118bd1ea1f06fa0e7dd751cd5f480f6765789e0a2320f544
z9a6c5d5222715c44f0a206b059e33f11d990edc4b0ab1c0f2276559871cc89bd7e2d6fc98451cb
z4acbad22db1884143759bc7e291db48a6e80e6a6ee81115bc17926d930dfc4f0b6bd0df85560f1
zbcb0f145a960cadd3af56d716f4d44f9c00c6745413ade5b8f1ab260b5a205e945454bc2d2051b
z017e3edda36122973b46d348ff92a72922694acd4e4da8fc0e1a1d30122bce12a9854db37bd9f1
zf291ceb7c609bff5b195147eb9bd1513ecd9dd6b6ef5f189da25f72cf712d70ddbd85ced5d19a3
zd1631503cbcfea6af1c384c7b50b5e400a03a75133bd9fd6b545b7c58b5c4cbd4c0b8116ff7f82
zef01b7b59e5267eb6ae42258e256eaba58ac23fff4c629010acadd6acbc906b2761c3822514079
z9a0b20fe727868d397ccd0fd72eef5f62061adb5e5c124a6587320a7cde4d1eba11a226db14b25
zdbf3f0b2052540ebb977eb28074af20426e005f0467c79ca9d161b6b2d1141ea304431bec2b238
z9de2cb5bb14e4881cef93153dedf7f4ef5dee7416a473a87c181b50884330c672d302361838b07
ze179e089caf49700dcd78a422def752ad97c52c6d1004eeab58ecf5ab435f4e619e6eb85aad8ba
z239bd38f9d20581c190d860174760dff9bc08d8b1b27991a97f2eb27e73ea3249637899afbd57b
z23a347c39dd871961712e92710838fd6ebbc29db5b0ff5a625ded421bceb55dacbbd4b2e5170d7
z56521639892f782e0abdf86a849fe4a10f7cf5761eeb6556fba0477e44b15594b97f6d955891c1
z238b2fe4fcd2beef32576b5e88eb52881d3e7954132630d82807062187d557888031d86a89b4b8
zb24bc571f5e8833772dfaa89230d92a8668e8eed14f22a187522dbe3ea7d32590cab9c3a313926
z7e05221636af595a311e7a775b8c8eb9f41d956ff3ec77e6cb7c97b28aa50437efe6c7c847cb20
z7b2d9ee7dd9e121178c958b4ca95b8158f7e619122d864a2a71e245438c8fb4bcc07b52ea5bcfd
z770ccf7ca0a5daca315e69ffbb98eb6be787c4b88e9048c9f1d7b7936036c8e2d54c9774ebf5d8
z09b3d24fe79e7298e2ea671b4d9842fd7d3c2d48684eebd40dbc8631cb68c3b3e36c16daa15fe3
z21cb9c46d8ee957e7396ed472d9add40b98040ee400031d4660b622e3156187b619e24da6a6be4
z40b3f43ffe1ebe4cca861e5f5000a68827992c346609d13df53f75e6f29125c66691b33ea840ef
z4d17f3552a745c6eb9e8aaa6fd1831c5353806347e126c9fcc6005f6fa646bb3a44974eddc5e4a
z31f9c5a5d46e757e28bd80508f21fad77653455e33cd3c79c1566201ddd5849a7158254f039b0b
z161f00aebcddee6b8ad3155df13b272700bc244990d7e3f3db9c225b363df8970758bb3f9b4d06
z547a7837ca07350f1e8ed0dbc122c28285e0e23a0434aa978e3ff271c4441b8bc04680865e0a22
z6342d68b75ab5d44ba4c59ed7bb381fadd489eed28f41556578c9b94d42cec8af5831084c26871
z312cdcd784f1b5370a652be1dd92d51a571788bb8b060cd9b4d2a1f002f1394d920ebb63459b9f
zb15d09a0064f6488c06fd1eb37a8117111ff0ce1eba530c09bf4c1bf68ff3dc26aacf39ed7ab49
z25b22dc1972e5be79285846de69f2cf290a3448d54f813bff0709d682563fdd464f12d23db7efb
zf8b232bc17a92ef4aea6ce21dfb53bd36aa89d60387783c8f0405d3f0fdd33b7aba69d1651c36a
z4396d5ec5594e50e3c97246df136a485f7f9d724503a157076578d5bec77ca2ec90239bcbe3ad4
z17561faa967137688595264533f6c04115a9e09e18d37515a26e37b28bf70ec49f425d6464684b
zad7f3ef057d81c95d0bd9a577f3ef526740976c651afab6c27b4b71bbfbc69fe434163ffc4022d
zfe3d43a8e19c5687c13756e8a61a530aecb696381390dfafb95a902eb7a2147e875ac0a24f40bc
z5e5a7b595310e1e4396194c060b9180072ae16056e704e4a6705ca3b70167a5928e254b5166abc
z03a46ab5874bb064ebbc612a6c403678bff6edc1ac52fdfef3fc0f1ac62f02c98cf41c7a336c1d
z38128270d17b70c43cffddebd9f9a49fe1c305180777aa49023ac498aba7e5096b7ac042756431
z00408ab10d4fc623097dd80554d1486b12aca8ebb3291d048c9fb8b3829748038aa2b182d55f2c
z57d57c53587a1f56de1dde589c86f7bff3f9267b6c95d671e1379766a030efe9b41d10067b7ca5
z1739c2e7c534310a27e1df7d633eb6f74d209e53db7be0c0ab1a9127acfbc1cfb2d1a2d4c8cf14
ze2bdd00217ea351c1ea3ba33599d7e78c18648a045bb6f8cab9b9bc6b13b1dbea2815274dd4460
z830ad98f0fecbc38754510273a45f0363a00e521d9aa4a87bf382478d3f91e5e206cfbb823d6db
ze6867e5ed2f35c84a2bf9047fa4ebc16bfae79781869a74710e54327faaef36a9d32f3dde533ac
z1802087d107986490a02dc7359121156a2869c52b10a73ee19cf5ee640ae2ab0ef0a92ab3f5595
z3513fbc39a29f7fdfd579eb978b2d56c6e6d73935843e06b709ae1f9d8291267dbf7a5436a9d97
z493fd300f95a954075a76d084f19d5d44b7ad458b3b253b898f6383a49191ae8abc0cfacfad7f2
zfaa631b35bab19069ccbbd9a63af6932c7e7d58fff253bb1d68822f392c88530154cccdad67604
z29730a9c5f59df98c50ef7bf7f80c37ddb1d5228e6b3af0f66c4d51f0e4105d09724eb301a1e55
z9dfcf9c8c984c4e3fb783a8996d2c285ece7a74c5914517d49786a9f8222a74dd463000b2b7813
ze98288a013ef20d1abbe1a8eb56e4cecd3dc1b53549216322ac5e42be370ec1f9ec659220bfa2f
z0fdd82e61879f9696ca9210278b68900fe06180c971ef5b64bfbd6e1f5568532c7337f0268e70b
zc614d5c5ccdb417bcdcb74a206033f99882a01caee2641a53e95f29d4b18eb4657dbf2fa62ae5c
z67e339966f8343f4d550bde010faa2a7988e1cd70ae57572bc1452c159b5fd336d7050f18511c4
z1f53cc305573187388a310ad26a1a6d47de69bf24948a6b2a3e9ab99fe94721f38feb9a4679940
z6d135fb58147e4e69f28869f8aa490532c90d014709c918be9d0992296a87ea107c06cb462c861
z01115b9b890ab450bfa4d4d0432a2e5f38609099c0184beb9118474e5799dc7084ce34d1b6e2e9
zd4e99af4729a571aa799e36af38263a1f7471ab0270e73b364be2680ccd87c60305e310b96dc05
z56b8930adc435fb87b70de86d276d81819a0bc5e9ac25c5f867fdc67cab2afcb1a6b177fca4149
z8ddcb1c74c881bb57d4da6fe026406431a61771a6ae932b2d78f2609527339068371c80a415500
za8a34ff3004751a58360c6698c73c8d52e7a912ba57bca40838a4f578a990f3f4e10dc9a8b1607
zd125b4bb5bb48def819334fb01cc3a6ece78f7d7de47ad4c74d36e24bc76cbd43df951c1dd78bf
z82b44ca4f8cd8e16f14b59c8cc72ee9a244806129962d17b28e29ab4f3b102343b85d8d3cbddd6
z876aef7876b8486ac3ab63cd592a5f74dd7d3583adbe146fcce3b3051cdd991629f8f9e441367c
z5ad0ebf2324a1ced3af74755a813f970002263f9772bb07d1c8b67c0578d8937ccfc32a044ad70
z48baaa511fd147d9c88f495bcd4130b21d07aea312b0ab702c9bb8253f4e8a39d95bfd916d0e8d
zde737a740e1b9932380c49340c2468e3e56d45a3cd75d77c206304bd1684c01464703183fa1865
z1540ecc7311bfdbc199d2750842f38df7a772f9b90e2570402d1ac9a55f6f2fe490a0d8a329d29
z2fe08d3395172222d5ea7e2ea8c66c6acc1812ae0b8e58cc34066862308d2b3b431c184351bad7
za22403a80021729a187fb439d35ca8551688b8cd513784ecd69b68564d51e853d13ac96cfe3275
ze1a2fd57a45b61bdff9d4a55085ff11cd21a6f3bdb019f6d8221d8ab20902c59102cadb35e9250
zf1713c47c4c7150fe6b5278529eb5b90bdb0be762adcdb860c5f445545e16613d7b40596105d85
z4d39309306e528e665ad8c57c3745f0bb1ab3fe749b216e8e9e59adf9474315d158996999ec3ff
zd11e9c551361162f876af09fe07d13945ef9bfd6319f5f22d7a31166bcdd67a17c2a588308d152
z42c27533991aca7d7663a9522afa549969fa7f43742f9c4706578f3387659109e9d715d62ca633
za3df34581e5d41d52c370259c20c3953c6591a0097d10da86f3c70e0258401cb5d1c70d05c1f3c
z3ab0a84f4c115d56d3fb53d315d4297d6a48aa52b78eec5dd3a8373517c930463559c7376a33e0
z3fa3eea103d18ede47ad995e0017d0d6865b6d0f50a20681629a9841465abb935298c60a5993fc
z77c6db163d2312b3e11ee6a3e765759ea4df3de894ed50db0dc6bd3add87b6977e415f99fba3c5
z86e3bf27a45cc0f9f8ba8858e9197b0ff417794e1d751fd38780721544d1c6dd392feb8e02848f
z1a2b1bf8255fea7e73212948272b1d2efc7b1beb5fa2d90e3b63a77b61831e0a3453f702eeba2f
zc96f1a185ecaf81bab6cd4b8b11634661079462de5f351e9920bb8e56794bf3d9c6552708f63c2
zad0a6f9d87c67cfa1fec672f4a9a68b2e65c4a90f87e378007f6653f566466071ff1aac113706c
z90a50b55f1a17ca1008946f3f787a19733ca575926f50924e0f0dc2d23d72b142a5158581f9e07
z5f77be9a342e24222c61db9c09006afd413d6177fd931b348d4cb8e29cf895e50e049d4b64df15
z568c25aa02853020ba6b38f1c4197da526c6464ace9381672b8a003e7e76380c2ace04a82deb16
zafe93276565b3b0f0962aa3d49f06b473c33e0ed6df5c0730013c2b0425befac786083853d95ad
z3899c222b5cb9615063573c3124907679824564b4cbb645cc58d8b2dfedad42e0b034bfd69c0e0
z82fdc205566b7cfbedc91f486577613d8ce1602e7b1456ceb5c9d830633beb1699aed94d4eabcb
z02181cd74b2fb3b0e9f6f80b04ac224f1f3162edf505674424c9d63c61ac4580c57228bca130be
z57d21053090c7bf7dc797c554313e75261c2e48cdb48151e2758d25f51974bf2433b692c067faa
z2a1cff5d69b98b6951d54e79ba682aa790e6b5256e3d51b7b82a5a0c6638023e40ca0d07ff73aa
z162146fddcaa202692702c2ae7f08810aef44bfe412370d1bdc10ab3ee0601edffad37fede5d6f
zab9aa3b05c08ac6782f368d7e0769c5491ad7eb991d0fde424f92fdee175f2cb8a0991cc90339c
z1c1f5c34b071fe1545a2a94b835836a63bf88b439017d8341ad034917a81c267c5b7d05bf621f0
z94a80a96a0741cb3a800ac46e67c97129df66510a18ccd9678848c0400bb2e6cf0451d63e0ee87
z3cc765b0fd60a30f903810fb4dd71d14850e70738a39e9d7b504b416135e5a617fdf294141d431
zba9183070c53182870a38ba12ec0a529591806b2a17111c3195dcafc0a02a0a0a36a620a02d9ee
zcf631ba09f9d4771a28190290a2ba88e2735c726d7cb2c492bee2df9e1dd0af19b1b88db326355
z12c72e254dd722f0214f438568baf0e038ae4e4036c9d8a8917bef674d4df85ef1d93b5c91ad6c
z3e816461f486ed17e18569ed5da9c971013ab2fe9d5493cf06cd574941b886c8f6243b6540d690
z9cecac164b049bd7ca66c2f29e2afbb56eb103cdeacad89258c6286685b0b12d9bfce7bb6207b2
z631a46749498575d0cac3df366f74aed16a4a02bcbd367ed45073c2c94bb5e6a892845b103be50
z2aa9a058f7cdee265ff6e48164c7f6fe584c48b1b6008eca7b038bcb4999d6660b43d912034b72
ze2033b1efae401a3233a3d833186e6a44c008f2a56ba5b947e9c833d9b1e62602a11c8af4be0a8
zf9f0fb73f4410023916107b3cf945ee289d5fe29750ef81b23297ea810346bf3392531ed028c33
za3cae4534c6450357720308be3e2e2a914dee8d77deff6b486c1f8a23693989c87aa0dfc823ef2
z53283fd311660af9e34fa2a42798c1c6d2dd72a8844a7074d31bfd6d10a83731c445bad5aa72f7
z1433adaeb85e9a5440548aa2e333073fd74dc9dbda78e8755802bf21bb0ee3544e060a167c7ee0
zbce5cd3532428ffc3811b970e9dedcf88bdc355fbd3e900f2265ae707a846ff07c42235e1d3ed9
za81a014e84458ff8b843e6f3f60f5e73bbc4d022922cbdf5067d5b0186d031763d73841a97ca53
z95ef991fae524c9f7e5b84712076f1ed81aafaf029e022e0120e2e25a9d050caa132a919c515ae
z55e032f248f4f4ba0ebe1bda485381de4aa44ec634f5c5cf60eb63df079650d167da1f8b9c573f
z77f5d70474df8a095188100d5bdc847f553ab6060b1959bd860f0e228c8bda8e4fa06b43fbe579
z5443f585672eac94f0fbf2aa7c2239b8c859dcd415213856edb7ca4a3be9d4e0e15ed37085f9ac
z0cb1be68c8370dbd26e93a4f0b2e27d3f76abd613d61188156f0e72d6444bfe36d14e12f6205ae
z2f9b7da3c78441e36395802c67baa4abcbca51b69201fb3b3bd01ca7e009d47c154fd81435fa3a
z43f9d91ee89a3c05975b3ecd5479d03e1327351e26e2c30c69c9a0e62c23fd8bd7b6fc0276d46b
zd4d0fb693d78df18873313f7ff4f9f6f0fe5f97f5d849a254171809b1b8df5ecc5ac0a8cedb9cf
z9f8a8ff531ab312c42a134121d7521e85edfd360289f1449da368249180982f6553fdd4596699d
z8c136763a46abc343f1c66bc9db984824f4f69404206f68991b4a9a7ec4148364328e68bed9f58
ze63b666b63c848f087253280cd266b38ad2029d73507288ee4abb6774e3225360fb5530ff7a171
za621340ff868e2e7a7ed665d0d4ceabfb4bbfe3147a9451f2e260ec3f58d6b58d88b775c47f43e
zfd4719d44e015628c00441c6a9b610a4f2bf08562de5d22be85393d131b50261b3392ba89e8e54
za32d161e0b3a06783693e1343d246c0db49ad531010025b227ea1e78f58ba631730f2e2fd9c516
za5bc6866480fca6e19e19f01d1542dc357fae1f80595ff9537d8bf08e7492d58329e74223c15bd
z57dc54d108d6281c2189f7f4453904aa61ccfe9fbb707c0c4c5a3fcd5af1ee0f1bd1d4e8e8e518
z2627f0abac3220766f2fd2691d0ef060acb96ad43495af5e398212acb912c5e487dc7abd5ec6f3
z38bb30e5f807e1cbd49936e0b7b5b3922f4b2cbe3df0a94c90e753a8b67e3eed2718d6495c42c3
zeac9af545199ec6433a64031fea72c6badc5a162b2e5a9c1d49065725bd26c00712ce237adcb6c
z786a56c0922016c6501488688eb855833a2e5468fecd35fc752462d99fba9feb006e9367adaa40
zf9cb34c1fd638ee3762928a6a04701f5ae70f81ce4c881974e1476de9e4011859170e960efebf6
z38c03e8fef9c53257e6cfe0675fe677f0db6c2fe98967b1a3a9261437fba8c8d6ff64fd452898f
z1442853cbbbec4ebee8ae6b26a4812d5f6b4d29a3dc75ada416f3f592bdf59cdbcc49e865e4a15
zfe47c4dd30cc95d4bacb467b70c569f788cec7df1089563bc39e7a1cbadc5a42f41974d960e0ed
z195213bb9a6a5aa78cfacd68f0314061d9c9113dbae7cbe96a0d4a13b49029c9686ee7c0b8563b
z7d92b558e7f1b8d4d016a603939e6e030b1f16c0fea00f0241b5d5e6202a11a399404fd6ca7f1a
zc56f75de55f5291f12727ea1cafb4027d60273559a8f992cadc9cc73a59b2adec8e39862793557
ze72cbba3a2a2937170415b0b36784c1dffe4b517c50f1099b0b17a113d296e8ffa6f6d2eedd48e
z2adde0fabae5242ddf4cdf3444b87e04944b2df5ab31cbe32af1e2b4f0a00b285f0bc3bf312c7b
z6cf749883cdde8b1f54d775bd9bfa52307ef1aa94c38d4b078b199fd6da472a80a26a4c08e6300
za5ec85cb7719f72c02b5ee9fee0eaadf52222fdfe9e76e57eae9371c98fac5528c0c1d633c39ff
zde1f2608e327c19d0411c065829c3c4a61725abfaec22779f01c47c90b932621568488f909bc92
z79950cad086ba63c33af44c1b7540d270180f601655127727c7e2706bb2910c3bf43014346853a
z2e3bb9d03f327593098e57ddce3c1da76151f275a7edbc90c72cff9054310210b4e8cd805f3916
z29317023b9659622bde19f8e181b6a5923621a6d699a0e7c388ac441f3fcfe186825404cd1b593
zc83975c96ea07b3d820d6ba524719153562bcef0c25126cc652a01d8b09fafc8e0743aed935390
z7325a7351060040a4c8c481546da73af5419a303302bf87edff6f9944f0c12edf4e8d8ab761e99
zb1566b9c20df087a182ac6fa883a40ebc706800c0ca52cc5183383d2d4561436f38f75f313e6ae
zf16fdcbc0bb47fe5a2facbc2bd450ca761e9e9855a85b939fc706885e9e26fd7728ec80d1b455a
z16d7b0a3a314f3782b5a848ce4531107d57ab51afcc45d5752b893b32fe8d97b110b8f760bdbc3
z1d9adf6f6a0ae1c05472a3d2a8f122e4b7f8458041c397b6bb6eab1ed1dff8af24b75c709d6341
z606bda32b3f20024da51ef10b3c5390402333b84cc545f078036a22eae5fa6d328f0c53eb753b2
z481fe9177f2fe51cc447b398531b476d06bffbd0c836a4524d45bcf3e87d74c9ac4981dffb7105
z94b001d7fa5df198f66409776131bcfac5e603068e291baa1e994bb014684fc814681301ef2965
z8556c6009bd47fff07da8e7aec772b785042d672912620ac8971986b1ce1c04ecb138ea18c521a
z1c84446f1ef9e249f942ad9db3d6bc387671bd02749d538c423f0413e1c16dc0e5cc20a7b89cc1
z1b1465feb6ffe6f6421682365305364e8b1f2bda084ba6f523f6a4ef6666549babcb99c568dcc7
z650992b791b2c725a8f2b688a4d33d36be6c46b503d2171cfe5871db09fd3b056df2eaa6423ba5
z2295989610279c15f1c5e41149310d491fcbe14bc96dfe38474693417efb9fce7d065db0b0f2e1
zc492e99fd397ef8170e108e6650307cdf4bc145858f70b9b321a05025e9bba390fed22af75ec07
zbaf14740203e2b549af369b49d4fbfc6237a9303cfadab688367e6a6fb076f160ed91e83b55cd6
z55365a97cb05ef0838ed87ff018ba1483371881b50c13292c076cfff721dbb60cbb0c6c9e26f1e
za263793319912ba222df8748f00806079e2936687bc8f17543ad7ee1eefa90a99802b740566fc5
zc76a9726005a560a8625c4e06fe851d0db8d1e207c35cdf7cabbd4e67ab8b9e5994dbbafe96080
za53c9e525918095fe75f0d0e94f2547e5ea034aae0da35a03010740833b65be0e5c512f4df5f28
z33412cee445f278d0ee43a7e194fd534073c08ddce0a7578300919bb1ef9e449b1076945cce633
zb3a7b49e71c495c51d5ed1b91f592235c5bed9de8b31e640c6c76f8f613c5ae15951e8d57b8654
z546719926873eb3311717bec854beffee243daf0a9ec1deb51ffa5149cc4d01c868bc5d5fd6091
zbb2a71795fabcd5b1f32126ee93bd602b38019754707ac6cb7a0899bf255acc690a19ef137f23e
z6b93efe941f74680bd841ec13eea19deb9a9f46bb727eeab033db39681aeed283cb409dcd0de7f
z3a43ecf5750704a5e612fb71df767d268f268dab4d4f5df2025d4ae098a1452f5c404a079ec5bf
z37bb193ab4dc9d75742b298b03b6280c8eeacb36b62e1f4be5df297b91afabfb895f314ada6de4
z17633beb65b80f2c01ad64c81844235bd9e29ec991704b1eed2e6e2efe0b8c7eab61a56e86c267
z67647249227703e526fcf23b4ccbbcc77382db237ccda5f1fba27a880ebe05b7539c02459e6596
zaa2fbce3fe5004e81119a55cb17f7ca82878070c0316ab790d580690c6bebbd9bb18877bd385f6
zf71daccccd2b6953a53cadf13bc685668a5837a6928a91c719ccc28d181e618eba6a77630383cc
z2d06f5b8012c4520ae33d897c6185a9ae4739470e56b09d7eb196002e7098e3ad7b14147d50aa6
z36f43b18f96a7e00e277d2dd7039d08e6e731270f5e2615abac0dd66c1c548dbfcbfc487df8cd2
z4d596ad56279ce50fdfa4c981f438a446fdbb670168ccf045e3420dda4b98c723aba34ae2b7e55
z5ebe325c365005f521a22df77058e06d3e797d143bf8cdedaca5ae82cfadfed6ee7b7a556108da
ze85e54828283ed9bac86114fdd8586e83e65e94705f28d1d2a53472ca798671027041a5445b763
z33c299566e3b2b6bd5130280a97541e9c19060d57d0cd1035010f3f46b41e518032ee5a1bf943d
z0812ba165032f92d8f2b371ec922218e7f7f8c16b3ac64e8139128b9ae54831d4b7d4d9bd3c39d
zac08d2f10be631ef43197cf93b343de329581207db08c2a7423c1c7ab95e954c247e1396589bda
zbe11dc9575cc938dd2c8b1db6100ba4d485d15857d80fa3ff710c20f4d80c377f1d86f4e769dd9
z7ab80760da47d0d633227e907ac19e82dd8bab833b6807acd309900e3e58f917ebdb0c9343a1f3
zb7da3f345fb2bb42a22ad86efc6ea18e08388c1fd7b1cf7ded1789e78d9ee169cf26328032dad5
zd889699126526df95a59c07da3c3b1267bd7744a16d14ac8cadd599c365b22dfeaad64d806bb63
zca712a92315a8116c70a9f8e1b7677f03c9231ee0132c571bf0c380a7c423a8b41fd86fcc4dc89
z261e85c0ff379f124f3b9a6f52f687ebb31650c3b7ba413ce78759aa82fea5314c1c3319f39ebe
z8349a9d4cbebe9ae8d5e617de6c244fa26f40bce7cd0202d8e9fcd1b1c3e0b8a00512c2c821be8
zb9538e41b3bbad414c895aa981b65e7ce86680c892ff234a909d324485a794e463bb89df7c7f4f
zd7a6c7560062307f9d3f2586fe7ade86a9cf2d11e40cb939d592ffae892d09504a4adcf1003cd8
ze07df730081378e9012cf248409c19adb5c9a60bbec6d5146cc1cbe20f49f300d89b8f6422469b
z776da44726f6412c7de7626dfcba481ebfb727581567b3184e7826e7324547ca36e73519efb5be
zb0a8c652475e0608a94e9a64e6ba92cbb8af9de202e4ecea3dcc52ef75a050c01c6160f2f75570
z6787ad9b3957f1072a1f2202ed943c9a1141cfd825d6585d2c339241b771f36d024338791e2e33
zfe14295cc75296fcb406fa3ec848e55f24514141caf28409e273fbe124cf8949f6089ba480a1f0
z485d4395599ce656b10c1360b8fc9e008ba2fbce63da06c93154aac9c01ff7c7da86204f12394b
zf3115a251d2d63d371543cf9aeea601c830ddfdf6964e0cbee223731049260088b5f242af9927f
z89896a65358227c6d5505652094b019b6f9496780c84fc8c5d85a4790319773ae6a94da2a86f13
zef175a06a8679e739763ed9c36a83abadd04b1af347ed6e3237995ebe6fc152ef13abaa99ae2fd
z6076240f3110794f3169a90b11793e7d2ac6a0e92e5783c7ee385098c60898cadd90d59bca3cb5
z00522f43adff8a247a7aa0e07a91e8e81a69f3a3515f2753692f02c5a4c3862ade6e3b4aabee34
ze2b9cd47fb67bd5012e4f8531e04e1426cc44ce81627df17d2230d207c51ee0b249ae3005a8ad3
z0eb6eb203598527019d2edb55192c44ef9959a12320c3421f221f4305c14e869a13c4d8d6e2b05
z8825ed38332603df51e0299a348dcb4c003a347ce555a365c68d4a9ab77e0411f081b23150943e
zd62dd22357537fa650c013568f781d45efebd1fc58a20b672c4ec2ae60c23c338e4de0ca0bfbd7
z1f0206b35275185ffc9afe84c8d0aa6ec2955727b36a6ea738c267ee2afab82860704ad615626b
z9b9c2e9e085d58b6a41e42baae86387fa49b20d0d0e54037ac0c4ddd4c84b82d6432d5a54f6807
z8e8f1d2ad0382d5822a859a6d54b4c1970705774e2be9795f95c8b6a9c55d0dbe4ee91276b52dd
z6da9e647b72ba6187faceea6cde448bb18229481feefdabb08d8e6703e2acc26a7c0832ff6f38e
zefb8d2976133cb408c3d834a4a91697f2ef2a2cc564c8a603174f1be4d442ac2a6b47e99a369e7
z73569a6e69628302c144766e462ee75cf35db990f9f1c8596fc383871390aa75759f6bc781e12a
zc64698dbb7661161bc44f706668fc5dc7c21a7ccd8dac0a11bb0a423f1662ca816724fea9bdc81
z12e2b641de1f883291abec920ff0984f0e19a937bc1964cb7463be5ab97be28e90cf1ac51be71a
z658d56ea3911e27a6c7bc387070632a14c4759b3cd5fc39586b11e0ebdf66fa27a65a8834394aa
z3a4fce464d533b25f38db1faee7d240c120284cb3df18405a7a9943c56924df0760f0f6e93413e
zca74538d126ea964ecdc7813a68d874253d9c7eebba47a039680b3a179a2cc0ae396424ecad56a
z180f49259a2ff039c463f9a474a9f85d236f8a87c806964dc41aac0518ec4b41804170a5dfded1
z1da682017fc9d0d1709ac34d216352bbe813cca3aac862604330e64bb5ce5c34b5bad5a3887efe
zed06334d8c0d5c1e6cdbc1591983980d4c07aaddfe26602c08eb4dc8ec4d16241f826612c7d775
z984f3ff414f3002f884dc2be71b03299e5818d5be148d08e9f52c318051f3fa4396c8798d08a16
z1677a414acddb2356195e6668431312c5d286292981204c2e069be5b6927800c7d29c2b72ac70b
zfc8a984dc18bc0bdd19dd136b1ee67bb106c8945c170503e3aecaa52508e09db76b2f4c0943ce0
zf95d2b4441185a7e9059f584f382bcd1e2349955da0cd4718de1b370fb913b0fadb693f444dbe6
z0c169073d6489278eabc8f111e9b3d827e1b509cebcc65507791b6e159d1da426cf22c18234967
z4d3f73f2b60a5dec8c4dfaa8e508d5f481251efa7f47fbb1a39f59fda2e5da5addb17752a3f7ee
zd4c0a13761aef4493d1cd4614c5c2b96703c83ff1c0f61a021fb6b322c5fb3f0b754813c3cf88d
z50ccf44f82f94d15832e9adb8b42567e56f4fa3c2f10f92096a1bf2d35e229f36485c081a85dfb
z6cc2387d419e08a1d7f4b5f4fdbe799fb7bc017dfbd202d232f44693e040abfb596d63c488712b
z74963850ee2b67d5abb10fcc1662385b4deeba64af38a4cd073a097f77245c69ea30767f948f11
z3d0d7e557b3eda862c61beed16469d58455789436173a2413dfc098bf61e03c89ff66a511d011a
zdcf366796c8f34533c4a1802a185bc3da554b37aa87508f8783fb03dabff63443c4670f8dd5950
zcec8730f016f04f7e6c3e0c54498cea4552905d6486fc21634aa84c4eabf08d1f506e33ea6db72
zfc63374ffd4c28321ec0ed8637bc5208f46f70af494cc3252171974e734ac0a96a4cb59f5843e7
z91d58962e18ca4ab5ffa066d3917d50a7db18bd84d2c0cb23fcbdb534c4440d0dcfef18446ae16
zd73d10dc1f69b2a0d61dc9a77c54b5c55c93878df54e27468976c8e8837f73ef09f5ecf68d28e5
zb2060c438976a4c87b1c366ab8bf950249918bb33b48a026c5579a180413f454f7948a21df1597
z8e24389538951b0d9462185adc9a73324afa9f05a89cc00fc708cdcb1aecd6b10b069d5ba45e21
za36c359975e0df3ffd619dbc560f1585c694dce337d0e47212da2df2ed3e95c5bafdc8a07ca812
z8cb29d2b475b773e1c8f0f4b3f62ab3413664a8585c4a2432d99624e267e3c5e7b61223c23d11e
zec5af84d46a6e6f94d8fc1a2582f1ba84aa3833b126f49b2d1c9199392e5f7cd8e4eeb1b7d8389
z642b0d824d914f7d0203b5c5058d40107d9c6a5761395e2f2d8b541b5b3bc60b0a3e5c04bf5b12
z3f3bfd0f6876cdff0231087035a0e28c9a7465120c79402fdac78f760e0d45ebbd05e63dc7933e
zd3843d63bdec1f3417586524f94663480cfa18c3df5ac177e1be59c09d02433629195a402af922
zb2e34fe8b35ad07ef301ed9452a9dd5c0e663bd39ac13088773264c55bb1dc395b1fbb23387f06
z0319661831c4f8fa7be31041db7c6db3555375567a419e397dae172ec8dc8cfb1c8251fab90be5
ze53bb2fc293996a5d3692c0c00510fa7d4b37acb7cd3eaed5c7191c4ab90fd3ee0328cccfd5942
z6b323d4cd481eec751d5b787df2572b8d8bec5ce5c600ce80da27ff77281c5919bb5a4a7b0142b
z8d260cb278e0b2485d9eecfbf82238ee31ab0ecbdec3fb3641923e6a12bb6a32f60e8744e7d38d
z063bf8d72e947e7bed968a33cd4371d7cf8cdc5f105cd249af9ce8afc754ba1478037cb798f45b
z1b01129149b92b6fd8b36ad8e4f3a488d22525b6fbfbb1cb8fa07195943d1b6e9d9c288878eb17
zf21ccf1aaf2327c0a2d22ba3944c5d39cdfdfcea7de534b4709aa0aeab91f7ec9e00a72aaed040
z3252eecb390e133607bd32d5a0f38421e718598dc34ea0f0577f1d1bc8065ce41c84121f1ac074
z26716f9a8918cd58c6e77a266cfa31c81191b159a81347d3318e6c311a931b621f98a48eae7bfc
z895c30ad4e3ef1303825de60884dd574e8071bc7ea88fe888e94eb0ed71865eb75d257be8af000
z2aa69079214ad0a9ef45f6b56c5f95f53e7bc09ed467d189bd9504f42b4c702c5ff94409b1f329
z304a8961c6671a0e5fbb3b25e49efc129d6ce553c24a7481cd96c45b12879ef5ba9138e5f98b9d
z79c3e07decbe5442b2196780886892c1d666d66bd7ad05b36510ca87d96e64ebeb880ce12c1641
z05e5e39a54e2bf10e97590708a178089cff32f34e4a9a8718121160e70c8b327c4854abb3aed09
z725aaafde3d80780851032a2866f6904f58ae8a4f3982fd7ccba79d52cea2a8e2a00ae41453709
ze07dbb32ae8213894f33198a25aca114c923aba68080ffe2e9a65bf99812ae580f5e48b843a0e4
zd45d625c116e2790e66739ff667d402bea59bff41ef3fa3231f7fd043f4dcfdfce5130ee704671
zc8a053ad46ef21e4724d338cf41d5ef5cf774c2af24b43bce2c5486f48e1cdc8278cc89c5924bd
z37cec1ec25aa8c6e0c017a0f48abd37713fae27860ac2de0f5a35dadcad5bdbe7aa7336b2a0be1
z286a826f1ec04364e29270c721b0b221370e024f2e07d239fbbb86d3bdd98340b97a9434504d38
zbe0a9818a5ea669354aec373737d07ebbf50fcd3a5db8acc82270aa2fa9a869ef2dd7429cb2fdb
z49587e0172632a7a881cbbe65faa32cc9f862ebe7e5b89a69f791a6cb54ad30c0a64aacbb02bc1
z61153630ad48c5857326bc893586b94fc669c7c5341aed2aae8645b49c4b6a5b021257dcd33e69
z801be58373793b5ec188ac9fb59e105daa4d1bde9e6001c9f2ff40b6ad1c172cbd1952fa99aa73
z7f58207072d67fd50d1c5a976fa5ae726d0872b29467474028fda9732c032b1f502aaa95f2f122
ze8c4dfe8363cfb36f39a257549822b014f32865d6abedcc78bf30e4f14cbe3560c4be2683997dd
zde975e451bf74ee8537eb1c2879371bce5d246e9590f0334fbd2ff63afd33603676fd91dc0da81
zca78e4ddddd6c34ac0ceafda5ca1c4e51a5b486733fb8a0d522f96f00bab89f5677d25c659b53b
z69c02d100e5f8cb607f6bedf1f7ed9423f52c7e450ee1fcfaead4d5e74827267d9e1c0f3638603
z83b427aa67080639a557d7648d4a28bd4452a2d05df28138230d62861597ee1e56961c4c9784ee
z9303cf810cd88dbda2b1585ac70d5df6315619fff7b3dd071f4df3c02d2a4b98ed48155f7b32bd
z5c13d520599aea6b6729330e239b444391834550f24894c55e3b02da868d27710fc2fdd1b48113
z0814db84f85ec3a7a8590f43f3017568d022589e172f8cdda55c38c91958810a665a4004c46525
z825606d790ffc5bd42717650a29278efb9c59affc03d315dd4e7de692017f7c62a41e2677882e3
z1b397dbf5733574283fa0f3f1a39303b2208e62418922200e2a7cbf34dbbc3064ebbb907a6625a
z7c540aea96cf422d6f29917958f974ee148dee3ee5c01f11525544bf3dd91163664a087da06993
zedf9deb1910918b6110fdf00bc5159aa08ac8dcaf83bc5510714cab5af8293662875c56f7c9f66
zd6e6ce64840dc026b500ad8720aa66df77233e4176b7abfe7c304d92e90486d8d2ded7e07668dd
z13f9c26c49d32b6d1ed1ccb6dcd75f27063bbeacc20f86ab1813b21ec52c09c129b83b6539729a
z536907986287dbd08f414ab6bdfff159d87e7a98ab21bc8af1dfe625b24a8acd877758cf819584
zbb1c3ccea4ca91a109adf78798605fc768bd3164e86ea1d520281f8da65f7eab0d97e615f7b14b
z7c84b5da507968e87ed5c8e7d1165485df1d9cf58d255c0b14df755a1b65e2b41b5960daa38b67
z46010c5c27e60114ef8bb3f579ddcd70a93ddbdb84f8bd55aad83a07904f58b8e5bc086e5f4703
zdf3924c05b77ad857f70ba407a7abd1b30ef57a6306b672dc1146ed8ad4ced57fc0ecdb0b4f40f
zd619c3ecac5afafeee52c4805b441cf300ba96fbfdcad701e548d874359c6014cf5530d98c538a
z3d99f0e0c96e2d6a655398658811b0155a813b315b1ae5c06ac83a7f208fbe7849760b275bb668
zc872b85086eafa6c6df7673fe91102c4c04c6197ee263692171c558929614c36a2f8aabfa7fa65
z4a602d43cefaace22d135d6acb20369c384635809c27b65213652b1a9c25fe0d9eb770506aea8e
z7cc3b70e126b03169beb0d43d05c3465a612f1f164f3be54c996e958cdd7c15c7fa1b051034f44
z553f15ab87331a240220d2e5d0d84c5ebe5f012e9961995cc65dfc3301c7ab3ade73915a6f194a
zb456c4c23f27ba8b9d2c6a5dd598433ae381877ca0f18dcc3935f51b2595e1354c4f1303e0716c
z63bf8a2d83a5d58e3717bf43ac87420a73f79e7fe9d54193bb4ce2e0e882845675974ad721ba9e
z2c7ad3ad1a019b58436cdfc650321c570759aeffb5710ba93107e6176c4ec098b415613ade59c4
z05b1754243ee5d414db209e758dfb8d0a5f96e61d01be92d9df55224a7916744cde1b1e5a34f3e
zbe9a36157c6dda87693b45c92b0e66cdfeb057d8b69b9a8f712f9a87f939621290d0603152dad4
zde926cd7c3b8d17859fa18e77f8af7b339099759093f45db64dc4e9f107328f107f1df0a868e63
z5edd695014df72cfe6b47335118bec259721e07cb9f50efdae571a8f1558e9144b6620f2465fda
z736cbbd98cf8f337c7753a776cf00615707dada62fdd63e23c6188a8c6f94b270f65054e06b5f2
zc741f84b1b2bad98a1e52e9bb058690e52bf11949d0105af54ddc7b32c9b64e9a5b96e77a4d021
z24edab3623369b79185e8756683fca42b3f6e173966c467276ff93b67bb5742198cf1f19a026dd
zdd3aa4097fd5995eb5dacc58ce3841ab48dbd7e91382368d007d6ab165a3c535d7c307256eb80d
zb4db99195cd4b3e23ce3e2fea1868e9fb2f304afe1dfc02ddefc46bf8f3919f8ccee9a73033f54
zb9ecbb008fefbc294a740e46fb172ce3d3c134e01a2b745e023c01b832d7bbea772b443d093115
z4e0cbf4bd0896787218d14fcb8d2539528ae9fc49c9c6b9debb205ea3eb2afa876a77a338c4f5a
ze1eb922c60d215126bb468de62d8663cbd914811f671c6cf83e2937f3d02e6d23fd17171ffc0ed
zd6c98b6d1731d39d90fcc6113580314e8ca7c5c51213e0d61a15cbc377586226307157f2c3b698
zaf7ae8abddfc0a88379303b3b3f44a36dfe38d0d0ae98952c35f792557e4933023b82a13b1dfe3
zc856fe34a174fff347bd9274c09a3207e5557cdb80d4439353cceb1f5d49dfcb77d660e78ef972
ze21acbaf8761991df33c7460ea1b3fddc23607e7e0183de0cf5b187d683f4b74015df9094f08da
z1f18540c003de14c51efac651202b0621a11a11aa5c572cffad6e525f932b21f6fa6d5b57342eb
z633b345e14b88281cb97119582e810d74506199ccb176b8f715e0aab3100baa8223d809ee2fb5d
z8651895089f87b7b21ddb616364fee2743f4cfeddab8c30a72cc471a36f1748f42a07931ec4832
ze800daba83f4e67b45f1f6c996c0f80201dcdb92cdaa3eaaf0be91739d1c638ec791006fdf30ff
zde1a6e6e24b861ba304d746606e9e74fb38a782470aabe2986f91a90a20f2279a61048c2d6bfcf
zd094d6905b4918fe649e4454ee924037067ddc9f2ba3b159121c8e9a3395378f15508c9b270eaa
zd8fa6a6df0403215be98781ae134fbb6b0f816b6168385ba67ef6f6361e17035fcdbca9cfb5483
z2aa0442da76b0971e11f1dac5691a7d9f82f65dc994775bec35aed31e6ad071b350839fa99eff5
z3a5aa78d3ca905524172176d052fd40cee3e57b5494c7a0481ab0cc59d86a7ece6b9bb9d266c72
zc25b37cb73efdba39514ed325a6fdeea6090d2fa4a8274ee3e381267350efd5e84263273062092
z3bd6e56025bf510e34a290d7d2886c4f50a74049bbffea7ac9311e83e7be4d6e62fa63905adf2f
z89837ca153ef860810dc3ed87f0eb2c9395586eff9a5d4708ca06f2ec037cb685b5f4d68faa8b9
zcfaa62cbd4b7b6f2d9836f429c4fa9c02981cfb81bbf1346d195ddc116fc92a918427aa733d257
zcbb99edbf6fae74e99a446bbb6612bb52defe926bb111f00210e30a8882cfbc8101db890d80a49
z3c9efca1cd88a13302d7c5808f492fd71843b85a33f88fd424003e72e02be81fb2a5adf69e621b
z11b5d0a86d73a4a9d4dfa36c64d440b0aa2a0b1ef2d6902d493c0b6095c230044b7bae2c89f406
z3f308ebd10d15c4d7b9f29c9d9f3c44d7c7a7ef91530bdf61fcb8190c1c9a74168a68288fadaae
z04bd92691b57feac7d079f88528091f5349c89f01a5a571ec1d1ba6af6b5f1a28dead381f4e2f9
z24551ff2492bd3e5997603672a83488163f7f25539158ba3de0c0294772ab57c28ecf6defa2f33
z1c7b1b6171e9bbdbeee9613cfbcde4e766fef6fdea15db9a167eefa12e826ecdeaf07c9491070b
z4c739790a466a3faf26971dcb6427b9cecd3b13a7011d2d911c1f6defd21d17b002f1e2601fcd7
z327ee8d04dc982e411aff547df8b60bf750be32f3ef26033403ee9548b814a947037ad2c9d8a7d
zed6618725f7199d1e71992dd07a0e0602f91eae0f939a994b396f972911ac764dd2ae85b540fb6
z975a1156ee3aecc137113e916a717c5d8df66c99100f46d6156b01c7f828ae838900558e3f91f3
zbd3c0db29fc5f4578e695bf98da5f16821178ade194855860e449fbb59747ecd5997436cd1991e
zb858e8f055112a9e06f44efda65707d66a97aba50c4838a452a839f3f8e427210320e0613f2780
z79082c5f862b8700ecbc017a86b6fdf520fd446e513031d320448474e0b57ee1fe15b2089af437
zc48bfb18069da1da399a2ef5a9ede2c83c56a7c4fdd8b3b0d5b323fad0931d0c69b3f4034d9e3b
z34df3529c4d7e71f9446bccdc78283118ebf834c5bc1f6028ef5f0aac6ad451ca11880959b4b55
z6fe239d91039de82c3c73d34b27527e21bffe5af4e8d839aeea4328b607e0b9d6d3167e60bdca9
zb661a4fb9a4736d2e5f8f9c941dfa8b11a5e3c35697d810eea6c475d07ca702423c3dd9512407e
z9c13edad964a28ae724e72ee013cc0ebf5d8b19fbd33dac5e377f56aaa4e38870a0ef3cd7b3d32
z8695782108876ff007649ba985b54bf521aab554eeadc6cbfe57fdbc0668ddfe36931211752317
zaf8eacb8ddfc5cecf07b51d192165568500d444cc55b407f02bd7302769770dc91e33af1488223
z5ea436408d940966f9962b9a39829a424655ea373cf44259b395e495259b6a6576b12d7c477edc
z0b7fb18823772d976451605238186b08fd907dcbf487ee04c4b72bec04d5e3cc5d0908f0f60ed2
z5e2011d1318a10b84212269e208124b6e861204990deb528db0cfad4b32915fb2f65e35b21d129
zd66a6a3073668f35f889fc975dd7d2841bb270b0dd6ca57176323397a897f9829dba5610c4a77f
z4066e45654bb70936e5df53acec9dff6dacd1daadf0558d32da3f980e49e1ac61feaf08f5d6736
zb42e4989abb37e06cb747e509413927a63daf1745e25609f95a68970b75b2e1f90f96acfb93f3d
zd698e50514500a277e172bf73ca203cc76b1e4a4d35d33e5306b2ec85881407bea86b86947c867
z9081ddc6e4890e6b7b1559994c0ca3a3fa10f3f523eb9382b392d43848de2c74aeaf427c011f56
z0ac40bf553afd225a6c541617dce6c07b4c2697032ecd132ba56be13c5f535a5315e4fb36757cc
z7d061aaee2097e42aed9b30e257219f749bef71d0e32d66eff09f905e39365715047b7fccd12b1
z80477d36b6df99e71833d2275506776316e5844484ae8efa0d6215018ed1963e07685f161e4a8b
z85ff2fd5312d7c3005f98aba8e3ce6b3fb394909d0114ddca22c368e7ba1dd00b4aa7418dae7b6
z4c559ece32651ddae53dcb9d86d686a949279a893919765d89b094e664e55cedcb619e012e3ed2
z5a59cd461f4698ca1261fc8319e581634613fcfb6b4c1477d462243559b5ed77f0f75a050b3ede
z147d3f4d378b102d53b5abcf572763737c9447c2af89d8e2422a7776c41d5da95a53173e0e9a38
zfe13514e02bf8d22c21b051d0e93fa02a9c919b9fa723f32ccc7972512eb05e2599edfac95cf0e
z7c05cf016e2104da1aeb53811881bea01d64050808ef5cf88421f0d0adf5f2abce1c10d6687f4f
z691917e3534c2e796378c2fc99807ab640e00ef4aa9f1c30631b17acfec304204261571427dffc
z149b35acaa0ff968914a0398464a20382b7d13ae32ae7c6d28b0637fb52e6de9ce09610031f48a
ze50f1e789de07b13ef3aa7368125d03d1bccc4f545155743b175a9104e7c8f09eafb837108a73a
z7ba474fdeaf59c362e84a64a7e19c7fec80e1a1fd3ac6068888e0708b49a970ae0717080796aa8
z9e961a2e2e90f99ad66581378da2ee0464dbd858ff9a26a46546e7f243f20986df45a0b08c18bf
z1c66cbcc2a4fd4ead21da656b15fd33b7a96b0c04f5838837198ce33bdbaaa2c11948e82400b4b
z24ae35f5dc0f4b689f836c5d6b25b6ea3540ef2e8da7318ced3a87a8bee7e962b608e9dafacf18
z74c12b39e95ae9ea78f07cf5220161e464752b18575adde776181e5f3704e0b479bdbe202d3c4b
zd91b1430e160e9e6507f81cc4af4db5c1faa079d1711f0f7f5b79d9f46b050999ff8a6b86c1ce2
z9e503d25b527df49aa3e61b489e19ada97da2d1381ff234c435f3824a2ec06aa055d5589e1bdbb
zc7523a545cbdc6fb86498f94ac8a9292e509e8aedce496b49d99d568742bb0ae2e188903b2695f
z512366d7b5625343b07b5b6ccc42487c382bf9384a69c9afe2c38e3a4577924fc91c73ef34316a
ze20d338917fd43525398c4bc9058e834599e33dc1c0389a8c4a53c0ed300461ebb0cb7865e9654
z0050406c40c7045d365f4f6c49abe835ca0610409471677d0a7e9b6bb759854bac79ff1966932f
z3b1104884215dc0609da41df30e48c2cc9685a3f70e86fc0f40492b66a79268ceec559e4110b7c
z49d241c273a723b24bad12bdfcc765ea109ca4ff2b5f328c61afb35ba4050e68cd3530d2ea1999
z89de4bcbfabac503e5f2a188419c2d6a9093bc8452db4ab5341266408212f87a5cefedd83a3216
z383afc55cea48f7d7b73031cf5a821607a1b250b61dce1f53957c9f9bf8a462b78e67cbe8ff1bb
zc956fc3743f01e93e9d78988311969e500585a8ab9017b5bf5668b304ba1b7d5ae2c83b56288e2
z892f0de57393735e48bcb57895df7f54f25c31eb06aaa4cadb0bdb770f097742ab76b0af0acde6
zb2b2e739d51bbea4551672ced45825c6fa54c6b42b3b0a7ed78f8db8ceebb7e5cc2ee4efc034c5
z652d1e832c851152b8f727afa6f1284de2af9d6710c8607b824c9451eb4f13bfbfd42a5f1ea886
zd76bbbbe55d94e310c8a7300fa748f2d553261bdee878545d9e9cc425dcc204317bdb9404dcc9c
z4d20d912f1730060447012cd601c88a143f9dc63856ddcd248e3aa8c05cadddea129431aca3ec4
zcf6611997ace0bc24b99633c27c827ea3962fe8d0d436a7ada899b8ed829b4aa4d6aca32d8027a
z7044e2cfb53edfe09f59c4af10d4b020825f31003f4aecb742511be15909c8cccc6a6a51b8be70
zba7ce045d20a465d919ab88e7e2e3282e3fe670e4514770e6d856471f2bb6c40abd2d0bca5ecf3
za1165a39f6af3ca55e3f79984126f664a07cea83d611a423ec0b101ec000b6270004da33b5ce49
zc2e1fee4fa2eab58518757f7c617767909c777091a77ceeb2e4d1bf751aac6c1c06ccd6fda2207
z9d23af4d448b4372a4b116032bb14d34b195b6fda596f16ee807feeb3e496a93c93189cd3a1140
zd9b77b4083779b4f3738ee93200d9d77c9bbc84568e50e39953e13a69b64f8cedd814f428dc9c4
zf4a88ecb01df481cadec857a81d15bb87777d2a8cac27f81e68e06988060bab19e42df28898972
z75ef308d4aea91732eb2de4ef21e04375bd86f7ade4b3dfa6025214cb6429424b54bcdbe565b8e
z63890ea2b02589f71d87b0ab617f7e31e478ae3c5a738db2f99d8c97bb8f990fbdc3031d78f3f9
z064e543ff7e5ac062dda5cc90b5832d477c4a3d452b197f9c5da1c76f3cd2305be3cdc35496503
z85c7f3ff16c99f6c4eb1fca369f7dd10ad360ff9982152dc23a6d4a3ac1f0ef366cceda95a8b5d
zb3f6223b42055be1fcbe92183951230589722d297ba8f6bf2a032e722d635f1f3f45c1d885cdd4
zb2d4612ce97910e825d5b2646219132f961d7e9d2ed1cd199699e66311278b9105256c4942b420
z8b6365b81de3681e2a7ff45ca38fb8ebe93b91c25cf15515bff3dfa9c28998eafda9421e1dc7d6
z24e441b0b6b00302abd6c370fda6e1068c57286030123f95adcec9801b9f56e2cf3c6d4aad0319
z0d031db73e7c1663f0bb6094a8248e17084aae2aa159be91fad23a19807e6ed4dfbae660dc77c1
z64b834737d0f3dc8809cd564663366ba481dd3c8f5e6c433e83e983ab824536ccb3f664f614de0
z7bc434c221b10647529d3ece8208ad17db22c183c631c75b12bfa08791ffb056e0cebf4ff1fa13
za3de1b7e05fffd7b866ab0440de61e10d1c760a7fde0efd366643ef800e1fcd7cce084dc38476b
z89a41ce7d167d1d6a08484d7854c8c67d311cfc608afb62622a4ee1396057b4ec40679f2c2bc4e
z0fd285c89982a2fd67c68e5a5fa5bd99ccfd116196a83f650729af0af8faa314bf86e56441b2c0
z5cfd226e9db0da2cf95ee9de0966cbe364a379eb8c2dcd216eb3b4ec98e9ae304eba7fc62e448f
z29553b621e9fcf21a25f184c4f28f4c23dea119bf64517466de03a6d965ce97ede6e85ae8c6f3e
z2c9cfc42b1f59842ee488170f63e7e9c3a43d83d5d0fc35e39ce3b3ad977b2cab6c36f1b9f69d2
zc3d500b510a833b0130558e43a9afe025272c23bf5b568598c18151ea92372ad49eb2a899c7990
z35a31d9a5b9fdb1b8fc4272800e7cb47df39d6236d95b2850f419ad72958e56e308cdca3a2cbc5
zee041a081ebf47ee0dd3e0bce3dcf6ddcb887be7f602bed70b83858b06544eb2763ca537791f8e
z22fadf8962125fb9496500c7ce5bb9eeb858ba211083ddbba545b96da3d7ca8cdd62217de9a6c2
zfcdd4cf6c8344fc7b1e46627b3c1047ec7b6f7e7bdb6afce2a195cd7321efb41f0bb674c4473f9
zabcc76a12c0697cac41152c7fcd84439e380e979433aa778893b34e74726d21656f76641823f00
z2f845ee5e627cbd5651fe6c9f857152ce3382c9f58da34ccf1f193377462d153e152aaabe801f7
zf81e5f27c4bd5b9c27c9135e6f3cfc88159ba41831521948308542a0c496cb5d67233f475359c7
z316c19375921484e1188912fa2560ccf2104663dfe73233f70170b3efd7a3e5ba4ae9ea01445cb
z081b21419afc10165da5876943bac9e1e0748202eb42ac18d91df03e92daa733203bcb1306c9e0
z44f7b528bdd5696b43ae03e71a26f574005be4c33aa1a701c73db9eeda73782fea1d37f9b218e2
z43f32bc22e81bc66d6aee816bbabfd6c6eb1dac0bbc5ea3e80b57845d35bc044fa31e43e275d6c
z7bf136c1ed4fbb1c22d1fa0f58da06e474926a99dfdddf930ad6ffb72d64906cecf09b444b4e98
z872bd8a942c4c6500c5802890974a769c4c7e2a5f5f7b2fa41d63b7df59486f23dc5108bc522e9
zba3f873d7f034cbe5a4c6d2f752879ac9d5911e50fc747fb3364dd26e26fad4e65c7c6c0c1afe0
z4dc5084f21faedb92da8252d620a5737c6a866dcb159bb654d08d5650a6edc249711f54220fd06
z44d8a8ffc6a87c49906a789b393e11a02db4e7f9f325b1f1efa38c6cfecfc56c9089e994619de2
zb1318866412022630f3eb51cb783ab5b781248ea356a7531e617098668fb9bd793f9578f294d4b
z4f80363d1b41037763a13b9985fad2e1622e4e2cf3c878abb3e92fa1e80142e0a0751c2c7ea14e
zcbb3d57dd92950fdf98066d429629f4f6c44a138cc618c39bb36067fb5031a28e555680170f4d1
z274b2ac91ad0c6938d18336c7396a60b1dc03107ab87436e079cc699255a9a0f9f2c5ca68d3f5e
z5edb5cca75bb2cc3de58deb8b188c8ca5bd11afd8b557646112f793d826465220fcadafcb9ffe1
zbb38c3e0c8b800b9cd5c52bf91796a8527e7a020a92e9758e009790d4bed02659e578d2f972e45
z2e85e659c8c995ac5007e9db25ba6091b35cf9316faac9888bae2a71b3fa79bc5edbf2bef55068
z7d3b68998c535d3860417f6adaa9780a456ce3d8d67c132da514e0411bb02460f716140e52a169
z1be84b5128848c0b4c429f8df9c032574d3915fa9b345e08ada25e76a34304497c7866be78860d
z23a8324b112b54bacbc9cd6dbf1cb6ed90db95f8f0f4f643182a9143ed4e92a7ea516164b2523b
z208c2cb2bb0069e3a4592b47aac6a9cbb9659bf31b8f243b67dda6d0c1100668b8b34b478c28cb
z5a2512f8f8da4fedfb35f58b633595185cadd01ed38680f462beec8f8ca45e80511cfb22f10518
z972b34205ed2a527cf2271a8bc915b1d1b57e6d05632bae59c4f706d5ce8480b77b8010e609c7f
z9b944717954025a02fa366da5168f41136a88a27fe6f8e6e3620eed015d63ea7bf4e6ad4bde386
z7e792353b2b71d068838aca66dd016e5b9cfe884903b86974666b9cb53419aabf78d75d3df47a6
z403d2b503d7a44452faca8456e6eaab26ca1cf0caed1794554eb054796b5a6ec8c726e9c829ce0
z55783571e558c1e4b84e4e80be8700cdae5e24e6520e9faff9edc5eec6d5dfdcfe595474634881
z8ef21b73ae8f42534fb70d67245faab7efff10e0b0741068fa58f643b5330e513a3c568c5775eb
z3a3a35daa8832563f22a8f6f7bf204de1719d4cb8350748947719addd18b2c0806853bd9e2db71
z36e03857d9a1d0627c46f8cc0bf3bce6fea7d282eedbf0d5ed1065db2d3a8d4de2c934396466fa
za820ef006d9af3203647e2bc33ada2f0b872271d11b8c5b620d9ed2265cab697efde6e422beca3
z2df22bb21ee9491082455eaa9161aa6c6a1ab03ba51f29b3f2d05d12de2337a10ebe597a76c2fc
z11ec354da6f674ff8a7787fa846673396e20178a447d7262d0723314dedc56b815680568229f7b
z71e53448cdaf81eb2246ec874e156ab1885f0224f6e543745a893eac63eacd287523e979d609ee
z52580fae08be29637ab6c63cb0eeeed5389c3b6a08caa7e1b4c068307709960603984f4594c017
zfc32c17d56e2cc7cb93494ccee5035ca755444c5ceed8067d15fca9866ec98570c017a17dfeb85
z608941a79f1ff2c5da10751b0c317d73606fbddeea38c2d2d22deb71361012ffdc4f9fbe410002
zcec08b3e9455f0be6f7e3aee3e6929772b9150e46b77aec74617855ce9ccd0c1dbe13cb95dbb10
ze3819f5744e04a08463bf9cdeafb402ac2138b4ba8f9afff7819b87345848ffa8d90361e223c75
za7b5b1202f487fc1c680fffa3521744ee8c90373b32240ea6f1799dfda6ea550e0d65f94787f9d
zea5a6dc2f69ce997a736b9d76b7851fe4acfbde744c7304a9e5c5b8d74f74d1e8e805fa9188fd0
z2a53153c36329e05ed601225d0b8c47e97e072a219cbb2fc0df154bea7a593f76f0faaa7baeb6f
z37d92b4ae5febb80a0a36a36de8b1e42a1d24b7c582fff0cd22c61c897f74e96629f5aa0f465e3
z55f64a1dada53c4b32e4c02c41f3dd05cf7f7d0046049d8817000dc08ad818e2424283bdeb21ea
z94abf3de11431d6c81c968c49d89bf627b6218279b241c062ac14db8d69dcd99eae5e03a8e01d7
z3becebc50972307056bdd5a180ed51abb450f151c99758a79360808437f405263ec5e82f7d9eb6
z691565fb027a2b41cc8aba524946e3077faf48effe19456adb4f97748dab36ce0f9f15c3a09605
zac424eb1c0115b1c1d1c24c6efe6bd7a16cf14932935f4f321e84fe978fca38a7ad43898096b8f
z66a7d7f4e0817e6048fcc7ebbab8188201140da59527a1b63ad1961a8985d111e5d0f32d4bbb8b
z1c86c81efcb169b2c5f9285db9b981827cd8d2f7d28845e11fc405357d93db9a324c6b53540d75
z6da2c97360b49974c00016ffb9b3a92f84efdd528bafa5d27ed4dcd555a494595fd6219a0c4e4c
zdc7ffa86bb1a826287c5678d702819aa100f93cf47cef5c1b2b5dc2abc3fafe79922e6699c83df
z0d0a2ed8a0531fac6fe8e89f0e2b6977d73d43b9f23a7dedf755c403e06d5cb4c07528dd378dd6
z3ea366771d10824d1d85d5727a07176f5297ed8e3a9d0b8dacd25868d81942ce5d548b58fd8e14
z49ea44a754e94763a638606b787a14a63e13c15b73459e3a659967d876edfc0b51f57057e4a058
zbad07d9bd382a9afab66a5d80edc0d25cb0a96cb7516d1380509f816b1fb197e5ab34c53b7cde5
zad8e5173e9027053baa0e10a9162957b22bedbd22a8da45053625c13172d615b122471d2373d3c
ze8db727074fb598eeaedab83b0869dcb70d8022b5109bfe6fc9839b35d480dd9dc984ecf45162e
z93052e46df9d19a305cbaff2bd29176914d22da123f319364d8d842dbba6b7734d8e627306cc6d
z3ce4e3f45a497356b222e85342408b07a3928183d78aba8608bb088e44dd608594001bf3bd30bf
z70e62185102eb19c48702557ff5179370e8875287d8eaad13017e6a00958e020e929ac2f3cbb84
z9e54f3ce8bf9a79ea10c6edb5d7e006a6f948a797240f2b158f659d2491af70b634a1951edc2d4
ze91f08f623aa4a0a95c0e83441326e8bee0633734e192ee49194ac9a800ab42d02e99bdb4d2870
zebf23490f09bee421f9f850b66d355732cbbde7dff1e27f12b85e1719b7b6d01fff3ee4530bcbe
zd8288be2d37e46d8f1b6ed312573395571f8c4e84c494565a22a85e8f2b5b94e0e6ff1bf3329ff
zd7a358bcb2a3257d1d4c49c01f9bbc1856864be2dfb10dbb4149c147e0fecb2b1c6a189a0f5d89
zba08406f591dbabd9f1de620ebf1df278d5f2555476b1f517c98752c04625d10d97a8205e94cb8
za9b6370589d2f3fc9d168ae537602af0d7be079127273cb05e18937ea34a5085434cce3be44c92
zedd6bf2593d2d5dead91ffc8adeb390ab111a1a9569d7ae40f2efed31f2615fdd72cf4fd55e7fa
zcb148bf3af22a030667ef1338fbedbe8cb327c4facc3fd474ae4e512be6027cb0c97b0e1f3fa24
z58f2f79d24eccf05fb499a97cb27793b0801175e2c0060f6d01d5e63f990e0713f9a02a804b55f
z23d61348b203d0e90d74e5e7b5e0395d78ad647100d691ba7ed1bdd0ef4a0c195ae925b8790c14
zb03a282d8108a1e5c0b7e8a8d17b4507eef4759377b6a6adfd3086433c272d05e5bef9fd9edf7e
z8acaa02a9cc88f82fa6a3b136cf0b0b53b089f23ee325b01c627a4e98c619ae45b0cd88901a42e
zd226c94eba58cfde60927d0cd3597402b1541106f2b2e0262494139d375d497f692cc9eb7b1dbe
z6ab3326e1a9d97dbca12a25af789aa15ce75458353ba5346adfe60ce08aaf1d7ac1cd0eaee55c4
z628db1f5eac615fed4d762b93ca1cff50d571c028a7c39fd779270955fd597af1dddac43975aa5
zf5b1d516777b55c1607881828ce49cfea35abe1cb709fa8669c9afc92392232e0a2bc22ad8454d
zd51a884bb2c587ce253286ff969c8f6dc5d65e064cf7d69916da8ef7b65599bc7b53c9678811b7
za21b34b78a80a49c538827950bddbe466a2b1a176fcdbe911bac942c167cbc33f9a5c9c2ae9b14
z2e9147c7eeeb166cbd16d9aa4109ac6eb9d30637e94045a2ac8a77cf27b3dee33befa9ebf36765
z69e3aa859ca97ac57d47f38997120626496d99fadd7ac770be3d560c492c54aa533e62d2b3196c
ze8c1f19af295550bc6988412975d8de72f41057d9d62ca3993967bd75e5268622bcb506aaa92e5
zd5d2b5fded0045c0aacb62d7c4ed571fc7bab1bf531523b977b091998d8bcaca821d530ec0c648
z2c5f1a8e3757bf11bb69f9d531028c1af6dc26440822e55f3cc0cd3a264f85aad0118d2efd7120
z031cabc78a552b1fae2f33cc14cfb1750088924734590a1a2bee3f4087f431a7b9d209f71ac420
z0e4b88caef9bbbdce32bf32d3064e036d686f63b6f3b6aacd37eaf9f1a5d3db570a92502018a28
z8b533691a5d6e5a493e77f18630e86430a65c7a4bdfdfa6959d734f0ce1b8515beeb7bc450c502
z67b3503de2775525c792ad7fbb6890e74f8b93fa044b9d61e83bc7c0cd9032c17275087138d11d
z1d7b8eeac6581d64c3f4492f0a040bdb3d538ea9f1e0c70f0a3c0fd4ffa17b0aa111f0f71858de
zea4b6c0976ee0211e4a4cde486ce8a25980cce19fb72989a30a56257fa0846570d8f87a2e1b200
z2392d7be1893624091ad0ae1cdd3b1513d2ae2e4c8a4527ac93c3d93d9b15791e2e5e9f98f9b01
zce84a623feb666948e8154acde6d7725a40f82501823ef958d8ef3d661b875fc5d9f669eae5e8c
z9d1eed571c7320990cdce1c851e1fdec0829ef353fe33c517bfdfdd18b7ef7b4bf2cb8b8b18ba4
z8797777f9b17d4d7d5367c0bad1d6483f75f2b2ddbccf33a37fd9b772b73810b0f86a65ff6cb78
z59c402b78adff3c40f601dcbec3c29666768ab6b71c294dbce8fbbe172a69cd3993cc37a2bbc4e
z4bd389ed1200cf274a67e311123f570e75ecba8dda3c69576f0174ca207418e0c74c0dc2e71fd9
zc9437f7783b37b09f9c7169e82951065d156da845ae66b1a5ebdbc09edd6d66c5a303e1b8bf01d
z1d5bc04d8e815fac6f422c4e143ac827024b99e3ea7b1a6cd31222da119c8b4f7db2ba7908fcf6
z4ad2142f1daf0f1c17e939d2520649cc95c98bd42d287267118ab39d075a762d22d9ce15fcded8
zb1d9a473d6b8334a401f4768ddcd489c90bf4a127e6de1fced7f6587be4fcbb0e6573329ee3de8
zf770f7e92d2f78cfa3ff08a518d7a73c0d962950f613b6d8332a5c1560b03a38ad9e51f55945d6
z91ae7288ae8e9a20706c406215821a2563f45080e5414ade2f5b2dc2b91f4827e32a9c40dda199
z193620e3840d8d71673aff3ad8e80575d36a588e092cc2e8d90dc66df944483853d50d93248b8d
z176cbacf026eb88131678db5cf4524eb5632c9092f3a3252417f2224ac5b7336aed53a10846a56
z2f301c5a9b39c97b5ad5913c5f5cd2e64662c053bea3d181226b863212038339ed7b303cf5b6a2
zc21152d1adfdc1155efc06cd8a51c0882a93075458bd3ab21c96f51013bada7f4bc01d95b43742
z19feb11566e8afdf362612162a94f279f3e3933d3c047fdbbe41ca69d4327ad03d0689f0b76f4a
zf7d4702919b70adef960d328963a09a6578bf13eda4659630f1cb4bb11ca5449ae399d86dbd380
zf9c3f57a92b4b3ff838f479533d0f4a0874d26cb8708a27420884f1b6edd4023f11072eae4d6a1
z16fb46679c4d02a2e1432150bae5704e5d8405a7c6b047f5b2a0d4de3d1df5dbea1edf0fd3ec12
z32ef509df67e72e9c22d073277b8c7b414ed44f6f27e04abd15d4b3182eb7a6882713d27abffd9
z79a521cb53d73532b055cdef14f1e9c1ee19d7fa2864f1ed135446fadc95625da96a480a116dff
z50693c3392c3a94106ad7488c053cc136023b8a7e46487338fef5632d2646a44710370b3e8fb7e
z457d58ad65c166fa9fdf73c0dc2f67f0bfc1360a97a0776a548d8f2a882ae8b33ef398ee0a8b9c
z9589b6434320aa5058e2c83c1ec6145d82e6deb82e83daa08fbfccec254c97a37b1e6f0dab0c6f
zbb92e87bcbc1086cc2d4a12cf5d60825813586f7e6940f11a73b4363b8ae8be4436bac67e38017
z73d5aea513a7f2a12c0a0e2b888089b60150e1022c7fb4647b474cd6496d36947755de3e67cb3e
z5cb1f192846f26e4c8f1bb23cf8057a7e1d0a063cb75eaca30299705148a08a14695ede07f1afa
zf1cf26eaf5d07c380ec65f82130b4708a64f2064e15d6e431ad3c22d258365f55bcbd3d33644ca
z2386176502c027e3a68a17d10dd57afe2da15dbfa66bc321c5943e19c5b3a3a85e15889ae18577
zf792133f339af05bfa8988dadec41c8bad685b246c3b512f1f212456d41c142f53705e45c78de9
z96ace1eae11e6b9f674ced154db2825004e24d59a482804e37b0fb5a9f16ae5e098fb032750dfe
z3c2279b998b9255038eb90b63306c8cc9ed042a30d450558f7777ce2600a92e736840d38959e3e
z916d02d85d30581cf74aa54edc345e5059198d2064abd2dc4a883435aa349c290bcc8413a50fcd
zb82b7f6389d2e4d5d0d9cffe5e32644f215a10fe2b202ef032efeddba46c3cfa581d8056407edd
z792c1ec1cb8116c69c2d2554dc579654cea18410d5d357e40f1d16a3571475b4c2e07ef6418502
zc1447c8646757915ff36903f742a41feae7aebee72a90fc3f57d308eabe119ec324ce95d6f7992
z7b6c61b0941677215bfebfeb9cd64586af0e84a2197132b95d6228c1d6da9d1192130a9302b2a0
z32369dba4c7cf513ef85d6ce29ebcb3d9530d3107e0623a1e5a0c64ee5f7a8a7f68b6e0217b216
z2f522779f080fd77c11133710bf1b98b8c64131c73e6d1356d90f653ccaef4d629ea8995f5345a
z26dc6ace789112d93a7311aca51f9a3132d004f15b313dea9a87b9798fae09aa00539e19fbfd30
zb75c0790334d8a2ddc2468b16506e48731f1c88269bdef4284eb6c7712f0fff5577cc2560b2763
za273508ee59526792741811cd8fe94d1b18ffa1229e5871f41e64a8098f6c349ff46bb693fb49a
z6b12b1b74ac006b61e049154d9667c51bcefe40ddf97812774fa9aa1d7cca5cba39136ec74eef1
z363257b9c944d617c0ad11dba8d5434badba0ecdbff634c2ab2d0b3651aede7ac88cfef44fb67a
zcd0e4d7f7666ebf38320dd7fe1c29d2dda86957e78b282f0b6fb1f3fa1ed85b6a86e06688fdf6c
z801b837a28fc89fc5902dbbcbd25b5522766edbe1ba94b45f9b5e3beccc251acd81613ea37456a
z3020c0866a63d1b72c29f947af12cc14ba5617b3bbc099497f6842a91a29404286cbd4dadb7d6c
z86990f02d3175c834ca0454769ba21ebe05544f5c4d68e9c1fcd7f109dfd08386907282791739d
z54f1f072f99c0347cee3307a38ba0fd940395bc90545fab5e0c7310c9c32efe002a5934cc55e1e
z238ee00949bb5a58b05dfc428105e7bc425ce05774c8bb6dd0bc845fc07dc7066466abb815da0a
z73b471a42b0e40258d51744f1b9f46f6982b2b6213e924d80074db18dab9c5155d04d87c780d6f
z39ed8bb372c44bcf87bfc4c624e46505a865a40d18f9ec1a1b8346185d224f19b6c629f7f1c552
z48477a9ce779123e2201fc95d9234392d42e94aad26b2cc05e4bf47c719541ba9b1c0ab5f1143f
z6fbd2949599a008bdbd0a18ccec5a2ffb74fc127b8f4d9f508b9c15e1bdbfbf0b1e5a9cca416f5
zf003159f829eb51e06bbc6434ad86060c1f66dae9efcc6043976102e56f4c40a7f167bdbcd21bd
z1344604e05d7fd5ea913da92266f33e4277d0327d455feaa7102e807d473e36b5cc741f13dc6cb
z5380321e902366d9fe48c6986ae8ea4f1268dd9ae2fb90d3b079d5687ef2c6d47ded2ade43e2f1
z0c0534a767abc99271643f17dee20e8f222d528f3a78e00c395f26b30852ceca959e1676af1cb4
z76ffc153df46b8cb77b5a1a1506995ca4679e12ceaa46768408b37ef8a941aeef3e5f43f57d4b0
z25a81cf7bd52055bbd5bee8e8d10b9bd84df1b23447cc71e80eb9eb16ec1cc9573b795ff742ebb
z4cb806ffbf1b047cbe6743201270644ca855b08ed55e4c38290b2892d65ea2b2b1b792c5563716
ze47cf5860b8786a790b95a6ef1b659b7f3a21144baf7e601d1e8cf8ccfa386214b88b493063670
z1a651b613389389e21238d9e29a6d2e0fa3d0e9039a20cbcc394ad54dd291786b6cff6e6604208
z2a072afc3fd40000ba149c9694bd7b4b127807cf6131ac22ea9ae792771def447e1fa3657669a8
z3b6de5dab09a1761f44290e38e859c471c8ed22196b472538fa836194b76026a5836a54fb50c74
ze7d8badb44f0375a3dc59c0b07ddfdbabc8ad72afdeed517067019ba3b4443a9d84b0ce1f66d88
z9cc5b46ff0e290bb18f0312e446284df61197087a768efd5f4b12040d7e4a3ca0f83e89045184f
za6b85b765e5fee736695c8d9b801f44c77112ae1beac2bf714399daa163c7da9ef7fc34d35a5c9
z01924508674be84a9b84f3e0a9156d2987c1f582da5d4da3c7b72e47bec0a3d0e2e736cda4850b
zaaa776db2a936a5f2e22f4e2c17dad8ce868415e3c0e91a3dcc39eb7ad004bb444b5ef0602dd3a
z683f2a705e286f978f5dd4d57c292d1604814d0af1a1916dbb9fb679b5cb8bc0e46872ef56ee15
zf18fd9707ee135d978daf6b81e82b0881b03c76180ac0021f05ded7a4854f7a18963ee4a4a8a17
z4fbf2f99703782628dff93600a47685fa0ef90ebdd8c399b991c772d52eb7d69d39f666f219294
z57bccf588ac1cbda20def7fe632b903a54d3ae4fd6c957c7f2c825c2fbb6dd5ef86dc01b7c0753
z596f9529caa8127acf95962b162771d2a8ce0a2c2e7ba4803e3d87827326e4e112c54faa180ae7
z05241f4c5704c0ccf2d8c3d75d649454c9c1af438fe98ba8e148e91a0b24a3aa3e1727b7b52bdb
z93be4fb58388dbe9b179b3c76ce8593d1f4e4fe542c6b287606e9c10baf2028494d267d889a063
z5d9ad63ee2e2bbdbb9bc17331ec05e92f695b150b634be6c87e9ba75d0bbb492be4aa40f4d1b0e
z88fb3e43f0a76d6363f2bcfd7f1dc041be3d68c62294b4b58c4cc6f964e7c451bb882290144968
zd83768a5bee854f3260f1e49c93905b4ee35f1b1cd3bc65bb85e36656b60ba7db61f547efd27b4
z7bb35a67115ec0956d4a98db74a1ec39f44d41b3cf116aef695d5367a6b09af897d61b66ac1b7c
z4fa2fee111cae73956baf7a9fe8b2bad2365f3cbcd603fce9a485f96472f0bb3d66f0d23770a1c
z378e05a3af9495c25491bf360ae39c6c19d25a36abad50df18d8ff280db8e3db2eb9115cb7846d
zd86b53a6e8119074ad665682455bfdc2e259faee0f4b59d53f93ffcfb3c2c44843696425543c3a
ze9b4bbab092857b3f029286d3281cf35c1c6a294132aa6897a382388ea1231e690867db5971e53
zabdb1b8b78d414757fbb84c7a6d88db4d409e2e2e494447755e2f2a23526861828297374ba3188
zdd712351045cb8883b9a8c304bc9b7503a445f415328a41c97c4f63e48007333ab06f8ec80ff8f
z045414e156a260aa92f12b8f154b0a37dfbed9d586a87a8acedc6b15afc2c688dea858207dd252
z7835b8311c44a1d57ed2bdb2c652c3b7452cfe386c1938e1554b322e18a04d6a68235c3405dfe2
z2aef75081c28c077564bd88cda9d339fafdcf4becdf1ff45cd9464cf55c740d930d31e4d3b46fa
ze19bfa19503646bda8e44b11b29f30ff195af3e4d8d24d23452ca0eba6bf4c6c4ed4c903dc55f8
zf9b607c2bc1f36f79da27bbca10fe8455655578817ea1a8fa693b8af0c527de281dbbee47bbf2c
zb24e21ecb42e0e8bfc75c67ff50b8b6e7c4b4cbb6f9ea3018060f6405fc5c1af2e74722396916f
z66c54fd9e1363d04530da42bdb4a042e41af6ae2c812b0a8d0d1d2cd05afc034693ba63f3ded2b
z22b71ddc984a35b01630cd2f431f0244f24e7039cd7cdd271a37bb0835d45392ba20d28e73d870
zc72c39752402ae07f1226891c5d6fc8538fd36d41ee8057dd38d54b9765bf1d1c0957fef232293
zd2e7f97866edc6dc8e86f1093c8f489d16d90542f920a53a702ee314748d9f3ef466223f7804cb
zceff63bb38be3b4066a99da3baedada64558e4aa559b6302be216d62c5a0932fc6c5ee4e21ca24
z809031cc9c24ddbf0c101a85b1f6aa2e0ae22d4e7b272551fe5f2f69d871cb9ffaad94ac8b9940
z124ac447e0069b07ef3143794792253e642e7f45c076270e28b26eb9c46b3d352b7ad0cbd84ac9
zf65d374ff6810c9bdf1db35083b6413426bde9db344eb19b8624bb813b11925358e91e0a380c5e
z410cb108a90ea002f268129848a7fa4aa48eafd0e6ae13be4a269651563c96f7ea3ec6ae00957f
z8fca76bc6387ff3154857d7584107c96f8e04d2acec7498eac87dff99f0cd97170274ce1f99140
zac80a6842b78b5a8347f59c74a0fc1fd0252ef0900e7777744c3610273af77da95bc0529c9e98e
z28fc864acc281c3aaa8c9d62561637d90a650c0b6b2a72ec4d2dc76261dc439b0a44b95e54dfe7
zdda3086cb8351121af8d99a4b661ef5d235f56b0c1b2f8eca82e237a26da2747bcb207b1cbe4e5
z071a11c540e0f72acfb54baf8d9655111ff079e2951bc52d65cc56e6dc31be5865398bae105ceb
zaf5bebb6862fb8da735e1a4ebeca7d0b2ef81f1585d57464fbce271201284d55e4cd3bb1b40bb9
ze5a075f36163e894005ffbe44f7c52a669f1541df5785aaa923af65f770ba5d192c92d4b1e9c0e
za2354e7cb9026a8defa74033e371a1b2583018bd0e83f30db9ebca8173b5ab58fa4c7b0e91b341
z7497601eb44471d4196a2cb13725d2ac4dabd0dd1d0adb38ff978677d8325287b24a226eb5de79
z229ff0654f4435f1970bd404f486454aff795ca0572306729d5a36d21014b7859898cd0cfa9369
zd3483d481cf1d467c2f965672ccae2a9bec3f752d48aa9a692ccb6f68a2fc24d38a8af262ac07d
z2c071d336f819ece7e0c5eb29832c6dc6700c452a63ab35ce6962ae5b4e864a5838e5d8642e7b2
z22ef04fb4db742b45702cb3ce2f84cfe34d43de1a8c4f5104457b1a575b1984815b879b180132e
zf35b2dbbb64c0bef591fe3dbdb31d6e46b619b9180d370f11727b132420e1a218b237b11c0ca35
z1b1f4884b0d6632cae03323c5b1b91391f11e52630f60e10a914d909b041adb459007fd93527fd
zc587d64ede16645bbf19736d5516e1b827c137b58098f3742f443afa5ed969bd113f1a6ab42b19
z0d9017d0e8aa2d20cfd0f1e7fb666f2b5740a2de0424ee0e14924bb40dfdd8a2df590ab1c7c368
z0dfb82793d0a7ddef167322976123b693a8188848acd6efbac37448a33598fb57125957c18c65f
z0244a18966a21cace1c8c357efe7f1bd0f4be4938e60ae982f05a4fe75f291e7bcffe1ae66e126
z5fa1c4c17d76e20e0eb20ff68331eb205d6f7985041be90883bf5ad5bf7e5e191c4171d4523ce1
zc1797f8c9fbe84627c58a26c998ffa429a44891a0fa18b35fa87159681ac93a2d85a181833f216
zba173e4d8417e93ad607111faf527cc8609ef10107c58003ab265339146a8319d820ab3b7b3db1
z0484b8b4cbb37793b0364bc634316e4737e9418592ba58bfd7c73685fbb00379340e67ca6afef0
z20b8bfb3b2b091ae5c0bbc905f815e1393f497715db31ce0b1be5d6c3295d4f8174624bdc02c20
z8089bc3d566090f10cac78b166ad6c9baebd90f97594e0c5be3831029da083f3da07b10127e079
z326ef03fd26153bb4050ca0fbfd3583f4bf33713048a0d64cca72d92d02674e7dfdf5aec191416
z1f9ba168727789109e50a19adbdeac07ea10e50abfa9269c56254d55af5397158af85050eb7002
z7f2f6445a3803ec3347fb2ca8e4ba8d0c93e57254d155f2b366bd86b99369a8688a1df7f1437b4
z9958fb0b21cbff67e71734c8008c6e9917e10e8d7ec76f492ab90a73e4012c807d8fc730b8c487
z876b0f36c1918995557aa7eaac11b22f3c3309d5e962cddb65854cde638fc5123feea65cc77aa8
z829a4a199a0a55c3aa66534d670445501e842dd91d756a4cbf172aa35c607113bb07e10f54d2d3
z5cd64a8684955cca6560f064d88ef19d27efc193bc5da1a8b6dd4fc56f32b8372e1f5b03c37478
z9ff7ccc4629e8b8b07db78f1daa0389085861e39220f85c6c5d991968dec65c83cae66901ccb0a
z16fed050a6eaa8696532feee8d6e3571461d1b57988ac2e51cd67977ded6c419eaf458ecb7558c
z7efcbb2bc77f10aab523c718371812b9a23817b701e4691400b114443cd8cf318a98a545785c83
z6704f7308e0a896e9429800fbfec11dfa1dc6ef51f129a15044c07eb76b2e166a21942219ec160
z4255a1047b66438bca256de801c350b40b4cdab92fb627a1ed2578f95620f09b585679c1418709
zde02b0b349c1f748fe069cb7932eb52b3aba7afd3e2b57bf2d8282b1d413f16a994be7f675464f
zda252d7192543e72a863572fe806a5434e8dec37456f463acb27bca0973bd7a2156bf114b63a93
z637b125013cc2dca38ec74f73a15f919a38a84db4b90889a78fbf5d7e7ec05b7ea1a8b0f25ede4
zd289ed2f438640ae615af72ba4818592f326f0e3f63d1a50aad9ab87d4c175ae5031f2b85bd7ec
z1d9f9959979f75c250fb32655a4af3686859a4b1b94b8a5ecb16f506a131ab62ed50e9e8789ed4
za34de40b192d9c466692751f4bd55c44eb5cd4cf5dfa8ba989d114510f1c3675de822dcc6b9019
z0259cbf6b454eb36dbc0d442d375358f02b02d43ff60369d76f21e24ebec5a247d439b7f140b3f
z781ed4342bec46a25701cfab5d4a19c51f520cc75697a093534beb4a67f8be41b5810c4425497e
z222f5c6b7d998f1b5f09905c03fd074105345ba6b605b9b7893cf7f99be0e2a05229fe498fb50c
zebc551087fc323dce135a29bf6e76177d3c1a94183b110a38e58451d32601772b1012d694ea532
z1feb5204304bfd3674658c95fea30fa98f615f86e697c81219df98823eb1d4ea424c5c46ec95f5
z0782ee95de0a4deee2c176f226b3a30e52d47ca5c4888883d42b1d46f7eba447c28cf1efe766c2
z6f29cb50a5d5940696ba434d327e819103ed7bb8b3a317af998bbff14a4bc761dad4ca750adf2a
z183d75baa54684dcc0304bd2021418b11652f2335e8251b1b247940b4b88d16cd943c910ad1540
z19a9256c43ba75522948d40aa9f6d11409be8bef4fee7ff592ce1a5f01d67b81da1db7b4aa0512
z3ec60a57f7962feba0d9e3a0ee36663cee8a66ffc19d3b6610c8030bd746ccaba25bdf38cd50bc
z4691d022239508c5c1e05d0a534db0fe66cfd5efc15f984661dbc7d2a2b0752e00d1a55d2d6408
zc8e2636a920ef8e73366448b0867bc18632a1673a0391b0c00992cfe6368cb8d259eecf43ee03e
zaa4bcd74f05a971ae37fc2be5be6d319694b71461f6ef144da114c51287472b1b3d7f4704e0792
za191d78c25dbb6fe02ae08bccb5fedb20ce2e0e2ed1bddc1436639692f95e77fe2ea45b0fbaae8
z8d70a2a59e03b45254766f6155c87b96c6181a5e98601730ca6cd60c301c16838182676f5a0eb2
zc496f9432b4dd0ae1235f25a44ab8003fc0c7d5d2e702181f4e91cb7c5eb70aef98ee9b8dbd415
z55f1f410d235d60cd4466b3958c2fd02923fee469e18ce70d1ab9446f34ed459d34c89d5653ffc
z8350feb9343e2a8b04ebec4f74f2c0f854815c93908ef892e5f4a34c32d526df1f643830c3a656
z87d249d64f0e439673892476401781a871457e85a05de4c83bba37cf955b4b0445a3c0ae8d729f
z0d0b7b7fa6b2247bc4ae3dbb82ea70fed1e1ac68378c883863b3614d772ee39c8624c37fd14b03
zccb7dbfda92d870acd9eebcde94e355ec0e735e35a058dd16d8b3cffc8dddb24cfb12a0f2d3e9a
z7d0f059dbaa05d940fefd82d8e5a6eec4dc3c2c30543ba17c82eae706bfe31bbe868f391bc7095
z7189254f94707d2e44ae60a95999a035cda0cd697ed2ec653a1cb5658ea773a9fef739e20b9eed
z1a635577ce4d0811b5a13302e85fff1fe87c4343dff7ca5f3a34bbce4dc205df6d7e4f35c1ba6f
zfd1700e406542a514c468ba25265cb0a17c438c1882ee64120e5e5219785b185964cc48f4b3c4e
zf6510bee2b774c595003e82fe47c2d3236c1f9491d4e81d9c6331d18084a186f85c6e3aa7b7395
zb6b9ae1d926d55c0d8fad209500efc495106c4a2932c0b79f8d3704f0bc2196b95088612d457c7
z5ff3fe6f973cf8627887d7a516773bacbc650e4e84a5cb4cd3902f78a85707af91ae2501dca737
z5d4944f0d17d5f16c3a5db0f4dfec68aeacb4eff09e190437a0767573e843327a6690e914797bf
zdb91967afe28fa536627c353440bae065718f7617531078d5753398e095790c316f7253c0f2793
zfc9edaa6326558fdb796a809602b00f230a940a414c118957328abaae07505249eaee7b01bb2e9
z403bac750889bff5b52b8beeb3b39e06fbe8f82eb68dc619bceb7ffdbbded950f9a265fec3d2d3
z71a12b67671504891ac1e8111aa7902bd18e0e2f79371bfcbda18eaee86931244d38a7c63394b4
z59bc6f6ad0097205566f8e32ddfa77a3396fc8ba0daa2c31815994e8de335caadb84bf3fd8e56c
z86e61439f84305a0f7ed2f65a3f241b3da45218702591c0ff3da8c11bc8499c10275aa668f7f4f
z540783d30812baeca56007cd75a42b1ea42236916828fe6a0a5a927783a72c438e29f40b7042d1
z7fb13b8437ad91b31a7b15991a9e3e29cd9851187bc05098075f9f783f1302b184e24968be11dd
z2587e29bb90c0835280f25f7457bb4844242a45aa36f571a185fc3059195a7193c0fda1639c011
zdf0401fcaee67e4780f39d15cd31aa7d30efff4c6a49bcb2521992ddf86e2200ec7a9e8a1bfdec
zdbb0ae30c9acdc48a7237125fac53d07b60455ee139e2b2f4e7859257d6d09754e489b6d3dc6be
z55213efbf5cd0e80e2b35f6b41debb3cc9f0f00ad4cac8ad9079fd83137d0fda91526968cdc8ea
z5c32c1b129893145f74ce04c05e9b3a4fbfb60b4a8c5d783b017a368b92a0c49b5f9b285ed58ef
zadaf917d0850cacd57fce77e00893a5a173b2a6ee3389bc959083bd2986483629a5abca2a2d6b5
z5da778a768d304025f07526ab002af94819b5bba4ce6e70b990a42a7e49cac71f0b29eded2d679
zfdfd84fb00d43c5c664c363c487909c90fb477cb279536582aacdcb4b696e59a5f7fc4e9310c43
z989a566797283f400e07c9c83683a688bee5bd6e1ac3938ecc58fe5f5f2664b58b983db8f93e1f
z0791a6257111c3ee17ce2b545d0ac70d2f52ff67577ad4d12da800b00eda73695bf327abc9a2df
z7ce0c95534f5a6512ec24761982daf5b485364719e0c9f3b95b71cd7a9c461f23f33d238f1a743
zeed448cfde7dac7744fa32d176a121a022c9ce219dbe28516a4964f4bd69eb92d61954e25d1886
z8c5a7bea78c3a4629b0127c1ab916a6ec9c2cb31781cb4c6f874b46bf3fd34ea13bd3c413a6bd2
z49f33cfc9504c8b9f692c3fb7a94a398ac271d1e88db4047ce42bb9e6e9c1952385dad306f36ec
z1de3bbe7b7a49e3d8fb9d3d700caf0e284df68bdefc89257741f7e158f522fdcb56c939e1b1745
zf700d57c112445334ae7ac69a0128b3a643e608ef92caa12352d7e8a0b46ecf09b9e1711b28b2a
zd82fb3decc04cd1e01a554c634e806f3e55f4e093082634e62a9a32c0591e8171d80c8ac41f3e4
z84a09aa69e592e2062b32398ed19a26fdd3741c96ec44e4af59be539ded5951475addc8b64ee0b
z8d9a5c9fc5bb05b04dcd3737914da5fd0d660f363c41b9885573ba2647535e6d1da11cbf3b1b3e
z0007bf4cb127b75182c86f0c0feb031dffb90f6f7050f7aa4fa36fcdfe9bce98f9621a0fa7918e
z4f851abdfe3664ad315bb65891ac3d1be131be6196e8f2d9062e79a3cc33492bf9a76026afa08f
zca73272f4eeaa88b96a8a4ff0976928227d0520a01c9d1252a5613ff36f6875774cf545b1dc23c
zdc4605962a461fb77e1860bc23067e72d12f53d3eb4a63a2ab34a9cfe566ebe246b435d6a58dc4
zbb3dcf978208c5928c99382b06894b34de6d91ec43c10984faed411db9c9ccfc6170723c0af1a5
z3ca4815df5b45b92a09c0a8ca547b6cbbfbcf1cf803138ed58b40f24339841e4487fdb989e3d80
z166f3c8754b01109a5006012293035ff80ef5fb13e001290e4452de31e826f59cc2a39892a8945
z193000b03198e06908a90700f993dbdd51c4c2ce08f6eceae35cab3395bf470727a04b339a27d9
zfb38cbd004a18022b6d7bcfe4e311483f247b69e5d17d1f3dfa6ecb48a19f67f2758cc4d404deb
z8bbca579f2b720365aa7dde8d1d3ccc6a61b008aca1fc986fe03a3431cbc4671903cd6fc1772e1
z121b4552f1f11f0d32ce8bdc164976c11285eea8ebdda1ef448bbd152569e20db43b76cb5658c5
z5ad03a3faa37e109abf0f3b7a39778e656ce5f8f5889ce38787577d69366caf0d433a948745ade
zf70c3512510bab4721187e51b634e27fc0f9e2c988c26821b6dd31491bf29da6e5a6b31ed6a0a7
z46a067d20164a33973e748857163a3e5402249870cd2a567ae0623544771766402a27421744c39
z46841e82a6476516561aa82acb6658c2b2ee483c67411a9747a59396fb0f33323a002902df7a80
z0436dba24464b9b23ca98775da535dfff8d7c3bdb958f2d10b1719bba1d596cb156e0072d901eb
zba99f44514d2e91e5d6ba82a07174b238e6c523256fd8e21ce3cb23ed7860e082a9c836b9d3cd4
z2a1aeb9eae0243a385cfabc3b8f089d1fa49fdb757dd7802a74ba8a469aad51cd63194122b0ada
zbec3b29a9624412ef629a5b89d0896fda0199f32f998dce394323b018ff31d30d512edfb9a70a9
zc18ddc4d5fc92dc9799c124ea73296c57161d05c34ff3310818f776ddd8a86a00126483cb9929b
zc0b2e0d99bf16b8a143ee49d1bc36ea388e336293747c38bb4456b2af0380ff6f66f6fcea787b1
z793b95456cc6e931c1f390275113ac27b22582522b234779dbdad76626bd3aba198867f7cf2991
zfdb444e4c1dfafeef24d5fb518608f5ed35e16470f6d0a7bb48a6d803cfaf286a523808015616c
z8e4866e61b0bc09858ea396e2ac9a4e6d3bd905093bb3e6b186f02db4e20812cab8601ee400306
zac80f2b9db7fd1ea7e3f80b1f31a5073a86003d937f4af9c7a1898fa63673541b4175c50fa4a58
z7c03770f88051efe74eb9facba9ed7be63f574566de74d10d6b598e53e96fc19a7ec9f2b7df417
zf03c9f57e170599a8cd1dde83fd9df523287ac4b01a6f4598adf6d53f86a09c455e77a9741c88f
z911ab5afb6e3abd4460d6f903d20fe9807ceb1fcd49920cba953d9b07d405758a1d7dbf6caa050
z5d8e45a971b143f7440abdd50c308b562ccb9997bdeda5a01e3bbc7cd9d2a6921d3a5d63e8dd16
z0d5ac9db391fd1f72535de980ffecdd69835ce398d6f503c38ae2a584d418600586628f813e524
z7b61cf04b30491394ba862d87607e1cbdcff573bb415b46bacbea9b9bdd5d7c44a2def0de332f1
zafc3a271fd9c56e6cc058d425fde9d6be73a81629c14e17b619dd91230666542426b40d146adfc
z815fef39855d976f6e62a35069d8759b6b30c8e8e4fba6981a7d9ec83786509e6afaa87da621d5
z719ed0287addef4202ca593e1d524d88bcd0d2a7d2716acbc774a6b16161b1b7bcbad40858b7c3
zd223064ce5df461d9aadf4fff8857b703285bd428e8cea336f0b29efa7d0c6fc1bc65d231906eb
z6fd2fbdac7e24867df413dd2f06a5388693b2ac9521e6fb3c030bc923b2c573d04459785255121
z62b6bc0cebe54af0d1800147113ff379384017efe0e2725a615f14e58e7a9de42ba7ef738a321f
z99b1cb027e441251ea63e6c0a908fff8e31da9e24c32b47b15bed98e20ce728e206fd5432705f6
z4504c5b7025d5e1dffac6cf0e74ce65d45768bc4b9f56b3c3ad44ea2f65ec0e7c3b6e136408620
z59f792c439b3eb92e5b30eee5842f3a9976981502a54c26590f338992f46dba450069ea3fc7d78
z476745218197b5624b5f4140d04f0322c4d8e34de66b22111a94ef095bdcad6934ae1e8e3f3266
za4e4c533cff923dac275cc5bfac19feef010907b31a27e9733028123415760629645bee36b59fc
z610aad8e96d72517264e2f99a2b16f6f142b763d1ce9b7f86ad2bf52b88acd3f3a2c1d69b5307b
z4610efecd2301f9deb8064596a770686c907554e1d71a8b8cd54b4f6f09c41b4fccaa8322270cf
z079728aa3b07083d129f7c6ec3eca01843f6f0a3830659362b01488a5bcd59bdfeef54895f28af
z6f1a23a09379da0eb1ab7ecbb48ebdac22a6e2ea7e3ed24daea05bf2ef4a8d418bb062d8dcb7f5
z585bf595b50c1d8e3d55f1e941b7ca801cd9e27853b5c84ffb0709e9e83b81ecc885d3d597c257
zb15abb26cc6625ddefc836e303cfc66176a5a4899fbc66bace253c815a812d7fc9128fd0b0c96d
z008f2782d00f47fe03665e5c4a9bacb3aa3daa366eb5e8d287734652073e01d57ba94bd6105727
zd3fd54f8eb4b4181d7210bc14ae00cddd458c576340ab4e05acfb95766a11d292ea52a3e35afbe
z348aa4746cd7799651c95cebb08b69745f96e154bb464dd23ea7a29581393fe88a3a2abc1d74bf
z9a17877315fbbb0090e4a8be32d6c8fac855f18d50d9175fa97a5011daee9df6222bd02452bed4
zd7f2052d795a8058e125d77a6b7cc882185da80baa88ba5420c25e0c6391baf076e811bd3a37ea
z2e54a261d8f3d69514d709f01dce36c4dfdf8f23e3829f1729f6958c343d6e9c793c4040afb7fd
zf0094e95185e703513e31d7dc66fee347b3ccf1fdc7e8ea9d31f20890621ec1521d58f6c8cb365
zd6501d64fbaabb024c3eaa048df5d5777940aa1f9f4fe43adbb5a70d82ca8d6d35d6a60dfc75b7
z82ddf78c94b45d19b0ed306afafd1db0daa4e16b4984c6ea7f4e087c692a6fd42e4d8e75e36a0d
z6177105b4e1421b91ac1316ea2a3d0e0c979c006e8259d17dfca8e2872e7c51b8a7b7d4d79a25f
z0aeab93df77d58c75598768f4a63116a7f61a7f19d12430c1454237d2e51996010b8e963b0cc7a
z61ec2e9effa6478c359b3f924ffbabd6b63b3a83e4f63f87ad2d4fded539d5ea225e96e24400e4
z2e3004b2de6eefe7d8d882f49bfa23c8af655f79c4e1989e1db793ca8dc7fc40695968542ed94e
zac8b245c9e3a75cfc84ae16c5dccbf8dc49eb835497a476ff180531fa3b5e16c966dc4241d3e44
zd3dc2a298954dea1571c4324e62ed3182bc67a88dc79ef6b07f7139fabbfb9e0249cf3c61b2fbc
z7bfc736053bf8746172240f9f34355139e8ab3c7bd19401119e5c79916bb6b7649c59f16699e57
za1d03994d29b1e8d2461e891ed832bdaeb26dcbb8df369e025794eab1c4d29b9624c235596172f
za56f9d2aea6ac37e0d761fcf999266ee2ad1f84980529bc005e1d6b49976a4b19775ff33f17a8d
z1cc2d1e469093d2e8c2a046bdcdf1ba98961df699057167bfaefa3126ace27da9696be15a27fa5
z0833f11f292a851bdd902490b8ee52f2086b23a4560cc26f2cb12689a19ff0f28fd78174d792af
za49d43e3c8f25a6b503b3e1eb178217b9a085ea20fd7628021890aa0fcb08f219ceec712be3ad4
ze0cb369e6957379a81c8a4752645a1c17293aca5b7c2c9d519b3c596cda8e61f0e2eef41cd5cc9
zaee053ee3d48875fc2729988b9009b66d301e1c95674dc3ff423f8229f3ead42ef67350d53f5bb
za2dd58c2ccda3b99c082ae63d53a69192b678b56ff1e33261178f383d0cca18abda6b97ef8687e
z89717ade8e65e2a70676082999c520a7ce5447a3e91b349f17b401b0b05a977aefdc1f477e8fd7
z0f02bf26088052fa680a730746f22dea7088200a4760fa233a4269611e9136a822be17cb39b842
z2abb785a5a0d471c0d450dea663f3b90f325432526bc39cc8af3d1c3bf6a019a4b101225c75e7e
z7c1067b978178183ee871266cd329028e3b859ceeebcab46821bbb6afc7a65664f4e2bf9f08b5f
z1fe1c13a0a853db9855bf52517d4bfc2100de0767b38121bed89e58a79c2a707a86f493270652b
zfbfa52b52f4dc895775c72c2c83dea43b088b5631ee6ec726922f3d707a03f146640cd85d9e568
z43392b295faaa0482d1724d322c744aa618c8e5607606333a6743835d3438538403c187cdbd869
zcb38ad94340d986bbbb2518c2794594db05e91c64091de9a3974144fdbff8d849c10e4cf889fb4
zcaad8fceee4263cce779f48ab4362a14d27ce7066a6e441e7d6af756a665540a958551bab4dfed
z0c0519c0c2c8e6a36217d568a3b6240f10d02d5383cf6481a5e4bf2e9e1d17dc9c262c8d5afbeb
zf7ed54103cfc82c0861a3a495f9a6f57a1da297b5a54f12a86462bf2eedde4189fd1aaa2c921ee
zdb6cbc562aaaef2bb51df03d50b329e2f3fb43fcadad42e223cc4c3539e3902596dcc18a68a416
zab225790af24c9c51fb8ef2fd5841088dbd85f20c63546cc1020abadb4126220a3a91b81c07b7d
z417dd097697c8ff81d894987125bf377f30c254d4d0eaa62ebed53bb6b99900234b6afdff89e99
z7e2ef9e5ed12f5dbfb9468c310d88a8d788f8b1fccd2e5dddaefb9a2bd5e1bae9eda9afc601dc3
z8a1862a9ac9163c2f8e3b57241b083fb3a8c3a4c65d9842870c20a156d82a08215e63f3477bdaf
zc1de87f708a676aba753e40f8d3fb20c709ca9b6b33616cd6fb2ccb63f71130396592ceeb1f6b5
z1c71502d2d43a534d9058702250fdaee37c0c36e5c105c7fa30c8bf4b9c26e56857e959dcc4325
zc73e5acfe0f99d6e1c3e877621f31bb3bfbf92285d10d46d8d52075b43a89941ba516a1433f062
z7ddc4af7f5a4c51c57d86b6ff17d5975ddb9b692766c0c97b8226e51fe5db748867c482044865a
z6ab364041a2f04cd165751f72bb1432d55f4992c7ee31e8fbccc9830a52be6802175eae1683799
zfcb5bc8ef2abd04b2ee6dd0f4100baa837f9211fce9c6eea2960e53548e1f73e50396e575cd448
zdd6883f07687bda28523b82c850c125e06960703f65eab2e029c63464e27b43748ca5a950cc121
zac3d3a1971fa6e65915f8a90880a56377b90f566f6f078b479eb4ed1dc06e04a7fa473b4d2ef3a
ze33fd56f93b19f5cd1c67f3184f39609e9d19bf11686a02bdf5c499bb41fd4a1c37c4271b66900
zb8da1e4eba5930b5b4396c6a07daf65f9400009e2cd90e2e1108612d4a3ca153332cd66eb18e39
z4b02bdaad822f3a22eff048c839f445056ccc154a5ebe9b03ee615228b4aa655174a3b3517cada
zb3b879fd395a93d37111a998901fe93a73ab1be681d8f01320d7be33b67b9758f868db81b9d99c
z641a2f38e20f5f552954015c8556fdec2f3895bd82d89e9aeb118db326228c158e7f0c9f108d0b
z3dd5485386ff5c16aa381a6b6739aca6e848567059b74be17ad8d62f7c9cb802505d0ce95923b1
z964d8189391f9fc1b1e058c92dd7c43eb2ccbbb7edf0cea162296b2eb38ec986e5c76f635d8070
ze3cbf9a2ca6dc1732067cc59ab8b0dd678f720f547d9b8d28e4a94eac38730a5d912d672768fef
zcc428350ed0e82d6cfb921e22b47ae38cf8532722d5a51f7df26586653fe789c3f8753b7458891
zd2ab480576dd2d5ad223bce1362e9d0fba71424f3ed7d773df30dc99ea662d807d99a74279cbfe
z6047e4e0e4e5368c7ec5583771650ddc0e370fabcb2e055dbd8dec62c782c182307f25b46533cf
z07e45c82bb752a9fc33d2f61366016ebce8c82fd6fc81454f32c1bb7122e8eb08fee893ca4a7bb
z19df5cc43b83c2bcd815b62b722702f127fd9b618a839cdeec813dbf1d73d3d9047b684667867b
z91fdb6e211ece154f4c23ba61ac381169021b14a05edebce8cf3d68617c0841d40550476818994
z50cf9f78a0aab4b5c9794dc87436336dcef5b46bd47fc4a031330b18909623644a4343a862cc34
za7dabf74de9009ef9a015fac072002b42d8fb61000c8fac39b93c437388e2a0eb3f62335cc3a98
zf7307cbef0598026eab13682410a41183e6797b93195dee09c84c91894fb22c95b5161cf7ad3ba
zb06a466915bd259d71994e8dbba7df4ba811fbec138fe3b3fc96fc1b14f8faf2ba39e568bf3560
zfba37aaf236dcbf39ad9c979b0366d85bfb5b8f3e6f1ac1ba1e08f45444f1079ee9076efd00884
zfe21843fe1e2599c886b9c427a78fe49c9123218d19198c31cdd69707a93e34987f4052014cd5b
z767a22a5b7ad80feb292e3389082d5430ff78c5bdfe92fe74116919cd2dbd17277db6e994cb419
zc0d3e77fe72089dccf1c0d1ac0eb5976eb8fe364cc37f8d013919a79d5b25e0e7e1ab5728b218e
z5d9fd0bf6b9f8bd39ffb0f6599bd19c6b2e8b023f257a8ac534eb57fea26e741037b8a40b18ac9
zc2d47c7ead4a373b4b97f8e2b33ff6e41373fd677ea4aa60de7c956f639c54036c402b227398c7
zadda3eb2c53a362ba9d2cc9ae62131c2a7304ab39e4fe0fd4840ccf10a135447a8816d02a7f903
z5f9c9916544bfb30aa8697e142ea2e335b047bdebabf95165f1bfd23a7dcd65b49cb49bed173d1
z6b28f7274be361d533ffbd9a7d8b5054d2f406da4b1c48d3c5df26cb31fa39e7fe5681983b590a
zed9a47aefe676eee2a9f87b5b0e224cce409edc454e9aefe8c5ca41b9ee20e8ebb74ba22d925ab
z69d8c83221c2191139b41234f3ab444e9f822df76cac3ffa7e448860ca69716e3a5fde4ff195e7
z48726fc084c0a1054b38a1f3c80a9de998ca4e7a13bc711f3e59e5a71856dd849680a1d550898c
z8be22d9fff4bb67bc2e9759a21ceb798503f8e00dd543c96d9439cf92d152a5e287e55a210b366
z05b7cb4ecfa47795b7da9bfa0a452476a4ba36271b14c4168060d130ae68603e92e89c8e05afbb
zdf6e0c5e16ca6f347bd5da601ff7b1aded4524dac500936a943c2a767cc2da749ad3dde244f511
z9e27a1c3d6e787da3e0cd4af46cd9aced2158bfa7776f26ecfc3c339792017b101f150c1fff63e
za2a85b6906170aaf04f11a578033461c3b0db89e3d03b3e6503f70a6d03fbd5ca8820760cd4907
z967a8173648766efa1ac950586c23f9a6de8f4b3ad8aaf526d0bfb80068d1b3e4ee58fcb900105
ze8a2ddd2eefd741729f9bba024e81af10668431fa20fb9cabf82f3ada3d3d9842143bf40b98594
z1b3771fd7ee3a7189d1c9bd3caf6684e2a406d16cc307796263117c2d05d42d1ce5ed3290fd3e7
ze08a5d73b1a6ff7515a5790dc14105905a60ee6201533a4aa49526f86c9d4ebe01cc253aa73697
zdb33ba2b0f3781ce039d9c8798b4d41dda120fb11512c3a03961cb6ab4a72914d573c73e342b23
z7420f0c115315a81fc0a5d884f7417da94db6ae9fb267bbfcbfc50e5b8167091d5e1347daea6d6
zba1d16392ed5d9017b03948b238b26d6ab5601c7045cc65c891b1c0b65a50216fdc0798f8028ca
z4acd1826720cd56261b79a963f30cd36cbaa272ba79a061ff5877558092445ee5076badd2f4c94
z5d7ca96eae0ae5dab7a313e0413b46eb0946d7377dd351bd4f31463baeb748c7fe0695a2f211af
z8b17d9044eec5909fd0f3223042a0b3c3ba4f6cb98db3e718b863dc78ee231f9fe30b00120484e
z5d137b23510e558c7f60dad8bf41761ad4592f90c314d6a302c9ac8350a4ab4406ce77f7b569b2
z3b4d9be1b1d879b351698ff58ea780729ec57c4163e5ff2c52f412f8fd67b70f74e9fd665f984f
z4a49823fc37afdcd7a16e788f0595695265a51791cc808cb79bf463af2fb127bbd4f49c534728b
zda3b1c6c7e66e3b1c8ee749cf26e90b83e268246b2642e7048567c4edf7d6864afcf1e1b3554d5
zfd7d5a2ff060d3e8f9ef2ec9257b0550acccd23f817669d7640840356758eb255d5fc7a06903c4
zb278428484d7f3e590cf63aecb5cf0bf2274c882a06173614736e55f3ffb4f5f5f6bea14860fa4
zba6d26752ca27d5ef108e28442625b1095a13328cf594f74404cc254a41a9977d6094e8ff907b4
z8b32ffbc351652d63e3c1fa00065d1d9b4d6a512487756d5fe5467bee5fe67609c29761a559071
z8c83c611377e24832417e06828cc6ae57912a9ed1495109ff59fcf7188633aa8d0c154cc5fb946
z4698fd701a0f39f451aeda46a1199ab6204175cd01ee28fbe884deea051e46e0ca3f1725fbc70e
z5f90e1f8e344514a57b6240ca1285995f04bf427c6fedc3f07e5b4ca82652b287107d2d33f3c7c
zfdafc3f521c745983aa1a206a415514772f3c40ff921dacb8b6523429bd39091b502069a0284d4
z01477be4b3a58817cc954eec31556d44568483e3cfd78f13493e599618adcf56648561d428389d
z27f73ae47d66349fc962f4e9393a6db22e31562e6ba7a20824f7b67abae2a2fe69bfdcfe302a20
z5534b22b498efc3ee138866c1d24f59f724f7f54d249dc2d5278f4ba2dd7cd45ab48f736cc3baf
z96a75cb64654374e63e82f940bb711db4c63184638152cdacdfcf0ec77e76e80997549a7570075
z2ed14ca66a105e76bfed39db2dd7536a267f34dc8251780301d532016581ab450763197a1d3ce7
z4259a201c608ee4d4eed2e22d8b0bd344d171e994b6ce06a36c66ee8d9883c7f30a249d9d40d31
ze1cf54bf39cd1fb23245fb32fd5ff911feca371c4c0bae851f0b95a983fe564997308ce90cc819
z487d6ae6ef7c27e4bba0763281b2ea28b44a5e213c14d1fdc80061c57daea7fc4338d285399ca9
zaaad031a19a5cd6b154901babe97ebd9afb70aabf13f33ff112fa872a662dba09a78b4a5b1f7c9
z9e5c8c7d4eea6480e19d032353bb8659cd1738d8160cb8305b1ec9f25f29f61ecca869b81475c0
za558d3f4850564134134fb9aaaef3fbc2a4a997d41388b85af9e40f3f87993e738eee14edea4f8
z3ae48b0e3e174514f12f4d9c6e15c9eb426af7be8a66f6a5b6384431bf5c39b544c746414cbb2d
zf0cf57bcc56f8227bed1055e1bfcdb4a93140fefe8b9e25d76f2ffcb044ea0566c69d749be0fcf
zb955d7632fe5ee033b3ca49137b2b33c16de1f91bea67e2ee532c423dcf2ed57958f7ac2dcea6f
z28cf6d7871c8cf808f3b0db3fad0ec62abd204554959ef2a4ec05c989d156987aa5fddcf3ac848
z97aa8940dcac1835dcf19448ce7a1cfa9dc01d53449cf9b6c665d41602ca76a29a60acbdeeaec5
z97b18afe124e9d605d1154e2d6fc3304b4871fd73d28a9ee1c706e4af96f47913a296b5fdf9ace
z88375cd230db50e955091f0d49573227e0432b0228cfd1a6c562a228cef99d3857442f04f03a82
zfa956c1b8d51c84bc23a641b3ffd3677981e3cfd9a26f1cc597e3a3f71f4db9e900eb175138be3
z995c20e44bf46cf0df602b137495f682177472dabea2ccf6568e5da074119bf27c149ffeb6ebda
zd7921f816f9e862bae022f6d10a592694751161c83b1bc481f8997c019b4819ddd8877c93289ad
z921ffa95898d9bc60a1f95cdebe9c0395369edd34b98d6c01264c3aa7957acc4d7957b9401cbe9
zbe85aef3923be0563cd6501cbe0627d40cf6e7a045db1dc214178845f4eda45ecc44bf9eb67658
z8f512434d75d1b61e1de4551261e538fca5cce6aeda4b46786f54b7a50c26fc01b38fe11a8e6f3
ze9836e984fcfb103e303ed151752b6f67d0bc5232ace123091e666bb179b6781f5dbf917a1b1be
z96ec602246f7df7c97d9c38edf050381e4f8b1534d6ce4c4af8b30a5c8256be1206bd0f4b0004b
zaffc219636cc578d0a195c57380a34c163e76e70f586c67ea533fff94162ca45c5042e1b51b22a
z99a5503b9b7e310cfa1090ac1f5c23ab3960d83e07d72ee9fed4be47c44fdf48f66ad478c86758
z5b9c1b2cd5cb377e7d774b6e1d1b8a7efbf7be9ecc7920ecb9e4b1965fbfeac151115d13cdfe02
zcbdf9abe4f3bdaa6f57a2ed87aacf5af9f43b2cf5bbfb7c175855e866ae007d319f3b835c49172
zac246d5241c024f51cd22e40891fcc633554095e6f91fd7c231e31471159a4208eabd57ab9b7b7
zd1e68be4439dfd93460f446b4244714831bb0505fb5a77cb8fbb040e94b013c014a9aefea12603
z6182da176af22ef2d6084d5e4d6e7c7dec006d324ac38a4dfd33c3fbde07a8d1cb521c9f7f3b8d
zac414be373e4b96372c6e77b8bbcb3ad81ca40c6dfbba95a425d21e3b3ce1f5e8a33a625bb7652
zd8c223f570434cc915927061682d26806504b194a1e65f3bb4c3378318fb6cf6632638b2f463ed
z874293178b65918cff89bfc3d6327824cf6a9a00bae572bddf7604f2ed2d87de3b1a76d325b019
z1e9ef874da49930004c4f1900f39be1de9003af49b41bc2d073cbb4f284244cb99931ebb7aae61
zee979094af1d5af9bead40339ec81a3b273f813c6e06ffc071d456f6f33366e1f243315b4c39cb
z34d18bdcbaddf94bd065d6e3db1b3d716448df6f74db674a3377783335a25acafa15cf6191cb31
z0438c03d91dc97620d2acdc68eda8891606d3360f202b96dd90af79294128e3eb83bd88d03b320
zf1b7bf3075efbe41f3c7c5eb1bf39f2792ebc243a13f484f1e8cd6adb5f78998a353da981cf2c3
z203821b1b9fe7112e90bf7bdecaaa50da01c4f7566bb7baafa9a093c055f77b7334a5d10d98479
ze357f1baca6c521bea94896a0514bb55f4876033a6ff53e32a66498b8137a656313dbbe4f4d7f7
z7e35a5bb3a1c59986cc43074088f6f6a99965f20474be86df96a29fc1b71a5268b44f3fe76e249
z75368a899464be205812845326dc3281a7a72432f0aeaf00e2ddb5baa178a8de4564ef5cbb8b1d
z6aabd92e8cae09c3b096b8583f7881c5126f7d4f2438f63d6e7330bb39c44ea51e174204f99a4a
z2ef5b2a6524aad4cf31e5c2ec2dd8fd8490ffa5dbe8fe1240415685d1030f0e3d7ddf351b0528d
z55d1d47a00fa9642195296beb11b3fd1f2eae8302199d672d7624634311f43698a22c1812cd278
zeb22a0ee67f122c1b7775ebd40477c532ca7dd1fbc4b917a660d6fe78f819e1ffbbf76e8b953c2
z87b9f6d28a4c64e33b0776896e7fd5bc893eaa0cd84a6c3c0b944430bc36e7c650c96473ae87b7
z2e3d518fe8507aa8cdcb7e304651087cb1f440b427be2017982288fea4a86c0778aa923fe5e9f5
z2608d496bdd1496680149b605b1f229614e6c191d3c65eec312d1707c86207214234a63225dbb8
ze47c8500ba20fb5e47b1417bab3d7ebc1c533b07c22c64249591a5e3917f30cdb3f0a1c8c24944
zd1a3d4e93e4fab12a4e2280c5d6e25dfbad483fefa330d2df2ec7c32276eef803c668726e79b88
zbcc26e829818f479c8514f446679acc4d2a3bf790a44fb06eea002c7e47a881c136d78ac3afd5d
z118d8c37a6c1a2b0c54a3fad98420daabc28ae083168af4b780c685c12eb5eca4496c2aa1632c7
zbf20b96d82ce2d14f3ef04f03f6e99a84fb3acf159607cd78cce918d1e966cd78a632627521f7b
zaf19add957adc59df6395dca4f51eca54984136ddd33a88bcdcc20a4c3f7e97c1595c70eab6f5e
z614fef082df5a94fcf1cd3c1d11cffde12aa112f30c21795798c4c3a41eeec684b3a13f347b29e
zc8b39f69f394f074fb530c4e7a59a42dec42a27f1ebcdbdfb608e228a126b851ff34e5f721bbfb
z03c7efc325248f3244aa5f530d3333b96c005357d7a2ab4f29798d12ad10b0fdc99cbae371cbf1
zb2a0ae6a83a0ab86c9d2f5c1391348173c9948c611f85076e9241185db1fa43178798dbf590600
z0b78ea9235f54030d722418b7c781ace840eed19ed6ba40d33e4326276733defaf18b60695e276
z091dd3d874c4db9f84b28e943c4705b7e01d2a4b0688bc25a2e55ffd4c53371edc66af130b0d56
z668d09fb9ec4c916302d35a788b9dea483a7f3d5dc49ba1e132bc33503710e0e9f929d35c4cf72
z538b8b3766ece48c8c20ebdff0306f1c5643d1ba66b7c142b41b8ad68cd4590c5c23db883a2555
zc67e6b72acbec10056a0ff4aa7f4088cfb28c026249fc6d6804ee67313a65dff1467facf350ac2
z4014ad50a5b9e2fbb8e804cac8863aa33f915a753ff00a5890e134af1cbd8a5656b623e6b0ed29
z3c8b878c749255f861745844af74829ac41cd599b2109150b109b3d9b8c7aa1ada65bd58477a3f
zaf05dad7bfa4c24c03466a788a76636245d658fbfa77f0a623f2b6314418f79acb37e518f11c23
zfd5ac600b1b34cffcd244d752348deaf8184242ed901e1151db0f4739edd33810a6903933d758d
zc346597904020832ff9913c1c49c7c26bdfa651ed2a7251c47778eeab30e8b142418c74a28e59d
z9eb7bcd0cc9cf7e8ef812e6c0e34f9cc6fdabe365d2f4c0d9000b4e5037f585df24f9f9dce4cdc
z47d295d61975156f12c568d5d2a4c3edb5a8b4bf8a43e1f18b6e2faadc721c501640f8b9359bab
zd9117bfe33fb2f288a39bff6035810c6203598037eae5e6fa0d3b1b4f88894aadf4f8e54ad4949
z2b49f6f26dc5122c9461a1bfe700fcf49c2584ea1a5cebdbeb111846c57987b01d3048007a9e47
zd4d612871dab68ecfdc48c8d65290b205729ec858999831f3cb2fa75dda985d64059b9d3852bed
z05ee4d01d917258e6b71f9fce731b7c96bbd98b73971b2a427895a57c921ca7ec4775123080926
z5597d972d1c977e77fece5c8cea4e989b9d02fa0b3ed9f7e86052b349d0fcedec67b01e8a9c8f1
z2bb5fd466b6a333b3fdd4fca66756c7af929f9379e781e32be3abe7f65419fd53905e274aaeee7
z75398496b743e1a7bd0a1c30c1f822fa3bbb5137bc2bf3e697c8a76608657398746b3e4f12b51a
z96aeca58e9d169c7700c0e70efc33cfb2e338986f07ff43bfaf756cbaf1997f72d0184a5f268c7
z9d52035fe8b0d6149a6b754b4120a403f0c6c467ad802975c0fb21b74b01989652b6151cc4b6c6
z5ec13f9cd39d2640040203415cd3cb7f97ee1f05561bcef71eb9d95f6cc22b59c026f3b0a0ed3d
z11ea56bc701b8c75ee59ef11b741a4b566cb8afd5e2e82f957837f69c36a81cbc30167b682c502
z771356f6ecedb0f85c53bb886b48e618117fbf42002cda16ebf5292139425314f569ea14a813ef
za08c568dbd581e956b9be24f84da9acae9d087150ead8903a2a3e79fe0026a1d19d3762322452f
ze210779de485abd6e68a7daf1024362becb62c5420f93fa91dcd34bdde21b572151885c029382f
z867702c413d3312dc58b4b8711f70df61d3bca9319e6328f2b58a5c40cd26112f1bed73be95756
z9d68b292b6a46180bc7c43ba6ffaa65e32bd547bf02c9174cb40caa22f5ab1317358c1e67a1ed4
z7f7c033195faf1fb55bc07c77f3049550532df0aedb68d6375a0b888b3921d1d1850a0004866a8
z77b882083b1ad2e3dd81e5254380c81bed0653e5d12b83d066ea5c75c664c6e427647b9c7f164f
zfa9844d77885de2b66ea0b80d6100013ab26a1fd6e337be72401f214c615d6540c90e81aadf2d3
zf3673f509766a5e41eb46c539732daad818197a5d4d2562ddaa858edf96b5672bcd2051f780e73
z1822e6a43c2f9b81703133fe05895f725efb81937a7068e58e1f1002b331f374f9bc478e17ffcf
z5cd4f13c2588c9d72802ebb52f3fbc853b3fe0ddee1b3799ba899bbc52aaf8086e59f078e5b338
z95d44a6a10a935a252c479715d8d49519f3bd155484fd9b6671c3d5e98b7fe7ae084090fd62ed7
zb6e92b65d8a9012ffe5a044341bc941230f5986dd021b2f7ce91a20e17aa3eebc8454a4f38f071
z0ebbbb5c3ce24cd0b8261a7c011dcce87a96cad70d6cd3a556f0fb06d4d51aadd88188b1b3ebfd
z89137ebe83c88a4a6c25fba7b4a73d93ca2ea42c4618ccf6018c9efa4480690b41b22335ccde23
z992642d6dd17686b1a9ca711316e0520854ddc5235d01919a7631956be727aa49cb25a2f660730
z8b0fcec10f191c356aba60062b5478a396eb6061309758dba26e6b9a8470028c1392bc63fc3763
z3df17e8929d6edaea3f0c96aefb921cedd6115546718efd2f8e7f40b67a5bfb90cbd2cf73a8b54
za5872086fcc8537b0d823a9c06f3c4c24838124ff978ec9dd6131ac0d26e0e95303c6e8d7f805c
z63b539985aa37dee0d7dc5cdd486694a459f8d145d520bb4931a6a2361246a9957e4138bd52c02
z97fac30982153c58ad8a1ae50a857761ba6dbdf446cb5252b8da884bf56abfa60e1a3c01523f09
zad5232f3f43ae01d8fff85d8ba056474c5f995b8d0dfa047175f276cd9c75d09a23c841536e2c7
z257632365b1ce998eac7e54ec8340a4874d2cff9a6d3afb9d03939dd60c32c9a827d94c46c3dd9
z1d4202853e494433f69b1f6dab6037b27556a97b27e44454e4fa4353c5b9b5900a4649142b0ed1
z0325b001bbcc2c9b6f244199503de70d1916f40602089f53fe5d7e08cd0bba696ca608d0a06914
zbb90a69aada18bfbfe6ff92af8422e044c9668570593f8b434785dd9727b24cf7b8ff53f6f2a17
z75c4c2b51c401969494eedb2c1e7425b0cecb9f44dd1aff2c65801d7323dc1b08428652948612e
z66cf04331a915b527824288abe1b0dbbb9decb6abd1e649b859c4fb00b7c15ea7f894cc1e6bb90
z1b35c3d676fc9f02dfba8c5df260bbf797ff8affbe2374212fd02ca5c4b7e645fd44f1d7f44dbb
z3a1bfc3a846ff1e113e89f0fa62bf65c25eb8ebd6c971caacbb24afcedcf3270292b977d7b230b
zbebbb4857b2b031ef7df212ce0bf574ab03df106528ba741c9cd0cc286416e01c2c25c1b41a465
z8ccfcc60d3d2cd19db8adee46eb6078e1d3120283af6ab7ae359015f1383b6990f24bed33cf9d3
z23f8250c8be3290e969fd67f30dd1ac56f35d6b48d7d12a93798a577400ada8b68d077562d49fb
z278a28b0f3620b410f0e381b5e4fd538aa921e158edd0f78e28cd89ee56b197aa672a2f032235e
z6d35fac1ef17c3e550b0983bacaedaf82507336228a5f071f50545b54d45b3a95c0cef19a831b4
z8e64f1ed6ed4f9af79e07d57aa3b0bc44b1dac9a976ac4468698983d83a300d8e0d318d165dfac
zf0cb354d1651de85657f50c3e13239dacb1f3fe85050039fed48dbdce14b8cb88402cb551d0765
zf99eb844e484c2dbd5bc2d170e0459e4950acc897d9b857c1e4d481eb6b2e9a9953bfc481bfcc4
za78fd673fe89f6a6bb2a6b36e1bf10f3dceecdbd91f8951a1dd422d642ae69d217e86a443720af
zf0e88ddbf8884834404f2d4425f2869d05912bb59c97d9df3b4dd6bf0308a6ecfca91126094409
z2c8ec64d49d31aa5067b0beaed93f69658a39934baadf583f4d939d271882c8a2679007a48bd93
zeb126f4aebbf1f25668bebfdde54817e67d76007b462fcfa32275eafb40244e46d5f7b33a9eb2d
zfaad49cf1f37d4ddeeba36feb0fc955fffcf1bd86ba3581bee42ab91be1ab8d6fd6b00ba1a0631
z3f2e4e8a9a5ca5845690592790961021bc30ca174bd537aaad3055289211db304ee8a37ddccf13
z2a05956701f1198a92c974034daf8e316117bfe3b20246825d3d079e700e00f7e0e4354453354f
zd029e378f8cd3b59a20d6f5d9f0f1090ecdddc3b611d21267f69450603711077ca536fc670e276
z046b804241f3e8c85f3c0725531518d3b97f9b25f63b1639993bc93f86d943c07a6bce134533bc
zf3f361b9d7d7ad543d8bc3d20718847b015ea11656276ca04a8458fd44747d8ee455149fee91d8
z0256851dd35a2e35b2fcc1f6520debb3e985b4c6380d46eb55d9bad5f1ba47854f1442075c05a4
zc8086ce4cd245110c90c1140d5f875a901fed55d2d5a45434a2c52825b59209539e491d97f92b3
zbe77c779bc21d06b311e5e9bcbf429ef95b8aa365b4f26cb405e5dfdc9cd62f8a25a117e508f98
zd4bfa55b7c8faed4060b1a2bb297ea6a31ba083ca10ea130475a17208df9c57d85745b66d65442
zfa65f1fc4e86f898b333630184f54d4673593062a56132e06dbf6183b76c3c69662d2fd9ecf999
z75ff303e3367def4be777019dedd118e9f47683bbe13fff80d06e80a69f991ad872a953b6742e1
z65b3c7feeb2c5f40c2802b3d874b76f418e3ea0695f3c3fa69323ea1b00ae031b547f4539da397
z3b3b85b0f98f800182f5b53656a61828cd9ff1933f21a4e5bf33d298722eb2b4434edea614199f
zbeb4897d1e427f02915fc11bc8b92942676d5c2d84bbdec6c8433a937fde4a684f42a52e9c6f9e
z76d86ffd6ff877a5a8e1f9decc3ce3c6d3450b69b4553d519643f9399ecc354422977b1aab276c
z630f97282cd418d54d9de6b1b48b4372c8a2adcb18dd949b49a7cb95836869b7689003ecba234a
z58177bb54b3283009cfef6378c9e7771eb69e963f0f4f7f8e9c10ec4cd129281e9b51dfc678f39
z1edbd4569d6157ce1e150baf1ed55c9235867ca797acfd6919ae9e3866971398adc490a50f7ef0
z7032c100379b97b4ae82063c62039a98e2c8323dbe5da064fc70d7c51510d682915df80de214a7
zeaba0837b517998ab8cb6719720e56a7bb8236f39e5a4af8ff5c422e4e494a1c24e16503e07f26
z772789bc00ebae45028b5bdaa7cab6d93fabf00534d1c24b53f3bf14ac191a1830545a7b476090
z00f3d3fecccfd92b4697193c5d8eb9d3a4c2f3062cf735827a7b147f52125fb64445631adfec56
z46025524397a3073e7aa078318ca016a5278381b92921491b13c88562e0f64987c8ebae3ac95d6
z257b83cbfd9e9ba52d648ae6834116e4af4e63f97ca3f4b2d0ab307e7357d3defb001b3ce23180
zc1100cdeb97d32be321d1e1ad425ec23eb251f6160fa82eca3f014a1453d8963ecadd9ecf5ccb1
zf0a86fff4c6e88bfeb909628d3de59bd4ab937a28a6b6416fae7ec674bc41b6a114a91f6d923f5
zc95be4c6583d2235a2ad893e90b26c161bb892adb7fef41c0b91e88625293309c2fc56ef05eea9
z287782df12ac6a33ddcb094052af0a7b19ff157ff8df9c5e35a7c31227d310130e48a55a4dd877
z3617c49c1a449232f75fd4ee0deba73adc9b1fa3f8e0a8932a1f73e6835923f598109d7a9fe612
zc83c25a7669284251be50eb794c8a86b454b31582b85034bcd4696a0f10aa8f3fd05e684164cf6
zc818d451824d72d7eb2e4988785c25a67ab60f3d97979356c552f1164115afb1e2cb070fbb9cf3
z7be91206ca01e058e0fbefbe2970669efebb3fe6d08a5a73fa71ef08c14019516e840c804e686d
z3732b6d5fe4dc2b4ce4d9fdbbe5e173bcbf0ffd5a9ee5ac5a028dbcff13e8af2541ea93ab9f2e1
z0a77ab5a7d681224a0b0eb6514e4c7fa702fc30c6464a3ccf27d274febb787f07d963239f46494
zf72cbe7001f249db9bb6247f5b94ce6b8daf5094235e5719687dcb3f9d1591b68aba3aba70842b
z13487300ff3bd11fbf7582f3d6052e3ca4d33fce59e48fc3622c3d6af09711cbe2add41c0b68a2
za7ab4875aae694ebc53f01f1098be4071abb612334df2c4689cfda4cdba96641e1b49f52439e93
ze3f7fbf96c84f1f2bcb83599e6f0ac117bf819263125f160b73a40446c4f792eefd83bf001e551
z507591221bb1a89979804d52b0df69243bb4e4e9df02b396ee7b7680f9c8a7f011e27f2234921d
z37119f0c060004ed641a61dc03e6f0daa6cc7287489c6622785bcffcb848675910fa1637a7ed1e
z273e52332b340b358e64037cd027a4313e59235bb1d8dbee8c000b789a28f2761dd5f988dd351c
z2a719692719e2f9253fa3545a3dec2bfb4db08248aabacd8deb0cd1067cf0092c9f51158985419
z3946e54e5d927f8789b76b43e2d238ecfa024e323380f017a75ee01a541de96ad406468269e885
z2aa39b448448dae52645f650ebed7c2c00851e3a8695cd387eb05882496ad13aff36a9c9116979
z88814acfe6b292d09ad183c4a49fd1b2df6cf9ccadb3c57969430a9acd54508b4b4fef0b970d02
zb8352db824637485bda4e68c96fbcb0b6a8f0cc58f78294b5e9bb96944d4fa8c9752ddf28bed8a
z24f488639775f3e860ed46c4df5a680bac9b2673f4ea78024322002e865d408d5c0cd1113841b0
z6b355139fe8fcaa14903579354f08e89f0493937ee5570fe15f09a0d1b49eea83f1c1db2554979
z9055a265120789b752d77c2f7d3032e4ad3bd25f6674643eb1060339c947d585edad4b64d6120f
zdc0504819c4627e6c246fb8adb98e5517534a114ac6b4822979b255d6c45964431bce68f3235ed
ze9ed669b92310677a042ece6e79cd286b0d2bd9cb2821c7804def2261af486006bd586d4c9d30e
ze767f55713b9eec7ee41ed0bafccf830d4ffa84ead232d45cb58892cde8552774f5649b73c084b
zcb37c3f121235c4c2b5d35643ad7601174ef7cafca0fb8bed68490a982cda172af90d555c1b6d6
z36765be4e2a4c76fc1caeb15ab6940ebe264fca0bae76cc349c8c4b9c5d25ad987fdc5f3e861ed
z645c1504d56d87e9577b82467cceaf6995a03cb118e29de6810de3f999d47ca657d2f4db845093
zcb1a4e2f0b01aea9b0cafab61fa1e279c2c1d2acc324a0c9ce09ee9fa7743dad380c18d5f6ed65
zf3cd1530fa98471ba132e8d61e443ffde77d4112b53d83c79555fc87212dcc71a88d548ca6a483
zb6260085ee24742ed8d48cd858b1d63548aa430e413c4529ae292d101cae30c79d81e47e1433a0
zddf8960dd1b95ffd821a3c8a764d43512b1f3a91a8ff6fc11f16affa85d198e610ce71453b9a7e
z6c1cb162ad9a7f3bb54cbf19c691e3b0829dfb879fac412fded6ddd6ef609294453b98ea4850e9
z9adef17ef78d7b2a3e1630dcde4130fdc65e81bfd9fa54fe2990da5ab864482fe466b122920773
zc5f8fb373c66abdedf4120e866855d6464c0fa2e6992285e16baa2da66f87ea9b306dc8a0b52f9
ze16a170def1d9507d310ca4a1bb65187929609825a24013f389397996728263bce09a74dd1d203
z613c87c318653dc25926d73229a61380dc184a82675e2b963cac88970d7ded2d883f8a2b960a92
zc888fba699f88d000452ca85c7fdc47238c6b0c3275cde2ac0ce2c3697ca3d91c06783263c3bc1
z2b5474cc20a87f2bb516f2b5d38cb8ab175b200bb8c7245c03b9bd06be322848612b26a6a123bf
z13ce1bb9cb2a02e0a5f13b32f8066570f57f58f872ae29b06d7fb17e08f1b0c2668288062f5813
zf527822125181d9aa1a44f1089e7653016d33953eb10c410814fb647ad64f4993cdcacc718723d
z6f04377ccececc76cb0d4e4c92ee8abdbdae52203a280e896c10955ad37c5368bed165fef42f4a
z0ecd3166a570e6d0f7e81c79c077dd2130f163a29545b6f46f46beff772b0d1b3cf6af2ff43c0b
z553535a61932f29ab247b602c81e9f43acc8c025c0bc9cc4efbcaf6a530d3c3cfdff56cf02dfa7
z4d262a4e35276122d7c910d28e37e35eb34ea45a47f077a4a2af1f4c34d723bb238b1bce1ffd93
z931560f38b10e2ce60cf5ea49b995fceab57067dd7f5cdae28935dff0b13055e9871c49523624f
z8f334721221395775fda66a7b69a7e6f4ed30b446f1c28d03b4843a64cb229beed9bc74b39b38f
z056151bf5bdda4360d378e059a33134dd5e141a201c3aea416de59bae8a138d318595ff7179545
zd349527f4b5af758074ad3f62aa4d0022643bb9d5a4e250481e702607f929da9bb6663cd7064ad
z6089a02a86d4de228cd59f1b3a2fa50e033828486baf07a5ae731c0937781c376087cccf5c163e
z42ede3d443186de4341afa07a5d2f1d402fa0ef88f28f9cd410e449cf8d4138554e2c823f4782e
z05a472168a31a4fb83f0a24ac49b7afd1214dc953d740dfccfd708e14d1bb704f9980f6aa6775d
zfe977b0b8e3304ac5c75e42bf9e818b61fadd3df20e61a9936717c553d89ac7acd9e51ed9daff3
zaa17531d591b0b124d8fd82aed77505825a1c3aa896b53c6e1a9c75d16475e5499def6770242c5
zf822ab012a2f084d6e8a3cbd8674623eac8a82c30250a72d96eed56738472840ce5d80d90b9308
z0bc7256955299ba0d60d88ecf7bd3fa4f3a840d50de697c0f32e02869c4fbe06623a5e104fbc2e
z917130b3b8c87f9cd620cf5673d3d628989b9609ed898a8ce64b54e5352ebe8e226faee89119a4
z7420459d410e801bb591c0c9d5d11de26752a7568ca2279b1b702dfc519a1351bd4beeac22831e
z9af6108eb973b070a81c2c77ebb877ebd166560855c2a05174f29117574101d77a6318b4c91069
z1510db78cc2e2a0f73543a3e540ad613dcdc05a7e522af483344dd47a16b202f9a093a3a37438c
z4b271fabb529ec0013a4278b1acd42ef46da39e5857bee751885ba71bb299278c6532b94dfde54
z017243d9486e237822326e47dcc9c935789d680a6ee2237b16b3187ff48a9cc4266d57ffeb261c
z99f4271ed52da7603a001791ece04a30398f14d03b7dd4ea9b7f39549d0a1697ebd4008974ea3c
zd3c07f6a671397a4aa6a79fb7b4138640885b7ccf3ef6b07759643dc18ef2d460a99b88a2b9190
z8d25dd9bd6e77c8b85a50c09dac73eb625d75bba26d610f34c36ab5807b6c3ce9efeb7b1975673
zb6f343a2ade84db294681665d3ea4cf2c50a256252e28bcdb564ce0b8f6c75f4bdfa27e297619f
z090ae88db739198ec1991d48b17491c0136b934558f65e0987a3a959fe9f62b47a43d6e2ab2c0e
zbc528929b4775558228cbec4bbe32aed71e018348cb63fbfbf0f3a9a9317f6ad008ac9b51a7aa0
z9019f40a30851b6e65bc74a2073d3f9155259819c424f107fb8a3f4e6ad4fee834f6c39e47d399
z3fafe4826d7a39971fe0b9d38b659de8eb2bda0d37afb6532d9df08bf74f726cc03e4b5b1f620d
z283cc3117b8a78a8bae2e84c73d1d0c33c14507665d100ca3eb28878ecb476c5331f50de1dc70d
z28c59cb186a3ac4646d197ca0fbe622c953411761373d2114c74a20703ae9f59df2fcefda37632
z837b54883ab828627b2ad225f855ba64ecec435a893dfc126f09c2f5234d53318a4492d5a3c03f
z33a0446c6891f5e2868fcdaae9653cc0ceeba8e7ed4cedea840af5295612fd1edcb5f3ba637cd2
z2e397f808a7f8dccd70a2e639e8eef27611bd500c9d0112ec63ae5c787cd6a1ca9d3d0e4815abe
z0f92658d2b36e9f0ad8f78783d8368151d8017b5c06c0f855c6087df5701b65105b65e432216dc
z7fe3c105a4cb7079a4d1293e3bb54909117415a627c350b96cbbcac3b924f590b5b643e23ee7d1
zc1257fed8e8a76b0c2cff36e675e3f3d4d5205f57a64a7bea6f331252db9648f825b19ca29d957
zbfa8cea4cb354818d4d5c390413f5868c33f1f50ebdcee078032e602fe97aee5f99f180054e4ba
z0774070cf699b4f9ce8e0895dbfb28d079eb7cac5e585bc062838007e81ff31f118c0fa8fab504
zd7dd5c9a753bb1a74e87e939e2e2a4316eb319e0cd3b69cbdea4aff0b5343306c04f488c58de7b
z94d441d4a674cf5e3c236d2e91b501d5d32f7a4b7449fe9b5a68768d9bf5610a97466207fc1b0c
z9a4bff21fff194e866d1da76fd3bf6e0b67fa35f532edd238e6b30209fe56bbf2197969ef4fd04
z0d12e0781d5feb9694044578f2981e75d1606d9048d592b6403f82a181d3307fa2b466a54299d0
z084c260af56012f0155da666035d2fb03c5eaeef620089eb606e0c6dc14f661461365759b9e99f
z728a5531f56ec52027f4b25181433211b22902bb734a5d55c96893c2d664512f071388553e58d8
z0f1c459d3e52118efade7e83e2ef2f881c766707f925e8e1d228e386adf1ba1f7323369e3b01a2
z8ed08c94981b2e3844547ae861b9b386d69f51f207a060e19e43135ae92ba3c97fdacff38a8bbf
zdcda5ae61ec014823b0667e7971cba2fa61e21654d7ee3223baf93d7ba55ab580ac87fa7d70a5e
z99b67db22f9a6878f448d79d569a7a85b79fd7c57e60011ef2afd60dbb32937b9dc411c0732587
zfb26aa1d3c2a28ec30e6566455c52cefc351a388ee339d25f0f889564c2cb3a4437276bf5b69c1
ze2e2ca0e459d5c73fa817449ec7f3ecdeab85b0772fca518580ff6d8a1b675e28cee38078a59d3
z90053260ab1ebf99683723630b7fd8521434dea4725cb99f848b51cdce57aaaaf77f83ab2e052e
z71d21ccf0c5a0bd82f09ba99a99b937c31eba5a5c0696eeb4ca3efb80519771c8af83b9482bd9a
z9e0a273675b14eb541cca431cf616450ce2554fcd3c0cf58b0d94047377ea20d685a986f99c13e
z0f5e7ed8bae9b75bf23cc0ddc03bc7f948cb5d2a0c0870efd4780699a84d800c1562459db3daf7
z27b9023b8765b32e3a3e98c8560e0357cd1fc3e92d717e5a1fe1d46931b570ad18186b3230c7ef
zb621cb6ab0b2c0ac8db1af005bbe119bae1d1c9561a650a6e9417e60fc11fb24e601528a023659
za06f6d2304ae2ca558689bf1ee65da06e2c41ca4e6889ca9e6c662bbcd3a90d0f3412c931f2e9f
zee53a78f974ee80c1118333a12ad876a4dab36b8b616a9486619f5dea9a78d6c9ff2e97dc91334
z22e53dbe8377b57ca61607165eeec5cc4baa95fa54a91a39dc2ae91c3ac39b15839b96e718f349
z5a621269c022800575404aa42d944ec90c15b1f2080e72ff8e21979754c7b046339c1012ed86e3
zdc1606fdfc431079dc0c5157f2dc548125286548bdb62589b7f2e51af4829a6a7d80b5e4b17409
zfd94f69150734655c8b6d791389519478769fc51002df8eff6ae871d3b402b36c05c1bac30e7ed
z9c2913fb7c808f8b02753ca21ef6931043d3857367a2b4dadb2817d6ea7e4fd32f142e3bbc761f
z7ac9ea9647680b4ccfabba798e2dbdf38a1207e5a65a488cdf23420b4dc5623542e561a199ae55
zfd47a188ec122273c16f2f3751c2fbd76df9b07e2c1d3cde78bd6242308cf2671ee4f9c2cee68d
z1bf9302600a284200220c3a0a1e569c83bd24a4ef11581250c586090d9a1d8b6e600e197f3dec0
zf33d6ffc75bb66ba4858cdb0a4ac07aa7256daaf83988003c0da5de1422af7573adac2f66683d6
z7ae05e553103960deb5712dbf608901135e213a40529025515bd1b1e7306a232f733f203c61977
z7de9f6552ed540ecec82112ac5fc0735a1808ea5b2ddc37e8a7fd04fd9bc4617bbdcb2c7e4aa14
z6d0f2b9321e29d7723dc94440425ffeb76cc0680fc9c0f5d5e2cae738b89792ad7bfc335161fd7
zb13a4ae2f365009d871532ffe98b17810e394243fe54458ee28c9ec39c24c76a8b990ea27038df
zac2be147a28f5694d771a508f9e3a336d468a02c7ab6e33865d0e2e1e17f46b33262162c19b2d8
z5382270039a470af84bbbf8d28a2ed8064abfbb2d48b095e69e9ae93f9b93bb92e63a4e3bccfd7
z4df9749983b25a4b63a1f368219f7990e3ad96b784eef9a0be1ec46a5c67e1b07c5451acd60a06
zf1af1680713c5d0aacdab07fc25f9efbb3d6bb5eba75f697b3bab32aaf20f71da1b1a2c255aafd
zf3d2638749b7ffb3053c1a2ed380863826e460fc10679950dfeb73f19626d86a5238a5223b9459
zd69434b6dd1f9a6b8f5ef0304f88fecaf11cbb8c66658b5d5edcbbdfd272c79e01911aee645f86
ze44b7fb127576b6e0610dc4f34f6000d848c83a053e723f28f9848ce6d65cd671289b6a80b5115
z39cf032415992d4d9e01e6278d59c06df23453571d00d527418c1a11bf0ba1a16fb59e69c6e174
z2076e5fc8d40629b670008bc424b2eb6deb0644b3867637df62e544587dd9be44fa7639e419da6
z528447c92b25b0ed574ee974c5590eb7bfb5d578ccd15efd962c131783f4771d5ba07b2b5a9c20
zdd89642cf597aa0c56e3d1acb970d20cc21d188dc838a0755110cfc64cc5b8f44bfa53b43fba9c
z6608a7e5d20a8b7b62ad6338a64dd239a8961f54d51dd05210ea43160ba8dfc8ab6d4fdf1bbefd
zc545ad1a6809ef5c33eaefd3ee8602f1d9c759b78551035b252fc9ae5c9449660afd6b625aef7c
z9c3189f156032dfe1a110139b4c0762515fa76c3adbb4b76f956d83988f4e9eb71ddec8091c186
z49180edf99d21cfded16a1b682729b0689b94f40cd5ba1199190e6ba5b3d0133c2957558949283
zfa154b0f15eab7b8316a346de1a9138986bda1e19bfaf67cd62d9c2b65beacabd8e5c216bf629c
z8c7539702dad28e8537eccd73e580b6f30f6a4a71020c321ed6634faf36b0f3f38268f7a872380
z59422b2d61f12b481863161977221bacb9c2f1aad8d59d5335e0088958016a6eaa49e3ec9402a3
zb5e1ac12f8d35a36b9c0e85e0b323205f78cbdc42c87418aae9dccb3dcd643d7e9b158af4b0021
z330ef91a16c8b289d0ecd793cf6bccdc1f79ef59a588c77af3f23d44c41ce67a820002c8247ff4
z30da28f17a59583f745e2120821c4bcfcaee7d6a1b0b8d9ebdbabdf379ef6e6521e3fd86f091e5
zb89529465d911b80752c06b60c27070361fdaa9ace583826da866d896bf7f2e8a76be3ff32a5cc
zdff456d2120c41eeaa25e6eaaa038324bd5e8d23aac9fb230b7b9d0df35a01578d6068865f958f
z44545b6e1706996a252b80a14a3569ab91b0e07b4cef46f8427794fc291528fa0b58a58c44b8b8
zfb72dac697594f491ce3309b29a71af8a966c4429fdd1661714d34db9f870df41c68bfe226dad8
zdd343f09a32117ac69dac8a43eebc1988f60026a44dc2c6f4c3f78c79c47f74d08c4bd3ecb8432
z0d89e8a8427fb2ebd0efe24ce175ec21659bbfe3b29d80c79571cf7ce40f1d5525ba46b749fbf0
z00ee302e3d725829028f57e924e982f951f18f04e0f03f49758610ccf9552ae3ed80d205ee2117
z852a06895bab7bc321b8edef054db8bcc61df6f0548f68cc7c0d102c238d4499f4cb8dc0a853d9
zdfcde8a827afcd4ffe0ca4b3a490e8ef7b527b7dd628d01284f0c4c6f5f8c1717576655d8e2a96
z11a04eaa5386d3b493646ac3be1950e1f736f48dbfcf67dc4ec67c12e432b0dfef85b888ba2ff8
z09bbc5f54851d8f3f08b3aaf4f2363f39eda49405a848824e659042892144fd2eeeed579204db1
zf7c5f769f68e95576b56fa6cfe02381a89bfdc42d89b24c280fdd5521e762d1ce40349232af8d7
z8d6ff0e6db0c3ab419a78fa3650b5c34e9107332e1e267c956f38411d91a8c36301b6b58fb734b
z72317bfe62ebcb478a25a88e5f07f4657705711d5884bd6cc3b2caa05e8cb2126ea985deb329a8
ze7c19f69d4272e688770e832a43bac6a802b723059310e09c3d45af32fd4ce2ee1e38dd23d61b4
z72047d010768dcea4419a225e3833fc1f3df82b10acaf50369b417bd28a8cb31517547a4c2910d
za1bfe8956599b6d41cb8a617c1d25015d858f9da612c1e799f38b974d43bc5aa6ad6d77c358846
z9a938262899d8e35371f51e0b16987fdd03193c0d983d0b99935e56ae89e47b682a952147f48e8
z09aa4077b8ceaf4f5cdd94a24ffb362a69673139263a7f31e3debfb1f6102061687d8b2775c7c6
z51845b1bc358af40c56f45443667a507e6a329b9658b0664271fa13a598d9e608a85cad3db17cc
z354e6aeaa27a90843064f46500a79db76f12fcfafcfa6f69d0a06538082510e230dcffe5bcbd05
z0673d0c272ffe86a05299e78eb5ae4d25a10948b3a51f5623fe12a85e52fc9bc8f649521418df5
zcdef6e57c9b14cba0aafc6549d21356f3d62b0f7fb0ccda2d87472e9d82c999cc2eb9cd1848082
z6000f68df5d1caff7ced48982752475e044e5a0a402a35cac01e2ad77961e76cf8bea41efe4cee
za697b04b02cdcdd38c0a127bafa2f4e1dec3150e9905feba5c8c9d6bc8a16a25344a9032a4896f
za13d9fd14b7ab5f3bd2b024bd06841220c803d3e35184bc8fdba80de5bdd39672b19fab79c8c15
ze291aee0a2f1abd004f01c897cf470c14bc6cccc3a865082d2079a34c2585e8b2236a168084f70
za40c27bfebc4902cedb44157294f6004f1eee8c052d1062e334fa9b4dc20bb94f03a99fd67f73b
za73946207c4ba63a56c3f3658431b3913b9cf6864efa978a0c1c5f0238036ddc874e8ed088e18e
z4ea19b0a220c17995ee07f3828a479bb361366936d01ffefdc673152f66f0448803f52d6edfbeb
z239041aa7dd79154576a83391f6cf6d3ada682a69311a1a4a3c8c37841c42a2cf2085ec31d029a
z0833b6c1d3492fcbb8acaa8ff870d8ae107e7799c949590f0c6aa7b344b8d4f66c4cd05df7d23d
z64fea72904dbb3a7db133ba666c3dec59d35334c4ec5859f35b1d1870ba9f6b6710ab228c75ea4
za9b74fa9da0fea6bedb903caeffcb5ebbe098ae6b2696e58dcde2d4bcdb8591d09c40f74d26ada
z838ed460bd0dcae0356ff177ee93f2802dc10af6dcc92aa80a020cec2bf87b05614964a3cf8189
z0850fbb088a59a7cac5f4c1d04701aa13f53b2d944768c38f7dd3ac4dde91fe62c194bd4a19203
zd0738cfc87059150a126e61688e2adb6844f1a40a256b176c9d91770af2993f4da3b272cc6f176
z5d88ee18ffe1eb0579ccb19d69719370e819f1281ced1e3b5801888ab5acf5e4d48db3fb3c0d6a
z0cca3b02bf02f4a57dbd506a4e607a3248573f1b98f4bcd1b4e659199e1eab284e4c2fb48e795f
z369bd1f48e518fa608fce712d9b28688ab5675da3938b08c8dc2cd8858b2ea617f0f0056faf4ee
z286c61b91b3d09895f55a4761eaadc486365c715fbcfc48b33927806e54bc64e351570d7ae93e9
z2004e153571a501fda002ef36c0b932d629de5b18e76d5c42eda5aa554e6b6ae31879804b6e0b2
z580e5be473c05b15154b9ac453185c09ede166b8ba731df46641115cad890c24894ad894a5fdeb
z8c1f981ae5008846b2a19aae63cd1c0b5f672f1604036ce15fe37bf0f4b9cf4de57015b103e1a9
z3aca56ee0ca5e81a940f69d6226de9f6a2095e79100e45f4510b652fcc6516417c4851470b7829
zabd7cb8c05598fa613515d05274319c30fa80d29cc67ed2f3c298e35b7cd7eced1eeee136d8961
z4e117f713c3c77b1e8f00c9d9f74e4538ec691b7eab8f3ef38fea35a048fce3c2c9fb0cfc6bd86
z8499c4ed7fbffdbfdb2829c24ab3ff075cc66f0b9c871b53fe2d5aa42f92b9cecb2ebff204768f
z05fc0af7d30b83aec1889da400447e3cf9824b20bb22e96db9fc8b81cfd100a01d7602c8f10830
z8b7366f1f9adfd9268c915fdf6b5e0b75cf4b89f375ca03f82a1bce11b53f2161fb476c2197d52
z5364372decb293d0b660d5c918bb43f8c8052c487278be1302f017a165b433ad8f31605b1f7d4a
z92a19a425c41f06b0d4d8e604a17e8758bfe0f65c32eef8c147f85765781ac09f121e101ed4c94
z48ef7e8239103c25a9ae6d8feb8de3f5577d48348de86afb96440086e1d2311a07b7eada39ee4d
z7cdb6d19fea2a633b4279b9b6143d26ab2c4e3919f524a5337b2e0776a3d346bd36fc74c85a189
z88c8b28475a04a85a210f16a651aab7d343e7523667437c7fcdad4bf4924648790c1fa5ae62484
z500acfef9b127d52513d4600f1b62becf5f42a99f6ca17b84384655bc8ee0d2e09c830923dcf29
zb7325faca0a00ee0c7fbab76e2e1f3e507df8970a7b9a108d0197aaef9b974b89005be2872caaa
z525965286287d561e6096f84e4a57b5dcfcfb1d9de41b055454b08bae13b4cf5f617f967f51920
z4afeea433ab7cd1070bcd2cedd19768258e7788210a1fbb95b0d57741af23f0a2700e735496ffa
ze8dee36193942c2fee13f1c076cddbc4d196ecb0fb728b9d43855eae23b7c5ed5cc308e4cdebd7
zc208f01291d153082edf5d4dda3ec36cbd05c5ac1ec3acfff97aee8f26a3c3394e49fdc23e5248
zc2ee3efda5e3b23b4f29ad6013f9c5154e9620a957b6a2d959a3e04db50b46d591be10900dcde7
z52fe69ac2bd95bd7d3c937562ca7e9511f7d18f329a29268ad7d378ad2906a89ada0629b7d7a8a
zff809eeb38071db90ceadd19cccf72dde231d092f8e0cefdacf460decd05a8df8f2a26a56f2655
ze0d8179d398373a9385c4815193e0348320439e1ec813ef954220b9cbd0ad657984e2e83c6e0e0
ze8721311c061dd62012483003cb5a00baf75997bdebc341be378a158bd86515eabe3f69bb9f0e3
zea1acca963fa2a29882eed4f5e495890a0c5ca96c4bdbc46ad100ed44d021df54fc2e7884e301c
ze9faf999a1717cb009eb5ca79cf6e06000c8dc40376992522517ec17aeab32459129f4fbcb43d9
z813d42510f05905cdd1638916714c63eef14b765af290de679c1aaaf78b68a05a168e987d7d250
zb38a804ead6abf173ebeeae1fc0cc9fcd99783151379844e243d7e0f849f56be2d2d0d8c9dde4c
zd5a3181eb254b1362d3f712227a429caf9292a33fd0036df46975928a220434ad3addfdfc17a23
z767a0708e3412f6687c340c0e74ac3b723dd83a6f83e7bf740950de01fffb0e909e0dd0691e885
z272eeb26bc29af17c71d5990e320e5d8676a201687d2e87e1a733d9ce3dd0dc781492e2d29f45e
z63b7555e1fecd7c77f037ad23e35074e6a8f6ba4a9a39a4c9f080b04efe57c97a2a867911faeea
zfa92d7bc843d284040c6076602185c005feb42c0186592f4e67158393bf47a85c14b201b7072ce
z7cf3eaedafcb30f8d99e153d2441c766b5bc4068df34415143fbbc2ad5012aad1f3722e42e4101
z290c2f7db7f7013db9871b04c85a3a48ecda1c1613d7415dd577c70ec9ef9cbca93ddfc83533d2
zdc634f845da2e58515a39b4176570df9e380c347a9d798176c769a0032e9e1cafba42480cc0d2d
z9279b8de9f8e688183488c041f781f8e398671afa05413e94ee3a4226fef590cc979509e0a5f0a
z34f39201abcf824cdd27bd1c64c0b42e0404eb1755c06cfa5a398ecd3208e4c47c8052fb68e520
zf65522083bc5abffaeb2392e394569e38e4990a67add47ef3e4e43c46173b8442fab534cf125ea
z2ad365f1d3de78a3acc848c79dda00567847325fc6845a99a4e20ddb620af12d9727f2548ff77b
z7d4379991c62540ef9de8443c4a62ea7fa55a7b7cc1d47255d9f292c751de3c3422c3719dd60e6
zb2c80a4f9c362d3a449f2edcf37b9cc8cd15f22f520e2e9121ea6aa35212b2a57e16d37199012c
z63daca78a6f53e9d3631c96f7408d90d941a585374c935bca832a062101f233d1c1f61c0d46a9a
z5c2c3861784dc02bd604ac7dab900c1a8a20942ac95b1cdf44d1ec6469929f945d38b7a3ac3a77
z9b30c06ee4f0056803c761c994dbe3f75bfef7ceecb3290573b5b6e5c41880d80e9fbf85799005
zf532d1da08c6ec5dc7dd01b975ecd6957ce7329c215626ff735d27b59e307e17c69824a36f8a5f
zc87fa77b4bfdfcc51e0f57dcd103352b900e781f0e74a91fd4c45acddf37e488c6adaad1d460e3
z36446ff466f24f1b29c9f4971fcd9232828d6d942b177344b7db010297f90395723be1271ec39a
zfe081cb82a0288f7c5ab2a8fa203d782549b19245ccafb92c46da9d8f9fc252643e48c1bfeac76
z7cd8e42fe39481dbf9aba8d07b64e8d08268b77f32117ba314802c883e5831bad218085c50e02c
z44d7abc441b399a02c1b6f79c2f41e73481431be4726636c23fa6f622355ad49a0cd36e22aeeab
zef73e7e2ebd0a72eb955dd2a0b56401e258aeefe88684ea6aa5adfbaed61aa4e530f49887c2273
zac2c6d6e437787964b30930dc960211dff064c094131474148d36f307893fb8fd2795a431a8a97
zc62ac2b4fbaa1448e2e097f0aea001da874c01686e1de188be553be074785fa3dc42ba9cb10e5c
za00524efbbe4a51dc7c8e0075ac130f5f12b855b7fdcbf0c584a62b22e0f21d874ac074dd12029
z806057f80159601274ada698d33318b57bf41e95b24465957007124360ff2e82342a76308b54f4
zeaac96fd4b3c314df46b074dcb63b923b48642530a5b27a4537776ca6963c06797267b699cfb45
z9e93edfe69b9cff7794e5aecd4162c8cbd8d7b48b7ec9d2d22da7b129dfe56b821333bca67cbd0
z0d8cb5156efbde647c1db0c5bd6b5cfaab90d0d22f099c1f912494c4e610f1ded8fcc0f96ac67e
zc425cb8a724d50af18840b72849e127a843246fc4b454a03b47fe4856d9718f8555b1e2f2248d5
zd9e4d9b09eab5871ca5ec5d770388127c83bc35dc17f4ae47e202c7c4cbbeb89f3fe1e96792607
z9fd1c00888221436a217f3c4850e02b1b0431f2a2ab22cc88df971f5665bc1b4167ffafce8e936
zb6b5fd358fef4238c95faabaa51ea6b68d27d70a8bb7bd071f02f737ed97e9d80f4308441f326e
za5f34ea175ffe74f7816c9d1bbc5f4e14615579f6871b96a44103513fb5aafe463a5d96c244f26
z9f482a5d8a5a6ad026a06f5c97d9368e84c378f1cdfc4e368edfe58b3a07b5129f990d4ef52eca
z2404c7568bdc9fc8f04dfb34d000b9b71252fc901f4bfbada07a9ea1ac3b4679efa26ec1476981
z1df1c358ecd8e7fc740d7e31b1ca0384f095d540f16ce3662fd37cced7faa577a3e33dbf1cf2eb
zcf696c223ad2f8c44342af48bbff03b8dbed6cfff7fae2bacb6f787bcfab2b9fc6d4d96f1d7e4b
z582efb3e03eaf755d78b4b6f258f869b896ba0aced9ff37d6befbc454cb0df07fbfbdb067dd976
zb5a051965929c39006385d2edb348b5a741147c781a316180681cfae5e53798869b8574c9050c3
z59f9559d7a72a03b02c4f1cb52e672a7059c604432abe7acc8167c0bad3124636d36d6523201d0
z7b32351ede6afc766a4ef250bb7ceda8e9daf757ef94d617a120ac389189fec4bfe7500b7b579a
za8b4b9da88d6bcf58946011ed9d3a50196a708beac055ffd0ed3d89944a56e7da84fa26abd6ede
z3585d8d8a485b235401072457d9eb192419a1f025a1ea585f2ba138c2889720b3eec840d964363
zefebaf7a6589ccad07ad281ae38f4ee12613c739f2f1a9b88abbd54509bbfc2bca4d41ac9c1270
z808d5e60c8be696714e447aff587e5599285186f93050079c11b6ab144776c3c1e29939c5417ef
z6bae47e99a27e5fe5f60fc46b67b0e56a88375c38319e0362cf7bac7132b5fb0205c9579dae1f6
ze2fb0bf0790698f6ee70161f1bd9501807ec9dd61eb60866dc596a2cdc59863161dc0976f5fa1c
z7980075aef0fde8c2037a58449757a0bdb5c403e67f962878014f5d770b514bd967a62269e6c20
z514f76692fdc168639914baa7eeccbcddbbeb5e49d46726ad89039433c776cdcc7b7b705cbc474
zcc81c7a917dfdf411f6f69c0803a1f8c9412e6da9f92e8acaa586f6568f50062384754d33dccfd
z19efe1b352442caaa8b2ed26f27bb8ac1cbd3d8e417da31b1f56165467fd9f2f04b36aee79aa81
zd3d1dc018d4b059284fc31c394b477b29cce997c31c8bd49b2b21aae95d9b06f2e8365fbddefe2
z326d56c39f74bae072f0bc75aa17bf5c2d1250a5dc6e11966902f101c88f71f5d5289d606805dd
z1aa1e674e757208d90e96709b4cc2d7a3bfa4fd40cce8dc701bfd1b1c66ced3e7a4d3baf75251b
z5910172fcd3bfc1b67addba7e489b7dac5c37d5ae2b9aaec0a1d12fe39bd69b29159e71e431959
zdcb5c929c4d1987fde9cb7ef328c5adc432fabfbbeafaa30ae4b3dbac69900f22c5f0f9b7e9a00
z19bf90cff21ba0e0ceb7c87fa88278bacf24d46a7239c8bd46b317c2be27d522a72c28c505f7e7
z6d190a7619ee1668fbb0af9f68237a229c0585d6dcbfbbb3d360e98a00faebcf4b56f448ec1334
zd1f19354986207db61c78a9b8a50d093bc6dc0f2e343d63e920e3bbd3f135cfc8d2e4cf443ae8d
z4be3979fc2f79b97dccd665de3560daa94182e5405b5106a0edadeab33f7d07c1df94fc7cf6ba0
z7ca77d2aca8686194d7600b8290a5a1b4f42b6511506f1eb60f594ae18f7e47b7df94f7ebb8f36
z531eaaa7247a169be2928201fae4df476a4e494030b27649273f81495f260c4d68d188b4ef9673
z55873067c57df416b7261b4e7d03d6d94494f45e78fbaf2a9877f06c3de43fbd89613c8aa774b1
zd8191b6730840e7580bb5a4786cee8e782aab78c070403e4c23e1aa1e66cb9691628a8cba4dae1
z90ca867355997be234ee768cdd4510cc7506e2f7e0592c953a020ac1ee606b78e5e31cce53c076
z4f51d556016542ada3f719e1176feea4b9bebf0817aed252886b45d35c2abfbf2dd24a352bee62
z13a28dc7ef70972680025445d7b6f458fe0b2f12fd0e9f1785edb72bbda9cc6b41a772a8f53eb8
z971de0ec09ac408518391b73d0cfedcb2c9781ba40198edcf7b94753a4fa6ba27641b96c1581dc
z2762b2132eda46468f036b559ef4121ddd56093aa617154b7d999abf0b35f5b93ba481a404a4db
zf1bb13dcff72a8ad4dc9f43c8b736550a57256e88de799ca0ed667a9e965767db600330391ce37
z46f75bc56286b582f0b36c307c02f398204226ad22e43bfe7616860fbdfe3a95e33e432fb2faca
z504fc9ba987afa110af1881ac7cfad854ad036ac52d2b14d86d4eca148e5e93aea5e91cc1cba56
z71de02a96ce3230db5c26e9097121b8b2e42345b25bc6b2c81a8cb3f5d63158a578e4fe3d5eddf
zdd0ed0a7f9f09c34ab227256025cc8cedc77475769bb458a8be1cfb87bbf74f30c27f08154399c
z0357daa4ac85e909b0c355571778c996f51b4f0f09cfefd33c91e848b943e35813bb17eade1f67
zc2d7a7e7d8ed35ec84d185fa5e178579b4e6356423b6962432d283431c1c94b813903251216617
z86c4319ebda677ae01b836de8b2123a23943f83505bd389224fa598e7c7d55edd01c54b19f600e
z6f739e6e2a28e5ea12bd01881a60584e003a8d5023effa0d665d3f6f41c5b20c5e188e1e203743
zefd28f1db11c58e4cb8308eace0ff7d8015a5950162b730cbdbab2fc02269620e7a93cf665d175
ze445d3f6c2eca2799d78af599744364693d2816ce04aba259f66bc8b4d582d09fe2c44be377ab5
za2164d80e2d3e259667ad50caa7e3dafd2ffdda39f162299bd7a858b6d37d81cb0ccc3beca964f
zc54b44f98db6c2bd27c68103e8b328927b937b719634e23c602b05ad14716cfff8a27d8db6fd5b
zabad351be2ef689d24ad4ed136ab247181fcb7af3633d9b912fb2b81e18ca13422016e608c3ba0
z2a79525eeab451008d32b6072d658e53ca85353f3ef8393b214ca7942ae4a02d14f5337a62b991
z71437d2e85ab5fcae977c18630b8b5e6edc41b7915f5380fa3e8a5fc54c7d890f846cbac8ac8f6
z906364113cc5666e3357f6b2954823ba69be9fceb0876d7426cd4c1787ffd7f7a4cbd71c7e65aa
z7de14208a9090ecabe866dcacb40a72a2ca97bc0009aa290b86af832b887e8e41d00d1140c0ba4
z5eb7f88468326bbcb189c668d1338e1256565e254e942da05c5786891968963ef4c3b52423adf9
z39d26b4147a8fa9071354edd6ccceae0f82c562b778845ca9de0c0892132dfe21b51b7a12962d1
z7a22b57df517c3647e7fe3d4d660b17dd6f9f5412a191cf3220d356d538d5ef5486d760a21d486
z3f02c15d096cfd02a8bbd2e0423c0c3267fda338271448a0ee84fec8724984a4a2b47601626850
zb3ed3adedc92cc807406ec8795a00b4258859a4f97328ccc606d4d3c23fc5838d45dbbbc4a9183
z25ecd85e3f91dd1ae94affd9ac1be6fd58bb9d64d54c97736ce2056e92627e3188622ad21c8c63
z30ef243601d095bc626544d3f7ba2d47645f5ac843b636609138416467b65ee8405eb38bcf8b73
z7955789e74290289e7b939a041e24e0bf4826115d978117203c2f11a96eff7225bc7bb1260ed98
z6ae730fe3d07dc99f10b0afc135cdd57305a350547874814036f2cf548aea808c576698c7ab666
zd03be64c4fdf3a9bcfc49796f10224492519f739df41bdb6a7075e9d303948eb81942696479bee
z9bacd1f8973bfe7e4873a7b4dfdc2aae4d314e31964751ada4035793ee330af91c37d813f42409
z13923e47a54c3b7f46400fdbade383f1f59c824fcfda6f37f50ac384c01987cb6765090d6e829d
z653750b8f7c03254f75a8874fb503c5ca49aac3a06e3c77e18fb1f3b664d6ee49c018b87877ff8
z0310302f5729dcb2fe60e988c3cb69e68820285c7d3f3b686f966dd3a4132aecb8f3abb03dc549
z32a1d54ad345303cafbf657714a49d2c17ef93f2a764d2f64ba2429478309ea190f16e859746f2
zfb35d30bc0ce320f07474a1af62aa1eed93bfd2395dd648b88c3335c64af0433eac15c681b252f
z07bfe98fb8ab944eb1a011b9a0e3ac42d880baaba28f4b5f7eeb1ecec1ca92ef23caa648ee59a5
z932f88e4240ffc86b0dbbde7648559fa13c622cde7ce82197b53ed903c564fa56f7154cb02f6d4
zb20b970af942d919ee989f0ad566cc508e520547f08ad59447c07bd80ef5123d9110f6e5a1a168
z66bd872fc710662e92b17adbe8a21895026f15680d94755875445830dee1bb0058112254bc867c
z7812897fd2571320b3f1a43335e35ecd51a7a7f94648b8ddcb93902c62ca7648d56c343ed5e7fa
zb6a6ea7ee0bc5af1e7391ed54a0fa7db7a3ec4e9c50a1cc3a06f91931106be80ec598a67de681a
zf2dea33b6c259a696b083a19451d09fe68ad9caf464589c744e182f7485ca1deaf8bf2618320f9
z564911d7250ef9ac244f040909f455ff2817e97198153cda8bdd2a73d37cff78c522df68eb46ba
z38b45e6992a85a65285dc381ce4029a3c894fe5cc1b458ec5df8786d6f2f9759e88632706037fe
z4c597c1a60abbeb439a743d275d8e02e75f0017202628250ded941e09a36ac18a3e5132b06af80
zb8725686acdb005db2b38c8c223f6b30957b6b93ab33d7e23fbef92d87ffb4270eddb2dc3f65ec
z0efd211171ff017d7a504233306323599806fa48887ecaa1aaf809ca22d823bfb936115a3bbb36
z0b8895f865157a0a592dde130ef668967bf7423e8d6d905569e04ad89a793f9572e7ce6a5a078e
z909c34e065319f8fb8dd23ed452bd97117074c6e59de389eeaac2c86d66239ffe7ea0060a13da1
z0ffca95f6dd7d85a3e3205646c54b2167cf7f8059f7a15343793479f641724b79bd7c49b26d046
zb6aca18eb5fa9fbb1c0ead5fa8d13a72df2130caa521c4680961badbeb80f7fb235e8e89f73e5e
z41c2912eadc10b2bc8f49f6fcf28a49ae688a6c9daa878f0cf358f2f7792726125f266b8e5477d
zc4e2bda69a5c36af61d1e6f9c595c12020b5a43962ac4903a03a76b3845f542a8c1b8c6ea7e231
z5b91afa4cb063c37c62c433771347a5e48828842281707e1723cdc76a0214ca1c5ce9dfb013cd3
zf63ee55462383e4dedf10c9e266cda104edc71b2aceb614fd47704e68ac290dde157dd7eada71e
z5b4ae82ae02905042ef191a9a74b9985c7b23ca4502c224e95d6b37fc8d3779cd67dacbcaa6b74
ze02282903535f6bab4a0ec6dedd5ea1fce389310240d42250077bf57283c43a08df51aed867c30
z78fa8999e04dd9c34293e6829243af15e9b108576559793bbeed45dae197b574a379774900b2f4
z218c0c147eb70bebef1e0fcc5b00523ce0e7e70060424f2fcf39514e942834a09ebb3a6f004283
z90635cdbe4167a698daa392cf5cbaee2fc914d71615b5d57eb5fbf525e636f8c1fd9a5c34271e5
z66490de426a790cd4050b41c27f07607d81474bbab959ad6ae67357d035fdd6028ba5758570b6a
zbbd07d0f00a496a67bfeb235fd1e7a70f29d3db51336abf4a8e825ce8d5b8f593093605b9ee8e9
z1ddccb61ef658ccb4526a158ef36b11c30da2e2448dbd2ce3e1b35eff86b9ab617a2d8d15a4bd8
z0489fbdf649db061d2157eb3adc3a42c87d5c6c566728c5e60447191e2e3c0d26f51d37f280473
z3c6842131ce59de1da6c068de1704c5b349a6e0f795321aba6d999fb669b39712e98967ec2d406
z38244b63f974ee6f3a3b59a7df07bba3552f5c60774f06cb0ddc3954141f7d31e502ec560a4b00
z7008adcd7db18330aa4d604c706ade939e05bf8366e1f0c07be1265bfe1cbe8405cc14b2edcb23
z9223870b7f295102120361db55dff04ea524a1dcf212a7fec53b1399edd678f341ef0c455491f2
zdf6ac1a735c5c15a97fdbf239d90514151ec12b72c40a65b8b91c3516721ac1da7af743b6001cd
z42e8c0f161abbbb90f6ad55670f90a80968af2279a26dd02a2de9573d79d85d735abcc5ac7b411
z993ad29275423f1e97d652d31011326469fc34539cb491cfedfd5aea089aa9110e6849ca8432fe
zd42533f419d36db3283a291bb7dcdf1b94e46231c20db8aaee98126cb2dd50d0c8a648c5aa7f3c
zf93d707b68c2b6c19b58085933c3cbb639790bff377da40d3169386323f0a7a364516d33b2d285
z9fea80f9f692727c796f04864ad7bd6273111bdd552c99a83ba8c0e88e0c8237bf956414b63b40
z9286d5bb95b347646af21540f1b1a3c43fbe6d96e5a2bddcfad81079f8b56111421ac0d910094c
z3ff9e24ee91094d923868c1648bfdbd89182e56d6bbab1ea3a14b8e093e59b4a65d6c8fd747d1b
z2734cd116207e914fc845862eab2cbe79f6c05e59eb4bafb2e7d34876cb51e993f065677cac51e
z3ba98f894667630d1e3b62f714f111f2a724bdd240fd9e5f79906e056cf3f4bd237bee76896ebb
z15497b58ec6df1d24005358205711208b437defdb6058a5aa6cbb6506cb1a4b49e55aa708d45ad
zbf7738445abbfadd31ec120ea2448f3d20e3869efe0dcb90bcf1b2d889f29354408af14d88b2f2
z41d688854d31a473cc70fcbfa82de728cfc7de6ae428d311a6561606e2a3ea2974872ca5959206
z0ae32823957ddcbce3075a8194d25cc7300eda105b461ac968d08ba12ec7475a7683802a57b9f2
ze400fc1bb2f530448eadec3810396190465f720bdb935b7e26dba61b7b859099d852d2503b0697
z2e840a929405c405887e6c74a55aaba3b1e3c2baae3ed9ba0786daaed967f6406ffae164e88c74
z164c9cd2bf6f5160a783e5455b1cd130817d6eb4f8b19f82093637e44f7d6b6ff0531cf45a92f0
z8311281da5b5c1a26bfa24abb2f9618df9e912eb3386d36bb9a890f7a0298cad25e49b17db6db8
zace455e2dc91fb6bff197200654e11acd60f5543078337f37a4f4d2e2d126fcd637014e028e081
z62bfc488392b2c3e937cf595e59d33bff8aa2464f6881215a65c7ed9e96c4029d43ef04182e5e7
zfa6543b7501d9b5b5dcb746921c79d9a42674980284494ff5ac681f38389b97f5665043f79e03c
z2d213f9510c97bd24cf5e667600516e2dfc499b51ac28bce1e9995f9f2f99a277e57190363d6bc
zcfe77dbc5ac3e50dd67a0bdb02518f0062c2d5e5e43600a4e30c01ca182cf50830a0107b1596ca
zcd8c10b9903e3c25ee05623400021c9207b20ddfe5df2e0fc6bee7e414068cf0bcd8e77ba990b0
zd162e66090508135b65bfdc7826002db7909c7051c11035ceecb86553e33aca89831b212d80b64
z746163711a6d1bd008379f09b6e7c2f97d0f2244a5790e4e5ea494f63280f4254f5cd0dc942cb5
z070f8ba2a35f8f550ca2c5412feaf4459c93a53ae4c2c185050f6368781dd2ae032a4e9a03628b
zd2b75d86f05d16d8282318d98ee4b8862ebcd3d969dbf6e3c94a65fbde1601e6cbbbf0d36aa44f
z8ae177242a2cceedc1bfc618afce137e78708c8a059a7fddd0ed75a09812f736f9b588db65ae18
z47ba6b0bddfa41ade349f0161346c0be841554931d0a8c79e95aac7ab2a3115276227b030b19ac
zd304e86b37a6de2d9d2ae94612a968a2a1dbe4e2285140a32cc3e1762bdce4228079b0d6ef807a
z1d94389cced25255f922c3071aa4baf145c39a57a4f16fce7e3c762d5a207a43c0aa1a7195e1ef
z277ca325c4e90e5495fe1a3919a04bfa682840cc64d765ae3c854e62bb968bde1d509eaf15a648
z4cec04ac5f1f39b72092231f0e58ac2010dea16b8bbbf15d5d61fea53d45bd82435dfcc4a10e19
z69defa3d56754f1d3c4dc9df7c6ce37a935128210a03354f318496b7e50e26929679042f499157
zd91177d2f15a8135aa7dde1dd5434df6610cf49bbab5647f4df67d377f173de435c3fc51f0ed5c
zf6c4eec72016b094210ca377ea01818c9ce99562876e4a82ebd6072a2470b332fb105ba067bd26
z4592fb4f29c6e9ee13561c325ba2494b46e0f0bd8e423e6852013f2aaa64d2132d393e0f604096
z02125d19318f8bfd47f31a7c343855ffa37255394674bf6566944e185fbaa2ac73ee730ff38c6d
zd435122e5fbe0cf71b7fd10f53e26f923856191aef10ddac92da200b1790db41597982285f07ad
zd8643cdd7bec3586422e9651a0ab509bb626986d18e7f9f8e1a44446393ce53d3f03bb56a99dfa
z281f614d4b7c7d1f69083ee8426d1aec0ffc9eefb406a65b42ef31bf6334c775b209485e598f78
z780abe1e72dbe008b2b2afe1b7a588268959a4ad69987677681796e11760d829a08f6eb92b7468
zf919e9f5bd6c9c0c7ba740b93518266f967b2dbb61e414596acff35b9ecce99a3b44d368f46b1a
z3598b5d490783f1088a3228e55bf6173401fd6cc1bccd14e08e4399595a0959bb998cdfe44f7d6
z0041fc5084291bbbf7ae6172a8397944fe622f29b22786a5667a49b68ae4e4ffd813e14bb28348
zcbc6b5de62c5e8a81a727538d73d3acfab18b4363b89da651a9d95dacd1beecc1cacc4e4645625
z83b8b0eb7e8bea022c7adf00d6c530e348fdc0a9b59e7bce5da194c70e21272318e800fe6de561
zb2e0a3db7c106b1a20574630e1f94451d6a2efa26644a3338388c2f0f2e60b402fb1e8d5b07894
z548cf777232a750816b761e81b96feb78ee5cc27461bfb5f97bc9b0a2029c11d191e09ec934487
z1bb26a48b780e3e15b2a33a138df17fbfce77e8d785c9022ebacfe22d1964c83fafcfea4755476
z0516a10e8d1be813dfcc8523908cbcdd877a5efce18efcf541e77b3e512f2ae2c63105f1b3f494
z1768463f337e12cc6e74e0a1446e8f879de85a8cd8989a87dfe5c3bcb2b1f6056de7e4e9b227d4
zed1e4a779c63c155de6a09bbaf53259d0e5379e84bada127dbbe262761072e8cdcc4200f158db1
z83e95a2c793efec4413e01fda89f5dbe3d1970c1c7f95a0df5a658914b3dc4ba0e28a99df5054a
zf93e5dcc7877fe6465c378c1278ca725f86df0d290e652bb360a6debe1bd55474305a496ed880c
z6fcd76927fa9b3704cec755acb93c7901cbc0dcfd83c7e7f7c157f44403ce6257162cf8160a372
zaea6965690b0f963d6dea2af172285358c1a7daabe584d539a08604b6304fdb7d117b406902d8b
z084daecc009f72780cf5cfa322290b41e027db8fd8ea4bda7e5ab3c4f0797a03a567946d81a167
z0a3b152022d5757cf50f580dc403ad9edd3af0a91b7454407d630938198ee5438d6c7724774f6f
zbb483a368ec13f560d024e936db074a68e65b07742daaeda4704ab14072a395c909a9a47c9351a
z0de5d95bbdc673b0162901f2f1e056caff8897dac1d9b58639069e1770b0115d3b5d03a50d6265
z7bd073c2fae82496c2abbb3cb374caa321d4bb0f675dd03e2d13d5d537d8615abbe8e7e4f11001
z0854544852193800632a498b9bdd07a12cf16692449de7feaa021bb2e5b313e232567c7397ea67
zfef2dc8b95f07b0be46bc46dda1ffa47a3d6d67555d86341eba7a47290e13410037a365b21cebd
zb61d9446f52a53feef9c221a2bb1c12ff91d59877ef58a8ed55aea6b99e3da41f12998787bcf6c
z9727feb265e5da4ce4ef83c3b1c960bd8050497460007afd3280cfe9f1cfe9ec40858734b5526c
z13d26afec6b5bbeac5046f4af6eac140258c446f36c6f95507b968feadc23ce7b1b8527afceb91
z39c6ed99158c81ff36d75ccc57be4213684c5769d4bff033dfa7d559c1f360219e9fd672c51c26
z843cb4824beb77adf62581571453a79e01c1fe5ac786fea4ed7f5888893aa333ab22066023bc66
z30b177bf22af997c7a29ba523de5f9c086dff51bb7105ae125adacd747a1c7a2cd38c85d76888e
z9a25ecc574fba7448f53eeef9946fe3deac2535bd5b61878252e0470d25981e0812e0078cdeaba
z1ab5f9e1b52cc41ad5b1650364f6ac7ea1849ecc2f42bbe5f7616d664abf534cf8a5f8ac1859e9
z6d6f1ed30b7b4d38e54d67492a564f7063a4d27e4e2ef7065ed90e4c4a3e0e5e6896f38b7b6c5b
z9011ef241152f4fb329a28036c2fbe98bbd2296343d514c4941872e6670da50721d4c94e7196b4
z5b83bef97c8fe1e05186dd15c7df3b6f24b241758fa3f0edce1d0ed43d0f2e565d9a3dd3b13501
z40ef8dca4b6256fc7604eed60fae74cb3a254175a1e0f18163e61c26dc97bff8ff06625d766d39
zd19ea3503a832468146287bc861f9f5c6be6c4da850f7ec4c175ecee56c00d22cbe8a34fb4fcc8
z80c838559b11ed60b38a1c074d2609f634ff5639b4c685897c136125fb6dd302e4ec98602516d4
z68bd243730422f46beccc83fa67585cd63405e3c193a85ca9affda84edbcff99047d82837536dc
zbb8616d664f6b23569667f6cd2bf9ed37e2ce214b7594719d78c411dacf26990118a395088a08a
zda32f2cf9a1ebf6a1d01cee2cec3e61756c7984935fb98453975d70a8e3d18fbac650a4532b132
zbab7d575f3d311105423f2401a557c2ab242cda4957827d2bfae0296429ea4c54a173b229afd6f
z43b884d32a87c257bd6ee37e141daf569fc25b08568cd246a466a7c4a6e0c803070737aabdb836
z5ed84990b32d687451fd55f580e22d798c9565fb58737974439057ba8f89e8ef4debcbdcff3a9c
z502b4b343f6c51dd47af45928b19022e6d14f3d4b1ad200a77a4f0a05bdd2f47b1fa37ac669efe
zb7a585ba15e8dad3443bc1d2cde306babe50a70c7acc6e6c71eba6574adc474da5c8ed8feb055e
z10d803af5bfa738eedf2b758ada3552d5d3f489ce86624158976b8dd2159c63f6c35c06d5cdf51
z13cd17a8e0dd29e7035b8a2ee38babc17d8721ff9dd84fc58515733df1e9129c3abc5a493bc055
z947d7a9cd779c7455c2af2470c240269c939b793a72df5c27b81c9f2e655883f02976e51b2069c
z59b99e5ddf8a364deaf8648975400e8b192508935316f8719fad6b678f9e0479145a231b09bfe1
za33317d8ac0dde4942c5c84b6ca8a7a4addf004e77e346c0d0c796ae35f1451e2bb47ae4061103
z2ad8417190cbeaa599a4ee4a854f66ee4f6b32586ec77b664a786d33910866fccd5ac1fbde90ea
zb9c5cad377ae0a81aca0020ebd96d8882088e52cf3b79b13f14adac9ba28fafff2f6a2b0df3a2d
z5b67536d89163f95013a3be553373083bb52a65104f9aa9385dcb96f3ff09a92accb4c8bdc0282
zdd951618af4e27df4f6edc8ecf814b71831581478dfb2712bfe0332f90968cac2eb469e9a30135
z3eb30b19f53cb2dbd9f66134c5091bc0bfdd020dfe18595b55e57790ec01b982730615a95b766e
z3aba003f5e548dbe1475ac509fae407e90ff3796962b4df447dc30b496f4cbe7c396b53fcf9adf
zd3f0cbfee7dfd21c24e96e76f18b9e92500f0f533420979ee518a3f027cae2ca21cfccfaa5eb1f
z5d1756178506005515e77c6157a03fbddf1a27aa42c23ce7c89b1e6e20755d7804409aeeb22de1
z1e7a8a4092b49aa1d89781c7cca7fe97077b6e17a93c89fc49081cee886a9fc8ed7f74a4871260
z5754fe457d2ccc18373fa887fa5165c656c6fb64cf55c38e90bfbd65c8b9738d34cf83a6059b95
z0b73ca5575a0a8696086ce07c2dce5bad3d5ab32acb4356faa2b73ae89589f1d170544bf65b39a
zdf08a03fcba2604c8eaf0855c26bc92a1f291c6a5015b8fa3365b3a54edae76f1a9745ba277aa9
zb3cfd96488584d4e6cf76b3c2deb53d32305f577c4b9dca201af7d038b0e0906a2898fc96ea48e
z5449f49814a4739e585af5e32ab45d771c2d47cd95d018671f35b243249ab8350d5eb6ca18a974
z210b9bef8d019d710556621b7f18712dd088a6b6fb2fa16dc4ea14c156a6874beff2bb0b10139b
z3a57cabdcc0f41da1f7bef4c8dc469e5de271e815d50be7a798602376349b3e377b5fdd891c804
z26817ccb5f26c33d61db198d4e7f3077896b3678f3821eb02ee1e656c24f0bf3d650fd1bd1808d
z3bea9ee52b65ee0d3dca191a728a19432957a858a5b1506dcd62b0775c544a7f56949d6d7d2914
z89ab9db50dc1b84bcfbe68e6c7b58cc25dda7d6f507fad823b80cb448f4f8576560f9f1449c7b1
z75167df86ecaf080d6306c1ec1fa6a7b164e3eea7c39ab1adb0334005be64808a3dbb08301d824
z20a36ebca29e3727ede0d644f399dc34e8811d65c5cf1eb659573d8c97d71ace43060f0cb7c316
zcfd866837d07d5fb56180042d5866aa3db4d97d4ddd4f1d4081f9ba171e4b05c9d60ba0e4272ad
z6010874f7668d23cc583e256a9524b9f817e66509347ee332388fe19d2ed501698bfe81f717671
zb7aff0894273a5e14a713f581afb1308c6b34633f5449ff1f01543c68ebd6796ccddf48a5023fb
z7d347172688dd61ee0ab9e2a0064a12de115329297f7684133ad31862d1deca816f715d1ca6f2a
zb49d2275fe4c7b8022db5a379b1dc28b5dce3ae004dda6fe6077f0cf7a545cd58e4455b106b600
za02099a73f60b00c335c81e51673a8045b7e8546e5e0998303727e6d5efb5c5480fac0abde29bc
z704391efed655628526cddb68ea626f4dfc3a692bfa8df12ef378849b052725af87e533f0e48b2
z97f6a15e56a5f269d256da0451d6d5018b2cb4d6e208284676ffabc2b2ad71d5df28417b08ceee
z5ddfff72190a06be63939f745edd07b8997f6f4a8a683850a9c2ad9280f5246fa31327db0ee107
ze32d09dee0a04edbc72302bef0b9fceedd48a5b0c1ba8f7a52a2d823724d4fcd5c42c49aa8ef47
z703cd5db7c6561ee13bd9e988480619cecef28370d88f0e2579ac83dc60c85fd0d0d4a681a510d
z1baa64a2edeee862871e431bd7a0d97d9c6c7d7ed6caef5acf7591c97a8c7cc2187e13669ef8d4
z8f28c9d810c6c67f4338fe2a0d76b9aa8092617144ff9592324685dbcd259860701d56cd29372a
z9a657164b6c5205f046156260db6357437ca094cc07dc92d4223de5244650a12e52b914ccd98b3
z337ba17a3910f38380fa6de680d2895689928383ac22e402a6e18bf831591fd50d101948079c96
za88e56e0e6b9cdf79c5e24039b3a6f3ba9c2a4674886b61b4e2f077e01e15851a5841332c3ddb9
z49db39049d1bb01643989fab7ec6a2de4d100f34d126e531a71fd79c352f258159002c9cbb3d68
zf03cb51429be9d2b544be590d608166f8f34fc62527039b8807fde3c9bd2a82d6d2c215440bfc4
z5e0b806ecf2eae4dcce582199d6826d284c6061924220f44392e72a3e9e6b3cc8eb2497359a06d
zff2d93edd984802a2fb9527499b0e5c93ca7c2eb4f017190da7e8da2a2d786e6908658a707ce92
z6c29c478b58847803639fa724a7fb81b73bfe326c752472c3a3123936efde2629ecb3321b5fef4
zf33a44a21dcc5a5a8df125d3af3954a45a16221abd2d2aa17b4c759fcc34d9d1888dd15a99a5bd
z75420511c1b80d83ae60022c602dc7e13d2335bff97338b533d3363d27eee276f7272f49e0fd83
z5fa24b7c07e8c57db159d36c55ced29891888e2f6d8697d5036e3ccdf8023baef2462c7154222e
z8f11a5dc931a5f0ba1862a0099fbd97283ba6fd2859341c3bba05548f5702cba384d29a9e3ff77
z4740bdb893e916337a7929b71df000789f82d7c24cfb369fd1e5419524480f65339075474d63d8
zd43310d9cd0bf050dc8e9691b71e4a5508972d39f01dbfcdbfd38c309b7ed2317edf8eab2d017f
zf06db89c744b78f3bb2f4e163910134d63048f04589b82f706331a889f92b8f4256390430e8fec
z5e2d3edf1324e4be1e5dc7aa5f3838babbcdf9a50c4d80322aa59235083de59f61026b18365501
z16a74c9962fa04311a678b69d93e891e410d3a929461630e4cea2c9f7a8f224c66ce20cc0805ad
z30e848b6754e2a19e67e421dd4aff353c44d151d460a6c24b111aca4820177ef86fa092b6785bb
ze8393233f24dc6a6e2ce828b8a8ac20d573a5e541f468bf8f21b77e62f4323bdef156692786b33
zccba02bfbd21810eef6075b0a2217fa15fc5c9d62e3898783c54bba8204c2ea8580c11d710b95c
z8be226f117ef7d85bd2501884b25989631ca159ae08a71099d2b45224a2a5d5834c641363b115c
zd5a85d9473085388b5415fd27009f417fef9f5e238ac4add600e1f202f2ea47dd4bb9fc89a3292
zf0adcdbc6276eaff57bddc9474eaffb384abd5e1b9c64cd122482ff384ed84b63b7618edd3a3b8
z10c11f90a51b09ac1c9913e9bf912bd2a8965381bd49822936ecee4be21bf46d9b1f91ac20a8b9
zca0033809ea7ba7503bad97aaefe79feda750947785df29ca9881140c180ced4a36b5b5fcf492f
z6df80abca994ee957e9ac9a9f68d27438578bb95d036d26f5f45e8adbe1c009d9934ef217dd7ad
zca392a395082a8434ddeb796d59038f907c7ed9aaa2944bda4976f50004f2a86b34f05018016ed
z80b26f686bdecd94be3d4e1b3c6f534d175977ff8e669e362176cc1db63875031cf8aca1ff2e36
z435786bf2a6ee13388755c1269fc8886cc6dff248e9650b8e21449e4d8624a5978ec843d2b03c5
zb66f01f899fdb13842794d464a460cb09df0be744b81736e56f8062cb775985161ffb4f653b0af
zb1acaee2d2a603abefa00b71b1e864dedf10c4235b5d26425bc7d54eeeb809379df7ff04253d61
zdd7e61219979f2b711e6474aef247b2c89f199736de83492d8ce3b935c8dd7effab977a792e38b
zff1a3c12ac70f591e272e4debe6910b5cf890d278eb44ff443566216d2f69c3007ceaa8785d28e
z01ead994d974b77b6ad9e15f688d31fb830cbd16c17f91692b0650a8312262c7e2093a601fc734
z0e2c7fb6975592536170e590be04dc0dfc743f23c026e95da14d4f6f1754fdf9f66875d7f574d0
z23b2db80c5604cfb2c88043418281feb77b5d0c63869786132c6ce41ac59b4d1118599d92053a8
z68b5e719acd38c32ef37b8f59e93595b6e7e11d36ae21ff8b90568f40aab46c57a127e1d39c44f
z83c5b46bda828b414532c3110a35633083e9a70600aed0c57d4226f453df0d7809a060b67e77b8
z5249ece8eff1f740ef225083463c5a106a7f75e5fa8ef6c154f257987607c2daeb90fcf339d7ab
z16719f480c5033a86d7adf1b44d20f910f9aafb089b60f9caad9309dc5599350f9fe526965cdb7
z811fbf7a1a6355bda0ef347b7a7d8eeb96367ecf5b90fcd45eb979dbbf026e3e284df1caeff132
ze3f7adf8f235dd0694911681425f28746fde0589f0155be5d8979d77bf8aa73731653320fd4ca6
zb272615fd0d2acb29c6cf823cf3c3e6a79bc70532b8c208b660aa5d6a9a246115c3ac4ab61ce5d
zd3fc58dc17d9e2d641a80b8661c4826660fcc02c969702f9ed3c8fa7ca3f5ba3e1b0a42ce2c66d
z4cf70a6b98e7984f663585872c8231bef9c6b2188bfaf3f7b0d7381e0ba19b7c7741d6fd3b38bd
z8f23e7574ef15877d6838c30b81a2b6fc8ba0d67ebc2385ef5f810b80e496e20ac25c3897c91f7
z6e30f9a4c69c685d626871e93dc3a464c51602d490179ad71df7f3644f993d30e7abe1a5246bdf
z44206e72947e3eec246778986895ebd25ab3e69c1acd90892046e6e58c21aa6f5305c67117b7da
z1fa24bce798985f3c0141c60dcde3bad4597afc7f0367020e197655ef144d1888947df50087aeb
z5728f486aac4d552c20157976c17e1a23025af359a3cbe9698489ac72e8d799363aea13318b388
z83cd22cbdcd327a0de965cf745485ec758ced29d1ae0dc7ca1644114531c205698981a4b47b15d
z7d8664d5b9065e068a61b28e57bc4a403d80268e4ee2cebde09ac6c89e68f0bbdf0414bdff125d
zda6acb6323647e60c3528038604541393d5f61f53e74c19daefb2bb1c6ee293f9c739638332008
z379b34c4de06106c63e1c93cb4085a56ac0d7f793deb970ac6499862134dc1beb91a01821fd03c
ze25ac9aee759a48decf4770612628ddfe2b2d2e2b3ffd7f7f1c3c436fb9413190df756e6977177
z3d2b2c55a2592beb5c56a3b53379909b65c36b7e0f76a79c85bdd64d5d22853758869c3a88eb1f
z90e45450957e8ee28c0d0938e9c41b0e9595d949c1c6de352c34d1013064a96c469a6bd869a5fd
z22aead2877c20b991b861efcdaf3ffd9c44a2ee02c1656efb9eac5d70233b4e51243eb92037fba
z209cdd598a071778611c6c6aac18fbbe0f8ba4c852cc8701f4ba9256f4d288f636463a52f0c4ba
z5213d6ce14d50a609a14c92e86741727a74b63a07bb97ead0a6d58649ba1c8ede9a1f9806ccb35
z32cabd8f85ff4bc1de78ed8979b1054a6af18a3c1624fe5f92bda9190f1ce5484d4cedc01483ae
z30e9a43b90d84fc6f63cc9ee4f02f2770fdb3cd00e9bc62b213209e7b8dd5e66754296e7247095
zbb75b2b81e2399e6d519a903e5833866fd1c4d1a94d929114e1dc09b35d48250f9cd2a18562c3c
z9a9d7bf5ec26291d421a01339efd51cb6115c623272912638652028ee8c19618b3f37a46054473
za0bf1053e169a8d6d1e0e4351792cc7739e854b51a12150ce8976b3ba9182d982745f45e31b607
zd4f6412c77eeccce0c8af3c9ee4eec08f388f7554163d41ebb3746e291f4ebe73fe023fded08b5
zfb5a47a9e258e0c0b18718948f84dbe6b10bfd9b81b293c4680a4ebeb1b8d9a6e6d1ce9686e746
z4243fb58b00013a97fc853130a92197aac01c4d544848468909ce8c0419612a591b0220a28d026
z40ecec06a65109470cb6f746167cf961bde04d0888358468498df4024a4899fc2458e2282a519a
z600caf089f896dec8eac5faee57c6ed42b57c938e5f5e9305b6259d73bca2eec7251ef0a41dc4b
zca20c3f2374d19398dacafdbcda9fc2ac6b909c450aa658eca27ed3d30f95ba881d847be91d605
ze72a41f979524696f5e54de79f58b64a0ca6e9286d74c3f007d2431223963ee3918bda1a9a02c6
za0461ab68c792456e5ced615818f5cf2ad0e7c52ad7c3a725a7171965df65b98d0e8c009768a28
zf3afd69b43986013f7ebd208afbffe5b7267346fb8d09def15388fd9959c492afdd31250ad06fa
z96a59d6f4493763c9c09b4b231cc49ddfd994fbd48480e844d2a4e753583424daeb7f4020647ec
z67cbb984f0c216527a7ca1385492b347d52b5220895b152dac7c47b797efdd49f4790263f93394
zba7ae252a5a73c150f241b03a70cc96749cd5aba2a1e8256954a1e3d4245e49203477f18fa52e7
za123e527e3d3678287dfdadf5a5eb5597fb8218838ede2f5eb2361336aab269f8620fad1481c08
zdf7ee116bfea48abfe0a6083520ac810e1a93cff89e28141c3126229850ebeda44007cda736d09
z11a696ff9ae144b7a7dd4aa3d4f19b864be3d8f81c7bff3d4392744da9fcf25fc0837f007670be
zc36731b0808c7c7763608f66a8a8ba85ec0c6424760cfbcc43afbae03588d88ef3b3db117af07e
z976f88a3e269fa08f2d50b4f59e4a9271a0c7f6368f1ee7eadb03eb72ba4922b3fda72cb236f52
zd2364fc82b1fe07d73a8a166ccbdb183913f1605a5990db7c08c3d0e04ed717b7a59a9f2e3d089
z62fb147bf88831e904ed8aae619f6d9a976ba1a63c53ce09d56cc9a35146091b5c6d25eaf1f1fc
z969f4aafc7cee5ca3c33aacbc575f4b3857d87a77f7b73c5001c8fe843d8d74d6406ca7a1ab776
zd9db3144a06377f697d43fc713d0f44a1499a74404b090905e36ecbd10f24e5405bc182f87e6e0
zda31d826d14147fad1ef65c8851505454dabef26eb8cdb718b60a0c2ec05905cd51b34b25c3b0e
z0da05ba9fe2916ad483c7f0a9f7ad622c8c39b346138b7365f40d334a2ed6e653af75b72335d6b
zbf475c7585df12cb967ee4b604461acc25041f76c079de4e347a1feac549fa2908179c7437e895
zd292692b97be5fde4763eda8d0dbf2d5664cbd6c93f387b6e79d99dc6bcda2bc0f02ce07a00933
zace09e8271b95df8c1922e5c51f0e157c17bcb3f37295bec1230d8c7ff350dd615cf680bf576a8
ze7f923d3917684a55b2dc24510cf92ccb9d7d3476c13dee69855300bde697ad0a819484be3b14f
z94b7fb8dfd6705f2f9e16aa07e390f61317c2c6db035bf1acbd52c466c2485136722a8761be927
ze2d6b4d0b48c21bddd9e050d6bc70827f6ec1754a9dbb88e2b2b3be2e4892ce784c6cef8c5631c
z8545c93ceccf743ebd63c5964f03db746f14882ee05a19433b8606257b9858504ac33d04e2ed10
zcd53a76c767ce386a4268c0571a20484aa451a5bd5fd0e63b5ce82399a5c723b22ab9c1a8c2add
z797b4245d6be39757f22d0370fc70661dfc88ca36d66c3f8fe5929e5aad742dc58d4d2910e2383
zb78d8d190e6d176a0d9f5c1d09ea4fabfa1ec4b559865d6e89e653cacb4a966058278a13916fa5
zd0b80aa61cc7e921f69062334cb4bad2eafc82a53cc2179f6bbff6e5057fea84ae2a3f2b9c46db
zad3beb4f75132cd452b8281f336b1d7f420583ef929de2d78eb77b41aa62d29087613b7904cb49
z446d7f502e9042adf2aea1e0bc5fca6442893bcb864b904b9a90f3253ace4a6903311609364683
z6e88922a8ea40ded4d5caf83cbf501595d8a3fbdb9f3270503f7a887a97c3b17f0afbc419463c7
z017d29636d3d8ea9299ea7c5fb023398b95e5f964c79f9141b94ef2f820568173fdc2b72de2ad3
zb5fc36324e4730c00b45c7414c407b855d427caacd177b34b4ec996c6181e1176cb89c65759c8e
z844f39b5c6506551957d1bef5c3372bc0c668698a3d8852a9793da22e3d7684a9fa1ab7ecc1b1e
z5a66d5cee95785493402b78492ce3d6e03f2241e641fb918b80b8d67fddd697a9349dd9107448a
z638352d72a5246a62232c21160db687397a82caaac60f63a9a99a8e651a072ddc09bf434be5c43
zbe05fe89e21bd6f2b099ab28589a7ae829c9e6f183bf68ed5243293169152cb75e0136aa349464
z46fd93c614804a8c568fc56376e8b0de9570c44a38b47624b6df7b4f488679c770cf69e499fa86
za1091d6d8fa5629ce8a6aee144e3e8e2c36b187d02c91700c75d40901883703a7489eb315e51b7
z64b7799af73b9a03836247288c6a159ea5af8070383f19234988de05ce7c15d64b53bf8ad3d3d6
z6c1dcb89aadec29024e158847bb4fac738970daaea4df92b852163cc6185142282d317555ebafa
z2c920a2cff28714374b3f408fc6e01b5e0d3e8fbcff81d536ede6a547507d3350f83c08e3aca69
zd419d8585fffdd655095fb6acde8f673d6b3ef29e60ec188d119cb7d37d33672a7488acfa0eeff
zc0208620a7b99bb596832321db3efa9d0f7b63f3b0db094acd480bcb52ce3a3f0db58a45cce435
z5b72678d0202d9dd1d9c8dd3190ff97fc921324bc3ee7a569ee6b0a947c04b10a28851f96df249
z0e78d4afeb4fdd3806b636aa86611e75b1a7e5a6c74bc76f09af72dfe40a9a7f489a36b0f89075
zefee0d841b1d7d6076f04e753b7b2cf3927e5f4a22c545e121ce0c5979140ece1e66053b787b15
z8298702c3386cfaa91321a98100b48d43258f36ffeddc13dc31f21008756013757f8712cac5c31
z906405a3fc5667c98ac569bf4163d03ea65d058d7093cdda76d488eb956c743c3c43c0c34d389f
zfc8026dba1c48f3ad6ec495f43f5424fdf7121717ea8014a55e805560ea8f6f52dbf872c18cd1f
z7103b6262b13616b4e53223dfafac36845ac6ba751dc8cb78c027a6915c8cff69a8b8db3646390
z4090b304e227cf7ed12c075f4c30564d097a4f3a373d45d16df6f7d7efa9f00cfed6d51b77cd30
zda2c52008bdb51aa40572e673b0de0a17bbc798882fe6b685129b1a6d2acc4c43ccde887e024cd
z73d945448afb2ef7d67250a0e8de53ec7d3c296cac8f5f03ddd7fc98342ffd222c6e9c5e8d326f
z33790c30b351b32a45a7524ea814181f4c6b9c43d2b00543616e2c109b45ed8a0e5aede15d8af6
z5920a985a0cc32fd921114f00b3272abb9f21ee416c412c07e58d87ac99d1b98b5e585fe1e7a15
zf92c23c709ac0bdb5314c090600b825a60ba0d8b6f1e734b079e80259ceab7e3ee163583eb9413
z7b83c34b34920e1daf06520698ab576fe6e0921821f584313ffa95c6de72313beecbd2313532b3
zb02dd3ca44609078a78e18fd37afba4a21d0ccb084774a9d7c275bb387c28faba2f7076460f264
zd45e1641ae82e9a5e8c738ee6c9d1bfd3015d7ad60bd4c423369d7de4b1379e2c7f93cb443d59b
z2a0693ffb91eeb20d7d1884c5f931e2700bf132273c4eba7daef78fb55a49da0c829e3c4f6b52d
z1c1562df2688864ad674fb4b69720aab35dc1d7d076dd8ff16fdf6567af1e2cb053a746f35f249
zd3f6f4ea503715488bc66f53575d931abf6ef19d3c8e099fa156cfd87ce2ac8b2f6f867089f996
z3b50dda54df50204b9e06a466b5301e342a1031c0a018b1da2c2e667bf46dc2a94c7eafb282271
z29cb55edc5a3b103a353820c1bbdfcf40c28274b10c2475c498a4314c1e8e8acefe92af40fd373
z7c2654f5a84f47f87b7d53bc2b1ee2aca898c88ee8a52754d3c79168ad02125ca4c9ce0594c176
z9828b439de6f32d6aa36dfdf4235cef93743466bcf1f5efa8096d4f73417834dd931328cf1c060
zf05ec7772c3d13081a70d414887d060ef5b461734ad4168d61e9a0fbb5a8d2e324e228df41fcd6
z4e747c2d6e2f0eb9f7b4dc2ff8abb4159abd32a839adf237c9db609981c1f4c79ea1432834b54f
z0406c158640f17d6f9530c2c27beace0fd24e4a6ee197964944e58801a108b46fc869b112a31c7
zfc4cba73be15891ccbbf5bff8454be70257a5b1be0e0bbd2561cb7ee21a1b07a49a45143866c2b
z2c00b5b64dafbecf93f1bfab4c5e7547bdc2402c8dfb324d22f7b0a32fc33d9fec514dd83ed959
zfc070cf93cd455df3a898e421bee9a39676cebf2e1c18eede19f610b6d6202660aca7ef16ccb48
z3347ebc7dedca5b1bc8e1383062076afdc07af1ba68b64247cd2555eafbb28cb124b8b4ff2f133
z68fc61b97b03245ee096ff8a3c108450291f8aaa3b024369cad8ca4b62b68dd3f84ab818da60ee
z3249d4ca692c55937380fa243fe2d4b3b0a038369f8c137ed5682cba489021933c03081aa72e75
z4762ee1ae9b41dc8f5ba115d6cc3762d9502cc8f2e4f504d1e7c3ac7e9e2e1f6a499c0ccc52d42
zccce797f48cb2c1eaa105f300bc78d928c9d7828f3d2471175dc3b9463a423674ce708dc611708
zb6e5f566bc7ccb00c6988f92028ce17620fd8e2a2a8d25afda42f2b1bf96644e532fb7c753b8b1
z017ccd3d825a07057224ac1d89c94d52cc4d9467f2126cb7da9e0d92622cf13c6124d980828207
zd9fe255664d493bbc8874766ebe8c31b4b9a3437eabb08b756a6a2a7c279aa99c426f53f21bde7
z421ebc738ffffc948f5333fd0308ab9cd7b1ded86a04b164a5820cc03c7fe2107380453689f1cb
z1ac3e42c85198e5438a68f9a940f2984d29b730d68e862b0c5c55b2dfd8a6104a521ac926f6db1
z592bf92409d4ed6ab16d67691b2c186a61aa5bf1f06446f17bdd49e6bdfb0cfd16e39fe8205169
z064c299a02c8e9f7293dc2ac0f15b8d3ba526458dbc671a527b081701eb736075b7d4dbc47e1a8
zb2947039de3ca0800e2a365c6ac8516da8646d939352185e645835efb3f17be2d169a64a472440
zf86fab82172dc86aafe0e2b5ae0059b8e84b88146d1a3d9d7646b5e3ed368b3661b9bd51a8dca3
zdfde7fc7fade66abdd4b2f9105daf546ab0f938b95d579e2521589b6826599eb89a9559adda28a
zea42714c4b94891d52594cb3371f17804fda194f44ab50f326808e025650b035b5282a96a6b57a
z33913126d3307c00c4fec04129bfa29301a98786831f4f86dbc1b20a22bc6a8f76b3be8cbb59a1
z376eb85d7721a6a9d0c8c1ab0bdc5b653200502dba5c44117b90d4679b4e22279056c510a9cdd5
zeac20e794238229577fe9900404d6a35fa36d719d36771ef7767f9c8dc36fa57719a96a5a8e595
z18a9d67153cea00fc5b46795381ac51a99c006aa488d52750cfe03739c01236a74cbc2e6791dc5
z8d861d1e419b0ac2be1e00a92e134ab8880f4780654440d4db06b41ec4c275aab440fee7c2a68d
z314ce26ec65406aedb7321a379777bdd64f9ecb31c0ef4ecd56d1df679cb55c6175569daaa2c4d
zaed57fee77f4b5d59c56a9e41fed25d265d1e9136f994c26a772eb0fd37fa054ad6b326a824c67
z47c7541e3e731e3d3652298d8b42b18857892241b294a95dc7062aae837060aac940eaa694a731
z1f72cab0bd65cd7e1da4196c80065c59f742549dba85b644b8c98fc1c1107d9bc2ee64de67b412
zb3a47c07438b734656405c2d03183949236db3536f1004837808b35dac8206ea93d36f9b3c9864
z8f7f99897e6a9664b7c4a187826b7c0c958dccae59a84208d492b394007a3b50de490bd945ee3a
ze63cb364c1f64c8b6c7cec940409ff46219779b566408699557d7f2e6d5f2e72908f091a833b55
z633bd9eaf1e25c59fb0cf5268a2ec15e08d5ae1221ce17fdd168ada2a872c93d5892b29f1e4e10
z1c692ceff8466ef752b3d3ac1e05608a4a49246462ebcf6f80717e258467cfa4cf517bb4484549
z1375154282cddd2c0be9aa804c1ee9dfbe58a7798ad808adb751ab81629d556aaf7b12d18dfa16
z6a2ad3775843fc15dc013824f9da6e806596d3580d877d9d70674bf46cbce612e714a64ef2d4fd
zaccd7877a30a8c340fdd3e2bf93b8a4257bdc970e4f532be49563fafce8cf38ced803a6dca7c4f
z87592037bc5bc8b5dbf3393578efb56758b5ed47b6b28a8dfeb020112e7bf80f86462fa373ae70
z455cdad06514dd069267aac946c6c3fd55989af9b8b32d6fbb5d74fc21c94633115ba2cfdb926a
z60605bd548cccd71a00321b2e608e84da76d76a071b97f805823634978cb2366682b7192a8c28a
z250bf68e47da52d161379d4919e8d6c8faf567569ffc278526c900e97a7e9c1f048d43279b03a9
z941cff93069ff557f885704806fa7b6d0cad8ace2e8ac59b2febdc5efa9bdd94ba1f75588cc46b
z0b0ca904f9d2aff74e6ea839dce14686c7aa37a21f01e44a46f574a2f5c8ad323efc1431b470e8
z9c2fe4ba23d1fac54a844ed83102d3fcf13191f932be9461c2632f5cd42750209c6f425f7f68c4
z9627d97ec1db8e230567fd081ef65d57c4dfbf5458093487608d2de7765ddd76b59c1bc0dbf539
zfa37c3c30babd440398d20f98106b25da6cf3a59f84d410fc95af80954f1490d91dc4ea6c781e4
ze34a79a648bc43c25b2c7f3eedb95ef68a369c0de930528e77d039f57672b9d123d31a1bb9daf1
z7ba44c0eca3583109d107a63aa3be6221d858ed3ee9d60b710d03d81528f22bb1751e11b69d7c9
zd9c11863938cb3eb109770698add4fb6525f943d6a0be87e81c602107a4a8a0c2a6a54e464ce37
zeb6d3911ecab01661b68f913eb1c32b7292f60c070e508d4c0e5e7d1bae04d7cbe8f2cb0232877
z58f913e7bdede6b42d81f081523ed0a8d0246d1d94f060aad371dd6f92cb93e6f71e6fbfc2b2f1
z48371ab669b15ed6c37b98041a62ad7400028da02c5c2c661a39de4eeca351dd54b33c626cf20f
zf08e7c467fd4518f6d29e0727b530aa2e928a00d125293b4d0ba053f8e85cf76ba59cc01a02b5f
z1325c3fc85a2105be3e0a74bf3950af640c16cad8f376be678326aa4a9a18b3f9e5352d920bce0
z9bf6a0991092346e74ef037316eea453fa3fa1f833f23feac099de50cd784145a54699a7a4ee27
z0d6f7097991c5568e8f26827c871cae07199304d950e1df77699f82aff6f7f2a1822e60754d8a8
z08522eb068a1c7d111777f3a00db8945cc90c3ce9aec92badf7a96859b1b35db541d2c005cedda
za3306e85d0dbd002461f4cf85639768cb91a5a3092f0d6228e1ab057218a14088494ea6521a665
z89bc8c31d947864cf6253bec52e7a18cc3d13b45acd285894ef97a0d77bbda77cdc74d4f8ff776
zc5bbe64ad9854c6c782d823f3783610d614376095b45d7847f307377b10a0076469d95973f5896
zad476b261d48cded184789c6cbe944bf61369a4f0268f2e19bc5e6b3fa0bc79114298ca99061f2
z67d20f653cf7b7abe3199e6c87c1e72eaf1ae186a11f9f0993220e820f96ed710f58b760d2e619
zb1881b874a2d788b333237bc8755fc42516fa39b9904dd9133087b078396b06f3c2490c468380d
z26676ab05b2cd90b72a4f283f3d7d453feedc73a99f7d82b585d28021ff61424ecd2ddc4605a72
z530a4487fa1f4b19f9505c970a2d0c229f2cd24e8afd7c1c69eea3e35b5722ecbef7682647fb20
z262e7c5c2daa876f10425351278b297d138dbf37e8a3c108cfa317bac1adc6218e66a4a115959b
z6e1e6c7189743776053e7cba2976c8dc2c440621b1417488956a95fb057ed56a83123bda4c0939
zb28548a1ea01a311cf7e422509500e73ae599d0d6ace77a6f60eabe377eacac8cc05158c6fc51a
ze83f641079c28a1f963963a904e99c0dda6a9ea912191aefce3abf11ba0848c96f9f4aa572e93e
za1cd211dfa4f53293d82568aba077eefc87c68df7f63c34b0e9ac8635c3d28a429612ea3062f1e
zd3efa74ecc648cb9261e2dfad812750b27ac8718e74876438f597ad13f23553037287671cd1de7
z45e6547b18ebeb2ff9031b469e0e84f2541566f8fe0f66c04351b0683f92865d53727af833edce
z845bdbef80f8db20c94f83a5adfb4db97d269d626f59b544767cf72b711f9c734d6835cd3a3656
z97d7e728c8d56b4df7931b12b4400ab65c66d3aa0eeeb65bc7d13bb3d749de72a5cfae3739b1eb
z08b463230e0cab555c38a95a1492e63d0ca4858293751f4a1abd63eea2a7e345493cbbb746e390
z468fa2331fc4815e9b46cee251505517d75a892d3bc0dd0aa78145023b2381e3f8f64d3aa08a9e
z5bff458b3b17676a9e997987a773cebc6f582786fd131ae121e747c2b4698483892d26327fe3e9
zae1103600183f75f33c08d94b089c801bbf27063585d1f0b7c387f6bd6511b41b38aeab3ea6493
z70e923f1026ac9f18e10c033871553a413956468651182ec3142035957fa4b1e79f2ebe73276f1
z8bd516e3c102c5c54eed57c8d0fd6a174f65a328e4f4bada8e6394a832286fc922d1ecfb61311a
z1b8a2556758877c6edd5def91483b50189c296d6dc5d3ff71f120aa2d68706d7a53c25860bb5c1
zdacc68a12fa85b4c21bfd7138d340023631d9edb094e12a60a056c51cd1cbd393dab097d5ae428
zc4c938ea73c8b1fb6e4a8d0794b55ad858bb64e2d03d5d9ea4aed8764a9aada24e4b845c45da6a
z7c5345426de562ccdc77f96538742662bac0ea24105e270eefd1171e07e7c71a6ecccaa2452cdd
z4853b983abc25bd9efc3020df7baa233122ee649e9074c8d9400eea002c73b57157ea562e921ca
z2f755545dd9713a73369429447bfa6ce82847585cb3ddf91a5078c2fff39c171ff53c4a6a8369e
za477823b4217aece07cbfed0b9f36950c293637ff788f99efb9ad79cf80b2b2bd37caeecfc74b7
z29086a76dd101ee14a1c298c6ac65397c59b2db602c3de4a94ee591806145568ab06a6763301f3
z113cd78ff21ba2d6d9f2caddb384054985636b1cb9b8dc3a3aed5fcd58e22049869eb887b4d017
z5ac081c11681752348d4ec333a3636bdb72d065cca2e21919c439e7e75a189d94beb8dbf2b1c27
z4f479ad006afcc86a80586ac8c567a629f3cf6009683c2f49b318ef928f13a912de6fae04eba7d
zc550b1f5f63eaa15e3eb0db3de553959796f6766c9f3a17374dc6ba98fd5f9f964f1084bf80a2b
z865507340675a877fc06d8145263b7e8279c9fc6d4faae7d54d8f1c07ef30adb3cf156319fc4b6
ze14f42a5ba664d589c6acdbe7f0b10a57ec572e57c10870af9b453a5a64899d6824fa4d124025f
z707c3c003c05cdd2d5f6217e65e067672851ce5bf23fc7724d68fd718638b6304e061534a7c5b4
z134fd9dbbc05c721409649063823209c7082b3a237d1f155fb4f2e0d50f2a23ed7eac62080f364
zea338e930ae653c98f0e0cb76e1e6e7683d8fc41fc9533162a4655cc77c075ab1c2200ea176d95
z2ef10c3ff57d93d9dd667db5328a2f8c49d88e3952d92038ba9528a28e8d574d7d98205795a62f
z1debc513413f4482b2ce3b13f46e86364f930f783f9124712e8bdf008b5c6930fa6f2828f5fb81
z9155b41703ed039a8d761523f28dc2afd9e1c59ebe01a62c0353828a6aa26d7486e8b6732e4915
z921f9816f05a22549f03668191ee12ad18ca52506b4733671953f210bda13775d9ddee5817c3a5
z51d4b8dc7543c4f547be1195a0cb4669bcfa570f66684ef1d6cf7d9565584c6d0513ecd510555d
z9f894d15a94b92d37a93c89e8bfb471e477ba3d530c87fb862c742644797412d97c18cf72689f5
zc821f1aa0165a440afb6391c9dc1839d8b5cf02554747fc76e66437cecec458c6ddbccc19cade3
z4eee0a3efe75fd4a952e350e9f0952eb427ae97f91231330b9d48fec7b6e5ab351cda87924c894
ze033a527aca36dc1c7e15351129887c524616e51c26ff2fb35b2c82ffd7a45019fd2d268e28468
z59eb6f5ed92cb4414e8358ab491677bc858add219de2bca1ed1004f189c2ab0ce3fe39bb4ca53c
za0263c247115a4138bb504218c97a6e329a54f2561d3078314eaa62c175a66d0192f2e6d49afec
z5f2155d853248a6077675cb8ba7469f2f2867641d77c42d472288d814960046c3bd3d73ddf6a4a
z4e25b9b4a18eeefad61ec8189a5d9b71bc2933863b0fef0b57d5a034336c3569e40f2c7b8d7aa0
ze6f7cc676d1248f6963a57ac84e950b6dc4127d1b02d8ed231b43a44f142d3b9fc0fde4f24d2b4
zc40b89c0bc4b9ec1984a31d5361a3b27d2053738e63c140a6fcd68085d908b3bf2ff986418ef82
z6ff4cf9969ee47023c732121f03502fe45c09a4aae3892af5d2d0f567e78f633aff52abf36beb7
z74f8219b036dfb4018da63ca798cf32efd768e3a6a6f3f15a28c014935ec3d0a12e84eaae0a35f
z296cd703232194d333c483b94e052b7f207e102e6ee838258b0e806d1b7fe247637e8d0d47475b
zff41fc5599bbfe68e527e98016ca9e6a327eeaa4eed24bbd118f330320f25dade83efec73f7e53
z2d2dacc7f3f6b81c0e2b5011ffae316f9a3be0fb2f1f31e97f86ec1f7bcfc9462c6b147382c348
z70d738d3435e097bb1197bb46a486158a4584ab06f06a6a4e4e8d10751e6805d9eade62e176e24
z51b67219a88d2ac0ceef0f7cdc1b1b0ce9ec02d578864bf8f2b659ef2f42cb23e775a3644df464
z816b7b2b6c027af08a0b2d15cf4941a28829711f57143ccc5d3082643372000e59051ac5c8dc91
z3b80dc3f09357b417d1941f8691dd0bfa93094ecfc93dac3824bd03b2232eea4cc919889a55843
z5984264dedd4092bc0435ed69a6b851359f3a4495815a63dcac11de2db628b1a7fe7c2851ed3f4
zcae23c0075a6ff804cd7a74406015b640aa50206b1a1511c47e19e1f82bd0db7f8629e5a3a9e25
za3720e101da7e00b671f99a3788271d93ac25e3993b68ac9c4a835ed5376a80de6b55fb52d31ae
z8ffbcc5814e539cdb582b2eeac468e693bd3e4db3c6216824675dbfaa250ea1959933bb07a1598
zb28419453d20aa3dfc2997ac93b66ba778e2c07716b00e57b1ad5ba2f60bcf7afc231a0c01d5ce
zac2ebd361450c187f77660df3714840d0b480f4365b42f829dd3e25bf38f7bf3e34917a5d468a3
z25fdd231049471cccdabed9fb79853b50e6b80af684fb60418f322e91d7348c57e2c9ec81674be
z1c6abd67d99e1c8d12776d20608edc6d18c8beebed87223414c3f22522bb66ce708ac91bad1d1c
z0de568275db70117ac1167b3663b5b84547468fefc1d73dd98e857dbe169c5ecfc2bb7dae1ce0b
z7cba7c10ffa88a4c21ef8fd554d259088c848a1a05c5adcbcb5bf8d86bd154af18c89072225ee3
zb2e7086a4f28f3bef961c86f232761d0e89c3a02cc283ad68ce030d96b993f1504a6d2fdb01ce9
z8dea950939269a07fb779264ffca6821fe75aab2187387ab170bd5c93e5dbc46bce9953d53973d
z91997ab88fc922e494892f1741b5272432757d7df5ddb7768b46c4fe8ffdce392432c32f59c3bc
z6880af032159d01fafaf0a1eb30896b4e4fbbcd086bdb6e1d58467ae2a1bd91a33b1e72aed77e2
zded6b1ffada70497117e2a75fbcace2e6c2e61aed670144dfd38167ccfc8aebc5fb432674b0a3a
z229efa588460a66cee463ecb24e0de4fe6fbe630ed53be5c43c4b625805f8717dc68f62ac555bf
zc6f4d66a308f81982048b9f8cbfce7c3267083f97cb6c39ab054b83a51ba59e8e8a5b912b8bce5
z112c3433727d62e1244dd4a48cd6fc5b31e96fb1a744946ffa32d13004f2e89ebcef40bf7bbcd9
zafdfbdd0650a6018d08a5c7f3232338123097e0c398ad46bd79b68c2e0a3d7244401d485123101
z8cea3e5e2a90d9ffd5241a8eb28b2e1613ab22020f61aca4c7826238f64175a7f1a3b354da81ea
zab34acb1ef3022ae4cfd90e4279cbeedcb785fc0b00bd38395d7b5fa90e8ac514930673176e391
zb3d4c411cb802b173768eb7191a53d56a667c485b29c5e7a9936bf5f35b49203eeda723ce9382f
zfcd3a1bd97e565ea54284ab4a14f1c996b781965f6d42b6e9de7537b6daa05cfcbf05e2d82d85a
z790ecb8db0c0be5f5491b14765b4b08533cafb50e7eaf2ee7e74b1d9b8fbba69de05d0e7a64cb9
z7d3692f6a278fa1c9b08becdd5874111faf6dc20824031b9a4cd0c3ec359c054bdc9d6f7972bee
z8611b97e549be058858b9c965b36ee3ab9a22333812b741136d9b68d354f0bf22ff74b3f9a83fa
z6e47b265919dc6d4cf257c1b44aa0b9e719280cae015511202612688b9211391d1565fc94c0476
z94f156e18909e29527070327ddc1ce99089a343dd83a3a738d5abf951489e59a187b1a4cefb1c1
zcc2d784c7144b1d08495061c13ce1746245ebcd1a31f5cfb53ae810437c273ec9fcf7679c4f6f1
za5bb18d6cd4aa170a877f7391e8f3eea025706fe52852b0fa6f82f76477580648d6eadb0ea7bc6
z69d01ebc9a80bb0cc4abde5601ad4d391b4c8a8d852296dd74eccb8146e5da5a470c01844a0a58
zbabe478e5017fc08c13a0cedd1f9d189e7499dc15fc4408071ee68144704753d309fa90468af01
zc57af574e7326e54ed8cc7f8c8f08383443001850904d8d69cf13848023bea7e90d525bf51a55d
z36b5bb563e55c3a9d31faaac8f97f9ccb54a9f2318c92fea7feef0cd0d0c848d6ae7cacaca40e7
zf56c60b1e7f41fe6c5bee4a12d30a1fa5877e90cc8f6ccd1a066cc852c0663e7f28958ca94215f
zde332aa00343887ca0590db57a51e11344b2522896705ef0590d49349be9728e5d41368b62ae15
z80ec5c2b79a6ac60d78e7536b74cace3e9328bc2d8f018f251b412e1cd3177b5cbe4a73c3e1cc7
z30ad921630bb6b157154fd9c19751b4b42063fd03f96a2fbedd28696c16be504c862aae5a37898
z7a290d0edd56dce42fb2c06c97642c55b8182e611f986eb6d9f0d1a2d14e1772b017b0df184a8b
z512e8de0123c51d774bf3cdf470a3dce656e4dee9662d29795f2f6ef5fc6dc87ce09fc73f1517c
zc066a075fdb4013b247c902ee665280ecac8b94bfafdfd0dedfaaa391351ff5d2f80823084f6c2
z65787a51e5e461bf8674163e560a8e748280f28e4c8797fccb005d52eca0b667c48a9e18f086c3
z5c6e2a73370e708b97a3b136eb5a4b6a8fe12817c9f32333dd2b9dc6f3fcfdff7fe8a9eea3f7f0
zf884cf5c0a6bc9b4609e6d3f0a6cd55c594d4c0dd9535ad4589827f430354d5ac795cd7d466975
zd5c7ae0990b7b61e25283b4ce06cdbfc47f7dd4e12076d459724a998a0c55af8f46f40c479cb63
z6c9bb4489eebc49440603bac9f1eaf278a5b79e2e7d15fd64f851a413f4f6a7b130a6f59d7c29c
z36de7a175aefc9fc34f0b119c146360ac19d583300cf672624525e9dd9451b93a1ddd55df4f38a
z963f0c498f44cfaa382e450f2ef849b2d009ed8fe554923a9af2e7a68945fb4c321f83bfd14581
z8784fc503f7a795b57f856574fd0c4c29bc3deb1088bd5c2c3351b7bcb29e2d62c97b7ff5af623
z3409d49d5489bf7245741ef81734582d2c06f15d587f10bde947e49cd8ed6edc63883c401ebc1d
z47641f6e4b681a2a4973595003d6089d9b3da3fc78aa430e93bc0ba52b561bc421ebc4ee56c28e
z49725367b7d045807bbe902f2c34a24d1f61938d826fa92b3692a63856798896e05c875023f6ac
z848cc1688cdf660812d5b5d14987ca807a56c650f50be24a4135d1f37ad6efdf1347c1c0af466f
z8881b53ac0b72e771f2e85c8bdb7df246f1c72f78d3b1c31f77cdb37b94b2b8249bebe84fc6442
z080087db36fb861bff0efbe7f808c521052f768ce56abdb4c30a4e875f5dd353635cb6f3c49f7e
z8419a649a6637f336e6b4d06b8c51f2f029d336b75db5c55286572f0fcfab2b933be9b0f908202
z9fa198063e754b206ff665620669a097537966761c436a4ce99c35b9894ac3405bb94f776c360c
z1c9a6d9c4de46ac3a79b3c2515bd8f65c415cf9b93b25bae1249f6def48357aba970b417e4c3f7
z67e0d32a2aaa85b30d0b675dd048246f7f7af5f7378be35e0a2c4c3aa8fc0b6cfddcaf5a2a596d
z8e0a55f0346014e813c40121f132bb69c8723a565bf1894980ec166cb1a6834c200375250c94f8
z2d8fa01e5d9e62803a7d935662bcd3f063789ed3380bb09120c7723db5ef5f13f8584d0e65abf6
z47e6eeaca7f43194f918c21905eea91b381ecf85d4632b385e69a60f4132228c88e6d9c78c9eb0
ze3d724524f11ed7783d9f6e4020a34a9c8fc7cb438e182f6d27e315694260acb99b5cc670b4f96
z98a7f7373c763394f924842c7a16ea15e0792a5331a0027fdd76a963fe6da9c7686a074dc81bd8
z1b362b58f358e32687840fdd0b99e9f0fe2ddae9750c9937aabb030be64fec489b423543c51175
z1af99c278b952395f4b2df1b21ff2d59d0058642b28dbaa31d52e1347fe31b5c222da5843f305e
z70bccd3c78171019ad87df114dd453f741543a2bdd6b04f23c3d2e90b551ee74ccb22c37dc7572
z39f85e463d0c4d30064fbf80a2198953cca44a08f4fec55b64deed72601280d0b50b8a3dbf27de
zbb58bf17dc9f3691385e147bb2415aaa4f3539f121ebac8538fd46d864ccff881da13efc60ad42
z4728fc340dc794323286787bc2d2a629ee8713e21b1474529f02f223c5c4612ec6b375aeda657b
z2d6693127c032c6005f1f506ca5ba8f8188dadadf58ec2e1706e20cb40d1c498608c91bc0735be
z4043c9adf7e29dadf6c3037dd8a1db7b5d74cb0dbac6e5a8047d6eeb2efdde848db1629388d4ff
z7d751ef7bd3f40ba76b79d8fa301f9474ec87589dcb03cfb10c46c0d01afd3c293f860d627f28f
ze7cc9b057da17c3109a131bef84939ae4450bb4194e4a47115985d8a80c36a5047f2b1c67ec8e7
zfda8521baee94e4957061e6efe0b3f4bcc2dc24e78f98770ea97fe780a3a45c8d3e37b20137f96
zd0ea7ba53a62aafd6e4b57560416980fedb3daad6c7a381ccf821b39d870a6a7e522c3fe033bf3
ze617896e03aec64d2ad5875b0d93d42612ce492175b5e0a277d8dbf96327de55da3c25ec6b3aa4
z28bea90744aa6f911a21096cf54fb99da1e2c99659b03994deaa7ea81b5c2eacc5b47327872be5
z62d9088a53975abd04757a712157675c7acb3d6cd49f2e762722c630f2a5f15aed32ae969e546b
za75ba592e698f851015a56924aaf42ba25d95eee1d8b848eae1eaf8064e2ae9c000933c5effe41
z9891cfedd84ee15f05bc5925c8fa0330e6cb6a4eb8ebd9a7a60624d875bf76fa050561cb821dc7
z0c4b072435054fa38fe9fe52de4f641216e599a4ac5a61d27cca8841a6cadf03c63a8212064431
z6cadc0267a3688edbc0010299870f201514786d7eea7d1c23193d9b82821e4288889cf51d5fd19
zab017211cc6c011797233fb76986c53917500136d2a09d7f54560cf859c9cfc8630114cb94461f
z9c455211f43fbcead36668bee3ae9878d5eb7ced1365259c9cdb4f2b6c422264f502880ba3ef3c
zb513484dea79a9cfb907acb38c33a8543453a6bf052ed30258fecd320b4531a8956dbba5d361c3
z3868ebd29077a2b43e4c7c615d4bc6143fd64d61ceef3b4afb7c56f480f666c359d7b8d0ba146e
z5b2d4023559209a870a66dad718c267ba121b4a75d1e037e01b16713754a62a6e60b607e68f62c
zae2388cb9bde3996d07fb6b08df1e6741dd66da7fb5351184035c46f9f285df5603120a0eeea3c
zab3b6c79e14efb1b14d5ade548cc427da1c6a887e3465bbf723ce41ee1d2d2672e1c8f29ea90f6
z8502c3d4b6cdd87fe82599ec39c1320272de02d573a1c139cc3ef56fcf2403ceaa7607c5a2b341
z01f33d30366c810e2e3746a5101837e617ebec1abfa1932bd08c9bbf5086f5212bece071232ac7
zf7baf4e381bf745325c4c067dcf4cf258b7948e734a0406f315ee973d49f0bee72431f55eaecf3
z485dd263574f6e8b747fb7a98c5bc5a801edfa7a0e9332aad4a9dfa1133d60f65fb73b54d72973
z3175f425261e0fbc6f03f009282eb68134491063ca000e701c1fda391af6ed8ead219746c04fc4
z9c80e29bdb1520a39fa1cb25b84579a341d50beb08493e57cc1ff1d5574d2852535301428eab48
z97da4502e609442c6f2eb4350fd5c7ec7580961f374b54faec337d68ceb7b68279f222e32b7a55
z70d074d7ab8a50dedb94e345e35b424dadba000617a9443d8a4eabdc3497def3431727736e3cdd
zcccaf00619b4530da60908ce57a975b1fca1f20d6e6d274739828ab196db712470b405ef7f5a89
zf91eabfc03841b7fcf1797074fa838d83f46cd3d01ec79402cbe1e5828beb4dc17063a78e1d0c8
z10d9c1decb5faa33e18dc83bbaf709c1bef23989e3a0df74a1194bb581cf558af77da95fe9e852
z5b4c0d0c463ae4db573387d77c0b8901cb697940e35b46561a25809b53c1eea5f9c13908eec290
z44f09d125f14ed41aab4e5d282b77161b11f648a0c5d93c5b1f3bce5eea38ab43c1ad51ce91099
z157a625f67293fadaea76e0549344be8768a588216a5faf118cd11dcfc8abf74288c402f23a86f
z958ef2fb6684095d4b70fe7c5372e12cdfb6add5509ce4d5e4f83b95f3cf36ab7057925c80af49
za42f4839623e70694a0460507749dfda0dd6f71a41bd5dc7f697f2d970dfe8698a9d77418fc586
z763ec6d05ed3f553c11a04b674c848d6f6ad5f0f0f6af23e9f9d937b164623e5b3ed564afd3600
zcbeb0e2e777976f5eb6a0967c16a76f6ed64e7f4e187c2dab1f4b1dd17f3819074b51e35cca6da
z89fd35cf230a6f05033a294c8cf16d0e02faf4a8ea28a436e2ca39d2a906d76ed7707dc0610b84
ze36867e71b8b6b7043978c5c8165082a4444ac467bf3ffe108face225d635b62b8a3c1191b1711
z6fc07b18754ec35a0ef55d01e4f6d0aec0ae119b5f25b573f06340e727dbe929fd7374347ca549
zcada4e50527aaf23657d82938ea38442500fdfcd2d46db4f74e106dd84ac9e86002df9bad6d1b2
z8e314a40f311b095832c1bc5f8d7f9f069e960a29064a8a316edd41cfbca586b89c836b87ce0fa
z33def22f6b2ad2cc0981592949c70a01b8b351e53332982de58da7ce1b6a7ba2585e229682384b
z1f36902213bb8e45292c5f0150ff327a5d5a10f3b915112dfa13b3dfb7fb5ba4d3c44de8b1e73f
z23f6f051c13fa63efc8d0960a2fe49fccb859ea4e21e8a8893359c9f86cc41188ae5e17e0a57ae
za8c60fd3c04eb279dfe2061d77d1225d9c71367dbe731b013009a100bfde8a80f4ead004e7bf79
z22217fef9f0088afa3efc285fe41595e87247e497b6b99ab4ce05a8819ee6074abaefdbcd2344b
zda2cdb99525ba4a93dbc3ae2bff851def1c00dad5e8a5097e1169f7dd7a10963a8a7b1a4dc3da5
ze525c712a77d4bc4383f21684c54df1d71526e2663c0d79d9365c00337e29d96f9a64be5b66864
z58406f3b298270445b34b28a81da06d25634e5c163552bb5d6fc1afe7a94218243daa1f41c2e4f
za89820a3823d6271cb5e0dd9d477f1ddd9f1928147e8219db640d8a9ead86e2e5890972080911d
z1128928e0669f445b9feb60be00b21818c8c97f63261090840a543b1f98b89412514b596621c8f
z90171dfd67d2a40adc6a0f96d71b038d8b46734bc0912fc5644439cc2fd35716846dba7c47029f
zad40fbb37c90ecad42ac0677e273779fd42cfea87af14ba025a73b736292bbc2065f50484125c0
zc7102a385f73b3e8067a0a8b1f35b860abd765468400ee18a848bbf3e5c215043cc9b8b3f2ecd8
z8a74d444677d3c86acaed6cf8dada12141ade1631398a21445655e39b96406ea7fac9c8de683c5
z483e1c68508734987e55bf826a40c04bc3f33666c7b40e0d7849516c61ad7563bfade0dbc30934
z559588165e6de7e2d8dfe521261028d50f7b572d99a7c0b7e9714d405ca852ef86a539d62dbfc5
z3fc88f408f186d4933b7ea1c738c9c500ca971c8b8ad1ac8f79dc8388f8ae39f085c6db8b5ea64
zad6a7286fbd787042368e2c76175afe9f4fa7c21bb715e15c3fbf2d29a149b0cdbad561ef1cd6f
zd012325dcf5f6b14f110874dc454f1a5d0ebf2e84b8778e1dedc6a6ab1e4da94aca8508119bb66
z45c37ae3ae40082280e63d97ee5b3869cab5a401c25001e1462ff06cd2b3fdf74653b1e328b0ff
zb6de9596b0f160295fb4e11d3f21d5cccda7573eaaae94a68fd1f1660593eba8902f10c1009940
z690b6a3b18f414461ea88df83a9f56cbb40e6e800919d18781a6b72699e57a1f5e2dd7ff584bf4
zb41d622693446d36ca3ff1efbfefcff8078935439a9e71675b48e25c74808590b895b07ba3a11e
z1a060180239397f6727bcb32258d1baf0597deaba836abcedc9a20127640c6254697884c7f1073
z26bc091617d9f26e67ec8cded810a5a484b94970eac20f19a07f7a58b726796570434e5524682c
zb7fa014089915e1d0d7cf2a1f7149e10ba62b9316cc722075e80493c54dc5fa62de573f984665a
zf3e505e4b42eeb78da69886f48321607642ef01d55546b279b89c5b0ac53261a32d8a9e477f418
z99c9e8cb8befff0a646b39fabe17e455f707dd91d2d3da4a1ce2f5ec6afc9475105b8cbedb2482
z2b5bf92a949c78717c1e7e55be74506f697b4de247a004cc602bc1a21d74172a3dd1c7dd9a8090
z6be89e6b6eccce66da2a631ff927efe47f2b40240b85d6ef2d0aaff7fcae80e46f456690131bc2
z07f77b08c24de3db4e012cddfa4e03f221126f76841b380c294a63e7982ede6feb5b08a631ff93
zc6e9f447236aaacf7a54e214c3ac9ca7264d68c2ded46e73668d2a525ebf5b51722ef300f22440
zea172dd48bdb8a5dcbb4c861d6ecc4fce0da90069ee1450f47ac050b187560f6b4102f8b3081d9
zf50502d2aa3a0559dfe8f62f3f9827161bbf5faec291e792832b7b5b0dd4cc60b6fadb8895d44a
zff8d6035a44263abe10d212fedbc88046fb3b7ef83bcb91ab53ea3c2409627f2bf08143235cc5f
za46d69ce563564fe7c5372a2b329656279cfdfb83ecd9b6ad1ab9b9a3d529fc0c7d15f6c60dc83
za98eac5928489ef81d17c5a04d10df1a013106f336f13ff7084da960b2c5b98c0883e270a73c8c
zdaf39d477f587749a39245493284ffc5da541344dab7a6731dc3cbd5fd1ef018596a20aee0aaeb
z7eaf5a5f8f76ca2482618be9a7f1564d2947ebd08ee79455e196289d976d89f3504448e1df5074
z6c3f7dada09e17f05c59285111ab16fdafac7934360de27736b936e6b6db552546fa67e6d4accd
z613416fc46d92064aeb32648e9f9affbae68f9f98c8960d41062f7aff14d397f47d531acb0f1e1
z838769e4ab8797510dbb012bdb6832c5b17412d9876e2fcc106bcc30d155849fc9a2f8f2e7ac54
z02f4141087f21ff2db892cfc3bcee914b7eaea5b4834cc7d0a0ebb58881977c991ae9ad01a1ded
z2428c3e79aaab9e8a75055e5213976647dc355ee752f75fb372362ed6ccb33d2a4ed0d3899925f
z99b02131f3a9cb805f18cf976f156b15af76c0ff98f31569b05ce6e71d2286937b5a21aecc4a60
z7f9de7c138519d1e99d6c0f09c0be13d0e61e96d0e47e7e1725f94d28500d6b9515c150c51508b
z9ed5e790a8132d6654fd5dd2d3a6b8fc67408a2738273caa6874fa4477e045beb61e1d75122daa
z2344022f28ce205002bd1b3df084a34c1dddd6d1debf59a5514a60449efc32864d517bee0c4f33
z29c778e42e7eff205d1f1219d1dd869ff742baf86050f32307d9583cf00d6821ce581f6489e929
z95b797eae69284a853555ee0f6594ce477c1d2940934865e5d3bcf77710450fb4f4469f0f513e3
zaddc22b288243e3ab480baed9dca91ed236448b36f33246acc90f9e08a4236a808d7995ac1731b
z1b2b8e9642b26de3366a342544a689350e7cf46b040f5065f125d096393ac0ef557b6634c98378
z701ce7169d0c9b90cb048c5afc8117f82d3315db7044f898bc4f2e69da6fa1adc5345e97cb34bb
z5d33f41ec735626e207d0b98526389d9b381801d9b7b8e3661954c6de02d35c1fda06ec3a13e62
za21f3f5da3c853edbded7b8b71fc72b7c24e120c78c939228cd2f18de327c9c5f9c94f4cd2524d
z77389bf8b68d0a7889815cf94b8349d867cb344e0062bf48fa87b76b4dce4160fc6d4eaa2b15fd
z63de3b16262ff03300ad2324d3fe91f8c7067a4d1db348598835a6d0c653873d3c0689d0c0765c
zb0c1afd8fe9c7984ef8c5a0c198f6c49a029381d1f1f64877f71a3df7d895b256cb622012fcc34
z76f13db87b47f1e9c79c394ecbc5d1f5bf07a4805b2602b35d02d52339fb3756a37230f111e1d8
z12b3fca9d3029edaa365b06f4bafb69fbcb67ef5a456ae050c3dda767074b09d65faac48d8a121
zdb1a03b40c011c5403835b5771530cd47a154c72c13b144d1634bff057112871cf2c0b1a6093ff
zd51615c2d9b57803ed6aa470f2618b1ebf9290f0fbab32b474e0699e538bd45e65b338f8a8d162
z5a0825c3f70daa3e32069f40528d1c005a9b41cb98308cd757178c70355e2ee7c3d3ec0fff6e5f
z6e8f2122971eea8ddf05ae743ef085cc332cb52043dba29b4ae83a87b64996b23fb515c6fcdbe1
z83f1eaf94c180f6199184f5a2f4e29cfaeef69a09be8aaff8b1830c6385a0702e2483082281ebb
ze4e72752a3deb5a506ae1c26d66cc009078c3d277b9673187a2030a4e9419366d3f123157aa8b6
z9fb8ce810c1b4971a43453a9d74da9487a7b309dcd289e0e96e7182ea33c1b6f2824d1bbe4361a
z189d52009a9deffd53d8cc407051b406faf513a4ddaf78d6b1d3a1da61da813b76838b72ce7bea
za777fa960e9e393521ec86b24e52c96d01a5ad3d23b70723d4002ef446b0f674535e087c8f894e
zec77b102c6d598a77fbb2e05301aa507e605004f89e8a5626e4ebc2e83e50137d6a8e942e9163f
za6312c573deda0d472859a210a6d8cf47d88ec6b94c9defb8fb84374807f79a7e48d36d3dc7b0b
z853783b5ce1af2ff8b260f37bf415061f7a4153a2fd80e8ef106c69c7a741eb67da46af3226ebc
z45b0af4ebf1c7ce3eaa2dbe56c09a278d94b4da660f9bf5473f32578395eb94d3471cd473137e5
z94f9bec096d88b71e3913bfab0021933205bb08dea5a7f41eeab29d17ae85924e3ad348230fa31
zc498f7c747529ce71016ce0af48ecd701db639489dc2d21e18c930e340aa683a33581b1071db7a
z33a202102bd5c38e6b06aff32facba2df89350d00feead7ff27f582edbb6192a5fd6a7ca770843
z43e05f923c3eb989ead97e9c0877334a65bcc18bcc31f06fa82213d96c3e4adceb00388a35edb6
zca3e0b46b13f3f39f740d463c83188a2a5047e6af1c84e577bc3e2cf9e42fa17a59765e705977e
z338e584d853eb9ea26d6ec50d0f5566a183a8c37d74115e5b3570c6b5025d5297307d7837c0b10
z444ae9ba7dd5c49c203606289ded448210b9a079c5b121754b00f5c6b430f7d1bd4e732fdf7e14
z0e74567355ea76354703b1b120e315ffdf3643aeb350431162875aec60cac863054eedd9ba8dd3
zc92638d713400cbb8277d039cbab1403a73b2a810eb3f7e82256dc6acb2de8cbcff496cc58106e
z21370cb834ee313b375871052339d76ed4639ce1e12e995f4e35c5786746cf8871428e070c1470
z0b6a92f7be102202651702bdfb055a6ae50bc8688998dfe3e24fa492db8f6d86f1716c82eb322b
z507bc9e48207396e9406ac98522c3b5d2cd0e7b519a2b8e7aa32a59eddde4871eaae00271798ce
z1194c24cc073104a279a8e4d36484e0263b13b48939f7e70d087b4d8c3e6155880b502edbe74d2
zdea900aaea196ef11f844d2aaa6c8b02ecf5b0a068cc95f450ec49d27318294160d43169025739
z8ae98bce81c90ac74dea44f712814d42a5edc50d346ab54aa331ecc606112a28cc1acbdb59dafc
zb5514f882209cc0b25040c163f53da5146bd394d77b1ee1436009b3c0b3694183ea809187c68cc
ze4205acb9124445b57707176d123348de3b9157295492e9feef26470ab667a78a167360c43cf5f
z9e956b2308b2ba0d5f917784dde7cd2dfdc10e3533b4cee9790ef42f800592e84873ef4afd49f6
zae4d8869f6dd899238318edbf7cece7d209146273dfd75753f819117ce8afbcd4f29c92e5baf10
z52ba7e166b0c32755b1cbc3f1a25a3f3edcc8a5e90422757ddd1fbe35ca4367dbb6c97b793b287
z33429504b1a283fb82d7744cb133429c0432962f6fc18bc6c5277fadcf5bf01ebaca7042b6c70a
z45c644bd4b4d63fb6c2891f220bfab7b635d1578a37bf2bc0884a17602f3558b5f7ac4bc0a5994
z96de6135dd90f4ce96438103665e0c5f4b62802a64579f0c3f072885a1388005b30e1ba5c163ef
z508d49cec7558f8eac706102eee6d72505ce76b40e513089db8347bd58da1462718c4a56101401
z71dd4025a25c4e2d54e7b8422d4bc13eddb2cd94e7a943e3b21bb3ccb5b1af1476e321ad2e9cf4
ze6870eb85253ca3ee3db2f5a41daf99a901b1d94efb0d5fa71872bfe67e3488339137ad1a703b7
zcb5f8969c80d262ff982ad7ac7651cacf30a9efdc801c4b3ad0c390e8824cfe0c841730e3902bd
zf485a6b8e2ae2afafe8865582b84343c69514c2cce02cd40822cdb173a2bb0b7a38c54f22b8857
z7c4facc8220a93f1b6e0b3718af6284b36e35b990df2dd23c762af73520552bc05fba6055f4cfc
z7909076640f3acc1148a6d9e664996d2e09b1fd1f7dbbc82d0863e42d5246f549b6494b3e2d57e
z243b9a0b25ff001b39734aa42aa7bdde655a28cda7875cd85e4869b2887713015dc9ffbe88dd6c
zc81c075074435b213caa4037b0a9d161aa7ab4ce92761c871a2199fcdda0646eb064ad97ea1f5e
z71c667b6ec3fe6e02da0f17101502b6dc84a31c72ec66befb5cef54a2c49f21b866c8e1ea0c175
zc267cee2744aca10f746b5102d36a70a0bc97ddb15475095b22408af77d8172a2d9d5d02b48e3f
z4f0962f2140cd5722231629b1fc736a335cf59851e62359a23251d79f36ae7a22a06d41fa9d22a
z2acb9597615f3ad331c32d91a9dc53054c3d0b1b5aa45db6ad527f822924a1b0eb135e1846f2b2
z2a0ba81bbd155c15d0f4ce953d0961205b0210fe4f34ef4741a1819c2d8a70e71f5568647f282d
zcc823bda458179204d6840b643185f4db1c42215010707d75d0ee2b91a974d6a0815e7787dc5ff
zd4a7a2259a13fc87dea30be73324781045c44ea6ace41a5b4fe8848c79ebedabd6964d91853f1a
zfaa2caf6684e4bd1147101bf6a9f82c39d5ccf695f998c91290750f63a0bbc3ff02079f2ff075c
zd002045a2851259ed4148e6642958c32c2932a3e3c3a507307d5e46fff2b5aa57ad25575a78bb5
z2b47d0b3f63230aec1de8d586d697009bf0cb4400d3028037a194d54e066b781ce0efde46f866e
z87d6509220d1699f690c936711ff2638b71fdcf1db3a4e13a5211de5d832e29e9d320e5da49c2b
zf348f2828eadcc548cd82862c25e843dd80045114dd8e8a90a9e83d242bce04254c08e9debc502
z5a898d4441f57448af58d3f53fb9cc6dc59e91c5ec2a26d62d9515c8e4af3121bd783e0019eb0f
z248ba4ed1905e800081251567344261eaea90186f681ed855b543a011036701d9982ec752b5d15
zcd3878bb636e2894d7f689797e98be586a5aee4905456f18ce33826a4b7c0ff81ecc3e4c50cfb8
ze5cc1c2f84aeba4ea39b5493826bb93d66a855dbd5f9290be4e4ebfca8a326b52ac4f75a1cf4bc
zd3fbbd8c23ad51bbc8921877f0fd71bf1ddfabc2832d90344af6ddd12e8143e65d4acc2e6a7a2d
z9f4c380c06bd840384c02a84cd307e0486a7eca9c657001554a31d4175fb215cff3703085d9f0c
zbd32d3160aef12f98dde42fd87e979e64360815ce7d650559e2294dc758e5a11fcc69041c7354f
zbbf042b02881fe09f28fd797fec0e0213d11a8676150f4cf7e79e14fb994f846cd382aa078166c
z07ea3607094f94876616d3e543b9bb090aa05952cff12c9aee61aaf7d9cff02a10b12a5e92ac44
zed1e249e7b18c535eb282ca1658a05a94ed6b0a182a81bd9c41441635968b210104042268f28de
z19b9d70a95ee93f4726e084e14f87926b45ba71ca7a8f7b0d0a17afbf7bc907fc64e677fd14645
z646cfa0ae24427bc3605a45fb6a9d7509dc7df7f8f297f14dcc7952b6510619d59fdb3da3d326b
zf5d69a47402686684cf7469d88a1966f0f8546893683bd828328014bf4a362e20403b6542d45e6
z5b0243538ebe47d629df55133df2ed4d8c7c0956033c9c5b969f294e63b3e6490543a39e8ebdbd
zb1b5b6aedf72ea385f72dbeca2735e0d2aff8b48490dc57b907297c315390c509a68b020b5d843
zad7c3f05dd917bfdc9c3691431e169ba7a8cff5c220cd856184f99657fbce42f4a70d4d0873a39
zfec55cda65be1676fd95dd1b69a71f04ee7f0ef3170918c5850a5ff1cbd1ef62130391613a44f9
z9cb9b045ab91d12857deabcaf99e052c51cde42a7440cba7f154f30a22131e27c04f41b8aaad7d
zfa6d5be44f6f2b52457cb9e225a131be3f1792ca977378dff01131a0672eb61720c5222bd55418
zf3f8cb7a3d23feefec74c1196348a02f8283e6dfd25d205200ab3965ec80ef75b6c3b7ea5d6d2f
z5e4ea02bddbf1160ed43a1a71e3757422372b42c2c1da8acd85a2083e86c6e6fd0e071717829e7
ze2a50cc28d301ef8a2c3ee2b8b194a8da4406ad8b4c2eaeb43e113703a0137010393f7f6f16ddd
ze1a631a592a1528469df5f49ebfbc2b6e0d96b40864447b697117c0762cb16094b72be12336747
zb56f701da2238d77030e7c5663c187bbfd5f1e850613d3fea2e33dccaff48226dcba47975e3540
z9831afb81160538cd336dc0f6601688d449e3d4572f4ea61086d70d291988edd480e46f687ffda
zfef03b1fcca89beefe710740065df8475a59913f6cea0952205e2c32edcd10a7dcdaff503ae230
z02fa4324e951752a8c2c55a7974e6b9f406be4f3dd7e62e1d3bd69648b9782fad8f6fe0a4f68c3
z23dbcbf78d9e8dbc71f46a52ddc7a816221a452568a943a85f2affe4a7c5f3dacfadf445130c42
z0ad6c8af63968290d43f00bb7d527108f62ecb974cce5f11179f13cdfdeaca13548dae1a81e1a0
z7250b779b22222849b749fe81e412f25d0197c58aae707dc409d935f5bdae20330fef716bff6e9
z2f4da26b0ddd8024ec39f46e04760eec9343748247f81f7cd5c88671a5eacdfad5b6f99c02aec0
z34fac956093bc3269edea3ceaa5ad74a6b13e9ee08c72db69a37a07e09574acf6618f0fa40f001
z907d4cb7e8fe10ae2cdd2f4fe237594e5e2e1b1d241235abfe1e5c65afcc9af7083f7a83def9e0
z6b80746bb73de23a3400058b734b1f759e37c2b59bb67ab2ac321d6b1543355b7e49b7b156a5aa
z18298d2ee2abe5b0bcaec7f5ba78d32d9c440b88f28539511f2ae6d4572127a0081bd18738e276
zd5b6977aafe476d5523318c601fa7e88e8337da7e9c31b4f3826853f476d805311814ec118474b
za6db848d2cf4fa3be26e6fee9f72671a8c96f9c775fdda93af8c9b899748586b925d248c56a93d
zc3504ccfc48611157aca0570395b1a92dc956fb97938578ed105e4678a1044b18eca986e52e2db
z500881ea99c711517112eee55869ec9847db647d18525e728cb5e5a7b6a53fbd3725e522043724
z1a567d292253747d13ff9689596f8c8f8632ba00211cf421bde21bbbbf96cda025a29182f99f57
z13b6623a39814a83ee016c0085107fcaa2e6d59ec01af745e5205557fded039ce63542828a75b5
zd387dff06618432a5dd0857ad6a975779d42cc953c2fba3adfa0b00c37efb8f04c847bed241078
zfa385a79855ccca14d698de248a9213336eef3951b7ef76bfef90681d1867e1a1a42ffa58dca35
z853627f33c065db3629304af96315a039c5744020b743de9951bc109656cdfd6a24ba2dbf6b571
z14880f832409c5a4d4ad3590ea1ce982fd3434b09b8fad93cbb5b54c04ac74a7ebff0c7ee75794
zff851441ccdb97fb3049666649fc9aa383bfc2e36adc978b233212b3ed6fd5f9391cb8f77e3393
z13871ed2187380ad460cfe9c63fd7782d939de13a3abaeae0947aa593c50accf8d03bf6105e308
z24fcd3e65f3d454626cf45ada8ed521d701a0c639b793daba8cd52583b1dd1cce9015d692add1c
zaff55cd7daeaa92395f8736329812de4936debdb3671b34422f5c339675314cb304055f2f51188
zc677a0206d8c7003ed98fbc9263e4028ec3483c9bb79b93bde176d1605100a369a23ff1b540f09
zf39326703007866452faa929e22ec5648fb4a3f8aa0a4ecd662d525546749a52d09220bf3a4cf5
z966b80e5040f7702d72327a69af51c7ab6401d7a57ea7d23ef83764a9b031e076ffe4d1b68867a
z62e1b065b3887d0fbf17d7eea4e24f64b010c94b1fe8c150ee040b199a7fe19fe41047232ad14e
z75f76672168570a364bf1271618b35b2e5355733fc77907a0b8ff2624914206dc0a82acec5bd69
zbf4ae5ec17534504744273540f2e8d6eaf41e8ed64fb2937c620c0ee40fd9e3d5cfbf68183b7ee
zba71e6b54a333e21c915f6195e6950ddd672377ea241828de21898ff1c7b15dd61636ec248d72b
z6d0811cf4af271da7970b311118b3c0374375e403295b03590f7fa364951758aa8e61a6541c398
za8bf3148cbee175733bdcc5e446e94f6d5eb77adb78905f18182733b0e69c15c607f4d812d20cf
z818fbba602fd14d37a3de48f4b6b8c02703828e4c15867463199c8cfbd8b7eeecb2cfe52975849
z83a6b67bcb6c6ebbcab16a96a79efcf5d363a4e49c3d162b22aae34eba896cadf64d776d384d57
zc18f3291ddad0eb230a24c27876a762bc6b288eabe846f43e970631afd2ef97464bfaf1b5ea189
zc78db8f1d1cf1470fdc7a3406baefc387bdbdb681c81ecc0ce4fa8379d87a74f8abbe6d57a62c2
zb66a042ae13ac225744d92d1486eeb4816453a54f5c41267cdaa8d47136e001b60fc100c07a54f
ze90d789d7638d79445117f5dbfe38c7b9c9a0c97e95e579d862af7c2f5ebe4ecffe383c7f7db7a
ze12c0f774ad4da8558892b477906cfdb009bb6a6924b461476064dc384f224969dca4a33e3f394
ze757f24ed4c9c1c3ea6fe9e8048c69a1751313bf10da712ca99263bdbc2524b262fe6d092e73f5
za0b9dbf884dcbdb5685e5df6589d796546aec85634bc65d5451ed68e8e0ac43fc16b44766f99ba
zea57c423dbe78bdfab239ebdfe64e495c795a013d59c8d3aff218168ae0a9bcb2c0b2dbd22150e
z30c71b18ec02a0aa0c96dab93fc8ca1672331a653d5784913c42399cbcedb8a41cb1d0de4be0a6
zf28e96cca9aed58a9a54f0bfb3f791c760992413074e64dd29e6737bf9481aaa9201d41e2424f0
z5901776935148ed8778fc4f4e7405b5da1229de30c3b9b5cf9d4942c065a59fe3739f9d870fbf0
za7a99af80f3493a9b506a0941972cf643586ffc4aa62c66eedaeaf722ec3fa72cab816f2a80b33
ze49406abd9655cf145a4301a0fcc4d25be053a17f1920008166fee1bd7fdb08f6dd568b4618e93
z2121155e6e24de5632d4bbe03f31b832a45bc8dded303b4a766d0349f2e966b6812faf939574dd
zfa15630f108e358778b581dcace61844a89b5c48557da844149d1ead2eead5bf7827aff1ae7269
za41429b9f5d5e6b45c81614a8b619037a202a6fbf796ce327f11306426d0b0f4bd4e709980ad1b
zd6df28397f21f2d02a31b5fccede8d5de8d18f471c2783337921bc1db46a204a54422cf9e4c433
z2818b127c2cb546fd41c368edc0449489cca4b09c17d959c5f012745ec227a238c482b1a086fec
zcaded3a216060c099858216c79b2739532eda9d21dc8b6da36c19fb6d89c39aed5574713405ead
z3a411649ea144692cba5f15159f00e2dcd9f9bf47830c96f32da57ca70bef33aa41ed8b57db4f0
zccb6fa59cbf1871dbc9319a258cefecb84fec61b58d11534036c024c35144e06fcb9ab42d310c2
z2b46c1d15b2ad19e45607fb5faaeac533fcb143378493b4626b80475bfa4de7676c5f1eaa04b92
z2dbf8be7d413136a272e48dfa988f3a02626c7a47f42a1f98cb35fda9cb147346009ce34a86ba0
z971297ad86f414bc8e0917253df2a2b0d4de4100cd27a803fea0ebe73a53f4a5682d9fff812ee2
zd54145bd25a0b504d7896776cdfd29e06fdd176b239f67038f53ef912fa5cf003c20367bd8a165
z6cdeba0987f729c4bff767cb4da0db8dad9771a68953e2ba01d0209f4fc7eb2f5f640b1355468f
z72b03dd5460badca89d20ac0c75299cb3a1bbe3e0ee475b23d0985dfa535d0b650d2fabcb00935
zbcfdfe7cc1c07fec7c13b967ecff30017e7fba7f9dcdc3b8f1ee5c8f7e5d29eb1a00a644747b95
zeb266cc62b87ef70634caaec9497af90b27a0f3b6aedb4ba827a5e9c95f0d6f576a1b98ba1a420
z62806926877584d549cad61bd318d6d8bb5ff8469578cf5fee8dfe3aebc30bf79061220f9adce1
z00ca17b72fc204d53c8fd92bcd69f13ae0fcb371ed1d09e9131075e060072cea5ebe49fe0289bc
z0d53a98ca43f03acdb15bbcf74b83cd331ffcb950b505cab0fc166a1c6315d346fe7b758b7d196
z70d28e5a9135aaadb64eba972b4f32b95c678172fba4e04fdfd8531f4a7b968f73bd31a16a2679
z6c1842c295ae4bc0597488ce429d88a9acda0b5efcf234613d3e4f96e0fdff675bbd25d3719b4b
z2272de1f8067ddf5db3acdb88975ea952c54bce02e9b055253e4dfa8ca0489a0fe36c9c16ff806
zf82e82ba887f2a8c27db6619c6dd0de7bd18a76a843c020abfda286b946385136146711326c3c2
zd3ebdff41659da220cba17fd3636fd97b37c5d5b5fc5ec400bece0a23c05c034f477670da1ba14
z964a73c2fd866cc127f48bd5febbb95c77b66cab60a9f5a3c30a9ebd9cf1dbe0847dc3c4a09de8
zbde61dc1becb33c96ee098d0db3eec2652c37e658409c7a3f16b60207809e8a8afde035be50f97
z913f5969bc2b201314b74cdb9dcbd3d2137941f6789683c7d2d6542e5473123a3b65c0ca2010d4
z8e055934ec789d399f6c71f590240ce9127051800c027b27b033306c5a8275c50fab32fe573c98
z4cffb64e849056a2f7a1220f14ef1b64ca2ea2b4827ef7db2c69eac54be7c5a4e0d79a27012f86
z75244d18f84b14af8702ee1ce2f108be4656e3a8834016438287968d09cee8346dad853264484c
zb10c897f3a6aa2eaefc0595dc385d6509a37ee8d7ae572baaeb6486bdf35fb39576fea2c0aaf35
z191a82ff30470b6fd0bcc8a50611dd1c38faa51f3b50ae4a9032adfdbb0d1d0d0cad7f2d5cf956
zff13f3e09d6bbba52235382e14344df14017f2d6afab685f6fc7ea3c3ff298b94f627170fd00c5
z16ed039bac1a81e8c199005b64b66ecf9872738960a73d50ee0f6788b081f84a458cb1dfbd1007
z7c05472e5edf9d1be61119034f5f38ee3ea5d2c1967b7beb9cdeb9a8eb8ae5cec4183d8dc70294
z8718ac0d769dc50f5238595a38b223a3d3db42b395b2e7fc3e9aeb70d65437c4ba878fde163653
z5a058427aa1f2822123b22ddf8ea8ef85bed405e589b1bb0eb915ade8c4577533c0e9df6fa4248
z013f4606f59640632e9d915d26c8b34052fd7ea105d4dbfe8483c605dd13fe7c58d8a6e1ee69c2
z0f405517793a000e94c576acec3bae83ab1ec6b8e5f4704b4dc2efd5032efecc8df723af72c88c
zc9f0941a16af1161a23f726cf103f76b853ad6e6aad20cbd380e029cb903d8373d7f7c1b98df60
z468deebbed42dacc6591d233abe5532b71b360962d8b2df7615b3aefdffd0cd1b16f1d69fb920d
zab6b92c0ee3cbd0174e56e5bfb9c09170d1dc912a0891e2c72380f2a233a811cc1f7ca6d907c4c
zc265d0e75f763bc071cdc55ec5c5daa3a5fe9995317e0c14ee3e8e70600e4260249a3629babd72
zc39bc08d083c7d2d9e8d4ac5f0e8719e316ae907790737b94799f2a59da79d3c834e4c2882df13
z7623dc4b76dd91ff4db475d4fcdc7eb3f8ba88e75be630e2bef6e4772fd1d06751479dcdfe84c4
zf40043771193b571f0b34d4030ab7f7bd4eb22093e95404d43c3c1a656c6c18499bce26162b975
zff524a7fabebcc3815d1f4afb9378cf53d0f59a4c9117841c31a7a5e425c1f0ffc7c42a5a504ae
za3e80df090161077a9485a51c702a0ebc597fc257c0dfdfbd5aa0aa0ba6342f230afc7d82c174d
z3c864cdd5b0a0427f44d6ef7e866ccd5b928ad3daf3265058e111d807359b80d20049b753150ea
z182d0906f6487f73223e530a55f821ff1d35d7ed5deca9aaa8031286ece489e163a1b8f224df4a
zace2b896b0f29d6d9bb7badd2a433d6ec99974328e9be46be0797788d49567cbe1cafbcc4d677c
z9ad16c39d3240385b6b88c7e5d7355497f8e7f8626ad549017d18dc6a0501050e557fcad13ab0d
z7106f05132e0ea9c72fc311b62cb25fe3ecf5e84cc8e8c3ba6ce759f514b208f754bef118a6399
z5286de19a653e75b82390a72e84a2ffa00af8e3f48c6deee7b74ca26b74bae275dd0a9648ff6e0
z4b6b62b267a7b8fb9650f62276459f5cd50be6437414d49b7ef48b2a5cdcd2c0810ea4e9722aa9
zb75fe44b70
`end_protected_0in
`else
`ifdef MODEL_TECH
`include "qvl_pci_express_logic.mti.svp"
`endif // MODEL_TECH
`endif // encrypted_0in
