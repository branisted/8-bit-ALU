`ifdef encrypted_0in
`protected_0in
ze74c34e226135848fe16db9ffd31815111b6d7fb642c521a3f628cf6da949865580b22efd062a7
ze90adae0e65e66a2c36a587d0a790699161455169ed55a01f2084f11770a774ec4c588039b380f
z6de9c5084882a40b79a175f5c2114b2b6d78b070cb806e1c0aa9258297f4687ab308bc470f0040
zb0b1de382961eeeaf2e279e1462520fc31c119af8f2b214846f56c2b3cd2eadbe4099496abff18
z15cec83ec4a77b868344aa20ba7360908f5c0de2a79abf8b3534b883bb12180f68b5d4beb444cf
z3fba8f13afb0abfe8fcc4294810f75afe452434d2d0f1166236c82f76edf1e12979f04bc35693e
z32ae028996dd85737a8f5adc1ebb94f39c940246e887647b64782cd7ab429b0544c173176cede7
z01dfb26b1f73408344a52b7e1f117f12bb9c8077b34876c2e6fdc085981637012dc9754765e1a9
zc512ce062e0b8fb16a214591f5c81e1353b900a611fe1f4886b57940b41b7f2ce99a7b84b04b90
z916f717e73bd10589c81e207ed77ec660a8cbed5b487fa50acde1b055c8870bd8676023f21ddcf
z9c98cc47cfa2d654ff1365d1f45035a045a66c5dfa82790502623b57a3af03bf0f0c0d35b51558
zb8b5f2d29acf03737a9ca2a053b7a8f06800d50b465c41b30eb585f62f3d0c2c5a43bc3904db24
zc5b00403e1023c01d567dc70f03774cb5f32042b7b5829588e293ddc99e016d15d352f50afa9dd
z2a950a0c92ad79f88f58f016849c522abd2e4c2249c47de2a58539f3d0b1f635178ddabf53ac1d
zd9d3b001c8e3cb0ecb91a31acf39fe413defaa195158c2922c483e2354abc16f720e6514faf1af
z5d5cad78f9d895145f6a9eb5c34f94f82c94a9b782d64d2270fb3e63dacdb3dd45795fb8857927
zbf043382a43b43fcd12cfa0b4c5242c993ad52d115489a6f47da000d682e105e84df5731c2ffed
z9dcc0e3b32e2288275db50962637a4764fd4f41302a7ea34012866dfb0962a233a50178ed5f852
z18b6ad225a3bf5fa94b0e649b2749aa72ea88ca32cac790d4e8abc2c5cbeb11ffd027bd8f104dc
z5a99cd91fa65443a6b6b7e144698128e578727a3c9793b57f1f838c5652c48eb1f43db2cb3bc3a
z6bb4957c0796004520e33dd16b2fc9a0a6c6c1d44e68a96d0cabcaa971f3ccff1311c92922b203
z2d04aaccc7ff78ba1100505d9f8b7ec611c067ebda30fbc1dea868354f58bb8aff297c0bc48dbc
zee25f47774418615d7b133373dbc697973cd1d5bc8a5e2b297f31b257ae52e931139364d348d41
zba0fb71fa9bf093dfd949809d3ec948651e592df2644538e83115b5e030b2a5ab35fcf675847f6
z92de9b7b8a5378be92df899f1f4fc5b23a6f919cc5d63cc791bd0375ae1749a39983cf217a0cf5
z562cfe476b211bd421a17dac25fb6ead72fb5e6c285e3b9c6637ab8a14534d434a64310573be45
z49c5db28452f17a18e14310af762825e5fa7c786ebfd2923c4611fca9b33bf934060f3302981c7
z0243b8515fa71e016edfb0cefee086a3e6c443bcefc3f96fce7be52d3e9d6d2371f69d37196f94
z176052e92a529b61e4b1a24e1381dc08a8bb767fd5f14e405437cc936901ad0a16c981d1d23161
z30f63f9f0c2873c5c8ccd29a3a93f7ca8de2fdd08a7c753a839d2adaec08d4beeb52e77a601144
zfda6e471680c1a12937695d0cf3a4ca8f965d45ae3f91965b6bb6bec41da2fd669846d80a618fa
za0ff364d043e88bd404f9cc650b31477ee564d63757e28ee8b3f5b5f72e8616ac8fe7b7e39703e
z686005ec36ccc7005399faff497291d3464f06997fcf90f288a4544ed8d265fa4bfd177324f57a
z4b0188f2137919741ee9552b139a84a1c44710c98249e8e619a4bd4cf10f29b7487c01c99ed7d2
z403b28510ceea6ad710aae4c5f91fa8878948419e7c6f9474e4969d031fb70f334f6aaa215c518
z7f35ee5b5b98ec505fc736db36b5fab845569b459063472b6168e905b39c1b3b6192f3b3e7b3ff
z7911a46d15fea85e153a85d25fe03c65a57ba9df0e41f79707206433d059175a0ce15fee012406
z158753e406a1d2407f7591439320b27d352bb77956f7e132b081d4d29bfc2e50e862afa8647c03
z9a080b759f754c5b84f42c02a6f0053f0c92c3b44c2be9bdab8b3db1d5e7c2a7c62aa9b9c101fc
z6c148b8fb2736e4523239cf49f91d75b6813311724d62448fce991f293a306ffb69b9d63ad6374
z07cd15327f36a129f0288388a81c8c88fc44e98644979a1d19258a006c6a8e24f73620fca0734d
z68c32041ca7a65e9f26f705ef59c2d308def098177d3bf8f9fbe65a30c0cf9c7daefbdfabccbcc
zbe748098fe4f24df2beeb9efec1cf60d6f912f83eb94fb9f19112ec1ddecf0c92ae496599854fb
z8a439bfd4afabf58a7ba34893d1cb655faca40855c869e289e5c94bf04361adfb18ec8a831499f
z6b55fbff02b54e751fba56c8f6c919379890b1d43ac2c6b384541f5d10f09133de29edd700ea46
z03e9e037fdfc1ced80c4d78b0a38b0ac27d0f84c1c32fdf0ef926494279074f60ae28c111ab73d
z5e3edaa997584fac624a4c365e0d4ec726b1966e43d0c1c035bad9d88cb7a84935d528faca2b7a
z83020d1a1c23b8852d7835289c82f484610cdab24c04720924d5d844dc345ae5113c0589b6d06f
z578670557e7e17bb68885d326581351024f1cc0c1635aee95c832aba6beb2566def4085b5ef08b
z493859a26975a73a808d37ff993d70dfff2fd932c8cbdf6dcfc2ad85e6eda5991030f74e1dd6c0
zc7341a5b9af593e5a2049ab48915c6c8936cdd833f9babbf6f6343919fc040fd6374c66a25fb92
zd2a06382207935db4eb92fcd55f4471bdb407cf9dde36d38adc38f332eeddd98b8d28289d1201a
zd1c86bcb4bb4049faefee40c1cd4431d89df039062faedb28d7c269f0072cb7e6b0dc54ada9de4
zcfa0c64936d5e4025a69a0c81753f90312009e61bf4ffa944d26d1c40fdb9fe277d4f758746504
z8ad40f7495f380a0645a8abf7f6a9ef71663221923b2fdcf49a6eec553810721e4159725d5d640
zc5410453c6beaef1518134eb7ec84a94647298d73f46af4a5b3c6f39dc836a1416ffa970124202
zcedb72201f49340cb9db7203a9acc895ff440d05f0d08c792754da18ffea9671050b235e42ea24
zf8cdba5c2c00440c66caab6fca350419bad2394f1202592b1f3bba0a2a1b05b4b6757a4dad8e5b
z48a0dde0b531ce76e32c68edf59eb28b380c0e0bf169ceaa8f0c9431e67afb6ed51fb48604c4d8
z8ccd1e8e2e05421c07098e8570cc8a0c16571aad5d4fde7d014a20d1a659075e41300f6f4e6d51
zfbdc6d697a66e02eb6976887c1a5341783abdcf835e0973680204f541d919118d76657f4160ec9
z9196139698285833abaa040aa85315f3262f6ffe55c36a170d8d57edbe770f61f2b87463440a7b
zb217d19df3f9c9fa3384f547e1a493a1102776b3135a27b1ce433bbde99a1eaa855e241c54e4bb
z37cf386aa7f43f767a3dd587304bcdf609cb3269931eb5920202b7ddf24ff60984736d26d849f6
z73df0522750d0f70e7cc31d54c99cd5207becdb732d128c46a3e9eca1b3f116d51e748b0e03bde
z6eb7b8ab787804cac38d73ea6f684b71a9d12a226d1cf20ee2f40f753931610f81ee9dc681eb16
z4d759bbb5c93596a5d6afdcc439a176be6cbcac0e12de334eb5197374c98906e681db788e6f626
z2a039b1dc79337e0e51455ddcf3abeff2c71e173d9672432a14fbd7624e16ea194ba9fc60e3cb2
zc32d1439e4b9d0c60970d2a069c48d542eef463eac79e83245205bb01b907796728cd158bb6bd3
z8502b86260886f4b7192fa625b4e18ea584a519adafe0c09dc8ff1015367e40c4869d3985ca4f7
z27cb1b70dd3793b12ba1c54fb6afbd0da7f028547dacd58034eed1c111c8912640d45e59a40ec5
z16d09d946878ef1d79961269e6a401994a1dadd30cd52f618e1c5af5ec257c8eda1d82173cb57b
z175ed014785aba649341ae5d3000e96c1798776818c559c74ba79fab8c1e5b55e38df5a087291c
z1e7ec712454dbb50bd6f158ff9595af62e560d237476f921d9747f3585e02659625af46e382e2f
zc5d7650743c8606f2d3ed9da45eb87eb344497d872db65e9bd029c8dd5bd103716ac1e68bcebf0
z8c395199eb7eb9e605629f6542b4be02bd3cae9485a81854ec9797d682461387810aa0eacfce9d
z960c05e0f23167b3393904e21a5b408a71f1fd328bc00ea1baee1649b098482a7757cbbe918e99
z032fe36e43f19a2070559e58f8e533cc088990c25200c1664078f57f4bd04320fe906780cd4d2b
zc6920cb158cfb9068cd3b67316178d29356f37af84465e8a1bab33409c08a063bacc06e5721059
z49208f24bebf3a91160997da50dddb4c56ffcba3704279a17d39829b95d134e9d0462110bdf5b8
zb353c75ada0555920ade8a2f40b437ca7450777ce9cc66e52a7d01cdd285da76c1c57728c700a6
zc4859ec9edbf883a450a0a5955cd13a9c62f73cd1075f381092882cfe1e5e911cb61860381a06f
z048ce271dd5a51038fe2081a84d4964a6a5755a0e47bb817a7d72a8ec1824721175c9e52fad6fb
z8a4bc6dd8f8ad8e04c526ef484a617bf84241466757bb6931b5302a82dae743c36af41fbf9975c
ze76a23dc5a56d49e401bf2b6d27d91b1777c290ef98dc50cbfe83a812d7e88f8777241a611647a
zcbb4e52b465b7c59d4f569222037df00c079187a7caa1776e88f9b9b19437cb89c5c90d0d8f4cd
zc361f75fb8e9ebab09b690f12953d283e99bd536ad648c8f7852f61c9a8f6aebf4d20f7c48adce
zdd69b094cd54ff3f229ba906e256f8fda0267e2d32417738b174431480596184d11bd084bd32a0
z52ecc2f782ea3ca0b3e187287470d835bedf4e2115a2323109efa00f61ce8305b9f1623a3f5cf2
z1333d806270d76e54dc90e0b59ec958a81a87423034a410e09b7e7882c96be2db878bf2ac17f23
z315e2fcfbbeca2fb17f445c1c5210680862f1fc0a04f44e0a290fb54df1b1d7dd9b4b9362c9056
z98a90973423c8677c7e3ae75051101b01450e71cd1c261310d7aeb0e73ee2bd3e9c1e2bdea6655
z5eb25572527c08f2fdda9ef995a65ba3aef25f93c159625f459f1fb47c040bc0d3f2b5990862d5
z4656b386f84ade38eb0144f0b7e477bb3177f8f1fbc2c6066d5110150adb77ecd0c8a712f64c3a
zfc707879866bf341e640718a21b8e692fe92b346f46c436b2c6060b0e504d699ec3c8ae0a14ffe
z25069755c185e0eb8a278b9515a91ff32ef44f04b6b504dd9520c0db351665650859a653bcad50
z252607aad29ff2e18d307402d733662d62180c614583c1433782f390639959b7228929c3dc81db
z81b401faefed21c977a589f9283aa9ee644b995bc3c9c6f699352d72f63b73ca0737cc422a7c0f
z571123754924cef2d8a6d33fa4f067ddd95abedab41f52ba22dfb895498ac167b93692fc2d48c8
za0dff9f03aab95a68f40d6d6c2d5c07b4a4f2db504c6623b90a94a67f74e6487d0fec8811c1e65
zf207cabeeb8a6a9fe1ecb81404377f46172eb87d99ece593b66d3cfdaf336dce56fec6f232fb31
zd3adf59a2467956c9b457322287bc3d315f6e271b5a3529a585d25b2d394630d4dde3c4bcdd23b
zafe0ebe7dce3711b1af5e8de8e47f54e69ed54dc56b6c7bd5ccd72b2791b704f2c7b0c6a943ed8
z78894718bb817f4925cc8c89c20ba03cbe509d8822d353a16064e021de095ee7adf2bb524fc445
z39e3e25386c5dbd012cf235a04f63855bb0b2364124f6dd2b54e844025bdfbfbcd3daee10af745
z395c549294841d4d687797a08cad435a0ad36255d4410c85f2c7cd334187adcfd24147fd6531a3
z8aecf1ed9ca0ad62f05075c50666f05b62cd41dc796025d045ff90b78a2c90f211e3d489e690ca
z16edeb8133c70f7138b1ecf7a8d1744e26f0436cecc3c138c46733925f72d295b251097f90586b
z0b143cfebdcf8dbd42184fd35f97fc85a7583117f0a5944f9d8e57fd3d61775d52759e91f3c7d0
zeb93f1bf77a0dd5a7309f9b79e534a646d63bebc7e93633f73626acace610e662c225d83ce7480
z078644235b8974f52b5844abac31856ed1a79de249c1491013a9b87ccb63dbd5641c58f9d34141
z343f2b581bdee1199da952864c8bb29584e9fb1beb64be6f642acaa318a43c72e4a0a5df33a009
zf5d868382a10044ec518fb89af35c7d0d97bba5fb1da483ab2efd50b0575b29ca0c32befdd4d27
z90e1338927202d90535a0d1cf611a0114ead4718c80dcb509def5d1d30811903593e1df2a72462
z2f3935c2b1c6db19b2d52df6616f94e81df9ac54a80c79f2dfef8b7593a888aca05a9e6395de2e
zef34f25d8271c822bf4e25a7a21f491ac5aff516e1b73c92288d94cc3be5dd096f3be0eb69a633
z7322ca5fbfdfda0a92aac266cb5803b1e60655cc104ea7cbaa6c2ee5fa5db9e937fefceaeb9c5f
zc5abcb2b51e0851298113143b6c709880b6cfb30d6b32060bf378599a3f8c69bb825020088f735
z490526f133cc0d04a26280bd2e850a6a709d8664cf098032d606691962bdaaa7541e50fd6bc2c8
za6f863eeb03e001e96e1d24ceca652c4aedeef95abab38c12fbf3609916f81346f25f0fb308f76
z2def105a145948b6f28615ee4047aaef7248a14a5630673baeabc9f956d6a428a57735ba032174
zb9c388cbf73c4f853136f06e3b7ce8fff2ec2d7119f66b90eeabea6bb3a07311b00ade01def7a2
ze2ed6f4602ddbb2ac78d3c354444ef82e7d36c3e72eeea9eb41096e3aacfee1128cc4814af507a
z22cec6a1f52ba5a7e524654914ccece01ae09a9d33622cc8e3d25a2bac33485a2a78e8b9008950
z2878c7ba00e897dca0467bc34f853194113f77b382f2aee75418e3d3c3c3556623b8acbda4deb0
z95a889aa8fe976ff967a809b8998001cc0b8be27a22a567c677a60932255fd9af6a4894dc5dc1d
zc2a483cb42a98efbd99db05aaed49e54024dd111037404049688cb6a19e834e38150e35d79c098
z75880cd76d6bd1fb7038cd1d309e196e29adad196ef89fd474d9abe599dcbeb8aa5f31ffc25926
zdb6658c22aebc5c88ff8c82cdd40d2a013f4da06e93b92338ac1c67014c917d6de1c1d0e485cf9
z5720da39e443988a6ec7bea9cfc29c4b3807b666cfd28f2c3afb14cdad953aa1edf1f85450b85e
z3cf588c60392683378743344d06d339f05db37168a91ff47b307542389a64336ba0364517e6396
zb4e54d99c700ef8995f764d941f698941f1dedc982e7878cf7ec056ab41be28d8b5b371f122480
z86372401533fd5673b0bdd595ba2e70294c501aff14c6dc215ecefbb28f40fbe80c653aaab01e5
z41c037e7f5b9bca29b35a2b490934da062d5cdcc6344d360bccf991e6c2e1100c09e92b8c38f67
zf55753a90d4a55310b54ce496c1211aae987f92d17c344bc4473eff8fafcd431701d909366b4a7
z242b90ea5ea9f9049f343942ab38b52b6b4998bcdc4273b59c96214f2154274b232b96b8d88839
zf68dd133ca574de9fd7f9df4f454ac86db453287521d10e9daab2ee97c0439a9889a22ac9b1199
z6579fff035a981496a7b45b571d1b90d248bbae471c1e15eaf2405080548eabf5e6cdbbefc6eed
zfdf2708d733091557839f033bef6f9ba70f04a772b3d2ad7672c8620e8288bfbfe068122440c67
z201d37806865f7d4d65937cc66c4d4f14b5f4b7d1b94e799fd2c9c2dd5d51568546a13e1a25c75
z9062fe95801071e1153d60498e9c815901c7cf2ed30b5a3b7a731d3729070deec0bb193e92f614
z6bb99c000e234300ec6a8fcf52d6e7567dc3c4df4f03db5cf9ab4a072bd6d084299bcc4a37899e
z1ddd546c8fac3ed8d8ac3de4f1530340d711f44cb5113f787d27603605b8de391384f257986bab
za7614c94f8b8af101b85f36ac48b1aac297ad0c4c42fbf06b647d80e5c3f06706bc57900ae6d95
z06c3612945f52b841ef28c5c4dfc97ad8855d3c256923d0797ec647b7ef9ccb742b49e1985f6e7
zf5273b6261d3e6696c0990cba1234368f52f516937c2965059fbb0d7ca17f93c9c5b316133c502
z0d80630b9a222d79effeb196a7e60d9a31f3fc5665703b79bede104184e944bfd324299c1a8f67
z55ba784d7db2d6fe6c083a7559ab680b615819512db7b6580ca3f74a43aab39137d91d04e86941
zd112415dcab16516d2d64a17c5b7d42902709d60ca781bf8a3093712fc452dd886660ac9203b26
zce1943bf6edaecba7202d82c212573c4a5c0324082f9eaafa5c8c961d07645a9bd1a8da4f07b39
z7729e7e500f5601b74bcf6703dff8a4d572262937f87b9af209e016076dc87d44a8f5d564ebdbb
z0eab8b2758c4eace0110ea4ac63b1c3b03cc54e662a42097023d6a0d76763c53bc6c0a7ecf623b
zafb765511022210c79b8f2fbb40dc5c8ba95f2397a60af5fc10c2997cf08fb277a3959b0b1ef3a
z17d7670b7e84e5130be211296a8950f80355956706a17d61def7715c778bad69a842075f33d3de
zd6ef65b9eeab5ea9cf41e0e606925536a3f32a7ad55fec62ec3d387491dfe33340f47973b72ad9
z9aa98e79a7fbf82e28adf85f57e978edf8780674010b026a0990a40dc252cde8e37fac45a42e92
ze60339a21091ebb5521a5816c42d03f3b729dfa226f63857fee7711924f39ddd935ad61b9a7cc2
z2df8f88092fdcc99149bb2fdf6c5ab4533d8fdf4aca2b1eea3f1d4a1b0891d68c5adb7a3a1fe37
zdff16b1f4f880a836206c5be3554e3feaacf446b74b1b9a456a327fa219599efc2a8888e411e40
zbcb7a3b75d522866d4a792c6d2b73fece89540496bbcacd58f468d41fa8706727d7afa9c11c38b
z00f84a92d7672760d127a7cf52e2beaa359496c452acf35280cae987681b4a9aedd32e4731416d
z15fb23cf4e6162ef7f87ec323d92ae943ddab3194c5df4feabc99f2c302713fcdedb8d5be490bb
zebad6884a80c4a452268ff5263489eab1af7de6f548e85950dc5b3f7a133045cecfcccdbf413db
z52324d32c58546e1290759f9c563d0a3586c40334c114503ad8932a8c812aec8942bfb71cebca4
zda67210c8d8aba44b4548308dbddd19c215e28886c181dae85ae48c175a898725ab65af9ad8f5b
z4291c94bdbfb21972277b9897d501fcdc38c4cc19837f820fc2945209b7498a42fa135405f7838
z9339e8b69ff37ab2aee53b5b0a2035e330da52791af2e46866185cc2df937e130842b8fdddadf7
z7a6e4e9b7df6ad6dae949b5ba3422a12e85eacb5071c878b65777a8d02be2f064d99433360636b
z2abde7cba6b1a70bab25d2d8d3c3a87cc30ad920188acf9ddacacb6b0cd8fb4d117901f19c7429
zdb06b7f43dfe1afa5e9feb13641e7d0080de615c4327ad76274dd8c73a2dc2ad2087a625ccc2b4
za1123d4137bf3601345f86c76684bc229e611f415ef7574728957cbb3828c42daf11faf52e29d6
z82c8469b4deb4661b823a2a5a09dfc3665f17ce575c530f67b81a1aca83ad15b06f3b66e849224
z604222983eaa51afedbbbd63f96d1bf47f6074998b0774d71fd78d01f522ef0154449d3915c336
z4b3627adbe584befd6509ac0f7ec941f40bbf9b3bd774c453b73d5070edd151897589f34c4e4af
z0491adfec912c6717f34954cbac418e847b1642d4ca418b1532ed9df66a25ebe85459dfa0f090d
zb9e99f2a5dfc4290ed05d48859b9a4348a4ea1751bad6b9877d5ece6b98792c3f8632062176531
za523fdf0978a0e24c127f604b8ec7deb05276fcb7c978e9713e38bca0dd8faf4f7939e4cbe8442
zcaf6520d5d2ef71447a56b28382eca12630e09208609e81dcffe09642ef60f1b6caa8866dd60bd
z1b8b05f25dd96a04b89f59b72321d27aac9c55a4b43b92328b21ff7041e63fd9f55bdac6ee2964
zba924b3245c52c34109052f54609382c47679477c8625437f6b9d5fe6eb02a7a57ad8cc30e326e
z13d6e7378c9fbc2157f24d54e661bd1a272c6385a262bf9538e64e8f554f0695faedf45de547c7
z25acc2cafd43544a721cba07ae544aec58eff00650fd74317c876385e394d9b2dcf9ec87f8173a
z42085018e233669a91bc442c95840cb3e54d1970eead4d88a234a1a0d666f92e389397ca24abf4
zf260d0784470b0c62740d01f2cdc71a1d40a8a6f746b3a7b82ddb29bf5c270f8cf4fda1619b48f
z5c3cbf5941df2a62c33b01d772decb2496f51e5265e047e0ca810e43f8ca08844fbe7ccff1039d
z76f926ff23cf1fe24c0458df65b4d4dc90795b0211f4542749a95ffa5c6ca31bb907d331bed131
z0f8072d1cd1bdaea09f5f37e155e765c3593320bd77fbb8db8d9262ed3102b640bca21beb6e9b9
z2dfe271b9104a58a11f7027c463446423a877749c42840884951dd66a11bd4d038897b818ccc55
zb74ad4b0fd9e9300f0f507e4dfc7c30e29b3986bf0d22c5a008dee471c5396dadc555664dc74de
zfa3928882413f92ccbf23463810360bcd7f0380d897258c361e9fe52b5e013bab2f59f47ea078f
ze75b352e736c45e0b6ef3447d62c99eefe797e9627ea3baac7ff77286ddc026460a977bbef168b
z1724e6b7fac75634150fef14901a14c872803a540550bd436198c878ee2d243ac158633a355b62
z19de54e004d2040cf9dd6fa3d9164e67942716c122e6e23379133dc86724126b9f455296c596a4
z8908524b845ffb27208ecc465a1c8ca8ed09bfd3e5baef02657412075b723fcde7ed23ff7e5ddd
z374c0c1c0eb527be704b440a0f5fc6bc956a06b237755df6bb703a772036ac7cf5c0d7f2d365db
zc90ea11e8fe4eb9335fc9a2b4851eb4074d9a2904af40b9871b77c6aec0005aaf708012cc3958c
z832cd62db14d3dc5d3d90cf8cb1dba1d0fad470e5972b21d7163d50a55a400207a4220eb6488e2
ze9dffba34d46968c39c3dd442e23af4272cadf3c9fe06a99eea4e254cc8005341de86257039d89
zab5d84ddd8c36003a7d6f581beaa8d16640b5cda837cc98bcb2f659589c18655c77426c00fd61d
z6393c2ba186793b11c9141e68b8b4111d8ab26bf483879722963f1096afdc6ae6fbf35da163e92
za7fe3acc602a75ba69883f6253e83c6337f698d6300353f9d80ce9906da8cf5aa462d1f90fc037
z9bddc014339e94b8a6b2cacc4ad6026eb4c4bc73c9676ec812b04402606cf4ec39b457091fd55d
z2f72f4cde8aadd53c83c21e112c2047af10b16b8d89983e38f1e97c44490a48574f91e0d4a2c9f
z7d6e60327def54574b10593ff3f082dc2f23dfbc6b9ad8e1dcd29f668734a5051e3487837024e5
ze1af82e60ceeb9fea7b21a46604c86e5a2467940cc3d7c456dabf68f9423efd423b8d8dcc5d95f
z03c2df8c4034eb8a0a1b44ba0b390478a138266298661097e85931f7aa3fc726fa1a135f30df21
z4a3dbc3fe5241ee8b2b8f98bbb7a847b1cb1b885e6a452c52bdafff982179038d775a0de3db72d
z25cb879112bc7c7d2dc0dca6747170c9fadbb695627177005f785cf801a9cb2e3a8b48a0b4f772
z3aa943b6d1ad54a176b77757d98106284dd2c2abbe8b0bf600bedbcd0b18ad3c596b4a03363934
z22b9b5dc38a11eac02ce0417c233d70e22b076964f7b4504ffe0e5782ee1ffe5336f0a423e5957
z94d4d2285e7b58af7ffb247cd071c736d93678e88de3f31b5bc8794fc76ea681856d2d3aeeb104
z951c686d46ce11526ffb199581057efd017e8cc2765698bf7e738bc2a13c9aec903a7d4f45344b
z141023bc3210b5b6c11fdbc6bbdf4e3ce335bccd770f12365676184f6a514c77ae74a33643e212
zd88d4b720a5dbaa672a15315646c98742ffcf5b22c1f7dbd7825b96647ee6d3a8564a0e9d0fd56
zd57eac7ff2c7b0d7c2189d4ce66361cb9927900a617673ca05b18f99a9f569424057ae005456c7
z5db4e662c56ed9e7ecca2508c70df08a3005f8e4fc39487ab94fc7e8bfc181b287006c3f69b510
z24569d4598b6b46dc33de0eb80d4996d3ae6d8d4ddcda3f146d99daa461c6b24bb0ef83feab93c
zc151fd9411c15abb309aba9fd7cb5410e69a6c707388345ae2ac4fe4f02bb3bceb43ae112ecc84
z7fe8df43802e3845abcc0d06bd422105ebf84dfbdf797053907ce112b0fa4d1c9ab92b99d10d3b
z3dc5bda824fc5bd9a103a6d30dd0207ea1e4c0fe204464af4a6fd78ec09413ddd5dca81927287e
z0f08f661668330eabe67d4f6c98383540bfc190923c58e898e9472a676eb29ea632ceafe7d6e82
z82facb809c0a51d96b91fab9019e24ce08ddd7cbb9ad400794338b49998a2435c60547f53b925f
z544ded0914294c13b31292c0a363ceddad58e11cfdbc832f40d2d4466fee81d94f8a3bf49a650b
za9e4b196405ae3ebcf99ecf43fb80162f320e0eb91b1587af5ca5b6d5a235d059da110640b6aa1
z6923671f48bf30e9c8adad4e579da24e3e1061a530aff4d885e22ab2143f0843404ddcbf147f86
z72ab6bead9a42fdb1cab507f1879bc8810c28fe402e624c1c2d1ad63c970342356627de7678653
zb61ffeb05d52869117bf4b0e67a61af5a58113616db098e78cef25ea162ccd0650dd9d4c6067a3
z3c7b4b6e1943f317ebecac0e4265b03bd1a370b258c0fe2d3a2d7efadea68d112743ce28345489
z347e37e44bab406349401ce67a8d45eb54e7a4c73a0846dbf376090bd6e3d6d33404009fe9a9c6
z92c6dee1af3fe18ed2e44903710d3aed0333baa325f6e6fe5cc343e4f548b0a6de9a380dc36e7f
z384735221c2c7feacbc7dab22aeb5bffbee6e0db6f6b18699fa3c62f5903315de4d3924fb46d49
z45d648e6ec32a2143e7f4d3189f1cb6d41b9d36e023fe85860095dcb9e316a6ccf9bb508798ce3
z34c788decc8e274ccc13295f91a731a851d85ecccf1569e97c3efb563c51e0be2735e801af04c9
za5b89e159aa595f4423a9782259b809d013d1aaa83f3212faadad9ea72ebe5ade6a3a7c6a62c62
zb1dad809a6d047c6ca7e480a76d1bacdc0bafa0f98eb280bfd6e8939b78e560c551b526abeca14
z4c27f94d6fc4028282438c771beb36a28662513d256018b890b4f1f171fd739af615e1fe63645c
z7c40306e28b025579ac68009c238e263d8d0d92510ee3d4d7003959906611dca8b6b2673055f6f
z1e6ae88b96a04af76cc063a51c92279599e08e28f468d3ccef7f70a5bd6297bd009c5b3953a3eb
z14fc6c44bab0d608b6a8935e4bc85ddcadd5a7b30efd283dcd0d8a8d941387352ab4877d96a888
z53673b080e980787a4f4621caa344274031bce51a25ba389665d4f67f39c3804dac6fdda9c43c6
zffbcbaf031f7c76137afe3d28b9ff6e7d84da4074ec3f22419580bb2557b874243a387153ae303
za3dbe82f5d37ecb07085ad6625b1393ac420bdbf2a33542d67599de6e25a23670e7bae8c639c87
z46d5e64e3cdb982908e6445e3e5191a36d51d8b5a99f681959c2d7cc65d5d2b43044e8a4c4fca4
zbfdb05ffe0dc8bdae14016e09bce543906adad99c7932f6be322006ba8e1d438c8907f125dae8f
zb0a91652fb05ebdfbae55ac273fa10f5902a52bb0edd1c9c1ed8c220e7bfaa896660376c06f10a
z7279577f6c383e19a905522b1704e91d526316877f47323c01258839288ea91e01f7bd9475d007
z52749da066dcd12a08981814e8119c325fd9c3187c315c8ec4d0b4b5c407a8b099e2a6fe77a0fb
z9f8122f0ec7207716c5ad273224321645368ed3b4066a39914101fae7e2bbfbed1bb1d888aa32c
z2480f716a72c0cad198155c8613d8d048908fda33c74f7eadae3b980e95842c5ef67f4402467d7
z8bc02ba1666a17f897b447d66c7492e0251b498c161228e6ebb4dc045cb0b68057fd4297f3d1e7
z5d25fbac12e6dca58806eb5a2ff3cd29f0553cdee56a9fd1851c332674509a9bc3c66c32b6c549
z95d01c3aef5ed6eb97e4c9c79da7cdabf20f711d7ac36621b31f0fc42f1d9715c2ed834f2f5d1d
z4d2ab58f7356dd6afffa5a089fcb69abbe13c5e8f1901ee530d4a3e8ec2b7120ef8f7d84b5af81
z79e931918d555ffa11f89597861202c89e29b7293fd6ec3bccc148cc4331b4a262dbce573ccb43
z7b0cbdb3029013142c638bde0f68fa1dbc452d4bc4081b0fb78975c86e6d390a8916b331ad26b9
z6c1a96d21b21ce13216317bc6a276e830c012c6235530ec4535f91d2dff9bbcf1d474b2d9a1543
z59ec3f0769ec650bbe182e66823d2a43d5d79bc2ef6390481c00009436406d2c4e4f55a13a1548
z2974d97448b2519e0f8fdf92728d107cc3ef24857ef456854c4ff1be86b9c50c45002d3ef1b9ec
z559e4b8c1e7ccc1258990805d53ba77bb9993cc6daf97ba7ecb47266b10a236ba5e28da61e8d6e
zf918d33776c3016902bceb03af9a4ea29ec466198b78baeaa8ab8574c59de9c6f205d6b118444f
z19e29901e4b5aa4846de1cdb0ea00bea4cf2ecdb8d50699793c550622f238514fa46a8a4fdcdcd
z941fa17caf00ddb5685795d4fd9a09964206c08bfcac6490ba7979f67e9ff473327c16519b849e
zf5de2cd71a3c46e6e52c03d7f255ac941f427f5516a4922834e05ef29f01ca2679703571598507
z3a856a6af4a8ca055dee7d72b1dc06d24eaada9e98eebf7c47a64ad801e4ced4ff6ebe23575642
z765f3cf82af6d29b9f2cfcf8f9cde56770db93129e2a5edbc18942e436562268617543bfb2bc7b
z759803cb6325efb145a1df9b8435b76df677c71dea64252e299d0e4cc7c27a5d0845cbe03ef7d7
z41632de969bf26f0581c9d58ccd12dc57c6217a2edb6500d21e3cc84d51fbea3491ed9cb5486fa
z4034155784bf3815d341bedf01d3079aa547c6d721edf47d5275943562e0938f1cdd27e70cd1e2
z9cd35ca543adc8a2b8dc7a74a94924e0d928e6b833f1849d916b5311e67d179bc6340af7926ba1
z7bb895a9c8cf7cc1a9ac9d1a0055ff86d0d572f5315666409ec433c056bbe8ecd3f7b42db9ff9a
z60741dfbf1bffcccabf0915a42ebcb5c3aa57fe3434ea9ee1fa7f254499468b7c66df444e97b9c
z40f8b1f0b31a5ad9b9ff39c82b0815f3dd5d518c0c62e1ffa5c7462ec49a558dccc54655a132de
z088c7e5c005f123b7b8770ff0301a186c152ad10faf17cc186a7f63977e753ca11bb2417de82c7
zf76c6e802ec0749647d21a684c2cc1496db2a5eb0db6cacedd7a002ffe864d36ce39ccde78601a
zff106b40c281f388852ca5bb80f2cb72c088d7a664b925d0cd9b93711e9c6d3b2d4839337b4ea9
zf37e97739c2cfcfc6a1fada676b2a80c96c24bb5cc550f6b6cb2a201c0d686351bec813d85a3bb
z3b4457b3e060d11c10dcf7b952c93407e90a3e0d6c970cc0fe77115165b57a32cd02362c05bd24
zbe207ba82c599ae119f8f8cfd8c4375372f469dd38d58e78448d5759f1ec48909cca1d3340949f
ze98de053b12d549a71fdff5643c6d4b5cf83baa79ad2b287ead6b7ea819a35425f2b877fce40d6
z774520997d634d41fafce701cf1211ae59eb01e604f00c564a3a4b49dceb802bc280af574e2b08
zbde7f598297d8e96654a6cf8ebf059620d1d222e49cae4f888c8eeb22cd5dc19488267696ef809
z95ef9943a88ac6648e81f2de500147f0539c76493fdee5c16dd50e4d4eacf25f522fa832cb48b3
z875792d242c51eb0397732431547042d623a6f5f008b747d403e9a94ab7e876101c5647d3451b5
z4455bf86ee8c683f1c9014c1dc44350eda77d16a2798dcf4f6ca12c8eaff5b299486feb5a8faa1
z85ef9f4a35e2259ae229bc7ae83d29a79da579d58ba16f3d3aa1c5e56d24d13ec7673d9572cfa8
z3230dac61437590d5dc0e594aa372e8e5e5d6b058f336ff443823cb351bd25228985b55fe631fc
z7044b3b5f3b058dbdc3a85ec0ae982ffcf82a1347d85c34696f8ff309e2e1bcf1ba86b03bee76c
z675e7a25c772a10ef2f22f9c61a433a3cbca4e065837843a47442beae3d3ad15c12e4ae133dcab
zc36a79e9490851577b1b94a6b2735b5c3b0ccccc8bf2bf397cfb200ceae16b179e8c08ad128340
z229d4cfe90005cc3087f44bc2632d0b06981ebf1b842928b9b1a7cc07b92b318ff170d51d330ef
z1bb45bd96307146339e7a5ae120ca3741b4a4b0e3e4f519b86b11b9d68a2608d768dbbdd019208
z4fb41546300d40f9e4f0ecf47aa619e648a1a9bbd3cc7e6c803fc6fb5c4daada62343f724f0e21
z74b3d30fac6b54ef3448d2f21a0966ce64ff84682c4e06f8c80a621c7cb259696f58980a4ce1ea
zc86d1a1f91cf6867d769ef6fca80c661467a43380bbf93b2c411a6460db0e635af9f9eff63660a
z66c9bec93368590ba04158fd536757d0b229ce35b27091db77458fe4958ce6dbbb81912b9a5f62
zaecf9d6616ad9212751786bfeff1b841b0692365cac5daea8fcfe93af69841912c498a5e2c42e7
z4cb041c117eea0b58f9976778c41201feca17c959c6ed28252ad2142e92d0da4bf7c391b5dfc8a
z050f0e6584f1437b9fc68f4ee474df3ae4494eab638c7908e633ffe83f11ccb643a6f077038a59
z581b15a923426d8d5fc73ead7185259691169a189416384a70c7dd467d5356b63f5503c75844a6
zc2a1c880b43a66b8022f7f16d8417b2f4129106f58b4aa56e03160b661a4b4a1c21b99412f65a4
z510b78bbe1d1018ae1588ab404c105348d7612af40d5916f8041f7c74c2864e8b497f765c3c1ae
zee30a307c61d1bc5754325c341b8866b4aa605a19dc8c174143796bc989ee4318db4bd8ef168c0
za42d95d30935054ae8ae176c342ee2b3886353f9d9eeea4a7cada01109bf8d7f76fb1979b5518c
z5e1f2207d8daf269636d0978ab0a5a6f7fd79f6bd5237afb8ac9d5f6e02d8f1f96d538c4ac0f15
z5703abfaa247ff7c6cd73c5fbd592f7d638dc2bec6dc7ff5a6bbd57fc2afd12f615a2d29a79f0d
z8cdd9b09f44bc9a346e1a6a64f10bb5ec69abcd5f50cdd07a2a9761a0446eceeb89a0b4d5590b5
z7f8b497a0e6494f426e0fe1503b097adac2573d3f0b6544311654051e553f65dd516f1da92bd93
z3d985fb00e53657fdcfdf1fbfdd6fe1fa788e72eb918085ad8bd9ee7476e399d267b263f8ab79f
z8107cad7bbc07cc1b54312b65412aa88e78102306353a96e7c6eaeab88b2e15b9519f85e443d6a
z2d47e0704ff17e825ff5266e3b8675967861fbfc473026d2157a343f52d2760905ede9eb9b5689
z7c8f30766f9faa381297f46c292a56730793cd42f6cb05d458757022623d4a8fd02d295a5625a8
zba5397921b6532f37bb9166a50860cc2afb2a842f1fe1dceec52fcf242fafc920f65207a4c0a93
z1dea0c23c67f72c32b277eef46158e96a934b655161ede1acb62b8045545ab7673ebdcb263556e
z7a18de48aec1c6ed093849ed7bc5a907e0f036cf958936eb8e16d3fbde042303d060f8c9a5e49d
z5819a95fd89885412027da901a792c4c7bb39900cd1c9c1b135df687054691cdab58036913da8b
zb068918218f43d5e044b13ecce9db1b5e07fbe67767dccba96fa006c57d55626803e580316c873
zbf03a63a18dca7155f0f0c9b01ddbf13b6021821b10287ae1ca2a476dac5cbca4d7e900fd3943f
z6959e0a1a87590a127c27de26da7b4e08eb66aab99f317438bb33dae80fc63de4adf0467544c68
zb8e41e695752c16b884bdc1df4e66f2c38654b4d659b64cced764316cc0115cbb7ff32cd58fc6a
z87ec6b47edf3f0751239fb1cdd8afc1155363895d3da7a4e8720428be188c71e68798e4a9f1620
z91a5d61e194fb00abfd08e6aa3be36033b00003e1175caeb8aac3d2b45c7e768859308985c7c27
z41e97a46260351699bd9896b120018c66906f145e1a60da58ca56f1bd9317008e0d7f1e67bdef7
zf7b7e8adfe02e1735ad0334095df956b9f2e64bd4ec6801bad101cea7f477bfdc3da05dfe1f2a1
z9edbd5de6adba1062e06dc80571b5ba86bf242b2a8edd94a57876e29ea3b44117f29a6099d7db8
z226f6932237d9dde77dcfa328664d44d54c1d0b22684304f4167bd633144ebc65945553b1031a6
z0c2e5d5eb5b110ed7536c33326a7f3d7bb961b41a1cc7eec6c1f4f311af472dded652213e93694
z65f6e54e928fa1ef548af63e619e137a1577ee240f44adc12e643619c51fa8cc0d32d281e604e4
zbbf4450fdde8e211fd5a00337daed6368b860c2dfd05593ad6299f470b1c0bf9ce5d6df824e449
z63235eb82a2aa2de8f35a5daf8987ca1e6b27eef4574cca5ace781c81094638749f5f41d3af2d2
z34476944164e0510c7d38e5c5f2b1c22cf678e92709c27c21796073e7125bac315400442899e81
zeed9a53ac1ef9358d88cfe8ee9c23033d4b472f9eb0f856fd2b832a4aae0923b1944dd1410ae8a
zea54b11dacbdfccc6ad6b8d48fd85721be4afb1c925800bfa0d613ab7cb05cf7f3f38507e33a66
zb93f5110a04efd492cdfc18e9c884bf0f26cc0463aecb90f429b5ef7e38b4abe9b97a5c1f91222
z677af5c74df51a9e9e9e9a57fab00d994b39b70af9a8de2eb5c3775168d720727d90563aa8d626
zbc3f7e7ee625a0ac88f59b331d62aa0f59c31829af572cd1723546e5a7c8d3aeeabe44609a6d8f
z99ec5feb0670b69cd69f9bfe97772391624a3de5daf0b5fbb39b19be11b1b7d4f15d31a47690f1
z6aed00f8753cfb08f8e2e3a0582d3d9adf9840d3f01cea88ac5a8c1ee374eca28874593e254065
z1d4c51de4b2830e00500dcaf018c111d2ed254f4b24842d47737df3d74a3c954f945dd35b80cb2
z32d0f60a148a91637157c0a021e49dbd0d02550cc9a4ba169c41d9c409e25089e888465633fd1e
z8a3af533eb973813c15b745ead310384574c2d953995fd81cf2eae0b3c0d75da96867316762e4e
zf7cbb5a389b8d40721ee65b7e7bd73553f2261547c661399a1ad03dd39df67b05376a90dc240f0
z1c2437bb306f6cb141fb1617e2b510b11433e23f2aaddde5af85e1bc72c963f497bdf9a4e17d2a
z9ac56966e1ebdad748e336ce7cc2ffce52b28be6eb7797ec97db32de1b0da3c4aa645e697b99ab
z935962fd2ec92b3fe6e47df1270e5556a7b6ba71b45b44e5bb2fb6c105a88cb88f10ba3e43a178
z9e2294c8638a32a50dee22ef47f9c6e110b2f335ec8f0f3f01452f71f8f2a52d0a7533e6e4e023
zf01906ec7c10d6213f75542916e6d47127071130e2e90b6fb3986184b7983af996242ff458f425
zc2991d4ce4716234a84df5bb3eb33ae2dd562dcf3527dcfaac304db18f7d84b550d187a0401f80
z9773fe9b98e6d88095a6ea2186746ccdc7bfcead82df8fafe1846c38a3b5b1188e3d170d086b8c
zc01e212d3c3fa0e566a47e9a10dded8b9067a212de9cb4cb15dcbcfa76852c1227c0e0e2f98c4c
ze754dc322ea429e2b983b079745ed0f51d3a2a6e621b8b747987bd7373e05ff278fe23da882b07
z02c477274f5c46ee0bffbc8e942d19f890e18f288871f91455c6773a52624cee5b30fa0af4a82e
z3e38a92cd92ced81f47472cf84d3493308ea9feefbdef592c9ccebb642642cf24be7473c4bd6c5
z83aa69b77e824a1eb7bc0bdfc9c2c6bf323dc4ed826e0f67208aadf0b40cd692ca92bf2296cef5
z8baec0a28bbe6e2072d5c70ea66a030f7673917e466b41ea1d5e503ad64a310a1f6a3815de850f
z326cb41ffd3b3d290ef3ef09f5d7e81a510f8dc1c93e8ffe7829d1a3eb8fee85d59aa61a295869
z067d60033d2c28adb15a6c0ad64751813a32e53c128d844dd05f101ce077e98d75841554e9805d
z8483feaa0d485a5d40c59b56fb6dc083afd35f2e3d07951968145f3c4cdd16ad0d4dfdea6badd6
z6ce6d6c82f9bd1f3f10f209cb0dd6d7b5838ad64ec00346ae575602a375049c2b3c3fb26a895a0
zcd82f56626a3c43c8d23e4954bb9884ae65f8296335aeb66eb7253eb4332dbf553ee26f90f20d4
z2df5cac488b32a05ded947493a917885a636b92672de26b07b5b89ff23dab13fcfe022891a6343
zceb7c4a4fc9888f1fa78ee6b3299d7506f0ccc73ad6e2ed7c5f3592d7092b1580c4a26d7f492ad
zbdf0afcd5e44cf7c2b0395eadaf3698140fc8ed706f1378d1e05aed9a0f8a6a2d9e5574b392966
z147e86f1bee0ec101cd878cc065b7a3997fb66c7b951f7f75468447c1d850d69b5c9a5b73bcdad
zd2b66fc3ad12ec752e3cddcef2626135a74720aa956de76adcbd8e29f4331275d83ddc1cbab757
zb88c3be2d6d7468642cae98e6f8ff596b5a31579cd60ef07ae5a16e56fcc7d954ac3d9a5a1847e
zfc9145300f608301266ef82d8ca482967e3e63c9b02f39ef6b57d7ce5da90097ab9b67ee0429be
z151aff5cdd8ef444de03b0060b47dfd6edf34d028821581a86adbc9a1068a54cf387da01de790c
z7465a9aeb8571e53dfa16036123f6efafe90abcdc0982329dec435c186c4e8ce9cd514c4ecc1c9
z0fe29e750f3242644cacfb2e7adcb9cf3c5fec4d3646bcaa867a61709ffdf95b6eca524863c1a9
z86176319ba798edf49ee561446c57d3384e7c906ec47b32331d4c5d23cb6dabb49fff5ead05765
z0b5f4e2987f27825333c4061819f8e5a57a5ec2fdcc6f28b32de67719425c69c055337d88433c7
z13fb2b6095de2aa7f214eecbbb6ec790ffba751ca675936f2b6c8c4ea7c7db4f66223ccefa5aa1
z45042845852b4b47061059534ab30c6e446ab9ced4c1e928c70ae73f3bfca933af6a23f6e99599
zcf1f77c73369c353478ed8993d2f029de425f1b33bdfc6fe0604e570a33f134b58c623c91efc83
z57bdf4d1ef70f024c600c8818ae00827f9bb9055c7e7d245289a5212bb29cde8f3106f89b5e825
z8bd47b991cc797fc1cbd8796ec50c153333c607283d9a842df11b19e3f8a64b11bc669dac12d1d
z73f33dd6af975fbc5158406589df9bebac9d7b97e63aa4b3060dcd689e3ad489acf18bbbda10fa
z863c69ac0ac35fde61bba8de497950f4f37f7e05ef4f074e49900117f86dc9f80cd9f05077be2c
z16e43445b42030eb383d352a83692fafe1e2908247c7321f7b01db707e0a160c0a8eee6e2c47db
z1bb7aea9c4b03c83f54ba3d13e16f2d08f094aa19d6837ade65547d6b3bae33d2fec671a4d2f02
z0891be8b81fd5741e348be778ce94eb28e0cbd3498bddc6dbb8670b1f7a64b380586ad482b2342
z9a65bd78e3fd8a9812555c9158072c51241283bd4de353847e4c9845a605ff5f97064c264194b2
zb627255e4967a569c2bacc4c52156bf66616cf3e4974894a7507431411a1cfcd1f15f96ecb390d
z0603e11b3419f293a442a2a6b7c1722a7e19473fc67451095f2bfb11d4122eb8276b8a38145780
zcd4fb6e8dfe79972cb540dd2149a3c3cd63cc3c45d506dd7f1aa12b9154e0534ca8b4b828fbe69
zd4e982e76d37546ec8e761607dbc3743f0c78a35bea792b3021987c15c4daf5282c4f78561c929
zd7f430b608e82591678491c80b7f0d43ff1f7d0ca9a8cb62e04e2140cf01fd3ee3d8dfd247e8aa
ze954b1de3c8826fcdf6b8a66cb13e693c4969a8aa73b7a476a1bfaf8502bff0b2f2197a3b7db59
z31d09a1148b7d57c33498f8e5cba2be9e56c45fcabbdf8cf5fa3d933497646791591c9a888392c
z6407fcdf6b144262c26cae1b5eaec3b21d27c0d978b427138a706d22c92e91398e910c194fa698
ze9c18c496f1a19452066562ece309c3ab6ef38524774ee3ad3f19107af38b463626a50129c5e31
z27ae7259caeca68df48510426cd805522ad5376cd11a8e206af0bf6d7bcb8d8f6f607a0b6464e3
zd8fe113cdb0222ba351d20c4a93a3a03f4714b3017e7f2076f79ca385e475f7cef98c9a333b4b7
z216c0b2cae52c2bf1769863022d837dfe02e62ed43e9a20ae2e2988b683df171b92c219a15b3df
zb156288cacd0fcba1eb7177477c79a2095ab76af1f8db9c3d749dd89766f6a33103f35e7b686ec
z32656f493005d3e553ee379e9a4d63f3a68123136dc7ecbf23f6874a5cb04599ef36ce4f0d837f
za1e589c90521946bbadbbc068dafed7b961346a502b612f4e9e184f3e45c1cb788d31a9b4161e8
z47dab5d90282b47ea2923ebb536b19736bd68fa531dd303d7d083091332faf2cf93372ec9be863
z067103163859cd9510a3a3a37dd90919974bc0c2243d8527801fdf4912b737379ab6a5c67778c1
z54626af17771ab84a359a8ea91fc156ae5127f39ece6305a347eb3e2acf60118e5c6ad41b22cd4
zee02f8216106b8d35b58ee6661ddb35c4ee5f7220d6a5dc653fd1552b6e75a4c1d5acd2a3e95bf
zeb4f46f55adeb5e31d1bd43f350c4be4fe8d4e55edbf77ea62fb14a990bd39759edf274db89104
z31f8e09a40bb450465ce3c247608bc2fca56717830a0a782f1cbd7092f91a290664b137060610d
za1a94421a1d8ac51244d3758fe2d6906b16e3830afd76a9b52585cef0a7b5ef43b6d0cee211c55
z70a3df941113d9f9f96ed666173a7c9998123a24a17eb243580ae21567afd83bd747b56d3385a2
zc0ccc9e489fd3aff0647782cc7a94d66f59e1ddf2f3f35bdc29b7364b820f519ec69c6b8de7dd1
z71a1437e009e0fe4ad96967efff642d7ab00254b0879935ba4ec4c3c87d89146572301f42866a2
zebb4d736a486d61f2aa752af09ea2d3e1355ebf3d1d0bddc37e1e43dc213ca46855dc661b71cd2
z6597a7cb0ec4dd69d6bddd5c8d08450c250bd441eba42c2ac21ed554b4117e6216b1e876ee4773
zd1ed0bb58c818f91430d55b86669f7d379c518f7493bb5055a7cf1a5160fd7982d471fea136ff1
za74032efdae252204d908181778d1b4f28e2a08a98bf7a078b81b86974b6657708892623897542
ze43116bb8c46e167ede21a07a7b28ada89328d929587842e61a831db54d8bd14126f62b9b4d849
zd764ddabf2854421eb7fe1bb7eb6aace27b63106909a784e9407051233d0c97b96d004180ad30f
z7ded9796a2f105c13601dbf7d8342ab0c2b33277fe3d8e005c7f7c3505f0fde015437d22b1a1e6
zf1b3819cf70c63ef5bbe88c847aa360778f0f2dc5898ca7e6d40cce6b5422910c8bf0a105bfafb
z1e0cd93cec4e72486839febb0f91a575251f2ea3d09ba523cfa10a1851b949d11448937aa5b828
z8dad04416b4dd5b1cd0b3d936ddfe9c764a6c2c07da3969ef9a320ac397cab437ace0824386c59
zcf08db60379187a1e476383d09db6b192d4618046e9b5c7987673977c9c205d96484e8f8f957a6
z9ec09cbaa37f613ff975117ad17577880f0a72540e02a30cb6eeec8262bf872eadf13a9b4870a6
z8c6ca8a0f6721e7a779aa618c980d42709b5a1e63b0d8c27418fee8d51283abc515d2315e34157
zd505f92b4d2b3aad060a70ec11cfed90d1cba2cd7cc45ea9d6bed1c023c3f121eb023e289dd1a7
zfa662616d617e1d66a5d04802d029d5ebfbb678c637a29a632519fbb1937801dd554054aaa384f
zb50e31649a4c1c97219154523e1a378853bb5b60386f364dc8cd8e123750a5e28335dc1d05c266
z0074a5b52c2e020993cbe7a73cba5394001259819d1b2e2f1c968c65206b3ebea763e903b44a4c
zf99665db4d6aff2ff1de206d8b50981d4e9263d49188a20635d8b003542c92e9bd3a9fb8e463de
z428b0d29348ca0eec2930bd15fd65c7e01892db613f9915c21a732d17ccd0333df98af9362ea3e
z9e9395d179db5330d5626e7b7216877b650509cef120164f5b5434ba9d007ef8ac7fc402bda2e3
z970d86f59d9f3d52edc03e06e17c44376c2dc967a8289053f1c5e30af185e0ef1b238a693f19eb
zf9fa132255c7f4b6cd556baae92a83d7d11b8ec920a6b091b41dd0ff134fdfafcdaaa62a76e2c9
zf2a0f5844e7569147af6b58ddb750c733b5cffe2fc94f1b4efc831c5c14c42cf41965bea94409c
ze9e32f95351bc118c4cc4a5016a515555239464bf077a0be5458ed6394a82be6128f2c112fe922
z85faddd47b39f139b0cc83f42262a48bd348cef7466a93d252dbb362b58071f8b51d07cf801d53
za4671cc8447ea9bb6b0dbbb29a59d6d25d2601f9b3e2f6a0bea97e45de0aed4ff8d582aaae7a80
zd615982091580623ba050932ff7708f950b61578789b9c1ab77adaac3786c9ef51f50fc2e6da1c
z3e14cf80d4406a01779ad9a25b9cce038fabc81cf721a39c0bb4d95612d1aface57433ff524956
zd8187a9456afa1e66907de62b4a2d1f48fca5f772ae5c41eaa3d75957c766250988596fa5ea2ca
zcc1cc6330141256d701b818bb7aa5f53e48b7a9fa5a6bc62bbbb3ed1561e2068cd3e1a327d82cf
z85346a458dc019646afed19317bba88d6592565cf431097b4a7ffd643dde895139cec0a448b3c3
z4ebc007eb8c31aa1485d4b81efcf7d7b6c68e89d48fda1e23e5b4004119b5d38a88b761718c93f
z263fefb1405efc1abad760f3d559b5cd65d4da696b1e80739ef60766ff0c9bdbd5608492c0da4d
z7a7449fcb517ddeca53c03fd5170b0335e2bc64cba3938de0a7eaa21f94129166e2147f024120b
z8dc7eeb7567fd2847303bbdf7eede4b7db3ec46a26a79e057024eb4c1035c4691bb7ceaf8b7b5d
z9e75bbfd8c7505614e055026f673488806a8f5fdacfd56a9d23f9dac6787e096a3b314d7236c4f
z208bad33aab1e9ddae61aa3720c3fcfa650dd3ed6f5fe09419d994e7c1f8d1a29a1e437f5d0573
z43b0693b8b0c03a10afa0a7ae4034c6655607fac586402a97d6a3bb5bc296a135d7c2e85e97f13
z275baf015755e12431418e8ef69ec6d9ce8c736253edcc36b8b2395967ca09299789eb5f7376d0
z7838a9c8c058ed693bc68fb09074461a0e6cc23e21854ee84ba76e19675b5412124d6ae0ccc5aa
z7dfa43d3aaf81693ea699e67341d5205b77ec2abfb1530c0ed8847d334b6457a466292562bcd5f
z86425434b1eb19bd7fd003d14f30faa6d1f940168e1df1403d62054704782812e1e2b434895149
z87c278278b968ae15039d64779aa48343cbf3742adaf056719aafbd818b2fdd17a371f38f6a75e
z913091f7e96f009d5927e73af2178a0a6b7b08381ae18ed1c822bd4ee22ac6356da60c6d866d7b
z276d0a2661a488e4940632010a7057db8a3d31eefea082a6548f101897fd61e4b206579a5c25f3
z977e7afc6808f728d8183faaeefff2b907bd1adde22f5acb336cbf3d0963843c66fead98e7f608
zf097ecfbbf5b88df0f7011dbc2933630af9ee0106191fec0810832766d3f9ec11406c4d5296209
z43fe8d8c35b87924de5559e06828ffac0b6c94b3e22c3540da6c01a79d4b7f7ab3075da7ba2455
z0ac4ea5ef60e030537af328353e9ad8f710bb73062471c2728b21fe09f1e132c896965e2a6de1a
z1552c3b4482cd0f06382419a2d9f9fd7e1ec0d351babc932e122131e36188ea9919e58f2c632fc
z41aa867a8c5533bdbda0ea1f8de62f50c90c6dbea37a1a7d1e9a6bb9d67d9910ee4300ec746045
zef6c5763e217202f79b6f7f77ac2ea4b35225c76494b96385208f487f00550c73fa1b48b4c0e26
z454ef915fd9211994af9294af50116a3d1d4f3e3eb5c6594ff5289fbf2a305754e9eea921951ff
z2f3ccabe3f5722aa9a866d6b8eab085bc6ea6e2c53d520dfb483e8c828bbadd56d59b7050d8c48
zb3c072a8bbafa9b3c45cbca6723acccebbd8821c28b26143875ec1d8f7bc58bd5137040d92f076
z200c4db33115a6d27899aaa17aebdb7a4dbace37bb5c122e375701132d77cce77986f44052156b
z888b3d7cfece8d07e35fd2732ea8719330da663950a44803c73f0f140a8200b1ae1dcfd3b02ecb
z6d39f21baf08ae5c6024a7caad94aff7273964dd9e13bbd9f3950118fabbcc7fdc1f924d489a39
zaa63327741793097aa0fd2d03e2d12bb7d4c71353aa5ce06e23e9b5baccf0821cf679e44edccbe
z2007c32949446f9ce8479cc83b1fae6c89c58a4dbc3c1ed276d089d92d5f4f73f430cd27b78875
zeb6f6cfd9078802bc3945ae2f45937f480242cab89cfe568973ae7490a3562caa58d230024f4cd
ze440d024010268bf7e6f37d8aa7a5d46990fb9a11c86e3d52e6538a1ee324092ac8482a1b73b6c
z7a1b04939c5698cf7d0d88f8acfafbb7631dbeed8634e6f567ce259302168b3cb296c54b7ff343
z4871fecb8edee122a8be1b4bb1df71a3d664720d85c7f4dc29699174e46b26e94c44ac723cb56e
z81068b375721d0e35a2b254b05ac1c6aad1401ce3acc7ae7889bea9aa2540591d30272656868af
z5992f5a41a53d2ee29da9bf0a758e0df622368b944b0e08fc88d2fbcbf03c7973feb2597a88943
z0566d60c3cdd987aad622ffb853ebdd34e4b6a23af1f23ea94b8fceb9ccf981e703d2b9bb9e02f
z03ea10db6ee686a0726f8e86fec1a00a9d2dee3a5770062e67face38ab76f2101e5f6c30269628
z226c2efe585f8f594882b3d22f5895739b20f15ff10308750f7557ddd3fcd543bcd4e8192f4a72
z1606ea4fa5ac011a7f7c2542fde18bae41434e4895e3466d30a0a0282dc7dd08c07583cf6d84a5
zecdab364e1e5774b61ee0aa63362b1bf84f12c572c7cdef13adaed434990223a550563c089d3eb
z95f22ef1e3c2eb6446954c2a78288e922e84d3c06f0dde499ae4643b485638f303629dada80846
z5dc7cef944e5db56c10e56db50af8c04cbf0b569732d2489a45bfe41687860898a51edd9857601
zea9fbeef9471d92e4162a3ea94db6e8d46b6ff01a46b0a6bbd1d65262d1714d3e59e4a00a5f64b
z600129f028b49f9b0f98aa08ee13a1649eb59ceb71f2d3cc448908f71950bc288aaf699f62ed9e
z7878586900b2dd4cd721db0eb9842af967099fb22f30fe1cd210a65035a273e2ec149279ed478f
z8e961ea14d8d94ee32b8a082a49ed63a8a2d8213c2af9b802305ef5260b0bade889369f4642e61
z323fd45339bf81f4208e1cc7f8d58de0204c048a8f7ecb4f6166d32ea8c5a772491d07738871a4
zf85e251052c64223407d4972d4a7923e204922a25e9c5e9145d9f8356b18c8b8d479176709c38d
z8cc7dd228289b481228caf86005214533079cd1eca32f0e48f9fab3ca614b2521e1ef199ee2a82
z3e68bf4a8d2f724d0d2dca1d3585b2be923068a532996c2bded4e6de1270f9856ba32cc412c1b9
z3398fd530787cc094065aad9a5b5e903cffda0517ddad7dec2b5f632b90668f5d57ada777b9df5
z2d154f7a652856eeef6f49074ef4ec0e263ffdb06ed442bfb91645efee593cfcdb62085647038c
z36f376d038e71d7401b43dbd95684ec2a2c84b10b18004c3211f2e585863521a0cd4ba7919840a
zc3cc14aab5eebff6d5c1b45a174fa150f8f9ed3960710c051d55803584a7616043fd5bcb68199b
z1c7de9677ec6020d7c947a82c5301f5be418f8097554491a488facfd866cdfb146d370bf689754
z2a1f80805e2e93b973142555adb698372e4af4a7d1b6aacd2e92828cbf5079cf6ac7e9424a2f35
zf6fd4f3afd7a20350a50eab07f347d8285f2266a5aface599779c746c580b194436d1754b2468a
z6636da56b5917ed3b73907b8efa6262755af6d52f5995e491f6011889d22bad97c12850cf96f31
z6bc68d679efec362cdce5ab59b96bc4107f565be470b7951d485590ccc7a609d30c0bf7f8b6a61
zea41de8b80926a99018014d1f90cb4e0bfc8a850a982389e4e71d55c0a9308f8f8a0b23f0e7e3b
zee3e662ac874dab6ca996160156369673087ae67e19aa5c5b9094982fcfe1ddd8d99d24bcf59cf
z04fc5926fc3842c155718ce322d7e2abe00351cd680871e7eec013164e4f55f065dc199e151607
z45cc035cdfd91630f9a1585fbe1c8ef2fefb55edee85973dbc04d443e5295e5485e6365406638f
zf8789c023d504eff0bb803d86b9c6f9c6acdc10c09b5b41344ece5f0c40cc575a5629bf3cfc790
z01af7fd082a08b29b7fcf25e2c4e5e9f6dfbb1074c4fe5bcdadd438f96982107abb5dbab63322d
zaf99b5b61a5c01732876fa6e6445cdda5b4acda60b704f54512d1277e931b0adbb669373a67a44
z41e47ac66827bc251d60a25e65fae60ea5cebbb9da048185c1ff8036a7242db48a050370d61195
z6e5f8478a5e02f8c741671d8e8ebe21599780d77b17b0a74a7b8b8c39511b52b7b1b10560461e5
z830e395f09868a6f05cc775a378c9b644ef5879fdc185539dff32db6be5d9ae74e9625931e107b
zb0ee652131ae7f1c6fcb5f8c20321350bb0219dda93a65260c3dcb5a5b2b55302b5ba349a5d146
zed581ca1cbfe70bb76782b5f6a8172fd665103cce82ef562c13167a1871567704bac64879c4362
zfb9151c5cd886e68b0c3ed13b3f6fc0683bfa7e4b680cb37e0a6b347fd130815efcd6005b35b8b
zdf5c60d10a92b35ef383e35b01f1a3a7ed05f4a71538bf6f7e1962ecf5bc5090a78cfe1d569b99
z4a6bdf78e3036f22be964580530e426e19f02f5b9d0e72f2861872b50140763dea9c7688a2b9c6
z425d31167cf175d178a360786c4fbf5c9be529f4cf05a966f9d70392f7c88c17a0713e2662a9c9
z2307e5c05c30245f3f6fc19decceec3175611f7b8c66c4f5d904db8bba35ce08a5177341003554
za7f2a53796fc1502fbe461d4b9f1af65593ca35038375ae9ba6478a3699310c34b9ca0f7e9bb18
z5344f98daf204242e42448836975685a81d7f7a2b5159cf5acd7f718b12703dd6c8dd558a961b5
zcd847952749dc05ebd38d7d89a1db6219757d88a4a1bbd5dbe435ed4ff2a301f902e95b6e11ebf
zda00436905824999758146b75bcae934f30e7c759264b22cfb4391c2a9bf5c8ce98673420c8a19
z799542bae43d33b02f429b6a6e111f7a9b3fd76cbccbe6752ad7fc1a97f427fc60f00449803f94
za8aa83e5b2a61b5bf76e7c9c654bac589c52fe01a17169d261ae89f41d917adab755af609fe7a6
z014707f9870602c6fef0d45e3fb27c56d336866ede34a73add8d0b5ede5efc71b3121fff12ef51
zada0b240943012e4aa361be788d0a8959d5729e03e4907194e7775b5d76a795aac793551b33766
zef82155dcc0fafba386a488332d65ec1f6c7f50d8438acddf9dc4be11008d349f71fe794ec3e7c
zd77238226eb9df205b96710b556ddce244ae0ca0924208285b0a7ed50b7b2ce4405d14b92907c0
zad87f33bcdd750017562149e65eeac21a4e19d36cc744328440db735b73688bfd8063b0decee7a
za89dd82b83d6b8575ef6c51c16b558b37f0561c41b44f6d228bd3d25ffe1cf01fa1d554a29c896
za8aaa013151242229e8332f4c4d9d30d11a4fa7d4a11c0810a30507817d342a463541894459d50
zeb7c82bc196e9d120be7e1b3a7b51c8ef5a691a557c229704d8583389d6ddf6e4eeefe69e2771a
za124ee7a186ed22e17fdddf087df2963b190527ed5321dcddfa1dfc4b027f204257b9f807d04f7
z0d8d6a9ad8971fa0d8ad4d27617f9fbacf13a8eb0702e84b75a8483f5cc300a783e532f9f48ad8
zeadd08cbb1702d36de9b48eedb6546013e03870c8db3acdba2384822fcd21028bf32efba5a93d1
zf720cdcd4ab91719b2fe9457afa55c2cfb8766a7abbe1f788ea6c34a4ad92e66441bfa22b0d760
z30bdacf1c40a5f4d105472fe5f1df9441fb46a6316e5b572bc7c4f6e9b48356ce31776190a3dff
z61bd3de348b65509dde7dac3a3decd786da0a178cb5b5ba4b4b7f65f68596107287f3722b353c2
z0bcfd4f41e7a13cfcc9ea5ab13b86a6cb0fb1e5e49fd339651c297711a5ea63529b6f19872ad99
z31ece0dcc7ebee194660676460cacb0ff710bfca407a4b7a58882f3b2db59d00e5447dee0e1ee7
z06814dbb95ace3560519d9dd6bb75013d89da3240521046a21302cbd83e0801c3004fb1e49b9af
z51db7d9a69bc6fe6f0aaf5565a403801cf6c696a038f440ab6be1a1a50cd28bd063c39ef184282
zf2913a2b981c81b57139d41e26bb7ee68b72bbf94a292f5af4df8fa27b3a659114482c19661fb7
z91b65fe115c75876dbe1ef690334d54accd3ce6d1e9707f3d11cd2033d17556bb8384a31894e92
z8beff78b5958261c11d329cb4c4a3bcf398d290fc5ac497977668e1060019b79c9b95709860245
z8a66c676614cb6b010b4dd0c3d70de139cd3ecb44ddb7ddb3b234fdbf3485b8c33976007158a63
z478370dff4d4f123e444ef1f42498d5c3ac2a10a418a99198ba4eeb51357937aa7e6d085676d80
z80744fec943e6bc09ee6b2335a90d34d51f3c7830bc68bf37ecd47ab38a651355067b381649fbd
z0590ff1536f0a1dd9b0a6a815fb7ab5e2e78d178195f119b5f0729f306f7637cf18f1c20e6d107
zcc4e066219d161be14cc9ac4fcfd8a7cb5f800c4e954e42a879e6d5449a3beb50760e09bd0196b
zff7f0833df71df2dc341d4672a01a71d9120773930a62af2843d22587a648e884c2f33896c1ee0
zed32a1cd1da1f1dd4da4c459aa30ea39afa48ecf054e826965aa5a4bcb590426485c968436fd8e
zea4e9e1c379612a66a565829e8cf008201566375068daa4193b173daff9adb20fd9946884b0f38
zaf934a624a82a94887419ef237ee35dc4cee5b2f30f297f5f5035f0b23f125c5d7957ace08be30
z95ddf92a885fe81d817da07fea972484f9126b65ed23a3f52b8aed9eee81f8aed06dda024b888d
z4ff6a1a0369c849a7d55ed35adf8d54287dbe98c2a9de9c96cd6db597bdd5cb6fb65aa0771688d
z5668b912aefa191057d25503615049a1ba70acb011493084948b11e91ecfffcd5627424ad42fd0
z3ce6095f03710fafd1e939bb7e280de246115cb3b835cd57d2e77f93a1aab4df6e84a05433e163
z3837208b22d941c9c258541adf2f94866e1c729c98b52045ea760cbb68ea57cb82480099ec7df5
z90b034a2bed58cd56a90796740013844f594e9dd68b43aaea02aa4441b813a611c3c29c64e9d48
zd03a6e8350264a18f69315365250b600f6df332cec194d68ecf58e593853b3314a573d9287e667
z5508a94f7800319ee12dd547edd7c3201a4511f8636344097940ad0de66fe1ffa4723a2a113b5b
z71ce10c92088957800f277c881852a2cbd19c206002d37b0902592fbd1b62aaea37aeb6bcdc623
z17b1d844f8b216b7632e665cc75162ba83d6de72d5471def11ee2f0dda09dcf9d3b876143d25cc
z115f21257cbcd4dc0c4bd08c1932a57ded050e528d38ab971f9f405964b31c4ee4745ee4e18545
z83c2f93c9629c828ce0c1a36849b77f79a50876c636c13b32c9c59111f5147b26b824a469c3b3a
zef4cf584c368884ad6b486f18d1af11433a1fdb86fc838070c8d59330d4bdefb2347b34e1dc753
z1f5594086e81a357c5abeeeb740ccab6a10894fd6f170acd8b5450cf0991476374b29f764e7c2a
z05f0415938b4e5a26e4174748439467fecf3ce71579923c61e72c7cce46dbcf06e6b9e038af411
z28022dd33d435f46bb66ff7ca6d9b616a3e2f0f47a74d8faa8194f1759f3473ba08e1e294ab86e
zb8634c407bb849157694e93b3c401392048f8ffa180edcbdd70d6aa84c5fc4e66e1f3b46c18a8b
zda0e8b0f998cf0318101371b2b99f69eea5fcc127b2d755c6b5767a149c46b99b6f83eb223bd20
ze68f571c03558d42da52b6308056a98138efa163bb64f1c9683540691971ba21bde5a7b370db5a
za63e378637867f865a5666723f785274f76fe025645202d147127e2371af7a50a44086f0bc9445
zdcfbf1ffbedda9d872375325c4771f2c2ee5b374ab983560d19ca19307d190d6e610f55c5ce8fd
z54adabc7dcbd581d9ac92f607db53d979d22ac8fe3d489e8d379dcfd5d55ffc1e16fa689880826
zaf7a3a17ca1ddc4a95b176a325f2d99a5be6565ac6b0debe4ab8e33e6c260e9aab3b916d3d3c92
ze58772996525e5fc3c179e02032a2a06d5aa5b0d0f17122950eab29658ea444aa13c8cfba014b5
zdcacd5e5ddbcd87a315842ef4e7fa03d5b7119e17fa13a1248871acda5161fbcc20dc249ba1cfa
z5095c2b7a5905353a1e19f55abd11bff1111125c510c248a6edde9b4547d6c44aa5ac87d3af3d0
zda738425d625cc3b980a3a0f1cdf89f8dddaeed1cfcfcb83ccbcc40185cb1469e8152e85d4d058
zde3da9b70e9095d69b0aadb30b387c3cb3581b018b2eca57f447b1302714af20fab727bbed39cf
zdcdd4d8a7b5c0f2b8cd7826ca12a103eddec4e6c8730699abd459cff2c688bf66fbec0d42d52dd
z0452a6cc9e12bacecb92c8d484b20cba8a06855e7bcf5bdbb467f8e1054eb6d531e002c6260959
zf5a97c8181a43add7762bfd70605f7eb1dd7783ce5c81aadda18c44a4b02a439e65b282119003f
zdc3b2ed2b8285714e65f9b3b7be564729e06565e11e25a76bc7bc8b8fe87571c1de8b58f10f48b
ze468966a0a946fbee1cf3b1cd3efc953dad327a1b0e6d1514e0784d2655e72fc312a9bdcba347b
z9a421f23ba5847f61bb3019f0e09f33b92b3752484617d0d563261c8a23b41602f1e7d33c46b38
zf984b939b6343c73e754dfb473674b30a08cf23481bbf8f158d6f9b03121640d518e69c386f5d7
zab1286d56357a30c81fa0dab2162aeac22a50127b9281ce3846c4b15e382694196cf384c0ebd5c
z7a4d9608dd58ff7e46f98c72ad00ac0b76ae6517b4b1eb400785a8186a3038d22d42efe8047881
zcbd8ea60902be89916c5e69f4fc61fe60e1fdde80da1d48ab275317b4518b2c1197d79b0026efa
z86342a0eb2d5376fd1d35f241c19e471a6c031f7395f0d23b282075c5a15864d87457003834b8d
z78003026a5c3ca21512f4715da092d19399e5c635476db7669c7d3b34c71909009714d4d98097c
z80f4290ca96d8a5b2fdea800d90193070e11ffeaf78a2821f451e7c57f9fc60d2e568067a36b76
ze32bf115a2710f76ba4c052dcd4328a5c26342d2d6c2e356ef2617319186023fb28a3ed27a9324
z012461c1d8712395038613e4d0bf20ccb77ca2932917ba3241e502471e28832c5d91e76e84e354
za856198a290ee9aca9b3b3616d70d710ad2a7f9b8fe8a7d09676353d7799386f9da8eb5d1a7187
z1b1ddbabdeb87534f127fbfde20e7056d0b5244cb2a8c69aba1c3d053e060e609bcf979bc6d07f
zd73df65ce06bd65d81b95d0fdce6dc94744e822e783dcef22c72b4a53486bb907431541914ea24
ze7a0954b4bc2d997025a71c62602926c7183cf08fe0b08b33981af6c4d823844486ccdb633fcf0
z16eb581533e4b06ace60e2bc55dd2243e0e0fb78abdcf9ccd7d97218f3cc766756b4ee7a68d206
zca59457a9ea1b12d1db273bfa78dad690a30811b7582dd8f900f9d4ffc5075d61cc5dc984ad43e
z22144d828834aeabbaa10edcc14641a93d9ed5976d060b9b3c8616623a905b5681733df9b5ef94
zecea604241ee4613b05d90e9f7643491377548875abef5411b194a5c7f71a0b7e752efbe199fd4
za2427dc118c77070ead7c3a3d00108772635e7718442b04b949244a8e2b306c9a1120f21eb6c4a
zfe2419517653bfce8098098b806321c3d392efc77ccb28604c00440db860cf22b1bb4979b0e11e
z51dda7e5e2ff0a987e714d4f7e9d75fd9fca46bb430d91fbf7daa16f7b8cde0b3a41864732f6ad
zc5385172b4087b69621b99cba450f34a5989f34cf3e82ffda212b4e480648b9958ffdb1d948d16
z3eb19560e346bf8bbff5463f948c64d175dfc938fabbd1184f2cfc96125054a8e04af701ef3caf
z3cd31e5e46c7f88ac962a45fafc2a06bd5c62abec196146118b8f8b35df446b47f65d202dc6fe4
z9719fd756e62369731afcefefdc8db2d5c8df1a718e660f281efb11c37d661d813487d8cc7794b
zbe476b71cd55fa896282e1f99eaa548235afade74a02e98dcab5a1948e0ad8a79aba0da841e557
z19c999908f016bf542684a0f2b6a31084d2e47c2a2e6090931ca29972131a9d4bcd02d8e8d44e1
z586c7b5ea5bc9d9fa202355dd55ef59e965ca9ba656cfaa5a4a5d573813d70e7ee15362c32fb24
z84ef2f1ee88382458aa595ec2862590f2e71f1b9b9bd9849fb3911dfabfc2ba386f453ad5ffa72
z1c051c9d8fcbdcc15e74611fbacc29079dfc56d7464b45f3c770ac702a44d0e5a6efe25b794c8b
z18689650db43cd8c88e6844e95e2487ea76e24e1c1481650a34a06cb02b4c3d9797b8579a2efe2
z6cdf144c39a9b6be413bb65ebde09070034da14f6f375e0c5271a9b8a6394d59a24506dd51176d
z7b87cb454b5d37113622bd862f9190f8c2f3e578b5efba68858c1aa5b828b02aca8ea3f2260fcc
zb8e18972a52f7741df3a4eda435179a3f9ee851312df981e20560d5366d8100a7e02168ec5910e
zac85195b58a45d69bcaead8f5c836dcc3b437c75beeb555b883810b1d95ae3a70c7651b3046ad9
z9e918a0d627bde619804dbb05e53b02e86adc3a5b61c5d92a79f88084354c829751a5924b89d48
z353040424ceabddc085f039378b12313437f5a2594bb7c1da7759ad9a7457380360a0830137f8e
zdbdc3c745b00bee6d5cc75c543b41b5b8f88afcf2177dde506337ddf6bea1d8f3f59c54403af50
z7d1db440eaa601ba3e6940db528d35d6fcdc7330945cf0f9db99be10419bb7530fbb7b42c8fcca
ze447a89947f99a36675ead31850757fe584d73e2b52c688c8c2cb6b44479ac522355af2ed541d7
z110cdfce6615c232a832e846483cf246bf387c2d0438295b075ba4f2cc109bae58fc24c25bdf8b
z15d10c7e56a9d29ed9dab55f57bda646efc943b85a3fe071e7c93e78697ec2edce2f1e84862e29
z2cbc9272cf26b91fd895464fd6a2a206a521c0372b14f4a17399495bb02f577840cf9b29c9a4e5
zad7830c8bbca5c4712002e2a9c3e3431876878213be6cd9b02c5b94363f25f56a1a204e3e046f5
zb05674274c21d94c1e6713f51eb492c138beec82cc0d6eb926ef36485dc21dc685581a48cfa755
z152b32e660035f24e065c56e7ebdc1a0abd3fdda5c8529cc9c13981369df625200eec0a7c3d767
z64244c16f2676e97950112e662d09b4f64280aec5ba4660b54b391fa7c81dbb90aa29f54da3409
z55aed3061efd15c5f611ce9643aa4526a7fba04adf8d0512e5aa8d1d8f97ece5d469b66f060a2a
zf0f2d00e130f238d06746c16ea93209d99fe61b6316017f3cd8d9f4851f182159865cf759c7435
za11e071678ec32c173b516df25b4890e44e11c24340388820a62eda5ea7af1795b7faccde4507f
zd0c56348ec4ddbfb7b473f963f4d1007c5db045617ebbb4338832357bf1366e5aa4debc996de5d
z3f4246fe6650ca25c43641d589a2a71ac5361607b2835d6d566a5fe5cbd6e81d13f9972720ac2b
z504928e0fdba7c131897d313b67e8a4c93665982fa153f6e67878a663a8b43bc5dd56ed60ab43b
z94faca1642ca595a60dcce669511c5654ef001d38994355c18177408f63db9131965ab6e428792
z0d58528d3366a2ddc8e8a21de16dc1f247ea09c3739e3bcecb380669320d282c7e8f8836aa7c9a
z2b6e59ecb7fa6a68483783864f46d2ef7b8b09344781f2c2908db441df1f5cad5ce5dbd3248a14
z7163fe9b62938c971c565b9590633dcd6fa38a7c4c3bea99bb8a9578b625d8341510a1757d328b
z049331d7e3fcaa47658097827ec33c11b36305b9090c8451e380cdbee644587c8c3ad696f1e8ff
z88e121a7056ece324dedb9385f079a03a0918ab19b0ae754f4ea36066cfce2d35d2fd385a9f355
z058dd491b0643ff5c1b0a359a6bf989845057d4d426c1129e13a94d62c939fc97dceae821cc9cc
za30e38718e56e731e75df55a3c703dfc95b775f4856f3728ad6aa999c4b6ebde09e7b8ce7386a1
zb8a2a7b682f50619844fed5e2db75ae2b8b7be0f95e9364ce0312203c9e51d0f3678556060c287
z46c471a9c6670bdd45f267aa6cc4b6176a6cfb1b5c635328a0a024234aab4b348a8c79f0f08f70
ze7cba80757743b8e4111c082e20077bbf5ff237afeed80ceaa04db35a6a87098e1f405f1f8b203
zd0503bbb6de4b611ab34436bdefaf2f28677849f4e5797c34e837dc9b80b3b2021d0ed756cf6ff
z37c808dbc4a1c82d7c3689ffc6e35234235c64c23573c3c4467c9ba4e30bf0f645713586da22f0
zf1bcfcf0b540a870b7344f79b7e45e994091a9822a60df7902029187d3d1d623cd4e6d135346df
zad1bc13f40bb8c60649cb4a0fb0149c6914cd53ae7e8db69dadc24a216ceac2b337e17e5c58c31
z219e543ca2abe3a86226d735e05f79c20db711581fc67cdb44d2002275f5bc98d2d57a93b10c56
zc1e31e4af97d16b005d79febe9e2d1276ab4f79f48277e30c87ec6fdef7b44af3765684246b5bc
z4790b6a349e889d7be85d96a9ddbd2ecadff961efbf776c46d6df97d3c07769f8d51d7636d1fee
z7741849818dda65c98ebfa5a28a3960cbb2c8455a8a22f8e73e47d4e6e210deec27dac0235997b
zb5d28817cec368228db584ef3b5bed87798d7481d37b35f05282ae1b38547bdd9f190a201c0631
z8e412432755c479b7ffa4638d5ff23214ce571f7b96b2ffee50f7e757f478c2de6458c481635dd
z10fdd10ce4c2a9359eddaecde176c1882dd54d68822077a7d6cd6b83be08f0aef8e4a5e9f818c3
z2fc38937965c9ade4c9e591a2aba40b61922569412e30a06d5636b1d86d8bb2a4df4e108d43c9f
z606418d1e8b49e797f516a95e29e6eb7b589e060961ccf116dfd2910c4ac413637d6c818a40847
z15d15518ab09bfcac7c25e4d5ae0714bb12ab9e39d95a57cafb0e8775799e7a60fc6240d991794
z438ab8db82bb4e91081ac4ca5f94a8e6911d60fcf35042da212cc44417897008bae1917110b66d
z98ec140bc4a12ee65a1d688c32008080cfd4e3e7ce2977a3f0c29714f843b3f9371e3ffb26ffe6
zecae2e568640e8007e81f6ec82838db6846ddacd6adaabe17d1b79d45cf1d0e4c52072b4e6248b
zb4e819ce092cadcf89331e511bb090d786f0e83ff9b706465475830c0dafa9b3ddae0510c2f4a8
za1fc36792e1d7ef4594cd71b1d6e2025f97373c8108c9535a6fdf917d8af02443f5b7c76bbda47
zbe96cad72e70f1f4025bc9d0ca01dd04fad50256270439c580ce4e0198201a9174c5201644bacd
z157e9820fef7a527558ca628f3472b420bb621b7522536329bbaf3b69b8ee759f7d7a1ea8ea643
zac8101b20810ec1296e24442ac6898010524c5ca1133c0693df07d339861a1c53ac52c1ce1c525
zed318ee8b6647e69f75d24dd11994a1bbf1fd54d0b1462c416c8613b56e6a672de31f30c3f2232
z6fc614e1114028785c85cf3d8c9a22d141ff87985299bbb127c2de5e045b412a78c0b110910541
z1dcbabc0f1435d0df53bbb15f54ce326ae5b6a0808148aacc538a3dbaa5b512c8b078bb5d2afb1
z50eafb41a2f45a16d789efded66be52b64dae65114540b5c386bd70ee5594b5241ce7ec9375886
zd0e6817c8f25fc42cadec9bfe8d51970f1175ec887acbb62569ab382363385edda830490f8870e
zdc87e85d2e782fa9a625197e5e00fdd1ebe6e74707e8587c3b0d56db8d6a9c31f1652d29c9bd77
z9ed5760f03c3df2bebac3966e6d897edf290ff44983aa1f5bfcdfa96854709e42c28d9edb38086
z4408f7167484457c43f3a076d7aed8334ddeeac5eecdec4dcdc21fc28b1bb1305d649053033fc6
zc9fc51e88f730794081a4600c30fd6368f8cf402ff02c9098798e96c513bc8c26730a021d422cd
z51106f84af6d9a402a6728bd27b75e3d9d74c750b113b2b3f697f65b74799830c1cb6cce63344a
z9eadc6e79731e860471d653e27d517ff3322d46f23dcf8aece5e06be9799c583482f6f8834bdd0
z038e705bf2d42af153ad6a5c7bb61166fe56706ce54c415b3a510fedc6ded2f931010e0fcd3c8f
z7fba5c6a42e54644627b016c5534bdbd682b9f66c2eac42500a7ac7536f494339bb762326a5202
z94dded69e9628e84fa55556447e9b7e31a394b23c89ff23522e64040314795c14501bf0bd0afa3
z9efc6ad245134e541431ac26bc9664a8581017eff5f65df246f113b7a0e4fd7c5e4cf0f99d3b15
zf5b405f763add0d689382bcc3b063c0e34c719dfb2a92f2b8eae8b1020e0edf60fa6e4a94965ea
z37c567ad48ea4a00f209ff286a5c23fd22a05cbca523b10cf3df87b17341e219362d9a47ebf1a5
zcc0a7e7f7bb7cc7516940df4ec2c27a81c6c1a3e71cc9071fdf7aa20824d981164af7f7e4b399d
z0a5d381d12a5bbb2d8da7a787ef9be51869af6f9db840a1fb81b4e538a5a311359fb36635d426d
z13d03a8619250fed0bcdcb38c29eb401c649b27ba44f93e6b441f8ec675f15162c9a875a18e58f
z28d1fa8a82241135a7e1d7fc96ae56e2918fd30fbb681abbf3bf1ba3baa35d8f6cf32b32824b93
z4cfbeb6ec2b854392004806fb8db78748369c04f7ea0938d64d4210530ba1f92db2f33cba57156
zc15211705ecad0347722cc36c1ed4c692938179015fde531512cb30b4ad3670ac2a2878e35d2f7
zedbdcd8b933025bdd9c3d8d1ae185a8b1694709926ebb94d5d23267d52a7fa2420e4910f9be847
z3375bc802e0c6527538e6ab8a8f37817971ea6b8bcf2ddcda9279544ad6920a52ccb2e8b4250c8
z56116ec659aaa32e625ae2db610f61a6531552f451103ea01dd1c1b3134a540fead1554c9252cb
zefe0ab0ab8be03aa351732bd916e175777bcfcded2c007b99d7ee9c66f61e2d0d5be17712de3a4
z377556008d4d599deb912999dc09a48a13b0a33d0458f113b26e2484262bc61811449e4fb20016
z1f4e2bf28e1c1c85d8a2354a1c170cfd32fff557af9ce4f1597c87de2b6d47b084b80c70a1ef99
z1b83d6cd2acd09cdefd747f62dc088a1067b10c26b964c4d757f5fa8631ba07c6466cc56fb8653
z82248db0065d6e7041759a6ff1c0f4b8321256a20d2872ec65ae291a73dbfd7d6ad9ee7956b211
ze0cb9cb2c158db24305d124f6e386faa26949b08234de837924914b94a56fd376a7fdef6a94631
z35c257df9005259e270835a184a4f155de4f2db08897ec488aeea1bc2b43ef0333ed773915695d
zab5a0a05ec13c52ace864a4dab851bdb033ffe2e9662abc642157397d28c2f291cbfee17923ba7
zd8ad80f10a908f495ab049b6c4f62de1dcab9469f75e105b874cd26c52e8179ae4735e5327245e
z8ef58d38350e40c4db4257dc21c41c59f7a49302f0f52bf828d7174f0db9936ff291f510bd2605
z031038655c1e096ad8f2181503c9bdecb307002491bd32cb1590586b3d8d14ee487353bf50d2f9
zd6eadb9dd1c5a10bf1d4b95dedd0b88d582d15f9fb53939c7fd697537dec8adbaf8e96a68c0285
z00f38a0116c53e7a7179068812e444e65e8a1e9f9c550e85ca20196e9c6cc8a271e614b7256f1c
zb9ee85dd5ba1ec9232151ce7284ea0a3ed51c77405933783ddd176ae5c7ba18628f9b25b40251e
z55c0606c76f5f8a81e07861f0fbeed066a8b5e742246e13d222cf9109f45eb3eed9447d44a21c9
za6b6b22b5babe6e230818c333da586336ebce4b3db034dd9a9bdfa72298ead175385a6cf673dd4
zedd7fc24469b05eec8023eed30d01f9e4698c8b93d230286263a1141b3c9eebc4c30cb63d00894
zc46254183120ee0a76e43b341e869d397e7b32cf0d905e2de6c8e7b425225574a6ec9753c1b4e0
za1e319c957955129e7ef231d0fdb4829f865516c83386ebb1d0ada670fedacbbdec6ae69cf5aab
zfe406e579f44439a0a135aadf902c3901fd73e5e25f5c0f55fc433664d9be57fd22db98c40b480
z03f5512511c5ed016728473cb8e72071224c41aa84a618ba96797882903bae3e0c45485a34b9e3
za9f44b1ddcded468dcdd2751894f3d12f260cf0ffa388496e46476b1316353f740b35ef84f3c67
zc75cf382a0f14fb36b10b8584b378043d4b0d2262e90d667974c4e05dc2b4989ee54f8c0eb8761
z96f03481a9a844b98cf35c4d24da511da6716b2b682447709aaf30eb838232e8b1bd6a7a2d6197
z31d5fddb835049e4267f5bc8a1921de32e0cbfa6bada7a773932d3bb4e1385c42df9dd1901b00a
ze9cf8fdbe55acf8d0a85268a3e11268030e00077b1db8817977bb205cb92b6874cc60df87be8a2
z51b0cb8ddd6033a74f773cc86793e848729b9f1a46783f0a55243c8588cbb6041fa028b47f52de
z1b6b27842b29934bf031f4d8f2aefbd7e5775847d9a4e2e84f6d95adae524dd66d96b51276ac9c
z5225426a7fe125d06300b7eb0a1a0cd1b0ca8eb62b7d7883d63c9344be9c020dbdb1575bdde081
zc63fd7ee0aba364f97890fe7fa05eb3c424eb2971bcfd521bd23cb6b88858639747c87b9f6032b
z8aa852b67aa91389e0117d0ca5ebb604deddb7391b5ed6a4273753c4e7b5ea0c26a7cc06860840
ze22d894f08a1ecc7e85bd564ef4bbb5f459f0f3c6c38bde9adb3517d04245beb0befec29ddba8c
zdb7f2b06c35c00db491d12e0ad4799c3ae5b3f370756479ff0720543fb22de4a7d8056d1699330
z60a23a7efdc5b989750597671ae556aa548b2158d82a853ad745e5c9b1955b02de0af228dead8c
z6592fd988fbe161befd4ff86edfe65ea9d6fdcfd6bb518ef376325eefba07dcae1a58b02a31482
z69341578e5f8e6dcd8cc8066acc20ea27b8c7ba2b60d987b8af4800e9b61a79ebdf2b4690acc64
z0950903e59a48e5f6aa29eb1440a73ea2ad371e7481f0070f65fef1427df2a2b9ee749f17a0673
za2aea52c917e71fd8f03fdb35b5362d1b5a234150ad2847323e333a9a8b72254e4d46f3ca07df6
zf88e26fe26af544049cbb00dcb6f209c4c5619d55f448d42be41c65e43ef5b348248cb02fa24d2
ze987e94a2646f6576b3b95aff283e476ee61584940bbcb74517231e204ff48c1bef994b5bf3c88
zb2fbbfe4a74fe88abd088a95e550ba81952bbccc30387357640dc7a8fee31daff75d9d8038b0bc
zf2b07ea7beb631448d2cd79af57af6bb15e5e841e514fc4856c721885b1ab37a6d8ef1f90182d2
z7f4fc9b64dd926349af7d0ae0af67f0ad8069e4801b56cbc3413424be28b99958d95f840b78be8
z60e38a6342858cfbe1a4be8afd7db20bab38815fbac9cd8685b59c7fb5fab6269f340992da9632
z8c1dd1baedccb0176530dedd79fcbb4efa77ff07e097b5c1c319d0fc5ee35725e78dea228742cf
zf8c6e905b278b73cb83d21c46a6e5ac0a2ed749e0068a6880e263a10451b85eee81d7a136c7d8a
zebc664760f2d0e79fcca5f5788dac06225b542d0b2feee69c8341aef5e03ae79640c3a43d00ae6
z236fa5066fc279e87a2871218aadb02d6e9f2689adfc1ee1d16a881ef04fee803ff5f4e809ffd7
z3e5a485829a8b91087697bbae9cfb96b0e26e1b29a1fac38fc6c587edf5a1b3c30d73b5c982a9c
z233543f40d375e570edd5b0a3bbf6196f12f44743239e56fe9096fe8ec8373a795fbed10bf96ac
z44256a6293e3c97bb418e7399d8fb7561f0ce7cb61a603baf49a392b93fc03bbdf061e4ddf4e76
z36867e69b2e3367a335f7af97e18142d267394b03160d484fdcd9dac6fa395304638992a0002e7
zab34630b3e28e37d7273a656cfd9d91b657fa4f18af3057c9073b1360bc492186fa46ed0d95523
z60c21e5b9d7c9bf1687422c66dd14863e8f9453518dde883464063ce87650fe976a9885a04427e
zd980015e291d309ae888cedc3ca2051ae0dd930208e4be259529da4f8e2e6c4da10bbbc8a7c817
z5f08410222e82436efa91e5f2801271e0f86dc7b57300aab32327d6ae0604efd7d7906e9f6469b
zd991e62ea68972e5515231ce1238e76ec876a8bf2e8954062eef8e71a902706d66739746b4d0ab
zb6397ed092ca6cdb2a303f0ad10e56418d77873f961b94404d76f21688b7de1cf4cf3805113996
z326dfb6e09049da41da594f3a11f5b753497ae2d2ba3578643a117f3ce12b3048fd8c35c6de80f
z8afa96a7b94f8088bee5fa1a3f11b9cc5188bf6b7a3fea04ecbfb5965ba5ceeea27a6c2ea61ae0
zfb18687227929d429efc522c35d18b4e819eefb69794e26aa1ae07be01868a98ebaca9e3a61886
z23130aa2844802e131d31458ff4335babd75eba37303224232f67e26d9859497c5ec53a78187ce
zf05cf9b494c02e704d7654c37e163d2f2821a99d0927a3fcbed907aa18ebae4a7e1b7651b185a6
z0b0dd32a75ed08facc809cc909c935b25793d0545add931e13542702361832a515330a1b2209ff
z6b11587327531147db90bd440dc0752ec914cad207cde77a08e18329736a57df48144a7ddd052b
ze5ed86836188ba9868e3c4f1f37f7e2a2e1482202a6d3e0ee651fa07b0d40e5f172ad86bd758be
z5b702d1c6c3e8d46510c2c684d64801b0eff2f84abd42c9f606a6f755e5592fa0e3409b658dd2c
za10a8e5666936d27343c39cadcc826d5f18d4aed7d0b9f2c992e2ef98536a65e981b1a60e8a2eb
zd4ac9965e3f2e9185939fcfae3d47e1c249b3e53217590942799a6828f1cb591152c3dbd55f497
z0bfe97aba5d63da2bd19e96d5f4403bef11186d53095c4eb95f2f1db88dbc9d5d97fa0ef85f1e4
z1f1755471ebb30170542f1c0556be74cb1aedefc18d9b2b437ca4754b44db11a5e5f5cd6dfedc7
z6294ac1fc560d95d7e57ee3298a6193f917853ed31d82b2a1b2ddec19210688bc7e83294e89eac
z24daf93259fd8d0966a37064ebc768c7ed2c8be071892db54dd6932f0e8a750caebc968a346762
z78015924695d93b3b5359c25d3b6a8e994282feb1295d846e365fdca36f6dcdcbc8eb5059a8e8c
zbb6bbdd5ca1404603b0eb73cb6597775bd27061b6b01512fda9c754c71a5a421af39ef231bae9d
z11b4b2fe6024ad4112c14ab33d543a5b0b4b09f91d5076435abbe0420419c522aac9375616d28f
z60ab7a103380e208dabaf63c147dc5ba694c15a0171027e09551906dcb696aec1d95ba44b554b2
z95b21e984d655625614a1b7018e9aae246f89f65e258220c73972535a355d5916b5369c7f71c8d
z9912915851f61ed1fc6595663083bdccfda6a5f9ac12c26287effbcf85a26a371a3bd73648b77c
zf996f33c35f075b6ab5b55a84ac8e42b66a4b13df823209e8805966e1703d48523b7787b567e39
z65b70513a790f24a73cf3c5bb2f89960722fde47223f8bfcc94d5125fe26ada3286d5e04fad1b2
zea0005d03c2a9d6f45235e7c8139ecc6914d3f55f8668f02f9457ff9756e27fb15a62e3af4589e
zc043c407e0f2f3b3df982280dbcf25297a96e265448e667b3c3dfde108ad48b3505a0039f67039
z2f6ab4db21ee20f6a34aa59ba47d6be2f9b6a72f8975fc00dd5e3223d63294899a5a097463b7f5
zea70af547bf4f180ce5bb551d8e23a1b0f1b51dd3366085c3d81ea05ff01e934b852e15307184c
zc681b7675bc5857aafeca75e874e955aa4fba2805c83bb1c4060d23ae4b96d60f75a4f86c2c309
zd81cbfd9198596b8dd6f377df633e54b7e8af14d74fe6272af9320377405eeaf2fb4e6622c2e30
z95aca943e4fac32f61003a5d1048dddf0319a1550d8d1e640ad39447cc2b2d86b23bb6cb9ccf94
zea1a6d346d5840a758cc4d43da244d050e970953fb7eab931c277482f3200bbd3b332e1a2aca62
zb3fc859ee7d7565ae890c10d7e08caf47c08927d42064211ebc35693f86623036207d2ae589c96
z1065c1fa1f974e460cebd7adf922597a053d2008d341208ab5fcfb370824f8c77fa6f4f362f0b9
zef0fbfbfefb92df9b78b237081aff23e531778d3f0cb21c097f1628718dff389d30e301683a5d1
z2d8c7621bc6a42172d10e5452453608e4e9601063391ee5192c64bad58974b550e1a59d382c0ae
zb5893dd4e971c322af12e334941b15a13c333cdb1c01dbcb71e69e0951f73eb976245de7332036
zaa6a6576e10adaf0ca1eba0acc82b590008de992e91669885f41c2456a5bb875464127383c1a7a
zfbda40548fc5a0ce7b539142f4bd759954092ccc84a9adf40710747b190dab8d9a8bf2706f4085
z1617c6f49e334c8e64b6fd3e9a5a18f2cfd54b986028e2af6f7618644988a5bc09460c57ca14e5
z0e70bf17d86f8c41adb648ed31e0a2d43f9a850c25ee1b0b4a7259f25cf424fe8a957f8d5fe7c9
zb0ed5a792cdc0ad8be12f3ea82e917d71ce564299d519569356d2b241c2d8fdf23e1533905a019
zf13d1da6bcf23c3b5ad8d72e428a30d29726e4544ee2412d8a1f74cda34ab85176b146089dd1d7
z187c252e8f1a83ba8df0dac5a9896cbe3182fbd9e18ad900d741a85544c52c6961d18ab942b7a3
z2d182f9970336dd38f7f9e4f40935212b41638e70c3f886fcf9026ae14b30032d563ff791bd423
z3768c44de3fe1712a2470781dba2f9cea06138f1e3d9beef2929fb8d8f0c9ac411e40bfa1fd247
za9328d2eea10f9b33a68f8c5734b0b07f30be8552ac3edb8ba9d97ef914971fead28dc12adf9b6
zab51b2b9314dcd5a07f3520b79aa248e5bac7a6a4687466e41573c6f9c4800684046a217d17607
zf2aeb803fce8d6c129f42765ea6851e218ab06010d54a29982c9b4343bba9af86f10dc149db1bb
zc6129e51c1cf0badf1f1188cf9faab590c9f9b2944c21792d9b9291d65e5514a2c03c6538c81b5
z0d7026f1310c3959abe52f07d9dcea793c1130521e92d5ec1e0bc65e4e4ab11bf5f57ea4515343
z618c9422186facd3d89fa7f993484b19c02be7daee8356dc924c4d8c506d0bc7a7ab566c2d4f52
z8a2ecb41d09b29ba8d40d73043a3a91844a9c143b2a62cac5faa285d29350db9c2f5ce9e715334
z839722e0c29c73ede69d8ff75f5a9bd250ce678bfbf45cf4389dab205fdd41898cf208a1285fc1
z62a299f2fb4f92b8de91ebbcbd6c5b07f7c959cd92cad1d0ab776f95cc9b9020ed04eeddc98dd2
z07d1ffef340d5edab09e2ea671f9c936a23f0463490727e35c82a526355250cae248d21bee6e6f
z8f80083dd31cd1ee14b1f8101051ca0dc08c8f92938a318cb8834b841e1bb263131920e15c35d4
z82d7a180384b2214bc025af6cb810ee91bf7a22c20f59a8287a35e68d19f227e33786c289ef10a
z93ff50a2b6e052bcac6050c706e7641c524dc743804ac8359e2e00c95d8e51d2e0e0aaae38b817
z6e050f39c934ae55e622aed41af6f91f11b081435d985ace576b208c4bafe034a3759fdd825f17
za56b0723a674bce24ef4083f492300bfd4eedcc22e75a387721f78a3555dde634cf8bbe87a9dac
z2086c1bbdb86d1566089b0d61f883adc8ea79fe92e36eeb9e572baa94ee64b3f66aed2f62bde6b
z746762e66e358dc97c09a26ffc612187db92202f6ed8475d894424dbb522f97df272cb19dc0248
z716134e70bb249a35c45035776e0727c1c3cee361a6f9f3b3f7095de1cdf556479e7be88a5ccd0
z67eaded82ae3319a08c91d62963b00f318d5c8105edfce74c2d673d818a6e03af978f0ddbd2a31
z8ebb6529705fe73d265699791228c4562e354f96affe9660678abf97431c9d47a53e797a9fed30
zb4b10d6465d628415a164e2d676e2db283447f6caf32f8703c4fc3697cb41ee16118f2a3af10ff
z6f439ae9a81dfc99e24adde0401d23c7ab83d5c3b77e0008eb9ba73e4be27682c631419e0f53a7
zf2b1162c84c554e5b1898bf0173de4c0b9903e7a0bd79b929731301521bc6ef0f43aa83adfb53e
zc711fa2f8be975893d3c9b8ee7e981d8ba2a01b5e241ad037bdcd6db4a33ddc6fc440d9b117b91
z7c4bc8f9514942d0b75418320b8f7334268209c8ec38049100e6cd8031a4cfbee934cbca7ad313
z90e6eb7b2097cb0042b3ba839a96ac7772788767af55c6af5fbe90471fa416c68747bff6700e36
z4841186b95c9e1354fdf05d0e046a3fa3759352983a359f3836546c406505b6fd23fe33cb9092c
zcf7a89ed2cbe0239e8e04543938dad3063fec836498702357123974f2c2953cdb6e7b9893bd6e2
z9d5c24944dceb031d502988c6b2327b0e3387b92305e55ecca22f4e6586073f94420e423294e69
za18b07ec905db1ed3ad7c904bb03e3edd471b67029c5da575a3f0595c09a3f206b1b1cb831333c
z34efeeb7e05e14de97ac2c0124966f4a429fde799583819af8aca59f7d884678ae85cf708c37d1
za364c950e3cb07b6e79fe87419550b8b1fc66286540a24c293af316d14a0ab0c6ff9f9c4c5d854
z0b0807f1abb1eb36c93d77ef27f67d55d2f287bcd7f44153faebf097fcf10c3e1e4eef7361d4af
z36102bc8d098b1fe2b40e65d9cf9322a4f9582271bd1e776c8b3956db30180319e0d213e87325e
z1ec6a33201b7920738a488701fc7015a6f86723c5bb8cd2bbd1a25ddacfd19c9fa0c5e292c9859
zfee7511ffe9fc1667f784fa2495760163c7dab6ce54ceebc034dc47ddc4087f32f8d72f55af83a
z96dadded61fdca2973718898f7e71b11f0f4c8c33d40e6df67f2d34487aaaba3898b9981b6dc60
z58d820b29148d5e8e4f4d5a088bd99b1e1245afea335101ef32b5925cb6168a69b90bb1185286c
z7c2d506e67edb3ead2dfd0b0d99d5c8ceea709520f9a3817480e2cb1e5e33687c07d4240bbde8d
z3aac49aaecb85fc53925fed50899f09c479aaf32068c4b991528f240e82cb5fd818a7452e9a3b5
z02d89a1f8355ebcf99accbe7fc743fe781f7a843d6a472b4d31a4572072eb8581626a45033fb94
z5c9210ee26c1243025a9fefebb771499d82e7b0ad04ba37a63c9752296d61b9c05537778d39b8d
zc16696f841f8ab63c111f7977d5926b739f215a5d73178e6b86f589dc3413bd527c3d3575d7e33
z0a7ac52e6969e968216adc95a99be9fd87164d50d412981bca07032cf2f44630c85068cf3a816c
zefbed3e53dadaf3fa728c208deaf976183473b5102e9c18e612235d98a1158fbd0b5ca0fd2e243
z3f091a8a5057e69490240777a276d775730f7b5c77bdf6d120d330a65ed79bd4178973c90e2ed4
zfa629c50971f6250174e7948b840c586e9185adfa9050d796c8f3c0bb8edeb63d156118aa80ec5
za17a36da96a49fdf0afecd4f5d7b9c3378b300d47e10c619f544f7d9d967eef0a3a36d431141a9
zfabdcb7eb540401c54619d18bb964923001095377bb061a0f6d250a1b7abad843ec94c4c4bd0f3
z531d4b71637f1e879b6892fa0126465f5cf8b51162ffa364e4a4c8c93703e0ccd5f80c1a1cbcec
ze2149753b07fc0c2ca3a129c172e5dd585facd29318d37bdeb707d35728999622ef410ce4e08c4
z934fd602c98d76e4ab8daf09a8035b1e7d2d9d15bd9f1eee67a1075eb5a0ac02614953737bba44
zb62d51a12ab2061f6cb46158cfdff925c0b49f4cd1168fc29f94b316027645c8ecd7f41e5e3b43
z37c3c1b69bb01e1380e771d7dd193c343474a7f16f4be6860b4183a492aa5754aa5dc95917ec13
z88aa92e01a120584689e5d59773d27ecb0108502c1238014fc7710fe2d9e90d75dee3997ffeeae
z94ff848a46063ad0b02b02e1ff121c2cbf6c16494b2d39daedb11ad82f7a0d1e45b42e3d1dfaa0
zf2da6803b7b6d640841488ff7e94a8fa89b2b5e3bd7c74726b00d7165e85e14593d4e323fc297f
z44bcb5447e1249c6171b273c2ea09fe7d8b9954e9d57abbc666c7651f732c4f1db68d2223d9c7d
z6474769e4f8a5fa840f5b26ceaa1a3b604fda433be4b6375c96f4115a85ef1875eb5cae49a6574
z490f063cf783190e10983880976f35da7e014ea8f68eccadd814176162b3bfcc6326390ec290ea
z0873e4bb5e559b18cc2972ed033c1f68a21902269158fffb540503acc247dce831014980bcc657
z24c141f1ee68700bcc5223d14bafaa3d3cd6083c506e2a5da411ae6ff32d57a151020fd7dd955e
z179b7b99b6f59ac54590ea8ff9c9540e998e1f20e8115eb8e1c5207ef1c21a32bb81058765984a
z3b22febd9d9fabf4552df9b32178b12444bb116ac2d9831f54938f772be30b17aabb951756e15c
z7b672dce47ff121cf4f7b1fd11f15fe955f3ab0fceef9fb511144adc259e7bf1508ee27f01cc2d
z5e3eaf84743a4601e3cdeb13ea24b378337015ba94971f366a83ff067ea777ddd4ab76a189b4ec
z984bbd4c0f66fab342344a328327458542b96d19a796a5ad5a1baabd6b9b6d939016b741e927d7
z5c792b7130d3a2435fd05d73f1415762a1610065e13941beac0ac95fabe255b0e9bf8abd0ed71b
ze50fd2658bf2ef63cc3f0e1ccb2b3d2dcd4e0f60d164efdd715a0ccbe11bfdf4262eb5dbf770d6
zd5314db831ab7cc4a4990acf985379db934c7daf96c96f7cc9961536a9f55d4385e37de7b64100
z478489c87ca1b11c8b465cf32d0ff84d8aed7b7b7c3443f1b242ab6b91fef7587b02cd5052888d
za564ac31455709a67a0df019f7679583f21996f7af80d7ff14ebf1e2e187bbb4744fb50879a843
z53cfdb1ff7bbc4988d1738c09afd9cd6f22dc6dc5f5bdfa0a969eaf84af2062f86a1ff162dbb8b
z863d895f34db531c8b0c78ff4537e4b5f972fec9237eed827c3ad566573444cc07473d5ab1444d
zfcec48eb84e74771c10e4ba5a8932f6ce7e161d687395afb2a0fca866f483480b124685f0b27d0
zbc969545f650b3f9ad990be1b89e7ffe033e71eee877f6cb6e096470990e3e5380ba19c79d03a7
z6c4fd77d743b9e9c5023f77936cc74394f879da59c10ef53ce8588d5859fdc6ea9473a3f6d8470
z6dceb187942cb0c5f9c41538399e3d88aac7cf25d11f75b5d2fd4dc3159070646442a2d2cf515f
z4eff0245eb761b42102834bc4656591e4975391019349f88ed94654d335d2a56a912527cd39365
zde6d43dcbf81b2e781834fb1ee1608cfb30b44fa248c9959767a7cee43a73385fb68e620179019
z0283384b340d8e83709f27616c6bb42556afa72fd1437a741f2b9c4d97d88e2cc4efb78e0542eb
ze49454d79546fc5651f25fdc48ff77b176f5054ac53f590d62f293490968499007cb16396299e2
zf1d7a03767bd9c9c812b9afb60e70ef77b03c200bb28e1277d5c650a0a511b9a102e55ea841914
z4a0f46a480f8f4bb2c4141acc093e8ecc6111356d58ca2ab4b139385905410abd7c4a3b552f7bc
z0119374c37b8399fa74840c986a42cb2b2031d94b08a0218ec67c93953dfc15892428fdf7c3cbd
z6733b221f9d4a4596838eb783b199bcb44bce55ce76d1b7223ae07f636140f1a34612f8e526497
z9101730f4ca411f173f6928f0bfc4c93a3eb62c711a2fe907e36227fabd8a443390bd76e11606d
z7746929bf323fbcd8b0ccfc3f8d7c83264cb184bfd316203947d96bc08d2cda68c15e8fa9d49d5
z10865253fd5cc7437c4c0a63e58fa746ce8065b0bfaef336c8e5fea6aeb803bd08920933f87f47
z06d0c511d577c13838550733dd17a40a75084ed16a512ed19baaf5d4471a80a7bab373f714a9a4
zbe1e1fa19cee61b5c4d6b4761a222fa5e08398a4d63e03cc80ea5d9721bbc5ce82cdd2d4d4e21d
z26daeb9b139a0caff127df71055ffb87fbd5f63390747c1b4d92ef23c8f0b2d9044afa64b1196b
zaf8f85e6d47a618cbe2dc61500b9a5bddec497179e123c3a2ef0978747e1d3ee6d31c9a5afca94
zd4664263aef5da764a8b143b7386e44f38823360ecd16e6eea76eee6289729e920a9fe4a3a92ef
z0d6ed79e2696bdbc16bc89908cbc1a90e24344b113f0bca8f96a5ee67e664510778faa36364cd5
z0e62389df0810a0769c4bcb944abb3bb3885c3f2b657694393e3b028ca56884c3185d2a3b74e45
z536d1505fff0c49da378d95e5a30468e9b85a3ecab237f221bdd2f57c9f21c01769c63f6ff9560
zd10267734aacf703afed449ab1bf42a8d7c8def91c2783e266370fd1b3136b1acc70c2fe12b812
z5531a9c1bf9338f9312434f459e190be1a34a86c43e5c34e83f6732e9c222705a1a66768321a07
zfbbf6baffb35081cd7d199df171280cba29fb6549170adbbed02481b086480963f991fbdec9280
zc18a8eb3bf4656ef4de11883f773425f010f78a00cdde8e2a0ebad13692164798abca8dd78537c
z01ef0ce2acd76b546a4639d55e0d34b2828e39662304b128cd5c093fa6a6e6b2cc6fa282133566
z858c1c05d537a444f012b4dae1f1fc89befe2afbce49f7eb1f4d92bc23b87ee5b30d4bc913e658
zd0b986a048428898ec3ceaca9837910d7ae865c2edfcc857ce457ad2084c348a0d8b838b184a2e
zb582ec79020047d6bf64802d54264c97294fa9637c360d2025341465808aeaa185a237236fffde
z945c41931536527bd4c75aa9570e2fc91100a69f5c9b0f61123fac0f8eadd9ccc5340b268f0d7f
zf9ca76538fe2b50c40aae1d5e58d52008c7d19b1483d593037d1e427a2d48e6c04162d980903da
zc26fe0c0af441a64ec04e7b00c8bd6244826023aa712ca657f7c851c5cf16ad739a84280715c32
z33728fb48c9c8c0f9e118196e36abaaa1a9d53725bad9bdba8280bf3118eec2b7b008345422d5f
ze7f02d3f884d6501dc6cdc6820449ee6484b367bc8095b033a65d9721e6f33382b63599f9e1624
z9601017e285e4f8607cbca0b51e37c068e8a2833f085d9e1a89670e39d5025a4c4b3c95f6d58d4
zbba9543c6ea2e942aa1847fd7837874b19af4750be2b2c44bec92121b9193b851c66a7041bd0c5
z0b06948d851d81de71fd50c8f143850de4fcadaa3663d2975dec070fde92d0650cb46198b93443
z8e6a1a3e8bd90e045e6b20eb0757693b3872fd2f3888784c3b9ca2d8ddd14706779eb2cdcdabcc
z0bf04cb7c71b59a0dda4a1bbbf2991ba8758deed2beec2dd0017fb0cc8ed1650a539bfff5a7754
zfd876aeedb87a64a9643b2f4edffc612f67346f4eddbb70ee48815357ea2bdf4dd28545aa22c24
zdaa98d2ca1010576c6366f6cc3cf6e84745019e5962323e80cb8089eadd80978ee5d291da4a969
z6d1ec74479b031016ad2b789ebfdcf4d114a3eb2be19f68642a2774afe3b1febfbc945a21af0a3
z46e9f2c372d91588a9e13a4da77ffd2bf3441b5979d089fd81381c02fb7339935991e17343ed0a
z92db01caf4f5b06914c1baf0c80cb575fffec0fcfd228b6157e9ae9472c7898d835d3d2ea039cd
z6d8c6e9c9c191f53c5d46014bbbd76ba44043ab3e0d1981f48954b22abe1d40ceb6105db7d3b88
z575ce6a8964f706427192a6564093faf5efe566b9129fbc44302ccbba523b2e271b69e4152ac77
za534b6fc6bbd54de76d7ab1aaea18ae7dedbff5335dd66d7bd5de47c997e43b267255fc549766f
z48f00113735e49c6727122d742250b6e4bc04adf805f65e92463635e356786863d223d6dfaf241
zb2ca671391c36046d172e7f21d942f7030f3d2adad067dce7877e0289e19459e401ee2b922d0fa
zb767f683255d47d6117287704dd1e3e091b04fbcb4052d0c3ce76beb8313f6c3fca1dbcb392d95
zcf29d39b7beed99265906a69a679d6162425c84de7a79eae5f962ebed62d563fd83e9e0c47801c
za7a7008697d9950bf99d28665aa0bfea004df5e4bd84b8097a79acfe9fbb4162a7f444472d7c4c
zf2249c70847a7b5fbe6d6801220ecc2d34cb4bc5c1a10331f5f94d62de99463dbe03c7d15cbc76
z42e9ad9d1ea61374f941109e7fa6925bcc6a7f19215d13722ad80af114454d60b4529564aee4cf
zffc515729f9e166e865badaff446de2ee7751d0b3b5e1352050951b3522b72ca9a76020064d641
zf533bea3ed1b13774bd49409dd6dd2fdb40e9338e550bafd6841775da2788e34a2407b9e4b85cd
z8a867372887a51d4a89ebd3991e462e44d1d466c046ad3210d44a59fb54c9f3573b11d593ee1e3
z876335bee061fd87e026711dbd6a77ac9518c41b5b827b5dec35a2621ae1b3abc8bb97ef33ee1b
zf8f93c236114d1873a53ee6c2fdc775975a65dfa495124fc978e7168363436dd292ce149741591
z69f93956f92718b5ef89cf68fb5465b599307d9e19448744be3ac9f49863e35b3c0345e9b83f82
z2b5bec2f0f3f5f91d24a6404947e84021282c2b6306ab96c922b4a0c2901a63d3b28d5a434de6e
z95883209aafbaf4a82818844bb8620faf27c686a5ad133038779b944f532ac8b7afe4d370dbd50
z377fd2c3209228336da11bb669748031748cf5b9c5dfbe4526886840240f126d78ccd13465d6a1
z884e3ac2b61bb4e0f9266efed59c2bab5234a7c488cd2d614b673e05f758dd4e39ec5f714283a6
z19de8f569ff13c9f6c981e2e6f9a61abd960ca475221ec1b22537a176c69560d0b446978f7465a
z474b5a15ad8d5f072c071fc8822dd71ea06897cafadbf53c9ff69bc2a31731eb3dd9d28031edf3
zf8d04d01f323d96e99f3033669cad26e7d7c74168f8534bd01baa18043b015cab152f6492e860e
zedd007d06bad3317614e54c9e17ce2cc91345bdce2256edb472f760c5ee56e77f1c37035d6acee
z8a878d9150b8dbeab24c5102d67682b82c3df107934bef67c1671c30ecdc584a1dd5f0c7a6db7c
za925544a6540ddd54854486f052211a68935d7c94c25e37e887af1b809eeafb1ca66d4d5101c46
z3086f0cbf1d20dd4d4d16de2104f9ddadb36f9be1262a631cc030c90f3da85b2606ec069ee7551
z0c67e992670055f5065d97fdeff31d337f24e79cf5892191cde60c9c5e68433dafc4da86973848
zbb4d64dd46d106aeb2069544b38b8d9405bc98277a3efb6a3bf328b7e84288aaa3ab8da7b8177a
za834e2ecd691b9f557d998be3ec9c3979a017c3cd2e246f7c985bc6d4c4e1fd1c8a6aa1508275f
z383361ff37c2f50a55ae89e4567e23b74e4db0f98f35d0f0be91b0dde52069dd58e0bc2ea3e9b4
ze8ba9d2d52d38c2d5f19b36ae6f446eba8c4826e2cd91e72eab4d1c6df33b11d1748321f4e12b3
zbe715c17401d7a81c7cfaee4d7c73d49ab9098757e9d43025a5d06f2091a5446779568551ac705
z19d8b2ba27505530d1094ba3cbdcbe3ea27ac4fda2aed7225002a5f5c6ef3679b8e67d87ca403d
z8eea0bc6ad1ec927a064f9ec294dece1384d92404ddd566a0b516b8a3dced22954f8f6b75269f3
zc85d2a586ae8ab1f0d0fbcd130acbe672141f5005fa47765326fe4e803184f33d6c8c5a3afb2f9
zc0cf2fd08b43571c149720c54b6b08071240856824be965ae501e517bdfc40c4d7b065380e679d
zf8e345b32d485c1c1dca41ebd6f83ba81b7821eac653bc89b3d1bfb6e3aae674241a143babf093
z26e1bcbceb4955af598b356096f185a529c0a184d3dabcf09d45f8db1510c9b9ecf3010add9e5f
z864973b923876152f46d0cdda5fad052c63d1c3dd73499ad9453b9807b9f2fc3ecfaf5a6c972ea
z47fcdf5b920dde7f23318121c729806f29193b8e9ad58c58cec4b8a8c107a0fcfd4b9cbc771c54
z72660ec9f71e6ebf484576cba507f71122310dbe1ef3e89dd6c0d76a7d04c5060f9278c807bdca
zb20534e9ad507e2ad0c399c25e653754b883b8b40eee97ab5e925e168b79c8a2acfc03508b9bfe
z3158f6806e44eae19d03ebee416f7525ce42d430994f08bc9b584662bb52b161f2f3c13039d8cb
zc59e15f35f7468f932d51fe2f158b82115f813e7a88bc76f5a4dd5fe3483e4d7e36bf0937e4fe4
z5dae5c9e2a6dec2731269f5d23119c12402450f5469ad04c95e0d5d6dff0ce229f44cefa0b7da2
z5ba9d37c0d3e44ff1c081513b026ca663582336275551fb495223b1c79e52401dd51825d43040c
zf677c871be64529773c186e16c2f862ae046a18f9a72cd5001b88219a7261a671f4ec47779d0b8
z46f2d2dfbc65ce196595a6346293ec75051f7cba1146e6c4220c348153c41f47d0b3deb181c367
zdb4161e7fad62896a4a3aaa7994b6459e24be1ca30bede0725866ca434ea7b99d46c5783a8fcb2
zb585e5f1364b090e3ac96b8ab94ce46f8144aef992364c6f49d4ab7002088e2ad0517ed5997831
za5f45a580e0c4289e7980d3bcb8e7fd7dabcbeb6c7f3ec6201318dcced5081e8288b81284e0bd4
zdb2c16552b4f7e7d649b93905d1a9e9269ac8d8b5e47fed7443035144b44f75c0c6af2f668377c
z3cf5a169dec31670d86129ccfb1b4e935ba8ad6fe200a79dba8173dd872870a3dd01e0648632b5
z4de3cae785ab050e84f60f9acc3c46b84532786a1d4e5580accc64b0681707e75b33974f300e63
zcb546be2f09fae2db85cd355b30df2b6caed834821e23117fbc85759b92269b5e7b6b9885197f4
za8ef7bebdc1432d392cb800bd29a79fef9181d04f123fcc59788ffeb61af1b54086863d62a9efe
z2e2db4926d62c1d55b3be34e500da6b94dca7bbacb48dae4d138c099ff46372b2b92f03385bdfa
zeed4ab143a3316a93d7192fb5920c2d3441d093fc9148634eeebd690ce7287b7518e1c9aaf8756
z7815c0022d4b1382272f8704ba7d3bb7d36670e0ebbdd906db9e69f67468fa425554ec7680b10b
z83e1e101c367c13f6889d04359c3f6a5a8cfddd50489037e1587e156325cd6febfb734abe86e80
ze0e93d94ba5d24a5d9ec91a6806c852485c3a9df6f1c1626eaaa9272d7c057c32bbb2836b4d827
z1dcc015cd0dff49716daf99d8a86a17b55eafbd6a53af833dea511a55a9cba45442611ae57a7fd
z8f2076124a4174b8e24923f874e4fe0850573e0fed3db8f8a35a044471191666625ddc6a84745a
z3c05c5f30ab33e1721076cef9b3f3702c451249f4eccebb0b8b15fc40ca431c278855a2f8d0b85
z55332b598cf0f72421a4ed55a4baebf398ba370f60146cf236e33754a7db7f2d7adde19765ccf4
z91119c0a6e928553cc946672d10bb48b75fe86114ff30faf801e10af1176c59b7e0bd8fbfd1328
z6a9e9b8098bd6ddaf8f1541c69ebb6addbac633d9528e2db69d98d60fbef32df0092dc6cf48bed
zc12fbbd4e4fb84022dcc5de67a24ff50e6ad6f27be1e4f0c98fa9af12f92c5ba8e147ec5dc8242
z675bb9f6cceb3a4b1ecf552b97951398612b3cf71952bb13358ad5df4923acbc9cfa7a36ed210b
zd6ceffc66a673c2745ffbe0a4379d9c40534cc41c5c442ac75869810f5eb8d929bf6d92f7eccab
zd7ec36777902dedf2b3e4774ec74b92bd46bce38074f29bb792e81789f697888b40f02ccd0cece
z7c2bd6e4be1b1da82b73a83e35256c4757441039b312a93fc63af90cabefa6642d205124c62aee
z57862e772ec400b016e7b35817a06ee824bd67a1a28226b63d728882d6dc9d008ae8f8c6697ded
zc2bda7690d33f1fd4bcafe401c462d85d6141240d21f39e30df96440b6c77130291caf51e444f9
z23ea65815b635cc69af9856f1b470c8ba0f4ab089f6153db18cb6c7d80e9df29cbc198aea13034
ze63acf8643e183299ff1054655f88b218190cd3a8938308e440dbffde1999d75c0760ce0d047bc
z99557dd5289b0b713576733b7cff1ade6fde3ea3f40b1fdf86d7903ce28fee2196e46c4c4e1552
z9d9934a09d372317b10b1bbae489f8eaee899fa946a39a6fa36e5064a515600c970e12e12cbac1
za0abc5f95ea02a1b2cfbe8025efcce24fe6cd928c1f0822567643b5870e079931ba252635a243b
zc2e20d3148f3cae7fb09b738137b1c216b5f2459f0260993d3c2d17ed08446d85f1ca219288629
z0daf813e97815bd210bac78fdba54112a94c2190458931104060907008a900bb9946cc2691cff0
z50bb0cdd0046f7debfc3514533196a86c226f5ecf7505cf613754b22cb2a35224fe23bdc94802d
zecce53f3d9f1b5be1c81e7398538e3673a490a8b52c582cf1c1dcccab3cc1e0e9c905aa40995a3
z04fcb6da9521eb91a645f8c02e6b123ebc2017ef33348a1d3155a93f6a8d5e8abdf93f3b0cddb8
z8921fc45de96bdb61d6efaf698481452dad28068bcd123b5ce89cb8bde0416efd31d5cf0b17370
z02f335357873f247ba2adf04eade991189f130de651be3aa5385fbbdd65843a737ef0eb026a5cd
z2196aafb784a1432506f28dd16e36494a228e47df6879b6b7a8c317dae7a72b4ccce93f1626bdc
z1abf366eeeede462cf14c5aae3d69a792853988aaf53123e161ad87905798d7544c6d4350b424c
z53e2f2dd5be9aeca0468fca4905caed29e28e64f6aa8773b61cd5a1e6d5c44ed9f1d9a3961f263
z0af67f565e440e9ad6c6dd7f494de088e5b7c9b63b21e6f7cd4cc38680f28affee286132e67a30
z8b27984d5f295dca9b2c85696be07bcc28d8d8b1c7cf0ac94b4d3aafed4c32bb9931d1a8538a1f
zc4c596d5bfc1d9892b1f2c68735c997d7a25fb6732839b6430242c8e0c2e43102eda2b2aa8ea1d
zab0da43a87e8d3bb1315f16e42adeef7fd29b451d9bb3ca69f010cfb56e72e83155f84db4137f5
z6fb019736ba337d7207231da64a4a19f927b8e5d1a00e2a95902ddd1dc781645b8e225b46df292
z6d22a4d9051e0ccad7d3ad6c90a8f91ce6a3f806b64ebca84c74ce94b23d0073740660bd86d4f1
z4658ef731e1f7066aa56cdc25c60aa31d53f348f4de9d67f48e5d92e5092b60ce8a6f9cf262ee1
zbe1e9cbdaadb97c918573a1158925a402e4f1e791bf86c3c3107b31e42bf4cc946a1924c8f376a
z20bd1b197221a94ad0c247340eee48521f536252f551a38e51b64389b98606b02e973a1f52d6e3
z81cc0a39d634be8e5e1e4f676ce6948197755095bacf7bdcd3bb9150c7d4cdd3301434de144179
ze67d2c62dc612d23e1b3ff69a1fa76aa12c1638563b6ad36e1d9e5303733cd0bf01070494954bf
z2b220be14ce67c60e75b82bec385d2dc420bc9f416815f5109772a808269bbaab611a108b079e3
z649605fb93085eba379d9d058694600334c01e0d4724dc8a1632fc292ad6008c98b143253c2f4a
zb7d2d0e78d844d616f0fae7bc975d0d38a9f4aad852695900fedf629fa1013a71fb290f13811e1
za8c0700e59832d481f94b328e966ecc37621c11f0d056f955ddd6e1d211a067755a2123d97e4e4
z52fab21b1970b560a7a27819b9ed111908c27443eafa34f93f8abbe49f3722e3a51bf737b32a5c
z46e890d6b3e7e56b388b1cfa13faa9eca20c915e874e291b7cde92debf36fa8496ad87a69327c8
z2f027058cbb0bf82d0cd1fd9c0ad9f7d398569d1e3630a219b58644b59bfcb145c02c15d08b485
z83fbe0d52106dbd077e92e9b4e91d0adc0ad21589ccd59ef5417525c6e1ebf86f1489311aa7b23
z0ec42f2af5fb2b1ca90b50ec84d5a6fe3d0f25b2c22cf5ef85bc25c2e6167877a1af2e49c6cf9c
zaca0e4b3b649bc2808d3799c1fdc6e905082de74f0f3f675881742a64b44625a93741e49e2bbaf
z01308a7a107f23aef5a8b432decb5eab1afe1579992d9e98b0d41d927a49c1675143d5e8f467e3
zaa889311813f53b1e877b325221a7b4c5e520e4c92932e791fe07166d77eb73b5fee32429d1b22
zd67c227bde739e644192ca686a806eabdc5091515e85ac7c89a0b173dcca82056ad3038d8bbe9f
z9a1a6932067706c2b3481b017ee0d0938b4aa01a02db0be34655998e193db1a38e282d81ea07ce
zd65c37e0b9de97aa2f5d66b3096e6743ee74fc6eb61ff5bcec34ef93eca9f753731097e0e531dd
zfcce1d910fcd4c7d5bb05fbbdbd9bc1d43a2be6d6116cccd3a8c93f79d87f01f8ebbf13f2f824a
z160c35ce89fb8106d5df28fa17292026eb4a3e38501108351ebec19ff8712ad45503e9baed63cf
z608ee0f423367c75fde557ca6621207189c28d67c892c09e75910111bb0c80ec1eccac008fa201
zb9fd4c8842a1ba0a6e1efdc05af28ef816ed41cb26809a547e82a738fdc9fc21a2c55abff54385
z8f282f68cb8522b9b8e228ad8cb04b73751cc38f8eae2a7907b6cbfe9f69c8305a0603bdad8882
zce92adaba686f05a54714503d72825d5f02cf9b2d3f1511a30af10de67beaee10ac2cd6b203799
za12bda0f2e36b90f3ce1a0dd353abfab97f60606f443a70fcd188e9ca976a67a6683404e2b4ee1
zd2145f1bbd5d940d4f610e04b33fe1c3fc0ac877a6c0109a68a9b9a022eb09c5cc8cf3d582b336
zb485501efa095973fb44bedbd30912c13d3b1e612813d2cd2f1f5b4b1bc2a9522c2c0cdaf27bd5
z4c7ccd4557026d9cbd1965bd14390bb624cc51422aba41997fe19e7ca9e4ef4dda750523f0d43f
z83e333914979c533487a3386567b65d3fafc65c9d730455c3dd92ad720edef643a7fdb4a0b54be
z82e33f7866c1f7cca7dbe5b4ee1bf580432e7573499a3825def40465bc4fa85059c0f815b6fc73
z78cb9459066f7968ed94b05e522b8a09102d2fb3e73ac2cd038dfd2e8699a8c1a6420097ae4cf4
z40c7093292552a9edb9c9f082dbfd83e05ea10d8c63ec6fae1fea9b6fedf311cc4d267a8f6bfd3
z432b3106a19186fc086436ba65cff4180db8fc5b22b146a78f58481a6af288a45abed98cdabe76
zfd37759223deca3d7f7dc57a745467fa29a8dff8ca69df8277f1fe06ea869d847eba50b4742825
z823e2f3816ec2b99aef58e874ff107b38562fdc9ff29e9e92d6cb729650088dfc89273aa49c99d
z2c559ad79932ee8ee3af11cc6d9fc6f4f5a937156c378d7c58f106e57d7ea5e53cc2085b34ed12
ze6a3d05e02ca39412f2011db8b5e896c8b8605672b11ff95b6339d1f0cce808d706fc8f24ba63c
z717220b3abeb55d86f15006be211f88575175be653f9be4f3e353c1c4e8112818eec332e807fb3
z2f26fcdce13c2be373142b555ed0981e83e59740dc965a2477ecd51fa73c8ef696751e5534a379
z1e819e1c3082c1375920d19bb2a5a27d3f2caa4ff592976738dcb9207b3a6049c6e8706e2c281f
z5d846e1e1c1509c855e9d3bf47d94f5a174d4196f0db9f770c24b7b897083da01b9e5c88cb0b9a
z121610473769a3c9b5db7950b43839b28a4b89b53bbdd9bc8f0f48e207c70d4e9e081a8f90e475
z9b2ab2f5ea105311552dc03776dcb41b01b01f9b1a403d720639399dd91d8fdc499eb4cb7a01cd
z4d0b115a9a130ad4b162fb646d4ee6ace73bd31345d5222de1db5b82bf3978590582b1fee443d4
z7f0c41886c6af089394db086370083c25eea1757c566e17d9c64698ffea79fc76c4528048b065d
z4748142926f8559c6fa39061519c7cb415e8cedcb98f1d8c0086c6031c3330f5385575584b0d0d
z3102109133ce0f586e6f901c4fb90518646990dc6ea8122fb5992e9044c9fcbebed50c0cb55764
zf2f2c9ba9f5d57a283f7b0bffc805cdbe3037f778914af1e5d237bdbceacd10f48da1cb7c307f3
zabfe7f04dbed6121435e45d54b75aef7ac40da3af30324dead4e383366f42ad1d77ab6981cf73a
z9acff4d7a517fd0e18f6bf7376ccacfcb03d1c1b42d3cf836e564ce39dc45d7d582fbc176c388e
z648a5d9303c16c7e3c0f3e25ce0ec32c3273fd54624c7b5d86e7e8c3563f586d5bb9eee2ef1dd1
zbcb061da346d95e7ede762607a8331e77620eae98c8cd489e705c6f2294f66f5a1e2df0cd1e177
z69390ac516d208bea114d7d7997d015447a86fbe073eff5ed1c95fd5409c8a642d3d5870ce2e4a
z966d30cca72faf546290de575697121d95a989db9419fd80e037a6988e72c24c25158c9f2b73b9
zeac2b67ac5c61dd08e473d5d33421fdd7c225d01f9998445ad0cefa038968f4da38a7a66ce164c
z7f936fcd213dc56fc108e4f68b4f31f2cc1c8c33b6280cd56a64b418d541e41f1d9be51a0598fc
zeaf7521307896a5056095be8a619ed68785fe911e043e81e226da00f1f81a491ac322709096a16
z1d42e42307af4647d97d4510504be5788e6e1941f2325ce1b64e15f3a0565ef73d6ca0f9e388ef
zc82ed442a95eec5192f8f5d1e671fce135d0e7415e210d21d1e9b5c6342f07b5a5946cf228e899
z09d988d9105a6e426a5141a3b1e3e1373da5d0a29162c0a876a5ed8a175de37a48824a10f10eb1
zd122164d565e02de3ca6286c53b69c760c77ad406d821bec6be83391d22df2a407a43a01c5cb48
z75ffc483b6056d99b14be82685a5635bf465c7d0fd0f5859fffe6461321fba8c5ebc7f4d7a94cd
zd0a8e093aec26563ec8c30e1bc07ded1471a018acaa0002fc36d0deff50c552fa72311c6dddf6d
z3721e4b358f15fb02cae2f723217c81ff11fd40c787da8f5e735c14217e744ef04510a762d1d7b
z99d75660a28cf8511fbe95bcc90a4724b42f4f28fdf9549711933c3c5d5df7748134a018104e86
z76b56abffabc3cc513c158540beaaf6c27c441fb56890a6406c5e2a3b2e1e0a625d93b1008c1f4
zb442e19d86f51bf431b73c5f4983a104381b5ff7667cb9d9057f21efed73933e7ea6fa59c3a6ff
z650cf508933a9d14d90ffc8060c23895f49094985d88fa00f6c8f0853450fd43a663ae457e6dbf
z3e8a512eb2132d2d9a8a2970a8e012b8e8c1d67662f2b56fa9b2d3072b69021f31b1af5ea6d0dd
zf8b630edcc976909f318a92ba0045faff188203f50c677c06d1d2d04b962c18baae4039921989e
zcb5e322837a32515d335256d05761793782cc65105e6979c2d7657b40b83f5e876581f65ec1132
z9ad166e4002fc2b795071f90f8976fa9c497ca9b32cd3ea652eddc1ab40f0461fae95b4b7d8a4f
z2c3fec9a0b99375d17dd1d9e6c5a731647463063abf5f1cd80ce311f168e00126911599885f898
z9f15767ebb83a9e6891e6b5270aea174bff1a5c11e72e98bacea2fc4c37c26ad5594f89a3f4bc7
zf2f77b28ec404c592cc5cc7574537343a0da6c78c46a0b880cffeb2d7c60a56b078b89c2d67c21
z865ba63f07096290be5b409e228a19c7a0261471c0cf9ee86b31c8f039ecdaeee9a113b16f7740
z1cd810251605016380b8427824ea1f36f040112816d9ebdcb535c7bfd26201f5e6e0c9cd420e6e
z69ca24ea6e4295c01a0fd29d86bfa79a7cdf8ec051803a2413de209f0425841ce051c02a2fb68e
zb8d2daad7879e1c627cdc7961d0863c4b6dd07a7fbee6613b77224154477c13f306edcf00ee9c9
z2eac7dbc3d3e28171b11f7124f133098be66c6e381be9d505c133b845bf6c024cee07cd09142d0
z7de20d72a07bac7f8bca76e8706ad05dd3ccd10138ee288eebfdd5eb57b24c71f10504474ee13c
zd5662755fee9e10de9f4a3fb57c5f812be874f1d1f021f9b84c6aca9c655cb9792d7ade472e29a
zdf2b42851980c7adc5d4459d46e5a0cd17d9b6d032492f286af3f971777dc353cb886a7f43558c
zfeb2ebeb9ffc66aa3c84d0c8f725cbfe04124375efe572eef0a81781c478f12597a068ec0a4433
za365ba47d7ca55fcc15acbe9cd9e121f40c65197c376f035438b5a79edcf94e8bb43e9876ca7d3
zf940464653aaec94cc13fe39928b310196eab358182d376c160133b9b93dc82a4d08ed8386b5c7
z12e86c78151ac1bdf623226fec4403c65badb278d14fa473ce3ed056f7f218756c945175a29e09
za939cf7b599f72dc2cb38366e012ec15402e954e7d61532b01270e3b7bef840f4e31276b1e9f3e
z5be7256d59b2de755522ec97c0e5be7885fe3c34b005e883d6a25dd47c75de96595b7e63ffe3a1
z01c85d06d981cb22bd7fa88ecf3bf6adebffbc5e153cc05c3330ead83f35d91b98946610229de7
zd9f4c35d5e2f3b21de43e84e0130d20f39a3943229357f310f94ae8fb5d5b8215c53553f30292b
za7ef4ab427dc4aa0ca5331700d46552f5f3149442d93f565db845bf650c9918b00c094969037c6
z398e798a658784036c1043e8ea29e7000c5889f242e3bb2b2351e64d853f3fa23d3715ff0b8a68
z59c0c64007db5cab4ac495adb360422fb4f152a7c5f92b44536738c22db17e73a1c1d25895c586
z2a9c33000f479fa5ca970c1db2349da68c381146114446078ecbca2d71c25f3700059207a1d398
z7b61dc807f2d1aff004298bf7e88ece116cf74fc46c0921fe3d8a640acb862db6281143c12117a
zd63419556754de51660bebde895ea0a24d0503bca9cfbec95049f3d2fdba0ddb4938f9c9a289ad
z14a2ff8860a5f3694a01f439bb08b32284a807dc152e1bb5b6c3c0f76c2757b19b0cf56f44f2f4
z57df22577ab5a9f7f488941dd7628d6e9dd84fa00f0f2883ec6033d222c0d843cd789690d5de46
z4dd114d5df37b5c22be0d9c3afa27f9a8305b0db7a11aa2d0d5aa544b97d434d9ea05ff3729c74
zbcd98644f3f57661d8b556ff46c5d5871d97062d40f953f2b68d34720daa89eb6c2bcd4dabfe86
zc95ddbb9df5ad79a8e32ed11b1760c125d237f0f833821e0068491becb89a0dc6e99fdbeb281a3
z0102c9de8de22f0e63e2d6f30c3e92a5c81cfebb770755e161cb46741660db12acef0d4c6259f6
z1422aa13b05a2b97dde283e434da7cf74f690e5548cabb8f257541f9dd25fdaeffe244e46c0c48
zfe4d1745db08b78d79a89bd57cbdadc995d65d17b42d75e16ed0df7b93b224d5e67a4038dfb4bb
z6dfe280f5b17390bf747fc6efffa2036a4452de9034be52721f89b2ffa4c3c3cda0af45a4ca2db
z1be7b351861834fa9056171872e19a69e047380d9132793a4993383c963a1244e9d746882f8780
z7d42ce075315c2cac921a646017e7d2e5430a40b0192b8e8c21dcf3cdc36ad0054e585850e31e9
z79d1e80fc6461b1ea844f7e339b8a9403b8f319267b54b8d7defa2c131468f181f3a29ae47a65c
zcdd7e9c4efbe5a93d680679fd6ad08b89908fb97a625fe6ac57dd081a3da70f40f44aaf88e617b
z1077f8b5e1d2a4a854c2ea94accae67072a7c0656543daf45f2a02373a1f63663e650e0447b175
z0d606255930972762462c807c7b1f9367b707407496763855bfd2a8a707e2e919ff82ba1b33610
z5eb3fd745833d6d5e2d74e17e618c50508b4e10589e9be4b3a32d8e05e0a52ebf9c3391e07372c
z30dfd44cb44fd57cfcd292fac8457698a9f80bec7f7fbd131a1cb35be7bfacb9f993af84d7d4ee
zea43fe89eef118a12fc980000fd957344649b5c94e0c659974d2558562c6189edc6bfb8b8e8f89
z0d615f760a08cd5897f920b8cc94058cdea9cafbf7cc1ef95b5146568b08118d9864e9b5bad44c
z5c2a020e0ffbac1d6efb319327c08f29b2b79228594492fdd48d134ae43da62a4decc921abbe7d
z80f4366478fba789eedb074ce3bedfd1b1405c1c691c767656e3c31d1e8ca4d439d3ed70e4c6a0
za202f8dbd06612a6eaf249fdf7570a4bbcf96a38dc6cee514c9716c6741460a289f62d027dd782
zf41f9f0cdb4701cfdf115a3e5e2d56dabe2223100ac24359e010208148a033c4330014e101603b
zd61f50bafe0a23d2320a8d0e06b04ea46f48ae907e79e9d0f26741fc4fffdda3ffadc7ced74bc9
z9ecbb3e19d6e8031139da52db8e706f9c1b6e6cd093d67aa4952048121416b857223569482cfee
z863ba9e5dc07e4a98dff20a67ebab2f4f262925d61b3141c5fee07d608d8db6afc7f3c40e22f6f
z7230b15d899e13705f04f9aa77f775c1fdbe306d2d16facff642da170795e9e5af0777526a080f
zf2261e7b09999af5077f78d2deff48338010d9f6535f92efde08d9385d8e13f3c0c7dd8a2f751b
zec91fe20c4525c266d4bfb8b36ec5e5ff86a5832f5cd70dba27a640b04a9885315fd07cf4ff93e
zbbf1b23839954edfe0fb89e9f773017b9218f23e1b5b4c716b52040cda15c7df54ec2f72f0aa5a
za8a5297079f06b1b0e4d3753d24c286eb9016239f07847b00aa0907a9b6494761a03a0ed042575
zc50479996e977bcb89627a9f8f7d615d46ad75f876416676d30f7c2d9167e4f292d0ad10ff9235
z93d88a0194fb37a5cdb93078d15728172c1ab7dbec6ad2a2a04069fc6b0edda83e87da0966c285
z5bc83e4d330d29abf6dc58fff3cc1e896fe43d56d170f2a345bf825ae7c9e8cff9a29dcdb4cc4e
z4cfc46acb343c2600a46abc01962bf031fcee05aaa17ffa7a33913fd7cf29f0a6b4a07b4c33723
z218da4feda017bcd1f545fbf6235c916a2723825bd05e51855f69fff4264fb243761797c8f2147
z03df3714f3d6c1bd04abf9dcb934c8a6645eaed7cb7cfaccd4ed6af7a56445c26f294e9e83e5ee
zb7db7f31dcc8f810992c15d5201468beab8f682363a845762f6dfa152aff12cc410346cfb58f0f
zc0f7afc90962a70c5694bf2b44278161dd00e1ced3e96fb90b6ed03417f175df7019e7aec799ca
z557e0026231dededbddcc2079623857d835d2fb3d718fa8e7a34884aec3d33b865f5f9a7e910fa
z9d049f76895243b66273c87f511bf781cd0a633a12b40dcd68908b4acd6af224131fde56e496c5
zc4f311bf88b26aebfc5ad9aca4926f7897a9db3cf5fed5425f3a95fe890b055ef6434e04db5cd8
z3139eb740ce05b90fca0d5e538195411c9d6e9d52267cdb1266bd7328b697194499ffc9f1f40b5
z77825d675588b0cb5ef6948ac9f950723150f8e70e360bcc009838c6ae3c7fd8f27b7b94cdef65
z74dbb6cdbbfd76db4f615c58a2ef1377f21bef72f154baaeea5efcbb60197e2c1addb52a48ffd8
zfa058748c37b72be95f76db0f88b80c36c3e5947292ccfdac5ef814954b7352a6ed81b97029d46
zf2c8668efd8864aa8c1570d98321864c0dada8396adfdf09c89ff3f0a9ea30ccce2ec63ef11572
z493ece2f84f8affe7e989cf1c497aaf9a1eadce5857a29e8ef7c56fe76d3112d99ec20f1b9575c
zc0276dccabb9005f85291410646df236a188f3828f6737c1b5252cbe5d97a67bfb414136458d5f
z8781ed58886d8f60b8309295d088892d901a83ec3e638f7cbfb8239afc4658ba5e9077e955c49c
z88803d9410d50deb2f9d7064346305825fb08618e1be8dbc8c1879f87513801d776fb52709aa02
z96bb2f1039658c484537a33d78ae486ef7e83d2a85e14b41da3930d89f4cf1e938983a914239ab
za495b60472c113073232bb57161e070815fbe6a04b2d076b056f9dd40e2c35da05f4fc2ce39690
za9ba45287207d9410605c835fc365d9e2b6fac4efacaf4509107e1dc9fd3edc259038662f5c1cf
z6c5450e558b9bcffe8af04ec261289462bf70f9eceda7580d246cceef6fe1099974b8b2d4b3955
zac6b978adbdfa5c9ebacf58f050580b411d8f351033f61d22e5cb4d56c9992fef369f0420f5785
z42315eb24f1fa857d8a9b067087d8875af01846dd29a8db2a8f0481c2e7ba6edc8c5e28fc31c2d
z9084f2400ad9e767400362b65ad1be62a23e7a1e13faf2f2ddadee21e179498e178f6575392aa5
z9c1ad7d05e747093703300e95ff8d6c64b919e091c4db686ccf413a6e3ce4dce92b6d590febe19
z23609cdba33aa7f67db857246d13edb9ff4c7be4cd560fa42a6385c72376bdc392c500989db2a7
za7c056babb301d0cfb78e3317d068b126de7ab12ac40745b84ee616daa06f16a995c7d8e9c0f7f
zd8cac4a2656b0fa20ba505e2b440cc2b57f4555bb73811bb74a3c59cc861dd3b515cb45b50c2ec
z47f70f4f6e527b979af2c0ecede1da65ae78628bdb42c4c3c7215385f0e3c3202a6f736b675867
zf667411114dcc971b4a93b7f168c83427ba743fd66f5bbeb7de5b742851dfad2bae505fc4899b1
zd4e409112241b623a3ce99b75f202af62f9506a3a52151fd8c3fb0f29f18b1297a5323ddf701b5
z0fd4978aa0b8f9a16bb2970d11b6b5442f8526eab0c055ef5707eccf4bfb9ad291dac89dd75416
za9c252d4e30dde4676185bb1a22886ba04a04f044549b80d9ea088e11f3d221e1e01214c973d3f
z63938089d4b6015e39f9fb5047a192de362543728a5b7382041c5c17df06a77ad19fe4c00f614a
z92de10161d97ed7120e2df6710b6b22ae35a1c191861f3c263501c228b02759c034c704b67877e
z4398ceaf392151c3d516963e853903e50d7ea87302790bcbfadab9b79a70d58089708d04654d6b
zf63fef3fe6c2e561b1da243bcd776cf5c1288c868c6904135fcf12bd0a2aa4a255e51f2a9a171f
zebca8216576b0e6f87f07e556603ed0ab814fa89807726e1bf653583657e3ee771edef881d9869
za0091ff1975bfa020da327dc82fed2e32506f0ed078c0417e9823a881f1c8367552b324bd22381
z1e2d6d966860aff8c0ff350c86b869a62a7958f29d53ba7062afb4544454a501bf02885b9c5585
z4179fea1b83c371b4640307f0d3756cd414d360fa4735855a18a6d7b0f7dcab7705a35da298374
z300c366720aa8bed3ae42e7ba7b01dc62d5386c45972a62f5c963e613a472f4ea812c13cbb7831
zac65f93e68e92fbec5c69c4c803eb084f43b0a7683f7cea91bcabfbabe92dfd2e6142d809799f4
z6ce42bda31929522e20a3dda000faf87d7a385929cc128a78f3ccf360de0a49416c4d629a913cf
za67cdc3e429ba192f5df85a16701e6a09edf704868e39d3740e586ab48b4e087e73a5961ad917b
z6a11e1f1bcf1d183651b78156a9da92fc0618f54f87df55423c68852feb217e2bffa3ebd435b98
z5140f72d67f8b255e0ef358b95eb8246ab4c37bcf12d8502546c5a6fa14fba6c211df552623f97
zcbb529cfd4098ef88a939a659f1a1335e9732a4af01bc770a4255deee5058cbc7e7a7eac7f8681
z46f17682f6cf76226271463a39d8d5af0ef2344315ea2671ff569b1af2255ec951f34a7f00a6d1
zb94cfcbb1e57058ae4a0c07020f159f40049276e2711331e7b06923e40edf22171a2bb882968f1
zf955825bd784a38f79303674496a6ce3415b4f429d68b5de8a2849de328b8c4a7b995f2c563ebe
z05f4baba6c0174f7a30d8cd8afaa42b6d2204f6be7fd381ef81ca6ee67f54ec2b780e88aeb39e8
z0e5d9dcc4476fb2a5b57a5c0f8d437e6751c4749288ba3f389c764ba146c031c0412179ee20d05
z6790b23f358b89e6d182e77bfebdf4d9dab4a9af82ccbd7512598b21d59e58b2ba69524f0e9e17
z9a9d62ee82efad0ce9f395fb4a4a252293fcea38b2dd07fe25193c46db6c4634c84693bf9b9771
z614c5394ad86652f42556ff48edc487abea446013373573375d4e5dcaf5eaa4d45950b12769634
z19416a3291db7f1e776c1cf46516f2792869fc74f071b1ec2100a7d9e68d0452a40641c8d0db3f
z1ad642a4539f5a4aef9920ac33844139b4816add3e7f9966e52c4cd2db1bbf9eba17b10e6fcb2e
z1e955569e4cf9437d51cbe6e83d6c33f2c9c93656c6128efb6d07ba865d7e970130ecc431dad93
z9f9726b1f92572dcf45d20d860f6e5b51d8dabc6365523d8254f1deb21f1a521d299e657ecc98f
z0ce634ad08464e9eea55d0119c9e3ea5c344aad96351190eee2503b1644f54714a211d40e25010
zccad188e6134b0af6fb0555a669936588c7862755ddbc9bf4195de4e7e538a4df73d874755ec81
z5a0b8ffd9b185dd71137b21b0fd2728f30d99495fef46d22dcef03a4f6a1895fb8277c0b397cf1
z7acae5b937c5f9224ef14fd354077cbfeb2eca6cd067b0fb9271f7cf152f378d509218a8bf4ac0
z07fffbd09030edcd3c7b42e9127d8f025be49027daa27a6f9f5e6274a239b3ac295e9c933f8865
z117713c6eeaef1e9dcad13e9231289d33382b7b03255420f767944a0c621d8f76a0bbbc368b8a5
z9d9fe304fd26ae436e70721fd9595574bd3323fadd0ed2f5f4b7f70dfa6d3cf2ece8bd65615617
zab6da6571f433b811d0b4628e453af0de756f55af2f5f324c1c7cb375863128fb2a64db0386d80
z278a23493940dfdf0c8e87c1fef6c487596edc70f1e74065eca9d5060b7f3c6c84bc1632ffb3aa
zb412b19dc3a546ad3dad7d62923acba926ca670cc214c40a44e63df0c75b0709e49c2bec3aeaa6
z9f4afd779ca34aa005cf60d0034c890bad4b08b6b583e8cf13af26248f0ddc06ec910779e38cd3
z92ff879be99d6963f97231e577257f91a902ee0ddd6a132f93ea252be35b1b9dccc10ee13734b3
zfa8867dc730afe54d45b0d9b9802716d2dde7182ea2cc432bef6ce573a0e0d0fab7d9e1bbeafcc
z8af265035891495682e4194135a43423c7a0eb3f6f481877c3d33f52e30caff483446f13a171e8
z806c537add2323a6bd557e1a4a55aa6f12b78f66e899b814e0bf6d87f671d62007b621bd1358d8
z995869a98a85bd1a4a1fb34547e508d192e605a4528c1ebade7cc25e100f8c773366a9255f1115
z38029a0cbbcc7a7539ec5547872fcd27300b360625737495f40dc905839b641d134244bba2eea5
z02a0f2e7e41bb7c43a43f43ed50c625ddce77f398ea47b3556a05a1c445e083837926c3712e1c3
z1f7c0f24ca789afe8cfc0478205a731426f0870bc14f7ba65d16d1fa88449027aacddc98b04e7f
z7729dc5174a8413400260c0bc4554caabea8c317ba48f28ab1b07d7af75c0eca7bff309710c5c5
z492c037f5962e3ba5eef39b2e6ee3ed07a28d5e41bf9487f195c2231698cb7badde2873b3f127f
z88f1bd11c0b5b22d96d47ce153ec0c36568f61f5631c181f56e863a4c4d0a07ae4b8085e2d4e4a
z7e7ed1fffb4945abafbe600c1e967ceaf3dc57b5e7ba40a2fa19b156ccf3f55ff47621808afeef
z2eafa0707a2aa20e3961dece75d960b9ffbb8c61b02ce831b9533cda12a10426b76104c65eb9a3
ze965eea8b4bd06969e522486fb2f69d9f441d00a78118911323924d3478745f2ea3938e4ef91c4
z58ffe00a27d7fabf63bf4c3714a14874c6c7e02ce2544a8525c30bcc6bd8cce2088ffd8baa4011
z8866efbdc3c2a7a4af9f9d74d6820800ec1aabc01300bcf169b788b904d171e733611c47b7d6f9
z475b098c601e84701b8389403d709a49826d5ce0d26d3866a17ae43367949b4262b1bc935fa8e9
zbb3d0c979953c3d02730b61b938584620d515e796ba718b39636cd9b19519bf47e532f66463fb5
z09e5619cbb2f421c7ca621c983a9930edabd498d6681172b9f85a40c5c2d2e2d03a008d68e5cc6
z1433f352db862870499ba0609f480621c85c49a04dfd29e9a17c59b8d9468e21f85b7a8bdb10df
z8cb6b67e47dcacb557decc13ce82d7cd7ae8f453d37c90670e31a807981f04613af6d043057a1a
z0d7fa9ff611bb92f143b50dc7dcb31f579bb801588d89e1e531bbf6208c654a0f8f0718159daf3
z758d2fc2ed8a8eb80ba8bae78f942e8c988cbcf123bedf399bbbcbb9a896fdce1ff10908a9d204
zef2dd48f0c4a2c776a0fef9ff87e15074561c68e49850bc5824dc4891c9793852b04a6f8f7b203
z7d11d1e02ad5cc4ad89a9dd591ef7848451fde71ac80b8812763c5227eb94e972c598c7807e9f8
z1ed54aac6deb2cc01c7a2eb3bdb38828369c258c96fcdba71da56a2b392da621cb3514515eaed4
z2f61563141f5fcbcaa95fc086d91861389bf13662d18b4d8e10155e76d328708f45bd89cbed4b3
zfd3575b88c6135ca37bcd513611ed883462cc8de445d27fcba82b05597848d0108c39199caea06
zf0dd346e598fe31e1a2ac45f9f937cdfd46c96b3be60b7abeb056238981fc879c7919cb2318b8b
z4c61f743b55b8d59222a56d5e63a21854e240dd5385dd74b189fcfe8b0eeb676c558ed5a0e896a
z7fd1454d46b4f7df56ebfdaafab236a2e22143b0ef138113d7cc4bfc70b5c00d21377a55dec9b5
za3e07639527c0f4cdf649a04008e34a42a88dcbf246ba203fa1af30ef73376ee269c2adb121a95
z831c99b0c5ed71d3f1a8974f1feb30e8aff8ed6e850ba9b759c8f4c2ea8c0ddabce64ce2ebbfe2
z310f1086fa563909fd6ca777f23671ce08f19b3abd3fb8b55363d8bd8f2588101c8904a1de10a7
za406af840d1a1574ff210eff4762facbd5b59a0bc5c13aa41a7145761b54336946f57ccccc7fd3
z08bd6ec4dcb17383634cc3d517bf34cf8f3263be1d19736a752b88cf5b35a42fe487f2240b8836
zf7ca9215d15fbfcbe2ca889fe633f572fd5792955e34e37cd02414a7ba4bc0a355c2d13138136f
z2616e9c62a9b44d8194877f49366fd109d1951bb2f946c455070fad1ea1a4bfdcb9813ff7649e1
z93f59f8decc7ff59f57c18bca0eb82ebfec30b96f35c87baf9eb086138a54e802a5185a7566ce2
zae9b8c4fe2f9b95888537ae50cd94bff2616ee33eae35718ecf144457069f81cd0908ccf87ab44
z1bbbc8566c279aaac63437bb7924869f8389a968142ddc025297aec81bb6b27f99b36ec3c4fb52
z818134bdd3d2a9b4c6f9197df0a69f89eaf43945851a643bae936dd9b96858ba6906774116ca91
zd95261a1318e40f8891e8fbebe34409dc01a86d23ba456c49074c91593b33488c60d1508b42fa8
ze8d7ff8b705e59b618d515001b9de6446ef964639a809e77986d35f7e8ebfbe6bf1f6b43abfd38
zc68a94b5d1407480bea7b8cd677eb89f42933ecc04e53e83ffc2fe8783233cba8f5cff22f0bd12
z88c1fccbdeaed3f4395e2a5bbcf322763952e996e7722e4ef196efe764cc20b9e409221b47edb3
z25c642fae64bac02cb6f80e2d61be1ed0a08e4e8dfd38186da1b42bc7c19252142c39bd4c370ce
zac4e4cc012fc82349ec45fe7d1a14dceef55ae566e8c97eaf9e6a18f21b25e7ea563bfb18a5741
zff5e5727d9ad140d3721e554bf6462c2dbbbac7d335a033ffe7513fb149fd94df8ad62c6c330ae
zfb310841e079c9ae65dbbd82bb6bf9f3b00a452ee12313adf81baf2eb23e4db7316421b5908228
zd7d3c0ffa53a1314dc423e81010fdb5eaaf0f1b082375b9b579010e492258ffa6f77aab8f682a3
z19d9b75408755c43d4a95a79f1e03bdf7ec4ec1a7756cd7fcaf481ab4d848a497132348af67ddd
z083504e1a4cc0262cd5579b11c3bcc363757463009e4f87c5ce07f26f5fe7790bae33546a3cf63
z9922202ac594e0841d296a090ca0f836b681fcf5caa9655608f6cd39917b325daca9b1ee2c7f61
z69384afa2858d7d6ecbb36516a2504ef2807ccdae95dff1db4b5f087bca9bcf66f3648e0ae84aa
zbb4a736616081d7aa46d5ba7807ef3ed16d21409d30bc5a341f8ee0841b40921a026f9dd139b93
zce3bd93c946d5aa8f83566fc105fa01782760ca9642535b58a5d66c7a0d98f652d80d5dd3439b5
z40b8829bdbdcb3a39413d2444d6989d7b6ce57019348a2dc12263ecefe90cd676595500dc502e8
z1e859b7655d53961ada9715636bc4da2fad80e2ebda1b7e359260dde1da313030f994242e0fa63
zf15072d2c2bb223a436efe5692395aca3526eb59b84b1fdc700e9aa36a13f0b866695e06fb400a
zdf1037085ebdcd8d80ef05dc0b6413893cdb706aba12a20dc0edd3777873cee4b9b0ae9230a5ed
z212ee5dae27a9c26ce51c3d6af2bf6e90fbf17e46ecdcf51bd61aba88308a24fd678a4a1c25625
z77529ef00a4f085d53dcbf95f926751173ff3f3cafc4fac789793dbc7f8ed20de58264d0e6d713
ze1e544bd78bf2d35713ad9ab6229238a35aff73fc4fbb3ebf29e214e1e339ca968aa41611b33aa
za31c27216226b886522384d34a3e9e406771d68604f47bc8d3663de784f4c2eed28b6ac41d4ab2
z3348a0b7da9eb1d0989f729ddf78ab491159051e8531589585995358089b3f65a124356dcc8331
z4c52af79415e1ee9fa542b5f247d61c870b192819326a19cb544fb550196b9a118a9175f912bb8
z3f1ec8a290cdbe15a95f40db10216160a163fdbf440df8930b8d0ed7870d57f679f5f4bfff5de6
z209648cd890303568e168b95dbb106f1edb55f062684d20333c58c518f356dc1ef24405b806c23
z78e23dd01452bd0654f8362005529c6991ba129bb8a1b883161bf85d611930c3777bc406f89b62
zae960c4bce1abd27a160e8907c3524bad13c3180eaf68729d5d63110050ffbc0f1d737e79613b8
z4a29c6148a06fe5f38af362f4ac6ef2060cd9c43ee3ba38f7b74dc5ef294477de60540f3168791
z60f6f214e1d0931593954188f634d88c7215682e8bc44d214d433df8e9cde6fe210f91e55a05f1
z6b06e3355315ca3f009abb7fe6b8ea2034f5da51efa9d8745729b607d38486fc16846565bcb4dc
z9ef218c3972c528a69c8084fc70bbcaa0ae26a9dabe6e59689255d8e39205f1f8c1266bb68c416
ze1f0f23f34c3cefe8d659c4410756eda21a733008c0c7337c9b258a3d1188c3fab836ac82c3702
zceebc60f343873081c4c0da3bd90ed6e008674e95dfdd5792a9ad689ac4faef90d64a4ac11c511
z9a738ccc4ec9f362dc63a1279986c31b3b1dbc78e5bc1bfeae7fe220268890fedb6844ca60e805
zd4364a919e34d236bc61f2e2bb5b712011c0fe2db1e7df815d02e6a670f16cd1b4a48a03f0ccbf
z9fa3ce16fb4024e8e03f663096d26f6c0f0abd019385c5046c2e12852a003d0a6b34ca8adf7297
z8c2299aa257f52ec38d1fe8f851f459a3074eda57a22a39994c701f52ba62768f5857cd1c4ba50
z8ce6e5ba0f7a43ea6be837287e9866ac1c7a7dd9f2d8ed8873d9e6ef62b755b0f6b4b09b869cf8
zbcfe9550815ec247b7aef10b372d191d61b2d7bada4c2969742165e802cf424aeff8310ef84c9f
zf6cac369fd0c101c0734fdbdb7e28324e3fb2462fc3b4b5b9005fff3c46b0fed6de5a7d508e60a
zcbd37578d5bc52a84d5e5093ab9b7908eef3f3e6db6969ccacb5a74887a72a28d5d658940e2f58
z185a696528ee6dcec4cd0d7acc45f715f0932a5c390ac369bc7c2a58f0cb0b0fbe8016ce18cfe2
z3b186796c17e538d978c4a5b623b2548acd4591493498003796dcecb3f8d86a6670bae0b7f61df
z54b8857b9c8b7ab37a4d408e8fc101ff9122894145f95bf67a138bbe22abccc3d0afca3ae2fd72
z9a2d6f708f8650feb3b7d0691aab0064cfe1f16c81565f39aaa6ce66f74558b811aa4721d44e6a
z614251145a539704c00bce548d81c001527a331ec1116b424a9af77e5ec93ef08d2fbb0ff8b61e
zb97f952c5f76f94ca5cff334a47e5276ff1dfff2f052a357d0e36a9ab48888a2b89625ef1a08f7
zc2a6ef4f1462dbb3a0eed8b6f8bb99418f5a8058395760ff69f591ddd98b335f648dd1a828360c
z46cad378bf56f84fce4be703a315b4ba7666cdf99e66e18b81643243f1006a6faf32342f49f3db
z4d2793155dc894dba266f0294984241d87f5f06767f85f76c8f1690bb164e246f371b7fee6fe6f
z6cbb70fc06f391fadb0cb88215dc7f864e5c78200730159fa69385465c65408163f2c5e4ccb621
z5cd55247910f69417ced24351e1c804f27e568f73a6c8a1b79a54df8b1ea3704d5829dba2a8de2
zfe98c2215cbaff1567fc3775e384376934c00f614c1217183f22126af710bc87bfd3a52fe9d824
z35d929c53c2cd8e2fea48df388a056158d519332ed47754b0eeb08ce99797e3af126f14836dc69
zf914a04d136b4135586ad54ad8e306524ff3d4b6415ed883b8204e68346aba2a44d5d43f02dc87
zfb0240808feb76f79c46b82e9f2a1862a686cc712aa6305e809cd18e1bf0246dad2805963b9fb3
z789c56c95d1bc0663b57ca90e26154105a67a617fc0e7caeec7b0c77944e34d2bf7c64b34edd9b
zd913f21f0baedcc77e7ceea3e09d13b62607c6593a8b3f7ce0a6e1873037a75456068bd7cd059d
z357811e6b2721e4c55413678e77ab62f2a47531b7233b2db94a86cef28e14bb634bae5e49b3d00
zec850ea3d552fa1db921e50bc5b2ff11c29afc5d1d1381619462042eb834af29940f98be4a770c
z86bedf7bc23834a4716515dc11355eb590d0c1c9f2a566c19f66598504717de6c4ba77ad700ade
za4a432bc3d6a6d4b31e853b0c0dc4a9f0c87e351ded8bf2cd00e84a4209cc449d2ad98df46fe7e
ze26ebd7556a68600068685435d794d40f9f28fdb345352cd6876803cef6fcdcfb5fef9445526a3
zba283eb6e2bf2d89b333659855bb5990c52b27d6eae502b9ddc68e250ae89a6670eed2870f672d
zb21f76cbf279cfa46eb5bbd4db2f6f221eae5385e89225e7381e03366f85d4ec376e99af500b19
z12ae77027fe1637f60ce815e568ed19c2b86f1fb175855762e24cca6003ae25da8186716de9a4f
z5bd966a4e0b894bc3b2a0edd71c92f81a9a32110a6a4225bf340374eba96fe470c54da7504aa13
z8c4b14aebdf2c58bdbae51c11332a136ab6f093769ab7ea121bd834d85ccc45ddb532e2695fef2
zc09093d43dfea520df40b027ad120c45d1dff6dd01bdf2350761c5c34aca760423c19c9fa03da5
z3de02c88d34a8ac41b57ccefbf66d1186bfa80e81c3300744c446217ba8ba6af9734027f1e52ea
z6a542abcbb77e01e194e664f5bc8c5e8fb8806ab4a439a3cbb12c5aa39de59e219702c519ec8d1
z71b912fcbfd3973853b4b2ee439daaf1b49cb50b8e932d2a5700c8dd819c782fd4da669f6a0fef
zd48a6e031ee372251bb851e067fe760c44442babb748a44199e76e86f640b29a7d4275cd61739b
z0da8d755e89ca28bdef270e8c130a61fb4e3b6c28aa09521fffc63247722a3dac48f75e31e8eac
z8ae0f3f7e605a7b783f63eb5cd6d068a52118a569a1aa9deb6562807829b453b30b4005519e8d3
zee46c420dda9ec010357e956a3b9bad76edfdc8b1dde1d6e7653e7ce9544823465df8ddf349788
z70aa5afbe40128fdb021b39c6e1b845ed806569f92f8014b5390b3eb2089be9545f425ddc7c34a
z16a80f84e3233ceefa341fc3228c746af64e7426d6637c4998a9b54e3a67d348bee677927027dc
z0b06a8211562acaa9f875b38dabe1dc33e1dd6343216fc086c0ea4437b86ed06057edd05b76b7c
zf053c6b8123ded0f3f0d4f4100fc00d8eefd17800695254e42f0dfee5b93aec28d97fe704b2de4
z397f4bec9b08a5c2a5ffb3c68647971b8be8875f9ffceab349d42eac2cf9780f4aad92a8d705a4
z270795f5e4407fd30f12c97a19aebf1b4501c500c65f369e01077803e6fdf7adcd0761a581e529
z484f242730edaaa55186f4f7a016d5321c26993abb820bbd80a1e69e2ed1c72b98e96f07e19fdd
zd20adad99fea104b2b7cb6a9445a2d7ae67aa960782348500918b38e1bd44117ccbe043442ce9a
z06f2de6562bc311727304237f64a557285f0185ec9a935bdcbd2ee50f841da703b70d978e2d78b
z46e288b148adc9c30635d3e66ed75c7ae4b0df3743134a0eca7ce0b874232698a13ae7d1b9861f
za3e38a6d7ecf3ecc7656f3840f367d7b63ef9f9470e7edc2baadc510caf302d1c2381cf62d98d0
z8d31544693d57eebb67128ce0c14b4bffc58ada87fae589963fd7a2bdffec836d3ee8a5ade393b
z9d7eb0db0e06f46ae523015c30d0a436f50d0a4685910f7144e687e38e7eaa20fe7ec8b3f84b88
zeee62fabcf34dc699b0deb4d81d9281fd3f34749f753b830916de4c0de582373b6ced52a67692e
z21125dbd3ec7c70d609e4bfb4d73bd6afeef2f921931ae6a5af46e7c5a9e7c22a5e9e8c2684fa9
zd06047dbebb8cd22e58b1665f3e0f096125286694e4f78f421602a91d863e3ca794bfb38430de8
z607353b2520304776dfb09acb5b7700c18642b7e458e6b9d9fa499b726d46b9e5817cee57bc8c0
z6cb144483bc3839f8beaa00f9a1156785aa1e5a2fff994feb1eb0b616b25f362d05b6338d6ef62
z48f2459632a8ac275a8e649cfef2f52bdb0ef0f2c8ccdb20af5a82da04718024e627475b29b622
zdd3686e968e19429cc47228aa7c659dca9da24db0dfd904f72a973ac37c6581042caaf1e42d2e2
zee3aa5cf973470fca361888c1f1929864695948c9daf3a8d85b6edb9e92fe3e135969af94fee4f
zaacabc145d3217c4d65d27198416ce20293b4c9f36694b463d7b3117a8adf653190f42f1e7d4b4
za2040a630f621501ca11034fcf712a2f44a82b6e3b976d614e44f0e24ac09d2c8b850fa28a8c68
za09f9862778005733fc1378254588ce158026cfebcbd4c5d235fdb40c7e1c469a51bba8bd2002f
z8773e1209d40cae2f55d4b1ae6e561be3b029e5d96c20850dce8cd51432769f40ab6a1df108d38
z88c3e8754e5ba2f0e472921bc740b50308783c11e4208fe6e79f0cb06cca06b61595f7abfa8550
z4c46e86c45160101a3b92b9d8e532a5946af2d36e4908b18912c2e093521ec17b8a9757233e9b3
zd6fa111f0dfc4d1234c393b42264f86e9080211b535f20ff18295f4795bf18942dc7b442af022e
z1ca6cb5c08d2df09aa1816b9397ea766dc7e1f97f8a101fef8d653ba380e4f007d48104877397b
z2069c9e0b78f1fe15652edd167b23ad087282e0ff6f7d03890b9476c40ffd312fe6f313f8e1ef3
z43a7b5330f6185e85a9bba000d06f426ce9254f3b33a786bc4798ff9de3c90b8d73fb1096cc6e2
z0e096c5c1ca5c29f34824e8d761ab15ac4556e8b8fe21a793b09ae5aac0888c8abdde4b6eb4d57
z04844dc695abae1e92afd81a7cc4b1dbe70fc0568fab04a7c845e542e4c4c426b6db4c428d0fdf
z64851dbfa52b1d6ab548b1cbd7cec68209fc9a979e17faa4c697ea2d0c4c08c804467b808b8486
z388a275bcd64f8849d33e1a5c3e82dc769dcb7ffcaa4fedfbff09fb38b92982c261574db9f391a
z5915bbff548bb76dd57dd26cfe632f1e31d7ffdf9a61b24c5a84eaee77609c316f56ba639b1f25
zfa0b2d1662f3e251e10eea35c405c5ad43bec86c040195bfa41884887ec7bc924212d20d0932d8
z98ce85fcf37c29457ece1d7e9b10c6216387af758dfa2260a60f8997fd096c29f249ffb6d031f8
z29779b99d4911065dd1ff7316c33909470581cf00b9de7fbcde92277d63561cf658b81383bb47c
z0ad657d68d0da6be7b574d12f2c33638c8d8ed8e325cd0465ededa647b2324ddc87e8d28bbd753
zc2700b31c2f05d4dbb90194ed90bc681722bb032868382adacd143afec1cbaa8aec76d41d2d0d2
z8b289b9f37bef4b26600209198948f71fac78a2a5b3e4c4ea448c3f186bbd20208ba4b74f17a63
zda4d9c417e0d11cadd53af955d3faf819eb305f5986b37faa4a77f6737ced5f960b4a88c1f342d
z303fb8c42d6c6842fabe6a5652085ade8c0f23bb71fbe4b14c4f521099cc68c925621ea951e735
z7133ec86ac1d8545a75540b1d7c6c6fcbd47bd0a315d28f487d8d26404f4cab2d74037128cc608
zbf20d37f8ea10ab7a02be3c3f9122370649b7ead417a4831753bbfdf092b2d2fd59836799a76ab
z7f6181f4b3e432e15b441b2ed14563fea41500ee53d605cbaf902f6616c4d54d120b1ad71c65a8
z3825eccf0958690cf116297e9b940ef71afb3cc1c37ac14165d5e742f1083306ca9c58607cf48e
zc190d5a26475750c208c8cd243accc376e1172bcdf4185b162b9b7ac9a1b4cabb356f0eb29a72e
z35156109af2903535896d6abfb6dd4b12ff5b6371b667bb2311712fe5c217d6889025d9f2b7a87
z8fca81956b3506ce73f7a17ee4e8b9090b76be8ce485acf2c828282af5e41609874bb6f90df9bf
z0d17d40ae331b6a8e8959c28a62519262383d28520c38f5ec234945b96318bc67bc50a80cd4dde
z86b137ab507a797d0d65a1cef520ba60cac934e1a79632a1b0e3b39169bb79dc129a0dd9c44cb9
z2027358c8d6010987934c77461a475f9f30ec5c9b14633032da2df6de467afb1f37619c71360a3
z46a08773c7aca71947d434173661debca45a9e8b6e66750005d4dc631715aa885751d020f568ff
za2ee38f2d0e9460ea54aa72d6b348a506885a66a7029b9eda538d24c4d78a513a7c95595fab93a
ze4e70c772e9dc0292d401bda36fff7f2e7e4d85e319692defd9f8a87a0a29ff1964bb9e8eb7dab
zecc5a4b5383c49a690be58c5ee640aeff32be3cf7f140c5c954424c87a7d0dfb3f4262ad5045bb
zeaf39d85d2f79bf1d9d5be7bf19ae0e5970f7625a1d64da155fb02a2dd5d07c316824cbcd67f5a
z322dd957b07988b662c9a990002750c891f979c1ad20c7655e64e7cedc90cefd89ca13c44f86d4
z905a5da1876cf33f0616bb699fab8e34d66ac390b5ceb3c3144086554182c97293d41bb51d1b2c
zf6cf559d56bdd5cdb9ab45b92913d48906db1831aa535e55b4989e8f212c4fa9f505f677cf079e
z98cc2e8a7d49d970ae4ac275061125d9c3179f239bab4ae9ff8605dc7526403c719a4452cd2323
z89aa06ba9af3e52b02f3bda5a5b09107fa5133dac4213834f73d2a3e191acc9d94d10988df1760
z0c1ff056a8bb1f8655000191f7005398f33d7b89e81482200b1874d40457def37a41c4d83dcfdf
zf75de499598d5ced39ee1c13460066064d2bf5ce488b6bcba67c7711bf6bf7c08262bcc10e44ee
z8e5d068f9a407881152ecdc5d74d5f0fbc676ac0937c273cce4f76b1162f2a9f402fce25e91c4a
z8bdd15ab6d2ad5bf4ba6cb42b73d09ef0b4cd6af2bf2db963b80425373f25321eeb4cccd3ddc01
zee8b71e6cf69f94f96ff23838622f77f54e6b234889bc3ea9d09bbe5a2d6875fbe29f87238e18b
z6323a4d10cbcca0c72710a852fdf4b5f998448299d4f93fbb6aab3653ee0aaf3ee369f242e021c
z61317e1301467333a1bfbfb2af9d2493e920e8c3bd4bf2305e930ac7f2bd6f67dfbf40a2a4ad8b
z53e7e3d77ad47de75c11f7615e110e05cf5b6bca598690d4dacba0ff6ffaee9a659abdeafed8cd
z1fed0b022d8481d08e466e8da72df2bdd0dde00a5468c49cef50eb9e69d429bb5d128ef4d80076
z6d3ff06aecf04dd5da9974e15346e7591cbfb9dfb4f562081c301db6983eb918fd4f3823b35fb5
z0d9c9adb73960754439018f3ba05d7107b8860039f704c23d1f51392f034cd44a494b62b3e1f84
z738b92647879b3fc7ca4ce477897741f4e75154ec505d7224b0a6aa3896eaadc9faac2955fc93b
z5f890bad54c84ec2c3a3b3110755d117c1fec38a4049948bfed6e7a086cfd339220f6b3edd7bf1
z4dda5633cefa1b7e030b69a33f094ee842d289a20f3db737bece2787ad32029c2b73807fcf69db
z80f035712a0d0a6e22c113a5c5c7e5ecde6b1374d760330d065edd1eb6ab03ee13a709fe595461
z5b8f04f77e3468c0bf803e050a23ba8484824f6903acbbc39c2ba1cee792abc0d4cf48e20e657a
zc21618743c27a703d3b935866713ba683343064f4026471f4e639be885afefbf1514bc28f1aeee
z2c52674054409abf96e0ae55a255d10a5691bf29462f9dbe85409b872efdef998901d7ba85af18
z3a8c93ed7d0519b1878e561e152e98369c039219f75c22e2d634810e8f5c1f0f516de516f31898
z6634445b75b7d49d1cef2d9f566c4d994e9d440447bc2924f88f070ece80b21b16329f1b7df9c1
zd4f05152d1449b845dc080755a67e3bd6c5857143a9ee08f93357fb8abb1f832f9216ddb54cfa5
zfc6b5bbf0c013147387ccbf3160e077c6e225241fefe5a149dc7e9a909c0645f30ebbc53b8b67c
zd09c9647fad22493faa033c820baacb20d9b28ae583f73a5fa46b0dbbbc97eb1a5ed38debd9ab1
ze325a8d3adcdbd96965f7e96f044585ef889906a8e2b3f817f7d93574bb6c8fcb31ef5b0cce84f
z563d55c59b0a6fed974d21d6882dec23ef78bc954c9a039ee85fa230c2dd53ea6dbf63352e0231
z60b7608c81337a29bb92d2ae737ef68edb002c5984df9040aba07d2b7156ff221a5049f71e618d
zdb15362188c10688d01f7eb24c4eaa267036fbbf2203fc9b70b96a4446c54dc3e1b4e935b825c2
za153569dd49c648212ece86d252dc7ed12d21b32ad0b1dd1d6da2306828433b9751cce1739be4a
zae09a81502bf00fdf3c416b1b7375e833a98213e7fc9352a9e25bb8ccf2fc8a5a9116ffe252ed7
z1f2178f22b9723b5de6964c8ffbd51609b990e81cb2be3cb2c70a8fc8e2ebdd36cf883a35fbe53
z62f62086461c33f39904b8aee048e685176cf8507b79da7105e6333722a1bd5c9c7ac5a5dd9cfd
z80db252031c12578e8d661b5858d71dd35b2e898dc7a744e73ff159d97025da51cfd85e3d33dd1
z9df3c4fff4df7130a03e8a9ff413b616e3c1ea748e62b4f4aaee8b1d2bb957cb26a6fc65978651
z80c36ef6f7e780a07024a8decbd2507d978e1b28e7b78e79cd62a15a467c068af55b66640b6fe2
zfa917d4d398eda3869281d6a9e06a139aefd18a4f56294efa0a401457972902979834a5e53dbf4
ze9e34a3bbd7519cd5297f1a369a6b14cbd9adb19c339668800084c879b0548301858a41876c1ee
z384c5a62ce486df4854311bd5e3d14d5e61bd5971153103f5a095f0ff46837d90efb813d087102
z2ef2121552282897b8677b558c91621506f5a383938c1e25d8d3c72f96986b6e11cd2d7c4c9c54
z20bca90d3309357c01a99f0ec952361e55faca6da6c991b99aede09c94086744aeb95bf505a73a
z83b66029ff6633cd5a88130eeb9802cb8ac9a556b1cf4a2f4445aab94ba4ed836f77ad7bbc81e5
z39f3b61e27c15b73b79f8c2ce34b79724e245c9838212b4df6216b0617d5bfebcfab4247955571
z0abb1b3a553ef3382b6018910d337f9deee875e89fa6b48c06129606176ec703d63126fe522d32
ze65c4ed60f3cc07f959f469096ab79d69e97e692dbec451c564c980764297079c09dd982f43b8a
z922ad94226d7fc5bf964a83faf9f7c10c226204cd85cb19afb1a0cadf2765bda891cfc8494833a
z4cbedb68c90d1400a981b7664118214ac7bbf0a91316ae0a64e0da697c5f1b38e40fe67896cd37
za26a72bdfe4eb693c74c815baf69aac920be6df458bb293401d37b2061b81adde7d193f117dc4f
z78531023672becd426fb6475979200bfce14b92e2448d8dc9a34a89774928fe4ad77774962ac8a
z82fdaadac8f195fbae1332bddf519176a3882cd6c1e2dbab5b475fc5ac7ebdd78afe0cd4904e75
z504d96428500460caf4b451706d4af6abe5ac93848265062f68b532906f7a66afea279dd171983
z7632bdb012d02b8ccb6639be62e9bcefd676a373d366535d33f0b4d8d01514d9b4d9166db0508a
zfa3499482dbd81b07bfb60c736add13f1b315da3ee8b9662b9c2d89336b035a649f4e6af06a998
z7f9cec77129780df4cbc4b63fd444041bc2d574c1725401983c0ea22081cd4aeaf2ade912352c4
z737adfee1c02f9759685230073c7db33ca5c457f1fcd5acdff73c40369757e7c02063892dd1ad0
zd592fdc290bd2fbcf388733e733cf24b6b6996e8e7a0a4e900fe4b3029849743e8d2ec6a75b6d6
z4df4a27c35b81af4bba67715acabb4509a0540e349467b603f439ccc23dfe2b3819c396601101c
z7ee031bfb495008e757983d2a54ffd6d7735e0c684e0be0ea50e262905d283e30ca37408ebbf93
z8f7ffe9673901fc57c2c95d74e9e1099a55e87fb4c06232f7663892cad2a925313738bb5fe03a5
z4108a8abd75f1097b0c31a374d32a01c20db4410fa8beddfaa63ae893165b558b45d143c09a42f
z6d3f2f818effc5ef45425da76c3eae6d0c6a539f47f7e1f85b6d921a97cd372b3017aa846a1edc
z919431208e5751322cb42ff48f7fcc77f702136dddfe8b17075693ad5c57d1ce9cbbe50a80cc19
z1e633b875afee7e2396c3e9884253fd7ef23211ea0e0d0c9ad4d6c339f1899f67413a495c5862b
zcc821eead38682ca8d290460f9c4717cc0ba775e2b11226029784155fae114b03f85573aadbff1
z5459f671eab9d40e8bc8680e8d3bb2d31f0a7ee819f4be752e1178a5b922ee578b77056bef9cd4
zc37b1b854ce15bd943fc01f42f18cab312bfbd9b311b0e6e39fc4b6f61d14de9efbd3af2838311
z7f846c61a112856af7776a078548218e845ace2a6223734e61dfe32bda1aa2ac27973b74028714
zd8155834c5ea7ae529bc1093f37892f575ee55e43cb7925a7c986b30e6b149aa4364761025f195
zadd33ea032637e3c32b8fc4a897af0df8b0ef8cec8241f718e24b585de378a9f63fa28552b42a6
z427f87063b63b37ba4ac17c9f47ccfe4e7285a4e63024873fc77e653b410f880599b6cb469a6a0
z55e241b5ce5a61e43e72617f6c31ecff6da18d682ab223cd7705ebe1ac311edc127f896416fc43
zcbd6afdf00a8b61624aa5d35720028d8b5463f1633d9bdfeec30c63880e68cc0d3d0269bd02e87
z85e6367692eecbd4ae1730a22f17e9f2a1b2787cc90c56df3bebfe6e771e99da75d505d178c4ba
z2ac30ea3d2e8eb7c1bf2c02ea37fdbc2ef3f7f88a4e30908f948a2e94fc2248142f6c18094389d
z5634b4a6bc3ba1f9d4aeb3be3cf406f15a8aca24395925fc8a9dd7574b49a123eb3862e588897c
zaa70b07faaee8cfb3e67dc189ee303529b1f8d5a5b91c73486ce494d499681c4bd5482f35f9548
zfeb9595f22c2ea5b6d36b21aa33a0501102aae9ed39e634a5591579e2c491f3b7aac405cefbf9a
zfa36967da684e53fa3adea909890c1b827ba26efd933f2ac30daaced6d62664194dfc479764a61
z3576c384260f069d86d74a2195e2baa49c0fbf16744ea9b81600e601c172221eeffc44ef73bcd9
zb63c81b422d225beb3962d3e02f7a1bc906a7ca3edd4b8b3777b316ad15f093cb7bd295040a37f
z0a9df50cf080a42cc28333828c4a5bc68c1a07d9f28052322dcdd6d41395c0c419ef3b77604cd8
z9dda5368accfc901963276ef36924087db4a00d0189cde82218a168b06e4ebd98af5eeefc00f18
zbc5fb471490e4404f71e6ccf4bf9de9b197aafffdac745f07ec527c14227ff0b3da49566031647
z0f7f8c3052a7047bf52ce817c1644b3768f1cf47d28860baa307245ba6fbe6eba20cfc0ef265ed
z6561e0c1fa4e2a77cc3e74da72ca081d8de0099af9eab43463a0110f9bf13d9cc4290f0eb5eb51
z0b86a78491df4c661f7ee59a307c658df2613fce4b42cbc11622a6439d9be029cdf42fde6947a6
zd86b464232e58f6f6df610ee4be1470ae6d095fd4edddaa05cf48478def27f1e15566bcaf9d44e
z30ca109e358326fe98575f3975fa11f615463347a8f1c019f036560b3205dbc5e76c780c56c2d1
ze6b08a6588da82b77499b5fce0cf35c38775353fa5d47fa333aa5880e5f0279333b869b09bbb8d
ze11c84626c00d7e187883315da9d722bb67cb7c7bcd1185bedade06091607b6fb4dfc1f8061dd2
z81590723f2cd65a4e024a173c139ee27b91468277f8395e785448db226185b7ba76437acf4c4a5
zb593b00f660bdf09e43a76bc91bc1b3556a1812f871a15faf43e9a98ef8237f5c02d961073c9d2
ze5fd4dd537c6710435c906e09673c03108331ebf42b4a3a693e108bbc7019e9653776cfa16ecb3
zf09286fe1a2373d4a9244f67327ac6e2b8284ac0617a956b1c460a11d960ab15224d97605ab805
zf1db0412bd560ecba3411331042c76f3f1e98ac9dec14e8a503de1bd34680c83de3f2cda541da2
z8393886f222dce3a1b66916a544e36c149a2a42a52cf54ac457d07fb2321d3dceedad091274adf
z0b070a53b9fd6b4e8896bd076bf936b3944f7e4e357e7fd26024325b424df97a8a1c2815e6c4b3
z7258ad63a1b829ba2a88e6ca6696c304552fc28303633d3122f167b4e50ba4d92b2937b5246c82
zc137113acd6a1162a03bfb14fb40d28698f3e782cd8f81b35822d6d860504aca3a6c705c69305e
z634a6979d53ebdd5583f6e959ec544b7fb6d15e444d66cf0b8a0d6a82127286fe6696fe576c432
zb078f3dcb606b4d5c51901af92f102966334d5d46f9f66bc7972a07e0313174477a38c968d7261
z0046526076ee58f8382763b0b19b8b023f02c60da87a3375575ae0bc93065e60c1d4f76693d13a
zedae711163b98aa4131e3aca53d57cd26bb00cc3e986be60effc7e4fc4f342e8571a22dca1505f
z8ad4a48d42d6db95abba24981d7d4a2d38f0eb970c633e0f41ccfa166f4cde48211537938a2e3c
ze9aea0d4e7bb2da2c1aa83db9fc837ff1377f64b24e881e50c69ce085e8a4273f152694971b08c
z59e637ecdac93c3d4eaccf10befacc8cac1d2a63e72193b6fb55cafa02010836415efa2f06e203
z45101cd96ee3dc4cc8d7c3d77c4a4cbea65ce19490980cacac653f06c6598f7d0c0271b100c8c3
z2c03a91d00d5baaa278f7553f2be0e74467923eb9ccf27e0ca788135fb7c6565181cbd02a0b7ee
z43b718803594167dec62a483178c1c888e30169872e7cc2522130348670c4ec6b1678055fba1ef
za9d9305956f0aad738cacd9023e1e9642fbacde652c6915012e874c3f6616039117a287bc04d69
zb387ac1a2cfd5b5627e34876e30bb0fc0cd2863f1208fe673f204d0c5c297f78ba074872cb67c9
zfa1e0bb625d9af1fa831f70676f3fc71c89d03d3f54f879784fba1a7e2c3e1
`end_protected_0in
`else
`ifdef MODEL_TECH
`include "qvl_multi_enq_deq_fifo_assertions.mti.svp"
`endif // MODEL_TECH
`endif // encrypted_0in
