`ifdef encrypted_0in
`protected_0in
ze74c34e226135848fe16db9ffd31815111b6d7fb642c521a3f628cf6da949865580b22efd062a7
ze90adae0e65e66a2c36a587d0a790699161455169ed55a01f2084f11770a774ec4c588039b380f
z6de9c5084882a40b79a175f5c2114b2b6d78b070cb806e1c0aa9258297f4687ab308bc470f0040
zb0b1de382961eeeaf2e279e1462520fc31c119af8f2b214846f56c2b3cd2eadbe4099496abff18
z15cec83ec4a77b868344aa20ba7360908f5c0de2a79abf8b3534b883bb12180f68b5d4beb444cf
z3fba8f13afb0abfe8fcc4294810f75afe452434d2d0f1166236c82f76edf1e12979f04bc35693e
z32ae028996dd85737a8f5adc1ebb94f39c940246e887647b64782cd7ab429b0544c173176cede7
z01dfb26b1f73408344a52b7e1f117f12bb9c8077b34876c2e6fdc085981637012dc9754765e1a9
zc512ce062e0b8fb16a214591f5c81e1353b900a611fe1f4886b57940b41b7f2ce99a7b84b04b90
z916f717e73bd10589c81e207ed77ec660a8cbed5b487fa50acde1b055c8870bd8676023f21ddcf
z9c98cc47cfa2d654ff1365d1f45035a045a66c5dfa8279050262529d2cac9e64fd27d9c7de62a7
z731bc808811ded9016570962244887f98fe5440167bd0088f2f049df882af501358497c3b28776
zcdc5426c7f52a851c35106bb93e16fff984784050fc808fad15da330f6f0607eda2d0e0e4b1215
z2ac5b11453f6b6c5c6b428261a64553d70b4ab9f1bc235c2ceff4f6e3b1ebe72fceb7af9adc96a
z694b4bad7241bfbe775016041d7caaa74d9c0e7b507ce89e8b01980415bfa35a8e346f54c548f9
zda8767c02ea87d27eb7a843f4cada7dc3b575fb5cede69da7a4701b2d725c73f1f7375e85a74e2
zdeae70c30f1127407402c955b283d7b9512dbb3cc85aff97f613d57a4efe57b3c092e5ccc5b6dc
zd04e277cea6810165bcacbe3f515b3d75051fbe8fa4af7e932d60d2b2a6cbc14783b996db7f97f
z0df4e054ec07012afe312c7c27fe5855e396fca2df20ec96282aa187aefef584e73225c3183714
z599297effba6810dbfe57acb29d5b025ac9a8ebc73f537d2977dc34b086017b79e71d435e90724
z58f8859c47b62c6b1fbee0ff19f88a66a8afa79b5c1920e87193650fc0cd3c6ab3d109eeec50bb
z55eb338914c7df8dad730fbec8e96d273894b815cddec84939381f647d6e3c4942eb7717872703
ze3f888408f4574b947406de74946046ade8314cbad547dada94ace0bf4ac13fb61e3f49bdac0d3
z4139ed71f83aeb75542b9c25ec57e9bfcb129ab35b8abcaa9a5cdafa5c33bccee73fc848104b0f
z751258809dae3de24d9a37858aaae417364b48e3cf9b58e5ffdf5a6b87f0e91dc867329bc68adc
z8ab348fa60cf03b1b0ad9f98b49770ca5e1581fc4db7d9507a27a49b8e909977d410ed44426c48
zcb42a72638c6df8505974a645ff2c8aba5542814be671de61b72334740fee00dab98e5242cea2c
z8f449709095ee26df77d7d833585b3998b1920d091a35cb4a0578c689ea38defe72dd2a036980d
zc0ae6d7c2bee1a8f68bbbbb00727803e1029f998700cc5f688c904bb946ea03e44239d94d84ecf
z251d67d12697411bca928da0a7f52b9c7834462780c469638836aba7e941a0ee7ad6acb3332f40
z525acb0f220959c7ca8a10e3d9a31cbdecfdd21991804b7be7df37ef272713c54e6e4e666eb349
z02f8eff176aa8b7282117ac5cf8a79c925948ec3944a539722a73445d54d14c1450f3352aa917e
z8c65e670a8d5020f5d9ec59a4f08a2fac14d62ccbb7d8da6d30963f13d020b4a6fa7e0934b8d09
z967199dd58560dc80ac6f0e1bcee7497202e99cd8b7a204801c4239574352abe5f588ad6cfb518
za7d248b7afdb43bc1062ee7c9451474d8cf7a0e32de2f4b03d9d67234715d1a0b4911dbf49b988
z4b20e32a4e1f1ea93d2ad700d41be85d79ba979280803c24b355606e8c0930d3078085813bc9ed
z3daae4ea956f4874a5563160ead3c34ff8023754ddb295eb3a9918686925ce455a555a32b47bd8
zaa5856a65989323ef1d7b6dfd7438bde6f87f8c536d386aebd052e7c4b36a21fbaa5435ac1e02f
z629eb3bca1d43616d1c1226ee58063166e000b0572dc97f94bbbd3245aa1b5c310eb11ad1f1565
zb55377b17eafeab0a38dd10ae3039aa0b8a66888ac8a2c16b4c64a965cdf19bbfd5d79d45fbb97
z08f8ed6b63b200507c32c77389b44f7592590dbfabc4243dba5f8e13af9710bec839f42e885f44
z2333c13ffa8e50c16a81a200fdb1b90f5085b2d74add5d0951801c0c88445030ebe68b1da1c3bd
zf1e6d12fab0df881c941ee5b31f5c68b81df8a8d336fd0a558f003483dfd467cf022d671b2625f
z055265bebd1d89a995d71c859b11500eac1415385238d2c1a930736ddaa21e097e100f3670fee8
z68411b4de0f4eb1de8eb277e886bfe0f6bbb683bd286cabc7da047ec9622319521767fc44657eb
z8a2194a3173677f946e003e8610279a1893a5bd035e8f74eee820515e4231ea51eda2f1a8378c1
z6c6ccce49d20caafe1b7c0c2608d9cc73ac5dd7732a722493562d5177a5d37cdefadd0ea87e955
z6a14d99bf65dc9acb33787c2015f5e4f6bbd3613a2fa7aeace44627a7f4e9847de3a85bff493a7
z32d09ec5d4c4dd4a9eaf83ff5118db9d381a8cf1bfb3bc4dceee7e51667c4b942e7df5f5110333
z4fb3efeae784c71bc8a303b5c5ec0424adc95053c5ec294af41a038fdb866d994d841e82230e4a
z309d46d978533ff09049899521ca599a8a786b7cbdb0110edb13a23a9611962af8157fd05da22c
z7b58e681f911d957d03d036c53286bea30133e6858f157a23cec4581afc2de121dbf0fd1fc09d9
zec21816488222da7cf4cae5af0041b7f266d8283c0edb50c4402650feac2c21818d36f804a4e15
z4c19c48e202810c9cc2365858ac636ed5c9b7c22e077cd7e8b5a5bc7cc2147b96f3c8246b4423c
z50a5bb3986393c1e264bc3ea70d2804c4c961aa7c3c21c93e1528bca418294d9d7cc588a9f14de
z7f381b438161d7038eb41f0a58eba0a0e21aec04adfc82f3ed9fabca1e903a9289711a8dbc877c
z07638786371dbc8bcad4e1ff117a4ee28473c6f7fa65440ce514c641c5c54212bff8ced3c11681
z4f8df60239e42d6c1046299327dde54a054ac790c4da27ed5f9299a27c8a61854fa7bdeed17f8b
z34499f6f49866bc317917b36b6af1577ca2d4c439a4fd7acb3596f627edda3f009fb0033984ac3
z450a2921d9f72410da425a51f5da8b2798f18945e6102bdb24d7f7866267f02215817e450802e4
z814e49f37580f8a554f9b569bfb1dbe61fe7fc8f2b67aecd932e66ac8abc392c4f1705c50bd63b
zdf4984d07be3ca179442c21dc7ad97c94acf8810e4c41dbe3da65c4715a092800e0ff8c748d8af
zf2e27c85e61d3043ec98df784d8e9e95df03d0c037794f93dd05b70ffdfb108586a4ea41268498
ze0902d9bb0f58653cc6164878a75bea51f8e3261f61511455331311ed0e12e2e84f5361a1ecdc7
z7e0ec15270e30e16ae6670012ed06a402bd4fc40043d6b0c123da35737df9a847f171fd54c50b4
zad29b0c34fd0be35fdd17dacb94b7f07c11caad1ddffac2e4c520b6cf53b6c9b670b99fa6ee149
z8bcc445d0397b71d9447d09fdd44df5802daba062b3e6d766ed9926e41c0cdb097003b3bc7f640
ze3f41f0a698dfbf3ff7a06e8a0964ab0436f238ceec9d7781d5c56ae4c89965171ab08c171f196
z0e44ceff13a89cfc3a11db0a033204691129412b91e1abecb31328840ce068cb686a53f73c1902
z4fcc38f76b63efda80308bddc3e00e4f8d0d7db53c4bc098bd1bf2e20dd80a3b5d959a07deb6ae
z1b45728b11074976241af18b7526961ab1683a08b7edf4d72cef0a16d6a30448ce609b0a3671e5
z2af623450b1eb965e93a94ebb3987734bd464f42c7a50049a0a48df9fa94c4138f977c55fe7089
ze23af3448e6c8c294cb399eefbce041ad3899b050e8931e8cd74105c6d5c01ffe5f95385de4e08
z85d80d2a3ed346756924983865b9fd85bd945a8f314416da8f080d43962669ac6a036fa77f95ab
z56a13df276c68519532ed1f00dcdee3bb5792352bc4ca270b3e73c3877a792bc57ed077a55e8e2
z88e91f102ddd0db0cd2132870d036d90c448a4814acd5994c856e9468bf3e9c8affe2e9d5ae9a0
z9e979a3a206b75be093b0971e1f2c57267d3eef8c15f46e255b518ab43c8e0364eba1371c93188
z6e0f84971e4f7a4d9d64418c2b63103f1e0a49fbf544f7f6ef9ec2fcc81b8d3ae07e9b36f91b25
zbc79ad3593817aa2e470a8af515e405662178d625027c4a4a4af2a22f454e94793bf4caad19e41
ze5100fb7efd054d2578e6fe21056ccbdcf49b952ecd5ad5f57add798cc8ae7d2a2d6b608fc91d2
z0554d7c28f59fb6e6ca88f29189c12afa13be488f562db51673807367ae680cd38d3a5ef9e07c4
zbd24d06e773fc2d4bda6cc8fdaf61a13d0088a5756e69a52b7104557d92466c89694dd72e1b380
z99ffa2727882e3e62e5cb48d4428a7d6e3ccf00eb2c0f82749b75e7ece99856efb96ee4b52f17a
z4525e79f5b5a222412c2335a7a00a7b27c6351da198b588bb64ceb887db8fa2b5300d0477c0c45
zffda80fcac6c7fb32a13d9f7cad3b76e4376e9619ce3ac0f3d7e7adc731cd217c2b0bc28fa649c
z7c9078e1e1f51146ee0e178c03bf2164127d2d6dcf991a813ee8993289d1e82db8b3cea0e862ae
zbb6bdd6aa50024755acf5c13b3f9ce6d49220071f8be6bb992310052ba369d7bbf3d866a4f48c3
z809084297d66cf3e1df6fe178b5363d6797bfb0883036acb8df585a51515be4270e44c79f86992
z4e5ae73313f689c3b1c5b15edd2ea2cceb939c6c6b30ab2b35f851ed6d20306bd757f3d544f8be
z4cdff789cf20b0078d421368c64b8631f25b2baa459cdd06421269e434d7d1eac6a82ab2ecdd16
z3e94d57ce5dfd7c043176ecd75ec7a21bf0f8371c932fdcacdcefed7d0fee1bc6997f1df2183df
z1cac556db7e150df86901733480d2355657e83cd0eaa1a513f75e5b5ce24e7733754c05289da62
zdad13d4dbae4e96df218a50319b410df7c7a8a64bb4c3b610d021c6380a6a0248e4a986b4c61d1
z567fb1adfd9c881d1d41b6bdd21d64fb68c7777ea1c09d904206969a9094dd5b8456b76270d6bf
z8ccc8dfb9d165872ef773a7b7056f5da082a359599d0fc8239b0788897c4b1757efbe27793335e
z9cc660aca83f82768ecf60e24c6338a182cc6125157d51688631beafaf982d917feb107c0aac61
z8934fc9f28449344c36bafb645415de3dc7f384867917e75fb2f7a440497f238ecd2b72d9a1cbd
zdeec9c3d21b6d29832fb37d25b987e91fd0ccd6dba1db3ee9b542fcff445ff7b742039eccdb2b3
zf756b398bc24f1074d93c6d32478e784cbe70952060f9d5fccd5f5e5eae5d2866bb4a0d5508ad6
z89de281d65570fb7e72368d3adda88a061e15dde5a6c9e745af0dcbd6761ae560a74452d9b5b30
ze5242da8be3532a03c0ee8dc048572f266fc276e9a0e2658d61dfb0fe8e803cb264799a530f913
zfc6786e86ae74b1b823a29f8ccac1233b380b21fcc85315a100739c9f2e15e0c81ad3c1fa7709c
z384ca07354c861858dbc9e228f4287848f40fcdb6fca6faa538bcd61850c6eb85af5fdb1494ef9
z9e5a3ffb73076f3251ea11af6ec991d6bb8b324e0853c7ad1be6c2cd7959de8e2e360d232b8b86
z4c7ea26ec0bf92c3b685f3f820673b38737dae592f6cb02e4bb72040a97b4ede429703b1e48d75
zf7fa94346c863229143207bcb7e565687636ca736f77deef6e3b6195af1f55c4582f00e8cc8541
z583f5221a1310ecdb8073a06d5b5add1ddae8a05c6279d64749959267ddf2eead2e42e43f9b3c8
z8489a91d155e04bb39bcefd388aedecfdd23383f3423fd19cea02583b4effc6dccd755fe0187bd
z65c2fa1431641dc876f6004b2adf968de877d0d231de901b61aafaf02a3d9063c3025761730b46
z8a96beb4a1434c22023368b9539946a5348ea013992a41607a74904ff1f80b48dc73777c8ef637
z6eaa679dcafc8d42f77b7e5a3677de04d108938ee912357bf1d9b800cce52d6cbb66314d56722d
zb53b50f03440c0b04462d24064e5b110f99f6cab877acd8482eaf5f448178a1f3e0b2a807cda2b
za1d21f378ec30ca00bb744be3e19e83b493900ca824a7894696b00c74dd9bd7b401e0dfcf5d731
za1b470cb5a7112074da1dbda2c685f1fea9797f21e65e0a54161897886b1194a030e92db920481
zcb13cd5aa2fd2a68a498e50d588b0d3b65e4f096eba43646ad70c5ee19ec8ec2906ba05f9ac799
zf68e7ce393dd8fbb287511bd961f279475d2c7f33ec599611886c8681c89d1245a542138001ced
z39409ac92cc62edc08527aa1ac1d55c31e2aae8578ad6fc26cf597aa2e217e53b11fa6ef8bf578
za1a8f71e74b9cfd45aa91f17e0317d0dd82cf0f945afd2e4acc7b1cea9e556ac3f83521e2487db
z917c014900d110744953f4a05bf1751b19c6e2a22dd9e84ec45bfae5513100c1164c9980106bc8
zd51716ea57e8bcaef1d0b842f6d63d4c0b66e64ff61eb81e2095633c42425a35e5646b547f9674
z3a380ae09f8d8e327dd38cad777941017a556cd377a3adb310176a25c3bcb7e88dbea6075cff29
ze1eabca027ad2336c055297c8e9111bcc75955ce4487ec1e14f5a77266902668e0c953607e5609
z769bc5161d48badd519aae0684d84d8770cf65226dc2c91a0bcba5d3a3238caaeab6b7e71083c2
z0a9ffef5152f587b991f0a48fd5954c7ccd4058ef5ee9dd1926577eb483058f848852de1b97719
z0e8278b996ebf339c797d2f24c47b354c85f1c1dfe3944102b12fd03ae5cb5efe243b4087fa269
ze280ca77314ae83c44ed124a2f5e7f3e6f18056a6348d0c90fefe2229d76fb86ad468be4a1a03f
zf8b7758420a7c8395a85ce3fe6763d20445c4fdf5c6598920c0ecb6afec065b06cceba12a7bf1c
zcd8cbac6569b11d92e370fc48148bfcf46126ca845eb002fb857e17b37a8062661c6f52a714772
zd11dc116c199d29fa6cfc6dbb2d928fab9a7d0aa4699649a5725616d62a55f8ea4f5736d0ee8df
zfaa92ceff894353f505e2e5fafe3a96abebf9db0b5fbacc62c1c28f6e98cfb0567ee85da5bb315
z88b26a08d23dfe5f8099377c5969eff29cae99a1f452f8b292d14c66a1eb593cb85092db3631ec
z9766f3ed3142d5f9322e66282a8d24e7e93ac10106a38f566289d94116aa4818596bd0377ffee2
ze4bba122e551b10bd56ab387f81900ae36660740b12351d7fcba421c9bc4248233fcdfbd9c94f3
z8340c0a9b4a53577e3d90ffe1b78fb78cac62fe4ba6ec9405562f49f5bfae2eb4e70aefca1d80e
ze91004a47850ad54943d48ae4bdcc7df4521c0e51185a8cfaf94bb2537bcfea8ebd93d9221979d
z19cc2c1d44a8d0d3d1cecae081acfbd152f42a160b194b003793bd7b33db30dbb830e9eaa40c78
z85be046b412283c704a8196b0ad308ccc528b4dcd7890ce6a50c8a112fcfb31d101ff166df408d
zbfb9d0d4fceaba17c5c6a8d9e3ee21e3840969845479831ed57f1ca61ba03f8b792fc0646f02b6
z423a4544eb2f724116d6c9aafd7ef015477c69b60d60f919e52cb4ab56083027c5b4c004f58acb
z0c3e7d365674ae7a21ee1bb44e1d968ffd8ef3ed63139005df002e3e2ee0a48fc5e7b20f546d84
z32b39bd406ca6c442574a931814e4caa40b0a3361f11ca47282631f7560b9f43797f1d5a2638ed
z19484c9d9e29d59bf1efc462bdccc9cd8f9e5e9da2b568ef6bbea6eebbbe72e5d9b1f44256df9a
zd81c00031a50361037796099e1ed0c0e312e95f711566bd680d5750f4e51d5808e285c05715a6c
ze7ee74e1fc1ef3277bbaac9571a68867ba93e5dd07c25d37a304194b95e9086ed6d2528968d114
zb46c0cf806ebd809cc8d065ba66c4266d90bac93a7c37243cc0a93029870d6aea7d046dd0c9ee3
z06d56730f15c9af6dec867c9728e35bf72b1d32af7787f17df3b39f153e7a7b3e440ac310c60d6
z54f03066a68f5e653a9dbb29df64933ada27c8a3357a5555d419d3c4fd29b813ff4b5851733488
z3621145889a8e8f165968e5a39b9a164ffb8bac64fc2d94fe72c575d64ab4773185e9af553af97
z917640e06c0efb0a5f834569b18f5ba46b01cbd9cdb1af6bb6b1eef759f473dca3b9201bed979f
zb814bdb06c9881cff359c0e13c6200ad1a50a34d81ea65156e640c13b778e253e3441a842764ce
z747cf57b3af6d0789f5f877804b38bf762b15d5ec65e3a9f827e223ed6d18f5fae7032673f69b8
zed7e29fcf22c8dfa961ec1963ef1d1147a66e3622011e4a7cab0d5fad4cfb610e643cbceeeafae
z2b3e00d3f0e479053b1d2c2e6160f50a9bdb7f51a49bb8b3501fd6a166c99918b34806ffe7de3e
zfdd91a9f7c1670c2ce64bd2602ed4d1d5237336b05d040fa139ca2323bdc30820563278764cf60
z5b893946e90f485ebe517003077f34cc6eeaea1cc449a9463daee1f24a6bbb0e93e19abdd8451f
z28e0964ef83e9de10ad1e9f066baffdbcaf4a5f20f05d8e33898a1df27ede99088b30db05e438b
zc9ab88fe177b0cd2a0567415f8bf5e010f95ea62dff5e5cbe9f5075df6c481ddd0ed952b53b7c2
z5e238c0e571e3e92190ac9dff6b47af48b9ee5ae5cb3569c0a1bb82041e617c418f18ba209f1d2
zd485bb37c7448d0aa4d61066d3eed8db1fc21226995f1082061d9ec2d989c64bebaa9ede4726f8
z509ee9e15e355f214acad808045b366a1b4e9ad93d14291387ce586ff6f94bd8359375f09c35b0
z3817691b1009d9b5b3d650efba4e57cda63c29963828aca07195157bc1aba94b1b94319b7cae9e
zb1c1b3b2f34b720224ca76f5c1f8cf770cda937d1d1d2353dc7c69ac1df7b1e655cc33b60b4f46
zee9a983419ca491133ce91e690e8dfe7ea8a37dbad355bbb91ce80c8a4497973d0f76835061886
z64efb1b0f6b26b9ba68f9f4ba1464a0f0b4f4b506dec309125db28bf0bf3d4430f78ecd4226b28
z1daa4f10b043fb7d5ca6a22439ccbc5c8651aa11928ac198401e2321fdfc3ad3c578c5d6722919
z11874ba1c89a18ab1711d9ee730710737d183b94f95b2b7aed8a6f73837aa13528a5f5a46f1efd
zc17ac2e195bb84ec5024e0d3f65b460d4141d426270716c4e15a6e24d471dba5ba9192bb566d33
zd6ff821b928b9eca91dacfac3acf9ac2d2811bd13cad79eeba70fcd4f7c4f1010515e8adcc1beb
zaac8459a46920d399a0e38dc9fb5144e4e17424115fd4847e4f8aa88cb07cabb238fff4ff83dfa
z191c2f944c3e29a0cba44a0d917cccf30a1abcb26c1fcc014351bd381a6f2d75e1276d8273edd0
z7a6f886cb8430e85fd7e55596e43cf9f1cacd5a4acd197810bbcf94ad62727e82eabe1e28e5326
z56dc48144f144cf1068280fd4bfb5f157c698eb87f7b20663a29c2284051cc45b0cd60b77d0d11
zc53e5b09c09bcaba89eecdc1406ef01358a8911330dea6b5642bffce734711e615f3b6abd7ca8b
zdeed4e9e8e862f40cab3209477ec8c1ca648d8d67234b14015c7472616ed3925d7c148741d8930
z3c092811ce4c9adfc05838b4812ca7e4c0f54c5d823aa45b147c345a77a70fd293e2f0538ed816
za084ee94944f97da085e37ebdccd0e5995190e577a6a288218a6ce3df766d9f15050ae91aabd2c
zbf7d0d9aa0b73e039a68968a056e687121107dc36291ac4986034ec63bcb953ed7309b0d237205
zac2672b62b7a3be8bc1129177ab016ae552ebf84067dd312129c880ade62f9a8aa3684c5736795
z912ec62a562bd3d6a9d886f351808f288b8e0cb1f6fb15d632424d688244a945bd0952f9bde264
zc2a69e927cbc3694bcb1f3405fffd37aa69fcc737612e84ae964ac5f3634423bcdc4617ee206ab
z54c4128ee01f76b1bad2896b96fc1c57e470fa377a05aaaedb757959415f07ae4a633cce26e7df
zca65239d16bf2a80b3323b00afe4f0b48e2cf3cd080cbce10a74252f4b88e188b720896484b051
z3392475347b1fb84f5488a1439934382ee664e187f50dfcc4435170ac165439c088cf1e4abd0fd
z91a60e0dee160a4394db439df9cce2af6d063d2f14925184bf4d53610cfceb694861232068f3d3
z5175677725347cda8bcd741fd6853ceffff106b2b91fdffc1991103494d382e965f3efadc434c2
zebe953a374772c8bb54c636285dde9e52f2721ad0b9a39199f7c484b63c4263c90d16113f1bb34
za779be1d49c89d4cc762177a94af68a0cae59472bcf59ff9a2ac788338313fc2beb406877d960c
z3ee1c83b61bab0cca57ce282cbff7d4bf88e2a8c4a00737d1604a6ab36a1507f2b84b00ac33680
za0509df38e8efa20630f595932239e5f71eaaea9bb086395715272b0babe2e9a383ab37ea0b19a
zaba8587423171816a272df60c608c8497bca914235de726ec006d96a725847fe76f6d507328738
z7931f3305d22d5bd834ba4e11c680b14c5c45b8552b11df66da427c1b74883ca78d943137c2cce
zd7ad796e2f2cc8a0ef6510e1b018bc413ce6401d08a182301f3b4499072f7c2eb0c787203ca866
ze5fa660b8f91bcd4902931a52f5c440182985b34547b42953c07ee0d227155e9c72379b1172c8f
z8757712c592bc8dd2bda41121ce475b46fb77c9550f88a3c6edd2bd33d9674dc1ee234a56aebc3
z21bafc421addbe06bab7f5cd5f05c421fa274f3c06ea3b1dcb05bb268911635f0d4c07bf738318
z05ad24a0bf4d1c5ca51eb1f667317b22066a1460fc6b89dd4b2d07d8b0b63c8c093bf498572127
z792d8bfccf179b605e0d3c2ef3da0e4279c2c51e9826ea6d6a558ab96180156a1bc835300264d7
zc691d52482b680528b4b500343dd51e296acf2448d135c586ce6d61ebac1b73fc14aad3e01c393
z83685acb699bb2ed2f029051e4ee0ff4696545cab6d3e9532a3f63049315c3c7cd7756c2a9ac54
z30db99824603da1a017a73033aba5b44a0eb57afb0e325055c6c2544075b1d3986ad3a8de13988
z4d7e3f059e195ce7d6ebd94b6cbd35d78b67a988bf2518906da6d8c9c7cc32f979d0267fa25f5d
z2f8cc90c941eef0dd31daabb592811e0b4c9c37fab7a0c42ffc426fe0696fb212a1ef84344b0ab
z3fc6204be3e9b02e486b8477b3c3e498a94d91afad217aacbd292fdd5cf70d270c46651a27cf41
zf4a6b08e3f5b6690672c1ffb792a64370c14fc0aec46dd44090f140547ea0a725ddd7f900237d2
z55fa768aa41478387f2f88e944f7897e0eddf1ff61351d7e5f4266d4d28aca574aea9010ee5a65
zee4474e273a0488dcc182a0593c0a1c2451639abcde42ff9b313c557cc67748e19c00cce8f7993
za5cc003d255b5842f87d0878ad8ee2acb9f8a1414319860e3917bb76ff35a76173e38e149e987f
z683b254a508b330ed298ef6b290082c89c214fb3704c781fe7a70e0315fdc06444f7268e39789b
zfd82b033e362be235a39437e54f8f05f63be1bbe9bbd37fa97eb01fe9f91cfcb5675212a52696b
z1aca35ee4bdc911630e1e5c9c830e2ccf3c74b2b43cbeb9a9870bbf747417213d658c0787fd2af
zbf836bcf8aed16f9140dd87faad30558823e18b9b1d0c5475c7c39e1cb9d0eebd1651d1a06f5c7
zef7384f98e802a5c5375805f85bb2c019e691cb79bd6280694abdadc72630524823f8afa164b08
z19d4c3356faee38d64b31cc50b4d6473c5e9d058e1f26cbf39431645cf242cf3b2c38f1b8dc284
zbf62f5ca7d91f36c64f45ab136ce31b3d25124ad4cbadae0afe3bac255e9eb0d5b3ee7ecf8b939
z9a24e7237a25c96c8350921a9273dfa98e610a929ceb1278d8123141e4d5df06fd30809053f082
z57f7ee01091d38f7315ddee8cae5c55bdc7d76a3457bf1b61fd0d03eb504e36bfa4871c02a0fc2
z62bc6b26c39cd57268577ee4cd44f9faa4dd0e1926f9ea6357c7a6eab179edaba8de3c80c4dab0
z91701cc508e3e35a4d2b9dcca10abca8eaf24a0341be474265e33cfb19bcf07a3d78e6ed3a8271
z12f6a4171917b04716936558597cb942bed6d0558f99ea7b9f56571bf37bdf6d960ab070ca1aab
zb0cf1e9e823a289c195251923c249af086716e8525d4eb63bccd2db24d5e68fe77ad7ed2e515d2
za63ae95515da59b1727c939cd06fb78208a138785ecd04a736ad929a01ebac3c5829db7f781929
zbc0a63e3d730f54d6bbe9e1b5db3f7d4b16e09df0c5c5f7cb34c016fc1360231e7ed11c45ce8e0
z44f912c0e30283859a285a778ada4584ca5e6489bdfc29b2e33c8b0143b65d821b80844a589fe3
z581ac86ab944ef345fccb8fc77852db62d4ee95935feca7c82b5fb03e49c4153c52953df265717
z09e7a9e47ac4a2eca4c4e0a2729d3d111ad209c731080189a101c66569b1de4ea174b371ecaa20
zfa8dd1e4a0d98f72ea9542d2ccbbe53765e96629dd8d8705e8a62453fe083231c70546042b4a0c
z4fffe081e02a3e62b49a09cabcf70102635f2200833cc56045d957d24686f5f9535f8f3f355e49
z71ed01d18aa405d26cdc2ffd0792022b5b220464af1fba5a2f970426f36c3b571065d7516edc70
zbdaa44e57d39c1ed3daeb60255fa7e8c7d0af8ac6e3305690d9f91824fa476f8d3677fdfeb9dda
zc9adbffbf67f09168abc8bc407e3cac85c48019029f0a91028fb85161d88c6e008a58a3440bfa5
z10a044cf799de770112dbb370058fd982b4885911761e2ced254a96b1706b6a8f9d1de41e65f64
zf67c095f40b14c694bb72353786b6031dd925064f69c587905d2609ee8bbfd47a37fc94ab305df
z8baa797f94551e495d6030bef4013f6e07a8c44b7139666d2c596882d377e8384c875e59a582b9
z9bb5b494ccac132f5bb45645a85e49be4b8466702f4046256774929fff1395f2513fa791fff4c0
z37ce81f92ea1b37bb1ba5d5cdb32fdf20b90b676fc8a5cc1d5c93cf7590711f7684963bba13a27
z3b49f9a8115adb0215737bdc3b502c83c7c20de03c44a03a6b6a54ae500e80c599c067b43fca64
z1567521a9bade7b4833572b83a6a09c47e8dc3d593564d25def245c8fd11d11ea4e852cd4df86e
z8f7a76070de793ae40a9f06774abaeccb069e57cc9c9af28035090806cf22baaada46f68076503
z768f5f2a1f48f753fdcda9f5e9d9288f65d4b25362095eea8a60c34c1b2bd315b3a4e431851119
zcafd3c29add771389789dfeec4a3d769472b9f77b4d7ba5de9aac1fa911ab157b3c4677c699756
zabab71d98e0fed5bf46ec4a0fdbfa1c11dd4566e53705c5115eee08b6c833fbc7fe4946dfcdd49
z91f3c6b55626a32d66ab6120df8eceec3a7bcb689639c4f66b845ab0728b800364967b8f8def76
zd8c699d27927754dc72c21c5897690dc21edb2d0c304bdf1514d359c064c15d908c22adeba640f
z97f4493edabd32e6207d3b8380bd1a78e171cf941fa4ea13f6caec04268a7f65faaf9a0c0cacb5
za03e163934ddbc85cc0366f1c24a41988afa30e04d7e56dfa7db75de244ff655a390777ccd0170
z871b39fd212ab5730984926dc9c74f70b7c22beb4b7ff668346f5408bd63a3fedde05c9f03b9d5
z35644ef34256f2e585972cb5bf272c749cb00b3992dbe7dff17d1ec591e319cc8ed62cc20d63db
zabe43896daadd4ec4a59b34f785a96557900035aec4045d8ca507c58a8d15303f2f34f3abe95e2
ze12a09bcc522e178da40b5dc5abbe1beec6f067df2ddfea0b0fb4ca55775383e908f6576074b3c
zfe990a2aaf99ad6c40cb2997f5f8e219de803dbb435b02ab57f25c52c681d03a35bd355d510805
z632dc0437b221f7b0ce9cd7b30473b83f651cb230dee1a60328b04f8563af8a4529f156cdd137c
z02260cb8b116c7be7a876bd01118a9aefad162675c28b0cd92546ab16b7a711f6c62d8f5dbf3e6
z50b8432281bdd8ad27ecb80d79bc355b7c82a5141b2a13e20d59153939ac0b1936f66407db8528
zd0b040f62da02856d858c244d069bde34564f69c292ab4a83314065672733c44f25fd6f6dec36a
z0e6f2e649f4b2862ad6a46dbf80cf193a94c812176959592a19671a3d4f4fbd8000794a732bc46
zfb43a3576c81d6d1803b79b9177bf0b71700036160cf94989fe4ba28fc5dd7ecf4d431c2d7aa7e
z46f91c83418daac0d8f36968cbd7a4d45c96fc6cee8eb83557c8b03ea44a2d6eb7938064bec675
z2d1faf1207a3ae2913f3235017bc035882d69e36e5d82b201828fc6ffd9f327ead214a2493b138
zf75f81d8bcdf410a32f046fd287376f1614294e797acddbd8b2bd3a412ec59b36c23849f525032
z5c2a95e1612cab9d49d1a1a9e14b22b0e71cb50521e937efe38bff84e279ae8a844ae518c933bf
zaa00169dc9132e734d9976883242a9670b846f511f8cb1efc82b7263a26997038aad8908f0fb3c
za4e9e17576441476bd0218f9d3fc0a63bd42def83ff3a5d1e3906285b905537c4047cc6094eca7
zf802834443763698208cf0cf601ca03d7dc8bcf7a9eae08687f2a2b99c8f37ea53373d731eaca2
zfd46be1cdb19ba980db935250110b71ee062b86d7f40910cf320a694ef184406befb0ffb97b71d
zc08110eff75a065a6228329361b51aa1d9f1db940cfdaf869bc51e635bfae086800734e29f8e80
z9c5ea1aee7d35b227d76a53ccf309a9186bf4032b0b27325d3c2bd28e0f59484727eef4eaa5a04
z8d21832a01d769a76cdb1bb6f7c3cb9f10fe192c9012c16141796a31049ebb739663a7f4effff2
z6aad9c5be413536471751f9d904498d24a7bcb16e3426027f82cca26fa84abf847bb64f1c2937b
zf3f017f0691436548cb41c9370052ed19f6b76a050167e9169a337c529641a5fbaffe8d89f5ffb
z776a33b7818d9db8a950bfedf8519f3e8c362a86bf0a1b5223bbdce4148c1c3982429ab4c1a030
zafdf31691a345e06091a0dfd16c1ce5847b8159ba137be3b9f2b0ed5129b816a7ce5431569783d
zfeeae35d82647be7d99d087a859300ec0d574347355647b11b38490013512f12ab3b66ee0e0149
z2626c4f66610bbd895be2a4e7f18fed93878e12e1a528ac31bf8814da52964510688a1a9b18b9f
zb009fb3b18a5fe775541f63b3f7acf7a00aa9241ee7e468f4a044e8ee1170570e30ed5e315d17b
z51bb961c9c1cca7e4a51720200a74dec8ba3dd1a402ff65cc0a28d4833d98d5f2e72f0bd19976b
z531ef6d991559e6894f49fed0b8cd2120a213a6d87debd61f09b901858b25bc0d043756121bd8e
zbc7eb01a4ba1db0c466d3e8597d12636df7ba634fd8dce704070611402f7cb5057ad1e61f7f74f
z1086dc66e9822572499b70741c035817fef19185ba19ada53d98b496129a91ff5b5066eff2427f
z78031419be657db592f867ed5df8b0b1f55b95b9812d34a686366a7ffc505c691ab04d65f1eb82
z19728f02d4792c31bb807f8a973393bef467cb2bb592e7eb6c97a293666fd580243bd54674fea4
z79ac1078b697ed2129502768dcd9288e122d7ff2986170f526a4a7b5209ba02b86a9e6fdebbc71
z1361aa1fb0a947ee44c300002df6c6838468bd072942e85191bc332a8d6ebde56dfa1e78b21b5f
zb156a7cbc0e57372f14a7206fb0fd85742ed3b2150e35c9826f1fed9f1b660c6d61d57f6fb7c4f
zae3338191bcec6209cae949732e4339b0e5ffa472e5e208fa94264f5157813a7712bcedb257aab
z85b65c15dfb9d590649a8a142f761629ea08adb08c0c64cf69b8279954189f06eedf650a5f0d6b
z990778a1fc3881b470f18f2dd0e3b0cca296ed00cca7ecda502c34d5754ce5a6a6eefebca7908f
z16e57b13b499a18ff4cfb286a6e11a67e949c566475024255320a50f84fe99e49a0fb57fe29964
z4c3fe2247dfafc1907b3a65fce0ef6a0972ac7004b8e2119dbe637278e4e25eb8155d42bbcca19
z523051da3ff941d08fc7da47c2fcfa16d5d03a92b87d43c750e7d9041f6b3060ac90b3f8d74c0b
z20feb0ad7a9950b1f341b8cb289dffb483670c7c39f1e8259714bf667808f3dc1e65781f40a515
zd28c6d27ff583b36745c0cbe56b6591b74d19fb89445a1697d99c6e2628a87dfa69798e2e9aaa7
zc0b9e0d50f3e02f49042da1c9693e35232b96fd810a789771dd388f5a9730e1823819a9422b866
z1cdcfdcf6a0f1b70aaa7114b154230a63b7bcde4ab0a59c204447f26fc12b67ffb2d986a34457e
z756c6ff6f07a614ceea8189fd4e767e11fa1c1166bf64849c0d36358be8bef214c94a75d4ed8a0
z3157e7e8fbe686f6f7a44601c47b7bd688ba9c34c8975dcf2972bde587848faa317e5f8fb43d07
z804040e81dabf3fce0f58379c68cef45776eb8a4b7ec6d3ab631dace4fc701db2716ddc9ff469e
ze1756f0287cb5cf6b830d566f09371fa7c4896f8c8bdbc792b37c5074284d957bfa9305ec78b46
zc5fedc13faa296925a170661e965491b3c468c7490986e2288d78870463ca219f65e768155a82e
z8ce67c9a85233ad3c00312df6308b4159828dd68f53cd223007ab20fbf5043929017a9dec04632
z8610a935b885c1339a90b3e51d6344c7ce03c3587543addfe4baf188ac3ac1419246c8e2b45d1d
z0dca3ba3089dc6783f9b1af9c1a097ec7c52d1d553e6fb287ccfdbef9fd610403358656c3a8524
z5811cd4feffea1bd33ec3d9b811dda75f87b6e38f4503de03bfdee9809686d99b9474ff2a5ce5a
z229e2485a5ef72de8d5667ae53dd55342b5c76d6ff8a35175b075095b7c87336580c3c343c2be6
z9c01d806134fc9693e6273f6c66ebb9722c572a1027ee20bca9beb7cba1e1accc425c5f6bb9cdb
z902c7095b536a423e5914c132d89e0111db214f8b7d79cc7704726126bc75175a73286571f24e8
zef4e399b0c62c6cfa150fdcf76e95d7900bcd1f059527a3bacf3568fd1d8e00408a2d4b0615cb9
z676adfc2ab355a6147c67d706125d2930122a474242d69a15b538b5b8ba286920533eb7081d82c
z2bfa740173bf81855747604f7853ee3fdb7ea7d4a130f67d673c70805b176cbf96f6a0738d5519
z4ed7adcd02e77f7ac9edc93e2f20fe36471512470dd747b371b1d37b79c552603d6bfcfc13d7a8
z713b3489451224b266acb30022a33c45566a24a484be5271b3c2b699bdd49a087a4a3118d7fc42
z74d70d964fe1d420afa630caad3ce8cfafe702c01c2543bc70318c8a61a110e8fe243f3bdbf731
z132b9e922a52e8b977294ac783567ef28329aeb4ae4b066b85fb1ce32a03d81ffe834349ee7c82
zd1e16d50736c75f9ab7af40194de8ece9fd5ce40008525e729d1b11c7807faf7631966ae0ceb25
z98cd4f00d77d1c77c7838a9e16131b8b5ea38eec8a5f2ab18d6daf095f2e9e7a9238eb19ef4971
z7becc8eae1e3df885e36513b04eaf41ae6ecba582a66fd3af7a5c1d39789f72c5b283fb7988f57
z25bba9210262715ec2a837b145d9e019e317634d852782da4d8c074258416a82e2c040dd7fc04d
z26f9e0a727651f8ab4d4d78ad2513501e5b3e45294e2565b2dc1c95a26c6be2a8d5afd5cd78f5c
z53aa06119ddcfc10ad05b94eabf0e576e6fedcdb0855598b8a1638ceec533e3b6ede3d893dd86a
z6c9d4a45367e3901ab375acf6046099a3f0344f44ef284ab8e622190869528ec85394c7ce69f42
zd91fe654d01840f62833223779ed008525a05d0e6d606c8e346b7361c715a19a56d5681dc71152
z6412d9532f78365aefa6f85b1b4c10fe894731f5af09fd160bc8eca3c1511fa02a3d82b26d8099
zee828ad269ebd120b649ba137de5103b3e724191194f46631cd77fa5292ecd551507f4436f7b61
z5a3f755cafc3cd683cd99a0bc7486ebab0b8662876bb0c5a03cdf6392e1f26c1484664e479949c
z0761331ca834796f63d04e72a739731c73dac70256aae7f34baaf98c5361cb273471b5cff83225
z8dee51b7040cf8e465800ef7fdd1ebe324780da55fcb9ef71b074b1074260f4b631a26a6879fad
z12bb2c514795714cdedc2f01edd4c1b7bf42cc5022a0c7a2f3e15f5bdd3789aa854563e12e5725
z5d5de7897930b18f31d4c8b1d96ab5a96f904004f3e493809c123c0c01a163f5828be6e36613ab
zcf1f1ec4beee4008622a20c67dbf1dbbd83f1d75c4f106dec2bb2f5ed8c8f54d8ec3add20527ed
zac2f78e70a4ae040e2596b9c0be94cc03195ded0538e011368206b8259075a9e8b9697c339b93a
z0e9ff7e36caf72fc4903740fff6d4eba40b92fb202066d604055bcb9ca0ac423f50cda69dbdcd0
z0921a29a8f4695ed045d1766d03369e43a090c729fbf9d0d66f7d4c9516ad1f951bdfc75c2eead
zbf885a4372fe241ac349e089e880d9b3ccde3616593db8fff255a48de0a90eef2f8ee9eb019421
z55ebb4116c7eea881e8b4557765570dd299795bef0ecbefb583e7e129c4ec09ec6a290c6b37ef3
z76ef916e1e5e14fe78e69926e52e35f6f2d1e1ba4fac204b61f28b2814bfbb9e74552ef026af63
z8b04512edf6112435d6850c9b8f686d12788c40364e74775a2f3247c15211423814d788ae45b1e
z6d832fba3ed5e2174cdeb87d138a9bed6051bccf3edb8f4e42932f5ecc8c36212998ef6d9f9b94
zd3109d1455bfce1683e0427ef39021ad8078c6f02fb85244ded1f2477a07912e055e1f62711430
z3b8bed2e9e8c502c33c565b6b16866bc7c89710521b6581fd1e81d5dc325cb4ed247d1eccbf444
z467aa482b7d13246b894a3d942472d6aa0471646d5f8c7ae933807c358977324468b36f57b0a4b
zcdf8b77e829022efbc83811aa3ee0a00e7202d5cc3fdf8e36ca4736fae35548f5988bf580cb7eb
zc8bf8a2ae76c02114fc11fd1dc645417e612d784bb9b660d42bfb62b95ce34aca81c7dd3226ed2
z73c6b84e59a872f402dc5b9266ac72473f593da6dec0f33e16b390b62245a0bef4502d7288675b
z289ccd7507dc35b93ee4ae5457921c6c14ae05842d341097c79bedce341ef40a96bc9bf7b27c68
z1979a83ee1e64b523d2aa426716197053836a7b05e3c70bdc22abdff9a955ad674c3cac258fd2c
z23e65aff375532279d68263b5b97384d07d145b41f245bb2e8aa953982c7be72a5045a7904df0d
z6e7f01106ec1ac3fd5cf411150728d538bb053e7423440907595bd4d9480619111cfe6bd37c576
zb2497e7652f75ab71494ba58b9058cad66371ea5f76e5713747457073cfe26c1d8b8732b3c258b
z81d9b33d21a87eceeb7ada866eee27dfb3c6a69f145308084cdbe42f81bc0b41a95bc95e21f264
z35364a9b1dfa1b9d7ba35ead80194a037d39c024bf6b5d206826055c06677bf1478782e198a547
z313e376cc19c9419e9ae0ce98b24f0e647b965a1e0d03427bab0bfb610e3e7710220e0df0a6556
z99d2c4a361e510c1f0de962e51d08739dc6240862781fe8843b1630bb57d5375b8452f40655cfc
zab3aed3972f054f56cae64c8aed4557443de44757f942a21987616e8aba3d3105ac9bd7142fd53
zb957dc671da138673ab8821d0c672cec04ad5b66abc70a99aaf2f229ebd1a766aac1505c97b32b
zd1e5779727cab30424f2362a793436efe0ca76d55f7c9225ceb4f3641857466003b98febe50144
z29f320fb6d7a78bb0b71827a456ead3f255960255e24df5f5ffa89c28b1b64eaad2035ad8446a6
zd85eaf94d046bbeb3616d8c0044a833408e08226d2d383ebb8057893f2974e861f3b11e0e73251
z55670e5a552d0d8f4f27e628ee5f6bc9fed55126fdb44a581ffa7d980c5add808d3de962487c38
z69e49f075d481d96e3258e310024d74001aac54db874a209531c7e79a394a60bad96af28f5a4f1
zaa5980782b1448630d0b1cb7298c87b095b8cefa18e91d2f56abaedcef5c03872209f28fc2979f
z782909a5dc4840c62b7944414c63d2a2e1829954f2937da5f8fbf323156eba0958ebbb88c401ee
z91253dac04ec50273104a92231031925d3d8d61f9b2c287fa04864e41f04cbc2e3a36d65481094
z6bfcac7d6c2b25caf707f7fc8b81459bab09f97e92a0df672797b91b0c5e8c64a167a61c2d66b2
z76651fa7a0e1374e0fd1c8c3255434efef8977f3f7ff989cd085bf510b07891a067f35f024e956
zb90b97d0416859e06e6e31fe61a575ef8b4de740c25e362f0ea8536696b50f6642b967a7f1b9b6
z37b883348d5adf8eadc2630ece88b4737db93fe8b8974093e051f196b6b55bb482e67f1e3d18fb
zf0df6f365a06edfd106df738c4c575f751ded99f74ca5ad90e0605505c1069e01ca5d781678f9c
z7f996bad67082e675e1f51106d5fe19a26912eb8a36d32d45cc382c432f532f9a74e16c4c7e244
zccf9bb4e9fe259d1e9eaf161e25abf17192a95f79216e06f800029c783edd87c0e6c22d4569c41
z80c8797db9cf7e6ad7473be0d9596640ffb203b88d0c7ca328fd73a2a4a54451c92cfdc4c036bf
zc0b0fc9aa027e9a36745c12832417dc1229c51312a317d032f4035dde07d19f0af1ac4a251c892
z85054ce4c78eabef7710804ce59687deac7de9418b64015925ce177de4dc7562a278a7abc1a375
zacccbf5ea777e9fbd23f35e6bcc220ba21f1b35148d37eb0c9204590871529611689ca061f1c61
zc72ab30952c644e4b2407005e7156094fe8eca7396b95826ecd98d9b42122b8605cf1ee984cd53
z0e1cdd06fdeba1ea7d64a471c16efb2fff968314c582e703eb9e45f6a8560ca6d386e88761afdd
zdb813bb1dad8e0aad56b262dab5c3eaca7a2ccb7b717b4d3e0311a6a29927b2cde7203ed9bb2b9
zfb60b645f8614fba1655c3d3619e3d3c0e7e30b3305bb6c7c4f10c8a219fb9124efe41eed0a702
z7c910b81f4d730eca2b74f139ede4f2b0853d961376a67c56129dd01729742e1da859db5043a2d
z95aa64e9296ce5645779db0a7fb385c4b367717485c7773cd81e3cec5ecfb0e3a263b9b7c5d3d0
z5a29be0ac2e8d343aa2aab2526cfd6b35154f70cdd2618170f99e8ea6058d5946a52e3d7ccc336
z6ae7c0b6b2f5860a0e82f370410c0ce2bdbcb236e624955983913157cc80d4623ce2f25d5b4233
zddb71efe1a3cf7c790735ad5df96fe332a492e575066e8b368c9a86b768d19f313db179e5ef01c
z4cabdfe3458da5c9c6624c40b6d5dc769366065736cb5275e052a7ff27ffe067969352cac4714e
z5e4f95dbcfcfae84b12ac9de1723e764fc95f2446adef2fc997d54ba3b03a0bc14ad7e25857c68
z5db1f7a7e35039b49462de452c366d2b1d2dac7bec324bb9c58f7ce70ffed03b788b7b00fdab80
z75019c1f095c3eabd4bde82d95a60b3b078c49ddec3ad83e597c27a0bc5642a9aae3a96f25cade
zca670e889f2f307874ae2e60e196612950ce51ac1cb7ad66d63faec85c66c8b2bdc0cafd8b54e9
z87a6f1c0e0de57e0d5a7344ee855a8c11e58816d10d4e5e9ada03a8af492099b3b104cf08c6087
z3238d39779958bc096e1e2c71d730a3ff43145701e5074ce9c1622ee9764e2d1cd9df94d49951b
zb9286d5c831bfa716e4281fa13033701a45023ac91c08e137145a8e87a3bf11f2a10db86d9fd34
z70e66ab94e575f24b6c4f029013f8bc47ec691bbb36e078da7024c6bd50adaa234f350ed6b2f99
zced2af071e6dfed959e30e16f00406187fd49b6e2caebdaae0e9bea6aa4585ba6e0066d15904ee
z402b438282760cb2c8bd75691cbaec0b77a953e3f19e098df88c3885f56ef1d72012838e775c5b
zcd55b1eabba87dfbc9a1ec27d37275088bfe0644b5ec8bb9345f9a08a3d3e4688839ee12f57b7f
z8fb2ce313aac5ffebc166f0d3892eb62595dfac4036346bc24e40c421e5160423b78a7f7b76fdb
z9320f1ff19fab2102cf28589109956a3ff4b4766410c18b63265cda942df1778e19db78ad04e29
z3c2111a712c40796e5a7cc7bb2f5ac4065fb0442ecb8025420120c56648932fb5cbf3f3bc8f225
z672f5faef47d2ef62ac4cdfa58fda59e001e0e45eb694d6de08417489ac3473df97c0144362bbb
z95fbaba8b76f14d789bab96f5218269fe4e33b7111d867a1acbd0e96774065cf0422a55b698597
za02c49ff2f75980e143c0749996a405be41beb89c1c44ab51a064ec99a274f9d526e28e992969b
z53917bf4466b2ceb018373093b514dab491e96370fc7f6d2d1fe1e4e8c75065265f57cb8b30513
z688ceaa518ead16e8aa12f25c9c7dd7c8ce72fa853ea90840147504159c95ea82fc8cc2e7eaa03
zc33fa5f328167a74cc007828773146669c19f54030952a73b02a0660bef0067e596c2df49d11a2
ze4fb84729ce1958e11089cef1d6253d9f7e7a8ab4c5653cfac00014691472a9c2b0b28e4151df1
z7d4f57df2ec3fb02e6d3b970bd73d8e5edb3551a0395f9b8c35cf102443d3014f69b5f5bce4180
zf0225385f7b3f27b1381b8a585a470d27c57f5324ffb6f23fed73958c68bab54fc2b2b46b5db7c
ze423da2775872e1588422e56834b6d005bd13b0b9fa4549c957891036274c7590d848958c5b9ed
ze1e8c766808142f367a973680a9a62c60d2247873610631216e6c9031c4e72dc0406e62638996b
ze0fbfa8e0280a8ac7343ec9e01fcdac2b5b654b1a058367195e0ba9b7af572e0ab451014ca07a9
z7eb00d68149ff18a493f355fddb9f9270aa19ebac5c025abd50d1ead00c82fb1b08a64c27ae0ac
z69b16297ffdc6a519c187051ad358556a59580e49619bcc75b546f102fe912855538b378b1d686
zfda105ddf66a0a6dbdb4f6e0e7b27230136c5f971d9c00be6f01483ae214d1902974037ca10625
zc2fd529f699097fc649421ae0814e87da6441e6b33c38f068ea62a00a900e8e6051a4fbfc837fb
z89026788b2063ec7a7535b6d359a2fa4f4796002391ceb92f9364a2ecceef013efc62683ee7573
zcab103caa76326a53565b801ef6140709695b6795ffa8db8e62b5f91cd61d8d9bded35b652317b
z4010695220003de211506f54ed28af30c284c5f754929f585605c8c04c25b4812713dfc3c8839e
zb5a5126237c6f5d22022e319d6925cb12cfdaba489451aebf1fca3770b74f4de8664ea7f6c1549
z6b07e85d2b5594b83818358600714920304768e3ef9cf59abcfc1ff93ca6fca8e219edae76c1e1
z8a956f899b7bc43fd573271ac6b95f1597bef50a2e22f7f8eb5df89c21e9be419e8651fab5ef57
z6f35499c6373a02ee11347f1a8ffc228e1c65f6ffaac33321fe9df52b5040951bcc8c7d234d675
z5479490f1320b283de7aa9d825b5c2c5967e78b595b8f416fc8c3891b3141fdae212e2cceb9e59
z38be836321879ccd072bdc1917aba997bab5db3d96ac6a7af7e69ae01aeb97ee87f5ddf5152a32
zc9fda50c150fc858d7a892b097217cf246fb3eb2c30b4557811a5bbe2d545376944833ead8551d
z2bb4c144a032fcf9a1ec448d79842177c61dc0cc9c6aee5be36dad44b005704106cb9f3d6f9441
z678d48aae1804e3da4ded427442ea5c6c17b36b80784473cea17e6fb992523e93725efaead3673
z58e7245f54b778c10262bda4a81b9c53213cfe516153fcf9c79db4ebdd60665405b89eafee18fa
zf8238a1a099f71ffa48254d0ac0a430eb5584d7087dc97531bf17f39ad666047b18b5a03d83195
ze27c715313450ea219f8bbdab5e138b498833db817ff9a19827b5d4bcf9677e03ecff58d55dcd3
z08263424e597f1a229191194b1a9c25d9294704fbdc84f5b7f6ad02f52878479531690f13c5688
ze6ecfee3b56d597d766bb8e4b7fb010a9490ad675904a362a16defd43d4257733aab572d6d1965
z96b39c4416d77502a7ebd241769b36e3be6a70d95343f789ac096f4ec93333dae44681f821bbac
zcb70c910102551ac278a40932c4713184554eca69ace23cfd229a558d27801a8f85395ac56644f
z10ee327806fe562faaca0fc88183adae07c2840f625c42dd53d4cd2d23a4ba59113eab2a06412e
zf8ccaf66cda198ffe4fda3b108a84d88bdf59e7b3f1216e4b1338ebf392bf29f2884130e6e867c
z4d1fa1c2d3c23fd7c437cc95d34e2562cc02b3de39b421695add9a49d70f64b64097b0b17e89e9
z86279cf87edad78e25b8a9b60c64f0b05fd9b46261306d0ea85487655de09383adb12d0d418363
z76325cccd0ddfbfe80a1ec558e33c9c9a49a201789c83444109f9185e7315de7e4d9fcd2485814
z6b439a83015f6befd27f5375839509bcab5f64e87f01800953d332e1e3198ef057f47164dcb6cb
zc077bdc83170962ddbaa1a49ec44866f53178d3732b7cc6c836eabfdce6ff945dec4846330fecc
z95eb8dfc8f544be5af82532b1f12a6709332ac43252368d1ad01e33b11320447de007ab1135fda
z097f15f82a9590bc3aa617a5d596fafdf20b9c197c73f64ce3e4bca7ade64ac121d47fa06f319c
za496a600fb45d97d87f593af5141745ba4094e97e34acdcf04f6d511f243e66f04c52af60f2bcd
z02df8a35960c688e1e3f7de2f6d579896e43d48ad06f8a6181c3b4d04c1c2b0adc26355cfacf6a
z796609f50f40bf8ce2ac42cd5ff4df0f797bdf4eb507acbcb8786319196987125fed235138d60e
z60dfb448129209f09cb138c87f825a7d7c0af45dcf3dfa3eb7334c75546f0f03f83b24a585328c
z5371553b0bd3620aadda3e13294362b83fc7b34e4c2339d64f9a457ee7b3caa27352d02a311cf5
z401a605da1f52147da5acc580baa08ef1d1cc8e5d3680c4326d1be3423cc654d2f73f8caf1757f
zd6bca4e628d9038e7865a568ce26deeffd1236bbc0cf1881f950bc3843d094e01cc0d68a5aa984
zef964cfd5b2d9b1c8a736ac884b751c590fcd5269107a34a8c7adb7056e253450942a2ac9e7ddf
z2fcc4b68aff91a4ae9f5be67f2e14b802afea4fdaf9fa844c2d27369ef94ff00bc7ab05fcd77c1
zf80eb70a843619aaf13958e519732a6bb3f6f9fde63f41d0fc3d9f35d47f8b5d4d964896e14ec0
ze026d28d2f9c856fdf1f42bfd64b6401afe5047141ca900804b0a0a573f0e160a310609f3024cb
zc2868d6f3336e8e982a82bde938c29b366d24fc0f3ec265e7f15026887494a058726950e844ff1
z12ecf5f453a4455ae42a5cc04710a3cdfefdea166861d2c1b3cb3a383299041cd39bc26338d992
z8b8a43f0c4e2bbe9616030f59027ad9902d98034364ade1b454705793a3d328612486bf717c57d
zff99c48159018f1e6e92d731cc3c1029d9613e98a06d224f025d17b55f72eaac506724b605c72b
z353a35206ea4f2dd7be7808421ed6fbb834d208de089e3928bcf9b8bbb007d650f2f21ff604396
z2d50c92090eacfc258aae45ebc297831e26818b5637dbc5eb1da03a288158010ba0a0b1e7ca701
zabf6e1c1643637a6ca816ad25586891044598655441a3525b26f929715e97b9ba9e21b84f718ff
z802c78f477c08cc1bc3a2ecd672b86e61e06cec224042b6ce573cb2cc6136ad523c27603e3453d
z66ea9cde3fe2daa11a02e374dc3b304c2121c3cc57eb33f94955c841294ae5bbd3ae417c80ad50
zdc306ba2656c6c77d1f47d8d6659df9bdc5444e8ce5f3dd275ea67436da3daf2ee2cb7c8f43780
z318a69bf4af873d2d411e387e8e1e202650bcb25d843d293dcf0472d19c250391c72c7505fbbb9
z8159d9aba6f90d8f3820f9719f153aef2e412848e6a12e01765b8dd02c855685365821c2f6d301
za6731bb2f2a31dcc5e5cf8330fe986af0437413cda10f5909cc7cd9535d588072f7df1faa02865
z772cc2fdcaa93eb500039f86d9141343adb0647ecc1d15a57663d3dcdf03ea6fe7c01a13963c54
zdd7ab10d55383a354f8f753db6c52524d333f50da332fbfb4fe2aab27707fb9312cdba2e7e8e35
z4e16596eaa0cef3e53fc0bb3200dd06a462e89e5760c69c4254b7ee2ca5c5f4efc5681218d74b2
zf3f7fa326f7e96f5998b019d09264c4da5fa2ae0640f098211ed4e473ecd5934f9290b11e8bff4
z1440f569717fea560c35e36a3e27aa85735e010260d1ff65d5bfd0e110bc13e93895d569c5451d
z2462640759ca868ab64999436f0ede7a1d975522a625881273cd50d2d854a7bae96757a38e152a
z24b8ec414f61a169c75d4c7c2b1c4be124311f4e028951a9cf8e080fdb25b4c631c01c8e2c33ef
zf32fc58137a5846f3f769d302dae3535f12cf6832a195de68ab119646ad5828b82196b489475a8
zcf4eaa3ac6a80c94feb2e92806b2db3d4b7710abbac7ce16d603eb095f13932cc9fc36e39ffe93
z04ab44f739db88b9d7362b640ddf7353ed52374794dfa43cc60dfc243911a27fa2e85eb062a716
zff6ada629c719594ce90284ae58576f1325b5d9e5ffe80c9abd93eff6883727cb1fcae2dfe596a
z969331fbcf6f44143997275e9640795d4583e4e8f94e26ff8d0c1b
`end_protected_0in
`else
`ifdef MODEL_TECH
`include "qvl_sata_monitor.mti.svp"
`endif // MODEL_TECH
`endif // encrypted_0in
