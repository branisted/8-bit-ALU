`ifdef encrypted_0in
`protected_0in
ze74c34e226135848fe16db9ffd31815111b6d7fb642c521a3f628cf6da949865580b22efd062a7
ze90adae0e65e66a2c36a587d0a790699161455169ed55a01f2084f11770a774ec4c588039b380f
z6de9c5084882a40b79a175f5c2114b2b6d78b070cb806e1c0aa9258297f4687ab30857016fc53a
za25afc8341302f0c829d94450c399b8ff9b0386c187cb854ee330605b7b59da379b1f26f488e1d
z36e675f0b1336408b3a1ad87d0723054f952fbefc8d5a33eaca6ef5be8f42bc59870a29a5cc9dd
z4fec09ce6e44cac279651402e7e1f590df88ce49ec26ab39f12b4a02855703c6f03b1e85c797d7
za357087d98e5b1f45502e45892e5823d6fa4b762932009620038c05d74efcea7c3fdb38901d620
z36515d0824367e48d1bc182335f158c262d396cada6b0ad58add4f945eee634c2dceadbfb5118e
z14969c29a743830a07124bfa78707f3952b96b0db7af7c9ff36f77137d8c490c4f79328328069e
zd7d5280e4f95742c9841340368b9764f0f80413adb175ecfbdf3c40716abca7b8cef6f7fe92ab9
z6bd2453f1aef7f7899c5365c5c83793cacc7795c269413f6cf0dabad14d40e9285afde8c01a47e
zb61893788ec5060288cabde8fb553f21b02eac61ab0b48ad3d54f4d1d76508b22f0c600861b5ce
zcb30ba708be817b1f50f59c0f6fce449203e7355c1be55b662fef3f92ba58243d81537761af8d6
ze27d7864d2dae99372b2b75bacdc0437a4f7e011d68c3487a89759e3625548fcc920ad06471ee7
z2d701aabf726859343208b0a543c73eeff8406febf277e3babff437ec820fb49d6b78e73bc2353
z884917487d35a6cd06d7d73ccff5f05355122888b886d1b7ae29679db6c9d2d7f218ac9728369e
z0ba3297b105b1781345d5dadc1077db50a0833d4730649f7637b2138ee147e4467e47d68c8e25b
z593a6bca87484aba5888b0d117862ed7c2676f9edaf1b7dff2a4c8c60dd9f44351e4f72dc5a0cc
z078e18bc1a3e16169dbe18fa92cf30976c736c34f1e53045f4ea0e07c779b0c89edd9128640419
za470c988c7537c955691824eeccec7b4044dc29db87904257d0cda47a378c392331eff47f59faa
z32e7d935c3f423dfb4b81dc647ebffeb4e5eb20af7a3dadb6c8c28af1cd13b2d1df46244422021
z08ffcfddd0595405f77411aaa3cb976db3deee12ac1d9957d2c9f9db27af1ede0c3a42b874893e
zbdfb4dfed03f6656c2b8a1497e95da46908e70237b4b661c7e12ad64d9481ce9229ffeba585c13
z7093f501dc87a2c3e79646199133e0d953ee21cc6fdbf961cf2d9e9be0f938368522253004c69a
z50b26ff3efd9ff1118b227c46abb2ba5820bc0e9687a2d93725446658af55a4ddfd48bacc1f1ea
z96c307e52c2929f482c753accdbc3cc1b5ef0dacbeba0ff4bf0fe9851df59e10c7f49d77f9aa3b
z2c907a2d33b61ac9bf7ee90f3ef2f242e7de85ab707329bc76a06684a3aec02637fd72b67c315b
z6f7d025d5cbce033bde9e941f363d450a204769871e3d4a98c13b2f8062fa1319d93976a9f4848
z13e4d2f7b4708f22f772242d494327e46a322cfc789447103ee132e8caac058ab50cd1ec83375b
z67771d808d80504e17fcda56fcf0e056893f4f911ba6f770739b4d0a5ac28351935a8cdf8a053d
zc65200eb84da471d85a1d1ce84f024484ce07ecb56a8135af56cd56beeb8ffa4a274aa67249d57
z27a94c8cf2514eba177c30c72c8a8d6d3babfb0ff43d27e13bd89c8e8f70e1a80d93fd5599d17a
z28ad7a7deeab8a53920129457ff701e664a3bf50e5ae8d0ac6feb9066eed6a9d606fda499a71fe
z96b7e751ec3acebfdd5e6893d038e6d4721d1065f6fd5b285e5747f641290a284d1d9eacff2766
zf38d88bb27fde2f64780a5454eb9d8e4d799f6a7907b3b7f2d42fb61bb2690011215507e5567fd
z8dac4f22a5e0a85cca75323de58dcd8a8a8839696b832cb2961a3900760e93a11af9274c916fd0
z012a617cc63a16ea8297b633e722525002e8602cb0c5af8a719777895c6e1903a26d074df2379a
z8b5c527ff74a591bf0d41bb7f254258cebcf043889e176ff06c4dbd55683b224a8df3526eb084d
z894738c33b308a97ca67b54ad0f18c777491af1e0819553fdef03439805ef6ea6fa8e2ad4baf7f
zb1855d8b618d2ec7f111fd868fd07c417f55dc16a8cf90bbd21dc0320c5dcd204b70d003036d01
zca710add3df23a0f5e287a3405e98bde3daed1a6f9380b406e8f1efccf5e98edec287fe9a9b754
z1a7f3a6dc4ed126573862017c736897f5d963a78d6b26c775a9cff1dc2156e2c20618d6f718af9
z37647117ecd747df97aacc43f34ae89ae8e9be39fefd8c0bca6927d5dadb32bd163e351c41eb9a
z0efc9844d79a2d42e8f86010661f5407b680e7cdd276b1ff858215bdd288abe1aee8bff917167f
zf7ba70dcdcf2b905cfb75a332b0493d3b8512e55c660d95605f65e980ee7d62ee5b1e35e277d79
z8f579cb6b3b87fe49e68db78af36c5edb59961b0819248269b2485333e757d2ce1db5cc75fe804
zd4f7de855cb12b3fa9ffa4f35a3a21f3a52898b6785fceda232a9dcd0291a85312eee695b0b59d
zc6273a4e00f7218b903c64a7cf756fc51efd19b630c13bc76c4a67b6ceb17f4fe650f1e998580a
z3c6e75d2f27fd9c42c35ec5e7d0fa057247143ec1cfeee47e178a1b569b82703c13176abc0f7f0
z881bbfb48eabf5c9a820a4ffcd16e6c4dd312e44257d7b8e0d8bf12daabeb6345f3db0495f92b4
z86cac0318e5cf653d339f39af08db8826fe12aace60ff1506695f88986d1a34b9014105826dfd2
zf530c063e75a81dc995311ba9b4157ad835b3f86b8d37d38bb3ad8a3a51a4c6166eb1b06f38ae3
z191847d21d1b7a370b7d6742cdb960f676a873fa65e30c732b34f8f3450daaba9dd8f0d6d85c0d
z1c09d827830ea24b9f27840e4e72f7a6067a1800b9b0d8e68b13d2d1de9ae3fe4ddf89cf20c4c3
z5acb9fb7c3340989d6941f7de18d54ebba072765188b8295cec6ecf4d0befdd91dd554af29af30
z261d6dfa94988c2b59c0cd1b4afc36c8b1ead333eae716391dd7221c8d86889b39b0b8793d334c
z2d4c918dcfccf6ca4ee2952f93d80ba0dfe3fd6cbd73c2b1183390cbb0a7c5726f5f3616f010bd
zc7df7063430bdc892523392c5442e5ce34897629d1fee83b08e5998f9383b0252db1cea72d20ce
z190fdd811bf92d0008b86c11e8947f0c0e62cefb65253e726a68ca14fe71cfa6b67ecba351ddfd
zbe1376d7de28ff354a86a00d19e6fe917b825ced8e7100ed1fa7788cb1e51d9744d41f6e085bbf
zcc45f1a343cb4d6bc2559b1cd35f26026d10039e8b9e1d14400b02cdeb2191df07d3677c8aae5b
ze4d0a240304ddeeb3104bafb6de74f67530266e2f38af583f91a7277fbad875c9b7d767239a755
z40074759d7467e940b50ab6050cdc2a807c33d366c527a262e1e0c2dccc29d9681681bd83c5f03
z32d759fe7b557fe2d3f17b3b57e5cc1e7903875f6564c5622982035b9e3233fc3d4be19a366935
z0007db01680a0bdc1141d27903c5dd38856156be37b177f71e5d26a84e0e2fc4161c2cb7b4376c
za4965e8ae6aa29177cf1f288875165642dd5b6c0453a79cc6bc6f0eb9a1d42bebd50cedfcd261c
z25a28fac4439642b1f48f4facaf526dfdfe137e1657ea84a05caf7f931a8407e53a5282b4f4f14
z2ac4fd8ad7bbc455cf13b3433f96101ef9d4db1326c047e0139b45cfbd5d796b46cf65e79e1ef6
za221e98a2e5cc3f244ba5bd50b94789ebedb4504a324b61f637e082e60a1615db34d83c1a0f6fc
z603f27e15f829d828ebd03a230718b816a17877ac1a576a91e75fadc3f8a1ff5ba8889f955e8ea
z3b9f0e489b6762a204e7221ec37121e8c5f24f36b49f50b023df7efecf72259928717b74987c6e
z05daea0d791615edba7a02fd593e4a59beb0edddd8fc079380220f136f39cd25b43753258e7f30
zb1733d27f3a04a8d73d67bfb3f233e22c2df0181d99ce63b675f26881c32b8d93c886f56acd1c9
z44fd58f5e151d96b3db5966f24c3ddd88c5340923ae47bf329c60f6c9658dc40b0a84455dea681
z82ba6bd6956fb594485d8cab3a45cb7fd69fbb387954c78c02e9c38b916dece701347692c87700
z7310e193ed44f8cc80e513c4e87c0231bf076c1f15c0d25ff4978cfe4d837b161ee3b4688f593d
z55f5ae19b02938b8d8c374e433239abdec2b4932635e5800a0a8893c86fccf11cacd6d1d9b6963
z36be7d625d66ab43a7dd874e443454350e8427a62d9e69c0fdfda16ae1ec3bd96d1fdabdf48d45
za0e64d56f37e694cd2809ab4d8bf63d88661ca894e8e1eb42641532e710b6d8a78014ce2588bab
z8a4297d756dd396ebaa32403daba0ec00bdc89b6fb087ee3103c8637a918363e0b99885231f5ad
ze992cc2a1aabe58b4ca189cb927983e7778812d28be5e1fde20b388ca696d0145aeed37cb5ca6b
zb4aaddb3a828004026ae194389415b3b3f453e7a461f728f354bd4840459e59c9660b6e7811e01
z4b53f8d3fdda1e395eaf2bff0b0789d0a0ce1b382ec0b93187a2af40bee743e1cd1d0ddee70210
z1b0c38bf0b52c640f745398a36bf0d3ea5ecf984588677a53f64871be48c3e86fe5c69dc72102f
za2b2504d41dc2c64d3f49330c4b2dbd490154acd6aac384b36df5c87c6827ace12c81b8ccc497f
zb19374e00d81b9fcd3d1fc82e06ef4255bf864e34bf1664cdef2c10b3d03f94b9acff82012a80b
z29ade42eb08576ca67b673cf7e2b316cc6d4da691b0c1577fb7e7d863d7602c1804a7f3a37e8f0
z5154641949e4341b805b8898c18dca6a0d4fd1757d22eec7e2785e158b0da2a036b456e019b4d0
zab1d520ac9c7619bf7f3b38a7033fd277490483c746c6ccd602320f8d27210ed126ecb569d2742
z945005a886922781452d21c5f1e816d9afa98ce502c1fc5d9c96ad21794ecc98a05e97e9279503
z5928ef8ab06a17e25c9df3a1f452499c3611c4cc3fb68522cbd9e96792042fdc6873a6fc8cb395
zd37c546e972008db10ef27f35ab575332854610cc79ef88d4ba3d0a616d3be386882c01a0c2e24
zf2a2c91fc58167d98b04c237116bcdc02468bf93f2878f4e2892a0f0eb5c41f039885cd70bf5ac
zd17a13847743df8d5c93ce46ba6703c8f921970bce6c5aa057cfd46d4f973602e72bf571c3fbb0
z224f2d71a84da466f71b084b9b3969f945b78d750eecb6d2755d50d82bad0192af3493f4c5af2d
z68a17021a7590f4a0b2ff4e503da289afefff654f42d1ef01f2d348d9f2326d4705fa75806add0
z748635511a81433b4f6b1f4338364c98e605c5417148f184d17c09bb01c22f4afe39021c0d9620
zb1fe5af44475baed6bdc95fefe907b4bcb0a58956a31d7427a257c9143cb14137a997d02727ad1
zdd620a2ad28efd5f41a5f9d67665fb8bb069c883b6266d874e98611e32e6e304dd2a883e4eb4f7
zcc02a046ff9122cbd4dce66ef6cdcc32ebcaff4d15c96f036403a4af4726a5b847192a70fd5884
zcfbff8c4a6f81ac75eb13897ada3aa7543ba670145836e54bdb9ccdcb89540706efd8aa4365309
z330dfd6072375c81de22fa76f2b5582b4eb10b4b932821b4f1fe543bb5e33fc8cbed7cdaa78ac5
zc75a8294d1c68a39002b3df65bf4d1dcf1a87a16a990cf6926c7980411611013e665bb52ec14ab
z6e92169df635f7c0d572966bbc9417143d728f792e8840bbe163f333d1c995e14efbd429f6d7fb
zb501e909c30c62894aa296f83fe78ceafa39f8d9dfbf1bfe11aa649fcca7619cdcbcdab9f7f530
z01b912711418b9d02c6620a77e4100d1510147bad8898bf87455cf3583d6ee8e025314b6b9f61b
zedda5d2bb9dfc826a74ec1064ffd09625bff3c5434f8a6c8b051196d024372a63b80f34225c11b
z6b636ee7f0e753840596dd8fb8c8a0a4eca2ce49ad63c283e8ccef43af34fa77ef3d1627dbd23d
z5d85b40e4bc6ff4be01d099e0bb304a52ea60de4e39794ed51d2ed8d847832922dd9cc191f9393
z3406b9b355c209fc81df4f0ec7e0a81c2bbb6e87365b870f8fff469ae89e7cf2a2ebf4f5ecd66c
z31b49b8d900ad96e3bc5438f4893ea0f7c410054750eabdcd6c531e6dcaca939a02f838343c62a
z32bfdd08981baec66613b7c75f619c79864293a6c95c0c80b5cd9468eb43d4e51c1a8451673676
zf39e7f520965b5830f572c4d61682cfa49c95374e3b3f78a4871a9417231106c6c0bbbce005c78
z071870b9d43b87ab1275e356abeafbdd0534062bbc6e6f93f59944f774bb2fb53bbef15d939ba6
zeb0f2e9502d94f23f3781c9a1d0d4f789cfb33ceb79d90204586e32f49c5d88c901797047c3eb2
z3453f2162a899fc56f36268a89e498c4a818605243cafe3e31388f58dbc24c0c10f5521be7e5ed
z7ce37fb25382355c1ee1653da75bace6c6c24a1348b8da4ac3174e2b004e97883ade8142d3b130
z33a3078d5a654acbeddd662f8fb0225e6b222a4baebd4e860d7e1c8dfbc8deafd3ed7b5657f3d7
z3565524a7184dab393ac45a3c479232aef9694b2a175ea864e5ab534feb65d25fe6839b65aa97f
zd9d1739973724944c682497ed169eefbdae6a7885ebcfab7fdbb733598a02e8a83dd58394ce03a
z7af488b4a07939dede7fbb5a1f90f5881a675c685219f2b58b680f085ea12dee5b94ed5b125c61
z92cb25fa38a7e5f780d668509af5df20e8d8ddfd3c99aba8554ea868c5f704e77f21559c10a7aa
zfd3e6e56edd1047839c90bbf1eb169ad3c684f89b6072fa1aa4bfe599b21fb9bb19444d856b08a
z3749cf71a39667daa8bb19d89c42af48a61e710348be1c2085865add0d40b0388b56c1091b6e88
z7322562d03dbb95f9fd24dcab81623063112739cbf044e3e7a7875cb1b9002e2c6b9f13e548ae9
z1a36c9a970b8166401937961b2659d0de368970561023a45f6aa3dae6223c6bc0a6dcf8a471121
z2f1be1f966d7a8750804ca92f3d86bb857389e81a6cfe2ab012003c1929a5cba243236a37650df
z4aa6dc96da28af635b9f08973d17ce3a9efe5c50b7d1d867f8000b5552341f210d1f07c6bcc29b
z68a043cd48e461ffcb917a95d95466f796438096e0839c07de35a0678dd3e0ef783f2ca6e7f61a
z842eb2ea99e12e7795c92f3e0ed184ce754660460f1c9805aefd15ccccfdde3ab5f9d1a8543a04
z8753592566f14e203eb45f93625581373b0f36dc99d938e0aead95b687456288d776e6f98003ed
z9e88bbea7d40387363ca9d9c66e9c7bd60b5fb1605add5cb03947ab0d7360c5f3b208224482ad9
z49654ab94cdbc176d46ce92d5ea88f824527f0c8e6ff752ec487f45ccd8cf5717af6af9268b7fb
z1d2cfaa1d8cd5bc42914258d159d98af45425b8bfd1c1923aef6a090a6b3df236ed9c6c119b331
z193a5617ef1cfd32a211aabb3c96672919c812aee82d53c6fb72d464ee252cea52c76af86840f8
z07a04de892d15db8e703f610ef450ab201334e16899419df3b03ab61b64dab9637c550c372b95c
zaf6bad8aa5f0175862e577fc3a4d56ac1f86dfdfeda8a889b2308ab68ce4120106533193d45c4e
z7e074a0f59bdebadf065fdcbd99087da063bd575283a69dc6f0dd77854e4d534c862b87356c6f4
zf32d2eade131704c3d372f52529fb4c54376ed3e9193fee69a82aeb0faba3465ff10c5d9233351
z53a2c031fa571a2e7e468e32e34792aa6df1d50226135d8460bc08cd79882a46261f7c54ef2153
z34e9b9f174fde5af5404c3cdd5caf48942475e6ff5feeb52fc2209e59f71a9cbcf819fcf7aea5a
z9b42af0e9c389438c8cf2dc394e80bb24c82d3573d066793ba8dc9043f9159ef3c8fd66a5bcd35
zaad70cd0e21bc54e0d271535d55ade6f2d90d979c5a86e22692c3adb9d6a144c802880c4955edc
z54ee5284118004cbcd3a6dfe28eda9b91f76746aeae3a22310442d3cd093accba4db1aac5db08e
z1bac1ded08eb14f11baad820f77e188f541f18db8e8fa492ae6c35edb5f31ba4c574ab7e1589c2
zeacff359432867ad7533c823b682b196ce8a175aa0523f0163f29de36f5c0dfe96ce8d0f6acb8d
ze34c2d2be7122c24ac1a98121c833d853c609d42039ed149602e0e09858530f2a7929bc329b09d
z826393101e69f7025f0a891ea34ee2bfa7805344ce9c6de46bb499b20bce97890b202c7b509ec2
zdf1f2ac209f2b6f2b1db3d2da024120f4c91bc8a83259e96d63fc5796710454ac78b5a930499f6
zcf3f1d87638a9654be20ee4cf8cb021db4cdfaeb3aa506d402018c8c6b66bddc36ae3b3599f9f3
z89d44742780a414cea104636e425021592a266a9281ee8401ffe81aa21ee8a1d0f7ab46909a52c
z9ae36fb92392a20cb5cf1533c2a971b07530c070503b1cd64b115d29f981ba68ab411b0663fadb
z3d31083e77dd610d239c754914a993bec675d4d292cef46f4f6bfb02216ec47546e8c4c9a64b90
z291a2deec638126c3014c90c5b9dfe1332483cb565d5f2826789b2bdb5a50f8378a85516b1d7e2
z6d2944a2064972624bda922ddf8b5ba2fb2e7e13d6c1a63a31dcf075d26a32dd939db5e25f87cf
zeb855733501d727a4bf0a989d93ca9502978256582c8579223df8b89ede1726135bd10be4db23d
z8f6fe5ff877f51fd75c6b3daa27b42af2c1b74775ec0c83b96808bf8e3376ad4c3967e3733a7b0
z997fd0676fcc9dec579f8367aefe76122aa9964071b8b1a0ebadf8ced62364d50959eec8577219
za0bf108ca6e1771e99ecb0b3a6277f26a9b681c4e185ca45d0f0a2b2d645a6984bcf912f078ae9
z41c6851ca9dd52a195bf4eb5d90087225509d4265166d1695bb875c73afa22beb24302d7239ef9
zd1589766e2ba8808417e381be69dac267fdb8410f51d7f1cf344c1538568ac9ef00b1341c56508
z20a9495506446408c1c746b4fe31676115405abcfccdb57ac9fba33b47047a764cac58d7ec4b8d
ze2c2c77423c031f742117393f1898d56c82a7d2d28b1f3977cfc16a6dbb56660a7cd95c7f0f28b
z76010cfdfcb8d365e86a013102c3c3ead06e07a3415d56a28d21326c657e6bbd6ada51a311588e
zaff694b3e9d1ff426f0fe8878793efd6ad6ce8abff1ae40fadcf79164ec1ec0ffef230b6fed37b
z4b7fd7627cbd94f612ec730dd0026137c13873d555685ffe8d66951ddee783bab2c33bee195e22
z6c677f38dc29c66cfc9d9dbf04026e423d87a3b60a39922b244acec6457fa909062339ebb12bbb
z2fa279f2db9dc8ceb19e60c2a57fb8436eadb9a9547e17fe8ea63e0b160e0b1468ea740cc54713
z5d9e851f541728f6fc71b9142c3d516079e965af89f7a35a38068824bb4f65bb9f01429b5c1522
z9b136017b4114fa8aa062880ceb5b8550c11df528a44970728d21ff0d494151d3fd103a58eb3df
z232ee61e0ecb4eb8df8b26fd5e1ce8db7163da1209f8c9cb40aa023f04b5fc806a29a6ee02fa6b
z29dfdc9ec06fcad3a454a0e4247e34f3fb2fbf0c39bf108f732c9a97caae95c3e75e9ac52a6ed2
za9b578f5a27dabccf429c32dcdccf6e1907ae95a58cec973ee85875cad5538d6ba4fc06ca67eba
z0e3a702f317eacfd12c35cda86cef7697b246bb56ff8d9c3d7800ee2254a71325e013155ca4660
z0bcb228235dd14c1e84ca5eafffdaa9fedb900c9f64db939df38ab63c65213149f8d420bae5dfa
z4aef44fceed430a5277e4774ec0cd9bb23f483b772a58199a2cef4226b8a39250273c0ec4d7842
za48b2b923fe53f711f301e656c6d3ed9246343c470c233a088f245d64a06078a2f397c565e11a0
za1e355579cd2565121eb6d71a69fe7b0f1ea260e4e14fe3563d901f63870b662345213f3729643
zabfdb86a78137221b81171efeae0aa039f5abbaa23e02f110f6a95ec5d8864d207b2c38290300a
z9df1c26ffba36f8b85b8bee660b688e2cd547ea106a4265cf0b3200e6a3e3b48fb0a3094e288fa
z9e497e541e1a633434641740ba6d37e93fd9445182d1b77fbcd36277a885258089b88ebfdf5f78
z318d84917d01aaa3c1be7609998c8d2e0e7ffef34fe70bc50652308d4d11069480c24adc237c1a
z52889858acfb4840bb40c6b76a65b498d40a5923e80b0481f62df1a7f946579d17d84badb2fd2b
z38a40da6c1cc6b6af091d34ba1ba238d09b473b89f31933a5038e7925846e604f7778aa5454f9f
zf778534127a30fbeeae914e7fa17a62a7e9005b628f02c7dd0441c7489443cdc413fb8449a6f42
z561e82e0733a1f70bb067f69d1ea3396f6bb31d3c39856eb3ea9676e29f567a31514dcfe5754ab
z11166eb781ff2e1b7ba9c117ac5956df166157a96aee0d615e0dbe4aca887832de2e0cf27a9de1
z7d34849a4a5507f97d47286780bd2e326e9ae839cfe1674777ff4933cedec8719491caba8c7fc4
z8176e20766b96e832eade10bb0537e5a77ee2313321c911e96da66619df3a8f0341300be99ab9c
zdd0c1a614cbb93da71acaea4ee5e3684b28ed0000e07a8c2def520831021ff6c0d7fe41b5e6f59
z48cd38c902f1e8157d0a57e59382768403e16f5ef6e60ad904974d85f82493118777bb38ce8279
z536a58b977f8c5ad51c4e0ce8ab1dd43b4f44e70471dc8d88411a6de9064ff8636d53279b69907
z507fc45e2da4ac98b17a78022a705d5a547d2f84f0749936df93d69fb143ccf8cf28c8c1f418cd
ze1f1d958eed8d99be6ac3fde3695a3f54b9ca814a8c69a6cfdf2019df98a450b9dbfe8c56d21b9
z5d123233228875de04681b88845d2a4c885d6179d13f8046498f631b93615536ff478c992fe548
z7a0fb014af4ebbf6e4c3bc4be26f21108d00579755838601ed2953d802bafdd640214552f2767d
ze208aa9dd94d7c91736291600f24ba2433f625f1531ad07d1ce914eb1525e68044d4e96e45d8ba
zc4ec8eaeea5a0bdaf74f5fa67a84f4433dfbb961a1bc587f303b4f4e7e6849c139ffc129d1c136
zf4a658d995765e99eea3599443c5d3d2b8bb6ef43c432288f219bab37b25b5d7454d426bfc8a75
z3ff8cebe28a1fc455ebe81df6437342d5507016e33a3c04922b885a54127680130e4901f40c1eb
z642a45a16a91afab45a5b80919eefade3f7200e913ba6376337b7b0c847a17796e0b8b29794145
zc4d7ef5306efd937e56218bad9ece1091b6bf18c6473a13ca1f95d2fee6701867256df3da0b79f
ze447e88022d80008a86ecbb260962a2e9ea697b9c51a474d03a41bc608cb563109e2bb5e2f0671
z36aa423472d79dc2b600d99696e006b236f2b3cfcf58df243686d0d59e1d8086a7c1ab0b6a0cfc
z836aaff44f4cce16be7813651bf843d66d969d1b1926bd801bee5578f027fe48931db8a5bcc6a2
z03a8602374b9cd9fc28a04539d42a378170df8312831adf339fad6fcc77fd51677aab3ea0341a8
z3b1c7174a486ed3527e70cd64ef031dc6ce7f4d88a0fa296d6e570628ffb2c156a84a2bacb09ce
z2648e41a2c93014c5a23cd9341e8b2f8a2fa6822f3fb44aabdb395ea66a772c4fb7e71409d46f0
zd02ba1d7948c20d598ab98f571e569db5a3604d0cf07426a21efd634b3dae6e55c2d49ec4fa167
z7f432a750105ba9e1ffffb9f884d8c5ee14d30b4318b66f7f3a5840d75d902eaa7871129798d01
zabf1d1e65bd32d7d1123d6d62d068951acf5436aa66dbcbbdb53fce2d44eb2850103a018bc5182
z0e06f2c2f6e0e69cd9bfbf29920ed47d5359d223f3d84ceba3b5339da98116f686d471fbbd8e5c
zfc53f5c36df711f2c6e889fc30797b2f88c20140c175a05e2280dd5e4e94f4b29554ed5f1b7314
ze51b2842260f9139b9255a0cbba90d0838efe7ffcec6936c3d75dab14cf0c80535bd1fa324b135
zdb27e3dc73de62ea682bea6d41251f3f97c6bb01afd469b4364b82c29b9d1fcc3f46457986290e
z7431684a50a1e596ecec9cdf231463d8329b665742d87b36f61732d8c5f11e9fb695443c93b94d
zdc00d920a6f750304043383c20995f19d4aea0cca76f486b1586bc5dce7cb31955f243cc823ee4
z0ba74ed62a6682596168b79186d8269ca287c6f5aaa760f16ff4bfc6515fadae1a78974c58ecb1
ze3afc91be09f7841beb80e307a4fb60381415253b77a6b012057fdaec32dc1baf56f3068ffd0ff
z39e88c3400fcb610e4b47eafac0cb9991220facf62ba47a3271392c44b1b20e52bcc18f1d3ac20
z73643fa4238f050bdd9506ea1f2cbc634c0115687b0f488a517df93343fb1d193c8377eff3a451
zfe31760bb351f51aa3568d08f23b25d66f2d6ce855bc8b0e9789ef5c2af05ffda90a2ccf022274
zfe5856fa0ad7d91d9cbf5ec9b7f45b39863e6336f7e31859db672ddc8831da3b20dabf75edde93
z8ce810306114a00f1fd8b4b7580a693d436cf1af6a412d3304c8b6f6c12323ba39b354b2726e10
z5fa29733a0eab64451dc1c1c3debdb7671b9568c8f76244c81e824e96250e77002aabbddfc7231
zac61d6599c0da773ada62c2fd0e930268dfb79125c1324a6cbd7ac89481dfd6b43044d4c7289d6
za0129dff2ae3b534fdbbaebc0fa0cad787446345ccc9529cea3c7484ab705f0c216762d75fface
z0f100498af0b967358f4ecbf29dad107f71b9b1b19f18a847befc31413d4f3ab2a7e7e23bc2beb
z8d53232739632c3b83a7bf4743fafed7963621f88b39dd695afbcd952d9ba26c0a97f0bc52a5c0
z5dac48bd3b2c164eefaa6c7880f742f3c53ccc14e0de294023855f231dd499f5a7952175964e16
z6a2a82494a12c8a933abb06bff72b468afa29159a6b59f4aef41cf00ffbbf9286223f43b2a3f63
zbbb2e58d74acd689aee30cd6be10dcf4ae7cba3e1f8f9fb94f63a9491185a96f288592ed7d6c1d
zbd6e1b33b4222154a0768d849c3938566dacec7193ba9f0d4f8bac0f3cb43e0ef763459f28e5a5
zc1ed458eee1b8fd75d5c74d239a25c889d3d3c84124277aed6c30cce53e50e1c172bfe68433466
zdc8b935b05354dd5258b7a9fd40ae4b55dae6dd784e9e445d99080d7badb6a941b8e20b3b4d0dd
z78a5b395b4b1c83e8c813266354103aadf0a7e21288a21983e77219c1814eb1a93bf8789028079
zc5a445b35e8c613cf72cc8afc7af03847a9e759ea5ade4bcdf7566626b51fe142d429cf85e21fe
zd307ebfd3c2375901331472a37879fce1d01bc977b01a436269d5dc2ae8f5ac63aa7d25c0c6da0
z25b4145933e15f1472429eb679ca134fe5ddaff7c4d24168bca4f795adf96a2e60e38ba6189af2
z1ee2548d6505ce6c6792fa3ede1ac41e161d8b93854c6a859355256c24ce15c68412f8d3a1dcaf
z790501e847f612e8af8fc391797b32f87ad77d2a459ec9ea484251024c87497e4ecdeeb0db3492
zaec18174af3d1f1cae3674a9fd9aebac9625fd2bad7da4a5efa1d9d3a6dff4b12de076d629aff6
zeb9d419180991cbc6bae8808d599ded863af1cbc438eb6b2523261f967c0cb8c8ea2e7c8de390e
z7216aadc6793b79da4d7f223e7f1c9be2498b86f999bb0a78bc946db665cb53bfd96ce688f0ce1
z6b57a197b87f5a3e1a49fec892f7fd52ff10ef27f08be3a78018be510971e83cf7505224ba0259
z2b0339d5cf78475809ccfbfe0e1876aa444da0879540c108163fb16b6642b17aac02b89c9dd5b7
za77e0aef6dc63d93e030a5fa6508531d16f6107d12aa2978f867dbb9fc359134833f2ef71c924c
z4c4648b5b287f62751985c68716b2c3b729cce92d6a75d07e9f1224964f62cfa6812463ff2d69a
z497fed12b12a4a3466be13e50d454af2f7e3619f7973263227c54c6d512deebc9f0a49467e74bc
z04ab64d133e778919dae328be0bedd46ebff3e098aa1ab0be8c48a612339f5d02f0ee168479d49
za4752fe53d485dd68b6e3e13dad4ee378c285c176c480a85656413e3e1e61c7e45a7affdf6a33e
z251af7016cb0a58fd12a3cd715dfb3813aae4075d01a2447b832e449b5ed99c4dca5ce72bbdec2
z1904787aa213b49bce580c6117a62b373225b333d9c8838a4d7a8e2cf82e305f11f52ea6bf955b
zc0b2127f4385af4e0411759c3968398920b5402ae67162fbb7a0b7c253ddb9a459bd8b9a0608d0
z701c0679248916f8bf0838f6cd93f983e561bd0ad3802ae0d3d2e9d49a6e63064ceeac1ac45df0
zc89eabe17bcb00ca60e92dfcbac13787899624bf3e7b31fb5abb698dff33a710ba5757322f4a97
z70962eb55e6b59707e9db4e2fd30d1eb122ec269adcbb59a2c2a50dc2e851de8bd58ce2236461c
zddd99a747a4cae756aa0e6b2c93130e11203042833c9c1933b84d95a5c255fc52eaebdab86add5
z908ad9fd1dc97f4492e043cc6c2f7aa5a2624abeb4787d3eb733796811723e48ce548439d00a02
z8f302b0a03937bc1cee86631d6512748be6fa616f60232fd18970430bc39309cbbb114d89d0efb
za0c3a923b161eb3d0fac7eecb22829bfdae3b50a08f476f981ce86d66b25f105384b2b3a2dc67a
z3f6f73bf2a71411355a07af863225d92d302c448ef527459dbb1738d9fca7dd28ae92a920e3f6b
zc4c12dc75230413ddbe9cfd5d0d8f2e2687335ee3e5dead4f6d4d5c7000809d98f057a249034d6
ze72d2e388c631f28bd780d49cbdcdda3150eb64781486d74dcd0cdcaebc8a41f8d947096292ec7
z5041c34a2c70e98f1e663b030c070da4b50e3a3be6934cedc6f1e1ae20a8784b5db9003ec50f8c
zdfb3902b22d8e644fd9830c7993a38df14cf40340dbfb1de41dcf188d51862cefc85c1a85bbbd5
z0d8494fcb598d9403a6caae10015e0dcadbd5f3292c71bf4135ff0b5ab5ad2ee73469bebe7703d
zd61a87b967cbb492eb6b72e0ec6f190c65c6f4c024ad4d598ba44758182f6ad98080f3c384a695
z18e6996b334bc01409d64ab7ccb9abb5a5661de5525572ce5cc95513d25255fcae30adbe3c67ba
zdca6cb468a277948948be3cea52ca00a4b8da95596c8432ddce94d655ebea929ed28521ee4019f
z116aa9f8433414cf2a0cb2b0540171d96ff66e4ee29b49e5e8a4107e53944219d081bada197a7b
za07529a3506636f126b222ea22c958ba6028d13f4a3f615877524efd62ddf9c52cc44b5310b9a2
ze420188bfd889d1a0080047ab04b654bfe8828f46b5d879569dc526f901eed2d83c3b65651c2eb
zc26d7b73764c577c2065ad90122e4f020bc4f5fb5aad6f024e2937e368ce7eacef8b797a359141
zd9fb2965119d81a684d2096367df8795634a9c1fecf52e1b183b3b6eac34ed8aa819c065fe6d31
z6aac37f1e88fe53ae357689793330aa019b476186e1ccbe7a13d78f6a77f3127240eb48752f7d6
zec5b40f79de49473c2ee46a2584358c955c470023bcec524edb26d7f42f649631b34bdfd927c87
ze53bf727788ce7bce941a25690f3e5b14c66b876130cb92b76223de3eb0eb76f0a7759ed70b9a7
z665ab208ad5890cc8b7d410695297dd53ee255d87563d82652b65778de94f19d9cbbe10b0e9eaa
z4db9624568f6cc745aec59990f13f5077038c9e923b0de5a40a63ccd343bb142876327ce8d2f3f
ze75040013a09bb1eac9077644f891d32e3b850ba99dc13818cc2c98bef7a3d7f47fea346587a8d
zc6a37c237c98db98178d64b5b57456e9e8e4903b72f66bafc6f6e38fdb997f079ce1f3152d1743
z3188dbe2f503034f4f135cc5d0af45ad12655e686440e900b4708b3b746a5d3a21047616ffd3c4
z57d9aaf2b33215667954e1e98eff9da75578f3aad7f9d46e23212d311ecaebae6a78ee256cd598
zd3c2b410c34753867c42e527df0600a80ca37e6129f5c44fdb263a86dbfb72cbdca8b59cf6bf6e
zb575b36170cb680cd837894594ca7bb1626571e28ee6549a12310ec243acc4f274078c239050f0
zc394e2b443ac708537bbff6e510b6e44408c031455f172309c06b276e9eee8e7212fed1f44e807
zebb0580cdb5e18a7d20840b25ad0976bf206b8c376ccb27e14d370f81920b8ac4723c4df5a869c
zfc2c32c9cc542be483a3435ecdc86139045f800b442df524da8283ad0d99d7b71d052909842466
z51c8d323dc019ad81fc9f8fa3875272e9640b48df3370435345d26d03703f9683555f49fe30f4b
z68b2a75df37f36db48da837ee0960a0a41cd832a386559d4bf91fb2464f8f188d797d41417e91a
zcb02ca5bc81aa6ebff8a7b248dc0fc0db8b239f4cef25000e56114e65c2db3b23c3f6b452af533
z9cc8e9d08c3d43b9ec5b884e8bde06107588f1785bb77d75ea20d6277627807566ddeff344aef8
z70958ff886179acf1e636d80e2d90efac772c73b142ca47d063cbec34320881d5695d4f32da8f2
z0a0a1a17387f88e9fd0110ad9d8b0f1a3fd91d2c7f4a57be7b1ff9bcc65d0e18956739f6ca0ea7
zf9fc49159f688717b5bac4defc87f2e5c71740db6d6522891694638576b2beb98d5a9b99170ede
z980a406d94a228fcb4e06506534064ea163dfd4dd34ea37a130c2b0f297b9933add7ea2694365d
z83a6e2b3edc9fb6e5c53f71220d6c65bc1b86b81a23d2dbacee0f8e1f231d6e74e9fcdffd4e94f
z14e71e35c7d9decca5042564334ab5f12992d8885e6858297e84c84dc3b2b3d69d442d490dd2ba
z362949f13d42f63390d22e14ea946d3437187210dafb2eee6998d8888773538988ed5f141a7012
zc106cb12b21f29b03e3ccc52f087c0d05fa26df526bfc19948d90f893c6224a95e2dcda13cd19f
z0c53f0a927a61b4de5c3e03635646acad97ea695d823d8c3e142ddaac9f75baf11a2572311fc91
z27c382271154d0610e51bd313aa63342f448e74bfce940f534d8989acce2610353794428baa7d2
z48a89a1f40e7c928dbe5476b4935919da9c478c9e6a82ab9e42ff37f70be1c7ceab568450445ae
z17ed369145ab2deb686ccdd8445925d83b6904cc10600e14309edb1e846c361b58668f108ac7ef
z6c2862a26be8353c58f1e328d9071d414aa0cdf3e91dbda20dd9b7fd369d17c9ea5f47eb118c40
z688a425c2c8cee0876856cb065261f834ef33a22a4ce3129d94c85515b344ff07c865bf051308f
z74a1bccdfd2441508adaadcda7fc0e55f24bfe924c42d9940cc73a5df23504ec8bb1b20ed75c23
z92c5b623af703a9afb1f5df8d97591e2621d25e58190482fca3574e6f467f1b809c8d63aced30c
za3f9a80c1ca99ce5638bacb92256d6ca039eade7903b7df668d52d9ca4b5c007996438766674fd
zf8f1fe2dfe936d2e887359da18a39ce3f3739957ec02ab69005c24df4d6fd4f28dd25f732bf48e
z4d40a80ce0bd0755ca743a737e5bb0974b8390af3f7c8245eb264d7dc6bd3b10e5bb91a75478fa
z51e94d1b0748339ea2d01b6a55510ded21df4ebdb1c49681c699da53c693f71a9ba5414e093c4b
z8b89f79af3689239ab2a7312f07e7e8fe43a53f1c9bd1da64deffd839d9d62cb31e424b1f8d3b5
z27d60711b52939468cfba577c0dd8190bd5d34068cdb033bade315867d22b3c27a79a862b8dd2f
z69b6edd82762fc586e8a29dbe9a5120fcff9a912c04a289c1bf81f651d28745e89e08ae7e04800
zf9db4de4e38c82d4be33b9db2dee33388c22ac90c941a95493f458e1b8f06aeb91e64475370709
za54c0fbf5c7bc051a21fedda2437c3a306910db710e7273dd8415a3cc7ba6637be49f7a61567ec
z1dd8d1b0da2ac766cc128981ecbe4f8ac58dfc9b5a070ef9f66b65921becefc8f2eb9881ae30d4
z12254802166d81c776d3448c423cfa32091fac3523c1af9f6a408ac26bbbd73827ab547b77ac39
z7858a7c2e02f2bcbaab0e57a4ae2608a839734853a72fe66b8070c322af49ab4b704bc0648fca8
z0ccbe5e4287405bb697beb9dec60e737be6951f7e97af1be58f60e5f66264b499c0d200efcf2bf
z1a7042db966678ff220eb54f0dd60e96a5f6f2574af531a104d28e35a73bd73af91ce520be1df5
zaae16ae966ae9d67043a4b45b3194e1727232d2089bb08be118c95119278b6193ab5d28da00485
z48b42b2aec20b53cc9039618f2b9d2c846267fd0aad6aa32cf2a0650fa154ceaed20b490b992a0
zf029fbae4081b31df491badcf4775f71bd901c7792749368b7be5430479a2630dac7b6241eb9b8
z5bbd8560005d10ee1d2d62bd1e998db024850ae4ca943aa733d618cf2f5178f04dea7e34eb9269
zdffcd5904c3c6242c1239976af0f08ef22538326f4da8825baadf2f46aa7c11b9902ddf5899853
ze4b0c820458ba99891e794731cf22a2a45f3c3fb28e95808bc1dc7b07638049580ed8c24a58237
zc130ac2d9a33a964a1c8955d30ce883574d57e95a538b1247dabf96187f6ffc10be86dc0667e5a
zf3af56e613cc614661fc3a902b7b77d0baa1c57bde59e4997ba0b134f99561e42e6eb04e9be155
zffab905a3fc8c375d82d2bc2e457e1adca04675331140a4892767bd1ed06a86f9e3e1656d8fdb4
z5d34b0a30ea1c4216a178af9ae04098baceb3ef5b82989ee8d925954aa3f0a530f94689ef34c39
z2a740a406304b56b3a1f76e07e82af3fc9fa66cd3d0ad1de521513c441974f3eafb03e7f064c87
z27c7b4bd62af901c015a2e7d82b39223609d55ae40cc1ca8bf4fde19c07e5cec6aacd6becccdfa
zaff03e9f5b1a875ec9b96d100eecf54eab7a61258ad0365d0b00012b6d6c39948db61b8ea79760
za17cc2f00552dddd38559f665d63b995dd73d68bdf454e0d9350098744d10f9836da78230cf892
zb881b81e86528209b68e87bd4eec07fcb03a180bd84aa215917cc55eb84c941d8270a343feee0b
zd8f19a8bb319f29e632785c9a7bb2972ca96a7d7bdc97b11bc4ce4a7121d1978ed84501538774e
z3f6180d858ca074ff7cecfe499cbb810bcfa29f6516f500953705c6346dc8c28b32486bc22b38b
zb2fbd5f0ca440998ca45bd9cdf369800ea24bad498a013ff8d346258c929c766377b9706652d26
z1e57d3c6c24523f4d46ec9458d0a94a7b1dab02726a9ab8033f715fe7545e14afb76ead516ec53
z32d4ad254beb37fa6decef9a9e2da7a3c30694b450f3b2403b184a8ef66da04290ff86a40e368f
z87a9981012b29bf0f3924115f194a4a970dc8e164696dda0f7558488987afb39035f0ac9ff8345
z6166546aafc2c88f27f324b12363d7dc4f0fe74fc4ab8a204848208df9703195ddde0c8d56cc25
z46646c4971c15f4a8f670c39b4eab5356e26a467d6cde4851e162597adab7301f992b9285bd94f
z1eff1b73db985e1c4c4ca4b2fda6f3baa79094209ddaa29233dea97a3364c384c10b376f09fab0
z7013dd6b4a727d7dcddf1c7f06a013229b03a8abe880e65a7444a337a30826dae5a6d6ae140c02
zb19eb0de754258392d15415a66c02381feb2877a52a11843e82904e3e4d6dd8e5ceb74e70d0b93
z69d797163f0f7674e9e4a900667060332626aa91ce8b6dd48fef18d78c9b03927f052ba113fbed
z38e55e65a9bcadea7a56e3b7607f10db4706fbdb6c7fa08bb480cfcc82832a60b4ae86778e2d09
z9e79ac3fe2bc4848ed09121a306d337e76646323e057ecddab60f82e0c7e860de8b4949373e83c
ze20fb8f807c466a2ae0081c279f89fd2a3f7a656005916eeae376154847371613fa09eb844f800
zeee771646652afde2e02d1b10e906190e2b35af5ece4efb72efef15c48d214754a904556c35dd1
z854386b3dd7d84e5737e4962cfc4237307c4f8ab1aff6543eb5c6c1e26ee7834381604e5490e82
z563673ab6df722e264018ed3d7418b5f8d9fef0732ebe1c93d86ec6281235347ad72efed038cf0
z02ac2ea973066001732f7e6b4a81772dd209fa5a5b84fdcf700e2d77913d6b8cb84371a2268412
zde36750aef04231cd2904a8e2450c769df1a40ad5920063c1565e73d6f34438cc4b2f17419798e
z2f1134cbc76be13a9c89ab8db33257e1d650496a1e42b06fe1b15498ee309bebf7ab9f9d8a8fba
z394bc205765f4feb7dd901e5fd4c6e78e64d2b2611956292f6c627337609bc7030769d16b70035
zfcba85d07baa0b35a150774a5214ad37d95c25bff8e0fcc03fbce10dbcc1678b6ae3419eeb0da1
z9e4b46a2c37159debbf68c5e35f2dd3a333d57bd48da616466355d35409ba45d31ee62c8fdadb7
zdbe4f5bacd3d37d063b5bfabd3bcfb0909064870629523bc6e3d8f71a886a0f3712959257c661b
za7205610ba9191762fe2fb168d6e39fb267ad9ba887cd028255800eb31825d64333ea8d70b5b2a
zc0e5bed1e6479fda42fe63511effcd2a7b9f86817e507cde80aae7980b5f0750713c61da6afa77
z18c55bc6ddcfef5ac3de97b86f533a073b2153ffb40dadd4e53e599898e42d3169733f1c6cb8eb
z7f566ab1fd06f6fb17dbbed0c465485b7b6e889a1daadcaca2cd6a9593cf6dd005fd2d9d5db875
zfd3f94c67cd5ee6bab0640384ec13a3278201edbc3bf17d034fabf3865846de6f9927b38460e4d
zcbd70fce86bce43ab22c192931f53fccaef6e58e4137e4db5ffbdad8dc4eaa12a0a1933a26d843
z46044fdfef77ebd73c25a72170135a44989dd0344a7a91b4d5261d1bce1771e93e19eb4d624741
z1929fdcf11eb309026e12afa5652848a5bfa5df11e3d7dacd26f1fcda333600ea98de448d6a4c6
z3209b686d6764564d7974f8f3d3defe44558776b18f521fd6cfc5faa401e1d062f7d6899efe3ae
ze92c5e73239e11790a418b340496992979bebc7b5aa7db0dd23028ac5c825c7d7a3497049a994e
z426de81fc752c8522a331e732249b41ba14f734aad684605da329abc15d319a87331524030aa2f
zeb7cd1d0d77ca49a95ae0ed9b1039dd0d4ced378066c012779d801f01b8bfde18d422d868b6f95
za9d02833f6d74a109a3eb122d96a54b5c8e950ded718e4304e8d638a959e5e30026883f8721177
z8745d4bcba3aeca89b2613cc6a0e5d358d55fdd5824bc88307e9ef31e03bb621f6aacc8e01b990
z013af12ad4b3285ca87afb065329bc4e9b8b82f5b6fe6d2d25d467adcfab7c5b5cf40eea85be18
z6fc9cf229c4ff8fbf29f537baf18020664e39afc1c9b172507cb65377e05651fe1f91f1e2b32cc
z7479af526828acbe1863d41b93279c899298ae20f523a391895ee7c0b3983f5f15544e0ed8aa17
z19cfe2365c53cfe84c9bc0aa24f0695fd51969e830f8dc8e6d92ef8a0b30bbadd24b4ad7eebf7e
z9cb294923b34d7809231de9527269d96bea36ecf020fd0d046b8d7b759af0ad03828b0f68beb1c
zd081f9774b7856d3a1d08336bfb40b18ff82af98ce7399551f6e88cd03bec97ebf0c2cd76903e8
z83197f2ea39ffcded6e2c4f58255dba6ff56bea8ab7f51745aa47afa66664a26ec05f8d94b0ca6
zb8a9e67733ea006d920c7a75b4237c1dde9884941e1b9f38c4d3c17ac7ffcc790b14c227f90490
ze9dd1fe604fcfd251ad6660d5f6d85982aed15f11a72c75dbc5af2917368be8157de100b2ee1d9
z59eed06f22ab03d7470eb20bb43bb9692252767696c7976f464411949081fa7ce46fcda6c8fe94
zef3dd017216fd7f84601074972a17aa1c0fbe556044b5ffbfc6d9ace1228e31d9ef03b344ef34c
z532c61fb2e5470713334ac75d58ba08043663aa7aa70640b443930281924300f79ca7ffd4dd312
za1a0633999f0e6127eb6be1172c3c9d33307994364fdde6e631c4e6b90fadfc9e237cc8b1eedbe
zdb8a84337333da6c018d3558430ca6166a1f27d10892c9ff30690faae0c96238271bc6e5f76be4
z018e4ab475a43dbadde1ad82c483a0f9c9f9cb16ed92aa5b996d1d494cfee6c81a7c37436eb3c7
z13ac03bbbf9a6aff44c9a66250049863b4b86b9ce130aa071486a58907781930d9895ed3b3b35a
z843fd5840ad87aa8ffee6bfbeeb594e4b8cd8ee7b2e9bc8984cdf190cacee33d8c63fdc3831d5c
z66e7ae18cacf94cc568e8ba58fae7c4d6105f179f289d8050f1e875dfa3f59b46b3073550bafd7
z21dc180b48f0b60c6d1bae678a51572a196ea536bb858ebf674d1f7f10dd9406a56ab5f8839ee8
z5a142a3d07081176c818cfd22dccc0b24a1c0104d919c1d360b7c70f2afe67e6c19f9e7b699675
zba27890ccf1b20c03b9e263d7ce3590e5757ca6e5abf9cbd69f120c7478b23f3a87d1f1e7eed2c
zca7b3a228b6e352ca1dc4fcc5c4cd99034ecc267b75096b7336ee4f5370eaa6fcfd9fa5334db7e
zfe0929f01e8972160a61b5abdd402efd4e7a929732a9a14e1fabe0421d30dfd6ea2bd107a5fe7d
zdb20a057e767c2d6bea6829f8a3364c784afc631933e54ba772da4e1d857a2a0ea19db15a0d768
z8191e038e8415768f271008b2e264231258367903eb3183daec111e43c744bb06548601460fdf5
za0ef841aeec2d865dd47ca42c46e24d4c564666145402650f89f1a3ca2186e89384a12fc4a0829
z823f66880dd82d12a27afd631fecda3569677808ba38d17e747ccc9293a52a81be34008030840c
ze4d615b54706c4cc2ef042314d47d758988006db827c7b2a42af79c01292e0d4a4279f12588724
z4ee7868acb1e0e964d79bc3e1108782cf958fe8aa091a15c92a06bb22e5530165fbd583c11f57e
z657eee1fc811915c59ebd7abf9f33836c6ce537803f9edef56e4f0014042359519d601dfee0402
z3457be7941758b6fbcbb7c77c380fd82d24f641648856caf71f74776def66de26209b3d08970a2
z647d3bd4fbdcf76289b4c781b3aeaae09d88c062a115ebf027bc000b18ad87d7c9507244574508
z1bf9d7e02d4a0eee2aedecf622f4d4d3be3553ee54b0f291e777ab04efd08cc78ccca9c4be903e
zb7b39dfbd8afd1e56375de2287a4a0cd20dc6295bab529f0d3edbcde4e9359b11d3e0f92fab683
z16b60a6da2e1f2f76525cbad1ca03585eaf477b4524887482a46f02d0c95540f82c2a7ba8cb948
z88407140e04860649c32272d28c1b3bdfd11b52dfa539a8ab0da4c48cb3709d9cc78bad8ed7168
zc0244f8d2d3c584cb37b44dab3709833640c8de63a57547332ed177ed05df82e4b07dfc1476815
zea01570b1fcb80f710e36e2691229fda537bdf219ccd304cc31aced3d23587c67885dc70ac21b6
za98f0605f1b667056f7db564565e31ca68244802bf75b51a6156c2e89cfaae3ebc26f43bcff9eb
z7bb51a2ca36e9974191af4d9ef0dbb2c25a47baad7924633434f1b2daf3ae1705a1535710fea40
zf5f213bcf1fe43f49a7c287c3b1dbd3b1fea3fe835e18a8991d68386793af0703c66d2857c7465
z52e876de8acabc2551a2eeac6d73e30a1ac2f36f2f80a664a6d5b66ff466ecf7f9693ef3de0dd0
z3b59f28e0d2dd4505eb85fce4141457bbddc9ef206e367af6069c7a923ca582ae5acc7351372a1
z9b56ea6186a409a626c6160ecc21cec3cb75b67bef21e016be92e9a496c370d6862a9cd645a3e6
z3b64993d7033ab1111ac4b3b3e2fe5be8d8b7cb70ebc160234882b6b9ffc5596a939e77dbf121f
z742dcba3723e980553739adee6a37028d756b1f5b937e4f82709b235c9533d5c86f54da433c3a7
zde2bec8452494316681a8ff90dc41be23a14cb073850f607c99a655b0d1a0a2c70c33b6ed27da1
za315cd0cba959ba4c45355ab66c07b6d268c0f987dda9948507a0d07440b8e3ac08880838f7fd1
zac423b12f972b652191029159bfa5928de838c0664ac1256107a5c4fc911af398a17f9228382db
z712f3913db93fc194ce9f8ca25c40d64959cbcac28a7419a36dfb4bd129fd4cb7d43ad51c640e4
z916093abb8d34eea917713eefaa3efe278f0684423de64ecb7c8414ff5982a3dc1f4becb7b3498
z6b4882c710534ba9e16b7617257f9fcf1b607eae0f0c80e5f07f31ca11b09c5d2d4d85a4755f05
z27f93e12b9c852768a42accecb430e4dbaf85e86b793b6102b680aa627782f4a9ed6667f70a64f
z88214bb8f30eef24f7155c29460c0851b7b01194ec02aadbc43db90ee006c0d6eafbb53dfe314b
ze1d21d380d43893d407a8805e4f646c0597b97ce458c9028119c5df7e3978cdc0d3eeff9668ffb
zd152e59cc49513266a4aa2a72c1650497070b16bbe39a7ea48acfd026c1d758ebb4155f151c57d
zba765b941cfff6d2575be2c1dc03e9c03a16b307a2bd5150613a6c4ae3fa0e9e98e9ae70d26953
zc3a4773aeee263e2c59e83a72936a00e9d9bb460988161ae8579b056b592de0f015ff7889c07f6
z543263a1d5e46b4b0dee98ac0b35f3693958a81b36b13a47ac37e508d2df81990d8110af265df5
z9752f8fbc1e519bfca3dbfc177f76d9346518076d169cb1389ddf15bfae153d2196ae86cb20d6f
zc60afa22518984eb616600d8d8a7ed93efdf8bd6d759bb4ff506b10e83fef9a709892261f947a9
zf5a8700f6a868ffd7fe9a29f5e6fe9d9e7e8318673fffdbde2b5537f84d775748264cfb236e460
z9d0dd8cac8a2d7404a6088d17efa6d55acd68d452091120c371fa1da07f47fef9b225733dfc861
z354e7ff4f31105f7ba6274e1857795c9f8c01a54ce7b4ad53ee8cbfb8bdcec997c981c8bfdd211
z56f8b2f984a89d35acc449c4c57ec6eb79ea976df6dc51437ee785f10fb157f4b779829e0e3d75
zee7bf4fa6c9d0324735c56bf23569dfe40ddd3399d3673ce148b5adecf03aac0f48e12774286d9
z2d7803896fed66b9b393816520f377b54fc5c027fcfefc8ca2ff8ccce3cf217513d5ad283f4c3a
za9ae68f1553fb7667f9420d0593f62aad68f5ffbc09e822e5ee67d14c64bd0c76b9f7c7b
`end_protected_0in
`else
`ifdef MODEL_TECH
`include "qvl_gigabit_ethernet_xsbi_link_monitor.mti.svp"
`endif // MODEL_TECH
`endif // encrypted_0in
