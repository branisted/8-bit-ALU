`ifdef encrypted_0in
`protected_0in
ze74c34e226135848fe16db9ffd31815111b6d7fb642c521a3f628cf6da949865580b22efd062a7
ze90adae0e65e66a2c36a587d0a790699161455169ed55a01f2084f11770a774ec4c588039b380f
z6de9c5084882a40b79a175f5c2114b2b6d78b070cb806e1c0aa9258297f4687ab30857016fc53a
za25afc8341302f0c829d94450c399b8ff9b0386c187cb854ee330605b7b59da379b1f26f488e1d
z36e675f0b1336408b3a1ad87d0723054f952fbefc8d5a33eaca6ef5be8f42bc59870a29a5cc9dd
z4fec09ce6e44cac279651402e7e1f590df88ce49ec26ab39f12b4a02855703c6f03b1e85c797d7
za357087d98e5b1f45502e45892e5823d6fa4b762932009620038c05d74efcea7c3fdb38901d620
z36515d0824367e48d1bc182335f158c262d396cada6b0ad58add4f945eee634c2dceadbfb5118e
z14969c29a743830a07124bfa78707f3952b96b0db7af7c9ff36f77137d8c490c4f79328328069e
zd7d5280e4f95742c9841340368b9764f0f80413adb175ecfbdf3c40716abca7b8cef6f7fe92ab9
z6bd2453f1aef7f7899c5365c5c83793cacc7795c269413f6cf0dabad14d40e9285afde8c01a47e
zb61893788ec5060288cabde8fb553f21b02eac61ab0b48ad3d54f4d1d76508b22f0c600861b5ce
zcb30ba708be817b1f50f59c0f6fce449203e7355c1be55b662fef3f92ba58243d81537761af8d6
ze27d7864d2dae99372b2b75bacdc0437a4f7e011d68c3487a89759e3625548fcc920ad06471ee7
z2d701aabf726859343208b0a543c73eeff8406febf277e3babff437ec820fb49d6b78e73bc2353
z884917487d35a6cd06d7d73ccff5f05355122888b886d1b7ae29679db6c9d2d7f218ac9728369e
z0ba3297b105b1781345d5dadc1077db50a0833d4730649f7637b2138ee147e4486fe0551f541b8
z43cb1f566ce4a86a39651786521e6c831c0a7a8984a034633d4209a41890c86668029516983a5a
z2a2918caecb85c3a38d21805a4b7e2da92879621bc299fa7b4555f7e1319c222d5509f48164b83
z9f45f9b9fd8b57ff2290408ba1dbf726ff7b13b8cbfde6de453a22cf49001d87d40be9d1294fea
zf8a4e779c301acca37954995d746a09bd36ae09a4dc137aca70eea5630b84fe037f3a7e8c9379b
z2e8a2bcbd28d3b5e7666c2a32f2ee20f9493a405aba267563cc3e8df277818faa7d622cd4d3769
z3d792e01df7dac144e0f1f792da35ff44da7b5199d4b1095b6e114fab5825bb216054616b1ab74
zbb026db66294329c54d92a71d5e70d2898078f64296784e52c9fb2ade6eecf23abf0f72b4903e5
zfd59834575526346ea56c16fb9ece1a8d53f60caa5b22c6bdf6369e1c0e5eb2ad9e04d02bf4eda
zc35bca74f64fc5edc71a8cf414582a6cb5ae5a15758c7cfd92c329c605df202899737b2aecd40b
z340393e62425c83397acf9abddf0ceb297283f595411bac67ee4652b7a0163b00d18f6820ae7e7
zce80b17d1b404abe49da62e124563f1100b061c8a738fc7db387c0d6cf41af46757e8c661841cd
z79f69f5af85c485edd5c4c16f6a1de8ba6f043349c173f8ec86ad2d0d069eaeeb1ab8143682bde
zc40ace2f4fb4cf66a28be7088e65a99e38751e6b4df85f4da0d79350737893a7e6079dc3a73401
z3445a8f010ec57f2e095062232fbeda1d47c5af597bc327711141704b4e0092e69b81e5a3fc464
zaf8d4474e55c25ab7da61a857a1c654823489d9e357c1e6690537777c83552b3f382ae49db634f
zaa90fa1c3f483502f190274544744f9ddc32e78ca807f909103a0281960c299e06b6fdb226832c
z4563b5d88f9d33120ce311f4ea503fd187a8db1011d9ddc4cefe5ac0f191144f32cb3fabcb112a
z1f63b80e44ed44acf9df051f5ba99bd16303553cab8f3e4f5c8617cfbb1f17d2125a41fd6614a8
zeb6c292e082201072a18d57f102ebefc0955549cbb59a389a21fe07f9939f9e50ffb432dd2fba6
z10988f60aa06acdd5651a84e0118e4c0d7cc1415ae477fda0e19b53dd5f615030bf36b846f9a6e
zb4f5ae08a2b8e62a814abcca7f02453f6ec32337b875ef93a13714583dad81a965a200378f3566
z6a28f86ee98f8226c3fa5b7f85cf2920385350842823866e264aaa4fa3d03fc56024cb10dc0458
zba9b1cf90144f2d2c2e3f53d16eb36ed502d0c297cb9cbf0a398907cbbaec0f824e2b7278d4116
zf9d766f2654f73c43f4eb810b3be37c606fa3f5944f5d0169c4356c0a929c4edf99f8b0953666d
z00b416b0a7a2fd6f4668d7d58da351f450c613469cfcc44f6687d845c2930f12d64602cf14d1e7
z013e463462830a8e345898a5cde895425b5098073d9d6a6e5c5fdba0ca35bea1db1ccd6dae3e1f
ze379f7d67b663e055057b89e0ccca5c59aeefaccbe0dcdf4366fdcd3dfc2139e5e9f69547092ae
zd1568584d7af0f61353f53452e262fce6edc0d2beab917cfdb675546211ddc22a2e89e6951245f
z84e9a1afa9271a8f443719e5495c2d014e076c1354df50924a90ddb968526b75a40b99f2f88f6c
z336887389cf3b0011e8616047e4ec51e28651d9b05d2eb30c155ef0b728294f8227b6b4d2b57b2
zfa1ec37aac9af028e2f281417ebbf32237696e9dcc793efcf959a573726f37431acb1050456241
zb1b065805299cac122dc3198bd5ba38fd54cce23cc2e6e65aa1059a3fddf1bdbf9c0dc543f0c05
zee07243fea7bfca3a2ba582ca3ce4ae097d454e4e0359d8094785af83717f797cf4079a6b603db
z99195c7f9ebf37b0ea1264bfa317b069a2aa6cdfa93d4fe6f1b6c1cebdc5cc298bca438aafb5ce
z6b953d0f6d175246d9ff697d56c1205ce821fd33899984c61957b70a7d634f67af7bbe37c3271d
z9cae08a7fb3b7026d6998d36f61816b0901678f0cb9db760ee65ed75f06e8ee58c4777532b8738
z40b566e7c020c64567e961469c37a09e12ecd4f9595ac471040757a097fa777348a0e8754a6df3
z767786941b955b5e853c03094c0b12e38e69ee590d4ddf0b6a649d59fb34534633e8f45cb7df05
z38d6ce75ae23e63b5c222f5c8a692dd5ed1580c5a607561aa988c6333c4f82e3e3fd111783b03b
z75745093b5a75fe0a7038207590234e6d036c4b20433d30197c63d25617c7a1786cb835349c091
z0faa74da192bb744600691e2c71814b6066e2d2e6adc3da1561c8f6824800652bddc13fb4125c4
z25d5cbbe8ad68af64aecd6eeda68e229d44ffa5e1b8ee9dedef5c3171525267e0f483d3ca6de32
z7047ca305f6f61b58e65f0171d94a5d86ea5c21722bf24b86060d6a0dfec8b811f8bec44966050
z2794521cb6a493aca7900bc11a72e68329e5a1a45a7d090476d6742ca20c5ae53482d2675d5dae
z3598f8bc16a187ded87bdca87d38a020c35135277a7f007927ac4ac4e3929d121f8337479ee180
z492afa3e6e242cbbe765358ff02131421a6d1dc227c4b4b85ab661c2cc684652045ec5fd368468
z41aff27e5a2a54b03bcd08275614a8676551854c79cf490b693cb968a435219164734d53ebf349
z9e2c4dec7baa27f89d0f711f986e1ae2635a15e0723cf7bf2f1c1b6d45f6952e4c69022bdc2d8d
z9ff3149f93cc6f7c5a05248a7a0cb2285f65f37781e0e00a7a8b652564dfe68a2a305d05783fe8
ze6eddb015c2c662d61f31d97a32d6569981565c40f1afc5608b118838d81058fa4b2bd3a28a536
zf9e23307b36e05546ccc834638c8114892b24ecd4b7eb5f2950184ed891f744d5c2b72c822a402
z97ccafec506a84ec296085948912c70a2be6f55ec0d76a36452344f69914b4c0e50afe1613a9d6
z2838d721cc2e87101f2f5be840b974f44729ae5e6d130b5599237f5706ceeaf0ba2808a79b248a
zf63d49275c66a3a90ac98714d8c7267b71e16e27d6fca196c94ca9b31bb75cd21e5c6af1f5db64
z755ac43a0f759c84a34ce12c0915a6b0baff1370c95668b2075e0326d9620b7a6c051a310828b6
zcffa6732df7c1f087d2de86337e29cf1bedf9bd33424993c1f43ede40be2efeb1d941426497e64
zc95e297e3784405975313ea1a95cb9b63c3dcbce0f2a238760b96aeaae7398ccefc90dc6317c4e
z4c12bfa247e37fb5c08a6896e0d7a4612fdfd26400db8095a1044cb68b15c6dbf447ff2bfe9d5e
z35d4be922bce9bb428230ecad8b4a47cf2ddc91864c10ccfce612391a0f4d65821a62b28633f13
z8759ca424f7d5c10b17403dfd245e97bf4858d0f35b9cbfbb1f73b24369c4447195feb3b1edb36
z6aa76e56dc9ad5882e7a89f7c3140d8d2d376c7526b897781c422bfb64eacff4292c94f3c32b34
ze53f026d831723c35ee5c5be7ffc1ed578dcc93a8e9a47628789ab7e95f81db9a12921899b3d0d
z21e3f54ea4907f01471ef5662386f957852f18691ca6cb4563e48728c9c0260ab9151bde4e961f
ze692c516694a8604f5709a40d9c2defcc589c201432681b9e8fba0c9fbc0da19a43947fed01144
z6ceeae9ddfb3695da863c6cf692ed96d07dfcada42922017bb12ba209801ad6dd94f212a9a3976
z162ac310c9f1b3d3a7dc8563ffaa78e4f4fe577d1d8bc562cf6f2c201105114199177c6f4fcdff
zf43ff4fda34236bde7c08ecc8fd2544489d811fd507113a1e0a838a24aaaae14ad2aeea564c28a
zf0bf6af315481177c5119ef6716433996b5889ae96917ee8d0ba77f147a7dad81f1936cdc51357
zffeaaf3307f48ef7c6d5f8602770f40c9ed6f367051584eb7a6c62c8bd104b03efb179c0daaad1
z153407be59890af72421af0d51a3909e66a3525953d288904adf9b42a501fac6678e11c497f1aa
zd95c258f97bfed240f5229ab6a0a3de0f48413b2ae3e93e4ed4a70f099b134b900dd2807eec0e7
z0c7c72044909a9ec02624fd329d98de30170db87e837fb30d84e3b073807a0379140aca41ba3ac
z72ee6683ef29bf4450d04e3c52fe036bf4b4942f179bcfd536bad17ff4a294e02d648236ab6c79
ze442a05164f6a62a260835d46771c8fc6efd4b9e4f87c2ac08cf8a9b5fb9352678c193dcc77257
zcc76066e82b334bee5b587c0ff3419afc8ca3948955c9ef1fdc9db8c3f9dc0c12845cc9f360c13
ze793ec78d49a7eec32dc53fb9a5d8f826222ac4abee9e31393604ef134ba5f48a4c5336df69738
za40a393ed6d3d9346ae4072d9cfbc4b16f6ea145b18c4128fc4f2673c7da7a19fb91ab7f1c22f0
z05e92aa0b41340f3b3d96de63859e7211806178514e0756756642f3a73756a6b42173fa3cc96e2
z23179e5c61d9f821017f553caa2d904b90140ae250d08b462b392bb31a87545a3652dcf4bae7ab
z2ad1ba992e30ec7f34bd57026fb4917efcdd745e0dd4ec71a6806a1419e75b0b14336059191b36
z49afdd9c99b2b9da439fe7e609b4f493d9f6738e71b3b5a68c5f6a6125263d20b7e6813674a49a
z80ad34d558ef41fafbe36807de6835935d53e1a2a5f31b7db13c43a6af669475994803166387c4
zfd9e5db7833fd8695af2876fea932aa065ba1150a48c02a07036ea1242f0a945f682700d7c28f6
zdf163cc82d0f3d60480a6c256c0a66b3eb8bd3219705de73530dec0f2cce730c7c80a5e737f171
z589b5181b701fa470baecbeb90343245d79d7e25a65ab40664fbc550131443ab7f5d16f5b84611
z65b26aee5df8598f46daacef1f91c0bd3689756ad1a7d0f30cc8ab480c8c8561d2e70fa59fe10d
z2520546a66043aa32c71fb62938548505d90fc20b343f7a080ddaa9c07f13e2901afcfd1757072
z849a5e054d05ef739db3d4932527280db360a93307d1239733bdd6175fb163366eb5d328fc159a
z488c7d721909a08cc66c28c69e87dab9ef93c1cc36c8dd7d92ff7ee2d94c89961356347673a0d9
z20bd1655fa5ffa78e94b41d257068c24cdafa36edf6990bba600e46b703ca6e7f6401998064d4c
zed00bc6f2097b01c3eb1becd8ba191c381e710b9a5bfec24705626ad94ade789c499506029ecd4
ze609579447b6ec21bd5358ac70450714327f2ea897c5c690b576f03b147c71d42d883b5c9c4b94
z1c19c625e6a1d305ed2d0d022ccd4d3316437996946d385a5cebd505cbb06400f20a349e6eae96
z2316bd031a57a6fb9dd2542d34413edf3d419f3b2cf14ad6209b9b1cbbfe6a549f3d16b456077b
z755ea5662bc367639519167ed2961d5d8ad4843b5fcc0ed400661ca1e639e49e101fc9d22175a5
z829b70eb8efa29001f3fe9fa2102322b175a5e161bec7126abbb6848b496c4b63d5363980ca34a
z1160e15013c09e6bd5c3f65ca2e5582e6f0668022b4e104fe02bdcf415fb73264cdd5eb7719cfd
z24c6b3fbf51da286d5b593b763a8699c6a57a907d115c9064ff81442edf5914c7496029b19e828
zadcbef9618c679531f2163990abe6e5d2da80ae9a7e1480c0b98c00af0ad796a1598c3f78fb7ef
ze43e2062d2aef7b731e7a4574d9b6f5995b92b68883cf9973bdb8d2c6cda082005393aa389f3b8
zee1320af8a45c39b516547559199ec4eb5dbd9b20389caf0acc4319398659b4465d833e6e6eb53
z84e83540497a835c776e75d1c5f1a680411e06618da8ba1a1fa0c39c78463c5ba6f9cf51c74b04
zf8ae667c03c1d15160a636cbf5e61572f8b07b874509bb2c01fdfee61b525eb3fda1472ff277a4
z782969cd48da0b614b8e1a86fdc2fc5f9f7b6f8dcf4e6d02eece6972293460ed9789a3eacdeac8
z931ee027c7d9baa14066beeddda1246df49ebd640b1b8f5577cc05fda55d72c45b44b35695f9b9
z01c1fe9cee3e4f7e4212833ff7b6d34d50b5a728cd9f57914f0f3a8a59648bb2526e1bfe019853
za4c16db8b495cb5793cf6b1d6194b2c5334000d962946c4484b073b55b2951e5c4b20b1b8cecc7
z2a842fd971abd84e88cbf409195243c10bb7f7d456063c3f5c41616660426bae481d31322dc048
z19d6cde3f81221d28e2270e25b48806d7211960ffbc363686a3f7a0b37120438e09c650d84439a
z20bebc1d27e3d1cc713fae990935a17dbd31509a4ca9721c6e803a550b28a1a64df83cf5b8246d
z7efa9096acff78db85cc549eb8bec29ec4108de9ebf1eebe6485a80e5d88bcb387e2094bb0b878
z21fb80f81d02245a605e4180424d3c0c21275fa3b2781fef7f1af41119058a4ca5c8b772ef3ac4
z5a38a7efa02f37c85ad49cac7f1f633702981393cf532bf09dc6a37541cfa886cef166d6301fc2
z0b008c90fc27e5e9c1c6e5c0ce857d6e287fd15d3e352eefd5e5037089d83ebc5fb67ed381d5a9
z00e2f75e1b33e9f3183aa81a27a4767d4ae772045800ba71c80cfdf5976e47ba4432c8b086120a
z0eb27f70f3cfa964ab63bbf8132754a5deec8baf744cd57ee08a99c33ad30fceb1b6316b720681
zeed90072ce4ce5b5b290714339a56f50615bf433dd3a64697000c644ba101ccdfd816709610533
z7f29bbf11ff8235f3defe8d1adc34e7dc95325f7408dc241ece66c165a7e036175ca8022cc9b24
za658f293de90d646c7d5c05824692c3d16a603e862ebaaf36f2272269439eb99408186482dc11f
z27460ab92c8c55f3acbb5b10d889c592acc5d1945b1f7fcba9e6c375d84ad4cb819f2a002d3191
z69b9332df1b3c402d01872c54910039a04ba377d703ffaa9a516d231d23570d8bc9c23a0f1bbe3
zf0bf85062a40eb5c0bbed797b349893a7c20359b5270d8a7c7d8e4096a432e834bfdb5135e5d5f
zba4491a231bad6947a7361231d300894a9dccbee20673592fa1e57bfaf8463c6db944d4b75968d
z070509067e489e1301e67351cc4c13adb64fdafec5dd8cc17158282056fc59277d330a935cb0c9
zd11192ad86bbf55d1f6d7263a8d953abb1d876e8e5013df10f14d6c49d7831a7af02e899c060d8
zd06bc9468d81b7605bdbd16a0265fd05fd441cc5f119ef73702ad18274e1fd7991c567300f9179
za1f07b448ed2fa559de890d08548190a421ef0949c0173595d4f4be08f87abc175943f8dc47017
z647efbe72876fde988b25ffcb723eb8e89a275bb7b6c9ac6c1c56a3c16ab534df81d0b3e2be24f
z4b5ee6e2f16624c7aab9d37f22f25e72d04958335765fee4b184ee9b11b60d3b8f1cab7e61e703
z9c0ddebe14ff0bfc6151302249f9e194fe72b655991214a222a4577d7db397b1f0c1108c724172
z51a4892cc86249ce885eb2313f4bd61f69a875eb33c7d05588f683afb81867c491acfd897a8ad6
zdfb450907a69713b5f8fd3b4dbf36909e9abc1475590fcaa992ee40850f67d3b4b8f8b78c39b1f
z8b15749ed1756afc6a12697b8351e4cc9d43eebfcf2e769864c8fc6079f1c43394a1005b76b23f
zd13f47ced5b2d1bf084df916f0286e2d1ae1ecf51b0d20b06228d7e760ae9ff2a925f441e6c16d
z6c9028df3761064dede48943b48fb69e89bcf77cd03db9c70d189c4b0f57404357f37d3b720555
zfc0e613e4dda895240908701365c3d99161fd8ef0824f8e5e2793737b353b4b35c0899c212ed20
z0fc7611453daf5cc650aa5dfff1d9369597a321abb478982a65a4aeff3aee5bee650e0383a0658
z8a74d78321c03f4214b2fd7daf53c1e223fb6508c80df6aa11a55644a20a62ff0356872e0faa28
z013d5d305db1d68ce9bdc67d9341533ce399cd2ceac5c4d38b2216bd8b179dd909661a3bd8dfef
zc3bc45e4484df7622b9e7609cb2e485cc6371462063e7f6bdc4dc3f390003645957696c055c206
z5185b21598f7413f93967dd436b8a978d749dcbace912af8ed5dec66b5fc91c2f3823efe0e0f67
z31728ee96276ae4b0cbc5bab5a39d9b4322f5e0d4c29bea1cacfbc9a646001538ab3b828ebf598
z035d7e652134d8aa1de2972958b0bee94946fae66d4f66efc05349cb9f4c4077174895970253a4
z6c1d4dc68e779ee806e6709db36426b38deff10434712462214170f5584b99561415a5080d632e
z84b6a26e0cfdeaf9bc3da117d623460e528808cad71ff1b69a9047b353162c54596c68bd39141d
ze8cb35ded49288505777f56a30e1e4071cabba788ce68e98dfc62ddbdddc33ec5677fedf9bd44f
z47512c16b04356b95ac10e1ce7c2674a05489ca01a4923e063f41793a34046011a7ec311c83d7e
z8edbeec53c878dce7fac6f49ed4aa44f24ed575f7b98bdaa3fa95050129c84e994e3d83b0349ec
zcc6f9c35315f989509ad3fc4639462d33f307ef778be7f4eed4577e1e97e14806397b3a6708fa0
z7f5170bf17f3f3ed5bbea2e65e3fe07b10571b3ca6a1a6130aed9549198f61aba3b42c56ffbece
ze5d22f2243468f26cf4054bf15d0916674fd75105f8e93eb158abb02924da390a5a1112acffd4d
zd2a580a4e3ffa5f31aa6cfd2706ec539a9b33961678e32c3e5627fd2613d323cc2cf2364656959
z09a2c493442830a8fe2cbf372b053373533edd7c8bb9e4c06f9f51ab28269a5cbce3d71a283e09
z7a53d3936fe4d14f087432a9eaab6fd6bfc13db934c8d2fae0dd1acc97a01ad8438844077aac5a
z8f2571f7b8e79520204fe292b663939cd19254686a6bd7e4cbcee3bf0e96a0984af4dee3a47848
zc7c6c799c9835484f7f322918395d64f615206943aac4c90ef630a511c2ed5cd861ed7f6f618b6
z3fd3f3f0dcaadb10e6a44086fa1ea3b7e2ac92013015078cfdae98091f455f59119b39eccc9112
zdbbd8f6b7eb05f09fec6fba9ea2e058c562e161c3895fdff22affdb965bc2af118096e439ceeac
z650d45063c9680293b365fd1f6e62e382e2535aa1c3d72eb66cd3672e2e2e0d9822272542520fb
z732c00199ba35f943e7e7b4b1e87329c2544d7deb341ea1cad54c440073373347c466e39f693d6
zabf7c56e99fe190a3ba684b32dfa6e6c1f1a0221851f0eb39cf82fa2a8f827c363ab3ee5d5ea03
z838cc40aa2123a5fd545b7bbca253e209e297a4727a07660c285e73a7b1f6c24948be452f220a7
z9749cea375371f5bda3dead875ad493f616dd026fabb874f1f9360759f5719baae4f00ab8daea5
zeb3f58d3f5a7e86c77e15920c58dfd837afa9e05b0bc4cc8f8b098773a8d4d65aa362d64bc3034
z6ae44137e3a19848b44a5ee9306ef8d7d0dddfaa16b75b03d5c1d4f5acb3434ba6521d7c0b2a63
zba523552021f781f38ccb7e55b10e92642390109a1681a37c67a15397eb43a06c383278d9080bf
z428529844f0416a10844f70a570515875b6acb73376f7acef77041bed3f86d15f9a4a914b15903
z56a06d732a5442d7696f2e9a8487810608f82d9193f8ecc05511dd6ac953e9c765085f12c2b88e
zb76fea022c680ca528d6e58e60791614b6c3348880d3b571570aa7cfd9773e0348dc14328515b0
z98da059dd6088987861dff04ea5e5016b2e0b6182aad2e5b8e1cdf843aedf0e74e949f9a56852b
z21b6f60cd2612202994b720a5869a45e99940f4d016e0292b35d6297252bcfaa93627fa936f6d4
zb20b55dd3809d5ccd85f1286098e8d4799845e10f8be8b72c5469929612146bcd860d80009d5fd
z8ae47b69db2afad47474a832b101e2505aac3c2e2c7701becfcfc4293beafdc338f88929e4cd3a
z029cc83cbb6be0ff5f4ec1f0c86fb1415a68e1e8ba3410a82d7a5688f9cc8193bfd87471a73666
z232de6d0f13902e301a25b8362fbc85ada896c70a4a205c8695faa8bc5dab1125001b36e16dda1
za387b43b1601e8033c67a2805b1e9af5e5103648b2dabcc88678df3d90329c09e92bb5f2eff85f
zb321426aa1bb3ecd7a68bfebc3fe38005804277771e7b1df353fc60ce31fcf2443d82ebad0c8db
z9fe8da6b527ee198c00144b966235a16ad7f492f4ec0e6ec55d7265bea3828fc0b72001a52a91d
z1eb1b545740d5ba4642651a623ff3cdf1fbb22fa8ad53a96c802175accca5c19c6b679bb7c88f3
z8e63f6d8b816f3e1be5ab05c1bea523bf331c10c76cbaa7816c8ba7bc62fbda9135696e1d9e8d8
z1e796b6e86ed4adcdda83d3cc2fc6537a8700dab656e4f84bd752a3f4d4347a02ce4464bbb0b97
zb79b0f7d8705ea6bb8fd14c4d4cc03271f4296cb71d7f4ea5ef6e3c5a6e3e55ca5ff3f5126d491
za7f5cefcee63397f7a86af34cef4b7cc0cf6b514d60dbec436b5ec8ef62945de37d5092c2e124e
zc863a9ce0a04b8b8fd0c2d421b01559eb1db84d9d6c1010a0cd4aaa0b80a159f34010d380dd090
z3dbbc68950becb066f9869523ef9fa22825ce679ca15975c142929c9486040ddd3cd961e88b2c3
zbb485739f9b781e4f7b787dfc6e4b89430ad7de5f67d7a8b7582d00c49293e2b459a2fb0542203
zc89ad7b2d82f12679e73f785c0efc9976434b542f5add5f9e22fc5880fd34b6627e32908238ec1
z7cb7bbcf58ee6f1f73bfdb94cb6367ea0edb0736221e5b85698b631f69a1fe5cdcaeeb078905f4
z73db53dfc497b85cc67065080f5b0b3d5aad39542d25f47a7f37cad2585e4b01f66a37516cf17e
za579c67cd50ddecc21e581c93d2f1d1bc8999183d08b376ae70c1c558c2a859a3a478574d534e2
ze42241f8e46bfe72a3ee0c98f76a6c244ff05f1409931aefb369c4a8f0ba1b8ae2d2eddc7df430
zc94f7155ba75781afd0c15793ffb5d4283f7a14a0b82cd43fbeea6acb7badd476e970d15053ff3
z601277811faf7dbea4150b49bf3c958ac443f1fb8b7c6dcf7ee5233d88edeb13c44fa93f7a5d83
z866345e2bf0ae9ceca6ea814b7f8ed2f5aca24fd56bf6ce2acb5c313b76ebbc207adfeb6318ded
z4ab38ee2f7bdfa0c4c4fc97b21cc7167e56b5de1873b2a791d3365024382b61f8bcc7db4d6f315
z0eb05bf6721cc38d74de2c75f978c1ee433af0d1c5eaadb8e89fd7024bcceaca2ba772d4743b64
z1f7e038e6768904781c1cada78006d6ccbcc6d11bf1c4b9dec0a3ba616344e319271e315736f0e
ze11041fef87ff93d8d686cc95190e1ae33b1755c56360e667c3b0c1cd56ea8fae3211b62255e64
z3f44bb0829f58b45acecbe2cefdcc33b4f28166e3dcb807107c58fe6ff8708f31d489614db706c
z403e59ec741e905f403ecf975886adb6908e25aae35516289d4176df40c482cff05131540b3fc7
z22231e9bc86f2745c49009b8c4f7dcaf66af24da277ef89b27bbd819f9d7f6f3591f859a3944bd
zaf9094c6b95b377fd15efd18c998483d4c4520e0248aa2a15538b97926111f0a2cb750494c6aa1
zb593ba78a0664a996f6626d15ed67302377894a6abacc07f713aec874f2bf7d840c87f476fabba
ze3adb83f5490606c2ff2afd2bc19cd75901e0d2c9ab00c99061cab77f04f8a39bb1bd1c68e8ecb
zbafeea9835e39433c896749a37172e33c6da2b4a8aec4b7ced5d15197649904fdfd46bfec9bfcf
z2b2fdbd545146be8bce5ac443764fa6aaa50094df16f8e376ba71d00bffe269aa7acfa82c739a9
z848e80656d422d1058a22105cab8ba297072feb7256e894689197f299f55a7082a7d60221ae8ad
z98aa92e7eb35677a1252f8fc94b7576c821682b3f394a4306ced0be0f32965323b7e11c8beaa7f
z91fbaa32d5e2ad4fe3959188e6e95b6b25fa7d817db78ef638ed9a73534ff109445280014c099e
za7983edabac0cedcfefd202f49e42a3420c2c63a2604f60c5c8356d28659245428be3ecdde1767
z1329b3bcc383279498ac9fe9c46c7f85584304e1da8d2d1e6c80f2f6ffe59d08292cb336c078b9
z21dd03349cb0898342814108d11ab41699e35cdc44cbe75ac798c41b7e5b65d59858738df78df7
zefcdef5f76554075c07707479e18d675c0a04eab310c6728e91a6ff5a9e4101aa0894e49d7013f
zcb55e6c0730527bb69ef9d7c601639b242db8b1d79011bd44fc8262b0b16ea196d010b2f7888ae
z4fe02a682ee7d1a653a04b7ead36d7ee74ca897a56209b5d9ff4c1940c5cbc72d533e9650cac8c
z22467f25053f81cdd2379173575c73a46f76f0c410a934a4a15f7d899917be6c9d9004946b0f74
z49238fb33da020515e7aaef62deb39c7c9684b59c7b0060911cc1e9b00880e031bbcf0f1475f7d
za2eb2e91c93a0d0c8134938c1aac4252c415a2d97b6b77185b5dcd460163e179f69ad4052284e1
zf8d939026c2511b7d7bd10b84284c7298dc6fe5a73da67a3651c59b12061c370d3c0cfbe2f37ea
zd2a97af549488c8cce3d3890f22ff5bd53affc40248f996d50f12b483ca1e7cbea2bc0ec241716
zac8e836bac3e4aa9c4ff6612c129880e2c471b36bd6a05e46d8c24ee4a67f119d9872f0fc458b1
z414e447aa4ecf1652a594361e7f0c0b19054cd7b442185673c8a319e5fcb12753fbc586c3ebf89
z7476cad79dd36d3e653f64704bf376d5a54a25f2562356adbc2256b7f6fd19c74e0f6520bf923c
z373ce6484e04c1ddb556c5cd4714b491f46b479ed302725470b48cfa81f1a39a1ef264ebd77302
zfc54b5e36e5c929d7a386236559f2fa13f89bd27c61b28277177af205aeae29b6435b942710a5b
zc7614e058e018c7a076dd98262c9963faea0421d73dd2b48b7839207d3296acf4aad68b889f11b
z892f87bd0313edc49243712152923661609264db4ace89a9e480712cb4793781ddc01622272293
zec3e227cae8e805d6b8f3aca2ed51431c1bfa77d2163fb83c100083dbba009813439ce929b578c
zc2f8d3489712d5d51e8f43da60d1c2efc9c837aef629bfdcb34f873468170fc37db7773290518d
zc494993ac515db52a9eff325f4b3513e28ddd322d149e9139473e42c2d056a0ffa8421470b8988
z146b64be1d54205c2beb669cf5eb2a9cb8ee1142339971f4b2ab8c4db0473034ae2729db8af5bf
z4455e1bab6823c916480c586c00ce0ed5a44a118e27dd608b992d5cd9189ed6d1d0da291867c5c
zc6744715a65148343f6e13a6020d8c5d62f0634031feb90884143d168bc607b136a2fbf85600f1
z6142adc1f57d50d5dcc672b21e4cda3fff813c1a3a42f9fd1145085f77f5252c4ed5038ef6028d
zed67e5163b20f9dad35ac47d4f4525619b29127df6cf637aef187aea0e3f5bc830c942439615c4
zf69d8db8912c1f542b6a009e74e45625b2c2aa1c746c3dfbf8f7db129fa9cd312c4dfe44dbe36c
zf1f0100b179cbfd27c40a216b104b75c47a775ac84d2c1de5ea857bc2e50c60aeff0ae6dd4884c
z3f46318c0cf403b967c3f3fe53745a1ceea55bc89feb9638920482f2e873b6b459ee6545c21c0e
z1228d85f624765c4381dd1ce3bcf343ed7b70f380d321ed7b491f22c1e22cc2bc2751493541414
zac98d9c18027c6fcfed5f6ffddbfcfcc81b18a6a78bd09bf09ddc7341bf871dd53dd4db6ae6f78
ze234b21fa0d8db47e2e35260abfd372af30db7e9940cb29640098f7f5a5bd8f63c36bcc9b867af
z8384c428acfc5d1a1e11e00a7e2d3708451fa5c36c01e49d1af57916fe4f272fd40ceb55bea14b
z1f54a993dc3538cb66cbed3b8a1c5bb6e4211f13d7a60f0954021fb24afa901fc21353868ad2ff
z4643d48ba10f706ea5c5c7164dc74c21442233221471754acbb43a31961f12c7758a159714b187
zdfbdbc78a92831be238b39447c3a1899c6107e32e7ba4a15e693503b70e053b5a37e2f2e8b69f6
zeb2f75429e3958c429b4a8fa158931f620e810dc71fb104315f07a15255aaaebe0f43def2f9135
z398ec457cb6a7d67c2105f3edb0cbe0100489b4694dd7727a14b0f4853351a4bb00dccef061c91
zb545c698ebc6cdae9f3f043e0250ceb67e68d66c71efc470d8ec1e5926f2ad6e8487c0f68c6498
z4ce4b8f674b025cbdd778fa4e5540949a07fea5826610fa5207763ec38f7e06c3973f83e18d963
z5bcf836b0c741b2a4c920f0703595ee25ed99148137745d25da3f0a052a0e50337f870ec30055a
z5d909a25b86cb0074e7d91d73fb24ef1184aa61a80010b4e26f29211e122dd3f1219a4f7ddadda
zbe626583ef5d5f5aa540ff3ae8af57b366c8820702eb26d7dd153407b98d0a9bf7e723bcd5a529
zee6dfc2610d7b69ce63809ba01c8b01bb5ccc4fa78e4a4045cc4d0707fddc76768b7019e2cd498
z5eaa86ad936e97370a34d675778eadeade16d9c4afa8fd6ed5018f87c845882894825e42d955da
z53ee21031706a5793581b5623713f3c16307c3754e9acdee318c4782e2c58942c697d4060c49c1
z6ae3a498c3210303a8b535b3963727804d990729e990e46666381177680fe8f0f7aa04dd875b5f
z466c6450e2b6140d925419bb184e5292e0d751a366875ade67b4432a37d857c48efe9cd97f49d9
zed96bf6d21352b63322ebc4000bac5b231380ea68e4d5d5398b5b578263d1ecec48a6c11669720
zfaf866662248cfa18c63bd85c323107ad265c644e108478e73aaf3d3042b7982ee5e969ffdb451
z4ec4522ddfaf9b9abb30115e63ae00f7a76e25a2b0488d83e3fa5e5f10058a90eba03b14ea2557
z7512e11189ac430923d5ed683810487c838519a4f42952b56ece0be8bc00e13a4efe043b035661
z8e669905a19aa9f82c6585f6139d193a482d6ab76f3476fbf576c365418bf2bd90d901c07ab478
z6b76c0278da0cbb6918aee25ad83d3aeb78885d83aaedb21130443e4c28a5bd669208d495b7447
z79a31c1f6cc94f26196b0052ab93aa451267dbf547d6386a9021fbc113b2bcd2d3ffbc7eeed3f2
z80166fd636b6c68c411148b6a020eab31a47c01eb790a243f4abbbdd42e2bc973a645a2ba77109
z208cb6334c6e975c1fb5afcc6ba92608f3f130d5068ce322f49c4e9d2e39547aa125f11ac24c51
zf7da64edb5b1625c28a412de1d5525f61c0f81b7623ec2b30f748d09ab1202b78960b9813854be
z06297751a5282a25353949853c3c04b7efad0e98ca6a5d229f46ecd7dd2d57c741d59f903dcb93
zc3e8a79aeb5b8cca342c247f2030253e40ad5590b53205258814dbd5bcc865a3b423c8d7d236b9
z4d63ce8aa616501d210e85587dfedf67d8384bcc6163a00a5e0a5a5ad812aae089c61044cf6deb
z2387c5a01b6888e58e9bff20f3b8c75dda96694e773d51c20c7a4e590ce3c3d5efe6ef7a8208d0
z7765dd52c797673804c3958089e8d154c9f95c0e3aff23c420af9b6046073124274cf2da64bcb3
z2ee422fc912172c88991dcc915674aa6e5c49c3c5e37f3ca89bcd44b36ebf28c05d76884c55af6
z30c5b8879994fdede79f3be22e3497a93d01546f8504353728e52dfb5578ac6e5030f473dbc294
z8647b79b957091ff31de4b4e6ac8034250b482d2a3d4127b77cc1b70e2fb71cc1b2526c79a3caa
z2c96ce602f21aae1207e6ba802eb844d37ead25912a8ff5392e7199c5d691ae6548d9871cbac7e
z326b1ab284f441f164dff22672609f9002e82f1f71c0ff44dd86f7bd9c9c5cbf2868c300857b81
z809bd349689005147cea8e36e48515c3d4f5fa4d8c5563f777ef8be5178c3378f9b426ac0075b1
z0211a74c9fbeaa778705f1c89bf3bd79d17341ca61804206edbce07d2462adc921fbddac274fe5
zcb3ea26773ef7232e89d88631cc2ecef8a16c596e67fe9660a85eac149769fad3f66f7ba7af773
z6c79dc1be4d3b3b477f8dd8f968f7b6ae2532633fb4b34be89d247129b3c77ed620fd8701c5beb
z2d29306294ec1089d9eb6ede727350f08d29d98a304f8c80953571d968e59b8bdb040d88815d3e
z1c6bf63bb4746d3f06a69829c115780bc9b4d1b3eee31ce8d489e23b48967d87813c0fa54fba8c
zfb596e45ade4dd9c2326719d080646932b2bd591475b8891552dc3962868680c5d6857ac0e5af8
z7dc90488b1bb50c17e9a0699e59a2ac1eb45626b6fd884ea285ae5d4857b42f80840fe940d3723
zb81fa5e085f41e22462981c7fad60edb19083b4da0f38e0cdb6b3793384300e4a2dcebc2838041
z84650185ad3b36b13778729c9e6dca6de0046b1103d5621d41e10c6126096536bf381fdec70c14
z2bf06de370f4af290c4e7028383b8ee603e282e0d3e51c9025c241e872e8baccbcecc5bda5ea32
zd89584a9697594071d2a1f3a02206e0566997564f6abc928e711d79360c82f713d0a3b502ebe1e
z5fda96a70f7a1f043f292bedb7bf1a88c7a01f3859462257d92bfa4fa18f08a26415538ca75678
zb353e62001057a05c001854c9e35f61c472222259e290157f7e38e8c5a99ccaaf8d3a3ba8478dd
zf459d5061afbff7360327b780d93e624993b949a16736ed2802e52b7ae53fd935aa7063ed6056f
z6bdca2ab32c35817cbc6aa9fcf110aeedb1e4d918909f7a0d766c82e3f5e86160e9a5acce81f4a
z964a34a5fabb6b10c36e6e5390269d11c133f17cc527cd3a20f509ef1492a8feeb8939da70e77a
z824805581bd27c522db288074f8829f76b040f182c183089dbf078a5296d2172a414f4e515f7d9
za664413acb6415a37d4681c3d64ce4120afc2c1dcd00594c62afcb9ec9ce379dddf3cccb8a6b7b
zaeede7a25c9d312d8600372af999fa3b5af0b58f349cdd878cdef891b6afc92dae94c1354bed3c
z1e02d3ce4b1462f485378cb98dea1c5291f363b3d16776c23a9326dbaa98cc7b334c4f66b4ea54
z4c7dcf6f3611a98b8955f6c735a5ef8df7eae286f7405cf5622ec29587f0890642667d7b92473f
zd401baaf0cd213735c7ff54377018ae7a0dbdfca6fcd4a7d1910c64e2d5a1ed4946d2bde9dabae
z057b09bc8493eeeb3bdaaf7dd5e0e16e5d0fb9d59d6a649a39efab002a4c03fc0bc6307ce7c370
zbd84f05d4dc23d1587853219cbc970401a00cb9a90930f3a41c739684e7ce117195ed3ca0ddde8
z098e021c84838e221d18e09fdef43e2754e3be577988eb007eb06229545cfbc3c8a7256f08cffe
z0f2ab11c7c6b3f7ebab865fbac9dae447c8764bcfb1b139ec515472d1dcb5881bde149b08b7fb4
zd96460649b9163018c7e3ee839cc6d07643f12b9f52de16df213e3acc564b1769be94243462112
z43bf3e55375cc63585a653f70c0d982d7de145a34e80417ebaa69bd63ecc044b3b53e544ef33e9
za3bc3e8797445b102740e07dc50a4c53d892f804e30a2609bb42f7f4882dd968e359471dd9607a
z6a629efe6cf62cedd17dfb65486ee67041b08f2799dfa8d583a18252904b90a2a05efd667f4c27
z53818370af16dc6b4c3de92a77a2c09224851aba20808a254ba76f8c2ea0cc45afb50a77ece65c
ze941d298241c3ced1433d53882245aec0bbb38549c6903fe53cabaf3c63519bf31fffeb520a241
zfdf8ce6391432b21a38ccc2c8cc2763d4ab8bb056aed900d901429cf23048abfe65d443ad9dc6f
z0c5132564785b050cec8a3473b7c77f49f2bd474a5d02ff62a41bbe86a42e37b11450f8838ecfa
zdd06d74a10c8193d7a53628fb2ca6e775abf236093b013fa2b0ce2bfb4063a399c6beca057a23a
z2038102b0b0d0276485c3b73cb9a42952e49564a7d0f0c04279aa6990607d10aafd0683ba20ee1
zc92225111b8250ce78593ecbfebe107b812dee13ebe16b19ee3cb3c5574d9fcc538f911f2bfad5
z4e62933778c9747d23d05ea95f82c41ce03657cd3c159733d432f5f7dc6e4c21c966a4ba6f68f7
zce9bc9248e791409268aa7abcb316d128b8cb60c5eb7b6bc81efd199b932da7611e812ef368688
z2798fe688e9629acf1fc39765760ffad57a0f240a4614585d61004275a4d2eb2508790ec9ab99b
ze6350a616d6b9b7dcd2f868fcf73af8eb786991dbde814dfdfd3975e103562635184228abdc09d
zcfeebbe74f1ac804cbb347524708c8f80b82a03714628844ee2e388e65ebc78ef7e679f3104ad0
z3b796b7fa8cd1d261577741fe57e7c2aef0234751b62bef849d801a63dc569049c9f2490287db0
z0807923c01f371735f8e31fe5a8b9dcc14580ac2fb134c9a7e21676364d68f4fad6dd4ef6b173f
z02a11d7a8389f09895d787e3c661cd84a937447a3a339c261f6e4531c0118a80b8e59334157672
zc2450154c952e9e0d70c2241170663b64665bd4ee7be624ea4566929e332eadd41084cf27af80f
z16a4e81d501fe75fa796f68c6a9cd2ebe8bcedec97b53e65aefeede72216fe183abf396015df93
z415afc6ae4ea8aa2c161cfbb4534b779fb8eb8051a7e007be1368b5b9049ab304a36ecd924f47b
zc613e2c1b8594a36a19c5580f2da65d67598259fb879b8e60c36fa86bed2f4ad1d5997ff217e51
z30781970067ca5c176e99831477fe956ceef61440927dd412a4ea11ab34617f84fbfcf132ebbbb
z7f1be74145673548a3ff0e6491e2287163de2864c081fbd0de96cb49d2adec26048481fc896e17
z8db3e4c374cb165142e0640ac46d1a5f2370c7c000b31163a720d28a2881755cf9ad840168d4f1
zf49e6702870ca521d6ecceb02b311e694102f92944af8e16e9b034308bb4c6aa867a5dec5b166b
z7d6063f10ea1722fd8eacb1341cbea60e16a0d4db9eb545c88b10bb87b4743004adae15e028f02
z46e7684ba6d3d3687a76abeecececefe0a186054b67c1ef94b763cc74912ad541ecdd6c75e3856
zf1d7b4d31270af454119cc8105d0f3a0926a5074b8dde4ca3e411f41105bdee22e70ec4591ab1b
zcf718b2b7238a6c5ade86c51fde83de46ac7cd20917b7b7c3120d1b07f77a1f4261812a7622e66
z71e1a19b3736c452e37813d73a88666e434c484b9d44a04eceff62aaee604b3cdc59180d6525e4
z19b5411c7e4cbe62768cc22e1849685fef1f74a99cb6ddc328bb003dd8180ef40760fb093d1e85
z8055cd752a5cc133939c02171a4f057391b3d776b4cf4852266e0fb30f8323b1041b5289a3633f
z67a7e0e4a15bd62f59ae3fa2870489ce4f8417e89d220471397acc928a6371ea476fbdbed8cde7
z3db73182966d9a957e9016a9e8d6eb88dad0ea7edbe0751c3184e37514e5a04c3217e68d9e0306
z205b5e1e6388fb33962cc1eac3dea90200fed0f3c762bb39ecfc015a0812e6dcd219f4a9bb5188
z7704701b31c384f687e57c65f60323f5e9017616dfb6466a2704a6c97513c1eb6c29a9e1581f9b
z17e6b3b8ec909fc1da152bac74b3bc60b91733f1f759a5585a3593f6a8712417b00e9487305661
z24e74351eb1ca6e377676e1de16a8115744c81700fd699bd6e340cb8e514a034ce226553948f54
zd248591cf169dcb0471f5ff07ef27d880e286fc126829b0add52acbf9f2d163145f56401cd2efd
z613194911e8112462122de54eff5351277604854fc319372cfbe58b10af378eeda57abe0066344
z36e0d237448595c4605a1895724f63cd57b42ec1c3e02f9338363b6556547de9f10b8a8e76f4d6
z8b1071adba41b74ff344188347321b6e31bd6f390e92aeda684be25bf44e8bcc7953b7668dbea5
z9c55b9cfaef6febfd5516961ff964b7adad0c59fcca79be3c12001f643fcd3a24b05525e4e0741
zf0fe8a1d1a865dc6009ab2e8f095662508e41ace8b0cf1653f7e41570d45dcca9d99b39b7c0447
z81e0efb4cc2eda24ee5cbb096aa2e53ca9f2e66331d9769743c1e59c9b71ccb015c4698e22c03b
zaf1760fa876c0c44310714bc1daf3c00c342bba750a03cabbeed6960665b8b13b0e1ff620d3dbc
z73457bd5ff5d2c1e4d050cd4c62674ddf11c28a413230082f8d8df50a90ffc0d5e6a590dcf6228
zd3538c3fb3d2f8fe843bc82d04c3f1f4552b8cbf10d38d26a18697b2f278d1d909b2276b96e20b
z33de00339b02a33a3bd6ea7ad20b01cce3764ca24d7e06410bad2450d8168326430ac35ed3bdfe
zbcf6de1f029500ebae05d33fe5f5599d1d310947fb5675f76b1610e03fa5e0f13d9ab5192eb825
z8c956b43bc928026ea48d5b96c134ea115b872a57b12c4b1f56fba2304f2375647458a6976b184
z25a7256b20b9685ca62766933cb92878ebfda40a28d8de61eff5d33f50415bd8ddb1bf28817c2f
z140d6a51ed2d27fd81ab1f676c8b3431a940d7326c740e9fba7ebb2fe98c102a86497b2c28540b
z05c7134f202fd4296e68b4f957ac13aa1a5527b8114018220782a7f9997e63f663d95a46985c80
zc4d50af426ca01290cc5441f371a86b678ff855a74ce88df3e3717b54cfe25e47969c844161071
z5d1dfc5b0d1651f73a663d54ee7a1bd84ff20f8c1ee2c0bb9fbcff2e064c073606ac2d69ded725
zf943ccd9aad59b794a857fbecf74eaec68f9c65b644c75d50e35b8daf51f60dba777df843840cc
z36fd7da38c38ca4e7a0c0a722098fa1f12551c88158954c929d918ce3abeedc0fdbcba3da15b8c
zb1cfcfa81ae594c5b729b97d250d93b1d9de99a8e1b2aa3bf74a3c5e7987a533a6c49a9faace51
z5da69bb5f64113a661a77a1f2f7dc0d8a69e893a20f4721ca844cfc7ff43037462d30e0779417d
ze6161d969830f21ba1cab37b8f8d9e1ecc95f316d3a25f24e75d2e6d8fc72fbbb923b88316037a
z146388f841ac3fd5d01386e9b0a476b0e69de5284bf6a47d8192dd317f907d2f1980801e567b3e
zb9e9e376e4eb5c027f11f59994417266515d1186c764de85575664a9502c518f74388bb3362f3d
zd60c5862a86e928132850b7b436322cf0c23e1e165b99180e8e6d3f6975ed9ac606e483ee9e799
z63e589b2881f98b784d8dcce769ee6dc01130e7fbaaf0763fcd2e5a3ec95b40fbcb55cb4091614
z316e2ca0eefef82decb2660430a06fe446394ca7d11f48cc1f43bbecb5a324e0121475a02e6e86
z8dcfdfe0d7ccb28df1d271dcb49b16897059d85cb87074140413b7ebc4f483ed2f409f0318f786
za8353a08a2c00ba1ada652c7630b2a323f9fb652008e355393cad4a1789cfe0376ed100f66b15d
z2ac9b8ab5c8f96cf89ed7522a943f5111ac202dcf07309a1f4c5f87ab17569dd100cdff2bc18ea
z127adf0d6fa80640e1e33811c1b86315beda31f8797bbc78a563ab19b73578c6aafcdeec69aac5
z434a32904f1874ea8167541b1d541096b1e85c32794c01fd68ebb3916cca19995e579cf3a9c738
z7d6854d815183f477d8bb10741dcbb25b9c5dff068ef6d1d927f2523457f3efca6c57cde2e3bc4
z79409c66d7a34cfe4da553ba2e4ad07533148625a0af155adef84bb170936ca696a322ef02d73f
zf3ba30cb9c4c3361a920905eb1b884ba48a22827d31f89a69b37f0b67ad15e1d90a306295d0c2b
zb425d794a8e868af8da1bff74394d9e5d3f549abff71c55abe3b5bc4fd2e0c37a7e3da33f7a5a2
z5800661c7691ff6af0a2ffd34b646155c50f35041bc75fc15e832b82cc7940c90fef7d02a93cae
z57783f0a3c9e229b8fbdaec096d11cc5d877dfbb1c82da795bdf34fd9fd11d4368f19d5e371112
z8b970ea6fe1edeadc426a023b109caa34a64439d02f65ee37e1a7295af0c7c72bb3c4874995d02
zfdcef065b16711f4c00d43a56de4cf4896650117d8de90885b8830ebf3aa766c90995441d87687
zdeba544dfe3fa6b17b13e1c0d2bd73c6358fed2bdbcd08a56c010c8f35e43fcc0d1ccd49f2db5b
zf98e43cc0cdc5d25b1c0fe6a815923bb12d4f37b49f244666aeff1b7487cd9704df77131486592
z2f5b8bdf1215fddca11a53dcb7aa6b623a2f892dd683ac265c9a218b0da487443e94ec14c2e7f7
z2fd1dc2e81417d23ad37132e5f89c1776e0408a444fa6406c9dbc5b1772c5a66449b92ec0044de
z7754b1a1e9b8b2a83a3f444a9b28d76bdf6aeeabd74674306135d03a36c32c1113608e67bb0852
z6901a194ebfad824daf33611c939754673c30047f55a2cd41f81644f52925afa498e78b01a3d3b
zd76b20ff9edfa8bcd5db573d4f0262a6b941004e1226b7b26673285c3811989894bf86ed4b75fd
z75fbffa0c9da8a6be74962f079a37b1c044e5f945502b2b855820571bb19655e8902d0376a026b
z54dd130cb1b414fb5c60384437e25d41828fbdcb5decee6998895402d5122f8069c8718743b947
z8189823970bd8afb131afd8e106d4eab3f5e3455ec598b1dc6d455628ee30b8e4179e4dd0950a0
z0f44fcda23f6c33012e30fdae6a7fab338b8bd3981f9fd1e9024ab302a116f322cd8df5ffce5c0
za9b2021111958e5e329124d77867dfe1d230cda6f73f07227a985418bd02a12e0ed21d8ea71b6b
za921360a54c0ab62cfcb530fc0c62066b62ba5aadba67bf5852be5557f947d9cc39babd37453ca
zd1cdf711352faad3dddfad1044a24438e9e790cc86150b8b6c58fea80ad4be5222b25285cbd7a9
za20efa355f685ced638eea9f4ea9dc51d3bc80bdd37c6aeb5992ce6e79940dc13ecae973d5abcf
zee89d5a641f1de37815f1e1d54136e376e676300c7b3a1975a75effdbd6298395dd5c473c4531a
z7dc2a303f30747cd669c53dae37b74c2ae292445899defed8ddf90011709c18e881668e687e8bd
z3dc33e278f6f7b066bee66dc18fccba0933508db94ccad4f19109e025d77125777f801034d7c4f
z215a7f096501038246ab793e88eb9b3fcb93b5fdf5406523377694cce53e1f749d07aad57c1a1b
z6a1ba10d9b0ac3f2a31cc043646f9c0e934ab8e6302b6412af5f9966509cf447eeef28e120ae6b
z93fef33a7ec6f9da3578535c0bdf4099656223578291fe0e33b9f4f85268cbbff6a627fd6961de
z8d7aeb48954a309a596809adecf1e7e32a8374cdebaac7fd78ffbde6679d8ea2f3ded3a75dc3d7
z8d34f1331741989832c54c2145bbf5092d47c015f2515da72bb83ddb71d11d90a16d8b88a1a59a
zf87f43046db0e6a7e45d47bd98fe0c489c44a2bca92a6321dfed689a7053d6982b6f6174e47a7a
zd6c111d443f075138ffe5f55fd509a5cb2377f1af7d70fe4d0c323bf33f5818fccc4099258e80a
zb22715f7833411a60ab5bc6880a6b4251556d1183176e3cc46da06ce089c267fe6605d915b1c02
z8cd5441470b0e0113b492691a2225844fdd837aac4b4fd47a5f1ae644c912e62b880b6d7f3affd
zd3eb03da1dea261064fd021ea6b4a1a3f42a68ffc2bbaae3643d6886032728f801280d67630a12
z685237d48e0903565762347b1f2decb99f86b66e13a463fed582924664c92377d010428022b66c
zae68a5e859addb2fd687a71ec1d0e212f9b96fe992dceda8f74befb6234c0362ce4abf6f8e89c0
zb9e8c119889fa4064c6a0f554d3c30bce41d78db6c8e423035993894c8022b0fabf81c3be2af75
z4e6bc22535259282838be61c64d6b890aeb3ef2a5612f533bc927c34d61aa31b096ff294aa7776
ze29e903d8b9e18d2b39ef5169917602f1b78d31e4845c9e199d824559548ffbdcb6fe0b6bbde71
z83356b104154cf871a8af4c0c74836348cacc658f44bdf24200fdab4b5810b527aa14bee3335fe
za62b519452e0aeb2d81bca0cd6d9517cecb49fb3c881b659666b4d81d17906bc7f103e9ca69cfe
zaf46f32aa5efe9ab28943412327f4fa1b24dbb258a57b19d55479deddc9605ff454d83dbc01508
zfd9a77119ef6b398b4075f2123d90fbb0e22c063aa982a686526d8b922df470525e24486aafea3
z2ed8b078c8f5e05477383f8a3cafe3620861ca6bad754411b02affacb965aef2ebfe6709385688
z0c77f153bcd2d9a41872e6c27449c6dfe0fe6fb5285c6658b5434218b69dfce773b8248e494142
zbba6b49c645bd28ae51d64eb24587c5272779e601f67d51b4743769092b627e02c176304f811ef
z0b17d3a4aa7020a9b323351f6ad407b138e74e0d4894a3fbf75178f3ee49020a592afc0151f826
z95400ac6647151e11d0d593b0ad2ee0120db8f300a1aec21ee42e4c89271e8d79fdf53bdffec64
zea256864ee37c271dc2ed6d7c411ad661cafdfa6a6e9f7ce9c21d3c2f3f3bbcbe0997d6b799074
z8748b9fbe1eb2422b3d904712a31d1ed94b8c5b5cb265571c400adcf892e14aa131ff1beaa165a
zd1231ea9f29ca4c6cc4e42c3dbb5ddecda9f7fda2809aed24f35c755b9730673a10127cc2dbf46
z420cb3a6e20c3a754dfbf30f5f0c07b49fc7d4db579788c5aa56dd7797644ae15a49fec81097fc
z892020fb8f9424b33d3223c5cb306d8a9078fb93073da659d1c4e13fd2001ee2f78ee4157a9523
z1dc4fdc68ffcaca6b03b79ca6fafa141f61410b927313d738dfbc723f5aae0ad7dd328b4fec117
z5f33e2cdb5523d06c24d412db44b160ae11067ac213e57874ee0ab2a690b44d3c48a65466625dc
z60a6b886b13af334cf93d87e3d4be233015524a2007dbc8b8dc6ac7bfe2b98489325d36ea9054a
z3a5d2a8662f61a6c6d26c8505f501f049a97da9e9b8fc2705379d919a356cfc41eef5f392448a2
z07b6b7bf3acfadc63af1d103cdaf6af6978322567424b0876338b34a0e5b001c082aa6b55255bf
z73280c661261bc99e7e197793f317f554a015203e2371851a4797630091d402181865308fbd632
z1ad4bdf1c5d08407fe440a84bd76c87460d6b9bd5e5410e03ab63f23ba74090e98373a532d1ba9
z001a161e337ffe361a511b91eedcc3a87b7f67a13a696e968809092951d0ee0ec12c5276d24605
zc8032757e1fa2bb40bd2c97391bcf82ac5d72b594d01f8351b1ecfbd1e7d4894397af0584ac91c
z9e9a2d2d7443cbb720c94898d5f5ff183829bf9f3d2131a367d397b7b1bbc45f0e6e638bba87a7
zd6d0f7e08a81ef90edd5c503e7e3cf9ca66df4b93d34b25a70ce489670b188a09d38877def223d
zef00750f419333b50345a85eb8f1fac6812c87e61df3c3e951908f409aa24660a2b3ccc48b702a
z1faafa1f24507b05a45f511d47e50045e0e73c63c7ea2e4315e480641ce95717452e48f58bd3b8
z161ead70bbbf0b004702177ad524ee35a2a33d3f83f0b54121fb1eec27650b806ca61ecbb73090
z9953e2cb64f430eb0aa9f7f632b05e098d9b02a08612358b6a30cd671c836b77791d6840c59549
z1e867461b3b3c916ceb00c8134f255d49ecc7e14937d7c23fdad2793999baebb109342b2699085
z9b05edaaf5a9e8cccf46dd1c719d32e049bc27c36d4b98379932b900240ed9a785f7c0a3747692
z81bcfb9e62cb8948e9322e01391b2282d7fadb7d8032147714eaaef98414323e4f9e7f0c9fb92c
z401db36ffa10d530d38f33e17f661c3ad9a30848832f92d00f86a3b34a0397078d6da21ad0db5c
z99b2c3774ae9b19f438776acc07c85486b14f6172bbbcf15c0053fcc25e672725832e32bcbad4d
ze3ed544ecce6a7e7bf0f4166c8bf7ab42bad395335c736c3dbccf6235d5b79c22fec15830aa6bb
zc59bf43d0435fbac1b3cccb8c7c2fb2849b423ea77be62e08c92063e59c02ddd34ec0f5fd951be
z22769d99d46d455eaff7b07e8ada3315b01185e81bdcda3e9cae802ef72f52a0986c326e089270
z09a288fe1f45a421402740b63c81b84a6d30504055daaec681203e885e1f81302cd68d8b902f2a
z234834a2da51fbc453a15fc1b43699dd76ad58aafbea313d88272126cea30c7caabaf6ec8120c0
z90398c89b1349ba20c5deff94fd57acd4b3f9d7b517a8c87179ff53dab10a76d5f02a200bfd5e0
ze3deceec73fad61f6693e17b30aa6e5031dcf58d9531848f898db7406fd0d64916a769b3a00c70
zf107c90f6a70eb0b0648d9e384ba4bc8d5312440c8da45e8ece6ea6f98e79a501a084cd94fe66e
zfda3c3fbfca0267da34ec05c6bf67d899d14936bdb14baefd3ce881a5438014a94aca50dcf7ec3
z6be96d54c009712ce845f3b8ddeff3cbb36c93a261b9bdb5c5b5023dd835ae7b17a908db9efc20
z091708b7c0c5cbb06543bbcf2f2dfdcc77784b37138393906f3968f085fb0246350a8cfdd92c71
z2406c7ea76be5e0242875e7f079e5fa76534648e1ecbcba01a1b155e0153cedfa75c9ccdb76f11
zc012a1999ba01b7169bb9296f5f66d4f3a7b3ab8c8f5d111cc20b35b8f8ecbe2290e76545f246e
zc16def919cd0dc9ca5b6fa29c62b36c95b4ddd542d225ebf8b63e86a6df00b91695feaeae8ce0f
zac03a58b68e4209374aec329499093ddf0e17d9c3edf28a25aaea257d541d5a50be63da774274e
z4b4910ffb73c68699403245e1878bbb4e66f6416e724ee1d64718dad1297a8b651447ba1dd7a2b
z1b7bcbc37f6374710426c8bfb61505b08a11f69b388b92d29028e2c6719c913d3fd720dfa5e27e
z2c7650bb7c73b69ce01db2666d1b61a21dc8634e925bab6f77e2e929e2565b463ff37568426b8d
z12d74e4f121b5019553de878859ae6a92e61abec3c1f79f633589d40e20d6846c2597170319abe
ze41b76015f8a056d5d1069de7e091e4e32e895925b71be914130aad4c72fae9abe830c20c103e2
za97a1e1073c0bbb986df867e82661e0eb61f29969959fcd39adfc247a7cd096777ebda5526ce29
zfce2822fa58713d6fe162cc20e05a7ac8f92b552622477de4d979c816949ec499e0cc39747cd81
z30a52b02736a88f4884a8606900a9fe5acf75e68e8089799d21cd3f73b98cd49f036cb65f91fd3
zfb6b523f96f61d1023405246b109c011d4b05926e82f418c8089e9be157ab7716b0927ad63db39
z6f58e1f2766dfe92e542132041bf16c6f1126464ae169d5536472b8e0a7e0eae91d66dd7d09e8a
zb94c7965d3c66026908d2dece639b478abe5b396c4a51670b057c560ae568071e92f8ba94de753
zf9e284fce75c9e50499383af2c22ce9495a3edc4b86a4a0f4ffb5618f266851b473b176a00c308
ze729517e6a4439926e3d2be3598940e56e38c7bd9b30f80fc6538939749efe0babaaa480e3301a
zf5a6340df74041992ba82d8295e22c816599c03a0154addafe5a45cdc5474e50999bd22d255bb2
za72300abcee6ab4712379359c19de34435d7266cdb5a30c5eec802ab108dc0cc166df7701c8e0d
zf22cb1ef93ac5394e6b09c007371e34f524db8278820683f5e1fc851d04181906f3601c385a027
z7226db9c373d29f3a2dea4648875524f22b8a7c4ba859e838f4dd8a24cb227cc3b8bca1beb7d90
z9bcfb80a2e7e3abe5c180aef022f9a1a57c2eaa3863847f08db4009760991ab04116a8396d21cf
zf68f4bb3b73a2cd9702f196b39a2a941c8ad712937a2f3ac3c247d87adac4168422cd66548c2d4
z0989f2c44465bb3eb5329d706ec30f59b70a3ae1b3113db80c94840ea3cb2cdf650e55a4e12a3c
zeccc897261868b605969f11d619de703a427cfc36317ac106ff2a36cd8f5592276d24401175a05
zb89c3e9bb69405668ea7f40b17cd2ca8526149fc1460b4eceec2364987a2b891e469eebcda227b
z37e717a4282e8f9f13d86422eb7a50886ae39595fe96bea498c0216c3ce4f3ebc5ea4c52826b84
z7e5d5bdc9ba8ce1b7f26b846fbf0f2779f4ec2c7dad6b4916cad070c9c8ce200b16a94ac74d623
z15680e5081e358cfb012a1a17a957dd666eb893a4472dc70d477e31535da70d39a9e983da4c78c
z10d5310b5d60a134116f0f7f01b7ceb4fb1771e3cc9516d1a3f05f3382d6d2ffef4996f526a31e
z2a8687ef62a98c5815d061f68fe526a22510b657abb8d2abd16b5527be6bfceddcc56e9c61a528
zac49adba50d020aad8d39eb98fd99b18b19a498e62df031e63c017b310858fe404e22652eb6c0d
z799c0b3f114ec0b315b709b276eaee34e8cd60a7b63ad22825fcc930e47877db342e8f7d31a69a
zef825e7fb18bd2d45d7e83e8634e3656990268c3f093e3fad723ac4cb47dec2696d3b6910ababa
z2ea3ca213d5cc7ba082859240b7b93f3c9a2dbca23e23b266612918d89bd14342c0e45b43239d2
z9c5413dd8a807ab1483873261f4365ef7aebe80a23d72811c3043803af9c1fbf095804831002ae
zfdc3c19d167c2712b8b39bd088229aa60503b0f20d1aa5557dcee72e76369308191d2c91b0cf87
zbd2b0705e3350d2980acfa6574ab638aec474b28aef2a22a662800ac15772172ae3d4e361f1fd3
ze36a8a50d8854a6652102a89c520db91a13ed08458be882c43cd395dc25e5305f64296b69a59c0
z6da54ef476ed4b5da95c906bd3e44ca01bdb7ac912c87c528b8825ab6efd5f9add3219393ffbb7
zdb59a208bde6eb4eb549ca891a5709b7115ad6a16034a0b0ae92b435fb6bc5159bbed42c25d1ac
z09afc43f583f9c25de652379ade0e0369da136426716fa30c872a1dfea25962366f36fa9f00fa3
zbb3f5cc085096e27c6a461cffadaa0ee395fcb22e88e7a1273b895f5a26f6e56fb7782199de704
z5e4d3b065296efd656a1582ef0eee98d2858c8653b81c90e2fcc4756d4e2185095951b84016d42
z0a16a22fa0a4d9bf8d1de79947b3ce5ad65e4d418b59b14153668efe4c08a0162b4636718ed923
zcc4394189b4b0cee8b4b54b805e1c50e67a078b3153a40d5214690e927de5427dfb55f195b2665
zf9f5401d0b028b1a55c34a0b9157b2ab9d303dc26b7ef4ac6373127396a184ce8c92b269283218
zd570ba74d924d2df2443bddd8aac7c8f3b5af70c5e04abcb88023acd7bfff4c694a0e0ef26d5fd
z40466b8889131211985f0f967080972f39a30e13c8ec149ee257a4c0b2fd8870ff8587419a5536
z3e521a97669dc7f7263636e80bc51553c4ba0615a583c19df9ab9f9f28a85573797d4f1a994a7a
z866f3df2068c8eb3431450307e71a31d04db2723463e3e7d0ee8f890b2ab488f9be4ff60c41240
ze570e40e9d8b150363ee242180949854528ceca24c9f2543ad1ce26f7d22c2273dc36877f5a2da
z3868be9f995434445065f04da23fbb7b71a7a64628dfb67fb0381f0957712b59d3aef41487a5c9
zbaf7e700f32807405953ea008cc80f1b7dd83a40b746dea99b8d926ad93bf0472c834e2105f5a1
z7c8678389275568d4a2933e8ee7cd1fe80e85a4930d63e11f8dc1aa2a4e920aa6c0d956d1fe211
zc571baf838dcd340d58d8f7fde77f7781111571a32cd2b49ea44cf918727a29bc12f88017d628f
za707fe985e045a1355281ca19302177434b46732f33f703cb3584e11c356d9a8b67c79c8923eee
z9ece88cb418a934689d397e64fa007912b2ad86e5f15be45cdf091a2960a3c85403396af9816f4
z02ab4a3898166e917261804d7b2b6f5237a5aaeb932ae7dd70a577cf57eaf2693fa56e3a61a0f3
zc31d0da0e0c915c05137b0242a7bd647cd1a919ec7417dc4f1a0d395fa7d1cd65a63cfd5e6b298
z2714e192b3b2c101a43f44e112d7658ecab22d3bc841bc92ed5efd3c96de1827b664f6d5f83184
zd373cdf98df8b6bc4d3f6b957b7673473184a5d3320a1ad3c981c02edbd1e7b9a27559e997c3e9
z93ef38aeffeb48739128f83ac5e78f721603615f9c42afc6e712d3d06b525bfb957343493c100e
z948fbbd86a5b89146e0002e1c85ffe6ad26e361739ac6c60be7582124246bda956322298585e26
zb03137fce993c9ef6ab6fc9c23871b55e1961afeb896d1e82396a164708596749904d2449e2444
z3321f478b82c0bf3dfb76a6229402ea26a77aad47307161ca3b848c0ec168f7c7db50ab5feca90
zeae4296f9e553b6bbbb16255e462ae0129b7d92af7dbe242017dd8a20cf1ff92f5f46f73db33e5
za90dc8586a4adb2afdcbeed0d90f0b7e10b4d85a9c6a5338393119091ddbc539d1b17530f63ad5
z7038419303ae5e76a2357f5912e27027c4d8cbdef02c15bd9367bc4e1a6d3f7bbb09d3129a80c0
zb562c75b2b505331712536aa564915421cd2171439985f79500d9b06b181cd7826d894fe9f01eb
zd7176dc42669894e97a37ae3c84622807cc436162a970ad7d844f4d2a3097716b3994983f983cc
z329ea15f265a188e52a93a3f41b2fb463e8589154485b8fa35d8c05fe582db1147b8da49c00ebb
zdf2147186dfce4488e07972c5af5508cc218cf91bdcc9673046d6c13450c804a8a1961fa84ab0c
z3c0a4b6374b0a9af00964ad9b4b63995393eda1e128313a6bf32b020fd24aa08bd41ac491ba9dc
z2bad8a11b2932ea22a46be2ddf31ed44d62ab9aabe814e9248b2fa162993ff51c047b7891ba26a
z4f7ece677e6816144d25f8566a17842ba842d065dbd76b719c127775ea2d72ee967156a2c5c2d5
z96b19c16f2e96715887e275a2400bb1d30c23b5e80a16c59a9da697b4f9f794cff211fe6ae457a
z007e068a51a5aa03b652950ebed9ed2a2016f7cfc0a7de2ea5f33d3b3872ffc8119ed9e7142823
z29eb7d5cec53fa1b23c2dad3b81bd5a6770adea50a63234fb2ef031a17495c60613d6e76763c72
z2cb4f154b7dd1fd6ff081ea2b5ac2458b88b2272843204880cd56749f69e8a44708fc06ba193d1
z0fe7d90bc0cb95f1baa2e8d1ee53fff1e44d92d215b38dcac833bb91230aee345bac3d3914709f
z79c9fa6638f330e867b190e05f9e8df13d8f77fe18684ae31d16259bcf26c5e9a2e22682b25693
ze91a4d08d90ceaaae3c1eb92aa04db794019f5ba4d128cf4832d792f29a0ae8228011d3ad1b465
z49aba74a65bfafc986a863bc9cdbb6bf29e0399069b6e8a6cdf703a312f2ec0ce3528971c3fc41
zb2af9a75cde05109088a6d5232a847a8adec0f18dac18415a62625816f9e78ee9ac065448b81da
z1aa67f2481f702e2a2f5fceb066fe49ef4d68a7856a0f262a449fa625c662ebef044ea0c9917f6
z50ebb846f3118fa71d12693c2a9b9464a38d0c67c4b65a25b4b1191d1f27d971bbf8a0f102a03c
z9807474fcd671a9684e8faa0d51fc88bede924b2d58cfa1f3568d7b4a1def9704161e7ee052452
z412bd2410069bbd2cb571bcae828eab68d3d3a29452f64b826412ee10855c03eec55f94b9f68c7
zbcae1efa872dfc1b596255d90dd556949470780b04686bd122d51c9512e0691b041a9db6005cb2
z3bd3b0251f11874f56afffaac17a667c8b9468e8b5ca342b3638f8015a51502a64d2eb978e6cb4
z7ac5590005fb12213eab43c56814438d406148d6f9f6e9ade00e857dc9bde801ec16b9f1c21e9f
z786d6c5a9c0e6b2526081e4a296a7d012ebb544c442f196251a0b1f880ae7b8891092e24443b32
z0fb5a1d6ea87c7194ca18d66ed9c6dbbcc4fbbfe98c2bd7aa43fa0a6ca0a73154add257a8510bd
z0e567821f46e6f12b5999393a063c309677a1906769cfd26506e83cd4858904e9cb9f7751636fc
zc4d0acb414104a1e22da4e356709f0a8c9807f1c63b768cde8afa4283c003e9960b6c3a60a9b6f
z0dcab4b9d05475aea2f0ebf42fde82156578ad4d1fc001b076478d1b5c50e8e39d3b1b3d62214e
z159c3f8a00f3cba419f914766227d50e3d05c815d50df467d0e13fcdc8a04725cd4ac94e94d5d9
z81ebfe81367aa4d2a5d72d84aa34399ffcad0f2ae33438a40695c6acdc4034b534a88b1b23cbdd
z3bb828b04863857ca9773f156b3365dd0fb7ebaf8f1ba8d4ba84204726fb1ac4a80834275f8ff1
z279608e989c339aab03a5f3cd3ae8ac97ea88b4dba468ca6bc7bb0193cad8e4607da3dbec0c930
z772d98bdabb347bc7238fd55d0198eeac128d9a971e0ee75fcdf8dfb08ccb9537c5ce52323b01e
za8374ff9eeb6ac4152cfa11d9f9518b789397ac20a66f07a04d2d9a9eb3131ef3428dff0129d0c
z4dfc6034f07a4d034ad644b85156b064f29e62ea515792a7a47e51e1cb6b25aa9ac1ff69cd4341
ze45cbc5e642f46aab68836ae0c014ac6d1bdbcc6c8b84d06febcaad4cea802f14f9100a6295731
zc480f201e95f37cb963e791fad9de74dc85de511945ec41fd6ff1bfc15c51de0c6eb02e11e6f68
ze1448e94c0fc5089fc105decf602b497e841d0695705a9614204074bb8e7feb06d147450ac7141
zb1d1830c821633644b17e0cc8cfa64b0401d0b27540b2cc245bb99e6fa54883b77d729d72b052e
za13f164737913057d9784ed07b1ccb8835c235a638a2a05fec640c233988dd1770bed74f2fbb8c
z0f1c75c24e9d4aaf47993374c354a215d1eef7fef7e57dcf15dfb65f835f5c8c2fb5255874dcdf
z613c065af343bc2103160e930adb6ae10cc926b3dbb62e20edd7aa042c9bc5266db217beb301d1
zd25a36b7d6db5822949870a46a371d66311a558f8c9c7d4111749b76a6fa939ac7ae3f39ed143f
z63ebb1fe2f4cfd18cc59ed52bab07484f47a9f26446d0c310f2e64a0b9090ee050092013525169
z805bc4961802c4faef8ad0560cbce0f96ff26f3580a2ce95a328135689ca94c6e35b4570e0b025
z0e1ebd11562e074a3e53bc949dc1c1d9ad36ab51e402ea7f0d5af53a397930760de3ec6f22226a
z4bbd75c0de351cff4c29b9702333907a4443b31c7757abe1ad9a26a572bf89a8cf6e71c4b329be
zaf7b0451d0cbf7279f0419d180b219ebb35ab85bf51b43792dc3d37cf974c890ee7daaab107939
z3eecff3b5602b6f9e030471f0e50794d9cdd642b0f9e1d759425db1bd15e43651ba0d664623d08
zb8683f0332369249845a04b057687c08290ea898c7b391b9768901d66847a5a3ab2a3ad944b57e
z2dc92089898038d76d955ce9d290814f4f8c4c760e1b54c9e8e5dda11554062e9f374c683bdc6d
zfca60e89a9af37ab18b3e8c07bc077e6efc155296fb4f9b89307d51359d1f3dc5e9b431a7fbd01
z92ee2c3d919a7af8a161640c310852fbb5c22bb137e2e65f3407779d03d9db6d85b24b19b92315
z96b31fdb2741d6c5e3b01d573da72c01d611087eac100ebf14c0f1dfb844489aeadc2c82a54bd3
z205f2828b7cda19619c6c73dc2742821fb7699
`end_protected_0in
`else
`ifdef MODEL_TECH
`include "qvl_pci_sub_monitor.mti.svp"
`endif // MODEL_TECH
`endif // encrypted_0in
