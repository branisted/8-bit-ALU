`ifdef encrypted_0in
`protected_0in
ze74c34e226135848fe16db9ffd31815111b6d7fb642c521a3f628cf6da949865580b22efd062a7
ze90adae0e65e66a2c36a587d0a790699166942afea5fb71013544a379d857e14682c5236087669
za040f2dbccbac59e8bb4ed6e90703eabc5da3fcb4cf9f80aa1298f4671fac620329c218c100101
zed6f713217a0741641167633de77ed77c2548cf70b6855633c380db97da98ee96bd521e19fff10
z0742589f83f1287fb5cb27df129bff148aa01abee5ab49e22511170fd96dff46c42a2423cac1da
zc3ceb4384b5198832c65e6b94b52b05b4487b3c735d6a007f05a329d81de71f6f0af02300ad959
z820755ac3bb2b166d010bf8bfdb8726b6a10a3e54ae6e789051bf1b87e86ef94d66538aa03da6d
z872502dd8e5c09af1526748a380d58259c52a2be1417f2224eea7574e4c3cf7da76c52b788f57b
zfb0006c6b9e2aa4d0ab6c54bbad65e202aab8b9234163c184166307cd81ec7c0c1a26398143578
z7e9bee7f42df35c319af4183f5a400a074d386ac2e0a2bf8855f12bd8ccc8e257b87f740006eb6
z31549d1bb749767b40703a8042aa7c7809a76a73547ff90ea233355614d4ff499308e2426fd8bc
z5b9081418146cb08fe1110fa8732194ca48dd3a4031f6c21cb94cfe63bb55ad6c496dfcc40aa39
z89e81482736ef3c0a1734ba94ee246087bf865249cf443767f6552f970ea9f085c2469fce13d20
z6e350d6f9c9f3576f5c188c4f019264336747603027703b8dfdce13bee506ba006dc89e1dd4d5a
zbba345d8401c694d8b9dac30a70c9c6f52c876ed5aa163beaa790993fe30105b49505dae1f4e4b
z15079a4e2633582922fe8bc280d2045f3c503d8e0bee7b2109e98e3528c23e87edeb04cdab76ec
z8f686dfdcf6dbb3c7bb28d022ba9e5a9e75ef6635b9ae86b67e250514e0532390b3c9eeed54bce
zd1827415d801576d9c80c20a2c33f621c2c8b30baa64876c747508fef5b6c6ad715c262beaf626
z71801981468e9f29a85c230f645996a10e53d2cbe097afecc50ef1eddb1b346060ea58a031e7ac
z9d4e6e9146b9963a2ae73025f0119592986c8ea20684e08262ac650c6e7ae82a12cc3a28b37edd
zbde9837c23fc5edfe72d861e1abcaf46ce4790c8679cf3a8a0052a520af291a96cedf219394c59
zd4d40f6b3faad0c5bde41c8a75a0b32b2fe7ebd18f1e34319fce69b85c712768225a0e54c99d61
z3f24d434a727846dffeb511f5f62f344d8e91b096b147a140377ca236dccf6256961a22c09b4ba
ze4016442d23581dce8428284c05a825c7a0a1ae1127ece8e081ad4fa0d9bb4f743fa5b5fa85575
zc4815404abf4248fbada016e84c59bb3498c1e5c35a2cdab84823e1a13e2def71058392fd82a27
zab9e87b5c1ef065203592f4513ce7bd33f88c8eb1734d0f371670e5cbee9d3c8003a64fc39f684
z08bafb38e021216a98f062209c148738e8f73b445f564ce5ab54d0e53ea1486494d3d5506cd10b
z5b03e3f125fc0da3c02872fbb45ff43ef7f5ddd7197681e97e25119c94ccbee35f11e02303b12a
z3ba6d6421569026556a257aaab0d7ec497a33b8979aefcf70126022316374391440004387718a4
z80675d0ecaa38d78ea61b825e6d36174b95f3516afb64649029700c82a8606206e66b2eb0ebdb8
z4b4f3b7c02fc8f2055c766815118f33e73a2c6d6d7119e60bf10a8867d45027be7deb60cfd6247
zf3092334e24a563b2bd82d14063a431a9cc24eb2aa32c50d8cddc245fefa185828a18800fd376a
z141b5460bf3b76fdc6f0e0d94598ff5bed0ce76e483d910ce72fcc62a5746713aba0325c7712e1
z56761a4291362acd5981fc3e5d7bfa5dad335dd6e772dc232c2c3dafb301cfe3016e91a9e4901a
zd53272cdea4e9d1b487bec5415793952851aedbafc22a4ab659de5c2531e3bf299d4808eaedf35
z683e96250a3368a7adfa6ea7245c144781d7003fa9bd2b76acda11f9fd3743b9c2aa405ec7deb4
zcdb8947a087322629355fc3c8358a53048e497e4b9d6b10faa0542065a39a6f0d1296c4c83e11d
z90a095479e86823cffe064e9027d2e2523f41f76115e70660f0f21868d9538acf142101c8427f5
z2c12cfc9d7e97bd8b019343394075b018c7cc38f8e1060d54f6799bf0853326afa48255b655180
zac92cbf01f6268d6aa980d20aa0aeef75639fa94ec0f3ebdb17aa976b32f31e43fa15ebd1bb599
z35f2bdc13a8f6133ff8c85e24583b6770f8b9888448af128a788a6b952754cc636b6ad215b9066
zf50957f8b2f262e15b96f052933f1f305615f86dbd5d40f3cd1dc5618d10435c27de9522617058
za698e26acc95839082a8e2709aba69362a9a3132344df6a1ed8d8f6e245a16e48bf6b2111f66df
zc13878aca91ba84e539ae8b31319104ba0c1bb090b29b1f309d5643d325bf129e453d7a39fe2bf
zea65cb59d50d1c9c4b81b677c038671142f2f9556ce2c597b8208002d2627e693c70d387b94e64
za7ce0cb7f86589028a766a1553a51ed323a1f1a60f74f5a2c1e2dd624249e5c68a226097de610a
zb1c65035f32ffad614d550344d63f12f4e0e11224a73e0d2eda653b86870f4d436a3f14f84472e
zce9bfdfc6956bc25876131306fbb96e7784889bcedbb845351678c3e5f916480a013c82e1bcf69
za813b8dbc195458fd04bf42938c94e2191a95ad3b369a2a42c49b808640d31e7c76de3daaa840e
z56e6f726a9ecd90e7403f4e22175b079e3533d231c074369703cad0ecacfd64481ed6c347171bc
z988de7721635a8942380eae51e98ac7a883c07df55a0b3962be8e3c54811baebd7fcf52a2c85f9
zf87ea70d407c8a66872ae4a77971f5935bfb9b5c44d6961748199a61adf55add7c6f3a4dae2a75
za2d93365864bcbf9029db5e326ebf998dbd5dbed77186b7839b34c7140246535a4ef45709a3963
z38e2a982448cdeccc2dc587833f705a276e25ae5409d323eb9a687c50e9ebd7ef6583b81e355f9
z9223fcf9a050938c06aa88b3d6443904a72b170c4d4e2672a065738901eb6cbc1d772cf43db105
zce6aac9814ce1497fe65e48f562f162bc0ad71b07f6017c215efcf4e94ae866efb9d74885d733b
z440efac35d9e138d2a59093344bec4a2a0f6a97b4e4ebdbf8cf80723314df99c5befcb0f0abbdb
zed8a274e1d2f0719c63ac25974c62778c26d646b14fb49ae0ae42cb366efc77c0a80656f2d7b98
z90e4240b25af9bad47d48bb4cc913028298dfe044e41f60db50af1105179fc3e99b78e0e51800f
ze6c3dd1353e81ad4a7c02fb29c3945463b2adcd8e7a215eec6308b8aa68c1f88df4b2fe04bf3a5
zd858b32d431a711cb17e930c319db026548c9e42f5ee2af026ea734eae4f43a84273839b002144
zfbb6cd2bde3d0468ea1d2bbe6323fae85098a73fce7280b1b934a01a4f922c4716838c06857961
zc1078a7da062146fe1719b076a723caccf9a8c70d2693528a8140fc0d8637643ea578d84b8213e
z8033a9de598dbfd14fd3c037a9e599b26238b99a6762514164aa53d22bb51f453eb14b82978d3e
z04cd9e3a688ba44c2475c3a1b7e6e91f50b7aa6304b12dddb73effc63f29604cf4f6569b3b7447
z557a767d04a84bfc944ab271662ec9e46f5afa64fbab9bc5e22f58c38f4967c897dc46b237f5a2
z48d48f27837acefc843bfaddb8b68784ebaecb251d2052bab3f82e6cde44bcd685d2113141aa02
z9ae30ad6a7541a0cb5d30bacf2072dfab165b06c4bce5205857c96db89b7df819e68c231d0f88a
z0aba008c15877ff3a691a43359cb150d8d3c82c7c328deee846c3c8d0f4b9814cdc817a3bb08d0
ze40c20b5953b7a8a0502c185e8ff70b23686c6078e3bfdbfdf7e90df316a003b35996b74fb9cd8
zf2e81c5850801903fcbd26300e3accabd5c58122ddc5ae16e819c6237299abe1875a849cbfd2c3
z7870613f450f4ffe38538f16e8e472a5ebcdd055eeb3a6bb209bb72fccba84b539d523dc8888bc
z075bf31d9f31d898b5b3e495f9273e31a4d716b04905eb4709804000b7085b10c5f4133a85cad7
z5a05daa3516d9220aabd030697057990b4ae873bc5d8f56df34a6a13c610dae1d87cbfc4ea4fb5
z688260b4d50f6ee09394a9973dc5e4ed86aca98d78878a039e91284186a0224038717429a370ca
z79823febb3b0142bf055ec47e98e13c3adab95086b0dafecf4bd514e2a546d5c5383e168cb9e72
z82bf47478648c1cddd17fb6d15561232088076ea608f19117d75aece133a3021a501e9928a7f59
z5b0559110461d888f7b495acd5469245ea614ef8d19a9e4b4eaf356bee671572ab29662969047a
z732a52fe7eb9d9c64a675b163550a2006ec4875c56c15e229efa7d75b6ad9a96b07d4b97b178ec
zed298a20e5e3edf4a19325b57b6e25bed9f1fd8dd524373f5504139a335f32517f34fc0a5bc46a
za2596eac4063793a41b2c6b286b6ac23e5e25744c69487b3072793aa80ac8bbf6f9883a3085a5b
z003fe5ebe76523820a13b08c64f4a0338d6e3f4dca0395ab93c7d571dd52f047f2b6570353243e
zd45f229f78c2cb24c32f496e5b7e1f63c79dd0f1fd43f814e45cfab6002393de96a228ac719c47
z7baf3b47aabd238a16711be42fd52e67e6355e7dc88c7f484cb594fae6f99d33a9bbd8a4355d75
z7f079e8fd37ff3f070d7bd41c249f4adf7a0cc7f7f648182189c03ffde007b8672a11de3b7acf6
z1681bd25db29910778c1bfad87842cdebd4e060a09c4f2925d2de09460c6b1176516e3dbb75f0b
z072bdcb830a9dfebdec2bf225a2242d653420f8e9f4c91384b6dc2c675d440d1cf855424211ee9
z64e7e9016817dbdd704407f0e68f6cb854113e4240dd3eb2f87e8cd225b0902521ddca8e6bc74b
zc000723f4036953997c96b27ba2f96feb1e0c55eb3fbb3dc797454006fc77e5e820889e9fbf9af
z808de40267a188448116bcb6fbcec19365922a7dac6508290e0f03c7c486790d02600c26b0fe85
zd9d6ed81df382fbffa3f52abe0df0f2a0d29b764240b1f038ab81baa114fee44722a1d2ae41903
z0c9dd6acfbb1a8b74fc45f7525def5bcf71007dfb94e7b617dc0aac608f5d9f83369e288f2ff84
z573bbed5b327b98a683a0cdc6c3f985cef2c4f389503cb7407813b8308134158957abcd175a1bc
z43bf63144e1f5dbb18947682c25ec40c65e97bffc224873ef7a5c139096fdd3d4d39b09075f9d3
za7fddbd1a24b8827f193ca5cea0d9c066fc05b4af92d52fbe1c982469721df55890cafdb172eaa
zadde9995067c0ce7b1ebfa0c973f140b04759538cf675bfc2fa8da67e493b1954f624ea490678a
zd83bc1a691e085de68410e1e213140ab481c28123e9239396ecd00786900b8c83f3ed95f9a7c34
z689c08865e9870952d13606b256423371bec11b33a92d0fa374572aba31f6fdb248d12d4a744c4
zeef9108cebcdd233cd9af51100c56b5810c27d94563b61a06d745f5693f9aefaae3b9730b6b711
z7c1073539dd9275d4624fd987eb2cf8795696db97adc8f69198ad00bb3cd283bb9a25cc28c7614
z7409e4ee6a23251dc1e99895b406d6920a633f6f1760410a0f0fc7df57d87cb9df7c1b410b3a4a
z30da035282e9adbf895b4f0825b85dde34a8b73987a4bb51d8ddbcfdb650b385a110439cfd67f6
z5f6a88717fbe8a46e49f8c4da1e9cb3f3ccb4832dbc237e1b86557b1ea8be0c5b04baac346fe8b
z3e1f33976e45bb236cd06d29d6aac3bf93d2eeb7808f8b1fa2f270f3f793d161c8e152c2d2cda6
z3de96ec02fb3f259b067210d472034dc2ac4e9f6eb36be7ba391c1cc26520c0d715309327f1df6
z7db4723f4116a3127d23e14326f94ac79746ef2ec02113aae123c8cf9d18f8f80c112b398906de
z645c37a0f7c8d4ea10d63aea9f117655f072372cb8d4695e43f2ca2a68ff158acc3f0fa713dcbf
z1f623bde3b4f8fa32b071b1bf6c806c3490f52bf237e4e118c361fbd0a3eaf633e9a8c96705ac6
z625933e3e4108eb202f67f94d76fcc7c7f9157221e35617b14f524aa9ccf9e83ff627860c2064c
z635b2d93de8550b81364d5c2bfbb2ef8d6737993e55d7df9332c866ab54f6d970af25d1b61dc50
z868b8a37ade1927f6931f27d45e07812bbd6cff827362db4dc9d3d4716204dd53bf75e95331a59
z8e6e319c0525e8e143dc9791234c94ccca69f6b93d39d095f714852a18adc097421e73f3eedc76
z30e0b66bdbfe88a9862b026782cc327ed6e8392d7164cdfb9e673e14f7b43e4c0b54bd8b970265
z85bb56a711881d2c308bdcb80f483d86d4fbdb7c1c955c21e738097cd76fee346fcc20937419fd
z883a738fb39b77bd1f3f566f0adbafb7e3546127a80efa5e5a006d4aa195122008009f0bad8fe6
z30e5a0fbd1006ae4d6655691f617b7fb40188a6367995b8b25917111f504dd4a06caf8de794872
z3df6758e381a16af4b7c0621edb97d7293ead8b86528118dbb1b0ba466515282e52bbcb4adb713
zad1f754dfb6becfba973a8e69e011fb10f2d9e6b18eed34c2b0bc3e003107f4fb1f94317831579
zd0d6c27100275cd0d3ea0a47a50b3a02b8d2d0f736fca6c7298e1fba3974f86efc0912fa3f29bf
z3a1685c2228fa02f0c64be301e36afd8cb35f79fc97365d32e9fe1fa3b40a008944077d2a45e80
z51a33357537aa92a77c60f805bd22c923d94e8fa8a9853e7c61ab7928e963bc1af48b470836fc4
z87a4338fc7fd8bc88646a86a376d6ac16ae7cf4ce68ba65dff5bb69d31bf88827ad15c855aef8f
z053c5e86735efd71ca72034596cdd79a04fe6d1e88c0a9e5736304b58265b1225c29000c5499c9
z3ecea3e60b1db253e8d8b7b6de81fc16a3612bcfe3d06c3117801462431e5ecdaa6ec764fe78fb
z89ed3abcefc51cefd0f4f480c71257e055552c97bb1ccce51ee4a45e1ebb2d00945627b3b309a5
z5ee72d336d6a2929c30e0f00c2298b46ff976b2962a0a862bb765c2abbde7e67efe8dc79528b71
z3b7794fe23d30cd237d09c0166164a113d0b0c4eaf442c79881351cf3dff94d6da1f9821463e29
zf58e41af310e5564fe910275aa388e54666ef4bd103aed70d8f818c804ee4ea4c093578cf9d888
z0bdd8bd7a7316ddb16c114e7a0a1b49f273192b350b582510be02b87ac05242d18bbdaa03cab9c
zc09ec87b4e2ab424a9c5e52b22dd32e222c4f370bb572b588b142bc790e3da76405c7fb3cfe2a3
ze8f9bc45d6c3979dadf45105039d50e728b238d5ab22a48cc9f27dd1bf3a65944ad9bc2ad58035
z77b53f13fa0a7365061285dc570553030b066988155c74366c1bc19dde5487316695a6e97f86f6
z8540016c551e6424058739d4f994a7caf827296b45ad4021f0d1ed56fd19f76ace750c293d3ae8
z60cac1d81e1ce68aee736b7f1fda66c5cdcc155ed3a93b3de825a96b00a615113deeaa7880fed5
zdcdcadc453c8dad3efedff1e6d299a9da23168097427f5dc176da83cc131d587bb20bd39f19f8f
zcbf84725deaa8d498d1b004488cb010eb7d8a96edf3f85ddae456943eccf0c9f70525ecbc00c4d
z6d025af4edeaac5f15c92de1f3677771c27410a7e8790103b87c4a15bdb950b31064d3648ec24b
z1eaac0c404c14fb82244b6a50a7e941def6cec6564b17730900a63fc9f25e1d376230d27709703
zc01b79087573c5d019a3934f42d1e3f14112312e8b6ca3ab80e1dcbf6edda540f6f7779572f0e8
z35437eacccb2f980f8a617e3b7df17d544d956af2249a40997dd7a12270bc7dca16378586afd0b
zdbe6ed88969020da0621aa653d368f4b16a9ed82df58a17a988bbc0bed47d53b3327d116503b10
z7b97468d8fffd28efe71ef43234537e3547efdcae1823624a1678cc757536f4a109bae28d448a7
z07146656d68d40b76c9c9d641f1638805bcb26be5aa0ebdb9fd813f4e7888fef21cdd18a3c18e3
z28791c008bf50b6b55ccba5b03be80d17008012b502d64dd36074331ae249db61a5c521a3927ce
z06af9c91c4e3c1316bf879d8c716efd2fef30b7eede91e2a1e0caa9c7619971ff9558c3dc9a78d
zee791194107e41f271f23504fd8607d944ed8985292932020dfc7e461a28a179c8df79eb34a3ca
zb71aa3d764e7f0b5725ee7eb7c09b123f710c295e8f207eb264454f7691b68d68ac02b4ef3c146
z3230dcd690fadfa2c657f60568db0953414ebbb733c8dd31b19306e8a5df1943e2c748a7b296f2
zc5b3a2ca6eedccbdb08ac6be7812d1c086c4a0238907897bff0fe6cf48c5b6fc1ddcd715d0cd52
z5587b769a527de228d773c877d3d8e659513c7282b9159cdd9c5e5ef61be4cd5730a8c7ce17508
z49e910e64cb203e69683c97afc02205b5c3cfac6bcee113fdf98157a68cd99bb2cbfe84f4aaf5f
z0eea657e600b839d29a117f9b5dac3a0cfac56dabbffeea608e510b3980328328ab0f0943f93e4
z18f95275428d0775dbf2297e7dca8b0b280210473650060f4cfd183fa6f4f8d09242db9795ba44
z4057e30588e34a81cd645dd67f53ec54202b6ccd66af4043b8820cb8bf7392fcf54db23d65f9c0
ze454a266fffa87bcfe1ed7cc64bf96998439eece6713cc1293ea5881ae6713d4864ee5fd7f3ac8
z8a8279a414e12d09ea42ea83c62b7b9cafa73f31ad425852c0b81cbb646c397f7517931fde8236
z3224d6796f47f6d293991fff0826919dbce8c22643d2d40b1d0643a1e97f2220c29fe1a19fd712
zc9a77b7a0ba07b8d49c1b080a8718b010967099c031c10a16aeb1f8332e0571af3b42e7ad9a186
z07be7160ce57848ec8176cea7d917655441e13662f20bd64b51dc9c3952d99b35f781ce8f88f43
z1763dfe17a812f8d87de9559a4b9040673e760831a51c745b780371ba8883fa2b22a7faa54cc0f
z8ccae959b1a1ca395adcecf5ee70fd055d2d3803879626259d4d3e20dd2f3831bc14504e6442c8
z8cc4f74340fdfec2aae89e5005cbd8042939465a22c1d98602d203e9adcac28fd868e4613e06fe
z0939fc6af729a7bfccd4f70066079f19cb46bf06f611bc32e5365ea2aaebe77ec77eafbc7b7b8b
zaf9cc21e8d681fe0e3fd5753037b26feac93c44efb0972af8a7efc8dec8a71d7b5831232db5ff0
zb5b96a530ae01d5b6a4fa1ebe895d98b199f7e2b40e417cf138dc695116d85f46ba642b20a1b85
zfa41fdede6e1ab52e31e36e64999ef689369f59d78d64dbf5427710423e8bb11dafddcb01398d0
z64abfcb5d8a5999c3eaa2beab3426cf1d12b813a801efbf05e3831878e253b94701647ec6b0ef8
z46f0279f90e080d485679897cab8265393a881fd34e271a0ee3b80d754c93b7042fb3f299064e9
z9933f63813d04a7ca867106f3e1eab6bf530aaa694c292d1c99393ad42f50589bb769a60b0d817
z45a1010100b82a1584dd87f8560b8bacb6ac8abafd06561e4cc91407a6a80575d7cd1e800765f5
z7dc2b25c92c0e0883d63dabcee64a60722196d590711baadd29cb29ced0180c253a2987f833cd7
zb393e34331853fb73a76b730bef7e753407a01aa42f029f3b1a63b216f65299d281b7b6f1d7c76
z55f1bd01a05dc690c68b4efc4a7e90edbfe18578d01501f9387d10c061c7fdcfc728a435a2b863
z1fe0809af22d6a278f8494389be01b30128ee51733ddcdfba7cbf92ff3469422a845d4d0987b3c
zaa27aa4153c9e7894d5269a4c17983a7f8c9c95ac64fdfbc939e4a86bd6a724bd7b572dfde1352
za50d497bdb01fa4d7f621f648ccc451b596442661b995b219160a595138e3d99511a9dcc82fa56
z3096084bca22c582fbe1ac6066bb78cc5517f30558c1db5ade15c1ec37e819b2811cc6bfc9266c
za9729022d64bcd38111548d6bd1be080df9a9d5f4332baad85a6800faa7fc3d39072672b5b0f9e
z62b308919e044062c1a1d1c460034d198bdd2bf852fef0c9cfd732b22829ce8508c07efe314aa9
z514241e7564a182e81b6d91455eb56d9e7ed720fd1d603d209c4933585812f5a727e7237dc99eb
z03cf7b79dca4c03d7463a408df2f8eb2830652a27e34d85ee658a506e149aba862ea77ed00c5b9
zf3bff9b49b1b6cb442eae8c8b64d31f8aa2b7edcdf8caf9043182c9ab7c9d7420965acdea63a94
z6e3a25edcecf1c891fa36cf3eae930cba0db8021ec1ea97d12b07f16a73d5d2b017000cac6f9be
z76a72ae4624c86e75b8f5ef0c3328f97e2ae905624cf9bff2688d2f4b1570ae70ab81e220e35d3
zc80266893f5bcb7d339d09085d794d751ebebee44c6ce05d3bd4d8db6240e2198196f858e71f96
zc2a565cf4ed2e3056c750a9a050967b8d713f54816c5effdc8a361f0d5c24b93bf84093fc9d201
z84741ac899f78123c785249f5f1d18f73022653202ffb6554108c545198f2b4635212658a2a02c
zc3d6131651ca87e6fc901596b3c07096994796f9f0b3d46764ea9b93c3bededd7c8b02f36a6e9f
z9a1cca854b434f77d4322c5da04b084c9c46d9ecde7bdfeb37e34b0f78cee37c22739738c1c3a2
zd0649bc1c2dd2b6d0f167d038b09e8b77f3a135bd4cf7c2d611a887457d5b568be1a861767f43d
z9b0590376f93394099e32bf48ac4f1cda9fb031ea3b08c1d64f85d1e55af33c7ba5fcecc3e9e43
zab2e319918dddec7d15c7e16e4bd382194fb585d4ddd906eb3bc123b6d816caf40a56c662e28c1
z00926c0ecac014e26473864d123a9880961baefd8c2ec5349ffacdbed52e18c919987f24039cd9
z8f43940e66a622b0e9aeca5b31ca4922a5c2de765c9308cb06fb1aec0fb0b86f84060edac29a77
zea932f4f1417d0d2d9d83966ba8aaf4ed7e8241fc44f5c5b96705787cf842b7adb15fbbb1550f6
z346a3868e1b1f60a92f63ab6296444023faa90272bdfce58a9831458eb21dd546d8acb35ff0e2a
z6bfa525d62dbacffe8276a1d7230fc7b467d8965f2344aeb13400df0cdba038cb302bce455d4e4
z169c804290280b5fa5db9f99f8929584fcbaacb3a5459a6c5ada53a0e24f26d1d5c71699f6db5c
zd782585d31e2843fbf7798d62d335d54da29561f404f85fc2565d7566844e5d03eaf345338b6da
z367dbacf3e6fa25d8b19ed11b86457eaea096adc6ca968acc7b1c18e910f4d752233364ef556f0
z43d66460dc0df25ed08a213625bda916dab2abf9ca8a2b6084898034a1b4e21d89982a0e30c17b
z562ebce3a52fb9f505215f3238c69a436798be0e6ab05798f3f54d6c4fae692b053cc721920f46
z54fb56ac2ee0f7769e7df756230dff207b9967e2b788e60d9a776334ae874d39ffdde0153e2d3c
z748266fd2136df2145f9dba4e805a11f70a364f04a37b8a1bd251e2a02a22171fcb5f2fdebbd93
z4332cc9b94ecd75bedc20875920175042feb841f7eb75b83b6b445f6093d57dec258db08d1ddb2
zd75c549f3011f93b3bd9fd59141e84c27eb06e28ff890925182fe0e7c0996af99f6543cefca426
zd17b889201d11312d60678d6a05136d01200db95f30adeaaa4a5260420833dba614c11a6386a32
z6a5006214bfdd9e59026251b11ee8f3ebede4724aeb83933da010001c3a629aaea3fc9722849bd
zec3d38f02b2266fb6a41a70ee283044b326abdc8d07728d65c94e0011c83e9e761e4e3f7676b5f
z44f934779add26201471718a30961ec72ca376e6ebf7e159b7a87ea218b3f21b2e6f885492b52b
zc421807b7cc14f6f595f4f91d20a6b6de2cf31d36a61959a4f9abfcb0afac97c76bb7afd053d4b
z39b4d492957e478f1a43088fa4c929e567f28a65c38d2abdad08b2f41fc15787f0a606a31cde06
zfeb73817b3a6b3a8558ff5267ee7b0ea048e2dc657a7d5b57114916d908437e305c1ad7f029798
ze9deffd837613a364801601961b945152b8da78b17d3fb4a7feab6c6da0c54694b49bb9c0ed10a
zfe42c3a4aadcbd749e2d2c7a1046c815a374c8e883ec4a452d35491652bbe25de36d3f13cd6968
z287faf0f960f6073afded3ddc968e098ab5d0df46eab8c8dbe46ec792df29e7ecc2da2fd617e90
zbd21e37d648a9f0557a6d7d2a94a67902d81518f3bf4f4b1b5ce0e08bc432b741c1d3ab5b354ab
z39b4aef91f156ce39ba1dc52e140e2a225a9a4d5d8f991939ff9e5617c02cae47b788b06b1049d
zc2746e543517ea9fe176c95eadbb683993a015498f1ba76777beb6db6512f5f5c986d2688d796e
ze4020b077b06b4948cfd37c6abec24e719067f1ce8af452322704f93396cd549802ea47a546550
z651e9b1451355174b2e3a1e655a2947d92a2f1fa9d3fc25e6192923a4a5fa72cb81806d68729cb
z3786e6f1164b632ed177016d3784133a03f2feec1a9f0e392dec22f48f3a6642641a55af22b2bc
z3377780fb36e801c49df0709d76a2b9a46bcffe26b1278a23ea7d6418f6d4422c8e73226fff193
z914585720775e1b4a9bae96fbc9127bcc63e4f54dd1effe508d11620ab4ab828eb33b819582357
z5fdb8ae93ff1307c6e11f5a33cf5d39275e2ba637cfc30f80f19f9c11c731cdfe14d0c7a4d4867
z9925dc3f17dc5c9127049288c2e965ea4f9e7bbfc6581c97c818d50409b2413ba1af6b9fed5bce
z5fb0eebfeb3e470846c4f55272ff03c5e3bbcdef8eda65b18df22eef4b643e2943bef33c2948e5
z7537559ac1618dedc0425bbaf74aaf8a8ae16c437631eec7aa8bc450686779d4eb58851f041dc7
z8f1ca8bfc3b9750f9736ec0bd2aa83c9f1af3da357503ae0425b1c9aa9f903cedf6fc7351c287f
z2bbae2ef405a9609ee7ab555d2cd9a49b50564f400d2d610f6bd60daaba6cc9aae01d71f51a4da
z95c44d0cae2b9ef0d70a2545a961e9b9cfd6ed97797be1e635c6bc3a0a157775cb92d75016e8b2
z92eccd9c8fddbc6669cb2ee5ba38f08cb7110faf90a2ea812c952a9325389b070d15bed35a9dd3
z1a9917871ee404512a4ea92b4c21d12114e160a7ebfff59b9f2a29b95a106e016f5004f0dec746
z5810f6e773c4b83862b5f84a34de34f2b011528b7f893fa5450b243aba6689828911d9a7af83d1
zdfcc4c0cbd247c353905deb8abf018d5c9c701880e481ccf252249a358ba8752a8b53062934c97
z5fd7bd22218788dffeb961e33ca24fe24b85c73775692baefb5ce6ac893d1a57058d56469a57e9
z5e763389844ba9ea87d6559b055019b86798ce894bacc2d852f7910ec4a0b6cbe3d93ebf897d8b
z6d8a3b98f259498a54a6866f13a2c218586be52c55ee39f1a7ed05545a6dc85776e4d9908d209c
z0a1a63a9d1c44e625c3364fcc487b583c21910b90ecb579070b6c4ac601a4259a893d6f5859c80
zd06873c05225d68dbe382c9410acdda4b2548eecaa389220f871fde9d35920b8d23e9e6125f4ab
z16f6e05d2ac67269c71476e0a42d3feda5e0929da2f18e44dce2f744f981e03a1e363c166e0791
zbc4b99e7664c1751a154b4a7145ba403de1e181543e9989347e00892c18e607f11c3386f72317b
zca432e6b72b9cfc9dc415c0743882adcc2d5ed595bd76e355de32c8efd35ef8c751cf27d8ce16b
z15ca914c613af9f3540a9976a54e831e404debc137c2494434d5646c424c17234b445f19e0264e
ze3ba2fe97b6461b1527ea630b796c7c0ba5809311a1d63f69127366451dc1f194a21202bb970b0
zeff2c2398988519e34002ccf15111e86ba557dab082c95a91d1c2dad394355e31d84d9af4c44a7
zd2255144d2e7724d243b15aeb961c1141cf9d219fbb16a82dd09640c8c8b41ea059e9bc048c06d
z51ab2292daa37404828483ee3503092a5ef05083ea1ca763fb65cef76eb1536b4e6afc52863d52
z9182dfde244ded8340db4f19978c4f717e59dec722fc733f15af3bbf8779099faaf2ceaae22f18
z6abf4d7894db689d0015fdf80e59cb8473e29025b3f99e2511867e690519fe08474daf20d31224
zff8edaef3bddc120505a26aba424d79577a78ebc356b916ae78694dfd60c3b91f4b94a7b72391d
zb703a00dad8dfa9bfe93f088b2fc303bb2d16b17045830bc8141a95caa39ddbce7ba9240611b58
z559e9f3939731369748d0043ff57495901d3d0d82db8baa287a76d8d683a050df035c3bfac63f8
ze125a14eff6dd8a916ee02f7f188574f0e743d3cfb05ed3543e536d770cc611b1ff2540093cb36
z749ba9ba88a8b06deb107f5cc8f77737b7a7fb121c60a36bc8824901c596086a170f9a93f6e1f5
z96a6b426fb7816cda8974bc2e3663ebef157f616db3cb12c5d6577431470f6f342312ad8dafd4b
ze9558e1fe409c03943c1cb77a2f889d21548835f7ea2420a36789f03ba6a6c2bfc8f527c03f30c
zeb9edd0dedbde6632d3b52c71323f692425160b6a2efcd09aa6dcf12f3019ce2df8a8cdc49eb7a
ze40381dce9af3cfd83cde468c8e541b639719729e8ce7992c52ecc4f39de80a016922caa9b5be9
z5c0ff6a159682ba5a18ca32c10baa9b6231005fbe3a2f3f554a0696c8874913e04fa70106a68de
z7ef5be50c30e542db375e165ab4e22c19aadb54072fe440c0fbb3abe6922ff98fff3442b2190a0
z95352c214351518306446f42744da2800b753b799499848c36ad4360cd4d7dc9229281b7543d36
z77dba62f3e46e9ae241c0bf1ee6893443ed0e41dabba72e051a6b50a8267821662154f045ca0b9
za725b8cdd81a23997e990d88c7d01f0e82d7c035d0eabdfad4b36cd891900373b50aafa720c149
ze44689f3233220531eadcc6688e377f46c9c3489ec45cfa23af3bea23923f6c8a8e8f0cf9fcd50
zc44802a810bdf8b9cc8ad01c3149870ed109ce1a0dca562f01627217dcbddcafe623d76170548c
z8fc0e9fe3ba641780abb817b4efeaef8d1062749c47cb0b0c7bace089d77d2ea6026f6a2955f32
z197136cdfb155a8dfa083be0e337776add880c93c8521f7c82dbea27aa0a6cbf01d7b030fd6271
zbd1acecbe777cf99d0a24c5ff5010565d885dfcb4b67f48f374cd5f5148e3f8cc30c66cab95133
z3b4ab4c60c4790455486c29070a87128db1007cd7a6500b3cedb24d36388d96c5b4a5dce13363c
z4a16f99e225dfdd3dc5650b0d8b694c54941b4b4cf1610fbce5a56e88dccb97626544d529daf1d
zc6c081fe37db22c63fe03123a90883c0b92432067b61486c4ca8ad9560baf016ff3396f20f7540
z621795f0b07b618b8a1b44eaaaee2fb1434ae4d0f88f268592febac80e7e7b660fe7b6b4f0ec59
z95dc66fbbcad1491004775474881d56118a0245c9537f6167e0503bc53a0d9b9d9e84b643dc12f
z7f7c67c6ad1dcdc317e781d963232a829f66eac5d31a462592bbc5921948d89794276180203679
zd831f21bf411768cd8268c75dfef9c979b3aaa46ce445c7948d3f9a6bfde66d7eab32f81cff3c2
z562aab5da12887a96584404cca5cdd1daac740fe1d02d26be060a0d7dc4d95a29947fca037ca79
zd772cc26a7742ef08e2cfa6a50be8c31ee270642cf9d74b3ffb04db98b5155f882d3531d0f826e
zb41ef1048681845723b51ef0ec13898763de1cee778d5199c277892ae04a2664291f221d4ebf93
z8581c31f45305776fc3966dee28837e34a15261d4af8a4cf319457e127b69526cfa8b6850c299d
zcd97d7e93317bacc0f95615c047dce5bd96f8a3d9d70c755d0bd3a1db9438a36d083641b9f95e2
z4203fb80faca720898713d8bc853271e3c6eec53c318c098c33a6f5fe76c50baa9cfc80065f513
z0f6ac547a53abce5a3d393a66efd6391e9d0fc4d5928daaa776ab81f5436edb92f5f190155e76c
zc62b88c8278fdf35c9c27a6cc21ac50d80b24effc9ccc260c763e1a512b966b07f5b9480d624d3
zd38ce83559167b130eefde1fc1f64eca1be7917eec18e40772811706b9f0184027948c2e164601
zadbb7191c2307114421325c3a3af059b9b3d87fba23e75328903c9fccd02d3b2aacedb776b6bbb
z6c44884dc3b81c29b06e43ed2e2dc2de90261b05415d14e47cf67b14e49b3a66571f75062c1a06
zad93fd75ab69bd46b467a5513b0c53c5707f13bc831c0bbc12184932538e86e5a00141b45fc9f3
zaf6685ed4109b6135bf20ab8f5c475bfe898364d36740a0417d370ca6afaf39187b151a1f83e01
za3dee966adbbc3e21e5848668269a43f27f4f0fb61887b809a75c9c6db054785c677e82148c8db
z64cf77640cbf699c98c204d01f8197d31bb4aab68a4af808e672dc885eddec60fa574ae957f86d
z3f0a2e5ae39461649896dd1042fef33b304f24ac9a338a20d91e30cf29429d9ecbf073123288d3
z1d0dd59ac52ef6fee23d17886a8a5a7a762479bbc56966f562386f84f84b37afe52085cad48f44
z11ed6ac560298ecf4ab1d26fdbe8eb5ebd37aac9844729e1b7c6ddefae78ffa11669209b68644b
z90c5baa8fc2c5a4749e86623b5d0edd6b58d371a007ceb9a606e73f8f01cd53ee650f4aa1a0104
z7784ffcf73c4e6a5b2981e0b8e3ac3631c9a2fed0d2733c9ee1349c51065e0f8a51c4d24eb2463
zc5caefbe8772d07fd89329f6e6adf6a090bf82bb5e4d1a8910177dde8fce2201fb197df1941343
z702a742a79bbce4c072bff3f497ee517a81e07ebbd12aad7b6da70744445c6b897b774b1a82494
zac1cc3ee26d59e02521f31117c87a51b796c29715ae209755978379911c275841bdf072511e5d0
zc5b0603bff88c3172d7f5a09e265098c97183f3485bc979081c7547239f2babb8a5b16d476e06f
z8f33241d584aa5f40096c3164f796079ab25a1d0a9f01c8aca88c1008d2f1874fe54113a172eb0
z9f26b75abc814911f9b7ca56966f5cc42f3e2a264a11d6b7499aca4522017bae675a8c608f21cd
z60e148bfc79629e32ae8f07b47d460729eeb88c63cb571aaa8e7dfb15a6c84dfb78057364d24e8
z3386e9b1d42b994513eef8ace4b7c82b2932f50f24dce1b155e8ca6f378c833e17074ebc21b418
z000b085735924946a31dccf82e5083c6695580c689a06cfde050173eeb53b35673f94801c0055c
z7cb646acbb944668241af2e26f226311a0fe1f3554a34861378b2eb357197452b4780eb653785f
zfdf8f80788de27f24a0ba15d5070a61ea0492399beae6e6246156e4b248ab9e37c144a10e12686
z9ff9b5d7bbe52d29eb63110ef32406f9becce76dca8496ee034479e1cf2aa43cabcbab960716a1
z0084f1c45041f0132f617db7e2f58b37ae4240263711738a10667c59ac5b912635650c826a5f43
ze72a2487d2a65cde08dd020e4717f1ac69c1b83badaffbab6f45a114cdef9ab66eef9c505c72b4
zcd9eef7ba435ddf82aeafe0523c792b684b82d2b818041cca93c856caf1d9a58138a3ca6ce4847
z0cb3ddf978ccb1f1c82b511128cb39471ee0982b239ebe9fac9ddc6aaa2ff9cfb41d630cd1edb4
z0627c739f5af09a3eeadec266ad35bf1abb71bc1c16073603cfea1630be36d8faf2bbe6dccd2d1
zba38c975ba1eff4ff466ecab2c65d73c71279e6a5581a618080ea3aa532dd5ff916e4fcf14c3eb
z715a34c6833619396eff3b6f2dd850958327d653896d1192340b6546203e9aa01bff5269897574
zcdce5b9882bc1aaa2b1a70bf499de6b2a2d752f6f38825e36f6db2874ed10a8c391df3fe3cf6b9
zd159c28a8ac83e2c96027b8d8f0c537fa7fc904bac893b80e89ab2eed77382551db8365f87c405
zf42146bac69bc4adba6067f6ae9de4659f44032cd62683a613fd5f3764bb4bf6839e739928eb0a
zeaf892342e7885bab0c17e17bed3eaddaef476ec9462451085551362c83bd027d2c6b1ec765068
za0414bf8f7ee5c82f2817da60c2b9f4b34959a6239f1a1016776412693c453e03d37d3cd0c2417
z060559c5890b77c72e66a840d45e532132e3ff7aaf32ae4a60cea1bb5883f7a5c1c08ebf5541fe
z403120419329e90f872957df0bcc85242a2595aef223b5718359cc251de32d76ab1f70b57497c1
zc0369e67931776d6ae1ee7455c12a50985a59add884921365542bbf886612b055a958483dff298
zd13f129d93f2cdb1db1498603b270d846ae1999e6f3b617d568e30c404dbbd7717dc204c87b523
z1a661fe5ea090f57f0921da69551baeb4d480946591f9c1eaa806a5c085dd660d7eef46ef5cc10
z436edc64d0c7aa05a7f6a7c84470e1a01f755b49aa6263d7f687c2ec029e546da104db1ed68bce
za7b798136281baa0298bd92910a9817fe2f71764910a1e5626a4449dffc6f78ab911f3815d21f2
z3a859f4921a947376c9fbf8c69edfe84c63654b41883a7a4904784aba6fdca084d8c708f32b5b0
ze34fc0b2f8fbe3dfb49c5a8e6096e1dfecc5d5c6e3b303fee6146bc5f5fd3408e0f59de19a68c6
z9ee980ba092ee3a05ca819b900d23b4e0a0505496ec37ce9fe66d5a12c473f9da1ee4f3805d31a
z362a26277a12b4c8f22b3fc95bd6ec746d0a1b390ab2dff7bebcfc43f48933ab1f955c1269eb90
z5fb58593df3a0aaaf25906d398d28f96843aacf53fb757a30e44d875a514e9132b26817b5b0ae1
zdaa65304e2f5c596a44a2c721fc7c70b717fd335989d06f88ec7dc0e8deceab59d814fe934b9b8
zfc557055249bea1f86f7735936509f20a7eef4b1e35a2ad14135b0e02fc8d42bef2a1e2bc74d48
za0b03f8534b3b745fd50e0ae54bfa7f86a4b0b1953bf0f29664b855c8f125ebaf74f79230dfa70
z178589963b0f0bb88a09a3d3d0db4628d0940a53b5eb95f7807de0ab86b50aa6d80dc8f63eaa5d
zd656aadd7f27e302f7b9cdad00e798db49aeda1864d130a552095d4b79f6290028300953c95579
zdcfdb3399e0cb4306a191b55b60c3755ce23ffa7788d5cb705eb5b13ac609abb5eab0cbfa2f6b4
z1046401f31d574a115f97f3b86aaa54d1c644a671feb61d1086272344aee9cc0ea349ba07c7a78
ze35e66d6c030e5c42873fad16c8baccc93ef5d7e101e548aaa5d6ce1279aafb29f3a95bbe49a33
zcfbfae4bd93ed7fd60c446c655b2b58c24ba188952f5157b07b08d901879b068b594049d43d712
z017949ded1e1423cd20aa5f7e83efa03061c29dc60060450655e39d37b77bc634ce5467e96d635
z033f773878737b3d89a94c2e0f11a4e26d52970da2d2f1cd032cb8a954d213374cc84f6e184366
z42c6db90a5b304fbade9ada5794e8e055c309df6eb91bf00cce193b4d562ee4dde3e592c594cf5
z9f7d59f5d305a0140e1a59691837e425fed97caf1585d4a296e5de98e439190173e88f67c1fd6f
z878287c67b70a3ef7c8a5743b18c96538ddeaf6e4edceaadd45f073a8580b61e16653429d63c36
zfbd7f02514c8c387130b552afe06cd7728f47d571ab08ffec52026631d53015e796ce374ce5094
z1ace4e17cafbceb8b8d58b5c620dee16ce91004fbda8cb7e105f65a8c9aead7bc94f6f4560f388
zab52254b6dd97a73e4ebbf4b9f3628a00e2effdb51032475471256a2f7489a79260eb51b187834
zfabe58cbc3ac751e83ae6f425657331aa4f7ec1ed8927d1d1258688d0f029f362c9be8964880f1
z157a5519f2dd5d609ad102ecdcc9997a9fc536b9f0add6608cc42084a023839f44f0bc98a3c184
z81b86c0edd7b4ded09e42b79620e74458ba376abf933118ac8cf1b501b67fe11ec56830d7e2a73
z53cb5aff91b20a023b057f006017353af210bf6333c0d32e1425d6421f7efb40fd2b277e5f1d63
ze5e3129ccc41b1ff11e957f079239b306b60680924725ed85b16fc727dbd43d80ae62f97ceb1f0
zafc840a994cd05fa4819f977850a8bc3b76ec37aeecd7759de1a5bbb0883b03ca0358d1ece5431
z8b776c15f987a673901e99c03e200919755e5e0b2065d4f617130aa75d9c364afe8aaffb8be893
zf6899a5a6e6c5784556222cfb0eb4e61da2c6c204d27892add004046d393d84859a2ae5c3933b0
z84fd9676b559a3e7eedee97442f3e8626ef0cefe5dffbebeba390492d6f24b818fd21bf96e56cb
zc1302fcdb889e07cc77fb94cf1a06b683f7a7c57ba55d5c46848b642fb79688dab97ae6ef8b82d
z8ecd4be6b5a65fb3c06b0bbe30ab6242ee2a855957b18ccfb3526ab819fba25ff9bc4fce18b36b
z6b237c22c6aa8c183aea8946a35ddcd302ed9335caddcca02410681e23b09cd4c83673969ebd5b
ze8047d5c01f7374df6ce219c4fca63cbf7bc079d572cd5742f94a078cad5fcb25d0e52a72c6efc
z11c876b93aa568062efa1db68c057bfeb3ede422d85dc64b556d6b01b0ac9f4f1a0c46e3ea0b7e
zec3ff4cfe00f19ef52ecbf8c4fa78cfa37083d6db77711eca2490cfca57936cb81cd4926903c29
za154ee43c271da7080e5f22e606dc6f6ff6fc6946963a0eb44f9261ff0985e1e9983c800e5d7c6
z9ebc28807a2e9be58a4fa91f3d9096c5e3e32851d9aec78e943b75e40c7b02cf896ad990c10c02
z3ef388a696e79cb1ef598aa9e73c84be90d2c87dabe45c10eae3dcff78301d5d73dc5542424f03
z86cbb3bc26b9cf16d40b785d2d94ee7768830d2c247e0089b438e0fb07ed6085550f72aad89bb2
z00ead960f29b1f29cb23da4818f70846095224fc777e7f4ffc50939f9bfd4d2e7cf9242dacbbd8
zec7d9eb75c642f3c71ec7f5e5ce62f327a75e15b9bc6ff9f187f4f9dff4cfa93a6bc72b896651c
z96f0f79cd5c83d0bf5102364715b31bdc90847084e869bb073adb9cda7b26d421835e90d6287de
z149e37985cd16a06c0729fe60f9d1538b993750046ce56165f4e7e355e2b4442a5e06e8e0912eb
z73176ab6f483813eb401498bb673df498266e389ca646552b6f24dc05f527753c961bc0b18a2e2
z20107dcfcd5c5a43a2d3463326ab011bda210adf5ce8422a2a79b148242a29e7d5f0b73b9623af
zb4c4e2dd6d20691985ba22b78e862a518fd7f331c06bdf4fdc247ac1f10b13da535227c4c57a56
zf4e886f01094998e5b3ba7e4ec83f9ebc46d939e5c27e2be54c33badec3b9f99a4a5fd68736a77
z0bdc59e8a5b6178b58fbb23a2de9c3366c1e3cb3f18d40bdce1eeb05757ec71537808ff92c388e
zb8f29fff9894ec804270cea4b9315f076c17088845223faa3df58f1aad684412edc38186cb1234
z6c27be08e939ed68b56f7407b38a6da3592d45c1e10a5536ca760863509f9921244f499efb9362
z7765e8146048351a334ad76512d104373ec74e607af0ceda6ef7eb9de07efe67936524f2265128
zb5df6df82949b38d86ca74c42d1c903d8f8b69f57ba646a6912f7221ea6c6e117a96ba60a6f94e
ze7c4f9ee048d0ec60b56bdcce38a343b9959d6efed236b9bc659901ae301552c2f3d006c49b439
ze76ff11b8eb7fcf13e29191a879a735eb8dd69e67bff38af0f95066b6575ff243f3710fbc3141a
z7f4402a66da01743d673e70e72c0536b7e851e2832c3f295df331f0c598af09a9179cdad016cc7
z68d43bb4485da147274fea19656c942537217a8f963654358c5c07ad5253ec9a199d0cd099fe2f
z5abb341475b282fd7643310fb8f6b48341eeacb91251c70e9fe49484bc2fc36bbfdfde45be6ba7
z6a22
`end_protected_0in
`else
`ifdef MODEL_TECH
`include "qvl_amba3_apb_logic.mti.svp"
`endif // MODEL_TECH
`endif // encrypted_0in
