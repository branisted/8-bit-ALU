module output_register (...);
// TODO: Implement output register
endmodule