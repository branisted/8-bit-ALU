`ifdef encrypted_0in
`protected_0in
ze74c34e226135848fe16db9ffd31815111b6d7fb642c521a3f628cf6da949865580b22efd062a7
ze90adae0e65e66a2c36a587d0a790699161455169ed55a01f2084f11770a774ec4c588039b380f
z6de9c5084882a40b79a175f5c2114b2b6d78b070cb806e1c0aa9258297f4687ab308bc470f0040
zb0b1de382961eeeaf2e279e1462520fc31c119af8f2b214846f56c2b3cd2eadbe4099496abff18
z15cec83ec4a77b868344aa20ba7360908f5c0de2a79abf8b3534b883bb12180f68b5d4beb444cf
z3fba8f13afb0abfe8fcc4294810f75afe452434d2d0f1166236c82f76edf1e12979f04bc35693e
z32ae028996dd85737a8f5adc1ebb94f39c940246e887647b64782cd7ab429b0544c173176cede7
z01dfb26b1f73408344a52b7e1f117f12bb9c8077b34876c2e6fdc085981637012dc9754765e1a9
zc512ce062e0b8fb16a214591f5c81e1353b900a611fe1f4886b57940b41b7f2ce99a7b84b04b90
z916f717e73bd10589c81e207ed77ec660a8cbed5b487fa50acde1b055c8870bd8676023f21ddcf
z9c98cc47cfa2d654ff1365d1f45035a045a66c5dfa8279050262529d2cac9e64fd27d9c7de62a7
z731bc808811ded9016570962244887f98fe5440167bd0088f2f049df882af501358497c3b28776
zcdc5426c7f52a851c35106bb93e16fff984784050fc808fad15da330f6f0607eda2d0e0e4b1215
z2ac5b11453f6b6c5c6b428261a64553d70b4ab9f1bc235c2ceff4f6e3b1ebe72fceb7af9adc96a
z694b4bad7241bfbe775016041d7caaa74d9c0e7b507ce89e8b01980415bfa35a8e346f54c548f9
zda8767c02ea87d27eb7a843f4cada7dc3b575fb5cede69da7a4701b2d725c73f1f7375e85a74e2
zdeae70c30f1127407402c955b283d7b9512dbb3cc85aff97f613d57a4efe57b3c092e5ccc5b6dc
zd04e277cea6810165bcacbe3f515b3d75051fbe8fa4af7e932d60d2b2a6cbc14783b996db7f97f
z0df4e054ec07012afe312c7c27fe5855e396fca2df20ec96282aa187aefef584e73225c3183714
z599297effba6810dbfe57acb29d5b025ac9a8ebc73f537d2977dc34b086017b79e71d435e90724
z58f8859c47b62c6b1fbee0ff19f88a66a8afa79b5c1920e87193650fc0cd3c6ab3d109ee7dddc7
z162107ca701eaf77ce18df51d1be11c0dd907a4d1366d43e0990f506187b3d9bd054ff243db092
ze701807474479b37f0911dfeb69e92838265d0284967e78f0d2051699430d6e5af93353f8a4ae7
z1c7984e0af29da5cd55d0e97dfcb42d4a71e64e6191520cec069152d02ad57291a620e755a98df
z6fa6dc8485546bbd2af18bf3cfd459437fbf0fdf80856bb76e4134572651e5be5debc0ba0a422d
zb22a56d6375c212b53f403b92b101660c31f60ef55e0f523e3c42b1912d207d2847c2d5f589467
zb0564bd25382cf356e2b913bffb723d2a5947deb138b8f58e3164cf9c4536c5892ee1fad6f37c3
zf49e4f9fb4f807a15d5e745c3f36ba39323eec5fc71ffe9c2295923faef30146512219c34eeaa2
ze903728229aed1a8bc81e80c910e5131f227aada86d0fa97e4d3c6af172ae7e3a4479e0b9c3835
z556c3569f38259c3c670e22a48b54dfb26ef9250cb604c9b079daf97d1dc43aff8ae811562452d
zcf99153f09c65607b271708ca9ec33d8f8641a84018c6332c9dc818e1152f45e185f5b2e1d9c60
z428626d8eb497945347ea0cfd65584a9fabf3e90d71649d944747ce8240898e92b34b704c418b3
z9207fa71d717e856dc72af751fd48c8b7a9bd999cc7ec6b8c3b2410a7a27e23494f36fe16a0129
zfed2528513fe2e7490a18f16dd18c6994f168ff9c1618ed1988ee35d7deb7d5f15e355ae572a4a
z8e34d5025d83e2ea4cbebd6ec5786aebb644f9a6eba714c39ab93986fa7bd07f3689763583a8fe
z2e52801874d0ab142a097ac722e5b21300004390198a0dac74bef2bd5a27a6dbd462ee7b52e333
z829265f172e2c947f6dec69cb02e490e49a6c72cf7541105357f59321cab4e3773a743ae7e12ee
zd5d9f6412f04fe26ce6a9894e1036938ae433dcb5494c814bb96dddfd7fd33e3746d40e1b3722f
z30578e0b8fc2d2f06b6afbbb7118872d75168aafb1ab995143bd13c6d0ac0a2fbf2fc5782b7970
z74735fb329bc35cd00ab488910cdba03e3534c11ff83920036bb0ef93e90aed700f5a212617bd9
z68c7106f4388f1224bd75a9d69765adef3f8da78462a0b9c4b55bccc8e0d69c7cfc9d40a034172
z65a07251c15285db4dfbe801c5585579eeac3766b70cfefe6b69d91a19056d1dcd2a14936d6761
z9a11cb2ea5e5c724490838a1a3331e459affc2f94d92fcfbf7d165b7e8bc2d7773887a9a66578c
z8d62ce5a77f35986542e53161921ce04b10e6c96048c00c610181eebe453e4552b8f44dc7948a2
z82de69e6189b77f52b79a0a0aecdc279dbbb95236b287e761590e4a0cac63515fad87bc1b94a76
z381580a7734cf4667d987397bba088780906ede296645cead64fa79c18a3c6453680652ad248d0
z038edbcced476747700ef83d0c3d57016b28203c727dcc4fe3163f6c156f7e66fab1a46d15f16e
z10ee88ce8e97b69399942d5f512bcbefff7203df87dd54287414daff5e915969990931082adfac
zf78ed2e45c6cf0983d59856ac92b1bce7c7de2db6254eb72229622d00109160a589c27cba58fcc
z57d8cd5436bd051fc117e9379a67b9c829091ec3263b33f1e4a2983693a66d66f906de10836d4c
zd5f3a1b7e6936ee45fff84fae7bb345ff41d1bc7cb41c0f741a5885225573eb757bf231f8c9ad1
zbcf70df8a6e22a4da296929310bbca371db5f6695a5a3b791c63ccee5846fab75d34316a8fa953
zad49ba43dafe5544467ad38225dd11313e0037609c764b85ff81816a05e8a41937ce1bf815a7ba
zff00441fed9a20ee1d3414c6739ea4d8b4593f8b57d3c6d780969a05f4517e9b371eeec4213c43
z2d9534e648866d9fddc97ae6823777c3b5dbbca8d131938f7b6796c8c241371876c271cfec8fed
zcf8247e43fae9d3308fcdefdcce7b7577c0a1c140c662b746a1af2db53190c49e08da867e7c52b
z70c45fdf7b5d224b2aa9a4c0b14bbf885a6151a0ad0834f9af7f92cb30da0fd25e98bcac87e9b3
zef050b573515f38278ef1268422acde306874d417ce98f140a7b0117416a933a60542458823db9
z8481833524f1964ed458e2c1f5bee0575ffe579761a47be700eb640a97ebae5a38c7d998e5d1f5
zde576d4c5c31cbf8e05fe2d6fe1e6fe7ef683d4c51dbc39ba3bd17de828ed6463e96db3c2501be
z1fbe690541615ebaa36340157d5bf08bc8c32a9e08074c67709d64fca14d843b3bf567c20bcd3d
z0a899acafeee65cadbb4d763377fe04d2286cb71d3de7ff25934f356cbdab6ae006fa766cec986
ze7804b447e8772c68b50e7076c1862fd7d2df121b7cd96ae60f892999cbb803f68fa1f3a4731e5
zf2c9dfea0777d74d64525425f6338bbca0a69682c68b346e893f3f09340aadb82d721605559aec
z20a3c27e35dd66f74852dbe0c6f6500ab0ac6e6748a00d514048a15fc2004a0a34ee6dc953da5e
z30b208567c30760e8e90146ea87c1308efec76a2485a6f611c5b7ebfce6f3a8a85c00b646405d2
za44a3463a71b12f94c97c8d9017529fb3108b2f176f692ef2cb32a8e45191fcc67293f2b11efc3
za7f2c307719340d42f5a0d0e94847a3c57f2b8818437b72c8d021599cb37400ab8a23465b7df62
za43a874d5706d14c84a399ac6ca3b2c7cdb4843385c8304ad1f35c3cb64dafdbe393103489c25e
ze573a8ca784ad8a6216d5ae2618a8b34245b076e1650fd534f78079bb241c843673f73169e8cba
zd6ab643fd85cf633433e1a083268aeafef84050027e9d746606c5db94ecb0b30dcc95337fc59db
z1078abe413771d680780f93cd1a657c49f86f76cf9ae365a7fba0af03c6e408c70f4ff6bd7d5ce
z83b63acab84775fb547d2336180bc850fd8e2c76ae38c46329ad141f5361220464ab8b6be92822
z28c7ca4ea48368f4ea80b99ce7e8fd6fc73f0b0898ab278dc9292ef5c716adc6a1df4742d5ebe3
zb442b605504e7b7842212014907ef5baa8a13ba82a1c23bb1e61423e645fb7d1eacd4154735a7e
z8c76aa00d63acb07c2b122621a0dc6db51e8737b77a32f90a172f111d045238010fd5f12f8aa04
z1d3083131867cdfa3ceea2f5949f08e2b3f34cc93a5b4cfa38906bf871c8352375d0502c1491e8
z2608f684cfd2d3ca5fb5101a36a0d640215f98c70228577e59c1283a23a41268dd979c6b978829
z4da777c7c57978ed33d758fc8fbe2c0271efb73ff562b63f2853c9d99bf6777ea21536ca1c7df7
z3d28332cc6d435b45c9d20b6c44e1ff9998deb40b189a33fb7ef3aa89766f6bf6138c6c79411cf
z8dfba846a6f443b44767a6cf849cba4a10c672a5821883dcd476342b8f6ca26d5c341a808d36ad
z5dc40998192336e5f583eca44711cfcfef4ddc016dc91e06ddd68fcc4cc18d51a132e7c1a97087
z0cd28202a4071a73a4bf5ff2a1b0ff151c7b5afa14caa3ea6336a10b14448fe78dac0061437fab
z532acc482fb43a6e7f2f2b9dbb05480f424a84306c90960033e935690699aeb23257c8bc6e21a7
z4aaf9ac8776c0365bf45c945aac07f796a1586f053842ee003f3d85b8297d83045c3b1a367e9cb
zf7288cecf9ec4ad3b84c6bb2c7bccffc0e72974a8e02f8a0323064f40537e51279c19f717d509f
z9975850aa70afcdaf96c89b6a6a57171b618700df24d7507a46d45448a1d2a16d5f01077826fc7
zc716e80f8cb4cd1330a1d9acc2e79c95e2cb0d88adc11f596eb38b97c28463a8ef1da2d240ee77
z9a7d82d6e095be5512d317eeeac636b833c5a5523ac1b3c9374d7bf7948f896694a7aa484eb897
z47197c0d4c0ada48b36a4c7269f0c335916a880da3d1b432a3ae31b421e76565ae310ad516c92a
z23f1c9197b81ec079e8ca9230ee25b1a7dbdecbc0bd27e0e3ea7b00d80456230932ab6dc423c51
za50baa46fa404e638205b56bb59edd69b7ae096c9489a1171c9a133da0b4e2babb3f54d3e00674
z5eb2aabe5c6a2cd02dbaba6f4dca7a1ac92719df7e3c602cd55ad207152e30fdba93d522d3ad02
zff63e1cd81d8e6b65b7ffbb95b992b1e00b106b9bd1252549ecb1df86a227075b5438b4cdd7b45
z0c2dcab3e93ffa00c7d50c774861933c6c46bcf53a22823a4ed8687cfcbfa22bfa4917c1da680f
zbcbf584decffb5c6b9182f01ced4264863b84ae6c31858070be7dedc4f25e9238a339940af71c5
z470e8e0d310025bff9d422a116b84d43a2e8fbed2a69ab26a57568241f0efc9cb53ed31031a069
zea7ac4300a0ce1890effb1048310276337d3f8cfe0ecb7e09e9589efbe402984d7224a2ea53edc
z5ab9d0583300e781bcb915d404b6a4569bced59ac68f52cb3e12056be1b07ec47d17b255105ad3
z8b28d8948fce7d5c86aaeb0f22f27a73db578de32949181b54aa5afd131f4a40c02cdd87682e06
z80b8d8632c8b2503f353c5b3109eeedc19cf9726e61f190aa80f4b2eeb9dd7481f528470708b05
z158e71e6c49bd34fa55e395c98edee8330755ede36fd57caac89845d9d699f9375e1a9d0cda7b7
z68cd0582ac08583da59ee486d8cee55f25911bfc388c0dea71289c49e5228e7f5c8ef2c653a711
z41dc27edc69d64e975fbe6345148c187d3c4c41a3798221c2f1480488b8d36b3c1b20c4d41d71b
z893cf786926fa28b69a67f4dbcb28dd8c2d2695c496f2ee76ba65748e425b3a3c6d8b260293914
z3a0ad7990ca5333f2631806cc88640d6de3e01fc784cefc7a40c5a73a1d5aa31fed455bec2aca1
zd361f9d3ce532b217db54386cdb27be5ba03c680c768e59dbaf807444105e5660fc364802d072b
z898e33d9ed38f55c59092706511a8b68ab6f46eadfae0f84bc866680ee3071f6fca838b282546c
z22625c84823a42e52f177c550fc6eeb6eb54f3dd1e6a4b3c88bdadbe736ff63ed19d39afea3824
zb2404007e8da2223f6ac289383d3f8b14e439fec1aa68652b6791d30ed2e13693202031a881e11
z2e93035601daa40d0bdce40837e57a4e720926dc34282a02f34b4833aff736e7b59b5650c04630
zd3b954df6ff25f7620af52f2a48162ac69882b0276f00124dae2a6377d0be46aaa9014df720206
z78caa9404edb81e7b6cba43feddc348231beeaee9e7155047a64000f345f6e49a1388b7b402f62
z44e6d673bc9333560f6f46adcb8883e0c616bddcab694991b9717ed1451a2d8eab8dcf8795b842
z0d4e5d305287ebbf57829df9e566d8483fac4ac0ae39bb95054fe1be5edb6d59a8ac1b04885b82
zb56d4f671a26ba5de8da412571b182806d64444c2a2852794d4ea21c187edd6902d5887e703b73
z7b582acbc30efac6a120e7dcc73bcac762f439bc46a1914e00ac581434f042e518a5940d146720
z523fae619b6335402903ce9542a4360f76964feb89de4306c95abe7035fdb0132a12dc2ac9adc4
zc28b9fb64ab276cc06b2958e8612b18174d2d7a3aad7d7ef682157cfaab6fa1d8a077476d7ae57
zeffb2766f3b857a51d6efb3b2edca1b46af13d0db22cec317fbefc8d2e5436949d7315f90d179e
za3758e48deb4f09bfb84b23e66c5a310f324208d924eb5b1c49a51e8da49ef6f39859179f3c303
z64d8c8ef39cb97a115028699ba1b12813bcc302497eb0ce31e0334f061f4e209ba110b6e475b0f
z9617d59cace5b6c39182ddebeaf30284872973487c8584fdd469127d30e0f95e479100817fc6cf
z1dfc4db5f81e4a4b9daab27bca1705ddb5888347a470163778d0ee1ccf970472a08ae0934cbcbe
z2a6265b3f6f15376a9b024df3885aebab2a95db585022b672070bb97ba811833a62ef674c0953e
z89fcfa166b3ff225dc4025c4d923710b91559aa46c5f95c85aa3f64ca0adcae604b4b5318d5c65
z848ee258303cff54462d95535154d0c923c5e0622dd728ddb468212d7f7ad3e22ccc3c28e62575
z221243ab4addec43f67401fc00361ea1ac13ff1920524044c5db8bb790804ab291b2c62dd937f9
z41516f39e7fb3119fda0b6f0ff7f324450109c1af274bc099000ccd51ab7c1f63754114e47f1e4
zf96ac20b78cfa1897aa062d58bbf064afc70bae827abbf3bff6a51470d7c2ceca0578c2642c72f
ze6b0eae0184d9240bbc6b98595ef14488892469bec894ba5e695d855ebf6396982f3f3f75d4533
z92fb988d675fe48afaa5c51463898ea528539ec7608de947894f415f372dbacf89c51430a26e21
z9d98813b45bdadd025c11a3fc6a3bbff59fe5ad794055998efe114ef1cba32c1a9fbec8294ab4c
z72ddacfc3d40bb68d3e47045ad229945754fc814fcbeaac75b0b135cde3dbf799e8fb545d0db02
zf8f3440a0bdb4f18fd37fc921097256b1f80c97d441469ec9147ba2765ecc3b02584c6956e1a72
z3bddb0b333ffd515d7b34fac57bb11ec4fa343aa635d769f2c12bdc0f6f6abc1d840110c90a87f
zaef793e7854bdefa53ff8ba36f30e7b8ccf0c6c9dec10b8fc2222bb03f66e95347b05835c64f05
zc6b7109b8df12fb44db4403bd8f17a97434b5828d9ec8b01c3c551b32c25a1ce91937e7c74adbf
z829558767cceb1753758477e03af8b7b172d23baa7d62d1486faa801506cadb42127bbb48fb74c
z5bf94cae589a1644cae6fe5a111d63d62067d32a652d41e59df03158a61c6f77f09662a65101ab
zc146ff744a1ea10ae283c83888a43698e13033947fdc3636790803683d6f632fd254401a3ef258
z7a98257393ea95907447012270937242f51795015191658254e418735e5b205b346c7557c7857b
z926e541cd872ef18dda286ce7c6c1a6805e14beada2c53c0251caf3eaa68f582562979a467aeff
ze73ccca4b9253631aef6f99144ea0536ad9a150246fc6c7c8cdb936eefcd22cabb2cf2037a6910
zbc1ad6c30400aa4004c8418b02c496fecffb36d1b569b09fcf874df9c3b885dd8bc0b1b418d7b8
z12beed59c4d0a094c0ec1e0f0ce9ad6ec9926d9c0686f8772c9afe9a40a94e2f1d59c2e423668a
z2e385a3e1f11e7400343d92f3b4ae14c8426ab684e0cdaf8514a7bebcd2da6ac8488ce1006db90
z8f9b42ff285a025393028dfbcb72abdcd27c30ee8695d3b361476541e1ce2c03b97b075885dddf
ze647492aff784e210dd05fbd1405e557a0a0b547fd0925847298a1d7d09c7333d19c377966653f
zd59804040140da467a156ee6d1be5892b9ab85dceeab76f2370304ce0de4d84242ed2c236429e6
zf97aba9f304ca2140626c20efaac593c6d153056586092e1a765f901268208039cdc8bf736173c
zc7bc0da36c4e125a1b141d4f3ed2a600a568f75678b22c7174913572a17309eea36d48b15ff27d
z5c6cd91c860876dc96665644ff01e52044fa4e7019d300e686a2e4345ee7b5456e7639d4d81a84
z9bd1e65fd1965254cb441956e9230bac74bde7dae9551b2b384b93b771f08163aa53dabb317f2c
z06710e31c073fe37d2b3026c9cdee306157b2d625c844879ea9ef5afa4c8a360ea3874bab8add3
ze96f5c1bdc066ddc4a2b986b80c81c64bcfd2ad80a9ffd48aa6e5d996f5a67eb18081dac1d46f4
zfa3d8bb7822df986606b62247135ad36b981fa0d82cc758adcf714884425ddb33f4c76ae275815
z3822cf62407a420d30310012388ec3429d610da6ad9e2e765833b0fcc21c78224b81d13276d924
zb7d3af7745d049fee6532f8e752a4054283f5bb78c1f41a3a3df0dac217df3eb396459f7ffc809
zf8e5920f59b2a226dec5cce1c7df68b8902ae9562dee0b510c03d7b29548aef604ad9112d393ae
zadedac0ec0a9d15e2a9e6c060626c7653db575fcddad2d05c8c8dcf7a2ce664510a782a0d8c6ba
za6764896dde932e6b36e2ed4f8ac79ef692a72976c607035bd8ebe592fad6a3ce518b95ba81fcd
zea2040ed2ce62c2dee6deb9c7725731a0d33e1a7f98adf560aac45108a6201a3aee8ac2da4101d
zd5a9c9943ed3f12784e5ad4dfeb64d74ab0b0e528caca27c4831a85461bfc85a2e2e4fb9add0c8
z926dfe3bf7c7ab8a70ca5c11fd32ce8a7556b21e4a5eb2885af495852a67294390627752c45348
z8940c47366e060d62fa41f8031f7b6d4a1033ba07b4f41c6688d3f84be37b23c87cc2918dca73d
zd3fa55131f8a5ed0e1eadff6c46d55f17b7145725eda6fba34724ae130319c1a3348bc0c154930
z722bb0afe286eabff3ac0f6aae4b881805df93cad2dc2344d18928b90d717d9f2215d49d15bed2
z591820553396cf3bc1a9be0c6986c7e6328e272aa465a6a3ebef8ddf718d97d124c14461f58784
z7cf53e6c1b132b14dda0e67ce557e0935c826a06c12bf16cc8923d04e5943692a8b584b5e76cd5
z9b4310f143c2cedd96ecc1c19946e4276212e282bdf9e36a2d38063175f3fc3630416de9573182
z247c9b5b661a16a8300489c3960ef9aada1f7523fcb321312391c20360de9304837eb6a5885559
z8d2220b8fcfb53e5ecb2104406614af8ec6cf0e6e5d5ccb07bb1a9f7f0ef3215c41246450b932c
zbd03df5835c8f88848fa952b3efcb04d42e0d0bf0730f4188642c659b8cc579630c4b5e6623eaa
z536a8de5c4aac0571e1dbec7246f1b54be19bd8f5d393b2712e621c19dc41dd0201eaf47736837
z7de694f8f6c31648fea8733e40918758ccb96234e6413219b5f752a19bb4492de01aa460b57950
z36105119ed7707fe4e5fb22fe75b35508569afb299ac521e7a941ddb971b3aef5a9a5ca7e83ac2
z7bf3807d6336d24402f0ab79b39d5f6dead757171d19f508a7796fd83233b61334433713f40e57
z987cfe1272f57a6ebeaaf388b23e22abfca37a92ba6de40f3c3c2672039309e24040a17a3ab43c
z867f5e7fabb21abedbb39cb7c6d782fa6fea16b88c20de3255839772fbb5113eb14419f184f696
z732e20f0970583a1f6b7847b59ec30b4dd86e597d83f7ebba9613a9e44f5f9136ed468316f3678
zfdf9da76b2f56bbb594343c130156ee4fdb3f8b7a132977dc62065493ec0755ca3b396b2667f57
z8cd5512ec6db80da6937ea748273136b4afde2e80b88fe5e6d38aed2f7f955c3e4c4794a8d542e
z5b6ca9b15e252ba859811259936866bf99e81855e4da985a935ba66e05ae741c1e2505332f8e99
zc4a302b5d93770ac74e96d6dc73d8b1ebd7c329828940245151e1cf28aedc8252c1b73c762e66f
z0accca64388bf4c9d705729754964e1632ccc8ed50266b8de12d20e59126d14ec7751c73fae8ea
z29f2219939363e68496e0e50bb6b1884fba9a93fa451c6c9af8eaae63c4388a16e4f78ceecf1ab
z5b4c8852d781bdb58d708f128fb651cda3fb045b6d2d347aee1b6ee2fca78a5b43a331ac235a34
z1fbfa23f35ecfea2dd4dfdf314d16cb6a812103d5a2d562665c6bbe533232bee69e914a0936f04
z24f4fd08aa00dfa89a71da1676ee495eb18a45416e453c7eb7cdd1ed52db15ee9790a494e57185
za7d517b54a3beb7e80254177e0819046d5d25e3ed57dfccfa4cb1ad2229edaa8bf1dc470648795
z6d4e40a41e1b43bc03fec427c1170b0337085f5348da45525cad8a3767d2aa5fd4ceadd09cb981
z49198d592aac6ef62acafc7da456d0769564f0136a9a6732a045d1f5896b3de854b08da76ad131
zad1db1d72b46933ec2539450c44a7bc3f53cf5a68e115bfb07e1dff4f27ab223e208b5b772ab02
z8a7585a13bd7bad0a1e0185e60ff15a491231af468a3269e867a74ebf73b555b0b1351be12f1c5
z8c29a5d61e4180b5b434d8baa5a4e9348282c210e13f1a515720ab5fee0a7ffd4be167a9bb06db
z36360611a0532abed9c698253224ecdab3b7620c99b57dd60d3f37f51807af6f9183b3d48f639f
zed09111873b042cdf063ebfc908600bbe3d649bcc5cc76f1eb4de8ff5afdf477ef049cc17a4f5d
zb84916a9d806a984689dc68771107bb0b6b9849c82479ab7d286585f5aadef9410e3ee11c03331
z940ce2188ced11c4b7aa4fd682109eaef6e3ab3dd712d47cf247f429759ab27668b1c72b9b1048
zca642f66ec41619a9630bf32a9aeccdc6ed688b735aaf0fa4563466aa21289d8710a11bb3f5260
z7387d27eacfe8b1dbe597a4c245bfa8fdc08a4b7d36d729b08071b6741651b339e6eadfc282d0c
z6788906e1d99c57d798578d7882e8255270c8fa62ae192946cc70ed14b6d98d61708a13539bad1
za23ecde11047ebeef016b90c8713d7e3cccf67b30812661bff1f469bb29fcbab26818b03d9ea39
z9007d9e9ce7cfb7f85cfd52c7f8a93ad68ef3d0baba956da8fbe89e31afa9d22e3d6b7460718eb
z3e0ea77931970d4611366979d16e6ea09f74824f6ea80b32a5bda16698bd3528073853d3f21e27
z1130456a3e1897ba5e2bc709f83f1261fd8e13da39bb18282e60029d828e0d16ebb1e1fc387dab
z622a1a54b3145f83f2054bd6147961cc169f64f4682ff55e1be0e1768d3ad6e09cfb534697a4a0
z076aa842b48c60628beedfbdb41b791262032e26ded6243f255d64798c9bbac5614e515b185b3f
zedb64cf108868f236b1c589e1edf3a470366f4f47123992850ef8508da026c0270ae5b28851ac7
zda59560ebdb7bd719092cc1e11804874869629943ef0efce99ccd8621a8484514cd59d062a94d2
zdff53b342e4c524e114c05d583bb793c0e747f58f709ba7e9f38886f884ba6382dc32344d3bbbb
z054a588dbd4f86f4b3163444aa6ffcd34fc81355083103bbcf9a6e1b2fc739cb3ea2e722c6c732
z7b9aa846d51ec16065195a34fa2f172110a98b7f1c6a104cbd8401fa0d7f3ce48be4adbdc510c9
zf84413fc210aef2257b24af61ca386515caa1754ee45f6d117da894f33d5d6d4e7783610cb7a62
z673b8bb1d4b32bc45a92d43e41b5f3788597b97133cc07e5575a65e87f4b6b772885b3e57843a2
za8b1c612cefe0fd1061665afa0d41a0e057c12a90e611f1f547655b38a4af033048a3502bea065
z54a63cdb94b4a16985bb3c8222a54f58b7210f2a8e482d6bc7d5105b0dcf6847d2bcebd64e2a50
z991d6f9c952255331937f3ff837d48b75481e475f70e6ad9153ab1467df2d0243b759cf24def6c
z1ec1e2971a917550f6f02dfb3bba71f3dea06c23a0b6c38c1ce03840a98a559704a5cf4039efaf
zd9cbdb992437de24326c452da6e3432cfdbdc99d0ddc6600a50eab97417a7073095414b8ea3e68
zbf6d40ba249bd2445888ad64b6a58c28a75b5fd52be5990b7763ea9c85a281872dafa3c95b5233
z9beb1347f699718634a3dfdc7295cf5b9cf400dd271bab18002ef19296c8cb7172bd4e5f7c526e
za29dd31ec25e6c204d7b41c83d566f18536aa07142d71ed5ab1c8adf65423ee2e26f5dd87b414a
zcd889e70f343126ae6769b584ba33dd0227d0ac364ea972cdae5928435c81d0a9019970ea187fa
zb1c001bb0e6f00cfea34d618800cfd096dcee571b4c81c69800089cacecb81711b1fbe192bbab5
z11f943335fbd6d2d30380d9745f025643f3f3d03bdfc4ef3d590da123a1842ecf82aceedc923d1
za3a0920520315030909b5d6a12c195af450569cb5aca1b508f3fc6328d1947579e8759ed6fc797
zfc7c8f144ec3ed769de6f891e8566df77d2789c3323690b5b7649cd26c05da0707b57b73dc7e25
z357bbb356860e4facc0328a9e7293586842babb27d5fe71041f115a14214e1780df3a7e7770e90
z6e2d8873ee3f8f874ac0e1e0862351ef8ca6cb8ff5f8d57cb392f9d7dd31727f7296381dcd39d1
z54de04a9ae7f06d7e72cd6ce2ed1ae46aa6f1946decee6b82fa398742bffa48dad10c5fd655b4a
z49107d7f6e6b30771019ea5dcc0bcc94225b4067d684b656a55a8e80b13a5e56d3564530f4507c
z9be8b3472ca0f99542475ce2d6230016df251baf64e1589bf0b1ad63657436282468a5194dc13a
zdfcf7f31af85a7891634ffb881a1ce42979355546e82843d80a67add973c47ecc6d9f08bd047ef
z8c250c24c6553dd8937f1d369fc455f40ed14e250861a2f970da0ef4f14026733f4235f4cf546d
z46153eb93fca1b17116d3c0612625073ae46fd5d9fdf4a4d7258bdadc128c5f8aecd4034e60c83
zc00fe3e8918892a7d9e85c120440757499d82265f79e9613fbe1ee83f009bfe160a4202639067e
z835914dff54e75668b50109554595c4833309f535eaacdb83574613bde9a620b1913588b8b1de7
zea3c07e91ff21a9b18c5d80a901eda9ae59337ab8f3f64535bae731bee02cb22133949fe0f5663
zcd3629eb669bbf6f5d9d0e3486bfb52402b0853fc7f66f9f363645d3fca34ab26baf96226605f8
z4ddefcc2bdf68239c84321e040721d430addafda1e91292c8c9eb36cda15d43b6dd6adf3ec0f86
zbf9066580e338b1cd171129290d38e2cf32e80cf389c989116b17e197035f5a2c7d814aea70698
z313482adbff8d21866e451c8d2e53e45c17489ad042240b930932d52e70eabcf9089864de88c08
z3f1590f61be5cb0aac0c73717451b10da4820db8e5f282ff806dda36452ce1e0e955746f2fb7d5
z28fbadf9a3ebcb6fb84484cf6fa7f4572f1d22d03373698ea396008ee9d4772aaca0e295366c34
zeca614ffb74cc31c7c19479b9e6e2c2d2dad4c9f37e5d42123669601bd3636ac4812129cee5cfb
zddfc95744680c5e78a73bf5b61c9313ce35656d3ee6fc9c790dad4f9e031f38e6bb9bacd6f047f
z64544d33c28072d478e8ba494f47f706500b5b4fa8ae46758669890d809704bdb5a16c51574721
zc454df08e113c063ad81e9ce98d4569b07d5ea12a5a6ea8729b0358bd7207a3594cbd1e5a10bb3
z3c6fdfa234d947680a5cf42411007002d5d73fcf2eb1ea06a93154e60d9913d45983561a58ff8a
ze450869c98c5c450b483ab0dab52e01ff23c2b77f6b630e2c73e3b423cfbb5b4b7317ad3a2a17d
z22b7a131bf996cdda78faa5010cc78966199318eeb8d60c38814b2a5f6248ab7937b897b811d62
z3c295aec7fdebec4143be7db832dd3b95bb40e9bf88442d99f7613ef446b276192dc3351d91bf0
z4c64a4a1797ec6eb516cb6ff43535ac61df8145110fc91480e398b54a666a9a9a74b6d1152d387
z62aae2571db16e36da08482b061a1cb25563a8b9f8d0fcfe2533e829606137e7bb80819e9d10fa
z4efd51f3efa2f09a4f7d4ca121101a37ff0afcb506de6875387fe19ad9caea591925afab54ec9e
z1fd6ddeff249635e733246b420fb79cfd94d10862e18f19e25bba34e6a79dbf9ffd551cb1b0d63
zb85540492c19641541260a15c5b774e5cba39f5c556d692e0bdcb21d01d06959b68af4b9cbdc05
z330b5a41489fc111940a902e5ed3c3ec5c8355fe400d32ace3ee739eea52996ff4bd19d37c5764
zbed7af6a2ba635136fe3f429b4b8c4e80039737eeb6f53970949a3b364740bc0b976bde17339b4
zce01afb1a206124a2d6e42ab15c46754d9d0723df9bf05a531b41e9fbb8cc6046e52007a43f674
z732909959bb419331bf97c264a36c72ee183cf7970065adb9e619a84f90b854dad92fbbb1d1758
z14b887a4223535ea14e3da3b1e0258e04d4f010120618e634596ed0432d1b523d8426772502282
z2013acce09b16d066159118a7d6aada8f4d0ed342ce36ed6a660e1577ae24a04f63ddfb5dcf35e
zf551a0efa042acca1c0e2fc69ef00ec78de1f2ac1f30881bc6c4771bc86084fb183fd7cce884bb
z99a9b72a212c5052c40f1de8ee9940bda05f854a4378bdce16c687ebb80f201734fc3ab8a7296a
zba821aa3d9cbeb9476cc9c503753bb7090a319b444147eebb2a9dd898d82ce2920a755323e3526
zb6a129a069e07d654b2ce185d6ca7c3c4c786e955c360559fbd92eb02fc136c1df3e24585b24c2
zf94af887b98431df10e08c20a4a5302d4ac26d5a00a0b33bf7a3d882426585f615891985674dc4
zd28a0c33398a97a42e4d2f2798f562bd60dd98137f3c566dd15aa8f19d38cdca9a7c89a79f25f8
z45aa59bb46ca51d41197dfccfb9269f21a74678828a3cf00920b9b405de054648aecd672c69652
ze548e7fc479403fe77a9afec71c31a5e26bcdabcf9613d40a53e52d0a2d7bed6c5399364383698
z66a83ca1b855a04b9713dad4473f12ddf6a832d90e46c0cd77ec8373fde8e8c98b401630323ae1
z430e86aed9e15530d4ba429f04a7cc9e963480414d6a50edd0aa7580a258561f05c7c92f107e15
zeb43846e24ba7d1baf759714e0e79dd06ff747979afefc6c053c319c0e4ac993949fe15952dfd1
z7ac55dbccca8bd0049efdb60cea8dc0f2e453bf8463ba29dac687d774c4308e553e7b61470896e
z87b7faf5834447c3288c3bf1ff7c1d887ea049da961a0c72e1c9766dab2d70d04880f4867e39c6
z9c56994bb6e96deb1831e1b5e7bcc832e07d7b4dc24e19b89131dddf8e6566178c4413caa20991
z141d62c991e153806a39ea66d9453d670c9215e815cf8a6be9424069840d4a149856dc6f016638
z3f3aa053bdcabc9ecf56af60510ac55d9f85bd88c8cf15b40d1fc69ee8639bed76111c8011b0a6
z18ce99b5fddc12dfc54548f491402c1628331a9d77b7b6a2f74ce14e233a5cffb078886e6b811d
z1c16288df3d96d2355cde639478aea7c86461a5777594113c861b74d3381225cfcc9315ab2c352
zb292d91d2a42fa3d9bdcbba98ac01a817f4451f86006f27b8f0829682d71563042dda7e12231b4
zc3e164abd71823fc00b5a0cc9767cb7e38b146fea632f10e765f06c03eb6d149e97d1a5b95376f
zb37201e57dbda32bcf422970fb5c1e662f2c0191740c171c156ab02fc92d904520ed3e7f25f080
z23eb1f71ad86c0ea4ef134e890bb64fe5dc299ddd7b6671e5800a7338a2efa36887cc8726829e3
z75e60cd1450e2ed4a736b8b8cb8c4bb058a053a936cde133801e68685c88c293e5cf82c0481f60
z845250a7c9634e4f9ee8562943a158aee8644ccf298cea35eea59522d99274ab0eec2fab95643d
za7298fec06dc0a1a438439bcfe3f51ca529d3f5a665386983fdf676d74ccfb9223e3d4e894c018
zbd7268362bcdb613b1ce19858f2e33bcb77414a6986d7d96234a0072513a9eb0bfad25e8676ad0
z1108591958974a3a27a772c3c5d5213aa060b6e5f96fbd6676a1d277cd64da46b929d8b7b7e219
zdce4c3525ad06a716a129ea01cf2c6bcedbbe760d46c05843d787ce988a4d8767161fa36c7b742
z747c53777c7a5126d1471e09eaf7d76e4afda7ea50cef78132661afde052c3549e7d669674d5fe
zdcb2b931402c60fdbc87b49b2db31b58d2e50f78cd7db16349c15737b7f970d89a4664b0b7cbc6
z97f1b2a2f7c67f694aa41854914edc5e9db4c08870ef507b26ba211fbce51db7297ec3687b701e
zadc0b18022de90a364a62da3991bc96b82f3c171b5c7bec6a6fe79b813b2c010f8c191e3555f1b
z58af14388e9070970b88560c755b9e4275e86069aa4af360ac18a310f6ca63f38340ecc5c64350
z9442869479af8f09cafb1cd3d3fa6566f8c6bcdfa23c5b407f472ec2a1ee05daa23a2ebc8f85ba
z30f334c563420fb48a4be2fdab6d159af4fab2f12aa6e7188208f3dd51b2f86c6ede025b063efb
z01380d1a2857a7f23a57718f108862f35ef8fda786e3e84fa46d4cd270c2e6e349081bc503b6b1
z0a571bf9ff0007cf9a606cbd0ff8281ad0be2c3e1bbc6c383239ce995b8e606136f89682a0d333
z89843a7ad91e14a2d9c535b1c53d29cf2e6872223ff0f8d8b9674cddf4495cf2bb5a209dada70c
z4b454f4a71313f81953d6345be0ddf1c08fdb40aa3934f15bbc9a9b73022c8e126480994557512
z5d035933827cd5b13341684c2e5e8b9e8f4586e8df0f6a3a41e925a83a1068874a2618ae6ac47f
z8e87d7a130878cd663d73902edb17daa2e8535d169144b33b55f1f182dc750151da28910953b2f
z807800547e7e819773ffce02d74af6dc2b40aa1cff80c913b0b21fe6034da2db201ef472129830
z42a53ae6b313ee9ce2111f2fb1c33d033679da113b366b6817d69acd28b85a44e57db17ec493a3
z7f7883baa4116652d29d145879ebf824c0a06de88e4b161a01ae8c8d2746f03013dacdd8bf7528
z2313f4b7d829f67e19685bc05d39535fa2b57025ed876743de14b10860cb6ec755d8f0fd510d1c
zc97dd5b73fbc91f67a6111167da963e43b94111ae6b600b13851a001d7a3b05ff7e61f7b67f9b4
zbfbd79f4dbe579de750422873df024d69541f0ca75e81f5bc3569e1896cb47fe852501e3ea0a2b
z69ec50303cf738bdb1eac4b739f4b2e456dcb6cec68015bc0fa5bf1a61953da41222e846dfb446
z4fe18359401bbdd8dcf3d356fd9e202b797dd6a030ef3e7837427a253d7d78befa7665a5964872
zd271d09e6cabecd291bac5bb464d07fbefaf8b512b2c5adf14229b316a786ea2a160b8c05f4c06
z24c0e1e6fb30e452a9692ce254f79ff8459dd03e48bc100358fdbebc58eb61771fd676fad9a3cd
z4a4f3ea2fbe9d41e777bda43c3e6eb51709e5cac79e707372733f218c0d9c1686c485b831fd933
z6c41f90a1d2e81cf7f49c1452582cc8a0b24dc3a12adf1f2ca662324cd87ebd0d69108058ff8b2
z55c297b817fdfb00112918985219cda5c2052ab26f98132508679e3ae0c1963b6a683aaa58ac06
z7ab1bfe762f0841799b547337d69172b48ba0e5f1fdffd5493c79d8dd7e7a03805bb2ce3141b80
z3523fa04df7af6ad2fa73e1250ede1adf9dd01a2a2fab31af36d13d404467ea05f1cdfdae003dd
z358b55093a31182114f02bb707a5f275c2301ceade41ef8f893bc7961a4cbcc89201c545a43283
z694cad3611560b9eeab8b41f3bf860c0c4cd5466857f620bb172e95664be2451ea901cf55dc9f9
z8a6480b9152a048fd808330e01ca2961dab085154d9d125ceac82cd3d813ac292d27b4dd09e796
z70a42b472f39aa025a1151739e9060e162c005bff800103792c1dc566c256530655a781dc9fcb8
zf9ed0c9d201491614eda61e1c14f7fb4494d8ff0f88db3035a060c17c62e225553f6f9f53e3702
z6272a6060c23cccbecbedf6c9b0359504f754f5f39fb45d64857124b38553b9c05b1692a599340
zd25bbd0a101614dd458f570ead3fba4bad28b3f6d7c56070e37ef59440ec7818e98b5bc5b0b341
z3353f0d9ae57b2accf4727970bdb4d6c15f47f2b9b25e18cf32af8cb286bad50bdc5b1204ff001
zbb9084e04078f627fb786d0568aba17ae0299d55163c332971dca92bba87170c43800432ec86fd
z30380105a3fbd5219082d4844cb3e72dcc02b99b6c6cda9e65e29acc0fcf73491746be62501967
z1a910e969d530b207f24ef867578bd9535dd9994e0a702b7f6a254993f606278dee68580e4a660
z22f5467ac1c67c087e6528bc29e3b123a19a3ac3a198de9f167bc7ad18d168ef8e11888286d750
zae13038711445dfa17485197283b682aef0448f537dbe7497935a3f21bac8ffd639dab6c2ff6e1
za0c3263259ec625a1787ce60d45a95a9069a14675ecaba6327ede152539dae8d0d01d03c2b4477
z95cbbca511b5138e61f0bc7523f1c6a31243093fb11db98b4716efd51426b5e4a59ac85e2b0910
z5fa0bb36b71681733f9110426bac9403ad3c479b902143fe451e74e77815a46c55d36fad402293
zf17ea6b3d3397d83657c38c7c7a1850ab2ee3573bb1cef27ed55767c1256518db6da14e0a73395
z0be1f4daae484a106584cc3e94207aa1ae1687f3c199ac14a0f74274bbce9018fe77c7af4a53a6
za92085717f1fc892c3907a72f51b4850908c216617fb394675401ca67804f3bf5a31ed7c72a0b7
z239a5620cf70b365d0390eef710ba82ec101a79af102d5f647071a5fe7964f898061f8a1cbf686
z42146548bee705feb5795fef6cb6d1682d007c78e45b9187578b7c82e046265088ed1595568a05
z9ddefb9db1f569494ed60fecb145e4429274663127826f809bbdd8371148cbe0f0e53f2305bc10
z2c39e3f2ca9433d64431165bd3d9488ddadf6c665d010f6e24e0b36a29422f45d90d88bc865520
z2c76f94600af1bbafe6dcd445a08ece14c8a92274b7d277cb59df09c883866efb4bc5e968ddba4
z49ad8d4ed01abbbcdd1a82cc3b645ee18dacc6e32f9de27cb7dd2cb6716ba4319bbb5165602708
zeb7f7d21d33909a0eaa68c68df4e8de13e4b02b3def895f1a847859ed3c8ed711c9d85d2d840c2
z36d07c9cc3dd1430de04006f375da0e099bdcbb5aa5118a7e39897a11e0e407dc64d566f65a809
z0c2a481584878ecce04b769ced7605c753a406c10aa93476336dd3841548d6a0370073218f1856
z31f2f62d4c7efe56656dda71c3a3b233e2f54f1985a93523a312fca85f23496300bc7d975a91d7
z35f7a59d9047a844ace613ff49276c3ada8747b5e40c9bc5c166d265bdc0b7895e068903c46143
z3995bd110ea134a19c29f442583b441299cbf01e35d8a0568c945d7c2af7eb06468b2e921951d3
z3e8841ed5f61ddae960af2205c45f96f482a50de7e0d9adeced97d6819e649e255f20ba8cfe7a8
zb5506beb445f1b034fe2405be9420f719b5e65197f6693f57cf99c37166d9d0850f53f34f299ed
ze79d4c01987463540dc2f85f13035ee38f3d365f9b58663ac1c5071cf5a76731177f19ba22db67
zb18473793752fc0379b5ceb441561b3ad35de5aa1e399fbaa3d3348a3741d19c41b6dcbb359cfd
z3ef03799e3c9d09409cecd96532957d161c9be2833f039dfbc559e67bfb2876e68487484662cee
z2d0fbe9b266ac904eca3c248d915b005b96013fb1a4497935922200adfe1dc12159ad32329acd7
z774c0c07428b153d6bf17086a8427d54e1a99982b0c98b796888e816760f9f42940460b9572507
z232e11b71844f64b8c90562893ff309ad297522cea891ba3897fa6d5a196f15498432866b8355c
z645f34dcc3ebf3fed5c283753702a4c5e2c446ae6184b49ba0e78c81ae592896d4451d630a2235
z55482a3ef51a8baa46bd51684f0ed22b4558f8a87f3fde61241314c63ff712f6e4d33d7b3308a5
z0e41057c03269ec84aba9a83c0b883239f86385d374cb82e68976a419e75f8b7fad0cf76911cd6
zfcc6b9df9c27e903351655a189cb2b14b621d92bc5bb32dfa19d80fe56b837d3416180255f36a4
z44188db72409aa9acfa17a95530083105a186492afa87fe3650da242aebda5b53636e34c3cfcf4
z6b51e5a256dfd38825056753700b66d1c79c0ded410236ce76956d9c3d01705ae3c997a0bb9ce7
z2303a4a5f5c6064846caf011d9e23ea885b5bac154e32ea33b9f57dcd34dba59ca63b8446cb877
z0a9d282bc8877ddf6d0263f0a1a26129c8dddc06005fc1ea8b7dac00ce04a0ab1891d2ba9c6396
z8d4ad7a443773df3950936d155847ef50632712638e3a6dc23d8a6245b59d1e32e737f294e4d5d
zcf99f2b21fe019c5341b4ec276e2cd63d1fe78888d279b730232d1b3b51dd7bfb61a385a78507f
ze9ba78d6e998b620428c3e8684e32ee210480cbbcfddeaffc8395a710a30c09acf42550a70ec8c
z665915f9d46a0db3fc8694990e58d9b958212e6b47ba15b95331d675590b1cfbaae5f4b24d9936
zd4726039da1f7c98e6a8b58758bf00cf37005031d8fe34833f273b37f2ff2f6723d05cb8612e92
zc773255d06294ca31b3ec0b94dbcd19a4e6afae700a9428a00d0cf8a4b6bc7bb106a5053bdbfbf
zfb20b96c719a3ade557c1fadcbb42e6ddd95ce6139e91c859c4b469c788022e14cb11e98bafe1d
z182f37a3a5f9302facc3036d8adac14935a7e560ca18ebe6b7500646e7b5f455b1d3c306fb7de0
z59e6f752d2b1c8950bff3425117d4f996032803631a43619f6ab61f5cee9fa28757e8e414710e8
zbc71947f6455690fb7dfd10090672dc778cbb51fd19074e69038c818904d5317832b1f6def0c1f
z66c4afb51b3584f95c8a8bae8fd2c933a9c8afc71d14347e904701cee383a8982b5d9cb4fb4f02
zd69eb8e6445f0c866486ed596070c1c070ea33cfda7d7b012550b8676e72f6950fe9adc05b0279
zb6a2ef79a9a16fbcf082e8516d0bdc1dd8ccdfc74e67d7588ccec6b65118a35a45231a14a15c7d
zd7f230b3579e510589b927a75a33f3b840c24339063e8969b8012cfe47e131a419ab5690fad588
zc330edca046c116b8b6ed4a8ffee18b2b5ca66b32ec185aa36d0d30e9c36e1403efabfd6001ab3
z3698ad647c92fc3152d62ab17d7595af8cbd397d5fcc9d933f0316e03f4fbabcdf709958f2bce8
z4cbe5e4de204f2f26d3316c595fc77e1dbddb0f9dd55756535f913ed1e009f3361bbb69a9ec0c2
z64b62a502ffc8263385a7a8f26a2a2a323c76599af3ba2ac7bc30d706d8702c9da8902bedc55a5
z325236fa35b947d479c1d6767e926faddd485c7ac293e925de6a9394082ffe40a8d9280c520d0f
z54713b52fab02ee1b5503bfc11a2dd112332b04da06e7c3a97d83f654355223cce4edbebf95035
z6f568aa1b243a3d2c84aa1ab7d5b2d3ff8bd8d9fa3e6e7a367a87b1a6297e7cde764e99ae9310e
z7483186c2db279441429881e7db381309eb3f63cb61e4485cf78424d80e1bb94881a2570126f6e
z46a9b2a9d8242dc0b44db1303d169bd2012bf9bd64c36fa0a2a8ee6d789399394b2b979cd369c0
z9f42f44a40e4bbd0efeedc0165e964fa8b5c7b0c298a2cb3716412509a8d0e26057b7b48efe00a
zf111b3bfed2196a3cf9133d9ce7edf48fde1c69d539869c0083e0a0111f5e32ae9358344b3a050
z6811e1af52e022cf53e85a67317db3e54311b6623f616a64547d56bd6a076afe9e0efd28e26030
za304f44818e4e4c6fbcd6335de76dae7190f9d5c10d37a23e079f47fa3ffa2686b4a041b5344ca
zd0bbc465994eea4f811b5bfeff3b7d2d3f64ce0b376b194bb9152decaf1a6d68637680e525ee1c
zd9bb93cf45749513272fdcfc37f193e16c803a309dfc0f07bb07fcd56b16504c8a3b1f828c105d
z8e45c7fd13eea2eda2d175c8973b161063a69e8362e12cc0f682978952d10a9d5817d5fd8e4b7c
zd6cfb94f09b10b30d5700acabe5cf2216f55ba2797810be2bade1f4c4c5991ce3a6dafd7ddd596
ze87a3d1ce05157a2366404d63d716ae6ed8fbe101d4a6e48b59494bb6f0c317f15fe5d08525c38
zde6a1e817e9f39a76c24c0bedc2c4451db9f2ee055ca2a043800a9b4673e9afe6da86fbbb223d0
z7d7f5475e180c1cdedf52bb07d268d121a7e915649c6d8a7e6bbb619880a4ffab84206425c6b54
z2fdd27dafeb4091d65488b51a222cc0b7d6befd25b3c2cdc448e76efeba318e680806898c5a780
z0eb692a3c6164731b28da902b15cdaceeb17051d32fe42dd9d0b4ceccaa095ccf9385c44fa69c9
z60b66bba5fd48c8868986b8f411149c00195d61e8b2b7544fd0e7848fa81453d98ba7a9db7f406
z720d1129f0f10a869bb25fd7f2087348d9cd2dc3c20033a787b7c056ee11be315a0add826d0855
z8e54fab8abec3c820ff1bd9b3add787bccc0ee7ff14985854572e13c26ae4874ffc06005c8e1a7
z39a14d78df83786a9015c55ae539914ea122123805cac7f08cd8d3def97164ccc07053765cda39
zd794eb0eb8d03b827b8a4f1b2cf504d3d69bbe4df19f072e2e81c7f953339840cbce180fb578d6
zf3df24adde616dc7972eb7a455a665add813a93ee9e22da4cccf659ecdd7d82645fe03ed8ec55b
z28e09a43801ce9fcc150eb85ec9dcd92d8ad9df2bb62e278c71e5bf60c1925f6711d694536d49b
zd47c4ff42b5c79db2d9de04087c4f260d21e153902ea5ccc8ea49b9a068d6a3e8ce7adf1759446
z3da92a8bed51d26724e409d626012eabcd955078b9ad551ebb64edcc73c575ac2962ec2e834779
z3d68824189dc7937ef0dffe5a3fa6bb3b782b0cd3cac54374098ea25047553c657af68cd616f42
z6b4455b85a4dd0115a5c31075774ed5ba0fa2b68d51259193ffec5e0e0c0e79b45f11f5f514876
zf500e171fe7e62ef985504932490e445ce42741c3e87e07cce397d3e119bd5990fb7acb1796230
zabc4aaf37fbb3e3389b096c42f865a92ca6070c63de5452ff96728feaaae9fefcd8db09fdf6fd3
zaeabe29b15c602710351b71c48a82b328069fa6281f40ecd4ba24ad851e92ead5c839f12a01ebb
z279abc245233ce16a95ef1802aa5943baf3327a3780ed8642404e9d16d7237c3cf6a7098c5b609
z43deda8e355a9a9959e345216e8be75fc7af8b50a09c1794aff210d4538d2627adfe70bced16f3
z0cb7db17ec59600d5de954cf090203d8763cfb1e48ebd5252552ad45331aa85e7f1361c6dfeccd
zd4bbe9363252700121302841fbf69ba7f498145dce44323d16e23ec08e87a38bdae76929522463
z051f1e4583bf6b3a5d90c1fbbbcd1d266c2d94252e623c7e2c9b791bf87010ec8b8adcd12357e2
z2f17a58664da824923c7f135d61a78f9db70a3cd0cc69029eaa3b6fc996a6176919fc837747b02
z5db4361177f2ed3b098993f8574273aee8a3bbbce188cdd640c28434c1c5802430bbec25ec41d8
z280840553519ad2407f1a8b866afd65d015b29abba8b3d6c5f1c3bb56f9c2fc9e96ca06eb21083
zf89fd76a0ae3ecadd70e42893a02770fb8706654fe35f992174eb3b7aa4be6fa64242bd15878a1
z67eab156fc3a92daed89ba8cb5418b96399282c1fbd4352f61cad7eb5951952b3fed33365bb3ba
za97c9c80aaa8db1991abb52ff77894c36bdfa142e182a2c4ef90fc4a090d40f266da534181549e
z294af65b601583ff607fe29c99b83e3ecc7d11e2bdba3ca5e09e8033542dcb08fb8713edeaf70a
zaa8c3eef9d12592eb5ad783bb078c41856ea9188e8984b58902d09e95b1eb5348ebcd9eb2bf3b3
z48e59e400ffee7a5c1f58a318233a43f7110e23f6624298d866420b0791a2cefbe1fe26d836f1e
z72b9d929fbf580065ad9821382871ddfe08008c7ab26ef5801c6a9575706e0361520bdb8625764
z906122ea4cbccb701e60d9c24adbec2b7b2547ea27ac595ec8bd0ddebc2873c71050f2f7e006e2
z3752d95fb8abaa2672996fb8dd0f37200048ddb639d60253a911fdca1c56c053f9844b0b8e2fa4
zf1fb59a1fc976973de7cfd74ae31d3572d445c90648697b9fc5d955bf0d9954db9e1bf5c609013
zd6393d85bb8e679c07631bb6da722889b8d9b8d003d831913ececa2f944f2d1e95d467d35c809c
z7435b962289dc22730b61a64d540bd1bc0a64406882f4ae1d012627714c80c9f7fa576b21cac65
z7a4fe8d84a2c3c681e442220fbcd4ce3ab89d5d8edf7494ddfcfd04aee3ed6a74fcae88e2281c9
zf2dff23a2f537465de2855c26b1dd1769c78e058502562b9b8b9aaaca25e4d5a22471718492d8f
z7ab3cc9a1f99fab8d5222ac31f5500b14c08b587ff96967bd8eacd3f0bf813a94f96e391f0ec50
z2593165b4ef70bd099cda573413110c8609906303d18360fb708f83852a246de1f617cce308f2b
z32285afcd7a140af2b152c395a9b63974a0fb672d19dc6885078f6f3cf15585641b77f984d67d4
zb1b8b32e53d0ba8c3537b742eb28769eeafe6b08f6b92a3b06e8df1face10d48967e44c7e7c499
z9f1a9efaab4a1e86d177a1a04c6f7fad72af4713a670b8c1b43246a9780b7f8300bed170120012
z65ff8e7620b714c7e56b63250b162222befbb461a76703b5b7404d19a30265a35059ebedafc06c
z20579f65a7561ba33c4f9b4af439423fae453dc50f0b08d54023e7428ba18d87c230a7a9c44f01
zb218a62b65537c02b165c360003b3da3424043dd21e277564215c710bb112e1da28c4f17a0e949
z9e138195f9f0236c38d27a4cfbbaa1c4064d1f654f34745f455a06375d0c12bcdf0bfc406866c7
zcc1fc195dc11bebef03e21da3d703eb2c734aafcad6eb19a6c994915d7e66a92567d2672856ba0
z912dec2315aae8fef51caa27e3112e63c5f8a63e48594f4a01611d9552b4575a81c3dfe4fa6604
zf5496e8397bf00f75f007a5c6ec06797c5912ad8fad5c0c7ecb017436e8c20dc81c1063db34b4e
z6f9aea96f35b066385c37ec3aac754eb43f677a72ea7bf01e5f8aa17e688bdee82311b6a5f64ea
zbecdf8dae61cea6fc6363c5009750c9d9940f9fd5cd170599f51abf420981cd5e7fc3c6686f5aa
z7d4deb61b240cf5af0875e6255f27727ceb4e06437fa745ff972d459aa4026a41b39092067aefc
za7321ecf1a83345ec7c603f3134d4b30cbcd2b95b2d340891f089126bf27a6f2d467a80ebe0e6c
z3724f932b01584cc6804dac62ac484f5fd5f989b4b2daf1405334d84fd5ea025aec6f380927a39
z257c2733c3a85279289dab4945479b7a33512df3f1d91c4b21299f066b8328688c41ead557bf06
zcb81a369528168438626b46f246e0be9cbcd13311e3b4c2787b45b0a23f0149f304efa01cdfdc0
zc1484f047af387b31f16b7828dcd515c8147d4a3924c2309d9c0d2e2f849ea5d7c38122f2f533d
z6b1ae3643000acd0878dfd544cfded070b0a2dca7cf85e894c7331eb95beded0281f56ca00ea75
ze098c24bb777f8b9d778a31ee30910d6b2b349a06f8083cef1d6556b1ece32d38989dd722de723
z63ff321afdea297be58614623a7a60e7462fa2b38823ef8bc2a7bb2f5cd609cdc1436a5d5546d4
zbe9c1d717d62ec450050f8442be401093b2995c0222b60e01c65bf3c414f1079b33b9757741d7e
za4d7e487a4502af10ed29ec07df06d9e8382b6b14f89824f501f211471f0892dcb00092e475ad0
z84767bc3d7be2c7b7ee4b0bf29c33964852656c5f153e6e6b623ba0fa6cb38c12ab6cc8d25d6e1
z3286bf024cf5ae13f234fc0b91295b81bcdd5feb90878f84948de40e8eb9b80cbed3cadeb17110
za176800d93cfebbf539d6b7b206b5e42d9857ee17aeaa23691c8835e300057101baf7218f81bc5
z63caf8767e6b635cd989bf6b34bef7d37deb2c127eb9f4a56db9d0dd8cdad9a55df9591c01e4dc
z1e5658ada787b299f349a5edf08f8edcfeed0c2786604d7e08267f9b9c3bd1a23cdb67043c6ba9
z1b16e20a760991681d37826258a42b9806a9bb6b6c25de320ed15a92464c642e9f4eb2f6dc05f1
z959d049ac5eb9103b90419675571ba1db6f98aa2b83dda5b9572807761a96f5d4153fe706be7e1
z994d4b4b113b1d7b2c849303ceebf0c67656225b387b8f6118f6b93674ef601b0286bdbf005955
z765e31832704131292e798f6e82683a668976a24bb9b5949b6b485e92ae38559c45dbd24c735f9
z9461fbe4e4a362acc646b1468795ce5d0e4a4e1d6550f8cd95f63dc8b205f61cfc37a7d29bc2e9
z408e564b07944ea6688772c3bbac167301c4ce9fb4f6879c9536226abc0fc65fcf9d4d84eefac6
z071be40e0b8baaabb1058202ef52a4c42c038e93ebdfe63f97fe31266b9cae2bb287e0fcaeb3a6
z94969c7e0a906b64ab96ed9d28f97a8baf033ef54dd5e179067993585cf4391c253c34dc01bd8d
zf421efa486b7f60191e90832a8e09649382705fae5685d0eb39c680128e9634209a03631eb1044
z7efcc4c9ed2699cf287aba2a7fa4d7ec594813ed58b9d0d4cd4333e29caa42bbaa8749ab9b8025
z491f44fb7b21442e025843627f0c118333f697f9b39abb55323d400f1445d2529d48e88462c5cf
z7ad43174843a71882f0ee2e39756d9351c368b39659724acddbf92b912dd58b27573910318bcca
zc10b3e1b5c3713b83d2bcbd3beb878c4c7b7a53ed144c0081f03784316195af4c16681fdf291f5
z7f98164626290ed70f60501425017e8d4cb0bc0a71ad4625face0ea4b32119781922beea9e2dd9
zf8ac5367a3fa0c6f81f4501f2e0b0f96e92250cf9697c7b9fa3d8e9c6f6f8fcc48056ec2fef862
zdac8f78275464836ab3d02acb3e1d42c8f24eb8a8e338ada108d34fe6ecc088faca8eabab9449a
zefce7f986949144819184098fe674d39d536dd243e1b2f2378f1321b0c6255f5e14f31ea3d07c1
zd0992e5c8159f787fe8428cd6159e5e4f726b48b29448e3d5b356cb20ae6d91f98c51d840e3b7e
z7f10dccabf35dfd3b239e1973d194e7b806af2bbd4dc5f4ae949847513db86283ab560eb22ad04
z39f1742c32f8ae5b50073e315aa2d23751dfbcbd80442de46f530e9e43c02a88882cb7044c65d5
zfe641911921d0a6bad520f0cb299651356c6b5813cdf37d8657861783cfc73bed18b98c64e7961
zdbec4f0ea4b9bcdd013564268b5c44ffb992300216b8b63a805eae447818effad57b9c361bca97
z8983a4ad14ef9567979f60de14e96278d5b1e82a034b2ffa9eb1d0ab6bb6f391bacaea3a774670
zc2011cbd8aae8f571d25f00a2b5a4255d3106e1bc0191885b6a9d7bd970dbf965695123e8b27b1
z20eb9e13d5d5f1a6efcee920d1206919abb8bd92fb85d734a0cb3073ba33b1d3e6e0b44474c842
za4e4a0a12cd795a73896cb3f9364cb74ea7323cffe56e1f4191738f49ba13f913b616c67335db9
`end_protected_0in
`else
`ifdef MODEL_TECH
`include "qvl_sata_sapis_monitor.mti.svp"
`endif // MODEL_TECH
`endif // encrypted_0in
