`ifdef encrypted_0in
`protected_0in
ze74c34e226135848fe16db9ffd31815111b6d7fb642c521a3f628cf6da949865580b22efd062a7
ze90adae0e65e66a2c36a587d0a790699161455169ed55a01f2084f11770a774ec4c588039b380f
z6de9c5084882a40b79a175f5c2114b2b6d78b070cb806e1c0aa9258297f4687ab308bc470f0040
zb0b1de382961eeeaf2e279e1462520fc31c119af8f2b214846f56c2b3cd2eadbe4099496abff18
z15cec83ec4a77b868344aa20ba7360908f5c0de2a79abf8b3534b883bb12180f68b5d4beb444cf
z3fba8f13afb0abfe8fcc4294810f75afe452434d2d0f1166236c82f76edf1e12979f04bc35693e
z32ae028996dd85737a8f5adc1ebb94f39c940246e887647b64782cd7ab429b0544c173176cede7
z01dfb26b1f73408344a52b7e1f117f12bb9c8077b34876c2e6fdc085981637012dc9754765e1a9
zc512ce062e0b8fb16a214591f5c81e1353b900a611fe1f4886b57940b41b7f2ce99a7b84b04b90
z916f717e73bd10589c81e207ed77ec660a8cbed5b487fa50acde1b055c8870bd8676023f21ddcf
z9c98cc47cfa2d654ff1365d1f45035a045a66c5dfa8279050262529d2cac9e64fd27d9c7de62a7
z731bc808811ded9016570962244887f98fe5440167bd0088f2f049df882af501358497c3b28776
zcdc5426c7f52a851c35106bb93e16fff984784050fc808fad15da330f6f0607eda2d0e0e4b1215
z2ac5b11453f6b6c5c6b428261a64553d70b4ab9f1bc235c2ceff4f6e3b1ebe72fceb7af9adc96a
z694b4bad7241bfbe775016041d7caaa74d9c0e7b507ce89e8b01980415bfa35a8e346f54c548f9
zda8767c02ea87d27eb7a843f4cada7dc3b575fb5cede69da7a4701b2d725c73f1f7375e85a74e2
zdeae70c30f1127407402c955b283d7b9512dbb3cc85aff97f613d57a4efe57b3c092e5ccc5b6dc
zd01018bef01fcb6b6afd138be37349905063433d6fc88423f78d0a5cd8c325dc906237be6d3673
zb87d9fada90e2c892651aecfcd04caae277f299df76d77ce870132e5e40888bd3b3b1b6bc6e799
z48a23782b89d176bd848937c64ea2b6938c5a6c2c52409c3721f00cb676ae49dbce756d647186a
z2d5ecb2321a08bb462a97b513b2f2f7e1913c836666420a662f742f4dd090636a3381f28becec1
z1708d87f1f0a00e76b7fab8e82c4b58a7479b0d3618edbc64d306b42be8b9498e21a252a9f7760
z4ddccf620c22105b64d3442eeae29848475b6321275c60da85fcc15cdfce58c0be67611b4ad217
z85faa32f1a391d7896ecd2d6a476653f33c744e342ca0bee6222cd817d247928bb48ab87008585
zf4c934887ffb02320d1f5e9901371c546d07491c6dc0560188ddf7660969a0521bcf06899960a2
z846b97706440dae0671d4d93134b115147c7d3bfbfec814d2c532f2bc7b5a866f7796e878f79fb
z6352953b57e9db9e47653b1e11547331dc0137729d159986fd727762f733f71a51abb4c40cde6b
z54c31b12df4f712a2c305b789f9c8c8d46984771a07097977cf132585a196985bb181add954404
z36bded7d75961463e3e276ac41eb95a919dd3f15d3ba1ce8c7f86d6b40597e5bb339c0a67daad6
zac5ee1863101a987222facc3bb678e491d899fb1eb431501044c2b2d35f783cb891ec5d5020e46
zd2ca6788f75aa91e62a9b1093a2efca24d5307dd08c6dddd7acfee5bfd4c2906f8ba35164346fc
z8d38f18585863e2f7b8d3aa32d2dfc1f4da86186443266a04614219ad5d9f8f6aac9e91c2cf60b
z7f8a858860e3bf81cbc9bb2155a49c53b4851dcecfd2c4b56efe1de06f660a83710e76f23f2f22
zd0bd217b24afe7b8ee8b016d1f156d4c1ca8c1c34a1fe24ebc22b7a10de60d6422c374930466d6
z56cbd54e5bf0cd0c652b9bcc268907004db8f51e0aaa235277b855f3133cfb60d1ae231f6ade4d
z0cd48de7e7ae52607b3ab6508bebfe2b5ee6d160dd1274b57d3b6201ac37d4a9bed038e4e6554d
z41138219af55863100d4bf833f81ad60e3e347f831260cb61f9950137088ebd58c0d3165264466
z222ef99b1bcf17065a01ac91ce5639387aef86de8c2dc191403d40545a03e85fca7fc901a118be
zf7f21e350c94f216e6168f5f1c6c743d0b4daf5dc683223a858975b483194eebe86ba672a710c6
z7b991ad9b48fad727a9de836c16ae386cb05ed753e8f6c33267d0ad13c8839b5dbe7e88913214a
z2e7912365545074d3e9daeed16d9a47c4e5d443f14048a4b26d8e252a1529ccea85cd180064057
z9c4bf7be906fe40beea0a0318100306591ac7f728581041db4d68fe11a016ac57da5655b824152
zce8dec0c29b429583eabdec51681b331da7b974f2630e93d4529ba975088338bfdb673e0a85fc4
zbe782adb7350a5fa17a683e3a5b867c33b9dbe10174fe867d2b94ead229863e34194db2f38db42
zdb4355aabc4eafc9b21eaba1a1c6bfd3c4f009552fb8523ece3496c0fb282859fa97b2900e7941
z405e00690e80fa337a36e0f3c6077d15ecbf911cfc2a7469c54abb1a27444e5ec315d4b69e8bf9
z5c64dc5d4b83ff426bba4080ba0ac8b2d668fe780661eb2e367e0d7d9f77419d46e8e5451faa59
z58dae9552641aaaafa9b6a0eb4227a7a8cbc1cbbc9db50de3cd6b3c76d49bf1293c96bb721eeb2
zbdc45eb75cf6c230f827acb5008a3a72290748e631898bbf59e022b631a577b86e5536f5c77da0
z18d78ce429573e0712552f23510ee8a5b699df73a2fd4db5f5f0e751b7803f1f5f4c1e6c437077
z16fa213fe64bca4d150bc0e27e5f55522cfbd687d6574df021ec0426a6ea1123932e99e718cdef
ze24337ae43e97f21c143fcdb8c462faaed2cae45746384e6b7ccc02621b18de5df2229e1b600f9
zd8aee9acc550567b0d00b087d187030b867ff8a3e89b3542f97965fe409704c2ec380b4c995909
zf41d3d628950c153941d8bf6d819540db0c02a343961f019f88aa1a3e56e530682eeab03c5d75e
zd23543a4ff45384c20e8d9af496f99b2c38b6af0158a069cda4e4cab1bf50d16e384baff2699f9
za853dd8dd504ef4cdefc6fcf791548436ca98882f17193d88c48f3adee594c6d63ce64584139c2
z7f41fd7588c26464bf2607e04e584e65185386c078dc0a262c53b6f93dfaef08825b2cd1675727
z1bd856c770ec393e8f6cc14ea04624d1385cecd4e7095b612624e085b989ce7e1c2d1078956da8
z6155144b94ff67ede507346e344223fbd039644007bed23433e5cac673e2e843bf525abfde7fa1
zb390f63afe105da4353ca6b34158c8b366b6e31a4a4acf1bbb3a59c4ef1271f234b9b018171e8e
z1d90f1e88de273efe94935e1eeba5b37c88c3e1c886a5c3aac0ebe4407c91735c6c24388867cf6
z976aab99d517f8a3e4794b02985618fce144c908dc47dfc1ad51da613645bcac9911b3a4b37f0f
z2d3facfa7501b312757e24a5f8bc2fde953bd7b1a0306d860446b0767087b7ad02d02d3d0836be
z98165af17138ad566a1841429f4bc5c77b364ebeeba85e5054b3b98af59d048998c844a23547e8
z7be70221f3c88365266753a728cb6f861b59a1fea3ce1212bf8af16a60514d4670833543180c47
z1ed04569681d565dd9c248175d000041763cdfde8b700bb439a3d005cb37953e79c7a589703f7c
z1e2d20f1c7349d99b1fc822ce7f9497c5808dfe62f38765ea375386119f21fb958dedea6d27c83
z2ac73f99df9b2699895abad6a66a368857856c1bb7b569231a06cb6c1c44fa67847e7f3a5cab31
zc48e7fa5925d2a238ae121b8d45ed9bebbf898c342c11ad091f617cc4bc1ab5e679dd8057d91ff
z2966b664d077f262c63f5e20f04f470995e2dcf8fffe9073af6b4d7860d0b862093f7c66be168a
z8c6b4fc1ed454fab7eef2b165f4262fbe9dc6b5437e546b4aedb1759d00cc77c5248df7ecb7182
zbfd550139d0d8cf9b97d30cb2d25f10735bb67a2d091cc5ae65d32e63903488b118619ac65e577
za5c47fe51b7c2ce069f45eba2feac3a2ed3d07dc7c1f0a03f230afdad57519164a78f9d3724143
z2b5ed5f2c97d8bd6c5c59792e9b58452457e5f28d70e968324b7a00486e7c2c8bb12c48119166f
z9c3555a106efc7218fd081f96bbabb443e97500b4b0f4e5f27da4a79def5d813b75ebaaf35d668
z45d9e4fcc0433dab32c78ab5dd7a8bd8b78d8f4bc24f7d81de1140be9641bdc402d8ec0ec6f127
z0df8d6e0ea892d3deaf3d5c78f932a6950425759457be43aafaed496cb7349f33fee40ba2d3cba
zdba668377dc8b4e13d8ea9244e44ad745ae2955b10b34f290b498ae2d9a6ee0fcdd4dc7727b8f8
z960805065a0cf1afb5ab71709c945913985c39324ac83cd22fa2ad43e7a463dc4fdf54a0fbc628
z9f509d8e7f7450d8d77edb2f24b2e7fabbd65305a40d7923dcc82e3f9ce692dac2ca24c3a71d4e
z9ae6309399fa6cf8b19891dfde5c8eb45b4400d22678abb10ffa07756865adbfe0bf049a346474
zeb095e54cbc9f99038fca1ec3407db77e3ad03beb78c447e25060d7fc8f19f6ba1c08cb035982e
z6bee464d92a0ac63504db5995294200f46137c85bf676a38f4f5715f6afe2859121a5bb568ca89
zcae4ba9e04437c71deb15565571578f5b7d6470ad80dc1af447bd1a562d1a89a9289cc764a7267
zae3aec0ae3dd66c6d623c3e6a99d4e2233a601276de64e200e26b9a1ca843631f67a61bcb30cb8
z65ef99a30e9044080a3f355e3b9da492ca54d358b1e990f9f684e1dda49d2619ac5fda165b0bcb
z0a792556344a48293ed946ec661039faa633cf9c0eb01204c9d4d2d990a5d8caf8027d0a5d4eb8
z1ec9538bca3e664ae4101ec3feaf416a23d4d7a71834830d5d9404076fbb4257144596ab4aa39f
z3831ad8cc1c336cea09987788710b61be5d3fe09a1a2233c331ad9db1c19d8997122d23c70d9fc
z325e00d248905f5b89bf05fb45aed952f765768925092c6c394bc2582161c285822d16357f30fa
zd8eb5b9ecd6f2c1b80fcf34ff691bf0a75830b6d3f9426f7019dd7add69ad53757f6d1cf91740c
z70fab5dd9bc32be66ff7c41721d560e5d8bbae4c2a1fe52fb1109113699faad20e17f81a677507
z2316202364d2555e01bbbebc8cce858600d991b98d2bd2fb51c6927ac0b12ea2d1f929443f021c
ze849db71a2f65f527864333b4136a69fd7967ff368f218e181b10c89f000d41e2e7e5e4e144f68
z00c5d4beef8d9efac3ecfdf5d2099c8debf0716fc3fda17dd04eb5a8ed9313efa721246d1624c9
zaec1352cd9a8109d6af0378060a2dd4e919b8adbae2f96619909fe403057fc09053fdab42cad2f
z12f18ab8ea8b178c6e8f0a7e653fa40f951349954bcf357557f8d8c559a551031759d5535dec52
z5fdda2c5b053d6aff0eac4fb85c5254d9d50b6acf0382978e81d455175f94966f2db14feefdc26
z92193bdd329c66159ac8a069f168fafb3db899072014f15f5d19ffe26b7e3ba7a58b49f22473b8
z13c124dc49c18f1bef368be38978805cad33b13d96316f378879bb87bc7adc8c23d20a54840cc7
z18370da2aaeb568d92faa9af65fdc91f4fe069b8bc316bf5f0262e283a21063fbdf48f02bfcc1f
z2265a95b7e0a33175c5930c21d5c13565f87162c6a345a8e21ddf5392f36fec0b47a2a13870f8a
zc51ac47598ec701d7c22286c408cfe63450ef0a7e5f97ba7d5076511326214940aba7232785399
z87b1b7af5f43ed776349a60598ea27906b389b69fcc41c143313fe20b573c552c51eb8528bc3b3
z1d3504d15195d18705072ddb0b6a928808e872ae83687140f485aacc0bc1639a2cb817beb1d4d6
z558b496e8327ce2a9729199797b409902804cba46691ca21549beb3e1eeb8f22031ae517d466dd
za589e887e06bd8f74dad8c972746506dd0c0e96ebe1ffb080e69e3433e6f8f025f86413bce80c2
z3a331ae24f9d52d737205e7ea3bfe9c6555b03c0961f859a2a3920904b727543bf85155cbe3cf3
zf8c3bfe1eca9f53a2ca979cea271d40cffac66d65cd6f719e8af1b7b1d0803e56921366ce39608
z5658996d05fd20fa454ec077fda353ccd2ab9364c7ed5978c191261f3c6c8036b7136ef6e0245a
z715c418c64ed93ad0058ff7953376de4e5d26d98f18749f7183117643a693d0980506b62967cb5
z02bd70071fb0dd7fae9f20d92346a32d355c56331dece4dd2d30bdab89c26f1a88daf9c7266467
z485e16c2bcffe7357f6cca117a7783b0f436dff433f903b100b6bfdfb6685438e5d9bf08b3b9cd
zd2ec3d84951413a956c866da6c879078f4b1d71c9796c0228de04e7aa5013f696f6570c4a47e62
z6b3e9c652d2e3ed5b93b596754fe2e28fe7fb846d059bf3726a19e6a54854804fc82ab047b8467
zffeee19c192667ab3056d497c7181dab7882fc1ed94ce91cbbac0ccdc30cd2bd55d4b38f5295ce
z7a77eb2c3b2ad7f49771862b102aad873ba51eb9992f1731af1f322570aa814b5d223a609d3884
z241dd4d591485c53e14b7e01d315ef6b5936644b58de7a45a3fd59a9287adb11af973b24d78eb2
zc490704d73d9071051a4157dc6cb89868ddf95cf0be60b19b0e0afdd1e5255fe3ace4846e48865
z6c6375001fde9a75df43f613cd78796a1564612a6ed11cc4cac99a0dae2766d3142f0a005206e9
z1a784a7c1f974cd06f5f979758cb0e91017dbf1c99f24c6132d396d1b220156d8150abe3c0d2a9
zb732ed1a175bfa7ea2ae5b3d1b417b5ef6dd797685f43e7dadac6ec989db72289162a7d5753e76
z2b571bf40307ac7c087cd684ed2e70c552a645a50f55dbe4d59d4aaa0c30c32c8044c3e04b0471
z50486deb9fbf02650e83ad956f83986d3c4e412d1e1aab190c281624711ba7aa4a5901458d3133
z6bc9b8fc5cbfe94f2e83066250708b9f4a5a30b1d80f68a35a75b147dc73b88a90b0e154902c1c
zc759f30323f647acdb002d8473371ca36fcacb085f513c9e6a182ead02bcb86d257a39f32d5040
z3a24b2e35f7829260d721b372485b916374d4e8d708ba32a1a2d4fafdd35dc87df114a3a94fd4f
z9e4554ff8c59cae3a13861985e38f3c1ced81f62c847a214f50d1544756f48cb8fd7fda70ece7a
zd2e46503290341176f8aef1a5144e2377bf0acac37b85fc5e27f9c1b78857a3926a6f50c1fc52d
zf6d1890039efd926a7bd35e1151e02f2542e9be13b279e7b4ea68936c159e49609de23e96393ab
z78418392ee55dcba7e4f12dc8849b716d92a4f12338e20697033dac9f7d64105eda9288b697cd1
zd3fd3c7979c89fd697b12068794052766b669d00383038704cc466bc5da6bc9189b0a93c76cd70
ze01a91f6921744ca3d88daeb799957f8913ee618ae2b0b44017f40faa974f8d8fcad763ddc4a17
z843a86c353266e496393356a65d88623e477e63cb3027e728dab1d7f8b4faa6ad77ed168bf4317
z3dc9554a5c5e82bcdcb31095014989741e5aab5366b4442f8f36e2d9887923fa862e00f4123ac3
z075757a09a2a7b75e420b7562bc36d0e8392f86b2a831c1e4107ad2feb3488a7117341628a0ffe
z754d8c842eb926b38f16fc5de9a7e10f7cda537de4512bc0757850fc5a8a717370d4ddfa82c0c1
zd72993eb176fe70d482277db56f7fb72ed1a862cd1b7d948606842e64e10c6af13731e2d78a4ed
zf3ac89b3103530cc5065b544539ce4d9581aa41c2c001557ab1b4dc45c9e0b07f0cb96dd73ddd4
z8c84ba0ebbc34ea151032e73a0cc24263cbbef153239279ace5bef9aff3f3435eabc3250fbd3b1
z555bda626d01217ca52cd74989525c854592178c086154bae478799ff50de1bd814806a8100cb2
z3a58c34a837ae4e66954c3055b6a014ab64ef5fcb010e64623a50238cd04327939fdc2f884138d
zefc8ac27fc602e1c4ece342a42e59de9471c89bc305d32f288bdcc6b98a79cd11eddf964bc76df
z07405043badc24453bbabf2cedb2a6aff4c265d5eac9cd921463e1629aa7696eb5c643f6b3595f
zdbf882c0e8707657e5e1e91e6a6f300ec06a4c2e33f9d86c071c7eb0157f8c2741da0e7c2e0d3f
z595dbad48f13f716129a142d17a43551fc62a0c83ef18b383a3c3a9540587cb79820944a4ff1e2
zc33c28598bc7b709ab9c8487927cbabb7cfff3e033980e5ac5f319fc9b8bd2d2131416a48baf3e
zd696953b68e0a2d16c6108feb2663d3e7666bce4508260ebe4259bac96828afb6e0d5bc3200156
z40d653f435d09d5d57c6594f50bc6ce06a166378df4cfac2ee04e320c80797bb3e2fc495a43b03
z5f04140628595ef1f5e62e1e1d95ade8a31c9e159f88ec3271b5f6d5b01450c49ef058e750b6b8
za6dba7c692eec715d24737b32aaa3b6b631ddf077f45f701498f08933685cad0b5debdff4b9a48
z21b28295d22e3a5eed90411b3ce41298af6f8a78bc8b4403c5016a68042a93f1ec7b8d19ababb0
z60d41192e61ecee11c3674b671cac27fbda08c0154372dc996e5cfe322cb2555b19261cfd4002a
z08c1aea320fc3a9704079caefec4668774f20618d7f37f48865b6e5df751a30fd2ebf4a8bf4d9f
z84c6503bce38137ac093342ad119115bd3efb29bb27fcb509446d44ef27cc17a610b4f58c19076
z0da58ecef8ab9c226e7aa7ad82c27deb7729076ceb512e34f43f2c319766dfce622dca77d2da2e
z061cba1b6ad0630d8b74f1bce564c05f42a4f4639c56344921880d99c41da646f8f0d70e6a28a2
z59d6222e1d44c4d6fc427a70978afad4b75fc01c843304852c3d8e10eddb615fe9ce39a305d69e
z7280edea2357873b0aac7da3f0cd98f881ca8b8ac70edf209cf984e125636a049eda5143fe75ae
z8198269a694cf4d7d3e1802d1dda7f2f3673bf27530c25f34cee89db95ed1c8bcf07325d22834f
ze6ef58b7d213314d733e75c2a98dd4398436cc36164d47f519a9f60b34cb4cd2a5a4faa90796ee
za08c7bdb63aa343f74debc029f7027943cc9fed64604ee521503c3ea070913003d698b7a0fd528
z320f4c79305b8cf7a02d619062ffd65b86ecc289d26b287d93ead2f5ab4f56faa6d17c9dd918ef
z94dc1a370cf0db7b2129b58a6d8e4f4dd981754c5822f48e57adc3e7c11f691329270b5827df4b
z2f77f3af33d2e1c04191c6321fd50c422fc1468a080d447a34e53bea9d1d125619b5d9f8cbf63e
zbd1b3051bd85b12c2e897dd9aa88315fc8a89d2929d95811ae612805e3a224e04ec528b9b6a7fa
zd83252d3327e24e582f2539646dba0196562a2ca54dea20517d9100c5556695343b1c8241c1c04
z4441b5fed9319ee1665ff8161a8280c0e3df0a69f29faf93941e0c8a4d956be57a9f4dd9851455
z8f6da83a65a080beb8c08b6aace28cdda0731c1e102c621da562c04a66462341f8a03cb2697728
z982ef6027dbd203410ecc10530036fae739be7be6933db69c2b3c62c5dabe9e254ebb8d0728ee8
z318cbeb7c6260e2557249b4c1960b090264ed3fed6bd92b0c0a962140de0d76878974d7db5dd10
zaba0e3bca66cd462a455e9d44d52dff9d26fd5fb642bfb312fa669a041ef53309ee0553454d4ba
zd27014aba0d7b904bb165923355189f4142153aac6270a1718416da024381103d04cc3c714f52c
z8491eed69f1bc439f4e857d94e4b9cd195576b6417a3b914d9e557e24007289ba58f30ad947b67
zc4135aa23a835ea967664ff179ab6d321754b1f927f0f05245805f73b7a7b0347aa43b0051ab0e
z2ce55053fbcec7cce9f320fffdaa8032c40296f425bed8516ba95775ef5b9b52a4eabbd486f631
zc48883f75ebd7e6cb3c54bb6e84b43d0a2be70fcb2103650e02d98eba5c694de5f3bfff219595c
z9873a757af9b8ca430d1ba82ff7dffeaceac1b0fb540676f9c0b3abe0ff373de428b6e55717324
zcc3e135d6c488f04c930d5be6ea361a7a76c920dcf492a5f1ecf19f9550fade2f871ad511b4c12
z3fbc5ecdf9deede9713f6f71429b8bb9eb32f2f361c4d5b1ac1f226ba6c6c9b200b377a67c3804
z76df83ed19c01677d3f3a704aea7a04b7755fb8ca76589b9f0fa75fcb7c05a7b704c311c580ee1
zd478420f60666aaed08980bf386c02e7c8702580e20c4b34e0ac4a53b5a89efa18a02ac7d397ec
z461c365ddf46b1df3ccf6b69eb810700f8715b05841a54e918e0ce3915a818f257d11bd5720218
z87870b0dc63fb80c66e596f1f1bc7e553e2d72603d7ac2ef9bee41c2d6e441445893b35bd485be
z8395c6dc86ab9b65a37c336aa44423badf7e498a2942e79532243f1be44abbb04765cff98e3c38
z8313e859f3052eae8ec4d44401184c7b8e1dd2deda7e3ca99b8efa28864fa4f66068ac169a4711
z9d117c5243436569bd67a01ab7731ae3d78d5b8abbbb1a11f288c17fb0e7be03ce74551b71a90e
za691f74137ae17b9e90548ebe3b09a645c0ba92a6f1bec664c85c571562cce4ab563672f963a78
z16f03ace43409dd90f8350d161b9f8a23827213ec5c7165d63856ee1608ad1ba2c9b7eed2a2558
z35e3ab83072d2e823121a5b2c1ed61667255cb8b93a84b2dc867bf3cf1c36644236ff2fe8b35ed
z98c35752495e116dc5e73b7398a5286dab244d4e56a1bdf91f3d3564e1f5732223a98f8baff229
zbe712156811d4aaf58d50177e7a10f88c7e53afcb67dae19727503899d7bbf0e1c8df039acf11d
za060de21560caa919417e4c1fe2c83dcf20ba31a29eabb39b52a0c3ee512d0f6e0596c4ac2e9c7
zacaf6d41b9cd8947518f7e8826160487a1436b39ffb17fdf4b54072e5c035fdbbfd0b7df9724eb
ze462ee04a998e0f9ea731da8e14465cfb14aaed39c71d00cc1729f912982a89175776cd12bfd8c
z28f976e5ab7cb890b7b578fca07061fa0ac8b1820dff9143471fa59175068b4274e4979051e558
zd866c3163d42ce040b811e6765000933e602ee5be41644a98e900547b0b69d0168c4b81865d7ce
z6de0eb653cccb9ca0cf4930c243a8357018b75f50109561d1b18728d1ed6d7dfef22ce4be91031
z9475d97d0f5455659658f75d1a2d1a082516627d266d3622a543379ac1702eeeadcba975b71af7
z01c4c63daf444be45c97d91a9041031191452a02881cbbfc361cb7dc0354c01fbb94eb06b29063
zf1346059104996afc6c85555fdda222c65938d94cd8b060255ea845a9853882badc9c5119b9256
za5721a03471de1f342491f1169fbfbe7080482577279ce78f678a7f5fea49683249e17470c490f
z09129850519f486be8a6a675c438436636ab67a465e30376bcb580d08deeec0da40dc8aebbf6c3
z7ef87455aa6b5520683ec7bb4e5095731063227513e3c641f556c50c63478e6463ee298f7df818
z3179f5277f8ceecda0cb4286519ace4133fc4ce249d9e5c8efa4c18a1d322fbf781458e86b8b32
z6937a49bbf8e986e1aca8a12f98bee45c074f6c2c9150b472e18aaf416852d2d3842d3ffb7f906
z0ae8561273f53f4ad60e70ab304e2abeb06c11153a029b13bbdd4a80fb342206e1ec09c3e3d8bd
z28e8786ddd7a7fe762c2dd471b2c51bd76371df2f6ceb9a500bda85ee009197961949cd13c3be3
z71ae095db5409d61a742a8b8f433dd996fdc3269f3888400a3e77a589053edb873c2f114417623
z83d8a43ee6b392d8f38fac813376f5e0525c2425f0ee6e47ea9f5e6461c8b8e12a746e0e28608e
z9f8637d937f284a637bf74c870af4a28855e805042889c4795d34fb6d75a32f6651bcf81e17b9b
z0be9c17efbd13a6c4dc0906aaa81cf20b2553f658325188cba369d8a721cc56b2705769ec07f74
z5d8ab1536d65d0bbf1f5d7b5eaabae90353169f418ee1e25b8ed8518223bf6223639d39174289c
z285c219cbc45b716cbd29730cba4076101f77b1e344567bd3136f6aff539204e18bdf8ea3c89ee
z491109991e35bf3c6be0bea9e53bb1ce372cf92b2f4aafb8bc5e1de336c731b038d30a9c78a82f
z35ef179d02c77fb389efdab1de7b8178d49fef9bd5f74246eaee4d50b0e810bf0f2926dd7f3dba
z7a1cde799f04d595f8380cf6f168d02cbf95f2f71df043581ac6e876209338f8289ad10ee591d1
ze5aba4600e194c41d96fee7b0d20f782a42d9d36298bbbbde50577bf978fe8b017b569f21858ad
z2336c9f0c89da76f8dc4b819f78e8e5d4f6424405221d1fdae2a892109c2079a798689c8db97ec
z6799129a97fa306498d7b5e1156e41d3fd8f973a3e2f140c7f55f1a654425816197d515ccc2278
z26cd1f075505229d8c67ef26541b7bbd7f5588ec642b6ba7dfcff52b0f7946f3c5cfeb665478da
zd97d4018c5660e787a70abba16949cedc9052b060c31d11f54944ab6014c045eb4f5158c9a7af3
z41e900cd29c6eb9953d36c29b9cd166318a8a157e3a6cd9736c5e94a4fc16e5082d5a17fa4dac7
z78309457c4fdd8c39910e595c9f3e4e5988a4101755e0abe4af199d3563b024a854d4cbb0e6db3
z286c3e5613813b81588adf6c1e714b3ce52f2efc4c83b6d8565790386abe10305ec2263d010855
z288ef6fb4834e1b84be623d84f5e0f541d15b9a67798ea16bbb51bb93aff233f405eeb4bd46b6c
z695285ddef09c79c12f9f9aa8aed91098c5fa4058ef9009bdbba3fe3fe2c9ef1378fb81b74a390
zfdc86c52665277fb75d92c0ffc7126f90d88fa19b719ced737cf71712aa4fafc215a8bad6dc396
z6c7c5b3b2dc9c532b3e7a5a5adfd642a14ec4ae6032626f8e9124d8fd5917247d0e1a122af578d
z4e887b465e18d443230255c607580bad7730b66a5c04448d2a100793597ac12f25cbd1a178a569
z7860cc774e66818e35fca14c7b2463363653704b954730175d57912dac2b75c649709e774148a6
zce9e7a90cbb3591c6ac7634d893a93b9589c2bf02b99abd139003fe698931bc0389a9a82625732
z3c4ac7cc23d796723b44f0c2d504977b086caa8fd730ee77659d81be303d4ec3bdd00e6697843f
zfa83f441e928342d5bf3d5b3c0b8fbbec35a8f7b81cb1b4349024354e3ca9c7e89af145023e2ab
z0242905422bfccbaa7e75f937ccc9efab935e10c2ed973fa193327d59446599f9adb2e03aeefdd
z5b051a7eb7a7ce12c74ff4caae0854d5958cd2850042ed1551d19ae449067fe2821c79ce789429
zd2c6011678e3d6c0360ec5826038818ef4dd7e425c1184fe7cc93331b575dfee72b452a1695cda
zb8e9aec102c570db975592c0c31863bbff4f6a34f1c279ec8a4baf5c368ea05b78cc49ccceebfa
z9d323e60f835f264d482524272b98687219520d92630dd91e13ea89048a61910c1120b6bf47280
zb8da15dddd8795c7afc40f1d136c9635de91acc16444b852f9d69f0995aeb8dfce9c6f033ba290
zfa4b6d20c02c341d0c89c8544b0c50ebbef4610ddb84b2d99cb65579edd0db7c4212d08e7573dc
zff7a156e91fb7c7bf048e822fa08b39e4f11e49037a815ee3f23282c564cbc102228c6fd8f890a
zf7695fdecb6161d14012e183a3d1a01abdb0636c7a51810a71a11c7dc442f319c288cc83dce6ad
zafd5fa9b53cacb05dbabcdf3c38f1dd9041cb5704510420b0617e0217764962dae0344cd9ded2d
z46e3c1afa90b720cd38badaf720458c520ae6a0035bd32542080a64cc58575ac36607558f46ef5
z3aa3c6bd763310d81e9256add6352fb30d3328fe99357acf14ba5a764eef998ebb701a58d54ba2
z6b5b8b2f5f907aa6399ea08c916c1109068a6291ee4ad5179595a4fd80e00379c6def56854cfd2
zbe408ce40a0f34a8f415e3bb09010112f031d434ee6c6db0d2c2ccb6b7dceed76dea95f840d916
zd507e66b42a770ceff8837d77802cb15ff458f4ea1e97649e07c31db569487162664ec7076f293
z34a184a50b80fd38f3e5523c7dcf35b7d0be90775c11750648ae3b34fc933fd0bc8bc61ec9b19b
z07bd3493b4731ef0a9b2b84f77dce6095e05d6b961a09c0afcc5189774c50ea91c9eb76e0200b3
zf591d6aed3dfbf5802494039d309de2f5579d12df9cc712f6ce91d261335fadfbd4df0563b0c33
z1cd64f2194039da3e1ab2b17d00e0b31f4e100503d34e775ade555b0aa4173ba4ba603861a11a2
z1a86f75e8ed346c8cdf9207b1500eb1e922ad441e555f377c71a008b89e677f3152c679710efd9
z7c525a543ee11ffe446d947c7262091c2aba484afd2443087c25e9107925ea84fec451c94b1cdf
z8b58927aa0ae118798b7f84f1f3e472ffc6dc9d6d3c1a19a6e5b3f907b56b32c233e1a83c9ff7d
z518ec79ecfd0e194fd81452406b396d49aa1ce14a4967bcc20d3a3b9663e79df7d063a515dfc0a
z8cda1840052e46fda0764fd595b9b733f19f20fd526dd95803f3dc9cabbc5e0b7274987cb8918c
zf5d3f4a640e60cac0569a0b515974895f935dce6938d325d891667eb307c5d07e15cea175d1c30
zad34dc02cdb8e20081cc8715ac7290bf506466636ad6190e3bb0e02a5089d4879257dd86464540
z1ec5c1d576a3cba0e3fd807d6fca92610b6b17192b78e9b46912ce274e2d998fb2f378f65b3fcf
zfc1b4ca8a5768dc6b061992a3ce62a636e3716a2b3d53de0e4cd08ddd0bebe28e25ba30eae3b73
z64cf8864eca69d731231eb207b405bca672a5826c1c5abf3fd1e20a9c33d5bc4a4c15352716c22
z94a4de3602d6713d3a3089af2e0ddf9863e28b2d3f9c25e6162b4b2ebeb50eec6c57a00571da7d
z9cf19483dfb504a48776144acc422ea1566ba871cb880aebca30de33ca805e9412a531cd250fa9
z408c9b8612079e6f1b37b615e129b658eee33ebab549f9b71f9e620298e9733d50e3b10dadec71
z8876b5ab213497f522db83a728273c634589985a564d34dce144986b53e2cea88edba1eba6067f
zc8dce1346d967f424a861624e65e1629abef281be9cb7691eef7d8a685fb3df9072cb87e30c853
za8695f62b48404da92425ef9cfe120d13f9ded127ee47334bc83efb22ea29501822f30c4078672
z724a816344e6174b8d61d7d960309c224d292c571536f94f5366ae3cd65c6a9669ec7a745816ef
z2179d42352978540c9ea1e4fc5d319da952b152b6a0b9a2303822c3afb2d04724804094f72f3a4
z277a09e2decee4cbba28a92d7efbc33cd109aad9942037b70d8b6fdad15ca0d2bdc1ea4235aa23
z672bc5539061a942488dad8d70c3a7e7384c8edc74149005e8a930d694a1b16debc84b4275eae7
z1127a95c87558471cc51a891ffa7836e2e45053f0a23eabea25203811515b3ed67abf7d7fd366c
z4ae6594adabba1eac2aa097c8d485553567a6a8817c5a2b535cc9b078442c71678e15df84ee49f
z19725a7c9684c45548a300c79a802a9542f777ead5ae3d535eceb2103d7200b4ea3f091053eaa6
zfda6889cce5036c5d978fc3ac4ad2a159c9ab72b9f1f749e9bac238812321ef31d3b364cd68fc4
z700b3f35c6cffd73f350055a874c8878844361a34598430f18e48de3cbec5a31590452f9aee3c3
z204cf6b3d020e8409207b9348f85b6791886a21c84a0083d1d423921e37d0a0cbd24cde450c77f
zc4a9fc883474c2bc1a45406d46151f575a6fab1d838a9bf5a4152b175d56a02e0a26a0b5e2a1bc
zcc6e3f1c16d1dc4511eac9bff72955eb69b4ff02651e82f64b95cf3dc83553ec0ba832ca8a3a28
z86e62976a2ec1f87a8b41af468a20955b3ea03f4aa9dbbc641f9d927e28c820a7ba24954f4178d
zea11088918b7e17cab6676d7db2802eeedcd21900ac70c94b0a221cbb26f3e7603ea187ab50fef
z68f11ba894cbbbf6ceb781596a2f63db1363c34728b9873da1e49ff7f8d1c741d8078cb110979f
z2f8beb865e696549662515de53dcd9f2f9225a464ec15fefa41de84e94233638d417a053a79137
z2b9b98a881eae57b881a9b55344b20e7ac8003d37cffcd673056c518799c79c9fd40315f5d425d
zd0f5b9fec67a532f7e8ba9b8ef4f766ae4a604afb28e70e621acec26aac41e57136606ee5ceb39
zebcd8f807a0acab6bf60c471f5e8b0b97cc4702423547c8299a5df66102121b69e82cb54ca1d8c
zdc3624bb50aa0eb0cddd2b2241ea19e11ab4a5f31a5de35ca42751cf9cabd4e94e3bbbb056be3d
z3b7ad63d079794b2bd3ba1a93808b96888c8b3b8758a90fdcf78935e5a7d73a3669d12dc793eb8
z01f2b4c22f063dc0e25e38e2ff7a82df388c75cceaaa3a047b4bc61462a47f80f8b2d59e1d3a17
z7586b8f00ba6542f7c7dcbc7fd62a35355e69d62d81e3943c7e2ec0efdcf5695fefacd47e72dac
z089d2a45754e3ceba6b34b9c311d6e16d91d81cf8a9402e8866cb873866296a55a774a9e8bacd7
z2e55655099b8a626269d2b02b2f58a8a318f9549b174ff0d302530456b3895163f87d83f840599
zba411d4569395c15d42e128929d499fc19608cec1e475d888afb33ae102882f62f68170c268060
z36be8d18a0e5b22288f86b0f8412b9b1bc6169bedc286ad3f877bee52aaa8b73fafcd65f0c79b3
z975da2c67bea64457eda3dc568392d02c8ce0f52f058c6429bb41fa87ce1cef2044173e9126181
z6e17e73a1b2766f22082a6971c7a14dfd41f98381bfcb12e14dc1b4bc639579363e609ee027ea3
z26d13bcf4185e36acfe3791795d4d1812815f2dae66cf88b2efb15c6796e2e3515ea8b91539d39
z7b44dbec03fc2d893a3e3a6ba88503a3f6525a148c7153e921f6a4697619099e2bf6885054e84e
ze880b241f26411dce3767839c10042d7782e5a821cd34a21753c592e0e372bb332d53a85f0c610
ze21deb946771bed017b64e0a5ef7b0a9e0c934a37a15180ed25874fa2a47b0f055b80fb5dec687
z822e2885bbc77ffc39fc92c36355ac5866959bab31c7578fee816d29cdd279ad161874eccb374c
z786ab290369a3803995774ac45fb1afa854d99409165e3751de72c73a1c999f67c3674e0b5f928
z1e50ad9f036b69df4138bd7ca774728ad18e33067374349b2f7a02bd079b3c969e7d33b9a7af58
z620bd2f3b9f3dcc38e00b30d1c0f0496662c805c23c97649d50ddc7ed4334a5b652bdc76a34e9c
z9977073a171069e1590668ab2c7f0ea6ffd782678febd35533367c63ac571fdaed05a76f445a86
z6a4e926530466db22c7366d24015fb6f13b8fb738d69612961904baa6ed665e57d6a06a80cfffe
z7f8273a025c94506faf2a3c0d081e92b3a598fb6ab17630649043038025ccd5c5ac36f9d956739
z1ac555ddba0b248f4ddd8c4b0c4a8ce881e5c3826a2baf3298ec3905efcb2e5cc4926f08295f03
z1681ae5a13297f5004a9e9343b8c9ff3f743b5baf46b2586588a34a34ebb6239096e52cd4cbc89
z3a23518dcbc03a7938e04a8735dd58aa00ba563e5dd08ce66608b0d0191783aabebe2f53f11215
zad7d73db33d036a74cd73387406f4f56d4af562bf25986da7658c6b1bd254e1653a55cf37afb48
z4f045d0abf072cb50eceb63b8c6965fc97640f2ea09fa06aefda9bc5e702c0844005eb54787bbc
zca81fc4bf702072c2487e6a682dfa1b16d4961ba965dd17fe9304de7f46e96bf839e49cf6c8176
z42a175056550d540a999c8077624c9482ad5d419a7276f3ad4f310c46daf87b095f54d2364a681
z40c32edf72dbf55175f3ecc408d1696c6f2ef77744ee76bf24875351ed8f27e590294eaf2a50a0
zf7469297779b09e782d558c988a3c5fa7f584f68433983372a9eb8bdcf8e9edc1d32c70870f1b4
z28ccacabc9e79bd58b41463800f72ad50e7fb5d3b383784f78beffbfd7989e96ac48b1be483fcf
zc72a762ead136ef758ffc67a5a32bec5d68853e7a4ef3721292698c6205e2cfd7e98c3f388a650
z6347dcec6a4b6fd8584550991f95c35e9df722e67c55a2f5b4436a6bb3324da5f2f6795e90f073
z54401a845679fa706c846053cc898ab2aef5b2b4de3f52f9c00598f8f59bcfdb6958469868a15a
zb5507bb5139250271656064e149aaede4ad9ca9451376194b4165d175e839d5b421c20e73d3dc2
zb9479967f4bbd86b56dba6fe6f11614f0f1371e73504c225f472da4c04b4799b45fa32e0cdc4ae
z220e9d1dc6f51917ef53908e0c707ebafd59d009da402f2b6a3e14096101284acbddb33df8ed8c
z566642d6040e1b26f3ecfe95f26ce30998a761489e8282aa01507b68be3f695d59d2d1e9372024
zaa7980ea68fd3c7e9b2c5d6fb998b9472527d701390a58e55e371dadf6a644ae34be63434fcde8
zd045ab5330517c9b78ed7cece74cadca360f155cb0371d6f502e7773aa886f44d995af70ffeb12
z9420c3bbfbf0c1a6cd3eacdb495a09aa7320520f60f41389602cdffc48d65c4d9f9fe15c33c1ef
zf973be73a792918817ba30e37ddfdf84bdf8ae1fb47a94c5184c7399faf3e7b323f1bfc59cb9c7
ze5b1fb2fb61ade9f64fc1f13eb3cd5513f9104f740345839fc8e3f910bf70339eaec0b8917cd75
zdbb623e510f9ba2430204a8fb8b2b6c21c248df6f83c934c98f42586728e4c1f6157ef29866f06
zeb06312ec494a8ade25e2ac71afcb757e95fcc98d5815efdda933b2f70538984a7b2430d63f1bf
z5c415a0ad22d3eecbfe7079aaf6f681659e3b655af1c18c960d0b44ca95fa3e8d6dc5b23cb5ddc
z84f7363c2b3436207a5310e2e3cf577c2966a6f74ea2e4d4af58c168d66437a665d16f033bea48
z13dbb429b9a1773fb2d392eeabfc3d3c8af6acc1b5d056dc1aece50adea69d2663817789430370
z972b50510bc247d7bc399975f7e4f937fd78ff8ff640e44e3a0d44c6575cf0543556557b815970
z3688da865c89f7ecce90bec006c6858f1ceda4b1d7f09e908e78adda9e8da69b7798cc9fcac210
zd2af3566cf065481e37ed86f29dc17efca3f4d85f631a53619085639e500a35448e90534bb1234
z11eec57a8efe57b8f039c69b5b9d99072d024b85a59087d7fc7078fe41a4d24e76fd92d36d27bf
zd501c5869a6f7dca669cb636e1a9aa386b93099b22f9424fbb80c8c6870f3d7cad2d8992ab3297
z8d05112bf72517c8fa8f32d65272d216f5ea64ccf590c0a1254d365cb0b94694a4c63f03722192
z75863b9c3d343212351e962bfaa213a3c107f9d5be41cd9617c4b4c61faef2130f243c0c6585ee
z5b0c1cab382d48742f8c97ff0a03793b2ab53a1549ae708b63bc79a9b7419b9311b4c24352ccd5
z4efde8f3a2b77345ef302a98b5bff6f64bbbd1988a07ecdd3ba5fa216908131897cdcbf2f0700d
zaad2bd908beb2892958ca4b96c9a26f58937ed064f738a6425c71d79a5f364c780c3428b72c7eb
z4aec580156eb06b1960e40ac8a05594883fcff7277cbf9f1490821736d74b4b21ef6ed337cf639
z3eef90d60ceaa0eef1faed6237a9293145e777223b8f0f26110f82b96ddea46c013a45ef575ed3
z6ae8a847ccb2e21412da21024c5dc93b2a634eedc6b47efad23025fc02c5a216ee85de6016bd72
zd39b0101d22de46c50343de99974b6a97d4d8424b50a78a4760bfbbae6081f032114723b8faee1
ze4c8d78768215ff3a88fe9723a2305935c119acd1b790e0a7c1b3cc60da08ecbaa95962af2d78c
z5148780e6f24c569fef2fb69a3b2c9d55d4b65cc58db4528a82be7734109f631383fe3b3355f57
zf2a4a07c2cd8851388a51d8c4a7edf13e9ef601c16a7ff5d0c3aced07545dcfab12059d86a5e7f
z7bd03c11aca5aff18a54152b086e73cd19d6dc81217a56c4ab199bb42560edf7e33500ddb7cccc
z25ac76e870989e19bc066f942f738ae3d3772c6048034a54d32288f7005d133af7f601c21f00a1
z4277c50d47c504e809ffb49e55e5a35e272ece91bb37240ed249f60da8adccc5bd1d4a6852fab6
z1fd8d4b3f952c5dca5c1df3f31807538385c6c2d8713b1f73be7c92f43eff41d61c600464e34f6
z929e7299ff35f81fe7ebd2db64a52c47b614eab4ed578475d62b50a91da59b54c46461f2036d27
z056489c2bde33ae464c9e31cea41e99b19b2470ccb4216cd04951f61d7676d28d5e0a398400fbc
zcf0155d8e1c79bc28ab6fca29e77f3a90e0fb0155b5591ef5feb825b36db62050ab8d8539ba416
zc8ff9a7d59b5316c4a5b4b02cbd6ae581f391739e63c358b5050114dec6c2d2dbaef3f03eb2e4e
z8c77d34992a9778f995f2e59bd758a462abe5c71045450e7c4bc4ede274a9163d89850cb278179
z8dcdb4f764cb94f09bd570e23f9ccae0725325e064716cb47cb289806391e61445e6e431b40370
z188ff2e8c7b93227af5706e3b3de82c97c8073cb3c60b6e14376bf73a5bb9ffdce43f92216e4f7
z66587a6eb6de23ace332a303c2b32cc15d0196c77432caf7da530c2ede58439f39eb27707cd35f
z0361867e4852b93627ce243d19115f8daa66c001b1ab2679e9292fa6a5342df9bb4649f45dcb5b
zc09a4487c25fee33ad4b950aa6b84d12ef6dc4fbb43d602a3ce9c72f476881fe5e7cefd9851647
z23e035ce717b0c401a028b4177987afd5dd68a1b6a14ed00f68ff9cc0d5089c88a49906d37cf98
z47c6d7154cbea24766879093aa761bc5cce028fad9d02a89b3b36ccb9ff19e89fb1cebb44c164c
z49c39e57999dab92a4cd7fba72d448d0b035c4df273887bdd355b23037302393054fea30ad7e06
z29ab48de6ca498e343cdda8effdec95de0ab08f8b4842999acc5c170747650c909eddb7ca097de
zb06279371716659df47034e1461ab8f000165c73cc0d0206477425873003f4b94f07ecd1c2b40e
zfd2e8b16c1d11550c0271dce0994d0ecb41015e21ec511ccef83e6971b360caf40908da1178645
zfa61cf79ac76afc7f6939d91efe59ec7175ae121250cb276a95bf80972970ff94402280180a652
zbf948d5551cdd3476f59eb50baf3065de0b3666484c51d8218f0678e24185f3d3ebab3088314a6
zcbc1d28df150334a8d0d7c5e2f625323d9cb942b84c14debc519e6569292ae781f785f97ff0535
za90f6785f4492ed6bf8431946e1107b4400033ed2883d9be1dfa80f040c454bac56fd3c35f4c6d
z0f92e0b04450031eaaf1cdffdf72fb4fce83693ee4dd01fc6c5ffb3dda9585ec7f0e3e80213227
z8510af602acbda49ba6fd91340339343b2cf743e1d5076e2e34db73f3fb317d8409a85c922c060
z727c9c84af25a26efa09c0c0d8ee5ba7bcfaaee9c623d3f2e709df8e707c144c57d42934e3e1f0
z4973216759928b5c19d2931db03f7dd38cce5775e118b194314e572fc663a806a18aefb3597748
z61816bc00ed0981c4e33f90589e19b3e4232326dc543c52059c5ecc857532fe36161621de5722f
z48e59889ab632c083415487b5469ffd226432d8fc2ae28b6a2cc6ee9e73e81cfc884d9a7e8eab7
z1fdf0172adc17fb7ed20e2311aad3746f085d5cf13042f305cce778908d6d5dab4402b3a5ec77b
z4532e2dc08db74da56add7ad4288960dddc48fd8504b4dd83b393fb6ee65e5d9e676f6f3abc56f
z82aa6eabaa009c2c73d4283c2db99c7ae1e560a3936e0cb6d6c9e65afa578f7d89bdb26fa8b0f7
zb3bd96eebbe6fb5076d385323c5f85abf569495b48fe006eb27246061fe243c6c5f6dd1b4dba49
z8b094443bc9000ad368fbd7451c1224171f20abf9e71ab80c76d39ccfa8764a9d78aded074963c
z920ea0c7a005aa3deb9923cf898fe8f0ef8046a9f48cb19d6f68618d51cde63f82148e4eb376a1
z484e0d9737554d09d2c7b4e381b6a1a1410833bd75f72b5303349565e402c81f2a74e38598f867
z82e9f8be83c1ef3a5968acde81e0b3971dc762a129fb338f7fd8a64fe68e29e95e46bf86301e03
z93059b51118217a738c960b8146f6eb7ee0e25d13e68a96ed21e9f46704489395911cb7a6cc20a
z82008d315054426e7ed8b3f292812290106b37306f0bf2ddea796aeab8813a5e8c6e15786190b5
zdcae914234094304994746f82c6ba39a35ae0e8fe430a576ca2b24d37159146596430be63ce739
zf922b67ef7095f92e49c63feeee64f9e94eaaff8344e7fdca0b7b921d0cfcdc07746356fa70e92
z77179f80ac48b4d08ae64cc62dab021e57d9a68c77d935992d0ef9626b0b8b829138d337392776
zd5e9cd60e807f3799b3e3ab4acab1fb3bd30168278ddf99a3b09a273e8b25b8da886a419e45b3e
z2cf173bb767004d4069af6e166d5fb5a7cd1ede194b9ede9c13832e37a184777edb014c7ff6c24
z315c57b2cfb402a1731375ee0c905c68213e297c59a169fa3a72c21ce0fb842e64874d295fb848
ze2644549a36700ff47be2efbb359692ccd7e59096371e3dd9b988c436e99972316feb03222c538
z5fce793e874191fa36767d7e2ec1baf9600bf732e239919027cd038e4f53a8dc34734548efc34a
z3d9014f2f10b97e22ac1efd53c8d4b9e233787ebb5f4bf8449151d3cb71d2c520354a5e0f45146
z273451334ee642dc83fb67c6f7a2bbf33bcc8c57d60fd97a4ee51e50de5d34e13c50af2b217d3a
z81ea02e4f7e5328510023fb07cdafe5b4891834839adbe8c05f5c3f4715461f7b57394b15c1eb0
ze92b87c72165deb83c7ccfceae0f0a02314cbd91c58ea6100c8b79bfb9727c575b497997ac7017
z3b1620a440f15ce14c98e03222abbbda6ec452ece1b01cc030eb4a7201d0c50cc18c450ade465e
z33e5a2994c9a32b1e19cc393880f1363a7605e8700aa61aa6de74f6dda85d1655cfc7e7727c22e
z82e97a65582f97226a86c1ebd22cbea5c50093aa03bb4805250f204b7adcd70cd94ca63d4198d8
zcdec602e468105e093c7c98656cf3f96b23e79d4fd1d55e1993d2f84db55a140aeb40006b11d0f
zae7dbea4cb8174ecf7d0c472910ef5ba6ff4b03bed295505c22776cb8045112d282c072c70a198
z2ecf1998d9272a946296c49b37af87319f535bad4e9283469ea12498caa0388c409825c1585d6f
z56607c3dd8fb9917218e414074025b9d3a622f3d4f9e3b44d02edce34099b28e6b73ddbdf08bc2
z60ecb78c764d115467bb098bdf76b36e7c4ca6b0cf833dd4d88fb5b40a107ec7e5b20ea0768958
zb2ef92120b92ea854f3190cf3a6e224d9269d5149f0d572c2d5fb0c32fc7fdcd888ecde130e211
z19ccd61bb82f3d40601f6ca85160f5a13714798b49a5803c6687753fe8d719e1324f9d98ec1d33
z2a7a647962ef9832baeffdc441863932af840819bcc692cace2e1cce0b3c44e63fd66566f24825
z945d1a324ced8d15654c00e2177b252abd79d5d19f3fbeba6f2c4c70c20a5b77a11a49099047c1
z2374bcb11bcd557ce35a4a3921432ec898bb2b069bce58289a7233803b1a31285b15ec5f4d7bb6
z684f9310fdc6060a64a836c5c8e81060c5d92b3625d307bf5d1cc799f3f3d1c5d57e29719fcaff
z4d0a56cd07393a5b0070429180518959a5056db064f429f1e5d99cf2f614085c6fa74cfb026644
z4dbc8bb71bde9c22aba088cf15d57c70dfd9b7eaa5faec859d030665a7a231bde5f8c35cc5690d
z6ad1fd439fd2f7909f02f3cad72cc2f5be99a53cd48771c1ce6ebc41b0df16564ee1e312c27c4a
zf8c88105baef9d49c5551888101d7eef3c613284a6cae44bd2c5c859a46d96335eefa1f944707f
z8880d48a6937b04c347d3276d80f641d596027d134f760afe2d3ad4e1e30b17aba43ba0ac57919
z750d475e5c1c2ee63490ddca9def68aaabc580da28ef930a48bc30bdd4f385e12bb85c2d61386f
z08610dacd18c62dac4c80fba83b013a3567dc06b6b05ff5ebda9a56a593290298e55bcf3e5f30a
z2ee0117311bfd1c9504d4a8237928f2ba72e8f183bea5cd77e30fbb0aec3a90116f08cbb8d04a8
ze8f659b00c5b66af7d4b1918ab32bb7eb218d2f912611573059000b30ebcdb67bf827c49255a85
z35fb2f604c60a5e3f55c5538c561a7a4e082e5c2ecf9e593a61d5b418f8d96013e4836faa2ff93
z58526317831eb7b72ac4467aa275be246350cfcc07e62ea8dec24aeb30ac4d3a389345493fc864
z8af41d75d3bfde468c8235906b23c2b1a468c1534782ebb4c9c5b04ac3617aac58f0601a4a03ce
z454b6d55414bfebcd1f55d7d20a68689ebac931391e1e635c7e2488cf5a2adb6fd2e61b2c495a3
z9d2b5fd5d3fda2fad435ef2057ede22b5ceda0f0dfd580e3c4af2c210b59f3a54eca4f798a56ba
ze1075d773d06f97268d9e0c4b2ed7d02fd74b724cb6a0963c64ae9192f6944e059ab580d5576cc
z6906701cc72a0ada9fd1ac574e74e59481e704fd8ceb3920f3d817fd8f5d9b7e4f5f43eeecb523
zf4435a5ca32cbe14b5c5534b1784db752a932e140ca2265c3cda830e7c2cf3208f83f1a9c24ac3
z6cdb48f79cfeba5c3d3f84a6ea3a0d9ed8c51c6acfed5dd82fa8a04008bb7282000150a7f98dfe
z2a2670dd87fcc9a35fe8f53c3d7984fd7839be168474dac47f740f3a0e9cc6a411373b6d6c285b
z20db9ad20d92ffec1f67091b0689cbdd65fcf4935f158e07f638c84296d50688aa9c81a0e37276
z117dd29ad55028eb839dd4924e6d6f4eca5dd351d5360fc718f10cd09a56998eefd7e207db8469
zff3f7a887a7e38871239d620e01c05745d3b7ab21c6219bebedfc2dd68e6d4f5ab69efd24ea353
z79782a065aa6ef1c482e0a887f715dcb865c199cdcf8b8b563f239be04d49ea0ab0fb0c02ad4b1
zced7935ee5a7260b1068edb9d340dcfb80efd1b177ad235379633a1aa8bbabaec1fdbbc6e8ee65
z8d4042e5e952131df5d08c6ea8f111d36014efbe1a30c14c1210e6495669e828d0de1180405a97
z29cb789fa8d3e632957853b5c1a2673a8c06f312bdaca786eeea88d95cf1fb18777dc6db26da00
zbb9ad97bd7eb55baf6a01daf8e31db3eda82941ae154cd229e375551c1a5d53af818c9c94b2c30
z45a21867130ec3b1a3c4aaed7bf15bb461e5af18dcc7b280ac513dc09b5ed0c49928a66ee9f833
z7349854a340803bada371d309e77c239bc571c96040ca573212c9677b3f5e299f2c5ca3d74dee7
z281b8b2dd8d505c126305a446b06c18f6e41c76ecd7ffbc01614a1378a4eba576e0f0829b84083
z85ca89fe78c4cd00ab194ac66bcc59795627b11db4e03f3849c1e133365967772750ea049ef8a7
z70b297ef689f07330f0f422c605f6be5d7aedcad030d127dde8d1a7c9989b33e20f04dc4e9e675
zebf6e32a827bb03c418e0394385f87199a5e6f2e259237ebc7ef2b47b574bfe6af5671fec25b38
z6b00c20fa8125eb2e7b909592dc1c935848e1f6a032edcabd66a87ca023e1b70e2ff811d9ae5ed
z441a517dcbf5b95906a75b8daa5a95278cc743167294d6cbc1bbb372402c92050fd7a98aa39fdd
ze8c7342cfbe5d93c110da03f6360f27fe44741d754f3b11e95d38394f231399d0a941b66f04a21
zbe76e34be1ece47c5eec57b985faf65deccbdba34c5eca2037eaa8bca147236ea9769f9579b49c
zfd14000d94d56ca7dec61ae2ab54086dbeabdf82044091f2f8eb097c729a2d1161bbdad66b9f59
z183271c80b200421488bf83868317a6879003d7ddaa244c57f12b35dc9354cd71bbf354f0ecd74
z868d65f58b7aad7e30d8de31d8de16037a8d2d6c0927e35bdd289b1bf949abbd8ac1b55b4a4e5b
za45610c6cd977ce4a02fa2c8015b23b6017d16bd41eab05d1029b90a776e9a898bc6947f36918d
z1165497b131090b07f18ea9c7aaaa481ba816b0aa1f824b0b5e8269d0f077693874e777bdccb6b
z4ecd17127ef3389e52e852a6b1ea0ba9e164bf25214a7872c1b4949881c18406f22ecdfdc8f163
zf92ec107f8584b7a2f64bd1d17a59ae1053fd83f9bf6077bd6735a5f9447184eb7bef2a5fb8b20
z29acb7b8c8de6c4ebc4aaabb193894d46312de08b2c200a54c35a97132e5c64e11426804e12a14
z3f79c2ca37d4b8cc0e0efb05a90fed891dc7593dba264990a16d86cd6097d2ac62d588927d314a
z2c1b02f7e213fa09ae64a501e6500734118cee3f3b3563d2a1758b055b3673f37205ab810b0fbf
z5ba670ae32e7a2bfd4d24a2bd0a1cf8f03b511fb449968be5f01fa77adaa4089f681738178d332
zdd5d8fe8db3db94b479846a0a8bc51f2739b2872b7910ab7ff0d3ff3820e53259a67277f30108d
z86c0311db9f9800ae9b4e7c15482c7522fdc58899a3a13f0425442ffe21176cf7d5d72ccde6e36
z5fc7608606d68226f958b8c75bc2b6358f55ec227da43bb222bd481d246726400fbf78bd223dae
z78875444265e77e8100b5a7a7050fa7e7a5dd74fb08a249c1d4f53c1e2510faa0b81dc830a3185
z15fdfb2ac213bdcc48275f741de2e09e440f89a4c957d314826b2a139f23d8650a902b7a176231
zc3490ec05c8cf606ec397042f4b1b0fc764a44366084cf29885c8b993dc45930bc187a78e01dbf
z1e9c7926c639a99f5fef9531ace62fb6989291436428c95f71cb3cf02dbd4b9b2801129211cd71
z7e93eab99c5ea78f847a22cdac8ba1b7fde93ce4e6b6ce7df46b73dee2899ef3f1c1c92aa80fa8
z32e99a72bef4640facc584e29bd62faf0e3c90c9ec7339669930f1e6d45c48d1089284f5e9cffd
z2f09a16655f8c85abe5993558e7aaee1e0e7f6138488f908b207cff9c9cc70dfc0049c62c00d61
z2f14731069ecd5a0fdc7b8a282ae3c06ea02995a5041a6e9a2c3fb4d73fd55925c80747120177d
zc006cbeae443037eb3a458b2f4200c695b5c2a80922c7263793f10bab0dce972c69270f73669d8
zc2ee46a4573759c169b48bccc72af8d91c4aabe7674e6187c5780ce4dd6f7a9401e3d9389fdbc3
z2dbc2865aac7ec2dd33a211c5f74eea65fcd6288f6f2727a936db6589bc7932b3b44187ba6d7bf
zdcc253de89e544fb76898f4cf254da4c8aba42617135f6664c7d5b27e5e588a80e7e8fd30961dd
zf5c38384ff089edde27341933bacb5c61b1a46d7e9bffee0f1f8a3d96a87ff4ba088eb46d4b3d1
z63849d90b20e59551063828d643b6d1efd448c0f9b93201963fa39065d3e0772b52c09d9565cd2
za84777e8d53d9cd784022df0d164e6d0531c71151483077461ba0fb057a3353e952fbbc9ebc21c
zcc618fa883ea88d1b6cc282c4b60d1f7fdd566f8c6ccfe0b4c11dc744bfcb19e26dd27558c79da
z3dbd37c59b1a93a5358a027e3d23053ecf2703a6b0c1b89fe100e10298d4751bd7f0a11bc866a4
zab351293cec3cf08778d3f8b26cca1b5d7f90b8330a5497777e5a4503de72a6f38482ebf9643a8
z5bd3beb7474dcc08a22ed0cc6552e69c34aea0666e0e7942d7840990a41ad821a4eb40c7d15516
z5a4b3ac9e004c212e2750e0b908a8e1c1a892fdbc8bbd3212438dd19139132c4901e7f69a7b1e7
z985b030898c86d239d3d6c38227c10686d5b864ff20bca88d4b1decbe232cd9fcb94d452df748a
zc75974bcb351b400a7242bd49378a966070feee6761f797d2f2592bb01bc10c36b99d55b482a66
z2858e1a82c3b8072a9dd7bbc9002ce0dda51ab19953e5fd8a459c0d96fd357f4452f5609ea998b
ze80ef75d5ed730e184cd8270c43e228292ae10af3821f2c6f3d817a9255d62962c652dbc798666
za3363256a0847baba097fe18d34c77bd9014138c732d97bdec46734380a2abe385df503b343756
zda0aecb9611b0ac718d44991211e12043168e37288483e60d2fcffca1eee2b4200b482a2601251
z406295e8a44b1324fc894dbb96fb3fbfe2ca7d9ede9429510c62b53f3b96f38b9c5458302c49ca
z635f44da827b6913a5a5418445e8162c412be6a6b2536b5952fa94fd945195e6c03824a0963714
z4eacf265798a9b0b8123030ff1fec29d9a366a326354f709c0d6b45331daf87ff7c56af7641311
z15f8a16a09e507d1bc5209790842b20fbc5bbf7d561a629074d93b481e83ffd558dce15375f399
z8f93f6a6ae905c7eaaeeb0959508e2ca3dfdbce8e1d4079dc24badbfa90c32abcbc8db28672d41
za68d6289fb01f098a5cdf764fb50c446c3c6a5861caa674c4c7e611c48dcc2a8609fed26c71b47
z256a2567e278aef833d64b8970e9eb65f9194b17d6abaef3be4ec1b2ed4ca3324dd2fe68ca94de
zc6f09098a957ae280264a5fa5c04d10f47ff6c9c33b3d12cb06bac445db0789627d1736c13c7a2
zea6e4324b8ed18d65514debeb50aa7d0679f4dcf8dbaf8db659b8396893aa37a607c9235592033
z61a19e253b91ba029d153fcb7f0cd8c870f1414355ef5dbd85476b832b09c2a3c6fde617fa201a
z48a8577715e3df665172ae2506d0b630884261a9608d5765d23cd7bf62ef418c47c861e491fab4
z0bd651753537d2f112b8cbcf16f5fabf23f15a0b015d7eab874ba2c01eb68145df00868dbc8825
zcdaa2b08f5b79672088d398ecd915775dbdac893c3fe2ddbbd4bccf3d511e97e7d6e93603f7c2a
z74d18eee7bc594793764384e7c1ef07102d2fa7f8f859f1dcac669cdc26ffb7d7eb91985960685
zf32b15199babd90103ccfde300326b57c81ffc91809729b7f5707c03f4e74bd4932f71ef9b33c0
z16d72afaa758cc9617e4064ef37229ef5e2c7ef92f051bdfa27c689863481022e4a73dcb649cab
zacacb352d25387d9c02bbf241690a761bfce3d29622265b1e4ff345061a7abacbe3d6ffaf21eb0
z44aad8085fdacf06d87c84b3d2d93b38890cc92d45563df4e4407aa1556a7e0f8b1583f3e73870
z8305aef5530a12ced3cdbc60bfb633a6613bfd566519732b5083e41ae82c7674fba9ebc9132d6f
z8b5a41282bc917aa4ba3e3243b3503ae4a1e73aae4b0f63f9c976471fc024aad79bb066817e7f2
z5650d042a7007aa144c57bb1f849c90aa6e892e858cccf02d608965c4cdcd99bf94a94d4418f6e
z05c6219f3bcba9813263ce7586bd1deb6ed31cf874b19d1e129769887a483c1ef970c8375ed487
zb388b741c891fdd5b6fecaedbbe0cc80a3ee83f034b5451c6c2034b4c7e5e7c51d9c7d427bcf25
z13bbf06d15812232087fc23e0cc2ff8175c376177a3098c565a583ddcf87bddc533bc940164719
zbec9d69e03affb3dd515d9b6088f13c01c2999c9329a9cbddaef2e3ea3209eb94ffe5010dcced0
za8585d94049966635b05d01b4e4021b1f90a751b998bbf0a793a010cc26966797d8096ab6ceb81
z55c3b93f0c54eeaebeb2056f98eab9de757febabee855e6463578379c3d6892f3485a4906b87e5
zd17c6532533de3ea9765f599cbaed815c247e050518ca174e1dd207c608d01436ba7799445602b
za843eb6d4510f682ee8442ea305192729473a4eb8bee0512328f2c66d634b8a4afefba201c367a
zd3c52c11cc996ccc21311472380a1e53a9e22e511608183fdf3a5e190055a0972f37d56dcebb5f
z5bb255467ed3be1ca85d309e418347fb29e8e7230792cde70baee986ae5ecec9c100350b3ea6c1
z2c6882bd3e55cb70f7e69faac7f06625e0daf7c24b71fe9113648c02f89749e2ad39d6d2798f1e
zfb28d52604809249c84a0ab7b8168efd2c79f47f0a7447a1ea89293643693c3593c07a0b4f3362
zd6a83e848935ac550659fbdcf1438a2946bdc5411e49a816b3569a62384860234c7ad64257ffff
zbca9629885654aeabf949c7848d29401de330ecb60f52f86d51e32ea573926f28f1ac713f1778b
za39a90b7e7cbed5c084ce3a9ede24dec0bff6258e6110a88c808ac55583dc57af24095aaa8dee8
z2f86ce4d15424d75bcf549a28bbe89716795263a31bfd13516322395c664d8e053fbc67fd3e1e8
z658f24aad94889be31934909f23c09e6af2e4c475c3a64dd451825f6ac4106a3d7712fee1987d8
z1e5b63ec3e9cffcf60f517ca3e81bc1b11263bf3dd094942fe7793149290865a6941799b1a54e9
z359637f124f440628a0fedf73ea7e9d265b86bac5a5d6c52c7ef6a27a4462ae572d946d0af27a7
z948619e2ba3ff04adfc2a58902476ddab01d966c7378c154289d072ec51b299bba12b445866542
z7555432a4b8276869dab7f88960a42d221b3de21fc0e3c850ef69a04ea1e388eb3c335aa3b8870
z064e1607721f23613c0fb36ddbd03cae447dff3c76f1848c06fb313a7d5f83ce888fc3ec9bd646
z7c5067c445f40f1f3e6f468562fe20783aa6bb8ce2e0c33faca55fc4df551d868c5cf6c2349b09
zce25903282b68f48fad9947b9e239e4cb87691ffedf2b42029940f69346d02b6b7af1c74109f58
z26333911cfec3d4ade2b4a56055e2e739f3605b657e02797e972c180bc87a97c1ffcb182eb63c6
z0e2e20ff9009936a232a8ce731a55694e9ace73cb1f5cc858d8dd5f7cfa075bae70f18d609f1d8
zacf4798326d114c2f53fd6b7a21b4afa7ae7fc780281805a0b42eea67a661e0da02b62ef3542cc
z05d04173cfb8c642c3533d4781e04bafcf599c9ac83659021bf53fa8db4815c601cb161ebc00bb
zf726978f54d3e4d5b453b210d614555dfee7aa797dd167b3721c463208622f655b3d0b54b6bd3f
z76b2780474887b15dff858ebbea4962016e363d6f49ac18483ed2c268708d1a0d247df6966de37
zf1a9983dfedf500e8785b484a4fa8573cbc5ba96418aeaf252b9bffbd8438dfd63a8b4e94d7716
z1127b2f11e4d4f1ca4fccfb0ce9b72b930df993242aa4c39262e4f98866657fc6a993a4201d0a0
zb4713221fef58adba646ac8dbefc7d08b80e5099097e7db725e3802a6c33d64a97ece73f031275
z6bb88e2ad04b097c8b5e030042993e38c7228a5ed399a462781fbd9996e7870c2f6dd0eafef1aa
z865b486d58b1a0cb30396d9786702d46565848eb5a5ed2cd45e95e1a06f7766b7701b15a9a09a0
zc222365edd183b1e1e5addc2427834ef7b4b4b094cb702bfcd1b5e4bd813a0ea43e8c8dbb8df5b
z0d1b6b68aa74f44b3061315b879115e1920f87c9d94deaea66c91616761dbcc534495e6a43e6ac
z6fd6f690d8c0cdbffbfb516f4a39580bd1d64836294f04bea1ff2e96d8a6c6e227b7536414bedb
z7e6c46055255755679e8a7579dff8a1ad78444b0a3e09a2b2f66dab0dd8a80fbc16780f8caf9de
z6508c8cd47271d831585c055c8e8fc60c8d09dfb1e5234edcf6280cf33f75df00f08d1ad9d9863
z1eb936377e4067eb6e7416a96fb5d79dbd16e7e198d3008c6bf82121d485b4634094c455cc4190
zdea131f5ad65359c7eb0158091196e72ac5f345b0483f1af285f78ba74f9671458bba6fcc0552e
z73975b9a30efe8f1d995bb8a85832576f1055d4ebbe0745214603e20aeccf73ded22d7471a5bd0
zda339d89c6a5a4cb99d69fce3ccd6377b84d74698752041ed7ecd535c7a841dc123c9794c3a028
z74f991de0a8b91b8974a61d3b7a7a933cdb299f15a5f71c22d4520e0c3e5b54c347259094af35d
zf737cb20e4abf02c36341eb009e40b52a1aec2f223356f071b33194af710b06ec26c089b085505
z12b6918f0aa966505ae751316598f897e44e3fc9ce1d8dc048261f65db5efc6af80ec9180030ef
z2f2d1db00c409a2bc68dae3779a8ecbf70a9025655c514501e7ead5d2a76dbac7a7ab33dee0e56
zc9b5401ee9a6d462b3841a77742ef00d2a3986076b99d046691ba1f811c2a881098ece161c29df
zd7d875096a108afa2ea441f0e278486c50359c688f250cb839c2937d1f6a8b386c970afbefb3e2
z68375aef572642e500b0f1a85b31b7e892ac44ffb1255f9ec20a720c081148a9d604e4313f7156
z38518ce930b14386a5214955ebbf2add8e67aae6c989241136f642c29058780f21f86b6436fad0
z9c93f0ad97b337c3ab649c7c926b927cba8ad0efe4e0313783e3d2a29fe4001adfaba10902e180
z72d44f4466a0c16827b61aa28111156c5d5c0fa4a4a13a5cccf4f096eea297f1399b073031d22d
zd064a66d4f2e8c00db340c1a54b31321fd1e90d94528b248aa27adf56be5034d5967262734d77a
zf3ef31ea175582ab4b71d5bc5b6cc87c7df580a66953d2a1cdb1636412aed0dc0b4c1bd1caef35
z17530102e271764afa56927d46b83135cfda4a03c8f50c6b88063cc673b7faae1d6e0c8c658bb5
z3a18a98586f1217a95841e9ccc93c5285382979630e70c29d80556b31f84a69646ddfee6da1512
zb9aaf53d1b36dca8c58bfd48e9d5aa8957757001085f1977a7edcdbe2e7225bbc2b0ca6b2fcd8a
zaa9434a23396db0403f14cea5a73875cf391460d11a6c9e27a5b701cf9444b3222af049cf7e0b5
zf8456e5a6340aa72d6f4a93e3638f58e414fc4db53fe648bcf283bd22111efb19a74d211f0ff84
zd59d65b063402274f740ecc7e6edf49a241c913f7c5258d7be3e960c36524c4a1eac10ad7fe0b2
z3fadbe0dc8bb093ba74c0929c82a4ffc2a9cdc6bde8ce18b5c91ca0ad7d1bbc5d1341c8e8befe1
z512f774fe202aca74d1d258a48a2aebca1e18706b22bb5b75454a97d4f038f75da3480a05c026f
zbcc54a5dc8b7a758e62b36aaf6e4836e61e965def49ce92f8083e949b494097da83273cf6733e2
z7f01ff8ef27c575992f5661e46c2c2362d8dcb955a08b2b2ccd940484bd040c8793271ffd64638
z5d3c1136da0d25ac8cbf8ec1c2ca6d673c8273d9111e10a11a911d8c0c557e2e742ebd9950f99e
zeb975102f3d3a3e3e97452384a5bda7aa24eb679308e35868451bf44e99b99fcfafa2f0f87be51
zde38934604a9b22550a8cbc2c91fc112379f316d3cbb1acc0305bc30fc700fd8384872425278ce
zaf02d41ce8ed098435b71b87e3d3fcac4381ac17770f586d245ff0295bf50a6b753d653f662dbe
z6bf40fe4d3a0c14e538422cc058754889e5049ecc455425200a69b558d5030544f4a8845d27250
z5d9c176156fc3a5662c23710c645fab7a4ccc6f376154921313506b7d3c0e509f5a6673f4b35d6
zd33f4a2c88afc1ba43c2168b70e092ead5f81c20ece39323c2395b25cbce430415f07ffd307590
z0c52221a0f80b9a75e17be27be139b776d63e5ef44a214c5873851b35ee44175afb3e31f4d7b52
zf7e909a87e1dc3b39a000265550b62b2536ad3e70078d7a914a4a94844e1e0fbdf0bcb0eef74d6
zae02a75d5a7bdb3e74a6f067a0642aac3b2cf622cc065e74bb52458967a659666adf7d06c0f004
ze402733cb90f710a267fb6081be8c498f500a15f142709b8e9242431939c797639bf0f928b8491
z5789cf5246b77dcf69e82bcf1b2cdd0ecc5421db47f82c7577041f57081a471593735ba41aee4e
za85d07540043a9890a91c080a2c07c7e84239db054cd098d5942fcf7bca1d1abe7d935feb95c16
z28fa91a8e884f9e6c417b85694b7dcf1b709675f687f98f954e2111f0939db7e093c2cdb434a23
z03d0268d8e9b0f754019f52fbdd44931a64794a5f316d2b07f18429ac38d020f183884a637f527
z5662e09aad21c8221d1b04508795354028ee549c565c13b94daf1f2d3cb19dc720bdde0670b07c
z19325abc60bfb915a4ed925977321161cb97fa84b91e52fe4038dd8bc5322c6d1a7f02e960704e
z961fa99b6ecd484856d7f9ac82855cd0bcbd5bc432c2c71b0a9acbd16636a97ee475df2a4cc523
z032442f687b59f39fdde10fe344e0861ae55a08d99aab5c494e1612c94aed9e6b224f6a1cf4bb8
z4d7178d438f7bdbf1af7f7538b0ba614c53a892f1d142a45b77be7f933b469c7acd2f5c9134661
ze25ef175ce8ee046553e2fbe4df40ccb9287323b7bac114095902c086a76e187e15f13b2d910c1
zbfdf0c5946e1949bc3787b4e576fc0df9d8aee04a04b2a6675fcad7484ab0f3003dc425f1f11b2
ze49f471dbf02fe30d8aade1c9b6efe469d033a3922f155fe54eef5ee9b4808723a231c0367e832
z3bc57d107080d5eb8ae790ee4487ba9cae8f5bf402f743e055beff1a8b08beb016ae5d2ceace93
z560f5be1f15ebfb8d11504dfcfd28f9477df8204aa1ec818221eae5f0bc384134f49a1c51eaffa
zbf2207a32844a59f816d26bc231338cddca9c2c0cdffcf877b26f689b3714263a1859babb1dc86
z716ef5095026f1d567084fd0c94a7f2332a34804902011bbc7fe26e485e64f9ac5eaa1035bad00
z5c94c4f1df3428b4dd8ee8a324b5ccbe2d8a2ab3ae71a26ddd76e51d3cb4a1f2f76484ab86c14e
z41b833f1c417943c7d72bf52224ecc530612214f2ef8be21cba2fd35aafe570a9f019733e86d88
z35812a6ea76a987da29470743851c133185b2691a085e61e3f029f9aa0e5a1b6ea112d838bfd90
z1c724e7fc16c3c46877916ff63de30e7e9a764ad46d92a4899eef394aa257fc16ac8258fc5f4d1
zf216ccdd9be8be15aa7a990b981212eecc67befaff7006d877b9d1481e0a975b818fd852237c01
zb0946a8b671d73f0d19a6864612429b1adad39d429b894626c94a089d996aecf507bfda586112a
z655009a30d3ac36e2f9c07b2b58491e48aacd890ef25b049d3cfec666b65911d355506b89b1541
zbd437abceb60271c0636c227165b40bcf1714f2f1c8eaaa5bd761cef22c251e10be5bc6b519413
z94a36fdf2d17c6b643c187606c9bd7012288986cbceec8c65b0ae4fe4b16861d1d50497a19dde8
z9bf15efeae5551f399be4b150af00cdda67d642b70ea385b21555981d99826a1ae220f7a6b790b
zee11527b2bf09d73a7cd8def44ee712bc0daf1b0e72989a0573cb7ebafaee57016598d4bb72134
za046570ae37ea803c3a9479b3e5f96330dcb0a038e9afb2c4737b3c64be82192c35591189c628a
z63d82d7d2de8fc078a9624c255f6460682d5cbd9ec90e8d0c971bf19e7f399a5abaa552da4a0d0
ze24ba3d69b86da2048173a776eb34f84858027d92411e076763ab5773d6880ae5d4556b8800a14
z7c4124febd6390a8efa081427ddbf8f99305ebdd222fee486b2f88c75acfe703486a121471a03d
zc3e1d5607dbfd9de3384f5afd04335d98d26b33279c89b74a12449f09d05870d8dccdd697f356d
zb0089dea99dbce550772741bbf412f7aea540909910bfac28dfd784209b6952ad5f55a7c9af351
z5195c4fce6153ad8fa268f6b623a2d7649c9524683ae67356fba2c1ebaa4c82f409d1038e17e6a
zeef52f6b15c97e29268b0309e12750f506f21d40bf56950150be790f347c6a9ab94cb616a92a7e
z1adb4b90be9ee0a4bd113f54694a383d182389e9d9361f0e4d5234d3eb1e2de17a224924b42633
ze80010635770f686c67d29d85b78f7953c213cd2a5539578d2889cd722dbaf27abd29b72fe3740
z836fbada025f4847dac7e9129ecda9852ad28b2024bc82dfee51ac1eeaaa0e8d55c31f84dca110
z6d289bc5eb9c1809d4478375a70164993ee0219b786c594ed50d65331ee1241dc4a22f352969a7
z0b4f0467fd9505a4be213fa8ea10acbb09d70d16231b1faf1229675247b9744e4f592ab23fa6ea
z1d2b7c8c1705812366e43e402f07f28e31ab46a510a374a10c32b525c8e0bc19100c76eb5dc973
z9035a0aebc79fcaa76958aa446bcbf1b6b4e2b316eb95e0df20674d6039158474edb17ba1b72c6
z2a7ad77bb5ee2e91c6a72228d6d5dd8aaa79f3958df45bb1ec933e49c3664963316d6c091fa233
z04705c76115815b4548c7080fa6895e9202a7986789bcad4f49f471aca20b00d9321d4942d27f9
z9eaf99f2fed513977f2c73f72906281dfa07d7fb196e43790ce7e039582733740f2fb48bb615c7
z1c4d40bde98e9f747a5b7ebaa489d3861d43045ec05d86b7bdcac4a370fce232f9d7d80602e1ca
z4dc98aca9de367dbbcc03154cab2c62fbaa7308b068bef374876c7b4f99fab4ea1da28753e1459
z8878c8b58c4276acc2507214460a48f6af7503e155ce9d9c3579d930bea315e6bf03807ca496d9
zda23cd928cad9f5261669994d3d03e92eee562963883c859a32478531da14bb6a5cacf52f157dd
z85ea5927b46d9f6b9e5d4918bd8aa15b8eef8075f5393ad442506976c1266872c7a06a3da56718
zbeef3c1075affe4f2aea6324ec5136084adb808082f17743c1a17e06838d4539e2b4c587fbc9b5
z2d1b5265e7bf6e2af7f293c7725558cea5a2e4c7966855f5db2babd3da6a9ad616920b64dda2b0
z54b5c94a5795cbcd0752b92f8d8c6e95e945eac41281bf393b70ac4ac431c039ecb308cc5bee37
z26e42ea8b0f14ccf8c4a33ace96d692281d227d75f5da85a4ebb343fd6fe1bee0c035717c45b28
z3247589c14b3da078b8a60a598fcd11a2bca34864352e47940128560bf3214a35597c129e090d1
z62a033861205cd8c4f56847f4dc0ae9963644da1c5399580b3429eb7d5dc681aabade726ed0723
z63d7e22fbcb1b45156a163431dd6b2b7689a547a35f98a0be8091c1f56089ac1a62b78e5bc64b9
z0854370e61a79c1b1380f79033446331237965e45b4bf1d429a81e0f9b69681f0691c43c9541d9
z6af7b369bf6b9e509f4d9a6b33e454e3d9faf991b3dbe1d03faff907cb109f5c35200d0256e0ab
z709a9971cb2c7ff52154ae0fbbe951655c7b28a44795cbdf0fce9ec776997b952226510a0fa15d
z9ecb091e217829937ccba9422da60e4e32ef9f640e9b65f73a95a34b08c3db7aff2dd8c49e330d
zf8e2c3b755a4917bc1648e352ebf62b6900b8e4b1ee14640b994cb4cb18397bd2474621a509f32
z7baf75c66c387f00855c083ace46e0c3409e6bf1fd18fbb67d6ebaf4292a5056399b6f20af3b7e
z009a530b89f5f88629cfee4889c692d0dd51efe9833f195a58978eb65435baf68563e297fe91b1
z37bc8bfd28fbe0170234b80b3e2f971ce6fd8e0b71a65a2ee8200944a01e3464b97d878078e2b3
z27004c15fe5e2330fcc290abd7adecb28f7e57568d2f267c2e4c2129709c0671b57c26f9f64c6e
za87f6f0a043318980fa983226f4aacb3bb95274961b772936ed325025ff6ce2d1ee0851dff1a47
z3c5fe3a3fa63ecba764a7161388ac1f4d138947fb158ac872e28d88bc0b4fd9131ac2a9ab3b3c4
z1702ffa8c1c821f7fce711625415e21a08ac2617d9801fe6bea0700933bf859d86e951dba208b6
zc6594801ceb6002fe1dfbd5c4e93571990c7a9680e88ba5f33b35f0d4ac71209cf3a4f0bb2e89c
z971fbb3527c22b438f309f0ae8c754403fd16be81ceed39d5a5195372da24bbbcf0b6c30f691a1
ze45eccebf7c020a27c12c63a67ed4ce8931971b1a3a2d8c05f5b654d0a6caf727003057af55931
za8a83bf98d6cfedd8d984d158399a755b325f38d0915e7e1411f51b68b9c4a25360bd9d2744da9
z42f25c6bebfe45b92a7012b7d1297e31c472366fe665349827ea68d86f151e0a509e35fdf849c4
z0a4a068ebd36bb30b8a17731b565ea41d444fe41e11fbcb6337dc0dbeefc83342246373d97c8e2
z5d9fefe6bae3e6dd064c833ddc20052b69439f426712f9f4fbfb32c4229ee0640c07175bd6df58
z488207d5a2ca46ecdf392ff61fefbd75cb328b368541e109faf8a3cfba654c6df5f29e4448429c
z860bfa6c4db27b7e22f1dbeaac253bf74a6bdcfd3b2792ab2331f5f4a8bfb3082c5df98998f2bc
z0c93208f0f41c47833caf8d05f52b5759aa668ff6cae8e7cf97f2c87798b335c0c92d930bfa1e6
z23f41b1d604ecf8799f36b3ecf3ae3bde73b2c00ff57b1ac54e3ed7dea710a9d497169df1e53de
zd6aa814f9957e9f80aaebdea712ba53ae41bd14e13e23f4ca7172d3f1e1d37fffc9ddf207f6ede
z4cac14c39b32fd735dda04b2dd48c50b3f250b4fa34de8d1dad9ed602a7ee54acb78a88e48e365
z155850874a220d0ffbcaa0b3afb1b757be95d892fc2f2343d2403a28ace23694eaa2d181885fef
zfbb701f3963a0d73bca769f889d12c7f3f282566b81b44cf86cb2fdb7f221b0d12d5b3f5a04e02
z071bb1df261d9d54aff95d5cec996d60c7e15b70c72b1ea1809e6c87c5c7e4085a09622ded2b24
zbe491c0f1f46519418f72db9b0d2f0a5bc59c9e65238b9c7f17f8947deb6360b44203b5af734b9
z8f542a570cd2806d446a36f84dbe7db48b8ce2d50d6546705f0014098256d8d180dee93de87e8e
zf168c3e78b7bf5414fd26a5200629ba2864354818c2a0b34d695b47fd8d410006082fd39aed9af
z4419e97ccac50e4d35b1e4e349ca2a1677331cc3a50247be3d5ac43f75a1e03b3cca83b3ff84cb
z23f0eb87031a662f9756aac6a1d993ddded6caef091e4498ff635ab2d665b0672ed0a93f014542
zd0519f69238a153191a1a5b20bec11600435890f261522fc654572e975f278a50b22fcf4fe3a68
z9e71d67a855f3b8a172e71fa593786732158c24667ff8b789ba10221d84dbfb4172b24d057abb1
zfca2186d3ab451ce55698a4f9622dd34ba61ce82e7bd906d9c7a42ec65d818cfef97f47ead5fd1
za3019583a397cdb47ceb758ac2be7437b59d8850f037844403f2228c16a949df813b5e429d9677
z101cf4ad1f5c23f2abcaa9400e1ff780a46279863bb13b18a0a3fce669ff827aa89b18fc6d652c
z3aa2f397d16949b770834dc4b381a139a816610b7f95a72fbfca4752b6a50ac72aece3cd665480
z546bdcef4b8f632067adfd7e727544d02324e13a50071ade4a1ae20ade993e4dc3b8aa6728cfce
z6681aa5e3b89ff2b653ac5f34ae30c43a30f377a99de4d5f8db51c31ab1f15268b301507afe3b0
z3bbc5bd69a46b837a9c8613dc5ff54ba5f9b4cb95c2b8e5706e9552a9d6816e4bfb6780e75fb1b
z6fd29435aa46132302461a1a65c508c73e330cedf33d9da8735b5a0ef99a97258a085895698ecb
z7063d19e0a9c8b35fa61d9e2d71e487ec07cca69ce28e6d2d7baf115a44eee717519a856c3fba7
z481db6b4bcc026e1fccd110e363237f9fbabdf65c76160cd7c9f2251d1d1f18a86b61ca9f3d17e
z172f5cc4ac5850647d96fe18923c6efe28f54db41960098797dc8090059ef99ad09081811383a4
z1ae2c01a4c7530f85495d047018b337286eeaabd6ea02f230fac82f4b8792c8353efb6df16f5d5
z7cd6e7fe75cc41641bb304939dcb9c4d45b1e6258655709b4e9d329ff56565daddeea43f0b68fd
z31897255ab107fba485f8a9820423739e199ff07364c8875c4b63462abc7364118a5128a3b0589
z528de9dacb4098249f585cd9351779140c1f8523075e086264ab468b3e8442c1958e70323c59d2
z819202e982de057233532fe86bd1bf771c1bc6b1c33676261621e76bff7a06975008cee19e499d
z929775e472bb657994043eb7792a9f7a1dab8015727236fa45b335087d6a9cbe5ae88d25a93ef4
ze9e249b9d51f5d5a408ff7e4895d7d29132e2deb43f876761fbf6ffc6381ef411767c407d913be
z2aeac8f5a1b7934f19a424200ef259e27127443cc5da5077bc4a1ca1246c75ee18699f74a27cb7
z91ec958cce13d76107aca03ccef168513cc382d2e38894892618675ba84f85be4ce1666700e145
za2a72d77c099a5feb660dcfc4c372d026f04ddfbd79e9d52056ae20245c0560bcf78614394bd18
z80cae9244c3ec2b7e8f9d8c2f1856d69cae8f9d1da5b05acba3684e9d160b204166e3ace118ed6
zff283a62eb5f3cad472c773b8295bec358ec00c2b3d6e902f4568f9b87e3cec640adce7be7ea96
zc08d85cf838f1d7ca0a1934984da03f56ec7b0257da886cd9d212d16d26b7b42083b022520825d
z21bbb130bf98d84ad7b64b46ffd409798f274129f35432f38556d42d9c3a15dd51cc2b99b0946f
z8cc59617f5bff20933314197d0729e321144dd08d7acc6c246bd2361fade3822506f87fe0d1155
zb8ecc01a9c2b02578b75c1be4d792705626187721c1023ad189dd1233f8ce038207e0a51e9534d
ze1d0dac9afd22f60193aa83a81d0c7e483e4adce8348dce4298b83b956ed4835e90e371bdd41ef
z85322dcb6205bf7182a64d17e7a1e9385767d1b321136d33d64576bf78a3395bf33697b4ef4095
zcaad6937b7870c4b02cab3c2a93eca00e22556229252c3098594b4e9ec11eeeafa31c3ea2c423c
zb2c7bb8bcef10c8a22a7d5aa5cf999982c7c91fabf8eaa80558e986d986e7528f3c2b2ff59c750
z70f33c8b1708c240ca9fce8ede52692dfdc9b680ab0e07513658cd80398b9cecc459685cf130a0
z10149e76e2b7caff712f71c3909d0a25810998eac67848237ca8f00343fa6301dab5d8341c15bb
zca1ee597e50f9223c654c51b12629f541ab018a4fec0a2dab6e305f3a22d16ecfadef6448a3b96
zd016b27f896150e335e7fe598aa669ace622853dbc524cbc23d9268627a88b24a75d1967d169ef
z0a219052db8813145b5cea3679a388f4dff6dce6ac641c7a6c10b8cc0592da5fa9433c824f1a5a
zec75a80ae70ad4e1f89f9cae3a8195b716198e27b63de96579b406e5aed7ed740e131d1324af42
z1b0703e7b87b411450261c1ed462fa1d8d1e37a5b734bd783d20f8217ef941bba46ac3076cd0dd
za67f569e5da1d1e835836a0f0b4b51880fca87284947651cc81f01e2f47896f299790ea9943bd5
z0d116e22e1d5434633fbe7e04ce6be196b61756eb5aa9e56bfbe1182570c3414f9c5d040d91fcd
zd73bceba47b986ee8d397aac68fa8187f3248462022a2d81142170074883d96257d34a2dce8285
za5ac05ee1a049179a6f6cc7c5644b089d914b8357488152b6ab7b4bc3490a84a88e12b516b3720
zd6731c087b6c46ab974462cfa5b869111902c0d5f262e716c23c073f5f3e5c80bd03245b233c96
zd6e149e766314fc6d4096763468220caf7be7604216dd52750e4a5ac1b3d484a06a26fade54bb0
z724adb1f57b7f9cd37a74e37bdacb7fe84445ff664cb669dd1dc82394f0963b90a57883e43d64f
zf8e5d477e7379596ee03b2f44ceb1c579e073881afdaaf45513109b86afb84b795b5d161699997
za1dcbc897f826aecd011fa75b2e9a8f2889de9b5780832bec060226bf8e8a544c00564835d2a38
z728590a40600bb80827c2d1d30c0815e139387210a64a343f99db315910822c6f07a8ee29060f7
zc7cf4652444602113c83d7071e2f166bd822aeb823b0e52b482a5599e8041ecc579790fe1a7621
zf4b3ccd51546dd292afbaa009d19f453839373bf5c7778f31e30d9e65f6ceb183822b78d83801d
zbd1c486b032ca0a5868620281138e63c2324ef294a84fb4a1a5e24c1cca0735eb1ef94ab8079c4
zfd6c935f36964ff0fe535dbbf5ea4f8c0ae0f84c99eeeacc4db49275d71e45b12595a32fa41157
z32be85222a50a432cb88c027ffdad3c5bd60bb95f4763a811fd0e8517081d2d5c4c7fee54ef39c
z574caba30b90045b8e751e0d49dc19a294e8353c26fe8f768a8d8522e06f0552712c1f50cad1b7
zce2ca2521cec367338a02d7a9177d31962fe0be433bcbb54792b2de84e83bcb056dc46ebd4d8a9
z070ec1915c0ba6a435cda5d23aaa7f936ea87e9a63ac8a428267b565890b8de384bb27cc1ad1d3
z6a56ff6438b9d973d9bf337200b7566998cbcb2144de87ad06ed139b584f495d9d9828fc275128
z501ec297b7ab198608f446fe1f20c5533947b55a5d3b4080abf45d673104930a2d3db56c168db8
z42bba441da539487f2e243713bd268d77624627063c21dcc022807944af4eabbe103f1a5e4e678
ze120433dc891b35e3155b7392cac816a7bb061675c439ef6ee8f3ef5e140a695d3a252cf8ca335
zb3040ca92fdea0e453bab2205a9b7e6fbf900f7f441d6829babfd1e0e66593af5d256d9d844187
z1cd4393cfc87de6c790e7eceb5fa2cc4ef95fe6eea22a5b3b26ea28f559498bc03799602f917f7
z358fa54a1513efa734cddafd0223d0884c456280d1cb0c8bfc0b4f6f2e866a32bf555981fe33ca
ze37df96d252e3c43b139b94cad457de078a9dfe6cf2973010f6d7ef3534e0565274d89ca147597
z8a0c90b03ca6d1538b1a67bf4e0c01dbe000bfea35a98a1cbc9caac282d7ed31b3fb042791b09c
ze71948a0124bb82bc6269b06789df8690c65bff11732158cadd6fbf42683999c83205e11a5165d
zc62cafbd123c42c6999cfccda74cfae23066690f34ae99a47089bba8d953b6c3837fe74ec47562
z59b04a8a90359ae195a456dd72e9e6f4bd6ca347526c3b90cd9d8c0e9b5e34dd77928469f2e60f
zf4eb5b1591d8aa00cbc5ecd2bb9aa60f7ce5bcb4f8612fb7e25f3de5a968ec90639029c3b278ac
za8201507e2a6f907f736f368266d4755b36c1c5fdc298669423bbfd1cf3586e3b310b8cae2123e
z1e5ee9a36ea42a9fb6da0f809cb8710cb000f0b75fd37779877e4186c6df7cb81179d150798ce6
za8aa63e6ba3f8a5c4f1a3464a34a66898bbe9db7bc61b2ee1b5906815cb0edf8606adc75bf7f72
zf222adc93dfc3aaff59e3d527f54c628b3f2c3caa2a24319d55e8725f5160e5f3d7d62188ad0a9
ze0455eb2a7e3d9ff378161d7a2f0de5c10a3b44a651cb006671d5b273e6a0986efd12674f69a32
zff410ae8596e68abf1b2bfc1a2a06475e14257610ee9b338e19b851a6d0705fbd51ee923463595
zd0812e828eb90f8fa3bac65a3ee5aea837d6bfdbba2ea3e35820c3ddf26e4a3b835a2e36478ec8
z5f57a20633b145461ffab4737398eb01b9c9e438bed2dc16cee3afca620a49b8f9d2287d708176
zdf4edf807be53cea596cf48291d36d9607f13c092f38b80301350bfd0b597bd3f99a9f8b3c9449
z894fbad4e38b20150fcab8e74f9718da92761bc93657eb6f81cb04300e5e3132553c4368e48981
z0aaec44ed89ea59aa391a9e146a01358f91282e944087a7e71c3ade6f13e270d66c445449aa688
z52f22314f8466a32a36c43b12da1a237ea792be48991229a68626a57ca52e971ee506ea626a34f
z9f03f20e9e4e4330fd518bd19561459077901dc50757c145a5646c3b4b0d9528a05223803a4b7e
z395eaf10e2bc0b15dd65cfd69fa8d334531bb46c64e273c405307cbf33b57c692906ef44f5557a
zd9255a8f7d1232fc8af3009eca5e1b977800e5ffb2f2859716f373451662087865d6a7f68308dc
z4aeea1c421d23f5d91cddf587bfb09758b3151f27e9793465c5017209ed8ebe8ea2f495c1feccf
zac404564c2c4404e6362e7fb96bc64726d3e758c26e5c0bad3d6deda1603791fe01e8bb47ae61d
z97efe733ac07d53fa2738a763b09ef3fc4d47aef86f4b84b085a2705147059a26305a98310baef
zb3495dfab24b0f14efa3c41261eda522db2cbf31e0bb5d4c6f41a876284d9c051b8c6d3425a8bf
z9d82c0d692c9efc2d1b76a37d4656dac6be4b3a171a67c346c511b899928bcdc9ef7dc0e586855
z31b2c5a8a0f497c983e8a527691a3adce482e6e95f6c9107764d6f6fdce1d9ae8588d84feba4bb
zfe9e697ef195c0d1a81dd7a46a3e3b4c10f5ea963dbef5464ae51da832790d1177a231ca13d0b7
z90543aa7d0d976fd4a2c46cf8bd9d3b01d522074ea75bb9149771d2e2b758d544ab0663b0564eb
z12698052e91d8b10230dfd79ec36fc9647ace52f1a1bc93c78982e4a24cad87b65fcd128510b01
zd6885db9ef78d6568af9cbfbc87bcdabb6a4fb7689a6f03dfdcff03507a12c893f3538b5d56c8c
z5014ce107c9db7ee13991acc4241df7302fb77b285b3e2481c6b7fd875cc520244deee268c878b
z6434eaa2cd54a1fd80b5b7e909cdbb7c954f862e92de6ab1f1373b2efcd6ef810a69e714cf34e6
zc43ac0442df3ba8bf3e04fba1f41d6e0765daaa5dcbfc4d3bff6f631341c4886f382b463415e6e
z90aefb9562962392515ddfaf45204bb37767f7adf8c2a5fa108f9a3e6468e968f8bd5fbbd7ab1b
ze77a431fbae6420816f626e4798fe3580b2c98b2310a3ab2b8c8e7302cd3e5a24aa2ec84010920
z381e1efd99c4cfaaa4287c224563033600b0a4c36122a4aa137be9a79fe54de6c2507bb56e1518
z54806c733d9f73d98734005aff466e1f54edc839a07cc431add8c3c6189054dac82e0c0a52fa9a
zcdc62207e13bb37790538cdaceaf0fee9080d461c233bf5604d5d94508818162d2c52d4d42257b
z666db141c9d54fbc22020d77041802087d61071935d4aa100d24b275e661b39ab853f5739a822b
zd45eaddab65b45bae06d74ef6900600bbc8485eac7b124bf30d1b96b947740d96a8a5ddf02babd
z9911846c5c3bc0e3f5ebd20682dcb6ae0cd7c7491e7cfefb128556f0a2e44475e9642597a16854
z6d617855b8e85cb83f4d02e8d286306808ce43473a5e71d8e699ab31d8a1ec4a09a0004425cbe2
z40b1b9417a67182aad4eed7b66f6c372584a74fb783d3d375a8ccca4d9d79781f4a684fe396bb1
zff7d4f3bb6e1b8fe81f3194123169e2bc51566efba200b4624d61efe9a3629bc6bd8169c36bdc2
ze5f2794d9129ea38ab38514808f627dc869f53d2969f0727f8193e9035f82acb3fabc81f2d955d
zb787136bac9c68504d98f86a399cc6ce21f62f216052f90fca6f88e1d1ac72136b963e299bbcbd
zefa6399f5f11f79e7e324827440b7b4422562ab0d40abf720992287719b7fcc0e0e159151dd957
z4c02b120507722951bb55bb601060ef93368327ba0c73a9d3f02069bf99a3bb009c27620fcf9c4
z7cb407bef40bdb5581f0b82b2af14ab8e6ed3334e2e960bd0423a65a0b38f33108d47c4fc7320c
z0827b08fc1a6cb7d9c99d57f61263dba6c9809ce95994aeb84f98529a07d4f4493b76f26a6ad28
za083e0dec9ab58cdccf797072821664af7a9d14b852224e0c90d50d7118df2fce8e5f3cdabcee3
z1f1c1eaf1d27a74a5e8943d0cfe240eacbda41aee09abb8712dc8f34b606fed301e9f544a8ce67
zce0ce18dd274aae6b538b38f643f95c9282ec38e5884b89c9898b1ae8facabf60058d3e0cd2bf0
zc1d62b4b40a374c6c5af57aa973db2ace972070833b37749b00825f20537b4061b3ba075ae80ec
zbbe9cf168e5942eb66649d326ba98c7986734cb038905e0281d402348cb774807cc449d9efc7ed
z673408c1d6b99703982d2edaa7b77a79b7a3b3798bfe5a361faee5698b1944d6f1067da71c179c
z017b635fb4956961f9cdbac7728b891067ef37f015784befed991ac89640aa0445d2051b274cde
z15c706f4b8643572b6948a3f45e35da6211dc41f4678d63db5bd2cc44466774fb11ec330ee8477
z3da381a739a79be6f00feff9766accc997a5b714ece9ebd9c2165a5af0603289cbf9b74db9bb64
z4c2abaf09907c8f214dddb84d94ed1d462c3abdb47854b6fc2928f50cc04d76a8cf847d47c51ab
z27d1c652e1af43852c3e7f6d6c09e98bf2055d476556d574cf2845ed8f3b8ca90b513315e38ab5
z52b5d4d14d8305f9973e2d065f0f00dd39ef8725744629cc840c8dbb8a5472f11fe96bdb917a01
z0ebad131cbf2998f7ab6070608994f021637c09fdfeb7b8c1f0d099892f95c89d1e6007924dde5
zb21c2d813c3beaca997e6dd48b2f8277b54b67c3f6928b01bf37fc1c8e9398c41b0b90a8ad10d2
zb1ff5f9689480219060bf1f66c1ce691892ed4aafcc614f1b7253a35b86c5126082c76caa55d2e
z3d6cbc1d52c62df4f5420a7819941ccac84721223955c831b24f05f8db068e1d2f4c6da1c2cc26
z9b733af6b3879fc4e78cd46ea6f73413018635059faa922a6b569d3d00d577b6476f42ea8e0818
z159204f7d80a42eb1009f030e2207150a4775ed86cfa5e01c0e25e674d2cdc2967912a2b44bd95
z2e6664691a984ab7fca38dd9cca35fe1ee116a3ed8f2afac88c094ea5dbf99acf5c1b5edca2034
zb7352db038d855d80e8c5f7323f7f921923c3750bfedae7e19a8e8aafaee9ffb7b8dd5b9388c57
z2abd13a91bd1c9b21b38a4e65a88e04cc7b2b2ca254c7596c8c187065f15fab882fd9a81d8f53a
z81d913ec2fd8537e01e994bbec1666127fe06de035f0b1ee66dc9caf6e6becddcf94f4b0143486
zbdb163b698ecc775980d24ea8cea0d9fc1fa54cbde853685334dec2ce8bcd6c679b5167ddc74e3
zd491f458b0174234327cbc8a8eccec17a7594bdecb66c24c1ec7c7d29563c17bf21462c5f4cae2
zfa1882810f91605e1fe53466dfb8eafe412670383ca93c97afc6b1774745c2760f5319d2fe4954
z17daf2e9e9ab4c8315f1834f7f326278e500ac37651708a5344683593f514c32cf2d0fc13d1fae
z2d56f496489d77f76e6e270adcbb7376ed557ad2a45f6d23380b698da44ba46325eab78dc0d58a
z7d33600387234be0661a546ac9000ef5be9d0b31bea6850d199a4f155f7e60bd436233655be10a
z593f345f46a5092134a18d939becedfac2fbb89afb20c9ee0a775a22c75ead677599a4ff7101fc
z35b0eb06a0d3fdd74e43f456f79c11abde154947e1c958b7c8e6cc9e0b1f0f1346d96860aa2b2a
zac34d885588ecf132ad2305515f7f349d15ed84e355709eaa7dfc774f9758070baee9e15c0f00c
za802cc2d9cd855a2ad444ccabae72be6fc9162b49f1b62bc6b9194cc26d186fa9615748335840e
z7499a7ab3c7103320fd97457e6d9cde544b530d9dc1f1a27fa4700e71a4baa7213e8b2f671f497
z1b40b7472c3de7cc5511b39dddfda4eb9aa3588bd0540e1efa22e3af22b32afadf77879a379bd2
z2fc816237f1a19e30ad25baad3ea37c7e2fc6b1bd6acd73b0d9c1537b588b282930b054ad2dff3
ze48c7ee459779aad9b16f6586b4e5eb9fc1c1e57203f2920d5df3016e52f5543b982b81e19d2fd
z91fce536f9dc868d2c6eb165d57ac6bb18cb931dcd1b4025c168fd5eed5c011a1555d6b8a109f4
zafec32c234d5fbe8548c9363af69c52b983042d14572dd4c59cce677a62fd5a3b153aff9dff5a8
zf90a59f2d5ca2fb1e381d0c7c6661abb4b4a1df7f1d00d31e63a4f365add582785c0a7ca8d50fb
z8fcc4caf849509aa9d3306afd4f5e14c4e80f419296ffb8b1202f1c2b6e8820f3b07f879807895
zb3b50160db871ff643e10b3471b2433c03296c4925c37137e1bb5115ccd0f68612ee3e7a4cd564
z693077681301e459c264926ed6e10d0badbf3f03a6c126e55f848cee3522aaf273343309e0702c
z41b5940d23c0ade1c3a85025ccb3f79446772e83f96d53659344c607744783fd038c6caf9fe0a9
zed7df15d0192e24f64e349781bb4607c38d5463f13bbc4318d1e49fd8edea2ab170caf661bf96a
z0a10a5ba1defff226ba070e7813bcdf51ddca8dc8c7c0069cafb58d0ca45241e522a218d752226
z9133ec9f1ec0e88353b7f8b2b098fd2e56882a4c163b3d9ffa264949ffb47048d136cc6c6c4319
z68339adb4f9b62410063826026480e3ab7e754c644098375cffb6ea34c8cfa6f43fab2e3eaca18
zbf601f028308303272170d0ef400652c58f0cc6bbd5045c69d36a0ff9701d05cc0198c49993749
z1b8e0e81883d91f88c14d4034824359d9803d5e5b7116e55ff85ef3708e307ac3725f6ead3e9a5
zfa710c2f031527339d558bdc9644ca3fea58983dd0c067c50b12ca760ceed25ab5c10562d4f6f8
z5d981fcf510da17ba7682e01651efba30c7394924ccb14909e257bd619175f22d4275076979710
zd1c2bfef5c6c231b6e0b8dc8aa585d6cd3587a0fe2c6b60b395a8197ab70fdfa97653d32d9a098
ze1395c6ba1e09aa1dfda13f4edc15f79cc7b2eeb68c731442fc76d7da91455e95e1c7f1eabad01
zc88931678c068301485d415f0880e824e8142a225a33c5993987dd02177c8515a224d02574845a
z051423cce85957d6a7c10d72c8a3d12ecb1e9937888e9c45ae6ca61957ebdfa0e0c7e786479f6f
z452383f416e5ea75beea855760114242254d594bf4bfcf299af4d069369a28581dfa912a3beab7
zed91a1d8704b8dfbadada9cf9d27a7065fb764e66dd8b2f72eaf16774cf86c0b6dafc2adfaf32f
z34617735338dcb4100473507d4124b86d85ca3a222215a7327c2713c8434dae6918bebd2abce92
zc28e644cd325fd728d7d8cdf140f0c6c2b2c4919e7f8e26093bfdad572594fad291546f8518e69
z7914833fb5449fe30327de3070f9ed6416ac32d139c198eafbc65ff910b980ac3db36a7ed1caef
z4089ef19328d81bc5918654859023984bb707db76f6fabeca5ab447c60b262bfeefd7347574b9b
zcb985e4ec71d509f98c29b5c0d94bf30ffc63f702e2341311e3553a98609920868478fb957cfd1
zfae74d43d4e72cb1baf5597d1e0a45dd64e4ff1877ef104a9d61c967742a79f338ee5066d8abae
zdab66f14bcee7a6724fc5b16e3103f7fe7806b3ae448f73da1beecc734abb99932e11ae799d3ba
z7bbf552bd5843a2300232db94d72e159dec4f7abcc07f496697ff4e801a109c296d6e82ad83a41
z422efdba3b86c67140590a18ffc97ee1257b7b447bf9be75c7cdc19066dc3ea5da304ba63bda61
z9d76414381fa9f4ea631abdbf5333f8a7657359a006b1578a4954c68a82e47cc64f5633397de25
zee2f285dfb0a9524c12a0ff9bc707b487517dbb4ad8089e0abb01e6196efbbe76a2ffc61457e3e
z2b6738723144e9d519ef0e03a50ee803ab3f269af3a47b9576199b98ce9e4275f6ae8b33b10494
z66b7f22091b922ffc7b6b5db9339a4566b99971886d662479203c3fbb8a80234146f80467c4456
za2ee6b9fbc938c1bdd39e7a666ddf0ceb701bf00ca0584b08fb441060b0bd50fc408489fcdb162
z1676ac516c54d0a5e7d245ca88316e0fa225ce0556c0c1f71ee5a80e3c0d7b99ef7df81b2ceb07
zb4c6ba6fc6a7ce938fee545efe5a9426d25e681eb6c0aea956c933b5222e2403efa618f4f65921
z88058d4d8e5d1c3b8b99d1808f2f79204d284acd57e2cbbad46d9bdb95313257824673f1fd9e83
z424a7b49d02b169277eb76cd25c2d484e8ff983f4047e8f5efb4ba12597d418c8edd677f542f14
ze7acce2e54e0491d27843a53ff96d009f6edc4c58f578268197ba57db70643efc73116ab3b848e
zba2c5dda2a5c008ebc4d61168f55cc56f32e8bdd6b0dfd7724184fb56310c430e4711442090f44
zbe249f6a5c425910e90aebc97111711530783f352037e27f67352d8ce4a3b42d840f64e6fec70f
z2a3a82c63bbf8223f11d15a459b6567e438c660b99a317eaf5aa877215bc50472f1ebb82a09e2a
zd9c0ed8351f7c2acb902924a531e5e4b18787487f4ff63b11ead720b3075f10e043d3ddd354ade
zc932fbcaa75da25e5d99c48420336d072c11c59832d285daaa6da7e3d01e2f7ef694b62f6414ba
z0316d8fbe5592a8e8033161a0726b06fa99ec4ca18e69663c4ac52c9c341ff81b81bb27c7e0de9
z6439dd6751d762085749237f2f227aff5475f3105fd18dd54a29404af2e388016c2f960889c7f3
z6137735635a46c6b2c31b43c4fe01230d47ccac3b8557bc5ed1d57c1970d35242ea4adb8f358ff
z1966584e70bf830a14a36a8bde9eca731b93911ed057158a7eba61c63c88e5ff3ef3aaae35f710
z7c659b07b02a3e3704218ee6a16159aa623417f08173df3871f7d42d5ad869fd83d12485a43f21
zc72f8d50648c8490dbf268339c3af6a621f98f6695a4c9b30252c538834b86021f0bfc01fc5e98
zdb0af4b23ff53e5d47a702a66023b5a14f05cf60648223f80c4edfdd463dc7327ac63415b6cfac
za4171cef57306e42a476360f74fd4b236eab14c0a9490ebcf79b39aa105b92c77db960dd4df98c
zb4642c6c9d1be4bb9c99214cd46d005c7dbaf6ae0e413dc47a97648d5ec966df99f92a2cd1cc1f
zddb01397faac1092a53b644d812bba9237c74ad6970e1533d744542469d7cff675746ae8361d94
ze2e22c43b148488fd3aca6f37ea7d48a4d6b9a63eee0693d55148225a09a3f75abea2d6c8dff8c
z7681628351af371db6bf5fdc034c57a1d960664ff86a7fe1724b01301d4a0b5b1882f800af57e3
z688f7aa731bd0267a6b6146579a5235fc13eb347ca6e8e24384bee1492c943b95247faff88c1f4
zb87895cb809c179707968f8fca578083a0820fa7d31b4beb0cdc4c4c03d567deea67bc7196d86d
z40d8f71dec7a4642aba4dd047c551bf0602524b11267355802b5080183f55bc41464c05e3f6ece
z821d00c87e087fffe4eda361578a599faca1450e76f567a77a25efb5065b42598e3970e4a9f9ff
z272a800bd7cab487c4f1b7ffaccb0972cf640691ac2fef2b6847065b38305eaece29452c3af281
zf83fc8d396eae9d5843499505158fcb495d744c44020c2e9af8a631e778319151542f578143fb8
z337fc9b3fce522ee8879d119419ecfa58977d7ae1b3d82fb196f98eaa02c24725366a7a24386c2
z5e9e69f6e30194a74c98f80f3f4415489d5a73cfe7bef855e0a12182e24385307db77b1c321597
zbde09d56614bd048cebf44167b4cd178db31219c714666769d70bbf4c1de4bf104f668348d5b5e
z5bd9f19555714a638e41182c840cefb1d790d2eb47af20eb55a34bce76624e3375365f4348e2f7
z5e7124a6bc359d8a7a93ec0b4e1765e665124100670953c79c309bd8cfe76f8cd5378d4324fb8a
z9d5275b513f26843eaebbc4d573ba305f8dbde1f5ee3a9a37322b5d3e329f37219d58ea1108b69
z408c6e2bae1f1587923d3902ca09aaa49565bfcec7f0e6ade9cf8f2698fdde49da5e2f93d643d1
z8aac16577d0a3452e3a82ffab0b413526a91400e38f734bb28dc700fa65a39d9350ca57ec620db
z5c8e6e14815a44f93c68be6c3db36ba06c69396ddec54ebe823aeef0c44d8023aed71f41803d93
z173ddf1f59da20625752ada997c6691ff160f8bf4ce48522f3f91f5267565f68ddbc27f6bc682a
ze571dfbea37e7616c81d41a9dff52a3d8e5ec5978a0edba1f7c15e00ae7baca8e0400024b35e6f
zb7c46667bc5fc860d3d6945e8ee0510a76d0d492230093ba3f5f35b282794bd864be7ae5c3db9f
zc0b912c6671281dda9a14703d8f0f484ecbe761f0aa4c583993ad0cd6b17118492f7a06b16f1bb
zcb14cd9f6007557ddf4e5c53427a23909bb57f2a87845f08fe338abcc4ee82a413edfe268dd54c
z173f88e2d33c797fd6acf3873aac46352b58488d1bbf37efd62780d71fa33f6c58a11af080c802
zb3086345c4823c6989aa0ced645a6712712cd37bc85fabbc990509c27fa26127a69dc79ee9b121
za72bfd4a540e92ec7d2b9583d86ce2d770d651b340767b3ad7879320c92fb70c9166068db11a3b
za50fa8c59c098a55aa3ad9385bb00a1ccff8f5e70ed112a020fe6c8a551dcc04e94a619dace738
z61730594104a88f70dbcfce4aaaaa48adfb5c5a252c18d49d933a1cf25a2d0aa3e0bc543ca3bd5
z48c5546f1adef1f80e4219875e954bd16d6fad7e0e043c61ea8b46467044660d22c97f9d12f7d7
z8a11163e6ab32d9873ea8e4be7f62f1ff4f9be3ee3617332e80a0566fa5cc866d8dc1cc23eaf01
z5508a1ed15f612b4d2303688e1e36b884737b2c7882f05a804e76d9223106d665c4fe3380cb674
z594579d1482aeac46ad75271732a53ac2a3a96c246277358b5634da2c65849ad7cac54a5dc8f4d
z5abf82a2b58917d1818e85d02b64573f578f81b1092170e352ad263380e79cd77d77f124b334c1
z9121bd4ff4692a069cb1af3a278827246b5ccf679bce1a47abf35efa2595fd6a3701048ecbca50
z99b5e03280187ee1177c284f8b7163ee83e4d15eb110c3fbab70258ed2cda91425b83f8bb7f062
z9222754c5e56a971dac927f9905bb2afaea4c149ed487dd11fd1ba2bae86d3e71872d348c36d9f
z813171e9db466f497310d3d299574c1cf778bcf8b060f793985781511170125c8f9997bc621d1d
ze12799ddf577cdfb8fd7c301bc947e61b786f4e6f829f483414106b4c80b2ef09b90c0d9ab68bb
z56528c66d4180df258b1770e0a4214b611296c76b771cb43f66d901eb4df76b4a0ee1d49db9da4
zdef5f4f35589c38498b9f838532773a261828fe58d5885884e6da81e25c5e4d0e9cdfd0964e3e3
z7d20c90f404a80f12bc5b4d4dee23395e5aee5988ff3d9627659a67f0a52a1c670c3d8fa63d6fb
z35d8a9edeabf3504b4e4763ef75820e969794f9a600c58f1ff163b39e058006ca160c6ab1c9a39
z9aff8ddf55a7c4ceab60df3de03184e38b7b7138c974488baefb9d7c5e7b7304c4d71f656fb044
z87cd4a259c5b2de518e52dfa81b5d982331f48d80031d92975e075ec708b0c1c9d62352d7ab252
zc5b450c876bb02351f8f02f8f92f677b5312b4847ad8a3fdffd74634c06fab3ba88188509e07b6
z56bd94eafa5bbd7bba499a8f1a8ab22db333672139f47154794234d414300d47fa435779bfbd1b
zec0e3b79ea78ce719b0c3ff7cda695b18bbd993f91bc8a056501ed62ea324d38e843ebed55f3ab
z28d6490fe7078a19109690330801d9018632d78dad4673610824fc5cc34dbb88ec6093b5571b80
z8dd11ba19f500de2bbdc9e494db7ed05ac5b035bf73dfd5d052ad91a44976b7a0c6a00edec2184
z048e9758e861fce904e82fcb99b5cbf0fee5f20edf374c32d15dab09782d0030e688d6067a5c80
z5e2f9e9549d5ddb80347e9fd59959e719c56d812656fb7496e1dcb6ad21ad4b9cdef5efe1d4140
zb62f5a4202bad16488ec1ba619fbe83e29d811931895d18b20980ecf08933e6016a41b1c93bfe4
z4aedd7fdbc9b73fb325d4be35ec13c1c92a07ce6124ce440e2e6cdde3a39bb6bbd18a0ee7f5414
z5cafa7fc10e8809766c4c229f7b99f07147839c8b54cb0d1b492f791d3ca9319492d51bd481dd6
zeb6323d84c421b77f6a64a5984c8f74c4a9093dbebb232ae4b4f1c50b1c61ebac4a0e6dc249f59
z1169ccbc6eb78452130302d2771520ba7a8ef26b85324b37291f2f00b084ffbde864522b294d03
z365155f16c5a49b52473689990af7b0fcf278aa8ed803c36fdc6ad7f5280db342864771745a761
zff555e824311a5b47eb0371228f0408e1d9e8a5c5eb64840536553406d084e58cc5df09dce9f42
z2c64e95503c8a26c8728249216ee00aa66cc80bf9b52e29bd19668c817b11c7816e1dbcbd625de
z0e157bf02265319181dfd8b17113116a4fcbceb6ec74f78d5c5b2f95cc91bbbc05cc2073364eac
z682e5d7981acc219b04cc8f3bf48c9807bc395bf3098140e23fe03482c030361e71034fc8d8774
z77250c115ae0fafe13ca11e6f4206fc428882113f112ce4eb3f18f20419549cb13433737d5a3b2
zec37229864f09ca7eaadbd900c56776188ac31be2136a23ef8da7911cb14bf49f3b0c038cd34b5
z888eb3ccbf450c779ecf241166d60991544bec935e1ea3c1c63ac368858c0d8e39da2449c2d0d0
zde7bfee7af489b023081b508b23988399773e4f7f25207e55f67a2cd2ad8e4f5f92e448e2c9c2a
z3385c1906ceb33c34ae70317fa893b92bb00e8fe04e9a74dad1e71f9d4cbd81d7b43a5e9f59f8e
z8752b9071b95656ec2a91b54f5614449f4439d35da004388f556fc43f2245e32f5a57240cc9829
z06ca58df47e3d27d801ce43ed0771f9e73df8bad249153893b770f2afb0f7c402e7c373dacf60e
z9acb1fb2960a3a0185c0f3b817d5612a15e8a1fca349fd149b418dbe7437d9dae0e42c5d9f6d46
zc7ef8b7aa21e7741eb5c4a37cf35a9977f4a656cd6f0af221e260d05e6627b03bf5d169ebfdd8a
za5fbe8c6e4352bf21bfc363364ef0fc261855ed3675d882592bb39b98c6aafbcbdb431cf2a00b1
z5fff4cc56bab274e552ad208bbb6431dee9115d87167022406fcf278f5ef449ba26c773cb5401e
zf86825afd5e5a6ee2bc7123ac92ceea69fbc8aafd5bdcc9c1a004f40893fae97887fb7cb087ad1
z2e82b6b6697710c4efb94080d5d9506c0625b78fe69c2f2b525e537d9fde4c475083a30ede255f
zafa99b8786038c597f7ef9acc97731e2c195e2530c338eecdb538b73cbd5d08bf1c224e5858395
za868f13be6ace9a72d3a940456013a7b2a24f47221864701708b36a64bcfbe8556144e3e33dd4f
zea246ce858ea5ee7adce54106f16dbde08c5889441b12eddd36b25a5c97671217ca23f6fbfdd13
z4e19be7abd97394d55809216432cc9df72a7b6106f7b2ff0e86bbebabbffcd119ceb67838efaa9
z2c3d3c79d4fa390ab07a59e5b60d275a25b7120baf76604908b1486628ad119cfbd5bbedb272f8
z36c08696e35146de7001b246ce368329c39f8b60a14e5a1d9929ac2bf3d8587be76b46a79369f9
z77e0c1588577b2143b7f6ba8e7a8a980c661eb68de826c72408bb3a6d427f4da8c4e934f3900e6
zbe68a3bcb9f3ea1e0a506c5b8f19e2af9c7f4bbbecf47781c011d41072e7c35f8799f9f1a3497a
z3ae088c704b1770e54b7c620d2ebfe41f5b6df894da2731651c2c06db61efcaa7552c90de5bc28
z19df88348f6c9e88ad704378155267394aa2d6cdea568eeaf402f8bede2559a0a024a4a606b78d
z77bccb4b3a47d3a5c6b7d6c6e32fbb0b4edc16d403a17b794f54b1603521b1cd9005afa757dfc5
zc21e3602511bd5eb49c62c56127dc8442b6ce8959bc232af995bbf46072226c94fdcdeaa9765d5
zd3bb715371991e219d70264b1711a0d200e7e90d40fbb945ad52e5e327042f86c995d551104270
zd1fc23eb94348f0ba4e58e1468c4b65157add9344cdbabd67cf56e4d41869c9ede2c8d4bdb3c4f
z0abca12142f098751af328023b15a986c8670a144b653fc9c6aa6d39d08cb83b5860d77c534630
zc4bdd9d80438a1f253d5af4ce79a39eb84ebb24282245e830abd1fda2dfc9c0ed00235af4aac66
zaae6ca896979522f9b4e62bfbe45ad439948f5116e0e671d8d00ab324ef695c05abd24c5e44880
z09df231249b4d1072927db2797f2c1c051d392001e7bc724fb6da534e03a6788e0fbb756939359
z464bf20270ac68ea5aa7260e8b1c33074f13c9237b6d315172a5b940772ff9ff055e1565567fcf
zaaa7c0b491a621c33db0885a662fa98cd4356b06e079d2619cfdaf0b42a5d5cba61b0001680eff
z493bd3addfd683d7ae7d67e3fba6a4dbbf77cb49164106872f7d05ac1e6dfe7e89395148642c20
z16f5a57c3a6c3c3f2db47651a9dc18773f9169a2c2e2f1afb48f1cbf691796b83f92d2688c4e25
z3c7adb8c225f936f31d9e118bad8a0f22704f416da26cba3c33c280faf3297f077bcb9cc91d989
z3db3d5e121f335537330402541c219bcb044439558f760791af6f616120702b653cfb402e84cca
z0b5becf19555691c295e54abf7e54c6a78bd77f98e131ad6172b46e923141bc179b8569aa89efc
z61c529a76f321f91dd7e83fd3934565b80e630bf00248703760729167a17c272b4fac12d1a5a5a
z7f07a7ae291a19268f1ec1ed7a41ad2cfa197e7ab5f80df88f5843fcc1b903cb0fa9cc80e25ad0
zd8b1f088e4fed42c87bcb3e491a8dacf666c9c50367d9f5392a7b15e9577d90cc73bcda4f52022
zb031cdc68bc64890abf2766add090653f487cfa95297003c89cbdd7e2f33383f8f4b1549a80c0e
zd8c376e3e6e7aea873161f007fa127b7dfa1a5b4a9412493ce51c02111f8eef57d6df3ccc07884
zd3d5012f1351bdee33898780956c198bb6b8e747224e10a34aaa146f8aedf8bfff3ce784f2ed74
zf3319243e7bc173ad6214832dabbe8ec0a3d263daeff812d728c8bc28af6ddc0fd46f38e641d64
z9fdcde1ed17aa6dfed8819b4863ce43d38f19ee50ebc955817554fe7a0f24c846e17f35e9e84b3
zbd92a345e09496e112309d8a54e0443bd68164ba65fbb7d4bb58c5fdee739abbb2609fdf967a32
z39a9d5a0a41418a9232a980d2ff45c86591acf6e40819842f5116c674db236ae15d19231c88212
zb6b06e362f8f35d6708a31485d357842479cae887d6c00af456bfcd2995da3bb0857cf7502538a
z9dfcd2fcb0b94f2a97c0b71e5a577a227c8d2ed23bb888d40241f147767d45c21883757d7b6cdc
z1691081be9e8f1e83849c827c645685642d758697f86b6632ba7d3a8f76a5fdaac3b3bcfcccdf5
z7ddda69fc617e03f0e7bd16cadc979745d793d7d8f6d8f00dc9606278668aac38cf24887f699b9
z3298c1420574fb21de0f70709d270cfc3b26f3833d727f75cd6d71dc0bc3a195237d623c9d5f55
z3699f8640b3d6018bd28d6a4b34e9db5229c0b2e5a400da4cda47109d2df3c03cbdf745b5e5f65
z65be83c629a283beacda1f340f25fb81a903f0b3e2b556665293b71846b76ab38ce5ece202dfa5
z7eebfedef12fa79f5ed42722f2fa08fa0f4b79da711f54915b7246465ae38bda6d930536e71ac4
zdf9ea6dfe2e1dd8b8a960b68c0e7fdb46403e94260978116d89aa49bedd536a9118846ba848480
z6dc2b71a63eec6f71c43481d5848acd78864e02a85fc3b089b962d65d8e23386fdaa534937d161
z799aae704df15e21f50c30dd9f6a508e8aa61dff44b0cb5deb5539d68fd5401adf32979f76ca63
z971ac41a38d92e9b103f6e1db76e5935549c5f914302ddbd772fa5ec606fe086e509e87b9be9e4
z77142c5b0b21c15f05151e44ec87c891c73149de63b4b6a42328413776b864d10654327b9072db
zc46c647f31576747345f59b27509ea6ca3086ce6a474468b92491d7f2a9b7bb12ef218590706aa
z5d39e3a7babb1942d7f0d3e0d2d116133528c3a9ff22824660abb9575e8e6975fea90d6bea4880
zf07fefe218952e0ac0c824a9e3333649d0b2e2d3d23d1b72eacab0ec1f96cb5e25806dfc669064
zb0b56ea691276b4371328f2eae50255eb7387a5aaeb9c67e8ce97721b7753e20c5993107863a13
zfe1ae35883bc0307f16a4c618125e6661e5260bde956aa06c888a0580c1229965f8278d89ecac8
z88cc5a457d6205319cb84ed80adea8bbab13725de9ee93fa8cbd0522f2fc22d0d46effa62d71b6
z571f5b02ff10fc68f22b2df3295761833080dd608665c46b21f20e2b9c46f11dd61618610a514e
zd3e1ac830a46911975aad31c5ac2ca96df96c70c8f20771308056305282b2f0dd0588c14bfd695
z3b62f6500cfd206c4b7ce27a7c6138e6b2cd39e9e5951bab28d52fbd3e1edf507483283fe7d305
z35f8804ec71eb81e19b616fefc7aeb584e29da138e941a09124ad67868607b5b475c7adad4982a
z938c684338d6afd51e9718c13aa60718c256f88fb53da95b5cf53279db988735e9a49de3af3035
z46e0f7caa0eb51a2c152b0c7a792a7b792beac119c6558cc565f5c4b2f475a372ddd5d3e601000
z77ff2ead960c1994cccf65fe99a6d08db861cee71627309706ef2e4141d500b21805debd2415c0
z5e10821cfa6bb2221ed02183af6a5d3c2fcc15dd720abd7d83dc96f311bd009a4c383e976f686e
zb93cd44149b6b43489753eea5604625f562f35075641cf13b9477dfdd9e2f8d7bd1e8a7346593c
z01d36cba9cc5a89bf860ee346baae3bea03773b4da52a239a99353e6f186c4a022c932b82a947b
zf9a8d349fe9867df26c77b91d5883f2c06c638d2584d5496b40b8e20b902795b76b08304f55a35
z003a83fc0a648cade9984507f8294de6dbdc447ea97b8c986ed30fffdba81701525ac4d117eb02
zddc3631a84a532cf4584b634e9bffb65ee6ccd345acbdeafdc8e25425c3fec3a66137308ca0601
zf0753e3993c0e3d3aec1f80f2c82f19446344dd64bc20a9a8a17525da2e186e9ff3dc797b27aa5
zc61e2dbf6d4f58e7b237c6e51f6d5f8cf7606ff71def343b142dd5debee956df66ba69bfe3ccbe
zb7fa82e15461e33d31f719a903ebc567d2fa33ddac49fc6ecafc06f6a8e55fbabaa371cd4038e0
z5300ed58abc3b9269397c3b15b768f8cf89021b4f889a7a7b7d3d9260d431b477488845c1344b8
z076e1d3d8550e352bb8704c4562344ad5192ca810175f7777d5e833f26c4e84022ab8f96856e44
zfa05ef4c536f5dc7bbe07f9dbdf94f65d50b574b9132edaafe7456ab0577694ddbd2e204e5f9c3
zae6b70c72ff8b9eec2db0cd09c1c8d574e5f312a814dc5314226d16f1e3a85332c1de41d77962e
z79b90b038e0f0c2c921a7c064528859e5fb0b29267fc634b881a1b0ae7c48cda80af240abae3f3
ze4b0a1b06fcc3f36f0411aa370c534d78457cd872a858d79b96938272034be092809c021ed1d68
z746254f03042f9b13da8c7930275b0d18db411eabab12c9d008853d35c5a43d96d5fc6a1cf4d5e
zb4d741e5c3544dcd47f37b88c5d996be58dcfbc4adb98b99d2d032de7d9e8bf3ac3394074091cb
z76d801cf0ea4a687230ca7ced28a9a53706f57996fec24962059a44270fc903c5591abd67c0cd4
z4c9c80e1d4ce0762cf222a918397696a9b4d4e21fc65c940e822d046f0f389c261420e2699dbc7
z0326ac2807b13f523222fc4a91ad50e50d363548619bbfc671a3bff5c80f5f85de4c1efdf1ed2e
zb591c7fdccfb97fac678bb7334f37aed307fce011244a5d3f98fa13bd60d1970b9294224d8a54e
z6c2ae5094fd73a607fa535b5bf605abf5879552c0d0877a8035d22ef28747538a8c72d4ff1ae38
zf04018be8153cdfc2ab859ba24decb517c69e62bb42c65a9a03753a06edd8b5fd235b81216aaf1
zb8aaf7a2402aee086aa6b7422fe701147e836615cfc3acb180a0788e33bca46a7b734b27398686
z885415272efb4eaa5f140744ccbc61543c523061b19862fc106f6a9dad914064aa01a8a1ae083c
z4d772fc019ef715e80739b751a7450f5093ca022a4e1779c5deb70b2d290af800e5520dfdaf81c
z0b94c783bd38feab031521d2804417713abca52a17ee404185bb8ab29bc2d92cc63ea34ba40404
z5bbe2055127303dbc6a3a7d01714c7fe3159f15b439add9ef6055c897408d957141eef555d7a53
z760321990142d08170c83ca7cf1cbd9c9f738551dc46652843ee8f2b293e9dfb9eaa90851cd582
z1e222822e13d9f5ef0f524d8c3232512a76bed50e4b60fdf82515742b167facf14857b3cda26c3
zb8fde3056feef67423aa6a88c898068012bf1a384307dcd3a833700ed1507e86c39cfcf7a382d8
z1dad66f617b0888840a86b2f3e12507792cba973f0bff2af720dc0b4141da47f2733fe811308b2
zdde212dd995f6e648b4f8049b686e11620599a537db4e30d692eaeb1110e48ca95a5a66de36229
z88048d9b348d5478877fb30aa155241c69276f7934ad79d69d9f5975f052b93e035b22b97da0ca
zeb307917a2058444211ef89feeae7e4552876e9175167528cfe9525511988510ff4a318587a939
z3d890a8c0d31f76bc34aff85560d5b16660861a7c5f0245bccf95a74c7eec6b9deaeccef6fae1e
z9375fc679067080b5f724c84374f8fc85446e729247cc91258e95d022c0a7cf350ef5b236f3d31
ze7a3ce9fdb517cca17e61abf21341c897ec89b0eb67fe41ece1b9d06b8a81d45b4c116f9f36b47
zae6cbe890d0684752b01811f42c840dcbaf52c882852db3d706a5f684bacc044da5c55c302a283
z28b43e3b10982ea4383e0cd795b9c435596f361f981db705c6841acdba32ca241b9f6a574d3a9d
z41dcd3b6d4d7a2fb21f032b69427bb27662d6f0d819939423a55eff75d0f002df663dc2ed49ee0
z4839d9e6275649afe2d5c10f56f2229754bac86b674c5384c869513090380f2c3a217ebda5c6a2
z4e8ca308ecf64794de933a0cca186a9d6e74656718a8618b211cd997cf423df18ed938d4614e23
z7d680d984980232ed40caaa900cee91a75603be712c2095e124c129ff4c9349558a48f4c1f16a3
z9558ba645f3a23eb87d4aa8bce87885213ce0070924c081a3d75ca41c91fb344bef7d373c7d77b
zb8066619b84c6bb057e8543a6b28b362d72b6dd3566a0eaf8a0679ccb3d5d8a60aa102870be68c
z2da8bddeec4cee0215b1e8fa820306dc72efbf589926a0464719ccf5213dc17385433bb40b5e0f
z55e56ee997e5c5e37c203a0335498ec8cb902af53dc1db794b9e9654d25efd079320d217afdabe
z2ada907244a052470965e2b5797ab92e6ac9d284ea2ca71d5fb90a123628d10673c6a2607d879b
z3c4cbec1b9e42b70e932762a52dc251f4d527a0c1e1cf2a1ffe880c82980c88a17b9a99504ebf3
z5b4085899c33073117159ec821c8d8ab5447d9f23ead1ef8ebf0b788c5200722c8a32ebe942116
zde175faedd7fd62ed2c460958f3f9595f94ec9264f472abd58c2da60d3398a20b505e272f4d823
zc609943889a3cb1a5300886bf64bb6627facd468d49e408094b5034f5e4d8677504e00a473202c
z841e681ff5dead079ade1425de00e7e4710a2e127f2e10ea60b083deb09ebf3585a576bdb9c843
zd3fdb37694e75ce8c462884ca808cd9a26d2f980613026751505242a4c88b6f054b828323e749b
z49a8bda310e1bcde8677e9245b70526825025a9c820ea6191373ae2d2bd909a59627c847134db8
zbf40d29717ceae5902c1b61732ffe96c2817ebcb5107b023b3b65f0fade0bf916db0ac47c021f0
z063cc7fd4e7149b86e2219baf2a0bf60767e2c3d8a3edbd0eff7a8264e7e1b0206ad06eb884151
zd5dc35c8f1a212197be0a124fe887813ff8bda604d7cc916065ba745a81502948bc340882daf93
z1a956d413414fe8c46a77acf21f8a04956aa4734799401520ed4182fe8ab2daae4ee6118c2f65a
z6283739e3cdb785fea989d43fa6bd9f941c424c0524e1d22413ed73ef4afe695fc9874f27d5fd5
zed8c3b158ac7f6c93d4bd0ed8138ba66f406bb724b1c3fd1616969ac012a8357f6ef65795ba6d6
z3cd204bd8c903cecfb8ef3fd3e84b084d6b027bcb63eddf50cc58ef20bd95265750cfe009683f1
za1777f5da6e8e3672d41248acac4ae7065b6f975817351fccbdbff4eccb1583da4aa79bdeff5bb
zd4d60b75852ed0c36c8723b894ed880e065bcf12278114826fba68a402f92c50bca85420cf2a16
za9405a4fd76f2fc62ecb71099e8a6840e4e1ca34fd2e30a7dbd543199f4328c5251c59c308d06b
za2ffb54450ecf32c2e8e8975525356b6b3cf37387a29bb97fa771916c1489563aaa762cda6d84f
z35489ffd22834f9eaa806897b521bb8455cd78da01444c7b8cdbf62e8a64ad3ad00092fabadcae
z629f4bdbfb1d8b8749cbac4c2963bc3684419d9217719a05f78ad57236cee1dcf273e30d248e0c
zcca62997fc58cb159d0f59e8cd2dc71fd0893f2b5951bb60bfe0cba993da8c5db623b81c287832
zfcb9ddbc0724167bf2661f8cd738b8057910254b515e732da5fae78ec12e1dab5e4b1366d381d9
z152dabddae7c3ae10dbba40726a4c0bd3518a93fe33fdf9a366f9f222b979330bafe0bdb0167fb
z67c467df5382a1a84daa03e67ab639662aadc6e604f57921aecd2d6bf9a1de11b0de57448263e4
z6ced6e78254556458ed0bd937c602aca378d60c303dfc788933de8fda7a19230e0db426cd6f87e
z2d5bbfa7e7a67038981a4044563029096e24d3653718eceb347d66f1bd243be03ce86cfc0e4ee4
zdb6959e7f93e9e4665b45f700e6ea92cddf9e2e2bdb54a742b78ad1f03b2912caf0a8d98620341
z2d4814403263766206358940e18ed7bd7a3b769a1668d5fdb59741c129880f7eb5fd07c515047e
z8bb4f22c735ff7803049d91e39d95b55e634cd5c8e8807df0442190b498a3717bc87d45c3c931a
z7d8b60dcdc31ff3db1c157f9fb4afba34deade84cd3b7a9838197b28ad75503bb222a9217769c5
z483f04fa9016689fdd589388b27689af781c32ef64f22748ac6b21558ae84c14be25ea41ad7c82
z2f575b4184ad35d3ed4d856d792aa72227c00777097bf2b9f796ccbdadc314f81e92d8abbf0623
z2956de3f68c2954f630d088c5f63836934519bcbda7452157a418c272f66610e7c17986e5f14eb
z8b3381400a9b15f8286134eae5667569e791dc089fbad5e870a627bee10ea5c7ec3a521162b848
z35c03a2ac5fb0d230517febe2e0f85a6f22ceac3c7385d4244ff9e0a10af657219452fd97b890f
z2ea0357d40d6f773d25e7e3aacec0d4e4068651dc93a5d574e555654a0aeece01e564ffdae85d4
z408027a5f93d853a0743b8ce04f6e3def97fa160bcdc59b3c46dac0a2dde89ca16156553168ae3
z69656238ee786e7635579514b8d75ee1f83610415d583ba6ac8015922f5690a93575018a42e727
z222b88c8803f69c4f282e938c50a5f1f9d16048284fa462ef8bd964229e0b104bc874199cc3a54
zbea86634c31cf3516311bfde3e40ab17595e38e7bc3e1a3722cec8ce7d339b184522e58e2408ad
z43039cbea9bfd756e7423162a2295e77b1263b04d6b1680deb403c16378b2059509f36599f8083
z17e46d435deb16786e078cae94e86314ec9503d029a4614bea0bcc86044721021ce4fcede7f95d
z1852ec99d690117b56a31cf02b1532542b5e9f12e272fa5c72cb78c97c8b8bc5bfea4a383cbd63
zfbd2e179975bdc837a88783364dd44e52a673a2bc8d432b8c210c82ed3ea56e724c9a731973d0e
z12e011a18b1defbdd779ed3df651cd367e16d19d6f4ffc61fdd33836e51ff7552db0a4f0343d33
z438da58c69d3eeac7138d2a5a2d3bf508092e0cb4a7b5d41f7be24c2595c39efdb70f764b9fe4b
z92d947d61ad786d9371c2c596ec67149c9301750f1441fb3e23b5fc2562d386cf271aa06538830
z2f6d6e0e5c5b4600545e9469ea0c03617d8ce79c0e1ff71048a1651b242d1bf331883064ab6fab
zcb0f8087fba1ce65f83e10eaa325f204d15d3c3c6e771b5249c479cbd6e0b76fd5552a3c044c9b
z800b72aa305c07f8f8263c774132cbea492ac7ec3d211868d608fac9403a96471d361a7dac9c12
z75e6f4afc4c9bbfa3d98fc070d0d64d028c15ef90a8c225743d394d3b2ce2223515207112053b5
za63a7da95c45c4fcf0f0df8cf0ed108ab1273fcfadaaadfdf462950c63145432967d18cf228b9d
z629512e02205928f74ce1346e94eb0bccc4c39ce397518a556deda0ec10319bc645ea36d5d42d3
zc3f5c933c6c2faa6b86942c5181e8e8c646991fdffecea88ea2e273bb9d5427bbc881e0682e1dc
z32dbbeeb26314ed87e84f7546c44c5a5a22272ffb8898943f92e3c8bb5185feeed3acfac60b1d1
zc56186b199db4a3199e5801709bca0c98f8095ae90876be979cdb7b9729969a6ed87ddf9e330bd
ze0c54b5a257fad367068479053f3a888e35ce44530b7ca55cea2e9cb9cbdebce2d0e0b6d45fb4b
zdcec51269ef3ad6f8acf2db2b0a24da2bf193db5daf4083e6392656e8479aa85e30f8fa5a71cd6
z0646ee6f04d45cbd9a845a3db4c7232c6b871af2d9e74b5d73bd058008e4930825a4cac3c6a13b
z45e3b9135258203b0d1db3a1e7c8ca0c5a8af5faeae3cb13438a29896fc08a67e24f26ea4f11c9
z6706efde333791b4cf33a9319bc05c712ae72ea4f7595e82944741a15222afa530ed8ce13d0a60
zdb5fe2751afe915837e432b3f04c080ffd92b243197634013b6396f88f460aba704d44600b710c
zda9815b066dd4393447fb8d2539525a7d730ae8c1b48ba91c0a4d0418c200f64ad736b0a35b44f
z3bc3c238135073cae5734b5c1b2593b6d193b610f73102b585bede945d6d51179bb92aae932a06
z1ca22d6325cea07faad0ccbe2291ef6506f8e5e26a54ddfb0534f3e730d5f68aa047b9b2c1438d
ze50785618cf231e076541aae26b1f1958f756fd62b62a88472a5aa5efb5450e3621474cc4c6523
zf9e29f91f64e163a166fde70680713721ed9e20f43480a3d6e0b8d793ab7bc147928093e9336df
z79d4316a403d46acfb996c907cc902976549f1c7f4d17d8f71ffdb6a4f9657e7646d93b556b547
zd202492c73575d427a1e1a1dcec7c9df7b9bc6bb2915a430d2a6c93a6f4844138e4de65c54bd2d
z67f84f7a0a6f7a13a050368cc61f4ea76a6da3806572e5d64d270fb2ecbcb401dd5a81b7bdd08a
z2b3d02eb0d0d1d0f7ce35adecaebd45c8a3beb8a5f6e53c6b4940c6bd9e4ff57cf335d81ffeef1
z5d7c79564fd896d790b99d1186187d53c4916c21b6c63e8cee75452a284101ed357020b29e3b61
z768b3a2f58dd3a990ce117d3157807129ce5bf452c4c247fa25e6c865021de81afed36ecc7ffc7
z96e96ca96b18bd0f77d9b9ca0faab2388914c24ccf3f7d3f7fac70d40f28c71d365628b3a00ada
z4b0711253f7ad34f07f4479d07a1a9a3393c443797189122a0390882792c751f8357d7a471f86f
z24bce629357f3eebe3d533f9d9a1fccb629c82b3ecb741806459e187186b44d71f8b894862b098
ze086eeb3888ce88f6ca1dc1e4a78906ce7a6466d3a5e472af2794b386fa3c22eb6ee459d8dbaff
zd09d4a7cba23ecebcc5ec29e576de989c8a3aacdc3a6fec91dcd361c5f41ddc81396e2b7e2e65a
zb61067cc53ae33c1ec1312e2807564689f226a00f8663a0f682e96a7371931a96056c478376572
zebde03cff6e02c18f6aef86f7028ca3205bfb25e383b3e43b19dfbb16cc56389767b04b5123187
zee1b74eb79d49689ac075aa309d390b7361245ec82e3969683d50dc086974af4fe468fc9cb95b7
z5bb24cec2b76153c7bf370bb435fbff44bf99f660cb37cc0d01769eff70e67454d4d0fd3fde659
z18d37e9d2f24abdead0b2ea862641925fb4da0c6f5eea8a619609db15c7df10b5c51fc6c1263bc
z5c0713b89fee3082e5d738efe61fb8e036fb18383dacdbd5be998d005e87fb16a959d45a7cba53
z96c942173dd7e3c110606c1bdd570763a46abc434c2aa1cbeaabd9ee0599828288e443e1c13ad1
z9b2266d22129b8da43ba56d76928780f2c4341446709717dca166280e4d31eb22416bbdfa4255f
zbb02119fa2b1139b7e617ec6fc63b0fad8bad34528360ad6acacc929e7f1de9dfdfa3ce4ea0e55
z101087d6474b70884023c58a8903768fc68e57362702ea51595f2285720c4e3e1582bd11c78162
z5d8a5f3b871528f9f161ef4230b21cc6c15af9ed7b5b73db1d18b37b1416003f22d420c72ecce7
z796b3a71f8f2231ed0319f529226595b0b0de1fcfe8bbaab95e94869444bb1cd6b8cd615273684
z11672702485aea6633bf8e2a6b0c196143ccf2b4bd88bb2341cfe1408f93e1ca7749b2d9cbf24f
za1189603ce6d22b9f535043ef45d995e5b8ecd69433207ce27cb1c96bb95db28b7d363f34368a0
z6e5d54d1d2a22802d5c6cac0dd497c4f477289eb4bb06fa93219b58f7f6d46a6a7ec3d337f0e36
za92e56779e59de6fca849da445d23899e837d20aba5e38b7a14e37401d7f16e4666f9bb5d03bb1
zca95c79df3990496fafb7fcc66b96305dc90037c05a8c0ba03944b35794b64f5b0c2ec6c2817f8
zad4f465129a1ae41ce290519498976a077403a6d4e61bb4f4b700a0df0f75e65242d7887cdfc5a
z5848fd2a61e4fa750452dda34456d28199d4493c8b42f803324477daf41ba6fc257a163d817bb3
z5831434718c9027baaf8e6dd4055c16e53170a68c18b34ba2e241c93d1fb87acf2d1ec2d26fd27
z0de80791c057aebaf072a6a6554440d331b696571b78a696ddef5f63cda9292a9eebb80a2e9c96
z4fc3ad6e98d3740ccd79af2e5aca6071edbef037ab789f5e92320c3a7f622b93742e48ef751739
z58261f1a4c75808046235da095f51aa21b8e0a20d9588d19352a36455ddb59bef9d433f684491c
z0b26f4d17447badde14d206afca9eaa3abd67f192b861c4d7d63f079b47b32f5f0accf2c2e29f3
zaaa090a1d1d7d4fcacd0c19fc0ccc9b69c861b2211c356ba76b0fa1632036c65fde2c19b4f7c8a
za60669f7e6fbca69a839efb84727945ee5a5cc61a26c36b05731c85e0888e92e77f3e537b5ef94
z210aa6d3e73faa8279326ef40c5b32505f4f09af33a8d442de31a1950f22f0c302ffe80fa160c0
z3d56e85c6df8155b8784e6f9cf14de634c339f2ee36d0327e089dc595a5f9d6cd08afe410e7814
z256c3e29f5b6cbc979ca0c0e1515d4644a15ddef7ad75e911cb158433a1369254dd364e80aba2f
z8585ad54334297d6523398ce804ad924b167837bf13d5cf54862430f7795299009ef5f5cfcc29b
zbefb37ecc1dff1cde986200837c7f6798e372edd18e0fa61e25aa809414f13a65497a3f462e735
zcd737f0870abd9aa047ba1e59ba9efe17eaac14a2c999ab15107f6ca58b1dcdfd7c18006aae7a6
z8704941dfff09690a34db8b132e592ad2679f5c4221383f8f776b84c29808ffae75ef7dfa67d97
z43201b7a8659e65efe48538337bbbd05a2c7cadd2e0bf6ac892f83951fc8ed0eec13c24a0b8c97
z3b25637065ec201783576be1f735587066f81de10d38ee87818269e328b5ba3d48806d5bae45d0
z5b54fdc8d448869dafd00e5d8688a5107edbe2e680a661fb47a610ec5432378523332dadeddfcb
zb2bf00e2506205a2a16edf71d4d98636c4f6b98beac0ad93e54d68da6ca3208838d13a7b7b0c1a
z6d1b066f32fbfdfec5e34832aad93ce0c3edae32e22bc7a8e08d267871c31f9c5c2a1598d7149b
z70dd804ac9ecba84ccb60c9eede2c63e82e5e3191968397476ecf724e2342bd71e3a38a9d45aaf
ze707f6ba3633a6cfb39bada4c9a3e13bf8026acbc78bd390fc22884937010e23136bac13a6201c
zdd95635d747ed9538dfcadb6888a79ab4b547ff9978f25f2bac6cf005ac36a5e1f58b7c770f40f
za5f5400e7ba1dda726bac8e86e4dc9e078a9011a750c682fc9082ec5f39f374974747c361c59b0
zfb45441b9dd10d385f42bd8c976e2aeac46a6ad0d63b9fe5f69b1536565a9c29d9b85cfcd34328
zdc220ea6935818068fa96d20475bc88cef29a81b21a2af46f30fae6e0abd516ab87d1138c2927d
zfbc8000df0308248b96062b6e310d756ce37355bac7d8bb12e784571dae3b9b7c6fa265bb1d56b
z0bb959c7ba2ce3754cb3804f2651a3928cc67f3b49eaebc33fec6905795e7a8e964d3c7bcd89dd
z5a94665f8a5c8ed103b75b83f19eb1c26da8d5361ee8abc3c9c7d1ae8bd4ab4aa39c04c0a5aa5c
z40c007a589159ebbfd848b57bbc9956d67eb146b6da53bf75b7aabf42b0fa8bd03f75e5297f735
z93715360a7eeae6a14f591f14cf3ff08ec1b285eae9fdfa4ef17979bc7a401cf85cdaeed5a41ca
z56be083e842955895ea7c87036a7daa269b09aa9e3ad812682184e62030766a71a835325e39816
z78bab20d52ee918e157e99873142bc7b63b068eb4accc1a916a1476823e155ddc599c0094d5c67
zed66e46fce75bd5f2a81967c14b4cb00cf1a4d0d3258464493c06cbd4806c760786730b19370f5
zf19ca97fdc068895cbf07291dd66892d44bf5bfec6a96f4da506fd6bb453ad4562585ccf201998
zdc610986ac2a8b3f1a97e68e973052d9575c9a3904e059673176de1add5a19b3938ec01d52e603
z3da9892aea017db1f2053b4a9d776d5ecd7a174974f19814d73104f5db2a97137ed4e4bb048363
z19c9a71d71c9caf2547c2bf661478405fc0bfb95c676e731fd2409d41451e42455cde0271ae757
z0fff70c457e6554a9559ed283c7baed63f87a0bf13b31cb703706c51c7cfc4923a398d91570666
z8e58c322a73a95191f946448a6b22064533ff0e5a7451995ed32af55120902334ae55c65670be8
z24649bf5277a30b84fb8fdc6f8b201beb79032768f12f7f3c8028b6d632841b9f0ec3bef3d5e88
z236086f5c32f64858e22ae5f1c4ad57f7c3a7086d2e189948754d2b56634ac99f1fdd1493b880c
zf57cb9fecd58483ccbf2120330b462da349cf05e98f0e87696030446f6bfc10d74d91d1278a632
z28cab32736da853dc9d0a9e297bfdf37ee710a342801dad5840406a8530919e0d25e33c2dad5a1
zf95e0f979513a6d670e8693c9965fced848cdfe4937571b87d62de856ce0038cc598cca2e234fc
z4122046b61b289beeb7c8cb5db44773e791a9a1e33e6a92b3bc40272a66fbee6cb5181387935a6
z5de40e26b0c826f246f1facc704aa7b55a7c1ebf77eac5569b9086251ae45592b2da4603dedb98
z2c0da45ab62f218a6dcefafde4cedaf32e55a24f27b114951d680e16ce8a2f5e236ec504467ac6
z20a6bde3bfc0a9eb4a953c4d5f56a8c643b8021263ef97c157a80e7c9e4d52d13c599ea08417e1
zcf1a3f8732c9fd40f5dfb6a3f7594b650a823f1b4e837e7a8207d8279b13edaa3f6a1ec0a9fff0
zc0380b762396f934143559214ddef1b146f8246dbbb7589010e4b463e1ab6970510e1e9219d62e
z262e0f9a5818f30b56430db400ec7722629523ace2d81bb4d57b548eb6bff6d9f33b68dedeced0
z8808bfd9100102557b8c165cc813a323a59ca858ad00498c4f7529c8df509599079427fb320f37
z002328efd3d636370d96bb5613d6baddf771f49ce6d2c2869df279654e1a5624bd9746e48c0959
zba48605ed8003349e647f40942ff918b209696845c1260a2a31663305ae42dbd686e7db4b20e9f
zf7c31c5d3f56424537004802b21ae1750752aab462b115d6d1ff992b9103a8d21ed70e87e3bf34
z3e9c66803ac257fefecefc5ea880d1950f779bb292b2ed071ffa8d4dc1da4729d4530b069f52a8
zbcd7d0f585f144a771ffe8a0a5ee877316716a2853be70a47583f3e7498d3481d95c136d52196f
zc8ad32aaab7a911952bf5ba5afaa514c962d2a8bf19282f50dab78e346798ca48868abf2bee6e8
z4de75e5c47bbfd583a015efac6a13bf66522d002874d89ac1cf671142aa6b3a27d09bee1184227
zb3989e6931e695934df5f1935c4f8bd33be7ddf0377fa39eb7b3edbe3c1a43ef7e6bcc11077720
zf580373e1cb57cc5356865414ab476f5967999d6de9ffe518233c383d17b09c7e7d0a815ac5c11
z130cc5fdac678ec28c8ae389a2028c93ba600eadd62e309f9d2d03628df1a27855012e9204541f
z151313151d98d679132c1d0fc422b33f04618d8f8f6ce01c4434288f81a93ced7446b4bb78dda2
z87af96cfdce8bac32de82af9636be6929299cabd415d03005b6c15e396db79e13a66728c1f45ab
zdc353576d658e85df13a2348bc2988aa53a17ef1ecccf3280d610a4ce7d472bebd53197d395a20
z85be2714823636a2c66272dec691fb9038dc4b73e66ebaaecf80c7f8114e70f956e27e85948aa5
z1fd5d07f92e60214edcfe1aa8931dceecc2369181792a5576c2e7a052f3d36fd8bc10c5188b854
z8e6f37fea9bed514102b914355f6f7b09fe210bf88e0cbd54d5f2b5560d09a3dc0d2a1ee68092b
z20b2429d03a1eeb72387552a8ea307e472efe208a0922b5df1ee702a45207bfbb9a885391fdea0
z3066c2818ecc2f75ba3857f12a76e09566be7146aceace679095be8efff2f46302e5fbfbdd2edd
z0417ad9e3ef5ab3fe6cc510ee0ff92a810a2ae90412c946901311d2f1ee060bd2c1edf2a68911c
z9ebfa8489404bba46d2943e46d8682ad6eb91bab70b7201648e74a54eba050213565a28cb2e819
z794cb04a6572b48f4d2733efbedafba98c67cfde8493d10cd5ece74ad74a3ec2e5d6721a44699d
zca6d3d0c3e871d7057c1b73d22233b68ee8dd4d7f0da492a0b08eda8aa90cbf570fb408f20c216
z01e1db6346e1012dfd550a3b5548da1c7f4851594ea41232974caf0dfd82a982edc230c1c5b142
zb0723825c2bbed2848a385af5b6845bbdf9cc3ad82fd373dc7eae35ab8a9dc6548dbafd18338d7
z6aff490ca22b30f8e27ab2dbb19f82ae7f1bff3d15a25f65ae9a92b0ec5afe7c98908ea408d9bd
z6a08b459a7c29bfcb0ae281e13450cf21a81d1732c55f1398e64c04351714ca075ce3707695172
z271c32757033566b044456a767067dda5b47b2e2ce2b38c2092ae4683ef1c4079dc94447c75013
za4ed39fd8857e14ed739ca612f21cec4be721cea58a8f2292dc89e290600eab421c8b240fb6e1b
z53942d5b7ba331a6d1ba60d1cf6815caa9787064dc6e3be6411b8d648dcbc7ef270ea58b05e978
z6240a1f5541d89d0d4310b95e0d3c71c342034cfcfb92f6ca21466569154f9aa37cb7ab2a8d57f
z2bff93dc3a2a6d23a073d2c029a25f4105f0ed3f173c27b4f76c659755ed7409eebd67abb3d86b
z12175f276739983d6f196000f6c983b942a49ccefec0c5dc2ca7a59e7ba02a87d95bfb7d22db9d
z7b01e85b389b7a66ae34c8d9e5c16097f02b1935de60d5e9921bb9e4a2867d2aae2c0d03b37e6c
z1835ad0fb12e2b7485845cfe2d9292bf2d8c93524845264ab5b5533b6a94e30331bc3b802cb15d
z55a9d62d5970a96715d9872bc1b8f7dc8f153963b38ba4b39dd511eca4aab4d95889c703dc45a1
zeb003534de147c9d77c77b306d67660840be22b14f68f59cefab55a923ecea80714712a3faf81b
zc38fe54cd68bde69dd4975b033eb260bf3829eb0677b88418b05c66f785f2e59ae9a1b96e35121
zffe3c95ad40a9a4fccf5b415d17e94935105af8771aef40685889151a041c34d3bd3c001897f8a
zaa81bed4a5b6268af48f084734dbf63cfcae965d8a79c33ecade52b0e1eee54b1e2be086bc9f66
z5ca70021df997dd3d26afac36a605d37970f2ed04f72832fafa2a4cece425caf6addbd47739a16
z7dbca7ea4041001b50cfbbcfbba3a65971a3bdc3773fe85f05fa146bbfe46ffcacfd0d7136ad64
z7ce131b44bff3549a7f06c332d527e2df2b7fab4d17fff5c5256d8b626cb55064237c7f1430ca8
z64c6889e4d43d0d6537776f4a00f15e0883a17d6401f1f32694d443cfc88ea3b2ea99d9a1728f0
zd74929647cf6d2ed7d7ac7d0d7629b5b9516407f0bda132b87fd284374a60eb942d5887bc478c3
z5f48e80622751b9f07d395662ce0a1b876f31bab792a74d843cba808585b96dafb8980360d51eb
z16beddbc75e4067ac3bb96ecb332ec7af38eeb8365cf66f11342bf887bf12006d2282274c2ecc2
zd67b14da35dfb2dde67610f1e613c23c48b57b4d80b1c5277eb10d9b97d13f7658c1e6979eb844
zadfdef6077acb090240f47f10cb0aeaeef971799f4abaf34612694b0103ee8c8d35513e656fd79
z7a2480c72c5e20e4bc490ab1e58f7be4dd8bff44b8f076c3071f0822dfb915c88ea4138b7ea81e
z8684434c777c37a19ec5cfa45effe8e4b34ca5bfee69d12809a9d0402b5f57888bec182324ff31
zdf45069ce5864d9175219676df4f44e76334ea16cadd35e2df947858e76781bbf35f3248992cb5
zd7f98fd0521f8ba378358efb04d853bebe88eb7265cac445e33730d5701a9bb5d44d511120415d
z3e8a0c8b5430ba2ee1ec67f49f9190f073db1e82b8a09ad0f41e246cbc59fe1ec9847273007148
zf116eebd224c32f80d3dc7e32fbb57f0534c8ab2368249961f02a3abb708a03443cf72abdfe504
z7a3afb3ee3c96839e95eff1061152835fe842b5b9febf37239c30e39d0b2a716589176578afeaf
z50de48fa71cfc2251de0526e427a77ae6b261e2c46d42a54acec5db535d893b5702577e31835be
z372df07b44fbec2811f5b46efcc653851476051bca1056d62a152f84796fc1a04db711a27e11c3
z34bf3cdb5414d15d9e0b5748a89b056c56b2cb9d4fa0b28a1f607fd6e9a0add69daf1d9d605ab8
zee6efa139090fbf8e2ac2dc3c4dd228e003c471cf557929ae4564e8bbf98aedda4170c81dd1bca
z342d40ddf9cc7ef1e514738f743effac4478102e90a73ef1dcbcd0c0e81d4b2e5b34184a428a9d
z15c42e07c77ff47e0a27c28b655e30ab4c6728521c644147cf75fe2c8598e26d518306e1ef85a2
z6e681fdc7c7846864503546ea008b084ce056362084b6a340d9844c3e91184b11880ecb8c43f58
z4dc5f0c17140bf89a61165aa3127612cc5ce02d76908498720cd1e7dc446c683da44dc9385b0f0
z4a9b21372d2c14cf4f4f5791652ab211ec4d8c909221ae5d085895ea50a8448bdc052417bc05dd
z491b7c59372e188b81b0500713dc74e32273b49b8a41731beed4670e75e675b0815752603023e7
ze9f1034e4c2845dd5446ec1640fc76baa719dd6d2ff0cb589b8d64e5c4159dd8f8aa8e4864708b
z68b213ff31823dd00f6da716e5bc384a8020b1545294fb67764f0abb35959492d6d2252982745d
z66aea038cbfd76f1b4600f1d708b20199a77381d50c2d5a9b14c41be4d52595b020883e093cc78
z12ba7b565358d880eac66fd4a63613c76a9e8a7426eccc0f0adeb564db8231ce9468bfcbaf4800
z3f72ff479af197520f21e9d941c1d69c29dd3008c54340d64a800ceb6748580645a952c25bbb7c
z235c003a8b6ac4fe2bfc4ad449918965385c205b33453ae9c700f6fe0427a02115837eacb13d27
z645b8e3a655c4f4520cac56f258c80292a65b6821ae843afefbd8688ff026dd8a78eeeece9e051
z1dcaf892dbcd311bb6925cff5a4896b51465e78288d7c25092e2cf82e2435436c45c84f435367b
zc2252415451f1a0490b2d265dddf12c4b3dcd6669aec8241ddc98429641b774a2507388b1a2acc
z0fff2d29417e16314a010514352b3279e2b7a47f16cd24ef2f03034245f7ed17e6b3f746764c23
z83acaa6ff34ab7e104c1c024e03cb982f0d1737cc2a9617fbd3074378e4c1097de07b1aa7db289
z5d572fc44b7f8b791b855377fb250cd9a1a3e62645d1a875fa940f3a8dc82737ed2256301bf1e5
zb4f6f34a138bde8588592ad76c5c4d75581de725625903789903d5c1fe8eaad17190e9b76ccdcc
z74fdb101d8478a6464fae6d38e6748eb636ba3e2277b0ddad010cb5c68d11c6ceba6dc6e25abd8
z6ca3f0402038118911a3e5254184f991976e4bfccf54f138b2befca0883891b782c787cd86ddfb
zc2bd30c0a072f95992f8fb505d6f666c87b62b55422c23dbba3e55f44029f5df4a139a0226edfc
zad601849c444ab9a8305f03392f65388f8f906cb87d889ae4c65356a2e7bfad31def544036618c
z1cd36a0fa47de468acc6c60aed57a565d28c51f1f48f42cb6b0ba9affd0f01717df503a0111421
z3ebb4c55b73e46b1e4f5d4715284ecd5333e53e5e760f771937bbab20f1fb890e76ec170561c1c
z00d368b86e085d75633397c6adf930931eb183c1ff01b9175d636e95b7de6b3295f732f87ce3a9
zfa253eec069833a64acdc2213e93019fe2a5cc4d5bf28391d145cc1b6d512bbd62cff2b1b29dc3
za4b1df486ae3bf3124136a11f985ae1feaff76bfbb9d5e1bc3d8bf742db758046c55fd060b9cca
z008854bd23fd6c028f14b73ac748b44a1733705b2c9e9cd120a675d8abdc99c224c8c3de1d2aa0
zffea8d37c0c8e0e829102ac1d6642b5cc312167c4ee020427e1ad055741b5e858a75fb1b00301a
zfb94cf5719d937753a0802c27114a4494c8b816c0ca96df108f6814f02f49783849812d0d51010
zb476ba275828824150bf663f6049e71d22ad077acaf21723f5fed6eb5fa429f3b9334284e0e649
z4f970a96a42d5e74b15a6e9b9374f6d862315c10bd80c65c306aa4acbab18bd3af862c62abf0a2
z9a3a999b7af2a00f4d0f3ffe93dfb990c5cfa7a980e2517e3e6f87ed059bc8fe820b8a35e266d5
z8e1954ece56d2a5ee32a1ea3cf60f049bc3a7c624b5ab4ec9a2c5b9f28e83df902888439a015d3
z9dcace55fd28848ec80701362a7b7cf21fa07a30814bbb69bf738b49502ad0f25b13bc700982d5
z4846d472027c1f9673dc9e8b14df4989824708b2978a6a0148dc1dfcf9f253a34160a761461d4c
z2cdfdb59b03096086586c192f1d32115642bf35363dcb0a3dc250e800c0c31b3c4eee12ca3e93e
z88fe5fa375d69466f2ff755f0db3f422531b2d9c3bc535f3fe53d5182ae1cfe52abcc3c445bb0a
zaff42c9e802c35c7c6aab90a2e734263ba8413a143e311a15c318bb7e35bd0e79530488dfdd00f
z44b326da2cf7c7ec81774adade9d4dab5b066cd140b74e5a48ca4bb3e916c6f8e359ec6825dfb6
z1544d89e43543998fe11b49ead37396fc97e497ca4f6290477d3721d6153c014696f4d9e9c0922
z4265ee310013914229e27b121d5b22eebffeca70175b1f672c9ece4d473beaea5111f249142407
zeef554bbe2c8a89cc2ec219c3898d3e9744a92b50378505609ee0a79e137916038a1fe160b6aa1
za892f678c0e9958f6f9ba622d1d84048ab1f8918cebf8174a8f9589f9b99f9e8cd98d3da23ceaa
ze2fd8a38bd2ae1d165d994990a94213d2d868aa61c95e9842eeb9230462e09262e859146a1eb86
z88c8e27ca5934ff10270c18ba62143512b3d7ef597ea31f0431cedc5eb2302344bd82286ba8725
zb71e2bd2f0beda81167c892c38edba606503e0b201e00445329a327587be74c8f66fb390679d9a
zf888868cd1f4cd16cf4e7d2509ce1ec97f3d206a09d02ce4cc9481714b65ad028ab96c6f3159cf
zb38c26029a79fdcab9ae7163588297b2c574cea3426fcc7b117252ec0024014c4fc9890be4ba79
z499fbfdd2defbbe4050d9a7711ef509177ff8f41d172fc03255cb39d93ec198032f90e30e231e9
z41dbc9cd91c76626bf78ed288467c91e26d448e683d69ed30175ce9723bf5e6af9a9ba599fed89
ze72246620820db6aa3b805dc6f7eaf5d3bb6ba31064e9157ed1b24432e9dfd762bc489ad4188df
zdc97ce6d9763a55e9ce0ea0b9508546b2c5a0e0db90380601bc5432f7fa6dd357ca1ad11494a08
zf0ca6b4cf778b74489753de7043edee7769da8f3a0aed1b4013375782c3ca493296f2b31aa1f10
za3184db78d018285e1f59d2ed1d3944a1ea9baa2b438062dc99bd94b2a17222159bf83eb4abcf6
z26a087da819f868a96d43299c63b0e2eb640cf9ebc1f53c52d080374c026e5ef8b909cccd8178f
z4b60eac4eed80efce2415151df1c8b3caf8adfa0117ea2ee701a4c120be8ee0114488d2aed57db
z8f0f51943c77efb6997f099f87d85d9c86c13a2a285f1083ebcd9e4fe451494ab51781b04e0679
z939a3d6a77d2580953a2857865bad923679f6edb317aafed46d4c5e9a4d90e41e567ce074b6ea4
z51fb276a4cfadb6d27af4f30e0a5c722d8272f46db7ab3e55be60a99f3688f66e27382af3f8d51
zdace6a04c88887de7c36d09d770e06a5258c2ac810b9d533d52341d877098d1acc48a0a21f3f4b
zd35c432f61126e0a803cf7009c332aa7bbed9c8f1f4fc258924b735df9062fc8dfb3eceb4f3051
z19a037c5fa64a01303770c9bfdfa2daf31065cbadfe28ca83e3dd6c6aca1a3bd4534f214e35365
zc303b5ce50afbae988f193b91d5be6621909954b8784a3b003da532eadb1c5a598cfc911013986
za2065479e2b9129d613cd5c5374382a5051dff45b24df7794647551a02251e183bbf3becb42f5b
z4d3ffc3eea58c6f69ab402e3e63a69a2f66feb266844796d69f70bfbfad8f4048d4a893edf808c
zfca16c8ebc11a40aeab5264a08badbd7cdcb5451c1f191a7bf39feee0470e47253f4c40b544d2b
z4d646cf030fc5c2c85b8875dd50b556d2848b4f6feafa74649f3854048b0fdfde2571d36624467
z5690af55fdadda9116b2812e4871619b5ef10dee190cd7d4b8e3ee2de33c1aea1d49bb558eec40
z9d05d764a9df8591f324ed755c79d992b376ae9b16f78a3a288b3f79f8717ed74bc474d49bba27
zba5a5abed41ff225e6583913ac6eaee879ba3ba739bf7fa6a9fecec0db706dc6cfe03f3da1ea09
zf07d43454601320fc62422dc4fb0141233a6c02dee3f37716de7cf5f99046962b3f8e04af1429e
zcc47f060e5b7afb8d2d96328d3062754b740d53711bb0c73fe0c9332d15a0c1fc024f3f2d0fe94
zad37a003bb8ddd63035b322e5a532e98e65215636d8fda37cdb53cb9ab5eb3ffbbd9103d21d3c3
z6ca934060e180a9c9f8f13cd85e78c893d4c02552f72c521c9ce12efaafc12d30ae34fa6842f29
z2903b9f5b5789bbbe9690b721be4f7f7c489592d68bc7edd936b82d0811fd310ba67bfb397b00b
zacc816b2a574cf731b1df2cc49944135e27cc1f0c3859731c5fbbb9748c77927614fa664ce4e94
z79729d51d869d1978e5988f35534e342770dd910fdc4115c7a6667aad8da2399b5f26d118a38c2
z40fc142265440a7d2278d4d4a4e0e4d1742ba09e42c0d2b5980e8cc405598d75696671cb2348a9
z5b288a603ca0e63e960457fbfca9a10e9d1020d5334d62a1e446d998973c6044458b42d904c015
zbc023e42c5a1fd0d14c963e20f65ab547f6707782dcc3a1e54a97584f22bb874982d3f8678c2e8
z0e45c2cee4769e29bf9bbb767be11b0792b3dd6dd047a3be1f23dcfb1b32e934a51ab675f4d978
z4dac483a0e91f7d407e82ec87eed12a3440577507f75a8c4bfdb6d4eca429e27bf5785ed94911a
z6ed7af825a7d6739e02a5c174be0eeb3975535528bbfe5555faea06935b7d1b54b3b9d858eb446
z095869abef6cc7da9ab086371fad228c1fb060a5d15fb3b5d4122a5b2f1c3ae830d477d3761192
zee95042d7ab6e9810a415279c2dc8bce01eb78cc0b862a65c4906e41ce3e72332d4520dd8c639c
z0ba289ebdbb225cbc6d2e6b3cbcb594ea8c49af41001010f07d22530f61c5e0c0a86c2115b2c01
zbcbfa8bf16ed0933cbddd62bbe96832ad19bb9a5e0e3159b1ddba24178db21576d75014819a7fb
z10656273f23f71e0a5c4e4d5355182c7ff56271a4ba55ef4ed52d771c3a14f757488bad3c97b0f
z6cf219db0a5f1a6f06b5cce69976e07c22c6e540cf3f11017a3baf1ffa0255e0e53e77f68a871d
zc447e20ef1bd669eb0a349bb43e84b0f2113f1712e447a67e11c6e63f4fdc585c375c188d38834
za6d41f0bf690924d811976722d02a14c2fb61d7f5428ca2701f849a8337fc89b24abd1cede99c9
z2710bd84855099237829a8250bd048f2ee5f1a2ab13c3b76b92729895d4fa72c2a1fc181860bd6
z4bffd29aa35782db0ec47a6f3c6b79438f22990e37bd9705e0fdd10b17b24ac39472f43a99d923
z508059c6188d0682545437b458492abafb23b22e7f21ad72cb6db7bb956040f032462f6c59a13b
z7c6853cdb3342d537e1ba3696b05c9c458c3beffd560f26accfa8cec3c55829c3dca5e7bf557c0
zd1352cb02270fdf61146341ffc878db66fb1942f73b562c9177602edd6100e1fcb08e044ea5108
z62f8813a25d72be86de9dac196ff86e87927dd7dcdae3bcdc87abbfe5d0ffb70632168778d65b5
zf8feade8e68e70297ba20012b34fed6a7083ea3ff139b8869af4a94c461df665ce58fc9fdb384f
ze1015ffe37603a50847ef91092ee012c4f513635c6a8d9ccaec4760552e9237839fd338fd9cb88
z4b943f8d6c34114f81b4a15e5049ad04a323b4d836f3ea4b4892c28a3f42aa10600757fb214603
zf3b1a5d85ba7adb2976cf244f00d2c7d21e10dc18579f155ce4c78f7242b53cf21e48d05b2ceab
z97dc8cd52c7552583f3d829472e9f1553554d72cf1764adaf7957c4872b7f54e77b8e5056ca92e
zf50bfb8ccea8dcabb80b24cd8641c84f2326a92fbfa245f7470d35dbfb40ce375408408bd37d12
zee5bc14a10c316f717afb8006e303059e0c5767a6d2aadce833035daa0f8efdcc8162e81828006
zdcd52d344d353737c542b4e5a82a3188ed4038019a0ac2feea7c4ec77d5e9a32efc5b3e2dc7f23
z9dd26046dc1ff42ae87fc8f7929866f0e8d56b9054984a1815fb8e8897e18bd5fd5b4a901abc4d
zd25c9e2366a089a98bfc6e56b3f6ae8c0dfeb6c72123bf99b9302bd700d2e678c4136cad79a5f9
z689601372a8d4d69799be29a1705a6aba5d5204078baf93c3e5f521478d35ce8110aa80a8ef13e
z8a1a538ab542cbca2d57803d1ef592ae236bd217b33e89a2ba93a3465cf6cd9366f2db2da9d522
z9ec79f3d00d6ef2cf1bef4ad51395b58a51d5feb87e827d2d051f86a0c4eea8e78158f693ce829
z4947b5bfbfc8bdf12711a8f2cefec205e5da868db088103db95c59b333ab485af0270a31b24261
z3c46911e9e089880c36effb911401d1b79d71ce78edbf33037b9ef4cf8d5dcd5dc91e7cdee0cd3
zae4a5293a02fcc4aad9beed356bf95dfaf88bc8fa06b33fd5c5f1baaa4ab3d0ff26320b258d0d5
z986f662416a0a4cbf03abd5b219eb56c5eda1b07be6d940c1b18b3cadc51675663f9d62a42b63b
zb2ab80fb30d607f99a3e4d9489af961a5d5d0f75dd9c71fc2726b8a0d4ca11adee7a1c90011f13
z415225e55669f825e9d766770a141876b3a3b34b957f77e8dda8990a4fdcb1cfc60da013614dd8
z0404c70928ee46f892fd207d36286d249ba1b1540963c3e2dc6e3112edffa3daacf4b38ac9ba72
z0a36845a87ba3cd6344de9fe48fad132e15ddf6d25c579bb930cf7fe7ff520e7bd5cc75d7c8311
ze0e40c5d9e6c43d4bde7a8971540ca202f30fed76a64f3a33f6e56d43fe8ff80795ad4fdc390c5
z0f9cf5d54934b61eced6bd5ab64ab70b79f47c48afca28b996bbd06211b7aa2d80d33ba02a4acb
z8a5f575e8a7a04220627e12a6fa69e716f252c0429716e4682ceee4e528a98e526f8ce4b2fcfbb
zed269a97aed175a370bf1b099c69f0f2435f3ea55aa8763dce150f463276fb86f0d2482712c10a
z77c792104c0fb7e0ec1d2d0d88346305aad6f39d186ded2d06087cd17c64e17faedc48cc037999
z1f2df571c4436f2c468d04b637a27eadabf862691e9a0da30d500724d875980e70341885c9f735
zbd9f993254a3740e37eff0a58806424c6764730aeff18eaba1eac74b5142be4639e618ee7bd65f
z0398571ef6cb36fa1734d8e18dc7be40becc32138ceaa7927f84f58a3d3e694e3ab37dfed9cde1
z05b40fd3d992bc44022a20cfb97a1ff7b5b7d8666b347d36eccd87a24a84c825644717955b8e71
z3b6957395d9c7e08c05c926b48b08a9cb86bf99ee4339b8bea3a85dde0322acec3a60ee58a584d
ze0d761f16eff0fb808f7834b2d2e08094105e84eaf5d5a2846d91c2f8f344d72661d3db95c9279
zd9d382f25a5682e52ebb4d18d9ae4dab7ab336b38e7efa24bd9f7bddbb46d4b55a1b28db314b13
ze7176aa8bfc8ce733c787278ff518a7a214706750949cc2ff40c18a78d2a46fe97046aa2b9e438
zc3e82c17c9e23a5e92f3cb947e6f3822abf6fc316fa179045a08b0c1875b4eac11b55fe5fa0ccb
z365b53a3bda12b26e3e9e8c1994b977e9a1883744dc5834f58fff90c9b571c060a4ab0b22d86f6
z8e12aac2edac4e9a60e3e53a0625f6a5a33f7a56331dfa14314fa317f523ac44a588cb1f8ad326
z600754a4192880ac12e2fd2be49a078c5de081d551dd6cf05e7fd87bfc818cc0a38beb8832cfda
z2d7b609a67fa077dadcac27f9cd8e9f9ebee6054378d57fcd789862be465709754c4acd4ae842a
z01dd1f5215bfbea01e8b8a1299ed7c110cbafff7376891afe210ac1738a4609f3681db9589e549
z906093a8fa1bde6243d9ee3bc6288adad15c612c0c5897dcc82b15b294a02d5efc6b3b3f5d41f9
zc6f4a54505e7652e617ec2e5074833fb57f9798ca010c7f9b42d06ba4875c946d7e3976c3ed6fd
z994db80dfb046374aeb66599684df9c9871deedf820c3db9e98a4729dbbba0236e329fb96939e0
z60cc0fa3ae93a85e5da5e341fbd47d8a391fbcefb078cb24af7488e2dd0ce7f987b1cc09f5a688
za6874babcbcc7380c1bc6f8ac37fe9aff2b87e097c068a3a70ffdc24b6b2932232c9196561d321
z65a76d0ed12a0f3f311beca91b21a3faa0a9f4c62654d917b960b8563be2d81a17e2bc9fc27b2e
z41467c4c5c0f26d57db08213f1b5473c240fadeb472271ab3430ef377d0b5959b64260388c9dbc
z8916b493ba4ab1612e8cb7a8b08c428a0a63ac4ebb04c664c732325407f3229ffa2a0dd47e8b1f
z4de6a576a3999f39c52cc2d58fd684a4c6fbdee6ce26d90362a6e95bbb932f63e714e4fc438542
z81f22242b6aaa0f4ea20e7b4bc57aad3c12380b9d3e82f85b6adca7a9d11f107d77fb1418989f6
zc8e342ff1a105877fd183380386ee4676f11da98989f65dfb8b2d87ede94bae38fadcafa1beb96
z63483b0a5d8bbbcf2f63ee6b16dbf0adfbfe5ecf02e1a91095562155faa40e5770951e555782ca
z740466431ed485993e6b6cb7cbc40a3d2b75bba08a45e7af26c428a1958780dd198d36208e604b
z651992a7d3cbb35fc9e41191747497aac63548489799580365aac9d37cd140fe8880b3d1f969e9
z7c7ef56e5cc5471484f7ab6ca9a879a763f9eea71a3e1888553fd75be7315b92c2dcd8712de7cc
z532da0e33d0ed3c87d31601fc08b51e6d4704771afbf92aebbb10a42ed163bdb703b9f2c02a7e5
z41adeb7d49ad46859496e0c28b55205f7a1577775e5dcc77044cfaaa8709b24b376de4cf9f9203
zee3e98793da2ca46cc095b88e8abeb71a412f8d37197426a361a8c892a2861a4452df2b0e478b7
z05dc28221353b412ae4f5426b258055d51366c62d5e93233177cd5e467ebaeebdc1d9bd30edcd8
z0d4c4f8aaa40c6b0f79096f37f0b1920b45298cdb4e43fe414b83cf217cc5f9e982f46a4973352
zb5228515ac15e964450c28676e67178f8e58f8130e1795003387061632e584bcbaa37c82c6d069
z87bda308820e01260821a668f486a875fbc6287f2fad55510b4947e75117e9d1f1e79f90a04c37
zc774027d6dea0a13cee6a73156f33366f30b9a0445a8751c16a09f82ee8f82add11512d486f1d4
z067fbcf8a583cf48bf62bbda3cd19eb996605cee663864552f25a141d4cdd3b5e97523e2558ffe
z11f70cad8f0c2e7e1e9603a390896b5c37b58edd177a3ecc5f75ea8f79fb51843a5b08cfc0682d
z6b8d62ac7edd1c7189c15f48565b0ce59d92b12b603f141fbdf137883e2418cdbf2b53aba9b33d
z9ba88a439cb051e7c1663bca2c1e09bd7bf491ff8c0afabf226d0913c6ee535a5fb31b4d2b23ff
zb1d3c33984a37b683ceea9fdf19bc07bb1a2d01a383b953faae069c4a3de4242a659c630194693
ze9bfd221cf8c888024b845ee9e454f7b7b571a617de7ee73ae5e1641e5d47835cb8e4ce3add612
z8709a507228dbab850eadf847f1a9dc689a5a256931fefe77ae647aa69412a086e995354377924
zcc6a8db11c3b841d7f85b74b546ed15a526c8a0bcfda18b37da7f9564c8dbb4028e697beb66811
z78e5f02303f4b1300ec1ac4625e3f5f0a369ed5008432d9a62f950434d03b91ca829ff8b44c8d1
zfc2fb66de3ab2be6a51a1451f11177e341e990615c7b4fd5e450a5696ed9ed63298d2c726232ff
z1d0eac1fd61dae5d2615e02ad3e84301f212ab9bf1acd085f973169ba407a2a4ae01288e53d7a3
z24062befb1b77158ad245b965efa4d1d3939278ae45436171fe24d0e8761630748db4e9f678bf8
z941ec7ea2d026b8efe58eba3688ab94328fa64a5cbc8a4f8936d584139ee3e2f50d26b46c52fff
z7a0123b3866bc071ff279f03a3b6686fd254e83feeb5aa98c8d2cafbc2a8d980e791ba01272cd0
z6050488e4a9ed964459f91882b820b379b07a441ad406d35ca04dad288e2debf8e1bde104d7c50
z7ad5b1596e8873fe0b11499933f13bf2d6abfc7ac7d9084311a0c37395946e13cc35e69ca413cf
z75ba91f5f9cec1c383eb8a98378bae14010c19c44055e47483525d5eb8e8aed574cf54f0a40615
z334915f9f74197be51500e87c5bf4d41737d9dd9e398f656a3efd459f13084de67e2c293e601a3
z67f37f155ecb67c438599c37f1b5ab6b3e88d748f2d54ea7b335ecd7b37fa03906c70c6862e893
zf32a069cb0c61f4d3ed743abf51712593a5ddd5c344d6a2eb661c36e5609cf48e3a4de124b4370
zb4625a2c447587af8921b5d072579c399184e6bc5d4de69246e6051f83c4204f70ca1dcf8ea6da
z2e2f2410b063f84ce72937e60dfe5dba2a728684f59614770491acfd26afcbb7259ab5297ccd25
z2227fb2b3c2ef0cafe04a8fd4242ec014abbb7a222235714e02b1010b6753072ca9f2dce28534d
zb29c8008cb3a7ce3b0d33da31012d9ba8f8123521d11871c12259b6a28cfe5b721bde91fd9a858
z3a488540526b8b8da4e8bbf7515a01ecde0e12a25e7821ba8667243c5bdb0f18344dffd26f05f2
z69a766162d405171f14bba77416bf9c0a635a02993e2a9876b14b8fa784f85da9367aead81f012
zaf46b6bc7147a5f6fe88ba49ce24ae5c684a7bdc5f6ab330ad68d5790011c009e6cad7ba3aeffd
zd8efe1e9aa4b5d4918dd337f3aab64880e1ef8a1139d2b291a9023c275eae907451d2234a7697b
z371cc5bb910f16de83494380efd4c8f1439b620648fd44380474ee386f68028397e025b18a1305
z560762456fc385ca44a2a72e0928995ca4db88287cb27c887ce6e9df354d82c478ac3e0ca2bcd6
z59e1b140189127497c1eea99509ce287f7433699f75713414295a2d8c8d2be906bb70e9e4c5cd5
z3b6c2b8d13fcd675cef074a93dfd740a490c253f4f1772c190423f1c34c921797ed7463f6d44d8
zb5a9cc5224a663696591993b58799e42a53885c70a5dac56614eb88961a9ff7bafe51ea8573018
z8ba5d3678b273fc9a25adb470b9d34df2e7ed2eb4e90d476b428565922773df734b3b8e858e5d7
zc91ab67df5c99c1c33b59a9b0cd9e5c035c91c24d930e42ec4ee2bbcd79bdc20d533157ecb2de3
z8024bfd3cb911f050c544a260692bf31753c83f8496e369f929a890da2b0f9ab6ab0db3b956957
z77857172874e9993794af29257dc0afc48655234f3a4e4e924070003c7b2b5a0237ed6396626b1
z7302f0af8fff1a3e6e7602183345c88fb9903da32983c57c72f117e66360217a3c8ff7be72db01
zf81f5518869011274d645b9d0f4a1e1897201b226794c43c2732eb786fef844ef1622bef164a12
z69649c1b686cabcb27d486aa43a6a0ed16cfede0caff4785b8139441a1da957f4068efb21699af
z22b3c8de0852b4860a98b469b94780d14777b642bf2fe0b541e049a964645f68ee9b3217e5f21e
z29f12168b855aef9b986eca6a3a65b0cbe773179d1287e2b5110e0651e95266e3518078754b59d
zdcd96829f929620374f1f6f23d19d84c83ba2e46b0048748140852d4fdbeedcb2f1c0fd7fffcaf
zcc2ef71f307fda927e40b3642afb286dc990a078b2544013247ae7312ff543d5c8c91e3c00b4d4
zb651774ad4e65472a0128f2ab4cba053288a52e19b835056cad108ae78701d654b0b5143bf74ae
z77ceb04cd34fd330fea12a39160983ecf6e5644c5e3ae6a3c9c783f73229fbdfd4273258b1bc72
z0eac3ccfa375bc4827c34129edd5b2f238d84d8a3881cffb57681e3462245461fb4729e1436a63
zddc70227c7eec90d18622e50f8e2685b98a5d8df67c1d891fecf33fa04aaa76c6cd4807529620b
z289c082dda3fbc29d1ab2c9f19879d150b6de4711f3c186ac14b23113bd8276e56d7e4296ba373
zf216154f9afde10be9e028690ec3d6d565145c27efdf1876c3b16a61f4f08985400256b0d22498
z8faba8786bfe4787f74ce8790a93c8cdb8f30d53defe3ee183fea12269359e9b3d04054a51b708
z1c4ae827ba023b1cc1ee448cf8452b381e3436e1fbc8c41f92ddacda61b37ef83bc4427c3cc96a
zf3eaee55b1f540bcf3829a629f7b0886ea92a8515f9d3663006ff8579844adf59162b0c6b267fb
z7d37472d004ac5a1d4c357f1adea5775fd392509417bfee8ae35d6f482acb8d2d61b0c2c42c499
z0f30be8b0e8e2e09734b0b93d3434583652f27610ba230c97655cec803594f53c576582567b5fb
z285535110f7840d9a3fda00a85b829abef1573a57f3353046eaa34406bd8cca8044b95bb66ce18
z9959f5e71078705391ba130db96b98809d124819296b536cabc5969197a4eea9a950c569197e0a
z2c7d2d8bf050207ec4dcd5063959c2e8c48751d3eb17e2f7ca73a645b179c59629c608c3aa1867
zfe0159889a708c0c15fddc264e7753e1b81f46b821572128e11d8198072f735ce1a346ba71c48d
z60d474ada0b2daf6ef50ee5034d308200b3ccfcc9be47b7a22dfcbe45d1497e2769ef847586356
z087648929606b38f8096fc398922aeb4a9d682ef3449d09e66ef5f5b3eb9fb8b37792fb6dd2497
z2bafee0c5820f6d7473daa45980e61890663d19c087ee517b36c28b5cd2bad16f3a68b5446f6b5
zc8aa30b284581e1a1bbe19bac4db74e778581cff7011a07b67830157fd5584e6d52a1df098c3a8
z206feb75f924f9668668dd2101f1078489f429abb27af0faba82e09202adebf257ad669974d100
z599043777710c83acf0776b7779f2e3e80e0bb8c71132f63b9d7dd391e4ba80f38f23c9fa57a07
zec0269ef8686e95aebe2dd7e9c3d8ee1873becf18fdeaaf770ec0bef486c0372d145be825abc82
zcafb355c1d305c6130b4d6bcc11bc4c1bf14fb15fe0ac43bcafcfda615062632de7a2ddcce7ce2
zce1055a4be78d7cb11541bb5b930b834c1f8f149d47b089725c01672449d8cf2f6c5daa066a694
z2b2d3815c0f038047946e784914c1fefc12ef828c7f0779f8c3b02d93532c4df59926ef7505f26
z20aaf23271d97c565f64ba4c59f3201f613223769934daacb234d80f1f4be3b9a4f9b526519019
zaec60c95aa36e67ec06e6daff696240210d2d19629c1f4c56a3301d60162ed4112d25d13ea1a3a
z762a67441beb173861937fd0024cbccc1d4538e24f8fa46eb552cf3c2096a2fdf517f41ad71998
zec02d5d4b8d2e65fbcb1f89fc0405090fcc2e9e0c34045d832b838a33f0386a6d1f3e117a787ae
z06a8d9a2f8359033857ed39efe73a6ab04fdf96d61ff481c55da1643f0a4bdf2644f6f1321e91a
zec4229c4921f5f77d75d25172fb382f1df622ea17d1681c93d1c608629896924d938ace54951ff
z29a87377a75d98ff59892e5a448e28dc1461b71493a5ef840574dbc6c01c91658fa36d79ff12c8
zf2593736f801320c66bca2d3ff9973d7b1f2a195ce8f27b47465927dae09412401851b7858b83e
zeb0c2fdd96155e5a9b570d9944b6ecd1f3ec39e6df84854e0645583ae6f5e7201531e30eb61fa7
z80499592eb3059aa6ca51b394ce96835f7b348355d6ff7617ef64cf99cc7fcd6c161356be8a950
z143efd80944bc3e377037ffe39c1ec1f4ec48fa6baf96d08c6455e8f453c273a528f0dfa8a5825
z8b61d5adb07a97b80392166f38321ac9ca1558bc2c4f8b2b0048d0bcdb8e7b9a25d84baba05eb7
z69ccadaee21d8ee3eef7ffd7e1f1f60f1916312cd3f179a865dd0f5c23e3332e5ea046a726fcd2
zeb85abd8168ddaa548e7134d3dc1403f63eb0a2e11baa826f775fa252c657d221891e0119daa6b
ze22f38da374d403284c5c50745d57344a72bc6824e69fb7c904acd5ca99462e1ced785e78ae3a2
z9108ea07f900a12d97379e5d152aaa62997c638b1f6694254b2c18e246d1d93b8e25afc8114526
zccf2c42395ccb134ee5b54a05e8b92304e1ed45d6502d32a0d8464e7db6793308acfc1c7e82b04
ze4d6ee3b6527c8a5c241cdc19618c374ff81407883a09d3d76bf4086b05055c3740a4360fbc1e5
z7446d8d287d893b1ca8cfc73aff5bf779ab559840c93840ea20dc7afed7b08c8ababf784f1fb6c
z5e7eb96e02c561dedd32e781c0e17adbffab0aab437a61fb642d969a4429b85a6bf34a42f4acd0
zf2140deda432158489e442e4207bd1227192ac599560fa179e339dd7abbe94d361ef4e100c06a1
z7609d54c00273d0ef231e9d42c7628e0972431b8a76f11a1c4ce641eab633e4c4288be2cebb3c6
z45a5883ffa6d01dc0bd399e760c624931f41237ff55da83dbf405530c4eb46e8e64d1ca09816b1
zc16f6ca810601e915a539592c4f56038ae7d352b20bf7fc37bbc35eb9b8306b30224c9da2b6ca3
z3e79e641a9f5c1f0bd70529c6bdabd5adfe1e9f59c334e381e4d74870055f728b67ab69b7e7e9a
zfb93acf8ed8d4ef4f74604f25f8b8b5e5bbb8292576dcec790d0f840862182bac7b7d9cbb2fc6e
ze5a88fcd6b40294142282af11625cccdefc44940c43cf622857ea8f8acd6749da53f44f1ac280f
z8291b08e3a3c68cdecac8b376b5e17717ef4b3389260e055b595d676379cca63e748a6443e23f9
z115459d009f6012bc934984c28eef6ea5a19b6705841ebf2932af7ea02d337742afce50a839ec6
z84982c05a25d9a28ad1daef0ee2597fbbd1709411a15725b012bf67c5aab7760d501915a2dfaa7
zc865563824c12e58d8a7b682556abd58dd641bf372910a6ff24ab5eb63a3a4ac52c84723040465
z472a3e2ba6b008f0a3c62eaf303a7ac1cd0b406a49f4a5db79c26d9f53daa0884be371a55d2c50
z9b5187d2e27ab6d036ac0211aa456fd39ef473a9dededa38c93361229e050fbd1376b66a3b75ae
zcca2b81ec6bc1d39e37a67785693388417fc229acafe7384ce89fa6cffab15323bea5b1e2df114
z4356dcd2ab5c74baa64d48eebf4b863b501d325c6fd7f7d7ef6c42bb7b067d37b7489ed6b89bbb
z4c736b5135995231c8c4a7fd20ecb99afba644f9845432c96ff3ae82c25b3914b7af1de7e82dba
zd0ecf406f5862acf094d6fd442258483f6da12d7fa23846e634ef9823b616b3d385908c10f7c84
zb30ffc1841e7d9d1194063b3f4df341e51402f0d4398e50904e4a82b9f36b9a748299ae6191852
z171a1877db5bce3722314e1878bc853d48dc9069018eb5b2e72e45ff79020dc0e311eae572cd44
zeb4bb4deea3486e55b6a2d62544590747b33d0f3d2831484b02831a3d154ba04e3f70562b2d3dd
z5335a1177e34d45b06f8d13ddaeaf2a962c8a554457c596c53bf9bb131dbb624953966004267a9
z6070dce6e8b7a00f58e28d4287fcd02893f0f603491cb423e4ef083e2215d4608c3dec90c08ebe
z26a131f299f628a8afae1f468964586602db9aca05596d6b9ece03ae07962d23b77d86f44c46ba
zaa367f90c24aaa0363ff4b16699b7e881ffcf3004bc68b717d5cf43ec5db2d9522ad217d243e26
zb0726e28d8eb4fec8be27a68bbf2ef2fe810fd310e9dbb638529812f9e91571ed5d3364c84fbbc
z8180eb7b58f920aa8c71477c46339fd28f1418d4d01db9e8a41e95cf4eae515f74c830f9035042
zf108a0601db781fbd24795865e497e819034e7eac42755cbe6755717bcca1a2114c6fef39df79b
z23ef81c53db6e08214085ccea83c88e2d0ce35c4aeafd9bf17d697f78c15d3945ed9cd6b2f20c8
z68977e43dcc8145294173d6749897dc72d940b0696a10b72e4eb3730775c6963e01aee8f453d16
z3a3074780dfeb80218b2cf6a904e2781621ceec6f2f64cbdafd590f1c3e7c5f2f9e4b70389e116
z120ff027c12184f26ddc16477c34e9b105af862706588c5078e9ba8bcc7d4d112be58e7db5f55d
z70bcd15b6407716977b86b4428406cda5b162088d614a5f470df47e79d9b54ce4e4a7c545d01cd
z2be22a9d6014ba2de6465eaf704b5671b84a01f5e01b3313f38b09b42da6f7cc49fe22f5c614aa
zf66f0ef48e13b230cb6e818b269fe6ad2cdc90b4efac37a0198562b615c04492cd7a1588eeb745
z2ec13e81301d62bd343ecda3701f4c44d1205eb995b31ffaddc1ace79d4147f35b73fc0c5d9d91
z3d5e91551688c676ab92a58e88363943bbc4dc80bc4529589080a932cbf4e6e7913f8fe8586080
zd2c42e428bb7e71e1a9bc71f4553a9d95b291a65a3afd23a582602c19e4ee7c5e3adca92d6cc08
ze6db90b8c9ca828a7deecaf605e13591b140e78ef185a5d6867a82c8102aceebc3d90790605c70
z7c4158e45f71671378a71ba11c3b07a7108b5a2d04d482f31718f295a389973cfef5622f913124
z71c28c7cc39711cf04741cb215fcf0eb71d2e89f1868b0e5e5a99dbf0d8393e29d93b6744daeee
z7e622b6e6043018509f194974c6753958ffe5d2020ad494413f7f96a6a84d079220dab58baab04
z969b76235ad94f635ba91b1d60ecd20afb9f7e129380fd5fb2ca3951bd04235279c622ea69b557
zc3fcb698f7d417da38a9b4581318f19ecfe724d67b084fe2d1a0b847aac8bfea92d9ac75c30ac1
z21b8498fad3c5da5799b855c1a8b11f22a236567567cd989597881461d08b19c9da2a739e55483
z2a73828e094cf45a85a77904295d82c8961e4ab218afa3f5827534c12b82929765487c526b0a15
zfdd23f7fe75868a36e655257ab4e3e7b0477b751b13bd4024dd1146003f3502b474f15bd726168
zb30815c04f619fc1645418a4c3b9378e7f6ab34cca18aba2091070a6dc4ca815b5241391ed9060
zc46f229020eebfdfe02f836560b5ee5fd3c596c0f1bcf2a8c9fa5d53435f6a3f14d6a14ecc412f
z88a7fced74b2fb8ba5eeb3d2d0d2aeff24e9e0f312011dbc2b50279613d1c3ac8606163fcc9c06
zd32605e7690509768f3017470e2af48091994c1b88c64a172d0ae11665244b191d3743f1d3c021
zdd030915cf846e3c0f687a163b7d497ed39c56ca7b3e60cc5b125a5276d35b08e30e651e36472c
z064cdd6959fe3ce6f828e480228c58a1c3ca2a376c3b85e054ccc635f1bf14532f79dabc3fbcfb
zcf63b6fbf64c0e8f663db4b3c05a828edd2d509ca82fee00d72a99120a6cc5e5cb6fa083cd6755
z9cdad4ed01d5dd8ad7d015d1516a66891ec2323d24401b173ad91a7b258265b2da395b28859cf0
z4c5978baf67c138dcdfccfa1681ba4fd03cd05c8eed9fdf4b5c8da7c7e760e35f5b94477dfad97
za8c8590a048a39fea2866a9eca5405a553da899525fa143e293c80447d5d2370ea371a2dfa5d8b
zeb6d533d1b048242bffece55d4ca1700d8a1c5f0dda40f91a842640ed0f57e55979f451d40a632
ze15e91e7803d466f8a57e3321f902fe6a8c89f3bf587bcb36eca427b8bf059a2a2430449c34ff5
z7a8fe4abe0a36284e1a37dad8773828cd24c484179d37a1d961f6d339d61b7cf7871a2815c0638
z3b9b44db76c20cd7a88fe1e8112df842af1e85d2757a11e103b5656b28a9a5c1dee196b5779ad3
z9a4e06f8678992ebcbe2d32cb1949d16bef1f971a8ff75696c8729e88d3c111009c9be2fff8e0f
z9fdbfa4d0bc1ca6cc78d43d435dad92e61667167722e7348d011310cbae7c5061054314adb398d
zce2b465d12984129809794e25628ac084924fe7bf5348ef3d44e743ec7c87b9ff20ee7dbde6d69
z070984c8dabad0ecb5cd2c5d7771b0c82beeebe35eb581ec8c6fec06051d4c31913f2a78be402b
zd9141ec5a65d5816e58b2320f6e8fbd0ee3e5c583f7c67e7a13a738b833f430d7e3dfe6674cb8f
zc271b0f32e864dd4e9ba018bc7cdf0e02f20da25a77ae9d0b5bf712c235898cf84ea17b7ccc2e8
z36a312588b834ede4aed6b6e807f59c10df669eae57af7ad65e7943849b2f751f8c998df1f8c20
zcd8d15109f76163091d0b1fb9a628557f1572ec1191946e18da2f8e1f7f8809f99169e8002a367
ze1baba43e0951e7ebdb9a1705d13ae38d44eb834dcd575f05d1d99adf3014b4d6b68933bc2743e
zdb894475c746f6a1fdeec74847e3ae20e9b4e404e2fe0787c2e5e73289a8108181712aff378ab9
za19272ea48b185a6193ca7c74eca851a854cf905a131d620898730df2f1ecefb9482498ed72c59
z004ee7d345c0335c213149be3ee0af243167486635971a6a43ee3bd66c3568089b8a7c37e86261
z45710b40fde42456e29ae1801c27b36835b775360193bbdbcab51ef0f1a4d44a8addd800df26a9
zed5793fd1abc45ddbd3a6772230b2d3d5090ce89c490cd839fe0ef3c72061ef45a17c5b2134627
z4dc1f20e3dc22d0221834cd07ce484c12aac638ff9ac9aad65e444fd01bd7e8180105689061715
zecc66c4dc4f9361b82a1a0c8f91768dec2d36abf098e706795c1b10058011a1e1f90af8f6b806a
z1a9e4ef4e86cefda938379dc9b427350b2c5d73efeb969a414c192415ddd45386fe0dd9fb8871d
z5f977f98da191830ec88d74114cc72eea4ccac3194fb67100e5ed5fb19a405c10cddec155c5bd5
z384abd930e6eb9347bb2f7749c329f0151033ba5a3e75e0c3cc09583d7613d1ff6bb33de14d514
z855da48623c325c2c2691e3db00f07fb775e03459266a4249e69f36a6615bd561199eb56c5c309
z91cda6dac77d68bcba425fb22a3b011935f2573b882a5f4e8590bd3c06d2e7c9dd278b19464075
z4454fcdd964d58e1274a1a0c228c906d709fa2d4b5fa2cc92fd696affbc33ca91b23adf97b1d31
z56dd075e9a2e303255ce2b31d999bbc8eec7d6961df1ea42e240847c4f2d0caef81bd7d9d618e2
z1aa9940dec9ce61beeede1375a0537a58fee854e9458f940790cc02218fea20fe4ae81457b1ebe
z9fbbde6f7c557b4e198d5924d6d8bb8be35f51679898e1d45649a78c86db46557ddec31278e88b
z5668654d7cc15d6262b4cecc0f1173d6751e1351ee636b40b503d921c4675b4a8709114ca62021
za3c0b02b3c54578ef0067bb3d68e4b952be643e7859791c4f7e7f407aa7d0a6a89f745888d7543
z71d0325196150f77a81359e7727662949454f16f4c81a3d7e937378e197a4309d04e572d2054c6
zc917fca5c58fd66ed2af36a1d0d9092b6739afa1f9969be6dc521eb248e6421225a78fd101100d
ze084b64b3e5a20f9d2a4d335f7c0894164f8d294790cb4db380929be8e105edb46c7823c69c1a0
z5038906c080e14aba185d101d4086e405f5b30a3d56102171773a7b97ac3bc5dd9df17c814a6a2
zf43da363be3965e2562145f6a2c6fcf0c8f62eda2001e9e4c51f47a6b06b9b9d2871bbbf3717e8
zc9fa660e08b65e4ba5d44fdfba29bcec3c63b188e4aa3641907c4e491dd002be8e7f47299d648c
z8849b84e43ab9a631ce584c57657eba34d8df3c7aa36da5dce07f13e7eef8b07fe8661f63b6559
z1c897619d5434ce8cf8ea7f279f07f6b6b83debceed207f4fffbed292ba20ff856e1341a5f7442
z6d32f61834d952aa83dae9f09699d45fc737f1e1c87a955436fff49eb102b44d77ab49d17a0d5a
z630b5b003b96da0108c8f62991230fe5b9f90f86a74fae686957d66867dbb9780ed9690d338535
z63a4a111e60096e8063fb682773b28cec41ee6f000c1317d929afde3fb9b1919537e90f13ac1cc
z24bbd1e1882ff91994486aed3ff2e94a969743ac54b0f7093590e64c91ec64b2fc2acff5d62e16
z3239bf8b1c4266d5d478f7fa7dd54d873d4818d8e5195053da4e229b88ce4052790a5f223d1e7d
z319553d11efcebcd6dbccfc3395f744520568dc03e95fb6fece73c9fafe34393d785edc574e96f
zfb67df193a68a733aaa148638fdb6652ece5f1a23f0bdf96da5a5b9199da53c5c2f849a1acc538
zc7b14cee5ce9f85927a8cce28391d70578e4d313e95f6d779f34cc00f9c8a33b3812bde7ea083d
z1214947d7b8cbf86ed202fc5ff2ac0fe42b0959ae974fe1f24b3bf0f17c15b56be4fd4b5a3136a
z001cafec0c1ccff528efb84efb72d38dc26c23ccfb79aa93a5c06f1f5a9d9ffda3c8e8278dfce1
zf24de89420eae5d3ddc045cefffac3d186cef437c6446f2e1d0f2adf77541ada5d924ff64a0e81
z523b752192c7e8d9acf332c0d87c2d5d459a23af54f36df7f2bd940915f2f113945e46bb07422a
zb2f2eb53aeb76e38224ac9ec145d272beae011baffd8fc2e995f2ed6c36dc46250ad80d2a31ccf
z3513d1cc7f9f4a67c4ea6ae7655abee702a10253ba4f4043e03a1ebbf1adeb4c80f0f06d28587f
zd232eb8de7578c35899b8c060592b605006b0b2e14d39fb2c2835d7526cb6c5aeb4fab0106d10a
z5317f493a4802402a9b9a3bef548e224e8a8d3b7fb640f8aa10e945ce0247510ab72f65fbaea50
z29851b11dbda7a279faf9c955a8c0dc3088c9dd1e7a63f2cb82ae5354803e2323565b8d3d05a37
zb494d3a019e543dca4825fc3e1b04d273f7c5c67068cd5b992b83bee31e6aac411a5d3b133b88e
z47e44378307248a04f89ded71ba82aab214c3a8a5f4cd8f5da1a08136c649da8b8a7e421804a2e
z5d353285e85ee39a9227ca3ff1da30866db71d145925e54371728312417945904a2854ca9822c6
zb7d544cda5a746b0dde8a57f9f3ea75b681ac5f0812a062b29e31577d787fc8e2721a8004a9251
z28a6795adbc1b4517de2901e4abd36cdf457e29c42553df201e29f22d4e5dfc697b4f0cb7bb4b1
zdd2e3003f774fde3603ca4167e82ea9fe312bc06e5aab68bfeb596fe94a46d7eb72b14b294616e
zc50f15acc796de31a73d61aa7895c14daccf04042b125943e31185ef106891e0f34d6815040d9d
z1095983012d4020ca9adc7b1e11cee5753e9719c435cfa85cfce5294f5d99fdb37279f482d0de7
z8b4bfcb9d116b0cad72472051b33ed5556daca000f90dd7ea4f194bc2193262684428b08ffcc28
z5ec5b9099390d5d75be3fc1f359762a660f6ff7e999ffd3247437db0213a1bf4c46c2be35e97aa
zb839725f30eed899608d85574041181ee79b658f31084c8b5d11e14756748848bdd180611088b4
z9db3a0d49d2944e38ca3cf194394e5aad94be3c0b96835686357c4d1c95997cf9a8887217fb94b
ze1d003c91563ae65effacc168e66ff0a7797352b2a155d765654e8dd136513c36b863bcc952087
z32940eaec27fa390a82a0373ed4c0fff4a894d1bc974b0be57922176d3a887aa566680b21fe4d6
za3b849789fb88faf63195383714a85f277095fc24ab2e17082695a73d5408b6db86aace126210a
zbd963a810a8f9a63b1b1c0bf67728ba428f04abd700c3223e9fac439db5f3db83b7931654c5237
z16a1090419da2ad5a1349ff54078389208a43c80a7ea9ab7d8e6595b6f11f65c6f60cfdbb82de1
z68ffdaa23f945fae81a6697357c6358039acc3469abebf75991423e58c3656c088aa4ca22f866d
zf1f681878a1be5d86fb62eadc161507d51d8325cb1db6d8a17ade869958cb57e605337315c041e
ze71a39ea633e7328111f83dc7a5c286287aefbf66022481d0721ff3c414da1ac7d768938de94ba
z9323b338405ca124b08d2cc8aab9f7d35d1a4eac8c5873ff0d23add1aaff6140ed5a916633d0bc
z0bd4793f5d749d1880f5766906bbe22200233b68eb6b020008834bda569e7c600cf6a9464fc4d8
zdd62e85a8d19f4b702456884e7b56a672b7fd7306cd38159a82ea78ecaace568e8228e0de4d96d
z9ebc6268d38bf8f9dffd1e7796aca7f82ee171b966ba5bb6368a3c50f7e01c65344ac5619080b6
z3f7c6fd408361173ca5c3211168d2b97a3dc99c694e246882fc58f9938f9b82663724b4b500436
z012515d1bcc8a1ba7f616f4bd980edcf6c834deff0ef7efb9550e801ff605608824dfa35bce6da
z1b4601f8a900360ee3e1b4b639b96b5d820244af96f0a431ab74a98208ad4e826066d89ff772ae
z49f8b1678c432d63cd2eb778c245694fffa58fda869063b345ab99b5c3e9c28e9ce7623c553010
zb0ae4e6ee1d182ec28e43bcad7ea68b29c8e0857156c42cbe433295b7ade5abac6b271f4a02cb7
z5e42d4ee5502d95e0c4a4ad4458a7c85da4d1d23730351135c2975f93806610d0e54fb8d1f17f6
z4f0ac3db74984aa6fb6c96f1e7cea91635a35103b76785a3f1bd1faf17a3600596ba161ec27210
z8c7472115ad4c4998cb6a973fad39b43ee19fddfd1e3f9d423ed088a9e3b1559aa07f61e9d50f0
z39666c7e484502b359fd5997e8a260c18ef221ccb36298d40d53766847a25af980c4948380ab64
zc3db6267d10b1b50724ad902aa53a83762def8d581701913c2c67ec5f171bdff2100944345bbdf
z8943250164d2dc099a6183eabe1975468dfe52f1298e4515935d66caf3b6f8a2d0ac9feb0a664a
zbf86be51751615e7f1c9d14eeb59d860f45673a7f7d81d3609dc24ea37b65a598d5c494ca0b707
ze77d4d69782efc57fd2f7223768aa42cd55a0f6444d7d220265a6773185aa0e996137732bca994
z0af5c5be2fc2b92c88f5a2f56615ab4efd0f7a6a9596c4e1703e7e9cd8dba3d30ccd044572ca67
zf3100952ef6a29cda0fa8115e5992d1b5509269725238602baaf78def36894ce611cb29ea4b36d
z2b676bc07561322cb20d1b34c1104a5b970c2f18087b7a446cfab9b1742dfbd155291a3d555d93
z9fdab2e18cbfe9c5ca2994b2efaccecd6cad2c7d15aa3ffb6b8c14544c0a136d0f90ca1430709d
zad5107c0300f9a7f9c29e61a2cb410d30056c7b8764057f07b2ec180037ac2f83d374b85d8c3e0
z71d75ea26bb331accf929279db1e4aebe2b5f6209b2e7e9b21aaccffd6acf26d6f57d9f5a57567
za81df14b6987361aa101be1d17d77dc808bb093c5b76f29691d0d516c5bfa53e520b22c7cd79c2
z2aad4d48d9025b3134bc359fe8212db09a94472d61524eff9c53006255dad75534580230c84677
ze19064fe8122521dbc6ea6d80dfa120143d796057c5efc43e4cf2ce1317e70b5c4c838855d8b24
z7d82490c77eea56b2499ae8f3b64cadd5a95322d3871e144108b6b7fe3114a97d21c9974856480
z60a5a62345f5e6ddde032c44c8f042340b7ccd068adb986015064c5811b13b3eac286c85610e8e
z2d1f54f17c18e36c9ccb28dab728018ad29ffe3f69ffe7a4e81a33aab8603a2c3d8e70494f6203
zecf44a86970dd2cea79ceee4b83261f799d7817a8bdf213325a85c16e4b02877ba0ef49ced210a
zb4e4f76cf98c6749b61587f7de910275fbce33e2304516caa4e3cc7bd6ad1c5f84e6b9f8df0ee9
z3a6b9cafac01adcea6e0d83148fa0e0f4558f803aeafc521dc9190cd14b9fffed1aedee2bfafe2
zffef5b87e6e7f49b4591aa3d5cf3f8b951691def8c095520d8bd17fd13fce545d64368f32f56bc
zc637ae015f0aa062a8c7412ac0b6e525e52df0d3027f2def082279cc18f6af316bea3e9ee964cb
z1eab52fdcab762474f456eddd3f39948ea5fb938bd58276902c90302ac2fbe7d81e6f9ee50c968
z600400ce2b5a5faa99e98ed68d72161a16aca52ef40a653a8f5d7de14a35d3aedc1aa12ff1a011
ze76a2ccaca22bf62c3f941941c19d6cc8bb4d3d2e203285690546cfdaf190e5c8f08869feb1b54
z929490f7e01edd63a32502dd3b99840863d7aa23682f73e76ba9141dd530e74d124822e821b2fd
z57db719091eafa6902e5dccbc051932b69e171bd293d1ae7739421dcb996a85c0f916a9ceb594e
z8f3ef889b8d0c318b653df58590c4049e6f516d10be0141a0f234c24c063389059dd4c0e94adb3
z91debcb4f57bc83dc56cf44daf61cdd3629b1dbb3abe555b319cfc2a548064eac48190bf1241b5
z6e2c96f692e7605e7d11d5fce87109e4e5de6cb63e21ac52db50bd01e7c9e1610d863b53a222b1
z08b22a920c356073bee89da5b996de77a1a71f275eaf788af01fc23adfd88714772e462714794b
zec712c5b6d7be69f13677f6ec21e8ea2d0c38d2d0533755885bf3b3315e43d01a4ef4d7cfad76f
z6e2842338fea6d84f5d53377ee0b01645807920c2abfee2f927f768fca7138f5f5f660ca061b79
z78f7b9a919f353567b5c1cf1c9d0b73581ccb437d4f71486d45455e51d091bbad56fd2339d76ce
z5fe2b446cce453646eca9b72516702cab01018862231a570e0fe3ba406d53903e0c6c74ffca91e
zc954e3893c19418da556671d9666f6950560853a08e8043bc8705d0c6e606b3d5542075440a320
zcc63590942ec26e7eee2477bc040828af5bfa1d74534eb86c6aab4a6639e627f8189edf51b8570
zc6333c9a4758faeb70ccd629d66eeba557937fdb2e0387a96d77a990f93e4b2c125d067297e5ec
z49a7641543d59e18c0fbbce3979d8382e96d70fc39940ba6981b850c7cde54395cc4f6e67c8294
zad2b4807ecedfca2a5f9cd6338df8e96523e23953ec43a09d885a4348e0e9eb4a97a40c14f7327
z3644d07b18254bee346cbb16471fc779673186fcc405404d3320254e5b1ecc43173455875c1083
z8c3c8563d29c064640e258e88bf687f554bfe61082c73c9d04002f7f9fa5da81edfa56997369b6
z39ce22bf96e03a8892a81feec890cbad486bc5ac88557592354b2078545083ef94880dd4740a0e
zbbaa50a84cb5da9f654255cba3a3a65cdf6da492c8a0738dfbc4cf283eb83ac844ddd95f200ec0
z35d27b9e8e9768dbbbad1cef45f27a594c842ccf36c8a0d46554b276d43fbbad74fad69e7ab654
z99f77c2e10497cbabdbc8b886dcc1dbb96257cefae82c0331b7f0c3fd214e752747d387c97d2b2
zf9817fc98f94f386c5ad1d1399bd18ec0bf950b421e8311609b6568aa540256045f54b28405ae7
z9b6417b8b2b9365e4bde3d32784680b19a06981399c09675a59556650c6b978fd0d4c6e54ffe78
z92c4c8ea8ff131eb06076668f40b361f43ef1d0658c56f2cee95341389cbc6a18284b51e39a181
z559b8e242f45b3d2e215168bc7bf3410165ab7313f291704cd4bddacf7048599c29c9d6b504e9b
zcbab089d73a77ab8d1961b295a2a29c50d3333d270e6c2116e4a8b815b8be2a707fad462b439ad
z9e72c16f86d861435093d110c058cccc85511ad83ff5d26b9ad31351d8f0a138b511cf97a67a28
zcee32594e3f9279081eda3b170d8d243429533971c751ffa384a57f363e0fbbe686593516b4956
z6c9a81a6c28bb57b96a8e92eb9c77234e1914e209977c13b4a91611dafd9caa17a7a48397216ae
zf5b0f8a95f065580d4fb666c226498e112b739f0c372bc5ada9f7de6c38003e33a7eb7c977486f
zdfde86de7d46e90c01ff07987636da2c62a572efd9aae9f8432915fcb28530297f05d416e168d5
z2a91f8556775d4cbc4922e7d1106cc120875c3ad0909df79bae26e7a50edc4effdf6a0d6daf2e0
z1bc13e0ab7bf5b9c63016512d1e2b99f346cf8b23963d447212909e1cb535cc2aea5e565f339ad
zb8e8e3b569d59fc5c0c5f133d8e871987c0c0faef6791dc7d756c6da63ffa2112a04af91577c3e
zf4e3d9d8ffbad1bc5a47f247c4cee703fded85e637a4458206617fce3f47cb8fde8d06f8f58131
z072590b05d66fdab263e3704678f83992fc8b55bc75a6f608b22de4b536e6dda94add4e65e3e3f
z0397f6a5d0dbad573d161d31858e432cd85aa77b73b24c8c89fd2dcf2058d631c105b5b05bd5f7
z85132caea2b5456d2e0dd5f063f32a726f69b2deb90571f0818e65cafb087ee5c9b0a609851233
z2a61310f6986bed34e5f0d950e23a9448a6b05e1b878eabc5111237c3e3571415577edc9be64c3
z207bc3883fbee162a51382fcb8a4b164f39c7176182ff538e17c7ac63347ef3110bf79e8219ff7
z1f83b1c98e6430565f7f655445de1f68ee41bbedd9482f6fb563f6ad9dee664f82f7da5ca21bc4
z1439001a974145e2803cea798cfde3714f4a67e2d310223e036cdefe8c92c6a32fbe4a54f351fc
z984987a3f169a54d18a02038acc410a2febbe0a732dd78df2a49638f1e23dd7555caa5229297a3
zfaf99865480219152635a4ecd2e7a23531aed0045c644c8fef0fd4e3e6fa70f6787f4f922c524b
z6604ba95c345d7263aced32d3ba030d5f13407f4b928d95818ce436e777860388aee270889133a
z67f559683cc2fc8d43673e749c9b8036076dc6961e3384324de3d4f81ab0d4840d3dbd3ecb4a80
z5b404bc9290bbf9a64cc899eb22d27b5be533d2f82d284f940adb25c715a6167807e555e6a0d3d
ze786c1d936ee32ac57020aca493022276a6e72fbf877354b7df0e07c2eb030b64de20223a9174d
z3faa34ca1281573f3ca9237efca631039ed2bbc37e1d9eb6b2e6e3bf074bcd97c01be1d5041531
z2592271f3048324d9e4b8c0e1b29b92fca6cdb29900544bacedf5b21cf2b98e7d8fd90ee438b75
z028f6c5ec35b2ba1fa3eaf98149d2efd5b6f15a08424ebc3d7f83867f227d5a65e8411279415e1
z4ab82d72d5110df61561b3c179cdc898fc9455facf2c37b5fa26cc5cd8c57db64d7470694a955d
zda56322ceb3f4a16a528c1b65fa55c6b8b12dcd71a345200273a7aaa7f5c9dfd1ee0e6b84e5e72
z1279fe534877beea398baae65cfa651d819b4e4bb9e3c4b0673d921fc5b2f5ecc16a2c4c42bc70
z1f8e11fd544dcddb8555f7ae8f7b2660147c46b6dfd42e259711c42c4887eee6c64c79a673be1b
z2e74f88a683fadf3110ffcb85dc0b6290f7285c52a908a0b495aab480473d33564db4d0f785fc8
z5f27872428623e20fa7fe23368468a8ea322bd62d377d023bcd94d86ef0bb4fa95620cf406ae09
zf6fac086379cf88dd1ad2a039a92f38b6ceacf86c8fd1b27d1a3cc9ad2a9d5709885c5ba1dc74e
za6769d7ca1f18c5efc2830822ecfd96ac267a3e764d5f6013a461cb2b2ab3ec43988895460ddda
z7e145a159ec6a4383efd37463ff84a4d710a074d55605bf4f98a85a10481f5a7143882f1bb7d13
zc5b26ae56a49e706d53b337a505644730edf2ef2952ac95d15abcb2afc7576e394368b1fc945ff
z75404e44bf36279fd61944d3a6348e6ffbd511bcd7fd58ba6537ad612b243f45398f9349cac444
zdecbce38f1610e4b1cf81749a31e847102c49a5cd16db7d7b91b110d9e28570b367df7d67ba969
zf17d90645fb2317f39285a6c98fdbbca621860ec68474cb55606fcd6ef0bb770cf666cacb3b192
za594ce77cb03061bb3c75013e327c3d3f44e007c6d97c36bad37708b670c14f00d988aa96b8b99
ze74daea0d9e25763d54545f91132d023f85318350f34a6fb4defc86bec618506b44338a68c9323
zccbd75547c754adf2a56abc11667c9fb21160826ff38ab8363398f90279e793b31e98e4c9dbecf
z7bda2a5d3df22c53f5705b4e1125a58fc34cf2f518f841790343241f2a48eeeb86a20c2fd7f225
zc3ca986dd5631cd844c78ca123e6b18e49576e7ffb7361b15e672240889fafbaf70cc5cb82ed57
z4118ccf0744bc23d66b4e23e1297a700b631071abcb70aee2db3d866ae1487af705663c8c966db
z47a4404cb49f7673e5ef69e24ef3a4459a6d5f52e8daee015fc877f1c01fd317b47a44413465fd
z9f0b95dde7629750a5a4578c219b3267e0facd7fb5f2ae85f04cf39dd9c8d9cf43ec5b50d0f975
z66d0cbb49d9c13ca93d78f936d3182b003593342d07871a1ff1c59b9259f3df73ad9d0d9a6846e
z3bdae9ac985cbf8555f47ba17ade97d40c6c62bc5402f68761ec64d6bebfc3a55da597e36b8a83
z7fc835512ce8104dcb6af334bab43f6720b4ca0dedaf65c2ee7e5eceea992bc3445ec67073889e
z7f6ffa3655b17172231766ea96df5b76b85a2884f72dee9861de4710dd074b2e595506c3d3d4a9
z7e6b92eeeb8485079cede4101e0afe68daf143ac153a207ed9572dad084d82d1febfbb540d88c6
ze2393204b0726e184515ce3bb1cb3bd1b7e90f9cce306ccb29ffacda4e49c875991aaa5cb9ab5e
zb2f24119228f6f4086bd88ce5596f0cd55d1cfbff0f2578a405c9ca342feaaa76a7e762a7590ac
zd4d57cdefd0ffc1b6baffb97e8e09a093a5f8efca31b970e05c981a1d0eba683560b122a221d27
za0c850231854c2646f7e9d494d0153336667457f960c07b48f7084c42fe10103009390ff480ff4
zb2670b8ce5c8c3d2b1e7e3e3fb35c1ec1cf37a3838671719778d31623f9c1a17164302506f179c
z8087a2ebb5c36c5f559c1350b00ce1aca460a26e5a3be1b628d5f4e6f5f478e94f34201f3d4d80
zab63d2d44ba9f0b999abac9aa46b836852654de7388965b3b36b6e0e72b5a2f1490c8e93557e58
z2ea7e95f305386815eadce82f53475f3fab4b0c96bbec1ff04ef65c8269d27a8d1ecea4d351527
ze6f9724507827f2db16806ffa47b0ff61bade1fa99bee0eb25ffaafe7a4bd7016d2818891a1e62
zcff908201ee7d2121b81d75800f2e1791c2f0eacc6856880754e983ddb2a046eb3c80d8044dfb6
ze735e3f70baaf627012d48e02923c31052cc1d8338e0c65be8f7fa38b14c99717cefbbdc077778
z8d9a801ae0586a9269a5561c1847c9b9efd051c44e5827a7c3dc7e27d573ef087b7f9ec9fb9771
zd5cc29b0f73bf50a596e8cf913ad2ceaa9d946b053cd0fbd7763133dbdeebcb8b383c077778823
zb599246e75e0c2206dfff30f095cf61c3ee1211e214bfab74844704d83cb92c086a39193e3a9d0
z45ea6e6c0d5012bb87c41b6b5531d2fa450934ea67bf0c64a7c0157d86e31b2327319d037569c9
z808f20ba036a4bb6dc357dc8f5ff623b9378b2bd9a076ce9be67e8e5c20ca29e87d312d4bf3faf
z58cd7b3f900b1dbbc81de02d3cc13220c028bae5015d6caecb268d59c303f0ba1bd84d1c244b95
z76f5eddea98088c4c3ab16bf654493d5c2b3e0a4d3f693a8a3b2051af380d06c57e1a744caf0e8
z90bcfb5e359c1d55ad9edee0062738c1c4ba971f2c3f69e9ac7a264b3e9fedba1d4fb073529958
z28bfad8936d65520d0dffeea9dfb5d4816cc4baac602ffbf9471d460ec30460bff4d3f44bf42ad
z1ee4e3543e5ce1308078584a49f2fce75d7e09752dca36a323078fff17c860a6bd9def8fb80456
z381dce440ee6fcb55a6a715bf40b75668d72cb2d197a2f60ca9d9c70e91650c68119b7d700fbe9
z186c37d613cadb3ff327e5de7dd2e534aad4c6a9902423b601688de99cca28f55fe08299cac34f
za43209a2542b906c9225090b2d1228c83f1c7faec9c85df07757b2ca6ed972fd7dfefd09d3fccf
z58d5db640a4355a54dd70e45bf86bf03af2eb63544ffbc6f1141d817b1c14c7b3750050b58e193
zda3db7cadd0cdc18a8e29a7ba4fd03a7e082d14b6abab90efd35c8ae23f2804ebee9543da30713
z2e2f43ad1c9ccfe957ee1b2220221a8617879e625a474acdab5851b944da5863eb77ef987cfc88
z14653b380e2685071d3e6bb518dd765baebe6b309075e671a88ecd11a5fa6be634fc55c06a7f8f
z107b24f747f51b7864828ae7cdc8601209f3217b6c038ee2ac8f0304f941d3124991a3e3c64699
z34b31f46e47b35196774d05c9e9bd28c4f410ee473cb9f11fd4b96789e33ec6f61a246311051e1
zfe7ea44a42d951abe1176f249c1f755b4479c08167ba839181c45c3a9e2ebfd516ffc00fa51077
z00cff07fb43ae1e449c0793ee55a12fc1c9c892ff403ab3b9af5b38b7b51ba7c6dc11de1ec1e28
z83b1dde726e6eb9f059ea11bb43e7eb11e353d478aa6d909a580d5c730baf8f494f00e944b51e7
zdc9a7cde1061ff64ce6cf7642fe5ce59ba55af20d4f6ac90348f9b9f07db0b316b4d72e27341dd
zd9c8a2fb0829e8556712965aa96da83967592750b42d9af5ed24b70b0630d5d9f096d5fe948440
z5653480473bf62fdca6b7c9f8e18d4989e18671570a51a942c6685ed31eb66d5bc889466434405
z2eeb21053b4e0dc7888f438035627ab9ed0023387ba18e3d6adb02802df384dc096c52a8de2396
zc768c21c94b3fa7dc6ee3f625b4699f3c399ca1634d9892e5aeeeaba85612837bb6c78dd965771
zfa768b742804a81249a03e6a27bc0cf769d2bc8ce4be1ac28c2ab011aa0d54abfc0cb256ba0c83
zfc8a5eaab74c995b8b80c3c0bdd9ecfdb9c59442b2b738d50ced96dd7bafb533b84cbe8bc16c03
zc288d1803b1fdde1f6bc35e56a5b3cc084258c614cb301053a05500d8017dbd831805d08efbe20
z92b8bf017fa08b83a6bf1b988ffb7c9d08c3d432232902935443bcf514e1e253cf83ad1576adcd
z804bd979ab18a4745099d65355c0d4fa2e3cc95bd493becd51c42442599b8d8d319516a56f7ea4
zfecc25decc27eb070d05308f698db4ae862e34aa0d961274d3503bdf2cc3cd962080b5b5c49f95
z2a82d4727474741ba90622f0bf5900e486f724b9efa8b02568cf106da1f0f0785e1b350f5712d5
z73b7d1c9f7abfbe9772d03c5bb93d2edbc7ab462cd22694c2263b9b34b15548a4f6eda63fd05a0
zdbe21acc7135a13be8fe74f0e6e93f671e743877865a2684200f4555d290a07360c45e4647d062
zc63285b306e2c1b8756a931955713abf28bc2ae0d5610ff571af595eda73d845e61cbbeab8ff80
z707f341006bafdd10dcd3e9f68325f2346d667dcb71a61904f8026a5cb8a77227d13307a56f041
zcbfdc25ed6fa559750a3033d813a7387474559a3e37ad413c3a1e513dd0df8aa9eac04ebc20068
z611192d40e7da1c18a9730b5701d19ee3ffbca0886145aa77a531f997b60f0a1be95cbdf2dbf17
z3c10b97cb17b12adda25666259b0b63d0f0e1d79c42bedca6f662ee3a55c58bd04d8bc415c708b
z06299091744bf6a6021fc68f607d6ff524a7bafe204fcbd909ef5d38bd10163ec2551a76c6b4e2
z593613a2c3d6c638c538272ad07336f0af952ffc62c674e52ebf5b552e9d414d5d128b6bc43939
zf0e1513486456ceca02b12dc6eb20152483fa10569bde89a7e553d2fe8bc07a702ff5c908c2699
ze15ef558418a8985569891f2a20a3fbbded3784cdf0c7c876c0f23f35c94509a247f2887a78fde
z96e5dae45b6ba181e290b7b19ff049397d06073bfb2d03ff21c06b9616734a38d38755ac22c17d
z9ac456c112c28ca045586851aeab445a600006ae82fb062c06a10728707c30e15b79309d6e0622
z639803d3eb97835b620fcae3b3aebce11c6dd316aa36f9f9159145777ad0009a7104a7efcadc39
z8c5b446a1ae1799af7d1b36cad56f9e68ab36f2a97bd7d5131b6d116f1124e16cc5a23a93999ea
z08c5886ac24c150d479492da4d7ee37e1a4889eda831c5cac6ba5ac607f5bcefdc4dd9d5afc934
z89a4de3853eaef3a3ae3c26d6b8faa37af588c4d6f1a4861a865b6c0ab5dc5b29b5187be9e8bfb
z5e5ef776ed535e2110e59ab1e7d44a4b16eee8331aa406799bcc1a88ec2be7693eb6c9776a6518
zc3a9d59f439b376ab9bdf65fabf9c1e0664bc767ec815d158ff16443412e6877a57da4e58dc9db
z675f90fef49fb4609b54f21d0360ad1675ce1e58a6aadbfc5b08f197a0a95375d77c69181b0b4c
z59aa1f70fc2a02c35bfae75d5abcce18d800d5788966990da4ee33e98c4c598d496b527e37e0da
z366dbb227a86e1b6727c5d07580a995d77d965fd5b4f34bfabe0a7e25b1c7ecc0b8989ef65e6f2
zcf34b2187aa59bf79670b9d6a51969bb2549b2a07e23d5c4acfd80d6b9790cedf0518866f23044
z30a69e81c55cc819eaf4803c329201f9c68541ae8e59e0f01f8a601b1d1e2cf7817fd2e4548d3c
z5daa2bfbd0d46092ad158aa422f09eeec73cba43c577fdcfe567a6424b605690684a0cc4f980f0
z2457e6399f51e449b5ec1e4fa7856f5fe6b4655acfe74d86b4ecc54d14245e04d5b6a4e6becf55
z7790a0628e5671b8a199e6621b624acd8895e1b7042a4d80478038317d54c63ede6d93107502b7
zd08b1e441894103d97a35c3c4db244ff97a934fe9ee068b01ad78d28814a4ebfc6be235d3724a9
zad92f76a9479adee4106a012ddb90a0acfe973ec086f32c8530ebb39698f59c368250eab7dd5c6
zcb197133c473efb724d6090d8c8bbfaca89ffa9f6abe837891f60343b413a8f8a226534521aa72
z061daaeb3ba290e0f443f36a8acccd921fef752be93a56332952d4ba2f019c1c1ed89399317697
ze010926a53a9da0a93c44d6b402aa5a304f51b932626f430223f54ab8c14159049dc59646c322d
z1713020096cb2be0dd322d75e7c46bee9b82405ef82617d8c92252ae0a420b3ae6d26222082409
ze953631667a3410a85c0299dc7dd392a03bb3929fdbbf59ae0597bb3c2e44bd871420b49fb1160
z5d370ec5059a51a02910c3b46bcc0f115e1fa63ba0c30b68bba631b4fb38e23fb259ee93573f26
zdd3a6dd4f62616eaa2f4d6855357652e978484cc36a41b6223643dc54cc795c755bafc1df584f0
z264ed5f393116e334c3b13ba7b7cdb0d3dd980710688a06867692f21f5eedce96186d5385181fa
zb240780677a63d90dc8bcb751d6f59a1fe297414a7d5237d7638d8f8faed80f288b51d66637408
z2007c889210bdce38f7b902e3b21ba30bcc6e9a95046da503135a27ac01b481ee2d670dd87d696
z3774372366c20404cf8a562d629a5942ca6ee40fc11a4ec9003b6c971d3853080eb34b74081bc7
ze71cb9153926eb0e5fb595152e5bb304bb7483ebdbfe3cf08720470659eda78a3cb8b36ac0ae7b
z3612db84157315bb5e771b70c4200f1dcf4f7ea49214965ec703da9bf442ab336f870539709d08
zd2c2a75272b66630496f0bec3b433a5d65621ec06158143a049e7ef6ff34ae94eac728913d6926
zfe13b547b66123eda672131e73d8460a643effc78c98033f7f0958a4071e5cf9c5476eb4d69493
z36c6a851a3aec2a32ba66d3b0497dc993f2165f28b623f15bfd7ca217a28c3687654a7f21c27bf
z7950ca32768beb7db3fa5e70ce5a83306faf00e1a3ebda3b91d0ba866372e4bdc32ae4738f6824
z37b7cc9c26de1aa5437f286bb317f5410f8c0da8d182842b6f4ecf892bb45c54a1cf8be527acb0
z0d5c12e1e9bfc830b2931fc685c1d3476929bf1124f3e5768855c8d6320db5743c57d845230056
zb6756992b41df35924a44d46c111d577b74b0b31f6d20a63189787d33b146b3db0122ba871c915
zed2896cd54912033957daf32907af136787e8749414d84b731e68466d9b4bd69fce7654e0a5563
z58c6bab15fc827984aca12d744a7b11d39591c376d1b76187849a5634d48e085a907d003eb2ca2
zd8c2ab3d5b1510abfc5b30238bcbf9829446176a05ae068041ab71889f034659c30ee31aefccf4
zc0b19a89e4307ac3e4e11c3e601b5a750172edba518260c7ed164b28d6e354b82979b2d779890a
z91e923dbce055c23a7603fb80de515084c2f076f2d4c0bd1b2620e47fbc1d5e3a562082e5c65e3
zb4be9e305668c43f3a726d5fc91ab1e74ca72c371c762cedbd75b77850f1f2d2e27378cdb28de7
z902ea357c9967d5fa35f513f4f6d8b3559464560e5a839ea6b1e586e5f6ecdd946502fae6b9fbd
z4150c2b6e3a8b9da2b61c60ec080702b94b278be2551549e61c460c371a97c2ce82018be2b71c4
zaaa134b5fd557316bdb6ce0761f26030961ce37495fa9bd859cd142e851650b8787d8dcf4af76b
z0f89e3201f6c5a2b432c23421523cd4ee35888b0c444075fa2dc52f2b700b3936bfec54fd9585c
z8802f244b1d089de4bf05c744af3e922b9414c0887cc131981ffaa5a4a1a0e7707d45e4040670b
zc43a428f7cd9730a818927228d5c4f3f1cf7e5af2e3d32ef4268c76ec93abc8e966e45d53726f2
z39bef1008ae801bef295ea640d6a7e48a9bcee95f8b8b9f4b6a6ab9fb54baabf1bef1656acdb51
z5454b7a7f19792bac1fedeb409edee4df32d09467c5b522760d58be3ae0538280f732669af1374
z97fb3a1536451d6ad879e8bc0779ea370d4c53c30090fd0fa0804859969aa8a2d038e484c00189
z735800567f87c463dd39b72973081787ddf91b929f9bc0630f538f7f65f1fbf4b5adc3ca75f49f
zf9b2b5b2fe497418af4ddfe05511604e7137da922f32daceaa39b98d598518db9df436cda747e8
z52a0b832f919fcdad96ac65e30ffb45b5ad485c80ae69f38099881ddfc475f391407e8f60b4283
z5051944c479e020df093eb6bef5b5426337a77f16f7e819b7b2a3921ef5ed32fd0aef6bc5101dd
z391627ce726aeed6a539b4373235ab62649542575f46c81263cb89de30e0ff7d8a95209b83399f
z33387ff13b6e3c61d9a691015cfa6afaf4f1621a87f0e51d62f10f5c1bb3ee91bae5c84862ad3d
ze1d8cdaf6e3fdffd221599d4dd2614e5e128db4155dc382761d72656055b1084992c578b2e1a85
z9771590a786b38c4cac9e1e4770432f268d34d9e185dfecb9aec840368490643ccd0af379467ef
zc5bdf0264e6bbdf73303797ce93ddb50203547d444636c33fc9c736974e6c786004e0051cdf566
z42a1e0a1a4512aa3980781f91c0f370134ca021fad71c7e7f9ff21aaff4a0fd908a0b43c1c4bb5
z943e3dea41948075022ff15dc199600a68d1483a8773a639b7b5285648d764655bc1d59ee0a43b
z6bef18b8335b583fe31f9107d81c2d68ecdadebd194434ee426a953fa7c85cd37a8b17565e7120
z909e793942812dd245fc3bdf9e0cc558bd405ee0cc55ef81b2f99f86430cf48aa9c93e9c1b2281
z04445c8a82f489fc64121048d849f9b7415da6736c14647052d45f73f78dafd52478aa9d4e14c8
z388a9a776ecd7acdc881b28361201edc6db243d835d64b3e0840994aa3a3dcaaf06b72d7f7da4a
z72f2cdf770dc8b0ff357a9b0bbbb01ad987e5cb2caae2ab44a093aaa0ba74c786b8ed244383487
z3a2d4048f326090d60851f9e10af93164f78812e962fdefea49c681983ade96fd660f5c23cc935
z15245b0d64c7265fc04595006a71fc912244c588a0b1db2ad7eb315deddf0db959e6a5e238e8d4
zb69d0c13914962a8963f685c22db4f9023d898fec21f102b85047dec254e943ff2196c2a579830
za119d328107d7891138842556ca448ba04a8d53390e4d524c593a80887687a88125e31ce5554d4
z0c60b6518a3968a6411a2eb8cce90b964edc0ff0a3b724c589a34e43f547210d99d378dc28393d
zb945649c37f76e5771e9ce39a3e273760e235e7c394917681d45bf7a00d2e1e14ada5d98e49006
zd23472bce1d38dad5579c733d6f084221b4ceb3a17a592c5ada500d674029510a3081a1f3ec8b7
z49405fa2a1526a59d34354275e5cff3ce2f3798bd08bb8733510b034e7561a84aca1682361c36f
z04be9d52c21f4900d7d6fe4cfbe9dbc3e9d7dcde5133a93df83ed1a6bc43c980d627b253ca142c
zb702f48523c200a94dcc4fedd24d4ecdf939059ccb7ec6b9945f280750d509ced98522e4094eca
za2458908bd382fa893ed0530a60627a932a18814e10df70397cd45e9ded1cf935801ad80997bf8
z0b363d7fe8a7f333ee84c6ae3d000c239cd96d249cb01806e43bdf447d739a51d4cb00eeff640d
zad5d6f18d1c986bc425f893af3842d4be1ab09f876a9b5ad742517ae278b200dc11e5e2a1c0c49
z52da4e3aac9ae2018f2cda19a458af70ef4c561edf46a1b93c833898f2a5ebf68e4d127bf6d5c1
z6796b4a4fd84c9f6953c3f491054f3a7eb9d25069335d74cca18a36bc1b200c7a5302e907d4426
z8289c5e92854936566d7571fff9198c79a176504c701f471248ff4632d020f070242fbc68af6e4
za71940abf88fbb277620da48f60bad5654073f3eab7807aea3b7bbaaece19c0614f5b8a5e2492c
z6dfbbdc31fb5105078305ea5eb3e59d926209320553a2a6982a95db4ac7df356e05c96749dbf28
ze7e5f47f5e3689e24d6ccc5f69c3fb78d4b2b94e2ff9a3fe9c55a995778504616194e717647e61
zb158fa262e09328a93b7e74b735b4aaf4a0d3187039ae0198b40d1029982d18e095ac1482c1fa8
z9e63ec0933c69ae0f63d22666e4632dfca90aa0e4e81c44678a1eb073e3899b3d59613b7f3aead
z648a43075ece4f1f1d6ed48845bc8ff5a7ed47bd3685e58a43f300c49a00f83471f794d6288086
z966f62c35b6159706908482ec24e1a372e2a8221d25b36626cddcebb9beda463bfda19a38d64a2
zff649f3bf3fd23f1e44e7c705dfadea6800192a180180514f5bb65e09145eb67e31b11c91f0d97
z82511eb8e88d8fb072a3040bcecaea787170ee5b00f4f8ce362d86ff11e33819a93271cf52acb0
z4eafdad0e50cebb6f2c2a3b127e2d4632261875b3d9cd74bd3a77c02245689a7d0cdaf777f9108
za0eec3bcc97a45b196da2e4581c46845a48cedaf7736c3f86e4fba679450e7dd814fd61229dd62
z93255eb84b15a819daba44b803dbb6f4aa336a8c5875beff226c3b27df664006361953c8fbffc7
za4330bdbcd836e94cc08b2aab3167d74a72777add0d1eee54a541fda149dd69a6c9a34fb1043c5
z1855ff24fc39a62b4897fdb9ab670481b10539101b1b2c8fb9437addd99f694483d81ca2db85bd
z5993a254f240a9246e7027f9e333dab42e5a37796aa84fb8b669ba9a3ddcfa738621014f5a70ef
za13830dcd262a185e0dd110467076a2fda6d9b998442322096275a605935e3cf0a4cefd6460ab6
z9996712a3b82af069ba5669cdb18f7eda1f43afe4d2faff50b96c052162b78c9ab8e69fdb4cd0e
zde4e85e16482b5ad63744e4223f42aab9af1410d0378e67b6a7efbf586cf38e91ac2a613c43aae
zcc804d361a005debcd5a423105d43fcf7db8a2b92f8fcd29f6d739b396be4878e51dc91a1444a4
z2da5cc477f0b80b73eb42abedde8473b3eaca50a79cc40b3d27af9de1791120459c431df4221e2
z594793aaef4daa052e8d99afd867dee82e6833657681cd39894505bbf2c2c84573fed868b801d6
z2802041edd93c09afa581670acf03809e3554237119601efd599a046ab996be8be7cb9eed21fe6
zdf99722748db0b1d172d5dc4e112c6abdbe040912c4948cebb4f4492fee2af7ba64e62af6740c7
z0a11db884544bcf4d53231d77fee340f24dd4b9a6f9155d528dbb5e8cde992258755feeacf07fe
z2eaf718b3118288038124bf5ce09464bcce9037d2b4e1e287f5b60d29baa618d2e1a9b3e31a664
z431313ed829ccb1368e643522d155201dd5f71c4ded0b8015e1859a0eecac52285dd2d9712f39a
zab835c38fd63775dfc31ff7a08e74ec64dc7587d7167634b0b1957fd6f6350493ea2fddd676744
zcde22d58eac39ec94447d474da06b2a56072c4c74d0f6916f32b0876ebafa2614a1e4100142b97
zbeb9e665ccae87141d84fd157e101584b2c4bcb23d780e7e91d7b05ee3dc40888f030b6dadf54b
z79c1dfee24efb92fc257c646716cf766cf0a00d5c664beb3e35075c64608c66d2ee4d360c31143
z38bbeb0cd1fbc2f39991684cf6515903b8d1a739cf07e345dad7ee3491f56564137298c5e34f3c
zffa5e7b9e4cf6e2f7b45ecb9aa3047b3a4a319fd3b3a88385be965ee6ba785d49cbad1cd56da6b
zccefb7b3e0bfe79b8052c8dfefe9fd2896eaf8ecf4ab838ce70a50ab8079ce6081fea4d5dab44c
z9856ca12027c908aacb4b78b5ef72d79e91e1c1bf1aa84db2eed317b9a104ce17065bd90a4efb2
zc153a2deb60bb4e3a468dbfd959d34e5317e0e1b7c21a6551d4820fba2701354d927056bc27e5a
z0861c5d2ccd7bc10324484b45cb852ee258d07ef204ed06fef5b553f24b3b5806ea2bd9d8402b8
z399526f671e4f477c8ddf76ec7a2b0935741e6b2a9976d442e6acbaee3f0cc0473e3a2414db790
zc02aedcebba51f7ca0f9261977372702680e1c81273aa85af004ae19f3db144329591b879fb9fe
zefe73860384420b6482a15030b31f4335c5f232736b5d4637c47a6d95b74768785730ee20384fd
z1f8d9adb15d04e91fc44692e7f704c6295b3bb2112c1829c2910c005e729676fee749707340caa
z06b6cd44e6304172722528c91fc84a841e41af93b1a76d035ae7710ba7065a6a8e43bbd9c4183c
z17f51d612101f719cd309ff1dab9e2419e2fba239ecffe6be93e315281e3a733ea21da32214300
zd30f6f9a30d529ec7998634c7f18e6ae87324e7325cb69655b9485fa5470615c8f02b638085827
zd84ba8ee92f82d7eb0d2db37f3c65abfac8d246bece26130219056dba242d06239d00e966a1667
z64bde82543d9cf383bc2331c99ebe6a10d329c2af2a5b348d731555336a4b36eb60e4ac14a2a8c
z732cffcb7a258255e079338dab88e6018573bfa14d07ec610cee50883ec87feb19c828ceff8ff9
z5f6800cf8c66ea4b59b1aaf172859df7d1a4037449c8f736c980fd9f6bbbdee66310e32b5f9c04
z889f58b26b60bcc476ee532113b754f119e3efc420a29338db35c4516e294b0c4ca5270606a665
z9aa327491fb60f3a66c91c5af316b8dbf1fff9d8cec743e903554590c78334630c17780779aa07
z166d1ed630ff219336fc3110abb82c6e06a7072cdc504b3dc4493e67f93f0ebe30c71e885b6c5a
z4d7fdb09813302af300e3a285a41c34728d2997caf3aee38231fc1048a1bbc97deed0ec0e425a4
zc0215cd74a6f181bdf3f8540bc7b0afef4159d7a1068f59d96e5612f3063b5a79ca4e52b0f112e
zf5419e26a0d6475aabaa16b588d856915c0726ddc6fa78be092d86288a27b7824e0342f4b90a4e
z28b4d79760701a7d1131e1f298ed90ffc47efbccb2f2d82f7bea2807860821ce5d1ca8b3aeed0b
zdb2b4b18750c4a1655a72b6bbd79556807d5a1ba9a0bda955d901811eafc764769c47b5e4ee1a1
z06e38c120418cc43e6588df9109b6c2b8a41f45e801dc2282adcb71a101e9ee48ea6c3c549cbc9
zab2bded1d332efe5b2224e23b9a0f68db33f4741a7b6fbd3d4b4f5f52d4728488e660febc21cf3
zff76f96042f1cf64a9468a4d7abc3c9155eb3d7aa31032db762c4d8c83bd7c351c39e512e4a2bb
z0741a60ecdc32de995cadbd34641d1c0bc9c82105345f086c9af66f23a498bdb896f4505b846d5
z6a50400bd59421e5f18d2182cc8af077aba84b2f919e491b08393cca68dc663924e96a98ff9051
z18f7fb74eb1383d344ec3ff285a7e2c34a09d623c367058c622bf18ff9d8841adbba94b2443685
zaf31634b5be177516829a5425e14479e3816533a4723820d2dc209b6289db0f2f8dad9b7cb52a9
zf9d3b16a2e30b995f1a208d564fea40b4374cc085ba19b3555d0e28f3d6c8ee93c9872ec7c45d6
z770ab6aa5eeeab1e681b1836499c9d03e05957a8ddb82599d7bdce673c7f670d2d8acc066e3abd
z4eb75c7a52a1a5fcbcba33d37b45718012b1c65ead787684d607717acc07ef06fdee9139e1ee9e
z43f8dc34a4e281b33e19f66fcfc34fbbf841552ceedaa2cee93779f3acec33e595c0b04dd88bcb
z72aeeb523752f6b35869e3fdb7339bbfd1688e20aebbc8d4752ee6489eeb8cee84c63072192bae
zac3a3860f1dc7cab0006e10cd8f8333a8bea5059a7ef9e0bcf4dd32278894a57d51e8e786f6c18
ze068f86237275f68af0cadc0beb34d199fb823742c1e96aba92909c996580dbfa3584add2ac52a
zc0424c4ea90af24e351a799fc7458c96849efe0a4b522e470edc2e001319f275676bf59e1e9e04
z3c8b0a447ca4f6dc9337721746b3878cd6d3a7be16306eb9b22f3e81fb9b9d2a81b9dcaae42694
z5564e03dae94fc7ec388a35ae19da525b897ee3c7b48f3a8d4ef5253a9c30a3b6fd4775dacddd3
z277cd1ab17fcb014261577527d43d6d4dd07d772834f0f1639da0e9277a358409ab8178a3c8fab
zd345a638edd91633f707058ace370bc82349f23c7b74367fc3747e1e3de3afbd1444e4b7a29723
zec24554860005b58e37119ec7d0144d363df0f243fb74559abaaec4182e733d77da4ee44ef8def
z9c84a33d474b0bdb6dae6e9e887fff5c39596e91df59d89162660caaddeb64c5a4ed5e4ffed00b
z54820571b0acd2d9f78d7575510b1d781d953efe800adc2467c8c77d82045dd9841c0c655263f3
z4a69b2d07730012a5725d09726c9b9e802306f09da28d0ea8bf6b1a80b73935df06bb5d40ed304
zc993645bdfb43d933fd56ef345af678664e9f6453f601a5ea267d3245bed15174f5e69d64d4ff1
z0169b15d215f345488a87a7f051081ec80d4f5914192a62c36cfa67ed3fe86ffb834bfd239f63b
z694f6a554008093ddb2e2c4b2be9944e075c6f50080f4baccc5887953ad36f17be505f90be4d2a
zf852e2dc3a8cebce8380f9ab390a0c306c8b3e0cf6932c448c30e62bd8f2cd068d5eb83ea65afe
zbb30863e3856733e85530230b7102946b796c5159792303f3a8379cf876d5065f6bd29df60053f
z24ade7ccc80765fee6de37e7572bbae3b75b598ad024fee10db6856dd798828aef1964f79f04a6
zac4626e90b9197b69df08b08be0c39d18b9a60d2ab3738b1da08f7d7a7299b249768e592b45c75
z947381b6b6b9c8f9e26e0f83229c044551c9ea2b460b2ace15751f7bcf6b0801e317ec974571e1
z4fb9cc503ae54f5a301b6a6891f8a90e73abe8bfe8669f8ae8293d382704f4336fb97ed16a4ed3
zdabd1ff9f927a8e22dc29c9e8444fe0f3a323c7800d07b766b6bf35d7d8ff9ae28523670dd5c64
z3eaba126c7e91022226457a93a5ec9c8350b1695a926b3bce7b4a7417b307cfee263bd7512806f
zf2b23e3a92922449af17904ec2334a27c4f11894f2a46f6fd2f687628447e4d31a978c158c1fd0
za619a553803274207af5849154f6f058062201bc8bbe46549342f04e602835e09908fa3c3f3773
ze76485cdfc51ce534fcfe5d5f5b1f2c94cd9d2320b1a9f84dabc79cff11c01cb766c321cba0555
z3b87a26a5f47a884fef028256ecdb527498f4d3742fc2f3028c9332443ba869f6dcf1b8d463b24
z0077f6ba700551095423c4105c56753d17c5fba3fa0862b398eeefcdb7b27b8a28bbe7141eed46
z1a169741a28272b7ea1c51620c7e0e51420108afe2ae7581ab3f1ddf3a51a9ea02e51b1a150d9f
zcb2795cd8a551a6993dd21a9118c5822c243140a355fb3003cb0167379d75d1250aaf8729a047b
zc01d08968e1fe825056b4f113f6e222e73773c674100b44b8fe23eb6b1c34b762748eb018fb4d9
zfac2463b601d86f4c776ddd34bbd215da5fcadb38ffc03ef2d3a20954223fc1a7db4b6fb82c940
zc5d9fbee5a31945496f0f627f8b035b0d5d3418d48db74dd07b9945ffaf02b836978c3aa50bebd
zcdeecc9ec535af9f61e98176548f5f91c05b17e41ffc43689fe99d4b54e747c57339ade6e776fc
zc003ddd715dbc885a8c4175427cdb6ef3f334b8958c88e572013289f0df91e2c59bdcd54d42e63
z06983efd469ebd61dc1a1530f1dc733ad993db9ea5431c936fde056cc0da8786d5340afb42e1ea
zfb0bdbdc6eff0565057a53a4cfed91b4853aeaf8f9ee30c11daa00fd6096adaa465b6fd08ee5a5
z94dfee743bb4605e546a1e3f44892943ff58dbee0bf3120de74da8992c31314c7dceaddd6b22ad
z942cf34c5287cd52df02bc2eed108cf2b5b25b4e56534eecc110426fc34185cbedcecaf58453bb
ze99c2fd395668e7b5c70863be6971ca462f5c28264cabd204428d9bd3d3e007a37674e278de7b9
za40f63aa9e8164afa9be3a5bfaaafb8715920d1446eef7c2b460ab7f83b065b09f1660e4712d44
z4a5be4f582d48df664730838788935af10165fd1d46d589e65dcc55c18acc11c0d1de38cfb5cca
z4b18d5e9837cdd749ae1c1d094ba1b28af8e34bc235bfab9514e45c986ec8e89238687bcfeecff
z1b42a5c38ff15c36aad3ad6233d10b86efaa5750bae369aa326822bca6287f0a4c593ddebbf3fe
zddbe4ba6b4bc9634fcb10a5ca2190de655e14760a80a6053e5cb4fa62fa95fca99ce9292b80187
zf394f6acdbb45e2a73fcd1cf0657d4553559c436c85625406b38834d8b6d2fec41436154a2ec51
zfb80055e3c4869d5c175f503917a627aad609bf56567ad74954e5c074460d97893e4b9ea4079fd
z52b7a4f5ad2a89a2aab60580fe8774970026451a5210581bc6e571b4875851f9103293390d76eb
zf834bb5d043f04d2474795decf63e319dbb85e78a75b9559c9c27d1cb4780eec45841c591e9ded
zc3c765d99c3b0c0791bed67e8561c076dc74d5e8ee3f77b6d07160019447ae62258410523b719a
z95eb5ffcb0687dd10a0ae9473943c0c299c970df01829e30bf3bea74a0a896832532126160803f
zb4c9e1649c9846ea5753c8eaa426614d73f890ea2572accbe80e29f23bccd14bf7feb8632491f8
z10000ae55da8e0903ef8176b2d2358a9a674f54acfe12a84fcf274e8c45d6680ff32ff8a7651e5
z534060546faf537d12b398cf0f882866cd789e80481cb52f1a108f93d2b972744b65dc5911646e
zac15caea5b2d518b7330cc29b4876395feea55a00b85fa5ecf3523115925011986010c1f700ed6
z638751dc90818cffd2e39c48e6d43d5f24a92aaef05377195120fa0960dbd799c97c5d7626849a
zfdcaaeb082fbf8098a7f3f75d979e102e644720e04a022b8fa2bd0db862a257e985f6bf4373ef3
ze6eb37f2e036337aecfade741ef05439a77ae4e159b9c4f5501fa69e2a7603358a297cb356358c
zb28465c7db317e5d5dfc7ac0eef7b17b18978c6a8fec0d369056650911a35cdf04a124dbad60ec
ze07ef14032b6cab998b04e2db2d41befa40d429787e324560ff7f5cb762cc47c21cabc7bde921f
zb5e77e4b3d5942c2b32c8cadd3e3b9f239b54df7bf1b2a1010fa2032e0ae52281921d4494141d0
z41faf4e940030ba527609d06604cec6f85de9598485ff35ceee36c34a994b1bf7ab53a9f3c7949
za075e405281bb8b0a30b6cad85b23fecbef22659b813eb919211589097972eea4af3fd7f200c64
z1a77c147d84493f0751fbdad83b7ccddfa7fe144c5d16b660942ff2c0441abe418884de282d1b8
z9679c7c5206d8738fa8edb519358d7310c5156b9b9fab8745be874b6a98992aea6cde6d0a614b2
z5c18980abc1fc92242270c42326f5b2e13343b752b5263779ae7cef76de5692ed4e2560954a443
ze6866420d446f2d768d6437313411c72c92279169ccba0be467b737f3ce76568af7e7b58c929b1
z410a7d46a8441f3f74590d920440f37b6ca2148ddc7d6b9d21b0fd034559b2843f99df2e5eedc9
z0d4ac535de34c1bdf903e2e86214aed28b907ada9ee26a91a7734433c1c44305dd9e0f3ffdfd2b
z27c4401a671c4a64bf89adc530fc2e4e5b95f15f7d84a6467b4791c548b72dbb864c43ebdcfe5d
z497c687d738a3e6903b349b6b9c0cf4ecc6fb40ddb7560767384b8c26c4e8521339b09c235303a
zb1a0bd87ed64a6abe899dfe8baf2cd03cacee43f17374d7b7067ab7da4402ed7ef0e5356344b82
zcac2e8f2397e89cbe7087099a093fef959538173ea6cff2671478a7284bb1b85dd3b5de1dff13f
z3e3518a42fe5a517ac5d7dcfa61970825dd3641eac4c6c3a502c1144641345f302cc1ee3349b30
zf82f584a4ef1e6eb5bd4560fb76813518f65b0d4765a64e0d3b2053142b04b17cd2e5901fbfbc8
z6a2a070de0e600d506d26c4f851a41ac1af9a4d39350fe73894a89b8649fa523f1e103b663ebe2
zf56d515a2bcc717afab3ed8195e36862d49ff33e35be563662db904fb559ceeb75bfe3e6a6313e
z2966b567e179d4a06e98d11cc21961e48b618bc72eae3e496ea9a21aaf68386511fe61a1bd33bd
z0e69aec1313996dfef2c13657917b62640055eac3d77ee0669af92f9164b8deed24383ccffb6fd
zd7da6c4ed9527a3bca31a025393bdd30ea6aba218b31e18587c3f41eb9cd68bf0578d7d0b40f2d
zfe500310e7a4651ed2ac18b75904b0268a6fbfe5a563684948776c3e628a089c57ea67a3432823
z0848bd4efc3cc0cdfd6b484c8e8d033d2e70c80075c9a5c92edc2a9e3bb384ecf6f93d72b54196
z84fe09a067594c2e105a99b104aaa1b39a36530b2cfdeecb7cd3accf69ab9d57e46b6acf11b8db
z2e7677d7c47436db132a1fd22f0507551072b455fa42b3c50e0901752689c55beff971eadf963d
za522ac6cf6d9993ce9e9c827ec9caaf9fcab615cf8517b39be566aa9302e5a20c23dfc1dcb7732
z17bb6c43534332197c7f41dbe93c78eff3fbcd8eff67a4040878f80e30c651e36c5bbdcf5674a3
zb2fdb1fa663b2116897e0537b6da5c2e0b4c896ba5c5a2cf2157b1c7a6b71e007ffe0434f9f44e
ze37bc6726c7dbb81fd5d1450a145814ecf3f11ac71a06b04bf5d2ffa807e94cd26c5f6df497357
z8bd0b3352c063a57bc4543a09bdc52daeb3e9bda73146722cd0603c5346b8b49ca17823d2a7d9f
z36af86976356253b50ff42062859bbb7e157add593e0f90c45df5a0b6a0723192a924218fc1cec
zc36329a2ee9c26c5a6b651dbe956f7fc0dc5d307e94397493395ac1ed567f198d69bdc31d09b30
z0c211ee2cee5759d6ee192e009b2643e100c641368af1c6667dfa9f15c7b24930ff00f6d22e995
z679183574fc6493baea78f1bd2c17729b26d3cf4b7d80471ac512aeb0c2e0a2658770504111306
z901b68c0cfcc13a1f73f7154825fe5623b387e389694bc87097b32e3d640266241d220400c5b13
zdf2eb98e15d83a6cc669378c9fc8d8365072b8471e8895c9c5f272b357657d9b980bc26bd66bfd
z0fbd4d1473a2747e79ad56b59e88bed29c66529c12a8bf291d301a994d2fee8d8174cd2702234a
z6b0d3e29428e8f7db2fdc229e48a339ee02d02c9991fa17896e4ce7db691b324e25839ee446c37
z8c100a64b3341570c03f81e15622a6f930a9706118b1b2b463a15c1ab17dfdcf2be587c2f826d9
z71110f85ab5ca6405071413b88e7e3c7479fdb671350086ce776222523d572e3e1b147e6f714c7
zb2ad561972fa49708d3f651a8e216953d84b7c4e53b0914b01db67555d90a1150ab713d6d91d1e
z69d3d6a6ab95f15c5cebf1b6171b561fdba4b6120e9ca4e0c480f468a7e56f518f7b57cc21c2bf
z977315beff5f66e19a0583147bdfbfe3dad6dbf0efd8252955b1bc4b1d5d5f7a295e9075a325b8
zbb74294c78a982cefbad9cd9bf8a85abb1d86bc173427730d44b3c8ea9262c8c99f31a628db838
z98127d0dfc8e757f43421c9a78187df85dbf2a92fa17fab028d091b94d79d4afa7b50ea70b4d01
z3b0c25d6a8afcd4bd9ffdbd39f31ca31de6e9957b0f1017054aa2965b73b7d889410bb034d1f82
z77d35ee58b0a3a576ff28c84ec4ed63af1cf31b9cb1a8207056018f309fb348b432c034f56d701
z2fef9c353e52c59f87f690f82ba7168bab13f2b7cc3bfd9334e969368bf69811c3fa242a854dca
z49ba4f40cfdf0d5ca9345fc931496c1b46f071afdfdc6fc0cceb9d28a4744117dd885084516703
zed5c4bdc735b8626da838f6c08bc931d3635bfe0fca4ca8f2667b5095e2742ae08bea26a9a14b7
z23cd145c3038c99ed7edda064f61e2fef7a671f017ebe11c295819ed3b72b51bcaab3bbb8c7954
zabbada2705f9c876236a17faf385ccfe2b37efcef2c994a3ff0b7d33a15b979dcfc1987232cd16
zdcdf5034a91b588f08191d2c066cbaec70b8fa84875544addad406118ca38fc6165fe9ca479186
zfc60a8c2d5c97b9c450479d208e306b139bdf8c32bde02d4ef461855a47cb1bd73fe4a60023b8d
zed1238c59bb37e47ed9f729cd117e2da274acd6de37e3e6e53a637641f000ddcf3dbcf586dc32c
zf2ff8f47c53d4562bcdf7764859530362158845aacd46eb707def060a8fa0d888835a0e2a13101
zb67f54ba85c7adc8ff94438c29907c80cbc26683a6c5bffc9fba07549541e60b40ae7852b06aa1
z90f3421150c1b3f1f86a57f6aa2d80bc080b0831485fa650638d60c0c0b7cf8beb45fa61bb1e6d
za1ba9baa1cc2aa579ad38259b9f7d5c8dfc5f3a2603a9570dc675e8acc8009094015766e1b68b7
z3f40e1303babcbbe4b1af27e58bbbc6013d5cb8b299371bc097da749884e6cde8219bdc7212d4b
z33d4d56b1a92a87c27494dccc7fc8364106dbe19b5004407fea7aca2f7186133871f66ff691f41
z09ee9d68b2d00095561398df0277c64e84633df51e3a33868af899f8c5eefc6ec2f8ede12c097d
z7f5fd9f2ed03450c891dd976acd1cd55b034ac98b78a5925ee335c774bfe184d061ec5ab077d51
z8c3a29739d336fa9d46fdacf02f89f0247f0a86a73e84a86a5cfcc85b7909a116b171fcbbad5b1
z3c85a9116dae3c2a2c92190470c9db0ece89552ce9128a444355f4cfd0b8df9329bc961a9ff0f6
z74e8ef43576bbfa17b1415ab7e9d1d24a889294ca339a3efcd3cfa0438c7ae2b0e71202afcc941
z650d79c48915a3c59ef4f256bd5dd0683c33c9a5fe5199b6e2c7ac9f0cc73e0df903738f1082ef
z203a3818223d7d76cca91cc1dfcf73f1d24a5073f858cdbdea0b782e45d7d14e9d94cdf66e023c
zbbc94198143c1a4d5b3765fcd6e4d63ed6827e08fa6af9b5ed59facdf07283eaf3c3201ad5a5f0
z5f37d11fd56da727511a937f631c7bfc96b2db4843a0563f5bc40f7e10dbc871be5fa4ac49f034
z08bcb4f5a5a00a6066c58b107fe3643e448a41001d50eb5ef02c4fe30087565330cb3c6342d977
z58020f88fe974657ba97e21af9a41a24bef7cc2a3cca95e6f0f2bfdcd9a3837342462f20f1c727
z598791de384c5297a3ec390c07a21a82c644b77b1f35bfdb78862520a0e6320546773242086168
z08fc4e074c21e5a136e005f15d3c591d8128f92399c5e1ce8b0f8ba047869e40592b6ac21782b0
z964cf383dc22f3c2b405f14b7220e684f571784221437e8b6b8aef29f0a744a6c5e0ac84bb7eb4
zc663c58ad41e9fadc8941cb2e7c364d22386df34b92d927eb130344ecedf8c497a3e2a9d9900b5
zc0bb2be58addb455f0269e8c2d94936593a9a257ac1ba322d339389d7e2e1479acfdb18276143b
z2a1f9d1b2c1d706cd7c2b11b1ad9c61f767a532802dc6811f1cf5a1c61c849056c8be239c560a8
ze9d859045b446a9a3d05afa06a06469b4e535e1a5768d64f4fd01bc856da5aefc0507bdf3c4eaa
z192d513504089f48bf95da22ab80d45198dfddb538d5bbe81b0bf49f210e6a8a5ac03a74436cae
zf96dd645afdacce24aedd3799b93f16a0e2287123acec8c30a4b2cfe44d528fbd21bd869d99f0a
z3f294da43c4d965469021cb82439b1c39a3663f34fb05d0660ca218ed8c2d9bba4cad52984f8a0
zcecdf46a5d80aaa39e6c98f65be8d05e183bac33f435fe8138db476378ce36f8f188d322df7d54
z554345f8d52a0d235cbf3b0bae92b9aaaac3f66d740641f489e9b36e1184aee6068d3fd15162e0
z227fd0685128b658ee23e461164cfdd46f62fa543f6fe0d9fb5de81922d0b8c755eb0620928916
z18411cb0ab4b862151b019b99a9976926d69cd7a2273f3651de6c52662ab61ad4c01b2c0953024
z022854c3985cc113e6f366ea0cf09de2095e8231c9438d5ab07394e3dbcad40f072b5a772d9059
zb521037690de2fbc7793e8c9fdcce99cc59e06c93f883c077f34aa3bd1fbdb769821aad0b6b98c
zf026caa555a9dc1287cee1484dbec9d69d208dcf9d83135220782aef5b142f5c3399c4cb90883a
za19aeb9e38eea493dc13f41ac71fc69db044fece37b02c34a68edad48aeeb9e3a6144b540c23c0
z52f5468fd0fb22071cc1d2f0ba15c4519f77b788d6427f6fce190ee74caf0e0c60a53757477b14
z775eb7b139b5dda2becb07ec79886d17bb1fdc01f7e69db08407f345cb9fee706325083eaf1b40
z0a429cd8fabaa1ecc35175cd456374164c3d732ab458b6f05888f5a4037c6af3f3708a0acc4abc
z9c20cee1da515788a14b9eeff0697c9148e3d51d9d8a86e8ec0eeed7d828e3c5b511b11a9b40cc
za1a6225c69c0ecdd28f308269cd38742a0eccb4a29f97e440c6e59c80885b6ac1cb8b897155757
zfd57021a5d38bf0a1f1de8ea58dc0a56decdb684dcc3bc00b77712d278576cfc76e3005970dd32
z24cda9283c06fd6300fc87907907bb2edebc9a921c0aeb7ab4660f8d1ad862aca32b281d05be13
z9b2aeca45b0af3d7a432f7860cefa2af40773d76e7ada6426ed8f30a8d9c7ea2d72b640be1d884
z163b6544c0e7d7e6e5eff306303b405ed775cf5be84f2b3bcbf522073ad139dfa85c56b8f58791
ze1ab7e75395b3598da7a9626b00b15e7ce8544b8e7abb940ba729641a6be88179de911f02df353
zd77d7dae3078baf57b77cd7a51e1dc70e1c658dab751db5a2d49a1ccfb759b1b1c20b1a05921f3
zbfb1205ccf3debda3258c3a36ec26325fff0219aec9041f820f3f14a816a4a87462b9d43729dbf
za2a601cd68a307178e1019d3500f8d8fc02a6ebfc06310bd2a492c0b213f496cf669ff80379504
zf3a50b9876e0ce827196925d17c92e54a388a0f44c2efab15b3ad459e6bd1e321218d5bb45b77a
z4ffec8dbdabe4f335cbf81fab49f81cf699fd17d0193c548b0f3aa348de41ad0b0f5f5e1765495
z27cc5374b0a6a94108fafe926ee8ccd2a39d95eed467cb4ed05a622310abaf83d591163492b1ae
zaf0ab3dcafc698df6eaa3cd2b6e2516058e623375d5f1f438da8161226f66242820a25594015fb
za31099babf4b79c1de0eca81dda35e88f0c2daba7438dad912b00595f07c50c3e41c6599ee11ca
zf136daa178a505314474d9feca2989cc15d177e21f94c10a8b9421a7fcb29aee5afb1cc1fcd130
z0e692b977bf75e379b1bbf05b5a1390029c04678ec8f06552a99dd3ef03b68d3b855f992cbdd8e
zfb3d7d88c27d6754a00a5087d43ba9a8ae7406fe8bfb72aaab3779381ddb2cdd82279264be6de8
z1774fcdcb28854bf3043c9e17175b6353eff80b7e6036569e4a2b18f7f02e60cf1ccb73e12e0fa
ze553f73bbd7ac6692185a868dbfc2982d85ef788e75a1d2c3c1166dd421bdaa592833299bf35de
z98868b0a1313931dbc06d7d9c3e787476201f386fe9e959b273fc7100564680994bed320136f29
za68529006c475e5089698c52fc26a897b13edac3f830eccdf692072d80750e27d4eac068852fb2
z526ad94170b15dfd37dc872d4dc51ba93023d1702d8204768304ca00d150c9c34db5adea4a984f
z427ada59f1ea3a004b2a7cda094fecbac824cd928c57d30054ccd512fd9db51bbbdc7f72332041
ze6674ca8a6e225b95e7fa4d518ff00e13063c4bff12dbc3d204947ed5d64b7f2e1155e576e31d8
z8db7333ba3e060c2dcf253df28b4cd077942e708ffaff96d9bb260749af9f73291086e753776ba
z02ac8360ecae66c23a44a02e1f7db3784c4b3d6d57a9a7edfb58ac895b0241b487407dfa8932d6
zb68af101e879d32c91c5103984f46df7198d613622cba3a9bd28b9f8b74be913002623ba3b1152
zb425facce0a18f8df2558a09f22ec86dc614620d5199f7724b2974f2a16a02b93ab5865cf95013
z895cadae1a9baac13b5c13a23e7745a89469e1d0363bf74d8f8515b1bd288fc3a08590443be59c
z6391117eef801c69a06571d624a6877061318f0134e3e718e2e352a1c11d86957057f1990b181c
za7e1aa1ce007d5b6dd0a47f404e7c5b96c8bcc88496d3e48131bc62f9d65ef95910fbbdd302de1
zfe7a92b617be4eab215e42054e19e1f7d75600be3e7c47b046dce1108e94fc5178a296095aa71a
z8ef1c89eca3b8310dfea7c8be5ec6cf93ffb640a38b0d144492828985d171f179525ab0307870e
ze81e6e83b14de1ff0ae1b919924aaebb88b6f473f0decfeb7ae589743779e9dd6a857bcfea1aab
z3f4ca97c47cde406713819c455541e82d538a9713e04e6d245a0be86c77128aa4d3af7eda3d9c7
z59c84e814f4ad2378f7935926bcaf963ebb7c95bd6ffdb8142135e2ad35034ff0a31372588dcfe
z51b1865b3563b6a42996037a6c36ef79c90e8ae93a5707d43c87e82088eb1cdbb3614be69cc195
zc295c97a63e87b2db58730b43fe740c4d9e05fada354028dccadc0349bbbf24d0f85dd6c8d78fb
z9668adcae3466d184e4ebd34bdd469356fac2d15f683c47b8b2bbcfc6f75323ff4513cfb8f4d4d
z95e8ffd2f63603a6ce77d1167ad4169b438912284c5764b20274f1302b17c4f667a098bb19cd28
z786b2cfd0d464a0a93c2b3d0e776de58ad2ffc51e4e7bbfe0cc144852a7f0b05e69b32ecc28893
ze7160ca140156827c10d1dcefeb2391f2bf5581e1e3fe49fce6f43893264ed4645aff479b63c98
z3ee29cac520ac5d3a229480441d937cb0fd0726a841a077316c7f8c81475edb1a9e90a07333aca
z925605919567c7e692f8e324d63291c59ed0ae7b7c62c61f5d7ed4ba5c7f51e07409d4334a8cd5
z740be31dad331b0732b7919d5ba02cd2e0d3b05db99e504c4730c368cac3ee13e3b71b5f2946d5
z4a02ad2ce1837dc690b4426e9eaad02ae51cd632d8b57914913011aac6fe70f309f88924814698
zbf74b15159965a1ae1a620358926aa48c8601d0a122332bfbdec5f8882ea7b11498290d98a3189
z5a80e912c734d3695b6924ae88eef15a45c9e9e64defc7b0e7bdda34a271cbc4557ee621b63b09
z5e18e9e5dd7d73102d9dce6b6c5c52999b5ba3d4f680fa93d5141375ebf03f934a192d79de9ae9
zce0759dc1cfcd7a61b8a0ba8dd1196a40801732fca9ce3dd2b90e8a3378d8395b733de69133a5b
z16c23ea14c97d122ad3c7b0329b06cb8de975e5e8bb1eb766029b54797101016d3b9df2d6e563a
z384bfc7a39cb5be270eeb3119db6bc009006e9f5dbd2425c987a879d70ba3256ee102c721350de
z350d6210a51dbf6ed35ac8c3731790108b73620df40172443aa3c4d9ca18717b484d5afb99c88e
zee7b469732c30c6e06adf97784eaa431dc15fb9379b55175cd466ba372a7e30b2b708b18cc4bf7
z856ab82e16e497a398476950a31cbf03b67f319d7e00bee3d4239ad62d96f93fe683df864713b1
z64bc813812c9a583230ad0957f79dc0073375b41af6b0e0c4d55f12fb4d6d8a900ecb9d0ddf17f
z74c6f5429213d292bed51edbb09aaf15434672254003f0d95733eca8710865fef01f6deabbf5dc
zc2e2757e829f010190c730bdc3c8a8eee77079f18b11bc078fa92d2fb1df3353fb9beaed18d964
z0e249f6a897b1b057ce5f7f1fe9947c353ee45f1f512fb226773379c142d1cd74c8ec28edb0d61
zde6d923835d2f2b3ad0b34b124b93fe01e2522f20bd56377f445c6ff6d9fb0b8c9bd48c4f86ed4
z1b9ce4aae70fc1ef5c04b2abfe334e4103621b1c9a184db81e57acc31da28247ad072e5f2ec83e
zcd009be14133e702e827335058185175ffa766dbe960f4097dc9060fd3419cd6e63eeb420e5472
z6e3f59eb3dd32fa83ab7e6b4327b6891dacd91bde9d0ed497cc4e6719ff54b9686ae2c9c727eb9
z107805102fdd2ba6acb59ca1cac0e60750c52a381b59286a35d433e63d867f7fe7f0dee67615e4
z030490f34b79df3c6d79f58b867aff683e426c420ed9f37047b3b78a9f2d31e16b08bcee0d962c
zf99907fbd268477ab5ded6bf9db3fd4077ae150a09c8c4fba48c0058f880ff71b407a90c52a711
z77f58798d821063315aac06c05e2c10b2cdd7e5457e2e4ccb0fa7fc71160562cf3989de1ad8dbc
z34663cf3b887333c49f005ef47202f0ac535ec440cc28f83a43cbf64e26c7d462374a6f4ab91bc
z7c30b4a1d28e3a772bbc931b56a3cd0ae81ab3e2f758d1209d4b5c19ce9f8bca1ba8c86f6162ea
zaa4548106e8b3289ba0c48051f598f88a74f5f9ce7255039733f8b639203328151c564734090d0
z6e859278a62cb0a399c655dfba92df11dd52484aebbd7825f789c598aaa4845428bd09bb081c19
zd6213419e3e02b85632b280598af1c5c3d7cc9dfbb9665be0a18b132a5789697c9260ca47d931f
z7b769538eac5a14945c17f7734a922ac474a24d7f7dcec1a6a92c8a5ec3ddfe3c13be9a6af9daf
z1f5c5a4d1f2afaa92f88eca71039d6bf8c10697593dde9e43bfe56baaa6d4134e385314c3c4475
z8b36dac1beadebbacad38fb1e141e319ffe4fb9b854c382f1aeab09e91f0644c0dc122d91fa918
zccc834843da9507cc778ed43cbb553a431eeab0e001b44de039c3de7db23d0d8ac67c82de4fbd2
z4156a4c7cdbe1d4c0f08a125662f4cf37326eca4489e8d44041ae6e2d1e898ab6de7f328f6365f
z770cd9aec0f1591a1c880e3d46f4eed6c61a1d282b528138920d8b0a1095e819e7a3671ea70c76
z45680a1afacffa7427c7bbecd6bf6fe3b3c3e234ca488f66dccf654db38607efc511c0211a5f2e
zb2ff8ffcf0af1a02a6f7dface2a6a10b454d1824844e0b14c8ba778ba6ffd5a16f68fe64a1e3a2
z86c63878486c7ba06a8ad78fefad9eafc68b6a97aef032742b747aeccb1be67cd7e72f49ef04ce
z81dd53be36d6f3c838d197542520b1dbbe6fbcfecbd90eb8d88f225d3d89af4b7f821e3a4582be
zaa05052305a4f93bd451029d1a44f068d906fdc4758eb1bbc168f01344bebae794ecd119d8abbe
z1eb0b844fd06d9d49944ba67a14ed24a017204900a979c7e421ffbc7278353153544537ed81883
zbe0d8aa5ca80948247bf59eb3736edc9dfbd54d1e607802476d1c34493882278d432c29c4ccd63
z4db281290e7a25988f3c235c92591b7feeda66d9998728225787d570e8172ce84e8710594915bd
zd4c1ba4544d34f82876c08b7687c03bb2c13ed6d5c06f75d361069d37382ba8e91d895a39dca74
zcf92fb3902e24b9d42b4745b247cb7f4dadd1656c8bb17a618573c51ba11c8d1459029346b3a1d
z659a0471cfe98fd480d1b62d828f1901c8be735569015cf9901e3913ac0a89732373f14a047c10
z8f3c5d56d47c571498a8a6c460ff3d5becef4c417e8d5d67e80f67d377131f7a09b6b2ad79e92e
zc4661e12c761540d0926104d88d14b8b08463072f41eeb73f3a51bbeb42affd05f65eb8c66b087
z196e753aac2026b88e04a30e51dc0880458d7bd6d256aa621e5101adfc35b4a7ca28a8600fe880
z0b0f0ca210711fdd1cf37f0d0d04106a9f5dff398de86a93435027ac7c0a72977b58c9a6962e73
zd140c7203a1ca7bf26e9268265aabf5e88763cc9a03a04663a0e556419ae7c2cbcd12eb0e409fc
zc9d0273f1e37df872142368c605cc1f26abd7c7202fbb81a32aac1aa0f7b830e79ebf2701f33d6
z5a1500a9c0c29906f98333a8373a8dedccf360482801859b8a286f1482bff077100ec9e38d692b
z0bad685edcf2a45893286bddbd5c39461b6d5f51e940c98f93a3e9a69efcefae4f27eb60bc6a39
z73b3fa2f0ebf51b2a412a62ded2482680a741fda6ed67c19ca07000fa63f519414a893df5c3f7b
z547d731cfa7f66d09560e2b4d7ee9b4369539e5cd565d889724431cec8e7b1b024ec1cd52a4e80
z7559907804cbf69caf8a949f2a46cb19a555ed27904a21b5ef775e1580b4552879084f797bec09
zb4bb594f83aaa62a0f3fdd2076461497250e19ff27d5a95cb062eaaf46240da3c533fb1063ccfe
z0f7b937630c197b741fcafb369dcebfa50c8df89951d721d6bfcf6f69e275cbd000e2f74d74272
zddb0058c162b370b91729f000b445197b6ec2715a7f393e0f7ea241aff7743925e9c0cad16d8db
zd4f51fb1ce6677dd13b7792be271789870e0282a05ae82f46e75a3eef0e81a7c611d7a7e420ce3
z67211e1231e16dd1ef9a23c77d70bb3be74bf4329ec9f14e56a88cc6a9b44aa6c2d9c8f8931b41
zdf12dff4861fcf2bc7184efe2a132c1d8d089fd87d81db65a1603eb1230815706f6268dd8264d4
zd76af5e7e5adb9a0615e34320c058be48cf72ad6015dbd354eb0e9a84f03596518007168adaf87
z2f5da5bb9270b68905f6492f76e7a8de355d1dd82bd464d6053e05174da9b4d0db94f42a1b2937
z69eccdff3222cb915ebf1c80602090822509c6d14f45a57966b0047e46acdea6319683bed1bf9d
z90bf01c21f9f4311f33b3b046e3803adaa33b20d98c562825301118ba86a6f09606e3bf88eb02b
zd426c186469599a720842128696c8832abdb8fd6837e1ced38fbf39ae62d396c9611561daac033
z797abc5682948a1d1646bfb61f955bf157484be92b27d4365756c87ca5710f72787863cee8444c
zfc3f652f6e7500be6cf2d3c22cc5316b234689274c203ab5861f9b21636de9e6b32bc0b5138005
z80a0c27db91e056624d744ecf3ab5fa191f20c673c30d1b2cc158938d2727eae93898297fb18d5
z41fdceb3e87d066802b25ca98b41e82eb101be9c1ca494e2857272fbf43da73a6132fe9757daa0
z52197528fa6b9898ed0c6f09a1c5afac4d8e1928da5e7626a528e33c9c227f77f1a2f932c7a881
zbe4e984680ccd2e3e29a37bfa9cd3e26331e793ab0ce856b75de0b9ce65fc62eb0ad45e411b054
z5eda3ebc20e9db2c298961fc8d5ddf87300e1667104831111e3abb9d2ca731f8e68ad86bd54dbc
z75775e73484b78a91b35e893a54e4c3eb510af3638beefe59304ec5efb14de0209e1136fea8920
zeab8c4ca7e0874b80d38c2a4daaa4bf82f6bd32d9f357cdba806a644540fc241d9fec8432aae7e
z7a8cfb1c836f7a03a930490c488af3af16b27ed89c897fa949c111cfa0a5effc30531f444af1be
zf85b1216d80388b97e2e0732267bfca25165a46855019c58784cd23203b92e41cf535f5822e02c
zf9a53d2e8fc9e455e36a44f62378058552128339c1b3e2d8b74c17d3a989a2fcb8f2fdbc28750d
z180274326c431a508b6da8d0393483bad03fd109010255c7e3830546301bf829a6fa1da1f8bd4e
z15d260311117efda2df70497effa1fa0c09fb43f5e6d0109f735bc0be0cbce437b22064f6b7931
z6fdab2ce48736091166f448054f729fc709feade7f3e9f2cadfe2daab08fba374d1c9bc3ab9e2c
z833b3fcda2bd11cce511e915a6b3c39981dc14b05f979735f7c1b6f66d8671ef5186f342aa94c5
z197e4f59f2a6e201e62cc1f44386e1e1d84c584eb28a87e540e128cb41a6a5c51b1ac7ec491943
z67f11d4d6091ecc16210f03c9ac9cf5d1666a9f5fab964c8f48ade7f6b536387f975ec15d5ea57
z1391ab7513cf16ea343eef895b086c3b80b82f1635b5817cc386fdbfdca70f97b11a4d5418143b
z8aca8cd6b8048f8c4c7feedfe96d80518583fc83c4116fd6e53dcf4a50442d1d5d2b545969654b
z72337d3436aa0a59dcccaaaa38a1cbbfc7cd97d95b1dede38041db5af4d3a4230002a0431ff027
z507015b8805c6eab04f2458908a07031586d262273f6a51114d2d14d6fe215c6668880322c54ab
z87cdfd63ff66f8dec73fa1329355227a74367c5333aa81f082dc91188a167ef1473ea0e2f34691
z2ee5310e827d3fe19999052f1ca03c584887bfbb2ce5290b93dd281fe52bfa9fc2232b418d0f61
z426d0c8123d370d379b19a5fa74a50408ff9e329097f0a546c1074834d7e0a2c8ce83888e0a817
zad747fd084e4ebe9e0d4665e17a4c314f3dee23b555345462841c9e39a9203852c67a809a4356d
z68fdf00584a1034e54485fb5ffea53bdce88f56fde54cfa288803c77978168528d3d70c257118c
z762058abc2fa43f22e7e381052acfd6df6c312959aadd2f9b42fcf51fb683f08f1a2b019efcd81
za81779d58c3367620a3d4dda3bf1636e59fbc2e13521259c25e155158540cc4f60b0b435874e4e
z7e6902e206d7f89ec7b9d0da20a5bd1de1fb2976215826bff35b8a78b90a7b8307a66b37f52dda
z661042f1ef48da6c49410df507595f2c8779b1730427f91988fc09514b497391851363e85107c4
z14af4453a542c2a7f81a6a0c11f6620fe57c56c7df82cbcc5e45b401ea96280fdda5c2df23860e
z6b7a5dc183dd070dbb8095fbc7e6ade6ff61522e75a2dd7a6ff901141de36376351f53a95e9bf2
zc68806a99a677a4ba9a278cb01479d5e8d3d8dd3d6b4bcda2303ad18aa769df145cc8b59a115ce
zd73c77548d060e0682e9b70a622181a4b604372f8f63aaaf5c0cd96302b77bba63ded153a72428
z0a16c209c24d0bd44806b03d518f235320d6ad8a0f94797ccdd26bd74ffb1c99d04757b74d4de3
zb320c766bcf83698c11da49b0bdec03eb45b736668d6fcd4271a054a6834449ad4b0a101da5f1a
z47d12b199b989accd70a482f27e891a76c31147a386e77fc92e3303da695d65d58def6bd8faeca
z9961a64b8acbe36c8b42f6dd023c82cd1af04461673eddcef2db74d96439dfb485b23016a4f5b2
zd0cb8a7925d2fa84f9b51e418f5fd3cfdb204d25658608010d257d4f10f6c855c47660134c0243
zade46e6e661ae115631e75657c0228b187e920811324a668eec8b00fe531f0774b3c4048568210
z7039073dae63a9e78f5430210afe3e003ba695202010995aeeeaea96f04ae5f4a31cc9fed67ec5
zc5b775e9152fa4f5ca5abc7655892026a8fffd512d3e78122d6dd71a540cb86986f8016f34005e
z26a46c5b90d634b9c3761555149b816072cfd6e91dbd633027889f8a79c44291c24e14ef9d5e74
zc714c676c4630de8114d3a8f218e1bdba6ab914def83d86c93e5a6f78068d49207546aa03a54fb
z0a612093f51fe9e6f137f8b9efb411a8ef802d7630e7f59737925e135a4770e8e230c3a3693153
z04564bd4e07d648906a1ee3b5657f079fd34c6df3be793cd5dad9f6012ec2ed699fd0b8bb68e5c
z7554af7540aefc16b473c6fddd10397a7990e6bb126e1142fd4abbb8069e115e6f2b63c9c8c4fc
z05bb86f7bda83ae8c819b12c4a4fb082185b6506e137591790b488da848d135f42febdc8206d13
zf694e164b357a0cfe8474e581956e5f96070297b1b00397fd0c4fc4066c8d74297546c95831058
zb4c04b8e7f13b3a75b785bc720f7d7bc32982a8228032c46dc9775bedcdca2a3cf3b692bf58cc2
z41863deebe9e6a543e10b4e539c5df046f1ff8dd8955823ec077921c207d57fb56373629ec242c
zc6d367af40f80b78196bf8b481e9bea1e17fbc5030829bd55fdc04ccc5273904a3e3e0e3af3ec7
z959afb71809992d4916ac87a3c5b39c56da4867c10f8142d430a06f350eb2dc6f8315e0bf477d6
z3ec56cd1d2ba844d9ede2555faef5dbaf794ad71fb77c5004e5da803944f6bb89c7f4fa9ba9295
z7cb98d6d1d538ae9305d95211575697bc9fe686358bdb28b924784e3ce6531712f3e2a17d2e82d
zea3aa2d87045afe42a4bd5069d36cd97036af6e94b6c512246619bdeff48ad9e13cea84c7fd491
z6c754615b1d964c975dcd2afeba0e7eef05679eb6b1be3072f522c48c66d0576add55dfa9c874c
z2bd6f2f556159b0d9e12a3bc629ac12a9d3b70912add78c8aec3ffdfe9160132534b99750eb025
zf518073c5398404b49c6541af997d97272031aabcaaa605e5b7cbc8ff6c62a2d1ccb422b021718
z751415d6c9894318f9268e4e74ddb405232a9a50aad3f7f27690121d9eba5548282efb0383c965
z9a0956013343f6af00dd4ae53bc4ba378fb80a69477bb71166fead86ae06d7fc3972bff4918501
z50715ce9207734bdc1df720009564afaf064b159f07fac9034a2052029b2d7e03ab1791fb26214
za6b56a51251d5db898cdef622a7b2baecd2827ecdbf546193be04ca7c6985cbe5c9ac4f0d86559
z472ac1976fc3cd923a6be32ee14c4fc24bb18726738ab0cde63efc0f6c9a40c830cfe90e3cc820
z666821ed77af32490d8fea64718758ed7308285cb102156f7c9339e03e690bff0dcd6d5a2d6c83
zf137d97660ece188bd6c1b864aed48e0a32fd56a1c95928a3ebf9f64b0f245c418ce43be6383f9
zd36489b0ef7d3304392f61667b1ac183c4ec7fc479fd50f579fd71c21fe8a80e2b815edfed3f01
z7515dc1c78f7a4f701d5e55767851a43b11c9b116e964fa24bed56dca33c891a5b968910be95b6
zb14e6c34193390a5bdb8a0435f161b0873528e0def4831beb49e27aa2150d67e1c6c3d85cb46a3
z8a4d629f674c40111802f488ddffb4fb7f3f927ec6ff14434de297f386f7a0b06d963e895a8785
zfcc3df0c9d2d302d06787b414be7391be7dd0aad63d9216a10cab78bcd7d1c2d7f8e5f1e3597d8
z6346c83a12458c7d45fe8559f6b85458970627d6c25cb2fe1b191bdac16199f593aaba9b42d366
z940e11168e2eefde69f9a55fecca1bd2b3dfc7a9315bf333aa093f15fec4dd569d326660ad6a5c
z078ba3833d5b3aad298cbbd73a81f9eafd84bc8900cad5046bc2a2c8fe97c71d783ff7bedc143e
zde6a8428c095a4ae27e10f8a71259817d20a34c8d5c89c827b6c2dd769c67cfe4cf62e40a5af31
z085a6e450f8cae4397cdffc4886a7e28093b91ce85c7667a9d5265e0d81ccfdf82f74d5f2e9251
z58c2eae79c8b70cee10a29a825e553f14e56c42005605e2d03421818f7e9d62439b3c7927b753c
zd0819d066408ea2628ca9e304a738b0c825a7ee9f94f375356f426189d4022510ea4297b9fc98b
ze311d25828ea024fbd74df30f92dddd8fa6d6dbf1a0d713e9c216d1287b6a4c3c8f9f2518dfb41
z2395fec1de7c24eee08374a85f648f94c7d4c7868917df23cb1240a035f0002a3b6f8cd0ba4bc7
ze27108c084463ba517e790e0a3b9977199745430555b7be8bec3afdee213df09ab92482ab79fc6
z09e6a93c5219e28273906f7d8e410afaf620a6c39c345874ef064450b8527eecedaf82c07eb477
zfb15cbe87967e2c3464bbdd07b111a2a751ea84c87e49b1d9dcca65dc1d8a9f97b35410889044c
ze27ab7c86d85fec3131d61c1c6e451aae9a8c1cef9dfc06036e235dd9fc1eaf1aaddd51075b177
z4bd944c05e43e8cae6e83f504e7f1cc2b10280c63c2c5d079bd7420a3e1021e8095f80ff64a0ac
z06be86988c15b09ce9cea4508af7c43e19d67361c5cb3264f9075c4b921787323a021223fae562
z87dddf057c6bddf751fd5c497a9babbb1f283b6dfc9aefeaabe7b48d3fad1ce6d2c5156fba5792
zd1d24459b7273526d3d044781bcbabfb499276c9481b202edde7f5610dac4f8c8f665bd5717c65
za206f6160d7596a4a17943329e533d0a9f36bcac80d7c0c218297fa15fb3d45a9b3d178555268d
zc722d012537462acf3133b900dc411300105a7db15283b527ddbff6ed65af6c7c9729bee2457f2
zd99da66ef60ba8dded83bae5f8b3e465b591c367ddffceb162fe020e4383045941ad5a000b97d9
z5c7b191b0a9fb100d45105f2f911c033e407d40875152f09a5009672b3eed68c44e73559a592ac
z7c6b050560458c92dcb37cbeaa167b8e220f07f39d34b70e9fc71592c53d8a95833d7b6d42bf7e
z8387b710379b59ed436b1a81c685eaa6a5979d748094431ae20b8f7207f97fe7337ee145c28423
z8b6d007ebeec7b2efb4e89eba8ccc23f8611ef5fda743bad2c00ac775645ed21be023876086fd6
zc13567d69bacbd5389146cad1bf538e120d17691328a29f00928bdcd17775b8ba4ec62bfe94059
za9a789b7fe610c7ff5675a8ce3d02237874173ab855563027afe740b1ad21e90c026fa3611991a
z876b55a57ce5bb6cf16217c3448e9e1cd7977b73514a425f947c44d65b752f0228205d236b2f4d
zbc5ab24aeeea41dda75f7fe19d40a30e268b0b3cff7c36b7ad5f91674f6563d965beeb86077c7e
z0170f2d929c92f0ac89c94e0aa938661e1899ef324af3da4430237043a57d6ed55d5cd66b24089
zaaec4bc2b7632dea812030a4aa283cf8d8e5baa71d68a25d30e71cdd8da51c791cdc82eb573dd6
z4bb0282406105f45eb5e21934c298224a17d2c3c699a48f82b753f3ed5dad6ea1c621b49908200
z48628caa3e175932aa63195f5f55ba0173cb234718c54b8b4c2b306f9d9f8af2a1b9f9981d06a3
z31f3a7631ebe25816e556807be92bdd4d3bf8d3416b33b8b8d24bfd3bd226ee8fef846dea24403
z15220df2823d8a1a362dfc1cb147f51dd522bf63876afa406d1a250cd31a3d53cf54c4f5fd13df
ze106ccb03d255d30b74deda783390bb6ad4a5649a5d0ff4a528fea40bcc6cc54718f14c1401701
z7f4ecf8b105478253de6984e108e891f5672935c0e3e49c937e22e124a5fb4ed24f88008f7e4c9
z026c17237e292c9d243e03be542cc353ed4d8bb392029705b4726ca522b9d15491f446d0f0c3a2
z10ecd8e7244b06493c068dd4f9343bc125fb3c9501dfca42287d99d919a82e699542c7a6556627
z473b1b7ddd4adca76072062cfbf381410b0ce588f93c0b6ffee47a8c57e2d599bdfabae3f940d3
zf4a087b4c39f316f11617e3ed1ebe3801506ee4743fc5b63e45c7f2a584d637fb4b85561747bc8
z57f073e4a6b5ec84f8a92200fa451ec3b0fdf542b3dcc65a4ebae9ee6cdd7375a43af00276a75a
zc8f3157aadd238d947daf09a5347254f50123df097b7bdf445b5f3b574b09d8ca479e89cf6c48d
z61db448981a7fd080f4eae21cd36905ab35586ea15a8899f619078bdc120939d62c428c9223757
zf7ef6cb4abf4d3785c4f31d5d80270b6f1c4bca0932fa4f7ad96b4125d5871c51f55b14a6adf38
z4819da89d473702ed411a83362e1ec93bae7a53266ac42faccf4dd005a5a5be7d9699b276711a0
z927f188da246b26a9a11c0f8eb432f4343d79d3eb4797e4b6bc98012a0aa382567ab898677eddd
z344d9ce08a7fd2d78d6b03256738f1af8239461085ed9a1bacaa9c681e49cefafb8fbe645234c5
z31daf30fc455112c81e8d6ec64ba20e4c4a6ece2c395289d2cf7f061b480c31dc0f053081f5584
z61ad396929f989019aba40efefdd4e2b0fe66edf79db2c590d06bacc3a8b7654d1a2a8d689b6f9
zb76cc2d6eb5cb92974c27f9cf0dda9457e9a9d07681a5c229cc60aff34993e103d992190d0c1e0
zb8e6ebeba8900f635f4475d82367672a9aec17aaf3e033bbf1d4c12b456ccfe07972b622b02a07
z9ecee6c10f8aa1a0220d6894ffb4d3d4289291a1c05f1e4fe698eac7e58b53f0c72d24789c0e7e
zc22dd65629a70eb8bc2e7b8cde51bfc1f70c38fabe4b886fd3d594df58284ba252497a4823e8e9
z91051a668688186812e37b8b65031cd5eff0e0b828eee7770dba622b1cd36e7cfa74dac150e6e0
z061892a02d9cbf43c9b952bbbd67083e25558a5aaa97f3ae6415ed205dbaef54373fe2a9f98b8f
zc9c28bf3186c9d29545c98e73105fd6d02c7da130c5a7ffbdc58bd455f0b21c9af14d9761b7c6f
za99b2ff50957d4032309adaa947b66883f4a5f8da0ee2e18d4650d7249e853bc246ec883cd5dbb
za32ea63990227d874a9f57cca27dda7e9fd48775d810a6ac64c8078e196828aaee8cdd48236fe9
z00979154ac91ccc77c4af2d040ea5aef722dd587479a4c24e949ec0dddf6de49435c6d68137d4f
zd3717ccf2de60dae5acb624b9b47586094273636a09f27c6427941cc864414660c0270bad62a20
z6fd47c9f90b641a4588888fac84b6a680841b8be309cc18e53ea84ede284d7ec7ba5055ff611fa
zd1bd50f4dd43ab6deb9b71ee62806edf6672335da91e35452a211c87e3e3d00873efafd8f7ccc7
z1c82a6ae97f6fc530c7bf139db7fb280eb4761c2f32d091ad1214e5e6ce13f5a5bbbf4c5750c0d
z3e28ed33c6f23f6728a0726f892bf2b66d4a07f8c34383b28422085c0bcbfc477c311d26786e37
zb099eef62e914ca4b08a679cafaaf4d250d51758d023b621abb137c681fd86f4addb5210f0ff45
z7823b2e49d5e83f19fa41674ca68255c88b4ac3ec8e36dff520706cf50faeddc3625634f5cee23
z1e81d0c608e22348f1b009371742cc663302152b929792771bb1daf11499cedd6427882e3eab2c
zff1e7480bcb7b2e0e5c83baf5947ba33176119457ad4af59894dfb7478c7f8953c532c9b4bbbf3
z705612c5debd8933c53f0f13314dac7b077d5ffa838ede6ef3011623f9a89d2c440077499060ab
z2a279856a859380345a864e7ea70bb3084d29de0885907fba8e4487573ee87cd89482f69e7fa7e
zccc12d27bd6c7f4493db4656c3951fa3d7beb4960b232fb62bf567a5b933b8dfc7f463a9808702
z10a016b3a21bc2a3a20e89f0f32a8e1790d527e20c465d7e66e0fc68356ae464cb08a59b43475c
zf1154bee843d26673562f81bab303ea58df302abec9e90b89cc126c82dad49f03f2de197c0db7b
z4810aef7545a169231726e42ab5f6321bfa012a3c26ee50b02ee084e7a7b265e488939a899292d
z918588217bd736a8793fe71d4ab239619c41e95e2b6cc11b5bdf4425192ffa2239c984eb66ac41
zd5acab72c60828a76a3da57befb3d20f5ba7100a85b82b0d602f289c7c9d16f6e8cd3c7372a30b
z21253772c881892ecb4496b05193e2bd5ade88947de12f50e11de504890cb70220cfa94ad61fa2
z683937f62ce08002dbdc95ccacfa7e1227c233a9504811e7af1cc52f519fec09067b0f44fca22c
z2bfeb6724df678df5ebb2e8d3134b408d0a7e26700ab30c5007105e9539a497933df0dfda33bf4
zd192a405823a0a8b0cc2d014d95c43b5340e27d002ad15b6a7ea9a429eb41923cccb61b36ad08e
zed0993b6d304a148d85fbaee2b03988ea4eb852b49edd27a0066f67f50eb8d760b6d635f8c6a53
z4f695973d5cd14f22a760719ea1ccab96e0b5976b6a92fa0d7e2c53ac1d8ad3fedd60c0934efd9
z93db1eaf4a44c5548d88e4e6244fe10cece18ed8dda46f60844a67e2960d2238001b9d84d9c60c
zea404a106b7af2889eb31aba8ec49bcb9aafc6d805448f4bfaafbdf5a4396dc3c05ed01c4b1097
z8d8e0840dfa37c84b1e020f46ad150e379a649247f495b7352e9d9355a33d9230a4b164df7de56
zafdaa02d5f06286e5c385c85114e61f36d976fe2f1947d7f1ea803b02601006f5eb8a39a2080db
z7ffba8efba4b07bbb474e984d7d5e21b3f356c566dd072bd610f62c3f08d7e77d2a4696dc44258
zaa319546235589879b245662e2ee88c85c9fb0e298df087974b81ff72d1acd4b03ebcad381f205
z34cd0434b8c264943fc07929133c46652a09b9b8f7c18f8ffc44b06bf44fbcdd90c1979ce3bb98
z59bee5550e0c45ff07fff8ef36eb3f72e7b0926b41d1ad9dc08d0e5575771e07cda01920bd1e78
z5d49ff4220ba453cb18a2138f7227e42b91e5a582f96d27bd00c61747e18e27f0ca9bc6a53650a
z583035dd02da4a76d8382608c7ba93567131a54744a9523ebf6ccbdd83d202785e51014a6d86f7
zfdce3dde30ef1336cac33baf1793cc523e539d11d98ebfb85af40f7df9a825d4dcb9b94bb8edb7
z45b7147b91f02028816cd85b07a3d17f864a3c8e657df1e6e18ee9b52dc388a6da33c98ba021e7
z262f8f41b848a1490c8922c3b3e3a821399b0011409a0cce5cd12c694d21f91b12c511dda5c2bf
z021eec7f13b145d05c3a0d41171789a610472711831c413bd8f7b0ae8f42c31c9d1757b0fb47b8
za36006743a0edb72f658a16ebcdf84203ab786d721272cfdf2fcfb485740614dd94012981ce260
z45eaef468ac6b64233023583be06fe3d073dc38e3924e1f6dab5c426c36bee8d33ccdd75310d2c
z1f8f43e4ad182d753cb6327bbe5aa272caae2613617a6dcbc2bade0f72f698db1c84a521ac0b4d
zadf3813201f7ec531f2da87d6c8a048241ae0763e8ad634644612b4564c24d7681204a59c7296e
zd7a2c9bd7df869d7abe0447b98513340ab2f846f6099d5fa66d797ba8b8f408ac71e44ae4ea0af
zb782677f14873269675870d1073c350debe90588165c40bb485bb4c7e8eecc30fe9812ef61e53f
z734ebed2d97a907162298aa26dcd34c0678653cb8bf3f46a815cbc8bfa1f37fece9a9664b0c0a3
z4397eb0b4e1ee7ea4e19cf26d793ba17a8eea1d88b7b395a9f17b8d6965ed2aa072e4db5619048
z181402d79e1c8e3b03371e39b4738aebc8095cf82c048a3eaf85c1cd2ebac0ae8d714070d8e607
za80a6a47d1d4b0e15b8df6230c8cf395db456c3d7d3d29f1648bdfbe47a6b639cc5ef36bd8e4da
zd1be56effe293d21d789905bccdc91f83deb4a6744e5b253a218ce33f095b9f760512f8cbbc679
z0ba2636f634a8324f05e9dcb2013ad1d0251169605d74d9df4a6ebedbc1c2b2935e4c92f335e62
z079f1cc0fbc9c9109b4d8077634eea1335626d43f34e50b9df546640669fe337712a0b2572df4b
z26cb58b27f024cc848caf0a84f44c13e72962ee4d6e0155029281d7669a8a9ce86ac9221f5830f
z7a2ee400a5f2bf55fce2179ffa0c26b5651df53e2ba25872a427a833ff66532a8002656b939976
z4c90b096cd417731f668788e6c3e448af65f856db7d049edad5883f6a7d9c022a7186dc494876e
zf5ac7004f9e06e5f793a77e0e0fa9c7c589856526b7d42f20011d0c940f701590997fdcb0c28f2
z4dff074c987a2354a579d808640dda74d8df59edba43a16277eda8f650c70c202cc7d717bd1839
ze23285f516cf0b1a8873ff1322aee11276ed1d5987b6664adde113c61a27e1551413884940ee59
z5fce889650a44a5cc514b4aa0faa5a2630e9bd90aafe9d61ea9cc95fc67afa34b0d21a26c0d71f
z8abd52ce6fda343f3cb8517f00a87d18ad6c08310e5f298b0a11c7857581142e44fff63e1eb395
z5b691dbfabb0f4f53884173926f98b0815685ef969633338eb0e921990836b0d421810dcf3b208
zbe22265045e4711b51ee0e58a90e336d5ca8c53649c0b3344c7335281b85ba218111a8cc8cfc7a
zc1c51cb15b66d51b77f2d70c7f4b307ed4fbcf2ed546fc8a513d1721c74754b6ab468caba6eb41
zda8713a7302a4a1737c95a46f969865d8d863bb94880c48ddda98b008ed4e7447541e6a2be8f2d
zfa6c9346c0ab61a7bab57c32fde943c8dc83efa82c5d09d660e53666f50800ea31c7f1002c4d81
zfd6a9f6a6b49e84c45f13a95f8440d40c6ff78ebe242c37e7577a803f68a6104d46a0463687dbe
zf5171b168d91475beb859fd0b44aa6a445ec09109ac32350bbd75d086ce1a9c4a3f7bcee220a84
z6a4a78deb2af84abc17d4d8494e7083f30488586f42f161dc2cf61390b2dfe5b2dd6e95f0ecd16
zf482b02187a61bc7f1e41dfe86571594c00723f50f4dbaaf1e2c481d58fdc8474e22f4088d5666
z7a611c9d9c84e5731eba11287baa0b2d2c3ab1012eb0915de98aa60e8840be820b801aea06d96b
zb1e6f9bf6d38ae5ad8f7a763a93d77e07e768b685dc2415b2df3b7ba15e5b914ce4df2c39340e8
za2440ac03d82f25d118b1e9d52b9295091e05e8490154f0067dc3ac7d949b7de0cc9edc5902997
z1abc40116a9fdf8c58a85d2998dfd0bf762914f16fa13a669bfeaf4021f9598820f4068d192f70
zf754b93625a152f466a585eaf2ed676483ed8b67d5c406d2d5f514f69376dfd2b858f9501a19e7
z6914e3e14e47123fc13d5a4dc871e1d05697cd4bb637f3d8b20e7f185d8cffce16babc4cd33fa5
z702ec558c8ecf78c7ca1857bbc939c6f1ce46bee7294098e739696b1ed22b8038d7338bb030440
ze0f8986933c0f1eef58da75d05269d30324c076f2187e5f6dc98a16d8b9d2b12268886b93235ec
ze631cb343f68c86a51e41e7a7a05213eb7b173077f75fe95dff5b04825f1d98939d8a694aff5a3
z4bebf40c391984cb9005a9ec51477514d758d2b898064d9cfad2dea38ad9d9579372f809e60f13
z1e5ced4242999a4bb712069dee9f440a5c024dcee1a7b5729eb56278be00e41ae419979b726757
zb5ecd691049cb031ce75cc7a3393b320b87abb2401028398d8d1ba6e20ea993929f83d901da9fa
zf3c5f846c2faf36b1f8d3a365df6368f3543176c1afc1240329c561a28e03465923f9129429292
z41e3dfc9f6d6da1e3f1f9b8ce8d5d83f0d396ada36deccca46f703bb38dd0df33df787f7a5391d
z1922ccac8880f71760d69ba28a68cc7b6a726cf6a57cd0a8810fd170dbe2bde0b8c62207961590
z4edd1f2680eb0ec19b03ac8ab0b880657ffdc18491fcf838b1f9e37fe18994de64dfbb79b9a676
zd345459f259033fc47f5c71284340fff1d554bf7aada266a425db360adc261387a901213c24c06
zee2cd589116db5fc3b15286644046450ee855a9334167ed3806d75901e2e83a4d0fd78e5f6a8ba
z8ffcb6f5ce3b74c75148329144a12b54b717be5f76fcfe3e690baa1076518e5ad97066989d985b
zf7ce118c5882827934b5479c75548aa97f0069dfefc5a7759abe45505913f45f4f8033cf2b05cd
z90a26ab5d32a0df5b2430a8dfd3f0d5f597c3a11e734b89a6499eda9b162576c9442ae20eb5bb0
z672af1208574447c46d337dc62980e0cac07169dac3bc321b04c528557e810f3a7f89ad4c6fafd
z3c32cb456fbe5343225b5f228701e9434b4146b86ea69a615e4cdf9e2f0d4a7ee6ebe730dd683c
z277d6b75a21c135b14388afc67fe0acef640cad92f650ef44606da1ca115e972b8e5b6cc5e9f8b
z219211dbf4baaa63862b5668f19f0f002ba75739e1b61df549c498c322cd512eb1d937d82c24ee
z8eca30a8d758f0e8e62cdb8bc5e910deca843c624ab730395b02b3535688ccd381cb3cd43d7fff
z368372d223cda6aeb1ad404dd5f6539d51d9ead8c9742231486527bf308ddefb46a0aa821361a8
z1aef8b045994d2b5960c029a6391c1ed15bc36f97dc7e72fb36c0c219303f963e28ba340605ba2
z37cd31cc8792a24e0cdb68ac6799746a252534a720f99f4120467613e3ed341318ce48bb15e76d
z9cf7bcadf45a1ee67cf22ec3606f3ee679f7c3542bac685c2365e3151a77bb4f24ab2a24bb54b5
zf9e1c8ddbd85314f13657f443f6f5c27c23355716f4b3f3462baf9ebd0ec463df7a0e1e3333290
z9edfd17b6f067c402d0003f53ad05c7a24c2680dcc9c8db0678b6c348043749c33e5cf8b5ac74a
z14cc5131825cd4c23c05f913f6456daf966c0bb1552dc2b338d41cbaea9805d279b1c7db4083bf
z1f8782094cec14302c907f8754a2130a0f35f7adb3881649fecaa5f5cec727911107a9ee4e5e61
z95656396cd4455eca49307d2818e676351f87d9328fcfa58321049363aaaa5fa4f045e28cd18ea
z28bde0bcc77df8a807204fea67dc5d5021bfca62080f9f4390798296791ddacf20bb54385d924a
z46e06267d0d7664da944f1ca0983f807c4d19b177bb29246a857a8bc3e219e34df239bd4b77824
z9a927034760d1003184fbcab9a03803c4d2ea40049a6ae7437520ddbeecd89162e101b3ac27f18
z660f3817153410fc009b0e5701e69af193b54d77a322954a9ea03886a22b4228723bf859afeda5
zb43e7c17632b7415c4f22c771825c9e59516c2f18289448911191d0b9e0c3597e8fb75fa68049a
zfd3cc8fedff221c6e1c53a069313c396cf491133045bf427b79e967d8c70fbf7e990345e9a7496
z39c986fe2fc252748b0867a20de3a1ffa5d514d61396cbc01aab053d6515e3086eff75fe3e7ba4
z013f80fa5e6de751121081809d5d697040c93d4db389f176a767337a83b319a7750e8e408c0931
zaee019289f5750cbf2844475d14b4831c1bae29931ce878a3f48402d479a2e938f393839a41e02
zda977b8bce18d1c2cdc2cd140f266fc7d1ee46e4eaf8651332db94fdeb989b93bd27c18216aade
z147aad1d94ddac732f3df9ac22b06c0c45b7b70b34b8fb8204a4573bbe671690b671fec78b468a
z5959c84b306d90f6b87f9ab81d39872294c19a7cee6230f8ad3c0a276d23a0aec00512f385092f
z69eb0a8386233d6062cce0e9d1ef18b9cf3af58fcb2d03642eef88ff4f9aa1852144880393c555
z35868fa2b787d6957bd74ca3ab886fd004663f5c9c7ab5d1a9971c63140f265f245798d5e2ff80
z7d48a702a7f07a366648d1363a0ff2bc031af8266fbd0c6647e3f9d6cd7a50062f0461b1727e1c
z96e0a33afc3225473baa345b3f6d79d0303b810f8cb5959e28ae4392aee664aa61bea3687d27d3
z08a85f71f08c9c71911a5a0ab4df6283a5e937f77bd425524a50bb245299feb3ac8c82f6f95c2e
z27f0cd3b9a78a9e82cb0ddc8f78ea07506c2f5ba04202ae8e2a4974fb5305f2c6c6bae04ee2671
z79fc792958a2b4a2548849d8fcba54bb0a0932e295f57918a993cc403651927d89ab0d9505d714
zfb099ef0b9075593469eb5d309927cb91600030c942f7251c5fe922bcce2f20603948edfd92a70
ze73c70299728b1e2907cd7a1d76d0c16b712a1a0b824924e5534726492ad0a7eea45a3d4e2ae2d
z84f25cf6582cce490c42ea3168eeb00645ff393c7c1b3d4e373ac633371f1f304debbcb09ac6af
zabf1b08ce519e3a7c06083acd37921739071351f56093586f143ddd2eda930828eaeabf04014b9
z3eea4edf4b706f4bcede0e60f2984984870c2c780cb87a90adc45e71985ce55927c5799e418f98
zfbea3517723b2a28839a690dd86ad5f3953913f9086516522f2ce74e995f85fd33e59a5321385b
zab4f2739f9c37cb5885f281eeb60b99dcf3ceacefda8e8aaef62d1213a9d71354fcb68ceb70b50
z5f6340e41402a96611990f39fbeb60af22c2e90fab42744cb2c5bcc5d14056af3e2c01082618e2
zf436e675d532b8eb4d51a9808609507019c483c1fc08261e6c3c081ed5500559c50fe23772d86e
z3d3f6074872a0cca4bb5e433ae06770b7e485a39a5d1ade26015b09d592c8b8e4bdd3f3613f475
z7c0ad13613f0ea42acac1cb407e8c859e12fb917b42be27b4d319c3a8cf07028fcb1fe30740501
zc40b944068a953cec25ff2cc93408043bd8a794a75d535033f50a34799a160d8360a2978664d28
z252f569779bd49850a9f7ffd4fdc3f7f6e1d2633510dd4cf18ffc3cf2dfbd6de0eeaac13289789
z80d2d2659b16b7a8cc72cf2c3546c01498e44bdf3119234ece3ecb52ab18ffb780a7881f84257d
z3688909742bb98b43b162039d4e3b2821419b09e0f2b2aad40781920ff090c2c5049c63ccdacf8
zcaed7894c89d76105e586e4177f58929dc2f536cbab654c28088f267e4d10ad61097a1d5d0ee86
zc56fd18d06d84593993ff559ee2781c1e9d8974f8483bb39ebc147407bb9faf68bbb7175510361
z720e5fa3f49d3394c1704de761624b3b9bddc5e59d32de67980cc153394c7bec0e689040df66ba
z9c74710630daf12ef27ebf9214bf4282b3af5926fe6fe6d24cd44941afca63e8d5906079ea58dc
z4a9fa695c41b3738e942288bfa036791ac332cc4243886a9c12e152bc684ac2a85189ced290479
zb2834f492dc66976779028cae5b7953ab59881c08e57eca8675ca5aef95ca26491ce75af4659ad
z048b573aa94ab0ea4333ffb6e99ac62db1e7f0e14229c90f1cf08b69fa1468b200e333e6669188
z7e5ef1299a0f226b99685d8779b920959baa10126baa2b8cbe5fa0841ae57f09da9b27f41a0e64
z82d7e8e4f622b4b64cf710bd4009dfde651d2505a00c1adfbf709c349abe54e5f4969fc7a8d9a0
zb3e4f0cdd747e9e6268dc820d0cc59b957abe9b1ce71b37f5c15cba76de0d8cf62055d5ff44904
z1b6398562eb90db770b039f2b289ac788e5d673544adc9e04224131c8019f24419f38de0716d68
ze09bd092c01257bfec1bca6ca45692558bcf8b7d889f890de95f93c185841f174d1adcca41b419
zcc53449c1342b532f014db863d982da286c71e83958b49e45f02b93c3413fc7f6acd840ff82862
zf22d1ba4d7fa1df0edd2ac62ac6f82b7d256dc257f8718d540ee19382bad652cd4fc0b6aab1227
z1bc97baca391835d2cb7dd4360a01ab983d2f1d905b96b37d9866d0fd4400eddcb43b756abf7a6
z115255b3b3fe175566be09005dfdb4f94297807e8cd114440087d19743e5254dc0bad559bf92b3
za879b6cc01b950ea9a0eeb233c9d10b933f3367ba74644a97b350494584d56bfdbedf685cb1547
zcd5c5503359677353713ec8e9bcf370bf78b02af09dc67f97c73f0a202e76648aed11e5dc51728
z5e5394fc05b4288baf750464139dbda05e2a07321f1639c64207fd40ab3a27d1965cbaa35548ff
z738c2ab5f5e74ed9d1c0d3da5b2b8deebee161cd139bcdc37aea305faee21b36959d40a468c5ef
zf5623765d83abaf276dda78746929b66849c9b9eb7eca6d559e35077807846e34d179933097331
zdaa82ba86563dd53e53fc4d3b7936e0776ab569853852a227e3c7942825020f5f7b05ac3239c6d
z3cebd10c4e23f4736dbec9c3814db043ce57ac5c1486120182f1a40247b0d578369593df823dc0
zdf1408e7a1545eb21f6b291b2aa4c359ec35a85674cb63b768028b8044777d2c7cff99863b219a
z2953878d505b9b06ae2f91755dc7e204ca28af58d02b669aca01e8f5ead79f167a29ade4ba37a4
z76dcd211648e288ab179e2452b995504bf7e72828977231fee0723cbfb65bc2d8d5e22502ff14d
z4bafb94cac276883a29a79dae42bd3ba6798b359a71dac52d95585ab19bf27140447084342b4e5
z465fdb3293efb5bafdc091fe5fe6a28e894186e7ebfcbb92ed2f740b5bcbee00f6e0450a733f8e
z85f2d54f17f5c9547beb8b064d31a5030f3bd36355a6f7e688cbd051261eb010d6185c08e3b910
z981d3c67761f167ce0b8db63e33fa938e6c00592040fa56c3b775283a82f7a0cf4869df0b19c87
zf3e32de8b25253a072b25b18b485f9f8b86fecae918974b2998e45b9c56f692add7aa5594cafc7
z86ba81b6973617350340340bb1ca49ddfa72c1891057c1842e384a5b889df70f901dc1a9283c9d
zf7541faace04e11555b5c441813151fb638a40ef1b08c8d7c9d39d1354fbbcf77af071e4f1e6fe
z6aa46b3d02a78754dfb665d37dc09bf90ab83713a9ae0872cb191f66b189de78a28db38ab80717
zaba89869581318219e5c38f2ae814cdb0461e3a78aa961306b8001129ebaaffc9a8f693706b504
z763d588b63068aece8064c4dd6f2d58bf38b7b8d3e042f9cfc01222b4729bbcb1f6ac0132e1a62
z2bfae3999428dcae291aba185a6175c26ea655c7d27162e41cb50adfa4cf18cd6d2915edc0aaf4
z6a65657f261220128b87ca188bb945c493a5386b7a073f49df255ee12bf5b2a2416bb07e446a69
zf7ad2fe28fbb1f42b64fc1bae60406c7b444acdc7b9444ace3b8b28e65f8c81cc12a01b080cf05
zeebdd6734f7c23dbc41c6a1ba27da394531554c07aa356f3ee9d81ecd6c21a3d54fa348f44e10c
zc3eb760c0bb2b6b1d6ab4c260d9585ac449b3b08385bdc284e88c6de7fec7246a779987809d0e5
z0cea0d9452a4a712ebff34cf8db1efe3a22a0cc4d9286656ca726714338c12634c1d077976b273
z0e7b3ba1f35612e98b3195e5224d6b734596472ca2b764012758b9db2095cd4e8c20c792db5164
z938307981d217ebada4c89748d20900acb7eb92f47376e253fbc48b2015f403cd7f0eabf5d0950
z2a3df07367f22c273dd901aecc93be42e0bd6bfbc3e46838144f4996cc807428786488308c1b30
zd696326f76974f7cb5c01375c1f67fe924f1e0685c0f7c7fcb5f0ee894ef5ee89709c5e8d7ca2f
z3af4729d47075e95db6e4f85089618f5e664effaa3eb9a075c8c40ad061fec71eaaea7862e7752
z87cb14fc4ed7255934ca268cbc510c4f6d702d0187abb5e45453eaa5c4e00ea4fa1fc791f117bd
z69aec4e3e827500be355495167c27e0ed68cd43c1acaced3ec7ce3c80548fde1908009e696f25b
z09e7f63327a4f4a50ea63a34ab291cfc5a7c71135cfb2da5b76246cfe51ba1012ea58cf523be9b
z69b8e3753963ea0099b192a2eb774ea90b57fcb7d5f5cb35b8258a898202d881c6ab4c54e42d13
z35dfe098e0d9e1d8390edaa26c448afdecb3a428de9f22f1e2dfc79fcae918fe099c97d95cbdc7
z1dc7f79c359100d17852278c6def31375dc9db62b0506fef43fef999fe958c3297f80cea4c1f02
ze0f1e2f4378fcfc80e2acc1050aedb9108f31c2f5fa9c216a1043a0dde669ef9b3d3953a394fec
z0cc6d0ffa7b2b39bb2aad1a1c0a6c6391c50109b89916d1a5782585cff299f19bf0df91a2661e1
z3ffb81e1d1aaa39a25febf37e72770704defac06ab77d3c653e30196931c27a3aa5a299f11755c
z69eba022e63b9ee5641a06c070014e19465fb79aea5113384cd64a558f28fb49b1d7e7e1ee7afc
zba4ec11e1fc0097610d6881b83684b8b4696213628a146bb879bbb3a2bb05897b5ffc491a1801f
z48ee699b80836598c69cd5e2a2b274403253c0654455abdc871d37abd60cf56a068926c2c40595
zae8a0e0969ea8137f216dfd47f62e2075a80b04f73942e83c004956d74d8290b1f6921de74abe2
z8fc36a8764c3cf7bad65607675c8afe721dcaf10caf376616726d7029689f27696abe0de93e8fc
z338a53f5c00d50bcc769fe6109b7d65bbe684796313738d98cf043c4149e74f10fdc96972e7289
z8dfdcf0eacecb628f8d3fb2570da14d955acfd2d87eda08749d486622c2b5b2b7357c1f18d220f
zf5a241d4040d0502fa3ae77e21785b722cf2296ee63d34d9c34ac9827af081394684fef0563ed9
z459ab410ae28d4501decd6686f25bb6684051fb6cc2b27807ed0054d95ab8628ecb4d13eaa9dc9
za43d45a02477f5990f1561aa8d229ffe15a50cce80f44a6fbb0a0a71d896e17c8c5e9fdffe4067
z70f27c85730de85fdeede377cd16e5b47e5d4718158228c25c4ec14fbeaef70fad064ede68006c
zb240f30d0f879b21403a086a781747d4a50064d5daa923c96c7017a0db216e9984830f3a9edf19
z8b5542b83c21a0678913299f39de1a83498499ed0886b7fe233b85a49e6f9e8d03b67d6526d99f
zd306363ead3d9e81335f9a0047c6845f2c29a6fbe9fca83bc559434e996e723fcc764fadc1b870
z7a21b8c1e14359f9f483277579ba4b85e77354216688fec6c09dfb028ac2d52004aad8d9e4fc30
zef2d9a7999b34b6b5a06141678e7fb5644bf8682a254ab966b0dca8e1fb48ab8a35324798a0891
z9608ded264fe6c4119c7295d7d6c34d4dfebd7460590abf841008dd54bf91d63becbf86dfa3016
zc28f4be5d55bae6d10f1687d18539660a8b66c06558059629e709b0fe22f0a3392fc7787bc9628
z435a0d605bcfd745dd8fd3729ee7a43642136b0e31a50b2537460a6d558366642257d748f83715
z8650ebdd9906415867959a2a895d854ca7b1ccd101a29b728bb34b68c73d5ce7d146ee0642402d
zac5a0a772dfceedc6756a5e7cef00c3e5d73a164c11cfdfcd419ce09efe3c5b0683e2346c47164
z648db558657dd9f2c6b09d5de91087843ffb41ad09e548e5306c9f6aa27fb224dd1a351d50382a
z0c0fa4c3f11623d42bc6842726abfb85494930f4bbcd50c539809f6c3bcd52f570548d0b028034
za460c0cd9cd591f0fe9c71a6396b62d686929349e6e57c68e8bd4c85d1c07ec198546cad2abb37
zc61327281609fef5e815437403fc4b003e7d04f953a9dab5b3c855c0bfb0e8b89f65bcb0864024
zdafc16055e91b4ddf24f1b8e10b73a8afef4499f5fe1f0eb15ab3f8aa49edf059a031a96fe9d08
zc9729b69192b0956cc977363a23ec739d19a25cfd074ae84675fdd9968f4740a828f1d9cadfda1
z56826416991114bb6691f93e0657c73585f402b7f41b4bd228f0e2b8b1934870bd1c4298f5c961
z250811cd857a43ed8dfd6e758d3cfa0911afa10fc9224d7412b9f6b32e812cde26c5391762be8f
z8a4155bb9a69d4e0416b394531ca8ab79041c0e85eaacce7d4c5e836fdbaa7e58de96f3993ed18
zb28131d5869e66f4c6bdcdf3417731f4d6053e829fe22c5a5d20fb2ff62791a4a4ae0e15197924
z6c0a70376c769732f52ea95ba24b94ee0b00b027e679a560a1d1e3a9339d265910c932433b0f3b
z370f7c24c070933f38f49edf304d8bc8cd78f9b52ae265840019dfc72a17c89b8836abff6da90a
z1e24feee0bd51b128bdf4ce96013a6a85d415896107c35d0bfa85b5b425635f4059b880c74678d
zb488690371d5985c94979cb6cd25c5df9746e65f4522839b91a87a8146b58256395abcb0bc79b7
z6565aee49e0adaefdeece3fb465a929e2838521caa3068a83dc6bfd4fe2b8463ff2239ec48d431
zff8a7eeb995b8597e8af52e1cfc16073e13ec9ff26cbcc45324f7e42298382ae16ce47ac0ba162
zceb05cb7d8e196f74fd3eab56831177ae46b42de95941bf35146a9fedbfbce534c55bfeb15a8e7
z08366a0f5c8b6dafe8d3a3d8f5f5f32386d4c500cce2ddcdd0c2badc6250bba38712cadb93c134
z7b1bbfb7ca5e0207e2b4e116d9a9edb36ecb01c9ffb1051b9e0fc0b41c0761b6cfc97e85f8ce5e
z985ed15b386abf809e8291b44afd7c95e2fe46f2fb96345aa7234d2a151e6ef4da58435f9e4a3a
zc622fe1f7551e4752b9e72b4240711236fa11111c8da291032b9588bd486780114dae264971ed0
ze03aa7023b595fc5c1105e380948e92bfca6f52dfc7e9776b483a5d45225d72c824d4ab8b40128
z790aa0b1dbc3932c88041ebd02e7ffd78b9be28a59c2dbdaf62e6fc2257ef81009ff62601e6296
z60cd7244b9c5fa47895b7df479c253d68fd76591b38fc05cc255c0c098b758e1ed59b4698e7c94
zfebeb424b6317ce841ebee16908495b86e86a53a842086e040f23c986d40d4b76a8ad3142b133d
ze79877538ecad4625c43ee957f8394de365f1d0ccb74bd217ef044bb182f4481edceefe18b61c1
z0258d79228083eb1d48fb85e02a579658c4e2fca4c04071be050d9479aef1b9fdc548c5160b30c
z8c0dfeefe2697d244b8288aeb0cd58af2555c570e1fe02ae0a3c06fb15094f429ca30201cc1b44
z2b2765abb76bf88c98734dbde9f9080f4dbf2e38f270372627391656ea7910f08ee5a5005ffd58
za22ba8b2bf47c3126b600af9f08be8a3fa849bc4869dedc837561d49becc9a49a9e562e77e7523
z059b9857a1325b716c31dd9dd0db73a3304e441e2f3ca087554859c898347a69d54fedfe74719d
z957d65fa881b61cde068f9a27406a4891aca553026644d4a60a2c353bcc4ea42a630d24a3be356
zbf92b18c77c7683d0bff654e71850d00286bf2235e3f9a76d049e65e747b095a7a4b6bfbbd0789
z50228c633577c0afed3336d865273d11fb21f3422d2e07a2557483a142340693516d7889313c44
z2d4de240e7edd23a9f73b8135857bfbf94d7a37ccd2d0fd1aaebdd9fb34e9120cb6e5f44419b62
z69107ed82f6cdaee00d83aa22ac2f46ad10d995c037234715c2bb3ce18385b46e01c3d738a56ff
z1e97d0b8b3862137725ff1b4c9e0a86644d2188e400323291129747bb49117c051b13ad0ee084b
zde980636f16bf76dc9bb0c4c27703afee2a8def5049db06d52650b76be6710350683a52a078b6c
zfbd962ab7db83d430c96cd42a222146e893f0fbc683ca8ff2e975cea5862714541dd197036d9fc
z358d73a3276dc0d3cfb1ba4166ee2fc1d8fb4e923f9f4e0c3cb1f6a8544d1752a23387908b3238
z697645b2d3439a030a3fb6271df0863d705b8b95f42cf777cf9e376356a9caabfae9a8188602f5
z89a01ce6bdac2ce293553cf97c1d0bc92da0e0fc310ce28f04bf309627e0103557f774cd013f6c
z520c4fec3c047907f5dc4d997377e1d65007a79373b3d3e6425d4bedb33978530479832e1d6d15
zf21035510cd59cad428ad697f38a0f314c5e03896562f0af06a1deda1a108de7c06e05461658df
z332be675f5c984c69b9d3d146edc4a998fab0d7d7933e2f6e1c0b9941cc774d755b2caaf5843af
za6738adc88576a8d2572773c1d657ca105bc460226b23ff2d5cd0361fb0204c3b5ac68136c7137
z612da8de37632a6fbfe36f10551f3f807a7c8c8544d6e84394110846185452ec3917d3ed457dd3
z34a149c29953e499906a97102ae8fbfad4daa2c060b8d613d3c3fc77e0b2215f17b7bc1182ab93
z06f512df819315d777c2bd054f8aba145ac6e0edfd72949fca2745a8efa2f57e68cdc1ef7a943d
z331c06207a826190811e54d594b30168c9f27790f078be1ac615c0c39bc74812e52f64ccf6e0f8
z4b67020af06d00d5f5735d1661bf277950c2f06491dd3ff905c7d5828f879d8170e82058fefc49
z78e8133ea98c2596c2931219786a845b400e3297cb7ac117f5a3182056e87c0c1fa2a01b9ee34e
z0785bd9ea305dbeb73c069433d7a8222ff38d9343d35942789ca7545fa33196e6b5e048e35a353
z0cd9c55547585d88b60d9be350c3550eb04717863e10da638ff8260499039cb7faaca49f45962f
z6577011da1d89ed740480dd8a4acf3c16780d53f8aa758fdf860edd97af4fad543fe1bedd8ef6c
z3f3e6109a029b5b08d1c7fcfa67665d22db6f9652f4376d9c80566a48d7b55d5c19faab74f6887
zba6203676d9b2f6e8bc34ba223ad173f4118b150e65ee3375d99a5418187cf3019b91eba072883
zbf23c075dd97b00772c2fb5e0c3bf84245d99d695174794f709ba722b7a5e221ccb06eff5c7dc2
z44b43697326dbdcedbbed7483ba88ce790d79d9d47c8bb6ba35be121152624389d65155b359eaa
z97793cffa5f16105e2d6099b82b362f24892e50d9c465a953f650395d1140440fdf96b700cb191
zc4e5bc1954f0be0a883dcd0884ba10e3b5f9c4d1c0d19cc775cd4f61c4b3c2b5945b471533e67b
zb07f2c002ba27d8ee02a82fc973ab28b0443b2f37dd9bd34323c80974c22b730d53acad20b7db7
z4acfe284bfc54dc5e6b293f2f5a85b861ae593bc2ee340a8693d96e091fbfd1b2100008cb79da2
z0cb35120215d4942f84cb2636e5c622ae871b5c2a1fd91870649dbfdb44663e50387bd31892cd7
z90e6fdf2f3ab816ebad234d93d02ba705fd455560a2ceea42831a829b9f946b495b2f7fed8bad9
zebc381a04f6fdeae1ec0e797863bc13f15d98f4b17d6c7792ec408ea200d64f44818e8e0513cbd
zdc52b61a1ecfb0ac3016a5d0a640ecb575cc5c21a7daf28a1c88837c0339ee3e3754d4d7a57622
zf52851c0315f4e39b3b358b5fc4088ac887e0ad9be12bfcd4f2a75a63bb22529e03e2c83dfbbf3
z234fd0e4b0bca5d71f54474d285d8199bbd4a1957efba330ae31fda47a8da765e0e1fb05e6f71e
z0698c4000e2ae65ad016fa0f09b1d532d20276602f926a635bfc6279f0104387d6a9837ded1fbd
z467d31ef3ad857d6377bd112d7ced45c3b638ef3245762cccf70d3648461246705bbd48d4f50fc
zdc36990b49e71046d799a579a9dee05adb8b87aa00acd1f35beceb773aee293a7604945291994b
z711adbeca279d6110cccdbd1110ff16d9a6bb2c9d0cf9335cb25f333b339cf3305e458dfdaf72a
zc254bc49e81539a54e6fbd35081590f50ea2c93a610b4507fa4cef4a1397b1e1bf374900fd7d84
z7bc4f7650959d51046a93b6e6ce26e1ddc2514563c20513969a4afd4be5e7ea40b226e241b1088
z8fd7381b14ddeb8b1b2413a388233ebbb30c38cde5aa5b9ac983e662d503fb21230b2090e241eb
z1e4c604bd0fd47d48f157c117de279ea19ec52b0a0d2cb5095442a90151dde55436118da3d5986
z4aba9050fa714ac84fa106b0ee8996c3dce21765794146b03bf0f1f054d34c45dc32ce24ecff55
za59f1103441fff9cd05baddf5380efa004ef16816fe42bf08d16eeeaa413f74787eec53090b8fd
z11145ad804d79a22b65081074a337450d44e6a20f3889508642244cd7d10b4bdc64e018f9c3a7f
z83565e5e7c9b0667f781e69d9912d763a33c30db7e87cc6b0422879ec295cb03d118e3eb7984d2
zd95a1495df9f03bf0f3b131c99192dfa98054641219be779bf9ac0fb564ed4e0b52f80dcacb830
z2c06860894dcdd8fd000b09aed4edb9992ddcaa32131a23bef853585e33ebc7f50977b59eba67d
zb8c1c2b183b23ef16cc53d5e3f15fc9f5be82536540ffa55b9bfa4c8c01af725ba910031c060c7
z7a224c3c0d21739e57435e1db895c36a2ca0a52a93b5ead56ebd7e089fb3e61dd01248fb3074c0
zbfeb3823b17a3ad13a18c1e831970833c4925f756f7db6d21e734a18f280c1b8a5b75b8384075c
zc7091b957ff8f729743087547df9f29329cd41eb4629de01c370f9e92c6606fea31de60ece2863
zb67be70028512abce6cf25bc74eceeb543bed791e597fd85c52c3cb5be9bdc3d6c93c4c7add692
zbe0f6a80a1d379c901d70aeb84dac2550b0e8a75b98abd6430691918977fd79f1bd1182901cd0f
z435bfe5d7db7a901c14978b2a0862e9359b26d97d3d4a8392e23e4f3ca8da20ee0ddde43aaf76f
z1ea2162849a31341568eacc5a385f8348a0088ef331a2cd41d1cd2c3fc7ec7866d53b5ac6281a4
z2c0fc0e89118edbbf614b6c6f9664900749fe1ab335d1dd2292740b503a90ec4d06a0a93be7aff
z15e581fa8b79a6e016164fdc4f93d19f94f7162af08b09308d76a85f3c2db17306ddd69236c44e
z2a91c02bfd40b14ff779691cd919fc14a03e5ba49dc6e817ad27706462cb5fcc488982b8b64c22
zbfc6412f4535b890f51a6c530f1ecf997c12bd4626319d37e72986e15fe7c20b4326fa1163e1bc
z5d2e4476282d3904f485c26c27dafab99edd73b545e72f93bcb6debb5228beca7203da8571caab
z8517f2465b96d7ebce91127aaed5fc3bbacf548c41b72bba09d6b19398ea5404cd7a46a06a34ff
zec0c890a442c6a0283493f2dee236048f092925b406c9af78b74721ec98c49611814dfdee71268
zebfe51cf9fe483a6857cd9f7176b52a6ee2f52816e8b287b0d96f6975d2ad6e54e7f274e00e742
zc7643182306dfed5c194a0c00f8bbc348ea5e5ebe6af468812bdaa857fd6043f3fbadba11d0b26
ze9b333af71c9aabc8b3a3a4979df11ab29a9f27cf4b6ac936511b67cb342bb303ce1b58916a84f
z35bcf98838d39f6d498668af4b9bbe2b347bd885b7e91d1d6e97277ac6c47ae0495b23020d74a6
z6085dad8d12ffbcd378f82af88215184a4d6d9d9f07f996595346f737dbf6492b21e9f73183fec
z7b650072b1dba8c31b5e1508d8ae10d71872515d3f199ab12d8bdac51db91e15999b0d6dd5a137
zc1c3c3e7d09fd48137c770f4547ba1860c6b73b3b012e6e27b17a325bca3a198045c39e6a93a8e
z773681fff6ef0fa2c0f07292a8a62bf2f5ead6122bf93358e1291d78ce7c300ac1878a811ffdc5
z81048fc85ed95a4c52fd7dc0914f1ece89e0da3db7aac16d8bd7d4d8dc1aad6e2b501f57cc1f3f
z510eac32e6d51e0aee37564f75d9d0826cb38320da22d55e44cc78bf8c031eb62160d0a456c80d
zcc534be8eac036f8fc7e8a1fa55bc23597e252aed098f5c91076543f978b4c125e52de752ab063
z368a5ee470d910070ad1661ab91a0fdacc7d37f73c6bf38c42e11cce5110056e2f46b92a97549d
zc23be5fbba0d4a014df3f5948f3b1941a46d88a0cdc1c689f467e7a3116fc1d6ead44de539faf9
z4de0a2760b764d8f32e18809c68279ebb08a59f68731d6207f5d8b4ff8014ebba5663f87204fa6
zee21be2dd6b9c3ac800066990e6567abb1054987fc7e77287375e2e52bfb89e660bfdfe18f6fd4
z6d6206eb46c13a9fabd80a337bb7a4b84216c93440c975039a3f9da9f9840c282802987aef5710
z6ba0be1913d6ca1f04b57224637f7617465f308e38c4ab60fd1873865e3664efeeef1fc93e3d5c
ze89abade245f99d17aa3336af29456bbdf26e5b2cd5eed48c876105dcf0b049b5c122fad7303d8
z93601eb36091e5c96e5da85984394eb5892b00c16789219aa636e14919581613f759c5c2c6abc0
zfcd990202007e0b71b5d6f4478571bed3ff3919f2d4e287f48bcab69af9028402cbac4c3670bd1
ze91b3f47d71da0d65220837e09f4a86250d052ba8010257b8acd6558dedd01397eeb2ff782b90a
z35c2df2143c2df1a363c26eb74a080e1bb3dd8f889970b2eb384f9cdf804c1a5d0439bfc9bb54b
z1f7273418e402427c21fc13286b15d75afb42282e202ee32afad516fac8b54c41b6e0c476575a8
z8a191cb7ec342bc22a7b81b33a91d09a1820ab9a4c7f731961626da359ccf6be33421e1dc65356
z72a4a9fb91133326fd928066d703047dd7d64c7efb04398849ba3371f363976f52a9133dd27f89
zb16a3363f93f78682e85132d54aafbc6ffe7d849f68137a736f45af27c319b1cc759d9d551a8bb
z4add0766f581fa6c00253e626c1df589aeb23d62046cc35869db2668fd2e57a2cdbd2a7f435b0e
zef33e5a29f58d649ff0d38e853f7310646f14eea909f07673f35e637110da0e84d24b30f7a36f0
zd72ad141a47571540d18ae9a3f9dc6696b3ff0b8437add97c0039d668a3507f127912452fc58f3
z738a9f69f727f1b862818d64c50a0e2d09479cde8191aedd5fe4499ad94baa26efd09c0f8ee1af
z47304af49561847bbb2271a252e32691392cf6a39a53932ce2080382d7d73b30ffdfd055ce4916
zca0ea7aa3ba11341a34c314aed72ed7b2e86a021a57720b979339bddb851f21dfc1adeb0055cce
za3d314c5900414e2ce9b286717672090f2a690123ee0b0e929f9b8c10b36db0b0a7b52910f476e
z65b26b6f7e06a81459550fa8cc7a6825754858edf9afee86d5910913625ba5a7d62af188b44b0f
z17be44598313f35f517028832b69497e420618c2c79cb6ba31099e69f2079e352811873c01c8d5
z9ff3ed4cacc4daee9ade2555c7f43634b8be4de33f23bc79ffd44af500b6717579c9922b7c9249
za09ec872529b91e645372e4b41f892a0dd4eb734d1d19fc233eb448b4620be7e7fea5236d1dec8
z37a85addd92fd772097d8bfd0dcd4f45e290030aef58a1fd2bee4ef5addbde7e10209706c1c3bf
z563b7b5491e74057fdedfb98170711a05f1fd207f0724a8d0c2be54881bbd570b7d05bd36dc804
z92797aecb8b341342edb4663353545cf4f3dd8e19708733557d58d566000c598b360c8f210d96c
zf0128467ee2badbd6e4ad4ff83bedea0baf4422461cee59170d6c3eb26288d82dd56012674e9f6
zab56dec9f30be28486892a9998650f161478e919f7c2dee049de2db574a31540454fa01c2c9f04
z9dad56e5ae2c7af7d840e0cbc801bce4544042e851eb247c4ecbc8c49c7686019ceed141a3bcd1
zbe341b49b23417e9ebf258ea714567f824c5bbc646a532003246d631012df835ae7b4589a4753a
z40afedb98dfdd6bcb45ece70bd3b665eabbd304ed820cf7c6fe610110d771e853f8732ee16fc88
z46a8f561e307e0f00e8c6b083d9ee6f51fc2383256439eb2100f058a683fb3fa5d04893ab3d571
zb7686ac2cf30dd837e8490f5921de1fb25e6fd3485339f135522dffbfe636f516c76bcc1457617
ze60ef5c40432d3324c75ce62254605107f64244bc16e96824d491d4f493ef4edbc311ed68371cc
z8a4a9a0113b5fd438acfa2959cd193f28e918b85c24154b76670742ff12572033553c93c09c492
zf7bc3e58675e662a553a61355e9a4373e5b06a87c715398d72e86c30112547af47c8f913660519
z07ab4a8bbc8b67bb3a182850152c68e17404105d229d9ca27b57df95b4ed725419ba485420bd89
z25b9d6ce3e06279b8e85bc1245f34889ed50b9479c489927b750cb8e05e90f8e8ef100008726e0
zd4faca758071325c7cfebc79d59064f449c9e915718bd57c4120311c373e0eda6a8abafa144882
z9581d4ed397b585b25ad7a96827fb3340cecfcd453181d5e497948b6b1cc6ca8a93088e3d6b7e6
z7944ca0e91d0ec1a0b554791d6ac7e2abbcc8977c22d55b663b2a8e2b7a45e11b0d35fdd64266e
z89358099fb01d10993738ed8d5e05052a0133a000995a7408f1bfa4ed7bc6487c9a613a4653b2b
z5d19934dea4d59cc479cce5654fd2e0d8da60fb51d220d4a6d10e6d7b6e79ae78808ef346634a8
zb77eae4af210c16e74e6300771328f067c6ce80dcd1fb320ee73c8d010d7dbfc36dcca83b5c814
z32091038ff84d92b67f7a4ecb4ed2ae2383c3d592ddbd9a6c99a5a15b26812b3699ed6dc661ff8
zebdb09f7971a130bf39cbfa3cd7da689c0e8045549461c5aa843b4545a079852da09a75b5e043d
z96a1ea53a0457ae640ac7ffe7478c01b21fa9dba00f171cf79f77a397447e9a70931b52d68ba50
z2acd26e32e1ec17628e0ca916a85fd80195aaa460aba8a61d295c16852b064feaca0d83f94be5f
zabbfad1e97c0bb7ae91dd3c682c4d433d757454382674c19a3a02dc325c2706c5c90c4d7557184
z27e7a9773beb6f96a7f6c5f985d734d630fbaed12920526f8543e87a27b908b37a32e70c5cce42
za5a31fe4ccd2a17f7da9fcd49a14d0b3dc371b1a96c030d7acb9e283a2f1f50df178c61bb48f0a
zb1088154d7450dc88a594ca2a73262f65207a1a5c50e91bee0d443a267c406ac1affd0c9b302b5
z04fb9166b30ffa6a0535f0dd95d21c82a04d9adf165767476174ad3dfd5c202b59e3cb0922d004
z5b0a19b2f637f48729d457aa7f648ba36c76978db5b35749785783d00e692c3a8fb7fdcc3b888b
z82cb83d53c62eb20006b02fafbec5efac49d22df47de9cfe89cb05606d65bbb9053d045fadb871
zdfbee9f9b97ec1f3a55556ce0ca0c5b574d9d00562b8f0ef1aa013ca2050b893038b8250458f76
z34fe3649223bf4a425bdd8311f0bc59a4bb90dcc3d4a2def59e3b8d0a4fae7fb0d055ba4326418
z6a3f9ef253cc45edcb0a9a0daea7209c6ee14f9a12f228d13b607c61019d55d75d3633d3744ed6
z8068df4cf7b35a87304c5ed30c969151ae3ce57942f1045c0209424ca6d2bb145e6f2a6a0bed63
zad294dfc55526ebd6e24371a5d94425cb0899f3b7d1fca0127607bf7b387b84edf494e3c7e6201
z526cff87216a6956792348e3c2b88dd826f37c608a1048a7b912ef8bee471e7959826e24f26b3d
z1d671958ee80e9df5d72f34bd30d410b4000037ea564a721db38fbe39017cb6cb80e4001301d0e
z0e8e5eb2149789d4494f84b379a68e8f81ce794066d7055abe3b06d836cfddbdda67ee8a691f6b
zebdd0230e48919aa9ada112c3a3a048252874ee511f805618ef0eef3d20102c933e0f68fe419ad
z15dab22d09fcd81f304be015ce6cd7ec963c056d4b6bb34de876bd0a48e73473bc7330c4b809ac
zae5502ef7d23c8ff4c60c9cfb069273ae1f0d8bddeb1e87112594bb299a148ac1e7e740f57093a
zd15c301f745ecd99fc1d749ffee2603bf778d7f00f10026c8bf89c31fa7be9cc29b5926b0cba8c
zc7656c1591b5a50a546e407e4d5f21fec439c81df9f5621a19499c2533ce40a1923340a59a69a2
zc63e7b8991e03765e01ea09037cb21c203fb0016e64f1dee9301bf33b4cce88aa1aabf89183157
z0d80b8bef0ba8d9113521e78d48510b4b1d9f7f9f19c82fdfe455e24594fe9c2d44d6d1b089eb8
z1c5ddd3ce39846d84ad817d4ad47446d6ee2a33c79f8ceae2a675580cbd307ab058789535b8ae5
zdf374b2bc61a7eff71303543e5f68e16d290e67ac0d2c67f5b808fcfeae3c95046e9fcb78856db
z42ac9be88f7a1fa3e546ce99b2d95791c38730873743f72e8ae954cab8b4c9f762dcbdaf7d7ae4
zdbc2827a0a0a470b46e4f2b63ab1d3418a17b43e0c82a2556c7e00eb195f1d4d449d8747f9942d
z42c55b8ed29b4b3251560509087fa2f24b6cc23313e59a8ed89ef2ca54071d81c0d8e22d03cf54
z2442793531a45a2a5a112eb98bc5d9a45faa06410c8abde0b45fcafa546c78d78d52ea07addce3
zf8dcd61c755ae3d3aeb4b3a1cb884c1a025d40e936bc14d8982e23f974363b1ddcb30919495e05
z6a994c423f89a30fb98cf223b0ab8c4e8b6ad8a224ca6e681fc374067bbf32daab497ca225bbaf
zf570d551ff3888fd0f7c48d9429a46d7934d588f7c915afca13621a2998e06d2913c5774ecbb04
z0bca8dd03b75db727312a8223a5e439b358196e162afb397990b4aff805f2a79b8452ef85f6c21
z36e5f234747c65d8b0d6dd3fb4e74dcbb5003518a226a6f757f0e6595fed83eeee9e95db9b2d48
zc5459bcf059683cc5833f2e1894f418761b197be5c61563d4f56bea74f0dc6552298832313eba4
z570b3ec2069df323386daa52d5c3ecb266669023ab3dc923e50bc00dd7c36011161046c78964be
ze31d0ac02d227dd14f5c041a4ed98f86319992c3537d2a5be36309af63ddc101163523544f3815
zc2240757913a6f66b4decc2e3bf452872cac2efd8276dd05b95e7e4847602419914894ef481bf8
zf6fd56002a2888b16d648c34497f67b2e745c9e78aae3dac648b8382f0e43256d983c14f5b0cbd
z08450a85cd966176b55bbc8b675e9abc4590a599208c1034e8e1041e7ec33a290d834c6be994fc
z8e4977b71f69f56875b5439a6e430cc8fab66ac03d93746863388684464289a4972c6de210f509
z1a8c3ca8a921d4348fd60090b2a855dec9ab38a9f5dd446bc6c3b4c7b42632eef6ff7672294f6b
zc6ec67fc223d9195936e8c425be60c186b8e0061a16fb99d01275873e448080d3ccc1bc609ccfe
z98577670526cc6933cd9a1ef88e23a24bde723422afbb796645eff5b5a2803f8423f23405b5bba
ze2df9c6b2e22731eb8dadce55cc970447a9dff6113712ffe5555d4b5e87b67929c9dd3333e2ac8
z3a2f9497cd2d0f5e258fb042af775060f5e5a992ad1161cf4b09527b6d3cfe80e243fbbf9c796b
z61c0f9a69eb4591566731a13fee28b9f59c66c341f06b7787afae54a787c0c803b1a9d29139bb6
z5403202016d4acab7424ed83a76660a9820d48dcaaeb0b8578367901f35ec400cafa2b4111e0a5
zb2244c177bed9c54ca7ada8afeea9b4f6dce1f817c88f3170846de3b22e4e76c7e18cc39fb02ca
z423f11d89afd2061ebba595e811ce7738597962b0ca45143131b8ee7e18295e47877260cf28356
z813e1424d0100a2f56910e32004ae1bec3f33f23ccd15ebfa78b226a87f2dc77434313f414ae65
z348588684a1f959e5d8df9c21a89fca389eb817727ca4536d3729ab07b59307473f187db9d8978
z839b6a9a7c2dbc4becfd6047fa4f0c4eb87d0c15a5b91db89980684e9e877eb0704eda7be51d30
z2a391b48eef6f573798e349ba11a2a4806ba0ec50e3e8a4ec5400d61e4ed695b0df90806f5490b
z943c7cfab04a5149b59c3042097df08ff050775f02507282cd784596e0458b5c7552abe1e29cb9
z8b83795809a9126117d635cd84e286adf78d008d1d1701d665db1867e4684d0ef9f1073c0a8035
z4de3bf481c15c6faec123e01f76d8dbd9874704f6c4890328aea0d925c389395db8640f10604c7
z3e52c7139ecba79df22c1a8384fad85e518c7afcf9104ad651506fe46b63fd2cb92387fb26dbe5
z9d3774277dc3d21939836f1cbd31d9c893f444ae3b1151b33db72e108cbb5b942745349fc31134
z4fbf63d2abca5205f8517db8286243ebbd593127c1ea2368c9ab83dd09f832af737de0cc8a77e1
zf0f971c7619b0ab6c6574697384ea87bd2cfa0155fcb7a711b28a1d7ba6aa52c9c40486a384257
z0263e3ff8ab9645fb22a1876629eb7b13dddf35b4ca29fe3398fabea719e5c6364f7e8bdb93bc1
zfcdfbf81ee57d5ebd58c32c6c7b3720e19516ad264e4acdf6e1593ca302a18ce3ffea36cb743b3
z4c6a3112cf4ea5611e5bb21d9b5a8e1c94863fb9a83a5bceca5f55de6ac9bfccb536d9bc342409
z3613cc8721422098dad31f5a0c95062a6e0d356a2a382b2329a618257f37c8f6ec3c1163d8c9eb
zd9bf8bd7ce4f1a2a192c73e9c4533d20ef4bbd5829dc9622a712ceb6e2c3a08f2646a3500499d6
z11b18fd5d67960cdc1e8452c6106556b5c77164bbd5d940297e9e2b1d612e6bf866f6eed9dcd35
z166757ce79bd0443c5e25a8eee6e88cbb56722fd13582db51803732f5f9aee2c6857e8c810c641
z51e94fc88e2714aafabc326e069fe25ea9d895010d1f4d0327969d6c04115f8c94b91b4401b7fb
za0fffab4503b63479329f43491502c6b6a26c1cb3beed9e3b771f7fe3bece3685dd462e1e1d6e5
z85c982cc6a647cccb7c78e81653aafc0be9637c74367f60f829bc0822788bc8655079a4221d163
z543c751214c6e509425ad58592be62af89aa33b24e7d98ae4d313d047be0ca199e8281cba56d75
zb7d7487ee1ef13bf4c6345f95870de7cf1f8e9b7f572e10e07fb61cd7ddde1f7b4f1990652563c
z8aabbbb83b98193b25d197d2105d46619534eb8db4e105e49e1c752833803163ad8052f41e2753
z7bf98af89dc0d3580a441aef499efe40301f39437659ca78bf1c03237f09029db2d5dd978a7b1e
zf5be74ce4e3e7c6d69f5aa42367cb2415e8cefc837372a513d018168fb4805f74fd1ee843443e6
z823a2d00f7fffab325fd1d620966ce8cd241780867711fdf7781e275ac6506e73065b86e40459b
zb66c74c03723547dc36c2c40df094b2ab2f030a8e5bc723ea5e5bb33e8039e993ba78de2946aa0
z6f6319905b48af5330b0937a9054aae72a18d211e550407b44353e4645cf4891bce3a599020df0
z1f75c74e2145049d148dbc5965a68e578f98523f1f0595a7e079963aa432ced71cc6f8f315cd7e
z149d120d76fac0479d6b66d6c974e99fc59660c51e4980e73a3b2447cfd58cddf58933f072ccb6
z56379f92212c10f38bc9bcb6cee8276ec0d4bc10dc19161b2e9ce3a887b259fe57f841dd08b1be
za42bfcad2b2893fc90d3644e6aa671a7d12222ac76eb09558d999288c3db270a7f8ffa7d3a5bb8
ze90b14094463973ce66f8036d3e0370d9449c895e91cd47d4ba264529b6d04a3567ae84dfae9ac
z733603a3e63baca862d9651e08711b9e4324ff5ec85a1b31e67a5ec0d60e320752683a34e97025
zb07e730d12f9f5044b00daf4a1d24c93c0fd1c949ef060dd0339b6f936bf2fbf09f2e6a5d7fd58
z54452f9597b046fcf688befdb3f3e3d2475a713d87df6a046b18023959ff9a0d05cd7f066224b4
z39233a114eb3596894b688c3827eba66a1174fda7dd5dd2de219517c90e77d660e88e691ff0c2f
zc5b4743a94430fbfb3baadbb24133716a2b097fb91439a9bb01e3edce21e194c3a4fb4de9ce5d3
z6f37f8c0bc275c5f9877e0ca7b62bff5c6c04788c433637259bc77d31d4ab2f3016175d9f9be9a
z4a32909bfd012db041ebb06a78e9c1815d0625e476945f5827a0fd990b94f36affbacec68e8af3
zf40109b05b4d71ec00c909959cf7e4def04e0f890273298246dd8491d00f92f2f54cb0d24e6133
z259abafc3371264cf06ba5e9cb83471988aa86630e518c86e1177924570b6aa9a45fa9291e816f
z78bc14b415d29757ee7dd6ea60dbe9e06847898467e1dc74e0a040bcd742bb9489e79f25ed06b1
zde0e2130223aba35f7f824949f1093cb066a57e021c4a7b552afb1c7c517f6bf75b93639b402c7
z9588b1816c547cd2be7b2efc79f46213348a3b42873b47ea20964ecc824ab1a9cb568533aa7aa1
z23df785181b95a0405b402328d534b337658fa215c036b70a2fcb4dc50a69f8f981eed0e56b4b6
z2da03c4c82e089f72382b78fd4e35483ae00ff285b2e1cfce2e5989d7fd405e43701fb1dd21af3
zc861ce7545f288d311e2d423172e552143bfd7c43679bdd65ac083c9310f2a49a066cf996c2dc7
zfb39a6be287c3f7c6b35b26eeb2feb6863e9d74fac8baf07b54183128fbf6481f48507a0bc804f
z6b84d2e2f04acec4ca1a5255cd99d4b340b7ef7eebe892583d70ebe4311e467eb3db46b65b8977
za28f58cc971e6a185cdb65bd68966c8aee5fdc2339c777ef73ee112ee9be2dde9af4ed3f634052
ze001b8364d9d6a92d99c041abb4277c080c97aea3f42bcb4f731e80454d322e09e4a0e2c54395a
z0e8ddf37cfe3f3efcfe9a213c92475f2d145e6a8b9b214aabcf489ef22d084f5d1d28ebdbe8261
z271dbc744ed36c43724da6b0bc993a7ce2d447a8c9f4e6d27812d7cd460ce9aa3a239ea3edc084
za64affd4ff404d4cd75010790fdd2e7f8678121d77820249663aefcaa79bb382eb016be1043416
ze4632973a315827fa678b47fc2c49524f9e69d03417e40f6358150086bbd568e836f50272f0dae
zb12997848ba34a5462aa192697d2e01112ffeecc9697f3b29e0ce3d2185f50189bb609e0345a88
z7839f6b4ce986f609c7c6349cb65a7d7cf2e4a3247ad933a1e3083f3791aeabc540acdaf1d921a
zcd57fd8c3f192092268e7afde6719fc23fb492a2e536b022d477552be067540feadaf5e749e36a
z265331b90e625828edc27151f7c5b785c5e239a24e6d783c86e92275b7b52c6b7dd370c8ecfd77
z0d46a9ecd0d5378977d32b7331cd138a4bb9a15cb43d555913835790bcdc1406ae077a80cc3d77
z609842d038d963cd03c993dab92319508ab6426b99261eef5784d63d3f4838d1aaf99f9fd63f9f
z04cce6cf9e3e205e4ce71773c4da123f2e712537ef26145f3ff79eb49890bb0dd005cffb46aae8
z69813ea6961b5926601b277bae9b43ee413ecf850501c49d3102dcd90b73d37dfaf0ee2363d357
z7d93af9973e9b8f8a07f8f4bb837ad4742ae5c4209ac068b3c96e91a0286af444e8572a516b0cb
ze2f6aeedd989022c31b4415f1a9fc77f869561d83499045ca44e0741ea245157d53a69ddc9d6a3
z8ca00c7ed711b767bd475f1d617ff303d3f90acb601344740d074e2f5281af39752cd45fa3fdd2
z6ad26b6c3c3c4be3d30024cd3a640b670720522fa8dd29c85bab9cd71dde3479858219cd782886
z1f18d252945bb834ee69ef09a5cef1ea530c82cdab0478109a64585805fa293fd718488c396521
z543be7c129d3c21abd2e8a1f0c49a968b9d1d5e9736c0ed4571ec55044d1c3bbb94199d89d6351
z2754fe94dc81bab7f2c34a4fb21e4d17f38acab4c9f75dcafb70040b1c68f2929b76907af53e01
zb83ecc3090f569fb510a39f89110d2559879b2b28f42d52f467646bfbfb5d62d2510912b846d48
z90358edeacbcb5d468f2f4b7798493097fe8c4d53c6f565bc19ee67ecb43d172b325a60ce52c47
z667aac24250d3fb67ca58203cba74c12c666686e459923b5c7e17c47a2d79d8494cacfa0e8fd2e
z0950d75dbcd57cc7d5493caa3bef41377c6a61441a280ef0170e940915ff733b09c773e3f02286
z24a2382fb19ab2ba9d0bc567a916064416518ee508c8f7d30e5ad05f31dc9f1234bd80aa3cd449
z85c2f8c5e2f3ff2ce6e3ebb676832d7fa6929ec70cde96acf67814d2db0adf7019263da7c4c57d
zedbef97894d6b2f3168be3f07ccab05f6679237969a70f1e904d7f0dcd25dce293e90d4227aa69
z7d4c10fa42fb32dcd5310d2f1d3a55d1a26828f7cf484586ebc56655475555e35854882d66df87
z1cfa60f6785072af4e11f7f2931ba4531ce7e657978c63a978bc966520ba940a591602b7832ccd
zad1f4f864e580e1076fc993be405054234530cf2dc3c0d0e1831e6619089db0d1a35471e7c7e61
z89e4318a06ebe48d920850794290311b81d943afc902a928793c96c856d978978ed8a7b5e7ebb7
zf741964a45cc5b00c0a4f765e3b261c30d8bcc124d878af6acc58df62a29c4feaa167b2f1b8b37
z4738419d4f574c7f09fa2c69566544a0bc0f7e10a9cbabd06e8d189a7086bfaf45b5e5fc2ed0fe
z7323495612f18dadd523a808bbed603e94a8a02b7c3c0c35d863cd3910401e5836658a16b5d606
z1573544cf9eea0d60a00fff2f8528743616a21cc47329dc3432c1ce16303892f532ee2e16694b9
z0232935c8216ba6f303cbdaeefc4125e36d0f9a456ee12a980820cafd610d81d81d225bf4d3d42
z711119d86dfa85e01a883969ec7568ff182969e9800ac83626957a2dadcaf6cee3a84616f75dd7
z068dd22a66c62022f49fe762c7279b4e6a9918c65d0af7ff3e1237f4d02bf05cda0c64ab40c371
zdc242b61790fa9cca35b02d9737e5986b8e7e218f0a59f79ddcbd3f3b733f0437a5d78e3a30fe0
z7c0623f42e3da2f76f9e3f6c5ecde2e3ddb43c99a9c54f1ac52fa67c7ebfdaacded4e623527c17
z7f598ca6727f836958143a7cbf9c87e621d70187aaf1d88b41210544d6106a32c394cbdcd18e93
z83fde7260637096a14dc23cbb460d21ea56d333b6b2fdf8b929c4dc736aab46b40d6bcb23bd7e6
zcb40aeabe2acb71167316bff774bfbef61b31f49e64a8767dad3bb9dab388171318f198a10a68c
z27eae7ead47fe747fb05a500fbc717a50c58c33f8d65814f6a725388b666bf6b10007b4f8853aa
z3780a04cc71cb6b054bc022d3404a88276f1ebbc50a8cfee3b053eb968644f2e51f6fe5330d2f7
za825bdb62c777cc03a3f424fa0d5b0f42143d0f1931cd90ab94bf707febbbdb2b95c48232ad6e4
z2cec076fc5134ec0ce04633bd435900cf27de39483a139fc11e015da32339999566b5121656068
z52d001ca5ad23a3a72ff5982d07c51d29898bf379b730a6cd277ee179ad76d7027e9f4b9c4d952
z58bcc8a4a002ad8b67f7ba7250446a4bb973af60f67bb2afad7cc0fd47e8ff784cbdd095c0ff93
zf8b7da36241ada318e61fa76e3f4fd365aa97c8baf731721f026fe2ef125aaa88e990d635f5e58
z1537ceb3d962a70ab8af6cfa5751fcb29566a15dfe5a1f2880041aba8e36ab187045683a594c7b
z2bf8bffc07f3fb5532a0d9ff1f457fbdc67b39cbbc1fa7ce6311c31f14a6d3df775ea97be6d429
zc21824f1c2c7066a56e3c3759a46763b422c2a56e09726ef8abdd0501f833adeaaefacfca9c25a
z621aee8e758a40b9019589c2d4fb9930dba3ca2890cdb7abc5753839c84e0a246ec51672e50899
z646ecb3a3a5608549cd059abbaa3d58c7c4af19e82e9d93beffe34f78d901bf036f38e182a784f
z1c4a1ed307e73dc9b10506f4c357b07b21836fa95daf87b51acf6196f4b5e3fbfa38344743e89a
zaf65822af20509d51aa0f41615f6d39209aa4c049faee29e720c00381476b82c7f847ef42a8cba
z9702458446f3478e35514ba6939c0945e43ede010ecf9885cba55a9abc7d9c880775968380b03c
zb26447320670b83c4ea62a10c6f2718324858a7ab8fd3060a6bad94cc753f93e6818cdf854845e
z5c174e592a27a0f855626aa945ea8226e0a5a6c9ccdeef6123425dc5767e595cd39b16fac5a529
z3c75a475e173b41ab8ea2381f56c755a9441b21e8e0da4f76b9c77ac0665f55b9f59b626bd623e
z62a6a277ffb8268887679b5dcafe626fd6434510773a674398197f1103ebc10f8eb65589c55c34
zb4ffd64ff81f1cfdbe1ad81c8b2dab181da0aed02dd456c6c796ca50e53653cc62a4811b928c07
z32cd4520a3a5a288f74f0a0065ef9f9a1532e5c1063380b03e35e22bcb06119da885c0682aeee8
zb78cdf51514ee31753ec8446d61f22e83270454da16b6b7f7cb9951f108ab84e1a930cd73f6d3a
zaf0a23605b7fa9d6e25f9b58118ce84117149edd9efbbea87f6189b004ef3166e55d6407d3e053
zc4babcf65d0265991ef69c2bfde2b5f7202f317bb70318b115d60166544d6934a55fd9914f3f59
z1a0d939a6337459d4c8827d83922dd442ecdfa0d5a2a8aa496e9982639d51e5e077de58f399ad9
z787fc6b456f6d3f43117ee4dc941c5343e9c79f29e4eb25a1a5aaa8645562f196da2cbf041811f
zf97a0264552481c710c119d0a40ae7a4bdc08d6829b84926b127ded467b540b56979705f0edbe2
z37123ef52c44428b4af55a02d2da8bd2a545b1721932ba0b6a13c244068644a78559fd5496aa16
zb43c89b765485fe5cf0acf67c37a71c6146e8d58822b2ab478db6f224e9c2a575fca230355223d
z2c6fbb362623d67677cb2791b5f8f56f0ce930f6f0e77084d3843a04dd4b542e0fe4214fbe0369
z10cd11d4cfc85879e2b9f344b3000ff377243751835e2dd0eff6b826c306fd820c98e65a6b8788
zef1169d53375cc574b8b65f52c5ad1a5b2024fff4352fdb2e14143f97906f32a1fe69e979a8071
z2ce09b6f6473d0692b56273d8ac7b39ade49cb8ea000324ad81d6bc83c3e71a77f598c72dd44a6
zca46ddcdf6965104364b5deda4771999d057670c6ead91530cc438b45959ef346ace4f9dc4c81a
ze36f15548c68f5501afb7c4e769ebc79c2ce06510a0d1b84c207202b11643c8bd1b5f459dffca7
zb7dde3cf136d52a72c514378ba25e2aa4cfa5e84accc8d7420cc4529a7c0b078b715c061d2861c
z610c9af48002f54e477f921c37157f3b851ab620bf2762699766bc09bf0e12f7a3bc15a31003c4
zea2ac5eafb278bc2d3878bda3723f3619cf0a5e96665665d36c6cdee8f9874cfd44f82ea9e77d8
z8b41e81b944fc9fba22e0eb94ea505b5aadbb85f3378c9d0d0201f74fa25d16369a765d79bbbe1
z79726ba4988027e250bc6a881fcf9589e809b1a22d5edddd9eb7728fd735783b405002abbf005e
zfb0490b41b7742475fcd7444f048b80a56f57ad1325fca081360b5af664f38deab2d80ef49ad36
z5ec5d73e8e1ddcd8c4b8350bdb159216d0282e381f5c6fc3401e1945d00bef0e6f1fe1dc0514d4
ze13aa47d69abe1ea979491902ff7650b15f33be34a10c72180956c33d43c10e1dfd19105e639ab
z0bea438aca6f8fa39947d8272067fa9ed1cfdddaeb28688090d85be64597547b25c751817bd874
zc9a62907d4023755ee01b3c11f01bec714addfaff56f9fe09c7ffc46ca8af5240dd546a42efe7e
z72164ec464165dc13ffc32c6b6868f30c86428ee875cb5ea5715398dcd8f83be2417f8d9eb3222
z30d08a8d09badddb163634e1e3adc31cf73dfd15cd0f20ffca4a5c01921e26137454d97c7823b4
z0cb25410790c5f9cf56cbc373a8e18c27366aee10288483b1aaa19920ceec6858b9cd8e0f7e7e5
z6f0d1e30e6bc15efa27d0c9f62fbf526f33895224e51b6d20ea57f94161dc143066cd371b65c18
zfc79fb686ea9f55e8a3733f583c83dcaf0cd24f051b87e08f2326b4f233e1cf66c8d8ae172c325
zedd6844ceec984eece42e5d3b11d664ededa9e6011676e0764540bbf818db0890460dd237c9a56
z54924aeedb6ce245603a716fb1d04cfe6627e2bd4c700dd46fc06ff478a2b03bb6b24a95e8758a
z97286862e4a061e90d46bca96dac31915bb5fd4f3bf10e46320fa4fd92cd558b2505af1c50ad77
z760fcfe4b8e59842a20b515891c10c10ebfa8ce6a618d83cdf5cb3bbc1f4bad99405fb5a161aab
z5dd209b2d47f487596e1e7abf73f93b02e1e3da189dec63168f3442684cda752962ec45ce25b5d
z5792e8f6f732637e579d73eda30d6c568e08cc93865b84d3ed9cc24385e966cec903dd67aaa7dd
z4a477dafc8cd2dde5911f27af89b80e25a2d6f565abd30ae934cdf3933e808b7d123c086e2749e
z579fe552ce0c43230906b7d4a3c34cfa8710a0ad208a9e94e06ae7be9883ff578306a45a8a6b24
z6198800d2f7790633bbb4f743bd7e5badc9c520a865bb2139aa172b772ac69610bfa10d27d45ef
z1244e5fe154178cc96ca19ff2f7d3760d776d9ee0b7fcfd4d9dd4df1a51d0cd67325750cca4654
zb90c56c55f44dda079e280b3bd525c95d2ce96a75071e7c03289626e24cd0f1dbdcb5605cc3cf3
z81fde03816a37dcef72111be0536e73c5cdb5ba47f9111c76bd3910925afea96d5261de7b3d746
z588204cd93fc3778fe1eb4092a2dd0cfaefe31459c0e193a1391efced72eb61ac515e3a9b9841c
zab2e47985d63063728f7b931e51618b0f2809f5f09dc5ab9f089f2f7cd42eb59bad119bc76f99c
z6caabfb5f124c68fe4f1841b4b09d9671cec4889327f9e484a327b7287b88b697b0015b8b41baa
z6e4f596d5d6009959d5551ed64c94c587abe794b4ec274376c1a153ca074476743916ea35507f9
z85c85a502e2ce0231a62fd9aafe5528724da14374800ee08824fb3fc645b0e660ec12c8484538e
ze2c17c90b8d223150afe58d2999d6409128db8dd317c05fc2f878130f1bcbd8682dc4ce021724a
z8b1b10b23a1885e5eb5ad541ed299ca707cfa6c4ceaa8848d49db248575f7252ad88ca10d05e57
z993801e551362421b6ad098e24644c5a0fc9dbcda773a74c889cfdd1148d4642efe6c1ecd954ba
z4012a90ee41300fcca368b62d7be2d1bc5d0c1b8c84e1557f88acb457fe951c10bd582250decd8
z81431d90affa3e7bc613e7582500bd20fcb94fcddd9a6172f2d77311beb4c23e706cc44d573016
zc3fd102400abae84fceeb86a75049ba2ae2ae8fcd3bf23e8515717f8f1616904631d24dd8ea2ed
z5c7f9c2e6f245a96a2a7a728776b46d4d597d3ce8ce4401bae90289a3b3eaeb1f741af610a24e0
z0291809aabb8fa655405ab7f3b190ac086cde73f1d9cb888969fa603e00f8b8492d00127945e75
zd2419b6dc713758847a3c9232da7acc4815162129555eca341f1d8cb097180aaad3e2395573714
z5beb6fa17565baaf54cf977eba465db6a0e35a0d06c4d1c1e866267c05ac6092fc323177ccfcf6
z6d1b5f76e0f8318fa586980e477ed5c05beb206a26e227365edc686a60bd0ffdfb3571e865f491
z91aa7c4aa9a48f98bd23ed21157b2b0eacca7c8c52c069d2d7581127605c40e71e269c424cd52f
z920f7c0b859e4881b55fc6a2b88c679da6c9cd6d5442e776b21eb5aa7fbe37e98237bfbbec7eb6
z5355b448513e23aeb362d6d1bb626cda15d29514292cb9efc5385e8f130f5bde8ce931655f0f7e
z204d77b7cf0dadb9cc5e1f354e95dd12a3ef437c4ea958b67ad2298f99ea314cb6a156b24350c0
z084b0c6ee0b8cfe0293f7b9ef9c3b0dffb6f79b69a9492820f95997d33d89ebfb11e35a941ae84
z5c2e00475ac57fdcad9478327b2da1ce0611b962f24f492454216040fc125e5e721c26c0bc5378
zcef16ed84c21e9cbc578bf180317e26256f35df1eac2442cb48bd847b03c7b1bc9c22c36762d19
z4b8010145ede45fd3359603ba6b4a38311e1966ce4354f82863c0c3eaad3a004f5343c69882d00
zac29a60a0b4f9a5d15c093afefffc8179bf490e30cd72603e09e55eed280cf240a324f3e2bb284
z3eba7de12a267bfd6879b1395602e8c802f9a56e9049930123fa83d96d3c2efdbfa693cf240208
z8f4a9bd1c6e17945b6ff231260895d5ced4a43223c9566b84e3295ab3bd3bbc31ae3a689df0f92
z1e3d5d3294064d35c065c106f06a70d64f6bf1b671341d50facd5d082d44c871b016a1b62fad35
zcc553ea1783bee2aa4546bd650e001b93b14bf70271b86c7bf1c9218f4137062ad49e0705a8e56
ze7f8cf8c5dbdfa2bebcbd0ad37159552c6f9a031567781e3d7a11458557759955530c5c718c8eb
z9b85e0876d3ae266bbafd1d097bd9547a06a1d7b40533064943576e97074e752cf7df657f2037a
ze3a352e4c27adab5aba0b9a82a30a9991b852aa11ddb32ffd8a577dfe3d5cc2e23247f606a7b62
z7f1709d5a8146f3cc9e427ff0b464df414a945e924d026689e4ce04793d7b12d977f6236d84a12
z55631b50d74144268fa1dac9a5bb52239ef4a05b8c64d864fca71eaaf06b70a7096ea80aac6e16
zfa424f2a6e1b7ba43bb92b33c957406de2838785cbfa66570d264d76aaa10790511b74e18b5652
zcfc9bdb9438f9f689fb3f58344cd6aa699a7287ed2fe52da64b4d3b31fe7bbb55bcebde806f2df
z8b8814ac5f96ab15214acafadb3d2349db5d937558c93d2ba27a454931a0fab2a29ebe0ba40180
z875f9993e12188ebf067b7d31c6cb8d9e2a5b86029f9594c03e8d60d7a3e71c489de9b0d3989a0
z7eae7c9480b5719c61cd15c21271829c74ed3ecdcb88b17923230d28c8957c7fb877d11d157e92
zc40a5c8a7b48c8e84728b6c24fd70965905ea4dac51f0a8eef1d7a46112872fdbe9773f5a9c05e
zaacb0f61a3a928aeb037b7f2258b3397ff53d88131ab6fa907abaff64485912ef6ac0cd678af74
z51a2ca6f8b8a1dcc30f15fbde53fcc1571e450b7e99a3c4e72c5d4fd32e1e68bda4c60b9406a66
zdd9a38133e2c7a80e8b766ad076b6d9c4dcfa825d4dd3b05d2331da44aad554afc67c231a9605a
z1e46df5047f3f6e911663bcc1ad1531cb92f05ae39af2ec0767e0f3611b4b2b3e8ded1839f19bc
zd82d21dd5bce484e6969787f07bcfb02f7bcaa83ab6cc57f372c34658cf96fa4eced83f8b22354
za3d6f5dedd7c5edd1dbf793a88f5bf532aad5f8f18b72c98f4370520a85883b301c1a7b23b899c
z782cc26e56c9facc20c0202ee62127d7411e88c2aca996351d1e23899679efa28729582a9bd638
zad2900d3ed550f9c47bcf172ae9e4dd7c6e10c4c0a7cec13431b3773bae03a7fd51c213d835bcf
zb7051cfcff99241cd2be943fd9b61ba18847dc0c0028715dfe465f26b6aea08f7ecf8b6c4e7ec3
z86f9299115f83ea680e105ecf327297cbcc199a50024f515197635b9ed836c6da933da404e58af
z78560fcc56152dbd2c68353817e9681fbcc8069526a5b0f261000e16cd1411d021e71e7eeb3e6e
z3b48adeeb7893feb84fd4dc2d612bcab4b8b92614a29d8dcb9f0f9dfe2b937e6db8d6511e708ec
zf6a12fce1775dd187b72190bf1a3c039aeb8c1acb4fe2e9dfa699170c973c8edc0b3212c1510a4
zf1497cf80062c04ba6c81e93a16b0a320ce5ca6d013f2a1c7f43d888a693877540ac6b977c5818
z680ab73739c96d009438210c661285c03c0f86b8f705ab75eb4c56cf1ecd06f266cdce3dd31666
zd280ca5a2e3f0707e6a1a645c96ccacc7bf05c04dbae99b4b333cc6471835e705a478ae68f6b30
zc85257c3e540669f1320e06e915628c7d2c3e43f85642f6f87f5422942a00ea7bdfb4331b8c669
z55794c578a3a564d09a1512c03f6fbbb6bf17d7ffb35f4100b1498f868404231d88f4615151059
z523603bb655ca4f48bf3cf468c5288e23c4e723c05e79cdb21c90b8e95eec495d68ae2a1e72d90
zaff109b3de440b6ca82bc53288ec2e6d76010d0b5b32f298cc06255e905dcc4226e7e75c26be02
z9c3d8ec3f503f21febd6fef6f12848fd465b77a1a6f1b25e732b2316b7629bb7fc13db2cee0f21
z83ef7f6c6bbfa43ac0d14cf6b65624bd77f7f492aecab87d4ed534d2324062449b74f2682b9b0e
zb8c41dc8b7bd1f4ae2ab22f3d156bf369a2fe2bf63b2201bce35b2229315a346f84eb7e99c159f
z2b143796fa576686c75b9b989010bd458abceef39cddafef6078f2182152f7fa859180dd2b0d28
z95a15262f23fee540e8de755eb6cf3382e40c5a654e8c3a839564b41a0ce41d95356303cca1366
zcd620ff27c806acdc556ce56346ef644f4efbec82ed66ac910b88c177adc1beaf5d6adab1b84e0
zd14d5bf010fe9a230b8e77f4e337025c0bf976122eeb730bb442e205ef2143b3c0d7a18ded8f2c
z3c059461a77219a27792808454a615c9da37338894b1227ce8fb3405b303786ed5d37b6ac453fa
z16f0ae6ef3ad7030f74ed10a7b749b69ac3d311d5adffe3a5e8ef6ca220e8779d72425c64fbdb7
zbc58a68aca11bc6ca1075493a4a2ae1321fd8d938ca5bb30bda806259699a167549a87a4810294
zc6b66d7b84c8f9788eb562dc57a33c9a3945ced443692cfa8e39bff29761f51ec7d53cd01369ee
zbfcf65ffbb1a09b1438541b4c2aedc5662814f880b971c9e92dacf5da8436b4fa3acfc76fc9685
za4ced6ec2aefbaa38b842e9b730de66f06c6a1acc54cb7fb39a6e218e2d22345d6870c85b5f0d6
z4cfef6240fbcfd30ae578fae0dc70b464ea4676987b0f86d6f42de6fbb81499b536d360cb45878
z4ab517ff53fe1a5c8c231d27b744a5e577c52e7d7b64c220c9c57ff7b0e3076c60a94430389f7f
zdbad1f19e18570ea0300001147b3dff11ed824c6a3bc739f1b3d6f284491c24c7398623e11c512
z3ea68e0009a7aef07154d1a131e839ac1368d045496871974b4a30e3742ca8cc51a0eb67022bc9
z22bab8907f41c20c37129a2094917e41309a2a1e13dacfc36c5197109ec4afc0ea69e5022f3db7
z9358ce67e2f998d5f6ef50a048ae8e705e38678aef85cf3104e50bb0f8ee01c4927d3ef78d4f5a
zeda7e9e4494f1dd66d3b4b2d9b8d53db27e4b3ecc001db4050b56520273fcce6dceeb6ce9f2955
za39cda46b1901f28857c1491640cfac7ed54e4f93d0bfb0e942810fd7e0cbfe89f89f57058719e
z540e3670a10006fb8bdad5c7e34d7493041f4e2df99671ca9447b70e91e13c81b7322e819dec28
z4224e85499099d8243bbca2ab634e2c3089e45b2d18a2131ef415dd1ebf61db2ee68e7aa6b0c43
z97148aca6e7260b6e43ef3e22d57d5ca7be047e8cd0c4bf1f598e6e02729ee4631d89cc9b6dd9a
z624244f763001a316fefa8d93e3ecb7a1e5c2f6cd65e875463328ab5d581010660e4293b94ecd6
zd43d4035e85fee1bdac30aa4d9b9566712b5cda307d2e20fbc0b5caafd3c31503f8c9f724d6911
zb655dad9f78d33138a72274a8484e01e22a0440f8defc4ab2ee9f1852bddefd4081220291071cf
zbb5000207b3c868711cb1a2fec3ce4bdce0a659af8c648b379e7ab60f62ad8687483c23e259071
z87ec1807c1e19d305186c1a5ed84f6c5bbfb484dd266aeb261f4301ef0f9536efa5d3e2aa9a8bc
zb4c0d1449a8106463b23627e5cb37807baf5f77e7edd6e5c03c3c35f47bc537f8742b30a231506
z6149f7a193b503886443e72074bc974d431752abafc54652682398be9e19688b8557d5c8ad6f24
z843c43b199cee78e786a5008b8a02f0d6597dc7bc06f5d51c18d04a3f70c007c81c7830b1b7ae6
z91016469ccdc35ac825b1db2b9aaf1108a953abe4666fa4c4fa7d3c6741a9d304b461e4b69ff55
z4e80446e65f3c0eeee044062ecd11fe7aec6157cadd8a6f9fc386c6422ba2d15eec8d011b9a1df
z2971172efd4db3f3b233447a829a6e8979f9a14d7ca3cc3b8209c6c15414fafd2bd33ff8c78055
z0e34bc62156494f6a9309e0d1f7b8b30aeaf4b734c0c03dd759aa733af76bc73a7744701961e96
z776ab4ce602b2e7a437e49c4fb84f30379aa67b705e037c38671c18f5c643c174389784ac12d2f
z9c86c3db17d5eab23ab2a349cee59833c50df9d3ad697f683d8e534a8daa22a1e5c9501f05840e
z5fc1536cecaf150250d434f8f97baf2d31bded59485823e1365b01b98beb68b0ccb49e73154382
z44b8c7614b8a8527d9d97517a6993373bd9005f6785e6c50ae8a4d5348ea9ca741107c1d626f77
z3fbcf5792b58cc60b62582d4c3edee89082ad22a29dfd0454372533d5e942f9f1f3558cb6b3fd3
zb32964274dd641716fc9082b666cef37f36e6fa58012f5661bf5d2f680e6950c0be34a20806093
z6f2f9c491a9b817fee297bcbfcab05e458904ea197611f9879d47deaa50cfba5519e1fbf8425e6
z6233ad174f337e5a85b90f9bad0cb231932a2baa69c73d41db7ef7ca8b1cb18635220765f5e775
z58bfd048eacfbc7b72c369529c33df29064466f3e13ca97f0a7d5686a4107a3d49fccd5a371037
z5072f9be05b5384f4f4c8e75a174c154d89508c43c91b0a6cb3df0a477305e4e95fd4c66f52a65
zdc449aa4c7e9194b357df0e591b0fc6f707b1072830bbffccc5d4c0f16929d7b4af827d02cccc4
z18ca559f2c7da5c6b2d537a5817ece28bd2f29f16dac41e80c2ee11f90f5d463eff22714a3bf65
z8c7c36927f0d6fef89079d8f1d254ff61e221f8752bc061178cbad2321984c0919b79ae1fc518f
z5597d1c25047c952eba6e071c093b0af94ed1cfd4f87ffe412b3a6b8eb044ce6992b3268a2d7ce
z780271f07bef0a491e32246355d83a178bc7c330afef20d4d349c310d860e86d6c5cf5d1ab43da
z3af7cf722802d17422721cbdc54bd3a4fdbd3feaa169e0bd8acd3bb95d5811a974b12d1292950a
zf6af530c27b29cd302d2788f6797199200672cb108443bec6d39b3f07d0243040b225155ee3084
z06037022aeeaebda66afc4fd713499b2b9c15875b7c9ef583e7fe6a31cd7340d0775675197e9f9
z58026ddb7febc0199e981bbdd7a9982bd5cfb4c6b83f79360667dc5461ea13a1a5aacbd3e7d223
z920fe594c1d5249d40043ea109fd3a4aa32b0e9212b63bec4e6841d7836e42cd9b666c11822e73
z1e081f7ce24c77cd10b4afa71448d99d7175df996d7fed9d8940f95af287a6cdfffda37ab47e0b
zba2c62463cad6ac279a67b305a7a1ddd4abdbca402b1545fe9bea29c85302a1c58f42595d0f05c
z7b6521f60ca3071df448fe98fcfa88d6e06a19b1a282e3d2a696df56511e529a71ea68b541eb11
za01ed320278c86362348d2ae0a6be4bdcc0ad6c6f16fba8003544ade0bc9581ae34c515810490d
z3c442d80a0edaefdc6ebc11ba68259490db54a80c2d20466da7be2829c28f7e3f64eb39cfa7445
z79248974de3ccd0fa73dbe5bc3abfdc56ffcc5a8f9e44b09e1bcf874c94c3f84c164fa6ccbaf45
zcf122230026c10a359786cb189bfb1e2b1563a45720114d2c1ade00968bb865a48cfb1cf4b0f25
z5638a671dd2d254ee9318f186e03fc788f0818f7d560a3954b404fc9f81fce846b77aeb08fa15a
ze747d4dcafba472584071fb6c3821cce3806cf8c57e8894766ca9fdc2c3b30776d731479e7267c
z94be26535568a1839e12431e299769333edac77cd02ca025addb6ec76f779c6c82a809d3655159
ze8fcd69393151284f0cc1f71f29ed302bd0f4eb8440da29836825b25541046042b1c06000f2791
zb3d22763883bfc33473d3cf6db7b36f356877e147137c6df41c847dba282bde11e276488017e49
z891c1535c8f805717f2c698c5a4f80c9e015b8cd0f62c126f132a9deb06a1eda644fe58cb24c11
zc7fbebfb57d9efe5beaeafe4801e04fda1911621819e59f271d6a5b12064dd724b2e03c584d76c
z2b9f5e289a832a88bb4e0025d7ca9c4801849c35862a76ef068038ae2d0070f97897b50cd04b5d
z764be96c0d6637526a459441780d7ca2672732c3b5a4885b52d01de0e62a5e2ff5cf58ebb45523
z08147d8247bbaf5bb557465b2f71f987989fe69c29a3cd95d17f13b2c46e24ff55d39a69aef177
zac81371b0b4cddf2d2001c49a2121f2941514efb1d5dd4fdaa3bc0a785c30965cb2936550c0bb6
zf059b7d7c198764836d9a09b0654264be33f3a75f1d160b859a703794b3248e4a86ea86a84e40b
z53eaa9b1b9e986001d01786ce50824ed430fd569f925b166d7352a5dbbbaf036c509af049d250b
z0c4222f74a583619e95923ceee2882087cef8d88b3a0c1cece9b9475dff7e92eefefc2b30c9138
zb129251c53f932c99ceae09aee276673447a2ba6047003595538afdba08d2fbb4935212ab577cb
z19946d736437046f97352dac2240a3b13c3a853745ff757d570aedf3b72bf63f7adccc4b290ad6
zd3a4c76cd2a704bf40a2a7a5991e971112c355462f51724381b6948cd21dcea355569dc7b5f981
z4703b18f5f63e3a86a0cec64cc9cc1cffee7f9e3c1ad757e50ea3b07a980f1d6698e117946a115
zacbc652925520cb7c32946df86d16b9c826c21a6539c7f4799b9859e57422bb3880f87f8c4383e
z4f6f896edd5cc0bf6f1ca6439c9bd433da29f721d75bf8ed4da0506249bb8ecdd6b263abb4bcdf
z01d9ef6f723e6bfe23a209d849028a86380e8504819213a6b3080bed74cb403f23bcb5abe91d95
z55549f2ffed4e4c40e87fd91740d470cd3a440270ae2f15cb45cffb4b1ddd89aed055fde94e4fc
zd4e5742091902504f2862548b49e0666d6e9014b90d228b3c01304c890cf58083a8848522f71af
z42bfccb718cef7f908dd8fb427dd4e90ed5339313d466b88ed4e130a8f7554477d81464c1da6d9
z3fb7742c465e46b29365038123592e510841b76e17c85b874497ec3a7496c10a52237aa9761732
z4765bb575f3a23f757bb131f89d745286f1192fe88211895610a40067dbd7fe74af85409f94c49
z2f1646b8ff8cab2b7bd0bf86c2e462219e83299d04bf331183383b5f0243512f8d420e02746903
z1a02dd773bd1a956f6575b929d94be7d190efff0c58129c1b79049920ee10882f1745624c00066
zfa56b9ca9e766364626abd13c191f0796f79ab7176dd3d648b3488a12ac360a988c5d95106a0fa
zc050d6fd95d6e4cb32a0e166109c335869d983df9ee2ef537a3612fe45b8d05497aaebcade8db5
ze010c6b96033634110bf626c88037683b933f6228cedc428bd06eaedfc96ac4ed13e70a692eb69
z13bec136315f4e17951b5f6d9219ae4c19c9c77813240287d4177f9a0d5f18d1169cf054a9cc0f
z5381412418bf969ba431b1562c600c10de96f30f296caa31e93eb6e97b2b292ac53cbbe16b440f
z28049909804f38496d90d07a7a5b095ba59982a33e4296e02c4dea5717c9adc83a7e58e3e81367
zac8dd6e112484fb52e12b8f1775ea694d32ef2604f0766a4b548ad48ed3ff64e7b78b36a6dec0f
z17b1b7f44652c7f102c0d532064bbe96ac944b94a59842dfb26879d7abaf3b4aaaa0214eddc767
z75b1a1e7f52c148432389e32bbe40c0ae0f54ee0b559963828f07805cea1cd7b0a86a91904cd5d
z92b92cfe761f6cfcbe0e2d2292fb4ac6b87f39f768906116dc9466319d8c39a6e7a4736241c88e
z24026576856f6ed1b3764c9a0b9c396986c4b01f31c0e82042c30dbb484b32413e8be3c910b954
z1eb9de16816edece2d54870a3a6b16e089f202a8ad55e2de0e636e5fcac5189e5b5c74c0d14488
z566fc8bafc6dcc47eee1a95bf8e18db86b0fe1368401df4bddf3b5fd1b7709e0373ec5e5e86c35
z1b8c51546145c81c2bb9c3135d83339a39a558f74e351f2b08eed678ea4b9948bf87bc41956ce5
zc6c1fd34d91583160e670154aae37429cef765eaac713744e45ccda931134c9c927b3f3c2edaf9
z57503f41781885e0dba467ee80fb6d4e4d3b208eb446fd5ef9594e403c8f225b08f92ce455d1b6
z663a45a39a2ddd435d4a213e2b5773cc0e5af68aa50ae42e09cb1532856d805922eafe6813eab6
z01b5f571175e9ead45cf8dbd1865d404adad183cd26494b8d85a08edc1c533ea3185e59b81a36d
z695fa9549db07ea66ded9a9f7e13c05d2cdca48380a89f62a6eeee666d2e4f294d7c27c443c4f8
z00d9302805ac4b10a56bf01175a14c0ba153c7ed983c812b683547ab681d1284be2c1687b0d3ee
z090dbeff4d3b627cb549f799c322955d6f49a70f802c415c4667684ab5187428a1119ff00c2b43
zb987c530972d045bc944ee6e0fbe4402c99e6121b280fab9c22e3ddf14284f5f40c390e8bed4be
z1242cd52c38e2df480647da1685a37eb0d02bf26144e85b8872db91cc9ee0ef21b67d850b27d53
z79dd63fcbdb93c6a150df225a367ab9cb3456bd7ecdad911efba2532b8a63309ce3a13dca8204d
zb30fff8ab6f96b91489d9dd4c09f2daa9252b0e826bc5e7e21fd27c64167d1c612d26652c6072a
z75539031a30caf09aa43d422c764cddeebdde63c1d9493b4a32473cd682d729dd346858bc213fd
z920af945b9b137b0c48ee66fe61e12783d31a58a4fdeaf4dd6e5e29ec0c7374b607aa177864925
zb7fb16c4ff91af9c0a1463c010f74652797fcf0edfe77da556903fe17ab1001d510fa8202d86ed
z1c74bb472dea3bb5111d62fc2aadf7cfdef3da016a7c798728bf8a95b6f614791b9dda218bf8cc
z91c22208130bbd499c70c81efeab6357b9239f1b0b4bc60ce41efd2c32a1027f5a3a787a8a27bb
zbb89e4c3dfbe8a71bf6624b3702b4e01b94f6d4deffd6a7dc9a862d827c9a4703711fcf95cd0cb
z4f52ed020d68b65f4c43eef840976d0adc8b37b120b4a157554c20bba152ad9573890aedc38d54
z991972282ed542793829d418dde7a8347b9d8c71a99b8bddebef0a55934ec173d23874b3e48705
z50db541f6380931a5640e33013fc3c5c65be0bb527b470c3f420c804a1aea0cc211c5f9020fe4e
z9c299e3ef9924ec119503d64446195c63947eab3cf1f08e284dcd6e2d92c1a4b8035032b9f2581
z1a5ec5584d1d75970235933ccd95daeb44effeb470f216111e93b263dae9c8d76d1a20fcfb9d73
zd81576bce841fa0c675a7a30c6af98d77cc526212adfbb390a8529a997640c1b559a2ceaf8585c
z7623da54c76ea1029b73457c3956d971bd9975003290ccf2679ef769d64155ae07aec61935fbe5
z73c82e37a946fa4ce4b4a289f1f3f41b2ab0c60ed34c2f360b181001ea97ad760beeed81f580c0
z9d4ff4a9584f86df6369cbd9c15d570961d4d3559695943ef452ff2c08171abce5787c8e68f83a
z6a132c17e375ed3b9182cefbbc38a5d3bbc9be844e5c6079c29e5f70de58c91b749ae92bcc519e
z42cdcab19ad6c229e53eae9a2232ed0436a8198052df10a2f8b5f77ddf6391c585af5a72b7e92c
zb4b5ba954823086575d20a435e7e764751c5fdd1d8286080742e578802a53936de696fcb31e689
zf3aafb57ccce0ec687979cd6d93b3ffa9927f85d564f683343f1aa022830bc2a8b92a1fcbfd24c
z496a64bb2171a02c3d0b8b9506b269955cb341df37f13ee7eb833073f350f9e9b809e508bfa037
z6f9b4ea77ccdf77c126abcb45dd92f5da348253b934d0d0a755031ab853544a86697121939dbff
zc3ccb3bf0d0e545e31f16d72a5e379b93dab01714209227d5ab4febdcc9b7adf54b6d42a7b4dbc
z2799770439e42adf695f107a8444821d258c27830bd3d35b6775278219690b6852366bddae313b
z2be904997065b9420298130da3888cb76f1dec8b02de54bf5e7747a6dc39851db7f312dfad63ed
z3fa4addf6988cdd6cef56c2628e5c008f47488549058b84ee0476a0676a13fe7016111392ce185
za16355ab23efb661ee042632123600718e5e850fdf2ac336d5fcd6571c8256990695b14535e025
z3a753f2a3cfaf036fa3d5add95e38781a46bb1243e755710b06dae63569d8ad09ffa569f3a4e99
zdecdac53122266181d42e75705630bb95b994ad7e60a7c14f161f35efd40d8d1e9c71eb29c1a8a
z137a703151bdcb9962f8aa549d9bb5812d5738d47ab716c977d0cf7aac54b5cadbc8c934072a5a
zaefa367e0b28442b9b7954a132f83a0d7ec0291a968a003aba786e9dcb2c8f75d453daa5d9239b
z0d4a4fa2f6fea43b51f6e8f2759347653aafc9dee447a0b3a62384d099f343bb8dcbf3be6337aa
z3c41ff318b7e85939f4b681bc6b845a5ba7eaeb6effbdd57813dec3a090988c14ac07d75e5bb36
zde64b1b15be1f5f7bc4eccd86e43f67444251ecd9e82509e1421e22657195424a2fa94618c30ac
z74fff52c813533e6718794f3b62a083b50eab5b1ecd5862523c3717c8220db33e28756cfc8bf97
z37b653846805f02c75ce853afe685ca0905188d2758274fdd167978bfe24c9f9900d2d55ed69c7
zd2f7a5ba8d6aae4a40f1521fb6b44f0088c1226da4463e2b37ffa1d41ce74cba7f0730be00fc88
zb6014e5a0dc59d72bdef647171d7cc1df197031e166f89e1c07bb6bb3717b15eef520a53d4e847
ze403894bc5dbc79b491550653004c622ac2dd14e34f739e78b62fde2a60bed65a3ba745708d0f4
z3f9e71f36988baba9e519e754c7cadce0683792421cfa3ddfeff38d7c86dc35978a1ad78702ce5
zbc81015b3cefcf22cec1638d7df63b7f84339f9e6c3f5908910b164905c5cf55f92efdb9c90c8e
za5aec69ddce5656ee837917e860a047f13a17207c87479e564729cf8ccecbcffee4e7abef6ae08
z2c386f880e22b2ea95ec132ca603e43cf714566922d87ea61dad155ad8e6d38d12376a8220f4c1
ze83ba5e5aae185db4954ff40459861a2936fc7069f1eafa9c6f54a60aa471d231f6de4ceb1a0ed
z4b13f46185e069b82ea9a41b5854e876b03e9508fe36f87d2f18cad49efca82e8eb29e86c9ac63
ze9d749c36748cc22f10b71d88c63a7903b5fb9495d865d65cb2fe4e9d49ac872363c9a92211650
z65eebce1b2ebe7d74e0c1088bca13b3a06eb9c51eb60ff2be2ec04c36c568a5865c49f6bcc196e
z1997ca9cd5629be20aaa71fdd00519e92e98dc3699c72f40385db786e1eb1bee2a00398ff15f39
zb0d5be5326c7093b0483c45f243524b07a536583e850420b9daaaa4d253614d9aa5534d0a62900
z1307ad8c1ea35cf34707e2098e6c10169d370a04f65abacf4cfe5cd8576de22359e29d5fc0ade6
ze3b826deb55fccaab2ec92c7280b04b840527bdfb4a712518a53b30a6a6498365bd9f008415cfa
z7a496fdd2866cb2cb68172fd4ce49413f2f49d17eff6b7b8bdc8e883681d8ba1e16f324cfaeec9
zd5eebae6a08d9229bc15172e009caf6503a341095bb40cd9d205f678a4062bc5f64f56c61afa97
z468cf2944af960922dc38eaded1cf991d1fe6df7d298d5b804b88769682f5c85473606468c5f5a
z0e0d1597f40ae5a3203831e81973ae4ca7bdc8a4777ad1a2b8efafbddab5e5b7b6cb69f9ce2121
zabbd1c5ffeab8da012eea6eac9e2557d9e60a5cbf39db6c96df0d008503c18982430255de7a988
z4e6c8bb9194aa765f5576b05ef1c2a617549863821d2743268ef4ad4323fcc35fd31a7b7bbc6f9
z563080574d891a4c957a4e9e269f5dba87e88809ff9f455bbe3d9e9fa9a1813fe3b438a9f9a0ce
zd16459193845b79ccb7e75137ade17a082f90e238fad93b09aeffde01e42225fd5ad644d458fee
z0515f4bd4ae85d1957b60c5c7ebb226af2732eb830da5af4b0af02d590baf3f4133e76bcbcacec
z07c6996d15dbe82c4ed61a147a3ab151b45c30890c9d5efca6008bb8466417bea8f275dde8d184
ze344b403d5afe43f940aad66973486910eea465a60bcfe9b90275219e0d663ece514e09414a7be
z675efd3df1ad4116c9d6824933bfd3bc27dd75f42b15e5e1630baa37ac7184a8818a7589fa073e
z3bf829b7f8a093c5d64434c3917de079bb9f3f8b55501fad4e23e0f39ac4dbc373cf8b0f41727e
z9e457e900b01a4fd61b7078b54f3b9109cfb788abaa18222e608fa1d83ccf192cdad6bd312de58
zba552b9988e04663fa115d2acb5c4d3d595715b94ed3d64511cdc8bd422b3ace2700ba47d2634f
ze0ed6fe12e15482f35889735b7f932b41b8a3b1ced148d450024dfa24decd157bd9ac1f985bda6
z44b814074f8f410900eca13573e4fb3c5cadaa052939f1e7d49425fa380bba0b6b7ebd196f1a96
z285209de695e5f948cd83b99adf1a45c295f90d328fcd81943fcdb3ccc482a5e7e9bbc3fda61e0
zd2b54c4e6087564a49d7f9b55bd9861441ab0c8c37754434ab151abe61848c4115a0859c84cdd5
zd7d743343f63bea501f2544e5feb9e8700a657423b8ce50952bd4aaa1974488fb590c24f9bca20
zdbd48782e9bd211f5d04b2df4c7c17d2bdd43e163e8450b600262ca3370a80296a10830f46db23
z373e4e0894ff6f97eb47e78d0d9b73ea150103781fd0c966bbafb02a84b2196fcbab2b56f5d3ef
zfde153504664090fef93752c6f182925cac1c00036ac03d8c877e5986741f98ef4995ea6673741
z3773802efe91a3a766e75c2ad3f352e3755a2c48afde4b85e273bcdca6e526dd4e811e70c19080
z030d5e2d86f8bad9b2fc0f21b2764f59a9e613f04942f81eb8bd1d6d861fc23ef91cf153b987ec
z9dd707f186a5becb6737f99584e526877f7df740856b7a6fda4b26dfcf04b3d7ae389f0d1bce5b
zb6d65445ce4af34acda663eae1e4c0939970a7e20e37bde5462ac876e4b9b42edd1c10b58eef22
z653a5049c6bc4c850ca49bdb8de027d53db08ca043b57fb9f73ebc1807f15c055b884f65c9f92c
z73389931ecd0be01548a45dbd99ba417870a793e2c143215c2356459c7ed6cbb7e2b856b59ca35
zbfc4029834711a6e2a764636a5cedfa1670a27406cdd9d45e42819c31ee630a29689b369f674b1
z786bf77a9662d2350e9e640f09ba8bcc77361394d6c170e22ca73563eca3bdd875d76730368010
za106aedd8642c919edecbb35b8046f687c1ac524c618095535dff7788ce26ec7539284eef129cf
z67a277cfdbf78e37c07b5449f0366c292371617f6e671bd08694a16158db89bd19984f62799cb7
z49b03af990b87adf736385c169684a24a91e0500abfd1b577c2d4202579cc521b187a4c43863ec
z46d61fcb3e116a092d1d0122834dcd82ac9235c7dda84a3bf9419e790e83a582c2615e693ba05b
z6f1fbe9d6b5579cb53f5bf478f645132c6dbf9a80aeca350176b9b15e164d19437ca2a8ebc396e
z5e9703ce948d7b6e70fe48f9097e92ac7292ba17a23e4a518604a8c4bb122fb725e9d867d64be8
z577dcc1b356fb1e4c11ead00821360761fd189f5dd39b6bcbe5b32a9c6a836972e943f69efa05d
z5b7f1a1cf90e2b0cedab50d1f5af1e804bf741d834e58be2467595ac148be198454800f59eb1ea
zee6cc13223e23ff16a5b2335a6e992968a2e25f99213cbf4d367f4e83e8e468161c179a4c5f20a
z892230c1e80bf967482c8642eb8aba428da40dedb24a79b83e5d52d28774908f4fde4af8a7ec4a
z2832a7fe06b781beee1be3b0e0c7dc965268d95347f6a462bcd6758450cf0eb37cde8d5ebde59b
z2085b6308a582fccfaefb430c8cc88ca5e9b2efc0e6e542076770973d2cbe1f63f0fdb6b45ccce
zd8361efe97ad16c6de926079097c39152ad0ddcdfb781ceaa085d1d43f031337f8f90a79b472d2
za1e54dc29770995b9467176bc833993578d54d6f171d8727bdc084cfad07b75fcc3e3df8e456d6
z30ae53ef1623a6f9984a6941310cf5d9bc8595ca72d221339e5f8e51bdb1fe3c919b3325c1d714
z2eeb6c7272f02962613bfafe4f05823d0815f622ec75f0b72d5f6d05f3afc63504a98629ceaff2
z923576e2deb126b546583afbd29a00bc261e1c25a8a42ff60715c4c62e10ff724ee0727a39d41c
zf215ef49c2efe3865fe20e3e4b08412cd2795858cb0e5bc5fe0a8edbd704dfd7b3dd8d574a4e1f
z3ec655fb4fcd67b1c95558617433edc728d5642d9d002f94a2fe2a9cdb6d000d9aed077785e56b
za6cdc63844ae37fe30f054241bd0c08ee1ddfef60856834d4aefe3e708aacc85e8dc3fcce61885
z27f56e44b950ac1d103fde4ff6a32a7d473bbb46de314d89b64ef688d978398e15c9682c128fcc
zef5c303134b722e183e1dd6e0243b4bd01455f8842e5668ffbcc091c1d2b96d796258d071e23a3
z37e4f3b355ea793bf3741cc50706629138ab24b444684fefd6cdc197f125319d92ae9c01405f5b
z0240c314b23ad4b4eb056ee339fd773ceb19f98096fb5f365d73d680c9194602f9d6750ce1ee10
z0303d48b68ad9244cf1d5571d80dac4fa4a1689b35ec4b764fc17190fbebaa96596412b5ca1ae2
z6553ba6c23934d88331bf9c8766268eb5292cef3c20e2b1df302dbe778052037f0f99c48a076fd
z7d6f03ddd79ee54c8317a6c2d268d27d5ae32241f551937c8066b4c70e2773563dd8c0d9bdf889
z16d6f000a01c42e52f73e1e2640281ee2fb1772775083394c987b31caddadee77cc3e8c1a67c5c
zbc556904a5c0805795e5b0170c90b9247015c8a297867363e04cefd2fd918899d6573335bde536
zc582000f9e7a6fa5f065def5cf70d39762c8da2737a15b0e22a41320525a0df0929369f9c24413
z85d07fb4e09fda69e82fd6f8ec59fc3de1a6cf01d3251af101b2cc4e3f33a993b49b9aa0a86438
z8ca9acc9f37d768e69ca7d52fde9d84ff774bd14bcd257b7cca1a4609060fdeb3c9cc7af831570
zc551e2710cb6070e1773094a29c0cf838d7f10e57debe3dec612dd57cd17f1d1213e4e0c6376d1
z836c456d8bbf72dfd4e96e39d2c80117db38fa534fc2970db45db1412efb9d8b89b2aaaee85d43
zaa630c630d299f6e9e55ea3d8af3b0e2b90a7999af41e12d2594eaa79c0a357a9f5373e42cfafe
z4b47a2423c3a3c7c5bd5ca2e9ad4ee7873f48725fb6e93191b84bcd317494620d816bcec1e2eb1
z7a94a35b893fabc138ee767f6ad656696e0133fdb93e6e53df812502f2b7d0b8d4f69f0d24111f
ze264c9aadb0d6a9ff2da62d910a2ae582bfc94afb7dbac285bdb7ff3c4d4aa4c7ed5f2e4e7775e
z10aefe659223561928c872e702eb8109bf33611cc85d00966830fa28f936ed3e78ab2d2054d7ba
z092febf97ab12cfd6319b4137906264e4fe5498faf5ab6e21527c7745dce4457ea2e2f8676b1d2
z63e6cf3389c3449d3a41ddcd6ea081358ce9d444feedfa48e8972b8f93c21494d2e90c35c3f6ce
z26e927ad6284855bce9a8cde7880ea42ec3fbaa47a171d34356cb22204d96aec67a79a2b25e0cc
z3f2e160cb89878f8d79d97d717b81d2908f855ae82a055c334951d472fde64dc046ee7e8607a7b
zb845a821e85e76b26df7b1198482e0e85aedeb20d93fa1d9681e1ebc42f4b32887895a8851155d
z145cd0eb9ce8dbe17a2184e9ab246c5838d86c3a007d7c144cb3401281eb339007ce271623d357
za901ba24858ae88192d5bf99861af4e245cc212d745362fa65d4d8e5239f7822eadb97fcb6b169
z593e7bfa1da72df7b08082320eff96d3bd606d5a2c78ecaca783b587c4b88dbb9b424510945eee
z1e8ec0fe7835591af995d1dfe131135f4c536003433c56f2986fa8350522394943e6b334bf29f0
z191bc929576a8fa3485294df69b0e927bf518bac11d71ae77d807547cac4412c468b6f04a772be
z69d27e8dbceb38c234c0c9b1cecfe6932250b39ebd1a4346892a41c3f0ca1231c20bffc760b0f9
ze551694d2d40b0c25676494849245bf72a688aa65b69ea7cae334823cadc7db8f793a3b97af0f9
z73e537c06b531cbe060c9f1049232b52bbc49933704e518980f1be865cabe66333dec2f732cb62
z5b1135ef5a4895bde7f545f94d0f7ab3c758e8c70dfe49e0b92d49051ec34c4b8987d8ad2872f5
za2b83ea404d2c83def178817e6c27747dfb066b3f6c3d0bac12f194fa92c2cd2c32a1eb1702935
zfa52d7e5538b0ce7aff7e5cfcab617de277f7fb947b625b99095827206a1b7a71948b5d0295eb5
z8d53ba870d52510514d7cbb270448c480d701747216f03c0eb8e3bfd4c56c8a76cbcddd3fd5b8a
z96f4c5c5041495e36ba6769a75ac968b7caa0ac60f804bd97b5341fe902cfc9a53a238f26085d2
z55f7ae630e785e719796bd7fd56e082fe960b4e5ea811863e90cff116a6704cbf17d79b1f7b34e
ze3a631d3e56ffa0c7b91d2da9eb8bddcb12272d655423dfe3178233ec56cec45c5d85036ac727c
za9438ce15e4595461760e2a527c38d51a395e8b4651b3cb885669491c87337818df64eda23b12c
z9c05b9646704c9607a1587dfc0b598c20a8aebf2c7c7f1eb4c39ee634dc2585f311725fe8ddc4f
z1319fed1f5c852e23d6343e2ca86fbec6b89b2f2508a23873aeae52469c3d7684263e90981d139
zc422d8cd6cea5ad6d1c4ddec868f0d2935e27121333abd5fd41640bdf353dc2ba8fd477187d883
zac523ac4f6ff7f1dd0af976fddd3cbb1a0ac942cde9a467c089e9eb8b014beef83ade6095b47f7
z6287cd9a7d3fd952e32376147040b18823839c6cceed77e0e18c8664290d917f619d378258846f
z7a13cd33702ec55b4019324d45db95c56822c8fd30c64be9197c9ccb55675bddaf8d5f33f05fe9
z7bef72a7a238b3c5f96799d29556d057643d3c3ddb813ebb7dc1e38ca83a5600170dcf0d5cd991
z582438276b1068e7037b5286e838ee0f9eab44f6a1d14aed88f9d209139a3df5557cb33ed9ea24
za84d6e80729bc68fbf8d43933fc3836c61cb17ba870b41091c5f8e6f3ef86999cbe66ac86f2cb2
z67e1f23b1d3de71d8d37494ec59e793dc58039b91918a3f52c020d6f821caee2995a7212363fd9
zefaac5713568e4807dbc09dcf9eeba314519bebcc849414950d4810f5611e05f19bd5b7276511e
z9fb85f3774a8f257359cbbd1963ed46a3e46cffb8bf19dbf477fb6708d4113019f06a794d29705
zf685adfe08d87fdf686ffc626768e91a87cc0570ee48bb8e3963a0b73dbca7f93c49dd87cb75fe
z5be907fcdb652adbae516dc6604660afd967597c9ee532547d84856e13a41c3529f47a9977f63e
z64dd67275281107a9d1967351db13f8dcbaef843716bafe53fc92aeaa38bbce5a68ab8b79eb4d9
zff4449572db6a3bf90d17ed39287a0c68b56a664c0fd80378c9400e70298ec066e41da61654fc2
z13e6fb1b217dfd4af227fca418a622bae180ebf61abf41e6cb3142c48bcde334bc9eb9927cfad9
zcb25f129b6891efb7b47a42aae2a794f9825fd160016eb6198956ab02d74a389a06afec7d5f8ee
z29dae0fa4691d5e378bf43d013aa86d5300143b4b32714e56bfa6560204f9edcd059dc1d966183
z256f4383591c13e630718f6a3cd13d0172c7de1f5a16bc1ffd43799befa375e9717337755dcf62
zfbc0855c769a0c1ba0d2a2ae389562e3905e99ff4e1309ef0f10db98c62bc2251b1eb0d048334a
za70c889fc08a977b52d1e1dc2f9e1327dac61e846f71f67c6bf648159a675a9e0e4cc4ba946480
z8c8facf00c4f6128c253c23eec885375e5e9c42f59f439223fde9f45789db7f8379d2b4b052d41
z5459e44ffa5031cc94c80cf3b05f044964f9e3001e17d5eede29f3ef269977216d3a9473855193
zdd5a3696748326af20dbb9e979df2d85c43aaa55562ca3a7f03b50627a65b706451ee3ce6c1ff2
zedce37bca2c74a3e4ca5f4ba9fdd2cc1bad2cccc09eb9ac24317399f3a0f503232d6f5a55811c4
zcc6c1636b5aca7c97a98f3673bbc8516246b856a907d49b84afc60dac6e39b4632a0f0eea4e9d5
zc8b6148e2e555dcc9478b60869413a4a608c426827bef366f10dc7098df5873ca5f028d09abfa3
z8359503a1c95eef0d7fe000a5518c1198bf11739e6105cd18a063fab485f331eea2b49933f1abc
ze7a08cf79204597ef44a1c5b20cf9ab32d48989e097aefe7b531a8c2f1b73172a1b7fc74bff506
z18a907698ab32a301a414e78f2798c08b3927373e933be35dd59f603aa4f15311f495786003413
zfd020db47a94d4b912805de385c1be9cdfd1247f6106cb753097a6827fb481b81a9c24986a0282
z008105b8020f8c77cd4530d6e0c85c277967083d2c5d1375b9bbbe73ebe7e036e6c6f5cc713c54
z573c292c2ca1e90e6e91019cb0711fae02e9bc4d79ffd9a5e97fcc04b43381da332a4a3749bb35
z1ecb55800b73819dae3364b1b83f5115bd70c6d63b0ff114d0391690894e19d5a5550b92e6a2c4
z9825fe9a4334e84359cc2d86c366493740f3132a066409cdacedca325a421733ec1d3c0464708c
z8a373ac1e33548f0810c01241159b353acc0e0794fc9a7eac344f26f078c992b1f55dbc1c8a12a
z7107855c4b2a7726f18a84aa844e906f7e866fea70b55ebf51b4df86537a43285d030da6ee111f
z606bf6d151af56d938953ee5f74f753d2da48e218aec9418f5844b07987a514bb57ec6a153014f
z1bb366182d939835006533b2d9100653c2fbe51bfd572a050448857ad1c0fd7483e6dc54a5972d
za23642332e67f6d6683fc61829594e96e4c48dc82c03ff7b4dcd44c1f4112e3a2c5bbeab25ac38
za7735f06f46a8f1ac81fbc62efcc541e0eb926c52175a6ebc10e957749e798bd326b53451d1685
z5cb9ebd13fb27f8e17b410b457c7d8ae2c6d785c55779d176a7356d928e59fcd5e12afda63fa9a
z2041ada8b24aa65f312ae753e448ef3baefd855902bbb28d47f0e2e8e86d24aeb18b3b4c6205ad
za1717e82bcae2bcbfa5693589d4364f9954fccfbb46547862d9ccf04aa06a465153e7f09154066
z81f61ecb8ad94ad182b956e8bc57127a09dfa3b65bfaa906bef84b35944ea45684bcc44ebe679f
z13e7039b7593129144d067a0744afe0394d0a35f163ac3e17ec11423cb985dcd76ac209b33dc15
zcd7471e249442be7ee776d47b4e17df9db6bfffc2b2ad1756eadeb6b4266694077f02b399f4ed4
z6dbcc27d8725866daea928fe336f3b131e9055652b2cb5fd2cb7e9d2430b57474dd439b51c9965
z0cb73aab2e318d3318466410abaae0eb498f8e7819cd962300333d382328878977da18cb718112
zf548a6991e9751a66fc736e43eec641eef0862822e52b7828149f1261645f368c8490d9efc66f7
z09dbc1a376fc89e71bb0e70d791d088a628e5dc8198417bea77cf0d872d8f16ffd3554e3b53c26
zf67782938414c0326d9012ee27ab973ecbb9c55605da8e32799841647f59f315a04054458a09c2
zfe68471eb0b7346c41b1dde9fb47db4c222d5c290fd43dfb38ced83e25810c16966d91af81239d
zfb2c18caa5cea29cfc6776d47be53a11a5ec9b12db03688df22f25de28068edbcb506527be62d4
z64d5ab5a7cc8092a2a94067379a9fbee647fc67c68a04c33f8b5fafddde768fa6b947630246c9e
z62b95ac30b38780cd68707862795f039fed5f2408696900de7dbdb23207bcc8bac5b79309b293f
z1a3e87b487c68d3de29a8cb982ef94678b5af5b6d8fdc069283bebc29edd04ab67a8bfb774a5a9
ze1e5e22d14f78de77460b9da0d7879776040f3008db8600efe1820c86dd6fa4beee9402cf59015
z78f04ae166eb2594e0c4118fa5fabf6ca15681b498085a0f03f92e8bb79522d8d3c3051e55132b
z87a7158588cc45cd702a2955df811d9eb84464ac8a6651910e0efe256e54e3122667a584487695
zf3ea9a8c7e7108eb47b06186ef4d64f30fa32f5928d93f712ad15525c85f622e271d4b147d7f1b
zd77a0f22b944bc61222ca281a4f2aaa4c27e6de8175a344ae0b7fd478cf7b419a17a160d2156e8
z85628659a3c95d4fbbde0d6e84fb77d2eda28d254f2710b83d19a9c7260de38ac242ae729cc929
z82195c1025a39af2a2807da82bb8c90c1f37eae6a948819ae8673cb8fcdb48eb22faacd1b81eab
z5553ad286b65859d6896abfc883261d915954b00eb3d32a92b77d6c7255a168da00129363da8a9
zd837ae4dcf741c895a648b3c78cae8997af80f15e839e786b57e3985b3b5b4c2d7f029a844dc5e
zdceb1be6b6a52fc2ceff52863af1228873ddde7792f0f5fdcf1a30e9ae4ffb6040568fd8cf4c1a
z138ac4335b168dec7e27f558c52a6d231c71f8e8b52e18844533bc14dbc6dd42cb4902a3e7e5b1
zc0179d39a233dc8faff87908beef17d1960b2cd54a4090ae177420535bdde8676ca6e46b97bf1e
z1dac7119230264f4f3fc0e1617e9f5ec7c3d8b3e36752b3bf9132c684a8d06da5c5e3baeaedbb8
z5c645d8a86d1cb9c99f2df956030b7354a31d4878826e03a18649f18772a46280c67c86df26be8
zd6324ba5e0891085b408970d27340f4263171d7741b323e1d301fc50339c520aa0fffdc0fad6ef
zdb3327d078d889909334616c11f3b184758f2d22974f5b0ef1f597940a573a726b0f9145c80a9f
z7f31c12cb2422dcb7fc7f9b35f5a007b852a977a04e03029cf6dfb70be44ebe4a051b72935436e
ze3dc43061f3530139047e134b96dfcb00d43f5986ba329332e333324e1cc1d60291dcae8cd9a19
zb7a35f7a1c3d44b36729e86aa0ff23f11872fcdae8c77c94cbc54cfd9acda459d6223a50516fe5
z072f880eb98540d61084786657e700cf01adf16d9e032aa0184e64b2f9d6168739e9f79c0e91a1
z63e6896d723001791c78f89c17bd67c2bb6d8fd07efb909370c2bffb91bc09a02313ccdf49c85d
zba09d399940ccf6ec59e549212b2cbd0f5c0acf95b3662f4df2733eeb24448ef52b984d937226d
ze181ac5bc7f2749c47b1d0909deffd907d10e4c504e062a907d74ff1546f952f3c1c0f3c2d6525
z95c4c80a971c6d7403403977bd2e99241c6b330eb0887fcfafc739bec8443243133e988343c59e
zd761acc43c2d69ca1286d32f2ec87989bf7fb2cd22e524dac0a4bc0a025e34ba579b3c9881a404
z5103460c9f296ad79ab5e5a3068f3e42fc0302cd5e064d78bc8c3de8ae309fa12fc28409d0e7a2
zed1ee5439104137b2e39994302600832145b83d5727951fc34e6acb353bda160877a258d6b67fc
z8f805364436171978e91c0fbd1c525640d2cbbfe1a370397916e5f71d691a48e27c16daef9469f
z46d35489d2bb0abafecc61128b219b7933afb08037dd17969edd63a00e15d44de9b1253552603e
z7fc35c8c4f7a35b3fa42ec49a4f8514810383b702299bb46f70510e48be712109ffe13aca65343
z92674f07c1e539b868d1085bccd90d251bba1bb523e0691dca00833f6e8a4c5420b57f47bf84d9
z18e7dd562d592028d7834bf88aa72ac318b09381aa004cba47cb5daf76ac0438b1e8e58e3a5353
zcb4350cf386f4fe57dee1a04f60a56916bd842583e853cd9af6650805b855be27ca1191096da64
zc5df8fb753e0859db8f4f8dee4879b029a30e025f74682c64d25c8b7ff472c0bcfce82ad56114b
zf7a3f5f5a894949f31045084e1b2ccd439c443e2a8f54da4f50ccf91033a2c12f8f7f89280a0ee
zbea069b76cbbf49c1be8c86dcc25ae8e7138bb6375a4d2995e57c87ee722b6b2e8f1b2090f637b
ze77e272114758c90bf01c916fdc83f777bd47cb0d38b5df6e27bec9917b9a47fdff42783a8f4d2
z4c80e7bce1cf2fe4b14cca45996fe78fb4ef90e73d268e480658f7110ec2c878167484811c29c0
z3010b06a5eeba5cffef7c034023298cc7cda5e2e042e2752bba7814aecbbcc6f74dd0de2838a4c
zb10138b80edeeb9a22606d3dce6cc8a95748c2396cc433ac4af6ba3155ee2377dacb00ba49541f
z6d79fb5116486de2eca8c7ab7c7ca9aae33dd4ecedeb948a7a7f4d17c8394efe2d8bb07fe51d1e
zc0ffeb18e7abc4e91d8f8813a4458495555dd7f928f7e50ecf91ef29a8c0bc17bb2ecd8ee1adea
z65f17ee78831ba72eedb1aefa27c50fd34b2783a65a42c6a8d9dc77cb35a5f05968f97c2535067
z955207d2cbef160fa52306a28dd6372aeb933fdfbb72ffc3a31313a146cbb9c1ff470b7f3140e1
z6df51d135f5538c255f12e09f3ce9d6b0f399c46ad3c5f693e7ed346c0c2cd3718e0b0c8ab9981
z3542c19c7bb2b26c16bdbe994b7d46c931505eabdf9059778e1dae00a6ba4b4b563f0d7611664d
zd7c6ceff976aecfcc277084d9deabebde4a829aa8da4d4181c02d64159a619db929f259d322a35
zf4e3a6e6860aad7004021f57b742fd48c349897751934a10f38ac9aed6621a77440307f47ac410
z428bab036da952da5af21644465b843cc5b163c130864cf79de994d0a301b34f97005f3c253a22
z5c600a745de976ff8ef6c65428eee47352f9df2921b260836e59a031c003ed773d4559db0c4742
z11ff15f6d634f946dd6c13deaf5f385817dc84545ce2bbdee1319c260d7228bb3d1874f443ec3c
z1a6cb8fe85134d41f0fe83b9335fcec78b005864f2357df33a8803181f52b4c827857bcaf63e6d
z1609f1a6b2e6eb7d9bacd386a4d0062cd02ed2e3067e9d8f4942a24d33897305b0dcfc0a4a5c3f
z6e838b7a8de0afadf2905bed191cd299510f5915c124e2b76e90ce2dd219f31ce7fcb26b2ff0da
zf110400a3a132cfe0e5c7bf90317a4e89c4c00edd9c853c913c81a9bf2233a7fca180665674b50
z75fce8b45ab85b53576c67c41834e66e835194638f9d1d529bb51592a9efdb6717485c61a751fa
z541dd86792de1ffd15762a097e7b9c6ab745e4d566ab77082cb8c841c9c40bf40f186362fe841d
z152c8433cc83fc0487573a2798373f897f7ae543c9ca178c0628a2c1923a1c7193a4732bacbf77
zeeee3ef944d3694ff3df75d5d6aa6eeaf333bd59ac99912f48e1b6faa6c698296b8331870b1ef2
z7424cb2449396b7ff2e5394e08ac1641b115fd86859f8fb7b487a4ce8c9199aa8cbe0507e10bcb
z5cedc48e05375c03abb842f85310a6fa4cd34020d3d262a9b434beb8e9149981b9c0569a26074a
z739b4b3408529a52cc3430fcd33a0a0fb756f95c050dba7fffd0c9353d7aa81925d5b5234361f4
z7ff79eaf3145fd2c5dd58781b9e5b51a735b02b3ecc28f4ce3a241ac8c137f25f2ee135dc8894f
z68320d773715dde3c08765362bf5af3be74d32dd110a65e725f8409bcfbd09ad0ce98100078ffb
z4705327c436fa815e9392e83e3775923c3a5c34d9daac6008a737e046747614cf5a9d4db18e508
zcda69b8da4e988dd3a859a478b3c274e5c691b137f99cb125edbfef9f036e255ddf0492f4ca80e
zc4bc276f3764f6b88e27337339a3e3f185d42985087315824831f7fc3551dea10db499b4dd5b83
z10176fb21c1f16fb560494e5f0d7d0700646019a3972cfd6146c94a095e43d5a0affb469bd7355
z1c4f52887147fe2c7b917e9b80f624205af60181160a4d44407381c2ca077c7dd2d466495589e5
z49a1f6c91a216d17b5acddb7545c775d3c3ecc66257fcafef4a12862cd5604f5b8ad4bb45b32a8
z5c24bcf16082f3d7626bbc18edee474a60d8ef94b3817be7b5f448a103e28a65fb540d150d197d
ze3216380232505c78b1dc660e35a489ea238df3a839ff5ac2cbf16775803b8e359db34890900da
z7e41cd9b2bcad21de2ece7a27a655f1849beebaa1fb7532931b5716ec1d29d50e2339fc7ac1277
z9500f9d276888560f8fe7723a4b0c1a370b7360ceb275af3b5bbca9683b5ac26b539ebee19e68c
z6a8fdb39dca7d8d2175286153f9fcc57aa9e3bdc776f14cabe72d63ac008b1fc8bdb2769723cca
z1b84c5d7e2239cb4278c6ee2836aa7998022b91bef4c2f47a12a10bff54438561009f2855c9213
zc73c6be4b67a4f4d61907361afe5a8348c97f03bc72149be9f5acad45530868154e99738854329
z87ed0c6cf4ad8d5c06539c03017af3218cf0cb97be31135d77d8233d0d4176c499180eed43515e
z5e4ac50315c86d249ed39b2e3f1e9998724b235364d492867d096d04173a86f8434a565a125d83
ze73b932b9d836cfa991d6de9e5829ca64a3dff721c431bc6fa82820f4dd6c1ff098d9a189e1f8d
z23a42c22d78bd7eb543d74af7efbeebf56254f7f7e7fd27446e6e917355af53042a07522e5c871
z57868dffdb6bd8b94c03c3f0b533f0a9e34cd41c59347c6af6bd7952b3c2f9384d3711e395e93c
z65d2e105b61ea0845c5c5ca3636d771ceb2b66946ec1df8cb79e36979c65fe8df1a041157334a7
z2e522515c354df67e1628f81df1a5cb3bdbfdb657445e57bd38550bc568c55acfb6054271642ad
z025eac3ba05b22817ab7efcc2936f117979a6245f8a0228e3e72c2f3aac972c9dbf3a021320306
z0f457453591e6057ada1c8039405c66c84965ab9a3dc60c12f4bc6fae70a512e2baf5d4cd5d465
ze1f8debcaf6b922fbb78a0c71cb04a303b04fa38c67bc29cd648fe19e1098075ed7a9228b8207d
za6d4f2f6be8802d2135d1e59d6ad80b0ea2bd0afaba98c9f987097c29aa677f01ad5fecc60b5bb
z739dc77582720dc05f888b777f6e549876d468af526ae7cba27aae86b50b0bb9fa0407aea1b0c8
z3c1d3e5c1742c0b033b7b3158d9aa46bc0583bf137ea905a62282ca8a9d96108be64e7022e2cdf
zc3f55af373a3e0f28498f977ca43c647d1aa841337b430255f7808290c3d4644e65261c2da5215
z547863ab7cdf7f33e4f76f665f454ce895bc1f6d971eb9193bd4e51779435abae994a8e8d12d61
zb42ad22e4aa56d57a589c741b6e4c6ba4e1935b4bdeee9a2537510d1944f0f519c8a35b5ca21ee
z6fdfe3ad512f1921d9037e333ab60c4115bc3ff240d5e00723ab57aae35fd14afb3932e56c71a7
ze0156041b74014f60d33292db6cc6d3e6a644a8e3335b3a2b29f72567406e58d3a8af32edfc1ac
zfc5fab8ee45d6aa86bbb1fcd45b70d2b0a36348a04e7f98f18583820e930ec0813893ad4da741e
z1cbd8b12d33ea46c7226c7ed50828d2c9740bed9e8469ca9886a9ffa96c7cc4942b05a483e77bd
z9fe5cc6d4c3cdebb63d9639a33779cb9db3331fe306d583ec517d33e84fc010f80adba98e2d55f
z0609396dfdbeddb5ed3cb56fa2e971408afda01908e135b1b84719dc717a542670a72be643d2f1
z9bdc83816e4b9d01595d0d29ae60ce41c8fb95d69f724f2f1018dff8d93c797894556e3ab6a6ba
zbf9aa95476ed835dab2e7ad17d158c960fbe24b0ff806f7acbca16dfa8ff1dddb4805bbfe8e6fe
z6984e0cde2f510850a34117a1cb205f19d13365868ce1b768927f79388a47c43027b721ef78258
za49afbfef799a3bfed7627f1c7285f2ddd89b759ebab08672cb466e1664837ced13c7991e9f02d
z48f9abff7f8967b7e732d9d4be2af6336e0aa7bae1d4f689defded09c671fbd60f0e9af8462283
zad0dcf93564e39e3448cb48b4657548684dc081350abcf27d655b2bffafaa583b012ef0f795b2d
z370f7cc3224963c85bb000dc6201bd8045edcbf626dcf1dec9b88de0ef72f7085f9f2e1cc15ee2
z749e4828495bf7a857887655a87df31d941374e4f13d8b5af9628e12e62e1f76b666cca360a079
z6daa2425d9718d8dea96efc854f398b45065f7f0cfaa30f13c8e673cd59d93bf71b7ab0140a76a
z238d523d5495de37bf0c274bc776c22b5b9c72fabd5b62f4563fd69b46bd1b69eca84f97129f33
z2dda9cfd3efcc40106152e0bdeb8f235393879bc07f7ffd41db5d087588a31b5609a9d55660927
z896a8ce83041dd6be2fbec13df0e95738bd6db22d80c45a775974a8954b0c0bd19926168109867
zd50e3c95bbd7caae470866c5496a0d83db6d7f6c12b686190b4fe70e8f3d4207b0889ecea2877e
ze9ac5e8e3020f9feffba53e3cba5b0f7d2cb1636c2b56a50fbfbc85cfb70efc0acb343b3d71769
zd64188ff3c08661246fd4d8070667ece2e7cae093c2eb80c3397031a8866fa703877c21c2605fc
z8013df53f8a36839ab4c3813d5a09aaea0827e3fbe76bc8431b917775c8c8dc3036d3947c41ee8
z3d9a90efcfbb40733526ffd07cb99d008298f8380bb664478d735e5f11d3cb0ae72d7315395611
z12fba25015738e89f29f034bc30dfd957b20ed8133deeb806a17af3d8381862efe19586aec6206
z3497e79deab3f168bd82757b5e69591a50eabe4d74b7c1d64db850b0366830dc3d39d33ed96841
z5b5c458b5d2b767c51531aaa79247bd07502f62b46badf400312d6a79a220224573442230e72e8
z8a5fefbb57d2c0439f05b3268ec369a74b1b521a5d225f5ded8ce0026735d9ce3c9f62e3c94d19
z39fd814338adda5c86d2fc692c239a6c602ebc18e8917fc5c373f78cf069f954da96f4489eb42a
zc0843cdf4209e34bb2340c739e30124398ef6b7ecb0fe37df84d6768f50e21865e06bfd3dc56b5
z3865e63eea99be95b15586a76c8eb902a5fcf179d6ccf74ea8cf4955dc708209d0d6f44a9b5c4b
zaa50fd2f8ceb0aca3f1f96c043b23eab9dc3449357933525f7256ab26e4b73eebd3834114211c9
z627a6d0459745e78461a6b8c8aa3c37e99dacc79b7bbb704a6a2993c2029950a163081204cd2a6
ze0ca32a661b6cd1505f69e21ee62dcb9ce7d623f0761f3dcff881696a12a005ce5fb7587b7d120
z8a0541292c23969bfae564fef867cdb043cb0ca0fbf0519c57cd69ef6c3ded037628980d164794
z66613bfbb2bef4a6962cb760d1deeb82e0e1c95b08cdb9ead97c4e796de4931eef85b87262e8bd
z0f0fc6fe7526901ea9ec7fa22b0ec7bffb346cff441bcc418c31393814d070ed45ac609502d264
zfe4176803d5220c803705c1fffe96276b62ff749d4077c2a312ffaba0834e07064b498de1ffc73
zf44e68bc7bd363c236bbb790e41db91ed462f3fe23459329f70699f5a760fce1d3e683a9a24f3a
z018d308f67bf7fb3e2379a593f8b18e0e55193ea2f9c020e8c404779d6532f560369b79d4707d6
z2eeafea730306e8b4eb320081e34ab7d72bb440a4a2655eda9646d1f7b19c61f695d051ea8cc42
z6e51b47002041fdb92c7683541fe6389658bc51654aa43d5ae34c19f1ad7e32b2f3bbe6bc3a04f
z3e9f442168129c717b1a23c250cf233ca9e359079ddf8213e13b8df31f358d9ed42f9616cd9478
zf3999a45e0e8a1ce5232e4f0a0c059d2b141961db86e0ebcc7974dae520b17c391cc30c95db097
z1b0556037536ad0ef6c449f424e2ecd5029d1239829d232fb29f1f1b949c2b9630c198795b40e4
z3656a8b24bc64c5c8a14b6a7f8d7bae39d64632d3b576318051d3929bb95ac8f7620b4a6afeb97
zd6e6dc0069acb8bfeccd4fe3db599273cc2628f6fb0e5fc746f5949386bb61e1cb9dd95f5e481b
z6ee9b1f65c2e70efcab9c53df1327aca5caf849c2d9e325c83d0ca449bcdd8260ae10499a70767
ze6c36acd6d6036544d177d9bd55ba42f81e84a33ad9c93b852ae6d39fb94aacf5b88462e61520c
z7a8a878ae85d32bbad1835b168d63ada7f317cc3765717663423dbfa708ce35f0e6955fc4f64d7
z33c0e586890fee57b2a469e10feee24a97c69b7e5f5f12e71d7d29d16a7b5523287f64440d5a27
zc5c5fb4f0f82e7e9390480e2b93485ccfc734b2ac999e0076a80e0aaacecd22e90239ed86792d9
zaf9ae28a7d5fbe570f9939348eeec1e2c4f0fc617a8f1d9f9c23d4e74213d5a26aab0aa86ec6b8
zb1ba2b4e80acd78ccd1c22fdad2e19af56092ef46f8cf13ab6e598c66d35a291da1f6a3f20d0d4
z4aa47c4c206457121bf9d0a865bb1cbba8ae30565d8316d20343a00d824fa48d2aea7916682098
ze7d901c23e29a896515c372559e232a73384f78ac39ce605429e2f7ed9111d3e337ca647b687ef
zd092d2cf6ac88733d018aed8db3f90e78fa07cf004cae10e59312c86b5697d332cafa1ded66fef
z228df37c4fab207a78b5c596c46f520e72d926d047d7b7cd0cd4a9c402b19b58429b508af22827
za11a3855b5e5d63a58d0579db02509441e4ab49d1244638216cda2f05fc854d1f5974f7c8e58ec
z7e3ed8baab7c3b600b42ee1acd419482f9f830c021e99e302fc61eeeec8a264b6fa35a8946f82e
z31b9c8c016f9e0853fe3d359d8156a94b441086fd4b5596d87b06beab479765bea085c37b3ddd4
zcf813d93b0c36b3c48d1d732df785aae7dade51cd9e6d36695e10e89ff9d157bef0e36cb7744dd
z44c345977963171a8994c0d16d1b955ed288c9f2ec4814097d8e7d529f3974947903d5e919295e
z7799cbbb3a4d30681aee2e58cb70150e4a0976f6b4a194bb6ddea0f26e905d1c174822ecc14cc7
z3e1a6e5dbd2525944d93f17b347283bf7a617a7116bcf34f07188c4735a39301a6547e53cd2bc3
z8e2855cdd0fc07772ed70e4b0d33a21fceffffa199d0f98b3e0a5fef760306871a364c762b25bd
z845cb4460d25fcac242eb43e5a81e5c5f9494690aa2d58671c9e4365d6a454f7d02c2b0562d332
zade79ad8631bb30ddbb2a057040e3f1e69495ccc9c192522ece4bf1786341f2e552bfedd563f71
z148890f32c86b69e9f84953a8a54bb947d331ac85e236f505158e0c8e3224893aafec0f878b5ef
z570ed72cbed79df9c4d833d48a975914b69139764323e1a4ba23fbccc571e546453e4fed9e825b
za9629be9315b9076e59ff9a1928e354f2fc6e8612d20a2b26c9ed6c60a630a3bd1e6fb81c343e3
z27361bc93b87093b871075e1080531cafafe93d93d582d44d6de4b03c9f8e71002ff68a6be0b02
z01de45b968e27c19fe9d5e8af572fa5cf7b02a768f670568af63a65761d603922125763a31658c
zd4813a11d1703d2f2e95461a1701619e9c04b808f7a871efe317a67b48d28f6cb76d2fdbae45c4
z79a2b2df7b220de5d526dec0ff1228c7b85fe62b60160c12dfa82415e420684a24e50f7b9d9e8c
za0831e8bd7869b4109176ab8ae3c0235f2c42275bb0978634f89b2121e1808b27a688475747518
z582c52bf076dfee3148c85e5ad01b898698a619185e7b02ac5a1e601b27ed10ff364a4803f30e5
z3660d05f5fbcea417272b710c02cc113fbf9ba427ffb8611dd4cb8da5722f0b12f5f150d41421c
z67f9c20fd45e5b2d4dc0368dad10fd965ef45dec40ade15b078b3f1d5d5f3c72009f9259b821a3
z8a3e960a0b334975c6bc6ea3646e20f8c4fbeb2a880f50a35b9104309f2bcc502f1f2f69b755be
z7931599a0c5d49269f3ecd8898a7e41daee4a9dee3aa64ddb8621cd47c1021528b15dbe50d223a
ze6b489c5c9ec2122dd8f8b3718e7ff4f7ee547e271e91fd84b6bab19b6ea8b2880c72a64c774c3
zb4b3c3666cec851e1d9adad44656bfad8d679cbd2f316301a574032a1dda5dbe0dbf9aaf0f20e0
ze9db46a5c74babefce3bb5d46a58529475b3030409ec12a498939f71838d7b0939d86f4517146d
z4b11e89e6941d78173e502aad3814dc8031e7cacc6f51bfb97040b384f102eed02ea846217bcc3
z9a5c070f9984d8d4aac2d6936c21809769400bf41cced3636803e1a581a96c8fd1f1474db1f934
z6e3cf766a81e45db9b498484b8e94942b144e971decd6f61f24aa26b803deff9341bad23e1421d
z46ca7fdfa17e6a08606406be1f9337058243b6d4b95c72b4d7bee6c5fc961581ed9d66bd4e0bf0
z245dddc30592762d5b12dd767557f309b4724426839c88f236c55ec549e2b7acb6eaca16de51bd
z7c416ef3adbfc8bbdf7408f03ed16f429f6a23a2d7bf5ae89409c0e53af6e3930bcccd7b07ab2e
zd06e7f6883c492dfe3e9d7c8204843627e86131f14c93640b922dfc18c0cc7be87c91ad5bfec9a
za388fbef8aa0bc45ccb1a013122d319963baa40222b0f68164fc2c9d2b8cbaead4a3d3c54fd374
zf62ddc6f5a1d56da16c1b803cee5cc9af6ddab8a8dc977e8bc40d2c6fb92df9a857bd03dde24d3
z09e7bd71db9493a686302b801e329080216c0f1167226b7dfe3777ec9cc203a6747050429acb7d
z13fa5ad9629ace370eb12f3a8280960e51b2ebcd821e32ef170752fe18bfa0947d73dfa014829c
z8ff71e0de27d96a0233a0d8dc560c0e61317f34b5e51dbb0934fcb6eb9407ab1b70a35521b7be0
zfe66bd48325c94baead7ba1f494712a9ff819bb9d162c5e99e62541225880f881e19353fc6dab3
zacbd2b5d81ad08c7e67f30f8add8d3146e4a0aebaf6876e150b52418c60a74ebcf1135506473c4
zdd8c757028f6f1cacce5a7613185011dee4051740fd8a7ed69a173b60bb0e12494c39653657bb2
z94051220f561d35d7e2814048e04cf30c37ca7dcccd31c3afabaf188c4e5d47946a2b5b31b926b
zafa60ad1fc0a2abc44ae25939bdfc17eb8e6687be32cc1dc96a9c49979ad09ee5128ea0b19d82e
z6a17b663150be26c8ef1394f252dc22421875e5a5f0e5a94024c8fded6002fdde14d9b60d78204
zc8878045a0151e1e2fccacd4cd4f349889854f95da0e8011d13f3ab355b0af9e4f107a4e54162d
zf56c85f996954b1dd9dd6d37a2ca370bc269123d3d1aa3677384a6e54cc7926b75221c883ca676
z687a2740d7085ec8df0dcf920ce755ae98777f27699003d0c10b3d7fbf727d0b0f36d661bd8b7f
zc50da059e6d543a1cd19efd51c89c59e6a5316d7db10313d00e3963ef483020dc6f1d5f023e14a
z6ec07733da3dcdfbe69101849baa764a78116a1279364724eb0924743486390ce0aa5bb2fcdef9
zd8f0108da18fb4836456d33c74c266772656afcfd4c347f15136a1fc2fef92b64f5189e7667bbe
z5cfbd57abfd56cb36be0e96222c7bcb8673084e057e381d20da0fc65107aa15b963e4787ae46d8
z99add20ddb00872f7128b309fd7508d0fbf3af450b68e135eeb9b8ae4dddb645e10976ec14d093
z374990c93f0614eb3d94c8e9a977ea5a9e954b3cd65ef73c10fc6837e7a19b6cf1555c1ee1b8aa
zedd78925f29db5d66f630d24a7e65faed0922fe9aa2fbf6517adde030d4b54d518d4ac69c37362
zb4e2912ad964ddc4f244d0e81513f230ca24e69aa9cfac33deb5fe5ff465b2fd73b5f6732bffd8
z93c0a52ecc0571462d5e720a6decba22fe0d1e1124a5b25d0fbc2fac0edaf2df1115bfa9c4b5db
zc16859fc9991fe60a0e091b89f9439ef85dbc84b34930f3eb4cc4ccb023dc3ae2793fe19b1c80c
zc73ac237806ee58990c471b5398a4d2a3e4f6c1d3d1d3ead6ff5854cda68606ce1f34465a99ccf
z6b5ac1f3d0d3ca6c820dceac5b903d263dcf82ee57597a54b5e654a667bf20f1dc959e533a234f
z552b8d101514db6c2c334573123bdd888a94356d17c1ab3286ff5e6c9769702ff73c547fde592e
za89453af20410abb91a8ff8d938cedd1781b29e1349185e5247288df6118d2552bc1680736a5e8
z5bfebe845c3d46b1082aad1747d191812888a3b3491e2714a84893ab93cf926178ea44f3b19790
zaac563038c087b475cdc3831c352e81d44b62cb6936b5a66d69428f33c1ebc2921fb66154cb17f
z0939044db6bdb2f43689eadf230dfd70147975cf12ec613460d7c6a72418eec1c03c694b4545e9
z702ce8accf4a89d55186c8d344d09f19988c618be9e0ba2b2599c5af631bc0fe45e6b64f41abdd
zb452202ff62fba6af52e6b4a0e9a86331a5d7027c1f96ef0c7c864809031e495012eecb8e5a4d1
z2f5009c5dab00c813380578b3e97407797429251ba8d6dd86da7909d3ef0850f1c5964793e04ff
z9d14d04fe42134b4b5b67b19390ad80613b83f36be42e1863666361e5f1d7d88a4925baafa5004
z71df852e28f1e639cfd31ccb3085f9e8879a9789d8e29cbebd90654974e7e352cdf6c84cec4178
z3abb20c05007fe6f99fe14470c3bf0d0ba31f825582c93bb20fee5a94a3172175b59b30de9707b
zf975681a3b5590035b5958ad2b6bf81769ea1cfc6a356bd7980df69b8463efb2648f22bffb8d31
z9c5e1cbf50a9ecb7c5d046be290b805b70219433b4fa28c8ce4767c5fb0fd2206c8342021e1ed6
zfe6bc28beea46e24bcbf830c023d2ff3eb7bfe966b777469ba81923cc3aba16c6a5b19130fa893
z61ab2e64a7593ab94df66caf06818d7480cebb24d9b4374f1b301b1aa286ed87d99fd5e42bc0b3
z6091ce19eed4e284903c875b5c664a528e0dfaba55a900923597daf42f84db24e64310e249e483
z36ba4f7970cea38c505158332ef7c43b555b2ab258958b4167f837325365f054b5949f71b57fa7
z1281799bc4d5eaad5e3eef1ff6b4f74ba50ea62fa113753ee27df58308ae98bb64b5e64a4f7aa7
z0f021f4b09084f7260c6e1134330a91bbc262ff5e805a6680ea8f2e7fef1eca9f9cfd08b577cde
z2cc4caec4369296062eb0f44be730657330cc958f6b4129b15e8f878418658e5bbde5d36bccf97
z4cd8d0a3bd0462f4cc842983ce81851c1d6fc84c75c8d2e2b07c8ac6945839f9c36db32679ed4f
zc6a83382cd746190b78ff9dd50c0291096b809018fef80772e3bf8854f388b1884451ecaf701d7
z055beb4bf8be0c4917d4ba8588473c11b6f9bb129881861aa0013a5021dc82f20a566f23d279fa
z662f055caeba629bb2ec168d82d8ed9c282ac63693bc1beb1d5644adee1ee789250482fcfa01cb
zc301df30319f26a5c95e740c6414e00b2bbdac581fe50018fd492bcb31837adcac47b28fa86140
zd30e42f87ea7ca19fe459bf8743da4068edead5743201415ef189f008792c96d6514591eb08557
zc75d19c29233275aa80bdfea6874d92aff74451a3e3f10cf0cc22274f5378e0772284e3772026e
z473ef1d224f0b65655a2361ab5e264f50bba1ad3fae7d113069c2bc741219971583e46358219ef
zd098d01b3c17d9dc2ef89b407832083d93450177870b842cfaad377a1d7f4e473c75d57d055fb7
zdeae48cfbee7361d449e10b8bed173ad5a67e10e2552372804968d78425e5ffacd8449402f1776
zfa85496ff83eda23ff1b346b135acb2aaadf6f78819ae9bdb599210a057bdb5c258b8137a1353a
z76fe006a42082416eb8425d2b343aea314ea4a93234d4ca15fdfb80820c38bf426813a26983763
zd3105cbc25900b4909e47794d9da3019900b132f92b30f3d0176568535d8c5ffbf538c41d9ffa3
z2ba9288f819b6d42aecc6111bdb20891ead8484d58dd27b2fdeda0f3ce64c7543db0b8699b12bc
z63c817227b25ccb55df677a2a1223185722cd9caa0fce97f1daf97b58050174686b6e2e213e5a1
z5b14870c2f6ae9de58665f2f5010a47832b57485433c4b69d62110970482f4503fd7ed04d9f0f2
zedc3afea7a5b7bd701f9e096a843844a41ffae3a4e1c6660ed7f7571f803669d03c3afd23f1468
zd84b0294a73adba6ab1b389dfb09db0c9e57cfc65782bd4bde4e65af4c19414fb5a6be7e266acc
z1441b8dfa2d6d30843ae9a0dc37e191c4e9294f081bf543c1d06898d52d132aaab84403827a576
z03bde2e50703cb2011f12f5b05468846afd7ae7015f9e89d50d5c9e6a5515c8de0a25f6b5f0ca3
z2c22963ab04819aa13898452b02feb9f3e9ea97258ab6ff07092f9f22e31ab90cc791d90b57701
za000a013f759b37ed43ff2f4b0d76d2c3304fcf5b26bf823878456ff3bdd5c59cdfa36cb7b965f
zd8c3539609f8a520c3b120581d64a46849995154e346e05d3650bfd1b20cf8b177eb8b9687e701
z74d53e7bd1360cd718132b43c17334857c7daa80502baf92b35e9e5b95557294fbb0678c3662a3
zc38416263e77d3b98fd7aa1007461607fe05ab23427eee7d70bccfe4e0f93da6867304a0d4764d
zff9ba157f9d1f0a4a3369b02b162d5bd25bb6c1c4b7a112957d54383c17bc7d20bb8690616b67f
z7dbac278c10c6e09bd2635da2cd8e85c295973ed1b025d27025fd52812ac226181cff11793cdb7
za6ba4053248384c5ca9a15e11ee66a17ee5ae16862d68d7d3d1d75954ad2a39aec41adc8f7b775
z3a2673b140432eb93da8263bf94a59db0fca2acbbeeedb760d3842133591232d9c904ecacc92c2
z627e1a67d63af3ef84827297a169da0037c434e6a46d6b99acba640f481bb52a498381726e131f
ze07001602578a9e9aded6138ec320398cdd9b621a7cc4c9fc01aacd12e628696953f6ea296860c
z337ed6e5a769422f86cba2ee8630b6fde5deb5b22c5f67946ed9c4909b0ec0610799474a01c97a
z4f5e34f327f2f21dddf819429f93aab4c706135e03de4a90b1314a7c92f9448f234a8975323865
z5cc16e42a5e95ac6e79676692015003223eecc9e2c59f3734e38aade591d964449296f2a4111a8
z9abdbeb487d75a5ca16066d634dd3ca11faadabb8782246f9b6d712243ad88be76875acdbda29b
z232228cccca353486cf56a7047984b5f7ad5185792fad2f234864c2c9ca7dc91b8e57506881943
z74c4aecafb8d554d7d2a21c53217cc415fdee09106aeace34f256316b7cb95d6f7fcdcfc0d5996
z22116cd3b993f191c4aa0ada84052e390c32a8f03c9d6ef3f791d912a9a9c3b413319daa005ce2
z7623d734506703c4a87e8fa0bb9b9f806471a488c22e36139e8c00b67cd738116bad65b3bbb79e
z47a984794ae69de0dbfcf09b60495f2466d63d33e50d5d3407ad7910a511b75ad3098e649f47c1
z57b4ee5233a7531a5271d1eadf8ef7ce8371f9409e4ec23f841d6475c0deefc22ac46bfe3d146b
z31488d5ab12893c3516a530942f2d9474365bedc8a8a8c7c0c692734c37c726e9e5c940b317fdc
z4fa1fe54ca685dfe0f013966d09a7820543f8aa51e84af284db3e79ebd216be7c09b58bb57dc71
z0e0603b59efa3a80b9a2e890d21ea97083d1299cc81287de641f215b0e28d8918bbf8e9d07e85b
zadd0e2ca8b42d2288eb5e311a7d09d6bec60931ec6852eb6d5b141ccf9ec4c79e52e4b02b09a5a
z11a5805880aa00827960d4ac0dbd4b8a1815b6a0bb09a57893cabd23fbb356280667230f8197b7
z246307f2ac2d02af1a1205da00abc449ebecebad492973d44ba84fe4ea0565aa48d4a00f96df7d
z4dbb3247595994f4ba34c3c738b8aa3b0355ece19beb11d19662a366ea182c794c7bcf867d4ac1
z230076cd0b862b71f517048a4e82d2916ba752241f0403a2af61389ea73eccdcbfd9586d893318
z16ddb427c08d29b749e9dfce7c5ceacc537dedfabf087569f985c7a0cf8e90f93142a673ac756e
z4e789c69fc21d1a98fd1cd5d200985929bcae3bee5bad232f8b353521022f57a4fa76f5d036255
z96e43fb442bc5d9bcb9737e3cac91430bd68a2a6c14576bea43ea5dcde786b0a2da5e7957455e1
zfb5e565a84d980528ce78979452ec554c6fd8ebee2a3b052fcbbc43ff37c3540cf783401cc6405
z0d6d976eac0245b117ca68540a6908e0ab6ae8c6767837a0c363107a7a38e38228e7a160ee44f5
z6e42baaa12eaa4ccc3bb0ad66e409761aea0ecb52fb0b45600e06d0c86d47be408ccf5b94ce8c1
z3db4fdc41759b14b12c5962833748cf776d1af164e37b54db7e5c70f6ef7f3ebff3bcfc539fbfb
z1f1637a0fc7fb20bb7359ba9fd1d47e1274d2c9e514dbc102e32e6bf142185dd63cbe06cb9828c
zd3ae80a511ad77cdb931d5637cbed0afea8cb8d073c1e95ab2cb078dda6a39bb8661142158198d
z8ea3b00322238a71ef76964e3385aa34395559025efaa359a41f557878cf34bfc2104bb724b3c7
zf111a0a91cd5b87b833c5e36d7749020341c314f63b6aee929b0616d1a7c939c03a724884546e0
z63da33011d0ac72ab57a22f254b763b96d2ce87657f04e0a11223ad6375df6e147c2bbf3e7efff
z827287be31b0be75448f5927de39fb96c48207aee4aceb596bde9fc60ecdf3ac3644e70cdcc0f5
zdf01a9e89806a0fbf4475da90e95f1726b3d3883e89fab6be4f463ceca86f2e67f62f939da2ece
z45e98424b252a02b7c4abe2fb10e36701d19380614619e07202b63d34f17ef725c04c5614cd778
z078ffc1d5b489f0feb47186dbc22d3e100da8d65b346b43926f86611a44f5fcfb0cfe783f6cd70
z08d9204b9ee7ad807f61b845c55117420414fa469ce6adb33ab08890089b0acceb671686bf0609
zbbf0794c7da16e53859bcd3cdf0dc04b4be3e7aec669850995b847d6c02a8f072e55825ede8060
z80b5c5948f52868a3fc64dc7a5c7609e58081b5b99a43bbd4ad4100faba91db08620c210d04520
z5ee04cee400d2dc4c3bceb686660f91f81020e8e49ce7d627f8627461a7f5605ec6ebc2f8a7588
zf8ae67e03a0b2fe1d900b7cdead02a9fe1e5ca53917b3a5e586d916eacdb33c7d4540f00650537
zdd85e4c0a18634e1d3464bcd05387e31c11f3a2c997a52aaccd784188bcd4fd9df2fbcd71a05a5
z62ce2c2a007f7c8a3f85afde0fd67f865c29fef514f411d8a313d50307147aaeff60388ca3848d
z60fd432412fcdc5eebd8a2debf2d45800be418583e3cb6e3d000f3a0a93c709071c40f8fc7f230
z88747d5ae9909bce2a563a692430b66d26f7717c6db2282bb217fae93065434d4d7e09e1e56093
z05d2c107559e14ec42118b6c48257bb4fffa8675b3f65d6fa731b313708cb864b2c7bbe4b7d704
zf9a29e69e7a16c680dcefeb2df25991a84e360f09994e0e284aa66d82b905a97cc5bde8921b7e6
zad44570874d47bdbe3a40b80ccd88b35547db069add1bbad84a367ca4c379ca4d9e9070ca8a669
zb7e48807fc2ad906611cd3e10d2465e11509be11692b823d312a389fbfc7a7cedb867ffd945045
za35583445b5c1d6fdd36bdfeb4ad2fe65d60e2818c726ac534a1bca4be32ef98ea8ccb7f8571cf
z2260ae954e84d561310e104bb577c03a14cedef1bd96474a3cbec76c467ec91b747e5c651c6ff8
z18b6cb48607d997675f256d59f85703953e70ec15177b8a2fd0e38bcddd2b41a1eb06c903a0142
zb9f18925b4447cba76b46f50ac97610d71d0538e982fd6f111af1b4346cbc62c60e6d526349ffe
z569715db0d842e7089323cd2b4ad598759a8faef1b0724fca905f213e8bd394482a4858a9c631d
zd6d982e8d0e073c6875589de0630d3404fb8ac1eef6dc47b8da376aa61722eccb6ad325d712204
z5de4ab11de10fac6f2121ce554f46c2af3010317c317c009ec784d58c18226f5bc348392768a79
z18020bef644c0d4a9f6389d34b3e633a8dd9741b160cfa68e65ba08625f319b28d2f050d835712
z0042b86f5493254e08e45e2fb73b681f71a79d6f42e00065a385eeb43e9e218d7043d82cef6899
z939b3f7a0598872e57d59f8209fd3ea098d8907196670bc06472b95cdfd0d0971b93a3d7829557
z9e6ea2bd6afa7c56baca4e676d82f306e3a376de587fc534352f639184610e67bc4e2a023e1feb
z6fd69b31a93662616b6aef481f5f7421e22f206337c14e99c472580acbc16ba7ba68d111ed9a79
zbbfa272fcdaf2f7df186e5d314f1c5c600ae89f6568930f9c76e0f33f91b1b35160cb425598f3a
z797abf1b6d9cf1867f3cf14992356ad38f00439bfdbc05fc3b01a1392edf246ece85c3ce2b7de7
z86307793604c1123d062d03e85048c9d5a337e9b7f04b83842291efe31ae838771d65def8d20e3
z6258684a41fea1cf25d2ef1de1fd190d8498134bd3361888e5f9e2ac480498af7fe16b88621b4d
z8be95371369eebfc790c9624124750e4470a986a2c730a5890b7ed370ae39f1ab5283e4c909532
zb826668d9e23e9c87d560c92a707625890245e98f2c9e85e82eb047eb8af9dd377f1c991f644bc
zc79b3156adead9ec6fe4906014b536d2e316658f0ab28de2a6a31d363e02b07007799cfc5add56
zd9d1a83c1afc33e65403fad831f68f7892415c8db739e2c3123ea473e682e7f2b9521c9e5ffbe1
zd40025f0af267fc64cb5e9783078488dc9ec7003498593a9720e1a29084a7bb59a373ff89ada71
z8d14d7f395b0455b59335db72be72144ed04d4fcb09bbb4e66c20d1a84fbb46be5dde9de306fc6
z8913ce02f913a5e0f11bf9df02c7e165a99446ddcb36f91d48098eab24c4bb6d1f2f90a7ac5c7e
z2eddc2bfc03677ce45153c0006c25ca17ad99ec3ba6ccc4d23af64ec109f2ebd2895da2e47189d
z65b39ea8387ee4b7cdca271cef1b969c15af9c370bcf05d9a2826bd4b19024cb5eb8c7daa25540
z0b9b6cca54a4d2bf731584e1876381e91d1317d6d7c044dcaa73576357d330ca7ce82097561e5a
z2a86f0e678afb6129808c286266e075d4dcc700a6ecda2f856154f75c429b35d5777c50b3c44bb
z59af4e6b7394c17e4731de283a2068aad1af483af1032ecce06c25bd59365ae9e101ddd2f974ac
z23c67f5f0b5e638d3cbe3300039b7dad03a42ea4edf32e9b613dadf09b4c45938f1281e5617c60
za0926bd22315adc2689a69744833b771dd9d7cd8520a0f5521751a79240e61b9f6d593edd0a555
z15893dc40c57c0926ea7bc9a81cdb5392b05176b9daa4ddc53485c294f122bed851bc5f10d0ab4
z3bd179e69371a7deaef239028da9f17768db8dbe0e52411bd2faa76996cadd35b13e72af5e4aa3
zcde5e77065e5f2a92ca3652de183024a26ee7d832243aa3b58cfcc84fc4364ec0d7f1c0cc7d34e
z1aa1084da150d581c1d7b5d9f84ef5fe850de936e913e3d2653646f13d15fd212a56128f35b47d
z3a8f964f93364ef18755db2d04a43efd8bbf623b0a25efa0061355e8e30612e28f3b1aae445b5c
zf2a47b80f6d567a17afe0b0aa3b67a60a9d5fca54420d05583e7b4286f8c25f4abd174415f0bef
zdff28fd36b7bd5f8fd87a095b6173ecd15f5a05e6cd7034961ab3ecd4a53941e5dff389a8db9ee
z8fbaff8690078552e66e01e1a9107ada92abb5211d2ca978403dd82f916c1426f17af432fd2b91
z37ca9c886b6ef21baf0fb10454621e0d2ffd930ecf883b4929ce49c61548e7bfe0ee4de9e6ef43
z054cc45b858be12625c14125d27f42c7bcd5a89f23a35b95165277f4402bbec33b82704ab132e4
ze2943272d00b5da49c04452d29d08745d991dba6a6af45b46ef74e07402e07742027770e3edacd
za778071805888d69a946344eee80d18ed702472545d105a776fd218d365b952de58b842e5d97a4
z4b8e62409cf5cfa431f9b24c5d0a8d1b3b84fbd6b629a094452644368f305101169f355dfc6ba0
z2f343021fdba269bdc545ca7a67672931cab6cc458195178eaf504660a45ded5ddb1ee25bd971f
z09f230111f0e4d8a23213fb7081e64d57814ca36b376c56e8fa9c9416865f07fe842c966c9bb08
zff3a996acf06381df7bfadcab0cca04c7e01d595166dfc1b203913cef483c45e64b2b8ec451a02
za64c7a5577e9f5f9bcf5eb9f0a4aa79f24d2d9644cde972ff8ccce5e071efd677a041acdef712f
z33b63a89008bc95fab7d6f7c9aa16702cd6f632d785744ea207ce974be05d3e24a013e4f3153f1
z45820b6cf2395fc86408c3f741cf0422b745befe071134934eba40b5cc5f2f74fd9b8c0fdbae18
z065370ec31342ce417316a9701cdbd4bfa7596014a3072c6431f09b70ff1466833dd72db805608
zd094c8d9746acf51ed14ea2ef69cc5a527b650c9a4d901572bd1443f3a20b3ff5c1c0bb8786157
z09085a2ab66d989f9388884bb50f1340e0b8dfda741648b5f7ff2c210687a6f54a6e0f5b9f1d42
z1f6e157fbc4ff604b9c322a232f1e75cb4ddca24a40064d9a46c57dd4f8214ccd7bc94d32b783d
zc06be0d934af00af468b9f21d4fc81be3ee9a2b8349477b49ed6cb0a50e8f65a567405e8cde6ea
z5d00aaf57b82e1527e6446c0c3f23830dbc4aca53929270e07c63d235653023ecfc1e4f5f80284
z3d1dd36cbf45b97fe08dcb0fbef3e99bcdbca09180a45967d8accf83a3637f1f054beee1043dfc
z94023d36a272d7e9cbe5b31331d6415643e0d32841f30424a7c60f1cffba8a89529740c2b6300e
z920787eb71b9c5d3d494a118ce1cee1b4a7ec6e2c032986c9ba2d00964ea54da6fecb3c69fd45e
z8a18ea75161316813ff13417269924d7f2a519ba98dbe148133ca0d1ce5858b65665cd9107ced0
z22bc53912dea91443e5b7d959d50b665da2345946c0cb54c5f6ecdc02492213b868d517ffdf8ee
z2d484ff84df1884fa0a8d47eca8598adef54efde09b52cba1f982add1cee99be10b6758490e01e
zcb3180678f16b9c76d16c3c8e0bab4d56198530be6fed7d68daa2cb7833e7eb34232d95dc2a120
zb6817c7c74b9fe70713808d2da1d1a24d2dbcfe16998b9fd724d2a04f60cd274e102973d9ccdbe
ze44fb5ee8e289bc9df05b6d4bd40fa3c8fdb478eeec51b8468946045b803a56f66f4b51b4fc276
z4cd4fa342015a89f01b528bd38dc375524d0033bc8d128876df2a0acca5aed01d4f7af550ef30d
z135d05143f890365060614ccff5a31adda588a1c44f8136681c87e0e64a2e5a44b99d16aab2a48
z33ef10f0729a21853d50ad4f051cfa0c64facb736c265e05e13795cb48b26756a449ad25e1fb01
z6a8283d5cbfe4a6388a1060f0d93b71f98b0dc9bbd3112891ea62283259c061db51b35fd5510eb
z6d2a9720ab606110d1a246a52233a51ad6c48db0eda96ddeab777051f4cb9ad331eea757e55752
z2f3a5aba17899341a2630a22572f0bcf48300a35cbcc2d91c113038166a5cc557749f3d9c9abba
z6b29c1fdf4ef076d4a00c117153c0be79cf0185380cf22063badd98e4d29c45f6a80694406cbc6
z59dfa71174687c669b578db909e456026871593a4a31bbbab106da358498cb68e80f7ad8000839
z1a07b93c224599a47fea738355f570534fda90313039b03f79c4e71d6c9b0b3f4f6788cca6e4e4
z272d60a11c9693e26f95cca529bc18c999fee0f5b75105eb7490dcb38ec97047d7024c5d6074ba
zc2d6895c45dcbc335b2145c3e8793c3996ec53383aa0dc542e6630f3fcb614206cae5666c9cb57
z57f12e3c3048860d6fa9da1477e2f2372a17e8648a48451d3f6f6d57062c618f53f6a04de936fa
z55f8826630a0fdc3d211b407284eb4c7463e35d50bed73e65c4cc97c68e89db3ef614fbb160f1a
za8eca086f60f1c0a52c9e4368acff9fff3930f9416915c6d1f8ec4510817be4b23400ede48d77f
z60761410aede5470d08773d14c8644c11e344df4569fd6a9e563a4ce8eb0230a1f27ba7b8b7185
zd9ee0197aa0215c408b6389f208eae8227922208ff7e6ce41a601e7347716552a2a092276d6fae
za04759a48d72e779d3c62272f96794e8ddd49536cf0d4469e2cecf68d429a5d42ff8567e1e9639
zefcfcaf1e7b6b89223a9b7817899c25a1adbb442c755688341ba0c171f797581bda6b7de16d8eb
zb9f80829345e6cde830a69d29ac9b09d8f0a99b506fe8f3cfdc4955ab3067e42394245e5780f94
ze324e1e0c4379cb8b62078c8871646c7cef4f9a60667646d7fa97b329b9f6869e1bd5e6e891798
ze4dc4e97ff42a6d3270c6198230aa56a9e37cf53ece1805dff1e753769be2961b72aafe62d5064
ze339c39050fda54ee45972b59353e73b67ae0c73fc4fea7b58743a92b9b634898c5b32e1c960a8
zef25da4f1230fed037901b4a560309f4ce8e0b642e22c70bf146f601ae16bf7ed59f19a65da3ba
z39855b25bee73e7370c9876f2d4fb2626723c5c3caebb195e85d96cceff1a4da1a01b4f3e95ec4
z9a3084befa898a809319432b51f50a5b53b9651330b80037f0fd799f57bede95f7635083d4c940
zc90b9da6d81fd5b9ec83b7eb7c6d0e988d60c01f773cad051cb06ad56801e1cd6b5262f7add323
z00712224e2a5540f40013740d775c6a1531eb3efa14217c3d716f8a977dfd8d9631ad85e6a502c
z07fae6d59b5840ee8bc3f4c59b4013fcbbcb5c161c6ac457be3d9f9224150c09b38845436820f5
zf28142afcbfa7a5f8b73a177759cd823b5797bcfd24ea44d6d184f5fd18b97e2f3126f19e8383b
zbb804764ceca966acf050ebb62aeb9b035e3287a8e92d104a181e0afa734f59f8db994016f67e1
z49e9414f6425e4e897d5a04bff79e3c5918554e858e76b2125989319c9f528a4df6ee83b8d9fcf
zabc3ffbcae2deb6502c81857468b7ea98bd6f85e67ba10a17f627939e3886f52bcb630d4c76f21
z1c3ba17fe30a767c01ba43fc8ab881448829ce88e705f3c51350371c9cfb055f9711cec7a9c270
z6e51beb3173dd0ba0827d8eb8be31646b4ccf3883940672f7e57ca6a68f4182cb1c462f687d37a
z02ad49738826d24734fda934ea2545b0ae7387c2366fd12367d567d5e1a8c1f2e26a3c7bd70c6a
z3911b491b902daacb999670f3051e8a0de658435e081208ec4f1e7ab2ad6c7572f12e425bcd69d
zd0546c130d4beff24715851e211d7304753e344616ad15225fa7f542c97a5e9d025f76044a3735
z0865ed5dafe34369f532446317da86b9440576bc25f347549bea61d1f5a295479f0f6053082407
z3984e3b95fff00cdbf11d57943eff034fd2c8bc30cc814399364034773d8a180035015e6bb021e
z1260fe6df3909c63c962037a1957bdf85b1e44e92f5b5ecb4f456d5eb3b13596fb546de6fc2fb1
z3c652bea9909478136eb5375a3fec3ae63713ddc551739e946ce8787db8bd2678a331ec1d66d50
z5225c154844aa6f7fe2f6c00ed481803f448113162a152187684f83578654a32882273fb202c74
z43081b20722f796e1ad9cb7d348c0a99a05257fb3901074bd66dfa709bf43782c0ea245e5fead1
z8a04479fa68a35ffecadf05f902092c8796f3a6c121325074fec9ca96441025d080408ded1186b
zfaed6c7a8cb511778777fe331faaeaa1c2d60dcd3d643f0524b43040ad2a3cf180ab82b899dd5e
z76ae1df6f1083d7d6557f05b6db4275fb861b599adc3731f1a88cdc224e91452982092d6fcb0c0
z2a01e0c07795771aa09dc23e914fc21b9152c7842016ed30f5d4803c70dd1b891f566740cdb86a
zaaa2674b834a875244e4102c79ebb298d3ddd462820e22e2dcb1acd3af7607995b32f4f968399f
zf15fafc4ce15dbb67e80ac415c80a179c1f38b991c74dffa24c3d32638fa4243c727ae655dcd70
z7706ee8e0d0be3eb6299dd3a7e28966894d2af3243d8bc1ca4c89f73d0838cd2f4ec9b399b027a
zccf83542e63f97c745f37ac633e083727501c73c4de112da4ff5ebab9092f6f680865f0a5d2dda
z08af92bae58bb92d6b7cb0f376ce5d1257ae70b524e63d8e02e30aead1e058b82c253bd57f09bf
z6ee26eee4894b9e11b0027c699c494201df7e1644c6379f51544540b1faed094c05ebb8b0a748f
z329ceba21b20dc5e1d0be4e0c30bdb020bf00557410bdb603d9a2e0ad772eaa309686292b24552
zb0d41496978e5279d569d7c44868257312fa4208b0b14104eb1f218894428c3dfe0a606afeb40e
z1d7d9dceb3eaf800f9660a009ba55452f35a6bfe7ad4943217d6252a47aedcfda61414316fd299
za4084edd098e606ea97484981b2114866eb6852384b81e7d64bf03693748e201a872552d6d4f49
z33962f5ce1156e8d51af76754b74b49737748a8c3b0b4ac442310e3fd7eb699a668f0beb2fe210
za66bd08c1721d0015646c7c09441be308211836a7f5cc309e3979b34f39411abad97506c0b3a9e
zfd2667416e2ae7db832f21f730ffabf99e9cb9106a344b8cb07df53423632c9daef0c985572d92
z6904d819174c344be809b6260734d07f75edf93d3c27d07e256588fcca3cf20e0244318ba0b071
za40c8fed1c1a0e7a57d2c55c7e613161e201fed011fa91c5b2a9e528f586b7502c81ed79024593
z6c337fec71433f65ce250314afce0e9af6c56dca91e617e663096422a5af57d872ea9df951f77b
z47d8fbb021f0719678adbb7e2b464cfdb90bed5737a596e094fe3ed1f42c6666feb61ddebe1498
za114a801c13b2c13303a9836c61c8a775bdea6abee8da84864629818a6057e0c7cb2b6b013e4ae
z92706d3ddb32ee35157db4c299044fa2f85bcb32c3ba9b671f924b44704d56a1fa18e0a5572437
zabc5659a7306ed217bc385088b8212ffacce89655c6a4439426ea1ed31445198ebc586b8dec94f
z7569eeda87b5eab8439e7e105f4d53520bc01a78a7db92b211869cf11343586026f9a4aa584167
z9be47a77b317388e61ec367346c92725b9995e74c09166d5aa4670779c87e61b465e153771a8f3
zad0973ca84f3b385e09519b5c87c6216cd23e5b49f3a5426dae3cdcba57cb819bd75b8f6d64b58
z96b19d71903fc61338a77ffc45091d83c38ab4b128896f8b8723b1f2bea14f449485fabbd257b6
zedc4dc871fefcda952d7bd0488e6e0da19eaa640fe8b60a53ca2abdfc5a2446eb6ba21d59d9081
z48ae5d81d113082624b6aad2ac13f7468563e4c2960758316b2e6d6b404bdb4134d8738ca75f12
zf229ea572e96f7b382fc8ce63c59a173f6ae0c86beb951ab5c9109625f8889be7c2fb782c2daec
zde27974d780f60cf4f3f88807bd27335355dd971032bf203db06093e331e05bec793791474b1f9
z50552cb245e13ec68d60ef13efe02ae93142b63cf8dce2497aa99c8d2058585c3817f9d0c9b1e1
z7fa06e2dbac307c8a56df48e51b3361fd872598259123c2c46840a8c4cc7c39582428e84df29e8
zfb5c211cf445ce22bcda9ea238293bc91621f6fa96a6fc7e6fbff8c911fd2dbe47fb89d2e8edc9
zf4e6c23f038dcee8545ce7de325a478220b9d8c253dc2de9dec2f834032a5eb7fa22b4053885d0
zef49b34b82d5dbdcfd060a8caca608aa61633790e4f23b8e0176673ce3239ec9f6297269a72aaa
z04de8d08c7e75906cfd789ffa8b275675afd04b80f64d48dd50569cf91505335de93424c58a562
zd3be6b4cf7c29221b2d684b9f5f42954c292a295bd01c1838d0291b4a383513a073b8c16d345ec
z2b31461cf32f927808b8a4c62dc9e996c55d9028949444bfce600e5b0579b0f4b012c56ebb37d3
zbb8daf218c5c1be1690c402c66880bcf45f5156bb0ca717e013f2a60ac1da891c1fcf3f27ee225
zc2fc22929a95dea36b22a063cfa9dbb3bae218bca16d28d4f446addcb1b7bc6553447128363358
z5aeb9153b192387b97c9a670dc585c12861ddd1a7bbcf1c4192d4bfbf76beab7208175d9059785
z355c50bf6fde4426ee4ef4b06798fdc81282938d68b35687afd3574a89ebafb30f7b8c239d1928
z57ff3de00ecb425598167d4d6a60af3cee46d6a10b850911028a65438aa3b9aa3747ba4762cafd
z59c3b776e79206bbab6b6077c777cc7374327202c2ece8976cec810b58b5384643f3b11f406888
zae9907693f67c64da01afef427a4d7ad6a8edd1247084304ee667c9a0bcfdaa8babea4a61a5f2a
zd298aa6fb2dd85618d459718fb459396591d8c3954bb5ea9ecfc0633f6b3d96695a34bbd91ef05
z639a49eed0c0013906f57a1aa537763461119d82aca5f625fdd468582b047c37a4f48640a8c064
z4496d397777c9c262dae7ccbb03edac58ee67340e4aac3c6596f5b176dd8db7f1ab091d775d5d8
z0bddefd66ebedcc2aac8bf226d34ad812cc292257a8aac02677fad081cf538c391e4cee2b49a59
z2248b6e06f5a5a177d0ebe38f32a832b3dcb33bed4440bff8194252d7ab2b05e154b5e56bb33a1
z1117dff4587cb8545978fce1428f3ca5ec63abb0bb648006a997bcc679fd8efb074381a159a043
z77f3d82dd3bc7bc40160ac311ca9cf8e177b34f437ed8cbdf9130968fdda1754ec1077c1cad4c1
z48c03095b66f0b3e3baa109337da9f40d43992a87da9cd56cbf0852591e461e9049610fff69b85
zd573c18d6317f55b16c8da444a418e47df52bf3353023abf4932a0d5c0480dee2ce60ca622175a
z4d2c51adfb46194c9a0a0d1dd07998792960ccc9b6a63529ebe0fcf769ee3486c1de835ff13151
z985ac2253be86aca8df5e035a141d883cfe75fa1717dc2c6e76cf81c8345b147f565d7ec7c7392
z7e16563d7f505e101c3d13cef62d3edd4b93b2e2feaef4d3a6b104bfaafe5bbea97859da832c91
z401d8a6c24ccb0b9fa3c9bfe214537965896da349c372b570631ad88e5d03b37f85c77598ca3f8
z4c5424165654ca121f248fec3b7a5df47709826ccb87084aed6dfaa43aa4e476a69943d13751a8
z6210d689d5bffdf31a5705e1567025a0b9097a0f06ca27689e95e34fa7415ce49b27b973c95e7b
z4cb4c51067428092524a405acd9978f263bd7df1b436f44875e55f4875c30e4a23b9479bab1c56
z6026d2724d8188c9a2ff0c996cc4eb8d98d68008ed30f6bf040e962749c46ca6abc47306380b7c
z67293d73ab65b8b5c5417b07b6980ff930124d70dcc1e4514585d2b24802a30f50b43c6358c0ff
z148cde28079ef71eba332083a92e0961a30f6a60f2f3e838a8bacfc22a4ce1b4f9c46c24e0dfec
zc58a788060e23182446ef1e07a311d93f4845cf135e65c2ed55521f84526c8cdff98be6f0fa0b6
z1888656366e08383d23e86ee1f9b4c728a8de6aea63d6405da54a23fc2950ed0e915b241602676
zc0e07edc8f510bf09d0646270db7c742d85bd8ac6a17cd2f77ea2e6e76fb9467e451cb04139bb7
z751ed0d53eb21c095529d71e7ba896a5c12b3d65b7b06689ad35bc752de02e18e365f69797a3e1
zfbe79ae851d62949be596f6e5303179f5c4819d2a26015a132ff0f4f0c67d28b16323c6c45ac01
z2e2a58b0e8b306a06ba519098ab0870e73398f67ed0c0275c1b6e66686ebc8c6f0ce6fcad01403
z05f7c7bd78dc7e9d7e6b5036f89b45fc743bb8d973db260b77fb662e3bd4d25a8fb35ab9ee2850
zbe25d5b475728b36131373c05c0681ff8deb38ebd030b4fc59e84e447391676cc527c66d69be10
z0fa423eb230438e9663d1fd42d45f2b53d0941cf1035c0d1fc659e2c29fae75da1df4e4376299b
zdd837c45501b08550329aa9c3c47160f11b55f04b7e8f815864e359cb5852137fc9250db6d83c1
ze0f89e0a2b2fcc106c98bea3617313254f55708afdc00cc91c01fadf904614988a1e7594ff4c6c
z4f7de69d452a8ccdebeedb07b459b87e7e973041f32d2743265fd20c7ed51f60c3072227286717
z4b7e479494bcf0ccf057d3312c81571ff35a0897cc700b2bf58676522dc31221513912ea657c2d
z8469c97b181c03d7f1f2c9be963aff9361d57f7e168e0191754aeaa0e708020d09912a866e3d1b
z9eecea22adab6ccdf720d6a12fc80ec4600471b3a331d6f9bf41a41936ce1a2661fdd382e6b88f
z8b563d505fe78d997135157c1cf0118719f533411debc907c9ce2b4b6ecaf399a454903fc37e2a
z527cf81e90b8324063c2e1f262e67ccca802fd3d1afabc54fc1b45257135961302d7a34d280489
z1e6faad78f921bc66dbd700903e2ad05464a311a865ef10d7b61c38332f3a9e5f0811cb811c5f2
za671f7b9144472504973a319fc0820d47f23a80b56aba1d61ec4a6b4cd7c1c11d5941fde051ca9
z7fcdab88be9bd12cc4bcceb480c209e21a2187314b8740ccab6a468f444261f979af6f1a6badbd
z87617cd7007bcfa3a9f28cae1e25866b4fa639dd0caadc8cdf2f9b31c0ecfeeb3e7d7459eab406
zc4d6c2b56fea7306522b3d827f25f7bfd07930356f9524b54400d9948638119e51665f3acad442
z3667ad74ade7ee752fad8ea984b8881dda134192fd6d73b572de0ae142d5f246ab699cedd4e001
z55f6e4c666309ff08b18beb825070c179fc542b15008f08a0e51e306692bf0c6ead27111f3603d
z9afa2ba8657feee486640c9f74cf23bb1bb62a0c6d07e3d8aa4ebec4d081448f57676db85d4f66
z3f97d0128e70f44760f25193798952b3fd51dea8349cd227b879dcf94f980abe4957c5ea542000
z769b6d246e9a8876f8d424ec1ec397b5df02bd11106a9bd184e63493750516d17144d26f91d944
za398326de436df67e6ea0149e2467f404a046b7e0f3ff0ac96e3f0b0ae68f5dca52acd41e5144f
z7c8c9d5888c61257acece2e953b92b514be72ba34e4cfd5b4742afcb37beaff4c140f8d157c79f
z4b3e7fa05a7f78555be4d119afab245f1ea0923a31b4f076d366e67e619cc8116dc5379648ec75
z1d3c9d203e96dd358c19adde0f32d93d42fbe76c944eba5775c199d9c463307160eff1ce7989b3
z1b196b70cce0a3906c9e5cd22061563482c7fcbb258e4ea8e791fe9223f6bcaa69c61ac86bb619
z1cbb282d64b497204eb3fc4a98db3eb6bd8f572e0b53eab4c8d034a20cf0b065e86a914b4b16d0
z6fc632b4d9c862bc9d454e3b1bf7104fe4b8b7b1f49901a203aabc17ef024d8dff660665ec3fad
z95bbb950ed8706687f9433d2853c44969e0b7c09c38d5263adf7133342cdf061ffb16251d2849a
z818d19a23f129796eef2019e55825a52ef3f945273a082b9363acc57fa3de95aee135c563fdd87
z9ef23ff0687551e597245ef834a756f03ed33cf3115f58914ea789879cf68b9827bb0e13a0ad57
z1ada45155899f751ff47676b79bd1e8652795611d9b03b10601352a939d4fc5ba52e8c61b6e607
zf3ed7538d7310b584d8ef84ec5756e6548ec11ff05cc43b0d75a67b66fb58c62cd253feaccd56f
zd474c0b8ba71b65187efed5d4e5d594535764e0af4e32cf1dd085556110db08cc4589dcbdf18ee
z4718b49ed6d8b61292a5161beb98b21eb758f9cbadd8ae0e1ef1cbb6fb01e7af33917cc3a9abc3
ze5b865062eb96b2954a193cd2dc3d3f203ce9ff75b87c95fb01013f4d3c9f846ec7ee8eecd2504
z7366cf5586be582898af43d97a02f1d6d4e295d693c9938a31e121202c18dee705f37e84024213
z4254ebfcf778d0a6ab1e584abc5de279602141ae88ff02966378536b4590da398dd1710d686191
z5f2a2dc126a448e861b1112227a165285402ba24788cf0aae3148d1885689c3eeb24b0e919fca8
z89be57bab9bcdcae8781feb05ebfdd96e70094484552477489f3da0e6d836368b29463c7b14622
zd6ddc5eddd638493006d1ac8efc1d873860f1952b295f7d29b02ce7616f6f4db72fa565a08c087
z957b938e37c28eceb70b8d7acf5fc55750c05af710becec690d82a606a9080268b4da4aca6b71d
zfc865dc20607be94ff1e4a7c9422c1b9651a55ebf2ddcde37c6cc16ad6c5baf271974b8e46df10
zaf92e5b1b417eae00a25ac973bb3ea805ba14aa116d6e6b54c996ea285674cf5c4b897d2ccbbeb
za259163e13ae0c8c22b7538e05ec9c35256650f95a5d9b9983ce65a55c9cf769a72dc39d5c9ebe
z6031d42dab69c8a7ed3cccc13259aa318d0d3eeb6d25750fdb694f39c400d7418481dc16441000
z393a79d43a2b8aecd78f40ede472a7d6bd9ff4771f81c7d9d0e4e4d1e3221a3b2d215849244fa2
zbf04dbefe0670f083d2eb71c8a7d20e64488fe05ea7d7bd7e8c368902b3c9a88a54848a8096beb
z78a5b232db366fb9897fa3e38249b74428b050292d8d6d53000b57ae3f5fb82b54fb8d2e9af3a9
zf35076c1e2cedb2f874e418f64349cc6bfb36e0f99b1a48da3bc62106fafc555f73d22c03171b6
zf79cfc30930ecce5f37751dbc0cb988f20b93335bb997f4c1461b0739e065c68b346a8456aa9bc
z854fdd1637e1c930efbec2cdeb3337e4a21d92cdc015226a4d67d719d506b9e6a49872b1d87aef
z7b0e485627e044c7f2e048d455d057da918860bfc9a8a9cb05fa447649d7a7926097ce7bbbf465
z0f67b270df5af594dd6ed0a4c224fa0134e889ccdbc9e36a6bcd3098e6fdc6cbd70871ae9b7621
z7b9082beb3dab2a335c1d5cfabf1253d6d69affddb4d49b50864e74d398dd44349b43557c37db5
z5ef6f65332ffdbb7650a4976b08787de84b86aa97d15774034732be0a575bd1acaeedbf906bc43
z2c3a8efcf322efede236311983d2177cab44948cb4515bb6facfc72ba7cd5697101dceb65fa5fc
z2ad0e36acfb8ddc14fa9541e70e56b2592cb8bee4dde3f4e788c6275a6cf058f0aa7a415921bdf
zabb0cd33bdf655c9e7808a0e23698df1c5e51bc1b56f8b0be0df436ef07a248c950795cd0bd951
z812d7fe76fe2ef296b03af44040d20b6c4ece72f52630f8c46982e6ad83bdfe61874e10e64fe53
z7cae7b7ac7b05fff20a1d7c6e030d7fd941cf7684f596ba75f72a8685583decb53efa7e32eaa1e
zcbbdc51c4953a2735594a0ef1d9866b96e79e76b70fc37cc472211d43dd5e1059817254adbe581
zf194ff0135ca04e3d605ec5390b80d631009caed3cc9e6438740808e0354fe02eb686099bc78c5
z3783efd01eb603b6620004cb1e053348b711036a251a18f4f686262d91caefa95b5ae3906e479c
z4ca8bbd489b14d9e99489fbdcc8c441c004576101293022befbbc02f999446e4544078ee8ed0c2
z9d4ce77968e506e6e39651388a7d56b862e5bb95801c7b80854432a2f0763991bf135c84509775
z65e7eda46c0789e29a048a8abdb0858da6a298ff89e11ee3a364c398729494e5c7532903372422
z39addfad5f23e728c763357523716d64df46b5386cb1dbdbe16a3418728275ba86381fc9ae6a68
z08dbab83acec6af465e7a018e1c968de0efc3894ddae32f828c655ec721d1e082aabba73b137f0
z3aab17593e09ec93afa743e3c469b3f2f6d320c58dd9310656dbe7d69bd13f88dfe6a1a6568697
z34ca64767d11e8d75c8dd4055e7c6f96a83062fac1bfdf92d9201fa9963846127aa93d04aae02d
z05d566c1dfea7dddd5f8944a0558003c84cb7a12b2096a0c78b78b7dee6a539da3ef4929120798
zf7e735b403cc5b0ea8e50c1529152a4e5572bfb0a904e959a173416602d2244ce2e26d8454d66a
z1f3b554aba149c030938bbfce1c570d25b8e388832ee225ff8f4d7d2eb80468521cda77dbace35
ze0bac5ea92ff5962cc02e985e0b3263fc4e832f9fd455ad2ac8d1b16d365bc30cb60c442174e02
z1ff38229abf9c07a8184abbce53debd49f00c75d63930e8c3699474bd2c065d7f34e0acc0433d1
zed836876bd456db7d479226ff36db590e8a6c7cd8633d69bab52854fc6d50d6261751ca0b2170a
z11a9aaa38bdfeed1fd1323d8d9c904542aa1b6c4ffb2786e4f6db0bbca77bbc3040f1c2ec543be
z7f8a50d230f9de67528c0ad3c8f8c40de1afaff99ff4b02d89cce344b9c7aed56fbc3525534e45
z1f2c7aa85d88ce30cc963897451babe1d00e9a410b6e6a09103fbc9d47f6f06dd8f76dfa3b2033
zaf513c7f0f263a17de89fde2458346f324ab45befb00ffbe6bb6daa025631fa30b3aa13b27b643
z9e6f8a7b8be30d7f6eca113ef4d3ea8a19bec6ec5d27f76362ff08c373990e16a3505a9d0c9bb0
z06be309628cabe9b6b35d53f096556d7787333255031f5986f500f1ca29c1398e1ddcc3f3c21f2
zbd3a9fe1ed4fb646b371566f5f13eff69df90d65995ffdf3217bb19d120711bb8fe50fa28e4b61
zd708c2ee62f5cfc29bf3268a0de70486576912de44e9e11834d52a1ed27a9205e323577b08da2e
z23e2034ee59d1bfefc02d959e2f64e847f9911b7d0f8c8491c76d67e7a12b900d16b6292c18a91
z82699c55f1be8918edcb9db5944f6e17f99558e119141d51fe5d31534cae2d3e0ab6bc1e3cb257
z41b09c55949f5f71777e6c676168347553a4fa2145eeb0f7b9ccdaf3e87912f48f757e7fc885b7
z0ab0092e1702ec431d69a23354bd686011df3591eead60d73880b9c520c6e19cc24a080736f85a
zab24f9bfef65d1549066c28ece457df7e4f7b7c47b80d8dab5f592f79245b2b6aab45ba8ea3bb1
z3e134a06ceb6a690d14ab7ed6133438f7620cd9f423ba306b4722039a3af9d4cb4f64909a27627
zd63acd302ce0c4cbae05f9638e562c904745e655d3171ec2af5e5ba1f618fb4912f633f8cce950
zb64334e4af0e66f78c99b1c78fb3e9694da8cc0475a6b6a619bc92e1963bb9bda2bfed806b9f6c
z63073c9130ba421c044d94185a6ee7bbcc3fa11144309390c266c960f0aa94adfa7427ac8d5655
z6aedf29f7131388e75ecf1287084cddfb9e189248eaf73babb77b9a589cffb6b497cc2bc9c4b7c
z5123b0df7b6a722399fcbfcca20f977afe174e2a1ebd22fb3ff07454723a8f4c53828d4682729c
z0b20f2846f1318f10a596d0271f51853dd6754c4f42f0a92677058dfd5659dcf8bd354578ab31f
z16b3a553d87488ff3cf44d68cb2af0e2e785b5b189ed2640dd4cc0571786b8d04bca1123d8e324
z1c91bb39ab6623fe4849d477f79e760ebcb9c979fcbe740f35cc693378e81bbe38f7608bc45807
zdc4f8486d6adfc237dace9667aa24c0c885a22dd11ce0f9830e874366a73506c6e2ceebc315635
z853f955447da6a47754f9578ab0640a5a2ed66e36d51ff9468813ee19a11e34785e1e70dc0e6f5
z7e4e656e0f5a435311de04bc8b1f0ffec352444ba79842881a830ff0dbcb4cd98c10ce014998e9
zcd55234de0616ee32cb0ec7099fa40ddad8a96e251871c29f2294278f11d2dd10d69b110d6dac1
z527db68451256e81156189ffaefde205183c5521dfbe01f457f29ea7b4c68657acd7f993a3abf6
zf8c947c873abdfbe72dc1e6799ec12a33c07d5259a6e5db283a854d93c7f2f93ee8278f0e5f2d0
zcd118f69c1d4e23bc5e9513dd027893c297af2e17fd592e8db33f795edd444731b78dd7e24fb69
z208f05535d85f486a833544500aae26ce995a1db477c0670b0d355892b8c0a72996140378b9a38
z5370f9ef3b68585ba9f851e590e79ecac0003e4a822315d7fda426190041909c01a4600f8d9f8e
zd9291f57b22fe1d87a09320dee3f116fab3ef46b0ebba2d3fdaee5ea7dca8081ac828f7ee54856
zccf0a0c0856c23645d31219a896c4d32cd24eae9930f9228a0ece95d46932a2598a45860f29ca9
z496807b0b44d6a9e4b9c8bc91d8aaf27c9d1ba33ca9f4e4c6a9ee9a19743afb37b5e42ff417c78
z9d995ba7ca8be62b26257cfc4795dbc4ab7541a59179b4e14d3748587b2bbb469e59ee63083caa
ze8756ceac0866223423631b9475b2094ab7133fed4146fee2975d88df4e433d46f5f53f27a44e7
zb6debae7a3864c770912c0277cc3f6146c1e1594926349f9616c13026605978a0cc74cbf5b21c3
z8f7a7556f298aa8fc16119ee34963f7c68fba5d72dbbb4fa64161d46c2bc14b7f62375a490e64b
z743d01e352543356a9c1f119bf11a75423520448c9de648e95ab9fffb36fd0a47cd547537b4db1
z04777229398aa48b61297aab1adff930d6c41c119889ec8cec89eedeea93f66b7982879e483814
zb971036a9cf98262ddfbea028b769834d75bb30e104b374addb110af259846b0d1284bee841c38
zf944c0346510bff39c12a77ea3c6c66c63766fc0b11236dca5397f821e0d61647e356e98e1b739
z9d59439e8b2e9252adea3d4994b69cdc81d665e9c066efd500d10a2b8835e9737c54e9ba550d24
zac429110978e1c1400dc64f6c1e027298eae5c1ef7484d1dcf684e8106efaacc8f775bdf2ffc05
zb677a7da495c0d2681a827273114875ea551fb2a3b881f3fe65b58476415291300c794c8cbbcc1
zdc357e686a4a42a15d0d876ed75121cb08880d77167b6a0a90f705708eb969d8ebe9a9f27035b7
zcd162d32bf9fa8df762018bd7671271ebbd329396862b629383897a7ca959d48b062fed8b5e0c0
z05f5536e6596f8d3cd55dad13e1e561812dd1156dfe4cde7db706de51eb78ea2ef76052b750dc0
zebd49cb18b3a9f5840b58ed4074d2dc4bbfb9aab979336b9730bd709410b8f010fbc51ec2dc134
z374f7582c51c5bedab1ffa65764e5e83a833bae3ee3024602722e5bd04e899d3ae6af5875e3f8c
z0f1e3683a4ed15a020a0549792d1f077eab5cb730e256389cecbc76bd34856b50c2279de7ece28
z27d0c8035714cf6f8fe869b2a1149040f422094f8e637e19db87dfc811932687cb6c915f90d5c1
z2709f05a234fa604e35578a5d99d324350feea8fb3f48adc665b88a7d2564956987ba2b26b27d0
z01e2ca0c4a2337334a6b624e3e8d9dbf040d523c2a59be093488959116cfd505b857609bfe2d74
z43d9f7fc4f14d662efe3459854258ce96c6f6f949ce371e485fddd1dd6117ed299a4140c4fe7fd
z8c79ee55bc602d2535e824337eff6b9c1b928576b74b490845c1565b58dd38ddc68d1beaab2e82
ze38fc28db4b77e963febf85008f4ac78914e079ca14760a7815fe1fd915971fd7de86e4ea053b1
z9c25dd6b4a7cf6ac9e6fb1272d3117e0c3a7bd0088dcdbde61b8fb75480b43bf0bda595bb7c2b6
z3222ea2aadf8e5d97d2289664e116a5736b5e302c8cdcedf15f31786416fbb6ec319d89fd26156
z68bbbdfed7094f87b50f4e42f44ea016f75c1275b0fbf923e4b3ec3d63247fe220ed32723bfd20
z57f39c2fc9c9358d6513ff6acc35184030e71157b800c84ce92b8443d63805911f1691236ceca5
zc51769a922cfbd611b8e92f732d08f7ae460b9e9939d1ab91b93def154702a45068dd559a38183
z97df80837815af9b0271ecb224423b4591941d67625dc38bfbcf5f04106de8700105865556f8bd
z3b8f454ca20228bc61209380cd415f706d2d4b36f6cabaa2b2ed5edf35f7b4005fbc02b822a999
z3c8fec34ff258c1b856ecd20f9544907f19bc154ecc1f8aad89ea45530c627b39f0341a58ac49d
zbc57c16fdb67c248f6d0fd9e1e0eb82744cf959f6b238303e665a43fda3ef251aadbe9f5415288
z14b5b83b6e1d7e13859069c12d2a1639f0047727309dfdbccff17d334bb54b87af37aabff409e3
z9b50fd8972b67279f2e58fb979cecd8cff1d8ae5885017c5ddc1d17f16dcd2718aeacb4e1d6de3
zdbed836372b604093a06949babc0a1036905de28b26203638724f5f010f3ffad7ae2061597913e
z8336544b7ecb1148bf2c32eb0450f71d1428b3f51f41f88e1ccdb684ba009b0fd37b945d26af8a
zcb1bd5bb3356c81b90be268ee2e400fa9b47da9855872ad32baf3260cc465de6c53e1125c05c16
z76b1a28e251c15efb3be6ac4cfc62962bacc40c3be11751b5002af184b0a9dd595d9c1fa681adc
z55f5fecd6a8e36b05a2cba59ce069b4e7ae6a1fbe2318922f30e29626b0863754685cfc13470f7
z1eb48422d324d6be115aa69c721b5ea186368001134e71a160b903b7a43cad9470801de7b6b6e6
z77055ff6ab7fbfc4a06e6d0acd72ea8677b512be88984fde2d6d723b6472f9346b31782eef2f37
zff7b8e5bfb082021d923bed852da3df5fa34bf21a1755d5b86574864b7753d717f7af73f74ba79
z2e289b6512044803e3f0460597a32256c8b17c03228555048a9707585f2866c921a7d4eb7a5cce
zc38cfa1dac38fcb05a9e59fb74544b7d81a855b3846ef68a0a749acfef69b7c6aad593cac04e74
z61cb0e8cf6f1e72d30798895cc58e970ed2b1409648af58fc890b90f246802c74229ea0c5ae6e6
z62759911e3e723af1aacada6806857664552159ebcdca911201c61291df6da14141ec3161b038d
z5e34eb2d387c2aaddb5a81aec689c1e5a20bb30968c7c972f61d5610f7e9fc80f1955485181e2b
zda8df89a7591b25347546ebcb5c8f42a483302b61d067334c67dd9aa0fdf43b8df1c4e42c10aee
z222f72b761ee937c2cbb23029f7de26c5a72784c5d6776dc7f57521de3e8cf36d5644d34af0761
z4e3c391bbd9cc23fb18376a1cf6ea23732a67313feeef68e43a8d961e7740803e6a770c9f51e11
zb03a091ee46cd65220521051b68abfcaed2b0874ffb16e6c20c50dde4c46ced841d1968a12a19c
z9ae4b337b85c1e483284d8aa3c5285e6a68960c8884e58f86bbe7b8af1e973c70ea7df70653172
zc44dac00ef2a3ca0abe3ff46d8fc62315d0fd5151bd341be6910b93b231f645e84b20a53714a5b
z72ca916b5901fb31bceac2425512b0e5efa23d4a3bc1b2b2dfa113d146b91c29657750596a5ed9
z56907058f18bda5c6d451e63270caac864b70648b0ec17adc8eaccc7be0cc013be60ce5bb7beef
z20b9ffe9fc02685495f8a2b43ee52a398504dc2aa44eac688571ddc3900b8f1b3c9108e480188d
z6399697043fd0d6122ed29bdf1de762f2eaa3adcae0e49eec76d954d01e8dd0dd021b481410456
z7713a09704f94138a703766b9db71505a5a8d84cca91d56ffec8a3bc6db7171e8e3a3bc24bde9a
z540d05a18771230dd26372d66456286a1a38430c74ecedfabc2f7bfaa3355787bb230a0e457e59
z84220872f6a6d1239088a0334ce31146d82328c84db39251f5a6fa883fce2bca60596fbe1e16f5
z43e48c2ed71108ecee6d063a055987c8df04140f967cb6f878d489a64363630cb299cd932f5ba6
z28af6f27b607a3e4873989db1477f5e3b7968d9bc0694933d9a33a7c1909d1bc3479a6480796f6
ze2dc638d4697e9dd19fccd9fedc8a4e075640c74a5c1e13d8f7c13c89fd3331854258a15e19dc4
zaab23d1247115fd5c78e9a5330dbc218b55a644be855bb3badea4b2591fc826148c877a625a400
z6747672b00d90637513850874bab2b4e750610df0775c4bbeb9bd0d91bc9dc47d7b2d940484d4f
z1cdc273d79af5a9b38645d21b738f869dc139ff6f2b30f7a6f12add9872126aa673f67731d86cd
ze4d5782c77750555eee5bf57c24e1288e5ba235940b0601c33d8aac10c6481970e7615d040602d
ze6ab255accfc4680dfbeac66e1c1522136770b1a33fa3f8d606a37900f6aa0cd3e7919161cea38
zb8f8381abd496c8b6342fd5c6cb5ef6c2835332a0ee8c952ac29804bd3bcd087136f24c4f2baea
z1b1034a4f525ac5240fea3025f25afc6d1a424dd5305cd10d4b8198ad4a7b89d81b8a538515979
z8eab25feb71b09f759c94921ea3123f2e01e397af23dd72e579bb40960efebd7185c651706b1c8
z25bcee0d81ca10aee7b92c54dcbdd6f5a3792acf3f3c508cbd79066a1fceabb2df6f6ccc1ea973
z8fad870e7036396a9cbf4bdfd50e6b96132387c24fb65e11aa72261fffe4dbaeca1ac856cd58ee
z630ce12c16093b3df74e75cb58767afac7e303babe6682d58040520e191883a66fdb4dbd154e49
z528117af82a3238717a359ab8ee4f09c0881f19639ce489be005713df142350a6fdb95c9bdba75
zc076b8e682602caaebead3881a37dbdd77ee5ef01eae8532e7fb31cf42be3c6368ff34514c5c3f
z6a2b4946cb53119e9d06c4b6c6231cb2ec73c1331e5974d617b2b4f999995f80f756dbfd2e6c5d
z003eeab833577277dc9c21a981895524499084f634d7ac035e7930d76a9f7ff380e6d9467f17a0
z9b622fd57e291d5a5c75a71da1519563476b453f45ea7a077b2edfeb5f936a376b5787b0fdc00d
za094a3557bb69aff80087743da85fba59151286cd7d55fe41953663495116ef029cf6ede3ee0e8
ze20fa005a69ccee24a940288af38de0d1f4445b533322e175311596e95cb375f34b4a509fc4715
zb9e74807aee3a0f1dca286e3e546123c0092fba24f2d67f576eb948832e5ce2e5a22c6d3037b6c
zf19cd8121bbffd54497013d4776197fbe6398195c007fc797be7ee743c0990a75091a77705f35a
z66f8a62fdcd3f9eed1b7388925bd9bf7d212deecb5f027c289a191b25a81caf55cec45e69816d8
zf9b2968a9db2c2fad69b873d36f6c98a77845e273fec47292bcb1f217d866003ffb7fec106097b
z8ebc013c90e3155910d7d2772a9d924e40b4e10d344f169651c5d53a5e9e66092e40e914e86a73
zff1b295b0d50ac95caf0f4eddd01bf0d5c177c463f8f9fe5d21aeb64b25fa184e7b0f0d43efa9f
z3cdab7950679f32aa7c783512a01e9007005bdaf9330f2eb96520fe116775e7a78131bbc010e2d
z2fe43f3415d0df5832fa5ea937de2383816560f121b2d62af9178ccca17f7a4de682b9c458a0d2
zdf09c012f77ba6352d571ee13c3c3ea5f2f614895b1c948140339826c25eb708653a4964bc81d2
z3160a6e3e0ac32a3a9cc4e6058e68b223e7e157d2962c2535386f8547ce73087fb0aeb3c77f294
zab6f19721c16d7b9a9ab77923c4bf848ddc565a7798a5c968b4a95dd2e3eae5768de2258bb28d3
zaa78d5cf16ab1d1d69978103dd1f1c1faf012693e160043c075816fb624f47edba391f9757ba43
zcb2dd0ae0a9fadf5df2eb9e76703df5f976045bbda0a12d8072e03b31dd83f690a28fffab32569
z3d9940fb5899e2761beef2f6eccb256de6e865ea06900a84b418db26fe28d906022964bd73b6e4
zcc9894152b07b417b31f8f1a6302e5ebbaf25a0dde32b4d142060c470aa530ecab29cb2b6e6f39
zff1f5ac3811e5118e788107693fec23c73f913215f3276eac99242a6ba4131f97befe132e88533
zf0e6c05e5e328e4a351f71e349361a8c9b1356d622e93ec14eddb9e49b44d54bb33942b5df8159
zf74ea7122ffd80d619b45c799b34e7f1056183e232c5ba6d2c9eddf25e2fe7a4d00e305aef61ce
z9a22ccdde9a2e8997064c9d02d54b4b18f1d1898c5a728f52f70761101dd8a78026f6a259d035b
zea70ad09645aa65f1717202fe1fb213ee8e3f81da23333e3fe68ea37e0c4c15bf1b5d4a09fb984
zcfee1761bcf426bb0b0a3cc2347c9ce531725799ca3cb1222c312bf44b7cc9b7a20b75aab2a3bf
z0cd7f12834f597f46b586612c4de38367a2c112ef969a086a995059497468c180d0e112710b1ad
z8fff083f22a1dbb40537f574af81e8b5758119fe02867ae2bd61741907f8883e7fbc0681db6ad4
z03b4d3df9c6ab5047d0ba339e50e495bc9e1141e4f64fca04e5cd2abb6df358237d48157299e1b
z8900003f3bf3d3445397f7228c1de155182ae988329a125944783a17f7c546f652929dec62eb38
zed4e1ee6878331b78ebccf3b9a7dc3aa25d4a5a440929ed4535d2aab382d15247e7ab9373265db
zc994abae1ccae81e90a46d72ff2af3458ded0e1785a64389c7e391ea3efc076023146a22048423
z20a446a7b69ef5308a59e7fd377fa4dfd7ac317330c3f22cea0fb50ef3674e9685908623296133
zcc2f3d6d8cb55bca7ce467044c849887f7415b8b53466bd37389a41196f9be96f730e8c2b73e38
z8c50e2ccd9e1e71c0b2cbb1c768287179bafad74d33ca657b0aa5c4e9dca100847d38a566bec99
za64e6363be946ac00c6ccc3204f7f722e99cd1a5fb36bd49d64c861c9af6c32dec04bccd7cf9bf
zcba0e3cf9c44ab4763852c53c7379a8a6c40227908302861eddfdcba875a944708e3c62a8cacd4
z7d1092fb862b7d655b1b474770e982f6698edcdefbddcb801b2bc6ac0b3e6a28ad01ce21c7bc05
zb0ff5e21cbafe8ca78c83b1d8a27761c0e209f7e3ccf322b5b1687adf251996834f75f08fb9025
z587575ad9f29a79f60be242a417ea215ece674aa95262c7ad81727c0354c1f1a5e7ae75475868b
zf1b070ab98ade481deb68a7a67c26f09fb6f2434676c2b3530ae35f319d1e0313e8c4b5276be74
z6b9349111535a1d206427bfcc6694e2da85959a6e4c6f9bd039e186d0399e11e981b05112ff0fc
z58f771342aac90313d027db47c38af82fd0b4482348cd7c4c4e4654450b4b2e5fa489f638ac2bd
z19a75fac67718c94bcb2e5f3217541926870a1dcc6926eb9ddd26708f75d3d091791189dbffd17
zd954e810e6544adcce9c6cb758689a2d1bd97a0232bd58c876b408657c6623f2928a0a80729fb4
z1ca3372487697d5666d3c2d110ac842c03cec1b9d22f18cb4e92db0b875cb219aef5a92f812923
za5d2ba3529928ea00fdb5fa22afcdf2584398457745a9c5687463fdbb73ecf25843b5a5ea93aa5
z14241d83dc0d4dbdba88cd8f2f5c6b5e4a12e65f109c2a8965d1b5d60d05e9dc7f018ded33f21b
z73bd02bbfbe8fb243d4060612662b27480ea798bba0ce0b6e0a357261f8ff6028dd6372fdb38b2
za8e0b1e458e35137cb040c50a275e90d109247ff0afee1106711eb2c4076d12b4e3a957f613fdc
z04ed6aa8af5ad81055430d66f7d9c260700da14acb7192a167bb812c326ed0b65e00a358946d96
z5b04e3505bd02efef2fbcff7e6516947995a3cd52f459f40264d3e8d39ea1747ba8ea215133019
zcea4676eb1e472c3a64fa9511d405c3c8b3c2ed1c1c2bbf2e6094cdddabd810f3ed25e116e15f8
z7f7d1a7257fee854cc5f2ab5a08ae052be919043b215ecb2927eca13237684d397c2e503512ddf
z3e90ae495cf9ca6f6c3766403a64e22546602a749539df7f819f62b2e320aac210e225c2275910
zd9fcfc0328ac1a2ebae8cf2b59f2f96df2526ce3c384c8a67b659f0bf6de776a5bb8a9e06358b2
z8a7c19a5d9048c72afc39fdbdb2ea352b605a8890943d29bb18f74d1c697074a377ff8543361b3
z357a19e3e2a815df23e2390e9238e545d04e87148d2b9b0d2268cadbfeac5fd76ddf551be2ca2f
z7d9f5b984bbc5af37b73654f83811d231dffbcfde5ea3b5b7faa7467bc1a3a1094a2d6ebe0e68e
z582a1ee18dfd137d4e9fb88e8ea34770479a560c111d89219466753082ba55313e1ea969ef664c
z88c767e8907ced60b6dbe9be72043f4ebf7ac9de9b233f661ca58c0fe70ed957486a39a12f4669
z22aa1da699ad3131c58fa0d3a73a97cc0279f974bc99700109cf4cfd65a4352a7ba1c8232064d0
z05455bc64ac4671d56ee874c8e2c518f8814cd9e6ac72793aa1c49b56bba71cae325427b0afec6
ze7d8e5b8d8c1bf1aa8e6c17b8d2c0da442ef6fb7d82f8920ad6589b171a27acac203f817f4512f
z57d5f756aafe96db8fdfe2e4dbda1ccdf50d2bf7a23bcf28980a681d0de2016d6921e18bd4d523
zbf8750cb7b15c243da7d16ceb1123aa25605c97de2e21cc1e08ecd1a343c6defbe43ab26121408
z9a5554d3e32b70b82b35f8fa63c7ae0134d7b6f4462b270258c3c1bf9295c38c0dac7974b69584
z457c59854449ea2018d6be8279f9b29bc4ebf8ecce25ecac823a89724a43b179a64c80c959dd16
zfa5702c37e41767e5ab1b7a0fed9fdfd64bb8757094fb39b39b2514ada8c944095dabef2b5a1a7
z361e3b069d29f91024886304db3ddd514aa528faabb0ef590c9bf9d2415ca1fd69a0d9b25caaaa
zd917345d66ba9ddf8cc70153e5eb6957a63d4f9cf37148ee1c646efafd365db5e2e62cdfa7c375
z998327de58a5cf9e98b249e495616bc97a128578028f26eb30cfcb708802d1c6759bb8592b1443
z8a22a16e3eb46c497daefff5c123e243d4307df9965b98d14c20b33ed6cfdd72af8646cf72d769
zb9c14c027ee2c3092037bd9f6561ebe39798e78085bcc116717b8e5a82503dee648cc4ed1c6a9e
zc1391294ee37951c1651060fd88d74070e8e39461442c8de85c03432ab76510c847f417d8da9bc
z5a87d9c2f1ece6436559b55300722fbeedecb82c840f0edd4f04e071af21dde7358f736c75c8e9
za14891a0c1fce80e0df3f446fa2ccf0b04a6cdf357ff4b389c3d4713a4c43f80649d3db1fe6062
z6d7a31dfe78ddb442671058c2f070599f20d25e8c0eba70fdc76d69ae8acba4c16334115ac9f1c
z727cf769463a12d9b5c936fd48958a868c309ac8f5449f430a71ac2fdd902f4d5af2df317a3afd
z460a7ca9c91ec9dce9842b583d6ffc81329fde400f0bc74cfff51e5c8be5f6ef2c89fc5f89f22c
z294afa47de77c7eafad7165d60f9bbe80e0196fbda56b8804ef02593210b020e89e1c64b7fdd35
zc613ca005a13208c3ac79c5d2a60f3d0fb164b556733ebbc62d9d9b761313698e3df380574e00a
z8b428402efaba3b3acc74b1c8da041c24eb93717a990854774b9d75379c405342bf741e57a15ff
z4c79f5d373897e0d7ee5db6baea1d5a391094f8d4832e809561e1d31697d19ef322b055da28171
z2c6df5dc9bec3992a9d4e3e8a05054c5dc53f7d127805445e72d94c120c2537423856732377ead
zbc4e30addc2f3bb3eecd646a39ae8afd6f3e3329a1465cde046621021904aff48aaa74ecae9ce3
z52d1a07c8bde64728a35f3d69c374712107ddb6b5759a21d07e7339e3190bd4a6deb24ac29a776
z8d8099ea0d3aa244888fcd73ee3f779a4d43413df2ddbe18829e1aae89b03daa6d917eb13e1683
ze3bea0435839a489922c8f235557aed7ffe4f98a050311bac14fa2adc86c1a9df93ae573baca7c
z86542aa24c83da0f3bfcd5e736ddc7c164458f6d346bf7dd4730ec026a904e6eb9757151c675a3
zae14cd742aea06959651b98c1c4524be9de078d18721c14a89b7ae89e17ac145ee261f027a1d88
z4f29d97df4d12f174902f4e348828ae6ccd42209fba378d9d3eb0573519e3db56a6e107c891f5c
zfff30a7c2e071f98dffb58c4501ef3ab30a93385dcb921fca894c55ab0d3ce604b2c70d92b1f8f
z4f2bee883f5f016d2ce8aadd1ac2e4d6be5ec44b6a9c84c9c76f52868971d3fb916f8acb43e59d
z6e1fac1aae7b8d22b00d52d874352ebe0609e1fd2e71a42f79e6c785edf103befe2eeaefedf92f
z47c152b1a79e3dd19490cc82dfd341d6cd3a38926bbb2d24f9d78d163128bdbde68683a034c31f
z369bfc44504bfcd23b78d3120ece1fca03299133dacd08433587eeecb3c2762d1c8acb131f7908
z031ecaa5fecdf4ef81ff3f7a78b6360f7dfee282418fd91f232431f8080c09d674c1dc43b3d9e1
z7e5fcde1c7cbdc7f62df696e8b1aceaeedbd9fb4976de833c979e38f9721c9219cd48d552f7495
z4533d58c8a6851986e22a276df89189ecdf9ad23775bcaa7d93ba1f65860a9f2a2b70121283443
z1ad0401c78ea0154f05bff46b3e3c18b88e497c3a8dbdd87d0f73850be231a4a7dda10d0b48923
zd616794273fc028ad41443b5e9f37b5b525c4e775ba17196bb17ca3f8c89c84031052d4c2df964
zf1c135f969883ccde740418f9534683fb798bfcd6494a2be03ad72ab95dfd53d72b7e335fe6140
zc9e7be4f4186f8cfef489ed000050096dcff175cdb5226279b2497b63d865ae0429ce1e83c8945
z07ac51f74d95b0be6bd3e80821ab8480c2e3a6a3c453ea0160fb241f0757b4fcfaa70076325443
z01f2b6556aac5eaf4c38e53f8c03d4ed5629358ef68ed748d3802c2e604ce003c60027475992ac
z1019ddb30a5126ad981e1093e70c03b0bfce02bb66c1f479443a87a7d99b4b15e7b4caf4d176ee
z4f4b9c67140e2c21cad9900875c938d6dee389b95b47334ad2c2010714f450e9799f9f1321ad49
zc808eb9496f6a6476a55113f1f1982f0139e0360006f5c5192ad28182621ce08bcdc70ca11f3a5
zd2f6abac4e60fbe1dc3b143678a96f95895218fd9e69baf1caf8dc050da2b96faaa1c4b4581de1
z88ea38d3d1479348d8acdcf2c9b789fd5c199d724d517c252c7d712344382d8920ce68deb2bb46
z279a468fd7a000e05be8194dcf833b8825353f91f8ebe2c64f0177e7ff5875cd2c596831c53e2c
z82edc1991efde2a3516bc81eda5dd4780d74f207b26324bc6b6afdb0180d60ad8e8a34894df0f2
za86f8b536467d47a4729443b458ad82db398fde70c6351d687bf1de040fa109ab02722aee17e81
zb5107b048be371b02c2ea9548b3b1eaf29b43811756b08c7c86a428d32387c98ed180a9d2d4601
z22fd1c8175aab8926391c356873c19b5ccf4fff4add8fac751e7cc4d2d482b2973ed594cc46354
z54d32167aeb2e315b3d9ef8f2b1913c653535efeac0a91ff597f22e69c702bee851b9aa8c3e2ce
zc5600949a00c9ff881120f31ca1dba6fe66868051e6802fe8b67ec5beb5eb76059b07a29cf65e3
zca166aef03292ca76abdd955b2baea6e2f08169e630b3ff7aa5004e603147cf079e339891e51d7
z116b73a27b68a1a53dabf2caa93633fcd6df56950173b715230184cd3b63a8601880098cd5940f
zd6b7836edf25cc1f903ddab78a8a676566fb8a52a9ea8d1729817012ba2b34d4166a76408b8f29
z2904c56cf7fb46920c3ec8b61cef366529daf329495b0578979d2d8d57bafcef33c0995ba394b6
zaa9bd5eaddac6132a03c2eddd8d7e20d99f4c1ffbbf2e248de868d954fc210a4190e9ef425de1a
z769fb849f58e5243e126ac2813b88908e888332f230c18fa07bfb8d99ad629a1e1bc8f4b64f0d3
z1b82ab454d89ef2ad4588155e8ab4183eef20fc0d30ca0a45c959602d2ca5f9f311bb965b8f69c
zff286bae4f3e5c202e9a8563e576e4a132806d892c700d03c011e0d7c446efc1234d4254f6c07a
z3ba23ee53663d1a186eab4a67b28971c35a2720189fc0916902a19a0551077a80e319da4116c5d
z4e441d3eac16c2faba9a0586e746550891275f9a48e6a33bcc87147645480eb68d3585dd5a3cb7
zb47eaf7700a58f44322817413fde040e1f8588cb6cf222e6f006fbbe30717741a82dfa233cde0b
z03aaa7464ce4caee806970d767be3ffba468ba0c8129befe14d2a5d762a34ea04449e337ec178a
z5dfac3f86d3d97fe3c541c07085510e865d6a09c29500f1437491ce536966b50cb046423144497
zf3229c8e31c5bfc56e6b52d19548a020d66f785e388481e6a85f93e5935b62410bb6bca957e376
z875dd6d8338435b9b954e7b057530519075097d9a4a610c304de5f5382dbffd9f7e401d2603ab6
z0c91a3ba1e72b9a65cf580a0b0c00e12ac549af5bfa54ec186304159bda9b1ba7687c03ab7e8fd
zbbbb77c72c272bf795402904bc5ef1195dd5a4d400aa44ef205d3a46cf47b0c0102ce562e90bf2
z75fa9fdbaa197190fcca13a3428ba06cad3d793d5559890b2cd4d449327aae3f1c3f3846f59856
z28900b8c29775537457bd3a1d84b9c790f752a7313c9ce3457e48530d6aadac177c8285262fe78
z159c7f7da43c66d74d5375485b21f442455271f41533395d32a8a925d07d45e0d4dee850f255d2
z82fc55a19175191937678f4ca0d159c1569affcfc34f0b428bfeaaf7ab0073f63223dc6859386d
zeabbe852f4f52956e04a91ae37e14a1670773b24faa4b8fd67eaf325039323fd41bdddba156cf6
z21ed6b19fb154c6da0f2b1182c1fbba1fd5744e4c2955a352e31954311ae100aa28835da234962
z8a42728af26f13eea01924ca080838d112052d284f5a7e9c16364a5868224fe1612a53ee4ead78
z9723230aeab9d995939fde22b239d11b870a0c2bfc8c4d6a89cecfddec918413b60e0809d80e83
z2a40d2d61c37aba042a0689eab61ca2f34b0a85cad44c1b64473a22f966bcc2b8c0503d0992ab1
zfe04b05a09ab33ca49d9e1de633283360475339a5bddeae6858e4902c989f66965e09008254523
z7017efcbb9596666286030ff79ca00dbb198e44771886216184f1575a281d08df9c2429b1c21c7
zc8c04b9aaeea70d297456bc318c99df01816a27f4e7b6478af414406a49fe5b1cd9ed6a7082a96
z9bc5d5cd87baad427fde3e65c7d3ab62971b1016df0a7f97c9f09abb4fade76a594bac072cd78f
z8e3d33bee6dd3721eb2fd3ef2804fa1df47c8f04e806c635c1579087184f1f1614ede7febe5b3b
z79f2f78a0779ea5e2d0ea4708d1912c385224a5341d2ba82afe379935d63e091ac0d4351bc8d9a
zc56df7e43b6a27f4fb2075ff671174ea84b6d318c1b1d090f1e62d82740c19f2e049958b7afb6b
z757a16f4e7c617ce7b12acd032e3c7cc196b864b4da116d67c92b328861bfcba47a64398fd3a5a
z03d798444ea2599c431d72b0b72a44479f2459bf9aa8466bd2a262c5460945f724f0ef43dc81a8
zb525af7be3d8291868f3c72eb7e76ecd9c8f299c5a0eee646bcb6c7a8223abb37986f885030ec3
zd4f8cd125fe163bad79c61b4655ddac84114e45f8c13be27cdb3e59fa2130637251fff4ac59e73
zd549979de71b1afd8298716dbfbe4539bf52e6c64d43239db2cc10ede3eced2f3ed5dba1325b20
z97b9cfde35ab5fcd8f0754e8e457d094061c097ecc6654b49471733b7043897a2a39907adb7346
zf744b41c511b6dd89891673de89a79a15bb7ea9693b0dbabf30b19929d18f9552b4283d19aeb06
z95d3491fc74b861ba27ea11f5855bcdc3620ba8b815fa524b7fca7d8a41a0aff85d095e2ad01a1
z6fb7453c0e86605ee25c7e99dcf09ee3d1179879e5e13622fc1fe4d68e9d4fca3d6fae293ef5eb
zfc572ce33cc92d775b16f5a5f9779e7fdd8b9ce3622b0e805fe977717788b6f0f1c596d228e328
zffd1d14188668803b95fc8684030236257cac3ba7757fdcf468b0b167f4c776c6047d215524c68
z658792ced6836e0022e3a16b0698f63f03f322ceb58177d106c0721df12dfccc9eb15989269226
z70d33ffc983ae639dcdb2176200f23adeab7aa45b5cd2181edfb72b430380dc4368d4a7380a9f4
zc0c11b580c893d59200f61e3734da7b1581d0f50f37ef3f2902a938953b9ee39d713ce4f442df3
z6e0c3c27630daa8e24d385676000391ab91146565141a7c4551d7f559dfe172b5f2b5da413a78c
ze5ecbcf8c79d55b5de0fe05fc58aaeeeb4388d9539af4d2ae460a28b316431ae7c7f8b56c6965a
zf8656ecc180ee6b78c772dec194f559398adc8c6bcbcb2f0ffd4f66d890dfecd1b08bc83f08915
zd6b26726154e01769c97763a48ecbb2338c3a592819e38cef6d349533cdbe3a1b9cf314c5678af
z732ddebc5116191dbdd224fa16d61ad8b97c4701861d9cf4ba1caa708370299a1ed77c8809f381
z9270cfd40b1fe3ce6d8e5349d95e3e3ecdcce257b43b7f66a18377523e666641ad4f5659cfc8e4
zbe680fc31da5dfcd11b7bfab6d07e1d95675afb45242a13f0dbc98cc64d6551ca4826d5ea2b606
z7969bb4980c9ff167ebf2440c2cbedd601fb6e42e36017a1a7e006f8b770119bc02b1741cd8c9a
zff4dfd53dad83892ab74d0cfa982bdae404f613e9be0c7f1038a099885c03e02a79743715a6ec2
z2705d1816370c015baa494dee1ed9842745a31575297cc0f38cbdf136d0d5cfead93026480f1aa
zdea8c82696321f4bfda8c3b67278f5d0755630b78bd068a6b3d9de73251f65f1c6bbfbb7cc354c
z6ba7ddf5758f1cbe8a994bd5582325fab9c912e4ae5881cba3d16f3143eef46ca38daab86fcb55
zbfebf94a01a95f579da93bf9ff6da64d608610e8d68b28a76b45a23460f040ca9c9861d3949351
z030ef3bf7ce0c23f114f185d8d6b0d90ea533fd03bca2fde1dcae9b6e9d5c97deb03565702dcf8
z509e6671c45eb8b4e7898668ea53becebc80587325e0a22ae3ade81bd851a49dabb85de54608d9
zc5a1cf7c2aea6f3a00f2d828de5c67d7e2ed99f7c302e9887b2eae0cef48826573c8d14a12696f
z11397e09eed37cf1cad998e201ec13c14a6ef30636d06b6b6434e7d6852ac13e0be8ef1d5f8137
zd50a692c6c482631cee4649d35e061dda866ebb4545db8fb834da26737e8296e7ccf0ca7d81ecd
z0c2b44ea82d99f5c38b0b79fa426d82a50fc9edac0c155963c0cb9114cdd0a811ced3878064cb0
z704ed0eb554d145cc13e9bc2f183a8615a086aae047479a43f5197ac47b35e7ea223c58b2ea843
z6e4e1308de763f9feb1fb0e62d5c12190eae68fa02b4563a46c4d345289c585fb8f40b16199481
zbb87761d8290f01d744f7f95c581aa3f5fed8ae0a3bad6eee7937ea0c554a4f1b47b514c440263
z99059cdc45b870e9f8796a97ea04311edf7e5564fb5e5934ea3c5953a148995dc84463bfc3c621
z0a87adde27c550af730be01bf6e1f5bee1558875b3169704e0937abb9a74bcc155c0e3d28ecbb2
z62140d85af5871654918fd826dbe566f07f54079aa87e4489d208e5479b9d53abae736d479b267
z3759c738fcbd1d2911c927fb4510a5d706fff7f79cf48674b51c21354107f0b57b337302939f57
z5ddd081958626bafc311f19c374acf87ac0de7aa2cee03ebd5255945ed81d138a7bd831d333eb3
z01c9c9311926406a8917a77a357306f42736421946506ee6628c70a6e39bbbf4ab21b94527a2ff
zaa7c68144907304370060042dc192e44784eec73a54f39a5b8149049fd1d01aa7fbe36faec7ad5
zd9a3f42430b0ab4300dd020fc62d76a23e2b2567625b3a51fee3d675dadd0db2706ce8be36a260
z018e522e013ce715c429e4ba46e32c77f9b2b5b6a68c3dbee4fbd6dbd62e5b4d160bad03c520da
ze05a5ae766a81208a66b82af77198a7703c756f2a1bd2c233079ffde2a99326cc17ea3640151ca
z47efa2d0db6c3f54132b41b7fc524f76c1bd35140e16f025e5e9ea6bba4c254e2fa01f9ed9546f
z643c2e72d9789c9ca4533d676c21329017a1c24ecc30d4077b09577b6bf2d28ccd5de8334b7ee4
ze66d7f41d5ac4bae0f2330c53f8af977b2de5693e56c2086c3dadfb7785f087b2ab2b7cb31798e
z5269fa5bbb45fed0ff59594309bff6a64fa1e34b307cfa3dd351e0d47cf23b2d7f7ac1458899df
z31dd01e12e75e13f9ff3719ff8894558a6dad3f8fbef23339eb1a1cc6181e52c789cebc84b5782
z5d0f14f2824fbeef68959fb4264c3d93ec88ce5ffd944861af10a35caebe14e7505334b6ecfe91
za428deb8007658bf16c8bcd8b7e1b3e4a43dd11f4959bb60121ab1fa3e00dab362b966867e0648
zbcf66f58e9085aede480c6d212fe04f8e7fa6e32400d1321db636eda0de8cfad92e9b2e9330e16
zcd38846218b583526ec5794bc6fdbf6430ebcde24896e8d9829b826db5abeb5129926456fd0a08
z368a228d096280655e6b513fbc575139aabf3dd4729e896d07e4dfa15ce8dd915ab68a544b1ed8
z6c03fd8fa9c131c1fd611378a3e8a35866d41b22176df0aa1b2419a6eabdf6a89c654772a11ac6
zfdb135130d974f865ca3b68c42dbbfa96d4da2dbd6dd5f282cd14e3c87aaf99e492ce8f8eda0eb
z10c2bc925df581e1bc5e387ce6d66553a4d3a517707f69864ed5ab346d629f7e12f62e6bd66f2d
z5e787a44f10636efb2aa64ec738ec67d18cf5bf355e0093a78444d1bf2594b4897f68b0d5013c9
z7ccca008de27d281b480510d5107dc31f153fc42b382ddfec75dd91672ad36188c90d6e8dcc9dc
z6404a0e49600f44c7c6130e79ac0dd1d02f34f46fe3ef903669f11857c0a65584fdb7a5b9a839c
ze12fd1869f4d730f8b5ee75406bf8edef4f0cd1e3b3e52684c107f7fadd1727d16bbf5ec0d5965
z22092a183324eae660d1d77516def605d4a2c1bb84a89029a2d23ee91bbec1b4bf6647ac526d6d
z1debb2b16c8575603d72d5c2e13270c7b82dbccb485a406bd1d8719b3bab3c95b229860e7cc358
z17045a760bb34dea1751db231f951f583a8e5560b1f6030e2ae744d54ecb4ffd2e6775647ae57a
za2d81aeb57aa6444ba4223060f8670fca96f195170a24839db640efa15860740c6fdf3c2256e3d
za6ec2583c7990848e4fb33abf16fa5214ed178d7191e814339b3e7a3e02cc59f10e0c7acc46da6
zc0fc04720fbbd83287ae5b958e433271b56dbd0b7ee1fa5d5131ea3923fed013763a8caf45737d
z962bd2e22c392892d9fbfee8ca7fe061bf507b4bb06ec3617966c36f58856b6649e0ef9f466a77
zb76ec10b21c6991100557d1b8f25efdb0c9b74ab061d39c28a9bb699c637bcdb0ce1a6753a2af2
z63f789a2176d6de77fd9b68853da4ceff3fa54b688142e3d66664ecdb68109698fe4640e44c23d
zdc082e0d576a171ca8d57dd8a9839169e672b4de7d51616ea997a3f53d053879b526d8db4f899f
z1e9d059d1a96c597e5c4f76f865d3843cc8c9488eb0de8dcfa4ff25adc5989ee3cb9e9c74ad358
zc31aea2d4b5ff885c688d32307f14f2db47c020231593e96156a6ab0ba66fae7a9c73f58691698
zcc05a684bfe3a5f3fd9c6dd8466c91d6a2f73fef34f1126a7354cdb9f7b97ae48ba47695909d9c
zed45e7b7889653bd2db9f5be88626c6491a95bcc9405f3fec690980510ea2ab9fa08ae5d5cfe91
zb182f45f92e1bc2b00e645e49d74b352066c00f1a0920d4c122e26015cc97ad99ea314b812e3ec
z8311f5624dff60c4f6d5d11137759a9d7d7067c64c7f10c7ec9437cda0c41e36a40023d757cf73
z3e44ba50ecd0b13aaebc82cbebb0f276c344f4beb7ef34e1bd9339ec7ae539949497ae67e27fe4
z625a1376a68d6ff1a996c97c3ee4912da33b9d75eb35ab5db00599b095c16cd0cda76a73cc17f4
z5c93d4909a2c0da463790b614f52b42a465872fcb09a0f12905bd19102e227246a91e8da433db1
z755092a5cf87438a092d8d44ff8dd19ac0a460f6f48e5b0dbb8b2553a87670d6ada041a02aa407
z8721e3b437848b76a0cff044f5a0b8170b7c59fb1110713ce8a4b2bfe63b6d791e64e7143f3691
z1428c84101ec964eda59e5c72c44c6546e7641b73903807574ec13b052a5a91fbe8346acba1f71
z121f8ad1246c38f19d8457d76564718aadacb406059409702bca7ddb3bf473ce45cfa400232351
z6af1d46f7015a5dd355f9a2ea30a5ee52564428e5dbe9b339dea3314ae049b24cc930d77d87cdd
z0e4a55689394b1cadb02a9673e8806ce4c863a7e56c50876c6604861a3ef7cbff16ebfdd33a8d2
z2b81ce2309726d0092365fbf4c8864a0370a18ba2906544ab2a9179aee92e7082515630534a1e1
z922cd9843a84211b205ebf1c13162da44b6ca0d1c102b5109dfd8c77df1718ca5933cf2549f8ec
zdee5bc699ac2f92bd3f3eb0bceef76205bfd0ce4c07ed969159583984e19ab81422caf6689abe2
z85c9e6cfacb92314a2cc56fcb7d8a12576c73bfe1eb3995352d6bc07ccc112c1af8224b6218468
z5ed6d9b51422e10cd9d7445b0bde6c3d2c68fd6e1589eb44f77442de410439ad44003fa9c23ba1
z927efe5787a5d9945535d6058e154f0f701deb0dbbd748a54a63833599745e51970662a5d2d258
z37b639323e71049e1daa5261392157cc3974f9649bc19d6a81ba18865c807f97ef58b8916cf229
z0b243b746c48875b09baa5cec35fe46b47a9c42ecd10f0e13a5d937329f65ba51e45bca47e4fc2
zd5b93ae1ffce11b326424c2116c60d55a7176ffa1b795280952a437761359abd40624512d2b4fd
zf09415c0d767a4220e69c4648b0fef17cc5bf0bd742a77635f2599817f1055a80414af7f2e1714
z4ca4a0c943d44f43684719377d09b9ae8d71047cd5621a270a2097837e895e9298c6a49595775b
zdc796dd58739b0b22736cb8f63159ed63e8b2872409e70e86422b6ed6a0f778b700b8b7bac036a
zb6d5e98d4d524c5b00d7b80c5f4aafd457464e7932803c201d35604cce8709c99e3be827099294
za60b284e7ce49f7382fc7506580aae2b192e2be1422ad44e6e8b7a8afe2c7f816d1aaa3c5d76db
zd29f5cc14f329716088c2f519609889f34969fd3b81ac1fdcd2d69e329f5c343c17b27ab1e1417
z167fc51d5255eff4e24ca87a126ace50eaa4a9ee00c9aa793c6f4f9ca5ba812d06ddabc4c3d45e
zc46b7b64484cb4adca286d078e0d1efe4716b9097abb6f56b6c0d52853d4b276e74a3473ea543b
z4bffaa0990ae94de3f75b2bfee0997a131676e64624085394e6f5fccee1db575c51a7436a6ce56
zf38d1ccada4c92d16d94831182eb1c80fc5f71234047d5d9567e7fa77adaed6e65d7d11ff5998e
z0aba6963b207e2fbda19c703f85c87db7dd4cc74476efba3b135dc2fefb2c9e638c503bfae9883
zaeeec45ae2dd568bdede35a35d19b57e82ff4a4f0bdb38437e84d032bf3bf6f090b158adb431f4
z406287901e5a77713ce245661a59638afa0070419a4f2ccc26afc62c638aef083b0cf5207ac066
z98c2218c7958b36477b08ce4f2bb1bb2c236e97794fca6a7b9f358244304229065f408c3c4df6f
zf23eacb477ae90b0345b4e51a946f6a23e3beb669ce821caebafd2bcfe27e408ccc6025d269ca4
z314d8d500469bee429b908e7e80466a54f8d4d2d70f5e578447e80e5a6bb568116430f6c79984f
z7bfcf501254d6e313724ea9c71ee7b5c87b33a69e24c1935fe7babdaa0e22c0c822b1fb406a00c
z02dbc3983d92233b4a1ed109030ecf28532f83116f0b700e5779dfaa3cea4e5e809a6551826860
zf34452c6c5537c722145807e9c7a482a562a55ad198d43cd195f6ada4b5b86ed6d4f5f6e92229b
zdd6e85509edb4703bdbf4e0a42157051f97102ca1f45b1d747fedd5c9f960084c5f744e428fb9e
z0c967f0edf99a08e81f0e201a304acab6e94912037faaf1c7b94f3fb1e9b8d5752e9fe7669cfce
zf2b271e8f3c3d1449692dd25dbed31e9d5149a56b782da71c63c809891bde45fa64091f4f93145
z0f039ece79d75366af001eda86e280047f33601e112672c9f04a1a19187436c86042f4c11bcfcb
z4465fcac1f6735ddfd0a31c154af45cfef8296943ec52f1bc698ba3ecd0971fe12e000fb0909fa
z2d23a49c78d08b67f63b4d78c12fc31ff55e58260bfff1fd7c8dba7b05f17bdc64e5566ead790b
ze1faba4700e7e06409318381df3c8c7e9bffc80a9723915e6a5028b8ca4ff2e0b93a16cef11943
z2197664394d889a323801a978023536fccf4fa02c82778ba000b14f1068cd5404241aa722d91ae
zbbb100c06fa83b4ff06d4f5d555221eef5c4569eb47ed85165294b72f22467b0bf06b59b844145
zae3815a3e456b339de8d1bb87dec4844bb0b64b538b79848c6868b69f7c6760a6eacfac66f5206
zfb9810fd67f22c8317753326e68685f14fe5b53a908381ca276a5d2390a82a7a25da5f3528786f
z3ed31c4b2d32a138a5ac22fa7340ed00363742c60e645d00569e2611de6c839566a6a72fbafcd7
z652ca4e755334d9cfb5ef0ad5d3fcd0f701c9fd88c31372159a48a817a61aa92c19ab6b0879efd
zde1569c7c459403aab2202b24d0c817bc8f33ea125cbac762f598940481e6bf5a2cc1bc03b0714
z488739c115450281d0014613a23f96dd686f66c584dd5d8724f165747854fd52bf0df10c7aad9b
z16e9724d955b1118c7fcfd1a793056b445faab7343826ede0e11627915eb15c67bb1692fb668f3
zd6285951a223df36f313db8feb12fac7009ce97d09efe47454a0ebf6a0b13953d4a5731183c39a
z668122c32152dcff64c4930d05a8e4c9b1bc7f3aa63007f3ba19afc4baf1009b4cb2916b5fe041
z15d71def45231ff2d4b8b50326e58833bc46c205f647074ca9837c5e2e66fd88f5530b0badd8d8
z21397f4534f975e1a6b3e60b6c8067af51956866bcf4acc6b0a22fcf6fabceb16df4887561ad66
zdf8c15e8bec21786b54f5d390614f5dca439a8183a0e87578aaac97ad65b3c8b40d86bfcbe1d36
z59769c4e4ed37b4aed2ccc456ab56c425a1bf55cefbf1bfcf77a7995655e5ee1f9ddccb3086e82
z84a5759aa5436ad6913e3a2893fcabd8bd5ca67dd1ea36c988043064da6c6fa54fb29c069dcef2
z44861da6cf38ce52542ed0c67d5d0ff382c5b56946e3cc99e2bd26058416ef61f7082aeadbe4fc
zc7655b400beebc413d6018a94a80abfdc3cc75b9e0de5223c61830e21258081ad962332027ae77
z172db1ed17a16f0ba321f85a1f301a03861917ae033743659394e6847e0235b1809b756cc6a643
zd37f20af57ff2eda1dd1557e295bc4650376a7a7a7df2c98252a20d1637a75a32444949c4351b9
zb6989612158c7cd3c25526a442011a6ff06d92e5a914639a28c29947234d3774c34555ad94bd0a
z968dcffdc9312788c93b71691923abf2d3ee18bf8ab1db48dbbed9b863bc18ebec49122bbad9c7
ze2dc66f82411fa5a043f7a84df90874c8e2f55c9c9965bd97d3c2247eb881181910bae8226b3fe
z836bf79978b11c1dc3a86d331ce5a84abbd442edbff4785b0978d3613e47c33b4ce2cc42897100
z13f83e745e8991805fd7eae87067528ef3544ee4c8f0091c851809b33a9752d0181dbab928dae1
z25e42675b33b99ae8f618a6c281e01263950ee1a76884368113f98309810ff7b66bcd5c580a352
z00fdeb7fdc5e37e75aa8376556f297a46f190a5a6846ef494519a9dc105fcdaebaa3384b3ea0a0
z27bd207697d7d30eda6669a18fa7d96da7c34d721ca9c1315137d5fa899992583968bbc8de0363
zce6a6ecd2bd77a4444ca71579fee74ca6a55629850d88b837711baf2768752e930ed05520b05e2
z521d5fb66b8250de07d5e828668058b9eed2a6d6e077375a4dfb72509c1fdb03ed26cf605f0632
z9a07b31bea61b5dbd42c5af00739df4210f021a60721aca6585a10e7fe43f8550d7ff0c85f9478
z32b78b9e2f323cf5aa1685a6057233335eb020b38f1b0b1c0fd48c517bc971a887fa478416465d
za9558d24c4657e0480f00d3cce915ad459d69fa22dd2476d210b768875e06ed10e7ce6017b6bc9
zb99be9c9bc3eb61249a0ea092fcfce80068f188e77f6bd5b5b95b4185273dd0faaaf1092a1c87c
z40b80cde5115a10c6cecaefae8bf4c91d1deb3af125385939131dccf03c2eb85424a4b30c980fe
z6effecb09839787ab789f38c1b2c48cd7375b1fa058c3c9cf9fd5101ab4d460b09b34b29ef3398
zb65351b601389f81182179386a1b1d6a910f3a0bca843a7de381295269bbfbda470a596d6d8850
z259d28b950bf91ca85826f85702f3fc2a9771271489947b03c4a21494050cdd855451525376b81
z34af7aa1ed5926540d7c9ff4df31a6c164a9b865a9f493042d8851a3683395f18355bec91bcca0
zba6e05ac8725ed409d6a30b73dcc57e99cabf7bfbf2fe7f080092daa12e7f1107081dbf5389a09
z1f54933837d319ea65ea5cd52059138b38ae534fc2e138eead3f7f21f11e631101eca2918221d7
zb3297cbd974d633557971c6df4a99d603617cdb643e9231e505eadd9fab804e860bb09c24acc48
zd0c35e726145f214e68546fe63c0d52abcb297698644b9049d121d5caf7421251255616f90d4ea
zf37fb06195dbf9adcb8e4827f0b9db72b4963fee6113ea80959a89e01cce9b27ed6c65bfa6afc9
z5aa81db7ffbe8c96f4917198bdd9b323b21e200f8be1feaa438d041510aecb7d6a75663730d50a
zfa94d52d8e6265e243817469d0a96a711dda551eba8e3f332af4433b2799ddc7ca419e7f6fe1d3
zfae33d4bcba9d534e16f84a684482bc95a12ca27f22f66a1781899392b1a5031cc68ec2ef18cd9
zd99d3703e4990a624ea3a5a576f07fbf1ba6a000cbe1043ca9dafba71dd09bf358916238825d9f
z4e6ac367551276bbf458752a93e7c637526fc3a8b2ca56e9f076b25d803040d3caf27b72875714
z0f3857e00951742a05cb0a573f0bb3208deff140bedc135f52612f830fbabd24ae520bda8b280c
z9c20e630a7cb46decc40a64ce2838ff6e4360d7f18ff690cc6d81730bd91a4bfa1cd99dbd1ac0a
zb7e8e481bedef427d34d36e9c3496991e5a298457f1334b2ff160aa4b77fe8f193566a8f03df44
z599324a5886732d5542d90964b480ee926b51bb25f8aaab3463cde63178d26ccb9a26e8d8f09e5
zd2ca57b8f98cffd3a33b84bbf4c0431930622269bd547d4a783e03064b1e9fc40023cf3724bffc
z7df8427b450b877f5dccc198076b283ed62e33837f7853fe239819f1ee12a2f625b12375ade645
zdfbfa20415a6d6b628b4dbac5f160bdf9c9f5ef757c2bb2d00359391b716c3f8bf94db143c4fd9
zc709f4b6c30753169d11c885e0c01e53aebeab97f0e93d67ffa5db9d7b91958d4bfebea4f4f389
z0554f572e2a290b0e4c9a3a0811826a3ded105a6eabd19860b365e51825145d209360722a545ea
zc97992792632447546949617ee63f065e9e999762381c50a01094a84dbe873a058e0e223f2b6aa
zfdea79f1e289d7a4527b7ef367d2ecd9d2903947cd6d26182f79e503e9cf1dac388d31891ff29d
zc1b25f101cbc6584ec8de2b629cba7b54dd85131af45e7f0556f7b81403d4e92cc797048d729ab
z772e00ba57777751395a8d046b6693819186d9b242147b4b24ae0be92a08dd75200fca2b09fd6f
zbaf8feee3098f7d97e680e8317ad66016177bee61382d283a7a2f210ba1ce8e92840bde1bfeaf1
zee36101d715cf9fd2d39cc472d59824a857762152f8e95d27fe71ff32d3fe60af1211ed65c5f02
z8b7522836acd29d5541b43b0a21fcfc0f1568d48b7867a7067b93957d7d34cc27121ae8a4e92d9
z3d4ea1f5d598f3e984e06cdfa9f877e84ec8fff9a3aa61d11b8fa77421ef5eee3c2b919a2be249
z9f38505eba91f6a7e355850805a435317cffde1100d0199c091c04a9c535557707fbab860919e3
z57739684bc11896ac99560bd8aef1c64eb8e60c36e125a8a41ace61bc368f67f443f69b320e0cd
z451558759c2644735ecb9675f79936b41d153fdc73b0b5e945c11607115307ff4eb63da989d200
z7b71f05b1c12f8be8287cbcee483f9020d4526958fb07e887b3e72ec4b6a10f702b7c1ee005aba
z2a6764c09e84e67e8adb0c40b5cef24cdea0c12ca873e8b8c6c10864c34e99a84f58ffc89dd3c8
z99fed028c111882e16839142883847db6b8cefc76a4e7c5204b4b4b2432c83a808b638b2ec815f
z383e4f56718b66845ffd616206ff4a23519a8b685a8c4c26d8c156725ade2f9b47d74f1e217164
z4925930ff550591aa94fbf2ded8e64137253bc8f2cbdf588d351977264bb398b770392292d5593
z04993212debd075cbed58cc54e894cc118825176b373a51dacd20db74dde3f7c50fa2cbaa7f69d
zb4fb2a894b97be0d259c4da66b53aca2bc670167881d67e935ff79bfdb02f8bbadddf20d17ff23
zd28c15f358465abc0175d68aa8fb18fa25f0b3124d1bceb285053b065b59a6864eda861f358ab2
z45b6faaed3f51814fd46d1fcf32b048ddb3e61729aca1c04181aade84ab12f105ec1a4510afc19
zfb8766bb2dcc6420957dcb9837a36a9c64b0a1e06a758c0d21fba2965fc42a9a6c918bab1ac649
z393bbaaa1f8a3acf48294a0a0e33f3bd90d36778f1862f8e5a854291018f7492c69dd362f092b8
zf1f21184907531547cfe4dcb2863e8a20f6d172ede72c5c672a3fc1636b2c65522f62a5ca4e366
z94681c069644b6c568607cbcdeffbbea0fb6c4f84eb5cc3f8977f5131a38078f82531c125d7b5b
za848fd3051135138e741faadcfe7c4ed623f923e9a4b0066437685711f7f5aacb4d1d687264712
z9823fb63b0961131fcaa4d7abe6f4ef82bc2f1a954a09452bf64e9abcd07ca435044f602ce6b25
z097af231b6ee56183078d8699d0b7858c68378436317a68badde07c2f12884fd311ee4faa659a5
z0e0b27badee190b1097e724bd646bc50e15b43f731535c0a5d853c348299376948ed1070b8b090
z2f8c7d4ceeacb9e8818f9d3bde034d7e944834c281e09281232689ab05e773ac87effec239436e
zdfc8774d928039589c55403abd6846b51d32e929ac7d2dd5c19a9c4734ed253c42f7eab8333e8c
za58b59ecdd69ea9eabe2e9198d5ff6801f45c17d7181787091b4b1f50f372c05403adee23b2b64
z06bc01f36d656cde8ffa9c2be7ea8bfc78d2fb11c294cda7b0f7f515c88286d0a3e7cf6a963ed3
zffd277954836141cc92c15bf954f6b013e04437b8b4c8f57bd6feea5819303b0bbd3f22e201b53
z1a6929567772222bbb542cda73f7053df2fe860863e3671d6afab4cb39b4e86412de7f8928c93f
z70208ef0dd25677e2b0163901fa25d4c4d15828fe1e5b935bac2917d05394096f4fda9c4b18c3b
z50cceb0ded70661051e64e05b1fde75d0a771a6a50f6ac9f2cacc535f7bc0a0fef35dab808b93f
z9d51491a2cb8caa7f094054e88097be9b49c816fa87f9df5491b82b9931c519f2125f8e47e8aff
z5b4ba36488a285e6a9eb17cd90a641aab51ea17fe90c59207f6d938527576485e7769539e13450
z052312523c49822e5a61627d4bd4c55b4437481944f3e88d0cd5cb630fb6558f085a40ab4a57f7
z8f7fe7bcac6b4fa6b38c9e8307e2115eb8a647480351fbe8f8b91f58ca5086f69b3c1e192f62d8
z6d65ac1dfdbbb6b58dc3b950b55deeff35a154fa3a34a1406704f04f0dbd1cef6db10c56dbf5dc
za820b018a3135667c91799a8c7106c299ec4e088676a2fc0c930815a1b4354e4bc8846b5f3b45e
za72f47854d0f5578bf1785339264a21bde6c4dfd3cb43c2baf932dd113fba6d81f207a516c91b0
zfc66cbb84374829690e5d4bcd000390b2102fe295b8d67f644f82bb8291235ffb70d9d47cec8cf
zf8e611609b1800d723751c2b3b8677d666f3571190a40fc42d493a46d6033c61c1a6caf3a83712
zbb6d7828686882605a72f7945a48b3691191bc7673f8b6a5d2f4a0c6075b78547ec938363a60f2
z38cf9b39a20eaadf8e7fe94079531a3202ef4a08581707f1c66cbe9cb659e55bd766d1676f05a5
zaf0d08d2c11390aba23431f69152ababcbec39112ed86747a1f1bcce025d74f5c87688d683cdf6
z782f127fedaae32339b2f66146e45791a0f7e3e2ec76ccaf0eb66bf6090914f8ab7425c95646a0
z7d5e0c8fbb5c295f78bb2915a9918828d550563ff17c6cbceec1293fe50da90bd809d6a8d91095
z0c15b0fa87e7365d5e60364e733d8b4fab4234b65c173f70035d67a75c26c3ed3b03dc3c6efe8e
zf05c5f85e5d1b3e64cd27ebaf80793e0c5e13416a56d8c091d36d733ae71d37cab2f20d824f215
zf68d2377f23529b0bddd38c265fda3591d2832183fa85659d7134668d4a919cd6aa775b5980a0c
za0ddc6f61382f8ef57c7e86803c1e076d92446fd37aea7b3ac51409a4b3db5b4d54bc4f0b92186
zab649438fc2be3ade7a821fede1c255a12b084118d0b3432b7c3d5352e03a2b8a4cf6efacbc286
ze1eb20202194d310b42e1b3cfefdaf10da28ab471d1188f8b4d962a7849d3663219974b0a0b4ab
z04de42ed995e99d17110f36dc6b022751a500094820fc32110a1d4c0157a17f6787ac51ded400d
z9d5f072f9144fc214761aee6d77d564beacd24c04cf28a45ef98574dfee428080dd3483d6dc4ed
zba620839862c3d5f1c83d07dfe958da956b709ed8242411a264e0880a8add6a573672e7fb21a75
zdfd0388196d4a6b58481559f64965bdc1332e34b025bc823699d903a941de0c2612118f4b08ba0
z34381901fe2e8b1c4de3549be2dfef1b2d2d385a9a4e25da7af3deee422288d80ecf5d91e55f67
z2c7eb03eeeb7058fc352be5c03c878628848312ba0b3a654bcfc4075f35ff770d283578ff1b8c5
z2bd000dab93ff7465be00df1809a6accff1a721697368c77e8511d6ee5dab59c174ca15fc9ed5d
z9aabeba3fa273546952aaefe30007933253bcfdb1dedcc15a349f6d4eb293d9bdca8f4238a7e22
zf805cd1b914f72b6bbdc800fbe643b9dc05e61e0eed7f22baf1236701de31553e26c6d4bd2c70e
zc284ee18d39bb448a4d7dfe21d26280fe9cab80fdb52ff8f0b1763236cd2a011f76607d89a170d
z910993c2215740297f39a069e2a3ab36852e451c0c18bec40e1d93d074ba212404ca822db641fc
z6764231334ac7bf53b2ae63f62d75f4a2cf0e593a2bc62915a1c9a6b2bad6bb5d28f66a76d9785
z9ebc5e5705358eb34d96674e422c160b3eb5418cc7cb9cc74f12e0202abb6b88c8e43b3bbe2848
zdc29294b3ea8e230c0d0f173e5dd615e5e52b8167a315c762188a21d3ca0f61d880a3437da59ab
za77b7011a5b61a2bc0f770b3e1d18f32fe66c75d4aa006d9afe47ecc737cb129135b6ea74fa68f
z52f14af7613ca53c29de310cbe82c8e69ab8958b55188cd07bc26f77f4173f3fbbe32b09df3e66
z22eee58c47785a70fed3dc7efc0763372f752acd61c4cf5c78828499ae37e09966f29653461fc0
zef61c4c0c6201461ddf0c367b1f3242eb9f4f14a082031b6af8e173a4124bca9bb24d1445af0f8
z0d4d7a5b569486757c97d8980af10957d52ef7d0f4ea19d918e4931150b95db33ef932ea4a2b84
z3244a9cc673aaeab4a4626a33425ccca0d3406d38001605500539032519c5fd37f41fa5e352c6b
za3fc283aab0c8f687e71c5c3c1d8e1864cc7f4f39b745dc0fdaaac8f630ca7d5d4dfe044fd2d3c
z871b354ed221b09b74a13805d05737ddcaff7ef58700cf42dc2e7c25c5d2eb366d80aaac637575
ze70087450e760e093a4e92c5f1e4a9ef3dff475cecc6bc13fae80625d22d9c7eb1b005552fb6c8
zacfd6dfc7e9786f5ae8354a00399d60f78f6d7e7fb69c80b6dcd750812c0bac410c377e18eb292
z24053e3561ba3f77f7f32ac7873cb88132219b73b616e62652deaf4c6d62a38beff505f8a51389
z4fadc9b1bbe9fce721804c89f5e2721331093ee9935815c93666c8f4aa6f51a0f44738325b6d8c
z97e6daa3391528828283b8adcccdecfce60c7dba44990fdfcc026eb1af1cb007028f187adc1c59
zc360a27886fd7867e8219371509c368e0b944dd8a09278e8df7e97f7faed92fe4681182b46187e
z7a65d42c9d1c2352732fb7935682831e3bea0db88343f1b6fa411830c88f388cc6a37411c5d338
za819f1e789492a60f5ab15d433c65032ca2bfb70934edb124f09961af6f25d2758ac4b49dea0b8
zd0fab7fcf442ec478238506fe0bcd49f5b52a2e0cf916e11b282fce9347ebd6342be6a58f3e4ff
z4cdcda0ee6b62c76504452f033256e92ce0a2c1bae6ee6e721e9784dc47e088316c424e553a202
z60026801e5f14eec0e39b204d01ed67b992a5396ea74769a53d765717ca66a3d37dcbbfe98c58c
z01b4cbb0d5b607001f544c7d29c3f1eb13723ab861a8225898888f413e84cdf96a9c4395f071cb
zb5fcced35ef3c60f1dda54b4528a08e3873e2f91d655616548e9ac676ec85df1e93c6273dd26d7
zd3a52662e2627744c72b75887549a54ed5e72dc8d5c0a28ee37890b282fbabf1d2e96a37a19a5e
zc37b1bc341ee9aefe2e780ddda6b7878639d7c259c72c2c368104432a8292ff731197756084948
z58b5e8d560dd84e0d82943dab4c6489f7f199c9bd69f08538c562a86ab07c9717482060101f12d
ze2599c769e3b27fead757b03f0183b0729982a38fc1e532d4a015571505c845cef19c061300c3c
zf034578e2c505768d056e1a6a5f58bc93552098687bae6214beb2dbbc038723418bbdbfd8fa748
z3012de5d374b70315f848171e6c64bd90ac4d3f2ea13817371a9fc61f2793c85cc70e0d48dde62
z81822ccd9b670e70707472b9b6de8ae9d133411be57b56f4e3417c981581bdbf194e2fdb185d7d
za5c2bd83fd7ba83a293ce636a84aeaa3ffa846a184af51f3b352c124a503ad78a7aec3535e510b
zd53fd6079e04e89a2bd39a6dcce3e7367d356fb7d0afe31fdcc87bc4310cb9eb4e215387cf8b9a
z4d447970efaf7795e8eab1fb54df8daecdfa7cd68d5ee251574debc6676057d0fac45521a1e15a
z4962d272b7c34a46e7b148a021a4beadb842a3cccf5f29b79389cf86c33f8c75975d1c718129b4
z9aa0e3aaec9e1c6ca9c91c6daf8f0bd3d00ce119dbaea5730446082f5fbfadd7243f92ec719e56
z47192ed14ba21db2c7068c37d80bbd5e493bac93b52224aa75ca0aa8e7c2b59a385885fc34c0e8
z16f996324da2641b6fa098b58be39b723cd60f3b318fc2166faea1d0babf649d2a331d6bb73e1b
zf756c417da34ecdd8b0e4694dd3c201685a436b8ce424f3b9ceed1484d846e2f87af9fd5b8a436
ze9c11608d3fc03b70386f9720cc0b8f55a23f6f696021d44dc074bd2ff1995e5a8827cf85aa92e
z4299d01a12f3b4758dc8eeff05a6f687e2acc96e3aa87dbb3bd98d8e650460eb1d494787ae6852
zed73c3a41fadaffef53c4e3999f48b565ba71ab2fcf462d3a9263a2722988aaaa194df934c83b3
z1cea4b46c3466c56e319bb7074fd2472854f47dbfd8f925d4ae89eb417f273158e64edd503d0a9
zb4a08502409d530832c3d77b82920ce133f0320623b0f873d4849816cf6e6ea77f298566a7aae6
zb49731c51e7d22d600af84252e9f4d49fc52b00b819a50e17fe128217c026f073eb0d03f30b11c
z5e6362de08040934e7570274a0320a5079ccae4fcfb8bb80a77e8d2d4cbccac175fca0c47fe892
z50aa8cb42504ef4d6056bc565e561cd40579ceb604a36eaaae242372c4bb3e7c91714019915cac
zcf344503bd16f9af06b369cd5d44a324595e7441a3aa005ac7ea6e4f8e0241f9a0fc3f60dd139f
z9ddfc110608ffc3a74d783a35a1f92f20f64535d698c56a42ced698c673b48a9e01629343ac22e
z06c04510111692615449baeec11ff7b7914d4a8bf51673f2ea201b3c84399b92efc5587b7f30d9
z6139bc76dd94ecdf63263bf83067cb162136721730da1ceb535e1649781cc498cda490e5e1b348
za1aa15f24bc77f76032551921db742f15b8eca149c471cda4d26b1a6a9e5f31410855f7f0fc087
z0c90f8c6f9054ce6ba33824974563da99ec259e064a5c033ca0da5879c0b30f47b3e471fdc493d
z185aec5734b659ca69b0d2bd1ab29987e0cdd18130631b326151c7ed1d1249bdc725eb414ae3ea
z49ece923c83383a7829913952bf513bf451283304abb8b7fec73027ac2f3e7725031f043dfcb0f
za740e9b4066952c931ced06803dc1fa9a01e3bff57e8f0d5d5ce0fe58477d3c463adc5c3267378
zf06bf71376bf7bc5e036ca2385719f8a728737f555d27a5638d3c08aa772eed5335a2cd0362dd3
zf8c1503e84c293c7765b2f98edf483c8c7ba2fc4b3008c5820bb18eef9eccb6df4bee3cc47a248
z315e4d51c56983c110aa0c4539eb1cc24749069ff8d276624e8346733ece74a563cbcf35071568
z5f8997c8b5c1c2b506ea352c2d279384c00516f92b22366a0bb229673cccbae5cbc66f6144f29e
z0397b5e0f910d960d63e96489304ab88e8d1fce73457ae2f246accd2e0653e6455cc5c7256dfcb
z74f5a265ad25a0bbc7b6efff84103c2b036db8a3f3a28a8f1a0d3c92e1a24638cc05dd5cad5925
zc798863c7e399b5f5fcf8fba4f1025b804cb7eb0ea7a82c76bf185123933eddc4f81dc531d0a00
zef320d5f6e25c7f627374fc1d1936c9e682b034117f7f2932cb4430a58c8314814a17bb9ee68ab
z13340f7a1c72d6cafb870cb701bc51cffd3b285756ffdff0764b19c9346d9123f1d054fa5c789b
z6e2c30f3939eafdbfeeaf1b51f20a794e2395138900ebe6906b8832dd3224f78e3c29656f0e2b9
z0835cd6444e0fb98cfc0c127fb5fdc72c6fc361c5431e73546e742bcb3925be9738e7325f3b792
z98e07bfced66d43b026e7c2b1b5f9dd03db588c22ffcfa30a453cc2cc4b425511e692598604c33
za167a7cf0b09a09f247593ea66a294055f6a86e85531f06d83f3c62cb0bdcc7f64a1446dd2f7d7
z2e36e564d75679a4cf7c0cf11f4cf91a0dec35b4e13fa3a129c16caa556efe6bd2202b23419707
zdc8b82fdaa5601df8bd0a5ea3dc86ad39c45b5dea3afc295bc1ac078f2c7d82cbd28ccde97c2b6
z6a274f2caac9b2b0fc91967b61fb0c27a6551dcc96c55b6c3db3714948a587ba844fa478981a28
z9b5f21e90bba4f6e557473de8415b99eeebdf1ee3242bc9d3fd7a48372bc818f994fd9cebeee07
zb964a36645d4f11300ce0f1bc244042f393572f912a99e6a1c3b427b47dca7f11b707090ee00b6
z2f8d7dc86eff5a4174534ab5fce3ebccac02e592c67cace328e2ace4ecacb066ab754375b30798
z391135afbbdb6844c4614f83a0894fda12e7fcb816f28a9c352c955019cbc4d45d148a2d460b44
z87b79dbc3481d7c73905863f6a9c35fb9693a7af9707bb9da61a1470d448a724e0ed28f08fd080
z7440b962da2ef405f2d58fd6f1a0e44dbc017e91d5c202e9a2ad95800c1013fb375bcf123c3d49
zd99d5e3233c97aaca08dbaa5fecbee2fd38eb2de4b4a7f4568c1b7ab0391b3732697701ab40aca
z0cfcdf54530e0d73264109ceb7dc74cc13e4390f04fddebd60ebaee82764e265764999f23ce0a5
z201303adc421d7c22aa55817f685abc1d91ec62a28577df50295bd066ecb3f846358cbd389094e
z85f138ff83c1651f7a87c4a0578c5c8fb1841da95d43e612fccf4d17b1a3ab3d95c7f7dc9d5531
za02c141953edae6582b5852cd18226887885746d391e9c4b64211961909d6b36c9edf4b4966e09
z9bfcb21cd846220c865584ff9cd15d6b2c065f6f5f2f6f1f37de552a52061e152d4d770d1d83c9
zb31a4c6864ae5269b2760c371e9255aef8935af490e05892551e9beb88c5cbcd8c65463a0e7f2c
zcec26263fe792217b5b4a034b8e341406fd075391b2e7daa1dae9c5161264f1106b4fd338697b4
zff8b8b2dc1cd21adb651cdb6d9bd5ac56e866643a0dfd0c34c0a2ac52fc401757b76e7c9495159
z1ffba713ce14af47f453170752e6270b19b635da8228a9893dc785293d4215f22f84ddf80c1689
z658826d08ac8ec13af0c115eca67c454f9461d07192e776a619d6798df447d333817a7ad15e9a9
z37d8d2c60b05aab187c6a681c9f3df133accb3f7d7e0ee2a3bc70780adedc7f9233c1d643c5acf
z34085ddf0c2f1650da70a8a8c2d66d30a5f8f30baccaa6883f27fba83ae2fa57d3fa80ac2728e3
z539357b1f524cd405d427811d53ffbfe11903e755fb8108441907786545608355dd19a972b64bd
z22825d5f98d6c79f93692e0a18cd403ca9baaa58987c6f65e2cee7eb57cbf3f0bbef8bfb24cbdb
z35746a17516956e96cab56a710ac3a316d3d923865229f98422d7d2b1e4213294dcbdd5f234c79
z6717f6eaff51d55d5e7fd43b76a75b7b9e910a5161f86725670173619e6165a96385ab06a40d23
zee7067b48ce4c10c458a4d4742e1196a93db01a658b6185eccd6aac4211a3714d90378c97cfbec
z6678352be3f84486aaa49256f9ca5c5baf54b8e9daacc9decfb130be944caa7922d80ba39b81d3
z98ac918510f6585941b7943f589c147de1ea08c48a3b5fc44196bb1632f51cd73c60b49c01b5f2
ze1a5f7cae20d4ed8339b2c51423a8866639b5b5ff2630b51d41e521a476647aa2bc05d7b5f8eb2
z7ad417c7c9354875bf27430400cb2323bee016fbfcf8f143e9ef1e0986096f33b556b5ae48c0b8
z5fcade641e1de292ed411c4d90f8a28c123fea0f4502bb217988b60355806d92b9d44250cfe8d2
z51e9d44a79d07c51d2e2a08d27acfbcbd83d25f7e2078651a3b7002ca19f4d6d8027d6bb824691
z4c728c89065e29003a1031c0be4b54167a56ac87fff9775782a4520a81c9ba216ac3a5635e0474
z4b8ac66d909665800cb25029371cf067b0f9c18c7ec2e62727247fa444ded3f2f958b7eb8de636
z7083f4ef5fe78aca198134cb938ed1bfa5daeccfd9f9d243d2dd00ccd5bd75b91e5e9b3729b67f
z3fd8a5ba9ccfc0318bb5376b82ce4c52b7be6b5ae2f3c9589d87074549130642788fc07487bacf
z515091bb4131cb16a8237d26c744bf30d30860f3434bf51d1fd0f578856d2ed0a94d08ea3349b4
z03a2c97a656dbbe13081d5ca41c94d29b7beb4916e5ec45c6d671ea7dccc0aca731780eba06b47
z81f771b3c612cdc0e7a5262d0238c20805eee0876b9cbd009423374ec68205199be4b21f163b12
zdcd540ddcafd7e3a7882e5a3b95e4ebe6be76aa15274a5eb44a13489e733a49fd47bb9fa03d66c
z97c9e90851d01495d8f3fa9d105c121c685460963baa932f501880dfa5eb12e353b65a0ee84802
z3c9f65402f679f504c137d42737f1dae031bf946fe0c9deab41a9118a14e9fae06ed7dff518b42
z9e88834cea6661644e5aacc2fdb772f546cd8bfba675327d74c7201162e28abd3dc634c03bf54b
z0f2844e800cdd4954c4a62560795732e727d4e52a25f36a160316fcdd66407d926fa841189acfe
z6df4f80c8803dc701abab1a4e27030bb1075397ff21e0c97a40f82a25e004a6b28f48ad6a03f7d
zffe58ff797ad9dfc2ec4579962f7461af377f64a9c5999873a2d13c7d6089dd487d00b3eace02e
z564acca970a77923430a246e7ea6fb99b75a729a9e7a16cb116e732f58b1b83680d6c65475f774
z6fd4384265e9695f0b0837c0a7c62548f9bece2bb4769a5b56ddf98d30152c20a7f4103349f774
z6387e2b98bd28b21da174569a00a9de1a87bae041e767f452c5d1c9c35b43aaddd4ae64786b8dc
za3f298ae0e0f8d507004490802ed010d3679f53075ed6da6ef0e773dca5d5e53fee3161a1a3b83
z29b17371c5164fdb01310666c6cf0562c2011a473bb03faebc63d1591e911edecb55283570aeb9
zc682e25d06d9e79d7c6e6d295e92a6be7f230952b110c8825f84067b6c381131657c01be7ed3c5
zd32169c5dd128f6103f51e5c8ecba95efcfc16696ceeb34d5d9335af10e659f0d50b2a2be1b030
z7af2417fb35a8480d6ead58307f45b44f95a2a077233dd4f5c7057184105755dad8e622ed384f8
zdd2e998f6ac5f5b04f4a6d90753d9229c7a4c2ef1795ca8888d1acfc2536f5755b41a1d272836e
zb277907b0596ba1342612d21b5dc57c433b7de8e97b011abe10196ed748de919fae4eb64e38658
z8ea54e96276919524bb82a046e1be7df831a03e6a52dd37c0dc9163f635cbc6e436f9b5f3af6d5
z09b2a8e5aff4c3d93d5a688714956bd88e758bce801c6490cfe3df567887587b032c9ab184186e
z16cdc37124dca50e5d41b2fee9e0db4f226143ebe2b649457e178fd7e011e5cb170cf95f0e7bad
z62ae01608175e9391365d702ac79362d372532337b027ed8bbf54de691ed43d0e7255acfff18a8
z528a16244ac021e3896680a3bf1dadd5581012db3c78c012042e3fd6fe65c7b885e3d3d48bfae6
zb64cd07f5e2a5f616bb033d6ad027c5f7250a7d3793b354def3f9c570b9e0615c6c3a90728802e
z8585458303e5a387c32b089ccda337c9db3b3b529207db6ddce5b769396059e4b786ec7ec29b36
z718de5a8ecc44f2a0987f39cd6f4db7d6173997a259fee574580a66ef4a69e15f62ecdfc8bc857
zd0321a51d0be2107bf1b9669495745317a0c0e593c919dbc6875ad258b4c82b10dd9678ec00242
z4d02dc8fc2aedc5286919fd01a8a1acc69711fcf36a7fe2c7aa5d980404447264429036788eb89
ze0d197005ba86af6d177e40730843f658c722ca78457941e42665f22f93435c7e3fe73657df3b6
z74a8512683ea9eec7e6af8f794510debaabcdd9de109cf1d05fc88d46722b08f05c9355eb69473
ze3166d4653ac239a24723ad77ac13c0374b3a05d316750f5858d84a04a6660ad9c9cd5b85497be
zaac50860befdc9f762db499b8eb73d2fff9e32526fe80bd551dfb01807804648dc75b813544275
z611e322f81b8f91ac8be0e277593251f6eeec5b1c4a4beb88f19a7ac9b40f6f1a290e77c97727f
zdbce1f1fdc383ab8e3be5d8eb91c2210f1cd914747fa2a4f8ffe08f3c205dfc2b2580268b89776
z66fb97c404a38f33a34c6804ea05574d0f35604dc1839ca9d6ed311fa8dc48d723978a29e1ee49
z13e17f4c1f97936142d0b43520a9b8acb3490e19478655bb33e1083545b77a4baedf91469a91ce
z470e4fd15fea2659fc01c66f9bf5be4e42fb7387e3c9d563541107a5fe8153bf99869e8d758cfa
ze378d86224151b58f199fe8e68545b2d04b5fb7fb1188a7f1f13692b758bf0ad1456a14ee7c63f
zc87201f3092dbe6d881185aa353c16bed6ca72d95ec8266969350c6f6ea7c87c71777ccde44399
z0e1504d7f81ff47875d3fd043bf91bf1dbe44608d0d8b4a268cbd4fba119e7d33392328d39edf2
zc478a08f0bd7b1ddb7f3ac5e9eac745be0ab49c14088a5916cafe432db1bdbff96139c86f93d0f
z55622952d306f473ffb4a15ac605cb73d6e0a93df97d127a6b59e45abb778af04d1fc443aacf07
z40a2a6f00a80f350784f7344fcb3ee522b544de82d40cc2ca3c08bf37852653adf8f3e8b145da1
z464a85d1e1d87261f3ba6d3b4ba9a2dcbd90461a3f7d95887293bb468e1d1aea2c051d43df1c2b
z822762c522cc441df597223356178f4a2a6701805b61f85837f72f5d56f21311facac6a06f7aa8
z9a0be45931868c83814978cfdf73a23f7cd986255cf4043e65884fa8eaa3760422dfdb6759574b
zcecac9522818ebfd8098b5da721f3d519c8d99f2db4c08d86b7acbce518c0d8c7f428fa33d2aa0
zd78d05d9875ff1b79436072e5ba5e88da7c90f388f4b1d7b77aa659fbc09f88010546c08007afd
z5127a89c7c82b5ed50ea57cf9921f358a235767459356105821f7d6784211104be51ad9590b507
z11ea4b8f7dcd53c187ad07fc1b37729b44926363f3316baceff85e1f8a6c6e49f652923b09c6cf
zbae13adf74be03fd988a88cca49826da8606b5a764fb6be379a9ac35434aae84b657bdfe49bf4f
z85c370e182caa94a110e314e5b52394337996705d42de99cd641ba4caa66ca26b02ea15fe62a9e
z83be74557e1b7f8387d6afab315d745c71ef0d7b671383b7d9dd62761fd468a20684f713037b06
z97d9c8afc879a577d1545150327fc1634ee99bc5d07e611de2e7b0240d74e3ec0beef5b4cb39c8
z0bad35d0265fc308533cfbfa998d5ba21394639816d0f44258be947525aa324104ad4f7d37ce86
zb1fd332fed9870894c31252ef77bfe753466e92ad308f3fd82408836834bd3528bda8400cfab81
zca4c81f9d64d22d3933f9d472ee4b0aab11638e15c96473d7d8e9344840d8c13a9a977636dcf4e
za0cdf267767ac6232222dd4b8ea42f58457e42038cf5d198e375594b8b8410fba32fab01cd1a8c
z76ac71aa0291cb96b4bc43d2d277d4a3f48a7c7b36c5e62e06f317351f284ddbe58a4eae73c83f
zb420126ad1c89454729e5fb53b6bac41b90b1d55741628e44fc9b3fb1685454f1d0d2c4437688a
z491f1d6ee72a3b79c321eeefdaa680486e493e1b5ecce13a76135156fa66024d3e9b641c01ee86
zf8100053bdcc6b1d610b56bb5c1130c3839dac1522872cfc746bf62baf9f475a62b3662d22c8fd
z6d770dfd654869eda206a1c3c5f11c0ce8fd1d728a883660a3b09ea7e151ed93aecf936141d487
z25e2fb772df8bddd92706dfcca3e535a65eb19007c174ca9fd6b47849f9a85733c803057909f03
z1994daccd6cd913285f69337fae92da9648903251387c8c35251a2aa105d96c2025cbd29adef12
zf9eecfc7fa947063c87a180e368807e2abe8e0ae49f59df0154ed45ea94bd790328867898a2ece
zdafe918eed3c4e53d5d25d9a7593daf488c2c4b9d2abba12105e97af67dcb9c800e13ae0cd109d
z99e8496120edc76072d170477b8f98de1417c1d1998ae20d340389aa21e359d31f27c8951b8d4e
zebe53a23fcadeab0188be6344694a349e771a0ff9cc3189a13cb09d76ae8047233114f70295fe1
z3a923095845b44af6ca25a85ba48cff33989acc98c38b6b4de7c91b7c69d21e12245888e3d1472
z1d55fb7f8d3ad1875bdd139909d92fba66c8385689298ee1de8db4f311fd057eea11e98ec0f37f
z249faf20f1d97d839c8fe155a5956c0b53c1ca6187d6270d68638fba3edeb975ebab42dcaa4d43
z02e1ee33c81c938eba77ea8239829a2ccd1420ffdf1d3f40286413c29bb278e5436f112e0a0c5f
z961f7da728fab3107ffbe6fc237ade1c8887afe2e762cfa33bc993c770224a53cc869905bfc627
z94153748b97704d33658cae00f6029aa0e96967657d84e0e15d1e742a4fff5942726b943014f27
za3906c8f4bdd61c65486fb32743e1027ea372572a5083d338a0382e0f48021755612063bd39fe4
z78c04ed85c501e8c3f80ffc2b270b37b8149e9e4ebe431902438d0ba1f709ffc9f4b9c62556832
z66893104f2fb3b04a40e07b9b63beb119741f43967a6eb6e1d9d3df0bdd90c38e090ef257b8a19
zee937d552bda2a1e68983249b275be13b4872700352d5b04f8bdec27670f29caf82c423e4ab15c
z6641e2f40ded8109f99373dbcb57d92d1036838a5825a483f589edf0e9809f2787fe0559bd7aa6
z95795597c6b9e817ad2db2eda1ea8340a8c0df88d18b6d169d457748e0199c43fb1a49ade58277
z1a3ceddb483dbab021187bcb8b7e3082f1965fdf9c4eb4ae9c3d0494c4f51f4a27e7bedb3456c0
zf388daca645c5c0a029a097b8fa9cbfe5b03db4f2b240c307e6e4ee7d6a4c718d11f9dc4011132
zf8c1c1d0fb7d3d4e329b5d2b4f46a4de7e23447a35da2982b026ac127a3d42d97babafab528977
zba5fe17dff9813b57f2405c67ddf288e0a457a3cb5e042212531553963406833ad9546850185b0
zf3eda982248b8a920eab6b9530197eb83fd6f10d11d0e893a74b73a4609c22e220ffc32e671637
zd33c9cc8bb29b6956477367be4a85e7aded0eb2958f09e76bed6c0bc3c886629d86bfb023b2432
zeab4f82cb333993c287658d956eee9315bb35064a4df0ef9f145962bb8c028d15d029717cba99c
z7221bca351c6be8bac758fa1c029acfa7e37000fbf870c4527b556fce77786c9cb32ca9805841f
zf9eb9f9c429df34c09079e3c2e3a49ab29c964a0b6e009f3f521ed568339da22099e19b944b032
z1cabda3268b938dca390795c08d54ecc1a12a700ec746186eaf46e34594d09ba03d1c57451bcc6
z1fa0a010d46ae23f48c430b4baefbf95ac13062bc1d418e0e111fe22d340323f5ccae1f3d894a1
zf27904ecfe6b5f6327dedbcc2e09caad85ceeff4e60af45703918cfca40d7f891a57027650f903
zb829df20cae87d370d618a4710dea15be15fd1067e49d6ece339b2fe543b16078ac6c315e1c779
z924d60f7479ad15358e8bbaf899ed17d94354ab961ad38431ae33c17969530c7e58d7e884dd4c0
z5df1796a803a0b7efcdbf752f5454fc67b45a9f1824353485c878962e676b8bacba91700c4af8a
z9d4fc30f1214b1831e85292c81564ca14545df2557783a0dd7ed1f4314db4d5aa970f08902d8d4
zbc6bd8fd0a7b637d941d8698cf851c6e0daa39823ab3197f59ac8f77ffce445ac37f76b03dafdd
z9ca978af56cdcc869cae5b4d558d5f8828874320767ed1c489cce4257f19a22f53499717331de2
z794e7c85e7f431abaf125ea524b8dddb54e3ab0eda15d8ba21381acbb2039173d3c607ae06b230
zafe84f57369eceb5072228f1f3a2faaebe34646b8b47da403a7540090798bef06e3784605fd478
z4ba6fb699511bd393ab3a3cbde0e07b722c95ed999c4bc5c475c17998d2474751ea19cd4e7ef74
z1d3007f590a17a7ecfb468bb91374f86c1bd4355be9dccbffebb6491a8428df0b1ed15575d185b
zf484dbc327225f1493739162c0356f9d06b5453f882738f806a32f3e162a3dadd9e9e07f262890
zefadf202aae187b6f66bc7bc5a2407d65167afa17f6372f100e47762fa7bc68f929bd80381a354
z26186cefa2183fbec807801b30424a19d2bc09dfc24243f4c33450e6a08cbacd81efefd8fa160e
z43e1931723e83ff09392a4416c784e248c683efed975889dc17f544760520b61d687be4260782f
z2f56da00bb34a8811934514cd4d0112d2b6006ebdb7bf3b8572b87b93a0a09e4d1ca530e1a91a7
z679448067fcdd249f081f5ef22ee9537e957495f3ac28f8e016b208a71b9ecb03a69947e797a4f
z7b859613331ef80da1748d33872b011b8f8c5748d3b3ac8faf9ce56514542c7b8d26e2905eed46
ze73c02bc10756d4759d1400876dc0916b921fc88af395f22c8ff9a8bb24b772393b626f70ab08d
z73e4dc520277be089bfec90a736cc6f84f55782902f4c1452b68e6b2e400979a07732850bf4686
zdaa6c7433d138c415cc163266c02d66cd4181c224b7f560151d40c4c6a315df567eb44c1a666ad
zdc084a0d27f5df274bf2a65cc487f36e5bea25a2bf31b3ab36dabb258f7542a4883ebd0ff58b46
z5f4d52377bbb3d6257d737755b9c14f461697f88faed090a5c01910c68105b0642d8b20bc57f17
z54c7818527c19644dbc0949042f37b3976e4b33cfc875e13075e733c3afb02384b236307c02e3c
zbd653c12670f76e357dd3c58dca04b8771b39b6f001859adfa12318b266de70957e0abe7974404
z1b6872886aa92b00826872bb1db35b3220e6f7f4e63231e4f59a5b2ba68a4eeb1add276c66d175
z589b676fe24f42daafe3e518b98db8248f8cf3108bf6d7dc8aeae6f7cb95e8991b85f2ad9c097c
z6a43cb8c838c1bc0c8dc401ba161dd7354900883ebab6ef82019d5962e30a0242071b78d558d4c
z9b3581ede7dbd8519c97bf11d5c63e01704ac629ab120b9d0c31f4774dd142cef827cb75fe9e2f
zcc38ef3072031d3e2dd0c6c079310bf5aa7b59d19c1f006077515559c1c7478d0fd8cccc54d6c1
zcbe8d12c8c9ec9b68095dcdf616b68ad811d394c372ff86732968c3ab32c5ef58cf622432579f8
zf827dec0c3d9f78c13ddefda9c15bc25dfc7237f5085a35e0ce5a8e13b2b83142d9c8c3baf2124
z192faaeb1b71cef6eb05cafdd67659b6fd452dbb6667882548487fb7e41330791792f09ebc6ed6
z6bcdfbccf2d2f10aa53699caf87da5c0e32e91d89314b07dfb2e65de3ea0030945136a93395dfd
z77c3d88d8c3d94ac2dae26bb18900c21799ffcd6ad70564cf6073be61d182cf55d2b45873d609a
z63aafa25138a2c78352baf6e020bba567f78c705b9b2d8009d5218b41c178697482589280294f9
z00e2aefe9c63e0673bc5dbe033b6f18084d1805a9b2e5892cfa5f59e2c1abef9ee4fc7a4e69af1
zda9aa7e68f21ce4076f027ecb703101a08dce678232a02c13dffe42395e3daf86b8e2202144dce
z480023fff23cba46ae2201f0383213ceb5d17921ca00c117c415c9624c7a7964af3065e2f601f1
z7d8479be32c9e31863b19cee137c96dad75f67f86dda81cf6266c0f76e91419ba38d3cf307b66e
z111c59e14185e1888f19a27397a81bcc6959ee5e8c4d4169819d851166fe2b75117ff9762df87e
ze13c762503462af50c2190c023509d23f94e91a2caafebadc47552cd24d4167fef01cb0a292f9e
z54744c609a245de98182cb307e527c335d38366cfe1b02ccdd86b4a2a3a28d3afe13d4df156f68
z24bfaf263486bfef90493338df1eeb5e80e9844c631aa29a24f30ddbd190b95338aac513a1f523
zcbc0e20f93372b696fa62eecf0b327328a7a693ff6332c99b4cee083c0ea39c8a9a954e965a828
zaa056ba5c861a2c31a913bc78125900e200f1e2ad6a88b76add907667f928116a240cff08974aa
z1ba353b001abfae823826de28bd6bb9b94d2a7995a4936d0ce1218c8888ff0ed4a7c39f964ca1b
z789cb875e57768970237f2b5412a626024d31c68657d904c0d5adb45d1d93b44511848ce8cbbe4
zcc452029f676a3058bb827dae88e866bf43d35e60b106bb02cb7922b4f5462d89d124e6280c7fd
z57dd20487322312fa2938ac7be96bab97a36d0d6c71a29e638f369951e7fa3f519aaf2650d7b34
zae0d94f057dc309be86589b50a4401341428addb885e9de21b0d1c37913b5871e839ddf93bd920
z0aefe35afaef00210aa206d42d1e6b91dadb752e23230d2247e4ff1846c3b078fc886119aedefd
z97e1f5f8824c72198411d6aacc62fcf42dbfc6b10208606c7f96f30d95d27021f50683c3e0a16f
z2d8710de4bc90e47a51f0f721b452239ecc99d792ef0cecdbbbfcadc619dbfbd509200ccbb8a84
z9e8b249e1ee87530a3f5f41679431efa53849469ffbb128f744f4e82b31b08ee7d2b342eb88db4
z7ebc4573ad2e50baeee37a9f566a32c4fc0fc4fa21c2616f712ceda8093e7e7315065e1a6653d3
z055ae97d91f6ed2e476d2406d4b0a0ab67d3b0352adcf67873d7853b8e001937037698cd08ff8e
z9f89d1e6847728b9ac2972d9a82f20774a83e8c1d389b77f3ec0881015d5eadb06d6be45197f17
z73eb873217879b9b75aa457013c8c304ec00c05efe695e7fea76267d5c6f44730be24fbb932470
zdc54ee7decd6da4b166781f0260ac16e84191ac609ffbbdb58f8515cd31ce6e9335cc4711d17cb
z39bc75da1a0407abcbf220c3049e10742610af0ae03f3f95fdc1546028366f28850d7ed446e3be
z0a8182f6bf5dc9af27a8dc342094ed37473893a9f862fd729f33542ef8d2e5ef6a234d93990396
z2b2811752f4f183d4790a8e8bd4c618d32e2c21747056d4f8195ffd5269603205f8df1e0e1d407
zeb7244e9ba156d34157626efb41eec9738fb9c8959bb742341a24493acdb30c2999a97d62abf88
z166d2b6b370f0e05a7c240b9f533a1fcac00815ae6c20cf6c424e750ed5ad96173ab8e6a499a9b
z2d789203148f82c64d58a04be054480951f4108b72c73c34f5094d67ce5ccbdc6201b568616619
z813232e15d209465c96cab0bae2156f079137c967e9302285b1952e571e5b02bc1129f12a3daf2
ze5c453d16b2a56b5a8cd7f2b5912500bca40f463b9fce274b90fb4a4e1442d2462d2502cc62472
z341847875dd85f10737a0efbd201846e7f56bc34ffa018d69bdfb0cfeea92ed6f2389113c5caed
zc70703336c70804a8a4f2b432bd887af5873f63238b9d638d0eb7a8515f32bc721d6a041fc6b3d
z01cd78866dfd7e06b03c0dd68f669295c69ff54f29f7b7825b2439df6a0cb47e9464ca62f8ad6d
z7a7ba22f83af939abb18a1f42dbb3557e384dc5a19789ad37f31455adec141f6cc8994165f7f18
z9ab15a89fc17c03962c79830f4defe3471d7d0f3e3eb2af406d02c498323b072a424356be5f6fc
zf2054938f2baac8e806cfbe805577357dd03c9aab4cacf8c29434611ee7b6c708b3388ab76c5b5
z872dafeb195c5a634c3fbf48538db876ded16554ce8a430396436e7121e074f54bf0dc2e1a3224
zb3adf7d93d4f34f1fa7cb22ccd661d88038ab0045321c1f99a41fbbee53cc73c4c435b49f13d71
z42bcc8612b1a693189066b928692b3022189a6203c1d028754ba8e2e19292e75929d7200500513
z6ea8a7a1c3d072e3c4185a5eaf9930b6daee369521225297de5b5b585d9d030d0cdfedc62925f6
za2ec96963600686b4b37e014cc529f82e0a4c98d8533607538e73c6deb7ed9d94aa1f05b4955cd
z7a5d7a8802eba544a09086137fce08f65b516ebfe281776bb5ddfd1e12e71459ae9aec201f1d48
zc3d731a2708ba127bc43fde47ea86d33c31a2546d9789b4a5485996f951481044e0a6de1b2f8ce
zb72aeacbd7a1746de6fc651537beac0e20c93cbc786636f7607eba3d631dbc7f1c1cf5a6966511
z02a69607f989b7222ce0a49cf72f387e796656a8d735ca1e02c43c0a4028d5c96ad0e02697ffb2
za01737f9103f2eef160a7758892d23a9e3d5f074239579f96a093b098e3c968d114a0f83846c69
z88f6451131ac7965c6b22a5a915a134e628f5f7421da880b8045a42d1ce218638fa17a0fd56f62
z7c9c152d8451fb6d4eb67e7fae5f31d91c2d9f3ad668e30a8358edc53a8c5dae4fca18cfd3cb20
zd94dfd970f60ea2e9a72d37f119c5911cd3a56acbdf81b9b57180c7f59926cf6ed4ef439f6c89e
z768dd65d4f9b15516a621724856cd771832324b12a3faf66a8a022903648baedbad1803b5489af
z396e39fc869201c1e2c75b63bd29d027024e7cc98b634ecae87dafc334d1155e2e302471c4bf8b
zac0ef126caae19289e6b83d9053cd64132e8207679b9de16917d215b78873e5586a4758915807c
ze15008d786919270ffae54b529170328c887fcefbf7e7b5dd7bdce9494bd232936c0d153fb1c3d
z076ae151a03c16ad88c399c950fd65890930781371118144c47199a465a179d1f1c601a1a0a2a4
z8daf1fedc800e7f7e27377cd9f271c35f09662b10d88ba07989876b3e5323846415c3a71c3af34
z3785c4e418b346fe7955fa35e9e53b90a578bafa046636561da08d21d185a745fd59bbfbdc1e5d
z3e18b37270ef6e3e3e1477d2d9cd8260b685b1f11dd7c4734cc23a6fa96ae92d3e7cb14f2b7435
z0b342e449edc4dc3836caf42ba08c18f8e4aaca88df27876aecf6695b18f825b453eda35cc183f
zc1ebbabf96407cdd4ac068282199159f99d96a3a6d228605864368ea8288b7f10111c63bcb1589
zc3e98ca7b89ce0dde35861a25dacab0c67cb4d818a5ae87ec0baca596ccfae1cf60fdc62093d92
zc7920f382abb0db8868153e655f166573053436651020cd01da6304553bfb16d783487c6860a43
zd7fd1fb595973cee73424a9b804f8dcadc4c13bf461036fd81a913096437c40cc0ee8249a8ceb7
z6d062eb40dd206f8bfe2ef90269664fd35fec3c5fc697c84630c25996de85b2b876e1a1b3138da
z658907ed4c08ca8a37278353c2ae5829d0840c578c3b5c584168cbbf6658fc48b84c787918bc49
za5a6b47de7d14eaae1633790995d3554c32c2e708181bffdb085a4beacc030ba2b0a62d4322ff9
z71e6bb164897ce8b27e8c53d835df894a8702ca028e31ed40305383d6381fd00e37ed576dbe0af
z50490f183c22d8d033a4408a1e8b4bbf863969fb99d650faaa9412ceb2d001dca536054194115d
zed0bc471db8959fe1a0d30539d083fc25d184ce0ab99f1c4f0b3d6121153095da1d4fa7f834546
z71003b3027f8575b464b6edd95b284706fe1e478505b5259fc733913150c8cc68d8ebe0331bffe
ze1628d997d3ce454c3bf905d5923a5046cf0b752d935c021ffb133f1ba7066118b36ca950c373d
z2363791564bf1bebb49ed31248d9401c6ecf33bf1dce5be76fcc53e379b5cf335788ed7e70f7d5
zb573900eee859d9fe9b9bcad70a85c74b3ea3e59ab3f9b0b26af5b110913883a45acb07e1cc988
z38a4691985f19ca2e7999ac72d973a145ae627f876b175f42df0e2057ad3820b88933d8b76e0fe
zb75b060000ea7abf4adf386403b2a88831bbbca3a35ae995f969bd91713f5d373dcd772bd87f17
z3f0509c299473cf17acdd5747e7efaad49eaafeb6fbacc20212e4bdc2348069a6fcb163a359fcf
zb201f35746684c519a94edd96229c49e7c8bd928299d1a37fa22536fbd59d13a87303c9ab99cdd
z279385fa460c8d4651489e7f0a9af117a710241303a9dc27f4a334ef864afc2d7257cdf4da5b1d
zf435587c8b0cb183321cf9cd8bf0ac15649d271c43aba7af67222b24d97ef7e26181c9926d55af
z14fb6b27652beb094aea574725a28b8369a7c6569f29b803bb0a344c38ea39be8a814d533f87be
zda883821b6c0fac762fa4517935471cf2b33a7de2b4c1c93900323971e9304dec4f7ae2f7c2476
zb3fbd2483cee938e8b7fabe7a21467d8e7709dfc8cbe6aab0c9c101b6bcc4cf275abeb5c672aad
z8022349a81a65e3f14f6cac675929f0f075c311f7801df99d0b1c0dbc3bed17b0176b9b7dff72a
z8d8cac7c481641732b0e46ab501e1fbdeb654097592fc0855f4eacb8eefb23b71f68f82f6446b5
z09c4f60a5f8c1d8cf211be98771978962e3a801112eb9ddbbbd1e7e432859476ef9aacdc178e1d
z3d86a662c765001fccb72a56c7dc8d0559958b1c8e865d3581325b61623bdf6831e69e272bd5a9
zc4c3df1f18a21d625a84ee587cc95a2f71fa0a1308a754498f035fc32289271fa9b04870cf8d57
z5cc51571e1e0586fee0d980fbad76e6cd420bda6f97c53bd787133ab15fce1d55bd1e78efd6293
z911f17137bb74b845296bd7811c4b591368ceb8fd58bb6067815b9e881c315d3744e34fd35ffcb
zfd2439319c2cd00cfc9295f9a738a1f6707eb36bb8f86978d3b1e79dfd291b612835d8f2e3dd1d
z45a2e6da46ea82b49206903e652c8879e186f09610dbd88429f03cfd9e50c3152acd13e6b599f7
z0195cc13db0456f09a08624b59371df5befbfe63adf9c0aa038d5a4eda0ed51b7cc0bd8b28cb86
zc9f47bd1e9dcc4a6310431669145886d4b1f0e00e88fab57e7a02be5dd2b13e536d3ce577d5c66
z9ae2c0484cce9cf53986f684d171ff21d710d95aef21f908132e5d7f3d5a01fbf9111a515b734f
z8a9c86eb63d67036195458162791ddcba5038054517fb6b5fbc77fb09df602ff11c52d00cf30db
z116604942de170aec11353efcce840a2f2d684300ac460039554741519c5dd28f548fea45daddf
z577181cbfbe73cd0c287a5a20834a8ef36fcea710667b580809bd99e692fb43f84da1b96e9375c
za3d4225463b4b6e16f828db9c11055869e4256c05f3fd3e994c81c5376f6da8476d94474458579
z2b177b82315706cd64a88270cba1d090163d6d6cc51c32b58733acfa124fca97d5d27ddba72136
z0b28b9a313f8d3ce536bf41e3f8b0ea8a32158c06e5168132fa4442739088e1c96c2c4f4dfc19c
za72a204d141cd7ea6347e3dd79b4fe7db4519721d877beb0142e26b200fab523df866b30129e29
z332b5efd26766b181cfeb33b291005ce0e9a41b2fe33ccb1f1b33498aa671fa88ed1c8d42b75d4
z801c46a46ea4d38fc87bfe3710ef70d4f950ac9269834592c19760441633fe0fd32f4b09f57eaa
z3f2c15135680eb28443dd66285afe0e994f6e661e9e11629799fb3d3868819da79e0f77f2c1678
z96e2125255021feedafc73c4923a78013f25299445ec3f3fd140b819c9106979ec53da6949dc22
z9c6675d2569ad9f53d146320fd8a594d82fe938c60beaccc774e46dbf2aa90426df097031e66ef
z9444580bbe0927da26090c3783a1d8723e4a61c488ea26500eacb59a3e0157c42146aa773131e7
z09c29475a4068e2c6d4523baa61948d29fa5651d5c205fd7e59aff90dc43c9b86ecd04d6932bfa
z9e7051f9bcf0e064efa4cf9db119ce67f58cb8461873ea14af0f737e0bb65c1e932523af6e4d1a
z366e4ae607791df0b8f819008541aba91cce0e48550f03691d8a63dc853aad38d0fbab34165de9
z7a3d1f459a8d36b5c2594c2fc816efd1dc551d3040a17df9a2b1135c7879238de99ec3a1fc99f9
ze6308a3db80ac329f586226ba95baa48c8fcd389b1fba4238fb55eb5021db7c06fa125e0444a8f
z7971b6ad6646167c5cced9646927bca7d3c46f0f86fada9bf7c1a05ed0ab5d2338cbe7ed815ef3
zc94e30ad9bb94ceb3e04906a7dd588ab1211c4f6b817c208aee49ae82cf76b2c3f6faa6a49d34e
z9072fa83d8287c8e6d6fa4bdf35bf7a09d7ad1a9f79dd2ad5955a6adff298ba3b233e66f3597e2
z168652002db18426923d32d44fee397cc8d5b53002a2b5aa793420de36168ac6d83aa299b68d92
z2d4998f78bebcc38a0344953057dcf7aff9f6011a1550fc4a251764cd2e34529957f152688cf38
z6f970da6709c892496843829e1aafc80284511396f77379eb5969e43016530103c9dc2ca8760ab
zd63bfea05e985b92e7ea95879bffd0970aa5808258232fbc12a5dc6d1cb53e78f49ca3275b2801
zdc6afd6f1120b6bccb71721a4506dae7f92c5bafac495331f524da75f18b0d9d15671ec986de8d
zd56d83b40beead205adf5b66f16d3c18a778259bb8a566c08fd07d5c7db5388c9968d1303e8028
z670c4b44f44529a783135ab8065559869ac2a601e7e257569da949271a5d7bb4b082f6b1766754
ze10ab19e941abcfd67811f9956cc9a3febd710262353530d2fb012a7ff20e3e53aadd254c4579d
zcb1d587f5cffc7b23bb62f0a0049b9651123a518f2e36c2f1090c0ba54af0f5dfa898002438649
z75619eae6a6e813b06752d9123610a78afcad45b5b1e527dc825b9d4dc9279c856a207202fd233
zef15e1d13036e057622bb3983af98d6355d6cb1e0c46d725a78d567dbed493a7cb404095b666e6
zbe59a5f085b3c3138f540bb7e5b87f75f36029e1c8a6c0c7d5a03a2ee253a0196ef7405648286b
zd8486c997f90c696a2386cc8072eb095232140cdf5290ed9d7081f95207d50d3dc8e475cde8ca4
zbf82585c2af4a19bcddb0d0715a9e89071bdb8f33821e60580fc2a860265c7607b1c4d6bc1b7d7
z3a142e8afc7e71eecca2b2f38b8c77b5c6d1b55c31f7b8dcdbdba3b4ddb9199af02c68655a549b
za05676af1136b453ae96ec56fcab605c9ba021cf86a664433517efe7fc7148b9d926896f0abb9f
z974b37bc5c7107848ce5963332d068a99ae51a1ad4676ae892c60607ce5eecef76cde58e23fbd6
z12877d36d150e74b1611d94200dac66cd7f1bf2d7fa5cca723050a2197514d9d1ad1cdc9665025
zc14925b6d82f6dc5c10452b3d03231f96830a9ce32992ffda6d8b2a691b963c91da5562a5c8b5c
z6056f3647b3196f95b0aa4ca9d512351fc24d405fc9ddc4057f53661cae50fd2ea262b80523d20
z662b3a7d7d1d4ae9181c479fc3c1d79a6394cc0ab7c0eb6fb0a416dd507bf31c4003db99b99c9f
ze1a81005f2c49baf6e679239bff33b6f484b7f7c35d3df184636bf99a646ebf7b8ce5515935492
ze04ced61318652f62d59d5bcaff2c7d7f819efa69541bdffc5e9df3056b2446668907c6293d8dc
zaf34d219512b492bd6e37e4167e16ed31c811d6d2246ba86ee8c648b1523733353e1a8d787134c
z0a95e8556665e4609cd2d75ba0a3674c9e380e49e5003871f9e7dfd926e921c8b24c6ef14b7219
zc6534a109c0e20a1691373fbf7edcc17b478bcf94dc601138fbd3cd9edf13138f46df9c4ef3f97
z8224ea6bf153e9100daa8e32e1b5d850564bf8746486f503f11fbaf996ef4233405ed54e548c10
zb93662ab12bd6ac710eea139f241915ba0a7f8e883a43e96f903745a459646c34808873efed4b6
z0fe958e53119611c19e92ae9742adeaa3911682b5c5b229cd2e75af88aa56529b363d56db9f091
zf250b6bb17852d501221c2cb5f8b94d979c6540cce57d66b5bf151e590150a03b2124784f80207
zc9353817b3e67af81345c0970ad5f9e1026c2393bc43c34943732de1a8095777894e5f72dedf72
zbc172ba10aa08e15dbf0a5d16edf3e72bb75c5b01f8a86b3598360455f57511fb597aa1e51624b
z4507dcb8d1cec2953e40bead6e333f7ec73012ae358e3faed25166fe401865e1cee7ef520dc549
zbd0315aacafcb104cc43479268b4756fa2863f4ce7ee42119415636c7e2fc7eebf013648af03d6
z0f5ae2dbddadad6d89dd7e32bfd9cf57dd6a8a98bc421c0d0c5fdac5f95282c318d26482897beb
z386343a789b2f8f307696b01d37bb5ed1e617299c627df9bffb2663a603dd796abfa225a97b0fb
zed7bfa10f2f92707a222fd8de3a0b4934017beb128ccfc82f99baad29f85a9278094c4141e5797
z7e61afd436b1757be894c1e31339c55883ce8768518d038a7c29635e16480c4582d3aa100bd0cf
z2ee29dc7e0ba16320760cda70298236cfaf1c9fc3bac2d29be1a34337581143551e63d776327b2
z56751f5694e8ab953148c158ae268d71118078a3e12a87516372c34132548140d45b2a8496d48d
z8576edd8f27459f7395e38dd8cceb00577dc4f36d2987671f3c73199a5bb53e08f40bbd60b9075
z4b15c80d1729c10b67116ce9e7cdf1b4ae0bc437bbeb86df609310db5ed1aabb40616c4e2b2b29
z84a35da2fc15870166c33ae1115d9dcdd72be83213e6e2b17a2e0d6d28240576991d8773b1785e
z6191012d45d0a3627eddd13e81b782f3d6c881546ee5e771e123e316df7f0e57e2ee52c3bcf908
za78b448494c289dc45df7a3a7aea0eba480e17f7e2f075920283a727f89889e6d2fa5e48aafbac
zf461773edcd7573692b07cc3722b0ddf7d5ea86016b21dd203cb58ea007a65fe8ee4d889079702
zd3bed46d211d65eab7fbd6e47896b24017331a5bc829ff47f49066267c9edc9d20f0d0d927f08a
z5f2005cb78d440b9d85c26437b21524f1963ccb7a55e2df1a84baf2471497a38acebc58a938ca1
zb5412174793e9e13c066624ee961b8079b94f900a8a812dee9d5115e3297a445edefc5b4af40ec
z79bab854cafa06474bfcff13198285d0d4c31db2d77d6d3f8b366a29a9f0da61d74f1e168bde26
z4cbd471278d3a4e12b6b9b0039afcb99591306b53d748a5f18778dd75b0e305923f8ab5d84a3cf
z564e058ba808f552033c68b262a95aaf2c07b14bd708938c452432716cd45eacacff75380562bf
z5783358a10b8cbcfa16defd2cf76b4347ede217741887899039db24f003900aa14e09afd219f37
z2edb47a37348ef2b3e265d6031ad53debff22ddc0f78883114c067eea696f855aa37b02a6bb024
zdc186592a8417e1a0d56361ee445c287e65401f2d490ba24cf1cc683d7a8b3d6936b4a26fbf998
zb65cf1ff33b1d59ad1b86169924d1895bda1582a12699fb942daaf32fdc8241344a7abe58284da
z9649b7cfcfe3b74069e0814cb5413c27df3a5c1d3eb9af7f57a74765b56d787b07673f3cc28a13
z9d67d8a06dc66c6dd1d5578ab69c727c73a131f32234c9e865a1d018364e43caef7648e0227f67
z94e3a09f5b865316e1e2a3412e36b5de4464a88870f9dffb9c17c11eff248ab50556f16c45bbe4
z2612031c91aee25a8b3475bf40d4461b5e99e4898db82310078dc6ffd4fdf063fed6693bc0d2c6
z5c8ee722ca1a5759ea99bef27f2e6fdd4c9f9804961a3d80aa65741d691f15e155919c2d8f9e3c
z34fa60e82e32a7923f8ca60a2b9ecaedd9b6e334524a910fe0ccb1270f43ff10a5b3b0ab34bcee
z4cae6c659d6b0bbb2e5dd78daf39c196c621babf5a10fa84a8a91e19cee79904a6e2b1db787ae6
zf8a293aa74c26a419262129f96f2f96d240a5c856eedfcae20f832c7dadee1d954aec9673b83f5
z2f436c73dac6d16e351788b65ca0cb472f4127e51e924119f4c96539a007944ea8cc93b39e20b2
za0af74b1ea822bba00210489dd3fde3e2f63e8e64ad33bd193d53962f8580d71a7d77ad233a7eb
z7038b2a31b448dc44eedcbac9a1f677dbc32f585bc5477ce3a538351b33d0635c5d640c4ad1989
z3dbeebc939f3096febe2f642314b5ee0d8db651bd80fba2d45e51c2a3b23363d716aba0d9a271f
z762e613932a57dbe5686284c7da86dcd8ba6ccfa7fb71cedbf61c0d269ada439d1ba5ca2a1d2c5
zcc899862bdb9bd28c2f502420b5838c6a57447a794eec77696b0bebf4d6055e6b848793e8f1a19
zb8a279d37cd6b8090340b2d039d5ebd17729bc147ebad87540743be841cb2a4282ce5486e1ef9b
z2b4c8ecfa04f7b5621e209c9af1a0b495bb24b3d38a34f5f2a47e4908225debf37145f1c61d671
zc6495f9b5b0f26efcca23daac6c902744c1855ad746f3935784664dc997f2b237f9936db863a39
za66be4fd1489880d584746a14d0d6d094df7533ee819f7bf5671a4b14d9ef3c36709139d2b03c2
zd513e7b5edb808bcbb382f6232c347371a8247665eb397046ed1102b6ff2fe2019bdebdd298305
z6b1a7fa15c1d7d4e93df86275c5a96c2f968b632fad0fed9265e12c8c24e8370f86cc74290cc43
z246e6d7da1c118feb760ff88c304ca886f3d2f49b078d80e829f07d752da61371c90b1c469da56
zbeaf9e526af63fd77f26ffd97597bb58f845b9ce6bc5a7e8c75df3d55c3f021cd7fc8be966a0ad
zc62ee3522224cc08be99a3585a72bb8c29a49322f6d3336a95d606ca96f4a438b48fdc40f3b809
za622d5c84101b68a3cb6abb7742d7cd705ef36ec5576dbddc159f5b8cf75f516e516706b1581c6
zcd94d245d7b32b91c5b407ca94647d9e6d2b6c3d1a148ac57782798e30d7f85cb103e1258ee652
z8f1dd482846baf6a0e46bc7d26adcdb53ee77b9a1300ae2d2544ce0049b8ebd99b751565fc079c
z1621d1c29a1df882efabbd6136ac2c3424a95c58833d3991b278f04b26c712a43e113e44bb8853
z3efe841038710969539fa1bb76da4a5ca812daee15278881eeb563f9e0195ce5b16599b566aaa9
z980deaa1a8374e5b9180f95363461ccb2a434ebfe9d90149de74ea1b4c14420c52c780aee699c6
z1648419a0b2cdde35bd02f80dff55924e1bae64c8ee45436757c534a2565b9f9fd3cc78897058e
z4baae841f76c25438ce47944dfbe6f77fd8027e11aded9c2525d9b7f0300a32877c07a48e6eaad
z3012adb9edbaf8b1c0d6c304eeb780c781eb5ac482c4b99e39249987bef8847fcfcbea63fa07b0
z2f64c9004774484338bf25ad98f9b9322409c51042b3ba266ed527b3a99c115300b7ead3f8e051
zbc523ae58696c52955df685191694fc5d3e070fdc5e2d0945008944f1ebf239bbeecaabd2851ac
z89021f60eebdb9f6e3b3fae482db61ba1ebf9b7c975ed4cd95a207c833913c63939ad49146b5dd
zfb4fcff102492cbd95362ed543fada928ce598964b3620899aa48343ecf3c1851a998ba2086fce
ze9c854de7f01b4355c81818123589b5e63b6490bef9a4eb8a648fa3213785f78bbaa4ca380af68
z333e7556f99f6017915ee56017e6107fa2e00c9f7f9568201622cd2beee5bb7e2e1b8413075b63
z5505dc766bc89079ae8d2e2e714cd47bc69a15f491372840bd5939312882560bcb4e620dc93864
zb9a7b3ff5037a0dfcfb22fb6701f9dda995acbe750bdd5b6727adeb04c3eb5967a99d50f2c571b
z6bfcd911107610dc8edb8026bf099cd3423635dd4e25522bbdbe643341334a301591ba5e848dd4
z9a8a1b851bd97e972e2b86ed684a1da32963688a215451c18c7f6d442fefbc0dbebe4832cb5bf7
z16152f0ebd60db60a505bd2ec662e9e0554e3da72ebda10f0da3f6e5de8c0ac53404a20eb21aab
z5e5959ebc4b601817ccf5eeede9f0db3ae4b9c208f8f48672ecee34e894e8d3ac3ce3ea07b62ca
z307dba715672ae9192ec76b9602ac1105c033bf283fe5bafcb061d2b8102b93cf532b7b24892b3
z5fa6d2900412d4135852612c1b03677f075d44cf746333abd096ed85eb58c473855460495ac7f2
zd87cd517bbb6e98f1bc6f72790e8748c1d86bbf770a5b5a8f9c881f0f5eb6815fcf3ada851460f
z09ecb06cecad6790a6447ef27f8805918677b611db97e317ba01c6e5239d088e740dda78216765
ze08fb27ca2a5452c5857d262b12c80f4e3b82a47c3d81fadacc2d5f65297ead1b8c1f91377f1ce
z00452ddf23bbeeeed252a38190d7090ed5c83000d2fa8ee50b5d7195eea1f028fedc2a988f6294
z6d1aa0a9840c7ee1eb1cf715ce0468700d7216f65b9517037075289449e126f151b58292c8bad4
z8c957a8273d5ef0df6da7469f770e490b90fbd6d0d88ebc84233d55f3d6a83d61a4b3844ec17f3
z16c69386f8dd051c6a139eab18f396c5465d7bffd34062c015e72397416499cd591ad1e2d3e434
z0a68971d1b546daafc9fc616cfac5061c8aa8ef583833b5b9b499097bd27fb4665de7c9cb93f9d
z0116e406452412fa9df20359f7645bd230d8b9f0bc98e0b04232914d1b1771db970e8d81345ecb
z2d69a11f0f758b9e76a900c28befd4fc50a07719e2b8c9c8b71938c99cd94e824764abd4818298
z8cbfb525e5eeb47eae94051e8fcb1a5916eba744304b5d3c78c5655fa117730f7ff969d1f6f73e
z1c9ca953d6291c03736415a248bf31baa0a807200b4be727567aee4f7d18876a4c403ac40fe3d4
zcfc637c7cea7cfbfabd55c03826c4fa1335f9dd1d94cc22ee19f2e56b61a86257d52614f8e74e1
za6d921252ce21f536fe78b5e5e6507492b6d5f5e3d5f01b6b56659cc06c0ebe685f5a01c5acabf
z3a650cec6d99f7d8d39b138bcb5f61287d942f4c69460e0be2a16bcf9863afe5e325e0f17d9d68
ze1bf0230474a0224cbac82fd3b911b9351ff79304a31ff0b3bb3de08b9689d1f963f0e460bd123
zf1c984e2b87bad3158dad828b0ee4aec8eed233add4ffcf061e589d694cdfa477d313009dc6e92
za8de92b78ee17b5e9149360bed17aaa49dd6826cd278f0e65bb7bf8b1688368f442e7c871273a6
z79419277800ada6a3727da5a0c38126dea16e691b071f87b50b2b576a55204a10a3dd7ec085438
z8dffcc5081fca4ed50d9f6ca3e7d2a5d502ac4bd29d1f89d503ec236d260c1f7fca8fdd40544fb
zaf765762c60aeff88da9470dff44156321805544bf1210e38a74a89775385b5ad1686778d46fc1
zc741c2e0eb49ea0b31de7038407c8624a58776b89605ae18164322cc0520dab2bfe69aae6e0abe
z8a4a3b84d6b26a1224d13b2ea702e4e9c344f5f1aa6977b6da46c4bccbb08bb0b1938f9bd44951
z5967dfafa7baed742de349b04f75a59bc9b4344f5715f34ef020b22d303cfa4cdea30d310ab026
z8b98c0bd37dc53eddb2a19702a55312b2dc65f5cdffbc49f15d9caa58b99d6238850c911966a1c
zdde67da7fdcd0169b7740a93d4ebd1f05d8e0cbeb46c5c885fe7287fb5c0b3925e638fb1ebfe51
z455c276f1ffbe6c661da62856f089376adad85c491f29f52b344f9dcc911eb52550ba5c1371307
z9f18714636d1b31202c3dca65aceb192a2a2834fdc76a57edae2b4896ad98447b69944a58895ee
z94766eaa9528b551f5ba11232883acb3996f3c9cdcc2fc8e600fe6e0652b75cb13db0ffb96829d
z7ed52cb99818b08e8de563be3b406bad2bb4a23ffdf1a5e11ba78a69f11a87724be0c4ebcf9bf2
zbd91d6a2cabe74973a59fe39c89b11c3e8ff4e21f09fa3bad7c29bb7ffa6cdafaff6574826dda8
z23eee4097937a63085cd4ec0db407fb2e3db05d9002663fe84d1c6bdc5c3bcade76b64c8e8effe
zd6f5b733b542a21b7815213b3145f3de2cfdcbbed8a5391b8c3f3cfe99014ec0209fda50eaa600
zb57e729e1c3768731d85fe3383e60419bdd2326d60cc9c9905d04fca677be6ed0c583adae49512
zc38287873525e26f3c658150d67d135e421f6fa9a9997a54d48dad32a777678c50c316077c438d
za3bc939c3d2bbc0e2b1043a9e2574efc12e8c46e350befe2920742aa415cd341baade4d2d13fd9
z35d05ba9a1ce80e12dbecf28c88b5278b14d72c0a5515ab50f52bb5b6613016a132edc7e7adda6
zc0a718cff00f33d155d60db4329fbecb3f1bcc2d50c38a9dbb22f200a3b4b3bf6abf2731eb61d2
za7f082d85511d0e2582029224124095ea91046c35443c4bb6b0ee1c005e1200450bb4b7899e804
z4c53720f96f99c680a1f4fcc01913ef757a3620ad79132aee9f9920a181312d3d1b587cde157a7
zfc72857c5f5b0de00cfef519f902b0d61667842e23aaaa4c6eb1e2317d1ddb37290afd0cd31b8c
z10a38bd7cee7cb6b8fbdafc325c77353534232c47b772d7c296a2dc09239acc2e3f4908aa64033
z94ed5d67d2e1a7873c0cbe14b1596bb1403d683c9682248e05e2227617edd34744ecf84f5b53e6
z9d8dd723c4e0330df962d8d1a286d6872e89cae71e630596fd6cddb2805699ea629d9c5a225798
z5c295bff0903a0e4568b283c27feac4dd9dee7da7c55bbce0189eb3540cb942a938a19e5efff31
z96a14e4b7dcb8ca40150a0af1d4f7198fc6347c5955deed7d061602663f746c6c9bb18e215cbea
z77b033db4e031f3fd13cbd7f82629608a255d46658ff8092e77f620391b4fbf584bccdd4a43ce1
zece4c4337c3833d7a9ba70871d2ffd71bfa6025154582789efcdc40a9269679a8cc4e8bf8c7a79
ze12e0ca9fcc2488692b54e385833c0d6d474da0a1336932c8d1a37bbb794258890530a3746c8ed
zeeb492f20c0d1c79d0411a9082fc598ec7e4e920a042df4013144fa826c66d4f218915160ac293
z26ff75aaa1d2bed4591444dfa85962034407ba60e3922b73c4ac378e2dbb8bdc0762fc32aa6667
zc50e410c2eb9faac6aba7507737644d144fc2e5bd8a52f05fcb3a3153a848904b10eef65f52f0a
z745fc713d61a2f5dcf3333708752761b97b9f17fcf7b935537bd7545f51d2cd8c133f67311da28
z1139e355dac6cbb0918b983595bf5eb01385ee2bf7052a8074a570573f473e3e13b3f621fca7b3
z518b50782d67b254fdc847e4de55ba44837e70cd99e1f0f2370eb0a3af64e8a34a63d7fd8b3981
z729078b96cc93fd30c8813bdd166eba8f9aae0988a1054654ac210c6719cbd26df3901878310b0
zbfe3af790ead02cf4c1ae41ab33a4a45ae4174f86ac6115203349cd7c8d27bb3972f145c471ecd
z87717f211fce12ea703dda9b1caa6624df8063542d3c9895bf8dd60ba223be9265e5b0b5c39d2a
z017daf2fd776426a09d33af27bbe475a438d1f34c8072ddc385bf38e669b59eb038e7e398ea48f
zc6cea998b1251f29b37b210eef22ef6e0959946607be0f0eb6315ceec7b9ae5f6c2d7950cf135e
z546d7cf9070a7c58cd6e43dac4663047cde8792187a83c4ba15eb7a3f44fb3fb6fd4e835fbad62
zb2b044b0e22e37aa3f339bc9ca2d03e7929b0e3cd5ee3ce7457a820da612fa946386ed74e0576e
zbfdf2999ef82ea58b7b0f64cc6ba43300db7077151fe02c55c64a217907dd04f7ce99ad05a6325
z28c326aac5ca742cd01fe9712ce4a68ac13bc6c3af7469792498ced6ef7bb8f89f19771b1d9922
z3f241b31bd2cedbf6bcdf11063819f4c30f0d1815cf3ee67e8270650ab2ce8a3250cecdce9d6d0
z0853b12e3fe8129136e09d35428bdfdc88e597120571c9694129c1c896dbda91a9e4057f88f53f
z6ffeb7242dea6885c9a2e0a9605c438d494553168a15f99ce86ca98257a7aa84041bf71ae69504
zde8de04e468c236b62402aa31b86dd0e9fbbac4af4e0931c60a48706f35ff5480cb3ff811ecaa2
z782dec0b293e78d88dd98282c8475f3ca74d875e69e3d5950f85985bdcb18b15c7c570dd5346ed
z472c717c2f4212b5f8fb72ca6ec19a7c708aed00eeba69637ebfa19748dc4c6e3807d5fe397c03
z4b34d3c2431db9a1930c3e13f0d2727a5026087c6e29dc25a02ba2fd8eb88181c3fe9ad2f68cb6
z9aede8b70bd5a2429f10a62ed9a7810feb75e3f11b4f574cccabbd9800e0bc08a20835e506ee57
zf6b8be91c41eb387b1948f4b6eb4dcc4052007a1ef372debbfc393fc42f40fff9498290bc37d72
z58cc8fb0805abe29ac04a1cf965cff4d06339865b2bbc8cfb6b9c48d7b88053be1e0e854f949c1
z550dd62d2c5bbadf4fc65e78d5b1728dd4d84d91a5905225b408cdd26a65817ea0730884280002
z73a3bb3e8663ff01c79ebb6de16316a41b56baef4bf31570795a0d08829863304ff23e8eaf9a73
zeace56a6c265bfc896c535618623c222948ab3d4c2af7cb55b41a7dababc3631e74d3d65cd60f6
zfe124dd334ae01c4c725ee0351387c878e92c2dd582de81d220cc21fbec2bf6ec0a59f1ed7c518
zaf29780e704cd471687e28807a78fe43f432eefe76ae561394843eccb5a8e807ba515138b2cd63
zdf89def5473c001e3450431721775c9f29aab5e7a802a5a56afda014fa90cd02ca5ec9996c40a9
z21b25d20040f539e5b38530916d16ee7514bd9c03536e55eb61cd8692108e241b8ba9ea17bb473
zfeaebf3953c9b1630e1de28f154edb97896ecb9634323331078a4a44fee8cb51f1134926f39e84
z5fe79c0d291c5e5410b5f98c6fa7481846d263b528411a5b310393abd7ecc82dbd6d54668733df
zb0b46625991149595f226a54b17a7291cacf6f90e9d331059f8c5f4c5bf8639e4ba71609d39ac9
z104ab1efee48e573f422a3b28a6de047ef49ad4aae13d04a96964d677b0d421a47e7435d296585
zdf1fc45e52cdcc55bb0d4ba84f765b101e55575cef326bb53d8ed8df29f8215fb1faf97adc9de0
zce0476c307f82508d0e6cbc1b05f41a72210cb334b47fda03536cbec462ac179b9c3c88de20010
z94551730ae106dabfe0faa780d435d6222be5431b72acf588a810847ce8159639156597f6dfc67
z21f57efae1a4a7afc4b517a5eea758e7fb5bf7c59969c81319087203a0cb5bcb1a489da1412a99
z9ca9eb8249d90215c149724d4158d922723f01618c96a032d58a92fd405402e199f63aeb833000
z79cda6ade3324bfabf8a8541a1b34b8d05fa1fd60b7266962f8a25cefeb3639462061d32e9a678
z09a7343a596dc5358e653e9907904bef4944929f4e7e261b1aa9f96c606a0ae7c2c27df9b103aa
z8109a55d6aa838e90a4285d211ac2a0fb466300ad9e8e1f0b07abed27999837be7ae04355402e9
z009075aa430e89522a769980d07d471c0a34ce813baf5f0b2c9cb51369bc8375b98879a7e7ff59
z9d5c959c0447e3deac5ddb4adef1df4b6bfacbeed69a961689b992cf8f6c854958ab2d379cafa7
z8802dc153b971870782e86723a88c0c080b412504c48d521c145561209afc453d39ce80b676a54
zd09158f734168a3c40512a065017a3b20c09331c4eec3b4b111595387398fcbab1dab819423912
z4affc3eeb30c0215c8b3f2c1b22564da324ba0e7b5a65f3383509785d553b0035b5fd8090fb1f7
z7daf09bada5b5cbe63170ce1fe04fdb149cc00f47005680ac9d9aa1b61f780679d1a31ba4e8eea
z7810d36d8dfceb6b11adc91a9ab398fb5759c4a5d10d73c0ed1b1cead6f27636b649fddda7d417
z927679f217db0494cb781dbfd88122655237526f53d2b3fa63e5c82277e738130df5575df507d5
z2d747abc4f82464937ef871afedc8363b69faea0b2bd34c146ce2772ed55a095a47d7a943c5927
za740f802bb8d4624c16f14facde3d20e8f907272180ac75c4974ff1416a5a963d852518a5a0ca4
z507107eb1c36756fcd622681956ee2b153f7f5608a33ac8cc60906577f0e92ba78b392a44fb19c
z534929c1181894b2dfe504da99aa0ccda5561b66d5304121ec1a636496639a35673df1b685b817
z3106d9e569836d1aa5d7599c8f024266977eb956b024f5e29d3c27f49e47e27e9620458a33f5fe
zeb9b84f5a5cdee3174ce29e5faef5626c1e996a2443de4ace21b3e8268b1fdb790f5edcda871eb
zae5a0997872468f5ac8a892091da4f508464e23e65f63018071e5cc26d3eaa94c35691bcd5fe79
z81c8af34f8d26fcb831eb72dbaee8bd1536ed11eee589015ee92581d709f72bdac5dd21235f2ae
ze4764427bfeef45156cf99cff6f7a0fefe2a6721065ccc2462603b0dad76caeb047d206f155847
zeefe70b6c88803ee3c953ab0ad17a2ac58ef3d4338bff075c87f62517829e1ac31446674d4e0b7
z9006d08894172a46800b209c61a12607aee00caf21bf4c482018eda1010c3e1c2b4e7726e54065
z328f1f75fa7ed2572f02e8381d51dc1682c51cb424664aaac7e332ab91fbe65f4210282510f307
z2270d1c2e56344cf19ba256cdb39108c15ea53fd4d3b9203447df3b7899a12852485318294a420
z038b1cf75f705e925ff0cc96631c8c77fe5c54455d371e097ca0c7d516a6fc251ac8e3cfd0f531
z41949e20a981455f1f2df5d791a26a83da7fb879b06d1ad44ab857b1790323dd2a093790fe2522
zb0a22691e3d414e738b0dc27838ba7c39d650ff183be43f5c23b63897eae8aa1978f4d6d6c5a79
z4b856471a4d0bec7a84d9ab8878d5e5e5cf4a3110e6794400632bef21d82e569655dd355123096
z4f0a3308d55acfd689adc66b7eacd316341361ed5e308c0f5dfae41179ec406ce20faedadfbe3b
zb5f48a00cd05b902524660d9ec61580055f7ab6738cc3b26bd7a0f4fdea0e26080a8aa8d469108
z793d48ef5ff1704db841dece6019a6df57c028688b96a3974344426958656a981d2e096a512e23
z83a3af6a775eee32e035758d8f16b02955c4934fe3a734ba8f20c95696ea39e220365d86efb4c1
z9a28798041c4f22033818c110fc4e39597e90070689b2db98553de67b90f83a5d05e541f85c89b
zd4a492de4d722627904541dc5f2ea1d1cdc04c29fe60a608a7d5690793b459dc5cc09f412bbef8
zfda149dbf15edf5c8900852d3dac09c76e7b3ae9137db52e97d998925d2e5dc862da19a0bee5e8
zf1bb10fc14461846df6bcbc23ec5dac297357eb8e1265e3c9a7c42cec615c82c2ed9de613dd346
z7221b2064a4cfc7b178450af9f7eae8a9a59c5d57b1b8cbcd55fcce0be49ee63d9d49294f4511d
za22795b43d36e4ff8363281330fa761f125723895250a567aca5468caa3345c4bcd9ef85e9cf2d
z27b3ecbfb9ccc984d440afa4f841fbc78a68c05a011c236ec3a46fc23589bb0ce8790bbac92b65
z7cd174c4a5c1983925d56e40cc2be0876f761d2e3fa037cfc050473875b827fcaf18ad6514cb7d
z1cc6fc3fba6d07ba55ea8231873556c89ba06f6faa79cc3bde2f3cd9b41c0b4fde280e0994a649
z89f5b56fb15a73dc46e1716d7f968462bb371c150136e176f094e88a11cbbd09744a28fa8026d9
zc3549821b80603a622d0b4fc23e53b0627ebc1e5d44d0088fbe070b273fa2a89a989d10860180e
z1d4d4cca26bd99c0ed7ac0f5918c4eed41468313cd52bef75b0bb97d497fcf11091689e63f6e29
z57cb7e2b4851e2fa7c359e934daf47b241ca531b5d7f1b1cba1952f235c47d0ba80b72ee9bbde0
z4c2b837d125fea18554048064b6e66d2d7c907c9b7ae7bc5a820d9ecf3757676e9a26a629b52d5
zeb94eed5076b830a2d01a47f74c3c47e501182556f26b1075fce8d1d07f5c01e650195ee5686c8
z4a5fb2880fcb5ace7d5dde8660dcd364e684e6c82fb23139b16e7d073d588a3d14a2cd78270c6f
zbbd1f5fb89a8d96799f511acf19029d3d617a734b9647586cec99bbaf06ea8ed769ed373341906
z2fd0156f22083aa3572a74934e58a1515678f98ab2db26735d406a02a8e1d48ad995646f6111a6
z19dc420da1a728ce6c25a7cd0ea5d5051c9a2f912f94da001209be25e9d1c0e25a813264617e4f
za6e734f8cbfcbe457dcd7cd93b19a14a44ab2bd5f178b17379bd8da816e9cf82ce48741f0c9f61
zf3b5a595c05126151c5c8ce6c2515f54e2d3314a809f1a877deac4b996ae955b513688f907ac7b
z140690186e120f6e279f75fd9f2ab18e37d3950094710b021703acc89cb76afe560b8ca8578c8e
zeddbd66cbd9a5fdad56591c1b5bc390e57dd145b983adb46501a37053c28245e47ba835c37237b
zbb06c6caaf8b0f5cadf4009f59144075d46a7068959cb961a606a66f3a02b1bfb6b614cdd41f67
z161d64e12b4652921929b24fde77ece4225efedbc7c538f5a563f60b7d1209c4596ae362286884
z6485ade1a1720af475c20a5f39e54847fb8311fbc4b43394798f0cb8652ba538488402c925f311
z07c6139015bd4fbcb4cbaa410ec0dd25df91a766ce91323ec3490f6d6877b0d667aa1083ace3fb
z7c55baa38e6cfe6110f9565efaeed7503c11eb39d73d44399995720784e53605239c6fae775fa0
z4a6e2fc530737c35fbb1effe5ed0f491468dca76a125f704abbd51721a4c4d29cb37761e23522e
z4793f29eb4343df466e3294a51e05de004964f068ea1338c00a11eb2f0b5f8e45109ba92db114b
z9271db75c3b3fa20df8fd34de53eadf67ceea225ffa4e5137117246ae93539b91e7f4caeb599c6
zc8d33c623f8ebde9ade446c7a51501b5657e354f755a06bd9b9e02fd481d13346debc91dc9a59f
z37f53233f33fa552b7e4b4ef389c6283dd4e90e7fc503060eb3a3f66966a498bca56c1f50d4cba
z79d6dd4dc563f5fc96ee40d9aa2a33f6f0b77ca99e4c1a79f782a6ead7c1482991fd05cb85c3ac
zdcc8b33757e0a34fcc1e0c8500a9a82317daeceef4b8f8e591e7b7a22c9f4b59f815cb6ccb7d46
zf90c60ba232a24b48fd548bfadcded17da85de2f42a5f62a3fa77ff274b984ff0f9b7dd40d3279
z7e139e71374516c3a8705e2899180b4eb8e47ca456b13ddda15a2f99011c2f23793050719a4da7
zd444cf74dd7d5eff4a39eca1215d2597bbfb1a6147423c9aec89a657208fe14e1a3a23a8f2c176
zfa7c089b4b52e6c5c355d9a76923324ff73bd23fd2ee0ca45f1049e9fe6fdeef878bdb2af02638
zbdafdfa04dbdb96fbb1aecaf3be090ebed03625b74b10467f90b194e1a2a6a272b4a8552377ab0
z95ea08b4d995d91bc46aeb66aac1aa3643c1009a1c4b4417af2c4e1c74266639d33c943cf1cf36
zae5ef9874b7e1f325dcacc9b2d2ad57d3a747029fec2af1a710f782fd60a256649e3d859351cb2
z2f46e4fe54ec9dea2c551ccbc2937d3427668af732d93f18a2083188503d4c80179e854d71a4c0
zadd5327f52efb9914e59dc189e5861af946aa8228fa34d98d04be2e9b399f53bad35e64481e293
zd5295fb7e6f2feb0f638528489f22594573a9b0f7cb431bce922210e8c6ceb3d6613f5c3b7c964
za06ee41b088aa5a159ff0a3685a0215e29498128edd0643c5e334e81c187bb70bc29d4a50b0c91
z0c39669bd6531efa47411914e19490ca88d5d70509ecf29b41aa28b676da7841b520896cba3288
z95127b4af3420fa784bdcd27f63f2935063b6edf79018c1e000289a61b9518c3e63eaa4b963e73
zaa469f5930e1e27dbfa1359f525639952a6c6486890d683a47814d5e96ef1a37b4770875125e38
z0104f03d7641d6d1d14f533c917eadc3bbf0344dbb1ccd87af368d2fe33da96d08561b57160e0a
z2576083206a4a628892f3a963115aaba13bcd8182d63d4acd7d769f87a799de2a2390805712859
z42e96db0d0b5829f03396864fd343a65963aed379ba75bb89cafad719f2860322abb19dac6ec89
z119069471838d70b37ce8e836c060ef3d99f06c472958d657425597ef4d6e438a2f50ac08d9997
z8d7caa3db9c5f834387252975bb870cdbe549ece3e58602c5c3b254c761be62be8b76229f699fe
z8d825a991bb79658c3370fb00fe91946016ffe0200fb39549f3749a43f8b2a53917b41763a0793
z88cf8ac85310e36314fd29b6c74aee2c9553b32919602bba5f62f74a4bc812f42334fd0a17b0c9
z7c5b419f61f59a9041deae143ff91614a2cecb0d3f8b2cd301f416e95a13f3078e960984579b8e
zbacc8b85f9fde522a2bbe3757faf8e1cedf8abc0f5ddf7041e31010cc3643bcfd4f5050b562a21
z3cb14e980b97b869a84fd91b4b3baa12f5f97dc8be00baab270eb912d403e714ab607c4eea0a91
z228f5802a88233d5972e34039e540d03a94732e7df85073da7aaa78ddb7d9ffda7d010c651a139
za182e1957d07f198c32c77d1d870e551604c43b95301feb7009a0b7566361c928a687b5cd18ec9
z9667e6767da1fbd2a1a9fd7ee1dfadc136fe668c1bbcde1eab172b8cdf4eab38a84d1c636b7dec
zfe9ca98ab765df3170bae7d13a1ef3e33db4369f07907957bd8977470bf98abe8114043dec9cb4
z5c4a1054b6d99e7a43a1d33080216a5b93309711a107071130611bf51230b4601f88b7d98cfff7
z3a902995b8da0605a1c81c4fe77fbb689ecf52ea3597c22e8c2ab346b782e1c101d399efe36b83
zfc0c4f460c1d02c49d18a041bb63819fe31f93902a8d604bf40cf932bbd60d3fae19ab02ea09e9
z87577bc063b71bb7153d6df9afeb32ba73365adfa614acaddbd82b44cfd5099e5a63de90882770
z04bb372476e6f27f2c777dfc987bfcf3233a7a180c29974cf5305c2d6c7f1cd43cf445ce54e1ff
z7b6788f96acc390a2aa6c492d11e13cc6cb3f14161ed652867af5f131ed78d90cf8ee7224f52e2
zc46744ceadda1dd2fa3b311f33a883220c59ed9d2a002017773d004218cb9b2e5a3b7e0a518e78
z490740f233caafb9f55d2b2f2de98a5f9fc8d893155a9ea53767401fe295848d72fc0a26ad4afa
zde31a48f4ed9c75a8f1e81ef7347229168f0f30f78ee7caaf8ad20891d1db2badf24eb5f2edcee
z7527eeaa9dac45b8f1b68f897b1969be7a5e51977d43eafb4d2738d48edc2542b02a297067da6d
zc1f854b1d535ee86193617df9eb323c16523b59c5ed2cc4f94697995a2dc00e79dba4ad0853a3f
z7ebbe8f42e0e3be2149e981be07d340ee3f77d5932f130be3cad92bd8a648290e6908aced59743
zcd42185e184d3a0a0fd88bca9078678803c7d8a4fc0ced02080fa10cff340efc88ee710738dd3d
zadfd8a8cceeb50d2758b168bd43dcfef0e4dd0a17ea6c0bb718e32731ee2aae59ae6e86235907b
z26f33014119b4b7b1b6fbdab980dcec482f02a3690ddb949f33fa730d697dd3351b6d7e8c320d2
z9400052ecd2c2e4b51723a7907e71f3155933345d4ed30217fe042685551877b1c5589a05db603
z197297e23b4394553ebaded55ab4ffce43b3f84c3875dd459b0ad2534ce3cbf1ec10a15758c28c
z8914524f31e871a58d6a6867901c5640117babd374fb3d158b40bee1f764d83ad25630b3dd3605
z30e0e167ce3ac88f6cab4fb6266f3293b26db3d3f6ecc3411a3062bf5122104eba8a19a49bfa89
z6ef1c66bc275a115a606b7ccfc1a54088a41d3f92defd45cc4f756eede67e0744d544a210ff0ec
z5a9fc1bca6e73d79c6626c4d69c7691ff5234dcd0751d6f718c44f595e1a3d029bdb2695c41c51
zdfdb93823e7079f2600447878190fc074f16b06caf11c951fb30efce8e59346a999c739664574d
z01f6aff0d9513a19418eb34a7d8d6b9222b830a6651276263eba1a2d37fea327c6923f663dc809
z9cdb50f7ecc57c42fe7566eee9e9029d0d0556f3f84ac1658aea05e9a307fbb6b822f2c47856b4
z36eb3242e48d3c6e8eb4319f4aecd4e8d797bc7f224c60f09ec58c173521d765bef21d80242c51
z6ad48ea700032d048f4baa0bdb717bdd40acfdf3bec9a771943cda2bf7a02d741007038d565cb8
z5eabb5295a05e97a9912be75bca7f7effb7c131cc5e226935cbb2e9a5806c8f51bf3517b1687f9
zf98a10b897ec2d01cd35fe926ca3f937c83891b21e9151a05cfe5dec54db13162c817f7819b359
z06faf497dd9a4d90cf5a41675363401a7294fe50a71bed910b96afd54162041d6896a15eef069f
zfba8a9402e7a11a9ff096a4b59d9c3ddeebce66b7175ec9a9c83c2122b4522c1343b34af02c8b4
z7a3660fab2e3e64ee144f14c51d8d313fda75fa22e66435cd7124f4b95cfbfbd06c4d9b2bf0ee2
zed1a9e511b86f65e248946bb19651c1b40f94f9b0257fff0a3fc920d8b5784cf7ea6569353b429
z6ce6eab12ab25702d8fb8fc78c9eaa7ee5087e1b456e59a0ba4eefe18390e790218c4697dc1fa5
z57cded38e05977faf4385c144e35bc39cef40dc122ba537f995cac8ec124f48739b4cab565089c
z5dcc2bf605a2654340259dc012eb7766791f40fb6aa1964d3257a78e0604d25cad223db2e4ccd1
z21f959283984c12d49457f846cb08ecd2dce11b0de846bee5bebd5e03e9eadd27108849c74cd57
z1274c67ca68c604d415859901b91ccbae42ca09f6db3d746f02a8ca08d36ae7d138573b9276839
z7e4c043eca0e32b4d2f9bcd1c668ad78025d8ffc691fee5804a88a535d5918c9a6c4212f065f90
z0e8fbda6f5d6526af102f27f7bc0b30a50b39db807a771c5981ed097475bde63ceb6cecfc0867a
zf4d90cb892aeb2d409fd7777ad7c3d43d59dc7ec5cc5d4e9d6be1cd0c41f66820477f2dadcebc2
z948ebea098287a7dbcc63e2a7237da57921b668d498d4360f84949b4683b2cf53956e7538cfc80
zae472a05f84bfea32a4237917b2f3efc126d944f22d55e4e27af5f83ba907bcdcd942b5f5354d3
zac507adc9f0934d854b5f53a915768c84e80d8c6ca86bb94841b7901c5474c3a3bd038581e3cb8
zf034e59f3c724382982f7fbe41123c73769be9c75520138fa110d71f37ea6280871e1cc364c6c1
zfeee29522f621210d5191c51e563766e43729f5d0928d32466a846fd4b755e858c6f2885d0991a
zefe018cef4f8a57f1821dfd78ebbafcc590e06bd89ccb0b073b8cba5d2e8055105be4a16661f2a
zc1f2dca3b9cb8d6acb41e68a8cd5ec4e7953f534c81f23ceac10da8a299df075253508eeae55ad
z6a7107328a6749088a305b24c88c38f23569618fd52cbb3247a653657b27f733699ebcaeade756
z61499bdb1acb8d703849a6694ef41917d5e4573ad83d7c5fa6e694f047965f63cc0272b4b23e11
z9ccd6b66fd5ef923c386442bc8ab9af5aebe6984f8f6c4da8fc1efd63f74cf18cbd33dc5998a9b
z19d030d6b29c5e96b5e77d9684b93a755c911996bfd7420293058163b72a2fc954b8e5916c24c5
za103f78950e7c54f486fa790b3287b4c5e70044b580fe0e3a49934f1950aa56bb524b48cdc79bb
zf48f7f54b9e23e311a2316a2f294a3a0af163a96075ae07fe45fd50b6b591e33c025fb98344b9e
zb1bde600e3be82974403985f234f647859793ccd69bb2937380273764547690aae8b59b0fe14b1
zaa3c9dff13ca7c780753f7daa2516a5f9f4a05b3970d4dc06b5a96be0a162180a9354ec572c2ec
zff74e312d2252278f01e88d0947022b806156fa60f5353194b2a20111317e2e1829c16efecb14a
z826591d9b572053aa14efed9cbdd0d8e1ad11faa9434e5771773c4e0975d2876b90ba90e021fc8
z7212a49b7573aa7cb5ed98bcb6fd88b306f94b37e71a98915a540fe1120c9e65d2db5ef0443ed8
z175a25297e1301bba432e479e8b0bdab343f29ce7d6fe1f18018d53e8af68ba0e6398dbdfcae41
z9937ca2444aec8db14964ef2a59af20587734f585f63b87a0fa49f04c4a93ffa52bb93dd5b443b
zff5628e9092a6262718efc3cd1387e57e1a7b9a0c392585d0eae68b6d6bcbd9397c40e9ee06706
z90caf9b4261c3ecd997882cf24b00bd01b550caad869ff608062b7b871d1c1d4aec30c246ba0df
z34632748d4bac2b1ea7570cb8f5264ac4fbb8d6670df031ce45c8abca963cd15cdeaf6ae914b03
z9809251dfa225116ab664cc921fe44535c7a343ab48147a980356e3000877136181708fac46880
z4fd0565879c090b20a442b80196e632557ea813cc7aec9f2981860253336fbf95e4745d153af4d
z9e1cbc87147f21c54e346d0928b6b2b31baba9cb7184be5c8ffd8f68b9f82113248c45d8ce8329
z3cf1beadcec83e2a3fc5dcbbcc058507f00a9e8557ee8da18a6545162de281f4d64ecf33921603
zd8560f2c7f6ee13661b1feece344c58800659f8e4104b7213a086752507569ade2f7fdee7502ae
zf6fb1b2e0a7c478a5cd76fd4b7428e16bcb67a457cfeb17a86efe2333dd493d97c4f9e50a6ec2a
zaf34b662b6e890f27ab22b37f7ab2922da0d79fe4064f6472b65f432bab461a4d94e32fe2cb7c5
za3a8fffa4f7449409b87160638c65b0708d99897ec9e7587dbe94c443c0884468c20e0db1b6685
z97ee9410b5d475021a2ade26bd0f92aea7480f0474bd3e22dacee8886c82561994bc9e61e8e1d4
z0ebbd6c5c098f7785faf8cca3abc01f79b19132d3c4ae9585fd6484ace9f34982586bfcab0b38f
z39a69df375276df79078bec3c21a8dde3b5acb4f9231cc3c81c5083880d001cf4e907e6c10b1ae
z0fa38a66d5c41555e5f240af9ce49e154026b241b4e7bad94092c30f51331471f608d5ff8a1cc7
zdd704a0cd4567bc91079b21560a7c57b55af4bdf3dfe4c948424bfdba827cbe7d9762e91f19402
z1f7ffff11b3457d225c2cd5e79f4dec8c173edfe0f40fd0a146fd96809e83ce562c0ab51dfa89a
zbdb5d233e3feb047720ec4b91265c553cc9f4a5aebc4a74259477e51d240245a69b2a4f831715b
zb2d7cdefe666f76a7666bc4370f21f2be233c43e16ab98a6895cefd4f5254ffbc61bcdb67d0dac
ze0900876f44c76e5c15d487e990081f8ee6b1d66b7d6cdea2242456e3c3f832bb9fca2648ad585
z64889371a255cf8c9f99fcaba011931b1eda8f34b82764cded71f7b3c542f2d48e56e5b3448c77
zfc23dec9b8a6412e7db8feeaf2db676a7e5183b02c3f60b4ff61bce5c1ca847cc24c2b819e6168
z285e6e266c4328a8e19f864eceecc607336fa099ba63718e391a2a91c99803a67255647e084142
z073e3e615adbd3a53a604d10a177f04f6d4954936723275c34bdc030e9cca056aa863d00469a13
z975598729aa7866c649bd047bdbc0dd59b9eb760f13d35be2ef9b85be82fb4a7a02d6bddb83a74
z0a35d377481d54d417e88db15d047e944143eeadc884edc1f68c473cdb3233c042482897034547
zf8bfad4267ad5c5ca811b3236a6e703a24d21cce397e7cdc167ef7c0065424954acca54fed77b9
zcc782ccdba6f65f416996713718c165100c48ce9f39d43bc360f34b218028bbc4ccb220f5d5708
z071a74e361ac4da5030c4b6103cecda040d4b5c12b0bd1489c6a2a142e314cc5e45e6dbed5da3c
zfcf8295fc83606f31fd38b3493d0d0397064bc5539ef1cbda438b3b94636c26e797b6e7c9b615a
z16b02350c6629ec7c2ae253e37d9d8473b118d43e5ff554ba9accd85ddb9b592bdafa5d148ccf4
z4780b8152e3b4ad6cb871c581a0c07a45d2250fd3dd58f1400fdcc5b521c1a50cc1f812232c7c2
z4612e444da9a40c31cab17b112957088c3f89e6640950a04f1ef710c2048e000ff156ce3a894c4
z3618b6c319df2419743f3d5f361d5a6324a12e97c41534cc45d58ee4008f62dc8b097ec5dde447
z5673591c6bb1959124d3c01385f4da40a04b42edc8db72d067f3cdb41af838ebd1702492dc3279
z57af3c242facee8bf567a816bf6774f4e3b8ce2369c767caf23ff9505fd7030640231eb373fc04
zb31d529e2ccfcfd787acd783f94bb0114c70b0d9c4e6db1c0fbed89ff3f59b11c5e75debb4553e
z79b3a6c243081f212d34da648aef417fe19795d6a7f4c75024b5d230bc9440b1999ba7488bcac2
z90ba0a6e9daf8dfbbcb1f35f7b1513b290480ea1914d5484ebed8b969345cc110949f180444cad
z47abb1c47cf869a82ab7a6d0753206b7309b378098e8bb675f86f553c0fa7a51c266eda8afb370
zb406b8528f599a9b04cf88840a1c686da772aeba4af92e5a7cefac0f92a362a2ad535916ead788
z50638a8e30c45d7ff3c1fb5b1274e8270ddac9d8fb54b50ba6e68d6f13f6dff53d2dddce3f2210
zcf5a8ed210d52d1f6c92a23897779ebf6750b02844c8215e7cd34fb597a16c40f60ee7baaf1eea
zd44dbe236fe4206b4226ca93ae53f0d45bb58ec68a1c9cf26bf914f6d5524203cb5dc96047d07f
zcfd4132ad80e869aa5a644fdd18cc7d52f239618229db45a5f7f05612c8f2de8c997cdd7fa2787
zdcfde4740cdb5d21a7e51b9f0cb1f4f6758dbb50bdbf995a7f1afca9b6c02608900c1642168675
z9f125592deede8e32505fd5b1a64140f78a3c2dcd80557132ffc3fbc47e53dbcdb80c784a763d8
za048602777ad0f634f71a376f2fddf57a15c4065c16030eaefdda6b51d1b5fd901a74b3e353270
z8b502dcec159c7d45232588d99172084887230a0d3cdb6ca1929392c7e3f6b83c00e6697ff8177
z8d15adbee5b0276565fe927635c5af2c0acebacca6d8c34c506a0bed6aa69910374104fcb456cb
z7989669aaaf681198138e67cfeafc15d5d5f9d643040562c33c2ba6ac5ad2e4d876bbaef603dc4
ze80ffdd3c3f6ccd590d01fd00fede16347fd11c138b6672cf72a14754253b91da03ca1266b0393
z9065ee0acb4451e1e56115dfc2a2536637c8004916058084093206e56a20cbf4015acc9642e064
zca3f781609401397e6df109e4c07c4303d4c0cbdbab64f0165eefa977542d11df0ab74fada058c
z02ba1bda5ef191bd34bb59342c25e6fb64763e1b66a4e9084a753d61177ea3ce17ec8f2a62c708
z70a0cd1d5378056b502cfcdac4d56a38865e577005943c88a879b5c8b2653d265113aa5dfb34b8
zf096d4b5a31edecaffa38e156109943c77de9aad7941828a1f5c099b28573ce37ce554e49b90e7
z9013e3e0951a1a672a7cab52f20f7465d714b2bc125f387bb4b995ee04983e1267edd3369250c0
zdaaa2660d5ac64130e5854a02229e04a22b9945ba97c6d9f0e4afd214a553b1c9e65c2ae86c21e
z1becf47059006d7be8d94b539ec4dfa794cb5c1e8fa1eede677b26470373c5ae3bfd703b05ffe3
zdb8b8cd6a74a91a4c31747f24e732a947b12df95ba2b989bc9f749dbff7bb35eeb33891c63cded
zb582927828b2db6dd1ab3b4800a9bd4135713da208ddf3c75fd3b48ada012c4512ebb848e45d28
z7174058373da622e163cea6c92ddec85cc3892feb53a3d5f72e7482c0e14f7cfad81581036398c
z68238d2313e63f57b2d7bca866fa03642d44d394ed360712b6b4b697bd7e27eda3dc74857913e3
z52ff84c75fc855bbe9e30728d6a8ea56de0be432aa325685e41024110b52c3648ecd0cf83bc70f
z10a85968b062c13c7d2ec2901c1f15b0835772fcbdcae3a3c83ccf5d3aac747608f5def790079f
za7ada7be0934ffadf04026be597202d93af183e548861e21b90141fd88d0d4a353ebd705372f9a
z899f1b20edcf63b265d4d12c675e24f727a7fc854f655b22d810fe3a9c6b1ec35a28392a3f9944
z9c958658584fa7d237b20a796361d398449286a3ef4a5b650e6b4d6d2f5b01ab9c1f830bc8a1e4
z62fed4c958b45308468391d1c23f817f21b8f8d457956c92d615b3fc946d0f697ebccca08040a6
zb1bd44c89569a43724b06adcbe0fe7750bda55d5aa8f925bf842a038a72e96fdf25ea0cecf6788
z8deb7e5c49c0c7e868b7b157a4c5a00b5abb88b38f4cb2f029c9ae1fdc22b583de8cf54ea75a62
z7394d0f3e75d28a3a5a341ffa4151a17dddca714ec3fe20c88c388ccb4230bd20fed582ceb668d
z79ffd6643e2b0f98410814f1989b85184c9f578bddeb90286f33e6d36e255490abd9619543fbe4
z9886be13954cdb3c7c7e267837de0a965b92090a9a71f72093e4e6a0147a426476ce3412c1826d
z43cc769a6a6b9c0056788773e931654ef3db6bb90c849ab7d91f6b009d8e4a8e01691513f4649c
z6c46cc65ca8499be80cd5ccbd4929255c326dcf22c86a53de003563ef67ac467e5107bf7029689
zabd04bc7bc16aaea8b9684b99b0ddef1662c67272e06cb8b08f7d0f3d2a658d68e7c1c75ed6f42
zcfad4c1bd970d7cc87bcf7bc35a47186009a8e7462fe1fadf1cb88ef9f11a8c7dfd7eafe60b456
za556a53d4ef3ecad65b2f31778f82179b147ef15ce18bc77a62b589f14e4c70bc597a432140714
z49e22da5a98bc6d9343ed3f331ed4a1f7e68796d380f0e7cc68629adc7a8006ecd958302cef24a
ze215221bf2eb70035c27b755ad0cf31cfd0e192f53ce34410f3d76fe8a504277e4dda6a1d38c3f
z02f97fff0e6b540dfd89afc8c70324cef69be6767847ae9f99b9d867c5a76c00504690d69891bd
z5c16c2a701414cc9525f17e4f26baed7c236e1cf77773704b700eb702cd2f75aa69877ab2477c6
zd59e989a1109e42202bf911477c971bdcdf1d498c90d06584f3bdef8766d82e92aa1c22e995988
z609c41ae10178f8240cf80f6c2e8deb53f543ec946a31229dc102f13d4b0c9a1f0ed2352192e04
zedf1ee0d0737ded72c242cd7974ed3354a60aa69cad8f5089329911c16797dc9194b26d87f7b3c
zf56365a27bfaccb89da48bd248285276da4789fad80c43637d1fa2118c59e821b804a7105d7bce
z55042824828bc6ee6e34894f01126d3ad329cf0934c7e7d8ac05f09f6fad757fb86c79fb433ece
zb9590b9fff41fcd43180e7c2bca2d2af943c6203f6fd15e72990d79a9a04c109f0fe0a662e9313
zc689c3829d1c5dbdb4833ab810e691621beabf2ed69e8758c07ffee6795c2326217a015ee8f8bd
z6954f440e5fe69f7ed54a6da20bfdc56f3ce21c8eb5e19a5f425cee76ff479757032e908a94ffc
z951af140d7983de82f6df2eed136b916c8dd8db710768be0fd587dc6854d96b43ca2d4c77019f5
zec8a30e904f0e2a44fc739010178cd6107b2f98064df116a24e4f4db22d9b384121986a3bfba52
z40464d3c1ca0b6eb86f63f8d26773b25ae241235b08535df2c9dd1a8cad3d1a04516f76a126282
z3f49fb324c3f36880b81cfcc3d639c16ba7d79bc1a950fac364dd2909c7246050f295fc4a3ea0f
z91261605c4bd6733324e6f8df94c1b2787f47b4cec194fc10bf4ec655d892d77d037a262d470e2
z044af6d9543353060b5b28486ff6f38f37721ff24a971e3537f028d9459a6367fe0e58fbafc5ca
z71ffc76aff1b03d511716e636daf909a135233c4ca09777989cc9dfeb04bd9b5351850753200d4
z507babd650df712e1afca1440cb13c4d5406a8011c6ff79a74fbf6ecb1c7a5599d970baa41f40a
z82bc7ce8769a04ed8507f2fbe7615b2fd9003c5a00f0c35198e083e8bde07ab60c22ec45817b88
z9f6690e5f0fa1a030062efcc5a2a221a3172085232d930731d36fe9b18e687962cf5508909ca30
zae3b6cbd461f8734cc4e4e1ef6d29eb153d1e3a0d5b087c8a0b121e9f4427c8e79974583ff0187
z38163cd9797097917af489cc2a4e1864e0e460371992cf82aa2bd83cb1472931889fb1e003c5e1
z598593b9c209474ac92538ac7eeb0db3fe653783fe17210237d346de2a3bd5d27ccfc8f8898316
ze877cdde0e637e6e8ab59ae19f82222990b37617db37f3a88aab736410b7ca265685ae35fe269b
zc6b58152d015890cf171308f34d5c9bfbcf6ffc0c9595cc2c4360527c9d36c107502c1c08c4cb0
zf58d720e4eb38cb5214cc1fb9da81772d9ddde55bd1fce64c64d4185c32920a9035d52163ef269
z46113c364c6174585980d6976778420185fc5218482264cff27e77915bcda1eb74581edd378cc5
z71feb40efb19cf5e08a1a51c0fcf89a128e5279152442301fa8f9114e5a77022bc31c249fe27db
z5e3f196923427c1dd3cf940fcdfc617b40d30f59803982c408560633e83d025f98debc3a88a182
zdbb0f3fcc63deb674cbb86edad30f0719f4d5be33e58ffe5f8a4d6e6710ee499b55352220cbe9e
zda027dbff1643b0f30c9a14b9f71c0e15bd778ce3c093ee854b7ac41f232f9ac761dcfc3814a2c
z7349d30d9f7e3e3d5946173bd0208d8b1d95a4adfde30568678cf1c96e0fe3196a59c34d6a5f1e
zc5398c604f521f7e9e95cc2eb02c10fb04ea19fe0af5b420754b6b204b2d6fa6ee26f9466b56ab
za325fc8561a23bae473baba409fa6ff40b7c644420730fa6f57f683c6b65dfcf7ea899600bcc63
z04ed85a22da84671ee486af8927bbc996b0b131353670ee7ff5adb30206012ec51a5823e44b1e6
z2e969e0b314d498cf403162928a6c0e82560a86194347e74bf6b58f7f176deda0546172375e5c4
z1b06d57d50f67edce210ddf1abddf5b21d2a0f88bd04cd2a98aec10e312e89247190cf417023e8
z7acad2923e8d87ff95964a5537f3a89e311c62030b63deb27b4c0c192b25f86412a294067fc23a
zc76f590db542f831880a0a4e8d0fcb8eabda20cc75c9cd4a2499ab65f6f0eb50b70d066e7f6d82
zb14d07cf281e35ab3192b2bfbee09c4d7cc7a58ce9f72b8bd851935f58a0d1478b1c8e9b2f215b
zc75feb4fa725f5b50f391295f5c087423afbfa98fdad4fbf05e2a0021ff5a56ef936cd1d969f21
ze1c7ee5d70956092b4bb6e53673be8717524bb90c7c4dfe6a01b3e0f97aae36e768d84876f87e3
z42e9626b405ca4195d48b60f4c35bf85b118bfae6c1414d23a3f3d1adb46d10db9471fc7e69653
z9b6bc6c6ce038c52155e94d5bb9cf54db3b04e91df2f180b9c0e9744c7db48494359e8ff99eb82
z7c16059f68633a9abf3ef48288a664b061ebba3049fa452f83ad01af357e1af308375394a572b7
z0ff39b543bd4ba2207dd4efafcea5d2ea170c6c80ce4c507c8eb488c0ff66e067bc8c7f2fc813b
z60511fa07b3233cdffd34fd03307adf7f5beb8a7e059df3f3957037ddb0eb9c6dfb5238793d939
z2662a8549bf2ffe97654300fdfaf4080844582f361e15b64a4054506ba4f9d087327078bd24381
zee1fc6359b47eb82de306fe70cb3b0a3d645987c3c21c8340d3f1a8de4927cad069ef8f8b1fdfd
z45a724b5730455702de40a2251bf75dac8bfda30cba5ae0dd50ba6b3632f7c64a8d244b8f2fe9e
z4edebec907ef6f67ce30cd3cde7b589db14471b931ffa063e25f284d3e2c26a35e020a0dfa7f83
zff759daa73df6a7d5ee4a694e1c9b833eaba3f3aa9297217ca883787460867b6f8ba3164bbd353
z35d838bd40e50494710b829f1666bcc855ee9e71ca131f72bb7987d3c6d2dcea057f7a00386f8d
z0cd988671a7867d5695ecc853de2b1ee384519a98ee225dac4fa9835f4d056bf89268c0199a3df
zde80b0e92fc374b0b9e37a43985bc797d43ed7761a13ea7e9f0272aae9450de77950e819296412
zea4fcc360c1043cd095eb4b4b2f279c87cc490af37953fb8d189cab96735ab66a29209e7073b3f
zadd3bdc744a6085c164987c069ec7831a43ff4837e2c21f83f2b769262539d2c3cf71dbe50ca1e
z5bb8daac1b9f49c198fea2a300ab03afb22cddb0f81a779e664fb8fe6aa534c6395b936c5814a8
z645b6d953e8b01ac383bdf605d8db1ce2b7524bc6386dc1edf412826eb1fde2d538a8e91c08c9c
z7d7ec7ef5a8357935813170597a4149bd904366041e28fabf297dde6d66924b55dffdd1f807e67
zb134bd12d501d6ec252b07757aa093bfc0a365cca9bc080f22fb72301f182550335324cf95ed94
z38def3bc1c040360ddad5ad359bafb9301b50e42814c5e2996a69564a4bf82325b043c126aec3c
z7291452d327ef0a2dc45d554fc92243bf02d9f18f69e39ecbb5ed7d55f6b336d0cbbca2bea39c6
zbd4432e19f120d4e245fd4b10c0fdce28e5d7c3391c4d6589b3777a0be70f0b09d5fe41a8fa30f
z29dcd222861fb961a19ad6a6003fb00712580a5e1b10acc978415afc3b633b22b41c40ce23222b
z40a6f3df9e3e748701fc08a21b2e852dfdc0ccd878006473ffe9244df87ee71c6f84395c00dadf
z39842feb1da5f1895584aeb857614fd23242bb5ee52964954e01c91029439651a7f17e21f82251
zb3dc9aa74274f358ce936e58510746ef087a1d077ebd658d0f3f2fff34f75d3ec8d0288152ad8f
z8249132b2e65937be6dd6629660d8fed370138079d0e3fd2ed364cf63e9ee0a881c3af7b5055bf
z883dd8cb5709ff82ddcf90fba49e64e6df226813195c1fbc0c5aba6b4a177835e5beba15247697
zc324a99ada808cdc80420772cd42a6bec9d2498491ccf022beb12a5202a90ea7fcc319e2cf2d5b
z735cf5e7cb35e1ff29c323911a3b21827c3dda8f48c2d70502fa18bd215a5aa04727530c434698
zbcf891080200182c0971bac817806ba17f189e0fe4c7986a62f310f48b8a6f3529c69e51ad7607
z17a27939220fefe4e3ce1d94b17aee221d9d38d04e628793625cafe2de5eaa2b56528e662b3f36
z2c1746e1d2025b38cc4bb5e10176cc8aa3ec7aee7bb95639c608d233ef13a26177deed0b0d62a2
ze516d70610480dd48730f0b5a84c2805cbf7d33dbe9a61dcb0cc968d955b3fe9c09638ad8f9a88
z6c3673c0cda87bd62ca057df94b673b4f9966dd8880177dbbdf98adf869d5b23a967225ba72b03
z883d55d478bd77334564e0b5f123d32076fd2867faad84f527483e85a6e7c4715541370d53b5b9
z88a83ce06e51a0e03b9fa265fe62b1975ce3d650626e1094850b88aea1d8d4d501c518e493ce5e
z636efee0a5939dc43033321176e685b43a9734e8ce8295b1015d2c4759734087fdc37dd4e032ca
zc66e4d8d2c52a1a1c3ececceb1a0fbfde324539f22caeba97d0668875f14435b0e0b5b0a29057c
ze747b53d53ab569564774678635dccd80976654be9f85f8b1992f9a48b8a955cbec40b1cffaf31
z92b6f151a84781c3a47bfb8db06ab4aa71f4be96c173b193c1b0c808b1bba83527c11f2699f861
zec36df919fef26685929cc22078f5b4f67c3e55b594e9d6047c374b4e18faefc76a11644603c8f
z6a7050ddb7ae7c09897f9c28dc2e98cecbb794aa8d11c3ed9a88f02fb1d029f63aa87bc7fa478b
zaf15a7b714f04d679f361b4aa5d04d370afa4fbde14bd97ee9c1c43031b8cb27e4d6a8e83cab28
zc72d825ecf340171374b60b25700825266f1a29ad86eedfe0ed9a2e4be1436b221dd038fd14734
z92519e31f0908d726b2517d30b4f35da093227e4b05f85e58f08a4b8ac8d77bfa0a3ae010ef0ad
z57d5034a2f1b63244fdbe68b9d2fa9136de5ddd269ded644ab63b100535cc0a8b47760ce3b4857
z91157009af15f521841b5b670fe8f9936e8ba3cf2543715a37232070929d65f0b5c5b8d0e19f05
z70698a482fe266c2a0df1f8db9bdf509e5e3a2fd50f950c1f259086a8e6c8e0617cc9e57b34e06
z13812a308525c7b6e0a27dd53dfae9742634ef8cc403f654c46bd74f452f9b0e4054c4494fa925
z9c535f8a871c0bd7261eb4eeae0db9d95089d86dc4ccb78f508dd6cd4cb69f2e4cae4eefbce2cd
zb09ead7fccc343767431feb2fc89fca68d4845bfc19486f628df920cea0dd6258a6f90a7c4838a
z8aec1741f83d401610c2344c3b51c0bf1cbada5395d6be134312a85fb7e7108ec5c6ca063a512e
zdec7f4a740ea796e134baadd08c2859cec05cf7cfdcc114fc0469b3d6818c280ea7f1c2e794200
zf513fd95a8ee4aa43ccf6fdd2da64a6cb5f4d096c1e18e88393219514ba65b654d28863375e222
zc1ffde57ec42cb9ce31a1777319a6c6bf02fea8ca736ecefa7dbe46e6475c4f200576fe95ba072
z78bd3458f7d79acc35d33875c4b1dec75825139c2179d634268ade0ed8baae65f897eb85eb6b7a
z8eb955b53f38c139eb008c7a7230fd791a3c99f4a832065c1325d6dd56d720e1e10c9df929ece3
z9b66066209d2d587888042ff292ff65b3bbd46c2e1b7a702ed78d153df142aededa8811828f0b3
z5df87976a361c43bd8e3edac3667782092262e0e08688c31cbe54d11452f99a6eb3c6a6721f19d
zd65ff33f4eb51d5973bd46268f71cae2d51a09f8f6a378b1cf9c0f804885b15da7572f7cc3e35b
z2d2cd7cda63b0669bc40c331332a3bf0a544e4e344b4945056b2bc1e9fb4a4991bfe1915b52b07
zcfcdd8424e3b8220b09b37a7c389c5aa4316a32421cd3cc511537210810266b3625e91c3ecc665
z5c1fc7da6d74ad109bcda4f4142cf6a030405b24f74b5db6e0231723eefda30e52576353dd72ad
zda8984abec0fe7fc4d5b465085e712064c803b944399c8249a9fa95a9c10d14e87e52129bd0f95
z1d610650dcb86274f38ae733cf824190bb5231f7b564bcf6824c9ca72f785a407c8d3dabaa6937
zc43c8cffa70ca85e6c4da94e6646df87ea744cdb1aa49ed0e8a28b88d754edd5f639d1b12330ac
z98c3af93590895732cabe964135594b1332279b5ceb1d95ce2b7df2fa4091597bb663ea4101b21
z6f4b17460a3ab9b902aedf4df6a89228999878a74aebd30eb2ec54fffa70f419b5bbf5ef283a94
za5ca06722414f4888188e7a190068f7c287c0071e9c09005973fed4669843667d2d18ffdd28aa9
zf0adf5983e45f5953b6d093dcc935bb980f3c56369eb88658fb2b2d9e4cc331bf4860f949b9ecb
z4a0ba507b32218722097bed7dd7e2d0fc4a2053e76fda1e5092cd9b46930ff2f4ae6d587be7b0b
z84a42be8f8d49b37764f37fc51c6af9dd119f01f540efc85e8906e05f0ce72317b81625edc2a89
z6c93c51edbb1b70b050d1f5260e115e5bfe2e19048843cb80e2d908506af3a3210872959c477e2
z4e493029272a19286a9d4e075aa17a0fa437b362ae973f6bab6b106ce46a2c76a01ff31295e6f4
z5e986ae66c402139b0764cb5e4bb4cb7c800350e91c0a029f2bcd48d9d2622bdb09f5be075c2c1
z511ff63b77ee1b6762acea1713397585e7866c3b5ed364870d8f17ffb8a691222d9fbe6023582d
zca119503a0ef5beacde6c7f10e7a72bda5d9378570ee4e9254850c7cfc4a9ce293eb18f6b8deb4
zefa1726055dab9ae15605cdc07724a25c79ce24e53f28e1d90cb469e35ba15df4a7394e7be7ae4
z1d97b852e7689dbe4d725c6b77859bf86bae361b3b072f7730a0e814eb308e384049b4dbfee98b
zcba01a83364a0774dd27dcef0f6dc4e78a9c5d9d404bb45518278deaa23e36dddb8788c0c6b19a
z41c5c825fbe09c242cf8dcafc31212501ab39b751e91a57101ee3d564f4640260e2f9b68d67f5a
z24a44af0a51bcbb1e529f7dc0465f1799984253d3fb30f57190830b35c82a075bb7d55cb3eb70c
z17129dc4603b5851fa988e45a72ac63acb57107a5e0d45a8a5449dcf062c281ec966b46b7a2bb2
z08180a1c8a205c5a9da7ddec1ed401fad70bed78358e4f4d59e692fe77087b76d103bd2a465666
zdf4c6b3ef086663cc6abd08deacf2ec085f0f357fcf4e7f1cf05ed0cb242b3c18a9c41b3306a13
z6c39d29d289009d3a5ec0640c3bad4008bc73c439b51453e3a31be797a1fd953f670ac9445ce8b
zbc62cac0918e51d736c2a04beb973ee594d06f890d67fc5b351cd26b6fe2bd492f02677c8b4802
z35c119edf39e32cf9020659c15ad49d9e47b4716923da19a5103a49a5df86e775f812ff467e198
z24bfcab2ac1d29bb9d2f361cd23a15a1dda0166af89ef2f92aa2b25fa3c94177a366f1e9c05db6
z2db22b512fefb6ea2b8a4d4b502669bea8832ce01a217ba14f1649937af2c47a9d9c71222f95d8
z8c4007ca84f649bdc2077598741ef10029ce1b2aeb7b53a27afca253f92bd3de1c102b14c969e1
z33c07b82dec58708590e8dc801617b7a842297355e0f56d233789f6c2e14010d986606d2347f7f
z9554717d4954f29371ec92dec5703dd3985fc4f63a038ae9208d72065b212519803360fa6b671d
z9daee0140339ddce090c7305dd7e4b078836ac0f415100f7c1766ab92ea943e37310ac69a07bdc
z2481a9058330eccda7094363a321868406835c002c2196446fedf9d9bd985af211eeeb67c4fb12
z241c81eb1b2f166df8d9f85adaca0c21e189eb775fdb54989b34e7c8241b184719d02ae429049f
zb171f03a4e5418a06120696773d10328746388563991ed69ce5c0c8c867b0329273885ad1686b4
zc938cd1ac4b809660f2f9d7630e653682c9b9acb9a1277e94b114f44f86962609fe8d069f769bc
z362c1227fdf82363e2eec71e1d78150052fabc42f5814e31d152f24e244bfd97afe18f58c52cc1
z7bafa32d7262743c69a3c872aefb194e89f3f6a53b5d6ea513e1b5f6a8c519dabff1ea512e11d0
z4472e2ec65509837cbc50f12931bc60e0e1fb23580e8c131cfb60a0d2f03ea1e0887d437504985
z64f6826533101e123679eedc5a16cf51d3dd240dc787514bdb2d7b83a839f799fc240bfa687efd
z139f9f5ed79363159d324db02b823ef77c311f6595d04c8d2cb3aac6b2f79075e604686f318c82
z2950f850dba71500eabe9c7d4c17ffadcd8df1e1af21cc2eafa5e07c47fbd32f471968b30acb5e
z791981f7e8ffe5b9a8cc2743cc03230748244b603e14b38388ebe025b66091f7b7b84c26d84f39
z7b96ce40214426969c939cc5a6969840fbc0fd62953d5a8a1a561e43a08e451d2ea7ce3c16499a
ze8fab2824f9fbc486fb6f3b9dbe299c0bd32c7db97b0a7fadb1b961b16fc0095530c899989397d
zc5150b8751cbf1a83b621bd0693b49aeed8fc960a70c9a97cf8a169f2e93efdb9501832531555d
ze6e98f004b2de55ae73d8c843eca6e28cc5ab1aa1a4548c2e5660eea2f436d5721b565515f82f7
z16b9a53fb6f2fbc597f7ed336538bf6b5ecb05d060c94d1589ee2e7ba9d74c4d42d0722f96df12
z4962bf017a1da62c87e55e11abe5b6ff80dd7105f2f30880b44fd45509aaa3487471858b64016c
z1a7abe1ede783cddad5906bbbae64cad1ff825b00ee2ff60cf56a207907b037b75f9cc9b51112b
zc249bd534c53f17c458d9e5fd81b011dfe971086a72b85e3dd94a96ffb23aea78387bc308ef3c7
z73ef6eddc819bc8bc976d8f8585c88b54a59171eb8ae2ff81ff42440f2dab6b47fb44b0f48abab
z31d9b5713587fb6b199d2e13d2b25ac5a6bc844c12c0e4146481929b20704213bed1c3115c6fbc
z2a90290d292e2384d1a15f5d0210512723b5d9afe7b6295082ef7f312499afc4b2e07e93fcf5df
zdaa2101814dabf3efdb511633a7a678c84735a97fd741399c57a3ce7220bf0cb25a84fa437511c
z039dca908a5539ad809f23523b67d84ef31cbaa1b52b1a00d4d255b48f3d72ef14a54400851939
z0623f1989b3d902a529fac5464d3c201d1de606957e33a104450aceb8a2cf40a93ff39b8e75ea6
z887ee770f6cfda988a1405781646de152969ed5d7faa8e3a1b33415ae56e92d9344c12c3000708
zf0f721a0119014c55ca572a02bd95d11ccbb06f124d06c81be736faf570d9f95e9e8df566f932f
z57a6d87ebfbca8d7e2ac26f1ca5715f2bdf5afa98d8249043cb9f27a13e3eab17bcd3f0580856b
zfc1593856f4ad940bea6d220f7715863ac78b6b9547ddbf2d0d489e361fe803d28138cfecdfecd
z013a0f295144f4eeff644447248ccccbbe8c0d236eb971280c2a79cd587b2180cfda2c5736e523
z54bb6fae052b81153a98ca4cc0872b2f8ca74295180d4e6a7b60b336541742e053db8e166b5260
z255f87f21b2fd52b49e0c51dba7ef67e556ccc22b25aeb3e0d0333bf9517416a6039df97553f6d
zb1cb52c581059b2c878290d31a81a8e651c5276edfb2eeac20f7ef7c12447af7c0b099c48fe3d1
zde310e87b76bff2211474a74f794c1525a1cc8720b6260dd0a2596a87b43f426550a714dd32a94
z8eef9dcc388e1e15637de6e451832dfff2c342fa25c9360cc21b2c51938c21ed6e20c36ba7377c
z42747ffe86e4c937e59a04b11e797bbe6a797ccd84573f407dbc651f6dd1b9f4701b7daa394c75
zd5a0b6f3f7614e5ed0343b7000ddfd915e53f7e34fcbcbfac3b9b031ad4cd19b8018ae91732fb3
z76ea91a00e108e0fb4612a54421fe20dd0ccbf9c948906ce14eb7a74e87b2fd5bfa8c8b705cbb4
z1690d211007fabc89cccfb4a51443234e99a00f91d0d24474b593105a399f138568e5feb69c151
z526aeb5199a7a20d2476f2974f6cbde295d10dfc3211d5d61fd0f16815cfe36264cb35415d5f3c
z629ec5436f915f7bb44850328f347c9169463a526b7209707f7e665899e23aec11afb6bb31d479
z3c7507d98956ee707b9c26c5c89761ec0c76b4eeb28257f1d1fb2e46da106ef0b62e6437512df1
z765e3f96e050346de648c3f10e3b0ad5e5e33b4b062eb8a0a362f960fbf1dc30916bc7b76e3a5a
zf189ad2da562bed3d337440276f76592e042392b198834631828064e754ca19ccb18ca9c221cc0
z608ccf0d03328dde956f4b12da51fd95dcd6b52232b4a6e855d0624d0035449b5c868ee97997b3
zdc257affb1e5c0b7f737d36b252a4fd201c7dd8b83e4587676cc36bdb5d22b7ff609e66945727c
z67aaee855df1c5fa532bf7459398093304a5775c404fe1095330f9e41f3dc8c44cfcfe492d5dd7
z5dbed3a7970c62cad1d946058f59e7cbc73a2d7f4fca37539fb2e37486adb1f550c78c5db4b63e
z6fe68a9a273e547bcc00b4327bd1e9bac88c6e6c00c39f0c916e87a767e5c1f0b613e4831abd2f
z8ddb8105490f09ec307c10ff75bee8646eee97efd993123b89687d1c21ad549c3f26378488e59a
zbd309ae31702fce1a1797955000c645bb2997872bfc7e1784c971c004a1b06566418c0678cb49a
z53b290d91e50babab5e8775877219485ee0531e2f3dc17055e8a965af38c846cc44dbfe289526c
za503885cffd47b025830fd9e89264950e531ecbf66ec42bd2d2d71f08761a8b0f520aee0527303
zaf639debcbc6fad4f0f90fda7ab484ab7357a263a13c099f137ccab30f05fab08611786d033163
zd83cfd8b14b874d6fe83e1b2f35e0e2e3ce34010a85857728ff72a2184ab5dc292883217cd4752
z9f6de902fd12cd04ecef17980542f7bb49e9f5bc18e082bbdf4b9dc4b790ab71d866eff6b9d156
zaf1cf6f427efaebbdd9a59a3948a2a29ea375cc0b55b2c43775adf5b639ef91e2d2337794d8fec
z7907ae739d3926b8492c87e9386e62ec22ba429a1fd07699bcdb2bf6060dfe36e9deb23dbb4be7
zb9e3319b5fafdafc60649d4778272c9b50ccdc0d7deee09d789c5ecaa0aec5768304ef9125435d
z213fcd11d37ba6f22a240bf43cd8596a0191ddcc8d180f70d707c8e67237625d21e31c59c2a28d
zaa9faede73b9233654b4fe81bad50d7f6687f872e714928e13afd8e6ff504fc8d04ffa67ba36cf
ze9a708a19be190f92df11ba38bfe30bdfd47a1fd9d317bdb5dd0e3a25dea9a2cbc98c94f1c8485
ze44d8f6295eae2aa01a98f562a563c99cf57de22cb9fc94889c77ae065a1775dbfe7a355734685
zeefef862a2c618a2a1f56533f5547139d6d300ff0bdce46b9ba6f583b2bf0f70e91775a9b06858
zbdcd8e9537017c42f07b5dc2f73194b76b8029d53c04d7d89a26e9cf36ad4cb6f29b15fa08855c
z22b66b56cb493dee6cd5a28f431e8a3e7ee526f8e741cddd10f9c31a224043d24eeb0b56a0d7ec
z875f413d9360ef0157a5959c8b20945e45319d4b2558b27b60fac5e724ec5ad7644b0db1965cb2
zb0761b69ea81fc5ef6fbd048b3034717e95f533643359eb69ea2de4f917c7ab32ee7f15c79c428
ze2489dd7889015f680d1026826db848598d9bd6282832845d7052044d617e7464e058bc8a93e01
zb11d0861906930781abed6ceeeb495d9f9d9d4f59644cf4e56ed676afb959168be20431b45d1a3
z119c19f101c1b1fc7a0c0c3ba898785999fe80e89c48cafdcdd58cec2c1f589eee5425278510ba
ze196ea3d563b2ae85eb1a8787efb66c92b837f845985c82e947ac5e3be0ffb17dc228541747f67
z226b56f6293e3a568873390f0d9a1fca4087c3f58fa29bb43c0df6f141702d75780d79c722a953
z63cb5eb67999e55bce008f6d553c4da169e71d2e4ae94a74924ac1bf68acf0b403534daddc0344
z37cdeb0d2a68aaa55bbe71db70d40c61f6a88c34015ba111c0282a8ec56b505d00a8ab5d6dcd2f
za8883ab7d13f65ed21a29c34c6a74354fd54bc5ff0a7c428cca9d961e6ab9ac9bde1cc0901218a
z65f719a3066943b4a0e389b77c13c07aa2c7f7658141a61a4efa33f4a2ac4f3b4135b032179ed5
z2da93f640c36633d1ebbc6ff31a4c902efeb0b239cf7a37131e5738698fd89806ad66991713b0b
z0e4aee7f3c37532048fd32c7b2f2ae2f91f62157f8cf2e5269b64b2186e0a09a3e97118d640eec
z47e124746e0fc5c2c5cb575ff10121b2fd82ccc3f68bf1ef176993e657653f4909ed4237bdf107
z6bda6ff40635ae37374a09b650279d9f5a825b8fbad5397ad57081bf8ccd7b06b46be414a4b966
z064c4450d0fd8cd4e721072b2de2b42118274beeb3accf4241465e02200337aa98ad6ec931a762
z5e8f495376c9c5c9c06e76235c6c1a32e94f246f2d1e7dafa82634a727cdf913b71e06ff7b968a
zce36c651b0c6e8d3c22e8967bbfb30cb39de9bab2b8ec6bbed728902087c24d8c4868e61d73d55
z5b345cee3560802ffe36d707669f64ce2d4bbb85f1c2ec4dd15b133f13d64303cb3bf1abbd9afb
z97c3164a0ef38f4d87568c6c439adf2ce834bd9cfb50b6a670c63ca7f039b1d2cb20931b659b2b
zec7019e135cde72c4664a7c72a987a25f2bd9ae913f30a8a792fb2d351a201bcf4882a39d892df
za031c8332d42699c069a8ae7f8739a0c12b74264836111540e29738b0e91a62601bcf256b2f48a
z9b25703f9a4cc257530cd5e9106c24dacb010dbab2e860428a754fbce3cd311bb4f6330636b66e
z588d36180328a4121ed773b9027d90e0de084c739ae2bca3e2d4b0666f1022c2d869d4d99cf04e
zf6f5b5602586f72898e297856ee26e0e5773b80f191481e32732fc7587b229dc370712b36756ee
za4bd2ae5bb1511e83a9a9ac7ac0e851739545d64c83d6651bdfa9d6dbc2abfc10e11b769785650
zcbec96d42df0863e5babd513f75f74ff2f4f0ae4ca1ea25b298391d85aae6f9f986639ed8ec40d
z1b91ebba8e93a050d5042f35d84de30e8991bbdb531e01f4113aa984736b4fb5cb8b3ee0f28d8a
z4838bc65197602773880d70ca0beb5db0788e052ef11ee28d9741f5905688e4412e6861760446e
z25e49aa7187f9f480b32ba81baa6d2bcc0c9659f9283a6d52fdc9a581765319980daf278e9718a
z92ed2950e265a5228e8d29b2b95124ba0ee194180636a751823fdc437fca3e349c8edef4c4f546
z3dabec0c2b3001d1214a0e0d25407a2df09f15a9c66b069d75abf1e315428ca4ba65794afa9cab
z529c7d44562d92e7c9e8e25dab19b39003caeb846370d6debd1187d1fda01bb6d790f1bbbffc8c
z6228eb8b2c6af04951896e86896115220c2d53f3c0373a77290c08f9edce717821b19380d1e704
zfeb462305adc46c91e9a9d54468faea617ed161f1524e95e1eb34d7d03fbd29a8fae5ce242ea3c
z5bd72ac52fa795a944f6c8705f4e0a5d1375f5916077747f9b5254d585457c07b9cf3a30ef9136
z001d36456c77b0909860a7d350da7f6f4923a4e5e86f3ee188afd313c25f6a58475c5e98f50b56
zb0ceaff38ae22d9daaec3f80bd43b0a11e466d36fd65fc99ea6d4e10ac659980560931ff219554
zec054f69332961f6d3d07bc40fc9f896013f6817aa485bee8c73ebb36bbfb4a3c4dd98bde95511
z2799e7ebae68be506614945e16c9946e5eec88e8a7f284e65a296f4be61373865a484021d3551c
z9b43bc11f5d09501be8f82085e59a4566427d5a6541dc9ed3176ee42243faf6fde1b49fa2619bf
zfefab29a16c667a3c9d89b23402b46a9542310d507811968586dc96c679eb5cc20704ed1730d18
z4c547ab56043f2853cc7cc26002c5e1648dcd371934681f833ccbd07030706de6efd49dab073b6
zf81a80bda7c95d85a404a8ff79290bd3e503531b28f48a6f0eec4500d8605b75a90539b21efe5b
z0b68615d3dc24d40df41e4f610f3f7f43daec48cc75929a914bd5320303d748ee06f13b5680d63
z50ec009067f7207e5461a5766c48b554198607013289b3c03e0b2aad1a5d665f20e2b84fe314fc
zc013c7ae79f3de34ca89d2fef6630da262c8776d412d272e1ffc2661b0c67c906b732fb08c517f
zbb6709a8fc56803049fe86081906d06b8fd6bbe8c6ecc1099650b11b8cc95f66cd15602a635616
z57036f846453249d50fcd93ef37117f45752d2461a75edd3cbac040e55895b58d91898945a2136
zd08fd9cbcf9988463c8be43af371918c5b024aa7399e0ba4b3f892672817427aa030ed56e3402f
zc41dc2ae826d20fb64799e1fbf82c02b9e8f7df6d00d721cb1f336e82cc158294b12e3dcdca33f
z9ce29d52beeb0d244bfae7c4d05363256659ca41559667381f05a3a16511d7735d2ac5eb420f78
z9acb64801b00160ad2a3fd303999809d8547c86b85f62a232e236218f812a3ea967da2631b2295
z1dfd85ed0dd702f90c53530308c3c85bd99a55f9802737d4bd1261ef4a94e48e2c978cbb38e82f
z4d94f4430bf837dd2b700b2370fc42aa511a28d018ee3a24aa449a686feacd811244b70ee47edb
zf150faa8fea5f0d3a4bef4b0997ec3af4e7a94eeef7a0a6bead7906ac41f0f9c32639038ba19a7
z9d9104716206e94488c83c821d991ae299a29877fa6745d449d95c9faa1b17b6dbbf8c7d2b6832
z3361968b07db17a2a36dcb26848d25cc235c7d7ebe27674ede5c1cc838a221ae553ff0bdc94542
zb48342cce820fe26362d5a26239f14d048258e82e73f55ef16aa907b6800f33c261e2b6e68ce5b
z3934afb311d39d480a65ed8342c5115557ad18bc6e3b07bae7786f501e262011fb000c0343c155
z6e5b4de0b3de86977286a4609a42332e032294b702be2bfd495d5839ecef50261c30a5cae1faaa
zc7ab095c7320625a9fc1c9d25835e3cdd0fd4460c681c4f4ea0c48958a3e2eafa7fbebe44f6263
z00504072734ddaaa24f3b0dfb8592824c38eedff04ac1bdf9fbd99aa63fac8b796144375676d94
zef0fa90c373d15c61ba25e432aef0f42dd9819de0c994a79af80eef497a733743b8a02f457f3c3
z6003d4ad53f596222e0249217ae1c55642ebde2d5be7d38ee9f7125b10fc1a4987160454f2cc7b
z01ce07ab051ec6e296e68019c5b4af06e40af02b5d7a222a134dff4061e5ebec5cc5f56d9d9030
za5daf77ae77437c995541de71f69827a5abd88b7c8e5a8b3303ce9522756bd6e96337906aaa4f3
z52b9f85e5b3cd5c168ae94fa1a96a6ce84f3be889c45b8ab42b8969ee52bf27f5e37cc465b4742
zd651cf9b7355df9568bba73861a51c76d4a6b18b1dba89e83f499360874d2cd8ff12f8bdcfa8ce
ze789cc08952e5c4ecacaed50cff13c442a8a7fb25ed128f28c7ed18059b30018aa10484189cce2
z5c06b714af9297fbeafbde976827e73ea63aa775b48daebcaf2b4c1179a7ef9ef11ebaa12a5d56
za4ed77ee9f76e838c900b9ee42b2e2802b0c3b561bff87a9259b2c40134e8aaac216bddeda771e
zaf465545c7bba7440bf4bd622e8a08debb610a42b46b1bb0bb20d9247da286ad3e1e54db8a642d
zd3a693564bb3945fc1530536cc1e5821c9818b5393331f47c50d9cd984b1788bd8129eb091ee93
zcff373bf7f0114047758ded44752cc5c23b039e3fec4cef5584d96bb2daaf49f8f42ee80f2ff3a
z6763dd3e71778602d694ed56b928e4a9d17ae2bafe7462b1b1ef00473b980f57bf8d4dcff77d34
z340d41b025a39389db2ce107b62567a5b22a6237b1569a937c5447300803c37799d139d38ef4a3
z34485a725e47cc41d305ca33b14699d4bd617466f586ba16b5a0b9c8d7dd34fc64cfe9c5d0d8bb
zf90c66c3f2376f6d512c4d34a7fe11a02cc8c141fa15b55ea0d8cb9024deaf9a318f8ec5c90433
z6c6afb091c2a684abffb9d48b7895cf4aad8bdfa99c0d7301a68a5eef9e7ecd493f4b384397c93
z6788e3b96500532271d1055ab562197416b0bbf8630585d282350d7355200b31b340bf1ccf85d9
zecf716f6d0c11666009dd741114b6f9f7144ae8331cf6ecdc8ec24f53c3a5dba78c1e5e7bcbe0e
z2439fee4d30b5c6402e4712e8e06b82650e08f014813d795f813e44cb6c6356bcf06c6c5c3049b
zd33d830670d9bbace6f78922401aec1fedda91f7dffd7d53c1e2e3757eecaff6c9f1b9f2c38ac5
z8bfe13901b8f1b3ae35474607a3c5f0220c81df43fa6d530858ff028d8c0c8402c646b978e295d
z5eaac9f067309196067db118d78dd3b9440bc9c1e02fb2518330e78a81d2de2e2ed903c268e66a
zae5ba811bbd0e8d89711d1eecce2b8c83f4f5a2d1b455af25101594a8fb7811a14fa0d64d4c93d
zc1d9a22a190a2f98d47d66025e4e92ccd51f7bfe49e5a47bcb63c20716487e08aba5ba937dbbc1
z26923e774ae191d881f03b7b6efec65c091f11f7793664178cf0fe023cd3dbc1c6f1e156142fb6
zfc05a79da344507129e4a82061d075b570b59c4de6546ba645c8344168a509591ca3128ac26762
zc873ba3706b46adfc99bf045cdd6a3555c8de9b7d27bd03188a51ff8547e0b6cf167f1a4cf9637
zb77551dd8e25672e2259ad3d79b9dc1db1e4bf9bc36be61b8980b75f29f0d9ef91e22c30b4bca0
z78be4b2bc2ae452e029232cce4aac1cc6906f17085980057c1d680b4cffb7fb278c21ecd85e81c
z5af103e39c8ed37b392a3801bab8e88e3bad76bf540e746551726d215c5b6585e776edfd52e94a
z3210e7ee04b3b2fef9b4c5fe93d455c87c3f893601f5c856dd95f3836dfd635fc370520f8a652f
z98474a9c21f2b9e4207ec22bc5f4fe475aadd4ccd1c26af571360a742033008c6ecf8a7298400b
z8568077dbfa940988908247611580527d878336ea166029712c4ce0785751ebbf82456410e678f
z964a540551c0cb300e94b8891a6ca654e7522ba1fc5e8ca57df4145d59f6a7e2377a9c81654780
z826455c8d8808b9b5ffa303757baf30dc1801fdd73bfa0c9018143295169fa2848dcf823a52a8d
z1e32c0df09adc7c22f9a76a9b4ef0235631a0a9f3d92e886ce9e9e1905c45611d9a748f7749e82
z56beac99220bf651ecd71dd0eaf2777f970a7017b36c71a693782b8d66914e5ec7fd6bf083a6d8
ze1d4c03bd2bd28ac023b3036fbd8377f11c505a110e08b795f7a3e1f92d15523f14dfce4c72434
z49fc606eeded88217de25e30adf49fff97b9fc4768a0dc3b103782f14dc6b4f5d4431e5bdffa04
zd7fb35563fe1ed27928ff3aa5e0fce70580b171faab55c60e2ece8a35e88053ad88d9c98ffa366
zfc2bad999ed405ad6ba34681aa6b3940dd580fb05c3fe80e327d2d080d7fd30fba7bfe4fd46648
zb209fe720146809c3aa210c9f9c1622dfcfbb2679dc79e50dc721f1563803b956195443fddffa9
z80d02cfc5f73b48839eac9ac84f2dc532f90745154eaaef47348b91fcc94ef4237bb2001f21b4e
z08d81829f2cb4782b9bdd84abc4d6e68456dc956d5d1313fb04aa5497599601c1466c9251d517d
zcbccf7569e15df003451e4fee47acffa294878655f92b4a8106b2586481f6a7916b5ae20e00018
z3dee84dddde42c89090ec05d6046c724a7cbd5cdc6faea530e751b12c71d4945bb495eccc79cf9
zf4395990187d557d6310d5bd13ce757d4254b1dc6aacc9e973a32bddd765a4b6edeb8d7b4c91db
z6675900e5f7b2a4983096f39a9ad2f6440242e84ee54952276db0bf9313f9d388e956d9f646df7
z7750d9f9d04b199fd924485ba2e72f2dbd6c5a4882258e6bd88d9b1de19353b1abe518cb3b02bf
z320c1a64d060d2488faab6e29408ee94b1a2c43f9b806bcb83a66a622cd5f3cb2eeb60a9a292c5
z8c9882041d3a6a0b68892c3c4a63fd2d55b2feca22ce7fe05bac93f9189709acc1e84cb17fc6bc
z05c9664857dfd75c8df8a0ebd5f888e058feab1308f79c3d2c8b2e03151f4386f48096367751a7
zf15157af39a81a8f1373149ac6ab621bbbefc42e949654d20b0774dc38e193fe5cf077fec11f7a
z92f5499fdc29cefd0707efe95cef0de3b2a404262981ca3bf51655c7ead05c890cbf476f500f87
zc5e848b45ac219120c190a52bda69f3a71cf974857185025f771e37e2a2028848a18d805916770
z0d92cf5619c563d16a2ff47ed13321940ca1edb0a8cf33c6a9b73de0709e0f22c034186793822d
z9db47ebcbd6bc7d5e877a1a739442cc26f702d52ca5647ec44685064e00b59c0e503cfa6566de3
z1de4be73dbe6e78cad5b9a7795cbbb93bb0a87e9bb99dd8e3c90c6f9e2f3a3c09a30191153d2ae
zb768acbfe38dc5742b388594e3acbd55d2d1a094d0c711905d6befdc4239aede02e076c06d4bf7
zf7c129ce420070c7b10e1c94d3407fbf7e21405b34cf44a6d0d0f8c2ca1c2bed7d09e1aa097976
z6f56cc9c7a009df9cbdbc34159f4a93fff0f41b9bba4f39c349910f573f353b917295fc07ebbb1
z54bcbe53255cf94526baadf7826cf300d610a3e87ec3e80e4997ab298ef69797525bbf8c09fa7d
zd7ef21a70c3ef33cbaa09b3261d051b2326710dcdccc8e0f915e390830be235328e2c699dc30ab
zfff387d97b14c09eae9227facfcd90dbd2a46b7110f9f4487cc7f6cbe4d3ce1b0dbc39ff4ae315
z2d690781c10c6cba1983171ef303959656e00a0a8a4b7746b2178a241c52c9fdb1aef7eaf988fd
zc0e05700785c5b6adfa5d96fba22cf46757ce83b76d2182a2538bcdda9f117700618019bfd6723
zba25769f5e064721f1365d652087dc0a3c586d26f30f80767cd43b18c61132467dafb867cd8d29
ze631500f131159eb00a4fef636e2919684fb8d2da43804d3f8f28945cd010faf902d11fb06f74f
z79ce637dbb041d0c51cfa0938a6e1d5d0c1ef20d793329cb207a951998b6fab14543238a976956
zf90ffb119a010213479fb6211a517c386927ea7a42c1d48bb3ab35d2655df2150adc01f14ac444
zd3867960fecac2f7f7807199e6556bc8cc37782641f9e010e1c4f781668dca4b06c7eb0a831d45
z381fc9b4b2286343af35a18e5ac0068dff41c9dd7bf7e6c29c67c3c17488415f9e33f7fa1efa6f
z52e20a221b6f37197c613ac13e17642be414442ab4957b5e39f8d269b1b0a37f1c2233cbcf854e
z4d8b9e4942c378610d426ec29d8df05c3889df3e3f9468917f86c8a99d05dfe6d91891f4d8300d
zaaaee2627cfe117d455872638947c81ec224664ddfd91a3bd467d436fb16e91f98348274d6d85d
z97417ce70e675b7ce8d682b7d305e17fe561d8e7ff32786de4e771bac71a57341fa1f110adddad
z5ad629452883fa5ccff4540c4bbaa6d368425ce6e5d9dcdeb807f7ce3e8f59dcb584e8a266cac7
zfdd5368fc68bbde0a49094c9c697fe32894a203f03087abf18ac9adf40d218a4ada453d5a3d4af
z53cd5fd36a81c1e75848d0ffa5f9859e1914857508d39a57e9e9a815f7fcac532c14862569604f
z3ea57bfa0d7d4a48d69259ce671b825052722b3409a7fa822afab1ec4e1da746cf44a2a19216b5
z7cc9dee61a79b0fdc03b4abdb9b15c3da316b925b17919ce24fb625a6da831be0b207a418fad62
z6b0b5d18579265fc03032ed4266dad9818fb25aa2a9db79c1a9b6b0f5ce5bac4365c9522755342
z7621c138db5aa65d759abe98a97b2e56e79ebaef7634ff7364a6b2ba60fb66ecba1f1980bf4fa1
z24be16b12e4e9faa50dec893306a4290497a7c6de00fbe6c2e2a81b357e9723db088126aca34e2
z6059d2238e98625d8aa046ecec3312b6e3715f972a07cc5e9021ccc88a65433e06b6a1b49cc13c
z0c1b1b17072fb30d87368aec32f3759c23c54acd2fba6daf8ffca0361f720ac0b1c066481a0dbe
zcfaf2b19c955104aab73e4523f930d1b3ff0b06677e8f33dbc97738b16d29fccbde450f5a48d43
z5106b20bc497fd13711fcf37e467e686497ae53cffc6d877e42a5353b97c90281c17dd6b34e144
z64929bfa1bc8f4ab87f9eb245d05b3fe4955da5c6ab1e026375ae2918daaa7650f6cc2465fa3c2
z1eddd66d4b4ed53d07e6e83f1d367d37cd8e499bfe8e13c58b901101021d3c0937c7d5e690fb9a
z28588efb9566b71a1c28fcde34f22cb7fbf3dcd6da014235faa83ef02fa420e65839d87602a154
z3fced59e670ff27987859461f17f6c21c6e77629ba6d64175f165b8cc15fa3567a6eaba459fc18
zebddfbc22ac04761e2961b57491ce007317e17151d0625d60687407c557ed0dd914cf2b9adf81c
zf92ec960b1c6f401692d028a7df3ad8e9658f9371a6c0db54055a2b92466aad158262794b8ec73
zbcbfd51260021e12a2872d96f9059237431a410ae67ca7539289090e313fcb0c258eae33d8f24b
z9d5d8eac4868d61dc18e9c610524afadd40032e47b2390949050d5aedd2ecc57d5f9c06de007b2
zec353eb2acd065b0919fca92ac348e377eb662e9abd0c9c975572c05f426e83372849c0c081453
z5060f3d1b1d72f749854b0e999da589083d3d1057b1aa48d042056a27393d271a0d0b6a69bd893
z37dc12c81c539af3d232a1eb6a92062501aee57d3d8ea54d16dbb0e318f8096747f9f513792c98
z2b7b3a6cdf42b6fea74ef8ec6fa29cb2f5173fae7a866c5c167542e1fe5d00247f5ba8c067f460
zf7f4bd1e4b029400ee225fa42a65f6af357bd74ff0143d49b2b9707390243761163ffffac29124
z16e209774c37b628fee9af69353a73a11edb07a4c66be9936218153b4c43e997e867f830ab78b1
z5273d268c766dacebfe8f769f22a1142f934694a14a3e799cb39e459c58bcac44070db245c28d4
z09f0c557325e379a2f3920350a0ced01e0ce967a379d8fdcdc8e052993593169e6b1c692fee7b4
zc2e4522ee6598f8df60f0eb998fb4e59da795489e30f9ebb27d04b7c5b42616e313ab7120d5ef5
z2f228ca37851ea219e859863561a26e47dc2024348217df54c42ff0d3b836a74bbd9eba163d411
zffe4214099bb3486c0deac17d8c493c9167dbdbf777941ee58c12a845c7d5695f3c10fb5c03efb
z8bd873154b96e87b2052864c7357a0bded8b030bd63cd748787ce1bacab5b0506b2707d9cfcd04
ze714c50fb86aff51f4afa8ce9e106895be59132447744f74ae081115d6c4763d32397642c65239
ze761c1d6833e245b08487ec93b59927c1c2021817f8aa616d171dbe5c3643fa0eee9aae518864c
z2e453356c32e9005cbd83d2e24b8f62179bb65a1d5ef8bcbafc8e61a11aafbbfe613064dc979b8
z210b225c3fe50018b1b21d9f2814416ddfdb0fbde01388a3391ab0c9a0a073592777a9373400bc
zecde1dc994f4be97fbb17b73d24d26cc9052c56fa284394d8338a705310855f0ea9b04dce879bb
z412f7b5cb05f11b186e2758286497813dee86052c43a5a398a95a0e57c133570f8e165c27a192b
z87e57c8ac5da6e8fdaf281e7491f3ed0712b6e3cb4b97c123c8e0c8c98cdd0a5e8abc054e7c85c
zced96a10380fa0597df553e27f7800a0918ec5a3d35dbdb497ee1f2052172993c8df14c3ac96f8
z19dd94f7b175e10362c5dd9cb62292eb4687352714c54f0bff2c7905e96c999af53d43df9bf9d1
zf6a7903f2e7dbb02e8a5a4effa6e9239d1f9e77994ef6bb1a26565df1fae15aa48bd372ecd900c
z5c5d234a985d4f1b98b08ed54bc782e0505c9df31efbf7b4f0c3176213241d23aef3a3a2ebc102
z6828f5ee4d47a3c6ea74164eb7e52f0588fab542b7c21078762612c8b36004b5f3b27355d09ca9
z986c9c0a3321296ab84193fd74d895cb4540aa3162a8db3c2693ee3a9651f60ba82c509d0ae669
z9924cdfa0d1bdc3a9f10c4dda15e85d963ab59d8e6274643228b751f32d85fefde39e0dd8567e9
z73be1ba4bd1a53a2a188602fd09dc616551eefab4ecdd2cd9f2dee6ba183e9535606e0cc3be8af
zb026317a547b3c5de82c8e15db0995b3f676086c304fe8d7634f9d605682ca031bbf8621dc7687
zb81d2df53a8fb0a6294b249f0405d0852aefe56e506ed87d735f331133d359ce8c16e70298925a
ze6b97d0ae3d882006279c8d009687deeb678b1f2d95035f8f9ef40772e22cd49a0d5f871bbe626
z435a894fe0db7ded6d1d1decc4f738aa12010051477df95289c6184e32a4433c1e48ca31b12e05
zad0d726142d6691d77a2d8f202b416ebe5b1ec6506076a3241956b91debcadc2cc71013f637f53
z5dea2314cf8e154ef1b84d0467c656542c56c479a6a8a0e0e15c050faa4ea4cb876abb9d8ad4fa
ze8978659bab2ba404158ad8aeb0c53af6ba4a0dce446ba09fd8a84334be445a50c29619accd80a
z7c4bf838f98359a68a4519d67856450db6dcb7bb85ce4fcfb7296896bcf11d4729da1ff9a75658
zca0bf6eef05bd4b4a8fe0d449f40f45edd503175777d04e69d00b8a2e8a8c15dc9d4d062e975b5
z150bbeb18e420298e68d40c6d0478b9504150e4cd6dbd86af10a146a0cd20cf9a8b53b89c15661
z0a9e7785584c6f4528536ba597b6a93db33b6520d835b2cecce3ea2a760e59bef962719b37f7e6
z6fffc37fab920e507d27dd096635497f7597fbe69824f334e72b65d721e8fdf8dcb0a80b791351
z81003c1069363b68cacb0f25d623f75bbcbeac6f866608716789b8dede214f1bf24a03bd29717d
zb04c1ce60e05b0505eb3e5e628a3f67eed182f93f3d6117cafbac24963c19a68870deb45249442
z25d28297a423a0a48ee7ed5cbf7457a10091da65ccdbb0fdfe432d83baae60e0ef54530e2eb4c2
z333b4ae84ddad4ca61183d81665245c63647acf1c19db9150ce95b2431703705962558cf20d8e7
z4537cc3aa999c7ccda9a8117596477385b5a469a4be98f5dc899e4554863eca62577a3c637271c
z401540882e7229a0a18dae545739b08e9e56dd236f69bbadc9cd634d58ba1223d075329c2e1755
zddd55b4077b7ef38dfbfa6c01ea503ad0a0c981a09083ba5a3d7ebd288e04eee0024b05b9089cd
z14c2384e68067413bb7fdfdb3bf25b49e01b32b4f1703a3cfbf5a084e307db250805bcf671ebae
z61be1e991816710026eeb38a3d79e30713fe905756573ac028f64a11532a1e15434a077f82fca8
z7538bceedd81bf759e76eb927efecf3b87598c73006a46ba71f74df325d00b69cb211bbdbcde83
z6552210228ced6af6feaf6706c0d44beedf055293d9dedfdd711182e75ea1064473bf2d998be7d
z4bd4e87bcaa23d2747eb4d41df5c70a052afc51c2c7a334be2b0caecf86a828d6645f28377c4cf
ze2e07f5e3d7f795308f941abdce1dd42062955f7ecff0e5f18c4aeee9131835d03e99de33585fd
z2d5f37ad8355f214db053cc56a3d2597df7d90524f982adba16306d228575605d161acf0728056
z6074677d832646bc26864bdb285170a6e88bb823d4d6e078365f87e85970a8a67bc1eeb70a82ba
zfbefef17829e329b595877259d133e84e1aafc9c1bb9479fc97e7c34d372eb2ed9c8675a18f1b1
z5fb66d91fd69b8f86f310d114b318223f092170357ae6f27a1fbfa957347764b53ee6d5e407816
z46f8dfac368e343e70a011de4f706e765ad1136a729e843a2f879b0b24b13c297796fda22b9400
z1e34ea3f65af1c4586628e58ed6e55015a533203164846f24c96ab0caac8049e4213f77be7fb20
z1d0bd74dccf7d1c0ed0ff09ca016be2c6c5e0588f8afefc5170a9383e0593acbfbcbfd3560faa8
zc734075429265306a0bdce3d3d347535a09b9ef1d51e27cba6e651fb546702dd751e521cb7f0c8
zb0a1f02e212d024933c2d4a9d673d4608819cae34cd740328a1132c89823eb3b4ad52732a6094a
z62905896683d91491697ef9f76b623e2920e3da92b8a8eb48ea7a96b3463bdf29c3114c57c1e19
z847bc175f50751eef4e98e9be42b71eea62a18f40f406282a3975284eca04bddd5871ff6ece70f
z60d77f105d708d712e4e0884ab4c4db5a6a9a7e85a17c8e44032657673236d62bfa159bcce1090
z9fe1b83ca254a504d5c2e76e1eebc93dee5b9e27e3c4d8e4889ff4073e07626b6df1ad0cda99d6
z6415a913fcfc94ffcecda23c7d8d84881b11ec78c5ea736a45617368866395d9b58afa90da1b97
zbffc712678b294cea6686af0e24e1d6578eb800b356387c600b67ad2d64267bb885ebcebace8dd
z61ce108a603aad6694efad30df620be1cce04a12c6505a7ea60acb054060fbd2ee0e6af2baca3d
z264657ba7a8754eedf3ef2d2916eed7850911eaca48a71289c3ac2d62b66df91c301e60eb60a11
zbcaa62dad4d4d9e864cb92f2c8c6778013d2e533d7e647c57e49f9d3c59960d876f44c7a5f0754
zb5b46cece28ba0699eea7a7ad6c517e5a01ce7a89b4e51a02ba1803a50494810dcaa5219e4699c
zc524be6221fceee40c54a2b6cdbc5a4055b64624d6e9faceadae1d6779ee36b5b0ca7f44ced042
z88b81ba15160736461591c0996186d89474c9e89090861e812de935ace5355b24b9d3a8b22df4a
z34f1e825279b48c75745542d961e2c76515b2098e8897c5c121eec1cf1391c5f9fc1762ed65af3
z147e5f00c78628aebfaaab6cb42a7d4273005f213e4c6744727c088892f0b80f2ec1a3c0f081a1
z3c1da98ac6ef01698f0352989a47d380014ab9fc62736e7d798d078a6e65d10c15c9afa79bdd43
z289ceeb2c03f62383633c701b796cf4acbcfc5ed4939b3f55eebbea39c1f939ca3a8087a5aca5a
z1f3579f74755130977e7442d027e11aeea1bc1e90aa5091b88790e164889f6e8b8775799650ecf
z2928e23426fc932c32d57df99c009f3ae7b8a35ce45a92f37fac9d068c5699e5c702c2ee13e57e
z1be0a77146d31efde5168d26dda5b79aef6a734024e6f7aa95d4a5874aca45133bf53445f0058f
z018440dab5c0b486efac14c7c3e3f3025896e290fb1b04bee1b9076df1b597952b0ea8ba1c874d
z84a476aeb9d872c007b2730c96b0d73f182bbde2f52e5c3642ece84b2b868246a5d8acfc0c55ff
za42f6f195bdc821aaad8015dbf911d1c5e1fc1e99833b4e1ce7001caf438876adae60b20bee79c
zd99c27dc096ddd51d46e373a59ad971e1998aacd58b18abd1494deddaac2586a4447278325c82c
z387ce6601ceb360c4997038cbe3abbd96b44d2118d4348033979a8b255c0189f639ffd7013f175
zfed63b159a28b0259e558fdf7c8720d2bd25a38ff30f34fe2d4676792803111bf846a1fa29166e
z354b31c7c39ef12c6a86c7a94c4786a9d2630037e266ca80e970d292acc6dd6cfeeba8d406a146
z3a6c966b16dbf1b085a6fde794cf967d32fb955570bff26c12603e31adf59dc287b9940f7f1afb
z8b9e9e13a83d90081859152e9b9763389876b3fc4589933eefbda1531a6673ad7f7c79a497cfcb
z7f286bb04856f3f849e36b5ec7feb2eb88b106797726fe1756beb4514697b6cb31d97ac03935b2
zf3be5a9a91d734f2d73859cd02d9fd004226c53ac45ba6addd8421c8f667c1186b75dea86ac069
zbe953ad0e5ef84c591a28f18e3d2572c6f242d289147a539a42bcac5bede78ab43981d063e49f5
z0d04603c6a24a135d4e9e6fae002726480ae344cffc95b7b1eb0cec8492b4b4a1a5b54f42a73f4
zab8ac44f819fe2e223a8cac4a3f93936d172effb9479e5479773b669042dab7b0e99d02ecc503d
z871c85730678dea56b6e0a30cdbdcd5d29a52f028b0e9d734b48ac7cef1a2c2c2f79769ebd0e8e
zb50bda4e7f54e749688fc910a8fecdd6a7dd7bebb61c51a25e3ab8e9393c780364109769168dcb
z3cee19b9528eb59482c33e871c23b5cf3ee6eda76158ecb53d16bc050e57d287237f4bb6817e0f
zefd6ab995db8d0d2e01dcd8407f0d3179451d8b070fc794709f7fd38d4089853fb1ed2a8ed82a7
z1580b75109f2670ca066b9c298527a1103bd7191145080389b8c98da21299fb62563a7883c1935
z4f93a65f2a15d0e3389afedb8183f2c37d33fbe7e4158ab47e5e7feffdb07994efd2d708b1a7af
zf4a3eb0b40f1337d69088f5383ae7ae5389dd624526317541c83b277f06bd668084490b6388d6e
z073e5ef2197a4294ac2d2c2aaca5f41ccea606d0b0ada5be57b6d49a1af9945c1b33d9d763bb16
z4ce4713fa98807fa5b1d84f57f0415cb9ee51b417a0fd98935d66007f87dccfcf7f23e72eba99e
zc759327ae8d38697b136b0f9201288ce463b9695458168442b493286515b0bb521e7e3249db864
zbb897fafbbbea0ae2c14fc4330de0c2b28633b8fbd65f8e371351246789c1f428f36204d95f1a1
zafd0dd03cbec66bb3c5b19e35c7060b436d8aa2ff72a2e70106c7d659d722e15e41c6ebbd6f4e6
z7b60ec134732bcf321af5f0e53bd2847a4abcec35cc34e074b288a217064366738816f70fe38f9
z49e49eddb8d5c6e00e8848ec8d5c166d9bacea2206b87c80f58b32168f19997303317b4d18c36e
z95fe95e732c743b669617e251526e3268b0583cd7e02977dc421248491eecac0adef336d14a038
z6add225f8854401e8fefdef9c7f914e6c2caf0ad26bcfdc9e247a5c8f0ffce98dc6c57a2c3c98b
z2355925c5c10ba108843e0fe9175d398ccd8b3324020aed95e3c65cc646d2480db34bafc6f2617
z84b04f4016ad4e873be0a383ab40da22639b83c89324b65104ef4eb36d398e68363da384013506
zdd4c2c8a0f8783ff8244d9102007e76bb27a961e1257571d0f6c9f1d8fce10541fa5c4594ca520
z855c8f34b88d0eedcbf925ed8e469a6064dd5d67484cdb942eb00c4255b3846a820a01ada4d553
z40127beaca3638a96313452c21219c9e475c722b439bf565bb29157ad49dc40b0fe214810dce14
z4c1d45b2c30825a08e7807183d657131525c513331cc85fffd22352e179d8c5027d18628a39f30
z066d27977d7f15e059a230a83ac1e77d67ee32b71c5e490b5bf024ef2dafb855d7015b26a9b02e
z5ae3a53c22c657f6481c57e80aca33257ed1164bd749001051531deeaafd3ed6006aa2495b9afb
z3b3a82cc4862f2a19f1649cf4526cae12707b290e725fbccfbb85e19bd8e57b381bcabfaa44ce7
zcfbe4c3b549733d33e8134fc1258387236ecf2b01de616f6d83cfb7add0d7c5cd35b2dfb3e748c
zd89a4280d7d5e79272f2f676614000565d0fd03a92c20571655d0ab0cae7e6a81cc595917e4864
z781ed010485f672ac72d9088039f855073d7b63fd3c1c618a34e79d3d9e09093d116ef7536c3fe
zef5e3f3c268bc4b489f4c533320e3fa9a8b7bc9b56edd09a2f31ed161e36a9589077b23daeec37
z6d8ac5e83f9b73f724f6393cec74715d5aa1db9a33bb4a1351ee35e33374e99cb29824731ce90d
zf86d735626de09a09d5d25787b90d47b2bfc03ea02a0ad583f166849ae8c0a9261172715c4a616
z61868216ba00d2333bbcfc56e968a893292b6d98742a0dec687af5ae72843641d9d276681781f2
z9bb427da42c23972bdd1f5a30c0f065c619fcf917b467362bb9142058c710bf59964cbe266dcec
zd57a4a089a536ed839bdc806210640e24548f3af625c2213bc055634aedd667f8f16edfeb4f374
z92f305611e70b73c6c4d9e3c9f050fdf7a160117125955fef53303cc5df0324384249b5b0a93fd
z1db6c7660f4ce44f7952317cc451dc33def8ab9a1b7f6ccbc204a67a3616efa79cfc9430e9f137
zec17f9b2540f831c5c927ecdc00d09d68d377ed784c5a06a784ec0a81746ff66534f5f91014f12
z5d1ff9307b1177fa6e8297999457646e2ccb3e66f1d60b8fad1f90cbbd41e9af60c0254f17f6ae
zb4013f38f5d61791bddcb6339cd04d96ea272c351a2176fc018b173829cdf2995e8817b09c877f
z087ae4fb98754aa0e219d78a5421460b004f12d53f71157d374e619fce8c26abefbfd5a60adec5
z1233c022e16fd774c4ad507bee530078e5d8a0ed6611e4b5babc16c7f248c6a33019e332c5056c
z80c7569152f84a537f24c3e90ac6c8f7112fed644d06e6bf60f54bef54203549643c73698451a0
zb749f2a1b982a65741a2da1dbc3607d9bae32bbef2150202029d6ccfc27c9453a88c8aaa2dac17
z837e8c6b8f736065b9e1e5c0c10e993318b7ddb360578f3ffbf905b39872227bece49de9df13c0
z9e6e41f7e968047253f42ae8d3f34b0fcd36a6f6e6b7c94aff1dc6ee9e9f3b1ccda761413d9b5f
z16f57d7dce09b5e8e46d67149a38030cb1ce6108d59330d7b5139e13e395803a1a77d809a85296
z06108d792174716ab7a36e6cf50d5681ba8196b3f621ccbf7a581691a09579662113ab4a296e7b
za57d2ade52e7f520b7b54e917b63f23231d941caee731281e7215858b6e3971d35a73f8c2e09b5
z7d82e345a963d3bdc08d506da5ce30e275759e957d532d40d838a74c0abcba7a7f0254a900d6c0
zcf4afbaa0f1d2a4f27e0c0cf7661023ce82545a8cf5ff86106e056ffcdd1ccf54683f81a3aca03
zd936f574d37f556fb0c64479dccf837444074996170036ea2278a0322e97737988ff416faf16a7
z61b55715562053b87d45e45d38db9eee829f7f63cf629a63e4107f150f25d3107b8706829ae5f8
zfbf8b6124ceedebe91da02079e2575ed915ea865878b54495bccd8f907f0f989d1de1229fc32b0
z8e8bec3f717bdd5d69e98095d72301ae9c93738175627742cdf916c909c3319d0ef58f14cfb852
z98d88ba304a7bac91de574966abd1ad80fb41e47754986fe4bfe64002e3b0614b967b2bad3b8f7
zff0533298afd751a6ec28f74f02542105ab8af0ebbab04664ac4022c5e9f33590aea05c4d34054
z1c6550b27c036732564601f9cee6171340c073f910ec58b4c5416d5100051f5604bdb6ebf4458c
zcb53b2c1c3cf26565493697579aaf1db581a76d248d5c82f33e350ee2c1b86b2c06916e9a6a435
z23b3b4c9d108322d7db0786df20a0099f4c40bfafdabd2746ea826e3a8dab5274f43aeae738cf9
z8c4349d59bb87323e5f36dbd4820575126c56297e4b6b9a91523a8101f2c2ab59a4d2db21bbdd7
z877471f842228b255fd49856408f873459ec4a772874c3083cbf1ee1b22e1cb384cd8d8e42ed6f
z3fe607e94aff9cd75407c5d41d8746e1271e1162c2768d42e4a4187efc6a861e7b1e0bc927c33a
zf5764f3e6e6e744d07bc90a0416e615101f280317c9357456b51da56f2b6d9c39b19626f2487b2
zd2bc98dd9c53521d42119567b82e2f4b153d35274a6fe6f2dcd9dcae73a18f22ee54b5f5651b78
z6daf3cf033190a38f3f6da2fddc5e03ca53e735fe94909b502f0d35939562d945cf2065eedbd3e
zf4baedea44e041d6622a08d60abac2dee690c502b372c498879271c8a53b4e0376b4515a185ee6
zcad036411d94fceebb42cd51a7a6bfe3bb3f243dcea3032e0df11061115682bc4c8737822ba2c6
zc9e9ef5f4e932dd1b8cca289d8ecc0e2eb43afa28d3487a9c7ac5a4bdbaddc4414eff965c21874
z35c5614451491483292da0214a6f030ddd644a6c94606ec3c586e2fb3decdf31edc8121e3ef5c4
zc2ea0af6f695a92076f5f03ff14e5e4cfbd96b9ffe83b2af17634835642ce183819a23f41f52d9
zc8eb71e3947ff68557edc63bb045c7dac680f028830c6dc2b0f5893956d9d69bbda787755bb698
z2b0ec5b619bfa479ff7818b06be6ba3f81c834db111858a73503f9e39a320fa38e9c0f0a45cc2b
ze90cdd8da19fe341bfeeef38768b2b09c075e16bdf78ddc63cd3256cff3985d2b0b0ae0a25aecf
zfc7ff6a60dcb1d3d17b73ad0690c523ffb661b29dc2387e36533c0ee94eea4912eb716b0ffa0e0
z2daed7a6132ad1560c33385766a6065cb35bec1094112697ae8ac93f19bfd911787f0274338f10
z0c10489324ca4e3c695eb5f7d82931a638f7e041ecc19d6d67268753cf3bd8e0603ddeb6f63b18
z7fe8e89429072ca29effd7b86588f49668cf11d6bcc91da6c42929eaa61d8c762c34789d390cb5
z2cbc25c7650bc17e6fb67aace60fc1bdfb2948f4f703836c75a60074fe91fa1d5d0bdd5c0717c3
z5ed09ab27e37ed5b0069febee9ad6c867096871780cbd225248c4f5aa5fb1826435931e5f912e1
z85739b1ba28a311c6faddd781e49db3cfbf330fcae605b525fca1ec1875bc5a0866e2047d0058b
z8ce5d98b450a585609ea474f790d4dfddda9b1bf5efdd86a3a359406df5bd5f833ef7a4740bed3
ze5014abe7b8190ace455d3921a8d225f9454719870c966b2626babf895638a193e07a00031daa4
zc510ebb1f5e6024d1bf7262c067b493805b45be999010839109f01a1636bcc2c586621b2354cb9
zda38925de7e66861ea0052864f087c649502edcefdd1f04948a1f2f2816b2cf5f0cff004c64eb0
z55f5d49f44379a458ea83fc920645980a5644d8ed68e4af79b4589682cb68e9f21c77114b0ac11
z3f55ec3eb24b2a7563254b94b2f535c213a7c4514f9aed8bfd8c142a75010f00f62195865b39a3
z65ec560b52e6d0fc0095c2f4892f347b5279b00ddddde1f84c3a84167d3e5ce318315f3cd890f8
z070919c7d8d2bb057ca07c3cfc992fcb2131edcbab9212fee608df6360543b38fe1abe74ec39f1
zbb1b707af745fc02ac4f774b5b4845af9af2dde3858f9a3fbed4a1bd11fb29a691e44a8f25be9c
zb23186e1bfc7a40fbadfc6546200eaa2b91cd14fd2de6e64dee106296542c151c0746f5f10c548
z75df9fd212372d68d7338f93877a1711e0b85031c064ad788eaaf4463e8109375437e5cf7ef036
zb05e3921f4926d3d5c2a9ae887b97c91af613b6136f838c774cd6872b511ac0e456f133143c70a
z01dc3bf022a4e0eb6b09132b360943f23804eef774992ff6f49152b252f14d6ff1c21d92a89afc
zffd75531a58d1f86cc1564c4c9a75a751d5f43adf1900785abcef5c7be9a1c4d3cad38d8c76052
z9def9ec502068ee6f45dbdc078763677e1db21cc74e07c1b77adce91c889ac885eb923b4d6a93a
z07e09259e0fbb557d2d933440940aedbc9f2c7d99313f5106e9c96577b4f63caf7e71abfb40f35
z803681c3ca7a59b6fb1e4dc5c55d5500c4ac26258de6485842e8e2dd4d9e32983c47b3427b1ba4
zef1d206866179afaebfcffc871e660a4d92174f224bc7ee0f9221b9f8c5249152db00adbaa5653
zb8dc1387eb88219999d27fed3990ad0d9863ac8463d2323fec8e372b77e64886920a7aa63b354b
z7bc0b6cca091edb342c4a121ee21abd849ade4643d406970aa60f13a364ca1601753685f34c6df
zbd35395c7919af08cd26424ca59150f321244baeefb2c85abcedeaef05131a2e0131f35ad96b16
z1daab51f7da60e5ff1e5a39ad4cab1d4a0a73de742fd1715a753aeff872488fc8844ca60b3ec7e
z64f825851f1fde8e801772d9b3af30297f4616c6f342f2e2f613cb1264288cb63205a87c55dd8d
z9cbea69147554c984e23cc6c15112f312effe01ad0eaf8cc8924460e75a3d3850095714a3f938e
zb00b36e79cf8410cc451d759df1ce4070b14b722e6ab3871401ce5ec30170aed4a48fde62d368f
z050726cdd2e20a9242c1922f18d1c9ea316094fa98bb98251cf6423547863cffb0844d691a8bb2
ze8149b3ab57a66122aa2813d73fa1e74d8525269d246b0c00559359851f6e6799af03d2bce5a1d
zfeeb493202d78955e19b0ef2b61fcedf0afc7439f966ba2b6c09b13b7e1c8cbc90171e7aed20c0
z4210a53fc594392d878e5c9ba5a3225db00e780a726ae6b4d27c0663a122f3459a586d560c8bbe
z8e10b8135542a82fdd336688fa7b03fcaf6c40c414ffa7a22dc4b9dffe8fc69cde69b71afdbe85
ze2670bd8fa24e5a9159ea4d059f4d32d599e4b68a864010ca8b94acd589fcf093f4812f2058cd1
z7619e81893fb4f7e4f3a930c58061a66296e10217dc207457ce21e61d5ae825a0b60f446880775
z4f84edeb95759bb761fbb5345b62a5f0329cd5e1a44ca2c22c0466356b3aea2fc43f8555224bd2
zad850b30d38afdd1a11979f105436e4d4d0aba3aead2b6b5d40d0e7e7f6d8ad6702ba782ce790c
z1a606232ddba36b28c674dc50844ac760d61c3ca53de50e35fc5918f36cc07b089d8274f103194
ze7f89ef57c6282d3b49668fd763c4448c8136293465916eba057f1e7051b099a0a0e80a31ce3aa
z65d554b99fc3de54fb407c06a5157762998876d1115ca2a39ee76e3faefd2595c6fa6c0b9bbd1b
z9fef22a3fa9056cd9790e80ff0d3f5c447dc3fc52ba94f2084b0146175e5eb74efd113cb789fba
z3c83bb7ff1efd0e045dbf80c8a14523c5066ef0df907eba9417c54b67abe0627c30d8ec6629a62
z46bc0d1190aa964694f1b8f286a906b4210178770a0729254b72bce18ed57127b88c6e2f2e0ae5
za669944d940c34cfb78c860d1566b7a28b3638f2db6ba205e8c07cf479e81e849caf92a08b6c50
za924cc0338a305638fb58a5dd3747c8e2e308e103895b2e9c4ffbac0a3952576e3699c34cbf534
z508dd7768c58e261d70f3b9e4d75691546301becc370398355829b92a9f2114b396e70d2a018b7
zc6ca01bce3d5bd30ca406ebfe69b2c0ae0b8a4c4697e81cc2c7f878b7fbcd14f2aad32328e372f
z89186a0bf1ad40af3618184b2b41d3eae0394dd78161c3d6b5265946981b28504dead8338e41e0
z253adbd58808ae0d59200dbd0ad0aba28611e798742e9b383c6b93301a7813ffeab0e5a699760f
z576e0c2bdb7281059da5650361c7e051da8180209492b77d44752bb8dcfc7f0d399daa96ca8a3a
z6f7fa846bfe8caecb0f1bcf444d23b9fdea4a7d827b87c1983ba755a2d830016b86f896e7aef16
z46248317e74dc43223facaf1425696a9af7c620ca40839c84e013a106bdda9900388886005d905
ze645a22b6e2e0edbce2879bacda3418a82e5a68359d58d9c67270560695b0f2619549af50b0f48
z6630bff5715765707f0a7cce84bddcd7096add80576ea1f47022e8a8b88ddc762b765a3bb24117
zb057634088d602431f64fa87a64d63e73fac33b123f31f911f3689ce3bf96dadc80849087ac397
z18eec4cf786a55c04937dccaa58abe70ecc3a6a754cf6b5f78732283161001b92642aa33af8d9f
z4d5b8927a9e5f2cff94171734d76f05dbcd22d0f75e3d21374fada359dc70861d5783766ccd8f1
zf806fdf520e9a5e91642b3386a9ca3e9fe05ae541ef0775b04a18ba63bb7ec7d9b0451cd25a18b
zb0190df73a58694f17937316ed7ad8ab56958710321e7445718e8d1e40da78d4cab2cae50f7732
z1c89e1fc1ceaf1b3c54d943e23360a2c914337a548fa3dc4194559c4bdbf7b48461fcb1cf796e1
zfdb326692af30c031cb03c4d97dcaa47af61c175437e6678c13dcabf0d46488c3a831e4d6e681d
ze895b57567e107bec44cb66d6649058ed788759252041f45b24d489052c46909355e29c1eed17a
ze149f4cd923dcbab54da3c7c6a0e1ba029e259c1a33354dfeb54eb408a1b07791e936f30544315
zb03a267dd0d7caf2109e12e057422dcea5e1e74004493f5e2904b272f6753cfb93d7bfa7ef8982
z68399a2c3fdef290554fd507d3c1fa4dd38fe8a0518df714b6db540f9033b02806d92a7e9166d4
z677867d578ad87da15eacf315ab5fbdebdd1bf0e5f7e7ce24cd7c4c2379a6c1b314e78cc334e25
z69abf3107b5eead0ff8302cc0f9339d3ec4157af6fd62a91a87997ee0431277d9cf877d50d84e4
z8457054ffa9f3cf289295e356262fa86c445511909bf272399af3764adcaf3f89c0d9e279cef30
z902dfca6bc316d95db578c1ef846339efd98e4bfc864fe3c89ea1df19ffd6b54517362ba134106
z327ba3ccecbb2a922b6802bfa9289f0842dad80f33d7781a4a21555ac2ce302ff6cb06028e6e30
zbda9faaef3d887ca48cf3d8b02bce1e537fb48b13702387cc76fc6dc2e5602a690d59632af186a
zcac3fb08870c23ccf9f008f4d71775289908f31e945bf3706f2a46e20376bf922f0848890224cc
z01dee81de86b696e493eff43b49e543c9e03db35101d77f9edfb19675576493f94f477ece384c4
zcd57d2e2e58737fbe6d6d12a6db96d002e2e58869e6fb8cdc45fdf5e48f99bc2936e4cd1006362
z66b4e8b29396c9c193ad9b99b83ea32690a09bef7f8f162555b1b504e96662c961e6a8d42642a7
zc665d7d0f185e63807df0585a083145bbd84a2430b8d8023bcf85837f4da2e3a69957a7ee3ed21
z934d499f2a6ae96bf0a1d56dee616be7e9e3518c1f8b4f911dc330d3bd2414fb21aacbbbcc6878
zaca7bef62ce4115a895853ab4fe91b32afb00a060c89832221b2e772d75a30497d62ba07bc851a
z8de962f1bfdc38aefec77862ab7f56145793ed5fcd13b6dda0a36b7bc9fb6f9e478ddf594bafaa
za33a660aaa65f32a62482e42350a2fd2a6232a714ca6ab61ef6ee529850b1280260168856935e1
zdba03452dfe4597eca9636216549d77cbb8ab48372e8d5362b95e3503b3447e302c4bcaeedb61a
z7c3aba2ad0c4b35f02210aedce0528a38fc6bd7bee779c3c557fcc772cddbc9419c497c6677077
z2e86c13a2a6d0ce0c46a81dd208b21f37fc50202efb0336026b60b108d5b50821ab77b025a3dd8
zc13e5ef4eaafc0423ab9afe760ad20e360a726dbdac9a77fdaeb1bdc74d3b289dfe494e903d3c9
z34d869f820f2c08c1440ede280f1bce71e0d8ec879e19dee20381a03cc094094e64a49b748a85e
zf5394e5f55eeac16725b254f4d5e9f550d29b8092000309438cc68946db50626ef3b087380b432
z3d5ceef2de89e428fd071434a95c386a3cd115582a091df4da9832ed8543bb1a9927045412a8a5
z4a210e244523979e37583a1d9a5ab1f117279f092a489b536f2e6d82cf4946de093b1831db85f8
z8d3585142ed7ade64d9930197cc0dc210bb4a4765bf8401d9b68e38aae2493acd6e6b0845ca9b1
z3423a8b32e4a94c0b6f960e13d8fdfe1c73a2fe2f94f0e39df7acf86cf2a53adb18fa82216e44a
ze6573e33adb5abe0fb2a4bd105abcc9712ee9b34e523d198bf7fd7f27efab1967d61a192cc3a2d
zc313f6e995da2bebcecd16852316e60b63d70703378a12b4edc832ba2a4c893be298c40ddfe5a3
z18750b8fec9e4b05e00869ea6b3510d8151f7b31088a7ad0ae26d50a31a2abc2d5a3ae235b1807
z540272e662ff13eddefaf3b5412a557cb9d26a687b9a852ea4cdb5681d38a5ca800df9f25f3f82
z1053a68130eb17cb29f54e3ea98a6c9bec77367bd529468301a89e0862bb59b2cc8c0334741e35
z519345b8f278a359d8ddff6ae6dee9fb334368729ab525f83995d909d63a013c7a28a076c803dc
ze0ea4f15763edaba4868b4c06b4f6247e52d47e87bcd4c880fc3ac5e200765c5d289bf8d612e48
z74479c9d5a9ede40e4879df1ecb6686e55810a9d76c1e27184a3efa27eea50ac39c6abe40d8eef
zbd57769acfc15a4e9b4a69b8ba0ff36e7dd73822f64bf343f80e9d847396cc2d45b4821f1ea28f
z203cb2672753a1632ad26a6aadca7fc7acdac69377ce3b42b1f5b02c5239f693ae17d478e1dab1
z0fd5655c2a92ba34bf0b583515657041c899b34d638c73ce7e2ab4558a6c7e0b76c3e7bcacde82
z287b45f32883edd32fdd46a7b10242cc831257183a5b75fb32bc3873304b5745a17da942c0be7c
z577eca49975219323280368b443d67b16408bd0cbb493df36a67e292edbeba2cfa0f764e4396d1
z0120cbc7a381cd810e0f61820601c38ce6445a4c4094a5d8f8eba735f9281fba63fa85548fc251
z3dbd9fafc47d211e19717002940c055d922f760f1a396e04d23a7f0b7970df1d1514bf6e00e7f1
zaf166022829d3f26ac614a8093757ff74c2eda41435f19b109edc854e30cae65a2929c2084eb22
z7697054a8d8b287e2a215edc713541e5b4d910bb54235f4ef706b70a32b82f66750ac0d9802950
zda38d5bc24be87cfd2b0ef2dda73d51e9603e987f20104d48aec18e4afa74ffed50f2fa709042e
z6b4be38fbb099fbfba8edc767b4fc4747dd5aaf4f7ce88bb1ba5173e6984498fef0aff02465c57
zad36a8869b2c306074432efffd3682735db3a02284d93b0f5637918195c6403038355e209a74e7
z5b00139f19acd63ee77ae3fc3db36d02f85a48b7e46a3b31f7be45268021591ca63282f60f50f8
zfa0872b5189d551baced38a77e0b69c9a4851f6c3a7240c461db038e2c36a948aa6887150d5a39
z2247ecf2ff6d0812fb73ab920afad46c44592296f5652c3f01117c2f9ab9a88948f193c08eaa7c
z95d44189b854e7c705474cf90504045803de30994d966fad5061980a47d95a8126712c6f98f507
z7b6030f5be82bdfb5b6273ec5888bd64c5c0836b7d760a58fcc90b8e951b252ab1b1e74186bda6
z27a4e1116c48e727f7c156cf577f3d420db834a2457263789b06bb10fbefbb731dcfb0810208f5
z0745d439deb7ab3af86eff622da28449435be4d43a00377883ac58e560d66e1523c8768c961bf5
z87598d715c79457167c2e8e0e1416bfcb27830c8d63f834df4bbc30b93d6f4034f578e86daf00b
zd7a2ebc85783c43a609c5b4a9a349cca325a954f25040b552cc421c0e093b70ec16b7efd4d5a20
z84e9c603f29ffccbe7aa79051c33da2ed1b18fa3408f22c1bd0450b381e388dbffaef4b6e90c1f
z686dc80bbc711a8572336af497d49e5a2c9b3575ae77bd7871c1cb43d79bf649979d9478cc64b1
z3c700a3c02cb09985c366e3006797d012fc1776d479c33477cc937f96789b8c1885e10aa09e632
zef908e0692512d3b9743cbe478913e732b8ce69035771b723db902e7b2d18c3d656009f5611786
zcf14c1b23acdbf763ea70f79acd3c25d9be4ed90925b7c95cf8d7a8fdcb3ea9bd11a3ecb8ddf99
z92a1a57a22c7f77114dc8b5f65aebb868de9c48ee276d378fcd5733ae724bfc5f74023c4f4e7d5
zd4b607f861c36a9e40d6ba5a2ac2fce176beb402a23462c34d845b608f7838db487f59c9ac3f2c
za83527acb4e285865e1bcd0f2991c4c008a5b914c6640c260678597f568020198beaf54a5dbd04
zd253295b35dd86663a58fa4a75f014da8c703cf18bcadd54c1c1a1748171f99ab3bef05e9e81b5
zf3425cec2c1890be4eeebcca3856b9c3083fc99ff520a57820b9c5a60754e0af0660bdd6b2a58f
z5e75e1a9b0b39c03ba5338379696dbb92254567c7803d3ffa502d855211ba6da4865875ec1d3fd
z43cfa89d9fbf9dd00f3854441aca0162d796068e0371d34a9e88f0b25131db622ec69e382b2731
z4f1555d854cfccfee0a38000a9100824277f4d0be437a0096e09a466c240866b86491524d4ba0b
z2ecfe2aa889deef9213e2bd99a2d9e54f50fb9a0d338a89d844de48c820af74a33ea624ffb0686
z1f2ee278b2187c8cdb2441e8bc85ca2cd4e63647f7b3f5190468cf6673f094422b321a367fb16a
ze04ad5ea408bbb4dc0e2608252dc077c603238c44c50b5a9d6e98716d630834891436abf2c48e0
z23700c13c08882120c8f1018022bf19451f10430d2edce3aa3d4b9c2390598981ecf88398a3834
zfe294c914977581b07e20a09c47f1169230dba40f1ef723930d3b80c223d5cc79b2a8cce62c6a3
z406c01d2fcf79c711df9c489c950b4e73f8f89ceca9228c3b67f3f7754de3ce8e54d71bd25e46a
z4eac583e80d8045594b3d6709100819cf28792bd33e7bd8606b4807aab371c0928bc1effab3f81
z5af8b87329bfd0d52e91d94c52878fed1424735b273d75cb698a299da6510fed8c32ebce7e64cc
z958452589d0a5d7dd5a73d3382d1e9355b63a58542aa17de9cfcba72055305c0aa7fe10271ca4f
ze7afcdd5f65e494cee395b3e9119db5e9292f86bf59340f2b0747d6438120d9acd5f8453cf2db4
zaeabfb19ddf38ec20cca1ad4e8be4ce5e16179d8b737ba7b78cdc95a1aaaeca381a16fad646f06
z622cfbbbbbeae32985db93750314bfaaa1b89fe4bb74205b18042e8ebb934ca6d4dc63a5fa2c15
z09caaf0c7de198904da396f17c56857e7b83636df9c601c0523eb4387a6669acccaa668552b107
z86ebcaac0b02e9586d636af802352cdc908a85e93c3bc6141919dc281946e4eea27ad7c405fc5f
z3e83e24d402491e7be3acd3b7f68ffba070dfcdab00a6ab1d19b767d0b801b88790dbc82cac24d
z37ea2d59d37f1766bb53747a7801610dcdb9497c98a2f17298936b5566ba8001277ce8bebfccbb
z4c87faab2b23c6552705dffbb89d99b0cca67cad1855dd44cc68738d1fa2b74d0929c599d3599f
z127ec61d831252ffe1efc2f6aca3a75510d83a16d5f0ea40a5d3e6bd52313b3aed87b712bd2a17
z99305bd866d4848c64969f66b3a875bbcc2e4ebf89a2738a47626a351f6afee3307f47515702c2
z12750cb4e9538977447ddbcef997bdb6d46d50afcbee017ca434a55f1e558cdbe1dfa14cced583
zee49e9ff1c759173239e5a57d8b1ab956109e1f9c5e36ea9730f642d3c8f4f3abca7bbbacec9e4
z3379e74bd46704510c132ba730715e3ac46e2464858512c2a627dce00f1ab2616f62a3b7beb81d
z6c327f7055c8fd7aac91f46571202e0f765a950641fa9c1023d5197167476380b0da5770e2de0c
z1ce49d1c13245613961959dcf7c0303a84c33fe7eed4e77df81c5c11ad3d532f9a714f933cd417
zfc4fc36016aee4ed5a6fa491b13ff6bb5e3db7a4e446d33a5c0cb81b53affc3abaaa7884e0f04f
z39e76873f011dc755ef332e5d4166619f141a6fee3913eecba8c01bbe6830eb487042139ff56d2
z9839142a67fd138edfa32e685cc0859cd752f1e5b91048efd2c28ebe906649e8b906d95521871e
z9d906ec012f99e01307fc72785b6c9b61944f52eb25b6b93eb6d38ae1b043516e721952621a723
zb54df7a30789f12a5076bb964ac5a44f3d891be6150621cf0268c588b1818c68e9742f0f53083f
zb334f72105d42e8da8935897f0c5e94ec559353baa9d7776971aaa304e7f1c9647920c6231fe59
z5807cd2153cf8b2cad11af1bcc42ab162b6a52dcbf673c31b8918da9078c790600daa9e5a68f72
zb02537d9b3bbdac7566f1ea08dee18e5f9f241f286e967666e6ca85b40b253ad6b0f8b604cfbee
z9b1ee00c9d6a5e9210e86f11ea7e66e368d785ab7e90220d0493cd9deeffd9151aa7bc2e60e1d7
z44854726a9352dd175c65f6b3c60769d0da9cb867e26435d1e8afc702d8c919cce58b57ac6a5d4
zc84e8aaef124c1e6ed21e54491e9c122c35fd7829abb38e93428e05eea5a1caa20f1a8a556c4da
z3640c96281915c0359b72add6c501ead348de48276e8aad02023e9b011a7516d447620c50dac20
zb81ed8ebf20a7f2ac83f12fd5b4a3f2247819a0960d04ab48eefebf4654459109e5d563e4cb1c3
z22bfe70cc82df859db2c1a20efdca305a0b04b88a6ce2cd6ef0809ac354be7019c83e685b2b206
zc32c0db250bd6d2f136df60681160f44ee5fe614f18bc1f1fc15ae23022fbcda4bc539b5cdfc74
z39269fa23a71f32557adda45304ef2c7f7deff5a238c5db6ea6a4c39385e6381281c265a6f04da
z97051408aeaed9d62b4e86595583263f1af2fba6469c7968609abdf7a4c67511fa7f5babf7aa6d
zbfd885629025fbf03a2cf0fc1f83d64bcc9c6f3a501a953f7fcfd287a77917ad8b3e5b6c5a227c
z29685e90642fe7f763cec43ace4ccda3269b0a654cfc1ecadfe33b5dad544051597921a4e54b42
z97a6d0701e298175defc13771b514179ae87b31abbb22ca7437709231a38eb2498b5e0c64f0dff
z7c470ec4c314476932470f61e5a85b4290f4a8341d380cdceedcd2a1a1958c07719bdca3030517
z1d1fbaa74fc4bbd9979ddfbd5a405f93780b90b5cd75b2236c90e1d09953dce75903e977191e93
zd05ee0582639e3fb7509978535b5944307414a0f5069d761e41722408b39d25779d0e89e860e84
z3d29813af0204b8779a49604676a831305c1cbf0fadf8f2079b47e49a496bdd524f8245f4c89df
z419cc6ca281b3b41a2b401e1edccaf3fc6e6f281afe299cba0c5ed88b534321082744b5a0d71a7
zf4f5f115e7b1a63eb5a996be195d83868e1541424875f8e83b49a1a6eb284dd6f5ee4b971fbb5e
zfa6612b241bc65875a6d60f55128a723d039813378a47f2d0fee7bd9c51339260bb88199d9dbfa
zedb404b94a335d964eb5156fe8c1151daa41a9b9ac90876cd3a98192dcf4d8c0aedb66d2c6f232
z642a63717f88bb643d0fbe74ac3838f405f815b981c503c2bce30ebf57daee6ca6d9c5c213ac83
z60b7c550ec84385e22c7264b49d9ce2508a990ee0a93430e8ca0e790fef184da3db62c4e37d541
zaa42e1dbf150a3f0d19b1fb4d3029aaf658d569976aa7905549b63bb14ae55b97929c604d9c069
z1f482c654b4965498ab03cae1d2c4f7b56f5baee1018082e167576629bc56b7b60164a04e04d0d
ze1dfc0c9ec35ff296f9f7d176e50e5f21e9dd26a091f3838138bfb29388ea7f59d0bd3a293cada
zfb23fa020615b271f39d6719b70411e968abda9f467b4e58622a38ff68b7300addc1ab577b5884
z2f499f0bb0c710b5a4bf8b3a4578bc9dd469d1d588dbfc734a00abf1a042eb70c1c8808d469fda
z7fbcb53e0c063b0c8d3cfd1a8a0f7d84e253d603d7b7e752bacc6328b6c7caa42f123e94cf52e5
zc77714dd6fef617d999d125cab3b4685c800e491e6b0716517dbf6d802cec1a75eec1b0886778f
z97093b18ebd387546d77c3eaa2a1e669cd6bdc70a8de3d3017c4ebe0c92d88d2f1f2382e2f21fd
z61793c2cc112a44fcd06b330557d2b24e4f0ebb544510ad69631cbf69412f3dfd18f7b8c31efd8
zea19b8a0bb6adeb0636d624efdaaeae5a16d5309c7e866ad176459a98500d8c14d00f34b3768c9
z68bc9fa5673ee3cfb830b37b1aa1d75cc32871762da69e4f36173de49620affc6721b7d3da7d8b
z2e40398ec188a4120851585a2b7cc50dd759cfd2b0bd8624d7759e2538a53b26ea5cbe52785a1d
zfa6fa4dcf6df112eaf189f7d2ef5535e4235bae3e8d555bdedacec6e9e868d7f65202daadaded8
zc2a8ce3ca350a3d7127dbe2ecbb073d4a13541adf6c8cf0a9cbe3cfcb4527f44e4fec2bfa27884
zd347b30003096e5f400e8e7f3ebcdca389819d3d702f7668b2dfc5a65cbc31cce5853cad00852c
z8172a0818885a46c54fc9abb38ef2744970beb57480422f155717c5bc0968cd4da663181387d3f
z508fecf54c4860bb4b8a7a9e2dc09bf2d1524fb1246e3069d2ffaddbff42550c537e61025fb656
z14bf68362a784f7c907855ecaa056f5d12d14d3f4c26276a2ab1c4605be18ee52d7f42fc2b1bfe
z25607f73e83bf2a1bf83d925f06745e163263eb8db7b4849b897460510e50da62d0a304dca19d8
z6689bd51c7c16e7929c34a9e525a8993b24dd91150d03a5c9aade9af7808273acb360ce1dc2f48
zec7e370714dd1ce225b8784a14cc3762bdf2a7ad11360571b32a7178314e6322de8a5685f1b3d5
zfa6a8dfcdba4bbb5d17236d20158726083451cdb106413aec3d329e8001def6f92ed8e07d35e03
z59f64a95b58a61c7e3d2ad9626f5b50747ca5be87cf6bf86934d3b87a55373943ca5fe31b8e1dc
zffa36301ae5b619d966aa2b761e5b37a717c0b6be5c3c12b1e5d6861aba2758f476a3dbeb068bc
z919bb5d994f46cce1d82f321aac1ad8bdc9059ef746138c084fa8ed45a72f091f12887e31bcbd9
zc2f7920525e8a4cd74a9b54c7ab1def5a7628d5615d6e1eb99fad4fdf7fc44c344cd0cae43e804
z345f0cece8bcc65b4f89fbc1ffc54b1e88897b555f8dc1467b1dc3ac3758ceb4c874470784fca7
zc0effbf4106434223b35593779bf984abd1dc5cc53818029eb317e72c670df4fd2049165ab5525
z9863a23825eb8fe9f0af5a0f863561cfd9db1e1a8e8e1b10ce435b102146de5bbf72e8e8e3ec26
z1b760cfdf49fcafa597b837e7f7ab283b02bb4ea0e63b53d84a08f3bb52ca6d2a101633f3d5fa9
z33dcb4ed01fc63d6ff658d0706dc05b21fba449744284eeff95c2c36bade721f374986199e9402
z483f43b45ce7a45e1a237418c5b121b6c9576b04534bdc871d1c079cd4e97fd816af2882035532
z2a190c83c830ec6c279570728aca43e65b4f34620d0b0bcaf9c020a9b464dbe5ccf4b3e5414810
z8333b0ab0eba082d222195f88f104062a72f371c4eb13bbd9a5223790f127d10ded5a1cbd24344
zaad896dafec2f444b889d9d10346ea99a61d65020d5ea40cbb7eeb191ed18c5151532203cff77e
zf220757c755b07eba6ecd94e304e62971c13c1101bc6cd458d061ee313b755b58ded4846e70178
z7ed3891293ada0d94e62c9b374f17e7c101aa69c361dcadf31c39ba198305e2c543173f9fe5003
z8dbbf6173f8950c5eeacb276956378390d68b5c66c1cc2f092cb876ca1db5f1d2c2966abfdfa16
z2858d841a2646b2c65c05ef37e2086b15b86761670e02a2d74c047aa5b2f59eca7140be74721ee
zebace2b56f1e7ed0b35bf772faeb145c0d91c15d539c20330a58ec639baa90cb8f15692f2b9455
z3d58e8906c85b58854d3d29bd0480708117c46973fd5e54f4f457c66bdeddc790f754195f799a0
z9047f36e0ff7bd8d97f5dcbb78d3a5cadc0ccd3f7937ebc0210d7a12313e6129a23e0966779da6
zf0f82f77b8543baed7327c9b8ab0114190900f1520923a6635dd8eb07b908ba06c1103afdfaf64
zaad4d0e98e99da3f1c68d3ee492bdd45c85bd989ecb841908db227ce9af847bfc0e9f6372cc027
zae6d6c14fa06ec1a7dcc93cb329f6fd072d62d0dacc141593f3c224e26bcf1a990756f72db468f
z19a858b32b1a021c25cf963ea749f2c4bd97cba4245ddbaccd93bf1244dad39524967e3a3adc12
z581f02e01df40e4a566dcfcd5fa68258996144147026c8bc23c06fbda505e25d706265c18a9b3c
z97b73215606f131a29943bc0ac0db698d07f48c2e663c2cc9a61e9dbcdccf451aeec0e59b380d5
zca3910c75735f6285bc79401c35ed944c24b708253a2e9618b8c777d83b99347123fe6c2bee2a9
z2554bcf564fa39f2f0e899ced769d643ac2bb0880cb319957be1b6882b3a8999576a99f1b671ea
zf26c98c0f79c0c07fa16c10e598d3c6d96a7aab8eb8cafa01d568d7d02bf5c18f428a25932a419
z0b79605facbdc168306dc73ef16264b165eab525d9ee74dc49f658f68cf018c89683dce3bdd53c
zcbb2cd6a55d9a10ce114620e1695b42921d6c7f68429c9a3d43a2832e650b17135ed62a9d405b3
z3b72f5d7bfcd97a5993695a6e9d25ae3b0f0a5b8ddb53a03817727eb9b898840ed4e47f94f2f48
z8aecdf7498cef8cf34305e9e65ba19d744ccfcfa09b3193c268fbcb82995e8486d4a8d0911199d
ze446f84d325640a4b4ecc913a979eb69c94760fb016b5989a5a1c2758baa7fea377cd8f9bc989a
ze1ee498f96799c95119d4c0ab0c056dad2e3b1180c94606ed3465a86dff36d0a3108999f5eccb0
zed9413406d76607f624e5dcfe8c513164609bf16f552e8b091448047f753080a304dcf37bbef44
z9cf1017c4efab3ec708db8f14fea1366d02fbba1053ae7ac6faeb5f0d9b7f79b0d8edf20be3523
z2356f549bea1238cfad4719020c1bceef08e2597f348242b23be265d88d5ad440f69eaad124a1e
z4fb3d54a714fa2278189d032c1b702ce880af46acdba9294862abb0319b0bf5d0b5a528ee6bdf3
z9bc02987366b5d18f0cf2daba1a51185c96b2a511e1a797e8f52257e0a1bdffc38d69907a70ef7
zf92b3a40e1ddab7f2b3c89dbf44755140530bc126a9e945c100fe33f28e87b631d5e44276ade3e
zd8aa03567c55109d18c6e1e0ea055de9fc6aa7a7d31cc152ad03628fa495b600899c46c68d13c8
zd71598e5b980ad1c45af6ba8c4bbff3d7e0e23252512764688fe254afeb0de8f247d9760fce397
zdacd6c337c3a313ce593b603bbb012fd93a3222b547276e6e4987c45617b12f32d7a9b2ebf5bc3
zfc6ad8d35816fc7b1f6d8eb1765fbe9ff96ca7497e6cc8d30e0549be1f189831faa4bd3cb8dd65
ze7e4e1e003ad97f69955a16f2090e6987027dbee76b5d3ada0c2038a43ad0b911ffddae8e5e798
z44b02ea4d8616f41fded340f9765ba6a5a347defe90c70bdc807062509eea736b68edc590f78d2
z5b30f00d659a5bb684785ef0fc9d1bcef9454a2b0d82d43dece34153d410aa8bd242d8b602c71c
zcaa2353dcccee04a9a9dfd7f4f02a1ed137925d12ce40219cc85083354d09c835811d4b9e9dfa4
z4e128f2f41a1320f08f01b3bd011bb9008858fece656599e70248c040294c7bd5ab7313d9c46fb
z0deb22f8ee578b342ad42f6278e5dd5ec5c74b49557cde39f2f31f2fd234f154ceb1e2bc4eee8c
za766cb3cde6a4cae6e761b5b9308315b54ba34767838a9a8843b197085e25b7f38f031a5fbf950
zf9c95a1c481c6da4b0a728d793549afc65b37ba7584680c89703065280cc3737fad339f1ae48cb
z0efc056bcf894f593d229b32d225ee711de949e4dba524f216721f3bf90bb761c4e11ea37548f5
zb374b87b0e68b0813a003a7434ef0f89806f531e6e8d6a29215345776b7b38897c80274865b4e1
z3b39aa5a1c51e29762d70a44d1c834c60905a88b8cb8b8bc1bf13d50d252e070296d9ec55a6f4d
z2313d47c36a6c640285e9c97aacd40262511905b2bac473d0211d01644b3694ca6675d6cc8ac84
zeccbc14609e3141205f7a6366202afeff8ac093c50c47769cbc57b2d1db3bb14ed1f279a7727c2
zf7433cb111d380947144eb8c7ba58b896cbecb74d7f217ccf1a48f536dcb5088485cc19ec5f863
z7e6b7c569b61a032072ac0c82fa73446b83d10f66588488507b0dabcca621b4265b1d515feaf51
z276b7091fcf00d9dce045adb20017d850f6e21ab40131bc31e7e56d2bde632f215bfd795719965
z1bf565a708f24b15a3bd6b10337c5f12d32efb7e52d0a9752135f58f5aca81c38d030f52439b71
z125c6eafb2653c0ab1b2153fbfcf902065e52faefd7e9f03497090f107c61d29b20f1dd2087abe
z60264751fddc32140a9391d30ca5ce8ca96a3e039e25dfacdbbf79c260667f5d364bc0a87d844d
zb37afdcc64de75b442ef93d71152f48e81a1ac11dad291c7f73e88219bd55a34f036531ae97009
z2856a800676e3e0e2fb44358c8ed5ca5bbfa1b5111d6b6d64a1cc01b3fbefe6c5209fbb9de93fe
ze991554f21efa982399a0c16a851ddf554f6ae57b320b067ddf7807123b9ac0441bab297a9fd2c
z38c00c2f0f79eae15163f3252893ebc44a5748986188ce6b5e6924259f28801f2007b7c24f49cc
za946f5be9ad7349e76ff187507e9ee92e6c5783a7fe654f2972d50fdab4701dee85b264e97c25e
z1d4270bd53fc5a1693721069f83a29e0f9b6ebf5a41cc1823c76768a8d6e6a002d9f1cc25e6610
z073bb24cc65ef04fff720ecb2b07c25a0a6073f25069a678408d9461f5a168e7cde1819f10c5c0
zcad32d903c77dcc42c569543ca5cf1cf98346bb3c048dced67816f25972daf653e9bc68d32c8bd
z59c6ff5b1fbaa80996437294783a85fd1c40095da48f74d4e1942619afbce07511f82563481557
z0a946296d642f940473b9b648ebf21db020833cf7d72fbce34e4f0b97dccefad8fb99400d11f94
zfbe4d0728914484b05873fe87bad6ab7c0476f49e019c3ada03a069c64570545abc811a279460c
zbb8487a1dcbe32b40fae6f7f3baa752be95a3b52d516d3902a0827b22f2d221cdffa805adcf737
z9215aa3925978f39333b19162304cbfb7a0f47af7e3e7865910e1a7514cf0998ef1b124ac4b16b
z8d3a8ffe385e72b6164a11b93138e2ccd463798085b79aaec66586c8fffe57ebf3f01ee4ffbdad
zae0903f0b0fa9d6b64c58a296863f40fbb627091209ccc6723875c03fc28fea4486d122533f841
zeb41e7127fbc810758a4ff3813124a334732d25fc93fdea09d8bc67d218c3800589e2be513db72
z877e7b918144bfd8c41257cfe719a5eef4abadcee7492359b5a638e4ea927e151bc6d62abb4fda
zd2d2c138319e37aa23327adf05121c02ff47c47ca57956e90d75457c79cc9eaec1653505408709
z5798299d3839fbf41f5dca1aba7679b92aba3bf4b8c85bb55d335f532e7e5ecfeda77593212595
zb7b1b2162ec9f6206c4cdf34a1d781672c2d306d7d4457ecb73652c9e926acf93f4d750793fcab
zb63de7f1f0bcd05add568ef2c49818a5470ccc51d7e73e8321f3f3c7fd1a432c4ca9b4e8da46bb
z21206c25e11d7d4f5e26908ea77e520244dc94aa75aeed90a89c369976e4da2a97e334d50beda3
z6615a73bc3b72a501dbfcc5690b0daaa105a960a9fde2c204c67fff1fcca9ead4a386f2df50782
zfa63bf9609647bcb7c3f76f0f21cd9a685ac2ea94dc223f7b2303c3b8db88b596b563ff0dc5dd6
zdb348a7296f15d7c8892b99d118d77cc28bc6738d58ead26a7e91e2d84a3641e2700023adcb87c
z60a7a6d0a1beaa5b4f849bd482c0c53dd2c32628512b37f03f745b2157590fa48198bf6996c8f9
z8f8a0367476b3004952ec76032958ecdea8598d9f82488e46d5054f825e09bb940350cf48dfed2
z93ece0e975b26cf97978acfcb4e4e8be3ae63b02c65fc6c6555d7a357f8ab8b3d8855968d2584c
z797c55ecf66a6c30d52bb1ce5469044d215596fca4024cb29f7a5011170d8c94b1c2362c783fc6
z65a2057da813037a83937a014a949db8098901f52ab6ffa3100bdb40c1a1a54d1ce6fdcf09e2d6
z81644fb78a04ec44d4a5d18612829ea339b72b779fd8b9a59592c69e64804ea5708a3806b389cd
z15ace212a7d4d25d1f491a7944ebe75e258064d392d496f40a92f8c35656a88c3b984341c79080
z3eb7521e8fd784750e66621558ebd74f5cfd8ea2857ae3a6a7473d52cd7144502aa53cc937ffe2
z2a3a666a7d1a6c9bb4f83128ea1af6b8fd107dd9b07852e2170f0f28bb970f25d40b44868506b9
zec38d36ce8137d600a67b49c916f0b399167f2ba663c3289587847919081a6ff3224edf48b6ca3
zbbf117751fc81fdb25a0810adcad3550fd7c9ed061257b5d74a81e17b0276e29b51b1b2ab1a8d7
z328f3bc9e00b7ef8957de66572c43fa32fa640ff584b7320ddafb1727233114e8a8cc2166002da
zb2dce5d61547df2ea5e5a2a173f743df93b9bd82bfc18babfc4966f3f676a38e97bd8eb61e5fa1
z8114178c78a968bffae9f6a198f92e3a18d982e951b87861297c3618c60e94413079ff19b61d26
z616437bd0d6c25aac74d807d0d0a2e088535edd356b6bdaa5b806dc536e7b68f61efc3a0b90da3
zdf3c6dedf9fc6690ae660ca613a222731d4973e16472da1ad070e6dc8d8cdf8be365b61d522bc5
z4676e2125ca9995ba43f2579e47cde2e4f958e8d4ba0661c5698d376632e9ff022efddbb87cdd6
z7345a7fb29596a1010b64e8ca9e3770ba58aa4a666e17e6da049de9c6b8c30b000828fdbbb60be
z3bc134a03f2cdd4b7a33422d2b90202f909bc24a0104e60c451c3f9ce44751e88e8a1c80bd93af
zac177e75b25ac0209b7da84ede1bb8795ba6390c933d89a124cc3be50ca02ce6e38143535b5694
zbfe942094bdd4c74d5062541774e3796188d49ba289d2b9cc96f370d65da10cfaf2b2e85ec9530
z6029bad4bcffa0219f6bb5aae9f695bcba3a57ee34ed84995666295ad77049b4336671838c34f8
z8ecef0aef916fa6cc31429303f4813ebb5907fd907b766d61fbd462c2257f6b3410c108dcdaee0
z5f8374c6429a9d664e2ae4c5efe8eabac98c12ee695e10c1474aa8babda69e277dba9ae8322d23
z746f69206c32f30855d67e9db11970f8303deea4a710f15ed462b8d5eb5494e58f559be0b52f25
za87e30fc8f99bac1526fe0020292d9c6180c2694641f71c1793e8a7003cc05990a8173dc5de81f
z697f8f23d4ce213e296f50383d71c7bed9d4bd3b4ac7fd4bdabc8720e1bd9f9f76d2750c826868
z15aa36d43692aea2a105acf41eadb8dc555c220a49b5c6b8428ec83db55bbc8fbd31287dc5d5ba
z3a267e26b9032466250ed6e95b2e06afd41c9438ae008a92ce53239c0878ad29d9f6bba49fd815
z19419e2862da4f291c866db0d7cf3fa0303b09afd469038c7b1b262abce1ccaa36fbf4e36a3149
z1b2b68195708d891ba13c37b4674803f7dccbf0f5427c905e258887fa3278ce2e411a5cb8187bc
zdd0d05fb317664c0205406ad55d065862fb98ee48aedfd7e39a1c5a0fc6752f9a8af60ba9987f0
ze09da2ea067ff6bf676250881a4840ce9bd606d51a3a814ffdb40b6b8bd33f83359fec34e99b73
z63318b073b87f843a6238bdbf7ea0d47fb0d9f5cd22a926b6218c80be89cf90f677f23e6b41e56
z7eddc8ff8494f0e96089a3f5474dcebf29c5bba638b1adc77bac75cd63e805f121090f6ef5fa0f
zad388377c91cd26faf209ed9d8c53f9a5deddcbf21a8c8d00c5d244a99a51f3ca66ce90e0c60b0
z0b34e08bcf116a5e6a31346bef0c73b215d0553bebb547ca1ba3e8654f5d39018acace81ea6ae2
z21a0dda10e3adbc6a6f56f6741eb96c835cfdb33571ec7d2728c4819e34534538c0c33480e6057
z33a9415be592cae7abd4319148c8e3a58780ec68c30b26e8c879c09afb1080736ec5deb6df2be0
z8c57f5ed71c850a5f5615f190800d3cfa8ddf3409150d1d3f10985c9356929a0b6652dc8be1395
z961b1f571ba774c7cdc31929cc28c9750abfd3a408a4374c4ab38c6b35344c99be88d8127f9ee3
z8283fcf531fd27963b2b1a9ba30fe3336382ff7e9b10ec3475abc366e5d433ddcc4614024dfc2f
z6100dc02d77792b4127860033f985c15fcadbc36ef1facb35e71bfc5642b9dd87cb68884655183
zdeddac646a8f3895005d856714202e7b1dda8cd121ddd365f9b95010c87832579f7aa7a46d55e8
ze81b56f2e73441d5d82ee29472e95f58d5cff2832b5b93af3eb215516c63c43aa1c6147f83ae9d
za2a1949049a20039bf4bd65664bbe91ed64906594ee36fc8fd797e396bee112b84ab942de38cb4
zbc1ac456989885a9ae02daf5942b1d9011c69fe2eb9239abbb85826aa5e59979fc406b85171778
z3f6725496fc40b5cbb2069bfa8fab93e7d363a9bd06de6629ad0bce141af6e996c487b716ee258
zdcc5351f7ca9def2c94cc4873c0e6acc1cae7229c55f312e7eb820ca55e9d7ef36c1747472f490
z58e76cfffff9ce1e628527825e5c90000de35f7d602f3c1b097aa0a71a604a2e270babaa78d528
za2acd5eba41b3b3cd1ddc36dbf5e001371e02fa452b8cb097f29d000afb596d5fad61b9a73229e
zad1100bf93d0d0657b4fabaae78fe8b6e5ee7473d69bfe646695a9b2452435a85a9af376197ac2
z8b3df3a2b7fbef7ea7814a117c50d51af6a14f2d2149e3e1fa4f7b7edeaab54e7fe898ca4cb72d
zc290e5c4c4d5928dde3314f46ddb13cbaadaa26beda2b8799128e3497f5fbab42316808e43eb3a
zfc596adfc72a58f746196d2fdcda6057c1e8ef6ecd6b3da090d7ee9fa80de492d2a49ee320e2ed
z6f72e79130d0542a50003386c9c315b65a7a32e0d9dc1e538a0bf7981a2f439a57798cbaa09a5c
zb7e2db0d0dc30e6cc439b895a8547e19e297e56a20e10f480d8ae8bbdb2f9de750cf9fcfdc6c56
zcf20c7ad10977d80df042684f8455e8c8fead698dcd03eb7a2ab29248a6e3d3701b0aa989767da
zf7286afc811623fb89bbda6bb5de07caf7f203974c948721bb221cf91ce104ca164ff585a996f8
z9b6bfbcc423415bc8d9662de7fd626d4271842c60055840c2489b9d1d403c78abdc0ab7f7f3b9d
zaa35ae7a6aab229fb37e30532c84d803657f6b4b5396fc5a6a87cef8749e6f082b4fe59156830c
z88b19087a766d5e57e77a3d4bc52536913134e884fafd51c19a4b894388f96f82c950a1541ae1b
z97bdbcfcc272ec36501b6419c7335561ca337f04c471426e1e226de14353b0094223702884f7f8
zd54ac5c5465f31216d2a671ca877585a01e27167a8d79b34711c92d2dc3135fee5526c292dde82
z0d22b748620683238852593c6c58c609ca14b1b282c6df47f6fbd3482eab2fc799c0111023fff3
zaab556703adc8fb6ce24abeb9eb3291fa97513e6cf4edd056e2700dad3ef7758ddfe641520a2aa
z7bca66728be8480284c38397e7c57aab223c4c136ddabb42aaa4977f09a4912e682bf66b438662
zd58f6c922aa75bd13c3e35b970d5d424b36abfca953b91a7dbc16fad602ee8de9c0ce6bf7f296f
z089028699bdb62faec354a64b45a5cc4742b55cff2183d2e0228ea9018a07ad905d912339b6297
zb74af156afb1d21af778ec69c848a6a541eea2cf0d9de2977c0a3ba2d22ee75be62174e2a2cea7
zede55c082c28f2802960fb9b8f45cb55d1bc673e6e63e8691f8a0908f3005ca38b2c95c32b5b49
zfc6c1720b09da01dfc9663d7efb18b1c3619b3084ad5d1624827201ce91d5421b694ad9580948a
z0c11ab4994887c03c6014533b0b6241ffd32d04cbe8c8b303b4843a0cf80438b3fee7526011882
z9891024c8ba4d86707a507dcfc6811c9b067e09147d455b580ba630a05cff0637101771db4065f
z5ef6726fa7994c23ca7a8cca7efb2d85d0493c9022b224ce5bedf7f9298b6a43ffa29c6ced293c
zf0eaa3321f7c64cd758650bdd5ea99c75dd357e7cee45720db682db31d43d821efbd485b620be9
z8623f73563a72fdca2ce073abde1ea68cb0758e5139e87b307dab50efb93cef25282ec04780876
zda5ac8c99a4f580cb742c917c6981b5990b4236faf9b46e07bcb90f3c586dd1ee97013230d9579
zb667e0c7dcd6926f5fbcfbbbec2fc679ed12fa6796036e5bb32ded5b95150d2c6e2e6e17d504b4
zef42882e44674a2c34af5deeb4354e208f64059a36b9b5d717d8ba4618d8fbd30739010091cd0b
z079dd08ee312e064fca45c449a5cd744b3d6e152264a7a1c32431cf2556948ee04f20fb3e6584c
z6b1b5216b79e9cc0f6f5af2be16b423912ee28cac88b38de242057feba8966ddf0666b05b84cb6
z31a9ee8feb3bef9f477e499c33baf52257e8833e2e1e573ae59e4e2895f87d3c5857a159018bda
z652cbd098e30ed904dd176ca2876f315caae215dfb29cfed387a9f983939ce1e5cb84b915f2492
zd71cbc162996525260310ece4206b95ab63451d7eed29a0eecf68131931ba196070f0ca34f3baa
z77f1decfa2dbf509c4e8318d64edd6ecc3ac01d969c19ff7ade1c400cba4db0cf7e5d16172ea88
zfd0d132d7f735c6cd1189216a5642a7d66d00e7409d755565a20a282ca0fabb3946508294c702f
zafea57af7c65982e7de41d2b0bac8326195900194cce8d28d317051a7b9153c79f64c2a009be85
z9601bda8221a7f4bba9d423e97a5ac51650c7ccea682361df6aa02dad02685dfe9634bad405e4d
zef5faa11d3853ebd6764abb6acb5f7c5f661b9dca478fc0ae4a0efc96409830b30ff051065d6b8
z356dac53e7b23f3c1c85dc9e122077b50ed25024df21fdbc90bbb7718d7a5cbd7c20bac6888127
zb21c891fa59d0fb5ccfac89f58a93db06a447cf3d0285713a7bc2f86cac9bdba1c7f7c88e4ca25
z2a1c621ee972b2a1b12cf31bd50c0b93beca3298efd46e0ba00d7f8407378f200dc681edc181dd
zbf4b1db1b07307f9444af3e7cb48a4d5c2c6f46aa8a8e0135aaa4f3311559101a2343b72a4cf53
z3871c003947d476311e1940040daf003c093c85f025391229e5f806efd0380eaecf94c792a3d19
za7c9e57ad2ec49a611a20e255c9df2c5d291f778ee9543d4d7d03db2655a2924571826ed4d7d19
zcc7a297f9f103a5af860bc9f2ad989b0be8027c090907f1b2039d076d3122d7013aeefc173da5f
z728d23591b6797848eb3964d78c2449b297057d8c7aaa96e98783149cdeb5897cc26cc4b67c8ce
zcaeb0fed6bdcef7647be5815f9ce23c208652742fa0cf2714e6dde3ae3d07918c8fbf658d75661
ze00e793a96eda45be03aea9b2863b4f337924cabc80a4d15bde1a35f03a4a1f4c4145432223487
z95071c7bf39c0fad738c87d7fa13ffaa0c43a3d0ecb8890302766c8fb49245f632b57959173155
z7837fd1028bbb7a60df041c9a67104aefe293a098934e0acc43e4bbe4eefe1a587282069e3c9bc
z0d530ecf26f945f924f352f26190cc75eb30725ec06717f8cd65f6fa68039daaa0b23712c00ca0
z61c915344837227092c4e99572af8ca85c17649cbdbb12dfcbf2a886690e50cd8ed86b8d31b81c
z65c0c8b69631dda6deb48672fba94467f90cda0126480da3f039d92ad78b81221aef291391c19f
z68a10ce0fa3a4e9cb21c1dce56a6b5cf840fc32bea195a28e842d6061c7eea2e8fa01aa60e4a29
zd309490c9bed4a46c0616a0cbd736963f98d4d7b71aaa8992fde32c27e6a48362497f0a8efd2a9
zb42330655cb0302950ba110064b42f27977b10d5c8ea4750ea87c46c0b1a9f0b4c44b9c2ed9f72
z3234327c5ba5d85afe0ae99a5cded398cd24d88279171e9a7d35942f2fc210b4e2b51df3b6f036
z716309584504f60e57f10b9db12413b9fe90f3afc181ae1a8f782dc6457bb49b7ed1deba22f748
z2d820cadf46c0e94f86e4c95ea2084a8c571b4e11e600a9c300cf2e9f7e74bf72e45f79fe9fbeb
zc300800a61ca1e9929afbc96a11734c155707fa380e58efa53e24301b0493060c235ab69e88251
zf9a128d08031a18fa1b2adf04da96521a790571256b6a519b1b106d5440d3aeadfc8d4b2539889
z8837f363c3be379920bc08a53393ee273145b6d7965f4be352a1626ae405c6ad8bda65806d3ef3
z8ab2dcc2a0382cea8f52c30a933b8813751729aac9d2d9d386093556c17ba73de34f51243659a6
zb7b3c2b3c6cdaaa025ccd21f7e189c584d83c01cd4762de2bafc7675b811548f3af0e168ad1b51
zdbc58e2566c6958da6039f68ead1fb341aee027fa65b4ec86bb89b811d05e687d39bc8d452677b
zdfd45034e1967301777b673eaf34e1ab67951c2d867c031d6e91fced6eb46064ea676bbd865237
z2e29be315482fbf958b34ece5355576bd5c8be6ae149808fdd9c4dae7c82bf6e55dfc201251b8c
z9ceb4768fd42185ae4ecc6b140f566ae0be4b70ea30d0409defd40f61a7063c71e879cba3bbcc2
z5d1475b0913d5fe4682afabc2d3cefe53cedb15106a89eee7acbb45fb778c92ac791063440abc6
z945b1b9d190461f05c49a157a74b0490b1984eb9d9e588a1ef856cb2b62cee650ff152ffa6a3fb
z3e98521bd6e799daa25c987655ea56fd6c5d0a8f80076c28d3534df07f7876ee29f53e9873bf11
z03e47a0ee79e77c42ed56f2e47fabc7f37c4ac867fc8387913e2948f9833d1820ae3e2219e9eb2
za82a8c4502ee8a446d83709e72165427191a3ab55166d14b8aa599ff42646d6793af279ee9004a
z4b9151d97f83e718695ee0d46fbac4eea45ae0cbf925e1b965a1f1a38b614f3491b8d4b10c373c
zf1dd27ab75cd3a175f0717782f97a9b9600f6312494980506c0c06a92b6df63e86d0bb5d0553fc
zd67580f02f7a775cba740aadbb3957506518435f52c441e3d5d75ad7674205919eb0b5fc5a77a7
z41cfbb735a097284779ee96f2b539d16467be4c59f659a7c9eea75e5ba6a6fd7910764d88fba81
zd548fd5195cb8980b8a50828c2e91c12c02a1eb7fc716dd6bb99241eda6d333ddcb96945209148
zdde424f03e3402536d0e4eae8f8c9847110e650927a056216f01bb9119cc528c82edf9206199c6
z65c5a4997b04e78d9b9c3eab29bcba62f06f45acd79cbbc9b0f186f04f1fc416420c525e41cffe
zc149e501ce31c699c6f78af7b710695a290eea21f446aaf4d30dedc6bb9d9e26517efc4055306b
z98ea54bb345c96dbac712a54c9e08c97fe1a4bb48495058f119216ab0ad8424e9cd8512dbbe5e0
z8c31f6905be8b11e4351f0b39bff33dbc31013b9797061fde80ed5c1eacbbb6f25fe343333e346
zf4bb3436f16f49352e9a5697e3dbfc2a9c1aabe48317a8852f270f13ba9f85899ea48ba876d1f2
z997969222846033b4a72dd88b3c6b3c5c269c8e8b47baefd5248b9292fac3cc4b022cdfd1dbdae
zca67e056ccb8534120a519ad4039ed66995eb6783543a83f3119dfaae16bbe46f0f468821145f8
z5350e46acf2d7e790d533d09b5de0dc30b3840ea6690b6bfc83087b91b11a1223b511be36f38d0
z9a4fa528cc887e32bb9b14b58ff50e5e691bc16d02fd1ffc6387bb38464c100f3405a761f2b5d7
z0e3dea55e52beceea0f1006be4e64c2305324649228bfe9c16e6bd189a2a96311e183cbc5810c5
zd90e7b79257630d2167089e00efb0bcdc1d0f602f77908b97f42ec9a2c9717d645a75d54e11082
z7160ac6bd5a926964ce977e7c3cc5e3a76faa1de6015590a592e85e58ac50ddb171003c74840b2
zc7ca9d477c849e2b4429b4f4f00f26ba9c39cd90624529d5f780fe75976fb61db85200fc2ed921
zb3a6986a009e95814ad7b229c917476e526392a59a4d56386e9fbc86d79bac798fc7eeb787f632
zf7ecdbacf3b321ed357e83d7574243803e68832f8400705108fbcb0eaa3364fd925c0bedbb9722
z714c169296601d80b540f21c281f522df399d3066b2179d7fab971e8705cbc5b1bd67e3706072e
z5ba6f4dea153cc1ce4fb2d7ae292fe0dcc8859baead28772193039deeb01029539ea13b65fe26a
z3816a6b4c7f594daeb1ae09a066a9e99e79027ab9c8144be197aa3ee03efe38eac7752089ec9ef
z66b565abdc4f62b7565f75190bad0d5361fe3f335f84e9894084fc4f0315e8ca7c079d30a47ee1
z24de017a689180259785e6d98cca548dbf5744645b5bc0dec6003ab975b2bd0aa26e390931c016
zcb7f945b30a2e6ee7643bd0cbdb0dc41d27120aa772551ad633af7d771ba8cfb3bb004ec55afd4
z589624c9810d2e23270bed9fe18e603338321a222e0c02ce8c052338e12de7a09ee2566edf002e
z7e266ce7761d053cd51b5cfa03497de0245e30dbaaca1c696db84cbaa2616c49325d4fcaf266cc
z5c86e065b2aae67bf6863fad29118f86b2d85e69ce3861940fbc350041d9807727e4dbe19c96db
z08614261df8d1222b3bee8f0c30af1cdd118ca3837fbea99200bc0c602b8ab92468c114bab2f75
z9c1cfcac83fc972b84ed370735b1e26faed125036d1412ff6a6f984e0af95f341bac3803cbc4cf
z7bbdf5d9f267413a4948a87a14ddb0f2f84d77412b38e37563134e5946ca68c76ceca5e36ca0ab
z51dc8b8c753c00f0ffde83a6d97663c878476402e17c93c0083056ff5e9e241b6a61d345ea6108
z8491e3674141f496fc3c81c5493525ee783628352e1d1cd09fff921b930c6ebea69f15710337d6
zb633cd451ecbb5c3487196c28229d32abe22c86deca16f80b3479180d1f8d946c892dcf3467dbc
z6d5611660a0466fcaa1e1fcfb31c65fd26af647063d9005a9dfbbf92b9418214e9b0777fe82c62
z5b4f88e1096e0e060ddac2793642964e47f8dca814f002b1e83270783c928b9ead4e04e12fe590
zbf3b902a5df05d5d7bbc5ca0d8978ee41bf3d02bdb9559743a336b3c375f610b6c56308b57081d
z393d39f5ba31c50f1649202b004ca00e395c3b9a5759b7e7ee7d0fca9d2f904cc1f5cf916a945e
z9778b29fdea399291a9ed5dc28caaa992a9451643916284ab0661b88135bcfaff6b915b25b682f
z099df67e0ed69b8b6c6085460788f509fbcddac00200ecba4bdfe64b777b2407de1cd8a24cbb27
z5c292e5e786d3933cecb42df6be85036703dcbb8850f6ccf23f8f8589f14390de5d0130e4314c3
zd7e365d721a13fa9dd318fed9400bdff7fa7847e07a37c30744a1bf7cf8324efe29fd2db2f84d8
z3dfa4bac3f555361d197431ef8882e1f2f3d505ad2588823b5993086a0103b61fb7cc60a059f57
za696f2ff7c73a77ce791e336e2a8657bc409ec6cd1a6016fd4d64a439bbeca4a4f890e38fe6b2f
zcfeb0202b5a6cad34d52b711d215991d534a04405c14575ee719889ac33f8481503b4d72efe1b7
z8083212b60ddce94a20e0a180b19d404ce1f24f732caf450488a6dbf622fab07c0fb22ceca7646
zaf28cc9b79d43f75bc04a9f1bdc8bd4f8a818730abbd04b3b4e16bbc0ccdc2ae55eec7a30fed59
z7617940a303f09d9046fd02e25704b25f45aef1fce2ae056a09b92fe13f74ad01710763230844e
zde42def9aec16c36d09564eb8c78cb3cace5fdab8328273a1ee83d1e3fc91a7d59dd836ec86375
z1fb5c33f12a837517d0e7c6f6f44936965859b27ece8a6dc87d8ffa07699957f2d9da8fd16f58e
z0b6720b5a6ba834310442cbe2b8ea916112dbc5367ef364f62d9cd4dd8a8f4ce33790b2644502b
z6a7529fb8b88c9e8320d6207c2cb5bd6a0244a1f07751df6108d3db147782af4d1d927c41df17e
ze5ceccff1681a2f74f60efb368c66de6b056b01bea3d6a7c93bcff131323d8b635adad663718c7
zb9eaafdcec6289d887180ffe0ce52214761165f811a6d818d1da3180c1ba5c7139f5138985fa5f
z1644a2b531dc4318c03e5db5e7587e244fdf82208462cc8252a3121e8d0680ab454bea3edf9710
z3502014735034f54f47844db1ad190a9ff5c39040d04ce9cf6795dd8d0a12019c707e8d0a9aeb9
zfff68a978c743810b439251c84747d50ce460064ac8f3b26cebef52b2a42bb1b695d188a7d514e
z7fd71897cca08a3606cacac82463c205571bc8c78e667fa1a105382ca204df9f8dcf1cbcba057b
z0a21ff5e7a410908a576096826fdc16d3b935169defa31189cbe73d1cf6649fffe3e2ff9d2befd
z6d746f394a864f3ff5196258f69707591840cf88d3f577e9667c74fde4461d1356c9628704ad6b
z884a9d087be3f3635073df2f2decef2213f02b7e0996b06438818f601b6bc2999f609a2e51e590
z3b4e19f697216b6fcfb0c5b84b1e303e7839de156005741b4cf00a35a700c22c5d133e6a44cc70
z55d6543a8bb39343a53d83fba09d43fb3022b2454fd4a725d18dc3870af22a63b8ad8497321e48
z26a5a5ecc37adc8c387c335e16eb3df1f3ecb6f908776f89e19db226efb42fd17ca3ede0471ecb
zd03303ab9386e5c5cdba70581aa164ebb109193dc3df3581c75068acfc71aa4df88ea2bae415be
z52cc2207cc1a7dc2ad4b10d33202699ba4cadd7410b3be2f70a3213ba0f991b96c493015255ef3
z376f866b0acc0e6b9d2091f75e768c1772be55f660fe3de8df13139efeb7014f5fad004d7f6c4d
ze08b59d7031b8e59e96c6eeb41076fbd22079fd71335ce43253dc46ab47c9f9c99b0d56564477e
zf5bb0b30bab03453c8c8b910943045634cf49624a2d3127fa28985ab1b94cba5548820b099a5df
zb978972a5c0e7772c27abbd2b474a2c39a8d8de173f36a6d5fb4593fea8f7cc9203a06d8f119fa
zc89ab7feb295ed943c5d69a6fa267405a4a0adb906349a97d07b8becad5b29507dab7c2a0ab6ec
z54fa6406d0a18abe6aee9451a35731379139498ce0d56794ef31cb5c1c8ba1437dd6ee867f2750
z10d8c6517d05270cc201abb2b52a191fedb7f47b4367572533bea4fee42c8a0b9bcee6966d0faa
z8a358edce85c91cd02c957997d17bb1da9a423c151c059a7dea28e048a1b31381fd1b80f9952f3
z603965f5284cf28a7af2c6aa89b2e553f3ea0e6f143564a604db7a5416b47232c65227f2c4b7a7
z563e899c0bfc4207c9aa26e5e06284f4cb9dc7495bd7794bfb61ad00f0544a5149da66ac2d8470
z557fa39b43214b10165fc691fa3d6073dcb5a75d4e651cafe9c1a43bc81e0ed969cc384047e3ec
zf29f91448d7a73b1146fcbc0713899a0f976aa1fa7a245f8a50f24dbf5d5b80b1c50c7ce98dece
z41292787ebf8327f7e0b3849b77e8b6a5e79cbfdae394b5881f0d3124ccccacc781c9cdabaecb4
zda3d965423ca1d8a74d9393e1f4af1c0a58d248d1b0b9058370cf9008f0ba732ba68ec7a7b7610
z2215183524a7f657475604575fbf7ec29b379f75b3bc5a242980a621dc347388a0fbb2e32f85e6
z1c19f020b575901dcaeaf8d4a82e89a49e6e4b7edd781c2e0d78e3369ebde09c6856ac453c1bbc
zae9f31e0f22519f22605f1cd114a4e3b6d3a43f4f09877bfe779768b347ddef521e502bea51ffa
zb59a53dbac2c6ca1a98a9908fa3cefaf3003709b2a75eb8fcc8831a13d37595c105a8556762f49
zd02353349b25cb1bc35d401c2a87532c7f10455f5c86fcbf7b307254de96bcf114d0e90650c374
z0febbdf136cb0267a9df504fe36c7ce42eef29f7bc4bba5e6c66c5050124da6e77906c5302d755
z8d3a2689a6dc143641c8cf8109b04416fbb4b6404f662ecbd20339c9af75cce88a5d5de3659953
z078877ac39513505c4c1bab3d2a9781292bd0e91b75e856b3b2c63b6b6b815c1c79287c6dd3775
z7dd971bd2dcc14e8b34915601d64ba1403a465ca976a3d5c2830c8e76e0d9162ceb1f0bbcdefb4
za7cff1303a3c940c9fcb218aa1dc5ca612ff0bad63c68c8d2d3cad038b72cf73d365d7219067c4
ze92af7077396a748263ecf9220a2532a9a3abbd6bcae84bc74f1e4af0f3e2858df4554b54db570
z32f71998ac6cc1ba356a2d4be8d1c018688f660c3ffe9d1e5d963c9127d9a5a109f2365b91ce2d
z92b9efc910fda526b6478c1a3f9714045b0c8edfc88bf13886a1caf93fe75e8f4cc6fa26f571d9
z04af1e4f1631e770e1c406b1899755fafe0c0a5b8da4397fc7a42d06fe738bf3cb99ec9243be8f
z863fe5c94344fe9fc6b1645da4895d4d44ba7957d7aa45ed082b2c61571fb55bf9a8d655bad68c
z8492f71eb6c6b96030ef85ee41ae80459165d1ad92e7ecef2f52e5b0f140c8834f09a8a2a139e0
zbf70951dbe4fb721b4d25e8625cbf9320ba111337b965925e4670673b5aab9e0a92af2d91c6bfd
z776ed9081848a58093f570f180371fda961824336927fdef021ec3fed75546fca161de73c837ac
z9ff8e25faf73dd985f26fdd13d63645b0a669f376d778b9508b1cf3255c2d3681486863d8ca510
zb9a16aba75cc69647ad0b7c6467e2e81d6e17875a8fb855dc6e2bc70e954a0db4473d07f5b9463
zc722ffec3cfb8a277cfd7d5fe17c59c9290ada16865384524de881bce3ba48d5f481d173e36e3c
zefef078f8eeffc47d7b0b9f0ca2a4fcb8d5f3aadfa0676bb7c1dd13a2af41af4ea080c12367c63
z34d426edb0db4dfcbde9ba27d539aa53a13dec12a2fcd05bbf5157923164abc77b31ceb982b875
z3b889879fab04ee9e2e7fb494a6f4e3c23bb99cb80987901da9773c3bb40ac3981af80284ae7f0
zab4639015bf3935355daa0c4cc7df912a57160942c24df92770058d43cd7698f96deb73205bccf
zb91278edc69d127f9c8451f32697f7f8e2ea6efdf4db7ba9d15887dd41c281e9540b46d63e1d2e
z6758aeab8541b22b8184262490c2ac38523e373cc3515cc0b9e4c5bff3aed72e0aeb46aef67a9d
z9f12760b9b78836bc8a9803dfdff8a219ec5975a8128fc63cc801a8656410a46b17213522b5309
z5ce483bd2905b53a9c70c7c8d642574226d11a40491e23a14bd969356c7449ca34330305e74552
zf88169361452e1cc4a718aaf42fa7484ba5e573946d12c2c9a5201dd9e5c3adec66b4c2b5dff66
zc66fb3e71d1574fdf5123a7e9d5782bc212428e4e3dd29e8d7f417528ef56c7ebe4ac77b134ca0
z1cbe034161cd3a1216e5f6239ea997586a49556b5e7dbcdb13469124482a2b6107157b80c560b2
z31bfd370bea76ed0fbaf12923f9c679c2ed7af4dc6652e7e4441acf6d1764c9e407d029717f63a
z3c881f84ed354be2a4a5adcc40051bdd01b32bd551c0645cab34aa282e950d81510d4e51789bf1
zaf00d0147b539f965c6e7b31adc5f694eacf9417a8ec3c72f30c30e9e95174a0f02b005afb745b
ze7bdc72036cb6b02095674945ccb878dccad2d8384b1101262648221cf3a9f5468be3327f0452e
z132908ef3d5c3391a2514cab0c8507dc07915b738b397c2b118666af25b2a08285ec77b01f7122
z7031dc126cab5795c26481bb7bd6b20342dbdd748df887242daf43782bf82b19f56de609e9a693
z75c6569e7de71b44be00ae0c6082b396919e3548bfebb6e0179efcd05ee682c44f2e0fefbfdbde
zb529d1f8652fea0c58fcb89b49920d4ad7c3b7825c8dd4bd7a92b6cc8a6a8ad411b4cfdb5e6fba
z4691d1c3237553a64dc1b687cafca60e0c728531d4703159ed794e84a3f0c3dea83baf92adeadf
z5ce080db4a3c206b29d289d4d7e4c5704ace66e5f73a22239c7576e892d2349443ca51580c6c2c
ze0c288abae21d273269f54b45e3e38cb6eec997b2fbdb481cc2451bd9ae85d588e30d8b093d11a
za11d80ec99b19ca20bdbafc267fa4380a9b8a7ba7cbc699cc045ea7f0445248c3391e999e4dcf5
z2f92fd0aac3660744d8b2057140b371975e21fcbea67586fcf3fc9d7ec582a1dd7ee48f77ff4f5
zff3a9750d70777ea6e33961d90547e795c0514aa89a93f502b62a13d6168485b0a93ddc2ff6f7a
z7f86feebf3f873e85f9f64566ed60310a0f2f374544afd2ad730c7f52e2734a7b8a24cec8fad05
z0d4b1bd195ca27c3c7fc720489906aa743baf9b6a4dfa9efcb785d0ec395dd8bafe273ab1f6518
z93f756b0c1cd29a7a2e40a460e11088d8b2b44735eecb9a1717d0f42d8f7a36db33ae6d1f018e1
z9de1ed7016c78ae92feeade019ea442e78f6ef99a0b938ebc8e6cf28f5ce44ff790a1c2a405b00
zfe6812d2988695874d27c726d75ff8ab9e3c435dfdc64cb80362f8ae7387e8333ae7f93a402e85
z3b5fa3a6462cf1ac8b605f7139ccb16338407f02a8920a94cb772abfd569c5317abd12c863e33d
zbfece47b6c5c0df4cc7195dc2704a3b7d7100b5763dabdd59147fe79aca59627ad2c97c756bf3a
zbbe7a70b50444981a26ef33b2b3b04aba28e66db1fb60ddcb6bf92d8359437f9fcf7fcdc7c1091
z74ead54897b24f638414b8f2c78b13c5c986d3b05517bc3cf77076e3b680d8949ae0c770164939
zbc723d8f25c2da34c9473957726fd1747c62869e1ff40445addacfccb9110c85fcc5edbc1a1093
zc33e227ef30546406d034d296ed4fe8ed9d0eb3056aa134e1ec9c421f9704bb51a4d13e0be00e4
z9e40d1c3b390f9acf5948e8d889ae91df6f777e0361a63b73a6785261aa1f63a8eec5a9065cb78
z91244f6387497253886f2ac07580833686dc04c78210e198db4874a87d1c61cbd5544708fa3cc4
zf749a97966c8f01d6a02b71465d63b23aa601796f0372d2ded2f0009a75c2ad83b7ba12778276d
zd2f79bd8c5fde60330530773df429cd2147740efe0306e70b43b3b032d5e5d1ccde6263b85ad1c
ze603fa01335e2c824079227728a66db365cc275b8ad629c751bc569ea18a6c4134241546f47bc8
zbdcd95b26a52f8bf35c48075d9d092b6e00208116a892823044918598d14dbd117612458a466c1
za247611b09a788fe892671a8310a661156fcf2f15dd48d1cbbd92821b5534a493b00d00978bf76
z145787ff7cf1df376cfc25b59356f05082b412e519942bc88c3805b42c2518f7b4aa7955e46247
ze1efb553282186271cc1144a84ffcf712ee090007b96919fff01524d3161dea785042eb1a521d7
za530c9c9286247321eb8aa610cf6ec3f4c9c5139e41a753626db51c0d7b6890a68ca4c6411e028
ze8d736a6ee96c432b527e6d177e5f7d7190f3d5176eaec8da3b860817ca23c6d2cdcba349781ce
z87d566ab4d7af2c876e82d36659d24ca90b363246430a651b3fa19c5f2e055f26cdea985a934b7
z7d0b4cca788394621d26857564fbd942660be49ae68a7824ad97762b6d510b199e0864aa1f7b63
z664130374fec13bb72a04618739fbeb472afbb0f30ef246bd02deff76653e453e9f3165db6faa9
z2ba1d9fbab358ba1e9201e101f1d409982d525c0fbe9298563c8582f4b3e77a7cce8a386a6bc72
z025b45a7c128deabba78877c1a75620c7dd96683fdd7f1b9ac0e0fc0730f3e982b7c9ec0c92835
z358a87f3aa72b8c16181839b970decc55a6dbc6ee693c2d68b948d69bdd542253bfef82c3eb20c
za95f8ab6d3657e0600a2b35ec0dcf8cfebc8adde7c5995b7686c1e7a82d77ea00a6b33b03e2b02
zb3d4642ed20df76aab2e7c8994513ba57da4f820e2a307714ed62fa89cebea9e893bbef88fd0a1
zb52658595464340b0e6c7b6eba2818814b8b73c51deb79ae84265bf1175ce3fa1fc6c0ab71c460
z6c8e40e11e9b2fca914392e70c96d746d589ca8618264f55eafc6cadd5a90ed8de0ba30f6b05ce
z6b8e524afe7fcb599b63e1ef7acd664136dcd69bbe672171624fa4bc37f631b4a461c9f0793288
zbf4d47fb335baf8cfb9f0427f8de46de592a6b1423bc209232af1ec672db9b77c76bbada778186
z8f1af2b4957eaf09e8f4758251924c37c7c3138561206b28d5df4108b98af0a53668f199c2ec4a
ze2a5ce703475bc95e86eb036ae2ef1c626ac0070164fe85cf70c9ff8cfce684a7a06d513353b65
z66e80bbbf65f8247b81dd141d09b7c8de6e41b7f5244df3ca52fc465799688cc84760d1cde6fbe
z4e351e048daa4005b3d17a620c813a4942a6d960502b749c03d90cd36608be6b35da97dc5b488f
z3e244991cd8635463dc2fec6cded0de7efe88ad7bbb7e2ff615f9aa74f8a231e1dee1b04523cc2
ze5db657f9f05dbe46ce4fe908af72f3b9cd713f3f4b04082b0baff646e9df73fe5be0d0124f9ff
z968438b92c21fcfb6834e0c36e2d639232952112d4c4b1d34efc1be2a2cceaee1bfd5c6b2d2535
z4a8d3c598764a25fc1674ff11dff3b6b7cd687fb2e0aecdae8f2d47aabfe1e562084f2934073db
z34f59df2bf44976f921b78aff0633ee1b639b1b5469fd62f68e1d5dd34d14dc54486da058acf3e
zb63b1f32955392f87305807bc96cc67a1b9b0bc6e2d6908e8d5875ba190feba997e3b55b98a420
z3576dbba5ea02b0a041c8ddb907d4ee7dfdc3d2787ca673c32e54bf983cefb10cf15a2c9034d30
zfba51fc3f9129118c34322b17e095314590f808c56f58af51a8e00af15adbf7a4f11a8ad8cc355
zd663573f24d10ec1942ae2476356fca5e58bf9315018d91da2e8773090745183ece3d5fb80c82d
z88463c627e6f40f84acc98e6077800706a6c2ffcac468d6300e394e89850076458e1e5aa606fc0
z1fc0651a391074760343e2fcddd9e9a0c3a57bc2fe09e57af9cba62e199aca7e3a9006ef635dd2
zc1c3b929bac6bebe60fffe8a8288a9e9122c22625e00f3b282dc8cd2fe88cea9cf45e72e1e2766
z5d778ea70f60c7ac81b529eed4700e5859223f4dcedc8e3bbdc84d868bd805ee7a91cb2f5c10e7
zcf8a8236f0326dbaf53bd04652b9402d257d6f79318727d90c44e3533a8ec7db52c2802a0bcd1c
z740b2fbe66f723e33e431abb391c9e73cf5195a20f340a7ef99aa938369628f2e18114917dc1ea
zd638a59a3e4bac8c031ff8cd14cf848631d181041e0c0f904978cee2e775736dea7d510557ef55
z77e2def3ab371821aa630a5f31e9c835eb7de715be8109141cba7cd4a77a782efe54f34c2e3d23
z55db0adf5203472e7299766c320dfd0cc309f82271a4706d24344dd4b3671dece22aec5a1cc66e
zef7bc329614324f4b73c7652498d0b5457ea83df9900f2846f5db5eb92838136f098c3d3e79d82
zaddd7d43598512b2e7849121c9f6c4382a2173f505091e6f8cbf6c461db250f66732cae9b06b58
z89ec54adbec8cedddd28b3c13c0455a3edb937642adf7921a25c92c251c37f1fb415d2d9c204ed
z31bd17d7e10b8131be42b510c84be23de994ee74a888d7ad22af1077eaec6016b815bad2a59fb6
z01881c07a4a145eba184e9e958f678d92b11ec5d6cfe787b5f5780b3b7ebae02373688307e5c0d
z0b149f51d0aef765db45d1ff09045482dee488a6739526f039731b504b40319dfcbce60f4c5cba
zf4f63de6047a94a19fc450fc6f509a02628e241d3faa29c508a3eea6c9db91dc2d0804be5c5aa1
z8a741922e49e80712a1e4bb9339874af6d9b5c2ff73d7043e4628a07a458090433e4a2de5b9282
z38d6975bdac2c92466c61375961a93df991e69ef8e69e9e2d2b485b27c05c007be8c121cd2fbbe
z4eb11d0fc71fe7e07bc8df2888c94333e1cd940b87b31d7b36802eabe4c42abe603482be310991
z372c9de81a31fc6059af2ccd7208dcb90d8de68537f7dad0cd49873fc0e59a20aebaff7c817e26
zbb19c31173bcf8117c981f18cc5a26632fe7bb4a802f9a6a693f3181547fbffd27a66cfd6934e4
zf3b5387f67904340f41a1a8f722b4191f0344cdd662011652157d938db6c73f121aff2d1497c73
z8e8f7f074b41144b85aaa50c4d76743f8e983ee6e41af9585e1000634b88dd26ba58bd74fa0bb7
z67e8ee6b484ca0a2bf1f3528e01e46d011472f65fa3f32a3e69f0d02489be8657a86f32f9c3cc8
zf30d68cfe18f7433d5896875f01ead2b343a90e64806382c180df948daebf96a03c1cb168684b6
z11e264a7ec9f3f2e592c6960f53e22164d0ac3e171feae496565afb75ed2c0ea3371361471ce02
zf2a077626e7f02caf8a2bbc6c2d563bfae3f07294fba7f964dabb748ce91811488bacb4c206c2d
z5d21a83d09e139cc232f98f1db60aca1527b9b7ecbfc5d06fed06246a14b6cf392cebbba69f827
z98ce09ce0cef6f336044cf94ee4b3a6d35641747348a9dce1595fdc00ca5f700f5dc154007c723
z532500becf4f16996ff6ffbef20fd6b53e83b60d38307bdf68f8054c1393ad9cff1920127be034
z1e98de4e98ddb411c170571b34c54ecec6247e24db4413363d94ee9be85c053569c95b0c72704b
zb780ae18b5056598962f3b213c66acf94809752ec73eee30852e723ac0adfc3ee7406d58568286
z5575f45ee7c13cfcd7ff29b578b396764c5ae7ac933e8bc24d5130fa5fc79bc9f9cd85611c77d4
z6cd66798d11bf80e8fdc1936c24baa96fcd0508a70ccf792e2994b512bf955818c0e05a9a503df
z14ff0165a7650e793d1eea8b7151cbce0a931c841ac04714f12f6a62f005a0caf9dde572514b7f
zcbdd31caaa452399e8a7ab9543867c46f46fa7e0db813e4487750aff59f0ffa685989dfaa84876
ze3a550c04192bdb70188ddf3bbc67b238feea345e68c07c7a3cd3baf4634327f1fd8074fb8f79a
zb49f394eb1d4982527e86043c0ae846aaffdc671734e3225d47c136c85281ce4c34db69f9bf245
z28ce13e555435ab214356a8e2e86536d9cf40cae4335795420e5b44c76129d2e7bd203fbcb36d0
zdb81065df3020d1324d7e7fbb1938eb55dc83a881bce12d9615aea74aa8d92374f252886d1dc49
z3ee86ee89bb4b343771941a839fa8761bdca03cddb8fb8331728d9299c5ccc56230b1fab54137c
zaa89306cf15d667577d9db004340bfc18082206892e01a4ac5854bec848a06c7fd4a1d85767518
z75d029afc69c8299c0a92c28c25f3f87ccd3510f076057c50b888d970d1e9f4bd5c69038c5414c
zafc60e3d26427cc48fcd1e7cd2d1df876a537c3b4c5f7b16adb240b31df4c1876f3a258b232e5b
z4a7b42ea59b91e33bd5b69243439c35d4b6abbb7218aa0793ab7da68b97d76f7db56f12669b3f3
z9de1fee3710f3dfb303f520fe3565eafe3b1e785b030ea68498146d4b88315457b92877e35eec8
z2f8d7f6be01286470ab8b5f272379707ff2fd53b0236344ab58f10cfbd5e7c38dcaa0a97bae2b1
z75bff1bc1bef980d58066b06ab89e33b04bb77ba99b3de4b63a9abcdd2b10eaf574619932a3bf2
z5914caed85a008de4c6c005f06dcdb546d97af845e206e9eb5dbd1fe8fd9a53ea1087d647996ef
za2d69e13529c65b38d8d502ca3be41657c17cf0a4b3297f91f0af2647ee84249386395b6e597e5
z15344ef978ace202f96abddac46829df0da3ddafd3550da3478269a091345219c8f27e5f67be06
z736434510647ba8c3517eda9ea0f8a2adae21c4cb05a33132c10812bcf12c3e889795ae07f09da
zc5a34c873a7f5a55a9cbf4634f0d8826c70e8eb8af5b6e3cf15e599303c091dc7d4c80053f1460
z95411ec443de06cfaed816e6c77a262b1095169746a2f8aba84e7b0052e9f945962cd5d482ea9f
ze48e601090bd6c195b20b122b09479ac3ecae18e133808061bff8a8ee34b56ff89243db3a7c0b4
zfa5a238ba0c55bab09c4cdbf8ed8740fb4696a9015d9f50e8f96f768617f35f6d91cf4b9f6ad94
zcf9e4cce214206d64c113537d07ce70c98bb90090c9dba8780572715f940b1c1f182bbca4908bd
z7e1a5421bac5a80e7cf80261d3c0949cdc670e33201232a4a701fce6b0e47d1b4d679839741290
z57bfb6cdcd197a2f995c489fadfe1ce3f181916a68eea4c2aaf22f180f5c64a417fd245dd6fd47
z940954a8f32d3776fae930b23082f2aa8d0cbd72b08224932b823fc4c9c4cb24e3f3da336906e4
ze98503c3adb9bd4838fc5c233a6006f3db8b056229f7fd5e91d054596c62ac0e4cdb05255207cc
z95b033db9707913a1176ce325af97e36df79523dd994f9965c940d4394aee95cc751524277c2db
z2d1fd25b5b930ec3b81545c5eeddab70ddaa20a246a22880d3525263831a9e15f08c4571959317
zd325d936baec95ea16facd571919d40bb60ae63ec1b19f3d85c185b5ad51dae1b1c6d6680d0443
zedafa598e454b9475ff89418b4522b81201b9a3eee1bba5fd612767654a562f5cd4c279adfcda2
zf76b7a267f4928520a76bef105803934168d19fb0b12222b27a0dd588e79097424ecba8b782dfa
za8a82e1b42c7a505a3de00781151b5ce7c726e77f46ba7a0984287c8c6fe37ca0b3df6593368a7
z75f73477a122107a4a3f0ffac7f52348466db3f4fc6a0e102e2f70c884e90469ca1c921749b329
z791965f4baf32a4f44ddee6a82942ea7612d1f9de78a766d02449d1c611991fc7f46b6040225b2
z9863eab04d01d3886d020091954a70c09dc2817f4eaec7441f75c88eed04f2d12a5e48e7596b27
zc3f96578e1fdc497e2aaed30e82336608a5c8fcec6ff2d9b5ea15e451d0f2ac493c63c9c223b50
z8fb8a2f08d55a27990b3d3c99f320190aae94b19202103e89b4a731834055b45baa2f26d50f169
z87846cda8bba4039f099d8a84d2bb9b7867d98b3e9f37719ef75e9ac796d9916304c967e998b2c
z3086d452e475fd21ae717983fdc3ad5e582c879eccc92508e929fd0e0ecb65187db55a15c85d39
za502671b02ef5073f9d127df50bd21e8029131b4b7f43d060e361feed8b6a8c6c0dd844a05b6aa
zdc9496466b158f3a9ab8e08aa1bf56298c4cb55ddd687b5c28946253a92b6508a8a9470c50c181
zb3e71333abf7858909e33fd9e58d3f17cabf0617fe8d5b5a00d85248a8713f6af9dd44cafb90f8
zb5b21b4c7dfb69a831cfef83f7ccddf093f3039f33dd5296907442341e3dfb1651329e44d016b2
z70288df70403c9a68aa65aed731e8c09d07a1be82e0f04fe47428c154136b20abaa1f343dc7039
zb71ef4a1f34e7d6afbc6bec5e8e1a491585779ccf2f7916d0488e03c9229367b76ce8532d2ce12
zf75b7ef36ddf090fa71e2382171200e6c8ba397321e0fed2d0f24e29259519d6c277d01eb8b7c4
z8549c75d6fcdd8d2b1bdb9f51a252b16dbcbf4a96b0dcbbef9059399e0ff8571ea73e61674e4bc
z72cb9ef4138e48759e5e854e862e9803fc5455993295ea3016977f035f8e75f8c00ef679ab2bb6
z12edf093298c66af6b9d099dceaf0da18d4c54e104260854fc90f9522928be240d4a8653d04ced
z5e928a0f7a519108807551b9847ed11e038b5ae76fc5ecff2c2a32f830fc807792bfbcc773fa65
z8866ebd47dedd1fa8ac5b6c565308b3997cb52f1c7b1d1f0153b6825a16bc600777200f87d15bf
z18862e36a0b86e97cbecefb301d4d574c0cf359402c8b2c7d186b42c0127eff0c84d5c5a2796ff
z5f7393e0b5204b0ca5029b5842616ec2cfa0d19a00d019dfac96a96620cca3eaa886f6d98fdb6f
zb4ba27a4c6c7c5692862729e001f7b43183ade5f5770b8d2679eb41e67e52815eb631bb17a1fc4
zd9317ecdd0df914885d7f67169f0ce56087d2d03efcd38e585b8a2463d346064dbbcdb8437a580
z0469a2e6bb3fc380b43793c670c5c5cb29df2eb09a38934199ffadabffa798f1a7c286461e903f
z9d098365fb21ac7c42f9ae03d7607ee028d073756708ead3271dbd4475eda3dcc60c05edb849d7
z7ea63f87ded5bb8f30d4ce723b1b87b7d2d2a92702c9d7c3f15a74b94ea633f12a15c6aeb7018f
z4abc9f4b2994d51c428c8727349a6cdfef44ca11beef34b2aecff2cdceb0180f73bc47b0587442
zf6262b73b6d75eb27ba8b1df15b768adf92d284656841a9765322be3e79d625acca8a762dc262c
z255809a32d7099c45c555462d574da5c77a7a4d4d89a7847458b68c331c6297dc149fb6031b9e1
za4434dbfdc4af3ab63a0861971e4c87248b5581b4fff7e4580382d83b888e775e72c5eebfb6412
z01629af5ef258381f4ff59184e9b07de4bff74d4a68c09ba7608f7fadb754b0aa15b2c7e90ebfa
z4dc54377aedb6c96754e8dba3979737efc77ebfe9182733113a1cc616af71370e8bd75b10ce15d
z726c6cc5e81685e0f94d97ec7795903a1cd4f82ddaaff2cf28f689c012b997152d3f827d18f7cf
zc8ae64b71bab6a947bf5c28a214da2d5c1917ec793963c9cb4af9376bd3b7dff3a3a4476c3b1be
ze05513570ba7c22b475e8b4a24d7f93c7291829553a30cd29cf0def5605cf76eaf2db0edc1e556
zf8d83510acc6a61dcee36e58b55c42f0ae1e21969bdb29b3b6a98f63871a1db36b83e196d86a78
z7ad1b28d2f78e8d39a8fed988c2ee166a35625d5877a034702216dd8d59e69267d693c060b65cf
z84b614412f12cb1cf7fabcf9990ff4d07cee393b348b8ce761f76dec69c280b1cba7c1a3849346
z1e01e52d96516c48981671bb20f6a638c45bcebac79caf18740c17fa9c7bb542603502ffb49606
zceabea0076a846f19edafacc2b07ecdd0d58e33ecdc85633f924500c10fced985fa6d47b2ec20e
z41741586203e85a6bb6980db06a0d58670ef8b7149396cf5e6eae5e0cb284bf8eb590887bdf5aa
z76966638bcb2a15fdad93cfb357010fa8b2c6edf39ec06f1b9a8e73978848d51988cb71c25725c
z9c188d26532c6168f6493e2bd48269ecf81a6aa6fc660e7862ccbbbe4fcebc6dc7fdca7e6d71bd
z18cd1dd986b611f121da3e33bc141a17423a45934c0d30838a847d37f296172155822267b368a9
zf1e03a38d2efc00effeed86839d76bf1a0d674aee851c8a67febba81129323ad8b405fd5c18c1e
z95236f3b5e83e852cc7a40c838c456c5e6024ad9caa1044cfe88a441efb7c351390394dfaa83fc
z8b451451e84b1c609f6639b67fb3e9438bab8b5db48265fb6b1849eb4788616191485f942fc9bb
z21226ca9e61a48c06b4b246cb34065f5a0d471217fff76966a96bafb177042a6bb5b8f786a8491
z6d5caff5f81ff04e19d73267fff633aede06e93a25bde30c8ecf3331773a2e70c3df7aedf40745
zc0d765ddb87519a80671e39f65546d7be98c05c2fdff2e6fa0eed704652fb69090e6962fed79a4
z5a86d3b91889ef3f7438068891ae6ae6fc7d76dc69612f4e45ad31cd5292f8e77c691860b615dc
z327c1893da17a90f08e516bc710af48da83f522f5b48317a8f40e9334723179886006f5be57572
z524585fcb775a44638f88f91fded91084f8085199579abc3288c1da13a7113d5f4e0ad78cca9b2
za7e8c810484384ac80b25bd7eaba1dad84055dc557f7a76347eb5fa74a7c8dfd6bb82f8e14cc39
zf62fca4be1dddf2740cded78c4a3b785e1b3805fd8ae13c2b62a2b88994df39c2bb12e2a9759fb
z225962c4afb867c679d270105183b2358153bab1cf2a3a45ed9f53ae8a97076345aa2c82299061
z05364e078c53459e6aafc6407ec2ca3bd63100ef86c7a0983309556c9db9baf2d97a9ad9e4c30f
z0767c7d5c8ee62439d0398b81a62a3b0a88e359d6ff075982f8d139dd2443e3521526b89b5595d
z677d97e2d9786195ada0bfe4e02f4d4a785779b7b291648518bdb9ab0990d46c33ce28a110a820
z7bb69b3af49cdc6f3958ee11873184e55c863e47eca615e36f654e6fc1435dd9c415652a8b84b3
z792f530e5bb7f6673b6b73abb92e429a66f2e983c7088d82561f081d86f7875db471624f780411
z4c74296c3252a58fe7b58d3af110a50fee3242873544e8e3ccccb2e832820c5ec9b26847f0c8a6
zc4542232d7881339e56b7f02b0f810be04e02e7b49064309cf203b677d15e5e899f16bac3dbdaa
z7adb9bd9fccb2ad2fd74a91ec22ecf81964ec275e573a7a347fea1db7dd8d4535af01a9cfed158
z264f78b6eaed38f0e2dfecdf34fa9dec02fb0ba5e38882727aeab0b09f62b48845e88578c0194e
zed0ad932a21df4e8a193153a879f2bed8c5224
`end_protected_0in
`else
`ifdef MODEL_TECH
`include "qvl_sata_link_monitor.mti.svp"
`endif // MODEL_TECH
`endif // encrypted_0in
