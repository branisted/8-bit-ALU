`ifdef encrypted_0in
`protected_0in
ze74c34e226135848fe16db9ffd31815111b6d7fb642c521a3f628cf6da949865580b22efd062a7
ze90adae0e65e66a2c36a587d0a790699161455169ed55a01f2084f11770a774ec4c588039b380f
z6de9c5084882a40b79a175f5c2114b2b6d78b070cb806e1c0aa9258297f4687ab308bc470f0040
zb0b1de382961eeeaf2e279e1462520fc31c119af8f2b214846f56c2b3cd2eadbe4099496abff18
z15cec83ec4a77b868344aa20ba7360908f5c0de2a79abf8b3534b883bb12180f68b5d4beb444cf
z3fba8f13afb0abfe8fcc4294810f75afe452434d2d0f1166236c82f76edf1e12979f04bc35693e
z32ae028996dd85737a8f5adc1ebb94f39c940246e887647b64782cd7ab429b0544c173176cede7
z01dfb26b1f73408344a52b7e1f117f12bb9c8077b34876c2e6fdc085981637012dc9754765e1a9
zc512ce062e0b8fb16a214591f5c81e1353b900a611fe1f4886b57940b41b7f2ce99a7b84b04b90
z916f717e73bd10589c81e207ed77ec660a8cbed5b487fa50acde1b055c8870bd8676023f21ddcf
z9c98cc47cfa2d654ff1365d1f45035a045a66c5dfa82790502623b57a3af03bf0f0c0d35b51558
zb8b5f2d29acf03737a9ca2a053b7a8f06800d50b465c41b30eb585f62f3d0c2c5a43bcc54fe309
za0852c3b0bd58f0cf3aac613498510a35e4db2f3cee2d51014b82a03c9a823a6d0e8cd11021eab
z1102200ec8f36d3b2327a0603b2b8770891f096096346309f4f1d017a2b3ffa01df84fa816d14b
z07cb3fcbef3b7735151dc11b1dd7bd809b3c348e19b3862ca5d1ae4b442631670bdfae31a99816
zaa360889d88d5b36c892526decbc16af2a8597da60c30fff84d6fa04924ae9d2fa9c875fddb856
z0010f1a04d62db18fe34f8aaf6d443b944d34c954e2219b14c3df7845df56c34fe447c15649058
ze091bccaed25587e22cd96ad67150a8ff074f547b1442c3297ff604013e6e9926ecbd133a5b115
z682e9648e4f6cdfd6b6ade595964fed0303e251a7b6ad6562dc26b5e9481bca600d02a73046662
z7dc344b4208c942998899fd0756702189707c09754319a6ee11e9fcfbbcdf4e1b502ff3a17a949
zff1bc3586cc63876d55108efcda6b85c302ddd3658b243e40a4d3e2682715aac451adc5b519327
z94f0f39800762a003d2c46c5dffaeab18e3ec76367a7eb83d1c96407c873ff1cf0534e9f484489
zf2a39170bef66c1aa7a2d9fcce66dba59e9a1727897e69606d011a915412102a63c867901b4f60
zfb7e5aa0f0b0747f621d634fba4139075a22c847da9b108d98eb77eacb904109d23e3904a49126
z2da72be4e3de8ab500b1c47c4778e15ad4e3e23c74876d19dbd6bb7eee155db89bfc890b9d1ee5
zf52572d2684d16525b766292e33e9efc702bc1391a6b809e66e13d07979b89fecd0683f6ce7c4d
zcac480c62e75209e46813767d1bf9f86aeeb9923b1588743882c3d1eb3b5a32da30f20398df4c8
z1ff926e69db27d0762829c1124726ec9c1ededbc2ad3083eb10636d82a6a35b40ca2a36ee40913
z947deb2c115fa5ad4778f61089be357306dfb6f322c8292870aedeb3b52ee0c75503321412e7e7
z085508d54cf1085b7890636618593d1783dc84abb3a9f28b0ecfc787ba342436d2aa3e0da589c7
z027f5c20087a868da71ae97d067bf29ee0fdf11173c7daf0177c1f86dae2aca4e92d6364102cad
zf7b90552f3b9ab5df8a8e7e7fc18ba0f17d1d7a040af49a3866e0746371e4073d1f26c7401536d
za82da8e15217ce7b01fc4022e58a7ee0dab36868d1db4abf5650e22fc63a0f8b6f1ba24c66e5d5
zc641d8f8b5301427b4d3d287e720ed615f3e9722d07a72239725da51944168226e9438d04db9d1
z2d8820160b4900dd113f79f60907b972f069be5bcfd7749f9ff33416c9b77a72cc20c23b02b97f
zdcc7806d0036b1c00893dae089e85847732aafc3577cfe790558f76f5fb9adc11254de66de37ee
z36fa3e6a81bdd2215756e0c8b2c9c3bce6dcaa6ae9c368cc000cf8fb765bc2093f09795eefefea
zecbeb20e4a95eccfbe863e98dff7dc3061e10e0d32bafa1399121ea7dba368f1b78ca9052bdae0
zaf0e908e25fac5ac3713d10d7c0ce4d1609dde1b8df6fc6778f32c11e37d6833f2200147017a0a
za6702da8cb2891ce4e4b2575ffe7b045b5ff99b8b9644bc6c77c6bff7c6f0ac84161ebdef210c1
ze81ed3384fa69d23d0a90e85d3baea95b9f39f28c5d8f304d3d7c0a9e7d1dd40254d39a507e0ed
z85d7b836f4dd821fe9d2ec7eaaa34bcb549f440aac56b26f8bc6a77d69b6475b4b5bdb3506de04
z9270b182d433772f4f0f77ee8527ac7ea0c1887e2b81768eebc32347b112ff74b6ce2e0f8e8b81
z414d502db19689ff31c571a3dc89d6addc34841b9a918df9bf374a37f4989eee37ebcf40c4fb2f
z09b0433ebd266bc3ad08e478a5f7af2a1fc57234911fd52f0c5f2a98989659792748d967e68cdc
z58b1aa42b7dff4c25dee2c503ab61dfe876e31d25c204bbc5280b94b8669ff5568107e44f1d622
z8093ee3508ceca7b1f5152a68ee97759e11a12b2d050c0ad43909d99c0954dfa45028a36e3c22e
z55fadc95da5e44837fd24437d0e2c62793cc5701e65a7bfee6abdb01e944a6a7a13693a882be6b
z209076a76f8895a830482f70041b55da3a8b358aa6b0c34efeabb942d08402511f94e915e0f099
zbc4fb2b34ac5743917759438e43a589933af2051c6355d27e9ba69d1f0e3841ba24f09f818a945
zcd055de7419ac0d53ad40110bf9f10509d3b535be8064a8816d72b9613881460a03ac04efb757e
z741312a3246aba4578c10fd90ede5b8d6f4fa6c5fce12fceca08b4cb7e61817fa975ad448a3ea1
z6f01a424acab64590362b3611629c957002ac12e43152ed3927bb6d43d76641e7acbd43a306d44
z2cd29ac1009b80f3674736c0b848eb30005561517bf5e6f7eafdce826303b72d9233276e74193a
zc8361c19a1577e42f8501af024d3275bfcdb5a2a5fb497733807c3a4bc0acb0d6d4da4eaaf8458
z44dd31a1a90b2b29e6c92b6ea1570bca8ff19cf9abc1865f91a55ee135b9c4af883889ba5afc35
z136f18df1e5c5e7311dba9aeb8722f57c7984a163ce6416c577d1057d9e8e7a1b6f269a923adb8
z9028e04688f4774d3c8b3fb378151c4d1015673c0ca6e672c82361c816ed7b63d13865bbe37f62
zb57efc11d5669679480458868bd92a37c41ae24ad6f33017c8fc05007233674b402e4e99e84fd9
z84d0b3e469d1eee22b21a932f1bf81d0f7843dad12a6fdcf72718f6189de5bd452ed22375bbb34
z63046f34049f14954bcf7b16003b7a3f3d1cbcb5126366684bbf827b6fdd380927cc17ec02575f
z55a293212af8f28da98e7387da12e40a7da9dd559cbbee8f3a5d67009ace29cc62dd0c8a31e1c5
za0f6acbe0e5a06669ca5b028af24094a95d6987362920bae3dee40127f4ca417032bd69c90321f
zbb2d7665c1b1a045da1a893abeace61f7b75fc70fb025dc01a095e76aa92fbcba27a3b461d2e5d
zc678021684fb4347245590ef4e0f488e104c8ea046f92a327e1c191fe2389150e8e0ce42abac97
zf3a6cb869793a2a14929c4d4f7665279408723a90b3afcd67c06a7fe6cbc9c06e42d9451560dd4
zb347e0d76ff155046aebc18330aca480a2b5243ed2b91ec001bcd9ec7c4752824cf63c85af9101
z27164bd32c5e6ddab0131ab6e3745a43540faa3a57830430200e82b1e3e62634a804adc05087a4
z01b1c3f69ad17eb50f3c70a4ea0f3d607bf543a1a60994dbacaa571b53a543f7633a17249cd74d
zda20eb344d9388cc8d017d1172fd628b670d567cb346d504009e72c1eab0bb034b732d1509cc41
zea8f7e5d14955a6afcdb2a0c1df147b7e8a6d20fcec57a9c4c610f277d5f660d25fd1630dc44f1
z697eb56c2b0b27f262d6d6237212aad32a7bf973812ae13dab725964d5af8b2db048dcb3ca7a8b
z8b0f5b29f6f98182a936e3d9d01bf4ca1d0b73eef1bcdbe592aa0a3bfb045f9d1ce015405ae9c1
zafae575b723af244e996ba37523c1e47614c0eecef8362c4d87bb5c7eec73df0f8a95a02e67c40
z0b87e5f50698418ac470ba709d95edaeb4e9f418bc54deda0018c85121c46422d0c53d2ac2be35
z088680b61d63cb2ee447f3302d4c684a17ebd6864f7d2bf0c7cbeacdda93bf48726700eed27ead
z259b37bbc9ddba42d26be37e97c4bd377e33704a151c1994c428c2561d30160d96ef12dc034e1a
zaa23a8b0ec68339c2df979ba152322e1d2a175f0d16ef30f4064255f0b28c6f02487986b3ba184
z09e0a96df4a873d98fd3003217f387bffb7646cff00cb5623840a218d948183fb7e6f757d06bf1
za40f8b7e6b260640e60a81b7279065c7d5c30460d991bf7abb73a853193ca4d7923ca9fb2780ff
zbdfe3c60463ded34141142eee8d341d8b4778b70ec105598b1d77897a29c9b5e2e049675847f36
zb077db2d4dd3e7577cf88ae39f58868a5ed69f170aa6a1139b366609c8f79e342e69a0af2f5471
ze64a94ac39862523b0d376d76e9ab4d6b34be5fbddf83b8fd54f22ce85e24ebecfff6064a3bbfc
zd7f5c1c4d1682792139a7811e520657d0367b4bb8a35a7a63dea5bb70c9c2609f8f6f7ddb63535
z5254e53b5f0d6b3f4ff48998eeb887493a828e77690ed2446db9a7e09bdffd80f30b8fc24e4872
z99df7e0cc4fccaf58ed1b10b012a457e14ed613e9d4dacd97d5ead1fa0bcd10d3c3521623cf57f
ze958b0d96cf6a79a19b31fb9d173c47d0a05622ab7433dd1cdb33dc36f2328f3aeafaa29056ac5
z42cb5723f495375b0953d4b0c9d69ebb3474e5f02fa12fdf1f9bcef2cf7968c4e672c52de3f93f
z9ae5938efb66c493f889374d11c2a290188c689e1535ef74890aee3e15e1a664c99ca66f629780
z239aaa9f7ac6500f65891dfac2fd146170e5b0fe7ae588785113a7d1ed2ef4c44fe4907f71116a
z192581460c6db9ddf42159929c701619b24020cb3f136f44709f8701bd9a045019518155f529bb
z4751600435e8bd019fbb86c2df90eddd4ef48d3c3924495adda72ad54b428fbf1015dbe6f59a30
z1bd429cddb7ae71a4f491561602e7054fe2160a92a25b5652a74f1816fa61042f740416e6fc02d
z4eab14ffba681e5ae04336142258d7988cfb1c71a9e0c7472660fc473699ed123d02c48df534b6
zd03dee323fb98e2ad0455ebf2f97581d8d7eed99b4bf98a5ae5f7aa51b35b5df10d3581423b51a
za9316cc65e8b4a6c77500efe8a91e97d2b8b996c9f475006353442b8f4442effdb2e8cdcde7586
z70e31fd938146a32ecb60f97c380acc338336c484f1a1eef06a0bf26f1ddec5ee81822ddffd8e3
z96d6b39e22f6e4f0c3ae5d578ed5a855c7865843f145f528a4bf6ac522026b6dac765969d61211
z23c4012d7d7466a3bdef0400e0590be2230761d5c1a7def7e40a21e359bcc4b9e45980f7ab1bec
z1e58fb19558600e67700b2cdc663c94381fa1584e6c1d9bf121e407507227b0acace8d22043b16
zec46aa55497d93052ff177a5c443d2833008c9c265a5fba8c6c6297b076b9f8583e00f0b434b87
z5af00322155768478926f63aaecf23ca5a6b4f20205aa4e739ba99223ad1a3c5fd0f2f36735006
z54622279907fc52669b096c666e3eeee4cc08e84bffb2424f4b6f765e382040689de1cff17eebd
zf54d2b781bd2a824a553978e6221e09f4f80b52c1ba687e15fed89a9ef67b7567469bdf2301775
z7935c0cf74ae45416d3afb3e4031cd2771bacf4c05163a209349ef8b0a7f17fa455012f59a4f03
z46c84ade48ee1172950e4c31d3263de3bb0d66e61a5afa3f391450d2fa6b1195f7d6f4ec8a2512
z5ed3ebfe75b51d2cec1959c101557cefa4cf7faef2915a02dd00103a1bb7e1203247afdfc3becd
z2aceafb1b32b647b1263d4ab9ca63bec520d38ebd06f15f3641a7c44122403cca581daad214e2a
zfe48eec07a19bacc257e33c7da3dcc8fd085ca7de89ce85a07dd2b0db5f62e6f2da7ec667141ea
z045acdf4afe18db271e33a5bc9802192d959e4ae1af6c70fe3623859dc6ac6de4c90ad36173e27
zc365de7ecf90d1aa61ac26a2612551139def48c6cc82f80e75e0f74752c4a8194bb647c0cd2fd2
z3a2a5daca18f4ad5f4bf2645ffa8073d9d3502dd62abbef0e4ebc1599a114a4f92c65d23af3472
zfd21e512a05f905a76412ecbf4c04a883ba15edc100198f94c7453309d5f56f07f774caa3e4529
z72e7dab5410dae655cf30af372cf69c710a01a46a8eaf728d6194f130378f59da4bb444d914798
zde1671e3d5abea12847d409c1025947de0bda920ef522c27107f4e66db660ab6956246d8151f06
zf80c8a03cb1ff54cfc707fbf65c8b5383634541071e69d8b1c47e4ac23889ee41340da98ca413c
z6bb746a7ef552fb571ca2fa555c00e1f8ce1b3ffe960bc945ac08af792956a9d8c6a9aa6fd7a37
z7aa52f095736455ced510ffb66cf6bf0583ea525611c4ac7fe75b43f9ec4b8ba3f90e6780ef333
zd5716c78c0ae88a214060511c391140abb033431653efead30cce58b4f7f63708ce1c82595201c
zd616deb3d969a873531034419f190c4b91731dd3a5171953e5ca39f1e936f001f6f8120177f645
z6a24798a5624ae9514f773da77faae9c35088ff431e4b049fe53de461917d2883d03ec46daae5d
z7512ff55ecc676dd01a87c701b370326dcd3a7a10770b506a7c0d922bb91957305dc543800bd99
zeed64fc3827e816f0bbf44c986d88752cc1fa48c55ebec4c29a62e2147b87636f37e06578dee24
z5450b18aff816dc57b81226a95e927978e7bc718da03f0fcbb11709fcaa03e6135c0bec5dcf8a1
z6440f9077c2523763510ae208d3897fcdec25e52d5f694ce8656b01af810c8ab6558a580638b7a
zdd3807153699a1f557e93cec0ff33cac375e29e74277c04374d921c8006b440910616a556906c3
z38be19db4f28e3596c1e6d6c5674cdf9486f1b860ad89cc4c29d5a5d53028f19b5eccc70f0877a
z8ce4d4fb22c78d3774b990a551dfce5a1809d33576b95b27c34d679863e6d90aa309bf6da6b61a
zc764aa133e45f3403d63fc72a94b41526437f7e68ab541a947f8238458223aa54fd0052b7371b6
zb6149278f35fa3ad497ffd50d59bab6b6fd6b8903735d11cc5885e2727b49cad4b42695c9fdc18
za90bcca0c6f41fc421bfab3f6157cc962167d88d1cd2ca8df7f16e19e4cd13d93cb83e9de8ec51
z2135debbcd82cd22c45354bd8363540d79146e49d83aa84dd23186d768e4e6cd3894de0655260d
z9d2d0a598439b5aac0ef9dfb11db50720247b00faa1ea45c3dce78fc809e04afbca58eacac5ade
z5f3f260312ec1227e102ffc2dee87d9626d213e3b0984eb574f018056d5c90ce6b0c433267ef31
z65e21b24981233c26fe7ebd99d80f48a5e725a7b6173dff60ea524190b926fd17cee45426914d0
z3937591f47f022383f5b9a7218c7a2875439c445998b2e65f151727d55f69beeaade982d674202
z713765fe8b31bb9d8e6c19157239ae0d1f3f227a473078dea8143360357c195b3e265808af5ab9
zb48e69c21f7b2123d4162b353181fda5fb99be29c07e47f59dee4533cdc5ea56ff141b1ac136f2
z60a13a3fdc73e52a740b3aa07c645d403bf57d2f8880bbe5d0a07bfa5713ef9c3a03f27c3c4352
za1b2c18dc60df3f8542fdbaf8033bb4980ac33b9ac3ae9e8d9b08c0f061af5083e7845035b2f63
zbed45a70048aacab67b859fe5afc230d388bbdb70b8ec08919cc63529704c2e96cab2fc578e5e1
z5901868ff99702c166236600d1e7decc61297cca1d119a3ef6cf62cd50b95cec29573dd4b843d2
z451dcb15af4f311ad76ea2f73065f3602e534a1e18f2282d2344ddc7a9b5ee1254e4e1c5f29a72
za4d0725aa439e7ca01e7f31b4cf19a37401544c45122f1a99d12d445a39415bd3f215e2c5daf5c
z95ac97cc71a5fd49380aded956039e82b5d5a783d1ee87a7ca5a6224b32589595fde5da859053c
z4c08f76995f76faf6bf30eb844f61b37fa958bdbf99ae6e86e2838fc1ab445b179638a000a49cb
zc869a176835bae53409101b04e259f78c49807eaefb13b5aa02e4271d5a0759818ff2e5627f27c
zec6b1f0aa86dfdddd70b0bfa3ca20579991affe0c941e6d3e2b8d8ce2d6650fd1b5dead93ae8cc
z3af6b45de40e899afe04108638bcca98aee5dbdc38ac12b87b2a8fcb9fa9a544bb8d1de7909203
z959608ff1ef5c26803bfc39a8c6ee3554ce492962c6a5cabd558443de345a7eb795be8ddf0304c
zf61a106c29cfcc29efac0dd60bd72f0127f678283cfc1b034d8ccfe8dbe138eaaf5848096f9246
zd8486995bdb248b5768df053900f82b125262e0ff815f5e8ac87c75fa5266f67e689c9279e13c7
z3b99c22e0c1f32b393901d5646656bc0d8e8882ba111ecf417f24c1cf446354cc07dd204f7e123
z503cc3838c2368cbbe2073fc20a3c4aff2ee9b60e55be5c43c110cfcb802decf2d3df3b6ef8cfe
zfd541e34bd272193755114ea29af54265c336f9426a1f201bc68387338837a1b999090666c9ad7
z0c301847885ae1936a09760f93125bf81cd60ea6271fc46e7af138c52641d352cbf99e95951001
z6c8ebaf854657435d251e279891cfa81bbed75f8c23b0005a697c60c0c9bb11ba13875e857aa2d
z66cd2787ebca76e0cc1b9cde40cd0e934abb2e8a42712d0dc8c95d54e749815809a0f69ef0b04e
z31b1244dae1de203e1f7bae9adbf19c2b4cd357940708e90363786c8d11059ed29288704d1746c
zabf084f83213bacf2aa5e7739a51adfb7fabe30a78ee69e05b81c1787f0f94f6e39b228cc27a08
z70eee9492f96dd6610b3ff961d135e11f0c9ebf91e41704fbf747164b001f5ef825402a2c708f9
z3d325ac519193f440d002b4c70c5fab4096a859c089253fa38833fdbd331e01bf07605a2dbc83d
z988917066987eb287da563a9e7b71ef5dacd854f68efd649d3a5ca1f059d61abae100888c6cb3b
z6077fce04323c08a20576209656c26f05b6ec91d20abf4dfc7ca9baf36ed7d012f10b91a52efdd
z712ae513a2e380aca7c772a22a4acd488d0e49a7a08600545c5104bf5eb56f27b47f2c8d59fca5
z0bc6a456fa96b9b9be787e86cc806b7427096d987c4410447ce0a07ba3abfb87ecbe24b927c411
zb6f9aef6e122f8c3987d2ac4c24bbfc48faae90fb422c23c22cd3ec4c6bfbee4f907afc8db150d
z31712db295795cc5d854d72bbe089177a1cdac89d7fe69c7089fcf7291fda740c91ceaad176a99
z610ed0729c14d034bcedffa6164dac2b24d7687be4a37eaba3daf76eda00e9b96ba83b49b61a37
zb8dbc5e6dad6a2f80ba794450ea4d9f34a560e866ce2748227a1254fa1c2da571c0c6aabe762f7
z196e265e971b2236f6637175b6b033ea8de0469661112f832b2fe7a7b8099a2d74e8330db230aa
z9816ae473e292f000c3e00d76806ce51e878609761de53ea7ff393ea2106e642fb1868cfff429e
zc9f33a2bdc233d1c7010ccfe7cf2123d976b1a3c1c9bd70d7ec78a7d14ba5da4c8fa9f065f5a0a
z9c674e29f15419dfde21bebfee81233b401352a272dd550e05c55230cc8c8f985ca46ed4bf5295
z5e1a7e53cfff8b8f3470bfa41bd25d71becaf30bfb4e8cc9efd86d0c1d87e1ce542969076a3d85
ze931ecbd773cd4b97661f7186c4d7482302f88cfd6a8367e26ca9d8346cbee0cfa01323c90408c
z4bd7d6349f61448272f9c007e36d69d97c5b107ebf3abcc5f351e6a20f5f337cf3d19171e8566e
z36ffb127bb1f9d9e4b46e7c0adb97691f89d0b7a7342b98e7520e074357cd15aef7f1282921a53
z06ed91cdd89748b2a973bf51091821aba8023e9f0eec2ec5db5dd200e6d73c9c326e0dae43c6b4
zcb976729dfbedb78074c88f7bbfcb40f3990bc67fda3c9d8f3d80ec6fd3b3ec515b6c3cd023f52
zf0b7a755ac11db6643cfcb3fd8a21255c08832615d4269da1b67ff2b5162d3da9afe58bfcda90c
z06174a47ca1eb2e56f432f1606c8d79481c55f163d88ebe7dad2beb7ec66c8e6e6a20f1be0a9f6
z33cb27dbe7074c944dcdb1d9596f56c8d2d7b4fce5d9443cbcd071c8ea05e8537ccf8b9642fcac
zf7d0467c45a5d13c8868b1ce2cedab634ee3d5d50561e648d95563458e44ce01651a2470570dc5
zf468dc40046afa5a499230c6f3e0b3063d6b8edf54d1aef5b4149e1ceac4451ae7cf1325277175
z8528e47f9c17400ffe212251e72f7fb9eaba4473c37766617a9302acc27c22a8df3657b11ec8fc
z9703484679b7f7b71da92ed9d3fb7083a8812071b4ed1db7daa34063872d74981cebbac2aa51d0
z81c7069bb5d1e6700024259e9b36bfc4bc952ca063ecbb10876c1a76ac8ff13b666f31a5fe62e6
z609e141c7246e151b422ebff79efbb2d4e28a39c447df01fa51863684cd12890687d6aee45eb7b
z05d522b6a268d7c4ffee1d555d1aa16ee139e211b38506c27be63b393cab43ab870fd7092abb66
z409853df492a370d33c721d7523b38b6bbf8f05442f3b293859a08340fa7310c9b1f97a4bcc1fd
z1587b0e41f0c1369ce274481b37caa5b5f0e5da3833700a834da8764550e4022b5e54bf6083f6e
zeb639c479ec64a3366c33ea26c421a859c908823495a4125e91f444b9d0c6a1551c72255bcd0f5
za21fbdbd27842063851e734e5be474b731fdb2941aee091a75975a6bc535e69c23f0c3175bcbd7
zfdcb42854602d5251591d3beeed54a35ecbfff431ae0e5dbcd350b552ec002540d36d987c7b3af
z553b6a2d561d01834a2b3cbce33ff4f38c2d20a899d66e840d8544d8c5f504cd556bd061209bdc
z77dd7fe8fa8a77ce0e4112076221a3f5ba3fc35bbd98d2118525568a8f5eb6980ec466a2f38db0
z349b73161816dbab553aea3f3207a671f88738b989610ed79cd1a18ceeb88a7d4d14530c1e4e38
ze2f2cbbbdc2cfab5abe2e72fecd973ef11acf58207f546e2312af20a67fda62a30baabac3f6654
z9c9d0858a09b65589b73cf281d3961b952738da9d6a0510ad1af0db78fd43358d6973ea77ce5b3
z5c269c644e9f22ab30cb9e44e1f32517ad8cf99a25e272c08be4e1a3365c7a196564a0682a246e
zf4246bf78cdc8d31f1242dba4d66c461f8b6447d4dc83877f1aec23f587477357e380c472caf92
zfee8196535bb37621db8d330cc5e36194050c1ad2dd8f01cf0de9be0ce19816007717b344afa26
z31086e16d78ea4e9847bd4b5b1f3d8189e26c6701c7f219f4414a002a10369cda9a13c4a9a6c5d
z0092d005ec8c77bb3de3abe526e9d5b65001cf7e3db08776bf54be0db79b30996676e52b8347d8
z942f45a6b079fb9ef65c7f0fba1f0c0e9a603e319618019eb44d09de37b3896fc246acb9fce64a
z7e59a465861baee16d249e36d6263396c7d46997afe15096ae9208193a169d545064f1536b7d66
zb475d2d1f419b16dc4a937fa9c5749a33592422fe42cc546300f4aab1511745728f8eb663f6c07
zd4caf74771c8d97d056fa598b61a7a7f8bbf2ca834c9b2d513245269393973135eff463b5e872e
z2f040784595114a7f179a0a8f94ab3a06d6ea77946a83105754195d96610fa50f7a314b5e2b8b4
z27296320b36f5d858b7d12b546876eac3444884ed21afd47a1bdef06cffe60ec96fcf741fe3103
z02683e8e51b7e8784e59349e59956d79d24de4d423a04271f69eda6997847b1253527a86752c0c
z73e1b4264a152a3f96efb4816d8a4ae81726eae4876b9e228e4b7f61221bfeb2fbc532f7439748
z08689c1b5a6590e1945d2bb69cb10a588f79596377ffd169d85022f44a8ed55efbe2d86853758a
zd9372ede0a8b84c9204c7db3a2779795e1458cb17953e790641d492bd20ce4cafa8e40440ca16f
zd2717a7d6cd219d854228409f49477e7a83a9b8e7d69adf5fc8f849d6c02f9cbb6aaf0f4eb4363
za86caf6baa846cc480a4a48f14b4ffb595a185bac8e8f90d7c02c180d4f8d7f060f1e7e05458be
ze222bd3f5c8be1d6d49c951d29a62a0c8cbc51a70d1201c90165400ee7808707c8f212299f7592
z3da64e6436174bd71d897d0e775f0e12a16b8e5f90d084875c59bf8c83eca55e7d4009fc3d35f7
zd9470dd6ab6eec49f7cb5a063b2a82fa49b088b3997d470b393c35a1d6c024475beda11f69dbfa
z5a6ac3350e56c5a22d2124027be5591f8bdb6540a68ed1db89d802cb9064616924228f77e51bb3
z4c4b159bf44659b4e39c248f7d8bf8b7a8d4fd2d365824a51f98d2116f204cd529f951691adb31
z205ff9a47abbb3074d66c45640daa842b516615acb95d0d917111bb9fa13e11cc2240bbe6f0251
zdfb35032d5dac2bd42ef3b7f3d564b615341246943b7a837566e5055e2975ae75d1b0b418b9349
z1e80a4c5d27dfde494c648ac3f60a61a62daa166aedae98737533f26758bae464ab7411bf12c92
zb0a14afa5cef31307fba4b255844190c8e5d2ac3378776455874d54ec9fd28010026bff11caa2d
z813f6fe055d7232ded3cf66bd483c3fcdb3c743ffc739a919bc124bb7239e7e4432159d825c98b
z0e3ffa02ccc95485e74373892a5b37395ae571cfc18a40a109ea229314be4b90205908917730b4
zc91740033412f225ac93cc543be90caeea212007d7d8cbe9dd705ee94dc051c2eb8cc2632548c3
ze49f08f6764f95b69466c1750f8c3b0e84fdc6747f965e5021a02ab71c2b33da2ec0a0facddee3
zdb61507e783372a7c95cfbf7dd6fa529937098e773d9fca1c2766da1c80cdf58340f821e2578c7
z2833da3a4388752f5df2222e79260fb7a30ad32f070e0fed51875a3c7992f2e2b66ece6c321a2c
z605b108e44c5f9712e24ce3ca95c95946d45556d4675688c708da2935119ef62f59af344e9bacb
z755ffed0f4575be6244cf0e023fa4ec3a39d11f11538f56207574881f2bb128acd4d1660ebeba8
z63a2a15882c7c57c472198d56f3e0018748ec3857c160e2ed69d456bad4e64988f68d561e9ff83
ze5eea573e6eec4f26eaa9df47cd182960f40c0f62a4ab30b0a0127565d0a60fd634846de61e2ef
z07c2f3743c41bd9f8fcb102afff1e12b47d8658f27e54a3a6cbdb1185d651d10204f4eefc74d37
zb62a3a1a34cb6637812753734075617e7cbd15845eada57c4e3bade4b97f2a1b10beff766563c2
zcf384850b2a14e140c466d1bceb109b94e3053d6483dd5af52a617f8f008ef6843c0c953cf08d7
zdb522d15a1cb43b2e57b83693905b0a5521f80f671e5b862e34086e2e639ce3ca02ff001288456
z398bac77a0513051968c7e7c8009e7a5b8d4ea4c36fda1b494dc912e58018245bd3488a166f8e9
zfae9304120edf71b7e846b50eae2a0566e0826c2e51abd216c1273488480cee3111077afb94bcf
zc72a18992744553879399aa3e4ee53b523916128da366578a419e5b0e800f53919d5446336cf45
zc98dae9560afdc12008a247b29153e9cf3db74f415ca5807dc067a3374f860587604f71b0ddca0
z010cab2bb76da2ae30a9a22f85fa7495bbe25df82176fd348cc5356483a4c2166c1ce3e9da4c19
z57b04b4ebc9d1dcd5051aebf2d49a5f3d160679d7149a309b4acdf701ad96171a27753f06bf612
z2f50d2f39bcc6f3a74634714e5a63f77738e8f55bcc3fb9fafb7e9521436cd562156c0109c162f
za4abfb99a4b409e7a4df36d3a0a1ee6ecfb2642c5a663a01321f2121a83e02fcfd4f47dff1d3f6
z0715bfa84a3bdd778029dcbabc5683cb7f474f45eb8789dfcd9be4f63193c9ac93ca998c95dc70
z5608d6f88a743a6d66c996c0388a3b0e0ecc5aa7354b82086dbfa8b3259bcce0cededd6fb2e1dc
zf44bbd607dbf5e6326ef55d8e5d306d721c5304f122bb0da21f577d9c4bfd3a512981f5b8f0036
zbfb6cc862ca7d1170a324d06b4581c92912878333db7d7e34e63cbb86b6faf575d7ffbaf22ef35
z3d9d42cd52eb637df67807357b6b4595f271b78c0b9aa84a9f7dd63cc0129b88812db910d003b5
zc010095028184cdc7eca708de15782c701887d399aad4c9e362cb2baeb2e7209411e74ceca939b
z54f6e61a6b17d3548dfa7c6b03b281cfedfc4a94f90256ab81bf893b18c93baf178b9fe695551a
zd17a89b0910f2c9c43aea268d42e47a9fe0349f22d30ff5196c754ba06a75a790ddca59926ffce
z7823ae4a514b8919c8ed28e4cc7d3670f6e145654a4e43a1a42d129c15ab86cf61a3103f921946
zd7777dbda4eec82bc0e6e88953ee5f0650b879af152e33c265d6989621fdfb13f5e1d50f99c53b
zaaebaa4260508f49383ad46dc7c6681b0b9340a9816f11a5054f084115d0d2637e79ffee41e612
z2467434a2c258f9ff8cdaa86d66df5f90f33258dc1a2dca6127c6df26424347f3800acdf3f581c
zf260141c5e12265bae6116678f4709da0127ebd187a02de8233f35a598f5aa0ab8f0a897f5af2e
z1222bfc6bd231023ed5d7f05b7ac9ea65e69f984ec821c4aa0124c7790b93f46f4c7c47d3e2d55
z82ee26794dc5faf0dab28c6efc6b6a96b0151b41ef155d7d4ce04ee661b385a1f55443f70268d9
zbbbb2780bcf13a14db0821585d4d7b2dcd3a199053555c19784a8d6c433ae72df1c1c639526889
z2fd0371bc0b7335e97195c4693fb9aec37e8cb2886815a2127c331863cbff509bdee7cf63f72b4
zcb6beea252b4ad96690d71d3634ec0dae62e279ed8a4cbf0633eaea7e974628179c9cd3d555bc6
z75cb6d0d037c61ec9f6f1fc78a460f9eb7253b926b04521dc8b506e1232540ab0a781431018b26
z438e1e34c76087858b307034ebaffaf3cd46b53ed8f83515ef0251e4ac1f2c4384376876b80159
za98290ca2343e8a7cfbab72ee284fc253d20243faec5e7624b8dde0330e6287928e9a12359e957
zcb98044e305ab654efc8f3f80b0f49fe7b1dc1bf2b1d8d8154ae1d7f7daa6997531e6328d4f345
z4ef127f55d914ad8d4cbb523adcc2a0723ebbc0f4a3af0cd2e08f59777c006beae400ffc5e5c56
z3df62c6d49fdf3634e6d3a417d62eecadec59065dacb76b3b0f6eb856cd65b08c5ca6bea8c289c
z9df4de819d42389f2570ef90fbbe3dc7b1df42acbe70a64dbf9f10874987fc5d2e0371a87122d1
z11875bf4139fe08ad6484bc44076328f93e68c2ac0da6d0c154cbdec4b5b735b9c03d76c7cf1af
z555636f983bbf9c46aa01637e45c40ccbad83516045e3668806b9f4dd6dc26ae3579b27a5e4065
z5660095f970a030d75ec34e728c78afeea321bb62cb0c6e4641001b5a12f7852ec700e2a932367
za78df7cffeb4aee1316be8d0a3d60831d23867f6eadec174532c7e2abfca2db657ba1b1869a954
z7552f84dd3744f0a4d073d5c8b58c26bf68a2e29e99b58bc9c73128cd1f409f45fb6b9b3e90d1d
z276688cefae6edf949a79eca7584c3e261ca730b0c8888c70c86e9a4aafc06fda3efddeb2aa75c
z07ec46773c4abdcc22aac904204c79275d8278c33a944f744e7ad4f28f8ee5b5cd58487382a7cb
z0ae042a6519818eb751466a53bcd535dbaf19f28ce26f983ba91cffc92207ae041a3eea7eacb12
z3853cab5883c1bc260302b942c0d18fccb9c4523b686655ab9260f6b8948849d9d34b9de7793ef
zf8f607ab396e95c89790daa1bc51642c035b2863963ece410980f8a6282410d1190018f3e46fde
za0d28f64c3301176c9273855819c6c6bf6674b955806166f0854f64b07d63dfe16b99e75629652
z965031a4b36b6b63927881ffb9ba6f4bc1cf6bccff36f449cc6b2515e17e06835f756b3ed26f04
z1e8af41904422636b16813de285c0558aac09057ecec9499372d7c8bcdabca4c62639024ec644b
z0b4beb5c8dea6deab1287b6da6e2d261a2d8784a62f86a30ae6207e8b5bdce378566ea86fddc00
z667489ccaaff808005c726e15b65dafc285c52ffa9ed47bf5765aa0c687bab11b260f696718b68
zc0a34090258f92e218506acea15983550d6536626e5aeaf9b5bd36d3b21f2db39ca9c401aae7d2
zaac329a79e71717250116847324674ca0f497b994f93ebbb36299f60368456ee7f844efed49c78
za4d5fc1d8893958bffde3f6dc3f3ab2dce0b0deb42d6ed927a4d8c89b281461a380580b901570d
z0f383a944bfcc190f482ed59a09d47072603f98c43b56aafd43376af19d1d4fc1f0dfa82dbd542
zb3a5e14ef3dd2b692870a2cefe163a94a13a61a0f71a666f776adb1d94c65d8ec11fbf315b4031
z53b23a9fce9aab889f5f1d03369fd9595043d4ac1f0b27141424200ffd6e1e77d109012624aeb0
z069e46f2907517ea930bffe7d1a703c49f3202f4ed37d16c63978287eae90f2a7a323adfaae6d7
z9913397595696efc211161d6c013aa1c6c4ef9fde58d32134951a93ae1bd43b0e823297cdf1be2
z06db34f2b107f43978c3cb36ced05fa26101e0e3b90f8f605345d817cdddc2da4b6d723e5bffe4
zb62af88b28ff027de58799e74cd4a64b01ead361a3d09bf4b8e767e768a1c420fea258a6fc7357
z7b842de8424c4d3755dcee6b12ee308b937ded68e1ed5e36764c4cc46c60b32f03fa08836160c6
ze5e412a945e2a7e2652ed75fc154742913c31ff46181320ae0539f739754cbed0d2c091826bfe7
zf68844e0d5be2faf09e1e5cd19d2310fc15ba63d2040b09fa8f4a082c3a2d30659acec5395ec5f
z3fc156e4fdd032f9fd1c8a34b8cea751a7e2331d25739be4a4719bc35e939ed0f4dde3b5b41020
z2e54cf7313c8d8f2213e8d0df70af6effe8dfb723dbc0e3a6f2bdde7834ee45106454c30d4dc8c
zabcf2b5027aa83c764e8d559abb8b6786c4b743e90273c26665c6de4eaeb0f764a8cb8c72c933e
z10e1446c1ef6d57ee2f73c217b043b5ff242d6e32eac2b60851755400663c6e507e9fff131d62a
z04c150b35d22121df5371f4f068b68eb93563b1aa91523c8dde722bd4f074db280f7aebc7f7dc2
z2a0279730b264df44c14b87fc78baa6bda906edbd2073234cc4c5b63a22ee4f668c8001ade202b
z38f03dbee71d622a99f4a7506465572eacd897ac7d2ba0da376f9ea67bb9fd0d8c6e9663f34465
z3fab94a3314fae9275897eeae3aa7467394ddb762ff030cf8edd5025e7815a9a10f2cd5d723f52
z29eaac81b2a0e3a0704cade73c6f2a78ac6c18a42de3e97b57479dd854c7b8edee1ff2b37c0afa
z6128d5e5e907e51fcc78dbcee72ba7510e9c9efa2fd47d67af848bc803671834822696ea1e14e0
z1a61ec23674ba6cc6643629b6b64e70cbef4ca73798c2c4058edf5415fa728d96ebe2c31ac00e0
z2443b540c5cfdeb52b978ee8a1e8d05a38e3db79661713275e1718498ca79087ab638d4e7be0b7
z5fb1d6608cf55f8ebb722dd5d7d4cf3ae629934be8f335ad5a16c6a7168759ec6420ef6aa3264e
zc865eebfadb7f3d347e73c930d7b74fce7f7b5a4da2b29f1389d995e56c8f1406e138ecdcc836e
z20fce16475df856a94c8306da16fd51d71118a650f2222b9154161abc8945f45416608b91c83e5
zf7bf0387701922fc5cb4c34bf4672a64fd3fbabc9b8764fe90b6b27e251425ee7510b807cb5181
z76f4b8ffb8d11f92c275b57edd42d7cbdfe96b7f660fec62e3eda81ea49f2d5c94a88fc271601e
za0e18fa6834d6fb2fa80bcfc8a1b9916b00246f6b8d3fd6432f7e920a5904cbac5387083946727
z09131e56891e433f21da6ef9c4d2c0a8e040f2a28c1660e6f41fdbe52e26753133a85f0b824b4c
zb36b4d024ca3a4cfdfe84ca27ed9a68e9e0ca837b4bbcf2e00469ec50d7e50a71c7bf325b84153
z65abd93d61f5e901c4d96b1ef1887fb950fea5be9288afe168641976685a21efe238d8720924be
z2b7e0cc380d6cce3304d44489c35c12f0f26483fd5476abb1b8fb8e0541fdad71e7ce94b32ed9d
z114f1421f6d70f6f1a9224a14ae749bf4565c2c9a3705f918309498f69bf5f5aa5e5538772d399
zb1f2e538f5fd522e349644d2d02d641ec511f3e1930e4cf080d56800e038511e1d6360a0379afd
zdb83fc2973b83aba0b29fd2ec163c6d4c382130f1e773476c6f23784b3629a86769e4150db1ef4
zd761c618f1a1792328369e5881f49d88c5b95a204cc7d51b7e97ce65e9a20736088a080e142355
z0a72ea3298b71960ac117b2e0c14ad9a11fee55c1295702e994b34fdc7705be90368c47f0f9caa
z6484b33b129fedd9752866c2c375c138f7ae060a2fb56b36340fcaa17e47e01b95bdf160a7dde3
zc1ee0a3ecdf75de7a306830f23fafcfd1edac57cba3072d3090560efae00526b30f5f2b67ce8d6
ze771cfcd0987423d7d71b6d1c539d6f38022632395dd0fbccdf7360fb8ae1b92a8dc1d432acf4d
z958cd0ae814b0b06c434ce528ed66cfd45c10074d60689bae70d166a0718f8f35cdc9c23259780
za5639d968878a757ca9a8e232c3db9e02e25b5f49a6c4f95bc669a365cc0b00398712edecceae9
zfb93d0430c161d6ee5e60cfc42d855447883fe38551980fb0d96a6f475c641c926b3242553ff31
zd64c7f23e1f9dea85a40865810e3758f4a0c95cad0d4c2871a84755804838e8879c7cc016b4db0
z4e96205d594f4a2d9a98eb089b24d628790efac3d0855a96ed5eee42d4f210d845829da3f77f44
z4e0c4433d5efd879dee5a401a54de7e226edd20e2d73b7b2bbcd16c91a02097f60c0075bcbc81d
z838a2ab26ed9b3ed2af9bf7ea9d05a886ddb4ce5bd35c762cdae13b36469d06abf81de770f5501
z5e1a207021bd26f0222db8f1f91069031e94fa3ae3b777204befe8d3e737590140c82255a7c02e
z52e1a90b6e3afc3a297408eb313f853dabd2dc27965bae8db3584b0e7bcc908ce3c453d615cd63
z80470fe629e0efff8fa5fd394f989ee1217042123f6e8c382bf4eee46e7965e574eecc44afb1e5
zee359d601dd934f51fc86a758a3b41f01902b358cf0a4703e52b9f44041281303b8128e5c99867
zf06f669f3da8ec5fc9d7babb0bcece20afb07ae3861b11eeeb53655f235a2887c52d23d4039286
z0b9d88ce9eedbd68d817136027149abf7d9309943e1db87d7c322be881beeace234e11514ffc34
zc1f204442a357e5069342a2de466b697661ddab72a9a2f7662624da0440f96ab0457c2c4146091
ze8c3edcc23db1e4da08ae49bf21f2604ba772a075c6618042eba3a595b3f58628e6f13ba8818bd
zac575d06969684fb0e088a4ee05b49ed0573f9d3632f44b8cdf9aac857fa607b97f51e748398b8
zc197f11d801f7530497a1ccd453444456b9856fa623718f9b042182f99e9175e3e3758fe889fbe
z07ced2093ad9f18ba246cf2309dcfdd908f4c472ccb8467853d0636607b2ed8a5df1f858b26f7c
z73aaf2e0f382fbb73617ac5e574e84ff5714b5e2f01c3a55569e1622c46d70e89c9d1d36dcfab4
za1ae9fc813749f703f8ea2498017b81685706c49e65e39c75e04afb35c58d23107bf4a995ba628
z32436d872adce0cf67ac92bd5a52d341627285123396b2f608c55aeb02e67e9b7ccf787dca5cb4
zb8958d64da42d8c8b5c8ed03c774f257660fd116c77cf78544c529cc94e442342d2e5f61c9d02b
z2678848c651d1ac9a2f72178459d8977697621ced9e24dc2ae82e60ff45971392d4b1706c1d5ff
z5b5046aaa7105ee2aadbc191a6ea3bb43db5569198b5a5f841aaf7dd14805cfd9b6cb3842a52df
z9b769fc008ecd5ceea830d22e91d654e22cd7d408ebf86a4f416d645861c0f454ff40eb091ad5c
z8cd58468f41420727de4dc1f99af5a1d1973e044af016ed1b0f398b2f4f3ef4aed76adb18d8331
z48e9e62d7cd514521259ec046ed4572d3413edc860043c279de843d1013af6de4fc0fbd5e7842f
zfb0f4cce1176d4b139e125390d529067bf6efd87dd863693fb4cfc5b17eb8d63222e89d5ee33e6
z71a3fac5921b007b26db52fa3bf2f5be35010486fd8b7102a002f56862957a1d2743bf7ba5d2d0
zea64c32c9f3cdbea33e79cc2aabb1465208769e72ef7b936c4e71aa67fa5cee350fcad0c8c90c6
z8f40999427e2c5b5957dc87ffc1beb321d07a2692c3273cb50d1c7c4eae72a53a77ce9efd696b1
z1d214809e2167a8e2e7733f356e6692b37174a3b2d5015c88f098c6219505ff388ae188ad0f641
zbe9be5a22465b102b8ed5d9f1ca6edcf3b1f36116187f07034966a0053e9b72c819d393cbd9ae1
z7ea75769a7a7bbda0f574642181b1231ad9455df3a5f3035a41daf94201559f23073650c2bd141
z67cd40e58d6433e683fddd68da286421b5de450dea2066c659f716efa569df8b9d8ecc6dcd8833
z2c83084d15158337e38e35b1ad404409ea8027f03adbc5b96bd70948af538bfee3dfe924482222
z19d1419298477914a790657e35910c0eff0169560286c4e734d36aabb7baf77b4da675a9345b8d
z21440c33a2908038ecece3774df3eb28fd974391f2e0535bb7912c36e334d31cf0e17cbe9dc660
zd9003a656b0e70a6435b8a843bab006ca3a4bbbcd20ab5e77228c5e4ad0bda22a2e9c9607a5c4d
zf624212af9e8486dcfbc8f03659f76568d980a855848414bf57656e37b33a50bcea772a8b809b0
z641dc85f6fdaa6a89b3666f5205b32d7665fe8d0b214a276f4d6d549e6f6981f779886c7fe3072
z844ba1a33688320321c2ee1082b1337ea7264424de6cbd54d17c08592b697987cce2b123e85656
z02a99486cbcbc70f78e9e2ad314b4df02aca0cd399a419da596bf847d12f9aa75c0cc01e4110c2
z2987a9bc401c084588cdd2cf9414ff644af89ba7c91898e1cb15ed4a2469db05d2d378107f6488
z6965cc25dc957ee824beb6c49e6987c324b165b292af1bec5c0a212b9b3182db50b4aa74fb949a
z344235d51dc30a01fdcc3293b195fdbb9f8e31d9007aea12b14346578e6a98e671ea77daddb1bf
z076ed0bfd2cdf02acc276cb2ac3b88830e20d430884dea20b3a0357c8612528efc266440a9413f
z5d8439710029038f8c113dcac352039c2132786663a42da1ccd38a5713ddd871febfbb3b331446
z5456e43ad52f165043c35a691399132d46cf836e36bd62a1800d1d804b17d902c27cf65653dfee
z9a20fdffdab1299d280a376417b28b5537d7ec24af4129516633867c604a26a2b41355c34db8b7
zb20453400a4598ec33bb18054835af0413174b9a5d21110ef0d7570d0e2f696e6c96be759d5157
z375c6cde5560b3a095fea52d3482e3bbd6b1f473552d5a97e8e810f4a3751f0f6c15e90dd4bc77
z7ab68fb093a96bf0264c93d61f670d3fd4ca6d3b672c1f1ce0b7743fb413e2ed0823e978e5d076
zdc4d9c3edc75c826e62919a4471026ab260ca87f0be6ad109ed79c9c494b577886a6b053e86a37
zd98adf1b1eb3b72b6739c1ef4c78c42e56eb4b0266e5b4251d632b6a8466d340a9e1cbc4bcc2e5
zd9cc17b12fcdec594eb7d5e4b47ac521c79d0f61a3e777a556928cd63a4a4961b0c6593f715532
ze954dafe3820eba7e69c36fb59fd7b5dad5c51e865b5b430c69aa9130f8a34686695118fb41577
za8d86c6f5fe9e351242425012e8844c48533ecf2c74abef8fc612d20f547e21b487778ce904de3
zd4ffbd1ddffb97fee5f30a31af7adaa6f356125dde696c5019e6efbeb8d638712bee18bccf0976
zf66fa3af835a1ff255f2d30b7ac54e27ad553ab673b4fc577b7d9061735879102bbe05487e27c7
zbc03e775cce75ecc687556a49bc629e6e0d00bc21e58180a881b943027d1149a4a6d33658e2585
z360ebafe131fe0fd94c6a2f52cdf8b4f80a00ab3a10e51aded6a1241eec935f3f329246427a8f4
zc2538086a8d63405a80e80ace5a668f6948b716a012f1e30c5789088db39c13abbeef8439692e4
zfcc4939b6ea75b6ab17558c0adc5f5c9e573c561e4cbb0df38936aee38285f9feec055e305a6a3
zab9b28d17d031b35a17ecc029360b0c70bf1ba83aff7503d6dd2cbf15fcd01b5b2c0c74eb4385e
za6c9e1f173508cd51ae4e1df6b4798627ba38d66381c982ad438e9641fa9001a6e48b075345179
zdd01b4c54881459c1032977ff53f27c8dd67c1ce6f3abb5e9ec24e3c8068b107dd155f730f4831
zc58f7a17a101018b5ec75d1b0807943cd1bb34166ee35a75e344ef5c34e39c6709bd5f01b2c23a
zd0c5353f88bf3f635bb51501f2f0be84262d7c4e2e4b94f8dcfeb47d70c7ab11b0cd55692e1b8e
zd0e663d7d66d1af44d102a37f46798f41b19ae507fce2dfc891187cb71e3f233e6d6465785a48b
z2d7b179a98f79d2f313ddad3ef79c38bb1c2d857a8b5160e158ef553b382a9bfb54d3de1a0b5c0
z180643fba47c34e8baefc62b7847e16f10870a4f8483007f34dcd0a536b89cdb0e1c0c50c27ee2
zd2ee865cb4342a8679272fba2dc2ecdbf257bc422fe1f9626243ff0bf3cfccd8703105473f1e40
z73154e2070c59fcf4957d0ee5c89aa01f968ec19c20c2a903f83bb7586ccc2c88332357bdd32f8
zeabafd7e05489c3d0941eef6ed67d6e4b52e015e5e94755a61fad1be3d89cc82a0713b617248ae
zb7c6ccb427d952492c4608c6b26ce86000c819336a61e200a7c98ed127de28d892293000a0aa47
z5b10a2d54230026831d10525e7ea50395fa4309dd984c7766a0c1391feddd3debb513a3e46897a
z0fa437292f682a0d09b7f6affd6dba50cef3cae646290a12c939ed42615cca38e662571ff7743d
z0c521bd044ff528af9570c030d842ae5f9d7c05b0b196032b96c9703d5bde7d2c466d5fafbe4ba
z87228c7f0052ab992ef31bbd049c6e272ec1be18a1c0a103c0fe52d7cf9d2dc0c8bc8583d3ad80
z3bc28906340f8892a6454382ced0f1b4777e3691f0b7f5aa1b3e3c9fe69d65ca57ebb741b8eb48
z1d14cb7f0c2b0c544cf17bb447a7c3c14d41497cf7d5e0d8e30ce5f268d45f2bbc2fdd283bdab5
zc851d544229bf6d588377bd6fcada7a78737147cf1ab39644488f8613d50c7d32ac75b6061db1c
zb7563ea86945e6d3fecbfa0c3c36d7d45d95959bba79cf44c464d32f265bc065ff065f4d3320e9
za2bf054b17e512d6167b2154a9af13e19bd5be76870f0118424c8e111284a46adccbb745872be0
z22b832ed1cef7be822084c613efda2b94da9c482c0b0ee6fb9a913d1cd2fbe26390ecf1e881be8
z076f0d164132c7bee8cd7b7304857528030dba910503d230f4af2fba8166ef894637d99950352e
zd665eabc54430281c596a371d388e553e00980068fd6e6f174eeb4232fa41af0431eac7836a571
z3fb3a7235135e86c8916391100d34cfafa554d0f4654adf2410fa932e1d51bc5f3b2ac9912af3a
z4a833dbb9a91da36592a8c223db138fc85072efc052723cb8aeeb593ffc0f9d42d0e489565d6ca
z4377d525f3eab345a579b6209d35626bf8464da44e51932b1362cf856d48c90964f764c0168629
z4bf2f7d81fa8d85324d0870485218a0890f6b132242f8a4e058b8d85bb88293c17a520bde2ac4b
z591ea7c9721b8dfac69ae05fbc13e3e9bbbb9a831f5c1796e5f82479ff0479690c2adaf6c1e558
zfc1ba11179a8435208b1ffc606f7eb3a17237f0f9ca6cfea119d04f714da27210583f0776959fc
z4d6d1b0edf3f34078a5d9367b91cda70798ef6853e6c3305379064b965fccaea54de1534800e72
zb9513acbf231400d446e0ee77121f2bf982630524090ce95c1f4cd15e56857b35d8cef7c88ecb6
z78104d10335c31360a248c82ca4b3207783ecc0ba906e219a10d5c4363c8551c6b07b856f51dfb
zde3d38b20d88297b0a6eb9856f599d5cdce4d0ae72f219b2d44494b0f197c90fb4d0c004d3e980
zf3c6da4cf8b06a630fb11fb23abba72c4c8ee18136a1e58371dcb57f734036821a82db75c296ca
z4b479516e0e2547cca79ff2e64ecbaf5ccc3e55ab3c803359b8e0c54035634cf8d86d6832151c5
z0d8e147cc91347bf73318c0dd42ccb7dda877828fb024e02956dffa15e12f4558705d95d2dd220
z7998c231227d84c827b29b86789e612b360599abe6b0e8d36a4b78dbb14f9259f372021c619567
z92fe90f0d858a19b39673e581dec74e2237336d4207ec0ba0c971b04d0ab706a5da53693d2bb93
z08882d48f65801d699c51c0f13d3d23450e70be48acde2a50268c037d836c63434ec028b8909c7
z866b73edc736f6e99b953d04f11592c1fbe6d1dfd657069cd23d541619468c05668a2e015ef255
z4c196979304e57792742fd60b2b9e7576b258c64c8754534d2377110d51cce153d0f98f719e08e
z1db1501bc6648a602a98bb8356d2034a9a2565f5b294d91505c5ccd061bea451b6b5589e1646d3
zad9c4ba0155bdd11847376854c9dfcff1ce1290480cddd3f869108792f4fa4c02a09a06d8ca9b9
z35acb93ddd2121261b16a1003b065d569eddca0f85d92146efcd319b2d225ae9fa0b105cdce602
zdcd0e45f7b0df46fcff51f6d940a09b09b90caea160f418fc520fe5fd8025017fc1e99f5af9a8f
zaf854bb6bff4061f847fd15e004999bd72e680737304ee36ff56c40706f9fa3d553e41cc7b7cc1
z4da5c1d79626bc7bc2ca4aebbe0ed4fba409f9a3e64a167324f90b27d02c01ce9ad6d12bcbf0d4
zc2e0a043d332ca194850194fa2a61486223b730254d7fec2ad1960e14a26612965abc0c9eb6759
z050a3b83c7710f87bc9d4249989b89e3d355dd0bd269beeddeb3c469b43573c9a40844ced0a786
z21ffea6a6e69bd1366d7f6a40cf111aa5ca98008b50a107e9fce781732fb061b3d4bcb1c53f17a
z71a0fee0477c5679cd94edafd5fb65a29cf029b7a5eaa8bc0483c7ad660640c178364ca9023716
z462a378d5d804e20f06789a6e517ea0bd0b56909494194dae95141204108eb65ed2e06bc673d86
z7c17aee59c829eae72797b74933c60a3fba6c6d5e87e70c00110ed2dc9c8cce53446cf1a00a2ee
z8cf9e8e8ec843d379750c3a718269976ba0a6a4abc6e6f8e2a4000595e6fae5c5ff57ad1c1a0d8
zfddbd3677418c54e94ca0f6844f9341c7aa5b82376f524779197a973a0b12b2c5618940cedb603
z4cb5ea9ef759e982ad52cdde9ad58d96a3fdd31eeb1d41f9b15d8a11d87be6862966f1fe9783fa
za9c15472222f99e7c33ff5fe28bb750817872c07b97995f9927c5b7588ff0e40a4104a13614213
zc23365c11e5bef47275b631645c509dada6bb46343fe319828f3f99562146cd657a616390e92ff
z52a5e0655b37bfcf1261757fdabaf45147ca7c127a94295ed84ca7f908de5d05d56301ebbea64a
zf756914c070705a533f974b92c2adf82a5838957f1c2141ef045391560f89a6e56a9911de5497c
zb61acd90d610df78d63b0c1867a584afbd4a0921f439d24a963fedb055720defb2050b39aed16f
z60b9dcec1270a7aba3a3b2304098df1fc960a9b4fb025f2c42c2c9b4d93715bac0c385576561b3
z4c701605a33b117a0809ac52b6824b5601b6b2136d085b080760078db161d522cb803934c73e10
zd319a0a42e415ecd290d65b19bc03719c8b23724958986708129f6e6b363fd8d0f5d8dbe044aa1
zf0ca214016aee149e741bdda554ed26561caabd20f5168d71f472581e00dcbf4bc733f483c25e1
z8ba7e534cf9568b9fbb0582905afebcaeac6e3cdabb94e30853e8b3c52e8311741b4db428d76cd
zf6270e40b0779d708b2e9ed6b23919c6a3fe5e38a6891fd49a7415db85260a287e64f29bcb5c39
z82a0278a38a6534b197fbb7d6943c5e43475957a99de407ec55b39b589e1e6231b76227bf3f1eb
zc24f7a7f25641d3432e2d1b9c19496303894888e55db6627973d17d872ce4c1150f9c7d9a13047
zb183949d0fb43bfced48fb41529faa60d01585370be353704beec4497691af7704eee3b4a07604
z2a4a43da2de9e0e939db31dac9674b75d40146ddfd20d61f4dbbd82f33a4900a95b36801f7248d
zdbffc5346cc515b09532607a4472aed0a917906a3546099e94d17330cafe4de9509485eaaa00ac
ze4d7e15a5cbdb6da51a858aeebcd8ed4abe048f3481878115f30f17c947e8521edd2fafc3c2024
zf7e9a27f88a03dc8fe18063eb181e710daf85cc96ee1ce20616b80a6b95958e788f0ea39573870
z05d1f18be45ccd501e9e21cd3a8bc5a33ddcd9ffcab1f89603c25b8670ef485bcf42e4a88520bb
z9e2fb523c1b9fe273edddb41816719fe5a41c2c71efaa60684a5732caf1aaafec93347d2a49ad5
z51fa76c4f19af4ba66a63d4c2dc2b351fb7af510866a5fb860f8e49fd7a8fbc983cfaa042853af
z0f878767f15f806c31be43f234fc1b557097ef9b4e1444b992ae5a1c00bb0ff5f9a75a9c501559
zd1d53eb1491b8f65cb08dbe64f4983d8dd4609dde3926a1dd759c9e208a940d83a5f441b0f028b
z785d29f5a202b6bcf8040216102c1d44513da375a285df38ed4cf0873e2ed73fbcfc3f221aa29d
z0a96c6a627faaeb92b5a3af8cef9daa172157578c409d3512b455a5796e8fba8e002e167fdff67
za7a77998fdd0a23fcb6dc216ef7d8b8547d2e8e9504bde3cfe4815b1df869e01bf51f8f7f1ed66
ze386955e6cd99f8c0a0575f09d2938ab82a42e6a80f71d3e8c10bdb598d3c658bc94fad9c637af
z5fc093c6c3ede7bc7a564720c868ecc6546626ece6be3590b3970b8e66978b2f8086d0816cebd0
zd9a858d4e7979b868a717a114d44040473a2b729e697cafa392446318c29d3743e874cae363f58
z4edfb84595dd905a76d7fb8fc8f14c210a3cf1ffdb6a5acb11da986cdd20e9fe124a860dabed85
z609240e22e9b21f4ed1eaf18dcfbb0ed09d5e5802d53ccbb06a7afa80295d6100e4cd082b7799d
z01deb6f2630733f08b8231654f7d68f7b355c715acff0a7eac5e3138082041b1fb6635eebb5d0d
z610bf568b06144471bb6a4887a14ec448bd8e8f70b54569ba30276305e14e8ea565fb0da1360c0
ze94546062e5b34b1cc13f7523d63d6d9d45cf2f54683eeb74074e38b60dee58ad29e532932bb05
zb1f223d9d7776d8729fb7385b23944ca0fbabdd3879527cf50bc2daebee3f707591d223c94bea7
zb2f7d475f27f1fe1df33783ab847dbbca1d59c20048f4acef17847a86a36bc3f7a8516598d7aaf
zefc4cf81ebefb0a3cbfa45cc11e0ef5bf1250a1fccffdd402a317cd3e804bf7bd7d71dee196433
z56e2819ede4462b6386c480740982af76f18761e21182eca912efd3bdaeba7b279b5efe2ea1609
zeaff886c69f62638dff3dfb009e9622a9d1c336f29d74f701607aeed77777adafd07b9cc52dfbb
z84d98714dc942d696aa17327758b31f0067a3b95d05a288b62c721ee26fd5aa2dbbf7eeb4137a3
z439a59e1bb287fe14574778ba3e7b992ba6d05c6536938a805e41d04a918011be5ac27435cf808
zc0a9683b4ea1cb05b1c7572247d19cc746f4dd4869aeaefa1181515e9ccf0d1c0b8903926ec2a2
zbd58921749f8a1b2ba55e77ed2b5690dd02abb47a113b43602241cbc80cf5e8aa1072291384bf1
zd5d2bb18a09d818c3a2ca5053d22dc703bac5604cb4bb1c34986b540da157512ce9d03d6703320
z0c7eecf49b2754710a107c8e6529a76761393ea71d642c65daa65971f1e4d87365f10328dfb332
zb79c6519465cf8b04e0f97ffd34cfe9d6795f8a630cef87f26898aa4a5414442cb3857342d9b03
z1fc5c5abdc99e87ba6e89e609dba04b1f735f037d21781c023e3a703c1ebdaafb5262bbf391e29
z2277f0fad42066a2dddf7ef07cf1e11f9ab879041741098f401066264ca1c952792cc7a12dddf0
z685f6a66bf2ea5820171b05ecdd543d0e71d6d95e1d8d33daa2dbad1c9b0262f94d3bff914ef09
za538e53e72821ae0a33d26b193d1bc522a3dc479cefabdc5493b5f6f6364fda469ce844edef5b7
zb216b1d008a6e2c53608b58e11e26e57d911539b986849053ae6df2fb537ea2dfd8d8fa3ca0ad6
z47ba33c99e72c4e2c9de563e4a0a045e571ee8a00d2ffc25e3e4e8c81cbbda803ee6b94caff6a2
ze9f1231e36808a13e31e414cf63ed2ed57d8221911230238f489132627897c74731464f1456f32
z97c5c3575fb6b3baaaefb420e4f339c5a6b33304bd37de8b9abccff80900160061b6cff1e79409
z0aabe7733cf3044c13be41f2baf5c520df413e088a8ca7b9478e721a1a99599e7b66f316f8f09e
z3572b4bc90f94dc2a2adb516edc42812f4fccddde161de16a91e6686e2a3a9aa4bbcbd35d67703
z3c257a65fc0ed02968dee1d5237057d9bca6e9b33a9474560c672006e02b2f6e00938670146753
z055151742266278859c9ad1d4286abefe3ab77fc3b74ee1aa66e6faea611eaf4d06e9d6efb3d47
z4ec274648e2f37ed760b40d294e4948d0cae9cd556d51ee7f31c176ec28b11fe948b46c0b07522
z8579d4545ebf6fe69848489c451e91ae96ecee09596ae4e8fa54c38fda591f29131011290ce089
z4167a487c8081e134aed92cdde32caac7dbc17e1c5a1cd59cd2ffcf2427b6ddb7ea3dc8e53078c
ze00f00c4cc20ea73e42413ebc2f3b42c8f6f73b447b4c4a7d24fc58b960d79f37709cec9890458
z7251c7e4a01282510bf19a1ad002165708b0ab8f6fb3ec28dc1e0609eb1e4584fd5c95fe1acd90
z9e9af231100437d167dad4604e5fb157d296c09417751a2c71fd40d1f140af9583643d9e6b97c7
zeae79838ff58692d73f526a4307a1333722d00e10ed9e7dd5899867100b5830edbe47c9864fbeb
zbe846da1cce8434f9c7d3f7a4bc9fb3242229ae83a73ffff7f81e8a6c3d3a8e8ea8d13f9913f9c
z70a94bf52414db8719c15ffd9d10d727e6bcf1068192d93a09d63596cff7984c8638881ae29e15
z0baf2580a174a4ea6488e3b86420c03559d759dd362422e1bf04cc5796f31d0f4489d0140cef21
z4e79ec143ef98bc9c04ed95a86f5999f66ca705ff8973bc5ee0601b7dbf480ad3b555681b5e2a4
za132bd52ca84463988741a4d5c6630c1546f8ecb9efa864aed8b4de727d6ffac11821c2e9ebe7a
zddf36dd5e4bec5340f09cad84b75a582012062dee8b7ed1fbf8ca1a4a2e60f6ac2506688ba3ddd
z611c2c5d43f4b553a583dafde68ee0d8d3b53b37efb0f622f71d914c1ef4c18b5e9ec5ba433682
za5f34573e0023d91279bebb3f2b3ce230ca87ad6516d8511cd165efb5d46e541e90a671664927a
z57cf6f818937bfb6c27295b41e408ab0bbb080d369e74a34b465f03f9c8cf4bfe041c950b9e3be
za2eeb4be03ffecf799cb170d1f6f1d134fb4a54fcbcdc0a0a85925dcf9101601bc88baf2d8d980
zd5b5459c1fc4fba40089d1c0d7b09afdbcd9f3701f46a5b2ac91302f02f5ea6f91559c10b2dafb
zb628174db0c6303385e89f4582500a925a82b63bab6bc98a1c84812eed47f6ace79a0404d163a9
zde21e8244e4fe4d0236abbc788857e9f00d3d1ea35533e86ed526a4d77d756c4d00b45bee8eccb
z56c982164470b5a928cc2e998c286db44fbeaceeaffa16225d283c687106dfdafe273f5f5a48ac
z3ffce453a519055a30a333afc22fbeebcfb0e8225e03ce1cb9878a0a7320778d9205287f03297d
z547432a7946428c40dd56c43326b8a2d1549222f4ebe81aaeba4cc18d14f2b2c80e7581ab9ce7f
z6737b1a32d20e36b4032005b409d4c783944edfba06d27ac9fc97aa7aef34a46682163a9c5b784
z05d4fe9c9bd3adee609cf73d4e61ccb811856c3f5212c4d3dbcc4c0b6f8e03df2c32c3a82a3131
zeb53e42a7f01334fd4b4ba38b59d165417771472d332987d0612352f6a549890bedb1c06013314
z60c35a8ceeaee96978d0fc699b6fc568b07665e90ceceb6687b878f42d4b5b738fe755cf8ed060
za8c1cf8fa40cffab688ea692ff7cfe5a3500316da0a434b62a4fcc4b72875af3b919fcae963251
za1da208696d7f81b76ac9acf086766e766533d0317543af05e41c5e62f67d9d6828984c5de2da6
zdea3bba822348b07782e80395fc1ca91b98c89d1ed0ab3d41ae49e9eca5571f5ca265d13827933
za1396dd14ed1759d94d2d84c0e00e0031555f745dba3a6d10f36a58f2083f738b28b3143183dc3
z352c24255403ee230727f0a7a8b5dd35a19606336e86d6b72024ff7d1e576ab16325146c290cf9
ze5e59c01c71323939c035263e37e78dba32e329c5b18b71e9adf0b0c1e9ad529cf9a7f33106889
zaed4a89db24315e009f241c7816924d82b3b5676736dfcfc1ed69bc2f41376ad130a8be580fc25
zfbf0d5c7c6d230b50ac0bd417844baed7f58bec48532890f552abe879e00cba1b607285c92c231
z7ffd8f70ff1fcf00884ddfb4da821e4ffb084497b208fe5477d26b3a15b42e1d02e7262460a658
z6a31a63a7573943ea0976dee1f4f1b11ecd37cf73956ae8ff98aa7f1927e0a94f0f092a51e53fa
zf62c6d672600d5965ee1c5fbdadeb2aaa70707fca63f8872cad635d935f0fd73a47c25fa079182
zb15763973cfc1566332ec0d6ae20265679196471c03ac1f29a0b2e48b912ccf9e4419d70a30485
z185b2a39dd52a581037b2f615235be7ad573a5cd3be8e9d870ab26b7d9348782ebdea18dfe3e64
z06eef10911277968ea75ee56bc9ab251c1c0c43e01bd8cb9357d00a2d955df6f6f99123c95eea0
za4295a6a05656451881ef7849872a55f406ee8234e6cf5ad4413c0423a01ff04fbe5781695e3dd
ze237fea030c34fc3ace797876c4e7fe011c65d61fdac7c04ac4718c3ee88792c68a3348165bb83
z47e40e8b87207ee1645b9ef79d9b9cd77cf5315467a584ef7c3df426248d66704ee14fa74af779
z5c1e81602bc734425b5d63c19013289faabcb0bd15d3f3d3c8526e3bd10b41d2a9d1d8790444e6
zb5f84bc25c9729583cd2be2a5351e739b1b37e0551a9e8855f5efdb1ed9d5b12dd2c78bd7b6a0a
z671f6d900c08763dd99ccdec00a42749cfab37f34c6405b6b79ae4296ec2ef3f40083719819ad8
z5f110d6468805003b3d6203f3de844d9e6f137bf59ce8a3f3ded942fc1e755403a83c34aeeb0b0
zbb1c9557a22ed6ba7e064aeab042e543495fa6ae8fb63eec2716916debece4e8954511f00ef317
zb3536d8857a0b8a28759f492e6fa88cef9de5a5912ef3fab018925f093f8455a32032bc8409fb6
zf5f6109480243c405460f246854b22ffe5905eb55b91510f8d48dc1292d9dcfde1aae4e656d442
zb207d6d82dfe6a7be19ea8eba40270a92c0a8bdfb2cc477a7895a856b74454e761ddb5a02ec4a3
z4a3f7c645823b425c240f70f0debd0854e877d482ff41b1cbbf52e0111a93c7f3f19a331a4ff97
z332abc667d64f1975d901d9708f8f9d9ee7eac65e90efc406d84fa7092228102adca9578a2616b
z4361e125c152e50aa856a44719f73138004a66f954eb512f9bad406afac3e64fd3a6281109e5fa
z98889c1d300d97087dbce1ee80dad938a8cf582f7ef32d23dadde6909fac694661e0f82ac71a59
zd98e227c7b4d4e47e41964d135f63266696fa914e89ccd827d7304de49729c262397edbc11e847
z5f2bdb9d4654604a73b1d3e7a89dfd2810e42a39261fd2e1929ddfd67a18ed07f1a85c5ec3bb4d
z0f7ba7d0bd90cecd0754fe406e4d2cdb8a0191a9a67790197a668e1409b1e4800ccacc06b4af6f
zff6ff053a3751e4e35ddc847c0085a19e2ab4d2cd43a8381cd5ac2ccdb54977e6bd13474c231e3
zddcb4eb86ff350635c2a99fee671ddcc173625907b5a17ae022e83fa5556d1339ff8ef81d42dda
z0051aeea111a05d45907874db1faee8ad55c4c1a1bc2e32dc96c61c42d17eabf2a9eb08363e6de
z371bf20ed509b77d25ba5049081bbadff5a1b9326c10821f96b0182bfe2361b9849e6d3124913b
zfd6a9e70888fdbda55b4ae961c9b4ba48daadfa23e36841a598e1aaf183add65c339c85ece1911
zcfb5dc0a01602befa3da612e7a95126166771a4a012840cf407efa33031dfc1dd2d94d053ad191
z7fcd19e1b90598e14c4e31d247ffce0eac36be4adc707c2c86f0424af720f0dac7d1b3e027765d
zc3af3d414f5f8a6515fc5a540a7aca6854d98e5fd28ff195239356e4e5c12fc4810ed88b9bf89c
za58c1c923700529473474b437e07edda2e0442c929ea9cea322b49371f0db8cf39fe6c7febf2d4
zcd088429abba49d117b3f1c71f4a3887ac8ee2b5885ecbe9ce0bed3b1381484b10479a89de94a1
za2953e527c27e28c143596733ef818b88435b7d27553947398f0a7f48bb8357619639485e10649
ze6c9018fa8ded2f1078ed7db70d526a3b128f016c6d029378c3a58a6c6f39b26a76393b023a44f
z1826207b99177287bdd579005762ab105ad549f777cc0bf3505b98add05d1a88cf0fa67af18126
z3671aee0db702e6e81be97373bfa476809581c9608f041a3b201664dd7bca99e19d188055693fe
z183523ced1d2c99d6ec295fed25a02a2d57b3602ec1c6ea1af8060c4a872922df19b2e14d2e56d
z45e6f81cdb509867bfa53a3ec13e10ccd1afcb570488d9c81cf202540f3981161217191902aa52
zde6acb9301f4860ec892fa2a290967f89cea563b1170745c90d5a26ae36f1485e9b4b1f062aabe
z7960318b013bbe1cbad25dcd634f2aba2a80df9f21a5ba79cb842e0f82b47f9b85d77fb8f15b50
z283d64e630de3c1bc85fcc59a34cb7bb7348e880b644f695c46ee274382148b1c89d45ef70df93
z92547c5ddfd83441cd8d1108ae3bb5896ce9fa4420520ab8299c26bb3f51d7bd6c3c2537be49df
za2f98b98a859a6dc3ecc6bc38539d803580e9b0fd56eba04fed81d952688c5abc247a999729580
z5b8bafebce5c156f44595ded3761cd2ab75cc2a974ce24a126e10f6e8bbfd30d3587d4be4d555f
zde2c1402a09684e9eccb01439369fd785914b6abab60b56aa9f7756ffe6e626d97774f34c24f70
z94515f39883044457cc680230e8f7795699471db01f3d6c50c5c5e97176e2a19efdf6370c9808c
z5c1ae8e93e312889aa2e91b4810f3a59f4e23073ded58ce52d21b6ccaea235fff1985a2e80b34c
zd217106530bdfb4dc27abfcd2d2b91739ca32a41580546849470da4bf3e3efdfbc29ec600817b7
z9af60a4130fd848c2e62f1cc7f09dd25ff34eb76b0d1f2eec0761aaa9ed6601735a10dd6e8514c
z0b05f360caa997a1dea6fcd55a44cf3ffa5b755a01f8cdf4f4713786538d0e5b089b106d496c72
z60c5bf87a8ed138a5980fff331169bb2fe165f28252c951216118ffdd7b277e4882f2523baea3e
zc7729b4510f568da2e6c25633242c27a0e040fe43ded5fc68dbcff5326ed8ed31fd3ad736bf60e
z0dcb32208fa1f6c83b85528128886387d089d85f10d1dcc7dfa799521a7e39ef8d6128d27086d3
z469eacf5f2cc4d536305349fa579898fd963cc30d89f5d89b0ba397966d5bb9bf4436569d93a12
z72ef07157b05d2a71f7040160cb8d6c555fd1fd8c8c870829e05ebf1a02f4a97e7bbd564952d56
z4c1ebdb9266d6fa9045e9a0c2b6169c97aaf9c53bcd5587e36ddb8625b8a43116c209e8146dff2
z044307816871ea454d243a10a1fc179439a81f49142b294657a49f794d86d815ef6a861ab1eaaa
z185073bf75da8ccfb27fa8131fc215c3e4e92c93a0d010fad8c46aa338de7783fc251686
`end_protected_0in
`else
`ifdef MODEL_TECH
`include "qvl_content_addressable_memory_assertions.mti.svp"
`endif // MODEL_TECH
`endif // encrypted_0in
