`ifdef encrypted_0in
`protected_0in
ze74c34e226135848fe16db9ffd31815111b6d7fb642c521a3f628cf6da949865580b22efd062a7
ze90adae0e65e66a2c36a587d0a790699161455169ed55a01f2084f11770a774ec4c588039b380f
z6de9c5084882a40b79a175f5c2114b2b6d78b070cb806e1c0aa9258297f4687ab308bc470f0040
zb0b1de382961eeeaf2e279e1462520fc31c119af8f2b214846f56c2b3cd2eadbe4099496abff18
z15cec83ec4a77b868344aa20ba7360908f5c0de2a79abf8b3534b883bb12180f68b5d4beb444cf
z3fba8f13afb0abfe8fcc4294810f75afe452434d2d0f1166236c82f76edf1e12979f04bc35693e
z32ae028996dd85737a8f5adc1ebb94f39c940246e887647b64782cd7ab429b0544c173176cede7
z01dfb26b1f73408344a52b7e1f117f12bb9c8077b34876c2e6fdc085981637012dc9754765e1a9
zc512ce062e0b8fb16a214591f5c81e1353b900a611fe1f4886b57940b41b7f2ce99a7b84b04b90
z916f717e73bd10589c81e207ed77ec660a8cbed5b487fa50acde1b055c8870bd8676023f21ddcf
z9c98cc47cfa2d654ff1365d1f45035a045a66c5dfa8279050262529d2cac9e64fd27d9c7de62a7
z731bc808811ded9016570962244887f98fe5440167bd0088f2f049df882af501358497c3b28776
zcdc5426c7f52a851c35106bb93e16fff984784050fc808fad15da330f6f0607eda2d0e0e4b1215
z2ac5b11453f6b6c5c6b428261a64553d70b4ab9f1bf3f153bd631387c118a296ca10cbf0349426
zcf2ea5eb241fa84c8ecbbf7180f10eb9ddd4966d421e6ca571b198ed195474578ea51160ffbd6b
z0f73216703aef2bba31d04f6d0877540c760cd2535de4136d5bd4771107747c34c07fab3aaf6bd
z67c5eab3938266c996e67839bfd448cabe88dac2c17438997a3ee0a0543dc656070eb3dfe7c0a1
z57e24e01799b1ae1652a0133882b63649084f8bfaa3118d2448218b5c4119ef2134dee0d7a292d
z80c07e69250e6cb0856a07c01efe3f869b070b26474ff619f1ee9676ce10b0179ed9855d8e02bd
z3e17bd42a654e974019a7ca7de85bfb3ac5c169726f832c6b918eae789fa38ca70f5115a2ee7c1
zfb52b503ce6ce35b7dc5989bd64a1623ecf327040db427ea1518177d8423992586c82ca8ef5783
z63913b3bff1336b6e3685dbd63eb482c1694cc8e7bb0121103cb3f779f1afdb33a5dc4caad3fca
z3ad61f9e6798c7fdebf82270990759ec1a4107e22a744a216da0132a2888c982add83dedd55b92
z473c98e970f0292cb4fd1c6ac764bf3440c9b1318f8d50bc16bd1ece42ab2031f5f07b6b7ed034
z152d8af907ce476029716b8636a467a9c888befa1aad211cc2ca016bdda818d13849dd75a5839f
z6756c38996bf1fd29a8013133e827e1284c5f908cbce9176d847fa4b906389b78f9e9e0343adee
z6c396694041397a7066b8ff8ba15acab4b0a8fca1cd59d7230893d14f43885c6d05745f6dcd5ff
z7b709857c385e6b3a44822e2299d67e0d1dd9b8a8e59d49f2fbc7471344d2e31253a3643a2d2ac
zc531ac47b48ba29b34a9b97ac839f2961ef05e9e569eb8116f423833b06a40d2ec125da5560702
z935b2e93f2d7b6fd0eba8d520de3e943ccad2bf09454417df7b75fdeb71b21ee1664ea4920dc05
z0e2c65b5d7ea0b06c1f6c7427878dd161f39bfa6d6e9db4341aaabbd1a919d9d59672f6d94767f
z65a75a6407f0fda0821edb1a0d812f55845dbcbea23e60d4360f619c9e920c2c23150c86b35074
z33a32c5b0ae7ec575f32e8bdfad06ac9746d1babda4322d4d98f9dd9b5461da30e9ce1e4e9e640
z301aa2035586dd3eabbbb8232856f3cbddeb4defb7b5242acd951c976b88adf29df990a5e477a4
zb27e44d9ca2b2efb77cabc8de060c57f6dc56eb62619ce08757dadf53b7863a85828b784bf1449
ze7b2394f82dac3520b11bf77fa430735f6836f2095024e4cb1d8be3e9190d3be63e0de72799461
z65791eca001e0351a11f794165295e779f43baebb74436a7bca277bae6c46695fa552409c0ec10
z919251344794ab9ad4838eb0498e675d28080a72ad443eb7aa949d94d3ef5ec26a82d3e0f73c36
z6b3f41c8d20efc11357a2c18d7b9d894ccd6ee4d3e6199538462cc70e292227e860613dcb08fc6
z38aed211500a33b19457a6c77a6d44f24bd16bff567bbb9db594199bb300c5be9762ecdfbc3f46
z0ab8f41c40f3613e09d140372e3f6a46609c743a06b86e702368c16178cf27918d854e60c7399e
zc4abf9a5bdf0c676123e38b04cb635c45d39ab79b6622976528f0f25b265839fa630f593819882
zf4dc295379e3b9904a233a3e6b1fb8620b5530785ef8a345e0e38ea0330a8f93cf9a5a7e7cbc05
z95c606b8772c9776d5ad0d20c8f901e52f8f928a581e0330d4981cd9a5722b69061d1fd0b74f3d
zf6b82e12c19dcd470c00f199a1b98f2c5713517487ccaa05c30b45a0d301db938f1d05fe45f0e3
z0b44e4b9162a12802f87f43db839f0fb03c790ff451718d89e6a84c66467aaaa98f2745901fa29
z96634044218ce0e80e14067baf36f5566a90f600e799fb1d0e09bd025e5c6be5aca351623cb582
z4a6b7e1ec885d37aba0b5ad5aeba9a688e9377a4aa563f4576d2432d66b8759d57e6057a282bb0
z542289ac47e4ed93e7bdf2b01de401e0ab91ee03ed554924b5eb410985dc0a4d0aedadf98a8b1a
zf823b605842bd0a2a1df959d601cf28d5caa1114dea17e4b5769a4628174b299f6471b61f854f1
z2c9e4b48aa3d7280c25372a9793c009a0e9b1fc0b7f1fc90796231ff83a9af176986316b93c624
z91343e9a7b4920f6245e196ee09573a7ea5b5307e76305139692215f839c152342248ce8dcef3b
zad6b98e5423dc6b3f96a59368deb15bb04837de37691214726a9b8678d3f3e1cbccd2d577c2f9b
zd19e35e103ec72071a5e3523c03e365114ab319029f694e0f9ddadcbee8511f6428cabcd922b77
z4c2e2832d943474d83c2b77686308a4f6a035f7d942efaef0953ea421c4e9bd8e90b169164199d
z1322e63a5d72fdb6d01dbdc3f8290730500386f9b4038f394257f65f65202dac42c2a34eb4bfc5
z812f91c9a2a043f1ada34b74bd39f01c53ddf82d16b08bfafa656e9bf2cbf8be25bddd5eb336bc
zb0c04153b98801384f8db31c2e10d80d457362c081b9210b0f5e0c431003f621febb64cb8ff9e6
z6708ee998515abe17a8be11dab279d65c0db545623bc63fe8e424ae581df19ddb433d42005500f
z15f8d07728625d480f9451f2bf58a92fb2f214f4add5bf35e810d903704df3f972bf2b5b18d32d
zff9fb10def312dbfc5bc84cc5d4212e57e98dd9b6e13003d748dfb95fcbf715550af9aacb6c16c
zee1c23b99349b532cd1bf314a5d70fcf338f81a011490b59330b800eb925580e74253fca9fa51e
z812ff1263404ab3cd1420e11a65f1202b85d6f07ef9780c738292f69495a6197f384a9956fe58d
zf431aa1755a4e7d83c28bf35225a4ad64310db90381fd27c3f79a745a423a8d526ebdb6d317019
z1163c3f5e4c582d6a7010aca857ca2eee3eeafeaec766ed20ac0c0b329675500c3779bcf4e6dc2
zf7cf8c2ca643a77c52e53c4c237d2a94e76322564f09a750dadf493ec522a8dc0e4487ee8dc8f2
z4b31ae6bdbaefb1130b55d9dc38ed7afd136f3ef8abe3d80751435b3e9de7f3412f1b0fc6e73d6
z6ea6fbb9c5363b927d2a959e217659ff5b0c624585e315e2fe6811856aaa2ec45d2e4d530f1eaf
z99762e0cdc199b060a56439bb52a0915092e846dd54c8a604fd6ab5d3051c40d0f9bbdf8c520a6
zd862db72f40abd87a6bae6edb09e1aff885eec73ee6a9d857c8f71e68783e64bb4721d2ca2b5e3
z62dd7d4554ed3e159e1add7251b6b1c579b8171f3c42e483cfc250e9a40e7880833a9cbf047b8c
zdf9204c90c97d522a1501b7f43c780d3eb3d27494c68343a3dc24318fe3e1b634c5b7bc4503291
z9827644d17ee1ca28b3371ea6dc287d2ae780655154d1a4b7cb9e8caae031db07a32d8c8ce08ee
z66268b6bd3dfb923c72b80b5b96deafe275417b60bc494a58b8f244c8904da850f4742c7b65f7e
z0e7d740bbd93cb666a677df004b4ca827bccb854d86f2428297e8aa802217cee1e37d272c5bd28
z9b484fee7bc037af953f006dba295fc52070c29da4210c90833426b6cd2730c2ca7efc486bd910
z5ae7e538772892d7696617928916143a69fc08caf58e3e9ea224390c73049f37b94fce4d38b92b
zd11bc15edc2fc57893250269eb75132be4555acc773796b4e56866673595afd73fb635b12451a8
zbcaf9b0dd73b2e74eb3df744eab1180d2d98f0880356cf8d99929e497b363eaa4a50080d227442
zba88647208f77a8717c9c0e4c1eb809a590a902e9437bbe8def62d19cdd4edd803fa70f0230518
z83e5a4671615869f07c3ac98485d7200b7a5953b83623329b25289611301285ae1698491201194
zc26712a991dc654bfe2c044d9a27105a95eb1d5bc28751f097dd2b0a77f069e74c8908f567297f
zf87d4c18f1522fbcf4e7891f0be802800d4b9b95213329e6e523184f3a1c16840f4630c03bdce1
z528042c0d10285756d8dd95edcf2e5f72850d1b505d697580b73b019094950623d9f2055795920
zc3970ab8c68b32a8514c80ed5bc282aef026e0c5c76b9a5541df523dfda8e66a9c6aa0ad934f3b
zf578b573b0a19f297e8f82a31cc5ccd9438105f632307f4be6281d66c86eadf176bd6eff1d98a8
zd2920376f99bc54f174070ae6c5f808d6619d1fe952a21cb08e679a9b98b159b9350c2e0add977
z27c9d4ace12221da68b965b1629257c3c8c942d78341ad530e7b6f4a5479976c9b08bd0461ec19
z27b5f080575bf84776ecfaaefc4a6e3fc2beec1725d33bdc07b026caf1488fd43ff726515ef48f
z87720fd81d104f1b902fa0799f84eccc6d967c7bb22a4f7820b206fc1c0a390a3323fbfece427e
z23202b41dfd514a5299be1dd5656c79fc52c11fea55f5678556322147dba305a9c2c2dd1a48535
zf4c0777cf5465838d842c66847597cdf221fb2ea86fd273e7a58d926063d6cfa7cbb90a7eb9bbe
z4097e15135e15483c5723bb684288290e16cf1e06fae21174180ad42ec7517c10a9a92c5daa480
z00cc54191a4f6a4780e1125c017e21ed077d3e6bfeb969444eb7e67db0f2988e60d3e3aaa64611
zddd917ab3af8647d4a4b534fb458c4ab7b74c65d61c6e1cb4954a5e94581358028f18eceb4a580
z64bbdb76e514e72c00880cbe429aebb360ce118ca83050e1364794fd05741ca0937451b2e3f11a
z302cd6d71077a7b07858f935cd19bb3a5c04b1982f152a69b4390aa66f08b81afa4aee3eeb9562
z60e1d9d89e17ddcb901ce7c668bd846b3270be4999bc445352c563167eba8719ff28341ca8baa0
z686084f0de218731dfa0b95ccf58f76c65588892cfad69e23dc3a59f63bf3de88f6741bc7fd19b
z0b79284e93d2f1f58cd5e04e327a6be755bd5a790c60c79817dbd5a4b2fbec0d89b2f31b2ba66c
z97e837363896047e5d2028d2aae6dfd3277a3c9109e81a72a67d6366d1813b5e5baadfbc721ca8
zd50965e91f8e25e73d9f8a9f1b8d47e29ce2c073105fab7e71599910c35df517f94d93ec39e2be
z1e3e9f9cbe8eaba7bdf3fd0aa0a6de61f15c784f69611f2f075d947bfbf19aeb2147780a61c3d7
zb930ef22bffc2771a2d6b5e415a562b6ceb91a18904e4f7ffe291377eb0dd6d1afd88fb154d079
z92d21ab8e9e57588207d77e388bb80fa660a4294fe13dc4ad367b6ea6464b75275aa9d1190802b
z2d1c220aa3e5a2b3fd973f915784fc555d71aeaa01cfa46fb1b8afe03db1492ea475a391b56e14
z60f886c930833ed7431e77efa5daa6b7cc8141db2da77ace7079da9cb0c5e772298e0343927900
z2146ff20ce6aa2e454e224fea6a987d173e9c9c8c006dc573d746b753262810b6d76c004a3938b
zbfc417574972068a1a62bf46ba5aa03fc8795e3fe41f8cbb87e18499c6d346333a809bf32c20ee
zdb294f7b92471e35f50ee41728e434e66fbee40051c58f90bd18a0e49b7e335299a7e8006f3910
z2e4086535070a5f75ef9eee36ea832973a4495406e8f16ac8cd16faf1bae9c4072835ab9de1d9e
z7457492bb0cd25628b1965fcb65cd5c612cfec27bc1a6816d6bb4a413d5591e26fba802fafc70d
z7bd5f5814625a1099f62ecbd0d30ea3186ad291e335bba09cb549a7aeefcb9c935501f829c644e
z370c96c2379e73e55715e4f03df7fa57916b87ba383b2d7dc5e29c47ad85a6893852fbf27579ee
zad912f699daf3b6f272493151626e5eca027130c14cb2cdfdcc37c0760f8111f99a41d4c5bb692
z3cfef11b60abf1e520dd52b60473689e896583ab09826c061976b46ff1d665c13e588c5696674c
zf324060f31afadb170579ab2734f76808bbe53929e3f2cf08aa887622df49ca814be9e8d5d8dbb
z659e1f83b1f57fa9fd6234b897081ea3fb078877e0a9448db06ebb587428b1f2bdece7458e147f
z06f22379e5338a2c86b584a55a2eeb857d70d9fc200bb60eebf12b73b739628f41bfccd71d8a7f
za635adc97e75d78540919f7b4c8e83901ffe148f07d59dd491dd2fa37930b85cdc2a3ac1e71fac
z4c7f21478df613f5aae21a54de1341c5b9a0c0fe3fed60daac36dcfd6482989e483c4e7a979003
zeff8875985b74560ff8dc1e1cc4e0fed1aa521a0c51134d2669fbe51b0ced886893c7fa35c5fb0
z5b7e672847b4d3fba88e243e18a4935f5c8ca3c15c5f6a43a8c8616b5ad7c1e43c62e2c115163e
z47c4f026cf4bba993acb21d0318072164e2df80f41349d342ab6c0bc2b38a5fecd52dac074d971
zbe4b8cedcf3368468dd8f8c9755e9ab5cdea7ddb7fdf5b714597d003c0efd11cd898f2a73e418a
z1a35aa776b793c432fac46cdf0fc124c24573fd67cd76a77f0cf687bb41ca03e8fe6245518db2c
z067c33d575164fd9b411a6d3306e7b6f8d09ddce9588c65a52c074266cf2ff73f0402af93e23ec
z4f32a91d7d814242decf22f145aa6e2729798c4a9f914b4aacb14b71483129f20c0fb7f4b5aa16
z10dd1a4e6916cac0b315e61422b6a32011c89af4cca9effb8fbea55d1bc93dfef77a03dae89d0e
z6ee8047f3cbe8d85137aec629ad0f52bcdcbc99e306be187b072efa1f5d45a6c2c925eb04cc278
zd75ce8da83eea39b812f2a56e8288b2ab339c651c79b65cfddfc90d106bba152a22fc453709211
zea735fb93cd386ceda04460ee1a6a4df92aa518aa346b379f9d494206f8f79e05402a90b8f0f77
z1db07bbd20be6648d27d8d740aacd2b03029e9f9071ac26a86f0c19bf8a75f3d16d97065b7be83
z6c5f2537d55509490b2ca2c069b425026b82e4c799549b0c7e4327457e3064b4a16e7ad6507fae
zb54d24c79dbb5f9633a67e7d312f2f428aab1688828720e36ac622695a259bfd0adfd1404f2634
zeee184d0efcfd56afb6cc191f18f9afb087ee4fb25cf2deabe03ecf656580055be8c4eff85605a
z889a6d978650ee48b77124f8dd19bde2a7bf394d0ca0245748c2e07d2b2939aabeb897dfca3691
z9df572ed50a4ee3d34a4b1028355cc6cbe58b0dfec2cb71175aab01f2890fb3d1e26ce65c0fb56
z8e6e49ad9b0355d11d5fe10cb0c731a14dda358c56e5bb7991237cbc7454665b8528082713cb13
zcaafd08a3656fb678cb2a04eb5230ed6665e77dc465c8f3607bfd049524733f79aa0b6276f60f4
z2f1784f0bfbf6e5c04b792c58e8dad362249761bf1325677f30116fd833205c720204ad57c27b7
zb1b068fd3e2b307fe996bff6550301d3642e2f7254742db339a5b69a9702046ff00969c1f38da5
z2ba77cd9b241aebc46d27c553701bf00d79d0dba00f0db4bfa7e1195cac6e2e8b4d6983e5c103c
z98f27e0e3864aa69a44f3f6f7da5cb87879ebd665b6765b4c49ec86b5d465677b0e789d2ca400e
z428d425ba3d0665d86704dd3048d213180436499ded3e813b4371c5da1d5ceeadc479af14cd32f
z9781f833253c672e5568f18baeb70f44850358b29cd38a4507f9b74426ac257d04acd5980401e1
z56b529f49382c725a2f6dca24b81a3e0a6467421117a0ddeb33f489a6e60fab45c3f6677865071
z2a558f82248388b93ff8a0c0ee0c5c9eca231789ed822b2e9a0bb7db085b40f7f9e9dd4046cbd3
z63872f42aa95d7af279ea55106a93071aa6b524c3061f379bbeafb193629d8272d7c5dc93be42a
zb6000c3b277a9e30ae938ef7741f3b7cd6170c882669584723442995378a0ec950a51c74d1708b
zf660bc0a8807aec02695eb0e31827ef770f8cee1f42ce7b1de4c0f81d89187ff11bbb43936d63c
z63918513e544d1eb96a17e8f2e3f2ce8697a3060e4c6841809d7aa2a2b5928517488ea66cbbc47
z0cde91d6a6f91deb737b9783b365fee4f37b7b1c19f87467ea1b50a7ade9b732da1b49a6bd213e
z69f2cccd1d0a4b482542c6733548344c5b8d9200438937db1e41ae10a083b79ddc0dbb4c837ded
z9180effddd64a13a47224702553791101137ff1944aaa76b4225d93991ebdee169d98c8b663363
zcbd48db048325c0f01e33d113bc72dbcb61dcfe463752d045ce54abf6975d194fa6fd90eb6f205
z8400b72afc6dbf0372320bb7b18ed8aed614cfb68ba7151470add3ecfbcc022dfb502061a3a7e4
z41a4c269701078d46421bc25820caacb7c5093d7a72bfad1496cd1f9fbbf5ad2a490593c5d9b22
z002e6362ba1524512e4eaa15190d6744f9a119314e6062a7065f8b00b9e1a9d39c92d9ee92bd9a
za8d00e83b12afbe79af301a9499fb21bc0d3ba775f1485fb9b5bf82e1390a3206dc29e54d5d71f
zb2e11ab1a62e7383f84640600ee56e09a26b4c5519d09c34fac028934fe2f4c862ab652935d4fa
z3ecbf63e75e2189cbd186bfb95c2c472cf68800e8b0a429b69253e9faf3b0bd0d2f190b2c9ca1f
zc91bd1cd50569b83d35b86122d4d88dcabcf6f1d24dc82f08c7f7538aec1929dade3203605658c
z13d7c0a9db8c878080ba75c67bd9162667aada1565f383f8b7a9bf4f8a3d33b5ee479b6f22a794
z958f3beebac85ccfe0c3a05c7d55262dca3abef6a537988a5082dd8ce2dd35dccf33a7551662ee
z426f2a68462d011f9fd9ad961d437f2b9867f1edcc3711bdda391a8d65163b1e7cd435c0fa4137
z50e5e034de33830a57e1c55923f21ad724cc190adb1c7615b05ee9fe449bfb309ff6f47ce645e8
z6540b1a920770f318a1031d58f7af14ead98af88d9ae3887c19c62a393c21b3c2622cb686adf6b
za3d8952b5e5c2985e472362d9b5bacef9477f9a0546d4da4f1e64c446350351117a52c0a6be2ce
zdf1ec1f923212734065e06a4ab55d6ec37c57db3dc61d8529598cfb62a3180a3373d5ba7f5a3a5
z51e454d61ee40bf45f64cd089bc9021748d23f4b30559c6c363b3ee31beeb00c0b604dec4fa3d4
z2231f323cf4141e7bc58b4969763728edab43d1e80267f62ea238ab5bc5a5a331188ff5321b03f
z931ce5583d3de351815fd1dcbc073afb7aab625f40bc25855641f0b880c25f32e65760f821c194
zdc934e55ffb2638cd37d21548b54ed856cebb9ef17dd07f8de61edc1a9906ff68f9b63f80b44c5
z337834754e55022e3b5b7f9c5ca6cce88261ec0829c9eac42765a9e8e8cf541b68630bf1cf97f4
zd0543e5ec15fdcbc394d2a60cb159651d0298feb95f428146d2d74f59df66a22dd2521d538bb46
z84fe27a551c0fb9754f578b1b58c7009bda1242b125f6a45bfd8f6e86ddf1b33f0923d28dbb446
z8f1a70504c5a21cce8bfa859f90de96bd6e36f9f3a68d3329fd3435c7fc8c52ca2304f2ce44778
z59c4b2d6cf2a26adb69ebd9b024aa3b4099a951908f7a30f3f8cee8faec07ec769ec650dbd9787
z08cd3fcf0af315b92f3b089b63592e1a5fbd59c9be29cbe6906cccfc24afd761311919cd31c84f
zb260903d9239e78bb7b1b46671c9079eb8db856b262913c4df4e9ab07342ccd8a9f4f3b58586ea
z6afbea1e019c70e746649435b1bfa0eb7ccfafad26fd4017595173801938406cfdf7bbe833c93a
za43ef6962d2564348b7909b3e30ed381ba1802dd92f9265159c14a64e5ed417436d7ff6b666973
z835a23566c2a4a395b77951ebff2677895692252cec47499dd47f607d1373f424f8ba7cf3e9077
z7e736bd395307e69cbafa95157d0e9f111be4e8a4cdd6eea6ca8d8a20d3acc0d02e4b9a7a2d61e
z9060619c97258400a70c0c65400ea3728328608ad84a21f0c589fb1e543d292b88e0bde6eb51b2
z240514027f6461d36ffd0106f267ef4b601c94847a926df8a7566f2bdb0a3b790bd23015e8cf9e
zd33ed8f23d762f043c493e076c39b258b06c69aa6986ef3300219ea361438a9ccc93baf4196528
zd424e2ad4ec47828cb542440ee2f73b6da120a2a804486a044a7470bfe1dbc7ba582f4a5c51133
zafedfcb32c151f3ff659a40e26f54f9230558bcbe2fa930917a049eb1e1b60bc84980981804922
zcabef86e9991296d32a9886434de3584678fe867aa231f2c7689e4b9d57294cd15ba7a8628777b
z8b113af8189516d9db5cd8bf27eb447628eef4216ca95d0801b3cb064bd17a36bc32d4e3df56e0
z3184e7273c5e568a66135a089cae49cc80d932365e07df3bab726b7c51a28dd87be4f78d0bf9ae
z971dea8a2e8772bfde696647e2614b714d3b7a0c35c5045d03f0d1023e11a278f4a90071952869
zb520963551c954d6f366f7b5dc1a1de5e87c25c30dbad2bca85469e2c3c5e8f2274114c7582b22
zf2aac57d5f38c6d59e834040e41ff58591ad5028c585787bb4b648d2842615bdadf7ad76b932d2
z7be9f98d8a0004c6333822c21e435f4b03e2bd1067d27383f6c03de5019edf8bafa243fa12d05e
z52f2c0b54e338d749e7e04031161e0068528602219fffda11b925e4502b1fe13ee68b99eca8e95
zdd4e76f524b6a4f4e135a28677cb537f44b67932f98205a0ac552fc04ea3c7cc9945e6a18b43c9
z08fc10c1e5ee0c87134603538d7ee4d62a8d43b83e661f9c861504b8fecc311b1038dd1eae2178
zc2e7a03338a930bfcb4efb02ca02976952ec4d7fca1f6f8e0ddca3e6434c4bf4c8a3aae76b6863
ze08db45bb14710d2b97ca9a4f01f8d6b5ef99a09a5df16c61b0947084d564279c766b8ba5e5fb0
z956658758ebbfed035184a06dff0291ceac864f623b6970f14a025f8e2abe4826a65475f7d8caf
zf089296dbf21410aa32621b7f6ea00c37f13e4f81d25fc0e5b6faf4f2033012ebd7d2d2f9a7ec3
z0a9e05a6394624b4d96b5d95a48bf4c18e95e891f7a3e12d8e96b39485b580087cd19781bacbdc
zbeb66291060b71ec59cd4ce1bf40131bb745e77920a3c01344d137836f219e4edc3b5f5a94476d
z7aac1f0075d00220cc5f983b8a8f283dbb23e2a9afde5d8f63409c6a226faa24dc9ad0fa853d5f
z4990df5e8a0e5843acd0474fd8ceac3f6caa1981af3cca21f9bf37c8559a250e58aed41e015c9e
zd7a44cb6228324de2a489fe8ef9ead3059fa28155ea5bbca59515060e6287722bb3e72f350022e
z76345d810d813285c166c7e595f5ff8b30dbd3e0f7b0c7766c4949e0c3a4db6a5c31d8fe0980cc
z45d2dcccae48c0b5bf72d6fbe75d76b6c6ba664bd028dadf603f78b2103d6794a143c1f99ccbd7
z72f623f5200b56bf36d527c00a3571ead84e7c3a7d764cd2ed856cc6363d64bef96df27391456b
z1b26e3bc4bd240107a1627127a0b16856128c5952832657e4834c35bd0895096831b5c428638b7
z357914f5037a107b1eeff66eca4f815632c2b7fc841ca4fd01674526a8f84f03dc73a73f73218d
z0f24aa5ab4448bb2fdff77d85162557baafdfe90d39ac32a7fdc9f71979a94bda97c3793f8eef3
zcdd77b0cc780b2b23c7e178eb1b7cd5ad358bbde4aac07df20a615b9755b7905a89104b23544ed
z8e80f2db48ee72b48cb5ee079ece4dfbb786aa390b065c7f11c77c6ac2b05101a8906264aa5092
zeaf88a24174d5e8452a14673da984241da88bedf0a87309b4ec8540987b213d1c4285cfc6e4ea0
z9f18e3dae23452f9edbb0e94b6542ea4e80b9bc8fa8d24cb1c02a7b8b75856468a15c7d3d6faab
z74d2d2764ac9603646d895b01d6dca9acf11dd204dc5e75a78d28c35919fce3a482c8593125fe4
zee8a0f6170e8a6f0b36000c728dfd943bf5b4d038ae7d7890d83abaea6f1bdf6331ecffb2d3d49
z8b50c73205fe658d35f6b648706c2a5d2e8a86c720946bd84534eea68574746a30e039425be828
zf2a7be2272a6bc536aae95c7be54f346c15429e7297cd43ef029dfe25f7af4d7d1cdcb3a19c241
zb4460f1d44d65c47a798dd9c7d736bfdbecf26ddde32b7f9b0f2222066664b50b55f11dd620427
z694097fb99929389a3c89c7cbe20293cc8c62e38b8cea96fdf2d9fcc93a12aa8390963e2ed9b2d
z76093b4468225439c82ca14445f4067c8469768bbbcee16c460d8b3a8dd66e100dc88e9dff86dd
z9d84b577f45688f20ebb2e416a8099503d63f4fca5153279c7236585801fb67b3aea169f881462
z80d9afa23a26eef7ef8925b4894208bc8926e7bc6283d5b80ca4193bab20be4eadcd80d0a35bdb
zfc71a8c910f75bcebde6a26fcc510d6f124e3017361fb664f3bf674ff2c5accbe1932a063f2fee
z77c73bbe049958af828e69bb4fd0235f1eb81707adf4f092d5c6bbc5a20f2c118788d4d581ac63
z86017b0aa4eb91846a205b2b9a47d0a50ab8c332097d831fbcb256ebffd426d6a1a445616ed676
z771035c8f018a3d490e74466300f30705f5fd29b1a4a9f987c86184f0258730578c7dd507b4799
z7bd5d8093e832c57b9c4639ac71aab4f9998ac044cb33fa7a6bffb371d200385b147bcc4c0111b
zdbd058c70ad93cb8251f999a188c97bccac1ed9814895ef69c6c8cb1aa2ad22bbc1b959d2bc9d1
zb2a1cc68b20887eb3a3373d84e2cd54905effe6bd7f1f30379951d7428aa1639065d8491483e84
z2fec27379455dc950b45ca9c64ff783af5569b59676fb1e55e4a4da64e45b1bd7578d27c6142b3
ze1f21183d48b1f6eb3912ade1c00e5bec9015a2d27f6c02495ccedc34197e0b28fa668a2ccc607
zd446ddc1bb32d3e0bb48676d2cf75eddf107dc5dc519b33726218efaf61d1095627b5030861111
za65eac452873193d9b7c23ecd522aa92296bd8cb6d0079e56dc8d233a12429bf3afa38f8ca785c
z58abd715db069e275f71d3c0fff9aafb4266d6806df7bfb07deae54e96798503e439da200dc761
z837e02f9e558fa9d290ceef62622119029caabace1a2eb5d71da229182d6051cc2626b87d58a7b
z4e15ecc1fd3cb4862427ca6920bc70b0baad16d7746bf7916ea1087abcb03751be456d807f4afe
za12887a0e2996060b001a88fe678b797b350c982949526893cba4bbc26e38e0348a0ae1e5889df
z70036ee647410e0b9155d35f087b982cf043f7bbd77c1629e382b885605488cfcbb7c573f02815
zbba1626dde342511f29debb1d86d3416601d479eb4956d105c5a02191a8fc01fe31c0e7069a84e
z033bb4670c9c52ae386f6c1ea06675e0a989b4df4f0dd86ded67d178578acccc1e41048ffe1d23
zebb45df3cc9bbd4a37df3bc0f00904076695066a5e35e7ef812b704520e7e766fe41a94e553a08
ze5c30315d7a0d3166b51de5e774096d7a557d5539f6ee5cf545dccc90b2bbb53b010018f498f29
z57993303a1dc66f6a82f49b9272516aae3c24e6a832e0471bc0811b17d258b131a05855d69071a
z768d750f6d050f095b7ecbf6ca674fb79d44b6592e18426c10b7f29f332390a54c71ec275ed8bf
z4477c8c8e809847783196fa65e34945b6201d010a769e2a3b303e44f50eb9b714ac279658556fb
z09ce19d446a12beef93af04c838fddbf0f499f87b465e7b810b6ec0566328bf0e0ea01c4ce2fb0
ze7a0476cf7dbf6d8b9279d2e46ae650260d988d45a4051ccb35d650c01034cb08a79e318c67eae
z60fc8396fe7613f7d8adf4c44fcfa57d14b2313c0638cdd12f21b09221e1b12518d336713d199c
z0b36dfb285bc18f587471dad01ffcda629e501c0e0e7314b0b06c06c647dd34303908524afef91
z995d4a7bec02aeb295ecdbd1797f4a62ed871a26d93abc6ae5511670e550e716538cd8613f0934
z37728ad2607fe9b57509ad61d888f92df12e21bf027f3aa34601adf67d7bfece606e42d681bb2a
za1b5c49a4af2f7a776a95b03d06ad10b432464538ebedd04170d52c7e5585ee9eb20d4b9f212ec
zbd14538c91835dcc70b29a619e85c97f07558205fcdd1699a032627300df4c695da09928a97362
z3f26636b6302a7b291734d8c6cfebffc88e13b804b0685004dd470b4c677fbe8346b99443f07d6
z4897b46e889a07065026fd519ae8761e091d191e26b1f5273d887ac9a01a242839d29a43a3c43a
za9bedcf10eb43700944e3437b2428a8e210b5019aed111c6638ad4f30a4ad74621926233acb9d4
ze246101e5c3ca7cbf1dd69da53aeb171fee388102b248f2ca7adb972ceda1563e5d4405889fa5b
z88a816bbad74df027a6e80758970acfb5d72f3a6713afeaca90ca03e517773128c907b5ede7310
z2e804cffc3425c0700029b61c4edce4aa97bfff053ba68b8432fb5aacafddffac45ff2360f0682
z163f8eabf1734769199a353dcdb48f57798254ee477c5df44dbcb3607faf03ab0bf01622ede09b
zd33975689080a7adccffd16329f6d76ddcf9e1ae7c50622401cbd7318c324ac7c395f3f424de43
z35f48df926092f7e229a28baf5d67dfa6d84fe9c0bb9f0d36fa7833bcbadcd0c26d9f62f642d1f
z7b1f4bf0a95dbd172d5fe067e4033a3fb863cb9f4215d2deaaa2a4996e544cb0250b0282227042
z30ae79b7299a8f3e0c4167f81f690bab8e4ba16f85878bc5dc1c4e4f4f49b58379619d50e9aa20
z8e7bb31ae17822815386b53805e1a71d9084d361edfe848015a04ab65b087139f5ffa38d703da9
zb6515270edb5fba251b61596be08bdc07905c3e495b14c5a4d1e7e41dfd106af698b23b82540cf
za0fd7ae3b663f1cb192a9e0b98a3532a3c9f888d01225a6fbefcda23db575416214acbf97f0278
zf0b683e77c9cb9548f89419d319e01e009b09e20f034db8fe128d9a2c36e3c64022f7ac3f58bb6
zae30a0a0eb4ff2c79b19b1af4675da02f3467cbf92438bfbae437d1d19b8eddec383c39778aa32
z0df2837810b7e3b7e57acfa62ccd3408d1253d8aa19f8a26bb72c065b645c732b4b85024f2ec7b
z1656a612bb2c267a5a62b241dd63de9f15742deb2b32fd4e029204ee6a11c8eb1e6656a039a51e
zb0e04ce426a8dbcec206080c0ba0e81a511e4226844bea15db488b5ed53ce599440fb119a80d29
z8feb90c289d90830601927076b7352fb61c216a3047a962aac3c49880fcb5e6080fc3e5866d4b1
zc72fdec65b5ca01677605b6682486b92b614744428f1c4b7009f9092a5e9860ee4ec34716e1a1c
z1050991ee0aed38d67d2e94d4d11568e63a96a2c7f821ed5940c6473b436639eb797bfbf1ed0bb
zeaf4a830530089255a507d578400b1a372bdd5875c852cf7fdda1896ce7453325eda056b97a6df
zd7f7a1ba7a60d27886c0735409bb4b7e3e1b51b5748ebb50df2b11a9a2eaf574ebb9d704d85959
z34422a5127fb4e9a6697062724a03c9c379bb831141a744a55f55026e5a599318e6135f95310c3
zf9ea903db928612b4438f0a6dccd03c58574b59b2d042e59a39903950279b967f7d0015df92314
zb53a3cc43df74e7c2f02458939259ae5a061156e6315ae0e7345655005d885bebce25c880e8f8d
zb2c7d61dbfcc01bf920c13ab8eba8525aba31d22090a042dc0cb5c62976ddfcc08571dfc6ed261
z31c3f463da44c8b928c7cc49b83083d917ded5676ffbc2ef09df0127fce16da2f177fa17ed5942
z035c87fc495c34b239440b33dc8185aada0ea178bf23908a146ee191de80f98511a106ef169489
z6fbc2e598d8e9149fc3e2c300527a64eca0e29732c6f3826f8b118a0f3072a80457080a7f90146
z516fd0ba3c93ded7300516daadf4849343ce27cc018a6ce9f364f1eb763a3f7f8700b6a1b02577
z404917f35d2abbda123ff3d18403ebbd4a7b2a55a58fdddf151ef394e6ddb045c8757d87ce2f56
zac681cc5bdb65d5af93df7a8ee2c84fdf1c28bddf5f0f3034d76266639cf7a35544eac475891d5
z0b4c5e48fdeb0b86a4f44da658216977384b4e0788bee9c6994afa94155f40971cbd2a20ea0238
z596b6b384a21e62bcb1b3654e279b5eb52f696b12eb43d0e6f97d9e7021464dd41de71d9d53db1
zfcbc95f7a249897fa9ce91aee30fb89aca50807ff97951df4371e1d1faad2afd3ef0bd1ca4708f
zf5f21d499cb848e52c0a9af4d35b9e286dca917a5b6da4f5450398590e58e057b39087f14ca8a6
z67dcdf6075ca50a7366fa66d9763dc8a582c9f8028d28470a6cf8eb1ea8e21368e1483826acad0
z34ac5819acaf81c7027c789b266e01f67bd19024e21219b3b99b94bd7fa24a81a9a361ce758c4b
z243a654ec0a7d3b743e269f2ac599919d2118135c9e782d40f6f78cd7e6b2788861b88aa82b3fb
ze767b2f04faf32f0c6cf89a2dba0d544b9b3f76246af40ff320786f30117b053d8e19bc84affbb
z679f9c2c66822d2c0c0679c3442e41dfef1c89838dd1aa42bdfe5e5640f39d27eb3119fc7cbdb7
z9e70a3c6dd9ea70e58162009b1b0fe4b355fab28f86cfd9d9de0e7430452adc08fc4c2c25a1f16
z9ea12322bb3017b29285cd53557b348f918c06aabfbf315ba3097597c075117d3f6db8a2f9d886
z4d9f078e4c94374f445fabc761db3bae14a4efbeca42a341f20c093f75abc3e9a4b68e18a16d16
z0605a386bd9e8564fd8375fe2af0eba57f1deb536de764b0a9d69d6f74435a81e0a43128fc68ac
z97e53d2ba38db939b5b4ba8ebab3cc87cb9fc0c632c23e8401cc1eb3382188578b6fb8ca36aa0c
zd4e67c09e1b69b53bb8017fe15bb966657421e2f9ee9a849da9be92c2d0aa7a5331c3ef7782269
zfdc39e83b787b8cecf8897dfcdbd0c8e29318561c01ff9e452c60b7dfcc5089048f381ba97d36b
z89d2eca9dbe7bafdb8c26212a8889d78974edce71b5fa9b96e9d97190350a24289d13570a664bb
zca03a82a1c8bd908dbe76104cbc06d38f92c8d6c1bec58f53ad0d8345818d40f80c5d80002dc54
zd4e8069c58d73bba3e1ee3abfb082afede8e42ab261c366657067754bb5f57295cde14710ecf34
z30525e7fbb84e2d99881d76ba7fa71045f539c39b05b1511bf9813c829aeab1c8041c8ee8ca947
z7f2fc2a45e32d4d3a77c25d802932b5e8732d771c489316cdc9e9e9dd2aecc3db0c1b320f0d0bc
zcbceaa25eceedeb47079a437e7a3aab57ee55cedbb71b16ae2af434d69cae011b2d8349041ad4f
zbf99e5afbc2b39aa2fa7d5aa75bb3cac6ec477227e114ec7491f20d7729bf7198972ae0c97d3ae
z990d222fa178fb0a46865e65f9f3421ecd7c4c1ff7676edf3b5161aee14ea22b9e6ff166984362
z5788f3bac739623fdd81d26a4da6b57d13bb3eea80fd7a318b9e0ea70c59740a77f960576904b6
zf14483ebd85bdeff5fe0fb9a056882b91a5690f7cf47efb1076a03b3b300202a5fb1ecbead7b9a
z0444012ff29cff76e6128551cf5482276fa352e27e30a551c337cf8cf1f07d1c85ffbe889b45c8
z724eadcaaa3c456d6392b35c5cd12fa98a15b6e24204caf3b953d8482bda622deb99fe1a5ffb9c
z34c2cccb6b9f4f334c9945725e055bd1f7052d1710bb29acd1924cf668b947859e4c89c40452f6
z9519fad19be08560d6ca88c30f0f1ae4fff466476c2c5eec21375220c6d4ef8d17f81403c3ead8
z5d45d2b9215d6d9ff8d4926cc14d3217b650adec2203ae87dae17e375ea87b2efa4b8e338bad66
za61faa0d0b435ace2723ffac49b6face7c87211bf682981fb9b2b389f4c923b838020056beb935
zefff3f6ac77a86868c8f126510ac79699b6cd5a818291d0651bac789d6d422a374a2673bbd0500
z315557d397f82e9a62257df04a44851303e720b6b6949504c5460f9a4d1c52ba3dffba5911a9a8
z7bf5542cdef36ea7a7b8415bc51850dc8da199d55f761a9e145723b32796465d51b924e7b1b6bb
ze06c67b522cbda0ab3f9bf91cb8c72167f644f6d6139c47766d1965fcf54b7e50c49a09f577393
z0a075a6932c4b136c366cee768fd150632e3f7d03edf7883b5ab0615d44f40ab2a1a3bfa188e6b
z26906c6068f4e9add85fed985e9d62436950ca0fcf88133e0443ad51fd7fe8624b9c28aae41e72
zd03ec45e76d623a11228af4309e811947aec14b9a3db618ec99960531595b7e89273147d4238a3
zb29bbd5873bc66ca8ea85c511b166c32ed7caf6f3b705682ca102c84d0f0ad093e7f1eb39b21f3
z6fae2e4110199aee605340090fdf87ce8c7540fa49e94510c17ba6a980be5dbc7406f8e11568d7
z911d550a1265eafd04464ca59ee57292cca4c063ba395973e89b3261c0925b2360fa4c3b9b2c0f
z8a4b063915a0852605ec74d855202d2dc6cb80d761a5de1ef5151fc25a68a67b66e733dda215cd
z8e39c4b8a3fbd23a49b9781496e3e5e32f95acf8ef05a3dc76828a6686e42a19b1cc6045e81067
ze3448eeff1b464cc2aa2295a2336cacf138fa78268bb714f90f71984820ac13863ff76a4c1350f
z8cf1a429205bbe94fbb816855472f39082dc9ca8e3a74a6f9907c225a88918f229511a903a666f
z30f70fe9a79343d5bf4ffd2c6ed65405c667a9820279cc86ba0b95f1e61ef27b60526be44d82a8
zaaf43d409d6a34d554df5bd82bbafe8338f05d1cd833c81df404a677aa7741508b47e6b9119863
z4a22c2706a5a12665f87c59a6117d635884e73b8291fd5465a76493f90e6fcff03a64a7c0273a0
zf248e4e7ef6708adff68a1dba55ec4b883d53d3235807770bdcf0fd1cbf31f536b96177de1e661
zff8c6232c7f4f1d3629d460c4408871d29d9e6646ba4d3722cefd68bedd63754cfa4bc453fd6ff
z811b4fd3c2b9afb97553b83464275b38b8bd4c4e755be8b28e0f8875132879773ed153dbdc32ee
z756293efb38c05f3e0915b6c2d99a1b4037078cdb87fcc1a449db7efcf24e22f1ac4e94060a68f
zd2f344fc994698afeb929020281837cb6151a3c05a9855c3da8de6e77986cb792c13d496339d32
z03986abd5b59e943051777360bf1414e3aa0db4f356f3d2618cd35d734bbfe256643ae4b47d5c6
z48a785b17397f0b57a7d12a7c501ef49e9995ae63b93b60b9583c70112101e07d42eb3d80534c9
z0b79ac17a17e2e60cda883d973c5c1ee1cf22484c23a979dbce58c38f34a805b993d157a2c1793
z566ae353231427571f8db88a95c45be0ceb83f8eb0a9d12abf9d23bacdff746243855621860467
z7be11184babdc6bd20a5d1f9edeca9de122b36fc54f1b7a2bdf8da885686b7b9c8fb13f09ae0a1
zd3bec72ade5183e263aacf81e86afd3a29230a118a4827cc7aa52453ae519df233c60303a9ceb6
z9f451c988b091327d8470c5e20d2bb2e87eaa3c57294f7ae8a3b585e3004ac23a6c6780957412a
z6cc8cdb2d73582c075bb0fa131cb683d02dd26a41c55d154f8f5a7f40fa6a0a62c40256d8c6a17
z2ba5e75311731f0b3f24f083a1a1ccc0de02ad56111b26f253ff927696f6ebfab349c09281a1f7
z5d62e80e5ea619a51f769ea9da237ce968cec08babbbafd3310063737855ec6c6bf22ddf8b279b
z8663563e18954af44c263979a629fc01ba989b9d222c8c0a116b7c5af1089df9e0385e92a7ff6a
z434107bace3dfbb2f68f49e0f8acc86765a4f772eb3d911b3c9b1f7cc848ab4638e31c6f877c9c
z39867205dfd1d86d48ef135251afb6c9056e4e196410d7736c6b8b5718008b693d55bbd873e424
z5601efe537a8a80ec6abc6fbfcd77c22e51f7cb423f6547d970fc969c9ad0062633130adde4bbe
zbe8da1f8dd9bbc754bd5a4f11ff542332689963ba2c4a048854f805b0736d6cf0eadecb3c4037d
z227feb87aeca4daf7fd8a43fe8d009ca71f30cc6faa861ee3a7f4421b6127bcc97c4b8b5a9cbaa
zef7a9150d2eaf3e243797e792f8febe259d4ca2dc79ddeb87153d7354c1aafef4358b3b64898be
zae8a13331310b709602deaf50895be358de173e1d8331c92e548af070f7f70c03593c41527e6e9
zd48ee727fd6bb13e5702facb6f884955c2edae2e5e0007b1f73b7e86d4ded04fd98208a9a7961e
zed50529734143f6c62cdbcf3449d9e849041bd584b76bd364b6dd6d60d54adbddc9d6beae2a5b0
z509e0b0f7d79675d44300c743744d459c2a72acf5eaf09f5f412187d92ae9667e89827eaf49372
z0eb76341d02679bf5b0464d1de0f905d712cc28f96c3c9dd3652309c16ce08b7d6c50f58b614c0
z0276cf3d975a164ea17caf8e1fff2d2690c1cb2ad37a892ccf58492dd6f281955a20ba4e88f3f7
zd6e9b6165ffb7380add8dde41f9bba2bac9b082000f0b76001f3ed7450f359588080d1f42cf17b
z3f572b879b877bb724464dc169210297c105d89a977a827ecd88a122b5e0b18783d02b6f9dfec7
zb2cd6c7048183bbc37f94d80e3b93c441a6ce13727a25a9a7dec82642029a86ae2aed5dcc4e040
zd2a1a0836de46fa185b968fe0c598ebe99152d897052399d3a3a7622d5c01644a1693a9dc64064
z17b7801b5dca9bf5477463ae3c2ceff4b6031af27fda47fea651f9408d74e7b60a4996e713bdff
z0c0abdeeecabdcd727740e19e4499207360d9549c9d84eb8600c429de7ca883145bab947cd79b9
z2e602ee8454015ebefc2f4538f9b5bf6a20dfc67483c7f50232bfe17b5d287d1ea931e3d2d73a5
zc7d69717bf0bbffcef3febcfe398595fdb198b0a1c4ff9a418f50c5084f484fdb4a3f913a26d2e
z108fbc30eaa0a4e3a2291a9fe15d320574c8fd9caad2db60dccb2ddad5c3a99c1e904424293e5a
z1fb93c3e782f895a9aa8ce4dcb48d99d5a3eca0c4a71ce3735fa5b212918ab46b1dad6b2b2d669
z302ed083ad46b5a4c91dad50bfab78606dac6e7090c2bb933090f030cd22934dd29a445c8aae45
z2ee32edaf45198eab27dbb42c276db5ef374f22f1db12848ccec46dac8bc027e366320a31fb8e0
zde80ed25ed2b5d6aaae0fd26d01fc68c074651e7dd205d074485d45a7e94137455650656370cfa
zf123d495f6d7fd78ad5d3e355760f0794211ae1b9bf9c52103b8bcd6e01ae65324530b90220f47
zad4413d3d32df79fb045df4929c9745dbac5111218158d53f12f7827b32cd02f029af934298515
z7d95a5b9d09ae9f31e17b50b2ec8e1ff3389a78b0d7ded5ee72e8b7c3aa4179f4c566c9b8c426a
z053d9786576625f863eab61eac68ac4fe2f9ad45c9ef3befe02c527bc8fe1262925105c34c14c9
zc634f5a72d96eb25d48e3970d15aea7f47db612f686a24ab6604678787dfb166f8e7f46c0bd1a8
z0eb85b44ed6b5f392f292da63030459920000beca233ed13e692b1e6441838ccb4a8702c36fb59
z97403c83b8dcbae855f784d8981efeee08a624d85133561e496f2f0581091dcd97b798ce8d8f3a
zbc0cfb98791d6e28f781d8250adcf7288c90556a2601f938cb8ce9e87c947e13d3f134cae7f89e
z1df78d4fa18a998e926879ee822384dfecc7049366b6006c0b831ab240e87bbcd89b348c498641
z2b61af396b904c276a3cea22037c1c4a3ea98501bc8ba21219ade636cd3713f0d7d1d835c93b82
zcb0338d4b3fa7a9bf8ff4abdad5caa387836c724e18277b853c806b658ec14cbc1ea9d38a0732e
z19d45e5b200c817e0b54465cd04c3dda71cb2d61b7ffb6de49a6569176043b03ec6f91b5827169
zb5e2b91b000a1d07d386a1118d42b646b3ff53247bbc1f415ed56847988a9cfc5f7a458ca480bb
z633a07a8822aaf5d3aac5ead174d06fce5826e670860607e750bae3d4f9f2a06b24da236d7da6a
z0e465197850a6d9112502a4a9ee936ae9483f557f441c307dd090988142d5ed83db7bf01510432
z114f9e4e64793b2a1b08f9e8fa3413b6712d5104d2c3fd966261e79a6668934698d5a2fb74eb7a
z1eda10bebdbb59348c6e6e6f1b7b12e07e9e4d4334c2373baa76c2bdc114cd3e52fdcc42b821a7
z60b52a447ac8529c36660213d0340ea9149b8b9c294506902b327c4fd9b38974fe5234e2a2d62d
zf34a7ce6dd8edeb35ad889e277a42b815a595815eeb21f4631ce1ba9c2e1827f9399ae7bf40401
zf08fc4eceb95de1350695f1611393fa8a4abc6a551ea6b2747ee0877556dd3b6996243a8143f09
z8a7ff53884163577b93a7385c03ce05fefa90233269cf90cf9fbc1c782c21994965b903f2f5748
z0b709f3c063c805dcb68a2c83a99ffff950fb846814bd3b4cc633f571a653b1feb037437048e56
z74ba483d64541e9bd0343cdbdd7dac79a488da1cd7a50b2fc626b81073318a7a6994beaf6e7731
z102a1e7c40c4c507aec97395edaa183211f2ed88e275cdc02ea4d3619f9087353325ba36fe7ac0
zafc18b9bb94ad93b35925c084f2fa0ddcb900013df66aee9f5e85d817357dc449c69a9f72d509f
z05072ec05faa9b4791bd7db9d9553ca47af49d4ff7021500232a74dc80be0a7da5e90f49ee6eae
z04fa1bcf427818b664ea350af900de6f48e46279315012e5ea82cb9cd08923c01709f829a046cd
z1ee1c778559e2d892ade870fb5650a8032290154fcf5639c92be0aab91b32bf4ac438961df07bd
z4ffcdd2dca57616f11287427f0f1461cf046be4db9dac47b955a8eb88aa1a1f4f242a90760a37b
zae919b185430fe62a1945e849f189b55773d8c59f4b707c02f1cd9182073ec9010c64333a27371
zf7f43d9416758c91ff81e001731b68ee6e1b42ab076e95b3fc2541c99d41a6854b28c44bfc4c69
z74d9f052c1aa0c1053eb87331931168706f2c0c51c0a674f33f9514d2257f2010d105774c09627
z5ba46bdf60e8a0f50818b36e66d3699695d6cb473e954fb0ec908eb165227786352653009f466c
zca847bdd0ba7b37e2253a98ac6584bd73f39ef36c8590ba80c19b45379f207b9dc187ba7a07b73
z96233b17b58f0ee37f0e2407f7e9a2cd66e0a531664a59ca4549626b149d7b5b6d17237008bb69
z84a64d3fb3f150d4e856998733ed60b29707c21ac12bdfa025c577fc77d34634afa1f3f33ca4f7
z6e959099d34bcf28f0c305dfceb38b4f6e1f93f1fb6da2a5894b3701fb52d4171c4e8fcc93d908
z8e869eefd7590ecc66a46bf444e60dd731e9580faf2fddae4cfcc10c52ae60f7b687685ed7a505
z35ad81bee77730bef93674bcda9d952cb45b15cea1c139ff118aade90512a0cb4b9f7a38c063a4
zebbb37cfa8f377b8a45626fb462cd27df459d312f08849ce957a0f8dc3db67268d28d9db6a46a1
zee846ccbf8a5973f01a019681478971ca8e9923a41f1d26f59823eb28979efb26a36db441f4ebc
zcde6d28066cc55ce556f991c63f88cb787c3d13d7bc274a137242b62f434f60eb48e0c1a0c29ca
ze956b3ff8e1da911e9d8f728421c69c960457fd1139f383f43cb7d331fb58d83fcc31a11078434
z96b4a115fb6907920f3ca04d5b79a49c728bf737c0939bc8c0ec262946d703b5171eb7475c66df
z221a3c3e18ec8264a1df61c4a847a96b8a659489b632bc966eee01b378d90a2be53cf7a6385383
z6678107d24adbcd2bfde0d660466e4adcbf5c9659be53d1698754456d7ff99125333a586fc06f7
z1fb3ae7c75c70d8ee30d2943caad69591a389e2b29d60a7f0a314e5a73805ed46a308dec94cd59
z4952f6a7ab6b6fdb5b86a5060dc607a70eaae734450bda165f29b47fe1afe7193d9d9368609dbb
zb26e1d736ec01b9ea50f85c28bcf9d79eb73e9bd14fdf03b9e34f7cb922d63b09851a5836d6602
z52bed082fc0d2f56b27bcca87b4739d5be9ed8c6f7270df2275aed0d9328020b4b3200f5c4e79c
z84a64df5c65284cd6415e3fa4eb10c1266d57072180151ea54884d1b9bc57e32c8c0b8065de221
z8149fbb1f0ba256e67367ef128dfd2535343d63f68a6dfa3f0376abcb77adfab0805740ab47c15
zc492cc0901f8a55740796996de7f50314bf300cc691efc8c878b3133d9ddcc31bdfe5c22e6bc9a
z9ab0906d72b612ef5673c3288fc40a4598ded6735de338494c4e4bcb74fe47265f17c81651f72c
z03d7dd402067da6bceff7b8e6472593a5f5279903249109c25901501e8e2b998a7950855c26dab
z73630e0f03bb33be28018a9e6d8d3e70cf5895bf96876b79697f6d62270b47a6cf569d7960fd08
z3192b17605cb0d4031c242624dead85dd8761c83fb54bff4e6fff2f0ecaeaef5f2998ea97ab230
zb5c970d9c9f0cb0f9c93e59fe9041fbfa3662bcf8d6c41749f5309248dd6df93963bfd3acfd650
zf3178dbc5f801ba328263afda12de1cc44ff5fc50af8b4ef6caf27161d83916a383aaba64ebf1c
z46447847b31ab354e69f432f102d97ee714f84896ee5d3096ed0cb13a1a4eafe31bc97bd7394a0
zcada37743359900378eafde1b8bcf1f8ea55c8e990c5250e05e1f87d6df2710603d435d38763c9
z09441eeff650fd504abcf046c330c7e639415351c78e79adeebb1ecf06d51712b4bc0d35c17960
z2d9d6572b3eeb3e4ce5d7d43e0f7764499beba1820ce3bd1fa4867d5a18fa616d3e1a5ba25bbbf
zef331f89aa1c705383f15cfb91f1b150a452e76c87f43a870c7e21ace70e7325541608dfe89cde
z0f549ad03797ef098ff10f16aeb9252d6ceaad2bce99440e859161a190e7f541cc9d339a63c7c3
zd16385fe3e7626ed7b25e03c17992c4db84ca808b1d18a6102763cc4fb777cca6acb44aeede526
z2ea23afa7757b02a2491cbe756f606e0d433e289f626d5e936cd90bd37fb5ed59296ca3ce14ffc
ze4998d4660b4a9d06779c0ef231207135120004c2efef44b0ffc13bd557ae3bee3f73c371b6f65
z03bafcace4fd6e36c30cf494ccce5c35cda218703da34d416eccc2994f626a85a31c5aa068ddc7
z75649e5626849f6df145dc802d7c21d4f99085cada4d70655aa8b34ad5db98a939265733ad541e
z3dfbc643897030a9550659bab7c571bd7ed4212acfb9242843884e9f663cb015b624cf7514e1a6
z613c8f9ded5aa5dbaac0b3302b1ff2302bcf261ee3d19ddfded5013cf5239c521f8c42ef9ccb88
z4715dd9679e6128eec6fcbef3f5530081b81e24bafbb40b1712ff3fa51a624a7e9e3ce19c90b65
zbba8d169e5a2de8f1a1f3a6ddb40e338449032d31b7412dea25d9e8820b5dad99ee57951a4bfae
z1305580ae190bc5a4af88f3409b9978aa6e120fb9a73d8fce02a3e5818ea6c74a08ec43879bc74
zcbbf72903d379f6110118bd19ba87b30be7e1215a202e2259fe698251809233fcee92b08e37082
z35223c50cd2cda75f3dacc13c81d12c09ec35c9e8e435d810825ad1a671e5d7c86ed45d6621f06
z38962fd25b3bcefab0feaf4211cb004c3eeddc1612d57c98d7a51bbafae04888c1b68e708d5342
za5f08a5628e9f6157e7543e099dc070a7d116098b5a46bde9bcdc8979c27ed4ccb730aa7a7f825
z6a052717dbf04a2eddf16e268b7d2ea4f694c83f4e98e62c6722a67b31598c111603ebce9817eb
zf266b64daf986fb04feef9d44c929c78324a373e3504088ec629abab2f761c726e48a9e209e833
za61584d13b5a68eb95135b64ebe603fd9eac5428a130944c4d57ae7215413fabe8618d8b9d77f2
zb8848a83a873f8cc7229727effa1abf576e58c5fd9cab1b9f6b7743aacf2d6d522ad2c259e325b
z1312593dbad4465a8eff0b01223d5e20844c57055cdb08f6f7432a7bfb5a8bca1fb5ed5e39ddb4
z91420cba3c2ef93aaab9a7e2a0b77ca57f0a5f2cf82df27f4cb6044dac913342e313feefa8e45d
z2866c833c1158beeed54da9f0c8056ce92c34116eea948fa1d8b4d603e31c1e4d1b04284e3a916
z26ef15aa0aa62ee27ced6342a7fa1dce141f3e3ce149c774a4d243c1160ddbd590b58f492be0e8
z9c743c1a493ad67141591e382a14972bc8aac7c7b15a54f2d9a6cb8ab9ce2b42e496c7e36fdbc5
z497e6aedee6c24aa0dd91073f31a795ad0725948c326b76f676a41658ef18177d032dffac61c0a
z7809e3d25411ad850a4273a80f30d7c8ba08abbfe348ec1a9bf0fffb99c25f3336679b7c665864
zb35f3a312a01e0faa1fb897849cc2bf2215e0312e5b81f34e3589ff843ee993e23d687147efc70
z5161bead89e29e4a033b2226f811fd7ede80d88c753df08e571f201555f3cdf918efa1d9ef6672
zdfcf127b6f887c233f76e9bb97d670ac9c40c7de26904d27183e6e855e8e5d9a23ce05e537c778
z76d6d493640d9b21276a252df3ec72009d6fd1e2bf7638d29ce5678abb270364a890cc9e9be8b9
zea5cfa8a242ded77e9d18686f64e74b436ae4f1a8ebd45170448a97097bf5a2c956bce8210cb87
z5447c7e96deab8665a818d0b42866cfab7a31d83350450b022cecd3c3f6608edf016cfaeb6d057
z83985688145799a90e4cf77a414f866b3560d5bc3380a88c66b1adadd78192b3eb5ab9ea9520c1
zcc85fcb88f6ed9f00cb67cf197b3ed14e917a1081a725b8e35a8462690a7c2d1f0041683da2fd6
za1434a31f31d8267e3eea7808f1e19c2ba9c725452d7a07545a32365a8a05a6de119d2e6e41898
z0230efa4378bc79f9df050c3dad5d753926b112ef11195868313412f7ea944b7443a4b1a3be54d
z93ef1854a15f52d68e73dfbf8e846682397292913dba09782fb06c45446b38b7657c884acaa518
z0014202186d368c80ab80c1e191e564437ae933a2d1dbb60613a7d1de25050b8d7b5b95d78d066
z52ae5c4cd2eb227a59d7c2ffbc33e70a6bb54098d00d49d6dac2fdcbe84f2f0b93d11b39612a6c
zc5e8d5fb17860f18edeaf851da83865778bea46cbe05cd7f09cf237aaa931fefdb99082eb235bd
z062691a1c6713dcd94ee36310abe5b44cc98cdb85982924445d34e08da44c0d6b977e9925beebc
z493fac73fa8b05bfc9b8507bfbd7a9a0e3abd9c32fae2a870d0bffb807d2b07574426737f84457
z6f700c5736adc8d71868ddab74b71e26630129476202a6454888b01c47b038a9f9dbb3b8a9a96c
zf452d5640a8bae8c81370d8a4b1e5580486cd0cf2a8a54cfb1b09a48f878737273d0dd2d4573d7
z27f9fa5d4fbe78273f172d5f2a3449a7910a593c36069527b115a071d5d611e43d955ef0fa38ea
z920412c7199ef4592998eefc2218ccfd6843239a6e41b98112eb39bd140eb583a5b93dbacaf3b0
z18c6f00f34ecf5a9e055f1305c6c5f09465822f8d547cc5d24a1f7b4fea1b0e036dd1feb987c81
z16caf5451ab41d8dd7e165a5f81b9c9ee015f8cda60078d95ce7aa3c70447a2293669442fea1dc
z8268979973e69bd4db21032cc2578f83f64e56b1b063b21e19a71cfe6cd25657f8e8eb5e564052
zc16daf90630c0e8b89367e473e6d60a168f5a0d8e8018d9b4bf5de39794faf4fc8bae4cd3f70f4
z46a1927a8c654ae330d30b2137581a35442ad7ea728a194d92fe4c483162fa28d040cf2bbb7f52
zbf4b9e6a70b25ae17efb25a7be93fdfefdfcdf93e65b2c5ee9feb1e939784fa0f0a08661f805e7
z799a15f644b4e7af19db957242df8c1d50aec5d4b55909159e26797fef4ad7d7aa5a0fd161baa4
z85719e2072c06dfe8d13bb0d08af961e86d6c9195244d85695191df03e5392e9a505e87068939d
za3fe7c6bb6cc0461c64d977534e80b8f39e1f687c1ebcf8323aef7802a1e95532f772646b45260
z74e69c5b1aead22fcf32c7d0cf6d76c4dcbc7248e1a41a92afe589037eb24ddf9ae856ff56c188
z1901dc209fd2b9af119c3a0db6b42988c630652fcc6299feb2baef6a3afff37eb88549ec0b01fa
zd5755f1dc1cc72addb67db6f2ec055f35dcbb551784d0b549b8dce6bdcffd30afed98ee13edcc0
zfb7223062d0e256502e35523fefbe0891cdc1f05a26e38d14ffb3a5bebd505c47bac92207428c3
z17b0e53c60c164e4ac9d8fb288c60c855c3f8e66e6ed1fa1bb38a583792fd0ad247adc3d1ec55f
zd9b60d72962b3ef2a971063679e61bcb424908c75657c20ecb31cf27780a595e73fed54c8b1c63
z77fe4c64af4cbd4f89585508a85459029e37c420959517cb06edcdb2fca12a9b17703c40b2931a
z6ae1cda57386fa9efedee853457e19816f9b120f03a071ef19d86b9c5a9f8c7d92a5e6d4f3c247
zb92dde49f636753cf1fd8c10c0d85264efa5ea0871a5d061344a226dbce80814a9e75a33aa7ae2
za5569fd423e6b8835ae1ea8c36a510811a2391223c12f17fd47a90ab0c5bfe826b76383623c0e1
za897c7736f318aacc2f4656dd4fa18647c1e78508c9acffceca1cd563b7c4c92441bab28b9776f
zd64a36419491471fd81f858a73f47a6c18bc3520d67c1eda7b079ba76ad079cb7cc35af1edc2c4
z34564a325ee6e939893e5152210d647e1e5a0fe8953b3ac14c054ad2fb5a2079e18b66c72e21da
ze676142cf24a40f41d7f2ad3918d965372c7a561ce1eaa074847a589c34a915d15124387fb5e6a
z12ed256db21dac3858e3b29b97e4ae9c9fb07544de3342e074a5589ee6f0a2ff63e76aabfe6efc
z4e20be44dce34506c7bef543dffeefe7c7f2200a96375fb2cc28ce60e7075eaf9bc04d0202e9cd
z6426d0768f750562874c23a5326f6529f2a8f29110855fbf6764feef87fccd59bbf0deaf98ea05
zd2568b50fffad2a31620909654c5f3ab52b3024da058542fe4a296944f081f1bf4cb1320897933
zd05d64420ca9038521145f54fce3baabb9abe2179c7f845f6bd9ae65710cece4fe715957ea7e4a
z4ad6f578d32af0cc9da717ea5abfc6bace64440cd633e96f11f774629345288fc42a830955513d
zfdd2bee45bb8f2db9cecfc66b795becc2defe6b877516511bd1f950ebc8edfd79dc93919b90b58
zcc5ef7f43acc29a1ff326b32acc85a994a7d906ffc0c458bda4d2b9e9e3d2484406b7c75d11bcb
z77ecd31dc795725a4558a5e16407bc4ca7c7ae5af13a109bf236ca57bc74cf5002fa4e46dce95f
zc82dad4180ed9eec2c1f6ef02f666b7dba31231ac55ae30adb35ac7e4ce1c5b37717dfc131cb3e
z0adef8d89d27adc3a1dc3b35c7ba1fd27bcf268b13c68325d94475c33bb3336869be12fa80b7c3
z449fcf531f4e21a829cdbb7d003f8f4c0d47c62b9de6ffc56364cc6a46bc99f96da12223cc8bd6
zd7598385c2db8b86f9c12e55d1ab5c612d09cd6983fa9c4a5161ec09de8e23ce1a8190512af490
ze05cc794cc64b7d892557dbc516e2192ce78ecf977080fbbf0bccfe946d78c9a54b7cd3c48ae21
z33f22acafa101772c210c951b296e404a5cc566f0f89191d5619a01511e1299c9cbbbd3217e599
zeae69a2aeb7e986fc66f812cbbb093b268fcf75aa491d36ed6c6fff56f7a1d36d56df3a52acc9f
z7f28995883aa2c0082720e301afaf1d1b66b8e483f41fade9d0ebc512e74c18681a3656a9c0b37
za74ab2da6dc93e4047e0bb8f9a4828cad005758115c58e2dd7c0f308c5e33df9102409f499ba10
z4523ffae37a403be21c3ff67a654657565abcf2b4b7bef0d5ec249bf238f31eeffc07aefa3d846
z7f9001bcd29ead6f63b891e98f87e7f8849a36ad8c91c85740043415c349be81fce79ecef7be6c
zb06e1c24930ed4eb961220f08fd5924c76382a515065c094a5184a52f0137502ee7ca2fac96560
z3b0044abda7c435e416ef19bad6b17cd123a0b11d40fb0b1ecc8e57807a5415c022b77a887d305
z9dc314071be91df842f8796c64183a6712a3f88614cbc9302c3ac5daf851a523a037eb1c89d3aa
zc8bdece4653ae210bab17d9a4e20e1d12350cd62fc3249ab3e8bb710d6f7034d276192fe4bff31
z3ac45f9ac436b10eee5763d9d970378a0290322e143551a29108cf3f43fd9ba523bc28eeba455a
zb05c3b261cec590610023a7d694c3edee205f353f165eb933ee0909627bdb83f7572e49716ae45
zc9a4889f9568679411751f7b3a34787fa30c0b3ac49a8c6d6359d0673b3e2008e7025134bd2522
z5cc8e48706beb3a6a656e522bf8ce494135d158cbe259f9f124bbdeb00f0927d9c4c47bb65eb0f
z72203e3be6cbb4dcd5d36ebbc7f0fcfe64eac42eee648045a809f927c2d7e7782642ea4f2e2146
z549f0acd266eb7822d22e6714d23cbbaee3b558f0c079c38c22fcfb1b6e5a0d0f27933d684bd24
z99a7d110fde0cd93bcec5d43e0f3e4663c860c24b0f01a36f0dd1cf8cbaec4fa3e4e680756be76
z9f433bfb90e6abe0a0f8d6bdf9ce03b4e37bac06f16178790973c84bd27675fb29d62b97a8cae8
zaa8bb28518de6b722496670059199cb3ce3914eda08f8ff3cf27ac707aeda1488b90a09e5cd3e4
za75b929c590ea8ea60735f7535ad42470c98f13f40a18e1c4af5898b0c15e389713c9dcb7d80cb
z39f8defa15ce4c9e615240cfc0dee646a1cc35921f3e4206811fd3bd776f1243d40d5a549b1921
za3c62f44df3f7b4da7cf2b323a2d6c2ad70363467d33a80b14b5838fd296a9f3e7c3f1f712228b
zf8bb6c483ca16d8742a90d07255b5853ed9221ea36c1d73c95cc19d3804d884a76f1edad1991f4
z778e9f28885e567867b78af7d6387573b857f23263325d1d3529f33e1c75648bd4506789ca0161
z7700b7e7a13e74d861268d8a400a66a39dc1598c5835a04324db272b304deae1c26c9a0889e13e
zc1a322ab6a55f8e894c469d90de49c8ee82f9efee26e32db4ce80bb6951d4def72c9421c3ad166
z0ed29e8ca01203c45fdcb3c2d6ac1f0357cc31effb436701c46969f052ed7c3b3cf3a7b2de34c4
zee4197b18e9dafb569e80d554533f0b9a5b3938f6449d2bd7312a4f2cc8a7397a008dfb532429e
z3adba7b7f270db27beea24d5080eec7c89db5cd5ea1509c9744fb24ff3d5e922e9f3835ce9db2b
z7d1066d270f1abd98f30cec2e7f413536b8876b1517ec6b8c0fe136041075fe356752ce48b2ba9
zdf9d092199bca00686c4067fc23b712405beb4f8ae851b2a6ad4f243f3338ba03bccbc48e33050
zcfded4dfb8a42a21b510635f038259b502e1e9865be5fdf74a108008b44909a7bd103fc961441e
za45621f6df919cca2c7d77e19695e11888ff615da8df50f326d3d93efa6f3159566109d5bb5df3
z853f46a9ad414cba09dbd1a665934909468623efdc4144e4447798129b297448bed836a1f2b2dc
z4ac4278ca7230d707e81bd1fce4dfd5d727d85c52b1933b8410c1c09efc716a68b234db4888a83
z99ac9d7fe9cbb0fa26bc00ea937af442b84071eaad7f3cc4cf600e56d06b3def1eff6724509d20
z51330eaa236a806e6ccf886682efa3af735b9817f2d0c9796db48a0937833fc15d4e8da5e511f3
z7344e5e90a5467d7a900b332ba5c5d0be890f8bae55de6aecf354cbc1005f7c85be73a223f0cb1
z10b0f61b4dcd3f836887722ea92b86dfa603091ab697cb7e73841973b913b2f1dbc21692cfa1fa
z1fc4d355ac963aee39bab2775cfa7e6076edda556dc5fa8639686b1563e1c5fbba0295e4d2bfec
za2f82555c77eca7106d82c64c414b1f7c58db199d664139af1b2b0b99c91ae63e3d577996dd02c
z238088ab559d2075ab09af21654fafe7ddfa921ecc5d3071f57d31d0b866d801197dc49b6ca710
z227ec63ec473f51879736971fd1100a7261104ad12608cc9a7557d22cae6273a3e4727e39cc02f
ze75140dfc112bf9fdfd42a23d376e4d3ca70875139b4d22b0a2f492eb8cbb24cc427093a998675
zb76e61725775ef785a1ed339a42114f66399e51d00cf6f30943a1e1b7cf76adeea9e4b0ad52c70
z16545036bb3911ae9e8ff92b53719d38fa0099386e05d50930a7457916d2dd0ae017cc5f825f7d
z7356605f02752ecec2fd6181495d30f17e41786557b3958bdccaecd53ff058536dcb582e86b8ba
zd73b64fe5766421dfb556bbc0e201a663600341cdaffa4fd0ac76025b811835178d46af0509f5f
zfbc8abf08d15981223659ce3ec9ab2eb564d8a0334521bc6df547caa290ba511f58d487c64c50f
zf3a5d6ad05a40152fe7cd71f45b740e6285d7c3f154a3af2673954d108ff596115bfb18365fe6b
ze9c3554537d59ea7552115a211eb3b0195f6bb01a6be7db7672fdee622315e90b3db9604dbb3b2
z1b1767902f61137a867129aa0bf7fdcf87046b709c3ba56b3ced739ae35c2b408b1a92966cdd64
zb2d1868da212c6c545a473362515bcf8684abcee449ddd889d595013fede2e5980810bb8a36d28
zea3687647713bfc6c77c97df4e52169826aa7d2ea53b615e311219432cf4ee0cc745854ea4ee4e
zc321272a7c7019a1b3c3abeb5f2bf9d67367ddf6f860f354eb64040e8ae695dd6fc4867f788817
zdb20e24777d6c983790c0211ee9ac73c545205b8fec59ac95638a229770bf3bc12c263b0803e9d
z3a81483c01a11e4dc2fe3736a7ac0b754bd53caa47677ba0b2789f9d59a1c444cf620d757ed50c
z9e28e2fb10b86a3b816fa33d7d2c43f3dcd76f7c56bb8008fc5883882a66cd3e2a5cd1f754b25c
z9cdec5ba0ac957252bb578329a0d9b3f9a076b32105a2c6d78654fd786d4c8f71b3a856a2fdf5b
zf61079d8c71ef0695086da3efef7e8b3c492c2e5e2c38567c1ab2a8586308608fd4fe4787d3fae
zc5bbab6cd2ed857ba248eb44c6ca2549a2a01e8e67ea642f841580ed59699204f28e37ccb2b9d1
z54a220d70c0d6b65f73a4913eaa937f7de453be468b6c006cd2005f34331e925fcb226771f6061
z62aade6a6549410781cea146676116091a537f643cf71b24ef6b950dcc427c1c1ff4871b467578
z760a42d3439600859f0c3fb15ff35cd56760669cecadb312c44c2571814bbe223c46dcfd94ce83
z40cf9fee7e6ef359cebc7e5d70368a2448e4754f2e555f6d78c6cd8bdba30309f5124a4d9290e5
zaf83410997a0a26bdb7c1815c6993bbd295eb735c1850a1649048f302854070e7c6d12690853a7
zb20c210134ffdb1f40b5739066e94767f752904eb5c9b7b7f084244e68254cb1d11affe6019601
z712b3bc6a2b78caad8b97ae26f23e0608a97c3cef55984248ab46b44ff0fc436369281bea86a13
z116319c3e926a6a6c0066306cb6a0ae9d91f0b64275f0177bb22418d8eb310160c5dbb05fabe60
zd6c34bcd20a29314c08c039820b591aae351a39cae1cee5575cf7dfb38cb8596242008b4ba2e03
zebd087796665b9bea58bc57b449b5e2bda8c3f2336b0117dd25a7708182173b60c4f735828fe74
zd913b17bc840e2815703adccebe49492fae760a1eb3bb1b73434301c5784c86423b87cf0c8301d
zf92731ac5862d6b8b71bb9c71ab4d361d18d5dc7ddc52d9343a9584dcfdc3f01c7881dfe8601ff
zbfc7ddc24a08f3ad7e913d0a7b2fe695bc6a6fde87c45925ba644d35e3e0a06ca10c61890ecbf8
z39ba06e900ae1472e14bae4522f26e12ae850cf44b02c0fc03074b06eeaf442f29579df1e9511c
zc60b03555cf483cf90584a3d82aeb21cb67981e2b2b6d21715ac7b4fc9cfadfadd9ab5befa3cb7
zf25c5e34df8efb7eb5671f3b0b78b1197b801764acfc30acafa5f9e3b49072830a9ac692e1719a
z63eaec3283a8333ef907e41e8b518f02b80600657a5eecfe57b3636b4ecd68c445d4a0776eb75b
zf798baa9607405c17d55e03a1405ea22f06f26fda99f5849324a89e461e829f42079bf34e581f9
ze51e8f280df55fc4e059ed926720881a6342393567a86edc522e656fb33ccec1872b773fb7816c
z699b9260638cdecc50f26a7b3bd1473be9722f36b37973a05eca203baaf5ddc136858d2daeea61
z10114102c77fb5e407bbe2e1b4ba5f81022c4b352d93c777cc0dfb6bd28e03833268b56162774f
za1000f66f22ce2babcdbef23076ead46f0229fa99eac694c4432e3f501378a4880fde423769cf4
z42ce40ec5bb0c15604af7c4306db010afeeb32a9f7249b6534524446c9ae9d0d62528ea9a6092c
zf3302682d3bafc66d9cbe72311a0d1b78b66eb07e42eb376de4420145882e4ac1898dd00fa500f
z16f9badb4f491ea0095cc56f61062c90a101f19d7fe6811a99d5481285ce45d5ef592a5bae3b2a
zc1866821f6ff946eeca143abcd3a46a862e2379d5ee22ed34ea0f0401678f6c9df7550a5ae26bb
z46b9ab9d5444e8d45a703b73278cee8eea02d5525c7f2ccfab4a299bf0f37b964b120509c55648
zcf7101590b4aa966798688b4d73c0b115bfdb845ae2e46856f4e86614604e6bcb0044caacfe61e
zce3eff3985064fd45befa15feb08ad78b210746b7a17111c1438736ee1d5674e80724f42da8737
zffdde7443a9ff97438e4f18b69347f21b6ce4703c71c0d68ac4ab3bf35f5446a3ad233a8150bc8
z041712a9085b646778b54667ecc809b95186a5fde57c4af554fa060179a34df082e848c1c0f389
z0b6af94bdc979664eeb3376b2d2f737b581a2521f591f7091dcbbb2a67d45daa83e16738763f17
zb57b2250381f47da08e2b12c838279095db90a695f9678aa111ecf65b9712475671a085e6f6bae
za3cad54e6c7186b9cefe99e8525791a87996d79ac8b28115f7c68b0dd30820c3b55a2576e9e492
zeefff06cfd088da14884e95c49acee3fbb57e56fe1265a9e80f5c07096c83a6489b6a94df6d84b
zd66dfcdce22088c6c980566927cbd0ba846f219b7266ab4fefdeb3cedc46c35eff551667819026
zdf9b150188f235b2b02b5353e371498b034fe8fa1df83583c64051493f9bf6b1ed201d131967bb
zf58a9d7bcd64d08605cecf3dc7cbc49e7e1cf7080a236f3d41f4ef7c04bdb37b9136f78462a3c3
zc17c55e9b8b134395ccd7d3f37f629bb4bc6656618e858431ff71129aedda5885f7d4a1a1fe682
z4f18fc6a2f9a30f0f238e73f935a2d84df3c09202ba0a667da2d98a2db19ae4e81bd74cb869a13
z3dfa300a027ff70b82c817a66203276f3cf6b93c4bbd9b8291870f814405f22473499f80d9ba03
z8d416805a35bd658e73ccca4f2040a668bbc6f01d9a4929f82b14e10660177d828ddffe26d58b5
zcfd55b00be7ec3640eb81081f2e8dafa2a0ff4dbc27cf448deb276aa2dcbbec673585416b5ca1b
z6d04e0ee69837aac9a2e2d31957a03f6ab0989b4dbc7f7b73b756c013d6c351e85dc04cf5095a5
z2eaacdc4f753326943d153e01a478de9766d779b452872bde5a7fcc47df99e48b124afcc8fb56d
z35127bd9ee2fc1ab1fb6d4759aff4496a5f680babfbf4fa902e3eba80462ea8b223548ccd52b8a
z6be0e5d230de44ce38d9b6d8ff10ca7dddb194d18c59b53d635c17ff735417bb65efb7da3ca1c0
z0930ef25c1b48abe1a5153d56c93a3505ba71cebf658f92317f7658ad8f70d2595206fe4233b35
ze4cad868c67a1629f9dd02a60429e9e6e5da78e346b436da90a94ce51ae268d4f167a2327c75b7
zb050f79504f3cd736c3c45cafe17ec633c199773ae36f6b4d00eb2f2a32f32a56367393d356af5
zebf88d6e5cdc5b1a8bb6fb6fc3376e307ce9bf7a3da5205842ef9457105ac1ced3bcf816008142
ze1214d47e7e80372d42d5be542081591fce72ad69b3e8a239479c115bdd0ad826f3efc4dc6a268
z7e40dddc34a4a46562ee3fc0a30a0ff51d11bf1c4dade87be6e09551d2496aa1335162b7ab5049
za8f51952053610c71d9d4cd7cd082a6d9ad0c79445927ab829756df691185ea2fb8718510e869f
zef72d77337a065fc15c6b71db39cb6fa4faba77ee8838fcd1bfe247f3fe0a59f8f7cd32ac6cb18
z58dcdef17e1fbafcc40efe1f6773a4c82b5d83b8289c363161c8232bb22e9f9f20029d58a9313a
z405a99287920fab247bc5bdb734a3818cf8d520f885da1cf4a0d99ca8b066d19759823bdb46f28
z4967e2149b59cb30503a62eec024e4d264f744613a52fcdb2b156229115877f55deba9cd0976fb
z296acab155eab31bd2c793598ef95a9de6eb43ec42e1659448847a0067ce3900f56f4341a63f58
ze82bfee2c5594388663c98bd0f3fa66a76c71a874439dc8e622097b9f227272da40a6ef88d5d59
za097cc08d9ecc9c09dae59692bea5219855c9f6aa93eaf61e1f675315a5696926643fbec0c5e47
z7387bd36ea5806c654255305f09e46be672b9b7ccc66ce3dd389fa0a2239bc463afee8a6eeba95
z959d3dbdf07e534a847c3932534164c8a6be3310493facd26d1717867e1a6d1f991c5647479aaa
z745b87d2c4106077456627828a9eb66d3f4170b8e3c282ab7e7baef0115752ca8f53e9dc31b858
z981f879ed2949ec4f242e5e37a2576a94049460077e0c5f8e696028ea8d421d6c1d44b15d3c678
z7bd5bb66bf195ab6edd75208e1b6e6473155364da8b1dddddce4ce53b4256f574a6751ee76a565
zd20b9d701240dcb030b331287053007c3bada68ea9831be0cca60d14d91ecce5b8a248fd14c9e0
zf52d64765e162642e1c7e053faf451a36a3ab2fd92e1c3437e7276f3069f0faf5f7b6b89b17498
z32967dbc924ccadd1b2c947bfe0add43ac2e6e3d7a1a85efc2f8f6f9fcd0bf5cdd0f67fca09244
zb9f0651035b335f3cd3a4aebb6f7aed0fa2353e8ba1daa0ce25487572ac2d9650c46464b8bc390
za9d64b27f7ad16bf415ab6e503e2452011b9a9d8965db9ce1d5d08283441a2596a806d7f8da071
z109d332d969505abbe0a82e2e0530ca04c7cd5eb33757cdb6cda81584dd09d470bdbbc4a8b0830
z410917fe4a15174b24187c5ccc6aadf7bbdb82733b7c33b2ec1e7f7fe83e4db094bd6bc5f4d0e0
zedcc9bffb4f4efa1dcbfeaeaa13b3b091c1d9d352d9818d0e8c31273f9d798c20dd59281a5b826
zec8ed30c17d86e07d126f2314619d6149736f4929b7d1dde78152b1b4ef2e5238725802cd246b8
zb491d7c0a404a6c66c0997513a141166149a564178738dd413621284fa0b23239446c7b2e44d8e
zd5742bb6409f9af3e9e823d96db1ab88c99af3570da4218df604f30ac40ef6ebad4af1a64a6dfb
zcd263b22907c50d34d9e2658f6cdecb0ea6bc640bc756b7bdf82df5e3640b799b293ecc0fe589c
zb6b179be6594655bf15e844d05359077899197c94d09b4ae19a22bcc080d0f82e1a8b1dc1a5396
z2b52bc25583e0f554986c0bc937586a88ba299663577246807e8981f898142c11d3201c7351f1a
zb3125ddb53e4c64f34991363667949ae1e082034fffb4c089403a8cbc7f016e1389b038debf4cb
z447e66e8fb5d12c918844c2d8dc0b0dbd3142eea301f4706197f6b08c77e87a42dc9177b8daf39
z236122e9ee14b38963c55a403ba6f1eba46f045976006e40f3c1e517b8cee6bc24440fc338604a
za449a2c55b22a530f26eaf3b6d9d1527f8253696b30c4884707f7102715957a97f4f87793f21c6
zcbe5b25add0761adf7f694f2f0468f55e80454d8c134a4cede5786bd6fd065b30baf9d0f34696d
zde9de9adfa521ea32bbdd499c428bc7a1b4e72858f8c507db1d738ee311761fd86a423c5e96ed9
z1b8bed41d9fbdba37c5cb1f5dbe879c6e05813e40baf7adcfff9b9f3faed54daf88bd3dd6cec4a
z769e9145ce8967b30a40f64056ab21c8013e2aff7e2733c8d8368fa2933bbfbb4cbb749293cd8b
zebe296d1de4658bb87762dd5f68ad2b09adc0f8a6691e76205bc96e18adbd59874ec88e997a40b
z10329d3ea04916362e1f7d8aa1213e3e8ad58eab560129d717ee4882d46758dc11948c40ececc4
z214d1847101d36b2a61e9cc7eea9ee43c1624d075f8c52f44c4a83439244d79eba89656bdb5e9b
zc5f1d5a82d2dc3039485a710d8de333a1684b54b12473510567203d0c271282e386b5c14c0e38a
zb9a3809e280067f140ccd1dae3302ac45846b21be48a219a5369a1f069f388f6e660c1f4e5ff8d
z8396cd3c2a64af26480a275d2df5743e16883fcef5d20061eb336fc81f21e9973f30eee7d74aaa
z6ddcfa9dcd5c52dfdecbc3624d0a4ef06b755226672edb1075e2e6ae7f31773cde6e4cbb6f0b7e
zc6e61b0bd88658ecc2f35ca6198bffeb905e22ff29902e2f8a1b42b2e759df715ededdbd740d37
zae76390a056ccdd522b5dc7120ea832ad34a0ca5e480e43fbe22fb11e79d6a9e46acd6640ade5a
z1352afc262d81b178fc3b432f1b17dc63de9ef325609f717f0ab073fcf5a89aae4121935e47326
zbca18d317b1b24ae9cb1de055ac3a5664d785fa7b236855a3e1b213d84e14d4663cbf301c6214c
z2e5a02ff01e2903101767453ba07473ef3807dd5b5303e84899aa590a9c7880578b789244a2898
za989c15ae88a363fe032071eca4536d74199b8a78ce9114056c0995dc95a70317d0919b8f01ea2
za3b25fb0265fea9cf6cbcfcad1781ce98628d0a4c12fc007fc88d2d8ab11c5b98351c8887e6d8d
z9b80bde1caa1f403cafcefe5d3e137148105a2a9c2a656052b00693a65b233986195c2e0c50eeb
zefe5d8176baa291c360fef4f6165ed898bdaf09576f992e5e9323e63ef4bd2274bd99d1831599d
z6f0ff0f44086603f998d6290aa9ca5302b13dcff73353b2fc343c3004c6ad26bc8191291503a97
z93453bc077840a629b39d08d2d9ea2c5ee4c6b15749d961ec026c1564d01be42ceb9ed87e17f26
zb8feb03ae1d0dc5872b6b9a28df98d7cec73c71e27af5c4882b1f82fa97f37172eb3363083c29f
z6f7b9b4a9a5ea08f0785c06819f5245ff82fc61805a2ea4572050c21016c30744f66b8049662ee
z9653388a53a15fd38310a6853dee9237031a84deb58dd0a8eee40785e19c4118e901d29317f3d5
z145dd4dd6ab36ebf24ddf133f992b416d4f720635e2cc0bd23dde854d5ab34c130f4cc855c8ee1
zdd00401c4569f7f01862abbaf367863d7b2509a158c4b757d1ae712806da48d812f16ffa112cb8
z770280e60a37d0a91e3efddfd6e539b06d70f3d248f17f6c9d495661f3ac749c6675c5f1af3bdc
zb61c7da122888a441a9e7cda07736f224989c4ef277457ed385bf3043024fce0d8fe4aa16ef2ec
z58ca8688c9feca8b9570c142e2c4d4d8f0aa56a0cefb685242d623ccba81216ed6e2249d0f299b
z95f47be1b85dd0c977317f3c150bd2e5f0dba3ad7598d6b52366deef0b6cac3587864d877ea50e
z875f477e0fd0b9ad9d6162575bce074f4f8b09a59c00015fb916ede99a210195f8355f6d93a6d2
zcd52609837462fda78d3995e5b3807e555d9599242cbf477f1521c4679869275247a8ee0bf9ef5
zcec7e5354de9d99dfff8779d8896a2814476a5d11035888bdc51848f1166dc5481171a3f8ed193
z5406031029c25f3bf234c8890ed0a024cd894f4ff61794cf8cc6555ad190bb6f307f76c5b3852b
z0fec75b2cb611af4fa70a907f8ce858143982a1177d61b8a187cdc462d1f0f3767c157ca626fe4
zaedfb47303350f973663d89e27e766567db2597c7da9f12732cc261c62d1d96cfd1f0e5a53c92d
zbd9e26736d6f5c215996a8be0874587fc10f8cb8027d632c6e01b730da5a39fb2c67874cc38089
z5237948509cdb12363a3c0928c38705e6dc2f69ebef0c8967a452eb66300eb03ed9c38e7127a1c
z3d7a91f7ca1e45e8fbdf1bd215bfaf0679fd3db7d1b5b048e93d8a7fccd7a1f8eb0f7ed12c7a63
z8a63fdd114cc7b9722593a552df98aae0c9afa13549a608c9d93c887084d9ec03baa27bacc565f
zfc52ffe7b8ae456c68b814ae50dc450349dfd8903af21fa59fa6d1146ee9c8f03ce4bdca2c7744
zbbba10d59a6c31852026611ef305e72cda764f14279f7b8ddabd9a307a96bc7fd311e96cbf5a14
z847e0a166241da1c0051c6022c86bf31813c77dd84afae91dd50858b5d0093b782095deb53a7a4
z70fe1002af69745f2b5152aaf451b925244af39da9aa48b35b4696eb21eefdb9f60328055e4025
z33739e0669933b6522c7382ca6f92ed20cb18be4d9b152c5aa7e0c69d461ce96fb7298f62fb2f8
z02c5ad92a05837fa045714347795f52d6cb5542f9894dfd9890ba1b1c49517fe8da1a3760c8b7b
zde1f4302aa859ec229b9bcde2173e8da505e6ce3690cd8018fcacc300efe9df0a29bb285f9363e
za4686aafc32c9c0278372c35978f8195d5aaf36e165ad577c52bb56e321889de5bfaba0d100eb0
z6c993919c78d0daaf06751fb1b1310d0f0817a95a1cec745353cab4011fee9220732ef962bf1ca
z4f3c4ed82c6dc821087be19ea07e04dc7a18081437e210609ef3f0f0e515dcda58dbae5ec343f1
zd041683aec0b60fba98a6818b9e8df81335511860dd481a2d519ef5054d0e033ee3263d9f79e2f
zee86bd74cc704fab9fb75737f4bfb1fe452115eec1d5e8ca06a1140c1f806cc02cc28cb1924c11
zd71eebd0e6ffa3a88ab23bf1d5c64aee6d3ac048be02f8e3312c9203996026ae4d1d80e1be8905
zbcfb3e7af08a67176c5af21e82a82fad885d8c48db96ba9fef9ceacf3493b0c10d704c9b8cb9f7
ze3bc10ec5a3f3aeb0497c4476e5587ad15cc1ced71d309bf2d3123ec45a44303a4e4b23a93b35a
z54a6e804f6a1e010e11edb9329ece03d88b2b67e598ed24f9d6b36709b2acfb61092e748d0a9ad
z4179c1f57d38a1abb62b7754e5c03844abecc3c5ade49dec7b2a0094f4858d2cd56f633f8324ea
z1602368d7c44ea049c421703aa26f9c1346fb1fceae5df3021b25b155ee7ad40cb0928838c8078
z6d5da978eb1e146acb4675b5e4df0d824a50d09c07b350983c2635a1f61a2eb1765761f19ecc95
z6ee93ff1e36a0aa36bfff2e32657bee3d1f2c46bb2d9408203b8e0ecf5c7e303ffaf3223efc299
z739d52bd870b102e31e660b5696a5ba801e5f14a313ebb31affca17a2dfe16014b709ef9ee6c0c
zb7da07eb2ea57f46abbbc1ce77ea39588ec9a29a7bc68084b5cdce72dc71423fe2645a3c0f3dba
z168dbb6165d86ae4217f7edc865a49844411f7fc935e0e6ab762ebeb196d2e8d57eb285075e396
ze05928c3ba0c7a92381e1f5931bd2707340f98e5be37b9ee57fdd46b3a1eeb098612136bdd7755
z2c4ad6cdaaefa68bac382e30e654344c49cac46877716a8714a93eb9a433b45b4f61e78de58c66
zd36b95ad6b3cc5d87127fc8baf1f468911000f64b0c54e5df97852d308cae57990b1e92de77504
zfd9ca819dc96b39cc5682a265bfbd8639c8d442da6abd3005c5188552a1bcdf9be581a159ead3e
zc73cd5542de0bf773004d295ef851cd5d10b2a6626fd1c90418dd403adc8fe8647880f1547b829
z84cbc08f7e4adb728636fbea10428cf932c30655e940f8a139693e5156b7ad8daaeed69db42008
zacade74f9a5428cc6cd0cc04091e2eebb20c8897890fa65abe09f4ffac2b164c0726a0179f6071
z21b74aa9bcc7e58a4cd999b1d732da8bd588fc99312372c80ea839c771a367e76f3bfb48ef55d0
z653173674eae74c533ad8f4a8757d47d588aca13a16a9d68114bdc751f34a303df4b54b16ce190
z827ed7a71de741accb31f56543fb9171f70c27efce0553e28e8aadac9c9548ef01bb0ec02fd981
z81eae141d9d6ff79b833d876d3f6d578d8ee2b5313869b94f7a07424574271a78f30ac4d190326
z0df120ce7014e6533427d2d65ce22c44cc42944c9625a84d5df31802769b05d046451e379ad9f1
zcbc0df3cb2a27fda7451e20e9e1d97614980ed7e5d57c5aada9a9cd25c40c87b71d3ac6e3176ac
za9011fe416b03a564b250dc159d56bae7efaee1688957c5c7e91a0096ea5b8f3dabd4a1ca91876
z9c30c93f58217f920508684d0f31c49034c70bc138cc7dc56ce57cc942ca144a403beb436e4f1b
z0a4e4831909412f4db9999df556e1a0411b0732829a4e56613ccdf77b78f53d68fe6309e1b883c
z1dfd99aacf71b1a2e845bb2a9ec783fc17bca567eab3faadf42056a1aee66465ae27298cf03ba2
z9efefb675f558280e8c2f3be35d7c1428c560a255f1b5100d0bfed58b1a4e477ded75bf9088f2e
z46b6949e375a395a726bfc77f43f30c4d410de9b8a8ec52148b2a86a14ddbe9cbb1d3a32eeef1e
z99bdb0f3d8f88d1e640f03e30f98ee8a37fb45545d136e6fd62fd3950914c8a43390aceca9f1c3
z946361c41c95cd275550ce28f6d9c43f491a1f5b0fa8896437f22e59fb4797df68e52218e20dcc
z7a8246c678723946036d8b9e20c1b3bbe706fc58b96eabcb2a903175499925314514c3034ecb08
z16de68a46967d42a8e1f51d62a0d035c82af6bf22167fa9e52c5c6d2a21173df174630c0c49ed9
z301231f8eafa7618197a6983721ec2efa3e9b4054580ec4dfcbd3899bd3db4c96e14dd31e41ac7
z158dbcd401252a1d4db3c11a2270c7940e2b702a6642839e03f7b0afcbf03217b92ba0d7cb59ea
z4981109d5a4c8e4a4e771362cba2dd7adc8a615b1dd434a7edbce12cb593eb521a696a1c5a1fb0
z176521c2011fdaff15e84a3406ec1b90f8cd1f61f63b47329a2c86a0f4288c6f7b9fbbfa1ebbb0
zdcb47b04488742033f23d7f060df006483dd1b9df03c73086e9f60789ef11aa1c684bdbbfb431a
z2fc5dd69d28bcdcbd7c89e49357a205b5416e9ef94f1ea9012eeea4a165c7c90619655a2cc3660
z15bc2458c93c783e514c4d972c81873b98c4668310ddcc485cc0f6fa7551d43655219486f44ef5
zab6a5fbfa77cce5c55f7731d5064e55b6efb7be265197c6d8e858924d1cdddf098bd32a93e9044
za532bde2e4ec8ab6b7fd823550af768bd858bb16dfee39d96a066352d6e75ef509c88ad6583c7f
z3b3c22b4af3ad14a65708c979cac7a8e227101f6df73333d231aa27899b451cf9f46cec16440cf
zad8d0255fcd096f5e8e3a160adfca6d36218c7ed5332078a36ded6881e80399be868e21cf939c6
z48825b3d4f15806d270c7da9cc646bf26563013867fcfb645627ca20e616fb6e17a72849c8485c
ze297b2708e7216c5f20b87d7ca2ddfbff6bc7ef362999ac2cd1c480a21d61323876ac1231efb9a
zecafb2b0138641cd000a9a8787d4f1715af91bd23b42b998b1daaedceef0c1b97e6a9be0323227
z47540c6a2abfd7a39791d77b7df820d63bdf496fcb14aae8962d95b084ce8216b0118fd7110974
z1cab2f997b83a2414fc0c5ae206c3dcac87c747b22260b6b92956b53bbde4517b4f59fdabee03e
z02861230ef51abac4135c6b1e40256018c84f96fff227688a7806d9e89648c0a28e7e7a0fbe4e3
z1377bd3c251dd1021442e1aacf17a27e5a1837851b22b2db4791497a9617501cf07d08b6cdc34d
zaa5bd1ff9dcfeb73303481bdeecfc99959eff81753328c79e4df489613f83f79912a3cadbd11c4
z9e32e0a63bd5a11b1ccad8914660808f79f813ce6eba663df0ecc471cd38ba8e0d4d5b2b2edd33
zd169bc4ba2d2c5a1f8d4fa07d4a60281ba12a040e7a2a5449d66e0291ad33e0a33cf96a36b36c1
zabcd4c8965c9e4a45439c0202cb16a58509227fd3a58bb707c149a18f8c55c42844a9f2742c71a
zab23f3c11345d6c93332fe0c36adb059df9ec11019d93bcc17b22471c40f9664cf49be07c75c53
z05d68036f53e34b0b8ab35d137741baa905667a00113ab4a1500d1c464d959bc5377dec4fd6b62
z8c204298b56d405f94ae8b77d56c6114ae87153a49e61fd324a808c0b604d5f85add1a70c66ea8
z9295c17fb1768c894ffab8eb284ffb8215f464d11aa8eb14c41f4722855987e8c777845075c3e1
z47fa606acc4964ab0bb44f9f5f14ffc131a383c5f7efdb9028135f161fa397bc00342b30107505
z04d94c440062f1fe963a1413f3927b2b18dd9fde7a4f1264f897fb24d37d9a6755d5aaa331d295
z27ad15f87cc6d94bc8f775204053ac9e00a9d856ce7944c3df789be1787518ce85c8ed9ea2f822
z88a8103373aa8149ffcfb0dd0309b88b8912a740c9986fc768fb1648ba45b7e0998895666aeda6
za54cd0672374dcb10ae2b129e99a59cf8b03a2e56eba53c5f01e007052b1311f10e3d5826d0f22
zd1b2cd3e09329aaf7e485c1fee789ef8221374253f20da219023fae63bf147ef86635f0863f43e
z88a224f960e2202fa9749912f7775c44627c5b3c18c64822a737970c325c8f4e8be49ca821811b
z68f758a008b4e0672aea0e72826e7e20569ff118240cd2f4cab617d4354fe3f0d37b47f7585e57
z144a3597a73a457ef821f07b6037b560f1916726777db28298ed6d8d0903f1acbca174f405537e
zc19e00ced40680e01076577270240df8637b3a0d3227d7e2060b8746136aaefe9d3cf57f1cf1f3
zca2f5a0c9a2162d999d89fd5167c189ce2ad978a671388ef22c371d2c7bafcce2797dd4b3ccad2
za25e2e286940f40b232b4bddae5a90759666dfdbbc5047b7a6faca3211892547a2e8346e65f704
zeaf710f5cad525887a1ce4b77475ae2d62efba9bf97b94fa67ab7e58884f9f641386019171da53
zd4f3fb3cdfec60958482223ae0137ea2a46c11a29926df7d04cae6d4c7a695cdb1bb1372d50da5
z7927564c58d5cf82af91b529e8468c47af2c1554a1eec5137350750c42a40253b42f464448d5f4
z96b9a38d3667e30282a128aaff5f0a35c571a42f2079cdbcdd731e717e88e838536a68dcc820aa
z03aac702ac05c857fc6dbd90097607c0d1adc1369b44bd5bb83a7ab195bf83ec84c6bd77a18963
zf9046e33ed1272ab4d663fa241d6ce6702f930c520ac70e8071976f50731f480b4431cd2fd55cf
ze6d6ffd3d68a60e47d28de31df396802e530624f56b1cb6c61d813c7a1e70e5d02e8f49eb6ecbe
zee2cf2863eb3676fb4595d109be8b5d72f7c64547f46fa98a86293c8c824b2ed089108d1a2b99d
z7e9b9686baa39983185b11dc77fd6133ef4651e7ecf1807b1bc2be53d90b99dce7450c87acdf01
zb6192a3d8ab0d706e66447275ce5b5b7f24194254740f976643667db8c6819ecd382df002e69f9
z579ef3566a3650415187faaff5e4a943cc4bc8f6a4c5faeba3528c2fdc6da16ffabd44fe59f977
zbd7648e4bc77da8d79f03ccda0ce33c901b0c9bec4c5c1df8a03d405a225e70b75e6df950d3bc9
ze3625150b9ae438c6d34df44febdd92e340d3679b19246a285e0618f9ea45072128fe28d1f162a
zde0f8a80a9da150c7f8d6ca864dbfc9401420d8a13c6e6fbb3aad391d81dd27a4bc95912da0866
zd2ab3a3e624611e29236e4b2c5ab7d2b2db6b2064a7d2c4612e9a69407ce1829ac03e44556f8d2
zdfe70c2d715ffef3e221481fc2fe4616d2ea6a7fc2a2bc64abece241e4b45b17cd0d04c4a80ddf
za3a5df855a3c3caa46b78f6a2ee705b361b0e83cf5706f4780ae74b43041b9a759195906ef9b9f
zd319032c74b0cc06e4b92628f5908d7cdf00f943ae68ed95df6f5ffa44b16520c286afe2c7b131
z593783f4cb167c7543c23e713a322cc32271b5397486cc12ff2d5e40a6b5a82705c4d606f1b52e
zcd7b94e3e05611ca237a360d47182d284c3484f259813b918eb206410c4730be4dc7c0d2c32da1
zd944a5e044a873e2a1c436fbcd17345dc920530ee146d3277937ff2845c82ff1449744c92a09ac
z9c4cb80177e70f2f1263b26a94862cbe4b9f2c4733156f48e913612371aae88923d5f226e8f80d
z20f50bb963e55ad1d6c7cbd9a2d29217ed05e1bd74598d8ea4f8f5bed1ad8c3a9db277fbdad563
z49570545de2a5d834eb7d0943f6b2aa0f63e2a543f7ee568ee03afd735d21626dcbac423502b23
zc3da8df098264b85e3b0d93f3214b1dea958dbaf92c778a912cb53768a8f116db264573a2f10e7
z0e25482b67bae2281106427c7a8526e239ee2f39c58925947553d7bc5cc8bd5eacc8d17d246266
z81e12e528ad7ac898ac17ddc7a2e66cab95140a8dab453f3530be2636f438343d544f578057f30
z5d73e13a0274112772c48a4308766dc6d58e5705c76b09115487b42695b45edd961e87aebead24
zfaa283a8125887999953d4128bd76b667ac1f32e600ab766ce54cc10896a531ea5971b8abf6356
z8c87bf32b73de76bd082967964897d2379e1a13483985385ac7d2a7b00431953b25767f3a75f6e
zc78233e8a0852dfc9737b4568df32f6be4cc881a948a7374343923cdd6816a8dcb9d7d37c0cd90
z96b55e58185ecc3b8bdf44cb2eaa9a7a60fb0c1ab571759d5259e670553ba26acbf0dc59e71a12
z0195470856d627b84c1b3de80cfdd6504442d95b29bff7873d6a4b0729da0d1a1f871d79e53570
z0e6fdf20fc5ec81f3f4c1fdbc82934c3cb49e5f3ae7335cea547534fa3d37a89b442d8ecc01d23
z9751a8533e443b0221f810da3e957c44eb715f3349eb5cffa7bfea8b0a1645d7f35c439c848af5
z0fccb4f43655a95c2201acdb11d6cb1420658b8dffc8d6b237710a8631df3d8109ce63331b8632
z5869bf17ab3cf09e92ef11531c4d812c46785cdf9f4e77fbce7ab221c2698aa71ba77fa92ffe0e
z507e27f6476f0fedef9f6bb3e38334344226e89bbf2e7ede51400b8a829c9bd4adfeed6f3a33d5
z035ce0992070b6111cc0a13d5470020e06822c0e492519ca4a43ed221c56bc3592abf223f068bb
z56174cd715717d4ce7c15f0b8b7f5b7cbadced7a2d1ab3aefc2346de49d661f4322cad40e687e8
zc3fee01e12a398050678ecc9550cbd786e023d846992d26692ddd30079484d32fdce3d72847056
z84d7e40fc0e95089a4e73f7ffbc36d564c2089d2a9ce2ef44279ba492eb7c093464e2bc047b361
z1a2d773877c6bc33af35c68c3381f7e03c3209bd8250f911407f3323e5ccba85552f83666e3f6a
z9dd2334596e155bceafc67e4461a454c2db65addaf6ab92aba681dc1201c9583e92423af97889f
z8646b7fd158134c53749fb43ce0c091cdc03b51756ab67d268ef17ee086cd203a767e699699e02
z3a9d123f5f8c4c27d2a17d19f6e7f6723acb38dd660ff05d33f2e32ddf942b8903854767d80db8
z9bec94146b617861b5ca9977aabc1f06dced7d9fdc18087bbd5c21e8f4a82b714ab2a867a4663c
zce2161d7f3d700857c1ba56de966d6f01c82471b8456b0a29d4417e2f4295b1e0c021645342dbe
z74cdaa0531ed322d063dcdfce15a04222892aac37015ee551f9a2b5def76b965515675f1d7a9f5
z2669942b893c040c3cab291d2a19211f3cb1563b74cc0c266582457f5cd40bce8867beab400f26
z5a9442caac4184b209f2b219cf71e0eac6f4cac1c87e6dc0904ad0c9d825304083705671a22f87
z110de871f3b1578c291ca498a84c5cc03e1f6b552f3109501c4d86145d80c44ecf2ff2ecd02525
zfc8e22046fff3c4cbc87e94e982dd99d156fd6fc12870a1ac7320225c72019787e0f43ffb2b3d1
zcec4b6bb0c89ad0ff1a971957cda51374ba956709bbc668472356d31917036d791ed9e93ef9e3d
za73892a6426077dc1c44731d66135d35d85374989aceaff7371c015bc32038d22d669eb9114cc5
z5c453711f92ed71098ce742f869a2532112292e5374529a6fc1a506e5c52fd89e30c75a9ebb6d7
ze0054960faa4ad0de6202031181ba55230493b14e773fb04da92785d2c0f488d6c7823bb24c244
zf4068570c10cc4ee95a3e837f8549701d67afaad6aa1aec8a9e5bb47a03292de94417aa479449b
z762a7ec984db61b767a08f0a5e78d3358cd346f4ecccdc7b860468cf0eff1d18bd1969f895a158
z732ebf097365adce3ee5212e2d26e3a5997696323166fdad2005a907df02b1f62e889be7742180
z33e88f3b06427338208d2d44c518998eca53ddac13233b6f504fcd13ab4a45e3e6e25cf8a0e4e7
z2d8b0ea7f3fc8d6ce265414ba66b9adf63fcfc934f9215f0743692eb18228417212b9aff0b300d
z860c8c1578a27ff00377435f650898bcebd76838c4076b3d0346af0709f4a72ba29458cc043b75
z79dbef9e1c52665cb556cad17b1ba81002af1a036a9ea3105a76ffaa359c0b581434ccc1aa0a95
zdb15ed4f55e90338fef22345eaa65b7c4339c0e6c9fb673cb82a0c7da07e3d4a82493b8ae3c4b0
zbeff124bee3dd80cdb45ac6446ee92de1932ce59de2ab8b4550c1b5dd125e8c3e4ea32b5ba0a9c
zb092a420b1ba463cccf9050a8881f1da84ee8c4ff9ceb8814a11e085744b43ac7f4235a3d95518
z8fc7d3b07edb966ca320f57cd9c014af822b3a6b613e38fc78207e5f0bc298f73d0746e2b16ba6
zfd06cc47236deee5219b2633216ea24a541c4728d6cdcbcf6393a168e8287e1d2f51718ff67bf8
za6f1c0411366d173c907d795696f22338b4fe53e005d8327aea4c6f046191e1aa93c2680a83764
z7da03bf00ac034ef11f826d47005cf1d01b7cb5b98d42e9f64ac0924d66ed49a920e7db71c0e22
z8199fb1429c880f688f75a4e658cc25bd6f621010e0b701f0f5230606d579cfb5275ce8585b2d1
z2e64a2cb70e7c11a93901e006e1ae739006b4bb6c826d76a5b54016893bc11fc76d4d0bf3abd92
z612870231189592f3e7fa5ef0a26d0c999c5d53b4df5fd7c3d2a74d1c3ea05651541ff72047f10
z51b282e6092e5be22802fcb1c942ef9ee5055427cb2c74241f81b6546e8057b3bf4135d4b27243
z78addee9ab54e0c520e37a46afa16ec21dcdf583f7d3907d59a5e760b291fa7b8563b425f47ef9
z78975e156b2b4f6d3f6a051d581b7412c66a3cb44de9d618a5d779417de1de8756fd26d2d216e6
zbe7a893c6700d724f9cb67ad3bdac6764591f6189b0d9c6cc45779b98057a23d421527b82f4063
zbf60d90915b878ece42b1a797e5299d0c8685e799a14dd32e0f4b956448bd80f7cb89762ee3081
z4df7b9176307c780b744dffe5362cbff9953412b566312f339438aa1fa5b53f5df3e5a40ecc19a
za02636015f106ddb0cad8ef815976298d3f53827d2158728d189693a7502093c19356cccd375ba
zcda0d2e34b008b24e301eec0fa78cd279b3bb44fe1eee5bd50082b4ea60eb99bbec4a3ea5157d3
z81618b878fb284d7a6b9bb03c5bbf5dc3b06f4b7fb7b1a47e9e16ec7ae28978ab5086f2fada0c8
zbc4843f139df62971314fdbeccf470f3109e94051fc90b27468f665daa19f36d0716987d588e3d
z0fb58362e27878a248913d9dc977bd97feac2c2c17e645f93ed5649f8cfc0953cde755acde8b9d
za05a25eee8fd81aa304b4d0ac69395b4e72ee64c4455ff5b3f61007fca58c9bce8d6cc66fef274
z81cf0a1c6eab8d4565546e0355201761fe4e83a38204eeb85cfae5fa94a6dda22ca555b4a91c78
z632610037fc65013dda57cd84757cb8b368a7ca6523d30b219cb563fe241ea0ec7a7adfa30e113
ze8c2ec8da9e5053ac11a6d3600c39e55162defea275e74afd9d5d9d43b906f9a8952c406740421
z76318f129f315282b73d5c51456657f2b9ef70edcfb3bc0a2c603d39be8451553ba3e7aa26df85
zf98ee927ad2c8f3adf635db1f815b51de71eb40e8139af111df6f3aafdf2e167e50c73064b1bf6
z070a3b28d1e55936d6488292ab06215f6d7e173a4c550841ecc05f4790d9fd72e9ee4cdeb026bf
z8e28fe59a50ac0ad5e110fa97b577a9470dc82318bb7676409a7872ce6fdcd19c4fdb0e616ad82
ze80508f9e69efae57bfa05e3dadeb39632c3bc1f98039e7b938971ba106ca8f39779dcbf284ca5
ze5ecbb79e1efbea47c2cda45ce5ef29ed8e46e8693a24ecbb8a3ed2529e6ab1e678e97e8f44248
z50a7dfa93ad5637f32b64321a00efeb9280e6cf7b61cf226371e651bf66c07f5dc7c7018e5b49d
z00978432b87bcb3dd9ae3f24aaa2c3bb5b2931ec11305906674db1e71d304e04b1f31ac5b179b0
zd4914ba63249463e17d878442c0dfc409d5421a56b06e7e97d558d27322c1242b25e88f155e8ec
zf557c9a2d257d32e0507aeb20b2e143f825ae8d7557082037b5ced606155a66dc947ab86bf5927
z08e4f018683fe847f911d7e51ec6ed41c24d86c574dbaab54c63325e1c82eee7b287551b66ab91
z38317af83e7119fec1f1c2823933ed40db8a1de319c6d747a2f83fd8532d034cac0613dc6b23b4
zcb616127180c0bb6a517ae5fc46083130f1cdfb00cb57d2bd9c61fae77a7bf91ca5f26fb1de88b
z338746bebb6bf8e07e6b689fdfa0e38b58512841ed67785535c0f8abc7cd474f3d9094369beae8
zcf35faf18728f8c932a47ea42f85b5fecf9c4ae8da4217b85036c743a606cf9e876d95beb21f41
z59094dadfc90575125c4ce0ce075ffd7564bd3d82e172fb428208466803660ffa9b9635ccffed7
z30508825358316289024635784155062f0b4efaa612a4aca458a4ec9f75fc68760ef15c37c5fe9
zd216d851434fd9177683bf71bd34204332eb0c59af7fbb07fa68fc694acae324db4fbbd931ccda
z298e907f427716565401ce7ad1095022dfc451d313791a28b519619b781d0604acedb10c792e3d
za1afbcd13606125de1969e9b44d2625d6449610b80d770878a1bc99d04087ec3bda0beafcce7d1
z1ea8e70ac4da352af5269c7aa6cdfcbffab7dd361c80ae67b406200c4c2d723e475dfbb4c00711
z50935190b0c1e475cec212882013021d01df53d4deb1100b08022c9faf77997b3b4eab30dd468a
z3f42dc6752261f2416f68680ff76c705dc2de64b7004ae5654d54f3544c06efce45588f5bab89f
z84f19224d4fc4e86c9ce1f93bd4413ae1013330cb4214441e0292b332a4fd3e64d24041cfb120d
zbf29c4f7e07dcbe0ad055fa5a5993d7ca4f869fdbcc1aac916f6f156491cde4223bfdad9d7ec7f
za6d9f838ac45e8b4cdd7a93c104197e0488bc216d23cdd65deb497b3dca8225ad89dd61a466d0a
z1bc13c341b8d26576b41e2f5704746d1abcebf679ecb1fcc4cf690e77cfea5fd1baf880243fcc0
z671fdd49dfcefe1a10680757bb013ea98e443c0abcb4f3509c91655d1895302eca3616f18ca3a8
zae024f5f0b0c6511f5f59a8a0fd47b87ddc8dd00cf1559e1768f58d0f2a3d4ec4af500417d0e37
z1106249940800eea714cc1d00c210329064861636c89e851f9b40ca48e614969b48360ba8e74a4
zd365bc858482f4fca4aadf75c24fa4756b1c861823c193549a62b989950005bc0cb844e1489b9e
z71895767392ce570eaaebddb05e3aa2abe58bd055323b74900d7b98a4c80bf4fcd5c7af8522ac1
za61873296007306630af7e1fca8cb0845100364c80123d9a3bbf1aeb4f797d91c80b6d20360931
z5c0b2f806f2a15a200eb83f4e3f7417fe3b45c12926bd1bb835352e46f7ecdcfb70291c3021144
zbc1b87837f34e2bf511f42de0548ea6649c7172694d3155668c164b441668de9a9154467668b54
z6ca183a6334925d720b84f0d9b8b00ddaac43580dbbf474f646e93ed66fc4daf372eba79dd1e2d
z3d9e7aac801df7b60531777488504c87ba2da86e8e2d4d73acc10cc2948a981f2c5c283f08c47b
z67561998869a1a5915515627c435fbd5d178dc6d1d695c54c02c273abc8eaaeef6668a9a2cdf1d
z99973587c124c3052ce7b6acacb70f85134ac3c8c2d251c51292fc84e3b1916c95833285b7c2da
ze6e94f97ceb1ef43be861ad300e85859bfa561a38d08fceea28400b9904c2ff8f6016085a4071e
z7c21a06c3ababc4a2ab49593846a147e00d04603d2cba85be10132ee41ef8f16453f78837e76ae
z7f932e29301cf98269b81d9b1302a1606bf6d7ade714f17745c6f47986a0b5a43839b64978a008
zcfb1a687f4d460d83a4867dd5fff4d7f7ea0155037a4d25f506d53bf4afad2d58ca1f4f57111a2
zafc3e589e1d28ebc3bb559ffb6d2d10321fdb857540cccb1e26bc9edd0200742bdc6007b57cc52
z2ef0c190376565dd7a5bae38ae76effa057f17267e2a24d18957df43f87499897b73f5c9284155
zfe7765d99d97c5da4fb5d306913504e1ce2953fdf9ca88e244b698bbab03d8873cf3c0c96d8006
zd9abf518675b87d94250c646a4f1750464aeb32a55c3758213e8c166e999384681d59f5b2cf99a
zeb95e34d2ac6dbc0be8ad17735a955192f15f8f4348b3c13e7eacf6973d121373dfe3eb7beefc3
z9f84511d71452aaa60319a4d55290dfaba737367b64ed865be3492d75aaee736c5d1db2cc4d606
z2286e0b81a77bbf5a9da16dea73e9ece98d14151738b09a87780cc238c7ccdd0f21f4f50f751df
zd07919b6f9f9ee31d6dfe7bdb5b5c9e7ff83244d7b528b944623a530d8a2fee419654fa8501a05
z7e2b31a53404338c8b7b78975d33d295a1ed27c920829065f45150c1daa86b0a69e29cf07eedc3
z76721bbf5a2a1278670ae166675238517baa0a94265f8436368f779e54ee07f9cf3cbe825c03dc
z10c1f07e478fc2f9bd9dba8a8d105ae6436d807fe4be6746f0b05f368ad40f22dbb67829ab615e
z88360fb80bb5bd4fa5ed96d325c27abf1f052969bd56e866680296a458d7c089b958928e7315d5
zfd8d1291e7c509128dacdf1fbf6d9d43dfb79a3f4eb5b639d0a45e4c74927a782f79971eac7d87
z18e1d20e42ba0b79755714fbe0c3c10cccfd32a51d76c70a966802b6aed5212de74eb84f1cb3f2
zb4271ec9768a8d2214e6a75b43e4eb57fbfe72a9791913154a5316f76496835b4f6fab58c2a5c6
zc319175d576fab3955d9f6b0d20f836d2677a1fdce0837a498c10a478291c764949cb627b4be6b
z8ba1c93a7d99c5738bfc8c8dddfb81e55b5d314390e73f9fb72c1e00b069e956ef9d2306d5a8a4
zacea4315a557016010e1733fb723cab4d03751094fe2a7b937e2eb12509010e78e9c4c4321ea56
z8896a3d5ebe058f5300ba0eb294c5d1e77d2820b7b79f7be04093a204c5950b298a091f88885da
z609485ce3de575b5f9c0457cd43dfadfdda53b1417a1ad70389232557638ca81a33ea9c6d992be
zca280b6bdb0d19a8fc2c70ec3b8ccda78222cea18c9dca6880699078f4fdc22d1255e1665b1321
z6120f5fe3053595b74362d68bf9d35b13d609001b9b19c7e3f0d72e7ac0b65f204a854f22156d8
zfa61137f21ba7e83b5cfd97d65c41b162b8cbfeda2c040c744ae74459c167bd976069fc67bfa55
z44d08c44879d5e9a6eb835e0bca6a36bba44259d5ebc1638abc60ee9d4c1d2f18139332d9c4f22
zfba75cfee1e4137b6dc4c18a85962a1abcceacd315d41daafd47a81369ff45107a51906d9ae169
z27700856e890a2151f5eb679490031628c0d63546d15626c803b5b1b97df97b1b30a1f69f85698
z0d9796dbf606b8e27227dbbb18c370913aa6c5fa7f770795fabfb5ec0f5269817120a644d472bc
z04aacdf2762bd0de67092a2c3fb7cb063a7cb0300033f5baa7537aa2d66621eaed05a4e7adb3c9
z41fc72f8209aa34078be5a31dd118b6068ee5d9278659dcdee3cf2270556421efc52dacecbf334
z30ab6952582488d8b14147a0a0068fe661bcec14c2e8c9b736140d69091138c1e7b0ce24749152
z84918b25cd76e38e7988fff79fee80efefee064b4ed12d4f29abddbe98d4fc6a1a2953e7b79b2a
z73e5bf86eed0f70f1dd6502bee8966ace1b1cc4c1f2a2be0aad1bf0694e49d5f994fef907302b5
zec0d7c06633f140803fcb78ef1976a93af065835475cb5ce5fcc66805e7a0161e508eb0719f2b4
z70180dfe6ef7997dfe88d2c25ecf618d91b210eeb66935ca86b16ee236d90df204dc50d5598aa9
zff0343f4a99c90373b363ecd26e2f6dad01922edd3b9a3c1339478c402f61bd0459bb84e0da599
z8a91904a986ee61cee7b044169f1cc4817df8ebdff5c4bf0a98512a9498403916fd5140c154c25
zd2dda78b1346e6cc304aa4dfdd7e0a1b97e82e2cffda24bffa9acbde6a45ede17ee842d3af7751
z285cfd0c51432892f54aba6e08cbf49ba4b4a7fd301056dd902d84258adeaded01723ad6a0867b
z674180c8cbd59ad5aa8e9bc782f9579527329554db439597ed0c5007dda43c66e0e56aca5d3655
z53fa57afab9c33de3291616f6342087c4561d31de14ae452b09bbecfdf6dea1e83b024e403ade5
ze1fff7b8c83ec326805dbb46a2e68c59823b78ab9e80806386e81b2338c51fcbbf21876570d774
zb63d685fcb73a51c7da0304975780c9a9a92337b1e2e795c9af7fa41a980d316ca034530c7fb25
z3966186461fd5624144ee726745aaf098365e3c26291f242f4e1fa4d3016399b01bc089cc62087
z920d3485bbe35e1f8eb46693aefe8c3f22fd3279cf00d26e70cfef0275fdfcbbd1c2376c99d52f
zd72546103409c2fc8f193c343272589fef482c9312df8d0086f74eeb66c01f98a50b70c7ea9a98
zc50c4149501f635d5c6f1cc188d061d51639d8dd4c1584302d206e86d660cce23959e76288b9ae
z0f869861926e21b01e540c8b751fefcb333146fe60d718d28b8aac73345c4bc02e0bf421889234
z663a16903a3f16811599e380d36c17606acdec6f7c95bf1e73871eec79ecd26fcdceb59674c8b6
z53f944bf8334c8ce474c06c459455d850797dc7f73705b188dfadc9968c141765cc6c48d661e24
z0007f9ec4092a67a73fcdae9381edad7907fed3264382d35f8524221c3c0022d31ad4dd7eea813
z1d875e3a1def6a0a6741c454c9cdd73735f1c8158a771d0081f9bd10320c9953974b9e152e8630
z431f3ae397e0030d6aaa4c6f82db2db889dc6fe45754b293843eae0a1c6473b9539796639f5e20
zb4f7ae4b3b73b74d58cb4a2cf2d6498195f9feb2e992bd66a06371b4d6bbe826b5ffbb068ccda6
zea3385699a798ccde37f9cba5364b5b489ee5aea2b05635fdc79830e93bbaff078a29bb17af71f
z2e3bde165b128826b9e53c978f377ce2d4e16117607e553d888c5fe5d34ca147b907911f156eec
zca1982ed71ebd2889a87b316b3d027dd596af9abd9304420669e91e62a4599090fadc5b930fd3d
z21a347f9edb7702cac8578fdf1d4599a418ca9afa5f5560a343c6d0a4f506acd5293ee3bd67e9c
zc2744738765d430829c14bf64fd95c5e80289d3b48b42db37a6e0cb8705abb8041e53a7a4ca6c2
z75ec91cd323167a8f2febee8893b0b31d6b8bafdbc606f94dfefe3732f7f0f287102238736b1bf
z002ddfdc399fa4e07ba06466cdbf210eb198747528091c135ca255664fa3a8b0692bcc5d5e1c36
z57871afc22794751057d34156671427e81d5d22bfc54f7552d7aa5d179da987d814933fbdcff98
zd7a9e4a559d9e3d60d04088f45e61bbcb682c6b25a34788768aa0cbab2fb7c00264b770f5ef4e7
zdb7f43d846958d19b3fdedecd52160394404db119700059279f4901fab3fbf24044e5d5e3e6b10
zdbcd75007c1e2e3275edddd32c3f0be46c222bc0fd357cc2f2c0b14ad4e0bdc2849eadb07e3d46
za6fc54cc768cfd27b1f7e3abca9a0918031bf118bcff54bc0cbdc37b800d56307d31d07b243855
zc23670e7c929ad6cffb89cf50add5c1fe8a45364a7f5629a953f1f29fc4f4effbb882844596349
z158feb270dab604433f07a0702ea27b44dfb1945a9de14043dc57d44d4e1643a74433618c00719
z2fe3ad74111357cc0beda13b7caf9b0d55e65c3244784c3223639967a0dc84157b3d798e15994c
z590eb7729fefe305381b90bd1d0c69202ef44afb82e1f10141bb66757d609ffe69dbe1a1224247
zb2783a93a043531012846cf4ada253c054e10e587dbacbe0258c5d25bc5febf6178947dccbcb1e
zef0d348995fa5e51b60e5b2507c60b1e161e835027b873c0e0b75fb86ee1b02852f752ae0d62b2
z6e80a5a7398ce401d453b9afc3d2eed9bde1c788698da3573650160b3c63547b9d109013d23c65
zbcef96dfc1c8d628ba362b7d6c68b40735c810908206e4ac44fad2e6da566d2735955cf5bac3d5
zad623d28cd66dad378907c634e846abf63206ed867cae5e46e54fecaef9a6e2baca8ae0d08c279
zc9e1d500384dbc2664b0e9d5946a243b4af6bd80445f35d0b59466ac208298a4644ce4374cbe22
zc47d6e091847d827f29fc3194955a099c51eaad265730c8596205e75e4ffe88c774a1a8689c94d
z6def3f70c6a984845331f9cca37b1caf007b80ee21a549097beae55bdcea40ca91b19479af6e96
zaaa64e821496f6c967956e6bbdd9884a185141707be007ba31b2680277ff24bb77f9a446d28a87
z2b1ccdb4e627612e549677bfe8285c99077ed2b6f098d0dd2f08c81a1449730e2d68bd112771f1
z0bf3b18339730c4adcd47cbaa00673d305e626a1f0befeefe67c5a7a6d0a5a740997394e7a9271
zdd10a3faf9b5780b646c20ad83c81ef22bffe763a42f10a8af51158a396dea4e09b472cb71d86d
z07f11f78da88c1cebaa3efb746fe9ffe88be9a7e59b9d52e4a2734b6f933b7bdef47d1349c931f
z7ea8a4c207f1246f98698dae21afd137dbd068c3997ab8243ae91497b0f2e07312218f07178bac
z33ea63a5ffb9faffeccaf7d79e8f312b01033d13c7c20a045bc8531836c6b6b2a21c2a92100a07
zfb3bb7ce7c17fec3f1afc13829bb5b402a72190b556d81fbeb06dea41a32e47b954ac0c8e27fa3
z4150ef0a39e0c803c1f3047248b1ea0b47ee64d0d35970ef1237d910edc3b986ed8c474d5a8cd1
z686ad81ac0f260dcd025bbc5ba3955dacee0132b434d54d63a936dd8e6a1f3bc766e64bfa88caa
z3cfa07ac8253f11447e04b89262b81c0a4ff2fc3422bcda79426270f26bc1923a53fac030d951f
z732a573c20543701dd27195697ec474f2a65cf2e9efaf64a928df94f9838522c64b232482172c6
zb541a506086786ac52fca8e5d25253d08a0b872492b7e7fa78c67b201181f55aed43c45fef1908
z93506b51c3efbf94c9a2462bb58719576c19f1ac371f65614200fa326736501a3e09c5256344cd
za5f9e983384d9d61a8596ee5fc15f6eb01445bd0a0d413340a1675b3b88c6c88434e002ac7cb65
z9a47828de11c42a0e53aaf579847ee9cb9a3abf53bf4aafbcaba8e4cf609a35939e7e7af38d70d
zb49d84eed5193269b53dcf38071db50469401984528c5be1eabb910bd9a9e6f0248fb9dd673a79
zf00b37897961a8fede745b754907b3d230088d14acd27f1cb7e99935875cbfe3739154b8bbd13a
z316fc62d2f6a2bfb5284476df9ab389c4260cc45ebd59798e6862bf1062068c70d6ef10c462bf2
z3fab0fb7fe9a30861188f71ad77a080e64d037f7dd18240e1c71fd5c112a8dbd6db2072a786a0d
z3a29ce8988ecd264cc0cbad9f695844ba957e93d8ee6fba09590db59370e2b1b1aabf7f3a548ba
ze7094e7262b28fc285f8c8bfdbf43781cc7f1f876e5d5434491488f2df8dbbe6a3af675f7f4fe4
z95ee1093685ebb8d792e939de084a4445ce843b7f4e0ef008e25548d8f96e2b5c5a1a3d6538660
z5713a3fded5764adf2f1472995539c1dadfabd29ed76dfc4948e33c1d24ead26d9dc8248ae7722
ze69c059c5271589382550f35359215f900eb57b8ea932c5101b5f11caf6edf922a302840e7eddd
z35a9452deab8c24fd364afd68bd310466ab26fb5420ac840381c1e2f1f0efca278831e25abec85
z43d7df5fb55f5ff8786776147b37176f1891fc156ce5fe215cf2a09236f4d3109a325e85b1d7d4
z6ae7175ab1fe768269299a6a7c23309efcd8f7072c5f2359931622e39f6e99d7600da1c81c7535
z293d885f3d497167212b0931678764e9d4a5cf14ced91efa5da1dac6c4d47327c98afedfae9651
z3a4b19e3ca8ba86ac7ae51596feaadcd7cbf76349974efec716dabbc505479602ce1614ad9f27f
z90869903f45b782b6149a18129f29b8c03ec093bebfea651b8905e4fb1f6a01000ec354b2a93b5
z422b922e00cbb60a1d3de3b511fe4ad6d2e9206632c30cbb830865ace325a6a188244d5ac63ee9
ze56e3019351f0246656675b4b86cf7f1e6dad572192fbd1abbeb45280f5c65fd020c77db764e2c
zb0672cfe970547ea4b670f927cdf85dcc5b71a15f196e24f35b2d6c65c17944e7a7999a3008b21
zae59431cb0a2ca9d41732f5894a48289bd8ef1271f4464d546e2430e37e87e0f6e6bad37cc09c9
z5ba89410c8415475a6367aa28b125f9a47a50570d42dfc6585f29bfcdd803add4139d4e464262c
z988e4be7bc0e0155e1bf5af2f3d32b3506bea681f096c54f8ef6dde16f2456f1244dff755466af
z24b27eb4ef5c46f64fa486550a353728658f0646e956d7756c03638f13738825e6e95245f2de1d
z836e754195bfd1c8f545c5284e2a558c5e0f6c5ababea327944742ddcf52b386e69966ab833b1a
zfd8f937e33808331b0e856204517a5abb79f85f3773d826ae626ef7a5df849182aa0de205b27b0
zda7fea1bbe90e2ef32c08fbeeb8fbc3437b7c54b9e06e0d4150b497edadf9df37d3aa7ac59ca7d
z224a68e7b9216ad5587704d81cb7b030be804daa1481a183168c828e4e9a80b6dd295c475143b3
z37b64a6ff1cb6cdd25f928a9fb13173d4a243d6c602c361ca40fc32b8575c5269d116b7ae099d7
zc548d58a779d15072e7eea426a96fdadc9455c94b36086d53fc68a20f0f5b015e4df48e7d7ae87
z722e841cdd5f5f96a75d1cce53be4c7169f793efa52db37cee303069fbe81660149f078fd41ce9
z6db750198d57127221cd8f5da8a11b23fa3c0dd38a9b1ea7824ef8ddfae6af6dc9a2c320ddf84c
zb9e1bf52c4e6cde8b81e3be8154253e5a759ac46068870763892f7626f7beeaaf5ea577496a848
zf2b3c10876399bd239718a2c2729711591e99abf88e99494a501312e601177aff7ea0b9844b28d
z04ba9b88eda4461d08233250d363f9fad6aa2a1f4e5ad1fb15ea215dba39b1da0a2e1645d9e973
z7dfab71b8c27838410069dbebce4328df6518938ebbb124c9c25a29106859e02dae648b4eb74e8
z0cf625a2f52270fee685a9ac973d30a532816ccf0d5efd0cf93004350fdf00e0e2ac34d6035338
z92fe417e869e70eba096e8bce82c45de780b3f4077374e7ecf433970468c3533d3bd4ab252ea34
zdb12a3ba45723c0c6bdf2679329ae1a9cd35c81be75fa2723052fc14ecab6aeec30ecc4a43708b
z86813710459e6a8b90fc5e641f494e98af855d287e56c07767ae696263fd2d8746d0f0f987787a
z2caec0c35ac851460df1bee876cce223f1c3d0782e11d3db50b5dd4e0268a93440d939c0b1f727
ze6460caa6eedd12a62756974de495ad67e835d242d3584703b65a7f227969b656511bc4134f31d
zf26294cf7e452c08e77a555297db7e65b9b08c917b9e74d24ef78a0c2c452a15c1b18efe77b954
z0dbe85cebe515fccec26929fd329cff76463a16d96ccc386b99858b443ae02c9e069d06d560bf6
ze027c8b1fb0b0a1d417cf2c9d4aab2d60a5c8af687a11f4639519154060fd9e9ec4f363b78b078
zd80632ad1c5a75f55e2c99554d902bd0e90a9ec3f985817fd1c42be649b1db72a3da255350cd42
z8d1820b633f57e350b07ccfd9aaa6792e084afb12196dcf7fd9ff361226f09416c4b82d111528c
z8ab9c1bcc8ca760d58d286c1a4d7f331ab8c3d9d2b7e101a308b9be5f7583543a4b222c0be83c0
zf19ce5c5319cefec323eeed7c7efb6db77c897aec3a54343090bc2ed8a36a2bb48c9a8ddee26df
z5ebeb2e80f6824114aa241e2707b6a8969c045947595a1c17af00dad70ef4ad625439364de388c
z78dbd643012496df5e4a580bd6da29e82530c85d7c83851d6cabb180c71765b30e54755dabce34
zfd56e573aafb22282639e2bdfa458b0e47a3e3166ba9a0aa32069a2b9cbf7e85118f7991bf1aaa
zb0db3dfd20f16212da239c03f10a5b0c605240343ec2d667cbc5d1f90396b4f860cfc3afa05f70
z6669fb44121b8c0cffc230ffd6139ec8d6b2ad53d708e99b5cc9a5148741a48947b37cc7dd0021
zf42f8c3e97c97c8d6f2f7a9f0e10960d26dee736fe130def50d8113341f4d89b6b57a52ed0fe7c
zb97bbeed23a968497676233a5dfe1cd481b5b71a4fa996a23c588a42a773466502702f7899cd6b
zf4e83e15ee498f8774bbe0c8fce9460b50e5c20485144da435482f51504d757d68794573c21ca9
z9d675350e9360bd4ef83a5d2d6e788050dd7587ac80f7531ad8bf2f0cd8c4cd9bccc27af4bb725
z348665bbfa963846040bcdb441d86651855cd972a38efc624be8d78b56f699eb714809ec78dc81
z610c58e746b6f1a1677790c7c39c067e083e007afab40aae7826d4cd9df1df29e01094701a586c
z9c4695fb8ed444bbd69f92d21ca569648da44be8b0e9c4f52401050bfa793c2a8c0c1a73207b9c
z153b9d4c4f83dad8b191001f19b2bb3d9378c012e72d3a8eee7eeebebb9c08dbac4bd1af370327
z8a14b6ea79642a1a9569594172a700581b8c9029120ef272f5ae7f5cbb636caa06d12e5aad2afe
zb5ef223ff6e45dba3cb8a3f7836a95e7d368b530d23640573a25850cfd0ce6d182e03877a18cb7
z129c6fef6341839d99dba27db93d1d30c55841ce6eb98c0f187c25cd22aa915e22fa3f1d3dfa17
z6336f4d6f0047295a3e12d46a035201b71dffb7cfd88e0cd535f5fd8e7271f15d90203508147b6
z629f93bd5841d27550ceeaa7a3870af403788909ed36fc9d28139bc7837fd9a3f49d6bf302251a
zb9fade9250eecb4956ef8a48850e6d29e98e8b962f73f8bb00ff1787b282e69d5fca4557f27331
z8e3ca58991cd05596747dcf0276030293052aaee369582457d56ab1a30afb9895dc498ef21e67f
z6131e9853c9d774faadb725212bea6904cdca3871f388f8c1ac3f18ea335f9991cdce7408abf11
za5983129ed3f46bcdbdd03d357289de92ef8efeb4473f5aa0753483674bdc032a04a7527678442
z9fa14789e9e4e14f0364807bd014b9f37ed40c84c45eb5a19b7496f66616d2d93ca0399254152a
z8389b7fbf14871106259123984def9bc0e165b6bef753646f2b356fc2a62507457d51edaa0757f
z6795212e7b97b1c96b44c96cc2ff5f3cadd9284c7cc5be6ef1c3ede36b9c40a9f764295e6d6aed
z553e49b070f538924cb0dac942054d3463f142cfac18d08e7092ad93ff04cefc3f594bb2cdd34f
z49a534a31b51f30e01b62e2c42764f4a59e27b1e8c059e7287267947f8970877a5d85ace9ed774
zda752b17efbb10ad79f8d51431eedce96c4893c0d9e17c1c4ce1070ace81aafe5746fd65493207
z22834617bfff15017f475f0d983953eac1a2260d60655902747b3a2601786b7f2989ece214757d
za4433a496559a536a45c6bb7bed90f04a3f45ea379a007155bdaca8d13a1942693a487a8df276b
zd5c35cfb5e5c0714282d167aac130df0c90dbf64b288ea666665725da33a667d115adeffffe762
zc858df296698998838c01b5e6895310df809d381ec19a7022b899afd7e19ca0fd83756b2bfa80f
zaaf56cb30f351542b0e4f059216242e70999ed2c3838e2791b0261ab0670ed40ea4b8e78f953f4
zb6849106637fb82589e7eaea1d0b6dc90243267b6b6ffd9980db1223a276af2577f21693a33880
zb43ef1b1feb65ab38caec20952117b5ea873c897f904f0261f41780ef895646139ae60e9cb0b1b
z1775cb3651bbe9f61fff17a3b64399823e67c80bf84a8e52aee838d186d0eb6bc8d656314186f9
z65c8d1cb009c361fd0f9a6085a3574d6700141f643a9dc2f44fafa8598c1adbae7eb5e57e90250
zebb8ed5e0100a6469458ab2cd83c8554001b632ad177a2d85ff41793f3713c5478e65c841d88a3
z12b5c93bad7412b78dc83338ccb9e035d11d9812e1dba60df2ba8fef37b7369969f7bc4737079e
zf4bc892604d35f38d70e5b144a9ba00053ef27849876ca7e7d959d7e24e56d1ad76895f00ce0d8
z347ab6c640c7d265c978a15ecb4b63e160ca2aee8d3504d3030647299f19f3522780e88a2cb540
z8124eedbd5b91559e0280c175b583e5716ba23f7d0121271a2fc1074c7831efce5b6f227579af2
z634c303d9a47f4c9d67ae6179a6c7f001d676f5a643b442c9844431ca6d9597842bf1f463653b6
zb22bd9119d9ef47f82d05defe0e1e76427bd5dcbf344b13ad4e89aa62bf107125304995935be2e
z401d1366826d67ddf20fb76cbcf6d4757015a5e738ff56b9685dfdb40e1dfa05721ca6e1b8d922
zc254b8900c0c99240e11e97f6cf8e30155cecbf1db2a670bfb6e6e19e3bbdaa94563fdfa1cd48d
z9d2a763e84c2c3a9f288450427f598ce400b4625236e48a62f7a1cad33bffad2a12868e4724bd6
z527fd52427a6cc6a85aa5ba1e131d0a581794d0c83dcbf0f7fa26c15e3cfaaa58b8bd1d85274d5
zced1447be6c05004b2d809479c9d8b7b9bc7fd813b31154dbdbfd6fe2f17298afb5911fe466368
z8b7b942449f581a4c45a20b8a91decafe79ba7f88424019057127f6c23fc6a197ac28b3ac82f8e
za157b47e8feebb2ae493fa5b69d29f7c365eebcf77d2985d6b30f7084026dfd85f04edd54cd9d4
zfe54ce12a0b06ad1189053c87e6192e6e2e4443b3584ec5f4f07eb685eca0662584feb0a2e22d4
zd8d56a2043cb69673524d712c159129040642a5a37e78306e50bc0e9bd9f2e2be7bf33e09c5cb2
za9513fc92888eaa6a07ea6274aca3a30f7ce3e91dba2a3e02423c51c37ca70c221cf2f2f62b0bb
zb0054a8803f4bf845fda48f043f330eee021784527cf6109e9c2d5ab163947eff20e21e748d1ad
z44a491188532eb0469686b54fb393899293620ffec51cf61241d0ae782ca7935bb54283de7b259
zbe7c77dd7b69f32d0f572c0d05edfa9c6733de36b3af1a7b2339d1b867bcb00f29b46a06b4d2a2
z7bd1fb39a134109805d95a7658c342e4d7457612df0ea6ce0f5b3678bd87bebb20f332113b4a47
z1dc10b647c977e79c7146d03f7ba11238ee2db3960a47618383ce3355e2192c6829129e479b87b
z8b205af64e893454f7e4d5249f48cce8c86cdabf890d4ee926d5d773c1f54a619c527a14676b07
zeeb9cb3119311ebe0f16aefe523ceebb9d6f70de78107c411cf9577ac9c753fa267d309a202575
zda4473a35f27730e1e6d361c2b7a0b9352178883b9ad66c0ff75d12c5fe0d2ab381f508a29d3f2
z60ba7ab0265dfd7b001921e3a2ba8379895e46ba4fa92a349d9bb1ac0d6b72ba9793c21032e973
z02ba15cf5e03fcbb9ed424f7619698a7b5c9c4c7e8d736a93950cc40057760098da790a122cf3f
z32fdd9c47316a447263667e9d687092d40405f97bff93bf74db42655dfe52f3bc9dc9d1791ad1f
z5a7ab9f0e4b5e923d285a18cde6363a8b29016818a9b6c29ac861fcf89bd117d0ea745911c1e24
ze47091a1e1c03323a95c0fad4f4f93662b2a208cfedafa08ea1f7b8640e735f04832be22fc4601
z08eac948f3f1bb50d81f8267f7166e9116621d5ff12e5873be57e647f8fec8e0c9256c939118de
ze56bab896c5b016bb1008ca00ea5df92ae9ba5ffcade9ed64626a2afb6ed6e7bf4d54e78d3cce2
z83056e647742f9cb7feca48f5513d6b86ce60dd78a15af6759273d2dfaf987c0c622208f3ee797
z7bb9f74fd788891ca8e5530c15804acdeebda8fc9533013f65fa75e153f55285d0266f48bd91f1
z0e4dbb1acb8f8bcce12eb6f5550c05bcf5ed77efcb812f30cd8328b25deacc1b7d33a2c3f98753
z12f703941a93eaa9616762fb12b1dd41dd8ecafe77ea730533124f2f4d13368e9b6df19ea2a89f
z9eb2c4fa39c34216f9924b0a977c835634695fdae413d36f32deb9c3b8789f9c81dcd1a03ca1e6
z6263333579d718c3d32e793172482e46865983848a38d71f23fa5ee7a44461d31a2c761e3c6e68
z17526d81bae909af35396eb3432a6c4bf61c62bd29fd807beb149d732577ec484c61c1a3b4d01b
zb213bb58bfb3487310114b903b46d994fb8afad2f6e14b0b1327bc4a64d19bfa8a3c4049de1e9c
z94ef2aeac6a5d213638e98399b35fc45a392d0acf202829a172c7433849a2617801d1938f5fd9a
zc2031f816c9bee1a40984167546d91e757b886411e626a4c07b5739be44e247ea522f7ebf95310
zb23a958a4157d9cc0b6968f0878c3aca826046df833f57db1798fb85b654362c27efe822bea92c
z3d0d11efa9df2772e593e14d3563fa47c5b618d14a4e095146b2621b4c01777045a96b32c7a9d5
z1a4384aa2309e965a0428a8253006b10df0edd922500716129ad578d9c07da06ac6ae496ff2696
zf02d9bf05728790df7f54cac9dd27afed89446c100f489b9deaa622219c3213ad901a6312953f7
za8d95947fb9c6716518fbb2abefda8cca3d25804a90a175f1841067edd433cd2d5b31cd2161e94
z4ebc7f903a0f1ba01acf776ae1ddb286744942aacb36bf76a3aa4ecdf92c60332910c4970995a0
z6dfccbf997ee2751a26fffa82f743fa30c0002459a2383e5394a7d850eb51eb09c53bcd2abac28
z27dd102f52472e70f2bd21a7a6b561ab41c5bb6a9d36724ef79bb5fd1e20908985c8a6895657f7
z50dcd4f1117efe17b642756363c78d54b57d67f651f4503e657b2d49c69faf464ec83b8f44177d
z99c665584de24e06c974805fd740e8b1a260237694982978b87052e5ed906416debdca31020847
z7972a465ff7433f8eac3e8f12419db50da3e96b0da1073c8629cae5423d587821c41b51a553d9a
z04cc805047985a54199626f9a1b7cd1490b3abfc66ef230ef573582cfa44827561b296c584eb7a
ze3a41b54552f226f291210cefa6f2cc5cc1e7922b72c9e851e97d4bc4f94bd157c5ace04ab6a03
zcdcb14967ae4d3cde78c6b1f5f0f751a79f67bc8509f4ddb4e5c5754615c04a02095e2be6ab94d
zb48e8b45a6130e2c544118c05504a19187c2c50efedeb876db362cafb3e60edc9ec37f3a990b19
z31ab467227de5a43e21e4fe96fbe0b56d8aefe65fc2f3b591c0a4c746332b88d35f43b818c7382
z2d0d0c0e2c32bbe6776abc804cd32c758a117cef139784e39349d676801d70a2492af2dc00e426
z66df736c6a019a08373ebd3ef42599d94c21f99aba78f38a0a4a6e76c86afbb3e612066544c9be
zdf6aad6556933f1a4696c226bd8a08446bd1bc10bea9d34f94168bcf26d9a828a002b5c2f23608
zb992f21ce9414cdb60a562f0161a97a4a213049e73ee8f00ff88a154058d48e2f39952bfccc630
z1aee4e53c83140b646bba3c14dde1b1b42a17a765ffffe8155c99f75053a42c096d6852ca84273
z7485fdda6c0bca2a5108b3f88d5ef3a8778a89a45270940ce736d09de847e6d85628e63b16762f
za96343b44e54dfbcc13adda55a67f5f6b62683a5437fb81e151b3abe4094c9260966ce572bbe23
z3a4eec6f111ccf807f86a47db5b48d7381522e1a78bbba76e39336eb450a45a38d5c4961c05c6e
z31f4a03d98b8bbc32ca888ab1f6ed251114328d57d2d4b82103fdcfd9583fc86fb0ee2587adee1
zcf2e0f083ac1af21dd69babb6527ee4efc5a8c3298153022b411e4eb2993e8f1fdc59ce504c30e
zeeb38c421c1a0a6f137a301df8c964f45e61d5cc1cda3d22f04f21acab5719b1410279250e2607
z48e5801c1836e6c589f389781a30860b609bfe47e7d7845b3410d747849345d53d86f7a9603005
z4ce07f58ca051d87c29e590599df06ddb5e8498610caeb7d300d17f3ded621180bcf0d661178fc
z85e14d9b653045dba707f2d8906f5f22db3ab01d037f8a5d4448d1ead11f08a82e4706f2927305
z60bccd678a2154bb1feffaf93d88f9e5c955a4ed7a5f232d9e8e216acb7480b829e9364ec31205
zd3fe94469509429d4d177eef7948ba455c2aaf243da2d30bee1c1039a02cce7cf35a5637d685af
za13b67fc00a0d5bb27d293cd60106b10b5857ca2ce113bf36a3620d468c5dd073558691e94fb27
z4e3aa3c7a4aa8945e1457eb87b0aadd3ee31efced93bc14b501a2b0cd087c79e08fd084a22205b
z18233efc6c0a347b7508516f75609bf5caa10790a3461acd8f4b4a68d8d8e5fd2175226675d9e9
z4e3b9ebadb84f761d6922529939c122662c5df3981c884807c23dab1f7af13d38b9f91fe00d508
z5914e28fa231ac4df2143c2c3910697cbb9979879bcaf96744c537726badd679f08ab3a54a75c1
z4886550f576178fccef7b747282403ef7dec255d89cc14b2534ff082296e8f51641d5ba014c668
z32c19b197b7ec18087b95e00fc20749dd8a024e4ee6771db208cb72ae580492a9067ec20aebd14
za03d8a1e6e02a7e0893365e49dad24429fcb1654d1de7ea138ebd2a9f5fe4ecc3d7749f0632de6
zd20ab90f7d90b1d0805279396a55908744fd0f364514b227f9acde090404fc6a450ad41c6cb6e0
z48cd7d112f7416003a300274e2787333ceb410b0e9aa62694d8c0e7b3d7118ace3ccd59cb682d7
zd1a41f407e390b9fc8b57f19267db7b38ecaab38025d2dfb37b2522fce6ce4acdc1e63167452ed
zca7942b6207db4e8d3fa93ca7e5ff36f6fdd1a1bfb54ef2503c385e96e5d0a420ac69c21dc5725
z45aaf7e8e4242e29bb056ff7445d1a65482c9f9fc44872b144387ea183e7c4654fa2de2f9f654a
z31db15da8a17211e7a592e52831f5fafca03f1b60a8a9f405edb27a106e23a9fbd12461e384b3c
za2f92ff4a562d81e0c731a0f511a47411cdef3b753ccf08de217c7935fb6e7a26c2810b90765a7
z18e3ffdd30d9e0c861e46448738814069b2b991bc922e1ceb4e411ad710cb05700f40379ce56e9
z132d3f36c81672f2eae5ae9593a8f256d11836d6a4bf7b1a7babd4609233035894300b04f9d537
z5efc1f601a5bf8bedb50dbc920b8c4010d26e011f06988807476d85c77d3d40b766d7b8295b05f
z714db340c5cf79a93a5ed6a9e4200318e94a5b19f08605ecebf64552290ccf6979090c2a3a7947
zd0abbacd488e02eb3627b39b9378620985eb0f0a2d180b8b2f83c0deaa7098d8ec89e2b1fa9f7f
z6b6c4f10acf4941b3d23d7ad13b3c30b90634b04c5c155f80b10d0d39592dbc2b835d7198c92e8
z97d32a36e95d25307039079ec11cad29c88c17e7aa72135a061401b50d7f4558d38434a1c77458
za23530d01ef08b1dfab433251c338f77a6b70ee9ee7924e5bce7aff4a54dd564686768da5bd3bb
z0a1901e54567ce706ec6c322fb881c148a1890ce5909f5c00a7db10395379dd45a02443312e30b
z45ab51a68a86a8060d61b4b4f4fa2ddb69a00ce7873d5384e7c6d19d6cef883ed47e2239b83201
z2b48d1e6850f13a2d8f23b92bb9485172dd85f3b40a9b7dace3578de12ba6ea8c451b48e9cc7cc
zf19e5776fbff09091f31b89811b362bdd63bcf548054b5a4c7aa9e5f0cfb8ede3c1d6d01c057cf
ze079dec2adc9e09f1f759d7bd3d5d685e4f989e993ecfc5629601fb46309fa15d750c5926dc957
z122f42bc92e46f83a62eb11d1a304c17ee1ea49865a5da257fb4500a0de56577364924c64eb036
z604ea983c9f79a0bf96e7fe3273184d510d8e06d729c292109ebaa5cd645f77c609fa5234e3e27
z48eb290bda1252f659a176d82e6198253385ac768b06b882fa2dfdf4dedcea19e58701de1cf1ed
z26947788984f254621cddca4bf58db8979082354f38eb3fd5e438abda6099e9f3110ff86bd5adf
zb78ed11837e6096a2a7fce6c9b23718f4971905f97c564e3465b5fd930ea984aa359a872ef91b5
z130fb34b930aa488dd01c0ed36d44cece3d7b95f9942343b6cc4e705d8b07124d2e52847b63688
z5ea271afee332eb54e2babc1fee4f7770606570b21cb62eaebfdb7fef3db1a28de3fdbab8139a5
z0ddb2a517c4a72c871a9b540b8dbb915f0ede0b6e864aaba53fbbd9ddf3bb0705a2079349a1539
zd51df828d80f9c38edf5aac823af2e7598fa06ffcb6a5429fcafa53693b5519a6acb07842998f4
z9e12955b4a55b259d0202279c42fd16785cbfee2b857edb75d4e22a696b2877a69e026fd2da696
z3f7a5573873fd83318039ef5eca75bd323837fad974be0f2554176051b4e67c414770c5dcc93b6
z567af1c2eed0edf8cb1144d0465aa5025acb3285a670c1ee9c069056ea49e2954b57ffcee2e9bb
z6305af4092005ef90e3e2f5e3c2c84caad27207ef612bbe176d58a386d952f85c4032a3aeaa35f
z17304c6e30518b703462654b81b77be12cb43270c566f002c3d0d396292e771fdefbacf346aea1
ze89127d2c705d8100034bb42d33aa8db23be74786b16c819314fa5a3d7cd506c64b5c3caa4c6e8
z9659c51547722abe9ad3a50cc92278f452d6544abdf089af686197373965600579fbe78fd1c322
z9ed1ebd561f9d011e1650c0e109d1bde2f2ce6ea1468f0c54a084a2ed2e4690575ec087717b044
z1eb5ec46480cdc9926d90282534996095a960822a8e1f27fc114e4905ab6079157f5514d64ff8d
z8a5d9506a4c90fbf3a24a6a082d4a74d5885b308323c2ed7f6cf5c7aabc9d0353faa363d1b58a9
z01fad5c9f15152f55adf762f5753a2ee5b03a286f6691d713904d27e57ee2a71422e4354320d37
z1cb4a3977cf9ad84de05a2797da7fcbb4cf8681c709b5dfc5247b85840a5c792333323654012dc
z3c4f7194e0cdc81e0749d24c045afcf41f0a930f2c8e028d3d4893669b8b16700c3a5d4ece2b69
zf6cd6bc4de0bf6ade42e65d1583128fc2ea7fbdddd2eaee5dd05ea47430ed432df92f2afd7c01d
z1cbb5902a0ca4bd1eddb284105d963228be9e4556eed0e060e1771873cbc2d755a00b042744579
z0d62ce6c0f4031109e6ffd844088acc8c7439eb69b8ec1bd3e12c7cd0fc30a14968176aa84c73a
z1d4087e24643da0b840b0978220d2de6bd32ec2dce498bf66d8faf852d6782f68f21604dc5f9b6
z4aac71f320c3402b31d69f9bfd416eb11d0af7c10a7255b580971fa23387670e10ed5b9ad786b9
z16d5c39928a0d37aac013acda252c654db661ed3c86a4ef74ceda5447add1029ae9b52641f962f
z9f1def19e81f4d029b0cb72638465b30bccbe3056e4f60e7198efc3603ea0c7c22278a50312c05
ze63094c7d47ea57c3ce40a19bb70635c2b61bf959fdcf5eb50b02870e4f0bd3dfdf10b02348c92
z055cce580cbde43b7f7117aa89ad8aaa6e77df2f7266d85e51255e1c5f235d9b519506467f2df7
zefa018edda53d9c487c93fad25203dd5e6e2328efdcb5f3c73c1d7b95a2be8b8c77f20f27a588c
zce6ad96836d479006c43b148252de9ae5bf1351719010a67ef453bc5fcecccc68f765b471579b5
z92e6d86754b3dbaf4ddc75f1324be5585843df93344d97418c51830562f7744015bed2cfd61900
z9e3f125892d2b3d7c5ff7788a27829586df7f5a227f4b459e726e4acf253ad66987d3896a70987
z72f28733cbdf537e6736e47c6540f0e76de161d2e57bd862f809e67cf70655439e40b5093283f6
zf92e0047b212943b1d36551cbc2f17cfa68209474611017f05499e45814e54e27ecdbbe0098aa3
z5c1f6d123d1e4832a11dc5d2044a1fd6f6698e01b379326843dd1735de985718149bc3b0ebcaa0
z2705cfb674ebb16f1e693974ff788b8b27b6359d07ed751756041a43689b2abdfe5262225fab6a
z4d6ae02299e92e46a293f42938413890d17bfa047c3710bdfe96af3767361dae31567e4df365ce
z50b269e6222a0e74bee1a70e526666dc0bbbb094ea73f717bca1e5bb957a0654a68564c3edb283
zdc5ebe496ecd2481658bb35cd9142396d8375e52a387f9585aaaa0b47dc6ec0ea9e3be3a829ed1
z7ba1abf67b94f89f358197769b02e17c421adf98adb8bace56acbc72adad9dbfb2bedd04a3114b
z70ba806c9ccd7be24134ac66946b135f75af37ef169dd29bce9ed5affa84e00219b7411ec0a93d
z74e570bf40a7172a777f3814d6b07a3119dc0b90134b13635c9ba8b2cc75fd7d480e8735db3566
z89350fec040abf644ab74def226c155d21c129aae381c6248e3557c7dbdaf56f62db513d8c2fc4
z95f97fd01aa130f5cd33556938d6d0193e7b28dcd35725feab4ccb49033a3b685f7f78b1edc90f
zf470a1331be1a100a89c462566b79dd991caa21a4507aa69f45180a87973e9c8973b63b8946ad2
zeade2fc7520ada98734169add11c7edead631b9c7d4f0004d91e0d6b8006b6a3652fc323d2d927
z91c947865013dabecb19277e5ff53472c9fa50d72ac906872cb041adbccb0807b51e19b2f48642
z76145300d583b59f3e6e5b663ed96cf1b602e59f11534c9acaa7f3c811c32eb31805d15961b8de
zf87860683c5620ca66fc41662cb6d66702bfb3f9e9fbe350434739d578ccef64b55f315e7dcb02
z8e7eb1806c37e752aa92ad164ba5501c2a232a7fda7d1746dbcc982187679ece7db9e6ab340fa3
z0ccd89457cbdc54104b7fadec02a0b2cc903be902f34fcf0074c902b4c4c596fe7e3588fb8dd85
z8aea6a1bb6e4465175a6c1ca5ee7c311e4051b13c5b501938a2e9d145278b4937f15ee096e8d9e
zbdf4e8ff93714ffa584366d0fb3eed72a243bb928b065f13fa292a151f2c4a0f02b15d83ed9d02
z5d0c332b71e7425bfe3980ff05dfc30ae9bf70c5c31fe9bd1bdb82d8b0bb7b1967be7fad31cb07
za6ec5df8148874a3148dd85a5feb80fad04a6c0ef63117a98a2e22132e27c9fda472be3e515e98
ze173a1d14a907cfb58623710ed7b7b7255244b455eac8901d4134c1e5b4596a392c07dfd505ffa
z1859b1761dd918d455ddad097e00c07fa97a83780c5bd99e9ea4e03a6ca353cbaaa5e91fcc0f7d
zaa0b54dae588b46ff2b77e39413b07f961a955e41662ad588ebf1d4bf3516f196f2e8ab5149f98
z41c58b8dc1adacfb7d13c1552a1d8dd59549f3df53ae69a88199c6a1e3a79213ccdf3f59fd83b5
zc0dd76502d622145039e451142293531d8ec48b28fb99a5258cda8305ab4beb48088d4950d6663
z404a98169250d1bc7c0492abd8cd7d8336b9e15c3dec9ba5d47e5136d668b88e54a0be22907a9c
z7e55b1f82874bce195f220448aa04605e0758239d7d95f92819cd902d17bb5081e4a998b6ad8c1
z35b732c05d78502aef4424f0cbee2949639fa583fd2d3b29486fc964d4f7bd5fa52a28e9a6f1c7
z9128ef2b863a545afb1148927a1b129419c1e3ee5f6eb7a731a5f19cca874dd4122321f573f495
z27ccba6f7a13b9a9cae5c7edaf2ed2acc2a2cf4f3de640de255224a98c310c291729bb720f7794
z0d478dbbb7b2c30b8b3eec439dbbb8bcd401e1f4a2a68a75ac0f2b6da3e6d98ab044de30178a88
z88bd179f535fcbdd6b4b1d4095e78864e43e604b96f449ffc004471a01fdf5494dcaf39a0b3297
z5c34049fdeb954771e2dba94663adfd03961d726e6235d3c0685181ea5519377ca9f89de95c74e
zae5eaf459104ee34de9ec385fe7fec2988bc7b46aec926a5477794be78726281254d8619f25a6f
z378226186107136e2357eeb57ab9729d3f7e9b3fd0c448d70a6a535b60763f265e78e65cd3d7c1
z4906d74dfd8e5ff474c1327f2d86acd2a0d7b50bc41d3803ca61303c1fb945ffe4ddc77cf7716b
z7e7eb9ec3ffc3b0da1965b5d4a645dd5b902ec25469146a0722e038d3add6b6c72c0085f36b104
zf3331f95ff8cca5db23c7fbcf7092af2bee45e2b3c64b795eada4faa0ace47e76f69f49d44e369
zcdfa4028a198b99f65cd64b11a01f626b4aca4b91a8bf18c1439c4dadf96219f70606522114c34
za366b8dee8ed9fed9f8a242da4767d3ba36fff807297cc46f25644e760d9f501f93b5e2acaefc7
z815ea7b8c407fd722718580e971bb67e8125fa887673253e509174f8a056e0509edf9be5c1ae9a
zf1df4246e2fd27281715559c44091daad53eec274a2fbecfedb681ae2eb5e7624a4ffd2a92ab58
z349ff4aa44575289d301815fd7af3686ff6c5b931649ee5fe34a703209952bfb3ed6d4a8a3c812
z535249a50459933ba636d2e52db1979af7f3e470ee969d9154bd04800f975a1acee349adb7f7af
zca5fdbd7c4b47bb9e9556097b39b71174c2df76b9cbe4c16ab0d475da9acefa7aba89fcb904a86
z60be1164dc3f8217a5ed0d113cde4956bd1743ba951e6f9396bc1cda28fcada4827cdbab3c45be
z37400784ab1fcaca755565da3b60fee2f8db0f868ae8cafb307e63901c42c727900cd140a178f7
z716421a51e2ef10ef651d5d18220a60b3386ca7c49e986736ab360954963a2d246aee4e45b3154
z72cbfc59a2331ba2a16030739d74015aa09a7072e2067bff8d644966ca3d6c522ef7f9b551e2a0
z43d953424674052151fe2568a8075d2333359fb091327ed0c2e0406bdddec5d008f795abbd0bc5
zea2e59fa9856dc3fa825ae424faa8d7c2d2111422bb71e26047ba9ca104c501bf01166cd30be31
z0b017b7c1c2b0640f6b621afdf385892663d0489bbb142891f07511603aff6c4c91a1136f8add0
z3aaee0cac73f94ebdc4f2c2d328d8cc33040da64c852992aed6b09d05a54f5560a36b4373440e6
zbaa1b84314c42a2aecdc114a5619631c9fdfaea04358128e66db1bc71f5044a99b7700a44084fe
zef57776237383c17ca6c188af5c282041273324c16e7234418480132404104d2c88a9b802c9f0e
za47f595699bf006f119d792bb5dad8022e74dc6db05bc7c011227524ea666de69378e4421af61f
z0230474c506d5d4fbc05d1ec5e25c54f15f20766848a261fa621fd769038f7ad88e7fe0fa75a10
z46b6dbe6234da28fe42ee1ec60f4d8265f91ba70fc181ca1fe19aeabd8f446a5ffd1c6019f24f7
z31a0727fc900a2a929a4d4e0169b89410b611ec35416c6307c73be1e73c5b8a5a050e5add85ac7
zfabc6c6f4d4eb6dcd6078745b73dec37ea4fb913e78a1cd29d2390a68c5e751648660eb742a86b
z645ba0b80ea3faf3b0a5b17b4d0a7520acfcc0f3fc90aa1e1c85d55c82585c297c99354294cfb1
z6d7da0e547b49946cb89ea6564663fed139a2dcaa66a5d0bd01552eea50734eb0dbeddbca69079
zfb3310786fcacda5df806dd28bad56275740231cf1758b60ddf4e4bc17cbbdff1f18b8dd61e4e3
z5d916f2dcb25ebc0d2048abb56fb861d06c015467f9eaea2fae050cbd739222ceed4f412caf04f
z8c20cd8be43706c9f459db620fa2c33e13bc39cdc952bc0c90877b22c8b04ae567ea8ef683a4fb
za7952b7d43679615903447bb74e6ffe07da6b57173284e7c8f73547f3d912e832af87166faba08
zabb6c0fb531f47325db631f2532a195ca15c43088801e191d8a9f9d527b7a84f793a0cdb1dcbd8
zcfa68c1f1c07407c30898d57dbedd461180fe1640224e61dd7f2febd5e1e542eeb420290f0df02
za84e0e6d8cc3b027b7b79672e671d59076d4c19d0351b074560cd01d11716e29ef74fa197ca162
z6ab080020d69eec2bc18f195b9c2117b9ca7c1dcd634eec2f0978dea23aa5885e4b8828046d5d4
z46fe683410f8b388d70fc224c7316c499c601ddbf65f25a5e2c7117843acf98387f14081d5f31e
z47d48d60c264fd663bfc61d2a211c8657786223628c926883de1682446c9d8fc7aac6853233b94
z6f4f4f8b645ecc3d3fd696bacd14a39d3bb2463701bf985cd82ebdc1edb7606b55ba1ea4f61aa9
z6e2008af9c281bbf557ed6248051ceb074263cb1df9ca5ce5ca4fdcee1998d26359f6475c022fb
zf6f34ac5551f63330ea51e72cb668d088425a407a6ee3f62a7e70795fd100ff94ae2def385de19
z9532f4d0f72036dc3e34cb5513d1b59ac01443acf4a3adb619fbd16760d7055b43101daa390067
z228304517dd2c112cf63ee447bc0bb2d7426ffa88f24c054bd946960e992e5e41335130fd9b652
zedde0e0ddddc6e0d3d418d299a34a807c45cc87e585edd95324761c8e5bdbb26c5565f31323ad5
z935e3bef28c0cd134cee6ec219bd4079fc2304a13c94abe664548d06d8169aa4a561d1ada8d787
zde43f65ca2e916fd0b9c7bce743ed6d9efdcab4ee6f3179bc0431eb62c68965a4a27e185f1e4b9
z3f0765886b3cfc36b218edacebc0963340fde7728996ddc72bc8ec50194efd1138e21f62b00fa6
ze3e0b23876d308ca1fdc43dcdb62f6499803225a2f55ad0ce8018fa505608e54e253648991ac1d
z86d8e86be2ce61226e0af6caf9e0ae441950d5dcb3b659f23ce961d2f147dec04ee5c597918248
zdb52c0f088458b95f99c4550f4e22c50764ed5bc1d142b56722262df620893a2008366e8d055aa
zca7b3c144552d01fe35eab8eec8554447179e457415ec0c840b5bcf567f89e8c9002d515415e90
z1f3ce0fe178ac445fa987f64f0b29259986499ff86032b691ec12fb9cdf64e7b4da660e65832ff
z0ccdb06a33cf1ff0d1dc7562c56629c3c3a4ef1f5d874e16522c0863403d83be9a3a6d88bbc05c
z59400f88c6229bdc9e0f276b07d4610472c76fbe31c8c89638e1a0cf5852c49f695516686301c1
z3033f9a3db5e1b0b54f5b2cecb62a63d10946ed5327179d09df352d3be3db17414f85f643a1da5
z6f9989e5d47738efb1a80e01fe484843c21ff224f094da2b6fdd81c7914dace66bb8687edc80dc
zc3858e5056ccea818a0e41e8d622b50d39648b1f632189b84eff018df2f745a19777fb5aa36c09
ze87f347e3ae8931999f5c49753a586b5c5d92a88f0e7cf3badd43effe32c1162328bfc39c60d6b
z0221367663d2684369522b82fdc570888bad19a0eece71091e6533efb53b1481d73081fd210884
z6ca2bee01e1db36ca9632d617d189b557956d6bad1bf94c05b08f36b49a46d3f4ca0040e1982f6
zdd884cce6636b0975b7d74685a3bac7be84e338707d93ccb2221ef87fca4faa8a3198938d5139c
z62f7b65b62771108d47e8ec1f560cc21e3f9ee44768f75a81f1e0a70cf6b2cd006fa48d0b5b57f
zef8a184743ed543d8a1e61febc5a0f37a02356a4358a296dae11c33950dd351ecb7bc07a18c7a6
z27e4c3eb9e47d95e829815abe189a201d272cc433bb366256917fd29448fb442d0e132fd4515d0
zd7cc42f2f9582615a49f678b0f313be6c8d20e53fad967f70d966ccacff60519aaf3048c4c91bd
z987f52e7b196b12de3be6337ee4f5277bd67b4ba679ce9298289b998dd26b59d422b7f9993a9e7
zffcbbc44e11590ae68f8058bf5a02065cdd727f878ec698c71cb676e7d799169e9a671c7c04ad2
z20383bfb3a3e809a5626bc17f70b7aca7867a898ba712364ea7b536352e2888c54e383d93d8a7c
zecdd1b6e5148360b4c42da021e56d0135a6269276e97e5b53f0714459ef280d4796c2c5303c8f3
z1d86ac503d391c673c4f6c0e67a9882bb5b075617e436746003c1d62ddff7b5c4ee8fa94a9b464
z10814417437f79c2c713d82a46c807448a6268bb7980c47984b9838d8505d5a0f361d734386117
za265ac2ec6a9f4e646ae65105c166a3c761b1e29538454b28078f645313c105e10b0fdb20dc65f
z00997005d4faa2a281089c7b871fb0daf63fd8e65e27206db4436ede78ffb4b311acdaa7311393
z78f0b083811c21566775afeffbb8537a52b7369a71dcc86ccdfe7ba983b1a9f583f3003810a003
z600dbc23a8e3a8da36cf4d742b71fd94ecb9b7775b42986d0fbea5736efa9766c7979dda52c8be
z06c687aca18ed840ae586f20b4a48f816b7787625d4e200baac052cc38c176e0192d9baf691788
z89bcc75c984421e96abb9c2bf694b4f5f31980b0084a19509f0111b24938a7415928e2b776ddf5
z862708ce0433370f735829703c56e2008f07d6246762088ef189d245a97082eb93d92f25b42ae3
z5654a5ce99cee990ee93ff49282fbb47c56f53b917a06d5beb72e8fa2c5f8f57d2a9f9d2b2acaf
z3ca8965fcad180dc77ec5144adf2d9464536f18baee3a90a32bdec4bf38d23591af246d7359e66
zecc5fee7063eea85db861a7ca64980647e81bb4cae2e3fb80d155e5b8366056a548f868a9bb5b6
z96666f9987435cf4af7107bc913a52d639aedf1f150ff9cbbcd0f2a637e5192428e1aacc2b7cfc
z7e384b8b5d01ea201f702d7c9dccce455a3914e351b2c9c66d494769a1eb5c1d91096842a51831
z77792a56cfffb025925e933c08cbe67dc8eb49e4b4fc66b2f14594672ca07353a93d40aa2374c6
z589c3ed817c3400fbaa1a4e2ddd73b7065afbfc09a71bab3a81cfed6f0c9d1e6bb45526e2cce43
zdeebcc4993589aab5427fcbe29ff904973b8b2a45849976e9d5b086102fd20e5bef6cb83fcb4e3
z3c9cdadbfdc5ee0641d705dd29651ab8116094d158d41893c5f3b12eb664477ca6989634172c97
zab3d49d3c756cdfc6763a15a32154f8637316357628a20568854bde6c4ca991f94f04123dff7df
za46663e86bfb7ca734c76313d4cce8f6d4ef60f69d53457bf2d5308495d334e93b1ecbd89b8881
z1065fe259eeb08bdf86cece093090d7f011f592f5985cccab64af9969e7810652749f07c90dee2
zb3482f897f82c75516c3cc52c78b8d65cab6b1859f5d4f91ae5a1e930f4345d6a948a959a3798e
zc7defc7432861a2efb235e0eebbc77292bad7e0efaac4595f290bfccdc3cb8397c82e728f83033
zd370cdfc8073d6e5ef61b5362c32f711ab8cf15d64e7a102d1b9c37b61c3cc2cb3bfe2a39c04f1
z839464d64d9b0e61d5fc21254e1ccea5e5499effaf917f01544f9d6d1160f4e3fc3a19d053a446
zdfa044570cd0e03b8ea12e9ac448841e84bfad496d0a40b5c0707fcdebc21039adbf35c8e51076
z92f4ebee84bcfca1c14818b347560993c26dc5c0e30557b9f304c86058a273a35a0d1efce33c76
z164e20d7354543a87d24443e0503caddd1c1c28f93c4b5e8e52651c2ab4c305df730af1305fbb1
z0c16675ba96b3a9dc13805126457c77dc387058207caee79cdb2853acd745be6b8a6a2103d4a01
z77993bcb8f32f07a829380f5498919bf99182fc9342e3ae72e38070ee4d13d33ae17a681c30a06
z3fb9b584b630ba45c26f84a6cd139196dd226a33564a2968c0c7942d7a6f69ddc00640addb7af7
z07359c2715561adc4feca638640e6f0497286c80cdbfb3edc19208b6caf28b04eab49261d57113
z7f91142bd34c1031e17d922b4984baaf821f6b696a6c8c42ecabcf5a845b1961ba5da65907094b
z796db4e9212d8fc15210b4813d507a18399ecc86928d69943ab630d429a0634177321ad972430c
zcc98aadef6853ca024b7a5319f6ffc80adc83fd0c23fb08529b6763b487d4d82700160129a46f8
zd38f2d36b8e29279d3be44f7960edb32211296df3ee76b7992b27d9b7c68e5e77224a6b3e7a70a
z2a0afe57ce6a4dac1a6384c98858af077d79f6405b559021be67d16450f631966b94f42f8dd33e
zba80a0165c872705890fbdc3e41c020cb35be4189771c2b439f038d1c4b4010072e42c5a0f7403
zd5b86a7f2579418b1829ef1a1bab5d573d371a66ea2e9cc0cc03f48eba355ec3bc1157e2d38f6d
z6660e06b8789bf4c5f086d77c1efce07e7eee40be85d3bb48fcbc6cd9b20e72021d6921dab98cd
z010d3791ead006e7cb5554f42897ff4173f2307b388ccabe71a5be9eaf4a2e211730090414a74f
z83ba0af9f7acb513903b8417f0cab5a503f3a68e3a0163edc108e2320d54ddc5e2d8424ad85810
zdd6269a6a7362c17954c5156b3d85b829d931de893257c5b6f0b35eba280c44e741e1a2531d1fa
z911eff2a623342a39103df8368153e3e8f75be8b84ff89b113ca806bd2f27e8bc7388322939f6d
z1addfdee6a5a94523a77ce5afa4ae8cde59a6544db880854cffdb9eec6b51a599d20c3d3c2aa0e
z9379d8f6477c19a540d3480c877b6e605e8687dc801cacd5293080fd05d3635bc2259f59f69edd
z759472c022448e3ce452011b1d22850a8510fd30f12e9d69e080c9ea4c25ae3c9a6944fc907634
zb982f43f17d60293a038a6ad2bd4e1a3b1f6f373472619585179a48e6a3f4b3c6e11582c551a88
zd8d5c4c2381c1e76809f4cfeb19f8b7b14f9312476222f9b1563ad865a5b03da3078e97969c2d2
z8a3813444ded7e4d5c57843ca82ee3b5c1b2891f52bf3e8952fcbc47d71f83d3589293adad77e1
z91133e294a4825ff3c68c4acc37cf1fe2f19a2e78a8de5de0a93830786572c61a90b20e820d183
zb6f1a4a559a20da2c5194507a7db019305a35100fa13f1368bf12b0cc613fa8f2ce1b9abd18a38
zba27ee19364467a8358300f9406679d6f789a7b9242ca28f85a231bc6936bc94df3e945f7628cd
z4bdccb4c271e7302d6d98f62cd3eae03e74de0f8c705fb0944b30271d341119d1b6a8909dd2b80
zc0e2d3595fb6c0d149320165bc012b2637bc6d992fd2f44680b1197c9374ece0f209fd28f89b89
zedd3efa8d25e33eb686eb64190aca6220e8672dd967396b5ba3b5181abaaf9ce5d78517b79862e
z4ff391c5f8123ceaf57d022f94aa0c8546ddc90038a98dd525f5018b4d7acc8e7e0283969dc03d
z651d71db8f3764e34f405870a507a8f1b4885418e2ec22fb3a8782cbf52a4f8f8ca927f94869e1
z840c72023e11b29613a4bf57b4fdd7c138374089feda13b24a703c19f4e784c5bb139d6b3b7eea
za8301773f379e25db12d7f66117b2088a2d91ea111b60230110b52c9ba700eece6ff0f4225ea50
zde3b0e26108ffc357a7bf43201cf17a8934fae76f95060b4dd9029ca9c09b795cfd395311ea03e
z9521f797777900957b40b14d09fee834c682bb8ac6ebdf75e3b5d659ce5f975fe02a4f256ca49f
z4e36b6fd7037e5c4473b5e0ea28f5aa5df4c81471189f9e2ee3e6d1b989b2904068b78d577dfc2
z45f4571cd4e1259ebb4fc129b9b1eb7059846b36be3b83de110831a4fcbb896d75f54d233ce933
z1b648719fa9288b3982247366f4f1658df89ca7970faf170838065b9dfa3a7cafb6162eaa307f8
ze4410837da207a743c5d5d72f9cb34744a0d30cd1ddd9a5133ed253275b372cb239b0fed6c2563
z58031f3a213b54d604b52917f6c2950c030246b5d4a011009ffb74051f40a997d5edda43f0ad49
z295c5dcbfe8d55e11479f5f46c256a6873db345f4486b8f9ae9b638c3c94f1cfa27f92efe446ed
z3913e787d1f0f20e77ede7f0da9e065fb49c24a0638a51205c03384f7a988cd832a0be5fb5b0f5
ze541e47f03158c4503bef71b11180c49619c8ca3c6f66e8fe70978759cc3cc286d54fe4328a440
zdd7e3f4a3b920cd3a8a2bc2cbd2e5ff48516162b03f3e994a3d511fb67f789e4521d739183768c
ze26d8d9886125f2d965682a4d46f6dbd4d750b0d9a32857d4fa5da96370fad29b1a68c37c28f6f
z5bb4cc2f69680377111ef97a7de487479964966e0dcff5b68c9cbf89aa67f2b21d598682c262db
z14595ae57efc14afefb63dbe1f9516658e0c99b9eafbc383a22a073f62cfee5b7340ff94f52132
zc4500ed0d9f05bab1617b0444c18d81838d5c9daacb97781cb547aba8e752d3d36f40f0b579262
zd9f53fab1c26a335f64eff7328160a9f37012d4dd1e53a2d7a5706add40a387a36ba5675197ec5
z4a255b7361dbf91dbadd1884602166fdeab91e24fc48163ae4cd062c33478eb9a1412ef5c9f5cc
ze42b06afceb2dc24636aac071a69dcd81611b59e79daaf978934ce49b11349005305e054395152
zc6f93d7357c4f85fecbd0da6545d8ad4ec0561e10ffdf82e56d605900d1161108a4838d26686b2
z7694b79ddb293045ebee0b15fe62940fc1d29d2c859392c2a6a2ce5f39d2a97cecaa034560c41e
ze12c49e8bc33151891686f9a5f736bb97c6db1d9ee84da83142963879605d21a4cc62ec7fdd935
z5e9841d6675b99824cc9ccdc76e2b3f296225ac1d92e958847c3f1b61a08c50a636f56211a7b0a
zdaa89fe58e1eac18e23f916451404be0529d419572977dd3d4bb70bf2ff6301215d78223269394
z113764191a64088fb4ec40ba467331cf6452a43b3bca433a74a824982c3182969c1ad1ac9e939a
z94551969bc6744a5d00c1b720d0c5182d12a7a43dccb6a1921f898e05a2f088816f1304907e411
z198bd4b258cc73b2bf06724cab93dbe6237cc144d447821a3b0895d7e9837ea9f1bed27ad10b35
z6f1f35f361146300dd18ba57235e5aebb7a74fddaa9f87e8877d30dc51910275d11c1fbc970659
z293b16cab6cde2b84d239072ca3bfac4c30e85f849d138078100239b382b83a76efa614f3be9d7
ze30b1c47f4c4d2e6b18de68b21940fff7ccd7357ae35962a11cf8372e2384a9c83bfdf992b2b14
zb934a9ac9af0fd9255679a939099f7bc7a16e4c9b894d57112d1c6f0cf6f5207b868ff6f255da0
z4a5bb80c5f454ac724ccf422c94912dc8ada7cb3f6269f9f7cdf2f792b0b0258c46f10bb210f5b
z8b896b46a85678a22e07e4ae6817989af8f87dd8d04e956d25be3d9c4e113536cb1fb131d9e9cc
zb48c27c3d04b88a645ba3a87b471926c7a8dd69c1f016af78640c6d2a616c84bdfff415e67ab6a
zc04eed49536c54ca4288537d156362820971c4fb029d6fbe4ecfbab7bc0e04bb0049c37439fcc9
z21f3a3b7286a5c3b2ed7181a32f5c7cde9c48ebe8bcf98ce2057f5727897606ad044c5bb1dd399
zb7f2ceb6c1e7c13e4a74d8d3166dcc66d232943f429444b6b278f5b06c584e00e72f4019b2b3ed
z4814dd5e86e2f2f348fe96e9e49b584b57edf53a3a7990c19528fc619d461e6a6c2a6bb40949f2
ze0fdd550cc01c271b39f74cce5f402de490b02db0789421114b48b9bada93c9717adbef1a620a5
z057bf422483a2c174cf4af9dc0f9db2aef295b9dd0c7a5045432cbd45440481b86d7466b67dae9
zcdf57233e7544af6860cec1cde90f7997c77637c6b56cd4a13e2fab15a793f949f869cd3cb6792
zd1b37dc47e6667f0c53d02b7d298ab24d58faa471c44ddd764883608e7b22d9e3e1b279536399e
zf3c8ff43bd69ada8b48529d627aa827db21ee199da146cd6b6a0b15c8c19e477fb0df72b4f4dae
zcc14a4bef95f1f19766b54e2df0eb2635bac833266b725888277b6e28ab602354a94aa3f1836ba
zae34ba5d7e4eb56735fd414b1d7e2066cb29002e29c5cdf53eeb2b0e4ad942db979bbac7524d6d
z50aadb47b1ea7334787ab2abf1741c1b0b358432000fd1f07c77ac1e9bbac12a6f9492cfad60ae
z670fca515a166aff4c8edc741f8f5e2b23b491349f3600108c899b0afdd2f185d2275ba85b0461
zef26072ea5ba3ba261079b7b440a3a02f9b18cc3c3afb913459f321c52ad8cdc7a90cbd949d815
z3a5aa1acc8d2a78023ca5cf7c47d6f5732bc6f9b69ee05a4a3128d083f31c82fdcb0d78c36ff45
z8f0c25ad91f53fc22ca754c57808d7080d7f87e15bf45fd95ecb1a1c10f19939e5b21adb9b43b5
zf0e484bee749762c7baecef5439f0a83033cdeeb286e07596bef5eb18e39d6cdde149a44ec7bdd
z00ff4ffae8fcaeaee3b895a8f203e93220331e1574294827885d48849b28c4d9dca0ae96fd3d05
z6e169f6f55984eaaf82aab895056d2ab57f81d44b6b1b348623b9a6289efe96d1743476d5ae039
z3acd3f466f62189c24d17d046034ce7aa7b9d5551e5cd26839b7e08d7557d750cf70f3a3a506d0
z622b2c6ab0de13aa211e94ddd38386d4480988038cf6ecf7ffbc32ff44e15f690362b47222e4c7
zd3d845f802f0287581214e33022ccbf52938fcebb4beb9844ff78174000d449d92a5c451a9e1dc
z9e684d40d72d7809311d58122e7aeca2a4a27fce0eafc46c4077178e5e637823dc10b156550a64
zcf7b6fcce82ff7be9cff583d98fa6df64eb489a94831d25e64e198e1af29a910bb8aac9495dd9f
z28c7cd8e218c8dbe9ad17e0903d9173eee2681279441b4eb8f6ce0887e580967ae4ebe29f639f5
z0de7fa9fe76ba68b4c27d0bcd6f8a130479e3e928f3235eb34ea415940abfe2f2d2ebb338cdb8f
z9c402d094ddc3be2d988b499a45f7dcdfed64041d8f33a8e37108e072e0a230b259da31e0913d4
z727f6636e86548f608c8b1425b42e25a58be2873f2657d7b95c4c962ac959376ca23a672e28aa1
zde456a5ee422adeac043684843fc7685e7b07eccc72321667792dbf609a44fb5762fd550b2f555
zac6330eed9ab748b309bd1a36906a7722bbbdd507904309842a413b52cf590868959cdf8a7d9b6
zd54ddd71dc094a8f939888557c9f2d288e561b7b2bf997cf89e090d9ce8fad5c5264b1d1eae6a5
z9c1bec62853516e6c23b57658e23aea73d19b5ce41a6ca8313f53544fa81403af5a0213139410a
z1890c9d73a089f50414e903d2ee60e5bde9f7b7ced44bd9467e1327d88b40fad1d452425f439c6
z3e554a7274090269c56809df3ae2848948333271b21cc783003c55f6aebf9fe208d7c0fab1963a
z016812c745c2547ef817d86559ac1ab4e612b998a891f7b753330898cb136bdc2dbc27226a3b01
z16b644f57cbbac0007c12193d6ff69be42499254fb58e004da75da056a2054985782520474bdc6
z1e9e6dbd8ac4db07d1b402311f5b0cb34a186549a5115d64465a69e68d91eef1fc8fb1434536d1
z6131b5b106861328854afbb8c70b85a8cd425bc29f73604883f7000b183837b77a14a0e9fa019f
zeddc2141d52f312f45ff13eadf2c3e672151bdad446d16dbc60ac0d4cf17a4c4d9dc803e59f9fc
z62e78a92605462dd69f13b1552c0a19cdc29a1bf895ecb0ba873cb79c585fbcb278194467827d8
zd431f4f204f43eaaac2dbebc1f57c071145d6bfecd432bd67d8f91aa94db142e427637f7b3accb
z5721c6a56fd336f61892137833b68e9ef781dc97357f07c7c668c037f49ba19ff33d206cb10ee4
z60939bcb7de3847422df91507c935d9e609b3fddb60598752778a7184e1175e17efda86645d453
zf6ac80420f25205c8a8baacd6706e0fa6fd6e4a804a55ff346dde559f712eeeffd324f56a6db0e
z06ef371a35d130d8ee901728221f7da4d0907296559f5b695dfb75e5cdb2c53d0a448f58c82ae2
z0824b8c05aaaa5189b4806bf6e0c32284ccbcd3b7e296f338655e44c747cc14377ffccf88a8700
zc085aeaa26b9a3fd6197ca316e7ff661a5e463a99ea89d12c30453a3c38f2fa31f781bdfee209c
zf399a16c6d3d2737de6c3dec4ab451cf2d9a15c0e3d23ae7851a1ea78be3211084b7d3c0f28705
z2adbd5667a6dff4dbfc8a91f53d4427f894358771edc1520c21400eada5e3ceffe6085a905483b
z8c712b17407482153bf7a219bf3546c81e324c899d984cc0ef7cbca187f76c70a95271808c5abb
z75f3dfebc362a598e29d3a2f8cbd2d679e857b93a071511e880cbcd927e808a226df0248d233e6
z0f708ea3379cf3abe8a384570a0164221477e6148f11eaa2c30223e045ec08a41b0a36dedc3caf
zb2f465007838e47ebf18b7b89acd025b5cf2a4b6a3f66d4d18f34a9358735d9e5ee40bf3a2c988
zc1943fb5e2fa051f6c8f91c138d1ee02e4ffb0a48ef27eebff7c2856d4cb48a4be52be1064cd20
zae390c4a18adf9834ee96683f4e724b96b681d4d8e9bae915611d35820f8ffdef9ee8f436d9a5d
za5a5bea56be21d81a1ca089dcb4487415a40f5d619f84c3324b430935e3b6c47f8cfde9cc06b8c
zfe7c6d6a7a1ab2de0f08c64261d0403105f6b0ed7f28ca6a31211620a20809cefcbbd9172ed163
zfad250e81d6802e1744b1cafd3113c7821daa2f3c106546a817f80fd67607ed87111cad1cf38bb
z72b99ff337128f57c9ce5c49534562ba6d686738f222517d706e50be3c032a629824bafe33185f
z750231a6a2579331e383eccb03462bed87a8c176bc4ee60e62a0fd918af5cf81ce22cd2ee4d172
z24b91867e9769a441c1726860e43241de44583a0d159378e892fed9428e5e8d28385447bb19ca7
zda495e7b3bc20083a921a094fb834c0af1103a71d112ce4e4595c4e35c1ef39274ca7e4a992e7d
zf8dea562ecbcdf26d349474571d10d9b81356fb4291b2240f3da1e3ee8ccbd5b9d660ca1a52627
z9ab7386cd23a40b7f3aa3b4e08980edb9c4c63253629efd36cd83a651b7566dcf38999fdeba56d
zca71b727609559adb5128f30602fea2f781b1bb03974c06c5438c208dd5a705027b89079f498dd
z2c9396a548cef0677aa0e1aff049030fc6dd3bbc3474733fb6bf522f7ec064b1fa35b045b7ec7d
z6f4a96bc02ba9cd3fb646f4026932b4d84f37e054d0a1fea1f70e593347aa9dbcebee70d6a2f90
zc35d778d94531cccb3399b8b42c8ee4b939c628b78b3be829f768406d471f32c38d0532e96cb95
zfa431c104eb0a13d47b1c0006228065775c2f6c210f50b77865006cb1b40140baf572c53c650cc
z96d38b07a660b53669edb9d6a88776f069465ad7ed1c22353dcf3aeefd58ce1c05bedbe2e48318
z12e33243338d05b4f0533278de9a2c8ce32fa3a97343233fee5532e6d438587c437a017edfab06
z5ea40358801666f08852c36ce5ff5957706cf1a1b4248edd532d1152aad0042857f7c4ea7282ab
z1dfea54756d3126ff9cb8bb7a08b9186781346cbbd97353cc1b01a8200e5cc580cc4ae58c27246
z7d2e3ac1368751ac04a520b1038adaee3929c4eaee92db9b402b567e80cfb2d8c6cbdc7de8b6e6
zb853aa77be5734e1a63abb00e452ac40b500f32286664ffb3433482a7957ed1497acdf6469b02c
z078c953122af2b6275b8ddecc99dac8e24dca955f20d7e1363f8df11a13e813be450b693225d91
z1c0ae560679c81ac6ae38c97fd991df5be12c7923e187a2d48bc2ce0584ed771b16023908d7d41
z4215057b20c50a33b3103868c3aad4a71beaf620b731f59df5d30a6651c3ff5cde267c8adfba79
za71c60db4f3b946425300afaf92a5da0e75685c32e08fd8d1151bc03d10e774a8696c30b01d74e
z7c161c10671a59486ccc3dd80bc365b8ad43714eb51e66aaa32a6111c122d6ff212a0b603fc823
z1ea4c71d03c51c1411ca7a895c400b8ec998311074abeb5d9a2abea8e689a71400d7aafb83e4ef
zfebbb0ed8f37803790a801129cfd458e159e17d9b96188c15fc418ca39b1b23a6e2d8eb4dad1dd
z846048a44198a09dd845de940bf415fe5544c7fb7944fc5203c9afd6bf1866feae18f6c8d83694
z725b3dd241e48c0d471b20312b7869243c1e6e830de9d2538529803ddff9b923a17f928f0e4a3f
zdda2350cd751947f643461b5c11fec05ab214b4e87262feed3ad8b5326821d093df4a5cfd1cb04
z25a7b9cf75e8bc194d5b1b0413da53d52d2fa099df317496b9b0b68dcef1e70226ed359828ae4b
z5b4c9e161bfab9bd9a013aed3dd53a963b0c452ca71553dd453904254cb85186284f90f6866033
z5fb7c975cece0e92e61b45693ebc4be76c86453c036f9ee021595e31cc4b807c4fa436c4c1f686
zad8a9e250222e8256b326f59f6c1561ad25dad73629ee294534fc7062e57ce2e448349932506a6
z8537796ded6a3cf1d964bcc6fe9b6dec433b1a9e06cbde695ff562c574fdd6a519dc26b3d94971
z71b75d4c42eb0d5f5dca4a32ff5bc9c682b30ac9d915cb82d11fcc2b95fb7ec25116200bc0943e
z2fc7c4d5f19246df7e0628503862b1203eb19af7dbf46c22a925f5053c321fc349ea7331369fbd
z0d83bee86b62cff77ee563e40ccfd2d4c9a16f3327c5abc38ba99071c7dc7405e5fb1fc8a57d1d
z7636aca75399a5ee7d1048297c40444338c6589e7a7a0991ae18225eed24f77a2e79c44c09c934
z5b0a5198988a1fc23c29a9335becdcd81d7b565e370bf47b27331445841194ff3722a8401115c7
zb1636079d734f2e813c867405da494bcb6ca92fbec593faf30bcc6bcceaf55afbe55cb54367672
za7f57ab32c6070ddd616668fe99f585af9a77a2cc84f191544be8cc59a6ceb7c8e895bf0710795
z06dc106836a7239621dcbf16ce694e7f50266d9372108cc243738c924c63073333a539c8f9f582
zd55ec89d6e34539c3eeeaeddb6e11e92e39b2acc5662061d94cbd66d2acfc6cc69f60bca89f1ff
zd19ad8ba38e69af1a2125e69e0e7f6d0ac12f5a8c2d1fa194cd5951bf14d5314036ce4d32769c0
z6059f2bffeac8dee9bb76aa5cb82645a3eae3305b423cbb539c9c399f746fde1bb975ec6bd96b3
z82d69c5c5569eb21b3f45f4c9f959d45172255f53835d262786db43bfb5cc44e645381997a222b
z9e5ff5d6e2807c49f4f24dee07b8766c26dbdf05049187bb7a7cd040b0e92c767baa2fdf9a46cc
z1a75a4c5381901c976ad91dc82aa7cde659d9a7e3109380dcae79952c57706e1d8e5414a400f32
zef692c319825e8c4570fabcbfe8105953e6ffbb4254f24b1ca072fb07fa138d842c62dc76c25c3
z8bb26bf722293163092730ad98fbf2d4970b886c8efd7a47015938186b8427bacbeb95da51ccc7
z2ad0a99d0c3342bd5fd10dffa69ac1d5a83b5d44f244613f656d4cb5c8dced54cc040b0afe0e9c
z9c7b8d04ba600bbf25e050d1245cc1ffa01905c1976a9913aa359d2ca9ff9a3acd922736f7aff7
zd9fd9a42ae5de5c2e3607a402903f95cc7e4a6577dba8e35371e9d5fb791cfd072b8858f2f4e5f
z6f897c57ee524e4e6c212d3b625c4b9ac32b31ae28cb0ddfc8cb3ec823d8f16d9de934822dea71
z3de4ad6b2a75222325291ec15bc5e1da9b865b8cf67a14a633bb8c484306474ac83306e795f00e
zba0afa88dcca0e78fda11a489214dfea435c3db16b7a0081a3782dd4a9c69cca361e22a84d193d
z1476ebec14537aea407fc6079b3587eb0e935bb20b6f033137f00668986fe8291e3730a5bd28b1
zd25c65c79a2358fdcffe70f17806c9f1bde9486db6860693a41a25ec6e21638c7d9fea634af8e2
ze518aca56f9693a675ca66e5127df18760a8831efa04ee207d6b82d92bb946962480c983b1d974
z7d8c0873b03649a5d5babc2f65eb04cb22696eadaaa227edeec3af03cd0c7a3571c14d87443f66
z00272ee012ed988815d909af14a7015044e684bf5f02ffbdd5d126d70a529d14704f41ce0d4f61
z8ceed11ed115761f14dd0708cb2ce6acbf4b364555165a06d973562cfa1db98ee198d39bdde607
zcb984fa8235342e3f75f8de8a7df8fc5e9b4657f40f607bf302bed2159eb4b7e5c7d727b066157
zb1e7d5dc1e45e680f26093e2805ad6deb2d996f56af74b31b40e2ad4f64fa208cb99931bb0da85
z1747f5e739c9b42253291346b18bf4f2723d37c4fe736721fdde5703325a9b9e929a66b05c4e17
zcccf63d6dd6f45d07edbeb090ee46418695c8629c9a3e3b99381ee377f3d98b92519d2b8cd62ad
z759ac12ad4856ba322571953db0f999cd34312cfb5639b2ecd3a2921178c61a147b558054f8bbc
zc0b9a796b37c9df4eedd45436a6e8d263b3c5557fdbc26421aaf5ecbcbe0737e424bbf73c8ee19
z689f5569bbe60a4a59d9586110db865ab21567f206aa7d694af8cf8ae172760c8c3eba1e255dc4
zd0e8ef065718801ffd1142c804b7f6a42390a6222fd73aa339b6148c12b3b6294c7f50023558a1
z0175850c9701d200bdb9a4ca848ab06c82cae32686af59032ecf3e04c056c2d62ba3210322db93
z1c7be852385ec217cf667cc548fe25c48acaf5536bf878e1c20c9eae13007f82e3f0aa08995a2d
z26c4f7b222d57a6f52dca6d2a68dd3d4f4aeeb241c67bef5917f7e46e4672c5884a41d22e32a4a
z54828f115cff890d148027e52a80229ae21b2c1cd1361e3d55364132173b680ce4a1df819524f6
zf9d2832a41f9bf2b87a27838f3aa83e95d18721f09ae253834fddf21d26cf6f0de91c3a36b5bbd
z64d27ad38aabc3ec6b6ba749fde757c1bc2b01e1691eb35ce3bf82a67cffcdc8d7ae4461532abd
z42aff59b38ead77877e4866f760406704c23ecebf681d3c0e11bf9d4692cc0850096219ca589d6
zd4ae48b7acb4b05895e18afeab81cea853261ad09ad62da864326f5a007fde489b8105849f0272
z961a5067dbdfc5ede6d23dc30bbfc3cb3cf1027d535ea8ea238a3e31bd06f02e0a55332b51b2d8
z4aa66ea54a3e91d000ef3da6897d9c6ecb3f2f40795e1888b4a9ec5133cf08afe9110997c938d8
z58be3deee34b7668f1865d589d9268ac6642eb17c71d1938a5cb4a20ff86dddb47583baacf8336
z748d12103ce288ea230938fe721db624b9d28d5aabd0847f68e10aff17a98a9c8f77698d362ca1
z47c179d0a2ea4a54a2ec896cbe3d941feb3ae4f67063efa502760e47ad379ac3fbdb5ea08cad93
z67ea5fcf2b8c96bd6e56b4a6cc191a1581029a5ffe26d2654d0cdf62c2d16a000166c415f397e1
z10878b79d8de1ef92338d828c73c90ab47defbc36a8312c9c06ced80bde8ab54cde7f5a34fe668
z0ce312674e13f268067f1804b75e143215ff95063852f80ef5c1b90e0ee614c4fde2d685c29c64
ze09175b2e61697d31cbe2c7cb01ed36dd8cf5c5055ea2d595548ce0dc2955cedc52d0d9a2af847
z41b6c435dcbb2c2c2f6057d3c26dc9a5444fff6ba247ed6d7608e64736261ca62438b408a3d512
za2c96e3a3bdaa27fa8d50918631262f06845707f485c89a5f5dd909187e378fe4ce0e921bad184
z66b6b1f13c4a0ad326cb812be3613844b21533d3709bc19bf34583d9c70691d33a2209c6bb0d66
z73ba52ad73e9bef82abbcd1082d3f6f4eaa2f7f41fedf71a13fbf37450b214dffc810c3b096e7f
z824425381c8127f75eb5b30ea15d160f8af912990101be6fd2680e918d2999138e3fcbf4f4f586
z8423c278dcd49cb61abbf585fe5375e0c28c04b34be107fba9500ddfc20556f6ed9ae38f4ac15f
z27d3614c3ca82f9f27915a773d845cd6f2f77cab631da194d56313e2f05b2c6bbca872358aa3d7
z4130ec1b7cc0aec33772459ddf7f2a62a62328e0924773852c10fe16a682660e9760c564e8ba32
zacd39de2695d6b86f198b6b53034e514c48d15d83deb479818db3738f8c951feee7180ba3ee062
z1068fa93c646d432d432a8e45724ae2c13130b7a3dc753b9f2f02ecdab81af5bb62585fb4e818d
z59f3b41af9f5b9e16a62f44be2f95167242f977305d9d4d90d7144309d8a94b3bcb89dc1042092
zbf545870f0d3d09c65ecf6faba74bcb184660491a5ef67167ee2c8f7ac0fdb96e246594f2b183f
zde9f809016985db822d65073fef913d2fa28417f259d5f637aad74f819d5637701b24eac68fcaf
z2e5ba2ecaca79de4969122389ac2a5d32c81086c46efe968ab3e1c3900adf06cf4697764b50a92
zc6378cd1ab43021118f5c2ef710bbc5a62f2f9287ae2d4a3d9b2a2c864839e1681e9041aee8f46
z3b6130d04c10ea73c9843aaa2f2286ddf269299bcb055e767d8df182f308cdabb31c0ce4ddcf39
ze16da13d55297625b3dcc202fb34bac048eb75f25dfa04bb884142ccbea119c655f1ad55d0bae7
z0b502e114819316d36f91f681383dd0f6d9f93feddbb947d848a6306d8cc30ca45fa5dd666eba6
z8f01230b5940c896647705559bcad7ea74b91606fc1eb201eb07dddc1a620d7cdb077f66b873bf
z58a186f82c91dbe5ee58fe74b6dbf0f85ef8b35dc9ae5f827f4e3c525034413abb22f374317d72
ze4136eab5268a29923653b35c0c50e22659001df074f5b1f651be3cb3b4f1b0998f4e1ab30e22b
z86607aec3726a771fa2ed26c1dab651928934947444a6c39526c8d9931c126cb45119e9faa4953
ze3d3ce5ac6ca6ece97f510c40970567c6a554149bf589ad57f01ce5c61e4ef8370471a5693f788
z3dd4cf7cf1db09a6d99c1fcdaff4e59dc9799a6f5241632ba8a435123801d50b1a4f28b5876412
z31174567c5a605333a7261414adbc30e251eff8ae813ee91b4f751676123a06df9747ded82426b
z0cdad304e8949ae6e42ce3adf9584fd8ebe5bab1d1395f5b7dc528139237f49d5e677e4cfb87dc
z2171220c1b84aa7286bcd51b3a7c40731fb636cc4a06c191cb935415ca2a90c5dd164efbabdb3f
z85c6444e17af3b06841bf0b47c34c40a19792abb3230f4894a65e9e3b1af09ec12e279e68d2376
ze67f00b94a9761909e8d47eb0e4b8c625f594a300d944a761e4720a9e08074cc2b4f1ff78dab72
ze4fe5ac71b6f673222a231427f6c3d940e00a845db9aab34a9b50af834cb0406da62ab5e8b6251
z5b86e1d379875f745005ad852547daa87a4ba5f50ac863ebde84571564b376d4c17f2e5923ff7c
zdc50558986f7d4fc5ca37f96b2cb7da72d34a5d8271b1974dff21bafbe5de9fa9401a2072a5267
z59d837e65be026490c86e0cb089a10be5f2ae8a90132aa90a7874949505c7186c21e3baf14cfd4
z398e23f2771cedbb3bf77625c763595973b39a4cb37c4a9bfb3ae4833705b7ebc98275c6b82a45
z5391b77027b06ef5e9fb07c0fb05e6b4dda61a2aa8c7d97ce9fcbaee47f0ef0a09cea6ca4ab2e1
z75aeba1735da730049282c85b8b33dfa9e80350ab728f150c9b5d0c0b5fdb66a0e43ed7c8e5ec1
z8d8e30f9d35539fc8cbf0f47b7064ba45a52ff861e79a03f63afb8a5ca6d979a00bbc38d36e846
zc437a7df166dcf0d2fff65bbda2cc945963437782a0443004d15987142edd11bcdff11302a2c45
ze31184aa913be6904976559c996b39d8cd0c92052b3e183d27b1127002cc667fc678062dba1c63
z932c50c55562eb15e93fc77181a7e3bdb9bfb55e6f1fa1a34d969e81afe69ed3a4d8f1bde7d4b4
z0798ca5418e111c187d339b57a834386b804f7178909d8d5ff4cb112b41fb95765adec9fee8332
z744df0a19f5b16a8b4f55f9096b8b5930b187f45fa3288715baf5a9da6c83c82fe9d9fa8114173
zdea5e174e5ea7255449fce7c4a891c963d2f22a785a049d61b41a9b598d1c171863f5060b73d37
z28cb66fbeeb7e2adc40f98b6aa4c9413e39ab45e9bf705cca81d4e906b38b6b0d9560c640972bf
z50ced98d8de1d1393497a7daa6362a709dd51868807ba2d33ea4e2c9e2cf64082591c3e3842666
ze8a28758db27bb88e6eb109661b1670c78bbce3598599c8b74911ce114e5481afb2f423be9ec05
z4a6fdf9054c5cd45ccd7ab442839635ba357e2429c8841c7a48152806689cfe45c626509c0574f
zaf1108b5b9bc36ec89750224b6c8935a73424902fa732196b9b602a68580e48e382ef3a43709e4
za3b0a1e139c20dca1f19c5f01b0e644dd821ff74265e0c2f74cecda21c592c9078f5f5562817bb
z492f3bc0855fe03e646f142366d5e69953ac183a6eac94f6d4224045c8fccb86fdc490d859f5da
zc64e8d5ca3e8798481c33a02a8536ead5c8bd301f67009b9969226d6373ef2a178af9606b21288
z5c54664e2350d9d7b8c30f8d3077a018dcda4dcc34dfb6ef82d527a8506703f6873725408c9d38
z53bb2f0e1505d9a59850bf568e8241c36eb0acd34b7f3e37650fc1b925cc718eb251a9f5af35a6
zee7f71501e992292442c9e0d0760309e4f7532ad823fa9659dd5591657597f5d694489b0faf6bd
zb4372b990f360ff422b68115902b624f3afc9a0815620b6093db8147f74836ad4c3b6389f0ee60
zdda2990490d9006e8eebb2bcad6a56c109573c352cdbd8b56cf42ed9ace02eb5a37d6ce615503e
z31b89fd059425fe4ba1cd9b68b0bfebdd4afdec32e1a8e8c2edbc2a73b564c867b02fe27aa97c8
z06885542b1ce18efe5af296ecf59f082ff30a3c9773fe472f39d94edd425dbcb7851298b191d97
z6c71b95480b3fc6785f3dd84731c5d5fec6f47356c78dbb0a53fb8a8b85bef898c7e2b5219cbd9
z3420c5c03f63c7dd59802602093d6bfcaf79f7ddaf0668e05a4bb6094a44049d54760ef638e2a5
z0949bec1525275046fe8ee39021dc2cd56b75b24ac7ec02763c025dbf46396c4506871902658a0
ze0dc0496b3aa4d077fb2d402700028b4e66f967f16e3c00cd290c3543297feb0506f4feb38edc4
z758327f36df1091457a2b2982eaafc85151a46ef5f9e4d6490eda362fd69225ce91db1e716302a
zb518899e3bb74005406606eb2641d973cee21507dd2f69024000273769f92153c59ff92f8863cd
z1f8983c7f53ed0e18c4d0dfa7ef97fda23acb26bb42e67446093099008d2ce9ad94895c2d38516
z57b06ee0f77f58ae7c2d37aac35175835352b84e07cf9a65cbf0b5faf84a56ca4422191441dead
z55d823bca939cf27e5b61c4f0b693752306211b4179743b9ab7d04806792d065dd051e54c179c5
ze29ea7b4265bf62c7b22e3883c991ab96326d04d98b1f60652760fdffffd7448381e0616955266
zd51bb37be533c2c3f94134ed260710752137ca71eb691ab5527f13f313af8de3fa7affddaa63a7
z910082791bb5b84add33a4ee9051784931ed39438f3eb8e7edaa039547b77dee0839e7c5c58369
zcd44fdfc4b8889f55d6cf6280ad83db690bae2eb365bfc5afa80486f2f333bc9630827f16a437d
z4f3b600d4a2337b16aac1b99329ae7efcf3059bc361876be5c485b4a435d0cb0be6b97b0b7c94b
z11c91aba11949761bde12704876c3fd3aed52f85ca24cd41bcc284b517b9e5d428b2d81546b301
z8ca61cdb7a0737e568983c404f708293268bcb62b4200b43b7271a16b95b83724aadcf22cb1cec
z20442add37c16c757de7e027ff3cfe7186e91096126d6055ddcb0815604decae3182c43a86e747
z515c04b3a953428fd15ead3eae15eb0f9338963f404eacc5d71f9651a712a14f0d56ae43bee5cf
zf5cdf6762805d72c37e69d4a3d0428ef8d8fae777b71a980124dce63ede5d63216f35579e77d1b
zca57da82e89d3769f341a02c16776f0cf5519a0a0d3d6a4f0202591d2415d908a28314a822b0b6
zd47fb5e0dd8abe8b7d1465951a8486d806347dbd6bb114f7e75d98e9fc1f402b363d07edebc028
z1218023bd206361ab182594173d1a97727c7437e399e314765b664a0fee59a1b41c2e130dfeb8d
z8ebb9d69061a56dbb37d30a1383324e120fa8fbab59f7d8d7a31eb89c31ddb758d9fd92816f4de
z5242fea012d3ef9a30b9f62db4f06a94026d5b9465f27959cb67edea23db25cc9a62452f453223
zdd0aea3172e227dce854bf511ad612d0019be7b26405d9ad1043a41c662d45315331cafefbd675
zf80122d311735081cf9d6734ec7481bc764dabbaa9258fccf05c7c07c815760b676b37a3f33008
z84252995272a1ce36906b352ddf298f565960fd84f4ed4f2fe867d3d2afec084d3d3bee18a9785
zaa320609f43d4effe29d8a93ba32ea56a31cf603da00456656b8ff06167ce202253a67be3a0906
z35e46f99d5b9c24642124ca6b488fd30dabf7adca1c31099d106790b941e8bbfc3e6d35f97765e
z96a4389109dc7c5fba86ccd02bad536577613f405f11895254b909f90e6df80431acd51a8bb541
z827129d9a8533208387b1617cf3c53811f3e1850bedf99272aa186385a31a886ef2a58143c2146
zc8d76a675d7798584feae176a49943572825bbe651a5b37abed3b1175945920a23b0d777c2b228
z2210963387bc78a8b99e16023a21350c80d37e0155d5810afab878c79d15aa0892963b4a5f0ffc
z4bdf88c4517af28b51612934d68ede22a0f497fdf37a33d15370c1228a06eef006c19d29858470
z1cc956585119e4079c48818a39d84b00bd954a92a96f385714a643ba7a9cc99ebb16fd48f3596e
zc5c8d6607820bc0e4a1e25ca9e65ca568fc816ee32da7d09732538853ac2caa0baa946052b9f96
z19e6415bdda524e05ebf3eadeef023b6e92d1acb0f1073322449dc0fbc9303a17d388ec472f01e
z7fe42e51d92d79bc70769a0a59156590c2783a32f96175c10b5e1e8226114ec4270365cb5699cd
z9e009cec008d6177f8381a24325563f103fd63316dbeacb87671b88a1454f1dfd6ada473b57136
zc3cd99468b0cb069594b380c3c5e25a1bced2d2fcdc98a8c13a2f2c0d960b1041df02df4bf5fc1
zee5e51d76c447171da72a23befc10fbae46c9075d8e8c08e95c3c3605403e084422a569e6ce27f
z9891cfa1b8a089035c9935074cb0c5e5768736a900c85ee77a6b1fb02efabc85f449ec0260a75c
z0a4ae5012edec9a33a18be895e0edec79ea80b0593e7223e8dd7afdda3ee03cd1a6311fae28ef8
zc2d1dd2bf34169aad888abefe7a0338e9174ef056b3770d8f0eb9ae75cf0605c3ec726907d87c8
z78f8dc2d98754599906c3a021087fea6149ee7ef5ed00a7035fa63f03644bbf5475a75aba89fe7
z21e8e81f86a3d038163a566a2455a6ae4e950cbb0e3e78dbb1ae79effb5591d06eb21518283a8d
z4954eb07790e4f9d8bd6bb8ea33b4dcd8ca075ae52314c1f6504a1ddab615abc312529274a45cf
zf99d507d98d3da36a6269c80fe9f0fc4bd4690c193b4a1b21080ac2da3005793a4330f4a1bb5bf
z911938147273fe93ca3b2946712ecc4ed4c2b05bb24cb5e1962d06185b59959c769bd5b356374d
z484b931ae294add10c117a5220bb7e63b1b25f4ba96ab02eef6f4e4c4e22d7b13e4b12d40cf2ce
zf70691bb2bea21503380cd2323105f2c505270dc805ad1bc2239886a8da149425e52b7ba2a93bb
zafbfc894d4da3f62e427aaa8f4bb445e9cdf2f98deed4d33594384a7d9bbc8a61c132766c863a6
z086e09f68b7b70a741ea1ad5e841b69c153dc36375fdd97a9d318b31631559b81511180e87543b
ze8977dad556c3b944a57a11caf1fbb6b0b6cda203336003ce8a244ddfe7811143462ea0c7d9e6d
z4b2fc4fb858656cba5ce68876fce250952700008085d64bfa32e1642bcc4639a60f60674820e36
zf2c82767153632294e8d09f93bada42162320d0fff156e5749f0c1cd87e73a9a5099226e1a6883
zd2b86d5918db1e342fc8433416bc81088a083629066f5b0533ed8f20f93200a2e49c8728d76c5e
z2fec583a7dfdb17d0626bd59cdb240c759bf9dddeff8f9d9397920e331f4bb0537b7cac5f7c8cc
z4227c0743e117b2737364646ebf4b712d6b94176b4d519908ac69769bfc77a169264b07a401b3c
zdc60f8ce6c53232fae7481c5bc6467ab2f440eb45ac033e25200c7c79d51fe88e17cd6bfa9e400
z8ffffa25be0c65b82e2e28639c7e109ccd14aad5954905fd3bf7c58c80861e84927b214638b75d
zc22008fb28d098a336dce2c218dec0b8e02d176d275462ae12c2133b0bcc66b09345ca3f99876e
z28245add51401f205b30c52886431fd8516013c9e8d614eead0d52173f0a713adf4e3ee95b0870
z6661c2f845900b9268d1e30174e27e30f92f1f6631731db137c61c254992baf560271a05e259f8
z23d6b548fa7c47ead3114677af431e4e08875c9ca8f51637d742f08c8e8db22c5efd04ef0c5c83
z45de7fd062835d00e99a5a8ed31118462a624099942760b77acd3f19ae371b5c8042158a2552bf
zadf27227e8ddd15a2c33765ac40f055b6849339864c05b942502f792e49f40a115a66053c6c1d4
z4c958e0a56720e84f23bc993430c35105f703cca8a9f3baaf05441b322de95475cda58219c7b83
zfa711c10ff9ab53c15bb8a5de6d966ffa86e433e9f48d4b905cf2cba4dc6911bcaa7f873d8814f
z6ed28ab78bd30509d36a38f9442fd93b82cd6b289bbed1799b6fc97cab2483e9239d69a730a481
z17aa3e2f475c90f12a840e8ce02d2e74df96081bbf669669127b1a1193522e67815d6da1f803d5
z05fae83e08fa6ca4bc80af999793f8492c401afdabd28d02d45a62a44899143b4dcff977b0615b
z14f636fffb6cce2e6f5db9bda86620d3bff33269890b8fe179284e62dbe14d4ad4dc9c92a36a88
z849ac5aaa4718b783a1f53c0552bc3112f4972e998da3792da27bb119424e64aabe2f71b74185c
z6d83723ad1df627382a49267bb0b2b1cdf6f89260782bfff851779c40883cc6144e72a1d922e3a
z00eb7e4f8bc4a8888c13cf2d44b660e7475077cac7bd5acea92b59bd39fecb42194ff27274a30f
zb16863dc8f4d5198504159d48e333bf03c7f524767cc7d0e1dc7f29e0a11c1de60fb56a8ffcabd
z235648041850870f32784e6c359d68e008c73b0b42d9aff539ae8efaef8d6c71052b284f0b69ad
z1aff9756bd48e1b2f3225e07159d6418c127816ac4b47130f22d40e019cff73dee74570addbdf6
z73816f986a0cf6e6d588c110fc152fa9a5e57a992c57feb0ed86884f03f9d4955900f5259cf6c7
zddda36a960f53b019fa79eff9bf0f32e2ab4d2d071f615686e1ef5575ea5cd82ba9167140e6460
z7ecc675b25b04a4f47657e0f7476a79db65d6f4e66404a0a22e600b9b9c8f96786be3b0096200e
z7f9d410271b6d4d2d12520ca55a5a80bf5c09da6687eda7f154cc7283fa8b8c9dae5d3936be968
z16eecfbbcbc2440f0014e4058cb3ffd6139cbea983504012affe1fb7e9e59489c9f0e254175a56
ze37b61dcf1b7fbeef66de8e3c430acc8b010215e540fdc08d472d41a3eaa4c9406fbb6ea1a111e
z9c6cf1f737ff7d3e284b0a3fc974f46c8a4cfafd5587ad344d8ffe47565b665e24d5b147a52a9b
z4f95aa8b3fec628f449dff0ab2cac2e698c9ae67fa699e29dd8252b3fd4a269bb292c53c2180e3
z8267947f5a5ff5d525a2753a8bb518aea8a0318e7e726baa42253666b27d9cca0ea33df7d3a8fc
zee74fd8efa5585eee883ded4d175a59738bd98a92e54b004be82d5f9b4bcbb968228e215779dc7
zf3b6a04f5d584c1c17dafa6acd911d61af2b5ff4efb50cd0b613dc3daacc9dfdf49576a2423d74
z499bcbfe93ed20b1f78a77783621cf713eb1d899a9c72b4e6d6c3e49b1d846b3b4fb440623fee5
za27d34e3d2b706845440f879db8b23f0df7cb36dc023bee25e5fb28ae1c0fcc070591818b5cd42
zf21f046bc408f80e412e18c0250240449e8d13f920f7a80c9294f3475bd63b3d8c62680232c317
z9d26c25dce19c7770c367a769b80e41886379dfda6002163744f12de0a413fb864a45c88a170b5
z66d5340c783f9fed9946ace0893c02ced73be4558d1e635fe0240e03676ab6e8d5e4a316fc3fc7
zcfc4907a81021c7fe899f8d82161c6b9033347cd4d602e083640adf5432f65409bee52f53c2040
z7cea94be4c11da67a1c894fb78b9940ea3fd314eb04f2487ea802631964e67bffa50fa4d92e7d5
z1f6b437090d44a2850dc631a8d43787e132f4b69e41e3588a19f5ed0815a13af3e8d279ee41096
z7583064482927540840475b80aa26f001873a510118bc8fb067b31bb670c41ec467bbcdbf37aae
z9c6185dbc71fc2e23e893639d7f7f4632d3a35b6b40b766b285832deba985fadd8dbe9c3dd89aa
z1f51192a2f724cbaa11025809cee01a38c034632de99d52fca9d469c38f8ff35e8f9b06c31b01a
z07fc7b634ba2c0b76a60f63666e92405c1c2f72648f847d3a966ca9baff7328d250d9299bd26e0
zf76680df85025a134193e6cb1eb0057cb3edf4f310453977e8755d07fe95c7a5ea9b7addb83c77
zf6e5a4b7d7697645efe10d70b8c7644482f4859ad5346f18c033015f469a395dbcb9576fa5264f
z87476fa991d9fcecd3e43e0acf889770eef8898edb81857ad1b9485f7d851b4bc63542b5929f6e
zbd904c9a9b5ef3fb6782d99fee1c7c6ecf9bbc05239f61c67f78324860bd8eed0eaad947bd91f8
z35cb261a29001a79daf4672581c4376cdc2cbbb844e4fd4898dbef541307299caed40c1cab275a
z3166fb8f3557a134c829f465616e348c016a5271bebfc56de12d29cec15732f337803d6258f653
zc9caf30e23a673f125709e3982acc78f2f326434a32e30bbc6808ea4146e4e16eeb8fa82f9edb4
z8413243d8937611a711877f88e815c783253b580ad7260df0f09a241db91778b1554f6b162edcf
z27e483a8402a5975b4f19a86da2291ab80f2fa280239dfb8cd149cbc87c3e4565e93cae8fc41ce
z39cf2fc5446b62097aa09bbce66d5ded5d8f57853cd020cc3046789cd684225a5f3d75621ffb16
zb60d49a691d875877628861553e9ffb13d75500c0854669edc888000835f0c69be71d7b7196a2f
z9fb55da8d3afa003491ab51904cc71d4deb309ab3a4093e162a16843c80be25988e72d2e6d79ae
z06fe6e66d5e7eebcd6b9b5f754e97e95cac9efb2b86ef31d33b92482f2139b2a6865963339367e
zd3f002ce3180402f4edcbe24c1903b4b0ba616b25235f0e8921153fa07c856c04eeb577d85f69a
z7fcceced4c4389c9120f9c21b3e72dc1ae784d6ad63558ab83fa36442b6cd9f20f186b5d8884a3
z30ee0fe9c9b96cef6401abce32097b1bc709e928a9ff252e8722d6d92bbe50ab9674afe679c496
ze3c4c8a5ab8b817c7411ba93a048b6807b6bc613d4df1df59f82973332b2370decc1b4a476e46b
zabeeff6568c58ea2841702f081e40b17a5850753de10f68bee6fd4430c0fad757ce579256c7e36
zfa8921ac5ff4688c453724d1ab39dbbf7a2741d0f249c54cc9414a0d0ea870d53e2fbbadd3adbf
zd6dfdae730f4feef304d1ccc680165e18c6a44f2588eacc4bad8eecaaa7b94e70e1fcf012d79b9
zc2e2ff7105958e2e40dd1c868cdbe227b84877d3859feca9a7dcd3bd1d8e84f7534557a1684dd7
z4ad2be594e24d626955145fc0fcf3b095fe087fc0d722dfa8657648d3b66d66871044ff0681967
z7d428d9b1e39ecff61459d1620463fa506aad233e9e28d4211c58dc4400d9ee2bbe4dd2cf98e49
ze24843db283d0719db8a9b299c45ed417e1aa889e35d6ed0a8916a14b4bc094224daef371fa916
za5101b4808cfeb19f733446ce05144d839ee45e3917efca2f4cf2ec731808048b4371ef47b3d6c
z15b4451eb8a8456a6455110f907365e0b4e4990308138df1c69912ddbd37a17577870d07d90e05
z1109ac4fcb08f8ea2858de50f8da4f71a736ca763db91813ec0ed739c79adad8eeb8e5438fb0a0
z8b4bf34b35710fe2df7323efe78d37ac8c258b31546c0ca9819cd27c913306cd6073dd9511c993
z2824b7abdfe1865e3786c1b0513d2b08bb3261f002fae054f2f8fbec621c90e4e9d9e8ad1a0436
zff9056b0cf9836a7a88a1c35676f4b9139df56bbf0f821edbdcf5d50117a672422098c853ce713
z4fecf26a2cda7cb372ae3db96b6a1268a053fb6332d5c29741691b75855a2bdd554b7041e9e587
zcb5fce1b9bf5cff4c467460e5ca0edb24d53729b026ed2db0c88fd8c96aff0743c0989c7574d72
z38519b8c26642e04a26f91a1af3e57dc2c7f9127856db6cefbfe196e4fc265a9933dfee918e442
z9334c51d99f274701ed79cb66b7f959b72c14d101535afaf934b6a21c5357d6848782832bdbbdd
z0a20083892dd2391021c6caf9e19b2217471b633fdfa8be3604d6592f866ba3a98109964429c23
z65abb772d0074209fdfccdf91b2dd47e62ff14bb407ad328f81bdf96651426cbcf4f51fcd6bfbf
z33b6fa61b091e16c5b935b15bd9fc4a0c877c4aab3fc796aceafa01e9bda678da8900153b5fe7e
zac90ccac38e358d93b368aa62b31b0b9b4700d47235f1b4c2fa8fbac17214f0783588db1043c44
z9f29981f40c1af0a4dc5a5b5c6eca29641d416deb2a92be4751b9f0cea3c0b58526ccf4f4ae8f4
z2c5ccd6f85bfc32641f95925ba02826017033c26668a239caf82a8612906e9a024f7c0f904b5b1
z321a81e7f83c4c656506f6e1795eab37e8537c669ddf47b300818f9e15fb686e0708ae9cbf2da1
z0ed92391b4d8bd2d1e6d2b10bfd4c30db6f81bbabc0bb175a44278c41884ded24317ae1736caf2
z1bc6ab26b3cedf317e4e59e043bc46460a4b0b63b8ce8d3170ba9c201d1c3167ebdf79234130aa
zffb4985940c5ff2a26bfdbb05fafef1428353a5f52ca77a718995e63a32142f0d8dd2c87b1cc05
z039efdf3b6cedce27c158f1f91958ce8fb1cb43c89a43c395988dd0ecebb9b5acf41ecfe26a4a7
z73759f578dbb7b835c9170c0d110f5c4c555d92036deb1dd8c5dff012d7542c393480fa4ee803f
zc0275e3c0b976204e6ec21a04d5a0d24922024e057f26e44c338e160bc51e95f1ca9827879d974
zf720fed861504cfd4b30d87291f86f691c592f7342e26538cdfdde8bec91a528fcae2fe8e2c71c
zddf8f0554294562866f95b3be0ca7218dab69818488195dfa81c0638e5279466ae2b347170c6a2
zb3467cb80c7af04ca049de3517b12357b89e755e392f1cc54dfd0666b182b813ce7e9a7c61e9f6
zc187c69d5683af17a215adf3fa06886dd75590a6def3a8eab6f818aa232937c3557c521dc36363
z5df0ecc4330efc6ecaf58b3499c0e1459552a47de781cc3e969e14fd17706434f29c0434a12f52
za2fa05fdf0823e32590abed8c0fb133740b67228d66b554a1f1db05e22bac61cb65e1c361cefeb
z3be99afb203dba11cd3a7d857e34afb8ebfedef245dfbe4546082b35f94c12f2f1f4476995a47a
z7ef73b86044dfaf39f40f8cb03dc864df45a33b6a4a5ae4f6eed8714ade216eefa9fb275d32b97
z4de990be5252e49659e1556e7a2ccf76cde1b3d9808d5b2c342d9a362fc2c76bf14e3cc32da000
z18007a995ae4ddbf1973093da2714d68f5f840bb31d85ffccf78dd202fd068e22f141b90b957a4
z956eacbc77f8e9c8eceea5d29229c69d527c0c53d2e1d947ac8c99a392e8e5e37fa08a0a1f38e2
z1588e1ee9c0c3b22cfc3a2fdfc898bbd99d7594d0b340b83b3acb6c4e757a20c6f88bec07adb05
z326f198a15a8bf5099ff5d1d83a68473d13508aa354dbf12df666fbcef3bb6f7ed5d9c6679abe7
z75e53689de7348ae10615b62d7a36ec5f1535ecb5c7dc630226dca47b08f0f2f0e9b0a81919fe2
zf1a37c63175759529f638d66fad69d6f25c9b73c9b27897f2a9dbaaf80c75cadc2965cd25d5bfe
z6d8b1cd94e2cc8eb9cff512cb15798fcbfe398a1f7fcf5375ebcd841b66873eef1a96d396188f0
z5bc6758cf94ef5965b1aa3cec07bbd203aa523f052ff7d452b768324107c951a53107115527eab
za5d5d8a3af8253ba70c47fc9572ef02486e20af35d3183eebf866e10fae6457b4ac291f2caba16
z193d6fa0887f89516b0771baea5cd4e495edf1496815adca563f87a1f56225986e1e5003ce3195
z84974e9326c460da5eed7fbde70ec7417f448ddb4c34144f24833f0a3b00e4d5d67971861d003f
z2a08d16e802e4c6cc2cb0d57cb16a13f3e8c93fb1377b2f64f3626b9ae2d44aa86d27c9a59f100
z844714c3cea3e790aa8584a0d124d019dd199a7b3f71249497f90f5d929d40a25b3b8f24fbdde7
z70dd530dc594124df915293619b417ab06999f36b795523392269ac11a23e2ee8fabf37439312e
zaf5a81cd94a327b7316e5ca59c216341bc4bab88d24c443917d45c7cc2f5e3e76784e2135deb39
z1961a1c7a3c5aa212c0e896acb075d01d41456c20ecb3d4761403a37d4455e87d08f2f4a2bbcfa
ze220ace70ccb3f2b583cb644d292edb9c05443bcea8c02ea9115fa4da5dde2863c9c92c272db9e
z7405ed78291a4f453da710146bad51f20185d537a813ffef49f77d879f3610888aa4e3bb9928b9
z8c39e72f9b777511761486a856c7d4234e4e469509215890293d1489aa702f9ccf733529470e22
za97064a6b1c846842b7f78b1fa9dd9576ffe14f45478ef76c94d7d3ae04a57333505406e0b7b82
zf8b7710c387eb0d11f935c639db1609ec3d26caf11ba389dd3c7b5b0877fab6db92dc0531ad569
z415c9bc938e2aec20b5b1c741f9b945c34da6332d6e998f301156b27487adfeae8ac7e99df092a
z7852c380d7b0a7309878ff3497277a5c63dc9b090cead3ba2c50810867b1d9630e1778f8141568
z41f915e554cd8d158f01b4ac0618db49149dc4c60e08a910aea8c69b95b2455c9740ef51ecdbc3
zcfa6241f51e2b17ce8eb83881074d9102581d519a7003812fed9fa63e72ade6c7d5e6963f424ac
zb95da8a05890ae508d4ca4e37502cf235c3a40a6bd35157ab9dca39c5fe732ede19a0bcf793203
z95b67e136ee2a33ddef2ff24212a70be32e53c7740e8e5c6b7072427f7583dde237ce09762e87b
zd264deb16330660f387f854f8680de3d2ead901172ed8f6a94d0ef5186c008acabc89362a4368c
z0bf89ee367993898907a7631a2ec323f4ba5e39ebaf5edfd84883ddb874f475cba664b00b31426
z2b2a90ccd3054403ecbc71693f4bd79b661165526c951d92420bd98da9424bda74e977d5861142
zee76abe00bc66e024423a2f3ce107968bcc492c80920f9dd784d36020bfa49a56b685a8e6d6a50
z25c7509eca7d2a954e51dec54dc3453d0ef1296ea18eedff5feadf484004dc8ffdca44d4bda58f
z9b72d771ff9243bcff77066c6192041b9f13351b29943dd31f7d6c3ef6532498618c03b0332f33
z04fcc8cfa38aa1c5bdb2600eb3793c0bc640476e82839a3e85fb25981b44b6428d1a9ed4fb657f
zba4539bdad5712a3005329665b5b607748a664aa5fae124970f0a8032f76b59a77e2c76eba6d1d
zcae579392706971cbca91a62272ae9b58ce94972e443e0831a28d494c56c1a57e33fb726e442b6
z6b84fb6eea38aacb1099ecbc8c701ce3ec4ce0dd5a58dfc5f0eed02de0033d3d63d0ed632fa4cf
z5f906c1761aad1ef955d0644010401f9e493de2115346bb0e850a3ef559e70ffa459209398624a
za273a3cce49a563637a150b73cff6fa34880f1a899532dc715c3e30475a3c8d05df3db262408ca
z3d815b02de65238506fbb88e8b5b6c4ebd3fd34e1424e11d662bd519800a5a933a7ecd8c4e6329
z428ed4a7325d73bce54dd49173746b6dea37dc55b4ae959f1ef1a2dff061e9bdd113eec29baefd
zc3ec908923d040591a3cc37b4c28c27322b9fbab20a16ab9fbe4a201558824236bfc9fd41a8433
z880cf622486b82002ada0587b7b1c46ddb83c72a644c3b58c8271d645ce4a96a77d68e2ca3ecf4
zb5e0a03b085b96798769aa92ace0ad7cf255fa278015e60597c9f28f0d45d1135d2550dccce5b5
z0df60c21cc4a856f045f3a971b207884e921949bd430b91b6eeca90c4b9c0db0d1073a2fcd33aa
z3b3822685d67a198aa62f49e09628bdd8a6b034ff4451f48aea4bc2764bb43871c1a13ca9e4b45
z3c750cdeaf31ac76d268a26330fb48bd58cc4e81949f46778fb7af101719f020a711310b42da6e
zfbf2319ef8be544a0b147577f671d6eabd59ae64de14397cb65455a383573903d70072d1bf6ef0
z6fe6324ae71ef9fbb48efefea79f051a4d8b012a13d358cfc51a7c56bbc6cec1472b9aca221220
z44efd77bd1f97ab355abb9507d2575e79412bc5be06f62e5c35ac75c33a928503b4a0b9e8cea66
z46d6dc3a3c07e73982a7ea95af484ce475f9dc6582b5195b5151e76438d531efca38891a23d158
zade4ce4fab4c9021eeed2229cb487a94c3240fda958c0b2057743e047c7428876556fda8aa8266
zc5ce1603acf98110db5745d714e14d29beb8d45298aea999335b06ad7262d13455d7dff42038c3
z5cc3f4ae4c977f69784bf8a149666a9e6cc4925b549dbc9193195c01dc660c8eb3314ff02d371f
zb2a55e51414b5b9cbae21554e7ebf50f078e1be20fbbc0060ffb046ef36ae97a3a79290e544be3
zf7b15dff290145ff050a8abf68ee4cd98f26b94313fd218be2b528326b4573c6dabd8d0169f97b
zaae5dae1215798fe27abd1521e971a15fa752d3f4a02717d7fe43d62084c61d63090c6ab04616d
zabaa78a839873fed121f99f6908034f991a47a5394ed9be1d63b2f62724084d1ae835137b35e0f
z9b383375b8a3a207b5d0a478a1afff8acbb39680d907367baf81f2b61442e2b9eb032747b584f0
za46bcb130baca8b41fc65339a57f834224164e318fbde7fcd01daeee35c11ccf52ee54a7979d5f
zae9a7c7d1fa1af56e9a377b5d105e46adb056562a069007683491c07996a6de8d7a9705eb3d4a2
z4efd8bbe1ffa88cb3f07bbeaa9b1b8187b0a9b4c4da2564cca19c3a25ff877604f6d93cfe82424
z84992f96cd0e15f24aa44457512d66c32361cfe2cae7bcd963d8048b094b0c322baef568e74e9b
z118e11f7058d3d5db5acb3b98ee564b1008189e390a87b4c72fe21ca42c79ee54f1020e19f08d5
z4d981b4d42da44c284bfe37d187ad497cc29691a450b65a34dcb9a6fbf9b1f3a659bb8916f8dbe
z1a475121960449d52c51bdd6dad9e389ffa05df2767b8b05b63f358be0330a835f18971d018baa
z19b8f5db759ed28186566a2834aec77b5b96da6b4af97e1eae0b160d1859eb0275f6b905f074f4
zfee110586d7a9c1a1b603f611b2a52349cba7d3e2242e941e47f275cc2016416a604b8d13103c2
z95b95361a267bc9bd2979747dc828cdfc7b8fdba7a309b34e8f9475dc74d13b4f482f042335855
z4c609ebad2b8039b60f341f39c1f93cad5ed4e6903a8aee660f6e7c6a40a25b849685b7a340cc1
za09d3d4ee82fca3cb57a34d6f2992070fd263645a2d22a2562820a344691efed7b46ff4fa8e78a
zb7ad0a5311242353f1326f4afe269dfc319120910706e50665bfde0aa6115c8ae79c47d66e590e
z75d8e0f63b7fe87655c01a05d0e770eeb74c11777d955d10e8593cf27a38d6e42876b5f9b4f5ca
z94a40910cfb6afbf70bcb771845b7deea2302ddc49e8ac2642ec6dbf4a2f05e4ac8d5028045f36
z2e9c425f32fa450efebe321b512161d20e29baabca27b14539ebb1580524e35d88810272964bd0
z9f6b3569a0845bbed75b4b398b2a5c5a135df5d860c9e97833f095ef2b29a8dd722d58146bcd9b
z5e9d32e8eb6b71f556223794cca1dae779fcdf43b0750cb3ea56c360dd56e8574d85e3dd641856
z929b759c36a232ce7b0501af0f7075de2aba85f6089326546e243c5e3e99465eac7e44a8b2c2ed
z60583b8843eb9da22069e96bfd7345a4c98745259e667cb997925c397645c70e0ad5fc76aa9e2a
z8d127f5edaeb558fa4310aad507ae060f1d9d6e2501844a95618b3ea0a6b287a6acd2a545e810d
z5de6db7f645f212f1980702134683af039c0be41ac21d37179dd441777be020d7abbdc1fe988f2
z9d9b66103e897aa29e852a7f2885560422ef69eb94d052b2c2ae99b64a2ee9f4d53a1005e19147
z557dcbcb16475edd6caab967ee61c7a662e783f38fd633c988275dd3dd711d791090f00e666b0c
zb5dcb4e0f11f5504caf6bc815d5f82ad50cd8816d31934c0bd272e38a3979448bea034fe79010c
z112f475a534a0eb8d1ae73eae3ef56f43292750f6aca35d09e72795fb2e53aef4a5abf4dc6e71b
zdccce1e82029a08e92dab00259add82b1055b954aa60f16abc14db81b525b69baedaff1fe5d50d
z94da36a37c7a17c82980520c125f18cecb080bebe1683976ca87368d625bac2af2a52aa1796411
zc7d0c27184dc44ff089abc434ad215cbdb029c9ff0dc7f5d09645078dde287e41f5224d5c326cf
zc7c386d42a8c0b22875d4f4920b426f1794d81caef5ec5c29b3d27304bc8c2872c3b560bd9084b
z4a9cc29a91a16f1ca4ab31679007fbfa73a53ccac9dc5a68a9c8af9230d502df82ee79634cc6ca
zaf749f5b0aefd264355b1adabc00f3592b3e935797168adc95ccd529ea335c5134baf40a2a3c3c
zb09fee4799e33ae22ce924dab36ff0cf0a340c6adcd1a68a5f93733baca243f001970be675f200
zb1a933d85f6a94526edae8360facba6346c872becf2fb3bf8753129bac255cb6e2a028f97c84e2
z3a8b857f6130033bf82d86d3ec15ff9f7c605c9dde22bea9d05abcb4d42d0f0644dac7efe11bb2
z57e5b278e1ec5d70e4ee7313f95f6bf1dceaa49b8496626b3ac721a743e2beaa9029ef189d28bd
zc3c0cb6fc914cd41c4e382700924bb1ee4b23a0066e8c5be330a5a4cca3e150e75e9e9a2e66dc0
zee8c336686c6ae2cf2fcba95d7d3301bf5d749c48893d9bb1d03542b35754099111a4a81cc4a15
z9f7e91a6b5666f8de4f18daccde49ff62134562bc4f508502b9e2dafd1f8b36721b6c4a0549dca
z2f85b10d33a785f8e1ec8bb17d47ecc03c859ca226a328908c8954eda655b7bc14eda4376bb18e
z33524588e68be40aff5fa91cf19837a82189136fca670e24c634befd1875c85df0012a4ff2df9a
z30935cebf138a48af6b6c86992bc7227d901e60a4879b2b56d7ff60b98b7a6f45540abfecc7216
z17fce7f388da8aeff916cd1336031005b885b3fb83017eb3e214bd48c32418545b9fd0e52451e8
zb06210909370ff043e592d9d0b790b1090a1bfdf7e984a869a2a74f4d62a3f0d245d2c6caedfe7
zc692d0cc86f9d4fda81e6a8feb25ceb6114e20792e232c66836ac9c3a347c79b5d67decdeeb38a
zce709a9cf2d26a6816d36144f85eadfde627fd64fcf423961edbc29104c91a8c58ae3046daf1c2
z9626ff0ca4fb0ce33cabe6452ab19695a420a2c6a9fbfbe99b94f014615a9091ecde01d812c918
z98fd7d10eaebe2d4c9c4c29f3de62aee162144df1bf148cc78f2d6e089bd63bb043dc836ece872
za07470426b295f9eb0a1640db1e25daebb41e0e240c401c0b15d34326053ca27ddcc1661572ca6
z0655cbcc677426ebb580bb2a6a78a5b8d8eb2cbcb83b87b7fba2130767d7228de85e39426bfb72
z7a81c425bbf1c2d837632d75902aad95521699a0b0e7924b1e0f86d429160eae414901f2f93289
z32dbe00772322e5db9c6f87e5db66b453159f96fe67609532adfe8104cb9a3c06c9c1ba535eea6
zec7bb049af81e7075d42522bd9b7603a082ee47bb612966a88ae056068be96bc8ae154ba2c4120
z7f0c2555f4806de43f3806fe0594a508694a9b0bd91ee05826e29305063e9d8e37d1fb321d0a42
z861d6fd4cc604a0290dd98104cc1809532a4d2a3a32e4366b1e156e9b429ff02770b8c63a85c7d
z94a360b9aa20fc3ab1eb900b49fe35485a510bae16b2c1324077e057532024410560884a4be4ee
z163e3c9231f5f6f9cf22e1d409a68f9d01e1a5585d0f3c05408f3db739f0cb4e2d9cde04f51da8
z91af0d0304e225882758467e90532220eea8bec34cdd2afc396c0a9e8f8d340d20fac3ac22f49c
zc5ce1539a27e8a98ce2b81e6fd3383903ea18348c5cc3182cf1271f36703e0bd144491692ecb68
z88a4e0b5c02df5a6547d5b11c6f6f4aaaf2af07b47b0c7a7d975e14ffa2f59c48d5b9e34d5427d
zc92825b4c2f7ebe2014d69f2df36681a193194a7f45012dbfcc4d71d9d09f8a9b2da31ed89fdd6
z46f4ff90e755508c971f87aae2ab1f9792cbe3f15a9f7e4895caad917d9d0f2bc8c9228d3852bb
z2844ebe91a9dc5660f103d657b94767c61f7fa5ce6965de99b71d6a320caa9cea9d2aeca2ec16e
z176c206355d1140c0428e9bb96c929c4daa0a09c17ea396ae20285ae667f4d549cad01a6041e10
z7a51100530eead3fc569ec79238c605efbdcf1eddc08ebe9e8b2511c9716b8ba3938e565ab13ea
zcf671a5cdfe73c3c0d739061f4c82411e184aeeeb3a5f66834d4ffff8d98424cc0329c361136ee
z1733b0c137f447297e7c31bd794cb2fd3f3d4544e03d2675967024da967f925f3a2df435127aa4
z49be021a24414b56c1bf41e01d734c7d483b41ebddfc4da10ad5d1233ade492b24c0d7f9ebd39a
z41679b92c319070581a155ae95065a8ad970b763d17c8a8e24c83e0248aec61fa61e8bdee71850
z29a750631644b2e22d6f28010a0961c6ba73323b5d15adf90a7222b189a48a44587665c3a388be
zdd8827aa316ad5f33d2fe5f05082441bb7eaba7f21f78a3ff55a92133b5ce0e63e54cf85e44431
zad20c558a73dd82fff503fa04da6ceff2b19f40163abade6867f8e39352a1a000149ec16072c35
z87b4dd56716975f322c0e430fea992f892077aea5029e62b0959e1d124ec234f1e5c7cfdd8599f
zad361ac8b409154d27290290a8614bc64e218d3f4fa765641bd43b7d520beb81b8fae44f029eba
z4ca7418861090c340b7e696199b4d6977bc948c4306c742ee3fee951c90b3ba19525087744ee72
zafabf84b00ea6f4ff7762a403fa9a840114fd18457d1356fb37dd41a3d9da532e17d3636a78a4b
z4a5dc58a625493c5a3e69bfc128535ed408f5f4050d2718d27a22325b99b6977a04e60cff85977
z25af07c61a7cdeb094ffaafd5722b2a36d789efed10eaed6687289ac932dcfc7aa04c97eb61f19
zbec8a5cfbf7fa4e63febd88e1813c5457d241da2dd19459e28aade05d5dc031ad6e92567eafcd7
zbb19f725a75cebbd3c160fee50aaf631a0fe4ee23975d6e21571269b1c67c919e7876820e14860
z1ec28d5cfbcabcfbac73787363574b8ad242790361ffd368b745a9861074e62e41e079d07d9d05
z5d44fb356cd5f1baa83129f1aff56ca1f462189a94d77efecc54e3179c03929b6e2fa62111123f
z2d58e082f7064573c0c9854c6682be53bfd767c187f014bcaefda81f880529eef3e7e07c643bd1
zc2183bd97b3c1edbcc85ef56598856ebdaedc82bf7fcb7a5167fe7881a189300a422cd8a672c29
za98ab20963bbed8f8631f1faa55ae494372d3464fe20915856560206bfdca432a8b422931561f3
z0a4640335ddb3d68057aa569bf156ff70e5d6219c71aeff366f3d7339dcc4e60c68271d4447357
z66d68a6341b4c3d6a43d0640fb4fcdd66a0fa9c363bf67b88de442be8bbf2805685b83d886477f
z5c03a7ff56a48c9c5126d6560c6ebd87f03e231721b16d4709b3714543b776ff2311b414ee3fea
z438407b5316afa98ccf24becdf8bcbad4f757e85c262c98de5d94bd0f1a3add37853c48d5326a0
z1afe10141b5640ebc45087b6ad7b2585880dce744beaa3b42b6d5661440bc38f613ad31b41ef8f
zf3d3dd6733cbf8973a897625c6a7eeeb4c1eb8d2858086c8bd5d1df2abe151a74ed12385d9e900
z9a8f504a648510c9db9acae7ef72514b1a02b3c090262406ca1a0971384d4e2b54613dc8ac106c
z13113f048e046cbd5554d388556c4cd945475b4d5142d110d6b817326d57c9729c940495704409
z6c62c29d724655ac6039bf2b97c8fe1f483ac617a62ac4d475d2d59f7baea7921d1c3cda796963
z2879e128c0357b07e2157b4dc2c747820db70c6c566ddf49a3da668f3ac4d7ef06ddc38f700440
z068b997e88d8de0f2e7d96b2413d039b9825e6cb22ab7e19130b5ddb565fdd20b92287b5e07c9e
z4179aebdb95424cecc3aed216a913e8c3e979b53addb977fd26b5eeab12e162e0ce9df847bb16a
z7683faa1b2b30ab5174a51a4fd29780e5f3f16ce9fdc814fb606d5f6d0cea8b037c464efb3bbbb
zd6198b9fc3f7f941ea6ac6d275e40977cc2c09495b012a1a0db2cf0662f06c73b4ad0b5c50d3ed
z96fc2cc9199e7e0e9e144131168381cf9bb5d18451b9a526dd9ae36f31499444429055ae4d272a
z6ec2342d96b0b9ec6e6668bce3c43d7e5609e93a9625790f2ef9d9ced9e4677ba0216886423b5d
z60965aec5d1caa097955bd43b7659e0a354e75d1e4d989bd99052b00a391cb4c35d7bfacd4d8ab
z1ecba9906747f24811a6e01d1a60064dca0dab28c4095615fd15e042fc154ceb34d1243576bae0
z7795cc8b384c58e4eba5430f57ece952a2f4f6b02e7f360e001d89983f2bc4628d3d7df5d10ed2
z767120c86d3dd43dc7f26ef8664bb1d2ace2bb6fade8081d118c7bee69cf7b5402822bba279e58
z542bcc63726f221c8864258337d9e2b681abd727e34502132e9e7623a8877c59aa830f4096535f
zaa22195e64eae0d7c25f43ee88025d4daf81417088d4537799614e20de2cb3e73702a18ab8b5b5
zb6195a70a11c291e4852c1a38c700298048487443c4181ef8e2c0d54950702e181e48df5cf1a75
z330ec3ca95cc74c28942540229e7d468a32532f81a8f126552ac95b01fd33c76c2619068108224
z59bde30e670e2eeeed644b68ee9d892580d2b3b632951ed6949eb4d94acb9139bd81f056f47c3e
zf552438dba574b26ce25322a569e1f492b7eb9714c0a7a8ab1f40dcc3f7c6a9870adb6e899ae3b
z4717a5c4ee82cff63f2b60ff4312756851a0d90f1ec5450658b7345d8ce543be913ad1ee980776
z69ae02c26bdafae58ca293550ebf4f196558d66e160a6a0d3cfd3322c223b7ba210c6c271f5cf9
ze43196d4f011b3d89b00d0123b577bef3b4a58939cd8909da99694dc95f5b13e123b408d158bd1
zefe7189fa23c7c6ec0c33ccdabedeedfed08faf9d9a8aab58738a0f4f37759544efccddf117f70
z0888b05ddb2414feac0db25ccffb15106be84912b4e63971dde486c480adb2ff505f266e2a8aa6
zfaedfa739dc03a9daeeb548ae14ef9653ef0417bb27fb1094ac01fda9b8f31ffd09f5d79a0c363
zba7038520a310d8a79b6154fb8e081ce10c5dfb5d8c53d33f2c5e5d85cd6df9ce1e749d955b578
zb721cbb8fff20978a8db7a55b2e688a8184750ef658250100eadbfc78624c1d92529da3f99e81d
zb7ceb1335f1d60d142980615a1b7084a14d31f7deddcc475ae0e302c8b6cd5129735c527ee5d86
z6839b935236c210f5b48e3d579ed770b527022ab80da0e3329ade3d11884402d129051c41b3387
ze1a098bf10e3b03cce1985b55484359b873f58fc2433486a815876f14e38bc368568609514c769
z7b22c1982da2ed68b0c5616c8712ada61b9506b0d0a65e96381d0590882bf236accdb8b10984c4
zfa685ce6f5acea6309c5811b1de58c2784ed8064fa9886375289774646d49ab55bbee5986e8973
zde91b9096ae9860d84a1a193e81821b9e9e00ad2c7807079a3c6a5d8a9c9b7cb8804278c5987ab
z8001ff353cb0c93499e180e58d9c73df31182e6130c4274c9d58e784add8051a7bfc574584e121
zc1e74c29eedc72c1c121ac94123d836549b6815b9f416aa4e8380d1d00f09878b0f9f0a53bb2d2
zd9d5cc6b2e3b805e07915851e4881b32ad4f9563c27acc72e8455294df0f04bd197e148f0cf423
z3a5371d91fbcb1cb089f37a7abd1ed6424b8cc0851db5ba8896cf03b1a5088a410c83a4ec9734e
zcea617d4f91f5e1c0f28229472a64d0847e2e45e9cdc15047ef2d56db817b2c9cb58f3f3573eea
z838c41c00fe2cdd2a17c637855765d90d3b40021d7a8747b7424706faba80a9e36e4941c146af3
z5e7590897ea5b5ef34f78fe19d712754d99caad41072e0d07cc8d4fb95aa8e8e6d535fd0afa4d7
zf180521ccfe5842f6a6eb73bfc2e5372101b54bd535a70fffc3580a7bc2028d54a01cb1c950af5
z95cbf91b2fa913655b1695fc0452ce7695247a0e23e0062d0876048c538c38f08bae06397d875d
z1aa727abfe475e4190e2560eb39be6cdafe067bc334508a6009a1bdd9c8e33a221ea8338803759
zfe89f72239889849f232efef8c9bb3a76fc02b34f5a99b5ee62f448ede7f6f1aac8f2ab4b8d08e
z86de31364efe4b0db471e17542d895d7f108c0dea97adc14ec6d1f91a197ecb6decd2fa096a845
zd467321a196b8e63beb3192cfbebbe67df80c6e37fd1dbd305863c607e981aec90f8f0eacdbc53
z4fde09ba10c2093f7436b167fdb4cb77a7ec177d4b3580292ea846a4779e51acf6a35ad81cb4eb
zd32f426a1ae4e5dd7a39cb623f1421d87e77e5c166fc0a53e76febcdd22a4fe0a5d8daf0b29fd8
z5ac6308b198123beb24171c0eb38b2ad4b7552edb709bbf1ed76e64b1f76e8594dda5ca8e987b2
zd7d3d97c54eae688c511674a70c78459499da49454624dbd724d20b32c8be7ea2fad04513fb372
z690eb0f15ab513b332ed4a7e1ae0267d32846edc4b8db1f62475c116f409b4ec797fe93cccc019
zf37f9ff476ed21966db88a16b43ea1c2b4d8070f13afc9db64c8755bf3c398b7d8c25bab2699bf
z286887abe73f05ce1e5a1551ee1df22f8750aeb9bfc04712a0c639d94e3c5b6209e788c1ad94a3
ze47034b1d2822ce6cc06f3664d73c12539385a30d9d2d518faf7fa44e43c6028612fe97374e2d8
z119ef5ef112ad2b226f5a636ff30e3ff80e71331797d0c2db78bc2bda29420983a4aedf1cdf0b0
zb8242a3df97b7d23f8af093668f0cc53d437d6fe51a48bb9a67788c02b7908f388caf20e287409
z2f7ad0ac0c0c5c9d0b0ef446f6b02f373431ed9d910e54954576cdc04647858b736a13455523e6
zdfeaf56b38328484cdad422f458468c78aee5884cab3dd7c4e8dd333a5d18e0abd3b2c187a840f
z66cbb17810d412b1ee28fe2a7e67393ae456e1ce66d5073c5b9385accc2d16c17256d77fde970c
z4fe902bc7143020fb885ef005449d29029fa67c64a9242fbca15b62130b50f40d844fd70ddf93b
zbd32ec5775a4f80c60ab83255df4f186d6c11bc458095f09af5e7109fbe7854f54d1126f6dcd2d
zc14d4bedcff6142601fcbeaf75fb1127f57452fce61b4bd012a98b30d8d9f2e6edbbb7938c03a7
z317bfbc5cf779f5146605f00a85ce15dc42d025c3ce3d5ef6fe745ba6f37d46daa5f768d410da2
z20854282cd347d051f7e2f8ce7f128dc3c06a6086c0fd5470eba04aa8b2816498d242c899a75e4
zacf286de184aa2b459183c23d1c1eaa66b50048752af293416dc841ed92aed306d90be7a587046
ze3003f7c9b9794d0923c51f57749a90566c73faf34947d37f6e737999fe8fce6e31b9fe9648372
z86be4cacf26c8d0b92df943eef159e8f97caa3c9bc4c9786c4089c5fc057fb2d8674a1f388dede
z3b670c353a229d2cf80c4de930bdd87984b18f5ee25e974ef432cbc3c3d21dc689d41f506241b3
zb58cce4b0bab18c56fdaa258e30f5f731ebd51a53e1687428482778f64991887697150954896d8
z9376759b70adc60f8221d68a98b9cb71f38becd47d8472bb4f080b0aa7b349c80adf5a37636eb3
z680a550c797a11fb46106345169a6aeaeb5aa0d706093b8b8d7b6864725697683b55641282f1dd
z75a3498fae73a1c508fe09d780478cfbe1405382a94820358b72edae1b2cfeff4ef8d01c776ad3
z220459a55dab1a3f5b73b14957fad657f624aaa405b4a69c68db955c4556f76e49dc720a737ecf
zb32a8720c3eb3b904ea819494f6fb8874a52cbcda57bce3144e7ce8fabc543bec93022563fa52f
zbbc087e206a4778c411a85f70bfed5c8b5a3e954ffbf28300c8e61dc42c3262167453306b5c99c
zaac70d9a01dbb0db45d371f34be5f5c5f6e8e5945dfabdf67e8c9a565d3361df6778eae7118b0f
z45525695fea6fd95bfa85015ea8ff764392034fe6b9fd966d79bbc24cbdceb27910f24ac520efe
z647299824edd22bf5c1179167b3fb11516568e40f4438dd46304b9eb2b7d26e4e03738a6638107
z30fdb8da0f6662f52d3a1fd24ace2017d9ba43750097e89d1275a82eeca8188cbe2ed0087be6f0
z0c8678c2e90e8986d81218eef3e36af6a7d92e70678e15a2fda44c0dd3a4ff2dc14904ea17edf5
z7400afbd5df2edec6b9467947fd3aed8dad8277609d9cecca627c7ed0755ceb9eb70324e63c4ed
zd0607aa9372bfb389f8f19563934ac3c9cb6d1f7195e00b7a276f4e74c768a69dfb831116a8bd2
z303f2a3498bfed8d9820a03e9f847a006d32308b95e5e5315e1b7431366eba1f4d2d2737b7583b
z843a247fe79898a0a5a9ee0308b4b453fad6612604e320a6c63b698cc903771a1bd30e57637111
z1a8da59649210e1d3f3f3554fdf5a0a3e08c51195f4d88abd0ff4e428e9c22e9d2e30e1c3bd8ff
z41eeba20291104b9b3a69a9b87202dab1c781eeccf64788cebea6f096448c0e0976e1fa3a69de6
zc55f5a5532fc9b27ac26f1fa7139de9fe001b39c1a6139b49d1d64ebe8fe06ec10abfcb6d08602
zfe5104260e7e6cfc9dcf4c6eef1965858fe9f8393830b1157b565cf38ad7d8c0be16001ae24b90
zb005ea7bf9c881f1807b2b47c0d9d5f1bcc622a59aaf48326baf2bd3ad88d8a698e4c610815a8c
z7611906a5c586af7880c93a5273e2500275b35933c8d386696f43af77fa0ee1f654ab1c53f0dbf
zb0ffbd810258b7913508037063d613560212aeb3073ddf21084b747f41237613f9a9a941ea853d
z92f96e7eb88fe9f57805ec2a4772f94affda24032009b8f4dcfdbe65ef386aa3f78f306c79c636
zdbd5d6693ac96f52fdd90f7be28f14f6dd861120ca768fa93e2830936895e52a17a51531ebbbe7
z4387cb28862a0af82f4bc709fd290b2e5a4bc2ab4bce97fb098e498da05c52e82c9b834ef31dcd
z6193cd487c87519418b68d65ceeec5bb2fec195ec5bd9d51f3434d09af292fa23042a4185bfe5c
z69c7a489dca81a1c497575e2f7a1f483bb4c388415ee593d99e0cde0f48d47e5e01dc1360debda
ze2d4556790d3053fc318dd09dac0801d5a5a198844f036bf9bd10be7883a71b670aeae3ca0bb26
zc974e3041fd21c2261adca895c2215718c5b7b86d29a141a61dc13ef483ca75d1998ad702dc7ad
zb4d441e952220a9d8f376b49a4427c099b60346a872dbd5fdbcea22468668aaf1abfcc05871f2b
zf4e56d3d760628ff127eefb997210a80513bc4f7038837961b6246571c440bec4e3277a705175d
z6c7d77e1706d0ce9cbdf615df6341b3f5b27d224bf589c4eea490def4f4bd8daef11d587336660
z72cd0a217391412ab86d442e46e86f40b1f1e604a209e9eb1ff9842db31fd7f9e5b4f89564b3ef
z146ae834dd3087796193242503cbe147015f84d0d3c2bedc821a1d7caba4dddd925372f8450980
z42b55a1189143775a4a146f2b18fec5def865b960b7cb712a77099ee543d2fb1eecdda5a09a85d
zeab01887f2f4883fc054d2107771bdbb1fcf481761ae9a0aa9786feee1761f4e0b21755d48cbbc
z965dcca8af277aa0335094aa7ef146d2128bf66488db13dce19f98d81fe840ef281329d4531671
zbad20d981410ab19f0a157b233e05181f224facf04c22b40e5fbb15416d905f60c3ee7e66a57f4
z3794471ee1be24fd6603e54c6179001c1777b382918eabc57bc59222b0f8ca72a4da7373b155c2
zdf1963127ddc281f7e75c3290eb911efc22848ed246d9ef4317d15002805f4d06de7360540bd7a
zdc87163b35f3f4c49e9779ad730d4d88ac07ce4847757cbcc8714b054816cca9889ab5c0580c64
z3bee301d30eb62b8871dc7b11ad4e7b6af2ce80ba014b06781888e4a1d96a608e4861b9cb1f491
z7c8865332c60321d68471443496fb7e4a9080fbd20be3c1b8381b59b892e7dff50b2db0e0d763c
zba10188a86b2d2153b92af67103f69e213a9ca0cef036a2bd13206a2b4996e28f2efdb253402bd
zb7fda26afb80654da2f45b97b562cac4cd1b79ab06f8b0facf53bd41cb72e101a51baf2a37bcd2
z0832f0447795273b3540a41110a6b95d9acbb22a156fed66b9ee02d8cb458bef8a712d2616550d
z227c4884fc9b24f95ed4e751ef50095be093684552cae92f7900cdbad9bbf45d40962173aed4cb
ze9b6ee5eb13efacc3fee499e1eb7765bb9a1a43b941a6b0aae8ad91517c424611a6b07cb3ed755
z20e01265d13cb39ba98e5a7b09f5dc47d969838067c9fee7e6c06646847edaba12b7027c81f537
zf227b38518339916b11b907c66672f47f72fe08b318c6a2013b3c5935954301f0b2b939f7cc610
z91e19be58cccda5d3d8d099097766d0c36096888967838e79f2b6c876d0a49c2fd69fcf98a29c7
zd5e11a21d2c17bcc4fbd9350b21a4df983ec6b9c338f08e293a62d04480ac30c1b39da8dadf3bb
z696116258cd7528dc81588c16290082166246335e12c4717a6f57275b861a18a47ab90073218c0
zed57e1f520d8ccbd8514e1b5d87a130eea2e5fdb53e6de7c5c705136fbf39211c737470482eb11
za6b3cb396ca0565c10a4dd0bcd51747e86e418f2938809466eaa94ed1e46f6ae45f15201f0739e
z4b258b0bde6ec4776a3232ab41002ea82ddbe1e7b526cc5d730647c22a9bf455e936c68a20b018
zeb14c6a8a4b6a00ead2a255c873079193e9dbdad9207be39c1f16a7f2ed4bad8d22a39eeb43579
zd83dc399c904aa1c93372597500288d9aaf95c7d575a71b1f2a070c04187f3549bd45482815c64
zae13a0d333bfcdeeb4085a3cadfe458e53fd0d4ddf58c7b032502f10fa98c4f82543fbd8a4d8f6
zf7aaee6a0f87cb5e5cdd31f192fdaad48bcd0238f51694cdfcb9582cdd0a0b9b1aa50cdd424540
z0f3acedb2c8f0aa0bd42b7e1eed1354d7ec8125712f0e899411e6c326691b09b4ee070f75545ef
z028d563dd8feb13473b7231e46472af6687dadb020de3840911e5ddc5eaab42afca8c2d9e33c3a
zf2936836599fda1cef7ac8610c2315c82f50b155e38e89d51b2b3b7250ffe16d9f28a7cfa9aca8
z21d9b14bc615837737a88b5aa11141e4938eef8ddcb71c59e01020a8d61a39edaa832a319fe0ee
z39c753b4162d13b32ca76f9b27f2b83877ab5ad470af6cf3c4fb6adc083fcd6aa27a797d588d42
zab77503866f80026d0e22964297bfd46389a3584f18cb2aebd6d98172b24c07ae75da61116bbcb
zb725398ab531925566bcffd9da2b2f011e52b189641f4b8a31d9738ce2742591e1e2de900c7191
z3ef920bb802585351fdf92d4604ec4b27ffa7ca2fb7cca3e0b61fc298e798be0bc39131987c4b1
ze1a8c8cb57b89333180675e89424ff063a49fa081951152548dcdc47fbae74a33d39422fd42100
zd22826275ec681e69ec683c79b24185a945e38dca9520ae78b2e75f637dd329bb5271946978977
z6aaa7f323d5a2574b12378d276568bca438b1691ed65a8cab50a55e6479121a401faae86f5c50b
z77ba5cf64b30e7ffe1a504adeed2688bf858e2f325f4c766dfcc730f1a241b63db45bd53556ca0
z12e6dd907cbeaefdc50d26534380d60bb55edee75a32831934ad6f3e17dfc7a13784d44bfe4795
z22d42385cfbea0919dbbeb1cd55102415a127dd2e60c5db970720eda03307b7ec1e3b7a2edf86d
zacb80a7a0e32bc566167f2d95745b939ed035e95a33dfb4e01242c253455fcc29f084d4570e8dd
z5a24e5dfe78d49a210ba9e191f3831e845a3e0b3a161f55ec3022571bc8f9d59b4e783fbb24cd0
zc9123ccf50f544fa0e42ac52d2aec138a93ee79528633d45c318a215a78c9da14abd64cefca025
z6add839f1adf411b4b819a98b995432819974f3fb56c9202e2c08ef2b170ad217ec82b10c08fba
z9aba83df99eab9886c46e17fb7c4fb2bff37f0fe1fe7584b8248ca56cdc61882f0963683238d39
z92a1754da1d916030b3d5a14272971c5f2278d8818938686789491f14dbad4db855e85d5998862
zcfc1c9c22f0ae3c3ad7bf43ecd263b6711faf36111fc4795d23fa6f1a427d28ae2b4e852610764
zad8d994417961c93ca2e6f449daa5b8e80e3b0e76aea8229181f40ef0cd75848dd0b6c02e0f6c5
z74089f0694ad7470e5ea906bd0c01e8e727066db5eda1711f2d1369c36ac86b0a4482882b407fd
z5a1e7947d4de9785e75fe2938b9b8648fda21c5328bf8b3439be759df027ecc4cc4471ebf7b702
zc5df0336970000263e8dc05f5b8c476055e09c0facc65e6df0bff71080b01369b3c604a91e2c49
ze9df2f679e87cc3c0d68e2e3cf8fde69397a0e330798dd28aa37e9405b6cf7300ec4ba464bcb36
z6c9100a5680c1925e44f24e529a99f0f81701d7837f758bbcf5bc66c4fc597eab6d9a141f77f7b
zf9d3c53251af9c73e9d9492f2f679e304e1fea4c0bcc4ce11ccea2b7bb8f5449827c12d5cae3a3
z9ae224191802045aad8ebba319e2f55bf9680a9e8692c9b21a8572e66f56efc60790385672005b
zc61c7b311e1bb6cfbd24b8c4cafb980137a63fd00c63914649f3a89bb9c64902126d6ac97abe72
z92f5f93e48ca80c97c2fbfe3efe81bc95a44e68feb0e17f8dcf3caa22c05ecea97c2dbc53146b3
za0f98bd8ba4a8e04fbfcd460083a71c6f6c77f7a82f8cc3f900fdc4c0073155913c730d2980af4
z4a7cdba30fe081a63a4d64f251f70ab3b317480dab07191654c20485918766199495e581f10937
z7da34af7b292615dac9a06c55124aac4656d0a217d814c2e70096a1295801b6a8015b5646004c3
ze43f3266f015f28b657a2e5cc8ece86d822c6c7d67da8f68ba0427af116036bf013d2d7841a585
ze58b2eb492806545273b23224a42de8f82d7c9712425d1ad97c3827fad537c083e12a1fc852582
zdd147cdccc25236e6e65e09da457f9db091b89e0b8f3eccf33a5a793b0c7568bb0027064801af3
zbc27a6480a6633412ca568b0239baf6b6ba861de486323605bde314fa7266958950f54a2bb9238
z0f3d8b4250783d2d18f158db1a25f404d074374d51879113b9095e9992f7f4e286c9cdb88ef585
zb7b6003cfb482650447a2b3c7985f78ecca5a0e69a87e2f579f13dcf05b0ddbf1c23b6ef5ef0e6
zf8cd8f7e2b26b65539d72efd32e87732215256a7dff7135d83d4f06e2051f6d8284f89183fb519
z3b83ece6cf91ee65730b2e7c3bf885dd056142a5057f84ce13ec9fb54015056b403dc36a7281a2
z55979607d8f9cd803a04777ae0492aeba246bc64f577eff5d7ba6791302a961eb6215b88bafc54
z3919e2a6a2c3f8fbeff43639a4a3fbb082b5995e81e990fcee933008d480f33bf3fe14d07146fa
z7760934ba80ba85241010132fbc13b6b1bd43ddd5d93767c9bf71d5cf0f5737841a4a3d01a862f
ze02cb03faa110e0e0d2fcf1f229b404b58c951edfa207aad1cf340bdee80abc5d0fcdc82c63e2b
zb7bc4d65bf6a19580c9286df1e4038a03306a945889b3a18c46113d94cace2e94f4ee8d9f189f5
z91765ba8338968574cd4830a4966191995c6234f2be88dc13cab169dd3b29cf21a119e45360ece
z675c3110770d4ee484afc0a31e4f0da15a65b3c1f9b81bd4c24359a0a3a30a5367b5177daa5c36
za92cd249bc6e43956c08ff8c7c4b6ad014297e98a05c7659f0766831e088437a3c95419b2e5bf8
z5512da128efb8633759f484cb3172ce7041fad2305794328458c3a0ee25130540d80d837992388
zb74c0dc1b221a5a741464a9ca85ad7b3f1b98a240805c3dd6e1e5d873536a164e3cb05c6eb2edc
z01742738f5040074a82a4e47917e26f3dc37a633bbb99a4415a7c6cb727d7e5a5dcb81442375ee
z8bbd0bb984765f88ebf1827b4d0f333010d86b0e6602eb4d3a344a135eb8ecc771c9a13a701783
zcf042cb59dce75d20286ff4309898e56b357e8d524e620b268b2192d8a29db785a1c8269389453
zd7068fe1a56a1beb20d27078c1c0e0b85996d7eddca8c840ce494ffd566320176f5253e1eac7cc
z6fc9e62810b4e61fa9e7c3f83d6f8f0f836f68f7554aed7d7e66200dbcb9df8c0d535d8d2f6aa5
zfec4e18a3a70ef9e382b3fc275c9d98bb3df11e3b311c7322b2016b88ceb17926d8e79f6923d94
z78e92f6f66f6bdde5276a682c4d404a52950c94f28543b4add3dfd4c968dfe292dd2cb5cf82cd2
z3e6f1462bc92c00a0bd11a297b04e37fd43d617b1878296807d09caeaffcaf589f934dc1c0be4d
z41855357556410159994168b3b5e0abe11dd5934f65f05fa06b96e18424dc2541701a400af730b
z8f81937016dea4f042011deeb54ffec1c6cac9e744b65cf2d69f38795f4cb324b065e6ad8f388c
z407fe9b23ea6a8f8026ac7c7e484050540d2184f03de1d9402e7283dd35b8d2aeaca061b6008f2
zdce190776cc81dfb59cc402dcf0515e00564d4ebaca296a903f0628fe74d18bb2e376289ce3746
z37c327b7bf537286e96ebadeacd4469116d024696e5576c032b4b85f06bc577a410a889a0d9273
ze9fa2c8c16cc0574813a2d366b291188c166d3763dcab20ae4b4f93ad16d53ac68244118382c20
z574a26c71d229e9713b4bf44e7276905c7665b22673d970c5abd9bfdd1c7a461fc8cff990c9250
z1371eebc5adcec54042cebe4cdc613114f769c30a2949017c819a4387aaa7b4d730ed4c9b973c1
z047651453de0af6eb8837db83461716d9828ab3f455b19561c0554555da9495e29c0f08c2d9ede
zbb6754c9ee6f88d8c5f24251b321772d52ad53774a17de211147f9b319ce93649e6edb3d3c196e
zf8ae399cc0ac25c4da1e85cbbcfc721c65a82940d820ddef48167dbca54a73712424ac034b27ec
z374d203b719f60421ce5cea90eb9bf32115eb8e3afff7f0190de850aec0e9d5a203581b610991d
zc2521886560e00d72f4c9de0de799c00c33e10a86921c28526061f78013f47bc960bc15005235a
z215c8e7e28e053957842e5714e66ebdc8f35257aeeb615bc5818cccff29084f3fd0b37f6b3189a
zc8ecebc7d84a80f3f8904ee68cb270595af77bb66930a9a101601d70205abd1f8c05cfcb0d6544
z18b7a3dafe85446c1ddaca03458721fd911aa8ae6a8a863a09422075ed6b4cfcddb7c8169398c6
zd73baa79c6e80f6a355ee953587e53c3899e032615518392087ad33c7c65aed3efd4c3821a915f
z231615d6075acddb5dfc457463df2d837e62a5c729b952ffa08037a6ba138f35fa4b4a4377fe7a
z3833feb185f4d7cda6716aa5be86290061b0f71caf4b6024db8025c9479b1372fa76480d3b242c
z370d4f55633d9dcd1ca1d17a6da7715accc0f4eb5d96f0b427ab69106c30803f6ee5d9833acd6c
z3ce4decc4420568cd14bfd1121bad8705806c4d81aff2fec32cc53ab7b054397a0b0c9bbe5bc56
za3699bc7c0e9657a63c84f53d4fdb7dbe32d7d405e7f827f4cdd243185205369082411efe0f760
z05fa21718d0f9cb78348e859723f153d67911ca1ded82fcf076264bcc8dfe51920b56126dcd32c
z1cc8a480cb3ae3f2e19b3b84a64dd84c5207a9a9798fd6511e70e91b640eea4f1a1edbe35876d5
z1ec43ba4fea76f0b64734af3ef331325b69c0bba6861eaf70775b39a8c7f3cf566a908856babec
z2b4fc10fdb856341038a2b6b467b147e42e7a670185f6c1988646716f42e6083c9becef86f9020
z75130e47b295926f06a961027f666cd325d034dbfa4f4fe2c9ee7531f4f830923042972bcc9d10
z24e5446789e69106268aea215ceb5c5e775788acc676448149189dd30ade291ac052ddca2aab2b
z9831dc3997c2354640e8fee1f1819ccbb5b5caec7f2165ec6a3df41dbc2ad9e9bf218b59ff4753
z31562be76439aaf03d7538f6bee84d4540f4ad4481de5df8bd3f517cc6d77a92bfb65f037de1b7
zec54055b3e17092ae734f8977ec1b7a3b2e0505b183faf6aeb41402d39dfc78e13bc18d8a5e4ac
z8b7f5da22eb40c2f9fc2c62cd2e346e5062ce771251a673a301b50f170616755155d0cb6be38f0
z6d2ff4d3aa4af008dd1751406c785728ffc84aa1ddd036a7322d917e2e60e56ee893ba9c5f840b
z73f618f71486327f698b0c052be678fa432b5f25ecf6656f0a513eb3a4acba65995796248b9c53
z77010902e90c37d89c385b3b7fc295346ee47e9b602a6e308ed30d6601a562f9c520b51edafe5d
zccc75fcf0f5b92db2c8e6b933ad8957dfac4cac52ba270e47d47de9982e65645d31320a4dc4e8f
z0ebb239cf27d5fac415d23b83a35bfa5ced26410bc5395db12f7111590e30e9c6ea19ea0443113
zdd83335b60595edeed7c814b5a5a2dde8842de075b417deb4ff22b2ce497480227c4eee7f16340
za0b521037a397b6da6d4314d374fb5915d838d461e25be9436586fd86a176945d8717f3a36d273
z7ded437b5e301d3830132cf142601ff4ff9ba189b8e129981fdff1946b1c760ba152553231d71f
z8b71886382f552d9a6b4e8bdfda73fd64ccff8e5c2fb98626e30122f413fe5dd8154ec4714f1a2
ze9de9f850313bbcee51dffe5b681e9a0e71297c001bf2911d324b21c06413d88acd9c781ad850c
z03b903f7e3c2d23c6464a7381677ddae35f2e5587e9307f107916f00b351ee714466541c858db4
z57fe3e0f0d4fe9597e51ae3c10576605af8eb2eee055fbc08e3c0f675f9b927a06f393642513bc
z6e7d17010cd5b07b4c7a97240a723ac33c73b02946bded1ecedcd9ac2d0b2b1252e83601749730
z994c78a05fbf9d8bd29c2b2fd61cba13772b02ffd8923235f64ba2b9fd73ffbcef0443b7bbee71
z257cf9926044764edc2bd8cda88c3f47221abe8dfc79d454e64bae0a677ac7e74248d71521a3f5
zffd368bc1ed85ab6df2ef5a22a5eb3fb4cab7a49a02eebd98f478d59953108e9a64f962ad319ab
zd72640b57f9ee40954d03af1846fd29e9e6661fedd5e66277e7c9f97df375be0af7f4fd5b74cb4
zc1aadac0a8135a3145b7eb5599928c11b63c21a7445165ab7915268ff7067824aafde3ef8ead91
zc09e0bd8428fd8dd76d06205f8ee68d2e1b7d7a84943d0ef7591921a2da07a42be4ef6793b3cac
zd99e2863bc02fb6a49ff58cc77f8464b0605533d9a6aad716905b5d3e1cd11b504b41ebf93ecc5
z826c9da98dfae55804c200204c448436b9885f5b74ea8f7410fcc0f9b4bfd0e7bc849d6358aac4
z1229c9fcdb4b5e4c9b5205b306ac4c7822e6f4efab58ecb036f4cd8aa6c376ae030569e1b4c107
z6b5ae6140f34793712f803d652ae182f51699995c247137e83b4d4960c088d8e38a4b04b90fcea
zc715cfc91e6f713bee66cd0c3cb5f6e654cc973f0456b15898b42095b3a41224301f562c73d68b
z7587f1b9154867fb855f9adcd01f1ea1da90907da2e4828d255db0e648a709511181fcac93d350
z0f1fc63a155135879979c09dd8d1d8df7a5d18d486ce1d244445a4f85876ba41168b1edc508ff2
z57fad0643d9b5f629b2a957b6be4cbb627bc7c91bc435b7ba3d5c4cc5753a9b898eabddf89007a
zeb014d431e690e37884116868ed69efb3e35d3ad42699cfa6f6c175ff7e3fc3a81564f7e266fbd
z2bb6d3f9d33de51ec18176699f0d32a5886f870fd52c7fb78724d70eca7635bb408782bcf352b4
ze38cc433c4853239f5b137cfe7abf3d9e67639fdd60a8ef335512a8ead148cd42b22a035068ae5
za8650497985cdb5c3f8203bb7f28089a72b8bf40cf9c8836b3a53dd39b98d54a604dac6a7f7bca
zee863dde5175657764b1048e27573b87b0ee1236e545b3b5883e9db80bc470bb36b86a55df0f3b
z1c506de37b7cf65867cc143d3bd7d10321f44181aca097ea56965280eaa33755504b08b94e0ce2
zc400d066b10562074df3d16905820281604ca501468c3ee6b5eb8eccdd2d28c6df2a1a6fe9a8fd
ze9d1b5dcf49927f7e2c1d6c848b368363cb85ca0b0489472ea35a24733dfa854ba252105b71ebe
zacc8f553fd4569548d297da3e66fe4bc95e71d151b6bde368370a6f5be755d19b3e61d04e56c6c
z94302516e923c33249fcb1fa38c10cf20e8a32a9764b15230ec184930b4eb78b90558a74f0fb02
z3af57181da92655964b06a3c7fdfe9bb5d0fb618d91e979e4bd3bb5022dea0ec59b0183dd60a07
z155f66f123ece522e340e67499f79c7cf5219cf9a44067bbe486d16bd751b5263bb8b744d95e0b
z735b89c7cd348e41478e6812bd68a9f3e5918b2346910b28ec053c0fc9131445376bed20516a4f
z3bad1fd3ec5066d34160e511e209abc4deaad5a29848f1ee99bb74400dd67fef729761c14a639e
z5067634bff699edba776a822f3d315694235f158becfbd95d4c4fb1ca3abee19d36ef8b525c9e3
z944d7081fdc352bc0e36b14e4b01b665a7e332590ec9736e480170a23d9c309779cf5d2b8a2911
zfafdfb67e80db25e424687f9d4100c604b7a9ee276acf795249d52d45c75767a9257b011e9c6d3
ze7f888d5f3e920c8aa7d8b37bfaf5979746526dad09b0033f0ffb52e9c171220b94f2b520afbb6
ze41ec20157d912e35aaafff827314f8b89a37f438c3b52c28b56d59f4815287eba206755c7d532
z0b1af34c16272b4e1100a8943b18a82a7d443b79f1ad3f759f9279185da47427a4339da176bceb
z0777e8e8ac3c409c550389df8d4bd7d9a8e68a9f336ff5a32f0dc8941f2be875a925c64c5d86de
z0677f9b65336df63b73de223503c1edafd428da1e2a4d40b9158d3f1e7c4b56f8234d38d0ec034
z0e74b61be0b999f5bbfc0eb924ca39a41ee4ce80184884bd8506e0902e534ae88d72ccc8a07df4
z97966a1d8d1d60e468e097918b41c53727183afe5c0195c54cd70f0aa3681ceb281c063cb173a9
z65e28441ea382d5cff7043fbb5480287ece2f900026cf3e303dd93a9ec03ab417bc928c3f0de80
z6c31567a4c667cc7306b175eef147491f163ca7f4b869f0b4ef79ae5ae419ba76fe3ff63a741e0
za5776b696717823d065e51005f1d8ec51ca623485ef836b2f90fce16a053c0006cb55194de55d6
z471da44e09b419138695e5c4f804816da363e3f2eb2cd2de52feb6515bded02b8e1162e4d89c74
za863a4938e194fc5a968f7a375ed59088477a4d252f5ead4630edb3b1a280093591cf1a0d3391e
za7fdb4fdb6e3498a79b1d006ed805f5dfbdb2fa3e35632aa02df0cd082f020f4747387f0498ec3
zccb2e3bb46f34da7b49242a055a8340cc7cadde888acd31de59ccd74f23014f5edc2506b71064d
z8243499386e81b6218462b41985482f52c11a9f3aa49a4e1d4557b5209355e6b8eeac89e271df4
z61c37b8cf5dbc03dfd9eb5fd1b9a4cfe58411ce2567b4681ca7e37fdc2c1931fd7fe99169273a8
zd8232d96b7e32fb3a40693774516896709757d4228d9ab93e46431f5c3e57f409480ac5e048c83
z5dd2f42380de988585f8250695a7f40fbdb5b30d1e6f3616ead541f67de19d22c75edd911af61d
zb5b8006d09568af3a3662df7dd87109ca9c2de26b7fb048dc00ebba7b695991ca47a8ede41112f
z34316c69b9ba02d190534cd5b0198b6ae78f7c6a860c8711ff875f12a189bd6c30638c11e53f8c
z66ecca77bec546a761f593b4fc0271d6baae9b8815da49f062e78a4041c92dd616e1dbf819351f
ze9c47194df2c0f929e66cb13a7b1aed79ef6c0eaa89c72558ed3b77ee930282ada273100db9ae5
z82160a02bb691f227ecb8138c78ac87903596b616feac35153d307a91d7479e0f7b58109f506ba
zde30a462bb37f7bbd266670b022a3d58148804f1581b549757a8ed8062b937e2ea410a9c4acfe6
zc7dbf76045c4749c28954290a7bcfc02d238a7b0f052802840f5e3647fc89f8cac454a5432e56e
za60ab3dd157c92a4b334fd5adf5675f850da89e4ba740ea403f370de4efb60f8d0d74b5d844048
z9fede2c6e2c1022f7212af9afa7689bce970463e642cc3c0ae77a6bc65a3e4ae11e1156c30d71c
z88e4a3b03a131a0e069d428da77cbf9a7dfab59ba1ebfbe5c5be2115710fa4425e751d916aa06b
z24c5d98bd2b9a4519595ecbaa3594121edff96ce519dfd7249931cb31a487d909394783185859b
z2f48cbd9ac0cc60e23e4d045a14deaf587a762ef89494196aa9686e75a954f089a4ce39ae1509d
z8e27b7fd3179077c4944953e073476054881e99db527f64da67f4637534e16184f94056bd56942
z3b66e95c546a3e7abc800f7eeddc8e049a09bd66524675be6644e304cadf0c04983bcbeb35a2b1
zf2b03ab29e6ed74b4aa8f38647a8e4b3d9a23c776d5d0f857ab097490be312c4ca18a59db6ebc3
z81abb2c75b61b04108f8867cebcaecab1d0379263cc51c4ac4e2a8df8687c88221063894a659b6
zb77d50fbe841bea3165535d0e12c131b6a01f1a59c446af675ba1c903471a413eeed241d76616a
zb64f13740ffdf33ba15287bb42db2ba23d36eb9e3d4a6af196c4334a6f3e9e7d92957b68851cfc
zf6fdac075f64f0169aeeba07ba4b6288e7c3a1a1ee132bbe00c185452d7588178ea36b1ff79ffd
z748d29ff060a06647d4faa9423859b95744d6df49e0b7aef42003c4491a291a4c05da3e821720e
z90e090610ade733c5e064a55b936b65eac7deb3dfd7d533f508b3e64b5f20e48f3e7b06f9d60cb
z9be81657792bb4cafc968df0e05b3cec4f17ed287b9b2711621b666dbab1e9ef566b1d8385f87d
zeceeb7e5b159d5be285fd600a57727ce523dcbe3eba85bbc735ac11d54921cfd31f7050d0199f9
zb06fdad3fa17f822d1959e8f7767a8ec5042f4a729942058d8c41d7789f95d393d07cb571fb1ce
z04051fcae35e38b5b993bc6d64be1a42b03532ae72813e218b2f8cb7c0380666c75c5c4c1f4553
zb3da7a5c4d40ab413ddd275ac3f5cc7e4014471f4ba91f04e4edf06ddcd1bf78f9ca5646b43709
zfa109887f23e1bf69121e79848561a653664678a28bc6e72ea679d68943ed71658f614b9aefe71
z095c246879c1398a45b46b0cfc3790c5b03e122e60c5a73d6ecec361d002c43ca3bfb9d1e984b2
zb0482f2c02331c8bd4869638e23463412ae186563b13f60036898c7d9eed82325fb5049490bab0
z75f195eb241c9ff0065fe0285de4a4b5e43039b3c65eca157c4baf1c4d7525f8ef36ed23b1415a
z29793badcc5736baa1046b784367956d78abb6ce15a1ad18258cef7371a4e2ed6bb7d226b30101
z8e33213441683dae35633c13b34bfad321df580709b0fbecebdf76311012ffe56ced90fb4efaeb
z15ac4a2d407d2b6a58fb0bf08fec0858c24ebd36586189a25b2b1904718334d4454dd9f3e497e2
z9687e62455a23491a8122f25971c9b24ec6de131d6bfd0b5c213372afaf6663e94e2fcdc8a5d1f
z45f1dd9efbb8350958ce5e57d384af162870b89e67555b1930692284290129948d0469ea138858
z8ba8b963397187b477c7a4f5186744b8079662a4399567d5d6bcd8755d85e8bedca4414d15f6ed
zac59a9977727986ca6f35d3d8861af1a518869703c1253279a07cf288bc41653e26f525779cb99
z6498b67bd109049300d3d7877679f97205e476b8e79a34b928266ef49a37bc8651f9fe8de57cb1
z0535cac066b7423e89d39f7e9d47eb4cbf3685ea2bf5f7caf11fd83018a44859eed4a77e3dcd22
zbb241d95b9d1549001e7d0ff6c2130de61d4a885f8152554f53cadeef05b6cf7aad74e9b084b31
zbbff73db35e9019781764d851c1e7954fcdc89b8e28d327a61a125be06757c0d646c67c558ce64
zd7b3c03495fd19397e3eb8eed87419563b3c63dc1be5131f5d8f67b20486a1bd1854e5af191271
ze302f48cb4e8dbc16110dfd6c85510cb387383589d8ce757a73586009509f2f0cd8b5afce51cfd
z0d3c0b8ccc1477234ec120bdcd77a6c66e4c2288db551c48211b2c2b0703e2315ab32e09b9342f
z75925de7455a6a4c806dea080ad6c61b4396f50c125ad3069de83a6c4e546db970a7bf2a3348a8
zfd67fdee5393cea1434f34791a7c08105a209eeb2ce0eb21dc8305dcf3f2cd40e60b290291390d
z49869eb089feba7099ba9d100b6dbb25d7d49815de64cfaa6fdcd8275d0885a7a6a46ee263252e
za873589b580584a2d64fd000ac2ce806d03917c62ca4905f7a43422640bdc15189a022f596a558
z6b38b040d325640927d2b45626a6c3ccfb109c2fcb20fb9546cee0c649bc802aebf9bc88e12c12
z936d16aef3cb8f726ed1cc5c3f4f95bd8d58f30425bb950665cdc59aae7190d86e48a9e7f64904
zf9db3a59347530746fb2de00b7d85fe53ca1fe3c8c85c7c4b02817df2e0fcbccda6b8c356c7839
z877291ecbecac69bf931a5c00880db4c7d666b25690ab102b0bb15bc685f04172c405b87dfc6b9
z330db77ab092a5bb9a18e95b3a0d5cec8fe9c0d144e0b9a680f4efc6cf385bd18b13ccb9b2bb7d
z57abcf55b19dd18b94819e4e94f6fd70ec1563879bf4f626eb655f2061be0b4dad7acffdf958a1
z793eefc4a0944ccef64c82576af1a801b4a018cbe918f6e3acc4a295af8d02ac3244776a0cb939
z1ad2b9748611056b6022ff58c8a3c842bd6c47d7dc4f1615b87e07c0b63eeaecb7fa916e229c96
z656adf6635f053e4b16023a0c0581f2b4f796620357b6870162d7173cb6d13858e1957116c9852
za09a08a26aa2a649c44393749a453d414f3c2926868fba38aec8d62b86a8485931bc4bef32749a
z529833ab3caacfa720e30eeadb617f410f5a6db42bcd62e00f531070c9413fd51436bdc5869b09
z6241e7abf1148c620da6351fb562d00e878e98349e140130150f80e0e8a48fa2fbd9f21be5759d
z40bf74bd89438d134fd3669529cb73480f3e2983a7b0042733272d7b73453a7d25fb2c498f5218
z3385a7690064b5eeeba5157f19dc23f2e2bbbe0701c84d3f68ac35cb66608d69c766327274a125
z7696304493f2b34d9e1a4fef3b6497305d941ca6ad25581b01b7833b26916ed315952c68f745e7
z82a2f5bd3523793a364e2432c48394846f83c764fd727e6035929fa7d41a2b921f7a9a79450ed2
z055c3c1cbdc76c091f976a81b1b28e2a964458b414e02e960baeda4509bcfd9db1d9eba478b7a7
zdaef90f2cee7110a821c01511793610e3631b597f4a6d9491c41079475c24672ee277762111110
z7ace21a97cbba18c16197b5476fc1fbbe36da37c53e3de7f4fdf7aa34247cff1a5809591c8bc47
zcd6295ddf35874d048dd6b0539895b3ffc19fbfc5963af5809513509ac4587112cdcc07866e5eb
z17551171fa5f6694e990f090aaf124be4f3cb13070a07f89b54509f1d8e8be1e6c1090bcc9f511
zc11f02380e7aee882abb59b7ec0f447d94bb00ffda3eafdf1c69bf68760d7e95d0b118ffc1f083
zfd4f6dd3f2f250b75543e572b0c41eda33a177723b5de9814247886a016a402ffa8c7723aeac60
z666bd2899950522591ec0ccbcb772f5dbc34fcbfca322424a8f327f250e9fe688a3f6d5d9f8b28
zb07b464406f15ee894dc98b064f801ab3901d3875c432ac118a25c27335aba533a3d489af393af
z11b9b2e60ad40e2ff08ee3561540d195d311b1591a873bb79b130ea92987e909f43cf02628dfae
z35c8b9a6b7af731910ed529ab9d9ab7fc2283ac7a12cd13d12ca3ed0d6a367cc2afd2703f9666b
z11c3d12ef190bacc5b155b33bdc0056173cd973de04d9c0997b406d3f3e9074c3e021fd6af7721
za4236f7c1954be62fcfe4f8dda8228c718564fb780e48fdfcd34118083befadf1d5ecdb884e8f5
z81185a6568ae0be3f655a18275a91fd383002e99af3d42421c409f7eb117cff5f87a030761ea27
z27995cb6196148ee02d7ed1bed3b3f5d60c6d144fea1b606a8a27410524fc3511f846cb818712f
z9f9f8122dae6bbd94355a0302ad6e74fa5301afbf9c06bcc77e8c00c973255629a040253d710a4
zc29f7b2057968109b7cf689d65559d941bcadf6528ef7a24857cf306f52a0f30ac5b13eea01ef9
z08b19ba791c0699383126e457223edc42287a78725047986e3be2636f07f42d1095db0e0cd0c2a
ze1644ccebb3447f2e0e6da42433d08aa71641d773f70f34e46e5bd4e7152d90ef51ba17ce265d2
z8f5e95e31cabaa72143341cf79416919097780a29924b1e188c052b941954fea1d222f1e077082
z028b78fbc39d12eeb484156830de0b38a3c41601a575b457dbd28762b80b4aced5552164b44be2
zd7ffe562373a57495518a0cdc58bf5a869fa8406cd85b4eef3bbcd8322f7b339d8146ed7a96d3d
zf8bfb5dc05e1d154797a1d00eabf111c468ce66f0b4097ae333cbf69e21348988d64b993d39229
z79b6a5c1d1f2a4adff51b3f3f1a60c905e606bf44e15465dd85fda9a25aba1cd944f90c87a614c
zbd417de6a2a953884765669d81a8153187b95bec8f0d0ba4101216f2eb9b6c037e7c9f49521f2f
zf234319273726ac67caff090a8feff006d64df70fb7b5b88cebba8d75d62b636413b75267e093b
zc3003de0bde3be7f14e80bbfee9b1caa4e4712e2472556e30b0c50f38f3589d390cce7f44f92b0
ze01703f0b5faf3398b3e41f0b4ede479daa75e5cef62298d6d27dbe0f9c6a336dcdc24e4034681
zb601ffd9660b0a6abbe1c7bbb9a9477b400c8f4732f0d440a1d043b14ebcc5a4902742178f6f42
zf6f4940ee1e8981a6d236556f1d6efdb2d59f5d1c9486cc91182ecb6388d89a2a05d41d1be2bea
zba0346b3dc63d5781df77828516fb6256168745f25da0b74f5b1f6561035ebdeb31aec5df61b6c
z61004d4b3a2e17d877b70fb1a6e02009e3c5916ce0d7f8a0aee7b678ce949991a55f3ce69797ff
z0b813efac20aaa4006bbd59fac6ea114ab6d29822b0b65a45977807d31f85bd6baed62cb7356df
zad450aee3b20f92d786866773a034247bc9b40b6ec9b89aeaa006db541d35e3bf0b381d7e4e192
zc378e6bcf232716fad8f3a87521d6a05dc4e2e1471de6cf6bd973f459155068ce1a7ca44f5ab87
zea291e7368081262445f227bb788c349f74090b0970d829845587cc918cdaef7dfa98990127398
z7bd631e21027f3cafeff027e6af90be90da49ca3b6f83e39b2ce932a5dc033243aa25416658dfd
z7f554717e17ec667330fd720bd5b47c640f13e1cdfe9ea74a9a583524af0aac666f6148c0f2fbc
zb4ea6976567a6904c01ed2cd2acc3b1f0e0adf7aa3824f82f0767f248e9d465011adff2ab4e12d
z573f21bdfa69a74037a3918f299a07aaed7d59469bff62f3acd0784e3bee6b08fc4d96e3720b23
zc22122782bc0895acfd2cf0309a7ac9cd580f34c794b2dffcf216324f86aafff4cbb606b51dea2
zbdd1d46d18aeb69d0bd1dde68fe0b084321e1f01c5aa40e274b8225db24c081eef9cf0e4291c38
z943de97946f6e0bdc5f252fed6488c133a42b06031463050cd197e8749ba4edc25fc70932181cc
z4dd72e1149dff617d651a167b2fd50fa1d3e8b0f47ab52b98d4cc55747a71c17a3bd09df43a344
z274048c6a303d15eb15b25ea552f1ed57b3daa41953f38655671e117768b2e701d96b4b63a8e35
z750fa40c21d02bc3d99ced1c8fbca65cd37e6e623b57954329c6d306e22b444b44fdf0072b4372
zc286e083d1d1eb35507c3b52b4300317ea6770a38736a8306258c126404d86c0f3814f94e4d02f
zb1874f4426c29de770f9eeac0af71f614c8108b15609a1f1f0d598499c3cded66aab12c14f2529
zd68f94c3cdb218620dd86e077d9465836e72f805d9ae319c3a81d60e4563e9265396121d96d551
z96f036f9a662f15a82bee6a1d9f8c1e0ca1d6fdfa05ac085c83292a61dcaceb9de6bd3ab90a46d
zfacfd9771b58a9fdd5615c00b9b5380b2489c22d1fad930d61c2bf85874694d086683be27c4341
z30df4d6b71cb77d6f9a8f7b5d27558de99ece6c103e57a878c86c972de1ec2e538081a37a3855c
z0f07d27ceb5e830fba973926fa61d45552cb3cedb195c2a70fa6dd1133e457a415abb7c87bfdd2
z7ecc1210617ae7e6ab49ff6bf39bf8deb183cb5100badaa54cab1e46af0802afecc5dc1a636ec9
zcef7cda38e27c6167ebda7e672d5676d5e354a717a656e43c24ad6181be6ae1eaa531fb91ef53c
z70074a4485d0a0c9b17e76614f5ef200d0e9aed510a9275857840c2211a98d9f50f77a6521c3ee
zb39535513204d295405380a26a0e5d25f42c4711119ef1c0e1ebddfb8cd53546340fffcec0b186
zb35eba3cfd8012cd816439d017e67f238eabb817a654ad05752e9cf586f3f2a86e8d35a0ff6364
z7e7db94c8dba5438316e07c503d84f377b8f742633316bb0eaf839bedc49650cb259def2cec356
ze73b2b1fa4bbd01bcda91884a9b90a2e199b264f35663ace454da455354d757c0cac297988ee39
z3812fbd0658b24163ced82bf9155b40a33ca76fc8a3fedea3e6ff699fafbd7d7a396294f48f038
z9f0ef1f1706f145d17d2bd5fcc36c82bdb2f41db124f52e07506f0dee3858b9454158f8cf5a199
zf63d6ab5cf43116bcdad0465776ee5a2ec3a18269f73ce23ccb916116f5368aa229ab18f3a98ae
ze8583cc9109a3490072b18df2d209b4bd7b4e66f331060aac6232d97086882e377d68e2593b538
zf85648e00f3a7965a40d6e189f5124887c95d73997c6dd8215503e8da37a7dca7ae53b7617d1ea
z54927399cef93aa2d5ca65eae2ffc30062ed41703660dd45acab866e6844c8badef21d8372c879
z7625565c9d7119b3007474554825c48d22ae272b5572fea5da908556ff1ba04a38d32c091b1567
zc44dbf9d88b154091ab8ce5c554033e192f985290d6c5cc994a01f9beaf916fc012e8dbd4b5a83
z7eac2a6cf82fafa0ea5867718c278e0cdd2855c47894b456acdcfbb203256952d1f616bf96a11a
z0ef0d69cfc187c6b81120d1d8d9a57af245331675c7a804274853d4a97ec638b389af7a153aba9
zae1358576ff8afc0e68b28cc0f0f01914faf5ba619e73e493c676f9c53240e2c0636f3cfdec5e3
z5b47c85bda82c39e7ad18da8c42d0c9c936cef9a9e8b2e0eeac9c8030b9e5490e101a315f080a1
zfb576d980a8163bc04a2d0b7d589abe48704ceaabad49fa197ddfc1b3b568bc1b98a65e7fbd796
z6f4dacfabb20af330d16efbbf084f9b2cda2b69974c241b0ab669fa37f19235217a4d1571fb2c0
zacb2f31295c555956092e08f5cb50af051ec495302dd05ead65ba9d391406e6634bc9ac425c598
z1223074390fbb318bd4a6fdd577ce42c8583190351a5e67b075c8e38b382dc95d2098f336a08cc
z470114c8795001835ba29c610ed198b239d6cd282c3f4a3811452081a7725db30c44c732b50001
z51c426516c4e3d5bdb21165cf0bd7b50fa3462ef67d0b7075cfc9e917c1655d9c06f20e68147fd
z41f76bad0eb903311b7217824caed72341bb985c17f1e56be126445f025333ab143743ca494e12
zb34737362852470b8abf4c4d3b7e747df61672ca00faedc971b7f78228bf2fa25187007b4e06be
zefbd3725135de89c26f4d9dd0fd3c9b59d9b6bacd2812629906c005f6a7e9258ed2fe9dc38b065
z6f5a4aab93adba336402e1ce17ed72de6b04334c0578fbfe0a56d81ff4491373b902aaab08a62f
z75c11d742760fda5cb3e4d4e454d3d74aec4523cf8858bba296d4a1550be210407bb90bc19a861
zb57883e2e553f73b05d26a819ffe77921e977c4dd3cfa04e50965b5ddf6b5e54a184fc56798427
z33c3fb646bbc2b07802a2013928850dc55e403b9b758e19fa25ec4c20840f29ed3633a246ee221
z1b27d74b50865060041ae2264540f8eae284e2cfb2ce3623b70f0f56412632638ecfb5ae8edb85
z269fdd44d54c7c64f28a9b13e58522da579811400604116b9aa6883eaa2c3ba1fbd0b90641251e
zdc3e867f599f3de41c60ca5a83075cc1a9f207f85eb0da9f60dc947f74adc41033b71531be8647
z7987048e8ee7de5c106f1c8e937195a36453e268cd04cc59a48bc536339e287c0e7320020aa9d0
z470d57559ca52713892a32e63a40b8116f2e34db37887124464a1fd74556c9ea0e25c4f6102987
zeb9134733681ebc1092620bedf3cbaba8b71de95c44602151f763176d0b3cda7631c8d0e555c01
zd70d9b7cdd7371463464b765c872df1d402999227c5bb11ecaa65547d882d91af41afcfc06d768
ze68af1b6cc1bb68aa68eee5c27b7c593e45e2c71dfb7d176663d57d0fa9c41e77cb703167359d7
z987b4c66ace3065c182d4ec6b1dea0a9c4d193f90b703e4a811a3802a57c0c06474ffb741ec284
z951b39a3cdeef62f41ad7686cf823460890759e668f4bc6e6b58961feb49378bd10a20f6ebffd6
zd324944c737f64f98a5936038d538f0295065c8da239745152e3a245e6886ff97eb17696c84425
z2d308e96a0292e341d3dddabb0ae807cb294743ae1c6afa044ed1e5ebe1f3a622b8bca0a61ce3d
z1bdafa30605b92088d21a3c2c0ef83b8836797ec85054042f34284559c280c7fa726fcfee54d43
zb9f19992228091899ed118ac34d25295c9dca46089848d8331e947027fc0b2d6ab10ea4e8fa5ff
ze0cb7029d86d49e4c20cffd4dc50f57c1fe3db3788a7ff70f4a18c9e86629efc45dee6535ac1af
z310682d6fe04aeb610a8fdfd4eea154d5e1808e3142a90164b5a5a176df6aaf77e6a706da68de4
z058e2625c9e8fe8bc38e08ab4f5d57d0118fd6c8d3b3589b76b3a649587d6929876419a12c2cc5
z9efe3791a91a7cb4d81803d231de12b53957c1d7a0b4c9a5caf8d2fd67f9a773b610965b044aec
z5ec47b28768c67d061f1a39c72493d2fdc9f977596bda61598991ddce274aa3ad84a6fc718dbd8
z1bce96b2df9667ab883852eb1199d1d8205403e336792b8b08c910da0dad6d73e4c61487656959
z3700d675c7eb5aa29271ff4bcbd98fdc4f042b8aa6be6988ee4223ab0f25c98052e4a4aca1a028
zb87d5397dcfa54e8d093d04547f92e814830637449e032715b52c3ed216c64291baf046a16191e
z27945cf7bfd17d04c7115b4571700a13b5ed2a0e370d1edcc3fac2a30080750a1dfb5cf01fd1f2
zf309468b69eeec6ba44d5df837eb21a2a2590b58bb5a7a735051097ab57d3c8badc2bda0154bd1
z2e3effbe0a413e78d0d9aae6083b1a4cc6d0822b9e58266fcd172d520d782f31ec4a4e4d37eaaf
z786148f0d1e11796c957061314ed5a7545105d1fe836a7b71cad6163553026dd093753e4089e76
zf5bd1ab8ff9ca4e17e0153cb537666c7f46b4bce90dff91b0585887510a90e461374597bf6b203
zedba38aff9e0bee2006872455c318b22a8a5fe172cd6146c2e91f00ab4e610d69c30c89f2015c2
z9728fd1c300d8a7495a9ebbd3fa1cf9730ba1c45b236c6aa641d2f13c2c2d582bd79040042074e
z59989b65e2ff9f2494c24316d8e5aa1b087af9f7066e34186ad6d3850a31703aeb0a689b0240af
zd0176f9bf896a13c1434ba309b75f9ca847ed6599ce879f68cf97cc829c57c222fbd0c8d45147e
zaedada5bc4b791ad3f34692fd6f63ed110aebe3a523d97d5c35731ec1e1da85121d1b4dde9cfb5
z6056f3914c86f1f4f77307628bfacde9f78857471d13a4ad73409c1918014785c34b40f47959e6
ze7c6dd29af146958cb60efd62aedb86ff29bfdbd73b93f604b8d120ee48549e88196872c908fe7
z3e7e6f536ea422cf3c597602770545262c74e02c131839cbccf3ad4a0467850a8f99e50f594cd8
z3e77b85cd6e878735ee5658b9baf69699ba62c7a91fd36640da9d219aee2f2e5103dc657ffb7b3
zb1e138110af36be3544c814e8d98f84f201b6aea7729d31050721dab2550a540663ad1e7ebb34d
zc581979b0edff651a9c20d906fa4a10f01fa6d95dc78a7b4d1c395a103a3bf9ffffff31f94991b
z559427ba733b7b74d314d2f68bd5dbd94ec352f8b096e205055cff500a11bc64f9346cc0e5baf3
zb22cfaeaa92195ca334d52d0b36ee13f609a4d591f3db3e3077fe2e763e67d72e9f973cf69fe95
z0ab07c44f3435814c3d35515c073b42cc96746c9fe6636d3ba1194bb8204810ea3bd6176decd8d
zb6ca48ce4edef7ed5d2f4977840abe6120945f2a2ea49e05e54d8d8e265f1c2f415239846bb99a
z709fbaf0c06c4c2b644e432066eaa81d16f9e8a6bca4657dcc0d70ad8e4e728a83e765b549d8f1
z58764df078bd35f6a97b44f423f895cbe2a117feadad60466745d98adabd856ff389925276eaba
zf5c4d36850cbddef1f3014882d2963d898af2473d5eedcbf7b29aa71efebadbc761a285f8e9e98
zca07354ff43950771080e8f65c6971920a3a36d04f71c20b593109a846b36f02db4e6890e31b5d
zd46dc2e5f2ffe915fbca130fea238054cd9771a2f3b86906f4325112078c05e092998a2f3f60b9
zef594ae90e221b4def0c880a201c357c79db371d33e31e9efcaa461f7994e681a540f11e13e3c3
zf7a49518f69e7750a543342e2ff2115873d2b8f1395a894ece796e738c81b658a7329554d28aeb
zad58550b22c460441b71288af220f502e46bcc512bd9054ced2438a9b6d7d2669e22b78ebda6be
z874c2cb5eebc5882bd14eb3cc3b7f2c966a6c38629b875958b09d2ebc5dc3e601b19c74cadd6ad
zc489004eb11583d4f871c7a7cf6dae400975c1fdabdc3a6d0b79f20f7a87b37936d2e20bd0ecdb
ze7d8b91dcb3c011c85d8017335ae5694aebb727798b5afbdad3a4939e8b2f823a685eeb7c7abc8
za38a68fa3c07986286db3ddedb4608d3dda2b2c09b0601ebc171c2a4e8a867008eaea85d96222a
z4b248e602ae4e20a143877c0ad1c37847b43d182ee3ad5854a28592d2842d898c479f89e93dc45
zc717aff09d1013ee51c3f7a1a4baad46bf224a9fdc1db97d1105ced61efc72f91b9171d2d5469c
z57a2134e8672413ac0c9a784bc483231f37a122d1c64c475d43c016898586d671790b18097f368
z615e05c3021b1ca957d797cdc1b131aa63c096fbea1be30ce66503deb5f54dba67251ab2570178
zb0a1650b706ff2d5c679823d322a38d32201dbaef33ea247ceada7e2528f5416e6d6785cc9e96e
zb9e222862d9118af2e286c2b6c2649b2189a55b0ffa7f0495c47e56f4e04673e8047dd55de4b07
z482ee201bfe2f19a91e46b140b3bb19441efcaf1cdc235edb33f098d96544a8074074bf94c4bfe
z7b8a289768b50158a26efefbb4e8886b076b2ea5b0724c492e506e479fc2f4aff9619a2c833ac9
z6614706dd8159c26f43b48e503f1a416bdc2c86d10697a3135cb6f32dd79bec3023273a477dfdb
z3a3c427fd2f25d80259fea80dd1942d666a00ea9311fdd93679cb4d5497d24f43d5896760ed02c
z90e1b5cb4cbeaf93e113368ff2ddac0da07448e9797ac830f6adb22a7eed025acbf4628594202e
z080fcf23991676553a2d0fca599f04945d25223ada03e7339003d79f99566476cd51686271f7bf
ze0fb81434b700a570b51fc49983a165eaacaea13210fd3277f5af5b7c8c3bf8d175693ecffcb2a
za5fc132ac9246f14c29e3626ed48b8eeb230bdd30d5cab210b34b5d64c97897569c761ab314831
z588090e02cabaecfed098fc7fe2e79dd6d5c1774bbae6140931e5d40ebb03e7d25957fb53fc530
z4c82533f040d161c830f2061f03f614efda8e7d2c5137ff78dce6d687b2b0f0ab054963a84adc6
ze219021a8aa21244c93a4833de55db9d94983b3f6433c3b04831bc31c550474f9e25d326649389
zed194ff52a6a636c33c7ac4b8c8a7a468763336baa78c8770f6e33a73daf7c95e672673d58a38d
zea3cb42d3232830ced8fb64284d6f6b59aa546c675536d183e018eb1c60d2c850b67c7beb45e94
z6a8033e641ea1dea89443b8afff3d1103158e7f2b52305050a9fdb8b4f58425312c4f1b42ae45c
zf8540677dfa6e26f2a8ae2e2e23a915177465a320c1b11ef876abb6945ff5c4850af0c856c5a15
z900826ad6d6635b016624517ad7bbad33e608399d8a07b629601738bb058ad53b3c150dd7bdb60
z43c7bed2628039d02f6a55b9906cfe4e13e4122b204674290e059a30c4a133f4d6cd72cc364caf
zb3412861989df9aaebf0a91bdec422eec27f43fa3172ec9c469a48cc85d734d695206c8b8f5e68
ze5c2bca5501b37645aec964435eecee2b2c49c1482c85c4079da88c88ad6b8d4d779321a58997b
ze1aa7325bdc17cd70f99f20bcd99ae219c55c24954610b831cdd8ac144d288d0cfc5a283d1ed03
zae23ddc4bf27ddbdc450e364c279ad8cc91d1c264003709dc9fc3191e0fec98012d232ab355efc
zade50b7dbeb80b008a1e20f374cdbce0cdbd89fbe312505e8693add8cddab4eb357f2a69d1b259
z2e3d41238fc403932ede01cd969345ae8626d83aa88e8695238e86a0e9b2bc0a281d1b3ddf5d54
zf0313e37cf560e0cf5e6f8c200e7a605c53243d2502a124e9ac53e5a2c7d217157f7ad33457a9c
zd4e9492f8d0c9a2701b2596d6e03f1ec87f3f8d3ceb895df657a79ba02d97b14f417595e52ca2d
z7c2ba989df7d1fe6e58f35c18a99bf6a4745cb438316d4ceec834962077badc1d2dd6e4bbdb44f
zbde1f6d413cd11fbfc197fa829d9f09a587caaddd3289dac1520c364ac74884ab28cfc1921c82c
z1b9f05a0fe90ff9fa63d2c95a11e3a1b1c59f811d099a731dd07c0afd501d32b2323dec323f05f
z6ab04d8e86d1c4e5a1dff6589cfa03e58fac48d5468511a010c18f5b2287d4843e2badd38a16ae
zd96e21bf5ee503f6db88f942fb5afdcca8042c91078abbdf353b4759a57ee9a3fec875bfc9c416
z6109ee2dc2dfcf012e5f005d4819022899a955dbd2657691257bf51e7d15031c08758bf5084355
ze0050fa6930f224c3793632ae9fdbeb3d99f398cb19f948cdf62a963d5ede78d465d81ebb9b3d4
zabb21976fe819d021f56477219fa42b7d4639657d0717f590a49c741f12f3a5b6a5b6b415167dd
z4afd2573cf2b1e762c2342c87f1ddeb1e88ef3d3524b5a1a63fa6bb8089127f79d1a9a97c54940
z6da5d7fd964c9dc451ba536207bd512b0b80f11cb57e03a6fd1e5d4b9345091444644534f350bb
z79ec21c4f8b78e18ef9a65774267df042982ef2a87bd1affad8580f3524996c292be2fcc172c01
z4e737c755b623872114867574893314ca8bec84b1e8576d4e7af30254597ed5ab1b710ab06494a
zfe9479bd2385c2b9238887bd4c5d3a4158df7a08a146c0ebf3e6cc104749aec8b66bdd67da6050
zc23ecb3d17a2c50a4e47614b9b8a433638a3c46bda8c03d24071c3cedc996d0dd07d577cc9b9f9
zc70997d309f9c247c1da94bf9e932835bec341ce64e5cb7deb3db11cde02145de1b38b51a82b82
zcc1d35a2eec93b6cab1cc16bfa62b3255ae46a6d6d31672872a827cc2ff83b09894ad1973d20f0
ze60dfad94a03a37721dba035d131e09ce72d2af398570a2f8d2dc2ee85a7ad7a501cedf4cd7f0c
z91288628aded5705cf55b1c85af4c07190b2b235d3dfd16db461895dd8385046ad3a71d17ce971
zf0a2d3ff3f1b2b8823ff4aa8e7ab4de5a1ec2c3d92d2ed2fbdda944fa54dcc0f4150e4dd255162
z6fcfbfe6c3176f72d16779b09ba2c9f84a24838bc85c106fc78f66055a9877f16b33cdb3166095
z7604b19da82e74465a45fefadc691c078ac75cb6cca03d71bf7df7f26fb4f2f02d26fcd6c270a7
zdcbd093bc9db26ddd87ea2b3224913c2781b29f5459885a136773ecfa3a8eeab3bad383fab1736
ze5b257d45c04dca04dfdd66ce16d8bb8fcbd56916c4e1fa28f43a21e297bfce661f0f71d947fd6
z49615568f250a372982d944b6a9e6ae9f2ae18ab595917fd93e082b2ea20c3a53f757aad806cce
z310966a0efe7a4ea2e45432167148e92ac8bb36798e81524d74757d492f54a88f481eb562a8eb3
zdd90fda50b0774fd34adc924eb693628df519f6de2402000a0fa4ce3aa551ffedcebcd368ec157
zff58a370bd7e3bba250779d0d05886236b84dae307ec675bc0f4439721606bac3552fab44c4981
z7842ec4364748f85cb68bf7108ac05e8128e215e0469d33fec70c54d940c48101e20e809dbfdd4
z015afe18f61ffe49e309ed954d119b1e5fa94216e5311dde8c160827865b7f5545b0abf851b562
z51340668995e8fec15aa27db6d146572be4ca6272368f20d46f7bcd105fe94f2c184ce73dab05c
z3c73b73947adf92ecbe12fdd54b65bc0f6bf30c9daa29e4b0cc20c807d732fc5cc7ca0bb3f8ed4
z92b9e8e54b21c606c04f73e10ac409ed5f641fdc3306352b3000b0895c234b49f3fa0632e7e059
z1fcdfa6d9622bebd4d9038eb3710f14a48bdfac5b5eb3aee4e986d6816f87db3bce4046a80b494
z659042caf70197ee4813a80add41b0449d89c7961f365303123b803a0a76df255e57b1196c35d3
zc46d1e02ad3ccbd058d18e0291de5fec2195e6420b1043d5e1c3805ecbd6e1684b6975d1c08b14
z34cd87979433c95f1c2984371f23837bd24d162c06eb8af46fa76116e6603eadb164594d562bee
z40e9210e94d33c07070b6f4b6277a3dbf9b46f5fa688e73eddee59e4ab71c9b7f1db85450604aa
z58bf793d0bb5bcce5d2b98b0333fd44b877649113655b2f996e516d94725b9bba5097b32b6975c
zd9b935a04b3104687985d98b4824ab56673966a2bc16a56edabdbea4a1013a00f443a15c767eab
z65718a05e5575ceed3b37ad5bded25e1287711a79de6a71afdb2f437e8d023617b3586a47b311d
zef9e5861db10076fed3ebde6c0f0786bb288d0c277dabcfb9829b20520b29dfd688c1378037740
z31d14e3d2c0f1d47f78935cb15cf72967dde6833208a1d89c2d7a1ae1181fca54762fae339744e
z0ea2cc4b01de9c4a000e0e90051b37c7f8004fec1cbabb946f483a18d1a142de1bb02b2af18224
z992aef7c120662bc537fba527870089c81249a4142851dcaa4553a1c9e706519252355fb90d2fd
z1f4761856fa561ffa396d29f84eff87e0c4d29849a55175cac2ffb074ffb601c9fd2fc42136bfc
ze3ea632f23949667728a8d57d9028448be6656ec33a919eb631dd84a1cf9a9100a782b53421311
za577a65c84f51425311ece49bae83dfaff75a48c54d982e711f26ab9f0848215fed0c4ba563af2
z85591b7260c77992b37aa59c2373a503c5d2216b1af96fe2fc17734aed600e9c4ff823a73276a3
z8019aa02ef68c4ae42086d254cf8fd14da5b70b986a9b465c5aaf69aaca3b2fe20818b1a7a84af
z799a73bfaef51a724aedeef6cb33ce6b608ab2df4f9dd4a16d4bf8d75d438a30100dbf7462122b
zeac4c58ad4e04d5711e6d1f65eeac5b66ef106ba0be8451604a4059ccd704de9f4572ff12c2a2e
z455a3646803f463267fd5cde9672b1a080ffd2e00d048784496749722aa80bcc11b92819cffee9
z02dc2e7fe6745258c2a35a2c4976aa1977f46a20afe320ff6d5c63bf66861c965a358fa6931a99
z6e80ea9d734e4edeb76cc76b8becec5c2dd6a605cadef7947063770bc89410a089da7c20298f72
z97ebcf8c9cc000f818e70054b06f7d9c43d5266d880fe16c94c6f1d8a8d1cc365ee5e24660a78b
zef58758515c24281a872e527b44a3989af92f62b1d38ec56ecf50eec1b8fb72bc57a1207ee0b76
zb7898b5dcb5ba0050dcdd0671fb2c8a9691d04a2577401b9cf7bff40afce04975ee90928718ebb
za1d34110a4777c0cd3d40ee969f25429e189549f55e8fdcf77473e05e7aa2c603f9f28ceb1da6d
z95cf1ea955d5052f67269fbdefb4386067ce94ddf66e46a43515df32b4ce4c0ead13f4bc393c26
zbe24839c9be2f4ce8c6ffbbb5e96de9482cd7ac68655652c8868dac03c9177fd7afe6ee1b95cac
z13a661df9cc2eaeca0e682163960c320f01193d21a8e7c772678b1c07a82434d0028766db7447f
z4c2528bfd965647685c71d8e1b892741a9469b7c98b2d493d33f77b6b82391ea762d9cf047b3c3
zab12fd007770b83286f3a1d16f83b6e5d17f48e46896d089e3f7074d027a7457cfe588f2c63621
z9369b43b55f3c64fdb2ac2f49a78e9e94b6949a361bda9ada3b6e58f15ee8353e625cde051ad99
z1cdf019b3eac2b29b9486c4452f8a89e417e12c5d4ea7108b0cb3544a17b5bf9a71eeb81b8d3d2
zc8cc86a7e7bd863982beb6e418863b0bd34327006c41d95526de26f00cd57946897854bcb08a74
z77eee6f5f193e3bf9e91e3ecd105a37e8eb4a0f83b7d38cc80563fd90328efc2084f106c74b54e
z9f1d36f855cbbd8439c40d91560ceb5ba945b747d6d5f55f075538ea6c5c931fd711b7f80a5d8b
z615e318db172080dfe45534870bd82b7baa4853158848a794597f13f276cfb1f7d4b10b5e3137c
za87c20670f692c061d0dfdfe3bc132ccda9df0f0c72b88b20781487691a6529bd505e8d8dd5780
za40bf241b658388a58aedaa92808cf93c55bba548dbfd371f3fc96612be4d0ee7e11448a389f32
z31cb78f1b669bcb84a1690c34e7bd1981fd3c20a351c6f2943d0778c1e65e5255b7f76e7fd26b1
z742fd667f38bb446f50d306a36ff969da4db068612191d0d618b65631497e88eaf74c97a33f4c4
z3e4267158151b6546cd8fbbaa1eddfef472db2987c06862d89a76749e63cc1edce28ca61637863
z86d3085fdab2c4b677391b2d45fd58af08884a1ef8f507feedaeb15c57a7cd9d6ebaab6728dad6
z9d4afeae5c1b1b1e190c58e8cabbd047a5b4fd92c007cae928aca828c957221517c0a196f1d7b1
zad17b16c9db57846b266554e6c4bfc2bba9d0f959d3b77ccb4af228f93212aa099c5afd6e8c272
z2a1b133af1b3519c5f3b764d170c8a4af94fe58f184a1bbde5c67cca897a5a7ecefc370484d793
z53174b4fa05135149aadb2699d32565e468e0813a114e0a07d8113fb0c103f426a42f7f36556b4
z520cb51e08d4e91a6c1475ac49892403d351b0951d2d29733a89c6f89596e48779c6ca5172541c
zbba6d91f1c63b63554de55ae63509083f0cca8724799387c99ca1a7eef576ee1874ae401b62140
z6580d2079c3969065f58730f18368743b9d9d52d84a2cf54a201e59903ddc25e46416d795ab4c1
za04ebc3c78874710046619725645615cd4062636e8d560b3e6183b7cb0b052170adfdb965411b8
z7e2792bd5ba25504207a233bc0cae8fccbf30bf223311f623a4a7281fe08170b8212f3726282ca
z0f0b3384be10a967079da436e4aa053fba6bc3b976128455185d2c73e9f3808ee0da1f85ab9835
zff8b3fba2a7762681c0d80beb0300a991f94e55aeb2554174f5b83f67ea95caa3b88d82f8eb051
z242c581fb1158373649bff718be4e3c787914aa910fb646be37caeb52423c218a3f6c032a533b9
zbb4df978798b7302f5f26861126c1fd52600e258c68a916632ac05b315de25fb7971d713167ee3
ze08ad65e224fd62d7d290d07850c153eab4585334ed8c1199bbc88b1a7a92b75448b0556e8047b
z8a852f942fb0cbcc30f1716edbf6e6caf8b3d443aaef2bdaf94d53f8180256e6b95de103b963a7
za86aae38ed90ea968e339502d76f4276275b350494b7935350ba4bdceeaaa40c48200ad0a6ab4b
z8ffb05cf29ceee4052f29bcf1fb0d1e311abfe344d86dcae66b9902d93e43be0b8fe5b00741037
ze748582720b245ede14c304fb4a212675bbc692daf340a5787ce46abffad1a054032e6a01138b9
z991132e97a16608afebe4d131afd1260dca3b54696e4cd9ea535f3c97f600e351ffc580b8c37d1
zb60db755813c0dabd7f572f05dad82b63fd6cebe9af90418f598c39837659b58c454d2fea84850
z33ba6b7809f73932668339522381a445b1bab6e723a484c59f2ebd28dc4a59a214e3ae92bb3106
zea6a89064f2fbe29b787f3b8db07710ec21a07f21ce502d99232cbec31e4fe5810d41e46a6c57c
z0f65d42846c771612975a6a37788509b5a4f687bd0f915f7b0069c703563f4efac05b9d7bf66fd
zb9741c1f2ccf6d8ac74d78308aa74e5f60744ebc20a8af342d20ea0032906ba15ad28023a6346d
zd79c155e139b6a325015a64cce147a4fd5ab644ec6b554dc23fd52281934832a11b69da6c1be9a
z82e38f3b7abbda94f60f8fe78a28c24b3e924d98e6c4f78e709b241d9acfd09c2e77aa85652624
z0bfe79c3309aa7f2ac08b3dda981d5be0e39a3a527ff018dd0bafc252b09b70ed67415f5592c34
zd0daa54b986d07182565938c5ae3f94eaa7de4bcd472bb0a5ca54b9015b508698fa116cb0609cc
z71e816d3ae58a19928139fd354739c69a69e885b94b9bf24830b3cccb479b084c78b257c804932
z7b3b8e7e64c4d4c6e05b37c5cc0afaf32208c43373c0fc7bbb34b84fe718d0df8e0f27101de1f5
ze5e5b0c8f41cbd907ec3f6449bf10bd684a4f1e612364503669255e0438bdd03909b1100977ed8
z5c7a3b20cdc882244ae275bfbfc952db0faf25d30df0869fea41882087053df1a84b73a90da8ea
zd915321b1a6d8e5f6cb57e8a16cb9f555db2f85fe2a126da0da0835c02fa26b0d3eb9fd233bab0
z0b591c9294446685177fffc6df2045d1654e71fe447ba0c67654be5a9f7bea59d7548c1e0c0d81
zaea156ca150ca179a5e1bcb4a85e8d65e22c4104f35344a811e990b41ea9e27254bc20f75d6d2e
zb2fbc872035a2e71f90ed3cd8ece65898ddaff7c0823294f8c175faad93228eb53df2f65e7ca1f
z93f879a1eef6cbd6a17d1c44fec63d31a197dd6bb0ac006252c2449c1a21c02f1003876cd615ea
z83cdaf82a84397d4789e847af747632e134ce2a9ad64ba1b0fc8678c4f7ff7e1c23919f62a4ee8
z49b8abdf48a33fc135eb997c7cf89141aa09637a342163043524840c3997077d6f4abead5417a6
z2e1ae6fecd4a02b6d89f3780c7fc405da41234781aa705851c4fb832cf6ee0b9ac17a2cbe9eda0
z3f34caecb085aa23e130bccfc2c404f73b3e48fb554b71d163b010bc9ef08bf03e0c55f8e90f24
z8c2c7a768eafead3015ec11dc8c152080daabc7979923b83f1b13c0c6a5f8fa82b120d2056ae2a
z39c29bb4d4dc6bd5684d818ec119d3d1f11a0a49bd9370d47f5e838c3a8fe1e015a45586bbd0c4
zb0ac91a0d237a4306458ac1685169dda44610bd07d122713d6025b42fb8d51bd017d4217269310
z7727cdafb324bf3b6daa1a888113c1e115927a16a57ffa9446aca107d57d53ef931c68a41f9bf6
zfac846112e91492038e6a05d60407964500a3169373e8afbf15a036a6053b052ea8b0465b00cf3
zac76b21d721dc3df99b7fb42faca5486b0e67651825d8e1954b2e24ba3b2b496aaf7bdb541a0e8
zd8067012131db1b815053335f982b623b214ed8965976373b04950754fc7d68dcbe0552783c8f8
z6d88a7f4fda91cc5ebf8766ed04cba52b3b0f007e61fa13f46608b19916d3b3118d447ec5402f6
z025aad6c155a647db597fe1ef2f089b1f1a96b245f0bc40a03fa72f0570c8014241c6a2ab0db39
zd32fa39dc95a6a02cb4b69e8e1784523fdcd0448344739a2def09ffd9e4071e43595a452fa80cc
z91e9156650d72f0180aec45ecb7b432e2deb3b629a0f8b79b3310e3dd6cd87f677dfc376c00c23
zd61b4f06edfbc1685207097c8e107b18ad3c5c22319d5235275787445c1c86715f8bd938dc131e
z48256b0cca060075f84aa7bc4de76258b35505ec885809797954a20e4f20263a03ac6c3d38b60a
z29d84851f676934df404eb76a2f57d7856a4790d76f9f08a49745800203d2ee96eee8ad67c8b03
zbe53b29479bd43220dcef09d3e62bd4eca13ff20adc1a92f3e89e86e7c855e732781e80a0a7c66
zf52d5c716a98f73680377e6d65bfc535e2f8ea8f073311e0f702503fbb6b1f13f7ccb3674a1a66
z537eb8e5d02054a0260808c05560d0fd357f8fbcf40d8d6bb21da5b60d663e0cd3bf729fda9d40
z85e548e24e0246423075222ea55d0763e885ee43c2dbee38b7021225e0dd031a283da65187508f
z54fc4ea235931db12f954c3c9dfc589158ceea8d2403e0efec744e9d180aad50bb8493ee8f3031
z565c8920389be57970a3c7bc9818c199517e14cae12632356ae802a07dc9cd886dad06770e7b36
z43335783b09005a58a94ce7ea2868d58915aa265e82d53527529d859add74ac10ac57f4712d6d7
z9761c83274900d6c76ea785f498d14ef96734fcc0a897b781dc2cbefe0723af45b20d9af18b615
z0d0f4f370f068f01dd759fe65f6a149290bfa41399b27ff51a6113df41b98bf24327b8fa760f2e
zfaf8a0d5c36e432dd743c421c3744e172dc7c558bc6b73a782538f05b634f6a747ae813be40fc9
zaed0bffb0369f3bc1cff778cbd7b64f410f437a04371f9d5980e28d01dcc6f2085dc420098e04a
z0f0b6e14faf63cf29dd7f6b5cd9860a4d31ff5c49461f39009b50e8644f35a241c46d74ee3586f
ze7b477f0546bb444df8ed0358cdd7d0f9215ad7bcfbd06c5d6c030e024a6e847e93fc98aef3a7d
ze0faa271a4c44d3d0edfe9dea7e974c6f9d8db2beaa0bb5ee6a18fc00294d0bfcb3d7c0b2861c7
zd4018f034e9f701f57b5cc7c61e12118b62e614a905454edbb676e27c79b6fe242094d96b81005
z1b7605d4c9c3dec28426b6ebf8e2f2466d2ae4787efae1cf634c1c853619e6986990250e17b9f2
zbd6145df9d7aba68c810bcdc8ccb3c7f907ebacc5e0b95f288e120a0864ac5f1cbbc5f42a6d054
z290e2cfd1a7487992dcae06c0eb8b5616a081773d827d2a3ece9159635d19caf8a7d66d2dd4597
zfd8556d2293374560ca26ba426afc84027b7875f0c196bdcadea2af991a3c1fb77c4e2be3ec76c
z8c4c06084c9f8e47c2686fcdd5d1cf282c4920736e5134144473735fc53261e33cd252e0b6c86a
zff18c59e68e2652a4f5ad857a3f2498867011e92b4e463e9283f16dd2749f2826dfe41ae43366d
z833b4c3faca1df841d432fcdcf5bceb30157003b56dac97b873a53d03d99dcb50a3a41732f24c9
z484f33ae1304bf4d5a8f251d94315e5d36f7798b1988338256558474c8bd7db721b287ae6c35d5
z355bcf7272e30bcdf9fbb87fe87b80997cf78d3661ffe87741d911260c5933e3e99efc2e7964bb
z7f4c07346cfe729bfc6f31d93038733f566895ad20b4ba9cda5c555a1a21c1178f137766327173
z3e591924139b0665fc9d48740a36d7527b45ea41fb58c31b3b1868a9fe8fc38dcf1a21ce1fd681
z629b87eb7ff251b09cb66f2a2e2954336b19fa99f97ade00c263ea9777ab86282798ecec32710b
z8f69da4b0f5dc67db79ca706364350a166497407975b033e58ceee29a377c2aa04816caa025b53
z5c892fc10c30308e0a4439b800f0750c6afa027459201b2489f8f451d0af63561b4e182e7b367c
zf9b68db4a28641a5dc7cce1177baf7c8e9ce986416b197ee3a7b037adc5d585630ec4bedf163f6
z80cc09a5cd3c2e5e3921176f15db9c6336f1102958b6a4291e6da67816965e6f72b30a5e372b02
z25a06131c80342d5df7fd27e80913910a5ac8309807a3aabafcce0d9fe111fa8f20222465d1e3e
z78e726a03d0ec9d701c6a56ca783c6612488d1553be1f28e6f127e79545f3bdef031519c86a562
za3f7fdbc0e8db8920c9b0f497e42cf07deaafb3df9ee28277c4a57f9751b9ec370589a198fd8fb
z1e2eead908f7b420bc2773ac22d3180627583d57c1236bb9e24258a9e2c50237aae0aa14c63a45
z6eab0eedcfa61eb23fdf95c8a5541d68aea4373b11b20b1d31db1c399af7c10ac25ba3743e5f56
za6bf64e9d4fa7cc713445d801cb0b6888628dbae5b2ab073358b2607a5199af41d4538fb419f08
z46e75bea59159fef98f2993a453349dafbddc486c1bade7aaa46edf58ff43312c5849f29f11eb1
zaba90737d3d407715ca5ee0f9e8d26edfc508cebfdaf4e672930efec966e12269d314489447a78
z4ba0325228b0bfb31a8fcb7cf714d21dfa6c892c2b3ac4d840313807f4bcc36606ab0abd4d647a
z972d9c04e56f38f1a608c9ef1b94743625c6eef61e9cdc36f57ce13df2b186b2d00ffd093adce3
z3e64301be04c75b056b6d394158f88ca2e2dffed495bddff45055452f2441866e91011def524bb
z08b1f6ea9594f6c50b31e235adae95bda64a843a3bad868a14ef91023d5d0fd58b70c8a491a559
z9cf480aaef46b4b705628c881a43e7f5c8f2fbc2d4c6ef98596747533a7817e0cbbdfa38f668d3
zd1f5e2d4a160dda063273ca59ba49309b338306c734f481c0e0220f0e92d7b289de5aaaa847694
zdc0dd86cbd9923709d043f2d75f93451610d705d96dfe6210267a82688c6418fb889188656cc8e
zf2d4255091aec86efae41c666cc9a05a7674f74fdd7fbcdd067f9749dbe8edf17307c88ce5d30e
z01be06b269d5b737e05f9b853d516c688ba9abeaf9550629a534b99e2a020e9463c416d5d85bcd
z489bc0fb27fbc0ae9e077fa490ad1fb961d71d4c8765f54cadfaa532287d9e839e2d85410ebe83
z93b8f23c915a51af87c858dd8f1ab169a26d2d32c2763fc955d1e5380891ab0e0b1b4414fcfc0d
zdb31fd2df96aa312bd36ac7abc25c6881fc79a95abbf06687bcf118fabe71b44263470044a321b
z180cbc649fa562eaa0e6f0142ae3dce4f908d8169e2dd7a64781e425563b17f0d15ea70a1e3f13
zd32b0412bac602fa1554cd385ad72bb4db8b4d335f18e298eaf26464805ad0db32b89ccf78b1de
z1f408037767d6b6028131ee73ee9b5b905fbe18e1ad4c91f859889737830df7824d58ecd82201a
z3ff921456c6f500a3419645f524cf5aa17ff09e46b31afbb3583b487c4fc44fe945c39c89db3c8
z8ba00f8895fe30cb110237eecb4a8a9627e9c92591f5f516f0242c1a8c2c2da11b8d3078653330
zd5b50314e04a44a17a679c7bd967d2bb6fccbdc9e9ec387dda4842517d78d09acd49e62afcfd8f
z22b1875e70fb35b3460262984fc01df9df51c87fff6a277178087486de90eff678ab266231849d
z274367527ecfa2f9bdaa746619510063966300e7dfe3a3fc6691ede27545366af8090c6083fa49
z4ba9c23c6f2e5e7a8af00f3a301534db7cf6d29b7bdc0bb0c58a152def2bacee3a5339e22b6791
z9022dd5a36166a8787164b4a55f6cea75b15ab92b49cdea377cbc2cd6b6deaeaa359068bb5e096
zbe1c5d18d0189ddb6e2b1a6758b9977a11ac7d71232c1b840dcd17b5b5490eec7472c96fdde25c
ze5a9c15228f9cf37ca5dde0012b93dac5725f934fc066a5a3d85284fc7fffd76d248f2cb14e493
z4d4ea10b3eab6f098cfec4b6f50535065cc2a4863416f6c9593444daa092daa241637eacd14408
zb0282421a62f1d3a455fa40e60dcf78994ff5eb99a2eaf40afd7f00cbcde4d7137ed63969f6f3c
zcc5923f4967196dd9fdf102cddc97b27b572ceedfa821993560e7c9e9c5854c6b4610396540763
zf02e5617de6f0e8b37a7606473fbc2735ae38457a83250b0e0dd8687932f238f21c95f7f89eec7
z9e7f08619dd590f1740cb3af9a2ed7524674f38ed77df24470c8dac02e6da0c07b2b664f82508b
z8b1540ebe5e910f4c3e6efb6855ec88868d5bb654e6922166a790908fa5ecdca00a4071a3612a6
z8300969a7fa1afbbaa852754c81314ece4d042c237c1a656464c8d5c3084c5055c1e25bd87e1e5
z234d84e17e6dbe7432a8194f08e8dc52349f666fc1a07d8c506c1efe89d1c0d37115fa41392da4
zca1c393a80b3d3001a71333d2bf4d70496a34c67278452d1cba61064035cec5df86ec7f96834cf
z663a35a3231b4402d776fda695149d6cfdf553a1a30e194a7e0a8f88ca4763bb085cd2bb31dc82
z1f8d05376e4f9ac2069b6acd88eac57586059d5ce8133732ca227a9fe4a275c390bf1659017341
z07eca1babe979ad131f9596d852bf24f425f452963e5a1f9a96d4750ac41509e67fe9aa0e67761
zb56625b25b6da933497d87ff9d754c26ff21abd2e7659bff6e01216726008b84185bda3bcee644
z2b8f5eed60810f49d4ffaa44a07f70c5a0b34d90dbdbc4e322bbaf312a198da04dc5d1a38dfe95
z1cdf42dbd0fafbfd456cc4866d2cc51410c056dfafbf3bb9f86ca544a87a876fa687a237abf995
z2399866fa61ff7d9129856ae6b0f774f3c024d62af4984048d0b46cca69dc074aa5a7aa5a5b73f
zfed1dabae7bbdf081cc7ae9bb4b519f1cff150d7734e8c3b63d4fbca10e9bca79d17f20abe5e5f
ze3962f5898462b3cd7b5252ba03c083d42d8c25b083edf61c0a9706944e67c037bb037cfd4f45c
zad28742a2d1669d94d73c75525fd2e856be0c95e9e131885054640125c0a9c0d0398cbf0b53c17
z6e292362fce910cc248fb05d3ac3e195dcfdeabfe1a97703df8ce46c5707b6eaeb7140026e3fca
zbe059ef286d4a3ae5bd7fd2cf960633875179b8fceccf5f049aab7764897c9b58d84bc6cc0ff4c
z6fa71fa07f97361d01319d8a266d04d3bde5472f85c8f8f27442c50f07e28b2a07c521469d6643
zd2002a8ab5d4e11692bc8c6f8b510539969ff957a4f36202935c733eecbc2c6aade387efed279a
zc28271f04c89aea2ba36b1a4014957d511f26cf40d3fc7760c4ba585801ce97258af1d1b1343b0
z6e32c488bde955dc1b5036135e95121aa384121e1fb82793c8fdfdb4983df75eee4e14364dc830
z828354c1599fd5c6cae306348b26c1f21a2eb0a1a1c76e6e35d6b2ba23f3636196d774b972171c
z5e003b4e072cb33c54ea5a35afb57fa7c0030d9dd0d745ef4eeb4ebbeb1290f738884927ed3ef7
z7bc6a7a26dc02a8186fc01758fa2e4b684bd8e3b971fc0ca6f39b21d955905c61cbe70b441eec9
zadacc11da3866b496765914837ee6ef8d0f92535a690b47d980cc1a66136e53a32cc6191775e9c
z6a91983132aff9d2e8fd3361d37301909386a9df98dd910078688ca12472661015aadf6f27687f
z58914327258880f1c27c924fce229174bf903f0a131fa7ca287cf2d6583c7f975ef95698a65839
z456cc350a7e528d4e1e76a559cee7ba8a420e75cd071e6c0bb069d12b552031174b3f4180714de
zfedb3916777ebf3fe2acd5277a6cd339aec74610103377c780e609e462291eed8e5be27fe02a4a
zbbb7288b28dbcdfcdefc6187ec87439c186a3b5624831fb3adc6b1be14450a848e053a228e2569
z41e250669b39bd7adfe75f14615f4fa05dfe891239c1248e0e518cda6bc75c2fca42654e2588c9
z050ee71e278f21f163cfa6eca927f496152d443f22a9b8a0123ad1190d0b11bad071d31ea2d648
zd1deda3ef7833cfc02e5c0ebf7fa9146fc4dd5ce93badfab8a93eb09234ddc7bac2049f75b44a8
ze70f59ec6e71d82c9e9015b770428e42cb99aa48d1a3c027ec108b1c9fa0e1ee96678c554024c3
ze8419b2c29e54c4c83bc7fb3bab01b095277fc730d81e069c2c342d0d8759db358f653fb359bf9
z12cdf921d4fbcc10396e7078bdf57c50cfa9da5c6c9752b6b9b962aba0a68c10a518c4d9313b56
z8ab02bdc84c5cd497f46a546e16fb574ba9860fd1a0c4561ec61df658d0d585139ba2da682aefa
zc9321f98d770ef26e9392d377876b1e9891483b857b1b61088dfe51987d80987c3c094decbe23c
zd65975e644b9f601e030d5207960dc5d3c0adc8f7cf013b0389f16e0334d5d9b6acdd1f6551022
zbf3939f66ab70cffa3f38aa2ce54dba472aa97862095a328ebdf502ba76f06a06b2fb583a736eb
zd3b18b3b940e25046867aa2ff39c52135cd3f0fd479850714966a6cf5a3f894f1d43dc542c5b2b
z3533b426bc319a286ca8f286a5b6132bcbe159e3ec06126e2ee4028717e202e901a1b7f2b14331
zbbce6278b8f2b277d5ec0ed8ca47e2ae11247d0492cefb9a9fa7456da31f26232c807cbc750fc3
z7ad6743d7a4569d4ab70d64dd509dd04abe24869cde0d021bd1467ac04da6a08edcb9f6006c86e
zd9b73db761f636359f3f57802b0e262ee0dd2fead5861d268e9c142341d5d6f4ddc8e48ee3e445
z7a3a4ca3d6e02f648c970b5ac0bb79079ad0eaf2acdb5b3f556a75f0ba63c4a5eb5c4f33ca5c2a
z8d1f9b45b9ff6eb0ad8829b87d5664352f91d2501c5dc9e98c135eb2cfdada3bed1e3581a1c3e0
z1e828ccabaee73ee6b82556eed46d58123d23c8589536482b0ee66d17db6db262def2b0d16fa2e
z92f7a3584a476cd3cab3e4a52a936ab27d5d339d5887e19a357ebb74c616d48f96204ddad55880
zdbc014071e6a798021ade0d0fd635e147d29d3e3fb9c18142ebe1224812298708137c48b98643e
z0bfa7fc528f30efdbe1d20df0173b862d2ae069fb30abffa7372309cdb2be5bda1b42519f9008b
z73ed0dfea47595124d184dc1f52fd6289d5afe47e3e98d4588dfaa3e5ec09875b87190f941dda7
z88cfafdd9dff7ea78ae6f0a12e9220f1751ffb9b0c70dd00a1f26f0cea42ddd6e67b5b8a09d76a
zaa81c6755d34ce05632207a80d639ae3b64fdc8fbddaf994543fa52402f987fe4ab6c0c5d9b7b8
z45471b857f246276ee88f445efc9d1163e5d4b04d8add5e948f57405b65155241d9657d175fda3
ze3fc3d2ddca664050fb6c561b0adfe69adce216c85740a870ea06f35e43ca250ede5b61a62f635
z3d8a413fe829e4443937655aa74f64adfd29f5d55650711b7a6281b1e9be09511346f603605887
z7932c1552d237cf99efc79903b6bebd6c5e1f82e2805ec90d060133728a064e8d6508180994e30
z837a3408150377a16caad8b8c8639f3913da1c1ed8dd898308b6e2ed9b289693664120983117dd
zd70e2fa01ade58ad673d18039fb533088c53ba13e3835a4045eb7ee09bca82a54de44a88f77cf2
z7b034baf13d9d4bb07139177762b328ff1ec913dc881040e2e73a5b9f228d2239195fd9d9f27da
zbc650b3a95c820514c62801eb071199db5a018128b3ec570daf4c85b4f69d8e23a574b93468d29
zc4471109e5dd4dfb648e0eb159970d75714e320132e78915c946c093d010997461cba5e778b25f
z75ec346c13273e6d9a17f592bcf9888ddb008f5136f320051e099985391f9efd0ae386552f0a3d
zd8bb8d565f8d5c8588c1379d0df96eaa3066494b678ee97a0ebe8abd13f762a60176f83e3405d7
zceb06fea5808816c8b403cab27ed9e6d061198a71ba4bb18e886111ab868530c76fd9d2bf3a071
zf749cf02d508c250876c9852685140654e56730dd9f1987608cb0a285335fd49f13ed718b766aa
z00edbab37b449539db5623c861cdda5b236cf9ff28494f01389708e14810b0c30894f805c012d5
za556671ee185c5b76b61af9fbb7e6b590a1e3e2ab4fdfc7900e76d1726468a93434e6d55a9a06c
zd747d324f5be884b16d9f5570576e13594efef5374c139f3ac3ca3bfa5f243e02c31caf4249246
z4ed147a486c788aab6382aee5496bdc0d10eef219bf1e9bd4a8d03c70de7ab2ae4174e714e9878
z3d7984add3010cb08ef66ed14be1bc11121ff460b584c122b56a0db5ab51e8a88209f35e63172c
z2d3bc092a14f394799c3b38bed8f8273959a12a0d54617242ceca3caf7e5ca98f352061d6291ae
z8777f62cff8c7c65b08f3652c328729a4259a086b356659c0789851e1b819efa03a82d2ca64ca1
z946fa089b396294a56d36d38b6edbc87666093d2871eaac539637372ef52202c68b945012e829e
zf49dc41b5aafe19d4a8cdefccf83a79edbb417a0ae9df3bf0007b1cce1a4158a8283c2f7504cad
z54349802ebd7f603d75ea78d9c3fe0467ca301b14c63fe0cab21f58686259305282471d221c6eb
z81a7b1258bd70911be41088045b84ba85e174cd2fecb76a9abbf1282131379605c097c4d063e9e
z8ade1f0997f89ebe8721d812376c12d5c34948ed37c7ec9a124a599d4a3961299dc0cf3d12775b
zbdf19bcdb557dea7ba73d2f7f004634cdb7edd353e5a034356096552f849e6e632deb05e1fd194
z4707ef7f99142117eff83c01a9fcae262a212e5fba2ee5a819704e0790bbe83dfe114aa89f450c
zcd90e410b351348e6ae596c1b087a261da9f3e4ec9522ee893d99cb7602a7c8f4a02a0d8ef70dd
za1020a81c2a2d4a7410d18d4b444eaa616b0d5af6bb26bb9ad96d16f422fa88bc6a6e208ef1a05
z6d57638eb665cc608c29f18904f4f0ebd83e03cdd01851c529b354f18be2040648b0a92d00a47d
z9e5a4ee64c889d18735e4b1e2a1bc396a0c89c93e5a6d125c5850450981369e1b86a2262010f7f
zd9dc40e29989a5f25e64e9e62182ba0c289a06a56bb6a085b6270ba707d54f0cea00ae20795c50
zcf02176cc2f5ae638bf81999db345d7f382a7a70ddb90bb0dac12ad656c56e7ab721ef6ba98f02
zf51c3b0f22b7182cc25888edbec83098d5988dbc87fbff7bf5d01db61defe5463b690b2723e2f4
z7fc27922f717c0b5994cf4eb85dea89ec733b65283fa3785e9e9ca25bc99846b3c73e22935c8dd
zc12e45ec0227d1a3f5dacfb16cd87c6022658274e5c4f842beed58ff9c46e1184cb1427025c330
z5cbab40ca3710687b872286275db62af75fb472a79b701762855e98aa4bc8354e24d6025517bf8
z16949ba9c6edf1aa04c682ee9794599443511e7111157dbf67b781eec63d43abecb71d2835eb68
z8425ca7292cd4dd8da659add04bbe644e928069e13936c3ac6
`end_protected_0in
`else
`ifdef MODEL_TECH
`include "qvl_pci_express_statistics.mti.svp"
`endif // MODEL_TECH
`endif // encrypted_0in
