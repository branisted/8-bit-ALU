`ifdef encrypted_0in
`protected_0in
ze74c34e226135848fe16db9ffd31815111b6d7fb642c521a3f628cf6da949865580b22efd062a7
ze90adae0e65e66a2c36a587d0a790699161455169ed55a01f2084f11770a774ec4c588039b380f
z6de9c5084882a40b79a175f5c2114b2b6d78b070cb806e1c0aa9258297f4687ab308bc470f0040
zb0b1de382961eeeaf2e279e1462520fc31c119af8f2b214846f56c2b3cd2eadbe4099496abff18
z15cec83ec4a77b868344aa20ba7360908f5c0de2a79abf8b3534b883bb12180f68b5d4beb444cf
z3fba8f13afb0abfe8fcc4294810f75afe452434d2d0f1166236c82f76edf1e12979f04bc35693e
z32ae028996dd85737a8f5adc1ebb94f39c940246e887647b64782cd7ab429b0544c173176cede7
z01dfb26b1f73408344a52b7e1f117f12bb9c8077b34876c2e6fdc085981637012dc9754765e1a9
zc512ce062e0b8fb16a214591f5c81e1353b900a611fe1f4886b57940b41b7f2ce99a7b84b04b90
z916f717e73bd10589c81e207ed77ec660a8cbed5b487fa50acde1b055c8870bd8676023f21ddcf
z9c98cc47cfa2d654ff1365d1f45035a045a66c5dfa8279050262529d2cac9e64fd27d9c7de62a7
z731bc808811ded9016570962244887f98fe5440167bd0088f2f049df882af501358497c3b28776
zcdc5426c7f52a851c35106bb93e16fff984784050fc808fad15da3306022d17da80d857bd32a53
z2ebc5737d466752dcf94171cd2cf105efa9c502d8d409200a8150244f03fba3a90bc8d5cf172ea
zadcf57f1aaf8cacc562c30d11230bfd4b456201e0488a1919517c8f4390b2a7a4b4b904dea5234
zc5fabe55b24358240562a4a4c3748d32e0a62d645c18703f0800adffddfbc1331e52ce31a92020
z0a11b00cc7a32d9cd8fcc96d850d6a7afafb0ff7b8dd5522938e682b6a6ef1ff504fb5dad69334
z247185f9503621dabbf693751f563e1eaf5527c14dc63cf6be2c35a203c34e03f8c8ca92056016
z889f604b3249950f0e5f3edfe116426da88d520d4ebf4181782a48ab23fa938bdf7588f9a30626
z22770d94031ec8c19d7029fcbc912962d6298796d42f87937f611a2e46eccde544622a924bd54e
za87cb737e49e1147a3683efd62056fa2fb31390f4e4349591a864f1298b32227ce7652c5226e37
z4db97b8cb0c346a2bd029ea81f3e26a63c4f2c8b09c802817db4d59a77dd84cfc4fec6a51c395a
z49d6940fe4a63f6fe2b5a1e77c53be40eee7261955299fc1880ba33c88905a260bdbd1cfccdb60
z0c4892820281521a45047932cea3aa7930ac38cf370cc9a3aed4bc6df2fbf4c2cf976591dff154
zba0d4c6c332ab6927d21db92426dae8cc6fc42c1297d14c609411f8cdba90c44f39c1b06abbd4f
z886bdfe075bb8cc19ee0df2d935037aa2d975a35da011ad652ab634c5f1418b7be7137aafc6fd0
z86bbdf36116deea5f683efc359f21a47b7ad383b8bef4e64bda0a28a529561ef7e55eacee59291
zbdd280d2fc2c9c4c7c359862566920ad88f7a547a934638e0a3f4ace20412ed10ce31964506ce0
zb40043e254983838d122295620f3113ea54f737b6673078bbd06635fede885c42940b3338e32f8
zfe1f731a924e0747372e695c62fdd39b6684a997fa75a9ed321bf0eb015cc6b5795daf3ef7c3f0
z618b4da466316a6455fd2ae3c44fd201d228fda1ab4fb1de70a0d39dd13213b2a7dcc049adb12b
z2d3ac36047a0d08d78dedf9986f9ae25a455577d49c76c6442791bea325a6d2c66dac96ffb0867
zdab7a6d25ebbb93163f40e791e6f4ab91300fe5cb7c5cf2c1515b02bc68f0b91c5f56ef045cf6c
z63de72155c8ee1ed388f91310038c3e93eb80f4b19ae88b67da3a27c0660b5ce08232c61fe4230
z89152232b268fd170bf9c46867567e0b1cb13bec7dec5cd93daa0ab437a32502b3ed8034e168e2
z1271ecaadca9dbd7ebfeb3d8a1ac6727de1e9db83ec81951f2c5412226df049c8e71d81b594529
z9c90487cc084b36726f681c2e37334e00134e9c72fa9d5790aa614d2851d34717f6ba6339fcebf
z97e18412364e3a71faebb0a230a2fc5c245cd63ce35c194ac60eaa173d0c30b85cfd1e2d8cf539
zb035408fe9179f37cb8ace35a98f15314e10d93ffe69f82a17cd51b0cb10ff83af20dc77ef3276
za7797c31a26410578e82c227312f72d02f8e1b711052ec7933f0c9847bc9cd0c37bac4ce94752b
z73a878449e90974daca569aaf5ebb583a95ed220b8c91edcaf83e3c56cb72e78f2a577f025d358
za190ee94e42eef3337026f8b8692cc525421aa3734e384cf27e549ce350a7e96811aa9e2099b14
z4dcb770fc6ccd9fbeff6dd343344e946814e4afeb5366587fb4159307868ea028b7badea3f87d8
z840b72f7c2c93e51dccb645fa26811d3a45cbd1b0f91292ca941dc24dd5861bf1f792788a7b146
zc850d68800d45ff866722ee2f33a622e2c2e79252d46ce6628de13b783e59240c510939ea74c66
z94b612ecd93a2be9f14770933a848605b12ffc97281cf00a9b82898676feac472fe36607892daf
z1985b158084412e01da4692ba76f35d68a28299551fffd4e315475f3abd21e866547a8dd9403a1
z6e8e7c1215c376b66e341b43eedb27d5b40ce6799758b7d33d4f4895c915f3b968836d3930fd55
z1b22f0175e2bc2420e120639ee0c6dc8ed96d0bcbef27f73b616dbc9ec2ca5bd08615cc6aa1962
z555bddc9fa7906e7ce22a8a606a49d4f0f2b4ded9e5e3e78505b9095edbfeda732dfcf9cb2ba95
zbd54d488af64129dbf11eeb7b18fa9659264955e37ff52eae8984e52aa6ea472960cb52b69e3de
z42908fe67d6db1e2e8dd5be7db26662ca1ff13480240fdb96bfa55da4bdd1081a48079b422c6dd
z028c8a5b9fe75e12dd4f27d7c52fd33c10311499159c97dfb900594d519cabff65c309452fd99d
z7694d1e552a43e202a5ec7df138e09513358623fda30af91e7b09f54b2758368bf1e63f38bb1e0
z51a6812949af43191d4463011b1e77ead2bcedddd97a076ca7d15889200a9c1132005b111b842a
z0447e7f059df870416ae5f7b3679a5d5f39b7355cec03ddf0023f02e8291af3a3677c0965f3b58
z09ffcc4a31f99c5d3d5da773aafd0126314bd6960d8a1277c80f39efdea02312d909f3b1ba757a
z23ec57c68947271a2aa2ac5587cefbffc78f086e055014e33f68b7ae811fad99434be8e2f9f918
z3929ec8d1968ec21d49b44c7522f69296ce13d26f925b800207bf463eaa861976a5eeaba152135
z8c18bd775c2a5fe75ae78bd2350d1b18585c15119d31e7d292273968ea5f20d63caad35297b111
z1ded6da353d46620db048db0bf58a5e16b649d691c0563bff97812006b38e21210b9a220815195
z04d59c7513cd1e80ab77fb3de6dd00c968ec79a08a43a090bfc95b97d1630637be470d1d9fecd5
z6935f3ac776f497fb2fb7d2d6c17f16be99b159ba3f587d74a10b7d5bdad8962078a3610a835d1
z668ea8014b859fed717764ac6c6a4258dd5e79d82aa14345013cc2d6057ba1f782010f4f1b14ad
z5b4dc05945e1824607fc6238af5ec0d52d458dfba92f13eadb8da5a72301564771f125eccc0304
z78993408a8e3f79121264d92f713bd9d2217c891de4ea49ccbb6e54f760fa39b59a5ca45bda249
z5975e30440cf021cd495f948d6c9a5e81d4269f47e28df0a5ba09322fc282a7b1fb2c48386da2b
zed75ff32ef1ceebe55a3ea6957fe11b1518544a90676996827158a2df239fa1d544aecfd18d932
zc79318992f5439eb060cbeeb15626e2f6015cdaec9b3c674cafa0d473c5b90f40b82f352f21b2a
zb9232bde298d3136ee4394f49e1bc2ee03241b3b95958a7c92a0fc63a23100291edf53152fc1ca
zd4c30a6409b526985bd409afa1215e29fab154aa3fe3e363af50042eb480585d87922dbd2321b0
zbae40b19333d750be610ac798164682df3bb6aa7eb0bee3a391011b8edb16f60bc2b9c7e18bc66
z07cb7d95a4fe53e01078fed074732119dfa12cc86714575006bb023b2868ba198274778490cef6
za086d44dec559b9c8c1538f17beaa41b002a095443bf21a037b9f6c66501c2a8d06e77f95f94c4
z0934453eb6a794ea5c912228e59ca2a09cc3ea3082b0aeb7369727a10d5d67ae8532aadac89938
zf021c3a6def9c7c78b2dff6c82fc3d86dc22fc0d575c762128180f835a9f669a04593e89609c6e
z7c2caf8af2e5fe9e90e0ca227c5f5b1fa396c44162c35449d664f15c5836900eb6830cdba16525
z71e47476fe4fd38770ed21bf7fb6c13dfd02fb21ffeff836d9f3b700980d029144ee35e3065df4
z7c30654d78ac3559aa3ce654d4394b2c59f212f678c487488b57ce2d9e26c3d96ac23c3a46b25b
zd109309286cc1a1c692909a34111813b97b397ed40412d2705eb9a548a67a4687436e85b7a0b17
z6d0d72384ba78c1bdb68f64d51caaec947f8b9d275a9de6eab01fed2213fc875fd3cf9b71ad6cd
z85b258293db37bbf4ee85a974dceef640898ca13521855d24024f684cea5fd33c51674bd8a6a22
z4508bfa5dbc0e23f5bc55ae46a96c919767b5b389adc23bac7a799cf5d3cb468a025d367c54aaa
zb8d3566c5fc40634343e3801c2c11da70a552af58bfeb4ec4a055d211f28c1b4e86f8160e5155a
z35341eadc878a8338c34450126b889861c89a02b9cb742bdb95a32197e60728e1125473662aef3
z61dcc12c289092cd33bd258e8e0fc44e078be2d22f23997f126c90c125e7943734b568f7e1da99
z6b729a93f3fc58a844e413e30a35c28cbde52b977b660a949392e8d11f8acfd493b6c4554c1f64
z278558d4336622372b477cf39d4d8862ad82ce8ceaddb5c19eafe30201ce98a0a60a8293fb5590
zd7b26fc7eb879d97932e10785963c67ac152e22e7df34a9a2465a44002e147c0e7eef6322e0d60
za6d41e5a7649a86b7a64412306e07ad1d720840c309d37f13c1fb83e7f5da81d319da741de9d8f
z5f2c2489259507e1f7ef084ad8f1b277a65c8b0958978ca2f7cdd93e4ca6e7519d0cde278443fc
z0f944f1a53014624254b73a031cc99f9aa47a0a52880502b702e14e314eda948e931621026c60f
z725e9dce40703c33deb79817368d34bff7109e4cf00693b040fca9c96961a597c8deb60439fec6
zb81272d3cccca38d7dd0ce5f49edf85d0d07127c52c505c17bf39bc124dcf8eaed675461795796
z985c89cbae264ff1510158e132be6b1734a152ef2ad9a1c42b461b6c26b80f2d960dd2e113dd8f
z26855ca1f7862edd295ace3ada5e7538e97365fff20b09186fe127f1fb2e71f55e825d5b7a3851
zefcde2dc0c05d0339affb49aa1098df65d2d44aa00e4bf2d544afe039686e3639dc9ebe1ad0739
z716583f505e309f90ad372b5b636f1142bae81960f54dee5cbb3bf7bb0048912c1facd92f7ef94
z80d11227624b6210f7c51fbc1a1daaee6d74081715ee857f9410c9b50cc631fed805fb848c1760
z963d7d2ba01d800e59c3dc0cbdd478eca07049745700a6e2ce1a80dbbcbf869a3179c83a36b804
z3d242441c073c3e2a56a00d6f1a50003a117e28368d1489ef28917a95c1a7b0a917aff1fcb32a7
z121f5ca2075b8e07f4dbac0f4f48b944075a76d7023796fe205ecf64c36999f4cfe32aef760773
zcee1131e736b092707aff6978f0fd7372c8309eb264ff550b395488820130862452e23172d1e49
zab4de00cd509f9c0afc8cce833d76508c2d50f14e064768e240d6d1d561f2501b56f0f30c7fed2
z59c810b993d1cb9dbceae7b2062c89ee9d768d954d3f72d91b3a026fd2ee7df10f3bc2f1057831
zd391330b4ed69f64b9db0765e23ff5458e7ca642fcd9bcbcdcc2619b34425a85a8a01239b6893d
zc36b635654fa7888d28fd8e086c542d3def081bdd5ba84cb0bbcfe400e9622e8c1ffa6ad1e1365
z6d6dcba9dccc674e28e18833ad64bf82dfd714199bae8dd8100c799931156b7bcb607d773fadc6
z27c0e11f5895a00d00ceaf16b8c10890f2f55a4b158d6073882e8efc01dd9d84f43e7db882bd15
z5e764b18a1dd1d906d27e067519de59c69589e94a1f2f54555649bcaab971d9b9974520c04909a
ze4de13628125f018732a46f911403712db02b1e6772513d1b186634e1d1d6afdb84d38e952a91f
z2bc56a1b19707560c5012a7d60a2f8c020dcc7fb215c4f811f903467cdcdc38abf27d40af516a3
ze835919d54cee3711142803256be95207e231c1d14f8ed3515ad35a82eaad03634b069e22203ff
zb2fec0b9f137868d315645858c1180bec31afe6350fe78c6d92ddf112c662bf57ba8a650171169
z96b309c135b1c4ac586bbd4339602b94a9071f4ed5a1a974d38fba3bfdf155db6fc9c4dea04e5f
zfc328989fc00aa1d159aedd1b216af08e8da7d41839299a0b3cebad9335a880503e2c73d57c6fb
z0bab15112103b3da72d68326cb82c5dd0098495dff81fab1ea27aa602fe7d5cdc185f79e483ac6
z819c2305bc7275c7788644cca8fa317292d57b224de1f3ca18848e70701531c205f87a1516f7e3
z7bd692b1cfbb33dc03cea8dd87d6a0230cfa033bac075c977fe75fcd1eccb0fbb17b69fd474410
z562f51f34aa28f3a3b91e0d34d312f68c3fc7dac069d9e5fcccf27a7050a1cd953ea795abd1b1a
z3c6626fe4935ce5a9ea9ff03515923d254d0803ba1584e490eb5ab413c7607cb45fe9130c1dc54
z7946d552a87b66d6f31abf381fc89b9c27f0b84e128fb906fb44e65ac72d31c55d82ab0dc4d87b
z252acbe49883053750cabf175f9418e27e197152f03acd307ea72b9a62399072d308c0d720df48
zf2e45889ab3cc0a2ce73cedb8dd141a710c3ed6f03cb8e1f3547291566e7c9648324dd0b36712e
za612278e3b2bf893f0baf4a1d8c6a90436f8c41e1f9a965e19f2f0a19296363bb293fa0dd4c8be
zd3d4516b5542f3c56048315229d10bf78e14d2e6d5ea6f8b14d3798553875d3e97acb5c2e6be66
zbe2d35b8653fd5033a5dd528a5ca5f0d1970dc677ada7debcfe91998fac821ffb894dd12903f18
z01d064b2233d56e7e3a7adfbbadadd5d1d57355eec0377f7577cccd2e0f7aae6355e1199a90a6b
ze0c634b285d9e72a674dc671a6a684c17209481812ca5a711dc16937ff9e105f3fc92db27938ad
z37a2c29a075fc36de65129c49990248a3934298bec81b39c94fff4fab9f9a98ddb0ea43c724026
z198b4414658442c850d128bb92731ae923bec156d1098dd672346fc55336391f21ec9e9cd4f8bb
z51a6354840652610722b2675e93e9550f4c627adf3314a13069e6ea2d6c292e3b959d280fa2ac2
zf1ab70fe411fee29c987c8f2589c486d9d37b591ebc87a1db938f2293cb65079291b350ca339d6
z9acc5e42040a9263a26586651e393d28a103a273e0c8241c43f45e89981be6d3b9902e3c733926
z8e0f4f1368c7f7d06ee87b4cc7e097d1ab284751bb4590ef044f2f32d29ec5c2fedb7792b04457
zf2a2a7bce2d924d835ef3f60768737d3076ad9122573df4e218e8b1d32feab6c4c9af571fd41a9
z2002db286c12855027a4e0292abf95af97d4f08a8da5441c838abfcdae94ade62d53b3c47539dc
z73332259a8f253af2e97986cb672e09ecec1f32c554e36d7719edb9dc8c208abacaa8f5aa0366f
z24d13d763f9f54541bbebb2f5b6542ff830ee40d4065fe9d946638db287b818682207d9680a09a
z31f4f4119123ae3ac7415e4ef15e42ad6febed2acad09726be33cec7c76fb19e4dda48fdb41cab
zf3b450a6595458d80ed927517e18b99ba6f9a028cfbfa2cddbba3ba567822d65efa1ccf0befd5c
zac9a9d2c73617531dd118d1bce188283590b1c57d2ce11647e53f64071fce21776367c638b24c9
z4d91496633d90f351e2c6f2e7837ab06b731f9e62676ca19e17d1124ee94945ef3b23c30f45012
zf584a24cf74b7cdb25611c8e5cf4f8101796104a017ee796978e2a11ea1aac83fd43a8fa7558dc
z61c83071b281571502e6a83f77ccfefe96ab175645eebe61789e9e916224c1e8631e4253c10c82
zc9a1fb341326bdbe3c950c2e7231dab16a14ce806f7f75935d32cc4521083dcf09cd21dddf3f77
z2b63b467aeabc8616a65b18146313d675e4bd071dabaa25f9fdb66105d4d728ee07ee7b4b5b09f
z649113878ec0001b009000c54c3a17eb955db02f68b3577c4ce1ae113012a64997ca07e139a5eb
z667f6296d7d4e8208fef52a7433db72d2b30b33c379478f480c9e6bdae6af56fe1b7eb3161eee1
zbd4766487b39bc6d9b9a949ce56ee453c49881fa3244caca68d27aef5d2eea2e4fca14376ddc29
z32e04548be87aea086aabf43614804df09b67ea374e05f7c485666148911d129a694a0ace4eb46
z11885f6ad8f2812eee7b2da842f52d12e40b7ddefdf095c3c99700f43eaa1415892bec617d3548
za372e666e3c902b469db3124499c53af6023f4e800bb846f9eb96d3471d99c1ad62a5ef1fda546
zb5022825ca64e4b4abf8853dc67b094d74f6dc088d0f0d740591ce50f23ce157257c995ef69fd8
zeeb466ceb381fd2649b7e5d985e5a9ff44c9ff80eb0e223ee46c033290bf6275694d6895a880fa
z12e91f99af60599fd1299336361ebed7ea7c5befbedd12440a7c70c81bc71201a10fe53e1d325b
z8d387dedc2764be4551285663b0aabcdbe8920192024a375bc5e032a2686b83c6b2a59c12e856e
z72b5b18d60a959c8d81b2130f3d9c6db25472aaf9b7400401c260408a5e4fb3540a4b3498bf258
z77b6c9215818bf26e722b1eeeb9032c36cdd2077ab9cc32a266946b53cf143ae771f34673fe5dd
z9338226bb514cadef959a6cb05cf531244f496d6b0c9bc6d2266588b14cb49bf7bc2efcbfaa48a
zebcdd62d143599d2c03e414d119e6833f98dd743848045d471a6c6bd0e0d0f6f5b78e675646681
z36f82e32e2916e60aea9cc0986150a3214d0577d27441fa64bdf283d09e34b480e99b9d89a62e7
z3565215ff74851e6629ed9a88807eb6e7f7472479cb6da566d9d1e1ca4625a5322dce18f407a08
zff746db522c51f6338bc9181178fdaafa273a306c06d21a25f7eaddf65832033d441401ee0e2c5
zb64fff0500544a1a502ce622c5fca98d55750f18641e226dfbc06f2a5ebd539caee4c6e6e4789d
zc51f12a62e43ee3002268f52a696b5a3e8889073b51cceae63a495e50896ccb4decffce65162b8
zeb9515cd676a0ebd693cb2ae27d004a64c1f23b7dac27bd4b00ecb5d4c70666b34b6f68b1398e4
zded2d4d1b84af18e342a1ca2d26245e4b08b1aee8b1bf1697df959324ba9d0d174f057fa83b03b
z82340bf20675193e82966d726777bf2ad20260d7d6d2c0c6d80d97db29c623c04f5924886a1694
zdf7f48dd1ef78b91c33c13e53dde158354a8e826537ee237ab71eabac649c8401c9999f1b67b40
z34689e0900374177b45b2df5732bb0fac79898a434cca7361114a78a2baa5e885101b854f62c99
zfc68ed228f587efc4b11fc28b3508bed5d30e3f554d51460c9d5322f23807a18226e152026b6b9
zbc9e7e6751d9773c85d40b6deded431c090f99e7a7eca428424834997a39465c1c8fa2c61cae01
zd516fcef365e5dd8b348a86451afc9fc6d0ad611d93b18f466ae3331c1b2baac8e063beead0384
z911a31751d158027887c845f8668c900e0629b1637671103c4ccce1eb9d20353d91cf57f1fdc8b
z682d6487090d08f50c2462d1ddfb157d157fb75d3b4070864d5514af2906ddf49996cb7ba9f04d
zd59fd515d3e4d31230bbd9bba82fa262433c70c7fc0bee0945d9820a88e6a0c62a2c98e1ec377b
zad97267dc75dfb9e9630994eb3fb46eff4a17be071912d12dd8ca457ef58c55bd301e4ed775ba3
z398cc72bf35888ea270e9fd96a9ce9ee6f21a731b708dd401eda4ee27d3db9de64b8699874d942
z2b89010c63b719a696b464edc0d6e9265829f6f0a2658b3c7e447aa58bd06560024fb942e07c42
z576c2f3133b58cd009ecec0f3e26439e4fec15dafc6a61cc6fa3f738d6d8c3009d97636df90abc
z79e0519f249ac27269496a7ab728ade3ad9929e87de7500a523ce2328d6c5c02ace6da701f8b37
zb5dd41d7e9dcc0bc1b65c03fe49b5cb0b2ef0f7e412c96230ac2d685923405863e653951f99a9e
zc73c683e848f364a20cecf751c641a637ca3434e6ba05e9dd5a1ec7eb03e8e0bb805b39495438e
z40f3052d0796fce43fba5f81f0206ee4989a72939c1ee642bb0c102de8bb0a7e57d7037f0f5bbc
zba36439baceb028748167facc27a6fe27220a1d3825cd56cb2e02299a32414514cec2244ce4648
zd74ce009b75a710fd2f6406ebc2a7533428e6232ce9d5dc79bf37be03e04ba2f780a256b9813a6
z1a2253577854611432ed28bd5ec71275fbb21cb69b002f9788ab47ae162ba6026c782a72311c72
zce1fad492e355fb6d6b4b95a552aaf5789efa21c8e775ddd7586a97402cdcc0acbd17b1fd0d9c7
ze175bff0ff658d084a4425361b20213bd3be8d401e8cb8ea6445e12ae032aa16b7bbf89b142983
z674e6911d77e8d79173d8363dd25fbf2fed847e7ebeec352eeeac830175881f17129dcf5464c3d
z727635d0f4c0906631cf8fa38f92ed2fd1db7563a425ebca878614a95b3e13e7a71fd96bf3e691
z12d64a7c79c3679dc4bb4b1f2bb9e328add775c573acb572e1ba746ebb04a8e0d8585e8327000f
z0b51830600c7c7451e2ffe8faeff510826751eeb7a214db9f0883a6f17bca988d2e774c2f0c7ff
zd825429fe043a4b7a0f8d2cc3e00363f85e50961f33394c2045e8fecb3885c3ce771d81ecaa7cc
ze4beda5df66b0cede0e22552623938f78cb384f7dc5a7a3d812823c775a1c2e5a045c29bdb7205
zdaad2ca848845f19249e11062f21bb7efdac0957ce97b39f9562fb7d9037a1e7a783cd36b21d7b
ze6f29f9bc2b439adf2e66246a908214d7544cd538a08a8f1a2a23da39d80f895388ddf97f1ac42
z012121bb7e8705c82ab891be77baafee541d20ae0dc0fa6872b57f2192fce07ea38f5ba5eb2d7d
za39ffdc5087768ec7a06626694b75b834f9d9ee82b0f76fd64dee62695307e389dffa7bf0dbeb4
z7d4b93a7f99cfbe2ed08fec236ec95636d5d2820c175b57bd993675c3d99ddf78c26090563c39a
z497fd6fa55223356bec9cf520c870682d34a6801686d0781d51645a93b227a1d08cb71c221d25a
zb7351b801b2a9f5e65aa623b87981f9eac070b0a3897d10f739d97d208290df799b0e492e2a72e
z779983808ffcff782f4e36ff7305c4f50e4c637c05b256907acbaf2d8bc0c999079aa66676fbc4
z672f1efbcaf6db0231780b33d254b222e2f1aa6dda5d4f53dc7e85dbce038cd9c3bc52eb12583a
z429c8798e9866151a3694688f5df7abd43bb0c584020c35ca210500f3fbd9648b296c3c7b85eca
z544fbcdf41f11cb79852602d6eadc051b609c0fcb507429d456d8c9cdf97b9f01ed6cfb823ac27
z117df650df1156bd29c60959deb02f6043db24d114d1be4aeaa391cb29a3872d9051ca98a703af
z477b049b55a3c0c54ce26b70142f6ea8a7407547b771bc1a842a2a9647eaf11fdde9e888363eca
z354876f0930d2d2678cdddf2a78dc52b004034af4b3891d71b9486a85be16d86b70291f3c47669
z5dd60f430a16fac90a5a42e4edba6c2587781c3fa86d956342ecdc488229443f9374a4d9f7fd0d
za195ead07446460bf68b49223dfbef47ce825ca9a792e3aa2881ec2cd32ca68630aef8464caa60
z36a918a08dd18f6514384176e1161e5b2dd494301d6ecea185f1583a3b6f80a0252f83cb64c464
zcc839819e4e73133ba7e628add0a6831c8a34155a4583241c34487f5e763ac5694b69d7fb4d2db
z84a71357f7befb7b6c7705cc84b20547609c4cc9141a4db5504ada3c74f445427437c8984e3ca5
zfbf08dfbb1185f98eeb050a358fe6470026da9669ad201540feea89164cda1479a63ebd1106458
z002bc7eff0f239f18d0c850d976288f8a89268acb7eee82dbc185228b39f2509bbe805014272c5
zc6d7a6c692ff37151a1906ccb45ebc7f529857fef411ef8962a1383785a7d201dc8543eb65b6a4
z12038cbebbd4eee0d39fce6ce47d06b8efb0fa2244a965fa54e7e061dd27c57b0253bc7e3aba2d
z41fbd84fa4000ee8ce440f7c0d63943b5df8a0859af734dc29749dd81e14072144c1be5f4db633
z35e51c658e8b289d7366871e650f87f7d0deabbacace6759fe1d2152bb3dcbc07ebd4f412dcb95
z6f5d5b9d675460754020b684590e0a32b63967e5fa77abe3ffbf8e1b91dd76d7fd76e9e7554e1e
z5016a2843cb6ab7bc3e9a4bf08f07a7460d24be1adcb1be041b9fcb2b8af084e731e70b3e47d94
zd3e0ccc3c4f640870e08c460a22a7fefeb8dd45f1b8a9a4a2fbd50c4ee257ca4a970c77ff9f4c0
ze934baeeb8749c92f5b943ab90bcfd2322dc0479d2a1cba2a4b6eb2ccfc95a972ed15488301f10
zc7d493f710d3ef54e0d3db937fc2b96b9ea550b90c9b978887a1067475e1c4fc0cdf8ce169ad53
z686056e684777596f6e2b0d804cb19bb390b57505aff041cb4542a96e066e07e1df82698a6e21b
z0baab029c28eb5e5e8b8b3c3620e8219f04f409fe67da4b96d42598798c4d49d1cad08a981976a
zdbb588186a9320a323c685cbb37fc85646c2dae8f2525f5c03118ede217b37d3a932f1fa1197dc
z5af0d8c405abe2eb36502fa332bcde136f2f80cd430d13a83f91e19b10c5327dc9468c4998f760
zbf657a2877448d065d4e94f8e579b953c2507df4d629c844f13879961ab62c06da63917ecdb19a
z80a269c956cdb44ed797a3a3d7784731ea7e863ece49d164ec9c1d519c18be0868b68947b88ea9
zf4281d43fb8556dc90872404bace53796ca945e1b77209f7f19b1c3eb1a6699cf1be2bb40409f7
z2c86c574761f8bc141802ca0f8ff914fb31ebc384bcd43d860c762f7b94ceb305bdd4642d0f585
z581359dcece4a166988d534d9de90f7569384808c1d9ae6439951b312925e38486263cc012dce0
zead21b474e957bf38d21169a8eb7653b315e87e6bf025d0bc8b31216b2d729ccf85a94719a9ec2
z015d2940d9c6f9b0e5480dcb537bf1c39706fdd9eff40642b7a909b1ead7fcb3dbc2a20b6fa36f
z8166a7ffb4a9bc093e52f6a4eec2bd2701ad06d4dffcacfef73c2d4d528c5c431d7b66e0a0bbe6
zb3e157a4a9aa7ed146deec722c3f763ff36d8eb0ff10b1c4212d3ce44ecffe604800ed396e2060
zf0ebbc4281818694ef5e0d5d5ad7989b12ad120f7fdc6588c5ae2dcead7c6f053434beb2b734fc
zc02da300718bef0d7de4e42eb360a148605d67ac2b54279fca131374b664e5f701c43138d18b49
z410b3fc4a14a2538a0c05cd66e1ac843892656b2d1b4fdac41d23374f8ae0cd636165b43fdb0d2
z9fc41fb3d916346ae967e3f3380b188bad033e2d9b1246f25ce99db8361041057ce219dcb6f050
z879e72f2097f03a03013f5ae79b1fa7249f66789acff100fe101cd95305f8aca0cc90edefdbf64
z603386b0e31581b868ec4878a69df09d1cf317de13868c5b74c64fd551fd1c6014f78f7f5d8f8c
za6ae41632fd90545110e038171cd29073051760e6d2fbeee8d746102d6a7842c0bf830ba75599f
zd08024e142767fd9a705a25a46cd13ba79fe50078255a1be65c85c6fcf76a463eb1e959e86e14e
z78bcdd2607fa005173e5aad153eba9c611a199ee0493d930ef2d439b9287264802b3eff09bc8b5
z37f4630bd33c793842c49763bc640f701de1f1de0dd60064f0793d132ce00084bc7dab196a2e59
z4b96cb15b04dfb4a90b3376566e4ab7b2cca93313fe1e605e5191e3359d693b0beb2604aede7a4
z45b67e0ea388aa6e048d2b3d1cb63f8b378f6e02e8fe2dc96ee36882a7c1b5d693ed4ebf651a9e
z45ef934a4f72f436ab1934a492f2f9911a1557594e7b615826ddbb8a5aa33e5a035ffeaa3cc46f
zcddd4a09bd46c9ecf518a943c828a043d07f2b2e9c19f35a4a90c4a25b2b999cf07c52e229e87b
z311ddacad23adeaa954a015cf7e4707168ed1e3b5279829deeb07388ca4142a0380d5ee5dc49d2
z4582908185e86537ad98be3a090efe92a1f08c77f764b644ef3a6073ef66c4a6b4aafb6af8af0a
z95269ff8bc891eaa878b5697e87706026a7ab06e1f23babd55711c5799fa21b173d9e25ac01e73
z3a5fd466449581dedc98c6e4b5c7e1313411ed2058d2a49715fe588a29fc220fc91dff36f2968e
ze8b3147510478b961081ee7d2eaa265afb57a18828fde0e52dbfc46acfcf409069c9a40725a7aa
z1542274086824475fc43ae6f889f6759f070fe34d8d3c4e30b637c3e0556385b2db5fa6968d8c0
z7ae736aa7475c55377e1bb488dd793e06a24634a1fdaf82feae2327bbaf5f4c9da6d75384f8071
zff78ac8f39ecc2950d612ca9538e72cf35badfe6d4b6d092a768beb510ad68808af5b6c73a1744
z67ec0a06c7a713f894f9431e277861561d3a816eed22c4225251d739e9fef4a2be9db116e2c599
z4be2b289f40267a48488ea116f4e4b954618ee2e18a31c5a7929884ceb453aff972289d4d4803c
zddd28999381e606fe634a04ab48dadf34f18132723981f4704990abc9fb599edec9bf169c2cdac
z2d5d600afdce8ac85baf5a4d8fa1f89eda8c34db125462dc43c74556269def5fcdf4b305d42d9e
z110ad69ee54968f14f8577f3b72f5a31ac805fbb65d8f32f41c514e89733b5fa1d7f2864ad0228
z14e6dbc5534dbdd4f0ec554a5995dbda42ed94719e2f7b7c1925c96eb9d9a1066b902469ad3270
zcfd3f82ee81b7c26113547cc01cdc47834d0cd61c27ae5c8a59fd6026237eef813929b22bfdc61
z05be7909e43cf02d5a1e8b66ca881cb8bfc3a5cde3a27618e1e554f083548197e32178d6252981
zcd8d7a8d0307dc5bb770253734c131b84eedb3c329d65a0d3c1920ffc9f34ca65d091c7411c3f0
z4a851b93a03cde1e361908c581ce38f65785fb0ae8717505e0ff84b09da404f295f55ae14af31b
z5f1ee639c4dec35370c09b37ba17ed4580f68a5d27432ab44f2bf37293208bd251a166fb9ee70c
z76d091a64967dc7f280a82c2dbfab38d7800d471a5c10e74727ab6649e101ad54c9266ec025fab
z567752661b209e3af9140a44cc2652cae38654c687ca05df9ab277573d5d1a65e69e97fb15d8b9
z4b97a80ad65a269f01b389e41798ddbdd6be6452b2961a6d72393684a6cae22eb9551d2dbf6129
z7974add7765e34b5c4f0dbbf0545f770dac7b165baa5558e217da081c1c385fa614f7dda484278
z0911fd60239790d21ff29774c88c92b7be039a1488e25ed591a43495f11b9de5d05e557154d106
za54ed1fadbe0876e9d268b0fa2015d8e6c40d7d33c2d6b7a441aef303089e4975e73618c1f2884
zd61c2c06709982ecf2de7723e6d32a8052e4ce940fedf167255fad3e4982f690bc8a4db480f3ba
ze8e037f585bc06d9b1d50e59064b09aa4eb6c1f16183d5ed4f70626ef9593f2a532df5d7b56604
zb5ba7da80fe1d1175fb5f8af5142bc42147bdf02db05901c7077cab0ff33653c8c397dfb473c4a
z28ca3e9b230a286cb98bd1b6663ab03ede2bdd65015638f481466cbdd3c1f52bda1f221d77309a
z58ede09fa6609cce8e810a90239923886e285e6c0c1e8920832613395aa7ae705244659643a660
ze2efe6d99ec002536c55d48d8ebe615dca2160c58cd29afc1942681675a3f53d13e3d8ea2e4f5a
zd33ab8050045b4b099f63cb159848b876033dff9624386827f5a08662d6c9b27d83fc1f7b2d6fd
zdaea5a381b60268d070a3c2207b8f39b5246ba9211cad4cfb38400afba381cec3aa3fc5f4e7552
z10eba9c93d40a32fb1f81283341440413385ee573fc73bd6ca3bebb6cf77f563c3d998c8261b37
z1467041e16b75346cbee56c127447ea9520767c81ed15f747108cdc37aabcf876152cdc2399284
z5d28146d0a46d2359ed77f59eac6c4afb7d3f8bc817fbd504b82f1b38a221afe2191b83fcaa070
zf105698165e7217505a5ff68f9020cfbdb2bfc11276765530292fb7cdd37b179b4ffc619308fd7
z6614bd0842c5cbf0bc9207038e70ca8339a084b83b01761734f822412214ca788e02a03bee60f5
z08c7ff59afa9fab0faa14f8e3a5d1003e9325d6f4e538d6bd1ce04e77b4b4426b53b217c716ccf
za9b7743c05bb239984391ca6aca2d1f32fd8d06387dc9ede0acd18e7f9b973c08a09e860a42331
z887d060941460c4d50e7515d7bd31ff0ea8bd1519f1188bf57ad43e654ebda6e0672e5793df68e
z89ef502be439c1ed2eee8832c7f36e7b663dda791b48c8c0d81e3ee026917de062a510ad82e04a
z3d35975fb5da52426f9bd1b1cdda3e64c3918ca55556d9edde32abe818659375cc87053d9d9bcc
z0f41e9543c7f2abb8d62865729ccba7310aa29a8fd11b942aa219b3872366bc7865fe1d9653504
zaa666758a5d1939ce718b6ecebdd9556590e35b9f8b45347ebc03d446c1901120d76cdcd34e914
z2014ca656d2076f2d64c51a70d39806394fc1aa90dd6cf0646f2c5ad7e9242be20c0a89867086b
zfca81e29fb87ac2bb436a44ff8fd9256fab1d074236f7d9de3bcdf272a7609e627c1cb8dcd220e
z0416c56417b4e1dec30d339e7a694a3f11f1c883d19674e6a2e2f1ac63b087cafb4b376d1ac5a1
zd2862ab65488005be6cf7da0e93a791fce874610053e89c413bcd937d20839f3de87aad91dd8f2
zc213b7edc01ea0d8e55e3f8463b37cce053bf25bca733f70aa6870053e10851a34e21979281311
zcc623f8835aa3592d24e0f4d5b27852573d6762dbb21bb3bbc71760bbca6602fd3450da136a304
z236dc879043e3ad10a11054294ca9579f99a20b24fddd86fcd72caa380bcf4502214da5188b275
z8c2b1f4e4902906162607800a55ecdafbcb7d8feb75eef903208c22b3ec0fd0c47dd90efbf9404
za17a139db9384636bd894e04028d649325d4a0d59e63602a4198bf52affdf0b7cf18bdc68a6b24
zdfd0ad25a08d251fd0c28b131cdc017e19619a20f626eefb96849249f7de0c97cd4a9b54df41a6
ze705e0340bcd8956a71fb85b17764a2d263cc7153d38d938512039edfc221f22fb0faecdd8f23a
z3f7b5a2979e1d30739c57bc0390f3ce56cc6bc1b6548bef560f2c5a28abe6c7cde23635319a622
z8ba47286820c6a47951b1a161b99f2dd501358e6d657936ed75e3dd688b72c7f7350b57d3be425
zf8824ab22a9d98877c403341d65d015a8280e595148cc26084193c5c02269415d250fff2a8654f
z3db5fee290de64c66e1844045d505a2dc3151db46483be779fda66682f93c5190511c6bd1902ce
z473ea807466f4dc47e01ba6a58eba3443eb8158f2307eb4704f8eb124cc9dd325765b6d0dd346d
zb552019a6fa284e83738b3d60357a6584145eceb4d7dc1c0583b832c7ac2a502dd60065428be84
z4936076fd7b18c3a87c838376957f863bf5da9021ba58ced34fcf180c6ff5a1edc78d1b9c1aea3
z3ff728fe21f25f6f800b8d1b6e0f6e4b19426de4cbcb498f9628bc69fd5eed269b99655c222707
zdc42a923b606b04951fe2dd8bdd8f6e8d9223cebb2b6ea701869ac57299ff1c003d7b62d032dae
zdd22e3092c1ac64a977024830f44c0728481805624b63b001de691b8afa2e5cd39f539384a2b72
zf07da50534fd6aad379876e43e6ee8e33d4d798c221a1fcde638c85bb338b29e1737624ae174f3
zf3294d03b31113b4e4246dbc807ac54fec91f13246892e2244b6f0aae3f109d99678ca53bdd452
ze16c9eac8924a242da8bc81b9a389ea20d434a78e2082f6320fcf5503021002875f202e0e0a873
z9d80b60a9fe885001e446462257a01680b6cdb78ef4e473e4a5540d79519d721dce81fba6d27a5
z1e0cc9094c06d33b497dc64cf186edbd9816e78f1c8535d358800cfe627f1850c193fee8a087f9
za1a429f4b94b4ab79b62e8ac0e3bf118347c3e597a4b9618b5b930e170c75e6ed40684629a4c1b
z464c8828ce62c02abe5b132025ace5c583e0f6fa3d3196a646c6fe882ca88007712fcb3e094342
z98f4092a2751bdf18fd3a6dfb0d79a1cfbcecc1627cf0242a0506c29523977ff9c4d5085482cc4
zad3ff86699f64a992844e56d0c3aaf033579ddb0ead4ca17d50a3e41829c7a36d800c23874ccc5
z4fde5fac6210f31054b8bebc72bf54612a948aacd8189d9137c426a617832d563f7dba5fdd29f2
z6df768d142109712d31699048ed62a7f86fe443614f6f960d881c9f30528b6a28a2e3edd6cabde
zc57613dc34c45a8be19e674bdc507d59272b9cc9d302ee0f5cfb375ac508a2cf2cc8bf5b06107d
z72abb14f3a1daf696e0dd5510c001b4ac94e346d1679bd0a8c26d05800b42e32102162f6f3047b
z9346f9a450020388cee4aa9fda795cc8e0e11c98d746c89336f763b8478eea3539c56fd7462d0a
zaed6c4e7911fe0e1f194dfdac8506492391eeabdcf494f77cde95fc31b1a4140058ae58c68ab2a
z94a57bd637c7469a3a75a53c82acfa77174ff3ae68429459f490f532f6980a1e45c34a107fc8b5
za093b107a0fec64a258cbb8ab60da229ea2efc92e60e88f88a3291cff7d35da4ec2a48ad15c65f
z24788bf80dccc2564221b95e1a03b8c063b25874957e4a2add6c5504f7035a997e9164388de121
zbc2874f7a7cdbedd4df478d9bde766462aedfd68f4056fab336b415fa95dd8acfa6eb4f8c3b17e
z62025d0fec038762d93f8106887356172b17835cf3253ac53379aadf9c0299dbaeeef975dafb53
z7c8866f9629a48c92f9953b95d640e6592143de898b651719703822e88eca8ccaf8665cb706329
z31454bb2a35bd015b30b1879a2ea0e4e9aea0b0b36873829d87266fcde5cc74f944a31ddd9824f
z7f779eb06963e9c108c745ebb8388ea7b5e7b147c0c2191430b072a2eba846dc6be8a0ab1c4e3d
z0f66c8122fdcfae94d617318211768a91a83ee0cf141d24db0a1344dd183f210e5932b6df8c278
z3a4e82e163473802408efb18bf290746a99f69a7a0e0ce029b38ca1082b92deab9a51cd47008ee
z3fd913e1e5f279fbc3ff4921ba03cc7b578f225da00a1695e7cd32a1b50d41fc7c6c78c8700ef0
z461e4855f53dec7207c41a37d5a86bf83bce81c8fb41db7a26d17de3180c3eb742a13d5fb6e659
z7c706f5391873ff14b7c328c2afc136ede16cd69dcae1ae8298e093e8f36c31714a17e4385ee45
z944562f62885bf40c06939a974b0031906ad60b41ac3ce7346fdaae1e3c57b72e4ebac024be1f0
zf4aaef4e68228da958cb198399adef0de659dbedd7d026e1174363746637203fdd4ff493adb1d0
ze64d7707fe9db548597ed6d7e6f3c207fa394f08d1db9853caad787ab8a3abb961e192974a35a7
z0855cc2587b379cd266c092ee15a168acc676cdae9ad8969b54821f36e990fc053b2aa5ae8e67e
z48fe02290e80773c2457c364c8d82b55056f38131bdbef12e91fa0e18c8cb0c88ebe6c9199f718
z878900a0cc5f2c67d56abf137b997d60a2841a73a5eae2d340c704224f95a9aa1f3aaba265a332
z65dad017d3b0c43c3a09db31ab77125210dc63d2820a9b095b21104381b17ce3555c074573daa3
z5a771594f274b465debf50c0f02875facb9f9456634e2b64375029c0e25411c6f33ab16a36292b
z0ce44236bf2b6bc9b998b6fca88968067ee0e77756dbdf0da00a75457b6026493d4999a4c15b3a
zc429f8ad9aeefcf99d68c090e1efff220a51ca6b317d935a518f4f36f3929a7904b40aa46d67ed
zdfe20e68f55544dd1cc6ece822d30e8570616f212592ff0ef279dc72410cb4d54804a482ba9807
z1543338794c204066008fd260b7237426e481ae277f6c2d8472dcfbe961a7fd5ebf7217a13332a
z4a52c396b0df6ad4142eba5252e188f0c3938cf9866884d8c2ad45332b0e7a3bcf7145f8d0d8ed
zc9339083aacf7beca05fef156519000c031dd8eb9c43e67779e18ba192c949f5d2d15fef9f1d3f
z14b21a205e45078893fffd3d26b29ca05376e503a2ea1dff4df8affc84d56910387b5cd9fd53ae
zfb7294f7965c29dba0724368a380a8e0dd4328ab877790c1bdea626d0facaedb178e58910f0f32
ze30859d54b7ee5bc3e60dd73635e3d808d71953f2c49da42f328e1c3fc419efca2d288b7010a80
z5d8f031b814fb3669111a9f0f3c92bffec88353ddac3e0f64f82e119e8c1381314b256658cc18b
z9945a6fc51044024c1e8bfcd86c695f6dfa0096a9ab177e7681f8fc1db7fc861110ff0fa01eb43
z09511419fa7c4a8d79a007ea18d982c85079149a632b05c526138055a2956e7ba34335bcad5ec1
z1215d9dcad493d97ea8d3084f5ac49aa7bdf44b4800d257bd2f26a05ae4db86bbe33a0cddc0eb8
z0a149dc2fde5a7c9f1e3a2e393193c28994441fe3920f2b5475e9ace30b6e4f2393b3b256c025f
z1314b569e8bdac8c27098e086d7647b8c30ac807ab7516a008dfa919f15a05f190206f4d69015e
zbb44b595be08aaabfb2477e8f10d6acba1fb2597a3ce224aa959efbcfe47a12abdf21ad9ae5ea3
zf9058ba58d8aa1d236cf3ee8af7fb608326348249602305dd1c96e68f7e96e28eaeda3f0b92215
z7c20f78931ad9df7a9e55443e279a16437599f0d076c5d06326d1b097565816a1202d53e97291d
zf3e14b414beef0fdd191e71b9d9fda1ceff0bbfed5b7829367c2dd4922b30826d05352b14766ad
z0151c2846d84bc5cbb668cf96ef8fb31647b5329782ba2d89aaca7d858c12b035bc07aab2cf1f8
za7c30f067551639961c0e2dd0ea117dfbe42fd16ebb46b625a2ff076005db42417ac4cbf2be0e0
z6e1da5bd4e117c6315cf503857e3c52aa7d2efcca5b8bdac7346e56efa6b94e2f72334fceb71e8
zd41eaa0a3bbb0c79a18938fa2d7cf862b98de5a081a99ae9f343cc8a44a4ed56ed0e263148c0b6
z2dc80241b456f60db5a7b5e203b94a632d12cdd254070b1f5e80e4f32122ba535c5c30eb016948
zaf2be730aef3dbb6f1c1c8b795e90f1b839e467d0cbd3848be2be8be3c9d9019eb4f0fd10f2f5d
zd9f4810a236fb77c45d6be0fc851f4ba7bd57bcc5b43b448aa476cdcf82c3d7c48e42aec31f7c0
z1424f58690f63124c1e8fb7a7f90260a963153d89282cd6056041f4bb8b42ce79e6f1497dfed72
za6c29cd7da99a86da47eb7a36c21de1cef95b88e913afae948254ea7318ad73960c06244fa10be
z2430a1bacf5412ddd63d5f7e81f042bb5b20c80f31e1d6a1a4da1063a55835acd16c422a5cc986
z8bffec388fe1167e0a2100e4a6b53a22ed15e6898aa44890d322db14678b00c0bae06c8a3a4e80
z86e75549422fee6dcc780016614dcf13b87d9bf291f50fd7a2c12364fae1e840185e328ed3a452
zd311f52310763fe24d5b57788130ba35e020677678cbdc1e51f6cfd2d93fd29f2f0b3a0bb43490
z4921bc9cd866ab7f0096ccf716305f8cb0241ef76fbe01ef0cb8316567d0941fe9e0df923ba02f
z3f9524d15ab2e4598057e7912fddb2dafc8caf3f8805e407ff9c89fb62146210cb82301ab5415f
z7c7dead1f4334978d8a8642aa5d517bbafd7669bcdbedda7829aab101ae0c97ed060a30dbbfe8a
z6c79dd2cfd465fdaa77ad7637877f6e98e9df1d05c77f2d5b9711107ca5b5d34bb8d9f2b74fd26
z44e78b7da655004b84c2b5d7c9c1dc3e7f4c762cceb09ef3b906f6437d25eebbbf6e5faf4640ba
z4b2ee6ddd1b3c2ef44d92d61b6ad8fab6d88d917880f530c48aa664b40d3eab241b252cf243806
z436ee74c544c899b6060d6f263160fb28039dc6b0015cea6fed5a24c4649f40680fde72f91d339
z354443b5f06805f7eb63081137ad49780742c26bf7cfb967d2ef530d97068d9fea269641219d00
z0e20ef3d1b06b4ebf571248f64c78b72179126f557806ae1e2a6c2b31b1a73994e9516c5e549ee
zf0b62e8563baeadcd33df3624b799473e4e55c630f929b40a963fd2b62a5d73d4b9ea031598093
z3fafe125aa814c41ca1f539b3309dc70e1564e0faf89a8ff0ee8e56851a77c7afed863de3294d3
z9786982665172b0ac7e19b82e1ea6241cd143ae6f1f652dca9e27ddc98d7dfd0b0ff55faf0e018
zae84797ae9ad70d90bd687a238d79759b5f7ef101790fb5cb8c0501e436ee868e8676a9f8fdf4f
z4f9c1b957e8327fb44506fb37a82f42da321bde14de03a273271fae5d421d3a96b262bdcaa66d9
z3a02de76ff1147dc8365736b36487949da1ef3dbc5011cd910337d4a2eb535bfc17e70dc719b0a
z1e48ab5cae12676af3f2f9d37888fb14624f518761805757b72d5a84a3a0ba58b934c8da0783b2
z7dfec6e9111bdcaaf5bcf6a18baae5e66185767ac71179a2752bf19f109b5badbe924adbe98c48
z7b01761f84d92af7c12805d800680607c47342752d7ade499e2a2d31adf6f47133c4b649e5e2d2
zeb7c3c197162c6ef4bf1ae27d7d638229daa0066c6648b215f12860665c3421299cd1aace2b658
z408b71d24023a5d4a65e5e22fa4247b2ec8a70d67287014d6c178e9be514d990475db56e70c5be
zea0197e3457e0dcac830de9a6536a796dc6615faf598dcc864d95640ce4a7817a8ed436ec5b34f
za472b5ec94bf9d73cecf52a058cf935513bf168602f9610c72611d3787646cb53c21cc2fffcfa7
z1a561ab1af61cea1b031c5d10fa3ac01241b679306ed6e6e212512fee20db5d1a4e9d031a98d37
z3cc5402c970d3434db6a15c69ec12114f76e9e1d962706851586b0ad1808a4b4673705a262d76c
zaacdfcc8ff92589ee5cf94c4de00215a6502d0f03e892d5e0d5929707cfe8469650a625cf14c9b
z2d4d71b20074c6b8a6f5a08bedf53c9aa10d3bf05972090b72c10fc7b486f91bf8c4cf05f49298
za1dd45eb156fa8b2d29e6b8c7989636ef88727b27999d97e4ca00c54e2a6c4698efe32b5797d71
z87f367586cc93eae34e31d4d3f587ac86481a10b71fd7a5f1d086c306f9882efc9f8e0268c9e08
ze460a9d65829e041ae9179617636abea2e9ff0a2419525a2d24e2ff328e459eee6c29a850a3445
ze5c2b609d950a5ee8c29853964e9dd723e10d4646e44bf4411aebf560d8563df1647448faf1de0
z7fd074a9f34cd0b082ebb382143e96e51db4921dadf2804809f110f0e96bd6da6eb2a81c857651
z84e7b07b9870cee871c2dd483c128375b096cfe2b69019cf03258d28500b7bc10760ffce734156
ze4939a2beaa03cd794b51dac45ae7861cf9ff24bdb49981e23d4807c17fd0ae8ca75ed8160c7f7
zdc9e1f6c55b0942abf5b1f2ca8023be718a71a30ca28f0a220d41b304aae42ec6b12672dcb4e42
za0ad558c3f908b290e4f7c367a077a5568c01366c98a3ade19d5dd51a683b48fe2a64b2ed87008
z2b86096a1f499286a86f7065759c563dc08c6e28b01006738c251edf26957493ff40ee32558029
z8fbc96268ad20f99eba517092ae9dd380d3c3d071415ef3f3783040a99c91efe7294f32d0ba770
z932770683da93633982d7469f69ddc0ebe3852827753dfc9c8cb2df922b451b9ee02acb6f22682
z38cf995318988e15d86dbfb2c6edb82d7ec765e128fa800300e86aec0243f0c3490ae637d67779
z53325d8ad50788dc2b196ef095cdc9922f922106dc82fb11475a8ccfe8bc8e2c2fb5d67114b73f
z184df37c22e15be18fb12e4fca95b24b908bdb3d74523e0d74b7c33b30e13a93e8bf96f2205977
zfc26306a4cb7a76e0d2f6372b5641f137bd3093fa30bb6b1251573eb5528a55fb8e8fdc139d012
z5539d1991cdb0424e81c573a350daed5f585bc1690a1334f2373cb56a9ffb7708f9180d2841dc9
z120efd0615cdbe11d3f080d4b93b1e284030209370d7abefcfbed4958a3be7b27d6a480ac36391
z3e01bb47a6f6b50587acf22ab398543e4c5421a97e2eafa1913b0df1bd5d9465f31f9f4a57f0b3
zc4addf775b7587661f72ec0421bb54e4040d2175ce54b154775e9fde64b3098deef25aed4319d3
z4ab7c945eefffd9593e0dde7d87832c6883d7946cceebbe0a076a8fce22232158e2dc65b05397f
z835b7f173b03b9e6fbcc5ec99a033899e24571ce2f27baf35cf8befa34bdfb1f28ccff27b552c1
zeaaacb3792d0f11db1458eb658cdf901a5424430c5a9004693ec17b486ac121b84662a9d02c9bb
zf6f7bff45fbec13805b61e7d1020ea49025617f08ebc189cee23e8657c9d2d8cfbafeef4a5c8fa
z75cd7a8e70af9a00b4e9c23f27769b708d27db09a4f24dee755c6a72c211b4a3aa5f40732522cf
z01114dd43a520afd0647421644407c3e7e822b06dbbdd9cbb397a99f4105d47554df5a67558351
zf025198a4b50967e9443125392a0458f4d9f7907c7e4419689dcf0154bd1e89b67ae6fbbee074c
zb9fbcff77873d2d3221fd6b175a72f23f7ba1ba3969a0ea57742121e17e8f69cfcf60c2774aa56
z9cb47de734384f350ebd4e2471b08295f6da6177efdff1f0c8ff2f0fba4be994f56be7b4884e23
zb16f60d170370ee89ba3a882e0894961dfd6a70291fa1924e061f1d5a7bcc7e43d1f37b83eaf3b
z1f39d41819b8910297530983d7308a999c001d1c7c15a52ad238042df2f13cfcb482d9f83fd7d9
zd6f8058412db4061b9bb927710c84875c69ba2ec06e231aff5140bf6fae77fb4e534d0c14d8be1
z8bba66739eea4e90df5a589696eaed68340cf6d97a83562392995cf11c96df608feee3ad04d522
z322bfeb6735f16c5cddbe2f40ae744cadb25a6a6b7fc8ba6520347602088ec5b4cd83d13047896
z9ae8ac378a4d43bd1dcc3c842da24815ba88220e03f9bf2dbcf4685717db98605abc3d9f8e8909
zf2a183781c00ad3db709792e27b181f98301462e0373dedbf534069d911b7c97b4daabc3e29017
zd0b10bf897d6829f5a4a21905c8637c3c61aeae922e3475790dfbf4057380a58aded77ea3ba538
za72df7837cea5260f2c808fe39786be264d0f04cd10c260a912d915b131f7388328f2bbe5b2b36
z303879bd051641a3a8185881fe7068e8d1b818cc0b63eb88a3e1bb7e7da2b5294a5d6559c84fda
zf99d5837acb70e74c320cc87a867a4605d20dfc7a2aa2dd57971a7820c6121b4be038c01f6b06a
z9cd3c0f2f44844d3f10afe72e246cf6d55d9a2cea585132d39e56db583819d0b542c1a8cab0e43
z1a83d2e971a36435d8e1459850ff6179385dec3ee1f237d95cb30347b65100215e78dcec50a5c6
z5e77e4146e824ff1a11e8483ff8d09fe5318942fe76c664468b8ecd482b1b2b63a924f1be7d4a3
z57e2fe5ddf64cb5e65f25e78ff46b510d2205ce1829c5c08e42a12e3656aeb8dcb8b730fb35340
zb76bf384b4ce466d5ae2e9fa65a5222743afe01ae7fbfe6ee99438ad23039171959f6aec9a18f9
zb78d38c8cd3b4ae6ba2c16ab99fc24df6ddf0fa49f832275c14378be115c0ce550bfdbfe9fa9fc
z9029c115c372697e6f79bdfabb352d8ed3b51b9ca73f5aeea55b879d91693aa5e9cf66e205bb7c
zbe9b7953f7f8ff42c507f9cef7e1c92ac994f47334acdfee6fcb2b1e512bbf48ce155864db1278
z04d30ae23b69d15e40e769a0c91eddd1984c7e352ad85d7ae7940d80ed8036a2563b961e0c56a1
z220222cb2e3c54bbb0db9d96cc69a8331acacac959cf21f4b844de646c09212ad77cd28fc1f34c
z3922adad03bb63d5eeaa6494e828947edcd822e86ec1249c7df7508476427e9b82825637d8b9f8
z60910a91d6c24c9e7b6c8176b736d17b3d580f4ec350aceffdcb94f4ea3de8778e56a5b98c5017
z39a7616784ac3cf92691eb9e96f18e0565617c79cc8230790d20d86aa0e2b31ab3701d1dcc1e6a
z63eae2da32f32a99945382304da03fc9cc08a27e60e0443ca49c934d64acc78a16cc6ced6caf8f
zc29bd22abc7f661fe0403c5bf31fd0a82edb0fe6ddab37374d929afb5a79404c2a86c1fc58def1
zaba09f802770df490c2433b4c2778e225bc0babac62a381c5fef480ff1511fe603b83a197d2c0b
z86cea5a2bb51ea09c699fc002ba1ffcc70495542c84012327bae40a24020e718c0900c77085720
z241998c95b6569585b9ca2fbed7ae4c58826040b34e80e89b8cdcb007e815cc67efe50cd3d5aa8
zdf0a50803000ffa9da200c1c7a759ec4efe32a20e98147628009eee38dd0f98ce35577fc180494
z3446632c70abee99d43b9b0e47d36e6d8fb0b4b4b32a25e46d339968cbcd441014902d28814f79
z401960fd067a236243798a827b0ce3626a2c49a51f981846a77098518230ec5402aa3c0e24428a
z03b8390f9350406e00b32c5aa34d76e69e9bd51f161184b04007c092761dfc8a168502f2930426
z494ed7a3e45bb5e12f2b5af55a1d45a80a4404d1b024e60cf46fd31680bbbf142d2212c855eb4e
z745e21abf97d569cf1bafa08c15c988e1bd7bc4a630602257ea0490fe4a6ffe82a57c04ff892a6
z364802041356a12072a966097b6d1c8e7aad8ea7b724a9a7fe6133648286780a69f25294c4461b
z5298774e22f0f8b9b02563084f3937064028ce0dbb6e9a16649e6a92052804f6f0cc64928217c5
zb13e4d310f5b818b4d9a02f854b9554e50b7675eff99c3aea590babbfa69f78b3aa798bc3a44d7
z3f12beba777e67b5ba3829c099f152920abc192b3304bd0dd96c4ea428fd276ab7eadbaa31457a
zf634809ef74bfd0110dd11b06eb2b988d268820b5a4d84d85bd8f5a0f6d2b710d63055d32b388a
z21df50a6d467a937d5e6fea98cff715ca08a8be2b51518ab43068f5a2fc93ad60586d9f70a6994
z99efb6a5d1ea9f914f025e4c2c569114200504061de8645df2e61a47f61babacd9d2e73ec52a7b
z1ba279c84d67dcf88fd6f259e6fcd6570b8c744fa6616c9d9a5224ee571a81c9bcc85ac4fef2a5
zbc9529ee19b24da1acfd351bad846a5d5cefd1913e6c92cfacd78294a04d627383b60da76d6b0d
zdb7c1b0c21b6aba6c2e54046844b3c37d7383ef74a37da35b995342d4e36868a81d2c12d5230f9
z50d75b54da0eca227d4b4bc687faed7aec356c2b6440a1ca877422a4a0892255b5b89eb3f0a634
z37912f7eb1b2310947718600b78ae0268aac4ac859aa96172f13a7cb1ac8325c821379e597fb4c
z04102bdb6baa7e5eb3263f6be0d579bd405aa8c506588d4c3a65c6cd50bc99e8f2bde329f6d379
z730f77d07dfa8ef7fd6bf069c3944ab1980c10eba01b6c279b9826151ca0a210eb01f928d738e2
z3d0e8fd1dd1b7be1192db523ac4ccd9d904f224b4a31ccafbbee10ed3a3aa5109d14d14fa469ee
z810b382a3673d5a5cc60f2ae137e6fff2a502bf19740f0964edb4713877b52243b86f6b22ff47c
zf35a8c072174a5d3984273823c1e5c5823dc5528252ff9d36cb2ce7a921f328e2ae4a3d3913c39
z7c406cac40708998ca2aae1b35f02ae816474723887fb3b20ff1b207e66c66ce5834ed549fe1db
z9984d07097dd1a6e9fbff6d94c614b2617282ccdc51f57c5fd8ef6d48a147766a27251b5e7932a
zb07f6fc066dd43fe373eb2e95f3c32c52745a83ebcd4358be63c989eea313dfe22c7feaf3ad6db
z9fe8c052336d462df9b49f5a59a2fa0a368093634cfd1e0f855d3827d59982eb8f2d011a9f5624
z016fd1d22c40bfe0eea9ee2486cdc53fca7430ba77e06815b602a4c251dedff1ed1ab03a4ff714
z6edc4986e142acef1a1d22cdfb3e043f39ed3f0892d4c3fde7371a62c00c33c6ad3a79f84900ed
z0aab55a5da724505efc2b4600e47bb1baf568ca91cd8b29342ee364ffebdb5a15fba8e80d6fe8b
z1d7e646f3ab92147a0b7bb297d0dcbac5a66880875e59b0ab70bf4bad1902fcaaf89c0338202c0
z21ce60aa26776001ce3e73f89f2105d0a26758742e08ad7a6d3e1999ebdaa242324138317b361b
z50cdb93be19193f658682c49599ffcf5ce8177af873ac1a33ea00a260a5d9f27f7e207fc201bb3
zfb64b2df20bd01fa44a12a67382a4f3f520adffbb2e714e5ec36f02daf8716c4fb7a996e26647c
zde2fc7f91c18db926018d797bb4dff334db3da1a6ef51e8ced0ca6c7bc47a03ab1efc9d02ca5a1
z4c58c55d42e40ac6a6b4c440c1729339bcaa560beef92aee88176754044a6e884fb6e2d7db5639
z3c54af13a752fad9152d7b0b67d6bcd7c0420f692ee695cbad3fd99244836a6a933c4c71d475ad
z7e03e6e3e7e881008b2caddf2e8598e1f2b190f2015563a775245a0db27b5772fefad9ac8eec95
zbfa8a8bedd69a2c4c8a6028bf427d39e2a42b9aec9008e5a566647f451b1b442f206fcf737d6b4
za1294e5e238625662799b2f0f4c24e153b47eb0b4701eb0be5c4567b2062f95d223d9973124377
z68d20c6445d64cccdffdb508eed1236ada737797e83260235accf9b88be46f90dad10f038a7b90
zbf3282cb8d30b2eadc8f9f04163340ea952a2064d87a45e86bd46a525f63d30f0404e92da4794b
zcd106794e9421d05453f8595ba97c36e4a7a0b95d5f6e64d5104ac9fb57f6e7479a5e119f7567d
zd4425beb61e8b7180fc8bdcc0fed4dc266fffa6865375083e547d361aedaceac5a28934ea67045
z03e8d3787f0e6ba359f71161320414c5dc4dc9a0218084d896d4a532e50c46c40a6e4a6ef980bd
zce38ed709429f5b6588e17461dc2e14b2f8896a92d695c1a5a9fd57376d23ea9c9dadbca702247
z5258c56bd6a9a875fc9fa592e182c053ab73cbbeec626f4aef969a838a14fd45bb540c9b2c48a8
zb7b4f1b92daadd297a3193e5ba399f56685b61c2ef3e314703b3f87d17950581ffead55ca08a81
z16ffc4342565cdb2846045d0e3b2f7734e767cdc94ab1599ffbffe8c581de4f408dc341b8272c7
z9f7ab5b3849ccd03b358a036796cba5d6fdfe01e8165294c2ee8b69b193a79375f54b9dcf5c2d2
z524270cb540f37108c6d98418bb8aa2af48ebad702f1d7b110d2970d49031bf64af6a78b5e7f58
ze85c7198dc385984e29894f793b59aeae7119c1dff6f4a21ad2e374904e6d920e32f9206208c05
zb951e3ae577ae70b32d799f2b099cdcfab8ac5fcb455788298b1f8f39059412590da5b1dfba872
z53d300d656f43e8cb54dd8ee4f64cd5ba65ac390b03d9c56e26756f3e9afb7ae16c04a7e1112bf
z5c1c870bb1ff62533b911aea04e0ff6ac7844a201696790968a85e4fdf6e44c00a441b32a7904c
zd2aeffb417de9ad9a9d21734682d886358dea692e45e9bcae40e508c38e1a2b2412fbf192440f2
z579ed2c6fd0ffcdf3b43079b21a99e3222b0c4a004ecd8545997b49369f6e18fa82c5b652a0c0a
z42994586fe4f8786e31421235b1f304a3a480adddd2532e2af81a4ec4e6161a4281eb7b95eba21
z27df04bdb6f4a1f32640429e1432de8971fb536fad2373f728220ee379891276e682c97406a2c8
z57868967b83bef7bc129ab80961a34a46ef5abbe53d5e5ba112d61abec6e25babe3d61e3d62bac
z6e804fe65d7f9d1883165328583fb14d04caca8ad122428a3a2d27c36bd53d55539561e9595df3
z8a11d712504bcb5d7ff09476f3bc662fab09b4e165500fe045fc2ae445e6d12ed0124308e230ed
z9e7fda392282c1bdca4b1503c1c7caaf2602a296d5e93bd49b446b8e555076fc06857b94129c2f
zd89ea302486f89c2e2cf6b2f834f9d19e8d79f7f8ee237dccf3f8b7da35caacee3700cdda2867d
z7bbd586ccbe1ad628f729a8a49b1b23c6012151e19f4b9773850c1820ee56bc229eac0d6da60f2
z091da959b5d7e799320bd57a210aab7f7c7b6607acacbe399369cdd1c6b59ce56a0009901acfb8
z5fa836af76a49064e23fcf783b777faac6355bf2f6d70eeb6022ef40ead5f7f374f100107ae8d6
z9d766ceb8177bbd1d45a7026145714c07ca8bf511fcfdfb447a82703d4b9a2af59919b3b232e57
z3bb9f5a704d5f1edbcf583c04f1d662e611ec85f270cdcc96c297b77e6e5e837ae803ee60005c7
z2a1c7d02fb84398dcc23658b095ac3ab9cc78fbeccdf020a8ae2ee79fd76a5b6fed47a579369f5
z59d2a032af82b3291e6b664549414c023f0b0263d6050957b680ba1b00ab4cb2dbc7fd126b51f5
z49a80c9cfc898022cede7e26a1a666f049cabd10468f502797420a678f1cf565349c4c501d4a76
z56a35faa2305fb16d8f913683355fb2aecb0ec03dc34f91519e9696d311aaa67ee42a1a60e8913
z28ad95dddb13402878335ea017c9dc1604b0e2da5cb5247d512eac9d3716db7a23b64d11a089af
z15ae26e9cf9555dd5deeb9d0f4a5669df8d5587f77cc9bb9767a01cc411462f985bb39b27b030f
z701f6c68a227044ffd482004a8a564df4aa18a06b0fcc8fb7e4fcb46907f6d57d3e92b5149990b
z649d771c0626fe07d5b06701713d44dd24277fdcd50a5f48df2a3c914516389594f30f6d899075
z3ba3dd5a640d353fd093af284e0e37f0447968a9fa81909e191b73155583a01e7346bd1fa1786a
zbf3e34b78d6afffcf1d73a33184802629f9bdb6bc54cf077b7762790f7f2f92385f847350dfde5
ze83020ed0d6e3ab08f6dea318e40fb82a87dd68f843f9e8ccd5627ab0943ed70da314866a8defa
ze8c2e000d59083cdc6aa52dc27c5f8cae2347094419ce399ab95a7b4e86b14b20cd3c6d8f0c467
zc4c1105e375eda602b98b8add0f32411451255143450c7a244a43a4538edbebe48604e5d1f3820
z51c082c0cdd6e485ce4e04dea38caa33d417b61c76e6197fd086ee544eed96ae702580f0484a5d
zdf5c6f2b0d3b966bd957be04022d88a3942df41f86f52ce2dc6b1a210a2b36443a26dbefb0e7a8
z5c055cb0b66c4c716d4463a1c6f4afdb0b80a7af89f66a4f41a7db10b2993e28a85c4129a8b1b6
zd4d49c9a4b92430a01310e3f5048687bcca611d28fa65159546bc2ff628eb61e76e5444b7d81be
z4a38ca3ed05a8b8ada50579243d68f40b8b540ac56eecdd03ab8f358c6e92989bf54761e49c330
z2675169c95c08c3f67404a2ba7b38b9145f73c75d998a565875467ccf7aab1f298a84c8efad2b5
zc1ca43a85059889c90557640696ea91236fcd6194c994ec09e496b97b20feae6d883ee515ba489
z4dde86aa7d3ce1b2ffec4bc6cee32acba3193a8fab2a34a2dff77647f6bfd05a8e49f14853dd87
z29796209499c2e008bf047dedc886e41fa791104953a66bf9c9b2b566c662df0e76cc7c86b6a49
zf283b2122eb44dcbe7495ef03241789b940138546c77ecf83ec04647959e86c73baf4f78056c2e
zd7a20efc5407cd3cb96726479ba680797d5243fb534c5365faf92fd6cdc8110e78295cd69ccbce
z5d975597234218682991cf77be4ba184e200ebc271fa8803b1a4b4c005e352c81d1e8068d4f8e4
z089f81b0961d7aabc86b3f860b83a4da882ed7dfcdd145aab106277ffd25039cb1bcbfefbd9292
z4e0b7ec5e927465ea0f36f36338514b1d2536ee514d9fbbd640c7aa3aa1db805fedc4ddac4a02a
zd55e3dee413e2b6422742fb3110290f20a02e234fecad4a28a6f11c9b83b16cf0c13d6e4be1ca2
zba05e62adba888329553f5c2b0506a190bdc2b80491950dcbeec6afa8c21aa1e68d3701a93ebf9
z7527fe4b36a689cbefbf0d1525c476318f32c1a12e079d6007676ac881436aa2e3497b00ddf482
z2d4fa17c4f0c4c13586ccfbc5c05dce06cf80a24f3f2d36d7c7f6756492d3dfe18575f98ba6fb3
z3b09dd5a1537f03384e21948abd42c0cef60a85bcc80088644abf99446a71b850cf4515384923e
zf02fffb2f5ef1a511d2980fb35592ea97f29d084cdae0b2b28d67eb77f5d92f0f28c59fb8ce519
zf4f94a37af1929213657a4fed00afa061d9c97f72de677ccefc162918107cb7a5c4fa8233146d1
z018997837f08f4e3c03052e669022f3d818774ca3614fbb4a45267782635550ef52455d3d4882d
z7492d886fc8f391b0ed827af8d30aed4b74ef72c483d9a7e8e0aaaf69e64c9e26c1c50a62308c4
z5fb6eefffccf926ddf359a9d11330afaf336b908d53075a47948f550f231f203f6fb7905228ca9
z1d1527a12bb67f0a4dcf04648f8ed530a8323154de7242a71ef8995b77c61a415b1d5eff543287
z14340b9d9d2d25b7536a455f61cac9db3a07af31f1419dbb9750934c4fe15797c8448180822d36
z14566b279f5d5d3556cfe32c99e16ca88c1cc5133fd50615c706017a916ba9f1df3c5a53cf82fc
zc65d50f298b5a99298a3e3ceda34a5da4d8c94b240f8dd3bec8302cb1bde7637b605a815089732
z38abcdf744f8a6d1b49e9f4765b3212120581d9d0460e04377397611af76ca8ee3ea1ece3544ce
z1656648277a46e0a94999076e09154e5202d317132a33b178fac51ed5b9c3be00c3a2210cc9646
z52e61d0fe33abfc9be997005db1f4872ad790550cc891b16ced51905d47b92bcb52fe339180251
z8d97845c3a6a907410b9419d78e4798954df34a3295e0d1502cbc604478908e6acceb3b89d2d46
z91ea8bb27a5bd8e32c2dde0b58df0af9a9d8ccf5c718f92b6c75b0345e51158a860d15cf37cc58
zbadcd203deb01fcfcbe922b4211389f846279b128349016b9a7307103ac5ffce6c80da808f9d79
z5e49a6bf528c1b237ed3e4e3956b8461c5eaa9c584433371446b037777f90df16dddfe9c0e61d6
zb2e63abe52c120bf7bd69f0107be32502b9b350cd97707bcb025f318f8066af8de49102db6a908
z65b31c29890db4e6bdb25bcc5523569b1bc519c833e8ba3cb713ab07e48a5ecaed06a3beb1fc3b
zcb30cdcddd9e2174fa0ac60ab0caa83739f5a0057abacee2d378016c736bfe08bc88d89d5ce801
z08c59856e5651462b6607312f1ccfa4434a4830f7b8ccef1ecbfc34a9083b2b71b7a3e768ffda1
z110cbddff2d10a9d0fa63041d3e6af1e75d396e1457ddee57d148a13c4917286347515fad5bcde
z4303a6ba78a2cc9e4f58385cbe437f48df7d57843342edfc73ada8332ef28304d545ab7974ce21
z4d2cf8e43e99774b057660e814ff1758f5b23b1b957e70898c54548d466e1330f98e95023ddff9
zbf8553032d33a2831357c7fce6b7143330c9a233c29cbe1b98b6017db58c0faf1a1a22ec0fdf59
zd6b324b76eb2be0c25d7065a5f41fdda30ca3e894e3c91ad94b56b12e13c72b5f030712b747f85
z1a752befbc55474abdf49235ed8a989bd1a83e379288d28aa81ccff20c9afa542f04da6ee572bd
zfa7d524822b9921cb32d611185927d57fe6c44fbedae4aac135863f94e2c189b75d95acff5ec8c
z282f07e935e78be66bced34f1428877332777f5ec066590b0c600cfb4e34b7a0affb23aa3de47a
z8a0a0e9fb202d5347e6084527899cc010fd167b5e5d07fb45523dd87f406d453c3433d5a52804c
zd0500bc872eea2a2f98f17178276609f1420adb0a489b33b2978a4a4a8c00edc8b53b8e793718e
z7903055f08916fe96ad9afec646beceedda22fbec9a50a27dfa749687a38e273886d4d6ef588fc
zc9e67f8e64cfd83139765d060a3949ffce7b985af1b4d7e3b57cb3d8b5a82a44fa2ac3f6af24b7
z2cf47c8457c80d6b8c63d3821fa1c3a64f8a2a0b4dd511128165370e29297d9649a5f9cb2b6835
zec1ff2808f2b57152d84ea1f81f73cd14b52d08ffe47e00c01dcea18502abd16e6e6accdfa9e91
z6ac78e26c2b81ad6c0d353692902cd18ae97a379ad5df9fc6e0c5ac6638c6e6012699c103151bd
z110616005af870aeca2120f0a86437156e11441654b234db4688d03f9f3261e73e37cde5f45328
z53b69ba335610db5527656ee277e6a53c0340445d7950a424103d67a0692ac665eda7b19e881b9
z99c4e3bf96135cef28973d8de09dcec524918a9657d266df7ac84fc494e90068edba8ca06a7561
zd2d600507481d3f7b33a2357a5a1e459c73d7dbe8192fe93030efdb71698bc369037da8ce68a11
zba32486c9aa2377e0af75eaa4f9efec398eed61cc6609061eceb5e24bdbc42079c240ead6fe4e3
z90feb25a275e50c1d9ca0720a41807e2009e6186f4053361234676a3c2ff393028564b49ce15bb
z692986a786e4e425f27aea6899cda6056100e6eff41bd8efe099af2d52ed60495fc12c0b9dbf38
zbcc0e93ca45ba91bf78e8d45f50300a311015a3e18721c28fa23005db4ee08ba7b5cfde31a938b
z856c69d390d17a9bfc1e83a648ce2caf4b952611ec79f0e86587000f522520dcb3149c8be6da8a
zba476e0d4a76fe27370c1bc89c72cea262f1e1420713a495b20e06e8fd0707a5e6589447b64f89
z4b5cdfd72ce7e5310fe26360d99a9bbed26a3c7ae70d14ebce628189b94b2ba1d5d783dccbc652
z7952250e2947f7a6bc83a6cd5848473febcfd61740f601dab47d4d788fbc277a43903400048b9c
z102b5b8b776c6654b8472bbaba061305dd704a5508bd365628f120c32c0b90b1e7f02a5c3f511f
zb76c88832ae36806dbabd051f038d8cde5c1215206f05895f4094ddb817f35858ff9936da7c4b3
zd7fe330d1830eb20bba558edf0299340fd1d140c960acf3650e17b9be3ab7e6ed5fce7da073ddd
z5b9e4035e75560c249192804d73eae29fa0db08cd7594229d15488c487d118e90619133d9baf04
zb84db75db287d66a0e688870b14df0fc8c092e486936603f2d8fc412125ccfdf9a01c04cef4cc3
z108d9073dc4b129cb8a13ec8d15da8989c64958ee16a68697ca4735f684171b224781538a555d1
z021ac1fa08997a18005a17f7bc63cae3eac11fbbd67bf86535392f2566af0e320b100f3223a3a6
z34e7c07470c44c9274aafa0f5bc1240f50501eb79d27bfb7d4342a89f87f4ee80036eed6218025
zf4c5620bad0221c9356edb2303db9c281bc67ff69bb3a03fa8f8779081500dedfbd15925fb5324
z5af0d5432a243818190d770baa4c524284fdf6f6ec12c5509ce83a6476b07af4583108f367e4dd
z30392a02c0f74b44cc571d9d9495be5f5097143bd24aa532904e7cef67cad004a9aac913d3b697
z727efbab9129bd6cf9618c474dcfe9cb32054eb9886987693d1e0c43da1aa7523320cd1f60edf7
z0875788592b32e19c2318c8a8e81c6fe6014e3a721292c399cf3b2e9ccd3db392bd9267d6e58d1
z1e67187b3af1380594f69ef980bbdbdb5af26ac7e2f9c41fccdd68a444bcc08156e4cbd6a57664
zf4456663008c8ce82de41c5c0ca7b7fa4db17653d1758190023428933b4a56c78ce7487f0f73f2
z4068a2b835dd7b05d6391fdf5684b9250d197b93a741880429a2303fa19f09f23c3e47fc6ebca2
z872152901d5315caf1ef315a9219da0bc050a98935751f0c4371ed636e3aba945d28983921ef32
zde67caf8704234776fb0d38812ab60bb3327a870b09ce720848bf924a860a731e8cd959d20094d
zf74be57e404494ab2f2e7b6d4f5ac461bcc15336ccdba56ba6a4888ac5dc1bcf3bafe451beec1e
zcfccc519c1325993865ada01938d1d97d1b26de8633e5558d8dd0e39f01359b69fc0b706b69db5
ze9d709d6c3e115dc0b994d85dfc39772d54b3917d28a4c1716382ee534ad01b5375cbcd7b9a883
zabf634277d70de982bde2dfeb14a343d54c9828b7bdcca0e22476aceaca5dd29f0785fe740aaee
z98185281c3f9d8f1fa38e6331fc676aed77c46df3ba453c3c1090cd88ec2e105850c3de2ae0a6f
zb66f176466e4c65a806ce0c8475c3326443fd2e4f3e47404df5136d0f7b81d3bd0f61da0b3eaf9
ze07415b0e002412ed5cee972014de66f142f4f0fa746a946a2920673fd550288d7c7a0562a8787
z88bf583686499a5bd939398bfc744dfb8f70086dadd7a485158839f7b9add628257c3349d61eef
z7d35222a049588d7aecc9ec7ec25429d9821f4c04c84f87d29c227118d2a60ab768a62fa3fd2c5
z91d8444b12d7a0c5489c1c5ed6e7d346e8ffd0f6b9e5bf7ef74e1b06b1250a84b417f53d465df5
z1796140e2417142a5f3950562c897ff2fe82336c73997f8739d33cebc9fb36c6a6e23ef5e717a3
z7244a3b22f897938602dfc8c9fa6b030140e965dd24ca5dc002a5a35e24894c1331577b58654e4
zdfc92a263886bff6d68d0addcd3a59fc2f3c7367347735fbf38d12eaae57981be4205ffdbeb35f
zfdd0dfc3d50ce8405d159d7df9c9c2ef4c64becbf4c5330d8e88d92dd8da7ddd34debc119f4bc1
z05d4a01ff81f3d4f5f54e4294c26291677684db059330b55e5500dd9b0b498cb740e4dc2ab14db
z1049fca5f98e68eb8685519c17472bd3ae9a665e8e092c03961ea332ba4ccee19c2155ef8421c9
zd68a3549a581ec7b9ee141c055b3f4a5afa1ff4ea10174f904aabff848f91c22f4f022f4a69c2d
zcb463758e41004515ce1827c4ecc74f3e7322e3458b3cd8ed8845f0be271d10b235b9807d0d494
z562ed2339a86697bdc530caeca8c351bbee02bf865618928e9adbb88fa2bd757620537d10f9c54
za4753b7992f50344865e7c404ab4c3e2299e972211bc58c2d0eabbfcb9b49b300420e4edb72d5a
z22c7edd75aa8954beae63a0f5950f68dcefddc507160f3c9168ce34782a818053451075c4b4d87
z08491a805da4db7369c0d29326444adfeb97fbc5a05c24fda1d3777849af3bd8fd30424f712c0a
zbfacd58ab8ee49322d2ff5dd159bd8e7e238ad257356f07d6a446290a77c00a24d67ac8f736bfd
z720d1aa0e78c133cbcbe8269f0ffdde25e2a96d9338f5e1ef430fc8f47f865f648d6ef239a9ffd
z781fba3e680002c24a0d9fbdc5e0411aa2e1ecb99bf3fa2ce5ab8a7f79704bbda2e80863c2eb61
zf12e2218053196c252db39e74f39cec320a954e363d98465c5e0c086501dbd08c29f74377522d1
zba16854b173c62b27cef4e0ec24b6e5560ec151ef2d5a296b9d295fcb1106f18cae2850df72dce
z127ba0bf804f18451a7654d7e2830a89697c12898f86b27bfeca34bb9e5efde54e77c11b10ccf8
zec58ec6d19c1a306a3f86557dcb77ae92a636f466356d51aab00ecfe2ba107bf038b54fec345ad
z2cddaf29abacf487027eec68a7f79401a7d0c115229bf59d251040879aae4e81b6a05f6cfcdda6
zf6149904cd481d515d8185ad6c8d048ab6eaa9350e54563843092e78e3cb30e85914be663a3b93
z1706eaf0b2f9ec3160b75e470d4922f5f3f89461ea92958b07b2ba233df5b77c7bf0e95b6e4dcc
z377fc34b2a3e27842db99e2dbed9da4902e56e4c22fc649fe235ad31ea3c9fc4235d77f7c6c94a
zaea6853086c5b0e8f3f7934dc8a44c2fe6ed77f5a31fca5b485544aa3cbf9d052fa4034b78e02f
zeab3902abffb073439a91a7e6e90509016b93c00f56145737d2be138282a56301413a5cf831c7d
zb9aa5ebef20f88fb22b54dc1dc40539fd45869e69612581852d1c5e725bc7059b0404b1f966099
za93a53e34378866d8437a5c2b77788e1b0eabbc602a6b547a43a09ac0a19a0832dab4b3601f439
z42e97638ca106f1d83116d1178783c3eeaeb6290ae2c4168acb65a51e33eb99c2a808c2a1323b3
z5b7055bb38adbbfcc90c56222d2348cc767aa9c0914d51c9f7bce81fe17340a46183123f4cb614
zef8d5a602e3c3aecd5cd04fc9e6effe0cf6f8c62f03eb55626f282800ec6abe3d4412fb4e17a3b
z153529a69a2e1a25dc525dc935bb4a1c23757eae8216365f4e3e9ff466547e7f9a1b3a39a1fbd2
zcf18000b09853aba71490003f8d00f99b935a43a8b6510d1a0d99f88221d9d23b46d661ad604ea
z33c37c9d0f84f13308188de630531e123d319c8ddd23d6240d0454ed76b3b39f5f65f66d162cf6
zad4a44a77ca2933875278b8011ce07116b223bedf03fb4bbc2863eef268c2178c97799425483c0
z9d7fb5a1587b382a3a1844db9d4807ddb6e77693949ae2b9e0b5e2ca4df7340b2951532e991af8
z2ad41112df0bb7dd58200f6acc3e38cf8832d8d53d41a6ade485bc4a3ffe3c1b379335961a4e36
z81631b6dc93821f58c3895ff7d9a4a70088cb44a9ebd80cdb558b7e020379b1fe9c2458f6c45b9
z41900354993e7d0f4be0d63d75402433454605f04787c5cfd1999de3df7812aea3c091beb94e63
z6e83864c7ba2deabdd2414fff849d736c8518c3fa735effe7ccaf0c536e070e2409fe5b9be30cb
z0f0d5647c1d94e03b5d4ef4959bfadc7ec0f3542dd8fd9ce250572ea7f20b99f46241a08eb65df
z498fa374f263653163856bde3a74fd6a8434784a6b183c9ae860530a15bcc0180c38d5eee757da
zd2a27a276dff010437765d5d16b17a730267fb5641b03e73b3e631a5da403b347e93890fba4de9
z3289404445bfa900351e302dd106b4f5b485008cede24d7caa50be967f61232f6d604fbae35308
ze28f0314f9eee3eb64b166e9c62ddef481034d239ff5eb69523385516b00d1731678af7861a12a
zdf8a7a889a8299b104920d0ec5dab287b3b031839954130e6fa11e47a84b81b0c648239ce2317e
zfb07f97321ec88b93822e6e4a59b6c1548ecdcd87f8680eadb54d51f1ded67d3080a04bc46b8cd
z486fad358157f95de22fd8b9b78e32fb440426f61ce401cffb4d1b6ae1e5b4765b32887a43285b
zf42ad6f8cb16ec6fdb1627a1365c849e0e35fc72d2ed9f7b035ca72e0fdb05ec46d516accd55ff
z01b96bc59d635cdac6d827fa8336e29f59886152495e2f5aea7f19bc545b6ef7c17042c83e4ab4
z23c514628976c372f3c6a90c5022190aff5431f55def44169df705db44c9c6632719a8aa56bc15
z9cefc6bd4db34e4e086004d7cdd91e4d0d2a6bcd6bf27f038766f23ffcc87f589749a06e4bfda2
za65401d864fc58e88f1b04f4a27bf4693011ca3ccc8821c5e7897d62f1650c3b09bf5891a4a342
zf509aa75081089d3bc5abde0697f57eb8848f1cb9582259d902e422c80468e2363f317a9d417a4
z5f62e2e5574ac81afafe241e64051d75aec6c264e589659e5632181fc9e999e4b62315a661579e
z7e4bef5340bc76f875e7a35f2878866ee25f9a69bbf8c2fc94a11883b6ace0c3e9e7c4113dd5cd
z53bfe632302eb7ef7e234d4d2d0c5793338f73826ee30f26ad7b3bb013897b92af9dd756988be6
z139ce0b7ff7bb07ac2a84673bb29adcb556cfe0dedab5702a5830e955a748a1aebd8cdb5d3f01a
z25cb8a5a161ce8e70d2489ea6f2cc48a38fdd015e8f98b8e844db3beda1ea6d100d534194b6a8f
zbabb926c885364c2d146ca86e8391849541a8decdb4ad19de8ee92d9942c62a77afba38188cfaf
zfaf7e9b5e6f67010bf318075d25b61a30a26f9e9421586dae45ba89e2dd35c51ace179fca55fdd
z91ddb0d373efbb0fa9ff847d75cb3887fb578904d224c318582d0d0f523b3c04d27a2ad7b91c20
z04913e3b0ef23eab491656407ed07f5cd063c608b3559022fcce3c89f28d1f021b4979d33a47ea
zc05bf108d268c27b8b39de55ea8b54754e549f360b929a27de62a2f5b76dff4ee58decfb0bbf82
z57478bf4c78bf3978a6786eb981542f0db8cf6d7be60a23f351707b4d0c60dbd772d80a82ae406
z29680a0d0c436a2baf804635ba9b1fcb25e3c07610b26038177c5551b7dd82791249aa00c7d8dd
z1d24f8b7325f02babf0d118838dd83cb30f44d12422952ee3ce014a89445cf520f9453f197a804
z0a97aa2b2391d07b85d272dccd7f4c9a4d5372bd1558afc90465171adbaf3853bdcd72fc5ca123
z4ac652b1c1420226a371fa8f9f70aa22dec23711884b17ff0716da4cd7a8d3bc97aa5983cdf663
z44bc188c8e22e8507f48e22e56bba2aa2232993c8c1183e31913b24c2a57325cf23898503a2bb3
zc014cd5e110296d2aa853f3267b0850ea8affa42ff59a95d3c62cddf9b3c64b2fc7faa1dabb5c3
z51c5993fc87e06e38edc037c6775e345ef03c81d2ad4ab9d9d01d63b85628a17c22ebc4f60d8d5
zdae02c2ca71cd0e15159da1209c7a889eb0e8c93a3c2650a2bf3f722dbea9d24713c64813bcc2c
zdec1b1c7f9c72110fe0b5c9d9b958be984fbfb233108cc172f25eb288a8fb3b379a3c6abee6577
za0d926986a532cd7b10261366b37b1ef00967ea6c7b4c896615d8bceaf43a97523e2d5c6664cf8
z5e0093089ad1e5e29fa0fa0a5b02a0890e38c9105e9e76a55a767857c44f5a91c65f0309a19bef
z3660cf2b906d53f02909d3ee724a9fe65a82e188acc90391fdceaa4dc0b75eee2b452d5a7a636a
zcf1d6442797d90550b08f8ca58f2d84ef955c6fd8d4f83822dd64d4e012d1f7355209a7d6c778d
zba67f6553d51daa2b03bc337be20645d3014729f7ccaae4f35d5bbf67d1f9c0363868179e3273e
z18d1fb8eabfa7122c6db04d98c9421403268e8e20fe1dacdcf44104a5952fa2af152b7548491e5
z725ec782bc878e20e940c44bbf5f8792f58a8b725b0459535fadc6336622e7815a0aa834ad5fbc
z0fee1e60d40abde94dcd7328fa916631acc3902e3698623e3655e29e5d1072dd42364b7a9fe3f5
z431a07f1d8297d601654bbf542caac0a95170509de5d5f137fb67d9ed0d618c696ca6bab73a4d4
z165d4ffb6d05381238d711b6b627cc177c0600a7ca43e92ee470552204e33f86b3498470caaa4d
zd31e8dbf305c52eb85b90fcb5db5b04c46af0060c8b3274261e377c90dedf0d016fbbe2d2dc38f
zf360c359a0dd2da314b0273c1503ce936afaf8b5f5e62a4e543008929ac7820185f2555439d28f
zd4e9c83e57cc418082ca68d0d1dbf314ff6fe8fd87282a568401ba83aa0fdff9bec534a24b4831
za51c504896220192cec51cb11f6bbd8935f8f9acbb252c4e076534843cf1f94e89c8e039c47bc7
za6fd202cf7ee99287957a10cb7b8fce55e98a196710561fb3269c349e772881d1d77bfa27072a5
zc29ad4eadad65bb65575b0d8df948acfe486aef0c127b0753330da522737d5a19bf31ed6f7ca15
zc8ae69bf2d75f03e86da610af5ad39c0e23b87108a2ae32de37f4a7867b0ae8105bf81a7e62ac0
z8b698e6027532ea517735144221f2ffc4f402174688b716714d80872ef626bead829d3054eb35c
zcb3674149ed17ec339468ca6cb2537800540693adbe6e88fec23857bf3ef03c85409c563a308b8
z43548e3be58f4e19cfa65276cbd867f5962524f39e34458fdae9895c303b766f6141615304e343
zc4e7409528b671517740f7fd90682f3ceccf6b46d43e7677a91e3d2b7659f879e25ba50c21daff
z5a6997746601e91715b090f000aec231b444dd80d7c3bd3feec004469530386e6e91f68b904baf
zd54ce61284d0f06672d7625609f38aa440e781ea094dff847a1d4dc8be741d08150ecd355151c9
z489a300238cf482986f5b7eb25ff93ace3f834a909310766808451c18515a2d9da2f913915cab0
z891b131625cf292a2df60e0fc4375216fd41c7b137ba2f3b18f1bec66f583da2cf3d9fe5eb2900
z0bce404f61ace24254bf6d23ad1815ff45c92a99b135bc40bee35533d3298122423bc5fe996edf
z3428ef37ed395967d356e6c092d1268001c265f0b3d7deec1a789eff4eea44939a9ee6bcb736df
z9eab1b19d4efee2d0f3517871b69e53b0e9a6c8ca878c2809b397562319e03f0f6af7e0607ceb1
z932324c24dcf964d63a0f5702b8a0b8bb0a1188ae3ccd9095bff381aa3aa77fb0520383e224b8f
z5f46c3cd689267643b092bdbe07455339583f7f927c18e373d61b974d417d6a5c445e5fbf96a3d
z78c17ae5fae80135de4492262f6fbcba5e80aea4a74b10a87869f9bb0a2ade048cf2327c560a5b
z4951afb3853ac57d3e3289355b84bd126f5f1efea809599ee3917a2dd344d3003f8075f007df16
zf3e9145e549f06ac21839dc3c2f59a278a4d818ea2004ba30f2bdd86783b505a52e2db8b8de025
z8c378664d2ca52285223d3d5fb1774ea4c90c73d8b169ed503c8e0447aad73855c8abb5198f157
z1460ccd50800925b84e4cd414a62399f314c8b11d2b95aa89067994a136ae45c245dbe94cea533
zbd029217e0bbc87f1f070ec0a07a0497260ee9a0dfb049ddc3a16b27447e311cc0d283bb8b6907
z03ff6b1796723d52a3e9d8bdf7d8f11a0a30f74c165aee824903c6e80183f2aca511a6125cdb83
z175a7cfe73d32d4faeb9d92ae3aafa175fcee9212f92916df8d4a352ef15e7387d9ae28bd3777c
zf78a8cd71c870a5e05d8c367e5a96d72271c4b0ccba716685cfdfcf68aff944385a531752906a1
z7bc3650ce378b70336fce863e31ceaaf02819b86a86d655938d6db523dc8e1344d1ff8d5b7a0bf
zc049b83912385c17a0fe1461c3761cded3b744d44efe2a3260a694e21dbf143d0197613f5cc7fb
zfe77ee406c4fed6668d410e43e05dd552902854caa4c85dca9842c7b27ce05b6a1ea5a62333b94
zc8dd5b5ff28d29a260213bf2d680d52e12e6f3151d0a9b83c188afc8fe5266c94acbd952ccd42b
zfafbc6856fe13b64f74e5a633f4fa197883edd91d27f0839d9449a304b64203093f4dc0d10ce3a
z0b13b0e1e09cf6075e6529d0442c316f98801bc2736c42e564f63b8cc4d7fc44ae4ea50ace462b
zc3e392e759217d4e677ec19d428c555d0b422a7372ea2c9ccbfe39beae499c3a4343999f1da9c5
zce8822a3ecb151d4511a2546c84348e27ab981bbb895811fc3bc2881332758f8dc903d522c5e50
zc7e83e7b05d11835b97831b55d0c56ecb049b8ebfc4e76432599ff8c54caef1cf89a22839f0fec
z35c833e1788b66b1ecb5a125af045cb1cd3a7154ddac5e50291db3a2885f18dd1cd422440bd631
ze29d1ad75a65473dad9f9d30ae81d094ee40c3ff0a1ab04a2b18272aa5c334965040355a4ad20a
zb98ca8e66d79c895c97f68e166677f246009eb8d7eceb30c3cd827b310219f397d826bf6071a7c
z840aa6ff9ca18d1f54a6b8ab122badb33461e8749c2abafce5ff347276014b67790899eff9c675
z673a3fc4100f2eff8e52ad998dee4e057fa21bed834a2f5b98d0f9b8be52b1d5ff1d9444cd3aad
z45e4f2cafc6ec3c602a92b69d7086c8e3029b7f76ffc5c92efce76191cd53969f4c7ea8d026cb4
z609a0b1272e374f6412c28ee03ab1f542bdda106a1e9f1f835112685388d35aa95712cf15b9055
za6c1796e704d1b9a4009b226d87abd9203050351aefdf3ca21743a215d8bcace1e92dec9cd5948
zab135ba7e373090637e24250bc905cc1b6112677df709d49755b3422b6b674995b2225527621cc
z378a70a9a05cb0401ccdb7233a633d5bdaaae302e3328914856fdc8d3648822f1f6fd449ad3997
zcc5efbbdd38cf9744c5b9911d110fb1be796324ee3242350988234dc184dd5bfa66db2f01682eb
z311026cb3d02c6c9f4510a7a9df766981452f516b74bbe06eda23c05edabfea0d8d1a0513a22fd
z336808a0ebb0fc2f56cf52e6047a257dc3a77fadb248a9649a1a7e82b4815a52ed746d10af617d
za646db6edbeaf7103a4f4e66e1698823fca4865c72e2ff9bcd09d59f42fec507df3b93b81afc12
z3fde174d802624b10665cbf91e68513ebf9fe789e044b4048cd3e01992be29d3f64d8e532f9415
zd00d74c83eafb7d1adee7b34760d54aa7c7883df62dbe1ea823d1a69249f04283572fc202ce0e6
za3a45587aa25c3ca407c4679676258268b7274100061a80ad040124a7f3b659834fbc134598aec
za4b245d7b19c5887b9575d3130321e2e42d1b7f1895b6a0531be020bcee00691d1762a568d5e27
z8e765de242caba4577c3c08d8f2ebcafc4cb28d6a6b8e8f687251cca98342131595ece7eb5327e
z715d103cf79b36937e78c1f0216c015c0262761cad3e593950852320390963a5f0cb34a636221b
z73e1096986ac1687d511a8839271c237ff176356ed5909c9e5683ce62e0c2c76ee29f77e2549ca
z91a8b2d064d73cf675c791f358a6df86afb2256014b3244a818465f74484fc4358c07535a28ee4
z07f4daf8dba60b9301b567c804180b38344a73a7bbd1801d155fa4a0a1e48943c1e81aefc97b69
za0050822c72dfb4c74da07e8afc30de27e6e4b49dd6e6f9f0fd735e01c71f16ab8d2fdc2bb710c
z929a0323a9c64e086218b5be351f379f506877e181e98061f3a61ce574adb34985bd48f94c6e23
z96dadef329f5af122978cc257623ff0cf62eba9f3870c838b187bccd2aa87ac23cb2cd777594d4
zd73aa1d44e0a893a29556afaeca9ed571f36ae371842edee52dcaeb9f86f48781d59ec60b34206
z700681c66d2d2abd44b630728fd6eeeb24b167b032831ae06fd27ad0e3e7d3f7e320c4fe6b46df
z6864973c1fec4df2231c218320ef6dae46e2d9daf7209863b9797552c297b36bb3361321ad6169
zbadadace6e1a79a51374c296b186f35b5ea55f6788220966dfb2732be5e9ea92e7b9821a3a29de
z83d880217a6c006e84717d5c954d4bf3bfc22346b1594553bdb8f3f45af653be08fa03cc5c8976
z1d6ed5edead003bba58d6dcf31d36954b86e0a4cad46bf8e172178dbaf9d65338803ab871ba52c
z583c87b60ad645a1cde78df7bd0e8a8bbfec2426406bf9bb98e31a19e16dad2c252d988a4d1a75
z9914b9ddb11e4b03a4484e5f45f04d4490834a4e445e6654b90ca2220d7ab95ff8fb0f7f6668e8
z1b622e7a55a186c7cbe95c024564fc24183736dce841dd1928c5e429d5d1c10295ce24444c3c0b
zea13d923b62d76b63c39734286eec868d2a751cdc085cfe501d6cf678479d0eac55e29c8ad86ec
z8af39f7d69f213286bda5d41009cb5d9f96fc1473c6f94b3734d9f17031cce7664867a494a8e4f
zc1b1ffaa6d914a708aff75c60201f9f49a08c1cade758f7a9d7348fe8613e9f47c8f53125b41ef
z9a04aec3512c6d962ece235a67d4fca97fc08c437b7a6ddebcb1da925e794872bc0066eab36319
z40fadb7e17e9b46e20e6eea76c3cac8dd96296ca30ce1cde3d518e21d5cc51ef6a8d0443c9466c
z29d4b0239d1bb14393517e41f8e4ce8763e520ab9731e5e639cdec748b4ceb366fe531337115a3
z042fa570f73a66ccd7c8c6cc0b773782bfcb2ddf65bcd53e3643d9b07b5210454ec24397947fb7
zbb67c698ad4ef3c116177aa434c577fb3aae3d5b281d51b7550f88d26440d7328a6763baddc9bc
z57419ef4cd73f03ec8e467252f955d5cc134a4fccaa555ee34ecb6186b17e6ec19c903361d9dfd
zcb1c759e4fb9e782ccdc4467492696a23145060efbde402218a25ee3a4a21ddfd8406e433b5706
zba3106c5e9e22b363f84c960a63f7670f480ccafa928aaf59a56f2df8459155605960fd902d531
z24de5ac845f864386a1986ae91d07f84a00b6c2c8d9fced259e392328e839531740533b7dc780e
zc999e547b05418e36e2d66655b4339fc401e65f0ff3abec188f4e5c494b6f05d06a6e1241d34e8
z6b9b686172325cebe30ec7ad1a01f84659c420bce7f17b37a9b02f4f36568532c03a1fca23653c
z0b5984ea714a69eab14db0464fd45ee84fe5c9331a53685c578a0e94028aaef30b283e53e575fa
z93867b8dfff508aca9870294b4ac80a9c429871b76f505e642b435b09e1fe4a84dc5ae77cbb1a6
zb002c9f848b6ebbf2d11efaf5d0cbb3c6152ca09b63efe54f5a23af6031a0c3437ba85323f28b4
z8bd46b0c85ebaf7632d10f926d9d50370713fddffa2b5c5bae07336456694298388d995be19f1d
z53563f5b06f4da7c31a179553fc24661040c665aa1a412816a00caf512475b178259175808f0db
zfa3b2ce045945eb43e788b06ca4d2c210b1a5dea1dc3403b2b0c196aee0775b1dfeb80187c2c75
z09407af470ac41304a2737617c0467d4052a069bf6e03ef7a3c7a5f2319f614d216b14233e6439
z956fd68f0cf1ed9ed22d57587d7c3d58afcd5b5f56a3212a771633b5026833c39c0244ad55abbf
zf1fca48fff951d8cc891cd4a4c0573638371767747120afbf52bf1bb4f8697b995089f4ca99b30
zc0295e6137f32352e00f598df556f697f2b20b9cf979def317a32b0d5e0184e3354eb9a18f5b8b
zbf963aab6bc13d74863fe5ccdfbb39522a6bf5243e67d7163472a2f150dcbac0b68e64d01338ad
z97e9b5550bad7d16c7609080a685c0517e19499d9f1e02b5abc0858100ad69959dbc1a3ba3a586
z9789ab4e46b11a299d5708933bfcb9959eb3a93e2ccc8a5b9023045251ca565294bac84eb7f813
z6422b79a96f2c44521c94ebeb0b4481535cd2d4e685bb960ed28abdb60e8c2e68f54e739a209f9
z8bd8aa530a62a101c553854f31b6183cb10f159aaf1829972501241af2fdef144ebe1ccdcc3258
zf42321f36aec2af790fd2cf0b996bf8152028dc1c2418e4b37dd0a17c54148e6b53509fd0996b9
zfcd87b93c8f901a8abb0b9c260bd4366f8d80c63b2b8ca6fa9f3cd226b219e4124d275e820d46c
za33b38f03628d5a49085fa5ae8bfa55dbfe117460a91d7d08c1c81e045e45805d9e45dd5a8a4a5
z73f78faf74019432250f87948f405537b5c29205b7da5bbc720a86a112e9e1a7822611c125d8f9
z98c05154cbc54ec2f06b81b9bb7715fcd5a80cf6e4caa5187a6dcf3dce39384e611b1c9a1bb2cc
z2f4d61cb3066f46fefac322a20a9a92aff4d1a5688e49be705905cdf6837462012d160fcecd38a
z940365b5a47038b890218fe789c71b50bce4bffeac2b99e67cf3288dc62b4e6d22efc6c2ffceb1
z3fedb0efe34c7947a761addff6c29104252af720a538679ec849e36e9ba38bc505396ec871797f
z42cb4f96cbb7794fccac50623651c29adfb2c9f234e21a2dc66e9cd172ccb4527a549ad133836d
z2e067729d5ac7272d19f1425d4ea93cf123147123bd85668d24ca4825b1285e8557766d9ea5281
z62d1c76ff15606e4cf2661790d3d8251c24fecc76d69760aac79c76e07356d40bf885ffcf1e238
zbe594c8f5b90096017b3936ab0e84b1a09f5adef483449ecb7027e727cc20b4e098d07e2e2f105
zcf991071357ee5f1053974b625afa763e840627f415b91c56a3a714a023bfb8f1165af3f448674
z74e3a6361ed8cef0ab2c1ef1f68ec5e0d4084106055de0f91aa7aa48812982bc805592b9ef53e3
z00b8c359216b7d7c2f6caee9ced89dee60228ac2a52f4d1c3a37f1948083da42800e9cfe7b66be
za185f1dd8b8e2175f0266458710fc58ae38d7f5f37b8b7803f48fc9e5ac916dbf43106e0dee7d2
z9a49dc1efdb7d48e7ac702545c235bb50dd23c69439e4e4018cf49de8f8ea026a9a97438ead522
zda4cc3be21ec2e17f0e53a7f08b66fb41ff29b261333d34ffdb99e0cd4859a4891f194f0d15603
zfb709b7e5b3cea3b7a2afaea67e540fd8cdce8f976675d9a7e74952e4b68361994642f5dd07963
zd587c6176d99751f865a1100547988c1f5a68d01b29ea1dd4ccda4537615d3c7ede5b35e73bef2
zb10d968ae4ed94c42c441afaa914b26749d85f5c6a03302cc107380237fd1dd0eedd18ecb09c1d
z795a0f92c63624061a3b7b8635b8d563f00b56dbcd8bedac96f2f29a669a4457f466c4741af3f7
za8bb986f353c936893443760edf0160e84dc6bc6c4ff66058b7c269fee28f821a9c86f558330c7
z95770977a08af13e43ff71d19d42b3e1cdc5d953b4ce487ed474e9fba93b3eed30250f8a197efd
z8e0ffff28647fadcc17a6292fcf3205f02c238281bf4cca12538b28b4a0186f42e23ce03b3e0ea
zefd85c9b8bfa203c4f06b83dbc5fb5eaa16aef69a9f117425f3b2089e8aabff40783e3124041d2
z6626f11d4a8c0a736c0f8ee81e759d1b5f92d79ccd6df09ac160f6515118f30e063895e6a5e423
z25e303fa767b8a35b123f860786902fc49ca6dc26e914712bc0df1d75f009af37a5806d01fec92
z10271ded5ce78ad3ec42800767dd080545c04440b3cd5d085daf71be0150a8d028d0e8662212ab
z42cd561a99d9bac371a7c130fdd1f4de3be41a06e72b0bd23e451f448876d2aeb0258606ca5f3d
z08c8cc61b41c7ede39e51329f263dcadabc9ddbad58a57c9802ecbb2fc46f072737f1fe38db545
za6314251639a8969ea435f23a3880c9952b9431d86b68dcaf4c11e31069cfd385dc8f95b1eb67e
z6814376f3976fbf0e42c573ad381f1c4fdbf87575a6d8c30d1f233e9df9f94df2aaacffed9f781
zb40368b48e26c8f6d391aa3fc454a298e86826d04792b498f4452f47ddaf430d247cfdc3766677
zd671577ee33023f0797bf634cdf7fd86d6c39e62bda94e5adafe29920962b02019acd0a06e58a9
zed7d9aa6b12ca116ffa548c567506e877c72d395fbc0f8508c6cf3571f1bd60d221b016832fcb3
zda648bacadc53ab16afe6bb31ed7d1def1d5906b753e4f4a6f457cd4b4bd11b869581ebee317c2
zc3b54c7108a13b6259712c6969e4f1f35db3a81bde650d9a11cf2c7e4cae307c4113be07674f25
z0d44f4bf8aae764d31a603b95bc0d065778cc59a9adffcc2a37c06cf90eeae4cdac35d61b40ec1
z75580957f16bebbf33ae75ed380006279a31afea5f0a5ec1c6e5a4f73710762d8c2a9b90cd1abf
z27ec529a83f2ee6d1f351e5d170529c65a74c1e2c47c9de222c17eaf2bb3998aeb366da20edd6c
zb5b6c30c4f66b50ff0cce239809c5996525248be110458dd3e5f98143acdeb0a0e02e5ae0a571b
z3e0042bbd7c361d30f5358065949180bb5f4cfde97e7d061fc24b5e40e116846a62a9ad763eaee
z109aea26821b35dbab3ef4a352bfb38484e2a6b5235f0a02aabf855c3962f314e7889761fe8f28
zb338c9e781398609f2aa9dc1257943669ac29a8b41719b878aaae9eb72d4a3977348f8a575f80a
zb20fd02e3ff2ff489b3c45b606baa36c811f08b845bfd7171e0cd3c71f8020bc3aa527764ea3ac
z9a611dcc3b093e66277440d0e151c38231ca0cbb3dc8b431a933292021a76c3ac5b83df2526b6b
z02c0136bb2910fc3db03ec35ad01a1753dc8ea0dd6f6f6122089b1b7a36c9be71108dffef6f0d0
z927a08fd537fdfbf25c877004ef10c612e7d6258eedbed3837d09b9e473fcd6ea45bf75f495575
z76e2df94070e21bd1619174ad08c080a45c8641c2ee1b7284c1b78270b2db97cdb360c30dffcb2
z011fc8d59b12d995e1335ad2515294d78271a196a2db1d551f0d9d4b1af625002898726df23fe6
zcd17b306f1ed43584daf93fcbe759a06b151239faf52a007a86dad445630033961c82e4f27bfb6
z3133367ec53d017a3590916aa6487dd31673c6af328c61c4ee624a15d332c3a864588c093f954d
z9ba3dac32a27e309ccfb302fe8e368d8b230a250c96036ea1efdb077aa71f8647a8381be250fbf
zd35b44da7bfe70aab2301f0420f92027563ebab270a56926d0cc740f0ced0b1d33fc84fc4242c1
z74054d8144f3c9065e6646800d3263e72cdc0be243ea70128880fa7093d45c648afdbd81558138
z0e5a0865ff4a3121773f2905e973082d85632191642bf1f1b63eb666590d6e34816f8178280345
z31c1a39d44e37ce9c6abd2f3299e148e3dfe543248dd4135eb89b01565a28ec15eb5fa43aebfdf
z45fefcc4d2d3d4be71df11c919f0c77f006dfe07ee9123687c1f426994d7c389737196510cbc9c
z511543f1e181c699913fde89c5a6ff83fb9fa94d1b3550d031ee8cd59e9a6e8986f28e02b208e0
z5e4286809ee0f29f649f8ad7c13c7e11d3369d2c0737b872172f3be62e40a44420cb6572c169f9
zbd02fc5c71e5f1d77b31e5f33ad6203cc979d59889bb6ca1ab4f0dde57e78b5918614257c40da9
z501011e78e42c4a0755369b666d55a53f482a86b698306fea5ebf4cf60122ca1974f4128c015b2
zeca8ad6d133712e845da8c40d83d594bed935b8ce1ec2ade9629557f3e58889094f5c6c3ef2cab
zda5961c4c09ce9302ae7bf3886fcba898dee3ecbc50bd5b61dddef0f4561c4d7bb05167d2e5ab1
za9e503e36dc08bdad21330d5d5641721a9d0b35f1c1aad0aa55a0f0ebe5d8951490696b2b48d84
zd67c54f8c3d344cab8c800f838726467a5930d85f7fdb61542975c469d214d33e996c887069e34
zd0047c7f91df7922ef3425153942f2c0cf0fde9a87ecee046035e68aa17231758f0c94e3153178
zf91f859dee65466b8faecee604eff533fda1f8dacb1a6b7f532bdae9b7828750b9161c2f122a1b
z4ada39271f4b6a45cb0303cefdd26ad3af1df845267379d2143a04c3ab9f338dd2aaa25f0f66c0
zf88d201becbeaff2422c88bd5f781811b15200698c28e7fd03fc25ebf5d9a3f532ea7dcbc4ce1e
zb1faf0b7e79abae68fbec5f77061994a73bb3da024ad6afa4662ff03184e48bc2f69cfecbf4eb0
zb5031ba12c36440be91a6c597a663992b7cedc9eb01a0d1998ac6b585c9ab9f6fa8da8ba894abc
zf0004f8503ebb0a3683acc38f6454f88b19bf327328fdcb1d8a2072e4677e77059f0d40ee514ae
z43dc98cf748a335689df5d24bc013e8770fd847e7d3551cf521bdaa3725ede7b50c48303b86cc3
zb33e583fd6f7b4385ff852e1bf38c11b4551a75588198a2057596bf1b26426349c824342533e1c
z8cef4c07a38ba8dbd69153d6f4f23363ee6c5cff16d20dddc6dd4c2536f3154cb1740e19a213b4
z67e3ee967faba5841771930a732fc8b1040bf68f498c656439575b0504eb3e156a51d03ee1dd6d
z258933f9428b45d3946798ed7c024d7adbfb4177d6d49cfe01c90098c31134c83c76bb95b3b299
z8d1dfea4b14cc261c625279fb6554a956257f23e4174c75d873465b5a5425010ed01f0b7f17177
ze97c8b0ca7e61e22cd976e05cab47f25e85167b0489937bb0eb79772296a3bd0f28a081fd92457
z9fe14b8c16e524af8cbc6cbe616e5250fe3160102a6cb779a8b3d9e5d701c67b85bca61297fffa
ze71f963e29309e54310ad7ad761dcce0c8104a25461d71d68547432cb5f7af3b32c3affa607cb0
z0303df9048a9e96cbda6ba08089841830b8aebb944d694964cd5a04cb63cb279c9627c836ae575
z5e0ddb26de363e65ef5145ff55671d4ca407c82a9646bab12a812c4c896eb93c371a6f0cb36e77
z206f307d9dcbcac7b13b6858b32853caba9b81dc3cd020c6afe058ecb16e21be6fa6f95ffd2c60
z309745418542a57dff55b7ff7f2e750f433f856d031ceea7de9c683873cdb44db8ce10feb57c7a
z695027f08c58629ad3dfd87db208b3ec73e55529055ebf8da083cb86c6e1af9b638a5adb81bdeb
z688bdebaccb79cebfdf967a1b1d7bba40fba7ff7948ae434b4f55650c2ab6c8604126582a82b0f
z91f58d2d43afe6ff018cc705d116bb3825b6fb53fd7f241779b80c4db6344f0e8605a857c33bd3
z7f308be7c270bfc1b20a9e90c36f6570c5f03f7401dba77346e0bf40bb7e4c2efe8eee8570eefa
zf41eb850db99b5d0653e290cd8f57773d18a7bae63415b4457a63f70c83bfd6a6481d94b85d8ce
z8fdf932e6bac56b81942730639f9d0f830558305f2249f0f9cec38db09f74d705e6de3d21803ab
z6dec6fcc2d554f283955edf64ca822f0e2c8c845aa2058e415594e8dcd9a1c7c773cd52cad4d60
z3b438ccd62871cdf01410777e13394ac92fb9733f0d540355ca884c1e7c84afaee89a31516d90c
z39be1c9d9816a0780634175b1d7d7dd01545dcbf0e18a22ea8ec12269c26c235de40494db271c0
ze92cd32ee0ed46285306249f5367e72bb5fcb3a51c641787c484168f1de1805d039ab505c844bf
z4e5e2f5aed4eabc5851bdcd7eb83e950d3efbc5a3513bc6ded78dabb80ebb8c0956d213a56407d
z370fdcff78446df27abc7d2ce12b16a6a0d7f7c0fc0108e36f362cf2237f9a89b70a50594e1804
ze5872915fcfd2e20c93850dee95ab279af39dbc69da1d428fc6bcda6dd974dfad52bc4b8496d81
zc7342de7df125fd184fd646bd8127a2cd9a4060695069e22bd82817f2ebfd9d10c24f74d10fe0a
z43cb596064be939d3984cfc7be5f8e310dc3e3d02c2eac1c8d5bd1ad35642affb82f83861c698c
z128fb6e1409ae398500b8a8a67f37472b93d0026541e997d3a29dbd719a76aeffdd3144827fcf9
z21258cd9cd72cd12b093e56898dd3f3afce430190f90320f17a0ccb591a817238f2fb32b8e8d6f
z22e0a8e2d383e4fc184d806d209e5b40a1de4cab9a80913d9a3157ce0b7273274444b80a2fab76
z7b25f69a5157bd5330637fb92f8ce6ff9e5e2c665e12d689c0699a4296f598fa4521cf76d7f13b
z58ac118c3eb4f6a381035344c0ec6323de8da5e615a6e2debe4de44206e5afe50dbee7ae1e0062
z08d0547de3fa4a0e6045433215971f71ea9cd6da04fcbcd9a1bef3fa3d6fc630f25437682a1a6a
z4024b40934108028dceb9b8563ebbf15a42a2b2caa82634586fb964ea9edcda2ab9a2821488d00
z12d26d89a0f3b4ae9aa61ec97a60d67f72c25e419c363a54655002923fbbcd19ad725d2173c40f
zb01ad6fae618d0c92c91e68da06af6309c5131e86e3f02e4c5d29ef938f59f7fb2c19a9a2a6633
z1fe19ada39ef3f688d40bdef71fbcc1b6787097324be5ac9474c7c86a436c004343120b19eb8c7
z0bd5afcc41cd3f3997aafc5772527f5a308378e6635ff44396b269dab0e6e0d6d2821f666ff18f
z649a19bbe4a53518db9ee7119786971f07974026211c892c43abe345e44980989c5936ca6f3d04
z081bf01b36e183194e436661b43fae1fda166b4a531493703e6f0cbb6f68e45b603077cd7ca8f7
ze683e313a14efafaa95a33b8d5678f72bcc4f4e8d7b328f5473dc9c92ea123642cdd5ed041245e
z925eb8bb20050a3e2842109e66d3cb72581e4a87e369c5026c515701d3f5c67084f4e7a3971820
z8c19a838eb7a4c3b3e49f275e603007398384247f85597483ba7e1363e3ecec6c53633cdf98317
z415dee8f38abd9ee52300a3c7d85cada32420ea95589b7190476b1b7abd4de4fd00db67223d999
zd6e4b28afbab414f5ebd50c9ca7649c6fe7c745486007092bff1cd2ca271d0a0453646df6fa77e
ze5ae248e54dab077abcda38a72eeef6a3e3f0db7136583459ce51df3eb437f8c49e9d3b4b03996
zab6faec775cb287b699c8ea9d661ca0d872b52a3e8dd3218bfdae5f171c1879e30b078dd20db8b
z83b1f4957089a96d427c3b7634c697dd92a711f289a88d77ade09b3ab1b852469106fafb9d6c65
z4c1d872b109669743410852af62284ef8806eef8fb3de953c58285c0361c13c068526f455a622a
z35e4e91ac08f9447e311421ed91562204c0bced43e91cb6ffd20dd84028b708523f3f8b22be1eb
z59ab5b6adbf0646a4cc1a3e4d20aae212dfc59e756b6f9b3836f4165c1ddf297c10516c94a2981
z4f98d8d281c69b4dda7622c6f4dca7482e517694c5df85c53f54605ba4fc12b264025ff79a2e6b
z6d808dd1069d6dcf85cc22b3a5d18a4650576605eb42a47395ca6e77222c1982e27aca6fac1640
zbacd4a2b0db88c6e27baa59d74c8c3576323b6b4c6e54001d8ce7fb1864ad77454ca2e78e625eb
z4aa5006dcb82a3b27cbb768b321919d463d75a93afeeb47cbbc8e30ca3e0e75a76ee2eee891a60
zc8112eadc29ca146f83faee09f0ade06bb9eeb8f79bd4e6c2aa31bc8ff838c8192a405aa229461
z07b13d2561f15ed31c8ed5dd89b1d7aa8074f0ade287e14e591b87858b29258a5748d6a0957f20
zbce769d586347a82e84c517ce595b5e60bef905a137610189c55bdf0d47a804e2505b6ad295ebd
z853b34bf4f23afe5e189b563ead38f88e358a1fb69b6027fed122b3f6c8f3a6c6ff46baf7c5412
z94f2c7e0a0d2882cc5794535dbb11cb6185b4ad2d11f1564874009855bf9020331f67a3940dfea
z5d90298d5ec1825e9a6381e8a001bd8c658b31912f2da7c7046ea554ff0904bb36054f39726cf4
z322e4d403da9b73c0006830ebfa80900ed3d8a82f2e019d49d3d301df8f54686776bba42775d8f
z513ba9572213b41a25262a56d991d274d78642dd6c4ebc9050052e07da75aea131b01b3ff3cedb
z28dc5a195733b10514410ebc4be838085bc86d72395c47a5027f5e3a3bd5e31aec174867b12c44
zd8b3598f10fde6b6386b52830ac975810179b53bfbe060a6cdf6ba5437fde8ba31cdde21a8d16e
za4e4a233b721e00f2c0d0d91530a088f79afc75f6d75d5593fa770743bc0ae81bae38a8aabdbf2
zafec34045157a460684e2b262ad9dafb0ddabf48ada9c9000fd71eda8883b8143683ff899cfb63
zd58e7997e789f1ce505de8fa66142f0f73604a395501fed409113519ab2ef6513c094438a1fa3c
z9e2b287611142fb5e9dc5d9daa394ebc5db51d69f53dd1bfc7169d249c9eb9cb71537e52ec9ea0
zea088b39d31675c9835ddececf51110788f90753ce32b0a5dbd4aa1a4160296921ecc22c050365
zdbf0002b990dbc255eabbcae078297e717f37da03bdeecba2a85a0b16ce0b3a2c80e8ee8ecea1b
zcbec9e772b3221f834f66cf15c778444897f477f5baf4b35488a522ebc63eca167302d92f64049
za1cc75040d782d561f33bfbfb98ad5677e259c3a09c88b89455678a4aa8b557f743990b1e697c0
z93faefce79507d763248231b0bcfed100642a17583cd4c4af40bc1973408d89dc6e79ea582531b
z276587c0e1f5f6c04150d594bf3c0c369c4bfc54baf26582199961437f7c7fd01bce159af27482
z28034a2495e1b200e725d4026682aef7ca107a097e22cedd115d867bfe16f72a0df7fa2b9ac813
z4b3ce06bba2a7e0cbd1524d78f2cebf91a86cff328df173ad6720eeebc07b816e13207a0beafab
z7c605f99e69a57349316156dbe3edce1a155116b3f493416dbf502e6c71de7041043016d92429a
zae0f2ab8059927a79bbb028718cecd97001a1a7049fb1dc783c9bd151cab178e8bbce4562b612e
z79f5dd78f69046add59db4aeb01e4f289aa4e542f55dfbb6a402d22f7941c69084ba7bf64363ae
z6b2501d2afe1333397974af3c7d933adf1acfe00a45bddc05870cfbb9398ebf1ee9c5b07eb6272
z353d75656dc0764bf5aaf65b1addef342ed1bc67a91565034f42e4e5bee7453980af3665e7ae48
zdce63d76545ea7e15e72ca37a60eb3b92a47f4eeab309e2dc61a0e58df1a7286744501a2c02f5d
za70ff1c793059d1319380b0ea91c80cea7e326976b6d8069c2d23a963c251a3f8e1ae3cab05869
ze5438e9f11745df314509afe7fef90726a30a485204c0bab8eefbf817d1f75c0f695164321a0bf
zedcaef9ab221ed430651812a2a1a33a6a5984b562b5caf9acb22b8b38576fcba8de9d6e4b6e7cf
z0f72069e1bc85425c69c344e0e77a459941695d929da5c7eab833dddecd2104d6bd6add1616443
zc35d56611028ceb83704986094919ac90d04141124e6c6219686296218fd8f2467acc16d9186e8
z4295eeb4b81f1a8baca9e6bfb8c64f4318cd06d8852ffe7e8f0247b99b63b00efc1faf17011cd2
z3611a33ab12e7a91c3651039c8c1311b394d734d636b147cfffdfd1f755613be62f10cd4d8880c
za5311f35f097680fe37287e1cd41db422e1ba2e2dacdff8731931783580d22926214501db068ca
zcf8e7f260eff2d2c51405c0f88e07da3929bef9d7efd53d6f877663e2f662ebdf3aed09e4de8f4
z7f5dd4bc076e79ffb47e7a4d5dce276b7ba8783d61cef22e6ad6577041453e9e5591fc3be02c12
z0b7fefa2445181761d6b3f33add6f7d6174a32773fd9ce31b3deb84971656cb9e4b08c9d3ec134
z06cca1febdc41d09b8c553bdb47b145fd7ddd92a77c058ac56c5d476c10f485585bb5f63888422
z62ed0b3a460c0354f4a666b9d37e8770920fd057b6bd6b2d97e29f0a3585bf5c595d5a1410a4df
z51612b5564a67024e5d30ff6e9ac37c9143ddd45aafd87047d40766e294faa98452d18dff16b39
ze5a32201597e6fd5ea47d6cb5c4651db6c9e5717241aa461204e1dcdabcd5fe127d196a810c3d8
z81642d6957e81d0f1ff34d376c21624827cb99ff37e6b57428698c127a9b7b7679fba27cd7537c
zfe25afd499447434c7d3154d7b0510ccdc7f418e86dd792c01d03cf34b66a967ddb653fab33478
z66b488ccacd8e6ae39eda797d943039092020d9bfa090fcd7b52fc4d4061086549b5e05e080f47
ze3e2b7f47224fdebbe9a69bc0b1b333f3d5536371a08329aac0c54960afe659353d613ff3ce6f3
z2cf73168122adcf0de01ee8da8cfd09fcc802848330db314d722569d22728b595823e9971e8163
z22bffcd4469432765effbae57059c6630716fa3654c94bd271c71a215414095c9860dd72df1033
z9a7df48d7ca94ec507f90209d3bfc7a328d2fd2e1a73b91c90092d04f27bb62965cce0c046a883
z5f73d4a1951347b81b2cf8a02f812d527100bbe6f9233db258743ecbbdf0e47778f77ee1612edd
zf2a349f045d6b894c9856bf69ba76ad2f1651dc21df56e7375907070aaeabf4a93c8c835320eb0
z3cd16ba61d01bc0bafbb58abe80a345226dda3cd3ed90dadb0f39fa4dddbac2e3444754d462c31
z2e6f11706a3fc5021cc03488f777f42c56308986ae1e6b3bed97312284842b2a14a66dc6244d19
zcafff7732d557896443f3714e0315b33f294dda96dffee4aeb204ac1c4249d043da9729620e3f0
z5f5cb90fd336d0a45d15446572bd2b3c801d2e75a9b813a014abbb21d0c487b3c8bad710a4cc9b
z75c8e05913f28b648b345808246fb7a18bbc88476b5b586fb137190e431df3c3e4ae308d140ef7
z59f68d44de30fac4b675727eebd2dbf869fd9479cd795827600dac9e1b1f0b9aa03af4bb2b03b0
zed364808585de9f6a754be3a541318542b17cb6ff6b8b68bd5625b4d78aecaa9b12cc385ab6b91
z6c9e1c7ee04680165771dd7d5d84c1690dc11393cc6814c76194f95d03e1ab4268840431787dc2
ze32bd4c7c524a6875544762b905d3e54e855796a14886ab0bf1951f9311fa58ff19ad8b98f8727
z5f03543ff54f43e2eaf08a46a911da1a66f4b2ba49a2c29b428a6ee9daba3fe8cc127494b817a9
zf70c51575a7d11edde12156dcb1a848b8fd392f1fa03202e559846c79c18664b9ff6665341fc12
zc0a1e48a3addc2a1456a08e0ce3aeb42d07f1cadde6f2c8e0016d68f4eba227b47ebe51835200d
z1964c39561ca14dc103f829ca2af5b27fd82c1e4217c032318f93846da4a28ca8771dfa5731f7e
zb10b25d868e08ea2b7108bfaeca5e86d537598dd0994c49f5448cecfce6c04bbc2bdade23fc480
z82904842e20b2349b5d32511c583e65926338c720d6443901bd0d755a3d7d7685c882a4b67b8e0
z5811f686af3771ffcf0d54712e69c7b4a69705bd8b33db3d3a552b0fc0004d0818a576cf961bb1
za33123c118859f1e69636e987fc3b0c2ae2e42859027b00580fbc2e1a46be94fefd9eaff1b86ef
zc8bf876dd5ce5053f6cac94e9724481a7521776ae35cc5511e6822684b28cd01c6382a6f58f81f
z35479d2f983bcb24562ec1d2ceff9055e5345455b0a18352a1c21928f959c9c91360bc00972368
z2f6f564d8acbdff53132637649023782c3c98b19101ef1bcc19e21782f9010942c1fdb0d36cfc4
z72380281e77dedbc93739fc5cd849d12357437aec938caf1ec1d0a07c82688c854b410aa7d863d
z5ed3c0547f135a0171bb7deb121279a3a29120cb3b6171fd77b79b004821d47001e158c65c58b2
z89f3da62a2fe12ee5ed7b3421b2e34482629112e544eb9002a7ae88d938e9b6a8edcc4c41e0432
za86e350088c734a219d001910ecc4aef57bdae6041dcfe86b51b815400f54e6a656dfb7bda9a65
z8d1b2004ab062787657412e5423f97e798b286468c3eff09d6a5df48f706ef918e0b4ff7abd011
zd1dbe59517312e5ef7bba8070fe5e1b85006d0b0646e7cdc22c5b2b7a6c971b3396701a9947997
z2865a94a12faa71e2496d05d30f02b054f303599215fa9d6e97fac76ed4af9900905ccac85e30e
ze779e965e23d8e76de442f0a8d0e520a5ff249a6bf939d144e72e25ebd53e98cbe221bdf4a4186
z524ac60a2d919139629f8076221cd92a9f74daecb498bd704234dd6d79f50754bfe7f7b8c1e0a3
zd925f3955afd834d7ea994eed7a5c23d113880c360c1168841385f53dcbfc0dc00c6cbcd99a80c
zf038114d030e10fcba236910e54181e45d54df0b3f03b25ce2a03330472ac134d4db92a3c69a8d
zd158b6f21afd46350f54c1835d5dca2245233f776b3b71c957ffd1556a35d80286ed300b478d18
z9b0a98e03a3dc156f39479ecd05efa607179aa7a5effcb3d61b4ca19b3a8cfaf7286c3392a8761
zc22860a8d3077a9a66c4d6c1448b172a36c6ad1f8d82fa90659ab02e93a72175f5164d9dc5c72c
zb26e8dafe9c37fe2788480fe4f1125008f9e94acb6d05e74eeff21ca07b4a8281b66911aed5ff7
z1f5f38a54a0a4d432e007ddf17ad4a5682b9073d4971311c6f7167392bbcb6770ba6457bad5ff6
z1a358c4fc5123ed9d4b2e720194799c08f1590195e4f9fae58df821cbdb408fe80b5ab4bd0559d
z00f4181a7cc6a98014c6dd7f80a294c8c940bc379d32b5e990ab390d1c9cd07e63df329437662a
z30f57d4d996256415c8fe68352f485156608085488e286ccb3ded60816f653dc7d6d630209fee7
z397e2b522de761447ae8cdd2d81d191cdd1376aeeaf504460be000750703547c95c78aa5e8ab53
z6bd5cb8f1d84c2989d51184f3082b1e4c67581b04d6e57fd2eb346826a745a98d6723af24aaf14
z2087558dbeac577bf9d8015b07a6e530bd6de3bdae53696cf4cc7e3eae0c4768346726798feee0
z537890abf6bed759e18b26546366d8a1616f152a89ae4506b31580c2b2e7418d59ecde49f0eda5
zd687adf0a68d8c116f994d1ea5bdc5a942d7467daad893a7c02a9e0888625d90a525946e64ca71
z5738dcfc80104fb8b4cf2d819412a097dace063d9a380e69b4bbcb38a48c6dbbf3469250ba631b
z191bb2cb496f6660dceebee327523c1e7c831092e7935abd3ea8fb6e81f4f49d3f821ce79348a8
z3daec96af1c073340c3d65241ab2a2db62380d2e274ab2745cac4b26f61a1721102fa615d93ecb
zbdd7ba91313135e89b4b8347b4a4045d2d94a88db85993a04f5511c6f961d9025b576418373452
z649f480e21fe8cb78a53755bf6fef1f78b0ce103d9fed651cad3a11f9f24dfdea1280075c6b010
za174476c23d4970078d4d33923df8bdecec9275213208b0c1ec7833c4a52109b66761b4648cb47
z3ae856d6b2ded47aad2bada8f34f4f9ee9eee91c07ee1b92ac6be0addd224a09f35e2cc11520f3
zd0cef2ac02f434d591d4350b0b552d3a3c4035cebe28021b96a4005a53ba8dd150e8e2af3bfc64
z21e67e342326b6639e3ea2ea8f045d05f426661cfa63cb555f89d1a8ce72e8ca44625e1a9af37a
z7fb131ffd303357996190475a5a0936fef3bea15a2a597f456ca59bb4da57765378d8afac8ab24
zc0dbfee66147afa71566de3651c97a0db67e09db42f0c800b1731cbc206441626def437566d718
z685c9792d822f9523dc0fc70505aec279a6fd208437376127b97d0488df81b914b2d6743660f21
zb872aeefbdc8b0e4d446b6eff80edc719c3d544e7b051b8079c726bedeb2bdd4d103b0270812e7
zc278c6c0a2f79b1f24f65d0cba61e4c1057adac51890054f8be04374e851e2c2d4e8566d1a300d
z0bdabbf7b162dcf52e1c33af1d8bd6d7c657a87124c161649e1890eb82e9f170c5e9951e8e4a99
z4e52c98c8b60ac9ca075ae79143c6327ac9be682e2dfdc124e5c26c92aa46718e12af556257b9c
z9a9f1bf4e9a7dacfb8270af956b8fec36da59f1ff6a24360029605e938f7c2c818853c6f051815
zcd495bcf4c0d430d7695c4c22201e18712fcab70d3b0dad135ae51fd25f8e230b1ba7d41b32dd6
z370fba8a5aecb4ac3cb1dbd83c58f31d69a91b44c9b5d050302f1fc8f16c174607173a7875936f
zc29c302ca03e70a17802cf362f5ecd1aa1070b755f2a78c199897bda3c629616b669b7cb73e33b
zc852d26c4d17ebfc87274108576ae85a7cce8ecc241195dd53d25e570f69bb7376d8a13c86a7ef
z83d6d0f51d12e90fbe70fa4bddcc452b38d32d5fb919dfce423b4c97b988c4662367c5885a9422
z52c58431764b97f96bf95632aa8a63d910e89c68f6f1fbf3290b5c536f7c76b43d2c43f7ffb846
zceab877eca82cf65d5a846f3e37c5bb4b1518ff7684e1e2d41814cd8142a3cd5237df2a6746cc4
ze4f8f50cc09941a2ef2ca540f4e34ab2e382017f69a8db75821f65ca11be338de78d9aac39de46
zfa630edef9d11c6c8d16844c066fa4b0dbfd4697a84f18829b5c8df8cddc5eecd40e96ea11c033
zb75a86c4d3af91eee66bc43a7dfacf0795f0515168fba33af927f545153bd19ad4396b472a7280
z12b2115f838ca4da0c1fc579b1a5c702d9e69b3eaf28148a7ef40dfdb91300a7b319ad2d77806d
z23e545e461f8309faef4199ee03231b867c595237dc27b7810f1f0e88970a24f9caf84c13ed3e2
z4391be3d7b9f9efd0c0db83a57c2e101bf33761d9f7a7881ec2d45e260772244975300c28bd44e
z00ca813e62ec8cf490b9d8e57ed9ab34adb18ab7def69c37df9188d6d5e767bc78c21d198690eb
z2f9d70465137e2fe9adc734daf8f95426e9baf922d1db013134abeca5800d9655f151870785d50
zeb6d04e21590922841ac03a73b74f3eaf5eca55aaeb3315028ca3761d827e86d65d67776aebafb
z87ba1fc230f684f94fa4a9e68feb5d81731afa4e605992d57e4332ced139931b178b228893015e
z337252cd9b055fe6ffb63134bad4f1e59790bdedd5779d53487f6d3f3fe6dc91c468fa970a325e
z97f411f75852ae1845e49c65b2669939eee0efebba8696365015bc128817ce09f229bcf52d69b0
z508b6bbc1bcd7f48bfe66712cf27b0037c8f415c87f913102772132b63732e103e1a7ab04f7c8f
zd2875801dd8347fd8768b7039d742568b70429842150c17b0667a25dc046a52a9aa9991f56a0e9
za80bff70686cf9e24937b1807435269ea167d037c839281c5808ee4e5c98e17777717b6eae6110
zef7b01129b7ca8eebf0824e2ca476efb9ba623e5f5b64deda94906e691a07e6a265f279a61ae1f
z7c16fa970e15a33b1db4206e6b3c34febcdd0f786c9d1a3682f4f11a31993d3ae5f2ce6b0317db
z1c51a3b11735f086abf5f69c0e9dbe7a3ffa5ce7d842f7fdebb4b7a09fbc39cc4c302c442de667
z961fa53b7885b4d91dd28668823654c07a6e1e460754f54fdb8d854d07f8c422cf726614ef166b
z6d3eb3db84ae3c351735e855c177f6f54054e9c32a1a54ea6e4baf40a96e9a598e72d259629d1d
zb6a5824e60b4fc83c9a4002e35f2239c20c9188b42c23567ab60706a697435c5516024cbc55196
ze8f4c9836fc100e315380bc0bcf56c554f079f1745e2c2c1d54993d0b5f960749e25ba880084a9
z440f646eac01eb6d9e2a87c79f58ddfa7218aeaad9b4e89006ded16c5b52ba8da3d74fe9cef7db
zb3ead271d6925d30880f0c2b203fa68e4d16debffccb58461182b39f586e06fcc606dc3911ddc1
z4a246344ca8b77198979da8a32b9d13cc714d29da81359b1a12196a4ae4777aac702ddef284f93
z69fa73ceb45aa5026f967ee7a338b51615a880309ca7922b07bf8493793492065edb9e9bd4514e
z53e6b4bf5a1b5f7550ada6c06ec2e6109ef8b3962a1ecca0f7fe097ca7841fd8d4c0626e584bcc
zfd8b69ffd5f7fb56939fb51f48938ddbc47abc2d669743fad1832b45e71512f941889f10d2f044
z192167724819c3ce3862a5cecf67f3cdc5adbaf578e60b42299899886c3d2f8f7ed4083b0480d8
z278536257a14ee4cec27389c37340e6ca5b8293eae499e1559269525010c7aa9be090c80eee931
zb27109cab54806503fd6c0ca2886e0b1864456d33f07b953c7845d9e95ea138103e7fd0995e9d5
z31a62005d321541411aa6142985a1d07adf704b56ab6cfcae35eb1c182323df7d7f60cd360b9ac
z645906374ba7832faaf1d9d686600cf5b034e1e041f2b3254561e7c5e095bb09fa717e80e44852
z4a850da2e3e363b93b8d70feb795d9ad01576fb57c47b67574309146d605583a75854d51225e55
z72329ace2ccae222b6a2c050343fb52035d8b67044bfd3268618e89f76eddd31c4d836e6ac0817
z3777784b95b517d2cb2443d65d4b9337a516010337a349ea8a43a5fa7bebbb49dea7f020bf3436
za06a196eeff0cba9d831131b04bd112006bd2de76fe5445808ffc16ce5d2a4f293c95cd0193c09
ze14ad5397f63485f2b0f4fd61c115d31f661d6855fae5e4159f5da2be0ce168fa9d1a27177051c
z3450bfb829b19fefd7eff61ad5700304c501dfb93e225afeb4b929a50afa4b06d0f2ec708daa47
z574255d7dd8288d2e96dd8393febc52e66a4370d8dcf18f67572ea9f77846d8988542327980e10
zf7f8114437fe64ce05174d28fe21a10bfa66a340523564eaa5080b88745e2c6e47049d400a441f
z24bc3321dd709d1571d387eb7567855d9b4e34654cbeaf8b838abb0417beef19d7a507d3c17208
z824ac7002bfe249ea6c859e7772c28fed3d9c3efa22aae03d6525e8b76d368a33bb2ee65f9801c
z7bf6ecef5f02573ea90a799c5ab428f17d43d51364c73ec5fe255f128a966fa223fcb6c7d350ae
zcc4c183d55f3c5149d73812c89084321e4807737263902d5a64a244ff6b5a3ee739cb527545802
zd30ceb1d98a4c2892d4b560ff79e5e13c6d7e2047bb00b8beeefd2357fb19cea476ce37b6c0482
z1b1eb1bac46cfc3e603139f16359a51804de945e2abea2f27e92a7161f1e47698022527eb2d6fe
z3d4426b4a5b6da1deab452ca0ef1fbda77c67de39a10067a8b56bc6ded89861533a48f29514c22
z55a85d619cd909743d274799828abe421d22a873de472220007a55fb12e3373181b084ec30cd13
z8e2bb4bc70f4f68792aeb83a894294daa042d06d75a995fc69cf5b2a5d8e3d6520c2f5035692af
z41fcfc2556eea69592e2e15ecfc766f9b9905436ac19d3a9506372830b87897adef2e1fa170d22
zf184c15989e04f596733b22ec8a5ce409dfd24035ad449b99ca785e5d87a89df0bcd226fbdb38b
z859cc345aa4b7a491c593f13afed3e4d42d25d020a181f12b3d003c711b4575139cfa8b20cc925
zf881ba684ff971f8afcd001f8ef74005d844f7b4c35e571719d100f6f4b42d057904eebc3a8cf1
z26d82f2cad9cf9de15fbd42470ee5b5d288fda2ab938347d1a60713dc39d34ed94360ec06e2f20
z82698b848321ceae0c89bcde66a9cf72449c338e366efc06a4dd748117b28a705b9055f4db0ae4
z29504a2f5cc2991fa0abd91ec955c03d4867b1f83f7ac2566d32072c35f0dc645a2dcfc7ca9c0f
z9ed311a28f8a98fc0fc67d8807660a8f1032082b05508e6ea6c763535386948c0368b6b6490a21
ze78037166d8aba8f695e077887d88b6a84ccbd854a2bc83a55d9f01f22f7441ede5287ecdcd46d
z4db3a6ac18216f43f42b48beca0f8e10cae6c012c7669dcd4430accb68c05365e44fa997443c8f
zc7880ffeb63f62eaa4dd6dc18d5de8966b5c2d354aeb2a0c89903e5b49245c06544d7ee8243a4c
zafca92243829bc1ee481cdf23688c0ff22e88f3650bce73449fb06a99dcd92210903e0d70431e2
zf34c58371b76c6d9fbe9ca2517c585dfdf24a9f378d76071a196b2bdb9f68c8193e035d0af673f
z8400d218097ede6dec98226cba8e125630e6b932333391b5fd00114594b0e50c567c18095e7782
z926397ec32b0cd768ee89eeb2289f0af6bc61200bc92b84591579bb085fa559e94a4b738e3ab40
zfd2c257295aac0b6e00f61aa681dc343d6fb55814d85c17b146dbdeb551a5c2f7edb9344514e5d
zc1e78a4fa5bcc1b6fbd5fd2e514625475b8b46b3e0cc716628c25f7d3686320f9b3f8ca271786c
za4abf51ca14a992bd1bc9e5ea328b64885abdefc9c382c974a2b880441cee9dd1b0d2ba40e5791
z7833a0e1538fff58cdab6e01f981f1f395182aaa2be667676a1bfbc223494ff867b7bdfa95aab5
z71e89ca32df91f62a819438b690ce6a1ee6aadd5beabf7807ad9234cf7232debeb6b2234b67d7c
z9007ea19674e1f9dceb5a8faace8d85b35c90b6edab857f375bf3e074fba981309dcc6e96c6586
zac1a76944e9757e931d6bd0aa3c1f4f18cec5a59bdaed72fc29f02bb417ccdfd756f5af941184b
z650f6f6f6bbea5f84a0d11a02eded5584c63d80c07adc503e0589ff0410c5beed4c47492ad1ea1
zc182f96b224b518474b153bec4f5b33a093d6f9c08cf2256e30cee67a462571789b3616f245198
zc81913447e2babce63c3ff604e1fb0decf76a2f6d157d7a3018e64fdb48618fc37905647cc390d
z7b98aeb7530250bb58aa5af811dcec8a0b0d2c5c44a77608dc1e9e6c290194b00590a1b79a94c9
z4e1c893339709899656222790a26402af5c2a4d8250225677be022d5c4938dc7f8e968b7fb7e12
z34205d001e61d1f124b88eb813e653b39220eaf3bd2eae5058ee65cc64883809526c7fb0ccfe56
zb52c744329d5c945508d764b42972bc4ed2fe768471a8e41a59ec745704540084c3f3abd4dda16
z8b889ea0efedae6fe8ed9d888b04c8f72118813592ca8093b9b4f76b686eff1c5f405e86dc62d0
z528caa0a5ccbbf064159b0d352b08af38e7a21c9bfb58ef09b18d8a3ec5be1593a33d21e8fa9e4
z6befc66904767bbf0d3fba6d6842fa1208271e5e5f52cd028642e333f06b97428eb918b34fa6e4
zde451b68ad469925353344fc2f10df340bd248eb9b8e67deab857035aa4a8159fa088a344e4719
zb06a4734749db34a53f12cc6af3ef9300444584f4d8e166c592921773c8685c66512440eec7191
z13fa1b97aec25eec85d2241d9e5f16d65c031f738aaf4c31fb5542d948f90122909df97c033303
z3935a062564529d0d98541f25256e3f28cae2358cd5b962a4f6d481df5b9420ea031fc236945f9
z815289291cccfa26099cca6cf3fabcba802897638b297aa59099be644eb6448d76475d2520ad5b
zefab0febc08b555e14950faf80145bb71edfa2fac6bb27d67d02c43e9c622b5c64d9d577f91135
z119e8ebcfd05d0ad65fc12c14338f8dac5e14bcc12c380e698411419562c4dd4fdee2c4e5a3274
zdc65c5c5dce87f423beb26273b8443e7d6652a77fceec3c2fb44c1f7c5997f3614fd2c8fd2da41
z6f8a44dbe0bb7b62cc2bbd7fc166336a7f1c20b4cf7b0d8f225a47e9256d9d58654ace2abd3f4e
zc784fd6aa76108c139f559f4563ac23e22a4baec33fca72cd0f68e4585ad96bd1292581ecd27e5
z774711feea03660c293a73d9c52b6888e1746923231025d6b4e298b6b4dd8cf49f269a94e21051
z62b73ec549f77c608f7e3d9a55f3fcbc8f912c23a35aa63447c58ed6255142a7210e2ac93baeb7
z9af6895f07ca21939b6c709db236fd60cc26290a5f670d7a30d53106951480c3a1b25565e82ff4
zf5224832eef1164003b921fa11fa1ce41e351755aef55a8b9e5ea63c462b2de63a7f66b0c327cd
zb339b5261a820f9634554905db5291f2aa62b33526795b0e9379019a160b7eabbd728ac3889729
zd22e48d33f2bc06bbe92e4ceecaae53849c68abb7bd7e12eb984031842cf9f8a7b2b2daa30affc
z0ad5399f3e801e202bad74f3b4d624da2b1200febb505295dcf48acc9dd2361996c2b2275d7198
z5980515d28d18802305141847a6e961c56117927578fe910a4b0ef30db336ec2a9675b1ba4e237
ze2fedc78fc7fb0640e86dd9ad2c50663029ee77a1aae85008792782635d60cf73500f1ad7bbec4
z5b3d80739817c93c03c607c87093b575360b6f2b16b18739d31632940256293e31bf94c89c796c
z9b14714ab84cd1623dd88e3e68703cb2ebf94f394b306f68e128d17aec99743ef7d636f25fb08c
zcf21e61d063d8deb7dbf780de97fae103ed68476c8b8efb0bab7c1ef09d482ebb0d16461d473c1
zadd9a93bad357e720290013bc6886600ba9429ae407f2cbafe87c115ce4f28631f5ae583b23640
z909d108b4ac87d84b2a6f58480f2c3eb2aa5fcca7208c4e68ba90786b761de00aab3545348d775
z49559d5c2a54f1aeafe906072077c1712645399c7c0b09442bb37d22b93dc3a4684bd8684a4202
zcc8b113faf2e1343798375da1133fc4ec911b5597ec562dc9eaae94bbd368d22c1f9686ca9b6e6
z54eace31b8379262bd0dc3666aef48cf1091a215c31570e1371afe82ed9c04537eeb8abff08606
ze39b1d4d9e75ee4e590e0962fc5957f9c7d13ef78cec4d8c269bc2d4fe3f36b163915cdd719db9
z287c9860f50d98f44b2ffb59f48d79275bf48478275886192dbad34e69a34753bf068b70b59e76
z389b50123726aa5a8832e2261aead170e3f75b1e283b37a8539ccffc1c92cd2133dee85d7b4dd4
z54adbadd9d79c12c6c835adf2c09ec3e1cbf89d209ec9fa8b7198b8b19b5a714806ed8ba5a93bd
z6e5a9e508135a3b2c0dad8d7e1837887b2256e1092642c17b229313ca7c50a61d7d41a871a6f7c
z33b3de265227e869a05ac7049f10d7e5f1860c334673643057d5906b21371229076233bee833e3
zb4741d59458377c0933bd642f4de0a3ffd96035c5ad8ab4673a7ad1825b396cdef8f1a7acecee4
z6e293854b9f53d187e7142d4fab863edf7866cc1cfc1aa4f2cf51d20805464b92f54cb230f0752
z0819cc4589a803149a73e4b99ad2ba3ebd13d7780653ffb15b9622fcd45b4c48f8512e28e68750
zbfbdbc410d86d98b63f9bb76fc5b8e16b666c9684789491fc42e3942fe2d87a8a883ec4aad77ca
zb80d48b40413c1a32044d1f6b42c06e81fc8f703d7532ee7efd6f42afa259722e7e8e0ebfb5557
zbd9dd624cf0edfb74ad5c3e519f71d78cf09b25996178b2c91885632ce55140754fe3f180152c2
z0da08ac0af9122f4f3bd44662124e95aec59a7c81cbffb5adc442997dd719ff8cdc454c405b4a7
z742f4710146a3624b243f7e7398272c0ddcf78e83def3a8bef2385f6bb95171f4ce051b9a76c9b
zb2adf61e0f74b546586d741f633af6188050a932068e32639d6ddc6ed173161f4c5e136c14c21b
z08f5a89c344cb39073b418b75b5fc49a2b233dc1ccfde8d57fed2e5565519c42abfc6cbf1a0abf
z6debea9ac4258d9fd111c83895deb2a365eb52f51c638316fabbda76be43b150e7a21ffdfbafa1
z96b1e080e15fc9509d5787654b83902da8163b13600313a8c991ddc861f568c1ba072566d6ba12
zdd8e62691ce873d3b82a120676e6badea928e452728cdf7374eea2f5c647c7102f401ac8c6b8ed
z41132aae2020dd61d633ce1a00f4bbe44e0ab6235a028352f058c892afc36b436ccb813c8708d8
z93aebe963f1805d96a509e588d4c83a415a813d3243fda4af00d9b09d8d8b83433246472f2d1af
za0f08c55b422f53c17a3c548aabefb26221e8076e717aaaa6dca5b585f571deef1f0af6c2c72b0
z889223de2ea30c02a6de64b1c57ed269a84f9e9b18d96441578c16e4cd640d7c3f01171f0b3445
ze9e739bd9c89ccbebf1f2c09b6e3d5bc77588bb1763eacfc946d2dc0cd15d26079577e6ce64a73
z5e34c61008636a062282895851d1fb6c3847b78b90961ea5bb6ebbf3ce5affb77b50de44a09386
z794f396d56603ea3433efda86b02000c34ae33d72cb22cbbe998457db46e64f9331b3d85cb2556
z3f722f90ef74da4a3d1f5df4dd6963b119f8951a1124dc5302e1f13d92b4c8f5646ab8641fba86
z640eefe66f9b0216fdc9cd1c17a932b327c6ca1a22d6cb6e6bcc7a38dc6a60c34d2030243318d3
z6e471b95e32d05462fb3d8e4f0eca887a26a5080b7af71ac33a7b3da5a3f71a963c0c0dbdef818
z9b8577c70be5873d321218831bd387ee8b3d360fa14b35f771c8ae7355244354d60210a485c123
z26d6de3a9d609b558d7edb8cce2252e1777bed84c45b7e774bea37a40bbe3d9378de2c7ecde6cd
z0f118979e1dc2ae64aa9bc8e40f1a3a8c759f58126368f06fdee229611406691b2efe7a12bfea3
z9f563b6e54eeee069637e396263e516a765100cbd8189fec755a2af96dde7c09b5aac7683ed9db
zdd20a360068373aad17b8b34a3f13ca4f7bb1063e23a7d37946a39697520a9ef6e27efad3e5d68
zc51407ed2a9745a26a331e5dde9069a2013d05fbefe9b0ed4578afae4deeb8369e739c4eacf8f5
zed836b693a7ae01ad4e2e3ffde8ac7e46f2008b369c00007a70c822469454a2c3110a86ada13f9
zcd20f5640dd490dd327733ee07bb7370cb9c8826ab5873d39da9ce2d4d4374093e3c23f872d08a
z165b46f6ddd38001c9bbcf5f40c6f6e5e6f8b54d763e404529877b32b55189a81acdc1c0f6f3a8
z7b1bf6389b49cd6b5b4792d31f316f7a2491842dfb966eed22e819dfe268de425e7617a60fdb7b
z0e4cab0b959386dea4ea6b409fe2b58331c3a24aed5d4ccc7bcab9020e8c03df645f63a552a630
z4729ef78ce23bb9b16591bc9ddf87ac20d72ca0de3c3dab98f847ca6ba58cb29fc0521527e1f5f
zbda6b5ad68503189f57fa69db0f9af8bff075b806b4b8751bbb980f50e7ebd924de45c980dec63
zb34b092df6d85bd9348019f0303c506a4b3e6147acdbd327188737c28da810b7c7c21180e162e1
ze50eea0491f2ba1f29431e90acb8a5ffb881320dcef7895db9df351cad3183756d5fdd4825425b
z8883e7e1fc09e153df81674f5e615d3c394968f0dd10dc6fd8024a990007b015f9dce668200442
z641f295ccfc61ec05be471474a98c465b557dbf09586bbba3c08206db24193f7af94c4860cc4bb
z5af25a6ce70896641977aeb03eb9a821eaf6aa3041ff3fb57e049167211483541029939c38c72c
z54b495171c1a70a5d0429e1f395174059646027ce13ee4c226d6a229b3a850b4e071a0ba786229
z5e13182957152cd2ccb147a7bf9dca902cc8cd377f3330c1d1a4741496904f4dd0d646d3667c91
z9118774fd5b328c7d38358edfed935f4d8e3266cc4e7adf60f87eac2505bd4eb39798d3ea53029
z85c0759734a3f0d0e9c4354dda2d16c2c56115f895db718a4349d358711c2446951e57db40733b
zd75871e3eef998c188eb4392adfe278c1a707563ef604bb089f43b9be290f32c8cc7ada598803b
z94e99c3707abb5e7afeea467698b915e4205f7f93354315024e4bcc297389f094d893a522956ae
zed56ecf61674278b6ffec5d7dd0f3f6002abe4cc59e45b42e7938391822071b7fbe26c7691e1bf
z0f733aad284cbc46f58b838c4db68c25ce5a01c650cdf6cd1e541689a62df7e19f475f42f7f5a9
z5183cb285eb2d74a003e9ea2a6947bef6cb2685cdcc8fbef3efca798d009b1eb4eccccf4a2429a
z9e361175f5aa83feb42d6b476803518dfe60f3e2893d5bf8555e34b629e710fefab6056992ca43
zab114dce241dbdeb574004be4d1f034897340a00783d6f5a8ff595f6bfbedbd93e5bcfa91c30c3
z9d9a4bfc9a562d069e34c6224eafdb59602a89279b53e226cab9d4988f18ee5e62f23a34b59f22
z766e3b4cab7d5de708ddc41c3705442d07e0532ff94dd2f1e006d6e9f2492565adc02c3675fc09
z9e040e35415f555ee389f4c6383012d1ae195464ab17dbe596d0cf58ac051c2619380853bb4cc8
zf3c555f119536a2128f0adfef0960c0b27e78d3feea56b613dadfc7c6f2af3377caf839a1d160b
z11606930639cb56c586a0a9789433335e9ea78fce83cade1d41b307bb97559657127fe7f6e4fbe
z300f97946e3e2eb40493f36dcd88cbb1d1a03acb5499882b7060b3e43e21251cc38c2671b9a497
z12ad3483119b5f6d6cf1278814100fc09751fe19ef2eec7be0424477713b73566da540066fb289
z74103b9ec539ae56692d92c46fda5d15ba1b1b4b07190bf76d6a2eec4fc486d320222c99bd2028
zdf4afbef74429778a3fbe7ea64f8e71ef2ea8340ccbcf7e31f5de007d235007a7c5aaa9727a520
z8c25f8943467e62397b3a7344f8be8e344294e4531df409588fdc8b26844bcca1b73e06b6d3ad4
z9a0bed9fa0d3f796918011b6f87acaad8877216dd746d0de22e31d9652dbdfe82c6fae14234b9b
z2b8b0154732aa11ec1edd4316793b2c83c2397e81114492fa8b097731f494e3f7e1a1d3e3a509d
z93af2920fd20159132dad9bb0c8043e779901a9bd93b5049b1b93f0c46ff3537dd015b8db5e83f
z2fa7f1db6cc27ebd689490e0efd3626b71b909c2e80f9167e5eb111e996e8f4531515e049b79a7
z552db25b250286c04eb92352ee2adc50eac30292a6cf61f4b57548d810fe745e8d703e45b5a21a
z2efc6b3aafaf1d982352944b6935231a9eb207f73e97ca45c3bf06404c2ceaaf20508a2b15e540
zba233c283e63d51a83e78a1099362acc1434177645902df2f0a6fa35ba81f347cf236ca2248053
zad95082cf32ee053b819839d7530d3331e3886843fe163a5586266bd88597eaadb537dd2d779a3
zb7e14f1a315347bade9b75a2a7068b925ef11c6070c7c2f189a6bcea9c3ee1d630850d07e70de8
zd7776c8b6c9b168f616d05aea0dbed79fc53f41f00cd7bc4a54ea320c909d9a5629b0040ee5dbd
z3773fc1ce1c1f09dd3032836e5788990e2e4cc94baa8256c441930445da316a5650911926b82d8
zc4b2e5d3561c06e7c63e8de8a2f91de2851d318aaf90b816f3342d4d2516f4f8a69b5db8c0f4c6
z7a2a1082f3a85f60fd43abf053387e15b81b712554a2775836d1ed2c752054c3e651b4ef8529aa
z5871c72f0b56a046612d7ec86403f86498be9703c2f54fc2edf1a3f7fc263fef99e8ca2f637577
zaa71f716f374fd82847025bbf595e58311184eede68113e24d11fbfb5144f7c674011386f6f5e0
z83cc23e7b05bbc92f5c6fa92754cda603eff7aac84ece7dc649d92771fb55b41bf8ae0d350b3f3
z7d294ea589141f059c788c4c44bc6102f6fec31208ab40ee185a0e2d794a1a3ae581678d0067b9
zb4b2393a62026300618424858882aa61a8e6f3f6d78942e2b9efff36a322c7b4e8e5bd01f83956
z7ec5b89f1169c3f578bad4c48f0de0a67aa1857ba6a7eae320a0af09f8834b36bd9d000fd71ce5
za73ba1d08937f607e51b9088dfc025b75371e6d19c731c4f6f9bbd1eff860b74fed23b093e0f95
z064cd5a9e95e46062e18ae2229bcb82b10ecc99e6b30afb59754189588a58bbccaa8e1d701945c
zb53cd5453422dfaa451883f63b16006538e47ab2dfe383d68ae30911a6d7c554aad6710ed43602
z3fe764cb7395f875f3b8d3a201fa533c461753159d5ac1eed7cc35ef58b71ea543d71f807de6c0
z00c323bd1ad545b69d257aab6ac6525d8a88b3abfd25b1315a5d562fe88201e1bc98705c65c9d9
z849ff384bf0c9d1962b213e5f53d2973666b768c2be9ac2af9dd63d062377214aed88700162002
z56871cb3a278dbf21b1e7c5c8abf340290a543c4c637216bd3b5158118beb716bd565e85350b88
z70f350b8886720211fc38beef8666168ae4f66760efa465a8ef2fa82ef3e15f8345f2c4b90fcec
z867671ce5ccf617a3fec5211bd2e9b62ad7974df56a347f0204735e3218666a241fbda34eca64a
z87bf8a31cc653c000db53476c4ab0a70d8933cfca1900804082f96776426422580781694332a19
zd5f0e65ff86739ddd4552fc4ba791e1de497d18f5c1b2d08e6b530c9ed970994866e71b281e7c3
zed9ba02541320b1cf163c5291729f341779c248a0a450862a707f56933cd189a9b1384246a8137
ze8d969c23d586234fa308e2ed58f3c094f58d1b92514bedc16c8ae4af8c7a0badf01f29ac65939
z4991861f481e4363efb5b29d0c8af21d2ce91420dfed48e6e12af6c3095c5686932f4befd0da91
z5b615aa52b8a450ea9956dcd4201ab55c75e3aa021c8576e95a9bef56f86572f29cce347ea1dab
z0b1a78c4f5c17fcdc02b4b987a27e024ed5ce95a491627896e6f4a4ae3e5ad358d413cc164a68b
zec66233235a59e5d59a29d24c324695d38d6c1329d328de23a6a66114c8af898292a7523914b96
z25a68ec4fbd477c0eed24d77c827a64ec342cd4f8452c1d2dd6dd6408e53775f870769db90f631
z383cc4cb7c9e6239a62f419a38d0093568e4384d6080c3f7c87beedb5510fd34eceba65979ab5d
z55b57e3b3512fc4272ba54695d21f97f831851954a3489862be066251f74fcaf5d9cfca826d727
z25f40b9d7eb290fa947bd3447fd26b032375ab5235b7dbdc1c541176bb18f97cd49643ff3479ca
zba8eaf198bc399d29437b15583b340533b6a8393062d956c3a4e053157aff3f7245a6eb8ee4456
z4153ee30dedbab9209a49691d0e3c5380897628aa250fbf986447bba8598369bb54e48f99b5e82
zc463baba5cb028352ff8f1add2e458a51f0dd407a2f178b63ab8a61f7eba9d349454b29ff4c92d
zb1b5f5e9446f162eb8aa00d09e903dca2cc12b343c788d6aaa630629930c946916a586b08acdca
z786ac67538381bfef1abe274eaa93b7bb33765b00ea1157ab69c777f740bdf9444e373a65f8a06
zdea2966a1acb4880012f20fe02bb13e56695a2bbef1a1621932adddedf679802bd34ab2db4483f
z4f0c2249e7ec34fbae157fbfd01afe275bf5d06c6d00eecb709acca81adc7883fddedea74bd9cd
zb746d5691809ef50c7f9ce849ce9753fea0541bd590a14c70cd896fa877381fb746843a7b90266
z82bb29dbaf528df74b66cafbbb7818ccd5531a878b73d4bf418ff5ad71a7180ca6e438d046d4ce
z54515c11338998128dbd9fbabb3c6eb5b7937317b1a318feadf8f2646bd6bb9437de848097c293
z2afcccfcd5a977ce9fdc06b4b0bb6d0c8112a627f52b793e7e76b0f59cb5378f43d3bbe52ea9e3
z28a97ecc11f5821b2d83f6533388e9a5626a95c219396417f0dc3ede4ed9b915272be6d68864b5
z83d981f33c47ef05f5f1251d791e1c6add2a9a2ef0a17378ced92825396c2dbea789dee29a2656
z978f4531c7856c46cc3ca2c5e37e9b3e3d71ce2134c9788bb412dd7cfcb2a758b6190b80a675db
zb7343f4714e72a7d6475d0a328e0ed173012dd39abdb17ec597d0ca2b9f0bb0c5d7e98e132a57c
z86d047d1c34dd1da62382d21cf0c7926a3872085baf072559d535dd1fd576037ee8187a132e1df
z476557238f4122055733fff31eefc548a27854423eb472a2d84d96e5f56e89a169c0094c84e4c9
zd009264d28a0f8a47ea193cb7afe3918eb7e6478f5f00eba03e94856331c193b8b70a1dcbd7485
z642b94a88e34765545f7014bbd9cd806f6bd7223ac3a5d5cca514f5641f3c1937be1398a9ee7c1
zb479e59f755d15b114cb019bc25cf43decee45defb1e51b850bc3267542ab820af4c6a8aa63970
z8dec623cd528bda07a71ba3c9cd48299d030594f26a6339cdec6a8cd1dbbca2b2e07477dad3984
zc4918ca572662636e0f7e17ea9181682f0de16cb7364c444640a51e97543807b303d53d5171694
z64924d4e7871bc044a03792bbe5a66156edd25d9a3e24cd9a8068ea122761e47e0ad642a43659b
z9e5ac4a5887e62e6c498311871aa709756fdc83e793f3b4be6bc7ca7bf4eedb772d771ce799201
za97b7df17a3c0930b4756c4480bc57ac3fb57cc99e98ddb503ea662ed3f62a4b444c9c46c7214b
zdd878f85bf7ed3d315e601c7af3254e4a1006828f43bf0be8f9c3cdaee0c5c489b72bf9f15114e
z626c4249590942238710956f9fe3b52bbf28b6c7c90621a6e9c2cc82050069cd4f1193ccac1709
z94d012eb5b281bed209670b83114399242c0a97ce101d8d3b6a794249d5ab229a3c057eca1b684
zd6c8266b4765faa0fa053a508baea5ac24dfaa65cfa1a001e16cd3acdae1c37cd6791b386c25d5
z5252d767a29333ebc5f34e6b05e0a5a4dc2b2f75e2f285865e397b134a69069fa7b4475fc6129e
z187925569403260f44bae16e04f5281c04f73b9432236650212b8ac30c3fb4e01af552231fb6f7
zff1c4f38907d2584000b4ff819be3048dfc01e284b98db63d69ce000f768f0480e8585dace839a
z430d8b7233eecc4d512ecd45f1cd1564e316b3a8ea30a6c9c4b555b927fab6e4e05c22a8eb2d25
z069ec774c9698aa9293269f108e836bfa70ad40af51e8998d542a0a468c12a657f2cf791aa96c5
z30fb8df2a677e8f7215e73dc07a6230f010627d8655ba59c97b84acc3342f883140912a9be25d5
z5b59c0f9cedb02a8863b9bc2946ec7b17559f268cac8e2150fcf9526382ab5d06d3eb351ae8564
zbfaf4eab62116cf18ee6413c967ddcb02375ad4b329f62ddeec0e0cef17952ef4eb50cbd2555b8
z5508a1030dc781c5a36fab40268488c8643f40a8f2a32f1cbe5472a18c2b9c004d9bd72e201295
z7fbeb8c7c06cb6793f49c52caa59e6eb3dc9693468efa7c1a5bd65e87e9db6a214a86597a9d81c
z844892afb3d395ba0991c921000a1a6b7b9eb526672bde17d1070e24830f2f0e3a8450a77fccc7
zfa19c75a5e5c7d33f3ea81fdbff033e5d3ad9e68cf7fd0126bd7e94e54911bbb36b49ebb2c5a7f
z42d9a28e8e9f2b30128a05a50d727418ab161aee10693a4cce942cf20e0c5f21adb6d613ed8fc4
z9031e7fb978550624de97bf85de3c9b6e1183b80bb1c3cc0d803c67ddb75b73cc98b76356ddec2
zb138688d5d22a1b4edcffb0c9689163561a5f166d2859f8c6041da0d5c8d8f64639e319ba72803
z05f2694ef05a732fcc5a154c8060ac0dc2389f1dbdb1187ed0ae2dd44e18f1d4015e1764646206
zc6d8810fb495422abf5fef50aae1e5b3cf15ec9d46c1551acbcb0bbdac79185b3999ff52ae99dc
z1e689e0180e7456901f315c18723fa00894063b5b6b6914b86bc61d58965b35ec66e8b9b955f29
z2e0c0550d6c8aeada02e222b36eb16150a038f6d9010a3c85357deccb9fb1143b039f48a49b936
z211bea062876e9c6d0bd257f15bf2a8f207f0ce6528adb648634ab8f3534a2ecfb45f79e0e2882
z4d80750e03bb88297e1b0380b08d1d30f4c553395757c3baeedb7541e49ece06a757b3e1a15d2c
z4daef20fb219db205acfcb2b7f9b96c8fa104b9c9926e0f411d67cc376aac839a874f3bd91b1a5
z67b2b25c8dedfb9e493e5f46b96832cebf490ac87c897b0a7e7bb5bdc777d2e09747eb1e2742b1
z482664725c06610a117ad26b3cf230dd68ff066fca886f50753db90b8a6400d5fed239ac4b018b
zacbc16226a17180464a010e053ccb02929672e00a26f4882ede1744778effdd79809d17c1c8c2c
za66c9c7179f187e5dd5eb1c704d0d2e7263e1ce2e3e44e3ff9ee20e267d204e0997c0cec6be144
z747c4d3f7c3ef2af1ca7c46189180c10edabc4430e2943725c0bfd5c2e2ada4a7b1ae55fbdfbd3
z1ad1e3dc0f33609b07981b83640ba2ce36e6c7e81e112a2db3bc18aa947cf496856f768e1d2964
z507000dd93047e16ff84c110e62a9fccfac1c0d6fae87d0e009209fa43294b634f1fca740571b4
zfcdaf4c77d58db7287b49cba7d9165827d7f31adda98b66e2fda63fe473da6230afdba7c93e538
zd3899d9803d7d8f0500dc62535edd0f69e21f13d576bc30dfe22a872f4caac1614076736f802dd
zcaf8a7ca7e8ad686278bc06469389c50f8c1561f2e64cfb01c3853ef0426a11723f6a1c99fdb00
z15f26f216fac0812515acc96771c4f98cf3eff3c299880dad01e45aa8001979e666885110fa0b9
zb5b185487f1a65ca13e8d7efaacb8ac547828c88012b6f7eab6411bce7f405cb23687818b71bd1
zf2704a3c3ebecd357b773c6ba40a8f446c59cc5646478544066e867f257e295bac494345933426
zffb5828da215025ee82f0056aceae40bd5b773949115ffe21a707fd99c8cf7d17b219774238463
z5243a525062f9b27084cbd48009a7d80e95d6dbb459f12d262d175061a14b368c16efd2ba196e3
zbc33c784352d796d2d272d8f6acf4a80ce1a152e1c9241e1439b97bb374a082570b736aee6f567
z84e0ef59161e3d3596a768107ba8d80a50af170833e876692148e2f4fc6b62d0e02873906affe5
z59007e0da6f568786ba64c6532bda88c4be17656752070d67efb3d770fbf4bbddff3626b1409e2
z67caf38637c1cdd8292102d04662b0a1a4f737d08eb8ea198be2a9a44ee51fd487d2f4bbc2c220
zfda024de69000509de8a51b6b3cc09f63ab49523a9e5f16e59535111bfbf72aabb0973e30a9b53
zc09ceefa8fbed48249ab76bc93c1955aa23f7af79c92b754ee9eb47f3454f7d9db34640caa9920
z53e553ca618ce80b5bd9e389e9b9c57f10c206f848f51996db5302f930d8020f5b8d939df429f3
z3437f0d55d520a7058c7b5a734ea90d8188b3af747bdcb8f013ca92f8c256e21f8cdaf275226af
z913e505e51805da05cf21ac1b7c237f3d9e2f70df0c783c8b07492ab7b749ba77cc3169d4a7560
ze64d72a9f79ddba472cbc211e201e73efdc69575a08539c02310c6aefc5d297cd35b810e724212
zd5d68fd72cb83e756442cba11c603b5d0223a2b2e9aee912879ece7e01700978281ff39da0e211
z6140bff20233a026978e3624453ef64028a83247b7a3cefbb7d6b43b6f6b2d50430742a484a0b1
z2bb5ff8da38ffc05f8c2a1ad37b7d67a1f151cb7cdabf2cc8d8faa8fdb6cfa7df057a49f5362ed
z8e4e8959f915a39c8a3b7a9c7de674d5edbaa9d6f2dc2bcb5d7c49ba1d15133c541b0f436ed99b
z47c4bff2b0495f175ca59ba6bad5c2e8e2d7bc794df9ea9b9a9b9beea5a6103eed1bbd759829a0
z479c0ab8db863b487ba95a2f96e70df8ed7251f176d859a35e6d0e575a4200d8e86f1eb1930406
za2294b43192b9501bee2cae3d874ae39feaabe5a9a582c317e858603f9b788748ecbcd8b4b8f9f
z28d20fd46bf131d32274401dc0bb52352c56cbbafed96dcb3002ebe68e6a3c421e3cc94d95983e
zce072d95f95233c02cb112d49ac07d57498af21ef29ef15593f02522b9e668588eea1c93807d14
z0a65c47d127d643d88b94760363fc611be45d1b45289560a890748f002e8756149088026bd074d
z291dbd2869f150c076fb5225a9ab229041fbbf38988e824072ba6837ea31ac1983fa0824eb7e64
z43e4e8fb2e25f50def5808634c15c2fc0355700b73883440c0b6ffb169604d788693bef2cf926a
z67eb47618910b8e16b27dffa98550c07bd2d2de3d45e1a4ed61544ee0b2ca0d256196402459d4c
z66a7eb4caadfd1fc2c0471d0e1f7ef524b3d783bca409aa4e7da4e128ca7007956edc2892e026c
z201b93f2e33df85122e3f6de562b443cb81ff55b3a4914fcc620c2bb81c673a8ff8e51dcb77ab1
zcf446ca5b1403106945b523ae76bcc83a00702f84c8878b436238706e292b2b3777e53ce1d6a8a
z5482dd5f625ac810f5d047dca9c9396ff1e611f1b722effe462c4f5bcaa750c15d8c1eef4091c5
zd99ba8a4bd0c0bceb23aaaebf4f89ebb9ecac972c911861241849123a54c85681d4071837f6e47
z0fe125fc6c0ad7851be39cac7da2a0bc2120fbcce9414ba9f5a749a8f2699607a8d18b78d58f6f
za8a0498a48dd9ca9242e8d87da4b1151139b6ac55a7a970e44e42dc59ac026d0a0d090c0b28825
ze7fc049f20cdc3fe04c580baaa7b6ff8a9ab2bac16fd9af045207253f60df15821a9b6115f435a
z9fdc9fa0d059dfd634db32644729ebf707396923ac9c3ba8e046078fc15d71baccdc6f6605bd98
z554d91f95d324b5c7d7f071565bfe4d1032214a4a7e09965c46186139e7b0574153a63e1e58ddf
z8374a038b4b863637bbcd50b1bcb4e152bf00ff89ed3102d52d148ebf94e07661357a207e089cb
z96699c64ae8f1c82c876213d60269c3166c12ab2cba453b131dc3d286c18cc9b0c923a3ab7899e
zd86e1a4b46ee29eefe1837fda6353d88a8927e1d0d9d82448267d7994e0e6aada040b18027e1c9
z4e18b05c373775c4579660532887f5322ef686b702d4703b95744fecf70dba0d66dc9f11c0dbee
z7e5d4eb6ee88ab53567148ef8d8795453762dc256e487463617c4cf4574f00610929d105ed3bae
zcf82fdbf3b857514b4f460bf805d6ce1cb4b49799975351c7feed160de7692b864e1e0e2145e43
z90b6aa7ed4a5047453741bc5d11cc5bd9e8aa7b710b23fefdf959e9658f8f4e14a8476eeb22f84
z6c859b3f634a84e0739c99b2cc6a93666116cbab65efe9bb21711b467e3e1753f54efd9903fc92
z70a9de49f01a1fe1b2bce012a22cedfee36e06ca634ff25a9aa93a79b4b03d4facc71fbdd2600d
z44c4a92e801430337943c32740191982a4a2e410e42e66fcd46d24a414cdb60709242b9e1f8068
z6e9dbb89f18c8562e7149d720f80c32ea4ad1aee8a1505d2ca2732bf9c5a053e883dc0ce64d34d
z1d2df245672db002e7851d7c7a32677bd374610f84d1c9811eeae5fc1bf07654ed426a41004e60
zc4a2278d793c3cca4dfe8cf191b96df505e975bd41b46025115c1afd2bc8a04d68099e1a280885
zb761ca3b203d64ff2caa9450757ef56d80e921eee8d9859f4df074b02b33aac53b6346c8585cb1
z956239990edaae129f9ee231e2643abad6a5a8e90652315e5966a5434145b71db73ec26125f6d5
z5227c29a4e04aa820d9fd6fe18f56e85cba12e0555089b938999d5701be155d67e7162b213705b
z3e232fa0bee75b5e09c72f2b76a093972b8c642db972139bc840f69325e04db91a9a11336796ff
za697001e0a0a7f73a20dfa3772223c7646bdb7fdcaef163200953432b0410f944ecf2f10539e2b
zf63640862ba427b82378c36424a5d0eac1f4ac9d7663406958c43ee0dd765179427c0b067e5b2d
z399c941db63ba14c9c6c4b3f4657d01911fedcd7b4d451b417a5b8694837b5431a891f35b6cba8
z90a947aff1b3565973fa959244720ca6d0ad3c923571de11b277f885a4940315913bc5bcedfd70
z75c06ab23500832ebbbaae1a06b32f25c7c187ef6cf7a474d133731dfe940119b64d55c82ed2ec
z2d7c6890de4d31bd32b9509dc58e94c41aa2b287835ba75671112210d9387cea85e78cb6e2aa63
z3048794abe16181749ef3acf7088f4e7273c1a7785de3aeec4019b1b7c4a56a4867016e68032f3
zbc29a26ccedd8928fdd47aeb54a5925125a328dba3c56eb4b13d32c625a4e5fa4ca22216870582
z123b1c0d4aa532340eebf4ff45d106eaf6725400f521e65db9e31c4666cb9245835f1bcaf20ea6
z3fa0d2290985cfb70268c9a8e9761bf3829992074561cb51512509c29fa0291b0d7fa944c4ed52
z17f567416f87054f0d7138e129a0d0fe4ba3435b0ac2033e638944e5953c2761e5932d41a73c3c
zacc5af1ebe552164251c08fb38424a7c6c608b682528e53f9c8890d7c2e6524770fb96a06bac0e
za5d36149d45b78f6953e26cdce8b7cfe13d144e6d853121c48a8190e2f6e6556787f72f2057bb7
z5139ca1f9503bdd487dce3184f0d6e0834e3e2ab618201a31228db95f1e4f239ce9aa1ba666fd7
zd13cfdbd662e62597d59ed6796252b6464ce0f2c4fd8742691bc55f496020fb76170b2b4d58374
z6bfac2cbf49b2e7d08774d57001d70736e2ed25ffd6a4b5800a54c36b08736ad8cbabb29d5e845
z8cc59e618db072361a39d1ca66716065a0540e0030ed12146538bf284c84d7d1a81ba5cdf87455
z5111b416b074e380f63e846fa75988a3cf0a6093e286f582a628283913b562e8517a079e3fc47c
z9766387da36f612733be90117e72650dfe03837d0ef4b917308746bdfc09f41b360ea8b621a617
z163de16b63d0a1a8970066359c68dd51053484d91705674fa925769d5c0774599f5d9e625f43ba
zc7559ae8a1994485b99eb7642e3e2afe5f7dcfa2a06b4c95240945ff6688dbe0b771c327f4f4e0
z73814856211666526fb8b6f62c01a83df59ad8515400e325ea43080b89d96f54b52a0962265bec
z31253d0269b40c23841e8fbb7ebddbcc41339c7f766be6c33357105aafba93c496017af67814e3
z3f56c2026a94dee807fa319e767f2cd78a76dbb4ff1d7c2c12fdc648a01d24125796e0b24f497e
z7e04a825290aa80c56fb98702eced9f0fe3af29dc2eb0cc0c647c0a91761ba9be4aa296310582b
z39b32ef2059c7cb788dc3128022ad48995d3024ca0d70d6d1cce3170f2ed5ce3bf086ce3f74f40
z11c38286c7ce80ba15fc55525b949aec17ab893bce282afe71c69e7458dbacfe60da20d7ed77c0
zb997af663e03f6804ea2a2a9ec52f523ab2d11f02514b09564851fe9ebed6af43d876e17c7255f
z30f88991eeddc9b80a3101ac289c4621f5e2e7fb3266266a022d4e0c4ba4938c95ad287b756645
z8f1dd86ce10a475874a8b3915fd3c275de6818fe37a2df26c2cdd16cc25d17ccbc14fe800f52b5
zef24f75a035fcd880e02192f906a528d5073587907aefb59d30f7b695a81be873e48540210a2d2
zf803df30e50d3570310557be7fddb3eadf61a8acb2a57be47aabe73589382848e1db34b8a031c5
z66216279ac53ec0f9dd2377abd0824604cef7bf3c04e34474a5ec69146317708427ce9e166655c
z7762db4ec4cbf9add52a93a2151665ff0436dfa3f4ac6797675930e5903b0c63e7fd69e771b02b
z92c5481321e9e07bbd91ff9e22e46f0709e741c40045da7e8e9057ec2a5281e42c9054e62fa3a1
z5622c42baf88dba069f91a8cc66314d48f470dd4df912c0bb656cc12ee81e9c7773c6b18222286
zc806b0cad1e15598bb561801bddb6ba51998fb536fcac7525b04f032b83e15a16a429d0719d9e9
z3cf25d6f9e6d5e641ea030c67fbebb320a6a57522c055aff772699a2e94e24448e0392e299517f
z8cff49f9d674b8f52635985f781b41421f0787d5fa5cddc0e6c445dd867c09e98883477b22ae3a
z21dfa3ab7b61a10f3a8fe8128313509be9dc16090baa6d5e3bd1516c21a6c96596a68c7d00d7d0
z5a46169867a34cfd77a552f4af3547ca1e2fd1aa532b93ec4e43ea064cc3c8eab294da9c94f433
zfcb9531c2189c2c31e0837d12ffcbcdbb9a074289e4cb6515d11eb1e78d45cbe096a92d92e03ce
za6ce8ce95eff3e8af4476fc39a0f73bd80ffc2d779c257b3d65881785db6b11db7c65064f6ba2d
z19f26dfc318b641a5013cf2541a48ca7476e79a1ddd9c1ecfcd1e31d68400a4adac87ef1a972e1
za7f42fdf267532ce56e5ae6d8cadcbb3f3e40bbb2e1b14c41c729e7b5f318faf9609e5416aaee4
z40f987c271aaa4e12b1b52dc146074d97f81f28905afb961479aeed7d65e8c6f95bf73034a463d
z6654e43e9ba3c9b9ca4d2526dd98208d1f80056b1fcdb0b464fd820aedcd8926187fab8a8190ba
z46730de27c96d597b54d5e108fbd9525a2e1ebbe39a2d38977b39a3b16180f4bf37d8600247ca0
zb8ca13dca29e28d862b1d2151cfd862fb924af8bbdaad7660de353f85a72c59b6cfc54c8b5fc96
z3fadb87f72b4c12bad34b2129e2c564aa170620710e0534e2bfb6304c6052510238fdd2c03a2dc
ze5e5aa903426bc16bc1ff34a99f59afdf1390b0e9fa3959b595e76825935894ae891a491c006b4
ze0df9a5cd11245ab8c189cfdb1e7a1e7cf4e77efb5de00dd8acad7a9f58204a698ad25ccda9bad
zc3f89fdce1fa95e0b46fc5b3c4454917936b99c8845864101a467a03096eedd3c5e0938a514268
z9c0b149f6d8b550a479b29d76b4cb3dfaf51eb66c7ddad762cc9c42b4309e991b0670f0cc41ac0
z19a3e445789c539bed03b0f71e9228ffb257a2a76d757c9e33a420d923b1f11768d5d59a288884
z23be0f5cd2ac7a193004b608e651fe24316a6a587bbece60547c14af8c3bd3d26bc03f244516f7
za0ff517b268e5dda2f0dfe67e572683a958d46d86d81d3519091b4fd3994d0e334bbd2bb67830c
z506f8a2b6e5f2bfb220b33c6e75ea0d91cd79fd5bdd7210eb87fd5ab5c2de9e003fdfe32f4d702
z533887784d12e2a2d887e159bbd9c858d10429a712c5d79716c978f0a93aa066f538e495a8d5a7
za3f528834023047a407525aee0cbbabf838ff7eaf396a228cecfc18646a591add632ae9e9dfc56
zcf054ba2033c280bddcd4cfe209b02f7a1fe05f62aab200a525205205eae30de46ea2611cf2ec5
zdcd6ecf101fc48124468438829a959988ef197eaca61ddfd6c40133540fba5572d7fb7c0dfd633
z5c13c6ac553e7c6bfafc5f2de64ef021184759a45e5f89a786e02607d6afdda2006a1e28692e50
z7bd2f1ae6f8c668955908875339a2d1640555faf002a9decfcef5a4881c10d55f1614fde4be304
zb7fc7072a5770106f03d3681696edd86cdd0ce5e36297719b03da590db6c810e89a35470c000bc
zb02f2af19404e1943652c0eee6646e927f86c923d200c8e795f2afe93dea196ab2f05a9f15c841
z33e878d9e7add2aca7c5347f2ea1d82a1546a23717ad23dac955d2a3de165d73ff7f98ff3ef77a
z4eecd5a80f4b22eafabc644ac5eaaf7f49685757a409f33003e414e710b5aa53c7ac0bfb0bd819
z1bbc0abd98e0c58db81b88bed9679462fe8262b01f7423c5599776da53b3076df875ac539f79c4
z76b028db744b02f75dcbd88e3364feedda21ea6c70b41686d8d2e5aff66745417a02ba5a9a4778
ze926f9f48f56b46e3e2822f49129d9a18df579d61f149b3aa8ff395e4e262e53526eededc4e513
z163a7a302d88c0c7f76509ec24dbabf1ebdf558afafaf2d14bebd2208ea68e03be810332e4ddaf
z8759bd43a96dd6a2763f3c46a278875872fb7b25fe3211dce31f11716de5c27f715c4f3f42575b
za84009f9dfed1bd70b1d1a4a575529f4a7318e5a61a71f170b07505515dbef0a14e0c3331f41d2
z8c22e6d941c461808c8a59bc3bfdbd64d52a13df4567577a938ac6b05ca6f0d1f07e2466b295cd
zbd02732d0446330cbca825068b91bcb12a75db1da7b17ca00ac3f5c4aa6e1fd7005f566a8b17a0
zf0f2164cd01906ee95c7d96a5608b73d3aea72bb20c921762a2a5dab9279ba63228a0fd2264673
z539e69c110f0a6d0ae6bf849c4b4bb2db507e1500880323b489ed705747ecdefd9af6b365bf819
z72e09188461e52f90368307286e691552101f308f2b26edcf4151dec7ecdd832b79de1d74dbd50
z6c1e6449e542c0ab2ac2311326399e22cc2669a4513a8cce14802a15926dea33df6d16a8fca653
zc1f2d3ccc3696dd741cdab5c65d3b5e3ce7a73a8b907a2bc581bb1cc322ea417729c273d315718
z27e44400be13d0bfbdbda2ac109e70990e32f16f0e23eae500de6575b134535750734b9e87a13c
z263fa88082a2dd8153a51f73ce276167d7c3815a4f782d1f06afe0487f4a7b896ab3324c8a6cc5
z550b970d85bfef33c227ebd15698a20ed7957ce1bca61adc47229e37b0b212ac9850bcdeb4a73e
z2240576f91dc2cda07478e63601d313e8cfbeec21df2f0582d0a74bea522d0985897b61b06c932
z661275acaa9a34ec6b86c0b77e470dd2bacd7d9cfe95081e2bdff3e410a3d3b7c5eadcc9ffcb8a
z9b4d1d27fb7f9ebb2a869e7a669a2c17668f7342479292d0fc0debc39ca79594e2e9e688c1cfac
zcee90b4c6912cfbe4b0ff0bf0e84ec8225c36fbaa9323d9b5eeda7e0a2d705e24866c9fc701c99
z1903e637895dcd97faf0dda448d00b5f1bca8ed1321e4a398c39c75069fbc56e2b548f17ffc216
z768f07d7d7501bfbb68f891decc6d5b1308f82db0d4e77092b3f97c76116a1f762ab25e2b7f6ee
zaf78928ffe87a4b8f10f8e607866c7f8146296b5181ef21c72104b24f589ef93cb0e26470c8c62
z6aff5b0183b1e0bcdd135f58970b1b6a5a3bcfbab384f2eb82401db1fa901d04debd0b8c8f1128
z4bcf3474d34cad915f0b4cdcebdc7408870e823a49e66f4cb4d89fd77b4f222920a906c7a83af7
z0c5cf567bc315756166e1f28cc40238bfc9a0301e2cb55f1e28a43fe02f02c5010ea753408dd7b
z19a433e909d8ac21a392173829555a7a6a067044142078456c919f4134a2da530096d9474bbc47
zda7fb5442646205575c06b5539d96851f8001d54b2ec72ef25a66a45d979ad39a51f6dc0eb1391
z04d8c95611b8b07cc6dacbe8f20ba47a7d1b1e1118a7a788c748f2bab7808b53e9c5fe84a5700a
z7b66581ea434ba5352e5ab5961f6fdd2eb48ae7285eb49b3d2c83dd7ca39bb36e68b62270fe28a
zf0618d6edc6c39d07c77eeb9255a8de688cdc1fe3b6d713c16b06a2e2ca9b771073f4a6d11946f
z7d4fa7ab08cb1fc57e98193cae54b12452baebf35157ffbb075cbb4fb1744c75449c3b8052b906
z01a1cd43ec827f51199621887e9bf830d9f08bf342982ac7326c5ded75dfb6c2af207a28a4a972
z86d93bb5757792f001a15a809ad9c6b436971c6587535ad31d50de92a9decaa5b922e660a487c5
z20ff089bb06224106c381b55fd8e0d51c92960c277c2da0a78d466475d0b70e430a148a0c8dad9
zd0a81248eeaa130f6181b368ba7458226045c820f7603371f663821b27de1bc81038b1b61b07ad
z648f9d2a8a07005182b8fc1593e68cfc59794b02a43e271028eee31fe718a0052c3a11b3e55ede
zef2d216a9851ec3265cae90fb6525b212beee65e5bdc0492e3fb48a70571a64c188ba5dfbf7954
z89e90a6a39b0ad4284baec4833481b38f51e8544af79917b95ca9bc96ad81a4f44c2600d17e857
zdd26dba1044f20ecc345407bbbcc1c7542fe8c663cd88d6a12e1ced6f848bfc6ed7489475e6460
zfb9871a25701fad8116087ce880da8242a0f5c136fff561ad0b47a32c4f37562f7d972de8418d4
z818753912eda4e0d5a372c3f4d9c93d549972c8b80322b9da6c37689fd5ab4886e5093122d7b43
z242c896cc4a84b7d13385fdcfc225e8a2969056d2b5da878aefbc69ab5db0e3b06f40b89e70f3b
zf5d39ca2f65a527a26760b59a797063be8463cbdfca70dcd1e12b47ee3417bc9edf39d19a50933
z6a27dd9eac559c
`end_protected_0in
`else
`ifdef MODEL_TECH
`include "qvl_usb_2_0_logic.mti.svp"
`endif // MODEL_TECH
`endif // encrypted_0in
