`ifdef encrypted_0in
`protected_0in
ze74c34e226135848fe16db9ffd31815111b6d7fb642c521a3f628cf6da949865580b22efd062a7
ze90adae0e65e66a2c36a587d0a790699166942afea5fb71013544a379d857e1468025bb8933d9c
zd1ee6dbf13a517bdceefd8805aa27c5b2bf034ff41fdb5715cb78f18db09b9b634b7b7bbcc42aa
zdd1c14120e2806248f14c78a05fc68e50d53bea922c36ef27c31db4ad6984f433b2a94bfd3d958
za6396c21b10f0fc400ee554f7094c3ef3f9b310aaa2ba11e410415deadac83bb0d3e2d41e573b6
zc9df011a4f49da64c6259120aed4ef52dbcf6e30c0724e64ed1058215310e6ee8b5a2da07089aa
zf5103a681bab47fb009f964db4ef98b434358d29eed12f2da156b5d6da599273d22ea2f14e9831
z433a480cafb63cca170e18ac267c5d0f91e2dc6fd3bf938aee8854181d4beef7d4023fbce03c0c
z9627868a1d6ca65b2da89f90ef23c36a99320fdba6bcf2def3d77fbd1b74a56be50cd62778172a
z4530c7937fa834737efb5df8cffbe067256890af6e6f8c8d0815ee47a628e8edf891c02093c763
z526977ef9f28942f76a8da5e13d49f3ab799ff4db018d35184fefb04bfbef0e6e6f7e6d0987a3d
zff7e86a714113dc471d402767ff2beafa5582a2e428663c6be68429c72ee464dd1c2a25956852f
z8c04c91347ae9311e2784f1bd6426b7c3d9a85e0287169f06e192a88785a764e2f37832536791b
z1c29992e354032388b3ba6c334baa9e156ba1da1b94ea07dda889a3dd98025b027af97d1cc534c
z5b13d6e8d641e07e91009d63740ae13cbebafd5280db671d877b65bf55800e3ea33aacb2d8fbb8
zbf1aa2e7dc62ff6c09bfa48f22b1a8ffe861051bbbce64b273de1fff221810bf910df011c45382
z0480525c46fb279a7afa7a80cf4be829bcde68ed434b1296cc79eb5805e73e8d17c338d9a6c0bb
zf9a3d9588bcf25d1336c351aa7637e7ae4e2a04da0eefcb1cf60231516f6323a22f3a5837bd05c
zf2e2b074727a0c77e4f0ab93248207682772f3ba811d6960b959852476b2955db65eedc25debcc
z0408f5d6bdc6ac0ec25ba1792d5d521e65f0a447b9917b752f3159001af3953a4afe4d60dc896a
z5f859cbde5f570ae178c9152c134467a437298f1124db38c4d844afa9376d24b82d10f42eb1e63
z9f8f3bf7cf793b7443ed016511cc7c6108e7d3da5f19e526930c4941ecf44319f21500cc249c0b
z62ca50249ef904ee17c2489554e68b32e88b53119086eca8f990552ee9389670ebbeefe9b2d5a7
z3c9bba727cb889e0d983800e9fc3c677eb766af4435e23250fab74d0ac4371a89c915ae15fe0e0
z129508d45d1d415f55123681afd5aa04868d41919aa809d57d21b26dc220cc27e4998d4a326436
z4194dd91084d8cccb536744d7be7c3a1ef00529288affb6c541cbba2247d497d5d9c54c75969bf
zaeaa4624663f29d3c02269d59a248cd859fb7223c93b2ae9065cd2c8793dabbe84d615e8e88fd5
z8d8209a55db15594928265b2593b1e3b0f7bd56f04e8f0e10c794cd79abd69bc19fdd784ae178e
z5612fe11afd986e1b4a5822d56232956488e0559997b7ef9917081168397524c6d006ad99f1849
zba9dab6ee63070825ce53b0b3f227e042148f11a2f100efb1c8b11c72c24fde7e27aa8f6f31bd2
z44b9932c909626b9366327480b0f531f4f87a0590b3bb8d929c77090ed781e92e1733d18a5314f
zba79426b619de631a7b0f1bd1179fa00dc2023d17488727127b1b193503c76cc4ac28b7994c247
z591ea4c91afd4cd84b483343cea3bc6185767268e6306bb03f5de6aaecd20f23cb06c2ad1c657f
zc761a4426bf68874bb28ed75dd4a634146bc91ac11f241aac403b1c1a9f9cb17042b73b16c1bf1
zd37ab88fd4f0827bbb704ed06c0488400b0620af76782480e09c2b637a8e1b1f411cb4605c668b
z2f8a89915c84d0c12a53d8a0d237e128efea99994bfb27513eb4c3279d08d23e2b5f9a48d6aa6b
z8b49ef024231211d0f734d9f6f1167d5f6dd74be70e3c85d0d52b42f36e6ba59d4ec06d1e2fb90
zac37d2c3213f25d69034d465b6a08f182cfe02d07f78ec407bf3b870818c9f51cb9d49f858d807
zac5dfde3b1ac4ce325597bf53f890974b396a7e288575c85e6138956a63a7bdfaca0da48413b0a
z270e7f5f19376eb8d50988a7c8c7a5a4a2b8da9707cc74331766edd94fc4aea9d9a393326f3b20
zc9658454ab28380361e649e666ab6e86cfa914391a10fd862b31aa8ffeff2283c32961dcd76b6b
z777095b67f4d443e27327fae590f62378e0c2212b51b17c08ca6e0859ca7213d71fea84ad90de2
z96984ecabf429190eb039bfc1cda5193c2d3b1bf2ae9ef0888b1bebce5a35189e6d3c0b39e476c
zabbac06f9af8319eed7c1753edc2d2e7e867a30faf2d02800aa7bd8208375a86ec345d56b80fcb
z46c385a7fa3b98cadc3229c3fcca6791bc53e33b7126aa6f194a1f5370aabc840123ce60051615
z2604b9ed011cfb6fa48bbff0723335d7129d1147372206c823d171cd9aa660a3a9e2720d6ac258
z885477497bbb8509c5b28d9d3112fb7caa56edb1a7170b33496eb9359befe9ba768fbc23222125
zd6d78d8080459ba30e92d1932543f237024bb3155bca7ceccb5d298a458b477f9296436bde1319
z842a7c2e2f6509b43b293eeac8449e21e3d5666d26ff2c44a94298d5b1672d4c6c8a8859eb9194
z807ee11cbf7919b30b2736d6f93c418d95c80cf029a83b45d590d6b56f740b8b285d845d14a019
z328fb2f6fa17f0132f24f30757f59e15324321b4644b1d649b79f3df47ee8596c3868c94054afe
zd284511a63ed6580815612b9679ffb0b86d9f55315c46ed560412774f55d8b654df2601a1feabf
z33571ff06a97bd8d5efef6e2ed7ca5c5ea28660cee20304ad3abdafc6fbe1eaddca4e609edbac2
zc33132cf62c2e85f0a226626d2768fd0987977fd43957dce9b5c55da02929116c2fce36a06cb36
z879693bf34af6713babb06e8e18f6a010a9fde73eca955727ea0ea855bb17c8f65a325278537ce
z79e480a23da3d05fa1014061203c6ed5d05c3cd8983058d75fee814eee030c7705c38aa6c059dd
zefa47f22bc6a74fa7ada8966932a7d4abf997c613d69468222dca44fa3ee4ad13c39e18744a51f
z677d8cf3bf2afd73ee4bce6f29c594faf050c14168585cad4d4e1863d3454827ddccfbaf5c170a
z5abe5124b69be848ab5ca1624ba3bb43c8c9ca4c402cabc4347f2325191677c2e0a3f9a5c19183
zd131acd6a74c2709ee120d404244f0e417a599e4ed68fa24dfafbac9cbfd4f09a18940200e985b
zf70a688c3384c4b51f6db899aaee9a56955d9fdaac5f6582f000a0586fd1a270c4ed2dc40136ab
z703771ebe2cee47ada16b952c722db7fd5d89ef82a75a3acbe43a6dc9912f812341fffa0f88464
z6239c6e41401d4070e5b4805580493e05ac56289b4322c71777e2559e9412b24e3490f92d25bd1
z81b610a001b15d5133ae328eb7a668d2bf33dc93178ee638665887efd00a0cf507e31eccc85035
zee83699add41aa5c947abfd1bf702f9aa05073c0c26e036df7208870a6a9c48613cd5a7a4fb2c7
z3f1a481c107f653ea6916db3f99dc2ea897ec44cac4a12603c0cee182412a635fc29f462b6e02b
zefbad33397de36597f791154fe6102a15e58b0043ee127c9455651d1a9eb23d0091d52f0b24b30
z748a988bd6d2b5f7e1f9aefab46443a76768d43a6694d3380caba61630ff631c734aa844d27f88
zfb134f82fcb93edc674add2f6f651f40d9fafdecd5636789feb55a0adb9f1f7865a0f60cb44266
za4d503645307db85782e87854924b302203eda87b4183df2c1bd6aa146a2ecd8e4926371af84f9
z078219cf8ba7613d6056465f5ccaed13f10948ec40d96fa32661ca0a4664f757332d3e71626830
zd7c930733a4867b803a4eb5ab33527da616d95a9057c3965fd21920459639a0b7c8a26d6448488
z11e9a0dc2eafa5096f618f483db5bf9dfdd86aeda6f654129ed057fa28d341df2f792a8cfc708d
z6a3de75352b42875891e8e43373370de128e567ef193547828f48656e6818903899c89fa238ef5
z7d339626e9aedf28127233e335ae3a9a27561d4557cc2e0f6ef406428c26ca1a38821ce709ec0e
zc5d07e1075736156421aed33ca813ba5fe523ae7eaca04cbdc195f37bbffd80507302836f99db1
zc1552bd204f70aacc6e91e0a57ef045dfdfb4d3eb2e03ba3fb615e91c297bb90dca008d7bcac14
z39fe7520b7edb0f4641f459252147aa24ba4891c4359301a6c6e6713ac482d1024489e2afab1f9
z5190d9afcd784ec463e6f7d35af661f2349a2ec9fe5f8757cf854b68eea84da29a2744ceafd3d2
z3f279b99f8bf1705e1a3b88d5bffd60f34a35f8cf45452fb9d96c8bfba13a96236356eb1b1a7a8
z50080b4e817eef042251a17ca25beac2cf0edcf50dee1e77ce141ac8992e3e0939568d45401a88
zb823ad7958fa48116380fc16cc5822749549e9fee721e603a41dd4eca000ab0e543cadc3faef30
z7079bc590ac83d1879b7f90527ca246698bb13d70ed80f6acd9f630c3160fc4514cd3727b30a57
z98e62c4e226b8bd59b4fc2ed26c754a34aec3cad5796d3ed383c7730d4f55536316bb5efabbf2a
ze3169b0eae88e7e8cc0083a31e938272a0bb18d93c912ce619ac8ffd8b986e673479e6e5c99bf8
z33d70dc236157698a78f6dd9dea7dba35625ad4619047e529e76f9a1f0ad041ea2c1e8a00a2c71
zb31f69ffbf11afdbcfb11d8e67d8101aca00f11fe3a3a44a38a79aa7fd9cd860ca9193d06a2df6
za0ffb8619b8b88ba0a9d47507bab97436523c33d00f550d5b62654e25593952e61e1b49ff7d0f4
za8fa3a772307bf723048693d9e689f7b20ee6add6757e3fdc974ecfb419218024406402b217f03
za23b43e8f85a3ca4475ba6e0bec42c235d7d2ceeed6eb2c1565b0370515beed81f7439fa2c458e
z94607eaf227a611f7ab80dc3f7fee5ab5581e6019af512ac2eaf34d8f48fc35f625924358f4f67
z512946d0082638ad49aab50cc29603a0a9fd5b8dad1cc5fa4fa6402b7dd15ef9fb75c8d18cec6c
z4c1c3d95f6a4d2de3f026b6aeb7cefe52e664e9674469f0cae779927c187a3f2b7d9db3c4c8c38
zdfb6e29095a63d4918cb7755d03dae587d34add091c70e6ebbcec6880c30b2605245e18cd1f6d6
ze0d45d1c73e60eb5d2f4cea3560be55f779fd136f867b7c7340129b17ed91764c6c2fbd1dcf693
z3b3ed4bef6fa68d3d29c9ae07b039c30210c00f2a5ff938728760720c74f07306a5fe44f73b662
zacc90325e1199dc57089cd35d17f23732e15865d68425bba4d250935faff7ce609dd8a0ef472b3
za933a9170a994a9d7157c5d5925eb4938468ead6a34da1c68b6d53416588640bfb4315046fc669
z87f8d040e60ff0422d1d84d43916f61c11e912ea007c41187fec7cfe543cb54ec8a7f49d4b98d0
zb24e93976b5769f3839bb7f761cdba374c043b1984b277504abb814b69352332b4c55ae44e4d43
zd56371990abb217297df54a73ee0db9e25f7961de146b8d054abd49f2d15a1a0ccaec0f4d92136
z58dd969b1566080851d4957b42ba95359d35c21ee96e458ac2d3882dac48eecd6ac1dfa78a682a
zef743a4c642fb17a346530cc3157ca62c6d39e029d2f5df36bd3f11616a29c6d752672b8f62451
z710f1b663edeef19fd7e8b01cd53c7c006d91d91e2a780302ccd7de6fc778ffca169e79aeb8f36
z6a500d614d47b11ab2af0a566f8fcdb4ce59726f50257e46222e5b6c668684f278dc344251924b
z4a58159b71fa6f51395d46e5b1df73f81353187179bdfa18f872e9b0cac454f48ab0fcb802e649
z56b3cfe8129ca970fd0bc75aeaa240bd6723f9f9babebcdc5d6ddaaf1e7293a111c474fe5d40ae
z8a0c68f9c2eb7172fcaedac04678cb6419a476c76219f6e57e3f2021dfc2048e90f881a1189666
z703cb3f6c7d8308badd97278e7ede5e96b09da603690fddf4d2b0dba9a52e584f799fc271f6890
z19a4c55a0cef23802b8cede2be43cb6158e6d9d72cda48884a9ad3a74094396fd797e376ebdd9c
z7464bbddab0461b5e5dcd8415cfd300d517a730675df64ec256c117a8c651e72263925b9a347d1
z14c4feb4d14e2ed89122360931e5249ee6a8b630a175739919761b3633877ed02506143fb2afcb
zcfea6811e8a516e5ee7ca36b68eba497a0f97a65112926611add65c5e15d33cc5b24cd47768b82
zb9dc140e09b088d4b291b20eb30903a03840212d1fbe296ddd8425c592b282625b011345263f52
z5d7864254c00bbef14d2055347bc59b0446b54a5f8104d57d1cac8997b2cb945247661b33f6d32
z3cb4148bf76c1443499d9a0d36a70c5be57bf1e972ec1a14040e773587429d074719a111045a27
zeb83af78a0d9caa82f8115d064937f3a98240a3a66e7e35b38e669fa150edf145a9845387baa6b
z6d8272397f130a21750a7f834225838256383c46a5c740a7e337c0244ade8f3fd1df72fdc94dc1
z63e280ef931a6b352b6bb494b7d32f69c717079d5bbda20964c5eb7c9017b29f6a5979c8052353
ze9b498cef00bc2785190c03760ca950ff659280a4ecf6eb70a67c2218d51c29a5bb325d8574e51
z2f8771703b559534501d43c3d2bab6b766c32a79eb4f2e361e5c39af13bd4d9d007b069a468b4a
zf3a053e68d517179e728696b4c9a9ddc3f53c6709ebefa9e730a252999cf5826d654dece9d1009
z92e73bf90a1474c7f5928b6b66a3779977fca1a5d9ff7cdcac942f776fcf1a71fa5c7ff22738d6
z296c5d6ad4426cadf9ba19497f198f8b5881bb9797db410611927a4a3c816d4e881a9baea49ee4
z763a2a07a7c5eb3f2a23765e788756d2c1ab4a83d3ce23b0355effa7332d836cd1ce119b7fa2eb
z4a176f446471a7ef9baf989e0f41eca34710601c3f444bba72f03f32d48f3075bbb75cff7fb13d
z4ad413ba2eaf64dc38876b8e717841de43d259c082dfc8b3b133f4ec276f485b58ae8ca03951ae
z02cd8c869d80bc6f22cb55c04384051420e9ef992e2790916ad4a76c4c3b5ba3630120a1ec1beb
z01cf8997038a5f51497d465c4ac284292706ddc55843dc4aab365bda0748ab3227fb46473463bd
z71d9d0693c942bb0cecb9f06e89baf57ad3dda72033ebfd6b628af78e64058ed799df66120105c
z1a3091f007f5c609847970308cbdc706d8b6ffd61c25d92738a9850ab7aba6c75b4bff39bf5892
z1e3344305e027114c4cef2f364ce0967cd2cbdc712db6d7305b07af7a2b83ce76dbf7a490b5b73
z0e49a37c00a3a6b4076cda62721e30605ec766f78cd74f6b1b2f911623624f3bc38763a113533f
zb6a6242bc12f7482cc36c8ce41f5dbab0ded5ab931cbbfc61f6df34f40831eae0d0a4c206f3d88
zb32749f55576010be139be466746c82c5187f61a5244b3aa98b05fd8a8bffce94bf4bbd6959c86
z689cc1901f3cb8ee3e1e62022c06572c9d6028522b2d45610260a922b9d1b237861be98d70d337
zd4852aadd6de8253064b18d01fd85afe30cffdb771bb5f5229ee0f903897833a5f28dd64575c50
zd93b3e20e1cf63718577d25e1eaa4c0102b0337c87ecd91857a52272ffbc6e47477640c24fd025
z3080327ce8f5784a5d9f3532c22f7f6a947b7fd2b68fa9aa9690e1721882ca27a49feda47b30d2
z3d737acbc3ed6d519999f0e67fecc480a20e4c222c9d53f265ea5ec3b92088574182386e43ce23
zae37c4df4b263b3ea1b98bd8b1af4c541c3a8082c0f127f1e10b4926de237e3d9eab5655eb8484
z26fa3da8cf6568f864e139a8e720a1018db5dfee10e9a6ae93bf5b1f99bfd1fa45520dc72d6795
z34f1fe1f3719418daed192a4bcf1afa6e2b8d2ed96c9de6e3ec64d5f8406d3fa8164390a8db660
z8790343b8c4cccea962981fc075f63f9c70b7072867e1da1bb2691cfb14612a721550ca38ab01e
z89404fd5b9bb61811431fb32eb0358cc4d8f9922f9f393c0e9ca28c59cb6ca233f3d5c14d8cbd1
z047fab162c4564871c0fe90114ade0763c35e7a859a1fedcab5a1800ab3141417628084727f180
za2cb3cd225ca74a8eb6364b94b11e84496193e29e33526802ea4133962c5283f8bbfd675624c41
z1f747ad6d6b52bae30ce5d96b8b6160ebecef0308c234e697158c474d2650db598a02871605189
z43bcf333b1b4500bb2adff215f137a7796ee0c53b32493e703267a8ce0a85e032dd23b642dd4ec
zfa1b221bdb075cf029f9847e069addbd7f86d609faf6cf3664bf89feacf3e7d1c6c9fb5f88ed14
zf58312cd13e2443d4d8d50590ece6057f01c95bc5ea84203d18c916ec33f5f9e4fbdf948d401d5
z06c4434fa9d7186a8e20fa2c62324e4595e3cb5f35922b3886bd01c9ffab574c636093cdcd205c
z1a42f1d5c0f4b13539e05523af316e59d61ad202e94d1d57a210ba9179216a0afb80889cd3b67e
z1b6265e3ea9ab8315c0a4088b1ce89eed8665d4ab16901b200ecd01094c74a40f72fc4ff5db018
zb0f96602c1612aa160f28c7dee61b3a638ad2f12788ad07f1798e62d23502c11fe43cc7122bf7e
zce288d358ca336893e47d689ca59caf239c62e33e00b76ce6a0b6694cb25603cd44f931bd98a2e
zaf2dc317de1f8b52c51f11418964aa03fc977057c40b04aaaa65a637d61d18059fed7a762c1973
z5cbcc8043f037c038bdc53ace605bb1a7497fe042af5627240f5319369386947b3ae69b90706e7
z47e8b3af2cb8aa2577700d51624123c0c498579f17236617be86a95f9764340f1833da3a74b30e
z8d7cc718ce89466f9254c5d0556bc4e62f0d2a1fbac436ee63fed9885af9a5f01caba6cb6c285d
z339a466c23b8cc6dac4b661fcaab0a3e49930b8cbc1969477633cd7fcb8a545ae519614d48c841
z3832d3adb5295ee6cdb631b7e6e7dd6643e93efd0b56a04d162153dd1c0422a843b2a6f2188d3f
zd851ea773b7f1e83fb504998ab4b75c9c6f9dc670763bfa0a063d54a0352dc1a91c0ddff1e3810
zc97a3c5b69f2c4c6c80a26a64521a2855de530efe701e5f3decc3bb97d0e6fc30c5ba4df0d3e51
zaf431be8e0e72ae2fbd0ea96d31c2b84f0ddf0c01bb581cdbeb954847478d2216d265efe869607
z4fd7fe017f86b032e518b0e66dcf5c4f87a7d7977602c96645acb099823abcf6835e7c1262b2d6
z44de3292264aca9bb9ed35813ece0da7ffd4613b88ef4f5830e90c510df9a68ffd2793dc531a72
za699f050dc9edd508281ac7b50560e78b91a16a81cb630e07090548f4c2bee21033b8341d2a6ea
z80ec12bf10a8e3cbda0aaf88b46d088706553e8744a594c594b7b888bbebb64352a20d167d7e6b
z16f4bbf346dcbaceecf9870a364e916bac6477b37f7552f2d40034139b93b5f9e7c05a04e77580
z906a6e3833a416322bc1caec3bc95f9f7bd92a99b9b899aea97ce8d3a2215cc33bc9741b0ecc29
zdd35417065aac19a3ef4493b11ee1dd6e8479a6d1ee37c9e2c6798c96757a3362011ac6ca4bece
z85fdadc2fae590637f944e26dd91df800cd3c8197d4492d28c007d228137d455e0227835225748
z12b97f01b2b58fa0f8c463606248946a7f11d6c0e8a95e2688ffcb79aae44b074eeea9c8192ef3
z87976a325b2e112ef6543bd58fd1240c35c7658eff6a458d4c9f9712f83b9dacaea3ddbaf015b0
z87963690e32b7ea8e9e10865467fffb2cf4bf8c323638e91a3369a9bce27ef49694b44bcd4148c
z9a5b4a38cc13838b5fe60661ad7f62ee64a3b7babd95418e64731ce23c97a4990bc01f9d69b578
zc9d0de46dc38e7085ec4deab9f86fd25d78a8189ce96dc2bdb2015c92b88a889db41ddbfede934
z7d11107091218e93e005216c4dd69af13639fc286714f33a0f11d598f38f6255509949898a09f1
z581675d1cb04a2316514a3b6b51443d3e06c508a1ad35c32d9ae89e9ed0ed427591c87185b85f9
z8a0c9ca19a815b81f0f8b02e5a730050c3b21beffe6edafa3ed4ea72604246137529fc351e305e
z09aaaee72e74af71668301322272883a602b6476c5b19d4089937ebc157d0fe9b9e1d9f30c73f0
zd1ddd9be561b9762329982377a1b8f1a00372f953ac3a196d0a28978ffa90769f9603081b009d6
z084fa1952ff7f97280eae961a5f724e2a095ca317a17906ba995f3070d9cb0e5246ff85ff2933d
za748e4b6f22f668954126fd8b94edb31e6eedd0061ce3a483b97cd799ab8e9675289b7149f9a5d
z9f9fa48e35e93513a1679c093664007addbe29219f585abad32b27169f95f79f10b6212a991457
zb229fbb2d6f538b86cd7cfed146475c192b8de32184e75cb1bbae8693821744b785cab465d3619
z9f052ee1e2b8aad6e9b8bd281d0cbe00d4060780cef76487ec151d6b918e04bb575b7be9a88b24
ze1f55b4f14f11a9b531aa44485f0214a0573f118e95b5e0fc23859985d5ec0e2c5951dee00e8dc
zb4d0ca07b900f4ebf1373c300be3660ee404f162d62f91585a3bde992e163c0ad02194e85553e2
z8c8d3c2778f8bc6958a5b99f28695305d1bb637327bd58bdaf51fe1fd79aeb0575da396e2ced02
z229997c06433cac53833711382b2bac11d0ef2bd3556c8df63c74891ca8dd75c8da6c5096b40ae
zae0024cc96f3e57d4a7b81698e7b21cdd0924d64027a643663e7d9e497ad32f21b448afc0d572f
z20daf5b759b2bd0f96859d397ad92840760d778428af4c50750eaa322ae24bf4544b5330e01038
z3248b67c3cd3c4f3949867d6d2f8cee3d464cee048deb6bb0ae482cdaeedef786a4d418b942b40
z178b242e89d87be1822280254f93326bd219b51e0e8a4df4a21978563b2e48f83a62e4274e56eb
z8345ef6c6a7327e306acbebd7a083ac8cc1bfe108d3e5925ebf662d5a3fd6f28862993a83abb9b
za12ecf2df0deac9dcafc666e9cd837a94fb1ab7e427ca9854028233beade6aa1c37c84bdf94183
zae7ba528b09bc7f30b7fcb9fb3a39791b449b3aa2b0d442db8ce411ee4dc29ca3ff53c824eee77
zc5d971fd5e2ef9bd4cd02f2ab1b944af8a0acae66d3e9aaab2d5c645b05780cea7db43901fa686
z9e37c0caa66c5411fe3c0996f1646fe082783fb085361c1cb9542d5d059ad4fca1ed9e854110ba
z856b851c1ec8b2b33b05860af43976413df66db388f43170ce7b3c083ccbae956650a68df5a4fa
z18d49c85566b2f433fdf8970b0d1ad252ff0c0c95e134bc06173abb8952b248645980454d45586
z7722848072d0730a0747e9aa5aaea986f95cef4734eede6cc2daa22703152b3163f53a369b1c8b
zf79cecf0a611e1512de2689a9669c10e254c4318d3b868b061a31c547cdeaeff1fb158a537fa7f
ze76ecce20c08898fc074dc6fab23581689917cdf9ed848105657e2bc8aa7f2f763131cb1fc3c00
z32f5af7dc2ad80969b9d2de55dcc257be70e1f73dd69393caa96de0ac72e5f6434baa8c53f9762
z8ad5b625ea63cd8a2de0729b93953c2f1511d52195cdc0cad0869fec587d0239514128cc84402c
z89baf0c3f7f1dcee0625fdfe8ab8bcc5a0fb98d60b8829ee7caa3927dc6c7d01fbbee3a255b5e2
z9e19eb4c73664fec3cc51a9e53bc9fb981b3cee785fcd88e23e749e895ae4d37062cda04b2813f
zd1a2881d12b5d6dba11f0a1cc66f2e81c209ce574d9b9e3a23a42f36dec9ef30dd05063bd8ff5e
z17f1ab3b012c5ef7adacb4c2b89f763983c573ccf8b2b6f43b67912392b644340d08f31d7d7b38
zb47e1aac56ba61ca5e3f599c8a28bf6ad16f1727999aeb215f0ef5d143d58e395abe8c551e000f
z45891a3249e881f15a15d8e9f0098794cd3f39a38ea0810e7df2e552be6e80a0e8e1dbf251d4db
zde93a8c2ca0ea4eb7232021be391056fbaccdf66600a86de697e86619915a17dcda011fb974307
z7696f7acb8948579fcfa8d1146843a69df86e24ba59f0c9e321508453bb42e23b70dd0ada43d66
zf8152982b739dc53512eefe0434d3edb6b89519a024447bb8e846554ee74aa9f44134bd97a31f8
ze788cf12c9014afcc254a8cfbb35726889fb2260061292a3d2df1027cd5b7e8f1ccedcadc72458
za4be71524b54d7060f5193b1500745e95e57c3ac252319845e8374acafe1e8d9c4de1282788eef
z92aff83a9499eb39176f6482974fea7b4c5e8eafb03163c37d16887cb7b48c05352419020eec6e
z4c8d705a62a098386b9937ec5f79c2e170a4e730edcdbf1bfa5f13f657314c997eb63b3b4aff5e
z5b916b26722959cc78caff6ee23fe2d9ffcb61be2738a22fe03e344cf8d962a94746520909910d
zabc0cd814bf44d6454664e7cafee404da6f01614aef97818a914fac90bfd14103b87d29bd0b38c
zb8742afe8ac26b6143057853458239f4b961d9680e579c89017aea5ec8f61b5961eeb06cb44b96
za19b4e44409b1105eac1d8ca6b06fdfabdd1fabe86ec09ce1542069cd8daa80b713127160b7b6c
z24ba878721942f35135aa7e0d0cf7ea73bde7c7186192c093ed9e7a058702c785665c195552d08
z4051d019be8521dbc2ed2a94bd25f3728ef895c951a54f5621cf66a8fb39125c078cf26b595f9c
zc406c1b4a64135e6aab1526656b8c863b1938e84d2e382c90db2f509c7d33bac35e4c67206ea27
zbbc25d20b6df1d634b47bebf2f3363696ddc0f1be3bbe9436da3ef0113b6ab92d28080ae017c5a
z360699d67ec7b0668bd1923a339f57e9a5d4ebd20e1e7c59831108b08162317bbc6a8d55b931c5
zd82331bfc29936762b021b64c95c65a3cb707d43a258f60803388685f661638bc9f55fde8273db
z9f3a3abde37af79ee62e39ff2a46adbab1509f820a3b639916e0699511e39046fcb5a92be83c94
zab0c6fe55f21f6f2a5204b09c3526fc0455282bb84a0ddb6189e33ab27279240e980720188a833
z95ed31c6f6f90c473ce6de6aa11bbd7abb90533883d4a3a27374c3dd9866918e2ce257d6fe5b93
z335780a0c85fb59e3c4e000bff5c975a09886859f6d09b46da747f88096d928fce10e85444ec85
zcb2fafcff8b3b25fd18b81380e344649d47fd11848f6aacba87819d44439fc3930c7716f62c7c6
z187a31b30ae0c2b50c9a0cd94c650e0fa3b27759e7054121f3d187a454f8cd24c6832df4d639d2
z8cb62072b4c46aeb3098e25c135f13593fe344a24f0da11e0009684220bdc83d216567a9e07167
zebe63d8787cc076ff0fe090150c5aa31c5ffccf09d8866a00234a177fe0fd04b39597b4a27def7
z002d9477430b2a2a7cc662f4bc32be3d41117c760ed37e9ae53644e2d9feb528a33764a1e11c08
z7965a7fe69bf2d5eb3ec8ced3ef7882eced76135c009881f6050bbe422cea5fdbc0af71306bf61
z71a2e7aefae740cb18db54d3c3179e38575900499bef86edac83d022d94a8b847125bc5e24713b
ze303399683b392daa5e2b11e243b9129f08e7b9f33a401a8d8efc275d126e739c181f401ca6bc9
z5f0fe7f585271200a032eee1901c60da7aa0b03304c9bc54813c6bc512bfae95848c0aab64f11c
z800d6ec20f199e0629d5ae436f4ed2a77b441a09092fbfb31fe126aa8bfe8d26793777edf48431
zff2c15c9fa3ce63def1c430610d6d97fe51a8ff5fa0b8fd008650b45156a3dbf05940481a2f31a
z034ac89eb36b008a4a1e216a4b61d5b8fb85f6cc12101f7aae720d2b91d55ac215b093792f9338
z58643580a5d0e0b0606c40804f962512016ac8a8d8b54ed5c2a06053e7205f31605d52c891e4f0
z03f1d306f2cdf87cd038809cc57ed4a8c27b418e6d32069d450fb4039c43ad6184bc246e6811ce
z1f8f7322526a47a29442964f0a0fe1fff29e8159163403df3357dd8f9635ac91b4bf6d3b93c3f5
z3d15e6fd3f51071e2c00a8d6cb980686bcbc2b74e14c9275415b3afbd811452e140df2a8e812b7
z347d95e53a8d73b1e22325b01c569736c77d9df25085c55dcecf9e51c3c33e65bb9b73651bd11f
z50334c055bee315bc6c88e8e76409d032a708c4cea4836b59c556edcbd074f0b0bda41c52de0f6
z702a2b60c73217d0ced6a500718e51f5381fb78df6abeca85dad4478a4e073c583be1368cc9975
z8e3a891d704ab283a2e76d61dce8f0a948ce28b898d9997f69a4f21514c78632ad2a22374bf7c8
zf137a4c0f717401d5b7c7c866722ac154ff438da5c87c2d27f42445aac6cdd86bc5a121f355784
zae4fd2ed6e967722340ef6c2582ceb211982b3ab12b4707467d2396c1e2c047e5a4c2f98c2af11
z527b0c3bc3171ac206adbfca0d5a1a494cf14589011e41ec5c94f304ae930f63fa0f683ab86eeb
z144f88291abeaa7526b640a188b534dd355b508ec16ea4503ed0d0d1a6cf23d07ebe2ffa15b365
z1a0e81c54bfad1712c8ecd6972cd3b22c6fa155c742e2178836a3373268aaae2892502e4bf980f
ze4a8332d1013e921e667bfcf096fd307ea0bf0b6daee9870410df484b76e649234e2a9d5b54322
z13d2249e3d59a519628bfe043d2835993f46dba3272e2d8724bb9a2ce9d42824f99cb17f80c52c
z107e7d905aee710d422fb09dc188772db95f978de660fb93ffd576af20af8a29cb30818662a5c6
z72ed73370aae629ba1d07f158305f52231012d41393289b8d500403418e2c545f95e359f419b2e
z473f55b025a67ee560b7515997054ca49b5f0b79d8912cb04324aec2b1cb3e16dab35710447963
zb3c01656cf02bc2b9b06ac3fee7520230b4825ca81dc0740c0152413e9924b888897c5d10106a5
z08130f86ef92be2bb155ed2006b5c6c449c6a66061a9fd083cb4af612d949685eb47a0a002da94
z1dc0d20e32a3380d0237c41706ccd02481cd98da275eb06053249a29f4d61b262937af4188b8c3
z94c2e1f7253e1e86eb60dba8b90fcb210d166f3ce7b8d95cc8558b1bc730c8d04e884d573c6d71
z929d6df8d6fcf935362f56f4fceafce45dba6b9b886c4c48eecf425151c594f4f78013c3255847
z18d3efb0d3b8388a07beda48406c5554af3bbde6438ab45d539c3a3f8b7978363352030bb5993a
z715f01897cc0bc57d0d12749f18995bfa97b22ebd6396100f2d3599fd619bb1a5dd4c1bac2dd73
z3481f9200ebf4908b62383c0d11d03566238d976398189b9ec7830aeab7860b9d8e1a166cd0b24
z890cdd247c4a04f9122f02f951b03a5d00f0d188128c6bc333949e24c14a4de55576fdacf4d422
z2cf860f4d035ed5b67cec10bade8a8ae5c25ab75acf777fc2febf03b955ca4f777db1c86ba37ed
z363480e1491e0b52773e433a20a3c659f23353d12a402bdc563958a3105a5c678a06d6277553a6
z04c226ea60082ffc4a6a924dec6f10ff5eff86217ef74671daa8d0e3ace0dac64f32e55c346758
zf3deb2349f60b1fddf8f405cc9595bd1f364bd64e0d3c50b162983a83c9c3562f172e31a28ecd8
z49feb1662e64a6fa4e9d2e1ce93ed7491ddc034c947cb54fe1f6696a43cf05cc61ea264d535a09
z86d9e72d9283ac6327e12df354a7c3753a770baa037bec7ef38e1bd097f5aa184524ae51112644
z9a993de3310cae7ec0e024345f3407ec67fd7f8c3514ee66150484b3be6c9f5b27c73378ce5610
za410c74599ffb01fca994893f64459a022bd4c9d7cafb59bb9f60c488a9ea90f5c6a814e1ed2ab
z5dbd6cc4cf143d2058753080b8d1466fb00aacb096a6e18035f7f40beecc5de475d745547bda53
z069bde73861795a4c4d0ac39ca938d4bdc0edf5597163d05a2fe6cf7c4fe3f2c6a3ba11800bb9a
z718d1ace6d31116a98182b3edd3d29603e1475d6e75d2853e04a1d30c7435375b7765082b17cc1
zf8d0e404648c50a8c4c4f96320be9b8cd2cbce5d8dda72c6204e2bc73c9aaa5e87798d0b56168d
z9e389326edec9be1436991a797ec83e9cf3226cf512a82aa132a1634760020222b4bf4d081dba0
z6128a9606aee47ade22fe2b208b90a6bcdea1b4e2d6d7088d5f94530d1b01a761b5a490ab1f8ea
ze3641dad049a729f00034b3fc378ba3fdb756fa79573f7e35a219ad2671cc570d9c15944a0833a
zb10f5d1b197ad1257ed28ff995168025bd254c2636f2d8b71452fe10852c239ec71d597e6a5314
zcd0973a3639e48cd87362226c9ef65b08b7b78df2ceb658f2af7aa45a6724ae7941dd85713d806
zfbd33fe55b81186a89ec57fe54ea4a2513fd7c83e86f14517dd3cbab3c183b232400da66e45082
za68dc1c4deae156f4602b3a35b04546fd93377b9a8c1482b4ef47adc07318ba16d405127743c19
zb47ce5230413d3242c5b88dca1a226a162bef1a5788e04beb78b6a6ea2fa9ec3286f49f3136e8d
z476ca57a6686a7d5f7b14128355ff84b556e81bb5ef383b70ae1dba0ba90b8956341ee42a300dc
z87e93723e6acc431cc60a42ba7204a3dfde9bd154344de38f4c98cd9691164ed7ad0900ff7e1f4
zc765bf563e2dd75d134bdb858bd7832a58515b59551d88df5dfc139eea155571454bdc4d7f1773
z7f37c0448579315a6625a1c2699d703e7f6f373c4fa5b8a76affb8d8338c8e205bc2ae732c1926
z7f75115041b743c306c016b1fc8c0ba0da424f2ff60f2583908db20f06b5ad94165d80e4fd9d1e
z9f31c8fd468a4fb7f245b63611b3145dca543eb3ff1405a56d7ab26851967b11e04884fae31531
z6c76421304b8f988bfc7fc5f2ad66a7f9dfdf965863cbc735128856e00cbde954659121b10fb1f
z52829bb6382c725191c0018b6c8515fb9fa9464d9594495bfa7772c0bdef4cb595c6453a774f5a
z6a232fcea34a8d6cff9920698a6ae3d166f5081696837fdce1264e52f0d98c863c77dbddd0cce5
z59b22d2425f19edea6893e4004f41b5c0c085c1fcd6c3d26b9c5687b804bf14a09f4c1301ab01a
z201090275742e2b84b21500a235e6ba43894d465537e091c45e8a25251f33f1fff5fcc31ad24f3
zbbd3f24004d1957506aa81b91ad556ee9926260d39662174137be0c18b5d499bcaf76d330ae02c
zef9962eb2fcb7116a99d0e24864dfe39784d56ab0fcf5a56c5def65dc5c6e95561ab85c1b41a77
z31f43e6cbbf3d7e8dac56175d4779da86cd4227a9dc98b8b8936474f24b4800c04926bd8d082c7
zae22e14104aada1c3b925db1b247a0959f71d6fe8751fd1310fe25392e27f1e7e0c277304106e5
z2dc8d52950fc0ef8e554db46b522c21975beb887369569ad5d351b264a8043df8670267955a632
z3ffbe9d3853ab7fbc1e1932a9800447fc46af22b6053cec367873214501769e24ccab456b66b69
z32bd3c9497e8de75526c9c0b1bb59a746f385c9d59cac03c0b2f96e6dcb9d27275132a20005968
zbf0a33ab2f8c67ce936dc269ad31d96de65b92422464b4908b7c24e2fc9be9c16129956f42f844
z5473f3a53659c801e80c595cff9dff5498196172660a50420e0f203b8f3bcbbf6ccfaaa93ead6b
z75bd42df05dc43308e8063be2afc6b22734fe10b5c669946e908f1e2ef12fde486273843146964
zc7a40b0ab83192e2a90338d93c79535927b4a704ab25fa9bef08558b89a4fc3805047831d5dd6c
ze2622df54c150fd20d5656826ef01fc40bef930a0d0adf62dd1c0697d07c30bfc1eac259a055cc
z8ecf835825f6aa3c19ae47241ccdd0f4190a03374ad2afaeca32c54dfa0e7a24b0df0e67dfb599
z7c61e9e167587c2ef36756229040c713cc50b9511d0743cf5835915e48313d8b9b9e44c11e53ad
z5b6fd0b82e6ebcf6a288641abe46e8fcd7e59915fa593b1e5a9e830c805bb51747bcb61985aba2
z25c7acf011bca4ebe89dd7d3c4717b4cef4cba3edf1df862b6d7457033c6597e09872364ea0bff
z5e9732fa07da8debf37525131af4315efd701b1007e1add9feb7376062e124cd7b407fdd55bbef
z72e9199c48ea7e080b2be531f664d6a0eebb5189a0ecee935be656443135a40b14f75f5464fbbb
z75fb4f06f1cb89c3fe90c95303b2c3f3be54831421746c60e5020511357d1198a8bbf8987004b0
zf707a86ce5a58774c4b63234af6401a81171b45c1e16e3f748418c5366af9ed7b588a4da1a72b1
zc27017447992e4dc8d0446bc535c4c02cf90e1102f6b52a349448aceb0abff6c1a2bf899e85ed5
z7832b899e231282acf5268084d2633b560fcd3703bb8eb591ce750ad6d8d419b11675cdebc5656
zbbbccba8dc5437be4274b38c3e0290b2ebcfb76a0ea2d4997509dc8754d9bb18f165ab7883a216
z317c5b7de1f25c2bd9c9d622673235820b64a888bdaf69dc1f5aeb749dd20b4e5666f8e2d7134b
z9b81b87d2c4b8b290524028d229588b96f6cf7107cc9d105f940cc50b6be7603204abb1e6cef9c
z35cf12612156e7c49ffa9ab9eb4a9d5ebd0d9b5726b83070a487262c664e250f2b47daab03b07f
z171e738e23722a3e95393e83ade0acee3532a4a515bf8b75cb11b6151b359a93f1abfa503b24cd
z623ceb867e017d8e07c059d8a5a8860ec7ef0cde634fe10de2416c15f8a71cefb9c2e72952c6ca
z8d026683ccb144de6c33284bbdb190dd2c3a281d3c969862431dd1900a730afbffa532cca076ba
zc5b49d3684f4c7f4e7d1fe73231211d7c70e6c50252cad3248189cb10eae4ff7a97db5bf7e1d2f
z24f037f4aa363521e9d4d28315c11b102a21e658006109b138d94d32bd0f6a80604fb7d2f9fc6e
zd16b562ebbf4e296856c80b1b3d55371d56b54c8541e519616e93261883b2675affa5c551a051f
ze347f0978e97faf314f8e09bc179f71a321b46707ee374862f594854e98793c50b877a297efefe
z579c65f169890b3052ec2ec4bd0aef9a83a0feb8bc4bbc6407b6326024f32f4e30631a504f1413
z8886dac6424a1a83d6a4afb8a2f84d8fe3318edefe282d521fa73a4f31d1898c4d84e5c66af3d2
zd057acfcf25657d9481669bf0329abe84da5dc318144113da08bb53f8ccf10a4b82bb958cb3816
za76f3359e0607d7cc5705cc3b1b8f435c6129d926f1565c97d6ef5fe0b083cbd8984215aceb33b
zc91d885686a34f6a144483180a547c58c828121407e3d2b1519914c15447360d84d21b989151cf
z7e2de17206548a4cf7b3153e0666c7c364dc7449d98f3c28798fd8ddc2dbd697c10cd8a08545a6
z981413d686f50441f1db2d49412702d280ec10ca9546e3a4d49e522c21c62f91a4a11f91b250d4
zcd3f319556e108d7d5fe5a2a4f1da81c0b901ab0e2f26ab365a3f2c7d93400e0dc85d5b48cfa21
z0a8f137a8189ff9737b95f21728bc82d6fa84a232c0d7717f84199deb06fc7d872b547d9edb3ed
z296e8b8e0b6be8dc5e56f5762c2307299e327a2e2dbd77ab7fd9ab7ab2925a07aa7ab10930cb5a
z11bedb677b1beb7f01ddd6ac0ca214a2e9fd1c825ce17f5ae7458423c715aa50bb2b6f3306050a
z65b541faef3b61bb98e01cdee481621e576c014fc0246774df2ad47f3c60ce7915a802377cf9ae
z4b08de36c4c168c94aaf253a123b501c0cd4105adc735bbb86bbaea7bb1987e041c2b9e5739985
z53a898f85a85a659cb14efe2724642075ae26c4473c6f15f18249dd2660a275e1e5ace18bc5f61
zd16e77feba7a8dd2dddfcea42347dbc54ef09c5eb8db9734fa19eb98d2f9ab9df012b73e740d5d
za7cb382b34f756b6da47d090ac6ee873c1787e53140df8e956a3596acb1b29fc0bb72eb7ffca05
zc1a40d24709be36ec506a16a34b83445c6870f7449a95355bfa122d454446327790f2a16ce3fcc
z677c4d3bb353e354dd687e603d02016764a7a996529f57a520e8c2ac3bb8c013952331965797cd
zfcac92830e8142e676f6075f8bfaca54efdd4b4414394e6fd5e3d152a34b48d521fcb5a3946b3d
zff42880d368f7b3e72a6a709c65ca4ce6aa276ec8c
`end_protected_0in
`else
`ifdef MODEL_TECH
`include "qvl_gigabit_ethernet_xgmii_logic.mti.svp"
`endif // MODEL_TECH
`endif // encrypted_0in
