`ifdef encrypted_0in
`protected_0in
ze74c34e226135848fe16db9ffd31815111b6d7fb642c521a3f628cf6da949865580b22efd062a7
ze90adae0e65e66a2c36a587d0a790699166942afea5fb71013f1cbb0be1cfe63975264f8dfa09e
zedee295aa41338d563976cd45ef779be1aadcc43f3866a5636f201c3c0e6f2b2b9b6dcd115781d
z9dbe6e0d28ae18919333fe43f18bcb318675bcb028d58970a6d57d633808d9f444a82aa62b4207
z749d58c9b3ff73e7ce028d31af66fd2846235b3438d5809aad1e42b8b2cbf7e6d520a2896a7109
z8c2b2c6e6262a4b40c3ebaf1514dbcd5b996eff2c5bc6aba1b2d745d2b14be60c6120c68837818
zc7ecc4c0e897c040dea618c92d39c90f3c000a6ce7b7ab3c718219d6d913f77320f749c40619e6
zb2f58d9466f35ea1d5ad718ac92a1a3b3b5aaf29cabd74b2cf4f3f2abab35e7063ef1db739df6a
z6107f7e8da614b4ca1966deb463cfe4e0fa56c4d18bca43cbe1f2631b9285c727030a7a4a55e2e
ze7d36649e0fbad22bc1c88b4f1c2df308ec006b358c1e1fdc0b1c264b9116a48a8f31504be627f
zb59c6855b504b8ca79a26bf58ab7a3ed29ba5401ab04acf2ce58baa395b722729d370131241743
zbc93d4c833e0c768e676e18ba0daf46196cdbf196b4db7d527f4fd34cef24989862b25a2884551
zac1d43d2a2ae0d5a11c70ed137a6aac05da52a98ec03a9077609b1dd81b09dd469f0f4c55ec874
z2d07887b2f0b55dac595d3d6ca31e1a9918f409d79c217feb108efbc75e9cd1d9d5310d3568acb
z65b0aa1f74b5ef86b53b874bfb44109640e479f3485aa4ca33a890e41b2dd86e68e75a1e00b369
z93e57b6b6df06266d8dc46ca1cd9f3f448f41a3543bceca85d040111cfa0ade839dbdf1cab2a17
zbf9abbeed57ce505a8b2d9817bee6807fc51c63e85beb6d5e55f56ca7663837becb01f7d360cab
z87d2166b70be29794a849fa18537aac25dab8a963d8892652d4c8d08409227be9f12ddc88ee795
zd902a857af5a1d8b1a4e87206909bb6d90ea645bd8b08f44bb1f23621e5e85fd0f700e1c56b2fa
z050c8afa93de9a3093b0183529913cbcf86aeb18ad960583d165c7a3dc5e99c573e7ea881fc9cb
z72c296ccd0830742f9af3e831fbb591b4fe9d63eb7c0f454f7ed9fe7560db196c2db868cfa27b9
za3fa467de62e4a090b19b63e334f61d546208fcef34f09ad549e19d690fad763096c3b672531bf
z23e3e74e7765b4da96960f490ceb47beaa039cc8c98eedf0657d21a561c88af16f4b815c6e906c
z748a5178a44ffe4963a8dd293591881a7ddcc7394eec365947ae4a40273cd6e73790376b4f145c
z9f35dcd46e72b44b900335657fe6dec4346831deade8b543e50d226024afe17d152a97c48b502b
z1858379b436bb4eca9ba22e88bc23f1083d246c4a6aab79fd2e5c93c5ffb38a72d31a590555b49
zb99c38d75deda6b98d05e998ba87a3bbc1ca1c43192a5afbb40fb6e78987b0ed608038f5a2397a
zd034a6e36b9b797e8dd346fbbc24f7611e8fe9bebcadcf3aebfbb1c24a3eb86200ce6123cbf5e3
z9e2aa856d077a5ddc71aca0744188c948a9d52effae73da7448be3186d69523abd121a9c927bf3
z8c9c3bc4b8cd622a4c3aca9fdc72de04f4abd1dcc4f4ca60ef588710e34b609bb1daa16ec67f08
ze83faa6a7ade4741f00aa66e279835b89967640a88210d001d9e44c0413b6f17399948b5b5fe17
z11e7cc58629f9226f97497f3dd760763cf5d58eee1fef59f8d85d44a331d090ee4658337a8bab5
z7ce9cdea10ede16902284009c38a6e4dc043b3f06a1577dc7a8f48d47a6d48fd2b5f1752b87fac
zb5fcd1675f376246a73456e2449e7c72679db357ba8ae96f97172bb2f30ecbece0ce338aa8d086
z26ad39b92f29690d3b979e3b21ab067067ba360410d8a35504c71c7f2770d3d48f3e2a5d5cddcc
z3f7dae940df1ac4473a8e246d28d413773e3af144c78ae029f2819798b5a614aa9b1a61c265ecf
z78577b1308ef69677ce12d6dc433c226fdbc68d827f9a8dad618c9d75cd1bccd439d9ac7d8e8d9
zca62be0cf5de17069b8af1a2206ae5b6d1057451b6dad6b67745d87d432ac76673d6837f6c0403
z4d79da7e87903aacce06c5e6901b6449120742e67bc357afb4c217f57b20ec1198cc5a933df48e
z85f6d892f518ac2d335313bec3d99b2d30a5aee0e049ec9d9cc3f8cf720ed401cebba8919b5899
zd77ed1950b068c6d806f26291299c5e97aeba32a2f68a6105616e759fb236464c50d54ead65df4
z24a9e0e510b26a067f289be43bf3cd49b318bbf5b1b54c1115a6c7d8a723afc48e6a025d830016
z1b6117ac65e36bd079fd7b069e8eed9376e915c9d9f42d39c9ccbe2df9ef67161cc16471e358f6
z6917c2082a9f2e9523708bd26ff30576b9e0a442a4792c677508b81b4ff33b9840d49777a79797
z20ca260184b165576ba5de02e10587d62d03548c50d591a985ef818334be994ad3dd5f04e6424a
zcc5b4c10dc7138aac39649a277041c4cc297d2f74cb855b43e3cbaa4ab344effdfa860632ba1ba
ze98af6a3833dcdc9960bb766f98b91561d899491174d1d0d2e8afdc38cfaed2244ced1f43242a5
zbed8cc5bc18b0dfb781745db75fc07a3b9ecc333c71e2dac92ecbe078c533beae4fc775897e382
zc3ab2551c0489ca35b39878e84881de9486a6e371cd373fba110975446d0dac4cd540ea6baab71
z0fccaf719cd516d4e232236537f83429474b9d73de315498f7cbe4d5ca07db4fd75e4233780af9
z70f511ce9bfcfaf0d3c2a061d6eda0a74d03159f3465963add84ed825761d2c43934617879c36a
zda9c22f733943a5f434acbd778d8e67adc67c16e432c1fcb189743cbe6bdab7859268c77c31b62
z806af367bbd97571d9a417dfdb8956191832393cc9f7400e3c047e09d56ccc327bf7ee5faeb292
z0b008f9c729ca5d08d92c4c834e5b0ae1739c1f7d3c1b16fdbd546da96b73666526f74be4f6222
zd03f6f5a3a4825ca5a5315ab9f8dce36b95a42476b007ea780befc10eedefee4a5caf30856fbd9
z25e801830a372c7c3c8c466d6f8d70346cb1d51e37cfd952d95ece5d0b351e179d7a6977cc25ee
ze0e05738d4ed8c0eca41d86e76e7436fb6c6a4c6c2489b44ca15b7bddcdc0210adfcacf137afc6
z76018203dec2fea8e68109cd63aa9f9c2b2ca00820850040f19ed7b6ca800e8b00ccffce5f0645
z9b42190c0d6ff3acb177d5ed04e44125b301bdb073f30c3bccd66931de3fa7bdf1693e4400113f
z05c0d252b3b531eb3a3dc83fff4218a6e8b3da029d3d2e50a78ab46b45c6b7a72522add484d5a9
z22fe28068f84a9a30b167cfd841ce66307258c0bf82b948ef45b99e58bc1eee979e52bc579cccf
z1d1de92ef46a3842ff5291d27f74656f5407dc310a8f5f61f90477235766354b3824695d10ace5
za16de1d313e84934ac25616b52291e3655847dad478644ffdcb952bd8195f7e34b9d8f88d0f30e
z503fff9e6bc99d33b0dfe23804c616504385aec32fb21f85d4e4661e8af806c4c85d9c01023f0f
z1e9bad7a54714caee1052af88e91afdcaecfcbf445f967afcdf4125a532c6721ad3ca5b6bfbcd0
za3e99354148aeef4e5a7edea33bcc8cea7e32bef1d7f43e277e7ba0d6714b3f2aad755c4d39eed
z2597dc180dabac3063527ead2d34153a3cc39953524bb4019fd367ea13b716d3be786af1ed47d8
z5a8a216e27151200a3b7981464569409b79a0b9896fdd48d645a062560bc605518d5a49bbc2ae3
zfad9e9b2f6901fbd9ee994845a7e43572d22b7244e646e1328275ba9ce778100e12b9da4709cbf
z2b9752d57f8af70004358ac5dea6622d886c9bb382a6645241710de847b70ebb6c4c352df58fd4
z9c9643392633ef6913b92a716963f3fda5041672ff2467fbffea4c9384294991ae15f1f10d3abe
z5411f293f2425f5cf1fa9e9d0221079d948c0f20e752848e076a00e766e1812a841a3c059c39ca
z0748a3fe08bd76a6f7f5393b3f50cc261a9cabee2eed6fee381e5e0126c3669dea0419e904a394
zc7362e45300e6507bccd24c22183131aa6e57c6c4807c164b7f3653aa73594c7bc6335ccc8f0a1
zd8cc7f4e880dd79157db728338c9985cd03f829814bc6a6ffe44d860fc823ba6946d527e3e6526
z753d81255073762a4a0672503423ada1be9c7b60e6cd148859bbcf59fb2ee44307957432f154b5
zda9ddffd5fd36fc159c8bdd19e8d1989a42d2c6a91d577f438756559c98bcc5d164a327c1c68ab
zda827e8243715f1a98c2a70e61f6e8f55e15be2f96c8e8b0914a6adb6ef2d5783d0a4f49b48432
z4d62a66c5e438d742530c50156bd71a48a2ea2fce0ed17b2008a46f1c9c0ab55121155c2171c8f
z40034464f548c3179ea1785a788abfa869293da7ce4338bb1da7ea3eb539b4f6b5002e7be5c41c
z4542eed7b1b4f87e4a4e3c88769e6c48de06b7c9cf5ee6b9ac5b6c4633cda1bdd4a79c48312e70
zdc97f9818d7ef46b6be535248f510f649a675fb9b7cd7cebfe210f9e07f010addfa69041bd7723
z369d970bbaab448c266597936c24bcfeb314fdaf32a52f045626ec2e6ec1dec51d119bb772ca31
z7137edddf3cc3c38583bfd68af2ba3c38924580527b7cb3d0537b6182a3fdf8ca5849c296fcc41
zdb2fb4232da61f5841540874ed6f394f39e1df86b4b21070e4916633135a212a6d2372c34e99ac
z77a62bcf5c23d6a1aba1b4fa606e031486923a2768717e8fb95bd630b2b5866ee6eb8318770d5e
z02d1c2b380a16ebd165accb1c566fa286a8ac67edeaec628fb25496ea20af973a45905ff4d4504
z11abfe16e597643c7b52ee278305319887c8b5eb750017a7d7ea617e61aa9f00642b07bd748610
z6d83f485c1b133c5fcede21df5fd2ab55c2c7a7cd2010c8002c07fda84e83e2ee635de699526e2
z8f44e495a2cf0319e3f0513a844c0135370f8e8bc464f7f75be1b2ee0bbe008c465e1acea65180
z2985886fc277f7663389a1a91d8855f1ce30fc95311ffa8ab4f9ebfa95e62603f96a343f8128b3
z4bb2f961e9569fc7a84d039e89c7d22887266cf0951acede079a6c2146cde3b43d770b934d9efd
zdac080690f1e883594cbfec1be70b21327ff57c0c6794751b61f77e2e4b16cbba33a1dbf6e7ff5
z602acb17f4b4f4ff3649a172ee4513d62311c42c9f18f38f55cc9f7563923e27bd00da11aa97f0
z306eb1b3cd4a71ecac59a44c340bf964f02a4611e131312dc98699544bbd741dad9405075bf2c3
zca29f0a6471c1f86648cc21dd5ed32a7b5663b4b7783cee2497774acc963d9a4d980864fe84e2a
ze5e0f44102caf8f91485ec51c904ca2825f44a5350cef0cc7e353d0ad79e7b811333ae2d5f083e
z77cce80a7f404dd731bd9481e04c0e17556eee69263797420c45f15365507c7915d7a618b0afb5
z3a8793f9067d97961b185fc341e3cdc2fdcc112a4bad873fcde48797d37e7d8a91847a78725cf9
z189901cb8b60c06acca3aa83c5938a52bd397a7a396c9ac5c500c69b9b3b66755bd2cdbdbe1820
z4dc45a34ee29253207d6d85f844a7739ae28c511bd7c9c036d4793aa4c6583f41ac3b6e79a2e59
zbc752d5a0810c63c46d28187f8d665630642030576fb881ebbc50723aee4708319d742749ea139
zcb11973552ad8074dd720ea23baf8e8e0d3b6cbcd440d7a29936f735c7690bad81fc4ee70ee1dd
za42f2fe46c7a45316919a6ee51e2ccaf430255192582c0d59d72bf8271096ab41ee8f8d7b63779
zad4a031044d76b23c89d3b732fb3857b3dc5e2fd7c7bdabd98ec74fb490f339dc2e3f692dc7654
z8b554d6f768c5d4e3c64ae183082f68dc53c044e6dfe306848e2f2cf5e86305f356533fc82065c
zbfa5c9c3311e0d83cf5260e8fa29771c5fc1367684f23326d08142cf6470eab8ee6ed9c32ea28c
z4c0ccdf259a0eedd5f4a112b2ea6880aecc2db4b3e14bf54b6b6703994f2deacbf6397fa7f18dd
z8c6b73b4e15c71a60a4b853d1713a9a7ef0d98f620d11fb4c9d88cbb7879c8c95b0c11363e08ee
zcc7f4a1e5c63815c1156c072742870e29ecad0eae68ef4eb537b659c64a334f5fe75753724a5f8
zcf45d656627807183a64c08c448ec506d7f3c151fbd658a6b254991ed44a3953ed033c2e25093d
z291e30bbcf8a6fdae5f95fc11a7264210427eaa1f9b517470a3eea9d47826ac39eb3042e61d771
z6731be9836ae8827801de45af66100138dfccf8bf1a2f75cd9bf16ecca73963878b83a68dfb9e3
z55b667621847677b8c18eb65025f2c3a121446dbf5fd434acc89ec98773d06af47b8ffde964c84
z14f8f629b4ff50ca6d78b31b50153d0142a24b0fef20078f0d803981fc82c59f20dda7370a20a0
z7e597bb57cc6d2008f60768578ec0c822d4171ca8919827ba2c2df2bfb938e519d1a50cf17c9bc
z2e9a1a0a5e153160bfb84a0001c2d50d1aa1bb9076d7c078dd72eda77dcfafb28e5d2506c0429d
z7f7d53e5ec6aab6f4c28dee576d53a91320e40e65391d65023758f9c06d6a4258e77b1e1a71456
zdf19eb3b48f52676f6456f36fa2e7e9165581c93393615ef01ec97e8ec648fd68a64373815bb96
z61ccc7748c84e446d78dd3a8f7315025303c2eb6d87a9f8e55fb72757cfc0ce98b3e9dabcd8fe4
z90c52184f24721fb53ad226ec3511de1f92a1e8044b370b01da8717c7bb07fb85c20f3255c91ef
z7580a7128c09edbc4991be4e3834dc0b81d9ff86111922599a0e046655e6913b22ab775ce36a0b
z0f2bd23ce718e39fd06b9120a528d20d0dd1dbb7b5f6a732a12c6a99750f0db51aa2cc12d00d8a
zddd51d9622572e820ab36268b4bba1d16c57650567ca3e21e55a497ae5a05b9666edfa8803749f
z8dfcc6fa5b63de3dc3695edb6f0a3910b76b7471beaf77172d356390152e10b4db36848702f22c
z0ddb04512630cad66070677617b70228f03af18f8326f4ac8b79dff03f6b2f3de999a44e91ec6d
z643cb0c88f474dd148afc1effc8a36ff9e8e6aaa23d56fbc11544686a6be424b0614bd4e62b2dd
za3f25f3f243aef9956818f35c4e616b219107bae39edb1d58937c291744046da460b665df83af1
z1c95e05278861c6e775f8ad9d81e77513a5f214158503a6d54bfe011319572772f62431632ba8e
z3f0313944f4df7ecee53656557fec92b88c9660dcb1457dd7be13cb14fd9e6cee8cb7519e77334
zf30bbe0e71a14be7489a4e93946c54d31b19ee569543c4f74a1456daf29d1c27ff237a21cf9b47
z963a39cfe5c7d0290802fec682ce9d67acacee832e46038c93c21e7cf2fa3ae43cb67001f967d8
ze43175049bd048b86dfcb7bb8bac144778e8a9746381503a449f84a23d9e457a1e64f396bad2f1
z88a1cb0dd4920e4e558bb866f450609223d33e897f70004f5ad6edf582cfee0f40b329fdd901b1
z0d405952a9c63bc9fdbcbff184ec965c8dac1a6c708176d7457f30f1051524f351cd3d3abc2155
zd13b5f21849163a20f3dfb3ca68fd6b827ef47a248ac45a5b042c7ddd8aa6d7cbfaa54945718da
z99748406a90b38cdb9d6fbce1e0e487f934f8186a5e53c6604acd839dd35488cb8b409b3143b64
zbf3f40df7925c01493175cb1d60621b0796df44925d44b1a47350a84809457d4816e1930554409
z05e76d6fcac70caa98f1c8ec9ffe5f5754e3e2c95aa10114fe290a9ef9375d988965a30bfd8da7
zbe5ee400dd5062f3903f8a1d19b2f229c9e551f64cd6fef0800d356a15ade6dfd9cc7125f9531c
zc346ffbef519067c76ebc567ab665392398fd1e5679dcca374c2fce33461207fd07f3708e2febc
zd07d6d8ee68fae7c1f74740f64c1ab3973e9518f70d532d5e4149275777e49b74f6aa51298096f
zbf906eacf05670ebd116e30f697ea603e916cdebbf47a92d37963c97edb8a43e8263ec58441923
zd7140dec97c1309ae67d89d97808d8363a03549b682fb2de6154dfbd4b418fb89b3f7e3ebd78b7
z07c8befdb4e5b47aadbcea68e5efbbed2a13f059fabe83e53aedcbeeec30da542c65df1fee1e74
z4dbf3e5ee93ccd2d1291329aa2818a502c24c8d7fac73ed87b0ecf22bbcf393e71e2ec275ee113
zc89fe057f547acf5defec98ba22016240ebf52926ccf06062c10d78d78e6b27f525b8126ba0ebb
z1d7e8b41dd77f5215037ef6217482fd3b1a0bec74d870fcb34c093bdbdccf594fd979dc04a5113
z149887388960f12c7dbfc930aa129209d9ec29b4b55c176b3a5efeb2ec790ef30f9da0a4b93c1c
z8656d3d6ae37354e6d8c5417a44c6eae36479cfce0be5da243c3ce3353189034d44d94f6790b3b
ze7e2ef96ff207a6c5fd4052a3cf177b4d31b5c55ffc3d972539e259efc952b33fbbec8ac87f952
z2e40bcffc4296ce20f4f394164c70e474b2b2849d60819164f0341eef4a3b22f9202150cd16821
z44e2dc8b3aa9455a627aa25e99b9e17df87d21a81f327be17006fdf2e062f4f2131d7591686402
z3ace260a1a5cfc70526dc4f6842c3082c7a5efa5aaf04d93ba08810590bc11d92e2801fe8ffe72
z9de9b68df8e050c59972d6f2d9772a6870c89494b7b237db8e576b62a0cb39ba03b8116760bb4c
zcda3d7b5ecf73f3ec9c3563a26007969fc0916dbf11d7d9b716ded88e5e6d697f7adec39e66781
z8b7a58880b641228d363264293a07a7201480795ebf52b4685138a6313ffbbb588e4bbb059cb77
zbd19677ee3c43e7081750e9a9d21162c8b46b64f5ef7fc64cd687b5eeba5a1938b2f044e45745e
zacfde23a282cb848ae1a8f8fbefd59f19728faffb8d992fa6e57281a105c3a3f3133a1879928d3
z3841e6d87e7b5560a8609e3f6a0d6cf6f0a802aa002e9252ce7b60a825155c71618b56f91bb755
z05d712c061a3a4a12a45d3e7b20b64f80e82bb964777dae63a99e29b523c4c58597ff96e412e90
z4da5c1d8531c5b78ba6776bf1e0d5c7daf7100a7d18c394364019aa016d0a8acef938eaeedd6dc
zddceecae6413ace32d1efc60c407dab13269c050030f47372e92eb190d2828770827fdac9a3f58
zf7db944fa458b1c071d54e4429e5533263be14f3e9d4b6d99499ae48c69b2cb1737c78143ad348
z97c658a6a0700bb86a8ed4156f2a0e16fb0ac71f7af6702c02df891ed468bec3fad117c4aa11c1
z6c2c50fa77e5625ebff0fca4cc7ae6a85d21a9c7e18029d24e2840438e4df159c5cbb12605c45d
z0f5e880c2038d973467f383a563acee5b0f7e2e370a5bc9e4cc9506fa4680123e035551f64a955
zc7e17df1a61674bfbeeee94290d3290fa16afcf0d982537d4c3b670465348ac2215d7c227642f9
z3aba27566f12526f5a792c7b7b35c9929cde0f505daf184425201098dd33e7e07cc2d1c01819f9
z350117d42835f48ddda87d1e72f405a98a39fb4647a57028739b9482f7c24506a6bdf47c943157
zbfcba30f1b3985c0d450f381d3d591e3c8a5de5ab0a79f389deae1e90558829ba0fece2045502c
z0ee54b88b6afa7ae2cfe738d5686b3ddbdb89ec91359a4c8db264ac05b3dc4a4bde46e607b7ed0
z1f58163b08c4c9a21f8f29d9c583dbc1112dfad913e960b0099efa06531b5b9974364f33844b42
zd7a7dd5947d2a23c2c66c3b847da5612aa7abdea0cd9c140238390c870027655bb622056992772
z6de11431fc2fa279d88f0a0a47ac705731aeca06ad1aff05fea9f3eafdbca1961fb7903dea0a6b
z752a55a427e29c41961fd456a4447d97e1af54de6010804df2697149716b4330ea311161101343
zbcc860166ff2b0b64b1cb3e59e2456709f51aa9d4ad13ffb38c0a110002cb010d72ea530c324e0
z796d789a5bba2460949d4ec5d5a990e0d7914db7cb39fee0e2d86c2bb20b6b71a1823d15b5b8d5
z7f1ffb759c88582bbee25b3f387f574d7edacf0ac7a8b4e97447f2bd77f106fd0fa94b44718b29
z6e9e62c9c2b29d0f5929637a991d222dfeb28f45121231afb3b21eb7642fa24dffa13bdcf79204
z1631a7ccf0d84fdc56d4d0c6d630eb34d6dff246405abf39ab7cf9c48ab3d61aebb4f26a66c551
z73b8e6fe5d3ff824c8dcc434bc4b2bde90a008d4475662a1ba75ec44ceae5cf40e0a0174a2faa7
z67f1493fb10e6f6bd1080637cc33df170d2e8c36fba90d24d24b875a68d8bd62a8375872917ebb
zc23581766fda8275fae4e080208d59d4b71895e0b7e79365a72b1363ddbbbd9878848d08bdacbb
zac730cd02003636e5c3d58bb8204d9f58386f314d253a1c5a94c3f127335f4f3e9b69580282e7a
z4687326454a5d749b72fffa15c6671ea46da0102d0b71f74b773304193ed715ee9a07ad9e5fcce
zd3980d675d1c826b8617d2f086af6ef05d0196f50fd36d9590368ffec4bb2635012dc9664d0bff
zc977eda6140298be567cf76b6408dde06aa2ec47622fa245a71b853fde299a2fec8c4663e1342e
z5d322fc76801c2568ef8159cbe4e031309ae1ef0afed977717cc1c8ec51d94fa7c4d9f47697b1d
z70bc5a7524464ff5a511e98242d59ba005d5acf1ae4c1cfc5363410d1563b416a011852acf40c5
z79ea7df0f4f0ead83bd893d6ecae9b6aa9cd90981f0749793eb7143970afa97175981ac546d523
za09e2e26c0e1d8e3e227e8da7e7a648e608667a5126cf7ed3b04f89167ba4e93c9aa91597fdc96
zb088b95af7f18ea7be2f6842f968a76d63996ff9d759737010cddf521801c8afaa66c76293f595
z817816953ed8b10fad80c9dd9c9ee2244a7ccb504bc57a9fb3a8a9a81048b7966ccbf4e45edf52
zd4dc784dcc1ae476802c95eb232bd8fa9c619ecdb7b9336714ba9a9acdb3fb685e6f39c8729dea
zd518aecbd6e4a3ef69189e25cc4741b9a706fa935f1cd01122a3d5568c88ed17df5f1674b109fa
zfe95bc191897c441cae615930c4adbe1fa778a55a671a95d5062955caac2b9ac196488da221979
z3a67575407ac696fb6f1394d15735194c270e4515d0f278d62fa46b4d2f23f0348a96566ac58f7
zf3e121b4c5fe4eb7ffc063aa57c5c9cef70e43091ef4e72e3c60e38b0b9fa9bbcb035dab70f9f6
z23ec8672f5c9d7919abc72f5958ba17733f50c6e4892278aef1b851ef399c6259cd4efecbdb2a3
z2303996a668c15db69bc21e959184f075cd66969d108b3fdc1069a75287460c5278bb8a8e9b702
z83bf78e2f33a880ac320acb290f698062d3c33155c904598cc4da0dcc60a995498e0c5851804a9
zdb4b1b4687b90d374820f2a187425502f7b75b8d99bf3f1a496a9b55fc64c1df0b00144f4bf74b
zf81fc102adcf3c0f610c036f24bd3d2ebbd5899ae3b9d4a92e6ec666d4f03e8b8b12be19eb9b1b
z2f9217f107445981cfe525b726fb319b29528e37f5d1fd8b7146848d0439819c7581c4cdc45469
z3e6418f29404fa1b4f36b22d91124da4f8940b91c9b6c155961f4162a65a5c1829b346e3722a55
z012a41bff54be37ee7b2802b4527bff9533aeebb38ced2c361456f1a39f99e6f49053510a808e7
z972a99d20d2b9505a3205854057410797d7790a4ea71b4c24b8dd4158a8c1ceae45a76198be873
z6fb9eb2742bbe0e2d0b0fbf7e38e634aa13d67c0f6091d551a6d34b532b5a83fce71c8b111375f
z3039d3ec857f432c8a9876c2a99bda7fd10c8d3c485a2ad7a4ee4cdea412fa374334f3e77ef2f6
za939b790be05d8cd84377dcb0ec87057ae7ca1dd102ee06157647a6c4cdb53b16fe42ba1fe59ec
z8d0947534ff046ee45c4be82bfea31d6e865fc12d2b5c07b7f71733ffdafefc6b05edd8fd821e3
z8ac73d182299fcb0a82b4d0a490a8774f15001ac73a5751951e766aae70f4a291ebad480073063
z623e636a1864ffbab96bab1b9394c58a9f55e7a1f101f5d71da4e286131ece4bed217f1448c182
ze3d8698e0455dd9c949cb843ad6b625127cbb25434cb3283445dc78b4e3e053110ebf42e19c237
zc829c5e38ac5172ec598dc6148a241f0b72cf6f9f6776fbb3a11d456734b19fe66120dbd720f96
zc3594fb2102075f88b5b5f996e5b62a3a18ff12399abcb95063f11a18e38c217b1ed6ca9b7db43
zce7e009eccc2682f731ee6670c2ada385fdc3484819a1a7fdec8ecfa27134ad4d8eedaea500992
z159d631b5010b070490160e8e1c151aeb82a15a93a2398d3a1e9af8750a7ceb36c5bf0f58921d2
zb5b3db78c296fcaff4a785a7474001966cbed4daa9e6b50dffb6271ca1f8067385ba60d411f4fb
zb6892da5fd444f2e8eb582bc9e76c359ff64f6c0639766b729470edcaefc21cf073251c9ecb33b
z6b8b63849bf14fb268d6f62c6e245d43e8356161018d0ec01dc6f77de12a084ea1af8c612bebd5
zf149e3db95f6da2d4b02cc8c3d293651b428ca4a66ea8f37c475f467c880727e835771cbf17024
z23f12fc9adaef445fa4fbe8c30b44ba7c62dfcbf594e69a81d4e698d263f3e1ed4efb13aa0f88b
z99fdf4a4392bf04de0a06da13113bc811a3105d33e5d3901c79a944300f35dc2b92c43c2d4f164
z3cd2a749b44bf6999248f8cb3ca7fe5cd95f2946b0d06f4254b54bf7c69e392df94e3dc26b7e69
zaacdbad8ac5b77e7b28f4fcb8b6f6f56e53d1cadb8ce7af9ebd85ba5c5ead179d6ae08fb74c2c4
z00cd540fd181872bbb296f43d4f04c931528ecd4882d0a6fd0c72b4107dcf8b0e136f9ad6623a8
z467f904931f995a102146ee21b725604d8630db4a17fc35ea40ec0fe262d4145d3207c431c8f26
z66e5b9659f73b0179682ee0a830a59179442bca925070956db281aae64820e306903ed39346762
z99ea3635e5f4141503000ce305199500a0a9894e1c6c1bae3cab8a4cb81f145bc8bd952a6ad418
zfa4bee1d793c91ea20e8340b73b64428e8b822d1965a924d299f766b28368c727e6bd958cda3e1
z397da48436e0856c664f52e51d1b26ce5c5085628daabe8ebcb08811f7ac73cfe9a90092bfb63c
ze57461779b86c558cd7e8817947b78c759945a203ad0a69829b96fc3f80286d01fb6a618b38c8b
z47d3b8159a808b59b8bcc05c4c59b183e6981ba2db9c69a5c17f4545602ed79f216edde86e7969
z8d00e6db2f148fdb27b42949b5f61c32b42f0e4e7cbbbfc39e51e315e6ec7d3be1cefc407cac19
za57f793bcce63e60a6557acc1ad502a3c5f507f471b7f5c130f0ddc6
`end_protected_0in
`else
`ifdef MODEL_TECH
`include "qvl_gigabit_ethernet_xsbi_logic.mti.svp"
`endif // MODEL_TECH
`endif // encrypted_0in
