`ifdef encrypted_0in
`protected_0in
ze74c34e226135848fe16db9ffd31815111b6d7fb642c521a3f628cf6da949865580b22efd062a7
ze90adae0e65e66a2c36a587d0a790699161455169ed55a01f2084f11770a774ec4c588039b380f
z6de9c5084882a40b79a175f5c2114b2b6d78b070cb806e1c0aa9258297f4687ab30857016fc53a
za25afc8341302f0c829d94450c399b8ff9b0386c187cb854ee330605b7b59da379b1f26f488e1d
z36e675f0b1336408b3a1ad87d0723054f952fbefc8d5a33eaca6ef5be8f42bc59870a29a5cc9dd
z4fec09ce6e44cac279651402e7e1f590df88ce49ec26ab39f12b4a02855703c6f03b1e85c797d7
za357087d98e5b1f45502e45892e5823d6fa4b762932009620038c05d74efcea7c3fdb38901d620
z36515d0824367e48d1bc182335f158c262d396cada6b0ad58add4f945eee634c2dceadbfb5118e
z14969c29a743830a07124bfa78707f3952b96b0db7af7c9ff36f77137d8c490c4f79328328069e
zd7d5280e4f95742c9841340368b9764f0f80413adb175ecfbdf3c40716abca7b8cef6f7fe92ab9
z6bd2453f1aef7f7899c5365c5c83793cacc7795c269413f6cf0dabad14d40e9285afde8c01a47e
zb61893788ec5060288cabde8fb553f21b02eac61ab0b48ad3d54f4d1d76508b22f0c600861b5ce
zcb30ba708be817b1f50f59c0f6fce449203e7355c1be55b662fef3f92ba58243d81537761af8d6
ze27d7864d2dae99372b2b75bacdc0437a4f7e011d68c3487a89759e3625548fcc920ad06471ee7
z2d701aabf726859343208b0a543c73eeff8406febf277e3babff437ec820fb49d6b78e73bc2353
z884917487d35a6cd06d7d73ccff5f0292fb3df6f439aded7c8bc5dd0187f22a0fe1ead93318eb8
z8c6e90111edd2a748769a8d92e19030b0323140a1ef01d3a257fd16256b12b03810bb4a4e82398
z2704088d587398546935b6339280ed10cfe93a3a5b7a4f04e0a6f073f8fa718c2f9190d76f588f
ze9fdbb73c2c6c983be7680e758043939fdd6803162983f37193ecbd51d83a9df901bce5c960f7a
z91451ccc98f8cc68bcf6283cc3f9b8b51e819fc5551032ae29e14474669999e5823f495289497c
zae28a8b4ebdcf6994f4de5bc4a011a9e97c810bc37473a1c49e8a523aa61750a9deb7cf32fdfff
zeb9463c632da84a78cf1a3608d612a0d34101f2fef8ea5d2be1f503fe59ffca705fb8449fe8266
zd4ff3b3a90e594935250f1ed844aee02503f5f9fb5bdaa30f12fa6c0447d9105a1d83a4a0a294b
z903b904f73719d885fa5903743c386099ff43bef2eb1fa8daf2613018e731e4428d166d1356b37
zc80f24cadada89e2f5b438bbce1d33cda669573a336c0afefc1412371d278c402780269e649e18
z88c6916aea8e688e3a73aec5dfb3632685ecd06fb0e4aaa88d4f1381bf2dbc1a4213d3c2d859f0
z341197c61d78e15c1de7a7b49da40463c00c01893bff26435e370b18a4c977050888d114184756
ze6991a6b4dfc2ec5b402952fe4ce176821f53cc284ff5be4c92d6046fbcdab1df78c149c4017b8
zd97342229438e161e2de89ba1c9f60fdd4f08ac05e832b6e0bbb5d3f1d4ac7ae5aa62083d72f52
z1b6c3c95a148b87175bea435b0effa305dc8b84bf55b6c5151272b582b27d962ba801d0ff05802
zc0390d678be337e406037f603b7bf50a4be29d7fee9781d65fe7ae7ac0355872bdccd20cce4a32
z827f81656f8c1fab3e628649de2f14a590ddfc9e4fd488799c9feb80d0e718c5df7db449edb72a
zb45b2a6d5beaac8a08e6ac96165ae550906548e122fdc6a20bf98e90a051f2c9506a41c02a1521
zca1f52c72368c23f2bd2af6e318ff0a4110be99f0efaf8b59fed44498e5eb7d08eb80e59e68db0
zac169200c9e107e92178f01883853c19f8da7229fad600e8901d95a93c04b142248c9776aeadec
zb2391ea73c24235b0a9c2b541a6fde68255e04e4a61cceaa7b17b744ca96b17bb636f3da94ba07
z5491e5198cb6e233d18177e1e29d53bdbff5bce4b9451c48aab634d62d7a7d235bef8fef0c55ac
zc3f06e051711ff5aedd3cb35729ce7a4bd46ef969c4f4e74f1e78198f1a3a666b075fbea147d9d
z632ec97ab88b2138c52d989aa8f3b41958edec72b264facb9c63a35f1c0dc8fd4cdaaed2bafcf3
z4f2d8872b1bb238cb028b7a68f8e45725ae958514440cdc5b502b9f2ec627fa56bdeba2541ce72
zfcfe2fca9e5af610ec0148d3b4ed8f52f7042727b1f88c61b9a110a4dbb7ea9b584cef7644c989
z9fb51b71f9cffd28d3896aac2b06f034b48bec34897bbdb74d11bcac376146671846ea4119ee98
zd05dc96c4128d516318290a1fd9054c4f715a968859ae027ad5414cbc9a34b9567cc868aa0a295
zf4d38172e6f7efe09a976c4656fc9676f1daf3ee1226981b896bc6a9522c66908696d0d6197d7e
zee3beb89b34d8a2b7513b040bf93604fe9d50d4e5998aa6d0710c4a41284b59de3ad9794e58c60
z576500d6e938e5c11c58252520f4b57f0fe7f465b23d04325ac67b71309194759f342d8a936a3a
za14b394d6c570b26de8027a1e8b98e6c3266b02476cbbfdb948da6de47cb269b4df7b05e2fe79b
zf55aa96feb88aabf5b06ce3254fee2b823c5059707a23187c9b835e8be12ff59eff32c0a050619
z21807e4894f773371c848f23105ca794c20df7e9bc306d165a31346e452a4edf0b4a9e3964f8ce
z3f78404fe7210ef28debe3afd569e830e78d0e82e69c6c5f2a8b33ed5c689dee64025dec1c937c
zc32ff84838cc9ccfee05aae537332be2ab031c5b16132d9b78b58f89e008cf8947de23ffefa40b
zec24ea8f1867fa26bacb3dfe77a87920f3980118b88470387cb88106a0941e007007f5a6b9bd9e
z0597018877bdf6811b45a2a2dbcda8c2923da14c45b4270f7b23a9755dce3471fac956e9c7b36a
z096a2e1c0c73de20964bd08a563387c39f35177d1c34630be0432bb327f03d0214babe5ce84f38
z8c4fbaf3b39e9130a58cea33871ebf27ed8f4645b816e9c0041852215b0bca935d88c50d8cb32a
zca4c9010a1928cfe317e60f856874f6ff800e88b1d74962e154307f17d4f5140cf83996549dd51
z4e3ed16c2ffd4b991458b21715dad124bc130114c27633aa2ef5213ed393dba4f2d2a2888796a4
za8ccb3d41897f5e74a374f8c1ba0e4d107eba1e403954a77d2eef4e4c03e31efd493e68616bb53
z6a6c8acd2a4798f268291598043c0407e278780943d4cab2ce02431cf341e53be5699e69820007
z9e8172a571ba0d462293a4bc3362a773ba7d8ec7f7dc72677cab93aa8e63239a3b6edc777581b2
z24b0f6229d675610e91efe1b55a1178352d998873d195fdc6bbdaa7d133d9a204a5acc0b559230
z33e5418e19a25b1bfc7fa1bd44abaed9db222cf29b3ecb2b923d12f888baed77025b8129a03974
ze71cdc7633db30c75553b804d1a5ca2f53417d431660b971f7b5689d2ab743ee3ec0de0f5ff9f9
z49f44e04c8d8ebde533de126fb64a1344e71c75795ca79b5c8ee012e4f4332f7574b7aebccc954
z5a97846cc24c6c1cbd79141b5960a7c4a0404e8a7cbb398f0f52501fa4f27d74616affa155898f
zfcfaa25c96813f65c983298cd1a05d723d61ebd13d0b063f4d9516b5fe79dd7a1127d4fde36c57
z68c232131f57d8fc9b49f6fd281826f4d1d1ede97871e74c01678b4a4ad2e80953e7602fc2c75d
z67a55a96f0cf214414d62e8088a93b3c521050da59c8392b07befdc5fccf359f9c57e5f54bf105
ze1b535dd0224040395ae2da75461d937200375b0c8baea9526b096f4d9814601ee7ade8b62d4a6
zd17efea42e541b83366061ff0e01e4ce4ac65fc3024aec00b5f9463b70e55e1959da86b2ff5f1d
zdcbcb46a70516dede72b1e20e585930f3904b3d221d3f6db7db36473bc5c9f83ef7b6aa89aab9c
zcef6947c7bb6e5fbdaee3a18794e946f7ccc1aa2bc7647aa5d805c694ffe1d7f6750b7242bda26
zd9b1d58a254907e31e54766a2238ead3d49d0ca255d25fd15ddfb7e0dbef173ecc246326e0aefc
zc92b4183808a007a9d060759547f5b652d102c218ef033ef33795965345b42dbd38a34f09fa0da
z852ce74f3e2d0625840ae1ee5e61dfd96d25958538749f8096614501500c95bf501dcf20b378e6
zdc4aaa1fe56dfbbdfb1cf2e40b28970aec247d3eca764694bc377329e4ca90a6f234cdc527a160
z69c9a60b6a212a741a1edba3971598b41675d5c2848446d7af14fcebb858a93d19717607d67c6c
z98be88237b89f8c008995c3a76a1cd3a941f22d4e60e58e8e4a01fd186a9bce4b0e329ca1ea372
z439f84207fea37b8e7a902d731e333104c556fe673e37f161ab0c2c4afbe96eae08ebcc54cb2b7
zd88db94e6bee5d33b7e3138a7b4fd1ed0d06222a8ad54d78241b0422abf431daab033a798a306f
zd2d589cb30325783cdaf6970662bb08334c6a5dbc634d464c4cb8c2647774509fb75624784674f
zc0ef244c3498b3fe346c49b6a9a34f32d6fb0a59dfec72235af1823732efc192bf9da07166d173
z73b16dff448ad9b744d7e8c8c1a610e6998fa2c7f1415898a2bc538a8d9d175752c237bf566f13
z00142ccfcbd834582d6a52354982d3773fda64cb509087e0edc987b14a7975b5a41aae027b3bc0
z7cc8beb74fa44716a02650cf837651e1be8411a83cb5ab281b6482451f4ff4386a2dab3e3a3595
z047d1df251c68deadc4394cf6454e31f313ab80dbe53c3fc64e82b9c0f9ad1d027b482f7020602
zb435960f6ec242174f8e2ac28e57de4fc35f079a87e072f40b545ec5f43c85d659bd2b18562191
z3e9c49d35df6a3fc47ae1a9101c4c63c2739ff5299c79fb025294d5cdb56080df7e38a5791bbbf
z0a701dde815162f5ac52525fcc54e291873db09ac23772767bb795a1e5d419aec32d497e08e962
z492fd534b242c2fce0a8691611f1e2e1c8070ef196248a53fea1325f4dfbb2f66900d6ce2719fa
zd290c739c891048d66c1e41ba4e98b88384859700c274113d3f4ffc5f166b4d300a02555af7fdd
zc9a78719c8d29b6a23d5c47a1bea6ed15e74dafe725a3e7cc7f90134092155833bf3a295b5cd96
z419b887397d1cc78d9c3c242ed9718ee5dacff199fb8b199b44fd4297fe35ad3d360b1b1826252
zd1c86cf66966dba2552cca02ce4821881814c03d32c967d934fe1ba67340154b3858006f0d881f
z71668e171afe7c83328c80677ae5f0c9423ea2f622a73835e42bd6dcad629a0f4f638ed6ebb277
zb2deb1accd693e92a8d14816ff80a168d67718c9464ad006994f5560a28af2863c698243f0fa48
z01ea44699a9d743226bb97ffd4775999d1b88a1b3b153d330853de2f912ddef43b699271e109cd
z618b917b4c3f1f993a3b1daec5b315e07941617dfb6d714b4d3b7805993d8421709d8a4db48911
z1ed259d469d625df53e319543d35790c013ef870ea968d837530a80c4fe45f567073a6b79ec68d
z93a86f1e78433cffa9659794ed1394d18c0d16dac23a5dfc22b8887843e03041d0f0f0c549f8f9
z9733316706f30ad90942590b5056721248bae496bb023071441cda29c8f9bfaa78a948a4474a8e
zcc1090ac4b8e4f12d2cf8468429d0abd109542124e7d7a2ae0ce6d22e2369266b2044296bc6753
z25201d6dbb3ed4c3fde9886179f70741a9188beaa38bb7cc7e7799da687eb9636130ced072bfd4
z279ce9cb4f2fce5de1930a7ebe3e7efade96927ff204daab8eaff90cfab37cb37e1c6a6af9d32b
z438a42ce2d31bfba430c239b836840c05675ecdafca2709d9f44779c545b9c6637e127ba53fc79
z191a59563419ce2212acd7a2f85f1bd24d20860a31f8aa715b38d6a62dc3309bab01d386d5605c
zc74fa754513968eb7848474dba814c0c9e0679205bd7905bec22c29706391b926efa0a0be65fe1
z8d2cd1cbd45bd583015e0ad0c6db770b25d33aaa7ac3bebecb507bf838d7554d34bdc4a668ac53
z28055c6f886c0d4fdfa081c3e64113db05610d24891eb8eecdf0341ac18bda1f3b6be85b9e6835
z017a8edc54795e1823679e580e123e33e9ff406dcce0af5e264d9c5d537d659e6536920c5db24b
z40bc9a7b9009c36f4749127b9848949cf215eb05ec4f10af8edc702b248131cac098f33b39d70f
z86698b01aa708bf20deda768550165c41cb4f6a246cf59b4378cc695824455eb9f3c532f948912
z487ae075250d1137516ee3f0be97ed3165c799d5044a56a54fb46f2262f24bd9780083e50be4f7
z1dc049242c11dfdc184893cf191019db135dba4cbe3069a60e804394ff768cc3c922c5f887689e
z61a53ffca4e3fa39ac23dd6fed8c75388b5748bf7e90c53e959a1012d6ee185d79bb0d7a338a89
z1b6c3054e0e08cfc41948f4601e0234f5e6fddeb24e7c873078b98ed0e75e61aab21486c46a016
z2bac305504e474f02cda07019b075714576b7d7d1684e85aa266fc98603925f0a563a6411e14ec
z356300a89981a2b8235ab186149bf211bb2351b8e64036db75141e362121f85019344fc93d884b
z1238b8d36bf2ff5c6d9ac7cb5967d98206d9dae43d45d944aa78a59a258559f2183f4d535987e8
z88090442ddd4d04a4ba95195899783f4e2b96228d8a9a3e29545c509ff8f2627c27411e1b1a4fb
z6d2b3d34f92695b9dae0b4d7c234e4fde83811d23c9250bce403db34d705fcd54468ac56e0b5aa
zb3a8019b66f8c43c8b42093c208d086a73d57572dac7f4831b277c50c85f2e96d13baf4d8267eb
z790d65b971c058303c9ea03320fadef565b863076d2342d6b00f1c65d7c8d5c5b7869eec6008de
z3dbdbbdede2bd48a86e99fd4c6e84d43f8018d42650c9ba38d890b582a1a6d78b7d4ac7d7df830
z1620606394d728a9f58a49acbe22b798030b604e3d90d429b5a015e70095b80a4392dd4806c73a
z7e71f7192a3771bd46099fe754d3a70b102f3823bd2ed31fadd24aa6a845d7686ca5f92359a2a3
z82fec0ceff85e24cbb4ca9acc379566182ec6ccdd101d0b848e3bc144e8c675a1c1100177d0f10
ze04b9f82cfc6bad902c37d69960f8c35affbb04fe681ca755f2d2f1b0f1c35ada25b93ecb93f80
zc42f2b5ba5c43630cd399c690d6ad12f9473ae37852c600f3d1a911c15c80c66bf495b7642d410
z941188748d7cde14371ffe6e03e0a806950f197c0c6de2696f4e010e201bf2589594d682c9357c
z5b6242592083e0d4b9a26e3d059f61acff97d416b0f52bd03e0053ec5eee62ff3feffbf147d170
z1ea1d2cfa656db72dc26f030e4dfea0ffcc5bcaf366f79d2c3601296e732f2c690f7584fcdf7e2
zc0839b3ba2e17048749941d440479aef3b96a53985c134608276df66fa373120d62ae2043dfaec
z8f711cb9eda7820e03735ac626cee1578a5fd0ab849304c58b96da0f7870ad7f40ed915007b3bb
z2a2c4c8a91764f4b3da490c4edf7e0d4bcc3aef5b3e466faa49557d4e3c50ec8c0620ebcc64f95
za4eac23e447df5f52f91b5eed9177482803178e072768b5112ebc860e164bdd21796c2dbc9253e
z6363ce43d0616b7239ab6130c19fb6b5ca6a4923b790a8f3ab28b57fc115fb134bf5b99567804a
zc17bab252e2c47350623964b4a251275a13c27a09f79d2b25e0cfdb14417017ac51599959e5a62
z8514cc4d7a4bb3c83c5e54a1f4991ccf48615c34ba4a1072b066f51a05cb2af37eb266578de8c2
z3b76ae0d4ad8ab194d86fcf20ddca54fe85dc6e3116996d82b8950e5a04b2c36b01c3ee0c8f16e
zbe78db6f8ecb90b1230202047247205075c54127bc571ce205136aa1388ef674959e214074d8cf
z010c4345780810fff37d806c3f0cf841b90d547dbdcaa6e2c3d929ddacf9a540476bd228d9fd60
z6b0acea463fb9ae742672bfdfb756366d575b85bc5a801924084e5369dee6469a56f82154c7d4d
z48c356cef7c0dbe206c5c434fad8a41c2462b2c6337467d32630fadfb204028388067cf02ec141
z87c906e3c3acee669460545172eadba943a57be0c883ec3fc05f776954996a434b840c9784116c
zc0839942c771d2b91f9654854cd80087af5284b6d2f4174d597af0865a119bff70d76d496a3c2b
z12b38aa71fbb966de45ac8086bda980eff39be515a0aad33b1ed85ce8b50c92e242ba77cc48d14
z404b5276257ea9ff349dac8d308740fc0f67cf4a7cb5899cce742b88b27fa45d90194d116583c6
zcef345a64cc05328f7b46a16c5b7473e1484425e042a6677b4c89519977cfc3523c392c8d8bf14
z96f14bf55641d57cb401d887e5fb2037cc29e36fac416675363ef515b64ab58170c0e800fcf620
ze388c3e65706fd472dca8c82beccb9388dfb5576cc9d87be1e6a01a8ac0b4b7a67057304499943
z69d07331ac1eb2db6bdce24196fb6e7cac34e88e14c499836bdb4b3edab9b6dd027ad77d88c3db
z064dac517577fb316025ffafc821f91f957c0ec5c9c13acf48400f661fbff7ee9aea65af3a22fc
zc89dd7dc8bef29c6bee18ac562395010ce61bb24be039774530ce626dda40cd2990f919c1020f3
zda34774f1ce76003af62c5469975d3a42138f1199e10f369df5585c89f83c4094137a75e9b5ef4
z36ccac962daa48e5cb8f886e355487f6bbc88a38794be7ae894157c8bdb49753de444385559603
zabf9248ecfeddaf31c4b4a24e57fdc0b3ffcd6a64fa3a700aed97bdcf28c8eaabaea50cb78463e
z7c03211f19752214d93b6274be955aea9e5a2d9a5f174ec7224afe2b01a122341b132ac7f90ead
zd8837f8a6965ce9a36f7dd70ff808a1f7ae820a8b26805719d40fe32c222c1ede5f93ffa78231f
z78b0fb76a037fad7f57d48ffbfd800cc7480a3c38383cc43704825ea2ba4b123db598deb04865c
z5be66306a6375bf9d51578b6a1f873c76b23d6611f8796f5e0efa383e6e598cc9eb0c1fc30540c
z5ce235395b1bb3903c16d0f8aea48be40543b0b5ab4621d71645951bd0790fd9b83b49e77a5392
zb03889e648502d0bba90ae3290d7699ee4c2ea1ec351c49595a4044f95d82311d8be03d7d51430
z6c6ab3c2609e2af7fe825adcf96afe8f0829833062c6905d25cef0e51087f04c210485928770b0
zbcb6234d08b0b9a7d9f9746b2f5e37a109841d8f6b627411c85a5ac71bc751b269b189b1167db6
z044f267708433118e6b06afcf01ad6b2d44c60a489eb5237797f9e3c2bd7689547b52883d1d713
z6f95397dcd4ff553fba6e416b6a52329d9334c3492c85a29d0ff7f0c33f73a62185b8ea6e89f9c
z177f9b32e712e9a901dac389596197054e7c2fa2face83a0543849c64dcc52dad974e24b07279c
z965d6810de319b66ded9d463237114ed9b33f34fe019685749f6112be368e3941d35f86855bca4
zbba9294a443854fa393d68684c8dab68e1a0e269f22148f4d1533775ae46b9154d7bf78453c1e3
zfb84ee87b2f4108488a29f30406f5bb3730e61ac202a1384a4264f9bdcc022aa67910b7b3875b1
z800fd01637262c4a2031e47a2164f9f1a8185803b4ce71618c935955fb18327538716fe6652dbb
z12cf97c82dbf35b7f68c2b33b5fee5831f4182eb17ff09daef8002618e53de44f57204b4a414d0
z4654637264ca9459b81ea8bcbfbd80786b507d244fb7a0e3ba9dcceec2ebaeeb208f34476d3eba
ze24c4934847e0797a8af9eabe2353f0ebdb1be7238a60090d3ffba97238f74e02af27ee0475390
z2d6ca4b8cde8c287c133adc66908c8036b2d6950886035eac42c18053030747f9041810b96ce01
z682867f3390d7d77a873e546dcfa2ba3ae11a213a5341e2c47bc922db461ba43df6fb61cc92b9b
z8b7d8089fa0137ee9ae9a647a72aacf50e99590a7634daf010fa368cfefe30dacaf02b7a313339
z7dac3c82af23b7894149d3f632f7083c22fe11a1171d3be47a3422e849c8422501b72c337798fc
zb888bdd344c04a9f87289824962fa4dec8c2a118c21eb55b1274b71f15df474961e0986d6f0f84
z8b6fb1febdadd95d168d2df98f87ecede06254187665485033ebef086adf00bbb9581622337b14
zb0cd1c281a51df60e7465c42bca6bdef823394b5b0eb491f1df28b7861f79524810ae70926b717
z30c77a87002817a9b7e888d19dcb586d3ecd1713559de813de9fb2f7e97e6714dd63cb839cabd8
z0e91b4d5415e85bf18ca92b1c3054f17d0f90b87cac22b5a6502ab640ebcd819d3c275e6d5fae2
zeaa77d09688551490e5dee22f5464cdda5f85fcf8a271127a8d1315433bb78c91c24d2dd35213b
z3eeac24aa07e0285469ff3ffb81c3579840db47ba679026677a6faf178c8692b14c36bc3876880
zd1827dbf986110283f3b34f0bc5ef58e4bbd3c5b8f913806dd39125c922aa4e794ed6c33e29a3c
z9c8605f4f687bc09301a3b746c7749466e4b7d3be00975d5718a7aa72b33104e308409d0f6eb8d
zec5dac9a07fef1677abef3bde622b12cab1cb3369124eb3789d5ffbce704b9ed777d68879cd1fc
z3e3e147564eb3b60fa839e3d9fd1380592df8395781b55c1f44f692e101e59b3e732a7ccdc2a4f
z27a6db0c2efed996a966e082eb00003e932dbabfbeaaae8a9cab6a5607c7cec110eac0ca96f86d
zeac1bdad07d03bccfa223150c22427c9fd0c3c1bc6496c2d3f53b307dd149e8d6b16bb6e8d2098
z6b5ea0144a49031ac4b342ba3a1b63fdbbc1b47c1daa71e42079be6cabb0495d3e0e4d41221e51
zce432aaf23603a5560b58714cd6d698346d32c11cc208a0e6a311a97a37d1b24cd7948ec6915c3
zb369e0728edc621a049174622f0c9bd1c3a493e9190e4d944630957aa0f3cfd066b8ac74cadafb
zf33f068f62e2f4bf756dc2395df7b22a46aa45a08333650e110a820afde6a0048d0575b2b4bda7
zc4b7bff5a9c2e128f853bffa6116a4410fe6e562236198385875f25e23a949d091b29cd02e974f
z243cd214ff76f1ca09f121a72683b77c9a4d204deb148eb757673dd03783a50057df3ce92d5c8d
ze9ff3d9b432ac523e62dbc2ff5a217d3ce93d23e63c73fe30b5fa61737c53d05a0036b0090ddee
zac0d60c4eb033e5bc1b4223718ea792a1bb037a4f6d9f10e186682df475cc4f0ec4e1b72fe8d98
ze4d107bd2ff6e448eed8dc6facf8a93435197e589f2dc8893a22287f5f1eebaac7f5b5fbad9ccd
zdc7ce94bcbb2d3b84256b69998035e95562855d04ebac0f99cad4d77c221937b49b2827c32127e
z28a9adfd13f4262c1a735e2c645313daaab1b3ed2a7b165e09a37d08f8a5b3cf746e2d02db62c7
z65c0f7121c0590935d0b5058e038df7b492d983bb47a039c919625c322d7bf107fb54bd81fa9a6
ze8be516a382405e9962504fccaede9c0ab641700f744465c46a4f23a8780c8805ee13cd41f584f
z13fb7da6f3f854d0f167e4b4d5ac63f0ba1ea8624c76b591dfb1dab0c6ca6a9d913f73339907d9
z69409f2d1eb4c48768fac5fa319de97d2044660684804fe3e89f5d3a781ca0f23745bc461d46ff
z8cfc5188e42066c6e947e726f88ca11a4f57d5e84da969e2027e29ddc449ca046c2d303aa9ebca
z83aab6e39f0fab40ba86b29ced62281ec47d3ca7b5981f9c54bdbc8b75926fa551c4a63546177b
z4735487167db0c204b7fec24750eeecea762a07634b7a2a7998cab045d9e82c6d491af88283170
z22e64719191db0496f0052612ddacaf85d3574d1feb899163e5c9d563320aaa5cf7c27d57f80fe
z29f68ae753ae908e87c3cf269a467b606e7fdbf081b802e664420ed62335550e576fbab751e894
z7c99f7a7ddea640376b7104e53213318bacf22d7478eff367186f888da2a635872b40fff4f9517
zb3c35c4ce50f202564b286d12fb377d9c775b94c10249bb48e07f6828767857017548ab8284d3e
zb135f82e2f1563fc19ea38fec95c92f38bcc932e600292f97320f77aad6719b7474f2f1743b69a
z4df5e168f40a8d0abde281165f38868bd15e8a90a050b149858de57949faaec3d3ed03b43dd513
z40e5f92f3a569817984602bf434281ebe967b6c5eaa510c94e8a2d76742b89fda9be3d4d385b6e
z143a625eca14ac0b36c3cf1430ba177491438b85b05cb42b44223e733c8bf0c55d91e1f8f76353
z747a5d8afdd6bf6cd97d130f217be5b66a31d66eaf3ba1fd59bfafbff18a00438f90b003c79cb8
zfdee5d4de1e79a8dadcf3eb5ccefc653dfc4742e6675360685b8f54c8d76e14a53f4b9d52d56de
za36e53c19990c533782b1815fc8c3c767bed49457486239faa9ef3dabb0b01008632504fb23763
z7da6458684d36bc818190aa97ed2d5d6ae2da0519ce0aaa51a77c05e44f49b838ab30e5b0fd372
ze956592614c9487dd01f364ad078bc05d9bbbd3effaf57cce809fc79d556604f7ff62012bb644e
z4f00a413e2f184dc2a06d57a7db378b55903eed6d1a3ac8e9bd9b034278f59d244e191ff4d980a
zd87dbc78eecb81ed1974143c3830376994ae0698b4f4d19aea758b92399f99b6e19215d9e080f5
z09791af5135910f517350d25ffffc61ab35f2cbf25c0adf4ee8bcf0d6605fc4cec40129805156f
zc3fc2f65907dbb0695b5415bbd40ea5efa3602e730d5dddc93e9ce6fa938d5a6a09991b8b17cea
zd685e436592553ea578093d9083f2a997dd9a075034847e94045318dcd25313025bc5b14b26283
zac9c8b566e3b48631bbfbe7b8d7692f4ac8a00114098f1327fa668db6498eb07d4ec757164ca2c
zbbd65f5c652b775562af6f83f00f5770932e7edbd9023f6a70a7e34e3e8291079f5fec47f31d0f
z40fc05258883aca1b4efebe41624693a708378b5bcee00445a6a012b1fd6c7128132e9984f9a10
z5b30fd0b53eca606d205d50bf085217952c347ccf4516eb0318bd67f2df1d989c9087758284c98
z703f1a72f8c99b3138ea4f758cbf077b3d3ace383734e8e23bed1785533c4fe4b8bf3f45961cbd
z6c6842962b992eea409e514d635f12bfff694d524a4af8841ee9503864d90f8c2a983978990b6e
z73136005ecf8d6c9c04b6763226a78347071d4b7b3c9b88a5b32293dbbf2a4504d8366d682f88d
z2e68b1670c74fd58cfdc1b522ecb536298de5b0e141d1b1283256c9b63556a1d3c1f0ed2d9afc9
z3ec28d06fa8689202db50c52943879d598df5558911e39cff49e382518efd858383fc0c0de6ebc
za8e20d14ea15096ae14337aefe76a0c05fbc9793dcd03ca7bbd2adb8ac39382e736f80a19c8b75
zbbbd9cbd1dbff3e8cf05891a59d47d1660568a231509674cc265c382196f0ee0dbc9452aa786c3
z30ef1037c1e7d1e5c585726bcbe0783e772500073c53704c4b4e04165658ac80705fff40d54047
z6352d2edec9cf0204acad1bb79006492d8a4d5c03b9a520acec3c9d79870ed7197212453a77afc
z4d0e59503eedb1e22b0be50ebaa027481d27a2f1db7cab70eed12bffe856c7c2f434c6d103fbf1
z538d8e1f4e0d6345442c839b4a673110f9b9df5a4fe3a6381a4a34b343e133b80ac93b6329e00b
zd9edcf16410e3972f4f4cc9f8c314ddeab7678f689041622bf533773751ebfc576b4875ccbdb9e
za6384a1a04cf793208e223ac710f8aecf4abd541fcc7a4d0ebccf23573578dad5de2d377f2e814
zd369113ab7563a36b5b962bff7c08055dbc1f49e1f949d33b1ea33bfdb867d179f7917ef7d4599
z7f4786af9a608993bc4e899d8e36eea2c8eadd0f671f6a3f71feef94217d3639fa5049440cb695
z6c5832d64958a472255459ca0c1876bde15cd2bdbec10237035c583368f892f9545bc550f4212d
z403deed467abb09a2d5b32764b9f46c36416c78af620f5494ac966107f08e5da9a59e781921e96
zaf248a3c79e749757c76c58c80677b657e8bf64015c112e985e6eba6e3a6ed0f66b37d29dfa9e6
z84ffab64810c85ad1321aafcd5ca65248a42948c84415af86399c22a7a301a1ca8ebf5c4f5ff66
zf76199575e7d74fec3afc573f7c21bfa76451c519f7ffabab3a4bfb08e244cea4ac5a9cc5ba287
zbdaaf1453e581103be59ea58d0f479e54c44add433236eaee06a97656bf58db53fa731218d61c3
z801da6b835898bd1e74560e1fb337e1e5667dbf4a7b951396c57181d774e76a146085a8286b976
z7da70c3f611014f4239244deacf06e9f94902e76a76b8bbfdc89e7425abb9f1867807489edd26c
zbed1d04992556a1d7313e234b2392ff3f382440a431904f7fb9a10a31d3aa9fbd1ce307ca701b2
za8ee0f73cd8aa112b94272b8b08e5907a46d905f999d0b3a0f0bff259cf123cab217899a172ff7
zeb4b231271cbe42d7f36b0cdc7c6ce5e805e62da2832a6d3a126136a1b80ade39b57a8d5837606
z5eac1127b6666cb7f2e760132046ddbb764737fd3073bde6782add1453c6f65965d850ad98e3b2
zb56abe45c2a06a82f95d765e9acc78de7cb18b883f9c822b49b5d19e79a68f721fa2dc0013ff53
z4961dd1881c20cc73e21ad08289316b5ea688478724a2e41f5e9cf3e27a9c2e7a9b073d839dbec
zaa99a9af4f516d5dd761655ec057e4f5dcd0743cdaa4790a595c60551c90f424019a71d76c80f7
z29a04945b7590facc649c4e7f3f23abb01fd9d3e6c319a89a71f7b07a974871936c42b67bc5571
z6dd41b664dbb0d92478404a8f74e767d968151dd02b15cd365c0d8a074e21e29d6e52fb75e8a14
zca5dcb6702b59754c54bd1d7da4e8ab362d720771cc55487c001557011ec1bf43acc2f67c51eb3
z23be4196fec3753ae7b9b6189699ef5d77a869450c3080af00482b1e548349ed99a9c6e75a98e7
z5efe841e39fb4f3b34f4fd80d199a5c111f8331c1b0c9c642a541d09cee380ec5fb1e1e862c0b1
z34a6a92766a0d0cacd0220dcf7d7a3ec209884e9f8a3a63ee1b4a15edd9f17a13096a1c8b2ab7e
z611a51c7813055365287ef18b50bd53d83199fa7c3709161d9215be6a8fb5e0594040f89211a92
z92f69d114041d9ad62f2184615e07a8e5b30a661b7be0e46096ecd93b3b622ecbe98de4e43ed32
z41d74c33c48d737f02c52786e00af0cb01d7cd1eea27fce9b472afcb91e5fea0c60c22291e59c9
z7f2937290b1445722dc2ff4c9111d601394a7e28c0e7d46b76c13be7969633b5cd2fe7bc513dc2
za434d620a5ae626b43f7e9719b91eb78a00875c837380d8205b429efd304de020a0eefe0c5d84f
z2341313c06f933eae855e90f383861b6deaa5c2bb7357dde9bae8e3a152b4de9cb9bdac3c6e66a
zc7231af24f728a9b7752b9fdf0a1fa89f3ba95a89e1cbda5561b19963ff2274f5386acba6f97b9
zcc6dab50409930501f1b22026b4688e8d9347c4fc2aedcba6ceab1123f3788383340da5826adf1
z97aafb9307a1c546f86e01e7c9314252f2edcff35315061242f4a89b5819207e605e7f38126f06
z2d01b04df846533a8665ce7d39adef7dbce05c4b2751b5c71483e14fbe6dbad41cacea3fede2d7
zb51ea0d4bfb0604c525ae566636a9d6bf81ae88517a24f7b3187b9fb6c98d94eba45031fb46745
z09b0b8e74ec8984a3cf94cb947c484141c3d9868222de48b9d31eda84e12b2d64f501a85cc66ae
zfdff7e4c14a6ed0378cb12f6ff6c8c2f887027c6803ffe32625345065d2b42c603e607127ff9f2
z77bb036928fdf858efdff8bb3f4dce6f4b999180adee5e242299918d37ced03509231d072cd21c
zc3dc9894ada5b73df8b861c4339d6dbcd94007c33daf5f4bf1206a64206054fd1fda332dacea26
z15989793b1835f1c790bc8faedcbad3827a26cb540070d1b4327962c3716a54a42f53fb1b71182
z7744dbb1a531284cb604aa812bd7efecaebfe53aa6a721d05947c57e13f95e29afe7f9e1b4dc68
z6b020fb182e0219a3dbe84832b806b4a0c074f2c803e9fd95927e7949a43993c3115d0667b3d8b
zb68fd4ca75d96a80f553443d45074ee7df9ab33924dc5bd4cf5566fb573ae93bbc118c61c49522
ze91c7cb3aa1cedc7628b806accb995bdd744502e69951e7a5bbacef043431c87fd8891d7875d3b
zd3e05bae673dc3ae3aa667928d2b61f4048ba44ee0858e89b1f5ce7037ffae6951a3535dc00400
z269dd723817101df91ecf505e6bdb7ca1bce7726b64c63f043958b82e30f265b57470d1cf1b815
zad9869f567cdf2902ea3851b1d8d807db46ceb97d0b593f3f42f09a858e352e66a43a3af256230
z4fba1f41c0d96b13f3ccabd61f69f8ab47e299ef68c27f444680c4f35fc1d7a18c315682e147fd
zbbc7879ad685887c44d015de8c5aacd5c7951ef74f5210f5ba6608e87f75da81b4cd3bec2d935b
z83c96e9b9a2d3ac834965bb5ea4d21eff0b260fef1af9a1c1e6a0bfa7132f06e641f2e23097ffe
zd528db13f656400f87cd7377adce1aa8bc0a77737160312054c4bdfdc9b1ae11917731d4a58710
zec419eea13b3090b578a9d800b9ff5cab3d78869aee84bd53bf06845bc22900183fa566ee734d4
z3b11bcaf7cdcf7f8ff2c573602cf5e156dcafa40a984ec51b4951b6cd77abced0a46a82437753f
z0be57b61c278a6e41b24935b7acc99642d26adf4b0acedf2f40b282121eacf26a1df8da6f63a65
z935b412a5c556eccd326419fcb5f9fed0911d03a4a3f1d3c76cc8dae6dd62aa04596e24e9bac5c
z707bb522b816ff3e911b8003b5609905f014017b5b9cd895431e5f86021d017b94af87d20e1f87
z63697f63211f8936fe960d09e0ea7d51c353ec7adf3fc2e4b5d7c33bd07b0893f2262a0cbb0c04
zf61320fdda4cfe3d5055e3cc43ffbfd861dfacb17563af4abc35a75890dab731849fb558406a00
z2007a9ce339c32c4fc6e8c93644bf282110b74eaafb8b323088340a6809c41652d93953d9c93f7
z4f0ac06d499950427a70bff963877e74132abb22458d34c7501e0d5e5253d59d6797389f9947da
zc3af9a57fe5fa932225f4fe38a277cc7feb063b5229595e601aa85f66ed913318e4dacf80523b3
z71dff4276c14751177fd1282d1f413a56cf39a0f4cc578f79e3248e90ae04d152770166d0622dc
z5d97f8fc35b143cd97c7f316213276e50c54d22279271c2048ad5ee45afdab5bea6449d28a7da0
ze1444174a2b107c5a06f9c338d77f45e78918145532193472fd6ff8e482c139d564d10eb65aa4d
z189d81fc8712d4f5884ccfb9e2cc1786ea8e6bac59ff5d08f024088844cec1f3721f3f8a543b7f
z74632a5896cff9a7a7cb14d13e39004b09c440faa690b849e22533fc51509a779c4b38ae8ff06d
z010a9c9b708bd8cde6cbb5e790b9dfc201b9c11887f6eca765569ee6384e401768e4f9ec1b9d12
z61b4dc210ceb515a664e56e253126836172e2fcc5ce07603a92a0a4b6437cd732401bb3afb4ebc
zbc4039ee35d429cb684b3112e0d27b1548ee84cc3aa943844332789c6c2cfe0f4191c79e0cd29d
zc7ee4889baea01286c7602b932f2bdbd36a45aefe15ac12e826f3ed212f630f0a437956475ed9b
z4d066058ffe94baa926d5112b62d4c1b17c7672cb900c817433b65c4d5b8d8fed39ed29d07571f
z068057ce6fe0e3be2f065d13f7203869fdc240a1f7df25b53eec89877d82bf53bf1acc907de5b9
z5881cf64e6cbd5fde28e41117f49892a0218b8de542530b9443e60de99e9f439b62491c2e2012a
z6b77a52f8d1fd10060e6d1c2b112c9743fb6a2080a59eb5ac03fc8a4b43f27429d5ea4404c22c2
zc5b89f4393c1407041f3f23c2f19001fd97ba2dd7812a2faaf07812d4d02a8ff00927a3d5ff645
z37722dbc71d9421041a84d39b4fd81bb6c8fc6fb9f606aaf40edce2df45a2e81181e7a7be10cac
z695213ea3ac55c664ae5563853a1014961e5b72c26e33b1053fce542a54072cf94dbf5f4b607af
z61be7b7dcae5e47973621bc4557964addee9a8f4033d0eb11b652dd3a13c74e02e092e792696ec
z687c03313212c71ab8da4fdcf412db37a8a1c3a4eda1a2471762015aa7181450f2a037a2f81a90
z77bfce0dac99f7691c4f66746bacd4057b7ebc236b91019b40d71429e197870ca69b89892b4f88
z0b2c76377cbc90b6f3f7f108da738acebbe5e30edd34b33ece1cfbb28535f0748b9a712517e0f0
z5f5e3a8d9eba7f613d12898f2df6ba788cd8b853ad28a768df76b04a39712804a7e7a4ab64c697
zf2bfd97c91973fa75df52b21dc9e54c3c2bca2a5afec332789e9290d2d142978be18b1747af706
z6dd04501e06387d1a9e6eda464012b51c99c5b8b70fc7fa24c7ea6b150d66a4e3b617c1738def9
z8f97da437f57ba43a15f910ff3c0c6f1839d78c167b4a872ea20e8e9ae8b6a9e9399f2b1150b18
z2316b175819d2d6c031c0f55e4031eca3a7b7e0419c096f4815a892c718c54980c044c4e3c77e7
zadc0fa851dcd03b5baf43a1873faa0c061b1910a3b0958715d40426a09a608023a967f47b1c301
zfdb0ba50c18ab4f405c403fc8596d9d63e46dcc361a3fc8d6c91a5e83346cf9232b52196040206
z4a80cd9838e819a6e759a9b2c3eb376ff184e08a60cb7d5e2f279693182351dc552a47dff12ec7
zcc3c45318418907cf4a4f604ba15dc4dc79d4667f4f8ff9b2a81fe9c11ce041899fcef1dd33d1d
z441aaa6508e72d908c0d09e25b0a66bdf47805fbb4d4d990cbf5c2477507c4c9df25803431f3ef
z0d8e22dc53accb51364838506fa5a64f8f108ba4e6bc02ed986906a351e30b82782e9e6f9a0d63
zfdf26cd4cec8d00f84b9ea17af57360ce513fdacac79715dddff84f6ffb6b8a6ebc677221aaa69
zda9c957ff92c158205142c3726f108653701d33b9ca9892de525ab9feaf0ecc3073feba37e0c48
zb87c3b7e12de61cf0edada00ced431d2e708e12468415809f6d95412394a72ad2c15732c22ed0b
zeb092e1b2f881cac23ed042dbaf02e0d904cdf80f0966d37e8da5eb67b8ce4516819585397a6ff
zdd1108716288ab1255891ae316bbd4494e2bde0ce0a96d8dfce81f6de1ffdc93cb08057198cd58
zbceb8d800213f908b6877adf5ec00b8594f26b0d7f2932f8b5efd901067f04b23581e7fe6c063f
z1a161098b830051308e7c6d045f2030e23793a2863c8ffa5dcfaa28eee303b749974f6b8b312b0
z9afb0ff1fb46e3225f382d649431cee47c33942b4dce258941d455bcbb8b1544b5b913c8a5138f
z40b640996441a4eba2d203c8124fb48ee30f1f7c07fda044771a95d2d8e4642d8a8b8afceebb22
z2326f22839829615d9b17636c849aad7f53e0d805c816c81111f804b71182d0b74105c1cdc5c43
ze80049ab507773201e279f50682ecc93ed8f70f25a5241b7487c5bac0b270ba4d1fa5809c661c2
z9a9dcdb34f6f158ed53a53d21691988d119ed9ba7b1562a8c08b5edff990cf538a131beacfdf29
zb916477c1bf41e37fd2c91bc07b51441db23a99c7c79f3c5292dae69eb75136eae00eca247d10d
z724a9ad94f194aeff65d9ab992315a7a495c329195fe97cc3779c8cf5bd0ccff602da83e9e46c1
z3e767536eadbdde0d34c0633a425e02478d7ea98585079f04fe0f486955eaf548c670b606333a3
z6b7be3d53ae8e3b11a9ded90f9f08a29cce53f598fcf9ba9b2effc7176f8f87e8c3b5e5e02a828
z49118bef8d5654c48a12745a70e16605e5acb64680ef2f3adfefd0d17f6238ceb0f8c1757b34b7
z97034eb38a0ba778cb5c6eabb7d2aff256d729ef241ab784960a3ff82d6a9912e5f2e3df232160
z5055b6c09fb3b1951c607559e7d1b9152f4241fa924f4d9e2312da4c002d90befaa929e8e2eda7
z317ed537080ab9cd98446636bfb31f4c26a8c6d51fe0841ac2dc347a8a2218398949c527946811
ze6e479b77f41206971dbdd35d2a211f8e99daad678e3342f4080cc5c465c2e7f79cc966f4885e1
zfa971a9370edebb08850c2c3ce5c89cc7085bf531183d7ac30fa165c3a171c2b0af0cba35d6f73
z22415fafe2a1f4ba27ef6027b50aa96edc85fe3c45d4b91212da57094b1e781155cadc5e9c28ec
z38695e396c3086d2cdd124d10781daf3fb965dac6702ccbecbeb3db80193100d51dadf14dc57e9
zd2d3a8257e8cdba785e3ee09cd586f56af9fa17dfce70b486b38b6448430db76841d47f1304c8b
zd478a87e460c515103386b108d152371091d59190d9dc7a38fa08620acfc4176906cb2a23b504b
zdf59c67784e55497f4c9014ab70ae43f12ee8415865369811e141bc2c79d9e361421d1df9acd53
z354e3b1e56604a8217245a8b12de8674daacfcd177c6d803fbfdeeec87d7251bd89fba12457902
z6a7fcd2b137aec7423686695f588d51477d713bbd0073f5ea8ea8460693d638a5434b9212651ee
zb9187ced98e09721da79d844ac1f4f770bb8e73d22208df57997820c25ae17e6560261ac11da43
z870a4040aea743b97d44e9a8e0a6a83baec94fcda344f01509f96627ca930ebec5937d1bea34d3
z92aa7c1db295e400e4892e02703a4c624ff50d219a225669a9b9c0ffe550a372b638f11c6ac52c
z4d20a392cd48b2bb8a0f148a15ad7b2286327cf0ec7f521a0c4a847ad77be3252983d6b71c72c8
z60e7eeaa85429ba770d9db2b3eba7526a6c033b9ce2ed5304f328d84ab79dbde8b1ca363dd509e
z1a7aeb0f12a991227e7ddf526323a45b1f706903550752fa2806b4ba662dc517191ec86f5dc9b2
z60285b4aa0813e3bc21242746f66a95c5553a05d963b8b61c370a791eaa3608fba9c1b72cdc57a
z23bcd42349bcad9506a7f836a1d6fe7b01e478391e7192225abfb67e9dbcf0c948ecf61ce7f25e
z29087dc5f4a427ebe3965ea1d3dc4d0478f93f23599a34837366cf7923f8e77fc6ebc35198ad32
z5c011b3a7bdb601b45d44501409705d9a3a8f7a92fc779b4e4ce862d18cbd354ce1d94f750d2bf
z07bc2770b960c45ef4e778f7bc2e7baef9845735980f125d60688236c120fb440adf16484bd6c5
z9c88a86996738697d2f18792386543fed5b7c43250fa71432284e3e6a9b927c59de8c8c75772b4
zbbfb812b98200371affd4bade461dc4b8eab570dc3d4e04ecf2abf712c7f2bb494481c674d6710
z1350f682011f2599343884aa1af0e2679f4f2290be55607e1428208967b4265ed35c7d8bdd3500
za7d583ea303ebe22dffc2b424b6ef79bca0609d820ca74c70ba211f724648bb3f2041e79ca274c
z5acc62a434a039c517f7f0f58cfbb936f8ac89645162ffb8c9ece26bb53b61d81c26068b547c49
z053e22be5d398e3c0d858c62603f77b2fd6694824fd99ead0d3f1742f23384d746dbd3eb9ea662
zd79e7165cd7f7737b2504247b0d1ba9d3e046ea5c7eae6138d8c1213ba12a670529cba44742e2b
z00e7ebd5fac78da48e8339afd96b560558845303d556de12094b3cfab5c590931b5aad67890b92
z8fe586e1210c261a964417d1dc6c51678b1942b877d92337a9a454d54dbe36d0d3b17bb86cb226
z0ebd2c8965bfb845bf71868a2c1363cb2ae131300b1831d5fa69679f75732a612fcbc9b69ff28a
z97f2e9f11d2a1ba7b71e16c0646344ff63e3c23f42e7c617dd91902b69726229dbedd993f03f45
z2ad1ebf472dc1c29c41f242dbaa1b22992c6424e751118ed7309b3f5aa0559eff93a3873ae29ff
zba0bbda840b1089adfe821d31261f64125af608c0b5778482fff7782a2e6ac512f0b8b40280baa
z29dc6acedd0c5d0e81da5b8b95939681d2f004a285a86d0a0ee6fb9ef9e747d8c5899a1d8936d0
zbd03982bc4cafae916c3c15417958eaac583669876516ebed03137ae37e72678d1ef832da7fe4a
z8eb73ca2938dea61b9914b02d905e281ab9d0f1f9eca05a1afeacefbc4ed0d12b32d6187a5ed01
zc76bad953adec860395646d12832cd3f003b8ab71551bf567dc0f9599e3b944ec1e7a39f2e36fd
z71643bde05a6f94b53a91645a77c1f13bc94eca49eb721c0af6f45ff0c3fd9a0f3fcdce2bb5c2c
zed26a0b63e4ad2885ab721ab63362d0d6ad83b6f0d054cb005eb36f744eaf3dcec0d303332cf9f
zdf3b6b1eea6f88a9d0571045e6e9533ed43d12bbb78c367d5111bb60d9ac84ca553aef1ea32756
z3eea39b1612c55b64511d89a553265489bc893770da1fbb6fa224bfd814adf6b6be99fdad980fd
z0dd94c706d132e19088d3b484409af52e6bce4b90ab820025f75e2267084b9fcae1d6ac80a9dec
z8f932f034d29ab337e41f5b5620733ebdce57a2e64c180bc7a93336e6b82ecad53d20da862764f
z466be38099042d7bfe8eb833cfad165d901b3e6788fdcbeb3324cd934b90fbec0908b523972ec4
z64db6ec2c162d09b31fa912bfc86c20cddae68b9234877162c9c97dfa5903ebbffd47f5ab2e33c
z1c864bca2ffd49ec09994bcc31213e09596ca0b25edd6a145b19d5d35d32287908c34b610ff649
z35923a8c9d1123c2820ce1244a3bd1e356f574914e255b5e3f72baac03c9d5d35c7ae11d9e2268
z04b0b21243be3c51d18840521bc497bca496a4a2dd8712bb27803950bbbd2ac893f116fb300c97
z9c975ce4a94dd0e60129d447096f74996c58db20f09ba833950e8c3f1dd29e0ae8c5c9dd18ce0f
z0dab0b7decbc091087c3df192c11878ddbe993e6207e50b6a2973c034a04a1a67fafa5784666a2
z86f704039f23eb6e00aff55beb26d0f47463769b6f14af7adaadfc350d19af9ca267978209743c
z8028d256bf5b9baa355fc1adf062dfaba8c99440f22e1950e7df12365b0139333c38d97536d779
z6cc006a5b5557c924b52e95cd9b130d45b238000e6b50da57eb4ade65731934b6f779c464ff0a0
z9ef1329eee04a8619f0a6b4d61a27df59e7fd32b8c79a67e87986d6239923c5ce0060aab94fc1f
z9f6d52b62c5be82f2f29cdb1f7a82cb503306bb54d48f9b39513c7ce3eff42673e5f6c6aa9b80f
z8ddce5d76495ed6f2b0f7c0ef90a51f12771d953420c3ce38855608658cdc98bc36a1bb8e5404e
z0ee9ce178c07eed603c1fee6220350cb5c2da872456bea8800d5cf6c2677111fd94826bfd2aa44
z3418f9dde1a5a8293c203812b499f2c4d6a1ab349d34b17e063082cd87714457a2f5dd79c94699
zb3fe16202c7b041f3cf4e9a2c282613f903c2dcea801359f1c2b364d28308fe10ba22dae73b0c1
z7d5cd6c4af99e40bae2d463740146a4e20c839c9e04c9f7a8738f8d75c6b30da874f4866a78f24
za6ca78a2685c9356b2058437f1e9376122c089a9f9529ccffa6afe2e8eb7eb8291e6ad652be472
zcfab945cef663991bb3ee42e6cf1bb39f7f5a459ffb8ac23dcc6a0a84e780478f9d81210846179
z860efc4b75e01d3a1b5dbc3a69fff89742c923eefead6a00db30a03aa5b1058b8caf8b8db491c8
z716e9fe356acb30427d95349ca5dee9d7192aad80eef05d54c7eead254b14c5959670b7bbabebf
z885001d914a8557ba17beb6718952308a8256dde8886719257463fafe9ddcf5a1a5fb2b18eea08
z9758556da8f24ef40cf7f828a784daccd97fd71e41e7720edefd682614653b52475b836eca3fa5
z66696f66328d31c20ccc130107049b9c84c1b1a42da714a6c4a0cbf0cb3494d41a81f4a12563f7
zf9894373cf97b0115e014f0a64144b8d6e62836a11ed3be8a89300096dafb1e56908968a379ea5
z869a02632966686fd5a3a3bcbca3de29d7df0b702e565dbe6a6787718cbf321a131c51058b3e8d
z4a0f7e159e64fc454f634f05bc3b01c715089a9e51c874b489d194513da5e6e682709ad6c3b68c
zef5f32828fe1a4a6bc6f17d26dd0a5070a952950eb06ff931c3a55665e7d2d33c71c3f3792d02f
zdf2361e58ce093a3920c527b6d9f1f71f986cb42237c856ff0e15852603af2df16fedb87292d5b
z6f82705206be89ff04db4e36bba414f81d1adef34c50243f5e9927e3e1f0369830a1cf98d9d33e
zda34aa7da2a9248412288894ad6132be10b9bb121de3850ca93a40baf59d1b7f68d127c93793c0
zf05bcea0e2382c8bbb0e99654db9c755bf99fed154683dc574014e44e32a9004460eca37a2c589
z88825dbd9646943edaae86d812ff8445b55d42b0362e0ddfe39ac420a68bcbc3b0773d1e1fb822
ze06ca83639f134fb9bc215b5b649ae0930c5910dd5787a70b226d970d99aa559e58ddd402a837d
z0f2b0063f159e9b3fd74c1fdc7875a19705892fff055eb3b1ed79d3a4b39074d31674b69428646
z52e5f38de81f74dc1f10c4d9ba0ea0aa2019ca815eda55c227ceb46da50b2ef0f3d80b7d1464e3
zf45a70c7be21b2aac9c12ab1a42281e8560f09d6e476ab8175f0d576d389e3aab4cabda816061e
z2cedb6393333d6119f37414ddb538e3a4409a4b6accc557ce6e7fb882c5c222043e160d359252d
z2bb81e8d469292babaa1df7375a817a84aa9ab1684f2ad1e8e2cd06a091b6937842183d4e76f2e
zfdb4029b9b99220a172189e37522827c2a893cc998177fe0d900ff749966d6e6ae9e1426563161
z00991cd5507fb439001a8c43bba106ba73b3f82bbe5c11423507e7c62219cb501c9b9e176d3071
z208581da68c8fff23088ca9d974747f722d15cd2d25028db414269465f33fa268d563aa6155bbd
z5cdcf3b37f50dfadf1f62f0b4de80d0ce3d6d7f1a50d4344cb77b36b425a2a94608b730bb61a14
z52800c00546b8eb8ea4ec28cbfa9c355ab587c582c51df8b21918bcde65222bc3e87be07b7edda
z5e614ddc0463253e778f719ee03b4c6ace2f894ace530664d18c262dda6cdc3b781ac2cacd262a
zef7903a2374c075ca8a3b99a9014713c6b11d0c7a6476b214db4a4905d8157ac6b763a9fb92076
zce3bdafd62ee7c6531dafe46d122e4f180d4eb1c67c9e8d486939deaabfa0a90a1f84cdd3fe0ab
z2169692807fb8d091cf3d4d2f536653cdb84c69993428cca7b844007e06b970c1df6469b990b67
zdc33806a5e7b9a7031a9ea3725aecf03080cda8cf0aa27f7bd559d2b51d2f444e1d16e1a9cc1bb
zb7a5b4aa73dac60eb3e5b5055073ffc6a965111bd4a1b0b4a6ea954547d16bc78bb138e67b152c
zb141133e912990e15c5be03f533b7774f38e138cd1cd87f2f792b00d2667d079ebad29137c997a
zcdd5765eb76ec4c9b24cd12a6dde963fa9419bb4bcea9987d332520fb32616a5fc87ed50d925c5
z52684bf736306543bb9226c9f7b69711e4990fa2cb22fa5ea5462507650d87e8bcc0d99aa8cc95
zab6820b2674a7c5c8195ec6ed957a871c5a84b2bf63b9c053a31359983f50b5aa8aa2d76b51276
z6fbeac7539ccd17a59e1bdb3b5cd21c6cd4eb28ca8c1a691a4e185d7e2c9c6b2dfc12211e1fcb9
z4a02b4dc665211af9d15f40ac131c267574f398900a8744c927c68c27d8552190122b7b06b05e4
z10e17dffd71667da562d8968de0a606a0983d3f3262cc962befdb7b26b9d51b46306ba9ef4cfca
z3559312533cfaabdeb69305ad04b0420d5e4519f8c0ac8432fdcd32bdc5d509f06eaba5e6fd5e1
z753828b0856935c468d161f212f6ceb319cd8cf1672293693392cce1c5c0d80a94ca15af929007
zddd250bb114036a58047fc12f371b06ae16bfbcf4fc2cac0b900d38915e88fadd159b002719906
z3a2c18a5b24261bcacd368341b540c27f879f6265614e6770c9db4e4a4afb038b4b6c90795223b
zd9f7596a6afbe24bb4088aa09ed5b5387a2005af5603365a2136dec7538be89cbdd555a0af7d9c
ze5a2243d44569b36c9322e6af8c4ed5f58aa82a44657adfd27211156caa2d6beb5565b112fc7c5
ze8d18dbdc2c5f1282829045cce855162aef33b461c6427ed03b20acde670aae7dc7d4f5c4e1939
zd0e878c8327a3ed4aba47025fc19c374543fa42917cecd76458befd9d36770b2a656b062ed7331
z618900064e0e9044e3c7c58e99b39cb1e50cc971a1ce64a21dedf041c103a2cdcfa14803f291b9
z1ccd9707fcfded740b0ce20d7ce856f8cda2590280e1a099b606b94344d6922bc8206accf9e918
zb3d5d0b9486627105ce9a03f0669c987c8002972f812881bb0660284fe4d224867f94a711ac3af
zfcd99cd48fc153199561c7f39d98481ba1786ddbb310047c52608b2eb680c93b22c06df35e749c
z07b1c55cb2a74564a2fc01fe4b25780e81df28fb440492235628cd4f05297ae69d519b6725d3dd
ze73dd0d79563c88d7a6e4339088e0ffa723e78ae6198cd79f34e6d1a56edb2a1b6fb6a2e049a62
zde8181e6f92d5ca365bee658a7b90f2e2a790e4f45b49efe95ca8c5db56e6b333453e071aed34a
z1a9449bf62a6fef1db44dafaeaf09be88907f88283855f15c7a6e1f10ec289cae80b35f2147b6e
zb84740cf705853c08d9d165f8aaa4dab71bc418051384b5ac6953a7659b566f8c9e10581707003
zec0271ad30b08d8acbde1e28bbf3cd6b8feeaaf83b84c905fc926687c7aabbc19d978c1dfbe65e
zf0148ae128674bdfd311c28deed87978078f8740b655564579da5a51b5ab8913afeeff860f9be4
z776ead93c90d5652f4ae90e08a78d338bd69825479d86e5a168f12f0e4dd29565f2f43305dc4ff
ze1e1485f7de92d1f1755fca3a296757297c85ec1891eaf6491b0878dd00e5912ac9ae60e2c5e83
z55068ad2dc7588a219a59c76c6b38d7d9f8e8bbc23102cafc4d3024e1d13162367e770f7539581
z171382d808e182fd73a13a549f4115d44d275e1cc41cb90fdad5cc106c7615880bf627c8047e3d
ze0deac97c67f0058b66d8d4aa74033ffcc878c8d768fb8644be81bb3b3df4a3c76753fdd7e63df
zd95f152f5c1afcdf6ef5e9b16522a182e30b66d428b924f90d1a948db545a3a7a2e6e9dc800218
zc8b9b084820a07f3f0b80a2704211bf00f1196ff3b9cab64d824dca042e24caf73916b6ab0c7f9
z5014bf0c0b4982b39862966a889e22313629a022312db6adcb8bf86a03842855211c00a966602b
zd6cf9c347cc169458eb335a506dea14f04899694e7597285861c2e8eff98e89f28b25c1fde783f
z055b8c3c9cfd3c1d8dd735fc4332eca04947c9f170cfb198b7c6eada963893deb21a5a1267b31f
z3179ac0b0a15b6269cdfb001a7b8049029c5feb0b96c5eb592d2ae845066fc780d1dc3a81a7437
z839e5ab8ba9bdab02b2274992652d548c0649b3e6b1fca28a5c0e5a4c0f9385458e9ed02d578d0
z143e1ed051978313e544275a85e33b66c16bd7be038b821c5442df795fe5f00b8cbd6f321637bd
z9b07a6f12bba8665881432299e6e7fa30b78a8ec4243662cbdd92307baa1790f60be6dbf84eb3f
z768a87ec41db46c2831f0c5eddd7dffde20dfc49abd349148af2128546c06b91fe1eba268b1aae
z431e52a3c3ccb4f2604711cc8e0e6f257259b1bdb2aa83c6a3fe83a67c2c86c42520cab493ef82
z762579e11c52dd1b9b2c001cb52e7465735f5918da5b6c0e8b46773aac8a9256684d6953e9d48e
z53c200432a1a4017845da988b90dd7cd57275306258a9a8cd3861cc5fc09e9d6772aaf879d4a72
zfd408dd218fd5cd67815be5d703efcf66474527a7993d5827aa595c11cbaba62b9408823a411d4
z73aeebd416da51e31bfbd4d1757ae37ed080cec9724463d9366401249f4180e37ac7d76f94ed3d
zf7ca2b9d13fa4e8ee3b44ff41cc67b4e40b6ff66d9c240324b0905c7e5a4637c82758ffea6d909
z0215c1067ad87f4e3f5f7aeb085eb682a933e43f0745222fc9e74d05eafe61299a72fca164bbd7
za70ecfc7a3df88c3ccc0f89652d092d213a7811f3a099107b95fa194eeb03737ab7308eee889ff
z8996a6b26e805a350dd7f1f4fb5226e04603c0d36ab5c6e8339025a70698615034030f87c7ba18
z3ea4bdbd4d1686a5b1aab41df527b8a98437e3fd5c5466da2af21221771593213feac4bfce68af
z3d4c4e22db6ce490d89c8c40a2d04308ee730ae4b320be20c910c72a5ed0839885240d1caef72d
z81e1bbaf0df72c2d6483f58238568ee9ed554d99247bb58a99ad5779de1f97382a583d9a9ea1b0
z2e7225569dfcd286a0a9b1250fda1294540d8917092f2ea2530ac76ef223fd84ae455779c04b71
z750c27761f946bce26d9c07e4e6cc5821cbfca5946927b205ddb049729dbe32db0582f761fd7db
z6a519d5676fb85cbdd1000ec962c536170f57fcaf995666e783ba62b5fd0ad1c95ba8df385f002
zcc667ebeecb8f30a35439d641892ceb10ae48838bf2a361e57c5cbd5e9903fcd255ef3152adfb5
z6aeaeef356febda625386c8d21fd20827df55225428bdf51346ad2a64b37ca8b25047945fc31b0
zbbe6bd0a6bfe3a3c01478c6a432585c0c3dcec778b5d17eeb0c56496c3855da6f9f810b7b7f39e
zffea200ed3c4c3489c5a636a845e155bc6086b4e7a567347fde50303cec9fc060208b2026e80a2
z7c6baa6ea32de95bcfa4cf3a9b585a9b8eefff762baeb9d713efef22376674b6e49e61c5e1585e
z07144538be6d515c04b0c4025c9d76d0f02ae05d7b806b9fa2a707b34ddae90a5409830b2564a2
zef08d8d715ac5572eeb6e8548ac660f4db5b5fb56b64b0c26b2c98ea96b0423fedc6697c34bc73
z0e4e6b183a6c4984ca81cd232cbf76b5b963a4f83ba47de3cea2c71c65227cdb62c7fbd96afe45
z1b41b3456064229576eeaab362918a93a1262f5cc97ed2c33d4e78017c033d4e4bef2cc6bc57a9
z26d98c74abf110e4f89984fdfff8439f1b36464ee1598508b71f19ec31e026b0aeef2bfbea6c28
z570f7cd54e24c3560303bf56ce796159ae14866e12c0ad9707206137587cbb4b277f819cbb0cc7
z76a45d07332c486cee916c01b23e73940dacdcff7a76c0e46510e0b16ea5c5254e06e4a2042e55
z3ea302ecc0f48aafe9552af8c7fa8289dc48afcd5b246b7de0944bd1b73898769eda0eb43b2181
z1d29974b7ddc7339e7dad9f6eb2cb8083c4d0fc6c582b188a9abcd385b84158d85a6f1525b85be
z5a3854ab3818975fab6b6c55559ef9b51ebc8275dc4e4d25710314edd7fdccd520c72eaaca9c74
zfdf1dc3040320821ccea9d6f46294c28d120c6a9d0c98447f27e412439317136f351f6c02e5372
z3fe7b023d1cf26cbdc46776c2e0f5b7f970941a7144680c9810b2d467402ff63cd40fed0a56617
z3d9658c029d73a1c8752b42613d685c39efe38370ea0f457aaf570af75fc632c67553e48669123
z206796c5865d226d93ddb18b58c7809bb0a105ac1b8a4d12ed4d281f8fcc53cb1f6958fd4a7468
za15ee5f22ae7a5abf1e680dcaf90aa0d085eb1d22d76a5466ae33c4a1bdb91ab226419fd2faba7
z59dc2206c20a249a7b0e07b53bd55a10e3dd805505efc075604c95dc01ea762985b0ab5fc1ddec
z8c544a22d1597591419a34c07a176ec7c306d4f68800f9ec6ede5886f977f1cec152e17d6db139
zfdc514847823cb0a4d8da2671b936d43e73565ca8bfadb60ca0457236ae1113cad5ffe5673022a
zcfba9af8b3a26d0907999b4c0bbb7cf3f9238aae906005f79c6fa6ea56334bd97f65dd4118a141
z222e59d785881a7313e091bbb3b7c343cbb669a3270eaf5183bf52a13d31912c570474df81d8e9
z5474ac55dbb2fdad002db9278a2f108aa1cd523819e9a6a13ab3e6667388bf8968513fc0013288
zae5a093e47af39c5f4003ee0c1ef3fc03ec45d160ddb226d63187288b606edfb39766ee47f5131
zd1314d1d7f5256c108373b052f9ae536c1e611b3ef754c58be6bd7ecbfa6f705c6f47d8d4c9546
z200d034d4d55634b8fba30fcc54604e386c4678578499f840431fd74450f866097136fd69262a3
z7ce482072b869b0fb75259092c3a82f78413732257b97233defade7742394fa39b9fcc928bbe28
z4a914c18388640ece42490605107130bc61896d54ddd83b0adde91cd36f270c4878a6510296865
z9cea330c2d083ec4c35cf487737774493bf9681ae884bcbddcb5215629ffdabda1d47c45a55d5f
z21a869eb2d1390f081cbcaf3a0a61a0bfb2cfd0b3c6362003ce0ff1770ce196a934919296e3875
z058f6724a73b904a0359352b371f7fa43282b6bf92343ff65da5f3f6c8b5fe3f8829c9781735eb
z9369032480169534ed591fea6426cba39888e98185dad1e3049084caed655cda0e5f145ea9780d
zd8c08f3e88b959eae0a5385d7fff0c632a7ab332e4b08483960befce7312008f0bc7834e904170
zfbc215bb59b9289ab748f7b67c67584563da96844ba227bcc5369859621d78ff13aa727beda983
z8b00aa3572719d9ce9178a033532291542ab7b2e1af75e1be5b7b77999c7309be22bb371658cf7
z300d91586fe1646d6df047b2bac7472a61ab44e8751ea1b041ec5d22c56c7280ba768b01e40cfa
zd27a390e813461ed619309a845d9342f278a3976c3c71c636fdbfa7441c5d30e7f0ef9416bc8f6
zf4a986b9c4c6032c67328f7da4f9ffe16b4d6d4f4bbb13ec9fb387e329779a13b6bd5262eaa2c6
ze5beeae62eed381daf49fd939675fdb1bdff9b1940cd02c6433a1c6b067e046f7b3aa742e9ac92
z5c633eb6fe0a11857c759d5ce2431717ab99f8b1e862e198161c1eae379f7a61cde41381808613
zdab2f6f534c9dd7b0e75f4247f471dc3d27207e7b5a52b60b2ad20db39ebed331234f91fbb394e
z0c66a71852f8beedbefdcc04b70de6a86257969092e97f1db9f553fdba562708dae2b7aa14149a
z6df56f8e8f8718add3f44c04d77ddc016f51a496469ebabc024c7852498d478ffab0ba1f798e09
z169704c040f534d0050e96707a29dd12f74fbfc84a7bd3d5c2429f4e84da74f50177ca0aab7be2
zb3828af71a5a8f7401789763cf96bd49777fbaa2d5888ddcd73ef86fb1de59d85eac1c6a835805
z4e5fb455edc04404423d6aa126e98cedf1b7ce6e4e73b9b0c209cdbab7186524a70dac952b0b74
za5f84e6ed0aa8d69df09243ab4d8e5eb424e0137c311791f1ff500c1e2be4750b8a091158463ca
z9cbc49f779a3248264b393539e91fe576427c05180aa880685f9a9d34aef3305af279f67d42f89
z8a0dba80f8e89866359f78604a9ab6ae67146246e1f4cc9ebd36529cf3091aee3a488b33b35e56
zfaa7f9dbc0aea40777ee5d6f200cd5ed04075836bddf4c0fa78b499b8c99322d6261d193e887f7
z15c4b1f534c899fbb12779dcff3d8128dea078d421306196fb9a576832599b4895f1bc1cf065af
zfc4d43f54e1c9a6da65af07b69a5454c794fbb9be502790c15bd21ff6ee9463e30ed442ab3e1a0
z0de416beafb738faa84e3e6c0ca11261b7386a4125d65be1d3651ea2fe903de7d47136762f94ea
z2c28aefa4b72d350223576c290bdf418ad54953e1058f8fb56a8dd9889e008ff3cbf0232505914
z42de5f325f3477f5ca58a204304258a24ca5328d0be5e314d325e2d022460cea3b6059fd91f4a4
z09ce94ac3d249e357a5f6131154b11688a208e3c8f32360cf51825ad00454073fd847433fbf773
z770918a0aa7f824fb6dcacb9b2057a8b9cc880d9e2a5df547cc81abff189e50546de112d3c129b
z688cbfc609cd62029bd777f1ce5f20f90cd3bef4592835d14ba93b0c06583ea86ece40ecfc02a0
zde6cd9f67e8150cd943cb4522f082e7ffe3d66055236917f742652233f3d923f5c9ce525fb18e3
zd9379e9739476a9799e38249cd41a924f48e3f721177d869251fe7a17697179506e14df92d7427
z43d3321ad58d2a7308caca4562b58c2997abb7b4984fd4a462eb9c4481265abe6f20b5560e7b7b
z58cebc4b6c37d98130f15a62874d2f1e205aaeb589ebe42d664513627df22b218a8769a3181a36
z03b59679553cf315c9f03e3faca60c3a91c091318d869f55a322822f78fcd3abf0caa9698be210
ze923918fb6b0a83f0d6cdb258240e00f6f99a2e165ffccda04447be4f7d73f8962a829407fa391
z276901f303b8891956b5205c9a51cafb80238aca993825e35c8787634881d830703f18cf45795b
z02308df08596e907184f2ed85cabc6ea9140041c3f21bae8f00b549b5d29929cd362c081b48d83
z463a740dac381d45c189f143b43355d455bdf6164d778cf972ce62392cb5328aaa2cc759ffa55c
z2ddac9266acce7b2e39758492ca46d100f27b6931f397cc9fd243249d23b9095337bab982ecfd7
ze19fe9b7b38b978166826a208175f632f5f2842bbc211fde86e3ba690116c0320617b1448ffa8a
zabb4ea275cf3a26c06200f839bee33f7be4addd4ffc0f5fcd447b1f53d3edab12d43d2e2448f4a
zff814df364ea311d0bd27ff95e508ac4fbc24e95983ecc6da6fe3cdbb3de8cba7b62e03fa51ed1
zb5599af5d692fc5fb79f98f89a3d206f04d4bd5b024dace0dc12c2f46d87463c12a1a9cf66c0b3
z1858e596bc843b7b44b4a14811d04398e33cb923717c88901a260b5941b592a9f098d44cd00745
z5632af4714793f7501869e50a629922ce9cbd189fa73933a530478bec8931e4ad4acdc792a47b1
z4b3f6ca1baeb6a0fec69a983fa5dfa02966b1a06a277317cb17173ae8645043648263fb6138ba5
z25e8c1f7a1aaf8f1769a82672e893057c08378bfa542584fba0d4e89f9bba38677145455165830
z0bed0edfc17140e126590a606453d30ffd222cc74a78a704f0472327888f9f4cdea1aff40a7be3
z8e0299c3c7104b3020d4c32bfeb531e2cfeb3509aa641ae313ff6d9979b7e356f6b97d2fbd7d1e
z0c55153366d92616a575b6b9b9ea46bd96d7f1ff36d9d2303080346cfc2ef78325ebac48a068ea
zbd1a5ffdcae0c8e89c1c17d8ebd7a97ac5cd35ef06433f8489ae8c70be80750ae7cc115fc4803e
z9cae531113f0115c6d4f6f3a7056ada178f274769b827052798f96da63136797fb70973247742a
zdf17160a0d220b43617351246482b212a51e219130b8c5a5fed38f277d921b643249e4e8cd37bf
za79f3e9acfa97cd4e39bba093a6b7d7bce8ad77f650fa61055f5135b82d1afd75973b5e273b18e
zed08c415a0a53db16e34d48b004c179dca97ee10fffb9516dee06d12890f0b3245e88d69ddff98
z64c103a45c7498a408f6cad213b69381936c6343fb73b25da0c687772ca38cd19f5ca7219dd936
zf9c321ed6ca68dbd9c3546675fdb4d1a8c4945e7277f2fe302e2d95447dd996f1036749c74ce7a
z2877191007439aa39ed76a1df30a29765bef86c7fff7de8c4f7a2636f4e47d98d846e7e0d78c01
z4ccb5e0516fd7f8a39d5d23862d3187826cccd5fedfa31f50db46cae4fd2ebdd770af83f4c4418
z47afd54f64d0fd01e84d7c3ecb80f3edf3c793a083f8d362fba1e899192ffb7d45782d1a72be9a
zfdb860199e6d8705d6890f80dcd3a63722fc52e2141627ef4b25076c8569450cfc9dc0bed362d4
z5f87492d95e6ea578e124ffb2029b386227748caabe39f9fa9aa55d1fc3fb8efe4f4b44197918f
z70eff240d92a9d81f542ac73e415de9a6b07d4dfd28219f5a23bcdc24b5b502c1c6eaeb86ca508
z357ade135dc9a8102deaa64695728fc481a309564ecd69e9481065d0f117b411eb595d58d7297c
z468367896b81842bbfa18fcdd2cb1003b4c0d59ad24d283dfe16ece90f19ed94d1bfaff65a3b3c
z5f475dc28158d6288b97c84ec24082a59046e4d7c0a8519293d9b4e07db622a33ab2ddbff16176
z61e1a692ee6a72b5965667597bf8d7a0556464ca6a6e3dbd71f4001c35090341e279f93e717d6f
z6150c62cb19a09a7a7900e9b79ae39dd5a8a2c3d43c807ddb53e4062baeb763f51f4992eeb960f
z2b751ee61caf22097829ba9d67e666ffadbc0e5e225c9d945f744d50b0a7a10001e2cecb7e2789
zb5795c98dca4d114567f680635271bc789b1578f757213c509a1ac4a858c8533167f3cc57c0226
zb75be1105f2ea6cc1de21ad692bd98b6cf13cd26cd037e395fc5e9be3d84df3a8c80c098112e18
z04f9edadb7a3dbceb6789541fc9de5262d52dc2459fb051cd6067b4e09a60f9544df2f7ac547bc
zc64f86d63ec4512ac72638e9bb2d76700320c8d249c1290af046c41d3c3eb399a85ca3defb812c
z6041e3cca00fa51dc593fdd9781796177769067c60e3a9f481c2a0261e02a2392fc78b0c42f3ee
zc1e0ca55b0b89004bfdd6e46d1759ec2d0c3942500c008a30a2efe550666963e60c7b0ab40776c
zaf98ba31953106c4de4a6ccc38e96f08dd93c00b3bdd173153d166d0f7562b3e428d69b3e4a37f
zfa3ce82d336ffff5db7042afebcaf158d7155f1bb52c1d2f4c5a43eb60324b083c285d356e5e9a
z14db9b00a39c83c9bff35448a1fdcceefe473a84eab2299eae0056ba074ccd6ce9c13a9c852a35
z0c8a25245b76f87451de38edb1a4cb7137781a1c8a9001cfb582b9c7956e2b4ff3adbf457940c9
z47921e925ce69fa4304cb54747b19bf98cf4a71dd36ff3e3e640563eeba302ac582c83f92c2d3e
z5de0c4dc4ca8e7ddffae0855c5f95832c42b200297a6fa8eb3bfbc800bc1e1d938dcb87103e483
za82b406cccf2e8c2c125f99cdf1dc35b3e22c97a92636e40c8d8408afc5dbd36a021b23863daac
zdf1e7088779118c5991e969a108edb3464d2dfd96e7b7bba0576b696761e3918535c3eb911ebc1
zdb00af88df53e813ff3d7721537937f344066e474e1d9c384212f4804084fd3ce93accbbe1ac27
za895d58a5662b57007194548bdfa821a3454e9115020c581c5c2a64a6064937e3a39a0a0436072
za3cc80eb53720e7b203b216e21225b64d776c8efe07e5f1447f4cb7af5b40e0d67614a2122b656
z80362d1d005d8cf059afa11d42761ad7ddc946357d0c3414fa28d03de79d188289236c95e01d26
za8668e3303725a8853dda04c8e5b49879164ce535e09c26d2f17a94862b7d5df755695fbfe021c
z52fe8bfd5ea2c7fa8cc9a401c12347335aac14161dac8fec43e66e1fc88134f4df1e2e133dec82
z35669ff4c73f40120b2660739131fbe72d8197b40bc04c38b9d14eaa1732fa26d2d4a47bf7bd32
ze5f402294cd2e017b29815ed8749938af9cb5afee952cff9026bad6d11bdcd03e790dc14716299
z45e31a41ece5d0825b4e9ae8a597d87a7d127c4d9ebee8eb08102c0012e43ea4217cb3448fb80c
z66db9413aec26c7bcdc4c83e445c2babd8f6b98f7c927a297b4ad556f183952f702e242ecdefdf
z5100c9f4340b85d7199b6b180ed3636da46bf7bd8d3f82df31a130aec447f0e2964eea2502ab38
z438c0eaea068a40016dde1bda0c62f9cd9311628f4f25e6637ee03cbf5eee8931d92942ae15a21
z262c7d38f2ba7c715ca6f72569b0cd817c1d8c3716878db2cc04515c4072ea50c4b17634892dcc
z5a22a854fbdbf794cbf21e4f35b00524759457592dda179035bbf12dc3e2fd1ae8ff43ef351281
z323cea4ff1bd1a5f9720816c0f5eb1a807d7ac12b119b9f4b70e19d8c4902f4f7447cb5e563e2d
z009bb8fc13bba3cdde2417c5952fe58ca9b9c146bbd24666312afdb7cd8961b043d60ee85ce29b
zd8096857b62243118d4a04a60e7715ef212f425357b997bbcd7eaac53c917d038fa5ecd118975f
z4e8ef29ece149b1786290c62cc185c4a7c7826b6d8f3de2d8700cb0b9b007ce692d7247b85bf0a
z52efefc0f492403281c15209874c0391b8a696dfb9c55b90ea19df2629d84a61527a4be6b68cbb
z8170cf82e24551d125f54d9ff60fe31288422fe7bbaeb8a580e5ed945d9dcb604a5a8f7f157988
z2f9e0e31d9b5cbb92e3917c07bf1dbef9b690743b43f449382a60f3891c2aff4ab7f10946f501e
z574643506dfc09d7e1e397c4fea6a60cc5ab7062f0b57edd5defbc241238ed0a604e30e432b7de
zecaa3964d9951d444ff3d01ec8002d746f85bb9edc6c078f86dcfea6a068d1b17a53a58ef7c650
z11bf70192e61b0dfa895eb9f2a1fc11056c8f89e1e00c4944f5365c3bc08dfad2004c594361f96
z3c4ffa5ea6debf264f274334ea9c9c7f1c3fbb9c221c017c64fa38279730c1af8dcded3bb5f784
z78c150fd5af982c58b2cdef14947093539d19dbe4fd4aae69b1c03c49ded3fdf9ae9342510b398
zb4127b2d7e10962fc47e7c21e021930fb12bab784f86dade81fb778fc41a324a3944a65a8d72b2
z1fedd52174087cf90d677417b66c1b4ee4239ab8e93795d04f624e4eaf6e9189a858f78555b3d6
z9eb88da95b811eac8ec98f90cd362f78ad3a3487b95d10899bd31c5e56211b365ba9d9374bc1bd
z77c1b30259e710069635f56662b4e93a9947f5f676fcfb940a6291d7ad5ef8d54c883f9fff0170
zf2f6e9940f7083145a0ad0e7b028433eeafcee79c139d6a8a84a046edf4b2d58006d15f350d081
z4fc12933e5ae7066769f95513c24f91a99b7b3cf6e35c676ed0b38f16f0fb48e8366656ef47639
z3c489e02bc8423d9d8e0eba00e35aa35491d5e2f46b1d9f478406f035b20da358d87ac814bf369
zb4fa2904e01031ddc4803a5ae765cb2b9b0b31757ed12ffef1a288e98072be51a0d8733832fdf0
zae3af0e443f3a909f4ff661a5932f93c703557c73e19d8ab6e8227e323b3a6c1b18144c4ae77f9
zd2b97ec856eb0dfbb413fcbf627d14a8c3e80b604ac3576f7fbc5203f27c89d54386657de21aa2
z361bed31c2d9b9ca05754c935d6588b59db56a8f212b14d638ee9e49b5c5bec8a86e7fdebbf42d
ze8967e3d1b74399b33ccae97846b3e4037973b9ca01182bff78bae628af57d36e9bcd8a608e2fe
z0dccc85c302365f72e9ab8af9037e9d4b5fcb4719202d523edb10ff22d96328db47ecdbe7ff027
z0e5809869befe652d44aaa58f3a1588f5586b3b4aa16c3f1e1d3fd9425f35a3e66f2057c214c00
z6b5bd0a3bdf4d31764e789945f267220a28c78cb1e8eed55a1564028a803a2ca7825f02400d38e
z4e60aa0607462a24f76f67f79527fb2c66b3582980e2a5c59966bb60c106f709172858b64e1f9d
z51128310f2a1a0240001ac93857e9d0e1df08129652fbe25766d8303fbd44ff976263bc89d120a
z6ab161433b60aca3c9e5e79bfdfc2476a38f1dd0226fd3da1635bce60bee13807dd38f451fb5c4
z088e57c1ca78a84442ae184058430d2630dea1397897410c1f31e411b63adeb4b4550634e7eff7
z37caeeb3d753dd411ff3ff3b37f2c58ffe974f172905826f1a14080083a3b00681cad2c3287835
zc9505594e2afdcde706b755eaecb55eceb779ce6ddc7831fa1fe3deb8cfc546bd5dc1982f9bf6d
zf947b08f1cd9c061b3d7df9ebcbc5818e15ca8c583203624c1998baf74bc269fd298df9ef28179
z14dc9d1105cf81036919286e92b195b796e25efd917b1ae28e63ba0877fa06c3d9918cb9a1c7d4
z3222a98584e01855fa340cb01ae4e146702e48ef2223859319c05d56debf7928cf071957f9ab6d
z49aafd80103244f1e2feb1c17621ee4dbc6f28322abc81099822bcff7bdca99e236780a19f7c69
z78176e7263fe1d37a51a28cace6bfc04458e0c359070f584c9dabb92c8fd5830ab9b5fb996f9f5
z65ebd8d08a5cca1c1f010c014406f1b5102fa1d166f71c3e796e28f36f14ddc279deab92b01528
z9e033ae1a9f40eb886ab622a161c5ce79488caf68e47b97d13cba34b583dfec86afc58c113c1a5
za57f6c09469c6c6860a1c0a748f944e6e0cba418bd6f5850f3ac5683f143461d96dacef752b1e2
z9bad76a332344f6a308f09777030f87aae60148673fc4db286f6e3febd944efc2d7fe3389f5609
z290dce47a9695df7309c7de4e8a4bef3514642878dd1ebdf8c460537c1bb6af5e5c6fd6a154390
zdb01f477aac3cc185a9d2cd2f148ac8b66a0c96d3109a91ab55d34895ba691b901a05667b8a107
z1b402a0777e9edcdcaa9fd9f67f32efe5916e820d7369475d027cd631b7811ad79b557e7dbb498
z94a4daa1c06c267f865c23d7796632f83148d39be6c1526ad6973ebe711b4f736e5a0f8a485841
z8cc2b9a19ae0a91361bd496a8aba4e069dbfee15798f189a5c333aaf230e0cf2bbd2d177bef92b
z5eda67cfcc2f77d9813586131bbfab1b0ca4b61ca91a927f076bcb3b39f6ab0ba56e28aaee4f4d
zd9205d91e155c6603c66267afab00343fbdf3d09841678c4f2f0a8c4a8eb9d6b674e31528c6b23
z1433ec6c214fb977238f58aa9362174646021f65532e4a3955ccbca9011c95b02ad525dad65dca
zdc23edbbad4eedde43c2485b3d41cd98d1cb67bc702327ee4c0f63a3b497802bb7964eb98527b1
z9f41c905c3f92d61ff0e58bb02f607a9851338658a11139c38e8b9978bc6735953566ca6b1713a
z4347fffba22b6cb86d0bd5cf76f231195532919a5550714483d58688de91162ebc07b8a716c3ff
z5c5ddc76840c68a34d4b06cf0c4c7dcc15937b769efb3dae7e73efc740d4e79bb3abd7fde37814
z683eaccc331e226c092374f5944cb704e8b47a5f2d163872ce0caf883b06b997fda639782b2729
z4bf53a2ff3a1a12303a3612cefaa981bc1f7e119a37f1eb77a00f9a43aaed54b0dbc7e5f559267
z72cb71086634aa592b76e0d342646ee73080aeeb5e1d7a7f143aa20e961575537456b929291c71
z20286a998c1573832408c8d20abc16c7c4d7c26daa3bcecf0b0f7a59dcbc273fb8dc9678b86853
za9d1b09db5208c8282c1edcc8afdcc46df0a4873dd86b0f57fa51bd5bab60a2e5ab1052e2732e3
zbce30fdef6f2794b46839921821cbec38a874c75ed06bd0cf18a718dad17eaa1a3d6ab5de7e2c7
zbd5e46b975a056a52e9d835094a964f0b2cfb2666378049470f3d039f9a34832e5041d5c641f63
zafb418ea27f0f06278b87b9a32dd8bad5e01474789c1e76a81f254aca253ed269e683cc00d6581
z4463e92c47976d0528c2b493d4a2c3376c281cf1b4af3c9d790f489f7cf416dd1955bda156ddd7
zee31a9beeb63929906dd7027db6bf6af3c676778e5009dad65f26099f62bf75e81655e8db93f92
zbb4a9b8f673f9d0ccfa068923d830b9381db124e1b5af9139886ad9f10f0650ecd36846133757b
zd2a00241c16ca10e1b1866f5c456f8fe6301020954ec11703f7b53b37ea12c13264c644bb7baad
z31bc2b7eed3cb6e68ea7c02de700e41bdd5b4d22c86637f9748d22ac2c4ba78351cff2e514593a
z5b7fb1d4a36053bb380df398ba8471c488326b53875adbf88a3cf8120775fc73d949d09a7931fb
z946f2090809e151206004a83f7763f9cdf30628e463a769906c81c2767b916437e9e500fa3e9e2
zb07ceb0c9c704822d50bd61b87e818e63e43f438fca4753a3b3c0fb2c8fdb76c6e5cc96dc35071
z99a79804089ec38d21f6a9301e3211fbdc240cb8e52b7b4b9521d8f29de1bbf18e1097963a19f0
zcaf22b5cbe5db350b813f65bde78efbb760a8c2ffa03cd4135780e4fbdb643ff1d622bbffca3c1
z8737ad1659c8d393a58b651fb8cdd58cfcaa6678ce330367d8af934618380865edd4691cdd77b6
zd02d257f6d356e9310e0a09ba483bf21c062fc5f771a646c955a0fdbd1bf3f21fe4dbcdc55d5f3
ze642b488da88fb93f1a1695f057cb31e1074aff4298661d60a57810020d88ddcea664ae611dd8c
z7836fee3e9db80a028f36c24a60adc9c0aacc2de4afac94c4f2708bbf318d799d76eb99fd445e1
zd5114ccaebe799909a10cf032ab05057c51a2d597cb59637964ebcf8b17970157d9d70cb601eff
zb72929bcf8bd373106c2bb23c973d4c892c8e5aa6bbe08333a722c139fbcd32eee538050f2a9f8
z624d8123e844cab4560f2f79ea5031c6a4e5b4af6d203cf8e8eb2fdba08de0cbe7f720175b9a2a
z7cd5e08e7d02c1016adf84f54ea1350cbf2d66e3bf8e35c8f48754fca4c92735f489beff184061
z32b3b0e15d9dfe54bb23e7a102393f98c45d313d808374213fa95a280361d0895968e2c86dba8f
zf000c1173a76097b96d8ae053239de75446745cacd9086a1ccd16a391985fe1f99fd10de36dc92
za1ff827f859ff65469d2e43752a3b8459417c0d49296b3db8897efac9ff65a38e46f4945adc3bc
zba61f8742dd256971f4e5582e5e3e9b787e14beacd38709ee02e7d5f9370b73dc0c714f51266c8
z7e17fdcf575c7041c123daa63459e06c909127d38b6d5e71176c10b7cac865a1aed6b52f481455
z93573c56a5acdff7142bd29a8577736c0da0161bae08bc195ccf3401465e10cfa9accacee4a390
zce9b87bddbc5fc02b3192ddf4426bae25332203117629d47c57daee4ea4f85df6835765c9b46fd
ze680cfe9568cb7eee938e15d6eeac244918fbb8c2e3e227b9761762c691319041264c5efb522df
zb9aaadd609e4f24b8af63fc2fbcd59248f1857fd788c087e653d527c16bb7340c320ecbb5bbbd8
z071c81d2c0e09eec7bb22282513d38bddc6dfa17e4c081a57763394b41bce8480c330fd497e722
z4b9d8c0ffdfd43d6f613a1a612fb94d19fd956d8189fec8af4a5e429ecdb38f17a8bb7b546cbea
z014d7e6bf5424f6dfb672ddf865cbe793d00ce34763abe95b4c0f6dc852325fd4c4d6a899a1a5e
z6a15c89b9a6778ee2804cb262c1ebe1efab3ce368cee2846f25b31c44ea05d754895e8f4f4c7ee
z8eb2bd09e521b9b2c8e92250c469e2a9f1e210be141b34637603f18c951e7f793268dc20e467ab
zde063dbaf2a5dee87066b41067990c873409b23a6436199b637517c61efbf464bc3dab0bcbc9fc
z47321df27f7b99feb3b68153435bf9b5d8ea871553c327531127c4be4b6a92a7d95dea9b7523a5
zf0df7702172cb8e8709c4988bb472a641407aaee79343e40183c2b589a806dafe9bb17c95025d4
z90a3c801d7dce5c83ef0e12d07b6c561d7c927ea832d9acc0f114c9f07376244a553f37fe34925
z1daa36201cc32071f0caffe7f240fa019e58d5c3d9f9d35c39be2e5cd8788fb161c152882ba86a
z5765cefadcb33795bc752374645afcc6248f6de195fd0124275301dc3dc14060b61bc1fd697871
z4c58d8e3a34b9e12db4f68fc994daf34187ecec0fdcf5517e681f13d626ea90f603d9b90eb28bf
z7f5ee60e7ee56980960a666ae393ec798a26112ae7ae35954e33b49f1680a6c720eaf65fbbadb5
zfcec038b7e4b8b2eeb1f4e8b9f1def03e92df158b8014d8bdf58dfc87762fb49b649509c88586a
z5e0d7ef89df29937eef695624f5ad9db03fbb629283a7807e09a19b26397e39f8745444bd67b78
z6e2eea2fee630efd58786e1fb35cf6f8c68f3d42191444bee763a9e4ac3856ec591dfc7b408687
z4f4d03140bc06b9d6258b8419bef142b75d45634bc8cf1214913304241242a2d7787f191338936
z9d4d25331ab119e400b8c52288d64595b8a9e9dda0b3453beba1f46db6aed0ce33b7df891a4f8e
z61ddc8d7bd691d21820bfa1fd2c8bf088e07a7e631dcb176c0b3b4868da486914c70a42409d311
z81b61d4be9aea81d2789219d5eb7f0f1c34f8115c5a8bbea436f0c3c1a3030088af7b9c20d76ab
ze09288084c5d6c019beb6492401d1fbbf5f9b08bcb63cff85396464b36e612c1dbf6bb5d86c82a
z046d332d4ceb2c8d871696e2f1aa321a626df0fc58fdabab02731f3a88f11c07877991816275fa
z6e3def3c9fb09608f3dcf024d94f75b1f172a04274669c540f134a5acd95af740b2b3ae583a650
z939e37e82539630b821d88cd44c4e5ce3e4a0b019d75046e3dcc060500b88d82d28ca25105bcd2
z777565787372ee83e18d931f7591f9e8cfb6e235c41f5d79fe1a9993ad585d179262eda0e45c3f
z0dc5d6fb14ae9eaf5cfd5dfbf49475e4910aa36bbfa1b161e48b79da80853592c773f898775f87
z79dab2ab1e988407c8a4ba8766daa4725a7d9ca5a1421332b9fab9076f792b126c4c35c26d4dae
zacef3455314ec55117b7d9dbffe5a921def02abf82c9427d9d7056f80dad4208bc4b938abe3013
z41955d5e734c18c4cb1742dc17ad5da5ea04d6030a02a372e89192db90f71fee7ebe4979851b68
z99eb37042a7d883877a67de39abe09d2b39e76709d0129d979a03054f317a42d763104795628a2
z843c78bb9050d2397bd3a3f488be0c0e661b1a604fe4bc6b83b7dd3ee176cfca68f547e333859e
zc708bbf358873be3a59e0a3b5926b3df4dc1231e83db41fba13b01d207d5e9815ecd53b5b4743b
z04feee9568fa202e09761b759098de47f58ded27b03c30c8b157445d1f2ed569706c6e9023ed87
z160720332fc6895dde77efc96fb505d26c7eaf7c0fd132b1897e4aaf583fc5f2d0234d27d61adb
zaf529b230d56650f197d2c1214e10cf4f670a780c1fd8f998cefc78b5cb10df8edafc339d4f17d
zae37d3609bf3599c5540553479333e4d5c1b4a5a97c028f1c0e96d9f456b564c84f1ea9505fc2d
zacafe9fec53ba83a8196f85746952e21fa15cfd341f59f74147b908a89f7ee32c5f45938c3e449
ze7fcbac68db6e1f31811e82f527b58fea08523f9b8f132d3a908ce06dbe2c0edaab88b48c9217f
zd966372b9c1365787b41753f3ef3033be27c036592e501309b6baf5d87f492d8fba4372a1e67df
z4a90d3d1af31dec6c3d425add85f57c5f811e3d539776a24812427a6ce981334b42f0a93f2e0ff
z50fd5d898d254fa2a9079678f545a249ee37ec80ec9f21103affbc881f0af8fc1bc3d9337f5c61
z6c7e96d844e8d1f9562f094f81000721b88dc9a740c5fc8936f956b713d513cc44a9e0a14f304a
z5ec9783f5a0ddd0d83b19a5c34dbfa08970a354c7118a19da278c122e270e763e4b247d5d572c4
z80869f8d5ed59e7b829db7718a72f21d6da96dab05e41c4764769584605352b2fec9b385f7cca5
za0241a866763fb38d0099603ddbf436a199f38151fc92c594f3896f823e5252a579c9ba4d3bb04
z02a15bf835e6fd971e6cf33fa4f210c4712496ed1294b53bfd64ec298bb2d985812749bb9a47cd
zced3f02cf3efb6bdf36cc06b436b5fb6a727258ec48f37392a50eb9dd3e67c691661b16549a0ec
z0e6531ca9c301a1dafbfb3d8ae1c3f3a9bbc47fbf27ddaabc36756a1b96738c6e6b17e97063ac9
zb58621b1230fe0e8b9fdf23982485647db07d63672a3beecd8cb6502c052646fcaf77250f56112
z59c46c36d58f8ae1192f233e0d4eea6a08cd4f1bd0076ab5d351600be150d567d481cc102b0c2d
z95d28a5a610e5fe14f40fb7393d86cd1c4ce2486d1d479e1640006a83ea9ecca94e3617461e3f5
z1dc3d79f1ff56125e75169f8166d784b7e2ace475d595f194fd06dd2b5c4c82fd5a943e74d8e47
zdc877bb883a0d656b53d405e9d9e5a02e653273984d3321b1dc0bbb9c9972cf03147ad215bc069
z0d52005529f4149bb3aec1756acb947e2fca2138f0c866791a03a4ba77017f270ee0e8f35db289
za41b5a2793d2298f16dd6f72d5b768fddc2081f1967a6a3c00a3b2bb334eef6302fe16cd5af8d8
zff846d9b4be032bffc5f8440330196b773bdff627ab52772965d66e827295fcbe7306859da8f32
z90ad1215ba80e7a5272864edf3010ad5960d55be285e721a6c5564773dedbee47185867177c944
z8802e71c5a61364294c4a702c639578b0e343eee1ef218a568d01cca90b7b23681a4eb4ac40d4a
z44d9b3875ed3aabc44ff22ae9689a00fec24bc89a78a31c1d628b761ba84a539863e8c14b2928d
z3c5750e4435f503046ec4db5993dbc73228a6b36916c19b6ccf82304ecc5cb93c1f8f77393ab0f
z83a423fee2e035308ac928ac5db402d65b3a418054bca7ca2d8c8c460bca3a7def6e316de6c142
z05afe2a3507852a4c2aeecf7a4b5110398b21687355822427d360bd47c7337e52505dcfea527c6
z3b741a8a7851b7f7bdd352200ca9629e6926048859d535534268df8af619d2c02854d19a5d496e
z5d8a304358aa4c3b86c1c1d54939be7890c5fa48364e0d107ac816470883b65a373c356c4b9750
z233a4db0c2c0050afe514599ef1ec15b0dc47573c6ee069dd27724f780112484d5fd24af3eb46d
zaaa409f592b9910aa559b5c0198e932a195f9faf530544c1cb9fda46340f7132c563f464d8a236
z4fb503a69f9d5f7afbdf61a8c8589fcc16b597deb7c81918c261e54950cbcafaa39bd8780343a3
zcc4de5246570022efb6cd4b68dd4298790de8f2380f70844f7012b1c70185babe009828147d752
z0757f0fb9bc1bb9a9f6d18b4b982c946548143641ee8e86e2d5db1d3b1d0724f97faba8111be07
z7326e8b6ccbf0df93c75353ca29b830c1177cf4da2ee75c19272bf2829410cc76d1d79d5e2e5db
z71a2b941c1003ede8391669748d3b0c4e48e169e64b927630d468802ab0605963c45cbd74df8c7
zb9591ddd95b8fb9775ea7e964e6b006001f251aa4cc8408f27846008c6fcdbbdd1b7f686e4d224
z2f162ff615637d67e84ea2e22f6f0cbb316fdeab0d06a004d3eb0aa2bba3d3861baaf92bf5ef78
z6f9c1988007e3a169e7ea9ff78266dda6a99369c5cfde8f890c4289e8e9d22c104649d2423cae7
z92aa4b641fd775b87fb784e56a36dfaaa5b13bf92e866f21bc5b65be3bd975b13d3f4f57d8d624
z5bfc30897903c0cf2eccb1191a38e337603f376d56ef066915c061c0347d5e42e8d514863642c2
z1d386d6adc471a52b0afeb7bad375571dbbfacf8c959121623c866a79d4562ccabf223d9f892d5
zdf223373e36d8fb09514cf499b327cabcd6970eb962ffc02b71f955a1d1648b130882791dff4a6
za18ca1d425cf87472c25a078695df0a8382d97f6f15397aa3f3047656f784febbe47ba3d353d71
zafde8d767b48605fd1a0ba28ec371c75668a49328b816c0aaa22630a5243f742d1ef1b1f538a58
zbb9abc3b92341fd56bd0eda793aa62f575796476f879081e3f7ecffa7748fcc5534438bb033985
za3e4d4f3c13d76ac5eeb69b1abac14a6a6d4a021f4dd0d8b5c247f3000c09f01a928f5e285863b
za71e662f529139d76a9c5dbe31d31d37acc6942e1bd4a2e25b8625f55bf6ef919ab054ec2a4e49
z55d3329f512c96035a36fe278508d874b4fb06f51b02c548a389b81cf252254f0a72f0d5b47827
z23d082200ddd2af0f24caedbdf6163c78bb87720fa4dc58734dfbc9d8b97e1c98bf090606d4e02
za6d734940a292a51e349ce7998da501f9c991df66aad559b9df48a345772360834493253b2f689
ze678c2ed66b206e2439656a510b980d632f677c9b5866f9f1ec98c56139773f610e684845ff0e2
zd3c1e68327f84035cd21e86bc32807e38a8def90f7dd8f1bd0c774fe0b46d5b9e238bb56db3c53
za3caf3267b2a53629e7799431a2baf791489cf59f8ed93391de7c2bdbc53f757878bccd4f01066
zd9e28c26d3ee34e41150f40364bbca9b98fd5229c748f3e8de6d70c3cefebb3ce2183963295716
z9114363beeeac94b74a75b88a53197fdac542c194fc457f4b1506db24aa91325f4b4886b8a6e54
z583c67fd1a1edbf40feda11216710f9250608d0deff2612c1a05c31c205d25ab372e3dab7f827b
zd204cc2942e03ea935d5eeb5cf1f7a9c48c48f53ff3f66839a1399249c56ba6176ce048221126f
zc0631678778821cf1b9507d65272599ee1fa3e57b940d77f43e84d059190c3f6cca63397f74085
z3073bff49ebb45bdeb3dcf356492200b020395af42f0d4e71a259798bd33e8246c3985259ee055
z6708f308ca11cd4d976e138e631b52cb9b0678bd084397d75a94564ee2101d98794972c84cb4b1
za4a9242865565b0ff39db1a8ed78fc6df76c0fcca15dd2b9f8de6386f6b787f52bef90c95ddf52
za43b06d5a0a4a214711ad7e7c8a6bbb1eb0ce951895b3dec646278e374833aaac191230569edd7
z1584d10d6084eff1c7c2629ecd39d8bb3eacc029f3365e750acf1c9ad499c31b0ce8fed894ac72
z4ccb062501ee53bfe6ebf37a4b3822d8b67a847d796b764569f2e9d2d182564519ce67f0b231af
z75699cc2bdd5f8b05ed698dbccc34703a00ab1c519a4c28dd304fae44708ddc2c9a8eb7b5ba8fe
za0eedb7c814d9996b4d40131c6bff1be73354ea7d8bfd6331933ac3a33b709555b4ee6d51b334d
zf85a34a984994ef8df26e25f3df7fcf0d06ad41b3884f84ba2302d39e061267287a0695087503a
z11bc8f5333089edb698356c8c189af9fd6bccdd7007d465f46bc597aadd071b0728e490e667603
zfdddf78a5c56c05760800c7c8e07af5ce95e10bafa8d864c4cca3a8681271a47b5cf251afa7b61
ze7b15f9d51bdc6a918a4a6c23cda1ef631cb11280f62f8efd9be77b401a44aff44b429accd95dc
z1d20f003bad22e78549a31ceb08b4e8e2e7bb6275ec033b44b2c3031bfb0eea1c4f6078babd5bd
z28d09e8d68ab3710337f1b4917e9aa01635a63245dc0ecf2d4e0c6cca26b853fd3f0e70d07c254
z26a1de7b37f98e9986e72999c799ee46a7f3a6212ba320ffa20b7bc6a0007bdc2ec7ebe65ee14f
zcbee030d5d005bfc1a7bbd3d057cde445054575003786435cd04660ba3d5e69491f5befff3c3d3
z584ad6745f78a2412f486f0e5a437e88d2ee674dba112d16a116e4fcf84ee73f29d169c4bacb19
z56ab6e044955a3586267e1d6011e9fcdddc9b5541ecf292415348fa988fe394f7d51bb6b488d27
z6ae2811608b44a30f657320674975d44a344ca1afefd569307c0648e6d3644585f05571763a11f
z2ec68379401f7cee61e8eeac20c193e798eaa2943dc18002fcc11f7cfef3daf06ca005c2627542
z773bf4766dfe395c9815639308713395a4cb6d9517c7d24c9d722048a0bc0f4923778024cbde6d
z59c2f4be8e89d8503661c95de82823e8a7c7e36e883828527626d429ff2e3f1cd61ce7b0fb81aa
zcd934de68f0efb70371eeb7534fed9a830fe3bc5fc666f9a24badfdaf3c5ca5d1120d02c97fe04
z630214f410b49cb17b235c28f1c015dbfe5873055143fd6a3378367eebe6f84ca2ca6d03d62904
z23eecec3b7dbcb392376163de74814c0c2b57390c455fe61fc3789354b1ec2f749d785c7341948
z87b420b0c41e374810136e7cd642c09f61d9208b8b2057a6885b51b49e998a88a9ebbe81a9f2a0
z4db55bcc3d46858435ea850f84904cc1332c07779f9aac99420d82d8c7b2e8bb5e2dd3c89993b4
z18b3478f44043d7946c06853bbcc2d84159c9c825e280a8c1f689e76f42be5bea225339ab5271a
z7a693660ebf3dbe2cfc240b6773bfe229c9381e4c32131b9c237f2efeff46a4520732ffb85d9c1
z5d7736baa563a5fa2c220823a89256e3234131ce8274668d884d52759bb578d052e0cf949b20a7
z775d4e6b489c3d698f4082606289da89621386033ab6911b6a18626d45d4d3d6a6ff8b025d9d63
z5c163904a84571329c1704a724f7fce8141f174abc8aea647621e3ca1a6afb72f40c14c159025c
z734532988ea0d58c5392920b3775bb9cf9f7cd87287106b8b33bd6193164540f3ee10565063512
z16112c86c8f647744cdb81c88833e16bd37f21f53793a7548bdd3d1b396e4f1130622db1b64ded
z71d6a63b84989ed4fa43648c05cfe5c6471bbfdd8478cd3f79e6141fb9358da856239b3eb1521c
z39073260253e3a3326ee96d00ddfb019cb0c2735e3f905cdf6ada8ad444f48865a1d5a0413ad31
zca6be3004773f5f11b1b3c3c11c8afc2cfb96457db8ecbeab270b05bdabe2e7ac0b4335ea9686f
z7fe64e63a795788277f8c710d77ad6461ba063c05798219186e5c8791a708b4e991be00741739c
z710b97f7aa69ced2a16fb0c934e3d8c54ef4687a727ae975912c3f28e9aba7ddadba0b52b6b3de
zfe7d66bb5e30e419ccdac5b8bde9d6d4bd5775a27d5654c4af8dade5f7459da188e2e8993bd7d0
z0ca5196fb04726b92adf06516a25da3c796eb22b2cde30df06ebbb147b87c3eb39eb84f63efa1e
zb098763dba05e114bb3f50e3565e2c12f539a16e84df0dcb5f20f14b6c396db948f259c9fef1d9
z63ffb378a6cca7410af248016a7ae8905aa78b5f247967df5d2d63239fb961bad062e003c2d2d8
z5cd3c453e455e83c7293276738b42d26ef3e14963de316f79ef81b0dbd9b215ebf5555b582c4f0
z460ce4ce3ee3a916c6d4c770e846b3526657007a534950782cf00abb3de42056cd6805f0a1c529
za3f329fef24f0f2321a63b7a2cce13462ec7f5ca52226f2036cac677fa2f3d90dd7f8925a7a330
ze02572bdeeecb8fdefcc7299d23b508474e2898df3cd29faec23942e6896c75f8cee06f909a686
zdabe093ce1c8c62430bb3c06c56f115667f6bf57ce14e01cdf66d1f1c3e5b81408db62889379ad
z0f5a752663c4ac192a6df419cad2039817a68cd91cc30d4cb2ec422687157e69a87fc8dd2df2e1
zbdaa022a8ef66384570a3a736f36da9c484bd32dfd5d2cac69294e50b8ecd9d73ffcf73cbad573
zfe92070fb6bff48005ec11d59ffdf2be27918cad90ceb4fa5633693fc7c50032456f909b17d1ce
z76f55b987752dcd4b671737cebb2cd5553e65c471f96b3f37811d2c0949317edfe2ee1a9f5a623
zb60e4d47bbb12caa1ce31993bc6105ee7872876816e4f355b2066c08541f57915bf33f90c86da1
z99bc71cf2d0d862b2efcc0dcc48688a8ddb7c3aed197f2b73fc542aee75113961fbe575152ba19
z42148c265045ecde7778bee506c0df525e318b9bf60025ad8be33ea7b4c6af67a4d1927132f88c
zd3c585bc67c10a3f7b827d9abaac8af1ba2b9ce18fe2466db742da14eb019e1dccb26576a145ed
z82d1fefc3ba3c34db3509feab7103cf0ffcb3d053fc2ee8275c7a246237e89d7540f717048107c
zf0db6d4af6f8e7924322ae945a97e0c5cba2d37cb4242c6c001999d5678bacbf73c4f53b722242
z87e905b573f531ebe2813d65d77eb1d347719836cc3d5aa9b25c3328c5cbd0455dc834d1650d89
z27aff7b5c8fdfc2c20a01bc40a8783e4ebe6586ade7f3a736b7536a043416dd5d22e95f91608ea
z3862a8969a4fdd20f42a25ea3472e59009b5b47cdedc1bd998aa708831c7a36c8eb45ca41ed6b8
z5b73c3091447fce694942b61fea4a179698b6be0c403483dacdc1429f7cec73b6f2c6d91f7773f
z1f99d8f5befdf2818a0e7459210c35a0bed19b6eceeb5ed31b69cbde8a80de5fb17a98df6c98f9
zfa0a6cdf148b36793c1e48431347812dea0b7b9d499a7db135be239e2e2f4cc6746f2e6aa8b23d
zb025adc0bfa00b32d4
`end_protected_0in
`else
`ifdef MODEL_TECH
`include "qvl_gigabit_ethernet_xgmii_link_monitor.mti.svp"
`endif // MODEL_TECH
`endif // encrypted_0in
