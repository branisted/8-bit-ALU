`ifdef encrypted_0in
`protected_0in
ze74c34e226135848fe16db9ffd31815111b6d7fb642c521a3f628cf6da949865580b22efd062a7
ze90adae0e65e66a2c36a587d0a790699161455169ed55a01f2084f11770a774ec4c588039b380f
z6de9c5084882a40b79a175f5c2114b2b6d78b070cb806e1c0aa9258297f4687ab308bc470f0040
zb0b1de382961eeeaf2e279e1462520fc31c119af8f2b214846f56c2b3cd2eadbe4099496abff18
z15cec83ec4a77b868344aa20ba7360908f5c0de2a79abf8b3534b883bb12180f68b5d4beb444cf
z3fba8f13afb0abfe8fcc4294810f75afe452434d2d0f1166236c82f76edf1e12979f04bc35693e
z32ae028996dd85737a8f5adc1ebb94f39c940246e887647b64782cd7ab429b0544c173176cede7
z01dfb26b1f73408344a52b7e1f117f12bb9c8077b34876c2e6fdc085981637012dc9754765e1a9
zc512ce062e0b8fb16a214591f5c81e1353b900a611fe1f4886b57940b41b7f2ce99a7b84b04b90
z916f717e73bd10589c81e207ed77ec660a8cbed5b487fa50acde1b055c8870bd8676023f21ddcf
z9c98cc47cfa2d654ff1365d1f45035a045a66c5dfa8279050262529d2cac9e64fd27d9c7de62a7
z731bc808811ded9016570962244887f98fe5440167bd0088f2f049df882af501358497c3b28776
zcdc5426c7f52a851c35106bb93e16fff98478405cb2c034d92a13b05dd6952355a8276837fe1ec
z31ed579935d1f03c8aed1f61cb6f74edabb0b099810d7bc07560d8599c70e6a86f124d46b24212
z6f7436923665fa4f4b9ca34814cd5e1dc0f216c9ecdd9bc4397e1ecbbac46671de6cba2b5302fd
z326344ef99372f0e53218d316ec3113070a886a09f7f3c491b2b14edf5c8ba6b3a4c7e157d1004
zf3558815e86434400eff349c425b15a130edcec15473a1e768cf805ab7876247c705be3327b3bc
z41d0e46f17b4e13cd0deb56f49b952dd6571cff90db4cf4245e0577e143e68084a3bdfdff7c121
z856571f8db959e9260d96cf692f0dffa9ab13ddf85f73dd9184e4df101facd5afff35758df10f2
z6cd940c781b541691bd94021a6df1475daf2c01ec564b6823564ddbbd4b45e6d9cee364831185a
za38abc72e73c45a6cf2a71b9eaf8caf5833e6797356fde956eee87b3b800c75f3bf059878c8b54
z777d807afc0fd7d069a1413d4079d66e51b8b554a8615576b5e4794a9ec84e906bca5a7abb65c0
z6bdc0a5eba61031a4b05bcb919f4f98619069d02433b748ec3c9c8195fa2a6c8b0aba45360af99
z6ae0d51c87961a8037b76c314a7e096f93cc86fbb9f22a9fc8b408934d1cb07b4e32b7e01d4d59
z0bd673c87fc2a78c645b2a08ace743521f50a6929c3828a438c8ee6826768da6cab55525a3c900
z4377e70207394fe01905fb4b56138174105f3b2081f58e3b7f9ccdc8ba8e92f0a04e9916f15bd3
zfbff59c1f551a009e56b8e651f1cc8c27491460a7b3cebb84dd82dbcae3e48efa71d1f6aabaf82
zd6d0c9689df53840e2e25a9d72f12d820e9ce940edecfd6287942fa0d78dc832c554165536d647
z38a1308541a02db19b6a431311b26264edf0e2b79823fa85ebd25aec2358ec664b92931fc2b21d
z9b706a1d586d5e68823cda348278d42c3678c8ef5dd375be89e6516530619287c62958503168c9
z362d62e33932908dacea5a3d682f9f5c70f1eb140f673eab012f103515f3a229e38f658885b8e8
z5886902e40fd1cc52edd45d0143b6848b5dc16ed45b4f72a52f564608f04e4781322eb523c0d71
z0f93174f0536e302cf2ea9739afabcdfe78d9306af2a187465555ab6caae9c51b69143545b1caf
z243968bc49ebca70d23b75bb9ba46f17f368805f297663652b86f8fa5b65a3c16115a4e061afac
z157b65cdc5583b20f628c4a15ec8c53e6b994d29e38b61d9f939815db341084cf778652fd61933
z1dff8b40f77ceda6d564cd6bc41407d2ce175f040f55960c93d1f9cc1e44d1752550381f85e409
z1e2b19599608652ae0e6272a9955765ec25273411499dd35e39a5e519eb8705e805999d5cb1b44
zae07ef5643db84201a2b8585e0d978e580ede8ae36d29b1384d66a56584428484bf715f0667aa4
ze7b47e65e8528b88397ca79a68ec49a6380de592a1dcc2b02253f39a1dc116e743cb1f832a0b2c
zfaa2666c240bb54f49ca6e63da91b4faf991de473fc020371b9a6ad9f33ac0bbc2e86b76d5b73a
zf088ebcf113cdd96bdc94755602364ff5e4a7f168f8e43e0cfe2bac0dfe28c68823b5781d844bc
z8169a0d787500e63183281ec8b507f8c4fd8bb5f03b5d6651c511f3c538d7340ba302e69810bca
z1ed253d8c3664ef502f62c0c5dbd1dea1fbc87b3aab741cc421758bdd189174cdd511c9fda0f72
z4fbbb0269ba25ef09e7dc143513d8a0594a11a499d1f6d9409da913f5fbc025355b0acd80347e8
z06a8500d851e9afd0a2ff2c21f64ec179e6b3971c489bb8c49e1ea8f9679050fae37db65ed260b
z92e9615a6da708a0ef9ad286e9f73258b8071158435d9fc9d0a4fe2a5b0784cb5c27fe1af3c861
zcea7e62c37642b9012e412aa43b96f22f0f3b3de2cf62197f51b668128daf9d99728d4af152594
z84b5d6bf015541565cf148fe3a13b124a7a9e9f5d81f2de5adb3ecb5f869e23d9d37d5a6c2432d
z573c2ab565ce7481cf1da25e0f139fe58c7f0f963cf197d7826c4fd7c07dc32fedbab510dc4071
z5fdc1995bbbc429478a159884285449d74ea2ea4c85d17cc43af4576ddda2c40d1c64de4ed65b5
z4ce75c781dfc25c5336f489eed5ff65d89397520c05ae10aedf19319009d1b1c20eb327b84d017
z41602acb6c6d3ad1a762b3aee0cdd9762543a7247402dbffe8af26b2fe3d44cbd6d15d4ca6ac9d
z6b6840b70df7f3556ec689ed47783343148b3a4e8dbc4b6fab2bf57f87faf5427321eab2803591
z1f5ec83c51c3829e03e93a3c04fa23e88dfda125897d708dd9a13c8a92f2790e629775691f4a62
z7f310ddd384f621de33d5420cf31a0e96b45318e0f92aded175a4c7d7321f230ee1d7ad99d6da3
za39ed3de9363f64b2107bba291f92d8a21a1123ce0db76181b1d1ed241113853e729ce3cfa0195
zb9841dd1c4a791beba94daaeb604ee820d7b3f8a1aa0dfadc75498f1696a4bd43ab3252912f146
zd879ab00b154de27dac481fef01a9b58fd9276460653fee76c51a70007ab9880da27c92b57d408
zc9a57729d215aaa488d13d6263b668216b534c24b456dfe937322f44ac9a625fbc97a25c355bd8
zd82edae12223be25ae363da9e3b5e880c8c52db694c3e45b8a1132aa0e3492825616fce461e797
zc13a37e98409737d511f7c84ce7db9d9411afccf348d11dad27da5ee2bdfa0e93fee9f4a34205d
zf66442bb454295b0b9a9fb17b6fac21d6f6b024b34bf26676b74f65e42cbc206220c536d31f869
z5f430d6d6d7395e3dbd5945a0bf05944fc5fcc2cff448cc291cb441b3215efbd3114a452e112bf
z97b9dd91bbba326a1a60afd811362351ebc99c0fc70ebbc7eb89a31e46d1c1da9ece86896c6ccd
z033b7c65769eb4b9a966dda26a715a476aa235c47c0f33de279ba171a3fd959847f33c1d680c41
ze054f8dcd6228e298d539e682c53c0c435a3dcb4ab39d2d69a303dc039816db5391c9b41dc491f
z489e2d31c35408729ba44669d7d3bf2331a7efbb8609186a9c3ac15c2313bc27556ab098283cf4
z4610d2d67b12d97c848c760f9c0e4ced1da592045e04e6ed12d4cda9653baf73aa41a0b1fd2fb5
ze3624573ec8471ac34dd801c84bce44fd4a2e868bff3a1b446d79cc66dc48349117fce88285f4d
zb7bc4712c8e9a1e1443656b8e5d74dc9fa7ee58160aa037169f6faf21e999dce952b5d94026f57
z0ded2a0262e17dd218a8d2f0ffd96645c43de9ff0da9b4b718614844e6bd0cae623ba08737a876
zc93a815bf27ce196e414e621a86c0ee789296be950a587e2e756e2d9096d70f718c2e4760157d5
z5b2056be1d9205c753b8ca73788de7fff67c96fc3c11e496eb38ac62ba3df54c66fb9dad035325
z4b93d2034071392b503b15d7d2537ea7ed1e40785b2b8cc9460065df30bf02bf45f1ebbe878eb1
zad6de9a39d493952d1f71198f5f1b2ff908afd8caea73a6cfe51e28155b82ad9dfee21795d6619
za18f6ade59bd6f28a2eb4d071c3e361cd4a22bd1742710db664e2463e435d5cacb7a9c1eb3ee1c
z269a012ac84f393c54e7a0665bef532a143f871067c5477c2c37687333b9b77d62ef97d6126c7f
zf794f31cc5d50e6f66033c53f28a0da1f1f76feda144cbd5a75fe1c9deeb144e99f71d732e0fa8
za20df4805ee276eca6f7dcc5df8b5cdcffd4870331ece446cf1b8f76a59e66f72340f2a1b2322a
za1795d3b97bb39963e95e5cf5c6e2fdcf165ae1692524fcc2d2b2cc1d5f772bbf1b4ef84f04302
z82dbeccb5cb7a1f6096682199afbf8638cc9b849a0d526686cd98ee11eb8e98e6cd9ff45a28465
z892dd86fcf3b553f4be728f27ddeb6936ff64a72251f00d0a7fe22809ead79b9d13fa5774c5679
zce893e91308a9b2814b968e2cb81bf90e6ac40a348f7e0cbfd8d93ccc6cb2e9606c5478802f422
z9b82e61949e62b7b6edf7bdf2b7c44ba701d325af1fb0d5d3194df906c68c8df1cb9f9158a7024
za9e69c23f6390d994ae41a73afd60aefda086ab42cbd2b54f9855d420b0c3547c33a9013ab2693
z9ea31002e94083a864d1db656d56dcfedccbadf698052040f00df796b4116f8a0f7ca52e3daa33
zc36553863ba9fab5898578d991a0aaefffc157c98c0384209e9d01bb2a004ea2a58ed9fdc455c7
zd9081302823edcf39b6fca5aff60b75406e1c38cb787c68df5f208d53d812fc410653f4e11382e
z63f86ec96f2714c8dbd2ca33bf660b3f0329f1cc6571b2db2fb8abd7cb84e5a7a163b637895655
z00dd0517f246b1c719afa5965a670cdf0469e073813bdecf26831e0079520f777c0b7440007e17
z0947ee5399cef637e3dc9958d63d8b51739c913a6787e6730884ea78791f90863aebc1396a2b67
z76ad7055a0325d26396399e8fe32db1eb0a0fb994059d74bedf0dbcef2dae43c6e1ba16db69ce1
z84b2a085db12e4e8f49d65c8c01cf82924fb07651bf5401b08643c479fd83e976f124a003b51b4
zd5b728269eed7632efcd8784a439ccaee4c4cd080832fdbc6a97c43e1d3307d91da10a592ceb2e
z3624535de38741779bf151cee7049d96f06bf0ac1778bda6c73642393a88cb1736bdb8f7dbd320
zf88b1f478fea3bfc86ac87c425ca368453635aab546dbbcab2aaf0f70d11899689e38a3eaf7ae5
zf5166c39c2980f5452a47ce666a962d305c5d039a2fd6ceda4ac55e44dc18a1101cdce1d558d76
z066e32980c49357992bda178b98382f01217fb033a25e64648489114c3bf98f9a74b5252fb6db7
z0f15e536045735f74e22f20d34bb61e01dcbcc1f0e5e148af9a6c6c8d911d5ef4192bb008af2b1
zf7f4c37270b200b532239c27b8e0cc3db4ae4b447f8bffa11f4070eafc54d90dd59a8fb38d219b
z6798f2ab95a6b5c843b4306b6a1396716f2b3b8f88e98bff5e475cde48ec32f75e5c5605a25e24
z6432344043ffec9a6fc3f2ab5dd99209cb215900215a453a7f651732017a80363dda11b46385b9
z95c3e75a82636e5331df9b795829ac29dd98dbd2c454a7913eeefed7d35a86f32f302c3990a150
zad3fd49c3af4250a51e5c3f6400db44924212a8b49c03620de5ea3b84c340ab5a272864542338a
zf03987b1164de8aeed70e953a279b42dfeb7dae8dc76b574a6867831ddddcbe55700616e99a10e
z5130395d3d64bfc6ca197b0442facc0f5054f809606f8bd2bea4033fa1026f110cb5c2c51712f1
zf6e4b1522c19eabba238065ca01e77842ffc2c9d07789530fe58556cc5af7af8477ada34b0bff8
z404c407983c99ddc9a27955929bc6e5bf57280ea964492c39ade9628332096de377fc5674ccf7d
z74b70ff8b6695d9e9943d69bdde560c92535a2e7bd550f4c45329e8f5d9fb70e2c8d95cef9ab90
zb46289a919410f920c6907daef7c870e571e94b1dde99ea6edf607eb7b1205c77dfb03e36e881b
z4a962699a6fb27b69f5cb67851a74d874b6ef574e754676f21a7e3b7bdd903164736dba9faf856
z770b289ff523febc437a0525199b613996bddedf3705398ed893386c82c885876ed3f6cec7eae0
zb0bbd2fef84bae1da7733ce61cdb840dbbc045227928410c16933ab510736d7828ac05428c64cb
z42151a00d6f5c79c39635826a3c0064623d2c7c9edae1043ea710fed1b43ab603c0acad4ddee7c
z375dba6dc5a03d785cfc0cbbedf6aa0049efb9e03f140a0c967843d982d242e6eac32469396854
zab2bb7b2cce51a6c5a7b0598497dd32f21e3516c2d4a5a666cd3ab1c7b917bc7498364d9bf2c73
zde68f8dbe66d5d00047351693e22b615f35cd6a467452dda361fac284f28afa53d54d9ba66aa79
za260328240058cc209c3e619bd2aa3ad5df7cc2f58a7e403ae3d9ad064d4098c1585e0453acbab
z2fbe3841e789bec626e4a8f18a389f959e53a1232bc0d3e70b40a3bf9383d96d9a9a82fddfc10e
zfddc9207143408e06dd2cadc2422eddd4a5b14e49c81ca3b6edc5beabb26506ec9a86aa523f6a7
z260ffa57820074ab9e0e06a41e772dafe757c39c6eef81789ff8489c72d3e90d7a98ea3d561a0c
ze354a370c0e84f4658c3f5c52fd0e72087419c92b317dd8ffbfbd58fc3b771b2c713bba0f5283a
z61eb1b5af3852e4cf61531b38362595439283bc5815fd95d0b20e3500e151d62ba1671dda2999e
za2c24be0d1fbbbb81a0a8706df563dd5722ccb79b47213ed8392440ba7e12254192582ea495def
z81924ff5a3a81384d256c9cb50e40497817b8b6c610a25e3fe7687261d98f45fe3d5a214b22391
z67edf479de4dc57ba7b68b238e7136922ba9cae68fb7354e94e613e7653136cb7ad9e1d6f70cf9
zbba8ff024ade5c167eb0c635f04a1554a9fdf91616e1612f9317457eeb9c60d7d10f2f6abe1ab5
z922e91a892e74ab71787732a15863b3607d0020980ea29b7d7bcbcaae721b512c959b75c28326f
z04b9d1098c24f21042338fc406d4c71fbb9437e776bcbd5676cf09f1fe75e6e11d82cf441b151f
z5f1a0bd0af4e2e277d8c681406efbd55c8094464d20853f2cefac51002834754cbe2f245cccc95
z870adb5be28e3f8306cc16a6d4abd36b2bc61c0b7bb0b7a2fa954c537829390f9eae3e751dba80
z48c6b83d31fb9328f2ae9186f7534a7c94ed006439fb711f4889ee22345ace329fcc2873d23865
zcb435f2788427bc3921584815b3195bdd26076ae2f9a062a5707d2cf1ebcef8ca86b5fec046214
zd0469cb21977888525b5f4b1509a649766601db66d1dd130ec4c155b111670d7f723fbc15799f8
z89eb94ebca8b49d0518ee32e34f2258a8ba7b5445b4b993bfba82990f787f2e4c95d72b31ca02c
z6a367e6e830ce9d71843158bc37641df04323ae6a8dfcd66547aca7fb50eca8a213d662e47477d
z8cb5be0dac78c39779075df85caf6e3266490167f4afbb54fbc301681112311d853b4062f9f938
zcc197e410460619ee642e36d0ce5f57a9824da319e7cdb00e7a9d2d8fbd1ecd6728944587f2a2f
z4b1f16a200246c8123b8d2e8c9344f4fca83712b3b2e4e3150316d774a0273a5bc4671448b8192
z5d8a7884f681e1cc758ff4995ec9f30aa412a7e15a0499e557a4c85d739810d46dd87d3eb16dbd
za8e20c4ea81ea7f1c613ec86f02dd310051181c58d4268a636ce502589519772d44362b8b2b16c
z5cbafc7f6f33d802234f8ec09d1c3d56f2a04f66a1943cb1bbd780bf6bb2fe58e123ed0535e01b
z04656672cef12751efbe64e0b74b7be0afdf92be69b5075c14deafda0da74de395ce390cd0d84c
z3ba339fd0ca3c25b7efdf452003bb00ed8ade01c715d535e6b18b21507c598084f0a295724fb91
zd481b5bfd71e59ccdf9163ffc0f88d09d6cde5d3f1763010b3a00743180f3d17dd7efd5dbde124
z8fc23ce706cee794337ca11d90b9eea2d1c8d6de7f746a7ccd841653217182d231ce4653e7553c
z47e8ffdc7b8a43bfe11e45b40e4f63787c695e3b45fc437379f6387928fe24c500ef7e9df31da3
z87a55b42365dfdb9530b751c7eda51e08013b9827d795a13682ae1264964ad6472c7f8f3783d1c
ze1c75840d61dd8ea29bb5b665778954d8841044627751cfb04101c71b45c06accaa148223f2599
z905907ff2423f2395b8154254bd873bc48aa3f2da61d7a696896ca4a2d63f0b638067b7778ec8e
zd3494713c6983b8fc065855c2cfa265bdc3bb278a54804ef08d9038ca6fb2436ae9478f2fd02c0
z1255e30c476ccab4a2d61420d2f57faf50836b36044f28de83b0388b558fc18253c9dc667391b4
z9bb81dd494a067aaa79905f37e33da772ed71563c8b839fb714fd03a3fa3a071d6265df7a6c4d8
zdf229172662975611c261a16bed9046bb8b6949bcea9680e4bed79e216d874d3deebcc3c0510b8
za72d533c80f34701fdde46f9d69bc4fe7777af76b1570f14f008a0f22e01e4335e35e0cd95d35a
zd6c27f0967e67159984d0045da23ac7b8f5d70ad6ab55d87359f3c3e4f05e3ae2f7b8f6c78b69a
zac7f465f12a1bcc09178e9ece7e83c30298bba1775649ce7d38b265a829f5990e2e2e15c942bfd
z49537846c9900eb4a6bc570fe3c95d7cff0529c8bc3d81009befd071145f875dd48af6ee168f28
zca8ea057e88bce7596b3847f1f8dcc0a60e7ffbf9da127364bca794fc8a1038b5425079fb36748
ze5e73707a199a3f40e4327e76dab62493870afaab72d76424d4bfb0aff4aac06f03a64c403b924
zf60c5ec2ab9cf13e4660fa7b27c6d94caf6254ed2b912b24c43bcac38444d93c059990ae4230db
z2c1d81463d2201319b1492914ddcdc60d9359c640f37831e2fc745a7559bc730b36378b9edcaae
z42f2fc7bdd123565b03cf099fd030f6799a78fd56913500c5bc5b96992595e16ae61c01c298890
za43f72f9c39b0769352f8be6503aefa366150599485fda4c611d01d6927008e1282a9e610808e7
z1ed68cc705c7ba0dd2a1ee06a5f54587f7841d74625810b543a827c082b2fb50abec2f776574d5
z9dd24204309e0220b92272022840cd89b3134fea065d894ed8dfc8653b3776e82305a399f2805f
z7145f414fa1eb5b0d11a7a30c9246d86d23bbcc0b3e01dd8934e8b03a859b52be2656a54a3edf5
z9c59a350c40046b6ef6054c74d31a41ebef5d763bd4f3479174a4ab5678797455909d6ac97c7d7
z77d7772d9c1ed313146ac7c0ea1a783c516e5b68b8d5b44cb68abf5824ef364647842e5750b11b
z23c01d8ab453d26e4efc15650d2d374488a1a8b76228868100b9f118804a56611bae22138dc541
zcc397aa3f31ff756f244ffe608c5aa716e48a55670805dcbd9df4a7c9faab6de2e7bf1db86a4d7
zc62b5e2dfede308c41a292f956941fede6dd402000b810cf6d519887d6dbf7f0e5ec4836b93c0c
z54befca96b94465fae75fe21fe467579209935b263cc6261f873a049269674bda878cb0cf75250
z041752c9f8e9de3aef32ae04b453ae9829e8fd28fc2c93f80d17d4769504156d47f8b474d91692
z1f216ae6910f6117250ff64124ffd60b690fd992d68ea3cb00d4572e2477ba97d5def230279c8d
zcf639e92e8a0274ecb7de88cb44bb9c0d1ca2c1cf5dbfdd380f2124e440b42c5379408c029b927
z0768fbf31e916e31a9c4806f16edba6551267bf392c92242dc951d46cbde6c93cfc83db8aeda75
z18566b80843543d81c38f5d6e45277e366f3ed482688acc2da1ea83aa8e3339f74751431c7ad6d
z0cbdc38d579e006950706738526c4e0094d568f12419c21f02b3dcb0b92795326d862c408dd818
za99d42a394c9d2e52c1116dea2370ad37c5c0073987d3dbc618576a27bf0f303b8cb93941950d1
zcce3f47f7253558597adc6b60031766935f5eb35afd1d1aa216138f05842bf89ca6c1e012eed9c
z27eb05bafe5fe980c0a5bee5bbef99b8b0b24370b761a5c35251c11ea0abc93ddf9807e6a9fc4b
zcf934e1e56830d0f58edbed4ebe4714e30d1334d3ab1ff7bdee07e9e942d6e9c6e1486fe3ec474
z0d9a9eb8926177f3fec01175534ddfa1ff3f8ba58375346f818be90e058c747d9f62fff4a0e341
z47dd1802b2ff039443038c96594e4e022a29dcc471f245be820689373b6f950bf775f668391288
zf22aa0832f8ffaa964d69263a70e36720ece18afe2f21736999907ef8f2d996fc3cbe95ccd0abe
zd4c413005652bd0bc0eed004cf014daa7fb973cf3d227df93645dbbed13a986bd289a6a4bbd1f6
zbfdced68a435dd06c68985c53fff9cd328390b8148e542bdf4bba01157bd81798a7c43cef2b4b6
z5d36be0aceb6b97220b661e2
`end_protected_0in
`else
`ifdef MODEL_TECH
`include "qvl_pci_express_sync_fifo.mti.svp"
`endif // MODEL_TECH
`endif // encrypted_0in
